* NGSPICE file created from opamp270.ext - technology: sky130A

.subckt opamp270 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 a_n7636_8799.t30 plus.t5 a_n3827_n3924.t37 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X1 CSoutput.t156 a_n7636_8799.t36 vdd.t240 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X2 a_n2140_13878.t23 a_n2318_13878.t52 vdd.t106 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 a_n2140_13878.t15 a_n2318_13878.t14 a_n2318_13878.t15 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 vdd.t239 a_n7636_8799.t37 CSoutput.t155 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X5 outputibias.t7 outputibias.t6 gnd.t170 gnd.t169 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X6 gnd.t329 gnd.t327 plus.t4 gnd.t328 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X7 a_n3827_n3924.t18 diffpairibias.t20 gnd.t154 gnd.t153 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X8 gnd.t82 commonsourceibias.t80 CSoutput.t23 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X9 gnd.t326 gnd.t324 gnd.t325 gnd.t305 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X10 CSoutput.t154 a_n7636_8799.t38 vdd.t238 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X11 commonsourceibias.t79 commonsourceibias.t78 gnd.t15 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X12 a_n3827_n3924.t38 plus.t6 a_n7636_8799.t29 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X13 commonsourceibias.t77 commonsourceibias.t76 gnd.t51 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X14 gnd.t323 gnd.t321 gnd.t322 gnd.t305 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X15 vdd.t87 vdd.t85 vdd.t86 vdd.t46 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X16 a_n3827_n3924.t13 minus.t5 a_n2318_13878.t42 gnd.t118 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X17 vdd.t10 CSoutput.t176 output.t19 gnd.t57 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X18 a_n2318_8322.t23 a_n2318_13878.t53 a_n7636_8799.t4 vdd.t103 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X19 gnd.t320 gnd.t318 gnd.t319 gnd.t237 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X20 CSoutput.t24 commonsourceibias.t81 gnd.t84 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X21 CSoutput.t153 a_n7636_8799.t39 vdd.t237 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X22 gnd.t339 commonsourceibias.t74 commonsourceibias.t75 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X23 CSoutput.t172 commonsourceibias.t82 gnd.t348 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X24 vdd.t236 a_n7636_8799.t40 CSoutput.t152 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X25 gnd.t317 gnd.t315 gnd.t316 gnd.t237 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X26 a_n2318_13878.t40 minus.t6 a_n3827_n3924.t11 gnd.t85 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X27 commonsourceibias.t73 commonsourceibias.t72 gnd.t202 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X28 vdd.t11 CSoutput.t177 output.t18 gnd.t58 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X29 a_n7636_8799.t6 a_n2318_13878.t54 a_n2318_8322.t22 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X30 CSoutput.t173 commonsourceibias.t83 gnd.t349 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X31 vdd.t235 a_n7636_8799.t41 CSoutput.t151 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X32 a_n2318_13878.t51 minus.t7 a_n3827_n3924.t26 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X33 CSoutput.t150 a_n7636_8799.t42 vdd.t234 vdd.t162 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X34 vdd.t233 a_n7636_8799.t43 CSoutput.t149 vdd.t205 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X35 a_n7636_8799.t7 a_n2318_13878.t55 a_n2318_8322.t21 vdd.t112 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X36 gnd.t314 gnd.t311 gnd.t313 gnd.t312 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X37 commonsourceibias.t71 commonsourceibias.t70 gnd.t184 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X38 a_n3827_n3924.t8 minus.t8 a_n2318_13878.t7 gnd.t29 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X39 vdd.t84 vdd.t82 vdd.t83 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X40 CSoutput.t148 a_n7636_8799.t44 vdd.t232 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X41 a_n3827_n3924.t20 diffpairibias.t21 gnd.t187 gnd.t186 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X42 CSoutput.t9 commonsourceibias.t84 gnd.t35 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 CSoutput.t147 a_n7636_8799.t45 vdd.t231 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X44 gnd.t37 commonsourceibias.t85 CSoutput.t10 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X45 gnd.t310 gnd.t308 gnd.t309 gnd.t223 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X46 gnd.t91 commonsourceibias.t68 commonsourceibias.t69 gnd.t90 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X47 CSoutput.t146 a_n7636_8799.t46 vdd.t230 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X48 commonsourceibias.t67 commonsourceibias.t66 gnd.t203 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X49 a_n3827_n3924.t36 plus.t7 a_n7636_8799.t28 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X50 gnd.t175 commonsourceibias.t86 CSoutput.t50 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X51 a_n2140_13878.t14 a_n2318_13878.t12 a_n2318_13878.t13 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X52 vdd.t81 vdd.t79 vdd.t80 vdd.t46 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X53 gnd.t176 commonsourceibias.t87 CSoutput.t51 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X54 a_n2318_13878.t27 a_n2318_13878.t26 a_n2140_13878.t13 vdd.t111 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X55 gnd.t114 commonsourceibias.t88 CSoutput.t29 gnd.t71 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X56 a_n7636_8799.t27 plus.t8 a_n3827_n3924.t35 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X57 CSoutput.t145 a_n7636_8799.t47 vdd.t224 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X58 output.t17 CSoutput.t178 vdd.t0 gnd.t16 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X59 vdd.t78 vdd.t76 vdd.t77 vdd.t59 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X60 vdd.t229 a_n7636_8799.t48 CSoutput.t144 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X61 gnd.t185 commonsourceibias.t64 commonsourceibias.t65 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X62 diffpairibias.t19 diffpairibias.t18 gnd.t123 gnd.t122 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X63 commonsourceibias.t63 commonsourceibias.t62 gnd.t92 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X64 a_n2318_13878.t45 minus.t9 a_n3827_n3924.t19 gnd.t171 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X65 a_n7636_8799.t31 a_n2318_13878.t56 a_n2318_8322.t20 vdd.t95 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X66 CSoutput.t143 a_n7636_8799.t49 vdd.t228 vdd.t193 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X67 commonsourceibias.t61 commonsourceibias.t60 gnd.t204 gnd.t95 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X68 vdd.t223 a_n7636_8799.t50 CSoutput.t142 vdd.t129 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X69 vdd.t227 a_n7636_8799.t51 CSoutput.t141 vdd.t205 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X70 gnd.t307 gnd.t304 gnd.t306 gnd.t305 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X71 plus.t3 gnd.t301 gnd.t303 gnd.t302 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X72 diffpairibias.t17 diffpairibias.t16 gnd.t109 gnd.t108 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X73 gnd.t94 commonsourceibias.t58 commonsourceibias.t59 gnd.t93 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X74 CSoutput.t140 a_n7636_8799.t52 vdd.t226 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X75 CSoutput.t30 commonsourceibias.t89 gnd.t115 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X76 gnd.t300 gnd.t298 gnd.t299 gnd.t245 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X77 vdd.t225 a_n7636_8799.t53 CSoutput.t139 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X78 CSoutput.t138 a_n7636_8799.t54 vdd.t222 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X79 CSoutput.t159 commonsourceibias.t90 gnd.t220 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 CSoutput.t137 a_n7636_8799.t55 vdd.t221 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X81 CSoutput.t136 a_n7636_8799.t56 vdd.t220 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X82 CSoutput.t135 a_n7636_8799.t57 vdd.t219 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 gnd.t72 commonsourceibias.t56 commonsourceibias.t57 gnd.t71 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X84 vdd.t1 CSoutput.t179 output.t16 gnd.t17 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X85 CSoutput.t160 commonsourceibias.t91 gnd.t221 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X86 CSoutput.t56 commonsourceibias.t92 gnd.t181 gnd.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X87 a_n3827_n3924.t40 plus.t9 a_n7636_8799.t26 gnd.t124 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X88 CSoutput.t57 commonsourceibias.t93 gnd.t182 gnd.t104 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 CSoutput.t5 commonsourceibias.t94 gnd.t24 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 a_n3827_n3924.t10 diffpairibias.t22 gnd.t60 gnd.t59 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X91 vdd.t218 a_n7636_8799.t58 CSoutput.t134 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X92 a_n2318_13878.t11 a_n2318_13878.t10 a_n2140_13878.t12 vdd.t103 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X93 vdd.t217 a_n7636_8799.t59 CSoutput.t133 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X94 output.t15 CSoutput.t180 vdd.t2 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X95 a_n7636_8799.t32 a_n2318_13878.t57 a_n2318_8322.t19 vdd.t249 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X96 vdd.t216 a_n7636_8799.t60 CSoutput.t132 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X97 a_n2318_13878.t37 a_n2318_13878.t36 a_n2140_13878.t11 vdd.t107 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X98 gnd.t190 commonsourceibias.t54 commonsourceibias.t55 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X99 gnd.t99 commonsourceibias.t52 commonsourceibias.t53 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X100 gnd.t140 commonsourceibias.t50 commonsourceibias.t51 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X101 output.t3 outputibias.t8 gnd.t117 gnd.t116 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X102 CSoutput.t181 a_n2318_8322.t27 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X103 vdd.t215 a_n7636_8799.t61 CSoutput.t131 vdd.t131 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X104 CSoutput.t130 a_n7636_8799.t62 vdd.t214 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X105 gnd.t297 gnd.t294 gnd.t296 gnd.t295 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X106 diffpairibias.t15 diffpairibias.t14 gnd.t217 gnd.t216 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X107 a_n2318_13878.t2 minus.t10 a_n3827_n3924.t2 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X108 output.t2 outputibias.t9 gnd.t168 gnd.t167 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X109 vdd.t75 vdd.t73 vdd.t74 vdd.t63 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X110 vdd.t72 vdd.t70 vdd.t71 vdd.t25 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X111 CSoutput.t129 a_n7636_8799.t63 vdd.t213 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X112 gnd.t26 commonsourceibias.t95 CSoutput.t6 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X113 vdd.t69 vdd.t66 vdd.t68 vdd.t67 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X114 gnd.t179 commonsourceibias.t96 CSoutput.t54 gnd.t90 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X115 gnd.t180 commonsourceibias.t97 CSoutput.t55 gnd.t93 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X116 gnd.t47 commonsourceibias.t98 CSoutput.t11 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X117 a_n3827_n3924.t12 minus.t11 a_n2318_13878.t41 gnd.t112 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X118 gnd.t49 commonsourceibias.t99 CSoutput.t12 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X119 output.t14 CSoutput.t182 vdd.t3 gnd.t41 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X120 vdd.t4 CSoutput.t183 output.t13 gnd.t42 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X121 vdd.t244 a_n2318_13878.t58 a_n2318_8322.t7 vdd.t243 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X122 a_n2318_13878.t19 a_n2318_13878.t18 a_n2140_13878.t10 vdd.t94 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X123 gnd.t12 commonsourceibias.t100 CSoutput.t1 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X124 gnd.t293 gnd.t291 gnd.t292 gnd.t241 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X125 a_n2318_8322.t6 a_n2318_13878.t59 vdd.t246 vdd.t245 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X126 a_n3827_n3924.t3 diffpairibias.t23 gnd.t6 gnd.t5 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X127 CSoutput.t128 a_n7636_8799.t64 vdd.t212 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X128 CSoutput.t127 a_n7636_8799.t65 vdd.t210 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X129 gnd.t290 gnd.t288 gnd.t289 gnd.t252 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X130 CSoutput.t2 commonsourceibias.t101 gnd.t14 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X131 a_n3827_n3924.t7 minus.t12 a_n2318_13878.t6 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X132 gnd.t100 commonsourceibias.t48 commonsourceibias.t49 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X133 vdd.t255 a_n2318_13878.t60 a_n2140_13878.t22 vdd.t254 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X134 a_n2318_13878.t1 minus.t13 a_n3827_n3924.t1 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X135 a_n3827_n3924.t27 plus.t10 a_n7636_8799.t25 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X136 a_n3827_n3924.t31 plus.t11 a_n7636_8799.t24 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X137 gnd.t211 commonsourceibias.t102 CSoutput.t157 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X138 vdd.t65 vdd.t62 vdd.t64 vdd.t63 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X139 vdd.t209 a_n7636_8799.t66 CSoutput.t126 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X140 gnd.t141 commonsourceibias.t46 commonsourceibias.t47 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X141 a_n7636_8799.t23 plus.t12 a_n3827_n3924.t39 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X142 a_n7636_8799.t22 plus.t13 a_n3827_n3924.t45 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X143 vdd.t61 vdd.t58 vdd.t60 vdd.t59 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X144 a_n2318_8322.t5 a_n2318_13878.t61 vdd.t257 vdd.t256 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X145 a_n7636_8799.t8 a_n2318_13878.t62 a_n2318_8322.t18 vdd.t88 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X146 CSoutput.t125 a_n7636_8799.t67 vdd.t207 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X147 diffpairibias.t13 diffpairibias.t12 gnd.t359 gnd.t358 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X148 CSoutput.t184 a_n2318_8322.t25 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X149 vdd.t206 a_n7636_8799.t68 CSoutput.t124 vdd.t205 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X150 CSoutput.t158 commonsourceibias.t103 gnd.t212 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X151 a_n2318_13878.t50 minus.t14 a_n3827_n3924.t25 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X152 a_n2318_13878.t23 a_n2318_13878.t22 a_n2140_13878.t9 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X153 vdd.t204 a_n7636_8799.t69 CSoutput.t123 vdd.t131 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X154 a_n7636_8799.t9 a_n2318_13878.t63 a_n2318_8322.t17 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X155 CSoutput.t122 a_n7636_8799.t70 vdd.t203 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X156 CSoutput.t40 commonsourceibias.t104 gnd.t137 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X157 a_n2140_13878.t8 a_n2318_13878.t16 a_n2318_13878.t17 vdd.t249 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X158 commonsourceibias.t45 commonsourceibias.t44 gnd.t191 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X159 CSoutput.t41 commonsourceibias.t105 gnd.t139 gnd.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X160 gnd.t287 gnd.t285 minus.t4 gnd.t286 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X161 vdd.t57 vdd.t55 vdd.t56 vdd.t25 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X162 gnd.t346 commonsourceibias.t106 CSoutput.t170 gnd.t143 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X163 a_n3827_n3924.t23 minus.t15 a_n2318_13878.t48 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X164 CSoutput.t171 commonsourceibias.t107 gnd.t347 gnd.t104 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 vdd.t5 CSoutput.t185 output.t12 gnd.t43 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X166 CSoutput.t8 commonsourceibias.t108 gnd.t33 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X167 gnd.t174 commonsourceibias.t109 CSoutput.t49 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X168 CSoutput.t121 a_n7636_8799.t71 vdd.t202 vdd.t193 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X169 gnd.t192 commonsourceibias.t42 commonsourceibias.t43 gnd.t128 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X170 vdd.t251 a_n2318_13878.t64 a_n2318_8322.t4 vdd.t250 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X171 a_n2140_13878.t7 a_n2318_13878.t8 a_n2318_13878.t9 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X172 gnd.t113 commonsourceibias.t110 CSoutput.t28 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X173 vdd.t201 a_n7636_8799.t72 CSoutput.t120 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X174 a_n2318_13878.t33 a_n2318_13878.t32 a_n2140_13878.t6 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X175 commonsourceibias.t41 commonsourceibias.t40 gnd.t101 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X176 gnd.t74 commonsourceibias.t38 commonsourceibias.t39 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X177 a_n3827_n3924.t43 plus.t14 a_n7636_8799.t21 gnd.t118 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X178 gnd.t284 gnd.t282 minus.t3 gnd.t283 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X179 vdd.t200 a_n7636_8799.t73 CSoutput.t119 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X180 gnd.t193 commonsourceibias.t36 commonsourceibias.t37 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X181 a_n3827_n3924.t9 diffpairibias.t24 gnd.t45 gnd.t44 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X182 commonsourceibias.t35 commonsourceibias.t34 gnd.t102 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X183 a_n3827_n3924.t17 diffpairibias.t25 gnd.t152 gnd.t151 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X184 gnd.t135 commonsourceibias.t111 CSoutput.t39 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X185 vdd.t199 a_n7636_8799.t74 CSoutput.t118 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X186 vdd.t198 a_n7636_8799.t75 CSoutput.t117 vdd.t152 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X187 a_n7636_8799.t20 plus.t15 a_n3827_n3924.t34 gnd.t85 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X188 gnd.t178 commonsourceibias.t112 CSoutput.t53 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X189 gnd.t177 commonsourceibias.t113 CSoutput.t52 gnd.t93 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X190 gnd.t134 commonsourceibias.t114 CSoutput.t38 gnd.t90 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X191 gnd.t133 commonsourceibias.t115 CSoutput.t37 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X192 CSoutput.t186 a_n2318_8322.t26 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X193 CSoutput.t36 commonsourceibias.t116 gnd.t132 gnd.t131 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X194 CSoutput.t116 a_n7636_8799.t76 vdd.t192 vdd.t115 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X195 commonsourceibias.t33 commonsourceibias.t32 gnd.t142 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 CSoutput.t35 commonsourceibias.t117 gnd.t130 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X197 CSoutput.t115 a_n7636_8799.t77 vdd.t197 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X198 CSoutput.t114 a_n7636_8799.t78 vdd.t195 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X199 CSoutput.t187 a_n2318_8322.t26 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X200 gnd.t338 commonsourceibias.t118 CSoutput.t167 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X201 CSoutput.t166 commonsourceibias.t119 gnd.t337 gnd.t145 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X202 gnd.t281 gnd.t279 gnd.t280 gnd.t223 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X203 diffpairibias.t11 diffpairibias.t10 gnd.t219 gnd.t218 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X204 a_n2140_13878.t21 a_n2318_13878.t65 vdd.t253 vdd.t252 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X205 gnd.t336 commonsourceibias.t120 CSoutput.t165 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X206 vdd.t248 a_n2318_13878.t66 a_n2140_13878.t20 vdd.t247 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X207 output.t1 outputibias.t10 gnd.t40 gnd.t39 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X208 vdd.t54 vdd.t52 vdd.t53 vdd.t42 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X209 gnd.t194 commonsourceibias.t30 commonsourceibias.t31 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X210 CSoutput.t113 a_n7636_8799.t79 vdd.t194 vdd.t193 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X211 gnd.t144 commonsourceibias.t28 commonsourceibias.t29 gnd.t143 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X212 vdd.t191 a_n7636_8799.t80 CSoutput.t112 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X213 commonsourceibias.t27 commonsourceibias.t26 gnd.t38 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X214 vdd.t51 vdd.t49 vdd.t50 vdd.t42 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X215 CSoutput.t161 commonsourceibias.t121 gnd.t332 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X216 a_n2140_13878.t5 a_n2318_13878.t38 a_n2318_13878.t39 vdd.t95 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X217 diffpairibias.t9 diffpairibias.t8 gnd.t206 gnd.t205 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X218 a_n3827_n3924.t5 minus.t16 a_n2318_13878.t4 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X219 vdd.t189 a_n7636_8799.t81 CSoutput.t111 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X220 gnd.t103 commonsourceibias.t24 commonsourceibias.t25 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X221 CSoutput.t164 commonsourceibias.t122 gnd.t335 gnd.t106 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X222 a_n2318_8322.t16 a_n2318_13878.t67 a_n7636_8799.t10 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X223 CSoutput.t110 a_n7636_8799.t82 vdd.t188 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X224 diffpairibias.t7 diffpairibias.t6 gnd.t111 gnd.t110 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X225 vdd.t187 a_n7636_8799.t83 CSoutput.t109 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X226 a_n2318_13878.t5 minus.t17 a_n3827_n3924.t6 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X227 a_n2318_13878.t0 minus.t18 a_n3827_n3924.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X228 gnd.t334 commonsourceibias.t123 CSoutput.t163 gnd.t143 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X229 plus.t0 gnd.t276 gnd.t278 gnd.t277 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X230 vdd.t259 a_n2318_13878.t68 a_n2318_8322.t3 vdd.t258 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X231 vdd.t185 a_n7636_8799.t84 CSoutput.t108 vdd.t152 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X232 vdd.t182 a_n7636_8799.t85 CSoutput.t107 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X233 vdd.t241 CSoutput.t188 output.t11 gnd.t214 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X234 CSoutput.t44 commonsourceibias.t124 gnd.t164 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 a_n7636_8799.t19 plus.t16 a_n3827_n3924.t30 gnd.t171 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X236 CSoutput.t162 commonsourceibias.t125 gnd.t333 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X237 gnd.t275 gnd.t272 gnd.t274 gnd.t273 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X238 gnd.t271 gnd.t269 minus.t2 gnd.t270 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X239 gnd.t81 commonsourceibias.t126 CSoutput.t22 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X240 a_n3827_n3924.t24 minus.t19 a_n2318_13878.t49 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X241 gnd.t268 gnd.t265 gnd.t267 gnd.t266 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X242 gnd.t70 commonsourceibias.t127 CSoutput.t18 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X243 a_n2140_13878.t19 a_n2318_13878.t69 vdd.t261 vdd.t260 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X244 CSoutput.t21 commonsourceibias.t128 gnd.t79 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X245 commonsourceibias.t23 commonsourceibias.t22 gnd.t105 gnd.t104 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X246 CSoutput.t17 commonsourceibias.t129 gnd.t68 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X247 vdd.t184 a_n7636_8799.t86 CSoutput.t106 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X248 CSoutput.t105 a_n7636_8799.t87 vdd.t183 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X249 CSoutput.t104 a_n7636_8799.t88 vdd.t180 vdd.t162 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X250 gnd.t264 gnd.t262 gnd.t263 gnd.t241 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X251 vdd.t48 vdd.t45 vdd.t47 vdd.t46 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X252 minus.t1 gnd.t259 gnd.t261 gnd.t260 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X253 a_n3827_n3924.t16 diffpairibias.t26 gnd.t150 gnd.t149 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X254 vdd.t44 vdd.t41 vdd.t43 vdd.t42 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X255 vdd.t263 a_n2318_13878.t70 a_n2318_8322.t2 vdd.t262 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X256 a_n2318_8322.t15 a_n2318_13878.t71 a_n7636_8799.t33 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X257 CSoutput.t103 a_n7636_8799.t89 vdd.t179 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X258 gnd.t78 commonsourceibias.t130 CSoutput.t20 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X259 vdd.t177 a_n7636_8799.t90 CSoutput.t102 vdd.t113 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X260 CSoutput.t101 a_n7636_8799.t91 vdd.t176 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X261 vdd.t175 a_n7636_8799.t92 CSoutput.t100 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X262 vdd.t174 a_n7636_8799.t93 CSoutput.t99 vdd.t125 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X263 a_n7636_8799.t18 plus.t17 a_n3827_n3924.t28 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X264 gnd.t67 commonsourceibias.t131 CSoutput.t16 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X265 CSoutput.t45 commonsourceibias.t132 gnd.t165 gnd.t95 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X266 vdd.t40 vdd.t38 vdd.t39 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X267 vdd.t37 vdd.t34 vdd.t36 vdd.t35 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X268 CSoutput.t46 commonsourceibias.t133 gnd.t166 gnd.t131 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X269 a_n3827_n3924.t32 plus.t18 a_n7636_8799.t17 gnd.t29 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X270 vdd.t173 a_n7636_8799.t94 CSoutput.t98 vdd.t119 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X271 CSoutput.t97 a_n7636_8799.t95 vdd.t172 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X272 gnd.t159 commonsourceibias.t134 CSoutput.t42 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X273 gnd.t201 commonsourceibias.t135 CSoutput.t60 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X274 a_n2140_13878.t4 a_n2318_13878.t34 a_n2318_13878.t35 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X275 CSoutput.t96 a_n7636_8799.t96 vdd.t167 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X276 vdd.t242 CSoutput.t189 output.t10 gnd.t215 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X277 CSoutput.t59 commonsourceibias.t136 gnd.t200 gnd.t145 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 a_n2318_8322.t14 a_n2318_13878.t72 a_n7636_8799.t34 vdd.t111 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X279 diffpairibias.t5 diffpairibias.t4 gnd.t120 gnd.t119 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X280 commonsourceibias.t21 commonsourceibias.t20 gnd.t146 gnd.t145 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X281 gnd.t258 gnd.t255 gnd.t257 gnd.t256 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X282 gnd.t199 commonsourceibias.t137 CSoutput.t58 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X283 CSoutput.t169 commonsourceibias.t138 gnd.t345 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X284 gnd.t195 commonsourceibias.t18 commonsourceibias.t19 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X285 CSoutput.t95 a_n7636_8799.t97 vdd.t170 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X286 CSoutput.t94 a_n7636_8799.t98 vdd.t166 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X287 a_n3827_n3924.t49 diffpairibias.t27 gnd.t355 gnd.t354 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X288 vdd.t168 a_n7636_8799.t99 CSoutput.t93 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X289 CSoutput.t175 commonsourceibias.t139 gnd.t357 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X290 CSoutput.t190 a_n2318_8322.t25 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X291 vdd.t165 a_n7636_8799.t100 CSoutput.t92 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X292 a_n2318_8322.t1 a_n2318_13878.t73 vdd.t265 vdd.t264 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X293 CSoutput.t91 a_n7636_8799.t101 vdd.t163 vdd.t162 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X294 CSoutput.t48 commonsourceibias.t140 gnd.t173 gnd.t106 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X295 vdd.t33 vdd.t31 vdd.t32 vdd.t17 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X296 vdd.t267 a_n2318_13878.t74 a_n2140_13878.t18 vdd.t266 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X297 gnd.t196 commonsourceibias.t16 commonsourceibias.t17 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X298 output.t0 outputibias.t11 gnd.t4 gnd.t3 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X299 CSoutput.t90 a_n7636_8799.t102 vdd.t161 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X300 CSoutput.t43 commonsourceibias.t141 gnd.t160 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X301 CSoutput.t89 a_n7636_8799.t103 vdd.t159 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X302 gnd.t129 commonsourceibias.t142 CSoutput.t34 gnd.t128 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X303 gnd.t254 gnd.t251 gnd.t253 gnd.t252 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X304 vdd.t158 a_n7636_8799.t104 CSoutput.t88 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X305 vdd.t156 a_n7636_8799.t105 CSoutput.t87 vdd.t125 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X306 CSoutput.t15 commonsourceibias.t143 gnd.t66 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 minus.t0 gnd.t248 gnd.t250 gnd.t249 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X308 vdd.t30 vdd.t28 vdd.t29 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X309 commonsourceibias.t15 commonsourceibias.t14 gnd.t107 gnd.t106 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X310 a_n3827_n3924.t22 minus.t20 a_n2318_13878.t47 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X311 commonsourceibias.t13 commonsourceibias.t12 gnd.t147 gnd.t131 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X312 a_n2318_8322.t13 a_n2318_13878.t75 a_n7636_8799.t35 vdd.t93 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X313 CSoutput.t86 a_n7636_8799.t106 vdd.t155 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X314 CSoutput.t33 commonsourceibias.t144 gnd.t127 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X315 a_n7636_8799.t3 a_n2318_13878.t76 a_n2318_8322.t12 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X316 gnd.t198 commonsourceibias.t10 commonsourceibias.t11 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X317 output.t9 CSoutput.t191 vdd.t90 gnd.t88 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X318 vdd.t153 a_n7636_8799.t107 CSoutput.t85 vdd.t152 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X319 a_n2140_13878.t17 a_n2318_13878.t77 vdd.t102 vdd.t101 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X320 gnd.t98 commonsourceibias.t145 CSoutput.t27 gnd.t97 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X321 CSoutput.t4 commonsourceibias.t146 gnd.t22 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X322 gnd.t247 gnd.t244 gnd.t246 gnd.t245 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X323 vdd.t151 a_n7636_8799.t108 CSoutput.t84 vdd.t129 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X324 a_n2318_13878.t46 minus.t21 a_n3827_n3924.t21 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X325 CSoutput.t83 a_n7636_8799.t109 vdd.t145 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X326 gnd.t243 gnd.t240 gnd.t242 gnd.t241 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X327 commonsourceibias.t9 commonsourceibias.t8 gnd.t148 gnd.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X328 a_n7636_8799.t16 plus.t19 a_n3827_n3924.t41 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X329 a_n2318_8322.t11 a_n2318_13878.t78 a_n7636_8799.t0 vdd.t94 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X330 a_n3827_n3924.t15 minus.t22 a_n2318_13878.t44 gnd.t124 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X331 vdd.t150 a_n7636_8799.t110 CSoutput.t82 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X332 CSoutput.t81 a_n7636_8799.t111 vdd.t148 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X333 CSoutput.t80 a_n7636_8799.t112 vdd.t146 vdd.t127 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X334 gnd.t213 commonsourceibias.t6 commonsourceibias.t7 gnd.t97 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X335 CSoutput.t79 a_n7636_8799.t113 vdd.t143 vdd.t127 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X336 a_n2140_13878.t3 a_n2318_13878.t30 a_n2318_13878.t31 vdd.t88 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X337 commonsourceibias.t5 commonsourceibias.t4 gnd.t52 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X338 a_n3827_n3924.t33 plus.t20 a_n7636_8799.t15 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X339 vdd.t142 a_n7636_8799.t114 CSoutput.t78 vdd.t123 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X340 gnd.t64 commonsourceibias.t147 CSoutput.t14 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X341 CSoutput.t26 commonsourceibias.t148 gnd.t96 gnd.t95 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X342 vdd.t27 vdd.t24 vdd.t26 vdd.t25 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X343 CSoutput.t192 a_n2318_8322.t24 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X344 vdd.t23 vdd.t20 vdd.t22 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X345 output.t8 CSoutput.t193 vdd.t91 gnd.t89 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X346 gnd.t31 commonsourceibias.t149 CSoutput.t7 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X347 a_n3827_n3924.t48 diffpairibias.t28 gnd.t351 gnd.t350 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X348 vdd.t141 a_n7636_8799.t115 CSoutput.t77 vdd.t119 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X349 vdd.t140 a_n7636_8799.t116 CSoutput.t76 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X350 gnd.t76 commonsourceibias.t150 CSoutput.t19 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X351 CSoutput.t75 a_n7636_8799.t117 vdd.t139 vdd.t115 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X352 a_n2318_13878.t21 a_n2318_13878.t20 a_n2140_13878.t2 vdd.t93 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X353 gnd.t239 gnd.t236 gnd.t238 gnd.t237 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X354 a_n7636_8799.t1 a_n2318_13878.t79 a_n2318_8322.t10 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X355 vdd.t138 a_n7636_8799.t118 CSoutput.t74 vdd.t123 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X356 output.t7 CSoutput.t194 vdd.t6 gnd.t53 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X357 gnd.t62 commonsourceibias.t151 CSoutput.t13 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X358 CSoutput.t73 a_n7636_8799.t119 vdd.t137 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X359 a_n7636_8799.t14 plus.t21 a_n3827_n3924.t42 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X360 vdd.t7 CSoutput.t195 output.t6 gnd.t54 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X361 vdd.t135 a_n7636_8799.t120 CSoutput.t72 vdd.t113 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X362 gnd.t235 gnd.t232 gnd.t234 gnd.t233 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X363 CSoutput.t3 commonsourceibias.t152 gnd.t20 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X364 CSoutput.t25 commonsourceibias.t153 gnd.t87 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X365 commonsourceibias.t3 commonsourceibias.t2 gnd.t163 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X366 gnd.t231 gnd.t229 plus.t2 gnd.t230 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X367 outputibias.t5 outputibias.t4 gnd.t341 gnd.t340 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X368 diffpairibias.t3 diffpairibias.t2 gnd.t353 gnd.t352 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X369 vdd.t132 a_n7636_8799.t121 CSoutput.t71 vdd.t131 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X370 CSoutput.t70 a_n7636_8799.t122 vdd.t134 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X371 a_n2318_8322.t9 a_n2318_13878.t80 a_n7636_8799.t2 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X372 a_n3827_n3924.t44 plus.t22 a_n7636_8799.t13 gnd.t112 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X373 gnd.t228 gnd.t226 plus.t1 gnd.t227 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X374 vdd.t130 a_n7636_8799.t123 CSoutput.t69 vdd.t129 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X375 outputibias.t3 outputibias.t2 gnd.t331 gnd.t330 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X376 diffpairibias.t1 diffpairibias.t0 gnd.t156 gnd.t155 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X377 a_n3827_n3924.t29 plus.t23 a_n7636_8799.t12 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X378 CSoutput.t0 commonsourceibias.t154 gnd.t10 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X379 outputibias.t1 outputibias.t0 gnd.t158 gnd.t157 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X380 vdd.t19 vdd.t16 vdd.t18 vdd.t17 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X381 vdd.t99 a_n2318_13878.t81 a_n2140_13878.t16 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X382 gnd.t344 commonsourceibias.t155 CSoutput.t168 gnd.t128 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X383 a_n7636_8799.t11 plus.t24 a_n3827_n3924.t46 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X384 CSoutput.t68 a_n7636_8799.t124 vdd.t128 vdd.t127 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X385 vdd.t15 vdd.t12 vdd.t14 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X386 a_n3827_n3924.t4 minus.t23 a_n2318_13878.t3 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X387 vdd.t126 a_n7636_8799.t125 CSoutput.t67 vdd.t125 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X388 vdd.t124 a_n7636_8799.t126 CSoutput.t66 vdd.t123 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X389 CSoutput.t174 commonsourceibias.t156 gnd.t356 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X390 CSoutput.t65 a_n7636_8799.t127 vdd.t122 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X391 output.t5 CSoutput.t196 vdd.t8 gnd.t55 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X392 gnd.t172 commonsourceibias.t157 CSoutput.t47 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X393 gnd.t225 gnd.t222 gnd.t224 gnd.t223 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X394 a_n2318_13878.t43 minus.t24 a_n3827_n3924.t14 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X395 gnd.t126 commonsourceibias.t158 CSoutput.t32 gnd.t97 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X396 a_n2318_8322.t8 a_n2318_13878.t82 a_n7636_8799.t5 vdd.t107 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X397 vdd.t120 a_n7636_8799.t128 CSoutput.t64 vdd.t119 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X398 vdd.t118 a_n7636_8799.t129 CSoutput.t63 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X399 CSoutput.t62 a_n7636_8799.t130 vdd.t116 vdd.t115 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X400 output.t4 CSoutput.t197 vdd.t9 gnd.t56 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X401 gnd.t125 commonsourceibias.t159 CSoutput.t31 gnd.t71 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X402 a_n2318_8322.t0 a_n2318_13878.t83 vdd.t109 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X403 a_n2140_13878.t1 a_n2318_13878.t28 a_n2318_13878.t29 vdd.t112 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X404 vdd.t114 a_n7636_8799.t131 CSoutput.t61 vdd.t113 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X405 commonsourceibias.t1 commonsourceibias.t0 gnd.t161 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X406 a_n3827_n3924.t47 diffpairibias.t29 gnd.t343 gnd.t342 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X407 a_n2318_13878.t25 a_n2318_13878.t24 a_n2140_13878.t0 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 plus.n43 plus.t18 322.512
R1 plus.n9 plus.t13 322.512
R2 plus.n42 plus.t17 297.12
R3 plus.n46 plus.t22 297.12
R4 plus.n48 plus.t21 297.12
R5 plus.n52 plus.t23 297.12
R6 plus.n54 plus.t8 297.12
R7 plus.n58 plus.t7 297.12
R8 plus.n60 plus.t12 297.12
R9 plus.n64 plus.t10 297.12
R10 plus.n66 plus.t24 297.12
R11 plus.n32 plus.t14 297.12
R12 plus.n30 plus.t15 297.12
R13 plus.n2 plus.t9 297.12
R14 plus.n24 plus.t5 297.12
R15 plus.n4 plus.t6 297.12
R16 plus.n18 plus.t19 297.12
R17 plus.n6 plus.t20 297.12
R18 plus.n12 plus.t16 297.12
R19 plus.n8 plus.t11 297.12
R20 plus.n70 plus.t1 243.97
R21 plus.n70 plus.n69 223.454
R22 plus.n72 plus.n71 223.454
R23 plus.n67 plus.n66 161.3
R24 plus.n65 plus.n34 161.3
R25 plus.n64 plus.n63 161.3
R26 plus.n62 plus.n35 161.3
R27 plus.n61 plus.n60 161.3
R28 plus.n59 plus.n36 161.3
R29 plus.n58 plus.n57 161.3
R30 plus.n56 plus.n37 161.3
R31 plus.n55 plus.n54 161.3
R32 plus.n53 plus.n38 161.3
R33 plus.n52 plus.n51 161.3
R34 plus.n50 plus.n39 161.3
R35 plus.n49 plus.n48 161.3
R36 plus.n47 plus.n40 161.3
R37 plus.n46 plus.n45 161.3
R38 plus.n44 plus.n41 161.3
R39 plus.n11 plus.n10 161.3
R40 plus.n12 plus.n7 161.3
R41 plus.n14 plus.n13 161.3
R42 plus.n15 plus.n6 161.3
R43 plus.n17 plus.n16 161.3
R44 plus.n18 plus.n5 161.3
R45 plus.n20 plus.n19 161.3
R46 plus.n21 plus.n4 161.3
R47 plus.n23 plus.n22 161.3
R48 plus.n24 plus.n3 161.3
R49 plus.n26 plus.n25 161.3
R50 plus.n27 plus.n2 161.3
R51 plus.n29 plus.n28 161.3
R52 plus.n30 plus.n1 161.3
R53 plus.n31 plus.n0 161.3
R54 plus.n33 plus.n32 161.3
R55 plus.n44 plus.n43 45.0031
R56 plus.n10 plus.n9 45.0031
R57 plus.n66 plus.n65 41.6278
R58 plus.n32 plus.n31 41.6278
R59 plus.n42 plus.n41 37.246
R60 plus.n64 plus.n35 37.246
R61 plus.n30 plus.n29 37.246
R62 plus.n11 plus.n8 37.246
R63 plus.n47 plus.n46 32.8641
R64 plus.n60 plus.n59 32.8641
R65 plus.n25 plus.n2 32.8641
R66 plus.n13 plus.n12 32.8641
R67 plus.n68 plus.n67 31.6047
R68 plus.n48 plus.n39 28.4823
R69 plus.n58 plus.n37 28.4823
R70 plus.n24 plus.n23 28.4823
R71 plus.n17 plus.n6 28.4823
R72 plus.n53 plus.n52 24.1005
R73 plus.n54 plus.n53 24.1005
R74 plus.n19 plus.n4 24.1005
R75 plus.n19 plus.n18 24.1005
R76 plus.n69 plus.t4 19.8005
R77 plus.n69 plus.t0 19.8005
R78 plus.n71 plus.t2 19.8005
R79 plus.n71 plus.t3 19.8005
R80 plus.n52 plus.n39 19.7187
R81 plus.n54 plus.n37 19.7187
R82 plus.n23 plus.n4 19.7187
R83 plus.n18 plus.n17 19.7187
R84 plus.n43 plus.n42 15.6319
R85 plus.n9 plus.n8 15.6319
R86 plus.n48 plus.n47 15.3369
R87 plus.n59 plus.n58 15.3369
R88 plus.n25 plus.n24 15.3369
R89 plus.n13 plus.n6 15.3369
R90 plus plus.n73 15.0665
R91 plus.n68 plus.n33 11.866
R92 plus.n46 plus.n41 10.955
R93 plus.n60 plus.n35 10.955
R94 plus.n29 plus.n2 10.955
R95 plus.n12 plus.n11 10.955
R96 plus.n65 plus.n64 6.57323
R97 plus.n31 plus.n30 6.57323
R98 plus.n73 plus.n72 5.40567
R99 plus.n73 plus.n68 1.188
R100 plus.n72 plus.n70 0.716017
R101 plus.n45 plus.n44 0.189894
R102 plus.n45 plus.n40 0.189894
R103 plus.n49 plus.n40 0.189894
R104 plus.n50 plus.n49 0.189894
R105 plus.n51 plus.n50 0.189894
R106 plus.n51 plus.n38 0.189894
R107 plus.n55 plus.n38 0.189894
R108 plus.n56 plus.n55 0.189894
R109 plus.n57 plus.n56 0.189894
R110 plus.n57 plus.n36 0.189894
R111 plus.n61 plus.n36 0.189894
R112 plus.n62 plus.n61 0.189894
R113 plus.n63 plus.n62 0.189894
R114 plus.n63 plus.n34 0.189894
R115 plus.n67 plus.n34 0.189894
R116 plus.n33 plus.n0 0.189894
R117 plus.n1 plus.n0 0.189894
R118 plus.n28 plus.n1 0.189894
R119 plus.n28 plus.n27 0.189894
R120 plus.n27 plus.n26 0.189894
R121 plus.n26 plus.n3 0.189894
R122 plus.n22 plus.n3 0.189894
R123 plus.n22 plus.n21 0.189894
R124 plus.n21 plus.n20 0.189894
R125 plus.n20 plus.n5 0.189894
R126 plus.n16 plus.n5 0.189894
R127 plus.n16 plus.n15 0.189894
R128 plus.n15 plus.n14 0.189894
R129 plus.n14 plus.n7 0.189894
R130 plus.n10 plus.n7 0.189894
R131 a_n3827_n3924.n9 a_n3827_n3924.t49 214.994
R132 a_n3827_n3924.n10 a_n3827_n3924.t18 214.994
R133 a_n3827_n3924.n9 a_n3827_n3924.t3 214.321
R134 a_n3827_n3924.n9 a_n3827_n3924.t48 214.321
R135 a_n3827_n3924.n7 a_n3827_n3924.t17 214.321
R136 a_n3827_n3924.n7 a_n3827_n3924.t47 214.321
R137 a_n3827_n3924.n8 a_n3827_n3924.t9 214.321
R138 a_n3827_n3924.n8 a_n3827_n3924.t20 214.321
R139 a_n3827_n3924.n10 a_n3827_n3924.t10 214.321
R140 a_n3827_n3924.n10 a_n3827_n3924.t16 214.321
R141 a_n3827_n3924.n1 a_n3827_n3924.t32 55.8337
R142 a_n3827_n3924.n1 a_n3827_n3924.t14 55.8337
R143 a_n3827_n3924.n3 a_n3827_n3924.t13 55.8337
R144 a_n3827_n3924.n0 a_n3827_n3924.t46 55.8335
R145 a_n3827_n3924.n5 a_n3827_n3924.t1 55.8335
R146 a_n3827_n3924.n4 a_n3827_n3924.t8 55.8335
R147 a_n3827_n3924.n4 a_n3827_n3924.t45 55.8335
R148 a_n3827_n3924.n6 a_n3827_n3924.t43 55.8335
R149 a_n3827_n3924.n0 a_n3827_n3924.n22 53.0052
R150 a_n3827_n3924.n1 a_n3827_n3924.n23 53.0052
R151 a_n3827_n3924.n1 a_n3827_n3924.n24 53.0052
R152 a_n3827_n3924.n1 a_n3827_n3924.n25 53.0052
R153 a_n3827_n3924.n2 a_n3827_n3924.n26 53.0052
R154 a_n3827_n3924.n2 a_n3827_n3924.n27 53.0052
R155 a_n3827_n3924.n3 a_n3827_n3924.n11 53.0052
R156 a_n3827_n3924.n5 a_n3827_n3924.n20 53.0051
R157 a_n3827_n3924.n5 a_n3827_n3924.n19 53.0051
R158 a_n3827_n3924.n5 a_n3827_n3924.n18 53.0051
R159 a_n3827_n3924.n4 a_n3827_n3924.n17 53.0051
R160 a_n3827_n3924.n4 a_n3827_n3924.n16 53.0051
R161 a_n3827_n3924.n4 a_n3827_n3924.n15 53.0051
R162 a_n3827_n3924.n4 a_n3827_n3924.n14 53.0051
R163 a_n3827_n3924.n6 a_n3827_n3924.n13 53.0051
R164 a_n3827_n3924.n28 a_n3827_n3924.n3 53.0051
R165 a_n3827_n3924.n12 a_n3827_n3924.n3 12.1986
R166 a_n3827_n3924.n0 a_n3827_n3924.n21 12.1986
R167 a_n3827_n3924.n6 a_n3827_n3924.n12 5.11903
R168 a_n3827_n3924.n21 a_n3827_n3924.n5 5.11903
R169 a_n3827_n3924.n22 a_n3827_n3924.t39 2.82907
R170 a_n3827_n3924.n22 a_n3827_n3924.t27 2.82907
R171 a_n3827_n3924.n23 a_n3827_n3924.t35 2.82907
R172 a_n3827_n3924.n23 a_n3827_n3924.t36 2.82907
R173 a_n3827_n3924.n24 a_n3827_n3924.t42 2.82907
R174 a_n3827_n3924.n24 a_n3827_n3924.t29 2.82907
R175 a_n3827_n3924.n25 a_n3827_n3924.t28 2.82907
R176 a_n3827_n3924.n25 a_n3827_n3924.t44 2.82907
R177 a_n3827_n3924.n26 a_n3827_n3924.t19 2.82907
R178 a_n3827_n3924.n26 a_n3827_n3924.t4 2.82907
R179 a_n3827_n3924.n27 a_n3827_n3924.t25 2.82907
R180 a_n3827_n3924.n27 a_n3827_n3924.t23 2.82907
R181 a_n3827_n3924.n11 a_n3827_n3924.t11 2.82907
R182 a_n3827_n3924.n11 a_n3827_n3924.t15 2.82907
R183 a_n3827_n3924.n20 a_n3827_n3924.t21 2.82907
R184 a_n3827_n3924.n20 a_n3827_n3924.t22 2.82907
R185 a_n3827_n3924.n19 a_n3827_n3924.t6 2.82907
R186 a_n3827_n3924.n19 a_n3827_n3924.t5 2.82907
R187 a_n3827_n3924.n18 a_n3827_n3924.t2 2.82907
R188 a_n3827_n3924.n18 a_n3827_n3924.t7 2.82907
R189 a_n3827_n3924.n17 a_n3827_n3924.t26 2.82907
R190 a_n3827_n3924.n17 a_n3827_n3924.t12 2.82907
R191 a_n3827_n3924.n16 a_n3827_n3924.t30 2.82907
R192 a_n3827_n3924.n16 a_n3827_n3924.t31 2.82907
R193 a_n3827_n3924.n15 a_n3827_n3924.t41 2.82907
R194 a_n3827_n3924.n15 a_n3827_n3924.t33 2.82907
R195 a_n3827_n3924.n14 a_n3827_n3924.t37 2.82907
R196 a_n3827_n3924.n14 a_n3827_n3924.t38 2.82907
R197 a_n3827_n3924.n13 a_n3827_n3924.t34 2.82907
R198 a_n3827_n3924.n13 a_n3827_n3924.t40 2.82907
R199 a_n3827_n3924.t0 a_n3827_n3924.n28 2.82907
R200 a_n3827_n3924.n28 a_n3827_n3924.t24 2.82907
R201 a_n3827_n3924.n5 a_n3827_n3924.n4 2.45524
R202 a_n3827_n3924.n4 a_n3827_n3924.n6 2.22033
R203 a_n3827_n3924.n10 a_n3827_n3924.n8 2.01503
R204 a_n3827_n3924.n21 a_n3827_n3924.n9 1.95694
R205 a_n3827_n3924.n12 a_n3827_n3924.n10 1.95694
R206 a_n3827_n3924.n3 a_n3827_n3924.n2 1.77636
R207 a_n3827_n3924.n1 a_n3827_n3924.n0 1.77636
R208 a_n3827_n3924.n8 a_n3827_n3924.n7 1.34352
R209 a_n3827_n3924.n7 a_n3827_n3924.n9 1.34352
R210 a_n3827_n3924.n2 a_n3827_n3924.n1 1.12334
R211 a_n7636_8799.n176 a_n7636_8799.t56 485.149
R212 a_n7636_8799.n224 a_n7636_8799.t65 485.149
R213 a_n7636_8799.n273 a_n7636_8799.t95 485.149
R214 a_n7636_8799.n28 a_n7636_8799.t115 485.149
R215 a_n7636_8799.n76 a_n7636_8799.t128 485.149
R216 a_n7636_8799.n125 a_n7636_8799.t94 485.149
R217 a_n7636_8799.n208 a_n7636_8799.t75 464.166
R218 a_n7636_8799.n207 a_n7636_8799.t57 464.166
R219 a_n7636_8799.n163 a_n7636_8799.t120 464.166
R220 a_n7636_8799.n201 a_n7636_8799.t88 464.166
R221 a_n7636_8799.n200 a_n7636_8799.t86 464.166
R222 a_n7636_8799.n166 a_n7636_8799.t38 464.166
R223 a_n7636_8799.n194 a_n7636_8799.t92 464.166
R224 a_n7636_8799.n193 a_n7636_8799.t91 464.166
R225 a_n7636_8799.n169 a_n7636_8799.t40 464.166
R226 a_n7636_8799.n188 a_n7636_8799.t39 464.166
R227 a_n7636_8799.n186 a_n7636_8799.t108 464.166
R228 a_n7636_8799.n172 a_n7636_8799.t52 464.166
R229 a_n7636_8799.n181 a_n7636_8799.t43 464.166
R230 a_n7636_8799.n179 a_n7636_8799.t112 464.166
R231 a_n7636_8799.n175 a_n7636_8799.t74 464.166
R232 a_n7636_8799.n256 a_n7636_8799.t84 464.166
R233 a_n7636_8799.n255 a_n7636_8799.t64 464.166
R234 a_n7636_8799.n211 a_n7636_8799.t131 464.166
R235 a_n7636_8799.n249 a_n7636_8799.t101 464.166
R236 a_n7636_8799.n248 a_n7636_8799.t100 464.166
R237 a_n7636_8799.n214 a_n7636_8799.t46 464.166
R238 a_n7636_8799.n242 a_n7636_8799.t104 464.166
R239 a_n7636_8799.n241 a_n7636_8799.t103 464.166
R240 a_n7636_8799.n217 a_n7636_8799.t48 464.166
R241 a_n7636_8799.n236 a_n7636_8799.t47 464.166
R242 a_n7636_8799.n234 a_n7636_8799.t123 464.166
R243 a_n7636_8799.n220 a_n7636_8799.t63 464.166
R244 a_n7636_8799.n229 a_n7636_8799.t51 464.166
R245 a_n7636_8799.n227 a_n7636_8799.t124 464.166
R246 a_n7636_8799.n223 a_n7636_8799.t85 464.166
R247 a_n7636_8799.n305 a_n7636_8799.t107 464.166
R248 a_n7636_8799.n304 a_n7636_8799.t54 464.166
R249 a_n7636_8799.n260 a_n7636_8799.t90 464.166
R250 a_n7636_8799.n298 a_n7636_8799.t42 464.166
R251 a_n7636_8799.n297 a_n7636_8799.t59 464.166
R252 a_n7636_8799.n263 a_n7636_8799.t127 464.166
R253 a_n7636_8799.n291 a_n7636_8799.t99 464.166
R254 a_n7636_8799.n290 a_n7636_8799.t122 464.166
R255 a_n7636_8799.n266 a_n7636_8799.t83 464.166
R256 a_n7636_8799.n285 a_n7636_8799.t102 464.166
R257 a_n7636_8799.n283 a_n7636_8799.t50 464.166
R258 a_n7636_8799.n269 a_n7636_8799.t119 464.166
R259 a_n7636_8799.n278 a_n7636_8799.t68 464.166
R260 a_n7636_8799.n276 a_n7636_8799.t113 464.166
R261 a_n7636_8799.n272 a_n7636_8799.t58 464.166
R262 a_n7636_8799.n27 a_n7636_8799.t117 464.166
R263 a_n7636_8799.n31 a_n7636_8799.t73 464.166
R264 a_n7636_8799.n25 a_n7636_8799.t98 464.166
R265 a_n7636_8799.n36 a_n7636_8799.t114 464.166
R266 a_n7636_8799.n38 a_n7636_8799.t71 464.166
R267 a_n7636_8799.n42 a_n7636_8799.t72 464.166
R268 a_n7636_8799.n43 a_n7636_8799.t96 464.166
R269 a_n7636_8799.n21 a_n7636_8799.t61 464.166
R270 a_n7636_8799.n48 a_n7636_8799.t62 464.166
R271 a_n7636_8799.n50 a_n7636_8799.t93 464.166
R272 a_n7636_8799.n54 a_n7636_8799.t36 464.166
R273 a_n7636_8799.n55 a_n7636_8799.t60 464.166
R274 a_n7636_8799.n17 a_n7636_8799.t78 464.166
R275 a_n7636_8799.n61 a_n7636_8799.t116 464.166
R276 a_n7636_8799.n62 a_n7636_8799.t45 464.166
R277 a_n7636_8799.n75 a_n7636_8799.t130 464.166
R278 a_n7636_8799.n79 a_n7636_8799.t81 464.166
R279 a_n7636_8799.n73 a_n7636_8799.t111 464.166
R280 a_n7636_8799.n84 a_n7636_8799.t126 464.166
R281 a_n7636_8799.n86 a_n7636_8799.t79 464.166
R282 a_n7636_8799.n90 a_n7636_8799.t80 464.166
R283 a_n7636_8799.n91 a_n7636_8799.t109 464.166
R284 a_n7636_8799.n69 a_n7636_8799.t69 464.166
R285 a_n7636_8799.n96 a_n7636_8799.t70 464.166
R286 a_n7636_8799.n98 a_n7636_8799.t105 464.166
R287 a_n7636_8799.n102 a_n7636_8799.t44 464.166
R288 a_n7636_8799.n103 a_n7636_8799.t66 464.166
R289 a_n7636_8799.n65 a_n7636_8799.t87 464.166
R290 a_n7636_8799.n109 a_n7636_8799.t129 464.166
R291 a_n7636_8799.n110 a_n7636_8799.t55 464.166
R292 a_n7636_8799.n124 a_n7636_8799.t76 464.166
R293 a_n7636_8799.n128 a_n7636_8799.t110 464.166
R294 a_n7636_8799.n122 a_n7636_8799.t67 464.166
R295 a_n7636_8799.n133 a_n7636_8799.t118 464.166
R296 a_n7636_8799.n135 a_n7636_8799.t49 464.166
R297 a_n7636_8799.n139 a_n7636_8799.t37 464.166
R298 a_n7636_8799.n140 a_n7636_8799.t82 464.166
R299 a_n7636_8799.n118 a_n7636_8799.t121 464.166
R300 a_n7636_8799.n145 a_n7636_8799.t97 464.166
R301 a_n7636_8799.n147 a_n7636_8799.t125 464.166
R302 a_n7636_8799.n151 a_n7636_8799.t77 464.166
R303 a_n7636_8799.n152 a_n7636_8799.t41 464.166
R304 a_n7636_8799.n114 a_n7636_8799.t89 464.166
R305 a_n7636_8799.n158 a_n7636_8799.t53 464.166
R306 a_n7636_8799.n159 a_n7636_8799.t106 464.166
R307 a_n7636_8799.n178 a_n7636_8799.n177 161.3
R308 a_n7636_8799.n179 a_n7636_8799.n174 161.3
R309 a_n7636_8799.n180 a_n7636_8799.n173 161.3
R310 a_n7636_8799.n182 a_n7636_8799.n181 161.3
R311 a_n7636_8799.n183 a_n7636_8799.n172 161.3
R312 a_n7636_8799.n185 a_n7636_8799.n184 161.3
R313 a_n7636_8799.n186 a_n7636_8799.n171 161.3
R314 a_n7636_8799.n187 a_n7636_8799.n170 161.3
R315 a_n7636_8799.n189 a_n7636_8799.n188 161.3
R316 a_n7636_8799.n190 a_n7636_8799.n169 161.3
R317 a_n7636_8799.n192 a_n7636_8799.n191 161.3
R318 a_n7636_8799.n193 a_n7636_8799.n168 161.3
R319 a_n7636_8799.n194 a_n7636_8799.n167 161.3
R320 a_n7636_8799.n196 a_n7636_8799.n195 161.3
R321 a_n7636_8799.n197 a_n7636_8799.n166 161.3
R322 a_n7636_8799.n199 a_n7636_8799.n198 161.3
R323 a_n7636_8799.n200 a_n7636_8799.n165 161.3
R324 a_n7636_8799.n201 a_n7636_8799.n164 161.3
R325 a_n7636_8799.n203 a_n7636_8799.n202 161.3
R326 a_n7636_8799.n204 a_n7636_8799.n163 161.3
R327 a_n7636_8799.n206 a_n7636_8799.n205 161.3
R328 a_n7636_8799.n207 a_n7636_8799.n162 161.3
R329 a_n7636_8799.n209 a_n7636_8799.n208 161.3
R330 a_n7636_8799.n226 a_n7636_8799.n225 161.3
R331 a_n7636_8799.n227 a_n7636_8799.n222 161.3
R332 a_n7636_8799.n228 a_n7636_8799.n221 161.3
R333 a_n7636_8799.n230 a_n7636_8799.n229 161.3
R334 a_n7636_8799.n231 a_n7636_8799.n220 161.3
R335 a_n7636_8799.n233 a_n7636_8799.n232 161.3
R336 a_n7636_8799.n234 a_n7636_8799.n219 161.3
R337 a_n7636_8799.n235 a_n7636_8799.n218 161.3
R338 a_n7636_8799.n237 a_n7636_8799.n236 161.3
R339 a_n7636_8799.n238 a_n7636_8799.n217 161.3
R340 a_n7636_8799.n240 a_n7636_8799.n239 161.3
R341 a_n7636_8799.n241 a_n7636_8799.n216 161.3
R342 a_n7636_8799.n242 a_n7636_8799.n215 161.3
R343 a_n7636_8799.n244 a_n7636_8799.n243 161.3
R344 a_n7636_8799.n245 a_n7636_8799.n214 161.3
R345 a_n7636_8799.n247 a_n7636_8799.n246 161.3
R346 a_n7636_8799.n248 a_n7636_8799.n213 161.3
R347 a_n7636_8799.n249 a_n7636_8799.n212 161.3
R348 a_n7636_8799.n251 a_n7636_8799.n250 161.3
R349 a_n7636_8799.n252 a_n7636_8799.n211 161.3
R350 a_n7636_8799.n254 a_n7636_8799.n253 161.3
R351 a_n7636_8799.n255 a_n7636_8799.n210 161.3
R352 a_n7636_8799.n257 a_n7636_8799.n256 161.3
R353 a_n7636_8799.n275 a_n7636_8799.n274 161.3
R354 a_n7636_8799.n276 a_n7636_8799.n271 161.3
R355 a_n7636_8799.n277 a_n7636_8799.n270 161.3
R356 a_n7636_8799.n279 a_n7636_8799.n278 161.3
R357 a_n7636_8799.n280 a_n7636_8799.n269 161.3
R358 a_n7636_8799.n282 a_n7636_8799.n281 161.3
R359 a_n7636_8799.n283 a_n7636_8799.n268 161.3
R360 a_n7636_8799.n284 a_n7636_8799.n267 161.3
R361 a_n7636_8799.n286 a_n7636_8799.n285 161.3
R362 a_n7636_8799.n287 a_n7636_8799.n266 161.3
R363 a_n7636_8799.n289 a_n7636_8799.n288 161.3
R364 a_n7636_8799.n290 a_n7636_8799.n265 161.3
R365 a_n7636_8799.n291 a_n7636_8799.n264 161.3
R366 a_n7636_8799.n293 a_n7636_8799.n292 161.3
R367 a_n7636_8799.n294 a_n7636_8799.n263 161.3
R368 a_n7636_8799.n296 a_n7636_8799.n295 161.3
R369 a_n7636_8799.n297 a_n7636_8799.n262 161.3
R370 a_n7636_8799.n298 a_n7636_8799.n261 161.3
R371 a_n7636_8799.n300 a_n7636_8799.n299 161.3
R372 a_n7636_8799.n301 a_n7636_8799.n260 161.3
R373 a_n7636_8799.n303 a_n7636_8799.n302 161.3
R374 a_n7636_8799.n304 a_n7636_8799.n259 161.3
R375 a_n7636_8799.n306 a_n7636_8799.n305 161.3
R376 a_n7636_8799.n63 a_n7636_8799.n62 161.3
R377 a_n7636_8799.n61 a_n7636_8799.n16 161.3
R378 a_n7636_8799.n60 a_n7636_8799.n59 161.3
R379 a_n7636_8799.n58 a_n7636_8799.n17 161.3
R380 a_n7636_8799.n57 a_n7636_8799.n56 161.3
R381 a_n7636_8799.n55 a_n7636_8799.n18 161.3
R382 a_n7636_8799.n54 a_n7636_8799.n53 161.3
R383 a_n7636_8799.n52 a_n7636_8799.n19 161.3
R384 a_n7636_8799.n51 a_n7636_8799.n50 161.3
R385 a_n7636_8799.n49 a_n7636_8799.n20 161.3
R386 a_n7636_8799.n48 a_n7636_8799.n47 161.3
R387 a_n7636_8799.n46 a_n7636_8799.n21 161.3
R388 a_n7636_8799.n45 a_n7636_8799.n44 161.3
R389 a_n7636_8799.n43 a_n7636_8799.n22 161.3
R390 a_n7636_8799.n42 a_n7636_8799.n41 161.3
R391 a_n7636_8799.n40 a_n7636_8799.n23 161.3
R392 a_n7636_8799.n39 a_n7636_8799.n38 161.3
R393 a_n7636_8799.n37 a_n7636_8799.n24 161.3
R394 a_n7636_8799.n36 a_n7636_8799.n35 161.3
R395 a_n7636_8799.n34 a_n7636_8799.n25 161.3
R396 a_n7636_8799.n33 a_n7636_8799.n32 161.3
R397 a_n7636_8799.n31 a_n7636_8799.n26 161.3
R398 a_n7636_8799.n30 a_n7636_8799.n29 161.3
R399 a_n7636_8799.n111 a_n7636_8799.n110 161.3
R400 a_n7636_8799.n109 a_n7636_8799.n64 161.3
R401 a_n7636_8799.n108 a_n7636_8799.n107 161.3
R402 a_n7636_8799.n106 a_n7636_8799.n65 161.3
R403 a_n7636_8799.n105 a_n7636_8799.n104 161.3
R404 a_n7636_8799.n103 a_n7636_8799.n66 161.3
R405 a_n7636_8799.n102 a_n7636_8799.n101 161.3
R406 a_n7636_8799.n100 a_n7636_8799.n67 161.3
R407 a_n7636_8799.n99 a_n7636_8799.n98 161.3
R408 a_n7636_8799.n97 a_n7636_8799.n68 161.3
R409 a_n7636_8799.n96 a_n7636_8799.n95 161.3
R410 a_n7636_8799.n94 a_n7636_8799.n69 161.3
R411 a_n7636_8799.n93 a_n7636_8799.n92 161.3
R412 a_n7636_8799.n91 a_n7636_8799.n70 161.3
R413 a_n7636_8799.n90 a_n7636_8799.n89 161.3
R414 a_n7636_8799.n88 a_n7636_8799.n71 161.3
R415 a_n7636_8799.n87 a_n7636_8799.n86 161.3
R416 a_n7636_8799.n85 a_n7636_8799.n72 161.3
R417 a_n7636_8799.n84 a_n7636_8799.n83 161.3
R418 a_n7636_8799.n82 a_n7636_8799.n73 161.3
R419 a_n7636_8799.n81 a_n7636_8799.n80 161.3
R420 a_n7636_8799.n79 a_n7636_8799.n74 161.3
R421 a_n7636_8799.n78 a_n7636_8799.n77 161.3
R422 a_n7636_8799.n160 a_n7636_8799.n159 161.3
R423 a_n7636_8799.n158 a_n7636_8799.n113 161.3
R424 a_n7636_8799.n157 a_n7636_8799.n156 161.3
R425 a_n7636_8799.n155 a_n7636_8799.n114 161.3
R426 a_n7636_8799.n154 a_n7636_8799.n153 161.3
R427 a_n7636_8799.n152 a_n7636_8799.n115 161.3
R428 a_n7636_8799.n151 a_n7636_8799.n150 161.3
R429 a_n7636_8799.n149 a_n7636_8799.n116 161.3
R430 a_n7636_8799.n148 a_n7636_8799.n147 161.3
R431 a_n7636_8799.n146 a_n7636_8799.n117 161.3
R432 a_n7636_8799.n145 a_n7636_8799.n144 161.3
R433 a_n7636_8799.n143 a_n7636_8799.n118 161.3
R434 a_n7636_8799.n142 a_n7636_8799.n141 161.3
R435 a_n7636_8799.n140 a_n7636_8799.n119 161.3
R436 a_n7636_8799.n139 a_n7636_8799.n138 161.3
R437 a_n7636_8799.n137 a_n7636_8799.n120 161.3
R438 a_n7636_8799.n136 a_n7636_8799.n135 161.3
R439 a_n7636_8799.n134 a_n7636_8799.n121 161.3
R440 a_n7636_8799.n133 a_n7636_8799.n132 161.3
R441 a_n7636_8799.n131 a_n7636_8799.n122 161.3
R442 a_n7636_8799.n130 a_n7636_8799.n129 161.3
R443 a_n7636_8799.n128 a_n7636_8799.n123 161.3
R444 a_n7636_8799.n127 a_n7636_8799.n126 161.3
R445 a_n7636_8799.n10 a_n7636_8799.n8 98.9633
R446 a_n7636_8799.n3 a_n7636_8799.n1 98.9631
R447 a_n7636_8799.n14 a_n7636_8799.n13 98.6055
R448 a_n7636_8799.n12 a_n7636_8799.n11 98.6055
R449 a_n7636_8799.n10 a_n7636_8799.n9 98.6055
R450 a_n7636_8799.n3 a_n7636_8799.n2 98.6055
R451 a_n7636_8799.n5 a_n7636_8799.n4 98.6055
R452 a_n7636_8799.n7 a_n7636_8799.n6 98.6055
R453 a_n7636_8799.n312 a_n7636_8799.n310 81.3764
R454 a_n7636_8799.n321 a_n7636_8799.n319 81.3764
R455 a_n7636_8799.n324 a_n7636_8799.n0 81.3764
R456 a_n7636_8799.n325 a_n7636_8799.n324 80.9326
R457 a_n7636_8799.n318 a_n7636_8799.n317 80.9324
R458 a_n7636_8799.n316 a_n7636_8799.n315 80.9324
R459 a_n7636_8799.n314 a_n7636_8799.n313 80.9324
R460 a_n7636_8799.n312 a_n7636_8799.n311 80.9324
R461 a_n7636_8799.n321 a_n7636_8799.n320 80.9324
R462 a_n7636_8799.n323 a_n7636_8799.n322 80.9324
R463 a_n7636_8799.n177 a_n7636_8799.n176 70.4033
R464 a_n7636_8799.n225 a_n7636_8799.n224 70.4033
R465 a_n7636_8799.n274 a_n7636_8799.n273 70.4033
R466 a_n7636_8799.n29 a_n7636_8799.n28 70.4033
R467 a_n7636_8799.n77 a_n7636_8799.n76 70.4033
R468 a_n7636_8799.n126 a_n7636_8799.n125 70.4033
R469 a_n7636_8799.n208 a_n7636_8799.n207 48.2005
R470 a_n7636_8799.n201 a_n7636_8799.n200 48.2005
R471 a_n7636_8799.n194 a_n7636_8799.n193 48.2005
R472 a_n7636_8799.n188 a_n7636_8799.n169 48.2005
R473 a_n7636_8799.n181 a_n7636_8799.n172 48.2005
R474 a_n7636_8799.n256 a_n7636_8799.n255 48.2005
R475 a_n7636_8799.n249 a_n7636_8799.n248 48.2005
R476 a_n7636_8799.n242 a_n7636_8799.n241 48.2005
R477 a_n7636_8799.n236 a_n7636_8799.n217 48.2005
R478 a_n7636_8799.n229 a_n7636_8799.n220 48.2005
R479 a_n7636_8799.n305 a_n7636_8799.n304 48.2005
R480 a_n7636_8799.n298 a_n7636_8799.n297 48.2005
R481 a_n7636_8799.n291 a_n7636_8799.n290 48.2005
R482 a_n7636_8799.n285 a_n7636_8799.n266 48.2005
R483 a_n7636_8799.n278 a_n7636_8799.n269 48.2005
R484 a_n7636_8799.n36 a_n7636_8799.n25 48.2005
R485 a_n7636_8799.n43 a_n7636_8799.n42 48.2005
R486 a_n7636_8799.n48 a_n7636_8799.n21 48.2005
R487 a_n7636_8799.n55 a_n7636_8799.n54 48.2005
R488 a_n7636_8799.n62 a_n7636_8799.n61 48.2005
R489 a_n7636_8799.n84 a_n7636_8799.n73 48.2005
R490 a_n7636_8799.n91 a_n7636_8799.n90 48.2005
R491 a_n7636_8799.n96 a_n7636_8799.n69 48.2005
R492 a_n7636_8799.n103 a_n7636_8799.n102 48.2005
R493 a_n7636_8799.n110 a_n7636_8799.n109 48.2005
R494 a_n7636_8799.n133 a_n7636_8799.n122 48.2005
R495 a_n7636_8799.n140 a_n7636_8799.n139 48.2005
R496 a_n7636_8799.n145 a_n7636_8799.n118 48.2005
R497 a_n7636_8799.n152 a_n7636_8799.n151 48.2005
R498 a_n7636_8799.n159 a_n7636_8799.n158 48.2005
R499 a_n7636_8799.n195 a_n7636_8799.n166 47.4702
R500 a_n7636_8799.n187 a_n7636_8799.n186 47.4702
R501 a_n7636_8799.n243 a_n7636_8799.n214 47.4702
R502 a_n7636_8799.n235 a_n7636_8799.n234 47.4702
R503 a_n7636_8799.n292 a_n7636_8799.n263 47.4702
R504 a_n7636_8799.n284 a_n7636_8799.n283 47.4702
R505 a_n7636_8799.n38 a_n7636_8799.n23 47.4702
R506 a_n7636_8799.n50 a_n7636_8799.n49 47.4702
R507 a_n7636_8799.n86 a_n7636_8799.n71 47.4702
R508 a_n7636_8799.n98 a_n7636_8799.n97 47.4702
R509 a_n7636_8799.n135 a_n7636_8799.n120 47.4702
R510 a_n7636_8799.n147 a_n7636_8799.n146 47.4702
R511 a_n7636_8799.n202 a_n7636_8799.n163 46.0096
R512 a_n7636_8799.n180 a_n7636_8799.n179 46.0096
R513 a_n7636_8799.n250 a_n7636_8799.n211 46.0096
R514 a_n7636_8799.n228 a_n7636_8799.n227 46.0096
R515 a_n7636_8799.n299 a_n7636_8799.n260 46.0096
R516 a_n7636_8799.n277 a_n7636_8799.n276 46.0096
R517 a_n7636_8799.n32 a_n7636_8799.n31 46.0096
R518 a_n7636_8799.n56 a_n7636_8799.n17 46.0096
R519 a_n7636_8799.n80 a_n7636_8799.n79 46.0096
R520 a_n7636_8799.n104 a_n7636_8799.n65 46.0096
R521 a_n7636_8799.n129 a_n7636_8799.n128 46.0096
R522 a_n7636_8799.n153 a_n7636_8799.n114 46.0096
R523 a_n7636_8799.n323 a_n7636_8799.n318 32.7526
R524 a_n7636_8799.n15 a_n7636_8799.n7 31.7868
R525 a_n7636_8799.n206 a_n7636_8799.n163 27.0217
R526 a_n7636_8799.n179 a_n7636_8799.n178 27.0217
R527 a_n7636_8799.n254 a_n7636_8799.n211 27.0217
R528 a_n7636_8799.n227 a_n7636_8799.n226 27.0217
R529 a_n7636_8799.n303 a_n7636_8799.n260 27.0217
R530 a_n7636_8799.n276 a_n7636_8799.n275 27.0217
R531 a_n7636_8799.n31 a_n7636_8799.n30 27.0217
R532 a_n7636_8799.n60 a_n7636_8799.n17 27.0217
R533 a_n7636_8799.n79 a_n7636_8799.n78 27.0217
R534 a_n7636_8799.n108 a_n7636_8799.n65 27.0217
R535 a_n7636_8799.n128 a_n7636_8799.n127 27.0217
R536 a_n7636_8799.n157 a_n7636_8799.n114 27.0217
R537 a_n7636_8799.n199 a_n7636_8799.n166 25.5611
R538 a_n7636_8799.n186 a_n7636_8799.n185 25.5611
R539 a_n7636_8799.n247 a_n7636_8799.n214 25.5611
R540 a_n7636_8799.n234 a_n7636_8799.n233 25.5611
R541 a_n7636_8799.n296 a_n7636_8799.n263 25.5611
R542 a_n7636_8799.n283 a_n7636_8799.n282 25.5611
R543 a_n7636_8799.n38 a_n7636_8799.n37 25.5611
R544 a_n7636_8799.n50 a_n7636_8799.n19 25.5611
R545 a_n7636_8799.n86 a_n7636_8799.n85 25.5611
R546 a_n7636_8799.n98 a_n7636_8799.n67 25.5611
R547 a_n7636_8799.n135 a_n7636_8799.n134 25.5611
R548 a_n7636_8799.n147 a_n7636_8799.n116 25.5611
R549 a_n7636_8799.n193 a_n7636_8799.n192 24.1005
R550 a_n7636_8799.n192 a_n7636_8799.n169 24.1005
R551 a_n7636_8799.n241 a_n7636_8799.n240 24.1005
R552 a_n7636_8799.n240 a_n7636_8799.n217 24.1005
R553 a_n7636_8799.n290 a_n7636_8799.n289 24.1005
R554 a_n7636_8799.n289 a_n7636_8799.n266 24.1005
R555 a_n7636_8799.n44 a_n7636_8799.n43 24.1005
R556 a_n7636_8799.n44 a_n7636_8799.n21 24.1005
R557 a_n7636_8799.n92 a_n7636_8799.n91 24.1005
R558 a_n7636_8799.n92 a_n7636_8799.n69 24.1005
R559 a_n7636_8799.n141 a_n7636_8799.n140 24.1005
R560 a_n7636_8799.n141 a_n7636_8799.n118 24.1005
R561 a_n7636_8799.n200 a_n7636_8799.n199 22.6399
R562 a_n7636_8799.n185 a_n7636_8799.n172 22.6399
R563 a_n7636_8799.n248 a_n7636_8799.n247 22.6399
R564 a_n7636_8799.n233 a_n7636_8799.n220 22.6399
R565 a_n7636_8799.n297 a_n7636_8799.n296 22.6399
R566 a_n7636_8799.n282 a_n7636_8799.n269 22.6399
R567 a_n7636_8799.n37 a_n7636_8799.n36 22.6399
R568 a_n7636_8799.n54 a_n7636_8799.n19 22.6399
R569 a_n7636_8799.n85 a_n7636_8799.n84 22.6399
R570 a_n7636_8799.n102 a_n7636_8799.n67 22.6399
R571 a_n7636_8799.n134 a_n7636_8799.n133 22.6399
R572 a_n7636_8799.n151 a_n7636_8799.n116 22.6399
R573 a_n7636_8799.n207 a_n7636_8799.n206 21.1793
R574 a_n7636_8799.n178 a_n7636_8799.n175 21.1793
R575 a_n7636_8799.n255 a_n7636_8799.n254 21.1793
R576 a_n7636_8799.n226 a_n7636_8799.n223 21.1793
R577 a_n7636_8799.n304 a_n7636_8799.n303 21.1793
R578 a_n7636_8799.n275 a_n7636_8799.n272 21.1793
R579 a_n7636_8799.n30 a_n7636_8799.n27 21.1793
R580 a_n7636_8799.n61 a_n7636_8799.n60 21.1793
R581 a_n7636_8799.n78 a_n7636_8799.n75 21.1793
R582 a_n7636_8799.n109 a_n7636_8799.n108 21.1793
R583 a_n7636_8799.n127 a_n7636_8799.n124 21.1793
R584 a_n7636_8799.n158 a_n7636_8799.n157 21.1793
R585 a_n7636_8799.n176 a_n7636_8799.n175 20.9576
R586 a_n7636_8799.n224 a_n7636_8799.n223 20.9576
R587 a_n7636_8799.n273 a_n7636_8799.n272 20.9576
R588 a_n7636_8799.n28 a_n7636_8799.n27 20.9576
R589 a_n7636_8799.n76 a_n7636_8799.n75 20.9576
R590 a_n7636_8799.n125 a_n7636_8799.n124 20.9576
R591 a_n7636_8799.n15 a_n7636_8799.n14 18.8093
R592 a_n7636_8799.n314 a_n7636_8799.n309 12.3339
R593 a_n7636_8799.n309 a_n7636_8799.n15 11.4887
R594 a_n7636_8799.n258 a_n7636_8799.n209 9.07815
R595 a_n7636_8799.n112 a_n7636_8799.n63 9.07815
R596 a_n7636_8799.n308 a_n7636_8799.n161 6.97387
R597 a_n7636_8799.n308 a_n7636_8799.n307 6.61699
R598 a_n7636_8799.n258 a_n7636_8799.n257 4.9702
R599 a_n7636_8799.n307 a_n7636_8799.n306 4.9702
R600 a_n7636_8799.n112 a_n7636_8799.n111 4.9702
R601 a_n7636_8799.n161 a_n7636_8799.n160 4.9702
R602 a_n7636_8799.n307 a_n7636_8799.n258 4.10845
R603 a_n7636_8799.n161 a_n7636_8799.n112 4.10845
R604 a_n7636_8799.n13 a_n7636_8799.t2 3.61217
R605 a_n7636_8799.n13 a_n7636_8799.t6 3.61217
R606 a_n7636_8799.n11 a_n7636_8799.t34 3.61217
R607 a_n7636_8799.n11 a_n7636_8799.t1 3.61217
R608 a_n7636_8799.n9 a_n7636_8799.t10 3.61217
R609 a_n7636_8799.n9 a_n7636_8799.t32 3.61217
R610 a_n7636_8799.n8 a_n7636_8799.t5 3.61217
R611 a_n7636_8799.n8 a_n7636_8799.t9 3.61217
R612 a_n7636_8799.n1 a_n7636_8799.t33 3.61217
R613 a_n7636_8799.n1 a_n7636_8799.t7 3.61217
R614 a_n7636_8799.n2 a_n7636_8799.t4 3.61217
R615 a_n7636_8799.n2 a_n7636_8799.t8 3.61217
R616 a_n7636_8799.n4 a_n7636_8799.t35 3.61217
R617 a_n7636_8799.n4 a_n7636_8799.t3 3.61217
R618 a_n7636_8799.n6 a_n7636_8799.t0 3.61217
R619 a_n7636_8799.n6 a_n7636_8799.t31 3.61217
R620 a_n7636_8799.n309 a_n7636_8799.n308 3.4105
R621 a_n7636_8799.n319 a_n7636_8799.t24 2.82907
R622 a_n7636_8799.n319 a_n7636_8799.t22 2.82907
R623 a_n7636_8799.n320 a_n7636_8799.t15 2.82907
R624 a_n7636_8799.n320 a_n7636_8799.t19 2.82907
R625 a_n7636_8799.n322 a_n7636_8799.t29 2.82907
R626 a_n7636_8799.n322 a_n7636_8799.t16 2.82907
R627 a_n7636_8799.n317 a_n7636_8799.t25 2.82907
R628 a_n7636_8799.n317 a_n7636_8799.t11 2.82907
R629 a_n7636_8799.n315 a_n7636_8799.t28 2.82907
R630 a_n7636_8799.n315 a_n7636_8799.t23 2.82907
R631 a_n7636_8799.n313 a_n7636_8799.t12 2.82907
R632 a_n7636_8799.n313 a_n7636_8799.t27 2.82907
R633 a_n7636_8799.n311 a_n7636_8799.t13 2.82907
R634 a_n7636_8799.n311 a_n7636_8799.t14 2.82907
R635 a_n7636_8799.n310 a_n7636_8799.t17 2.82907
R636 a_n7636_8799.n310 a_n7636_8799.t18 2.82907
R637 a_n7636_8799.n0 a_n7636_8799.t21 2.82907
R638 a_n7636_8799.n0 a_n7636_8799.t20 2.82907
R639 a_n7636_8799.n325 a_n7636_8799.t26 2.82907
R640 a_n7636_8799.t30 a_n7636_8799.n325 2.82907
R641 a_n7636_8799.n202 a_n7636_8799.n201 2.19141
R642 a_n7636_8799.n181 a_n7636_8799.n180 2.19141
R643 a_n7636_8799.n250 a_n7636_8799.n249 2.19141
R644 a_n7636_8799.n229 a_n7636_8799.n228 2.19141
R645 a_n7636_8799.n299 a_n7636_8799.n298 2.19141
R646 a_n7636_8799.n278 a_n7636_8799.n277 2.19141
R647 a_n7636_8799.n32 a_n7636_8799.n25 2.19141
R648 a_n7636_8799.n56 a_n7636_8799.n55 2.19141
R649 a_n7636_8799.n80 a_n7636_8799.n73 2.19141
R650 a_n7636_8799.n104 a_n7636_8799.n103 2.19141
R651 a_n7636_8799.n129 a_n7636_8799.n122 2.19141
R652 a_n7636_8799.n153 a_n7636_8799.n152 2.19141
R653 a_n7636_8799.n195 a_n7636_8799.n194 0.730803
R654 a_n7636_8799.n188 a_n7636_8799.n187 0.730803
R655 a_n7636_8799.n243 a_n7636_8799.n242 0.730803
R656 a_n7636_8799.n236 a_n7636_8799.n235 0.730803
R657 a_n7636_8799.n292 a_n7636_8799.n291 0.730803
R658 a_n7636_8799.n285 a_n7636_8799.n284 0.730803
R659 a_n7636_8799.n42 a_n7636_8799.n23 0.730803
R660 a_n7636_8799.n49 a_n7636_8799.n48 0.730803
R661 a_n7636_8799.n90 a_n7636_8799.n71 0.730803
R662 a_n7636_8799.n97 a_n7636_8799.n96 0.730803
R663 a_n7636_8799.n139 a_n7636_8799.n120 0.730803
R664 a_n7636_8799.n146 a_n7636_8799.n145 0.730803
R665 a_n7636_8799.n314 a_n7636_8799.n312 0.444466
R666 a_n7636_8799.n316 a_n7636_8799.n314 0.444466
R667 a_n7636_8799.n318 a_n7636_8799.n316 0.444466
R668 a_n7636_8799.n324 a_n7636_8799.n323 0.444466
R669 a_n7636_8799.n323 a_n7636_8799.n321 0.444466
R670 a_n7636_8799.n12 a_n7636_8799.n10 0.358259
R671 a_n7636_8799.n14 a_n7636_8799.n12 0.358259
R672 a_n7636_8799.n7 a_n7636_8799.n5 0.358259
R673 a_n7636_8799.n5 a_n7636_8799.n3 0.358259
R674 a_n7636_8799.n209 a_n7636_8799.n162 0.189894
R675 a_n7636_8799.n205 a_n7636_8799.n162 0.189894
R676 a_n7636_8799.n205 a_n7636_8799.n204 0.189894
R677 a_n7636_8799.n204 a_n7636_8799.n203 0.189894
R678 a_n7636_8799.n203 a_n7636_8799.n164 0.189894
R679 a_n7636_8799.n165 a_n7636_8799.n164 0.189894
R680 a_n7636_8799.n198 a_n7636_8799.n165 0.189894
R681 a_n7636_8799.n198 a_n7636_8799.n197 0.189894
R682 a_n7636_8799.n197 a_n7636_8799.n196 0.189894
R683 a_n7636_8799.n196 a_n7636_8799.n167 0.189894
R684 a_n7636_8799.n168 a_n7636_8799.n167 0.189894
R685 a_n7636_8799.n191 a_n7636_8799.n168 0.189894
R686 a_n7636_8799.n191 a_n7636_8799.n190 0.189894
R687 a_n7636_8799.n190 a_n7636_8799.n189 0.189894
R688 a_n7636_8799.n189 a_n7636_8799.n170 0.189894
R689 a_n7636_8799.n171 a_n7636_8799.n170 0.189894
R690 a_n7636_8799.n184 a_n7636_8799.n171 0.189894
R691 a_n7636_8799.n184 a_n7636_8799.n183 0.189894
R692 a_n7636_8799.n183 a_n7636_8799.n182 0.189894
R693 a_n7636_8799.n182 a_n7636_8799.n173 0.189894
R694 a_n7636_8799.n174 a_n7636_8799.n173 0.189894
R695 a_n7636_8799.n177 a_n7636_8799.n174 0.189894
R696 a_n7636_8799.n257 a_n7636_8799.n210 0.189894
R697 a_n7636_8799.n253 a_n7636_8799.n210 0.189894
R698 a_n7636_8799.n253 a_n7636_8799.n252 0.189894
R699 a_n7636_8799.n252 a_n7636_8799.n251 0.189894
R700 a_n7636_8799.n251 a_n7636_8799.n212 0.189894
R701 a_n7636_8799.n213 a_n7636_8799.n212 0.189894
R702 a_n7636_8799.n246 a_n7636_8799.n213 0.189894
R703 a_n7636_8799.n246 a_n7636_8799.n245 0.189894
R704 a_n7636_8799.n245 a_n7636_8799.n244 0.189894
R705 a_n7636_8799.n244 a_n7636_8799.n215 0.189894
R706 a_n7636_8799.n216 a_n7636_8799.n215 0.189894
R707 a_n7636_8799.n239 a_n7636_8799.n216 0.189894
R708 a_n7636_8799.n239 a_n7636_8799.n238 0.189894
R709 a_n7636_8799.n238 a_n7636_8799.n237 0.189894
R710 a_n7636_8799.n237 a_n7636_8799.n218 0.189894
R711 a_n7636_8799.n219 a_n7636_8799.n218 0.189894
R712 a_n7636_8799.n232 a_n7636_8799.n219 0.189894
R713 a_n7636_8799.n232 a_n7636_8799.n231 0.189894
R714 a_n7636_8799.n231 a_n7636_8799.n230 0.189894
R715 a_n7636_8799.n230 a_n7636_8799.n221 0.189894
R716 a_n7636_8799.n222 a_n7636_8799.n221 0.189894
R717 a_n7636_8799.n225 a_n7636_8799.n222 0.189894
R718 a_n7636_8799.n306 a_n7636_8799.n259 0.189894
R719 a_n7636_8799.n302 a_n7636_8799.n259 0.189894
R720 a_n7636_8799.n302 a_n7636_8799.n301 0.189894
R721 a_n7636_8799.n301 a_n7636_8799.n300 0.189894
R722 a_n7636_8799.n300 a_n7636_8799.n261 0.189894
R723 a_n7636_8799.n262 a_n7636_8799.n261 0.189894
R724 a_n7636_8799.n295 a_n7636_8799.n262 0.189894
R725 a_n7636_8799.n295 a_n7636_8799.n294 0.189894
R726 a_n7636_8799.n294 a_n7636_8799.n293 0.189894
R727 a_n7636_8799.n293 a_n7636_8799.n264 0.189894
R728 a_n7636_8799.n265 a_n7636_8799.n264 0.189894
R729 a_n7636_8799.n288 a_n7636_8799.n265 0.189894
R730 a_n7636_8799.n288 a_n7636_8799.n287 0.189894
R731 a_n7636_8799.n287 a_n7636_8799.n286 0.189894
R732 a_n7636_8799.n286 a_n7636_8799.n267 0.189894
R733 a_n7636_8799.n268 a_n7636_8799.n267 0.189894
R734 a_n7636_8799.n281 a_n7636_8799.n268 0.189894
R735 a_n7636_8799.n281 a_n7636_8799.n280 0.189894
R736 a_n7636_8799.n280 a_n7636_8799.n279 0.189894
R737 a_n7636_8799.n279 a_n7636_8799.n270 0.189894
R738 a_n7636_8799.n271 a_n7636_8799.n270 0.189894
R739 a_n7636_8799.n274 a_n7636_8799.n271 0.189894
R740 a_n7636_8799.n29 a_n7636_8799.n26 0.189894
R741 a_n7636_8799.n33 a_n7636_8799.n26 0.189894
R742 a_n7636_8799.n34 a_n7636_8799.n33 0.189894
R743 a_n7636_8799.n35 a_n7636_8799.n34 0.189894
R744 a_n7636_8799.n35 a_n7636_8799.n24 0.189894
R745 a_n7636_8799.n39 a_n7636_8799.n24 0.189894
R746 a_n7636_8799.n40 a_n7636_8799.n39 0.189894
R747 a_n7636_8799.n41 a_n7636_8799.n40 0.189894
R748 a_n7636_8799.n41 a_n7636_8799.n22 0.189894
R749 a_n7636_8799.n45 a_n7636_8799.n22 0.189894
R750 a_n7636_8799.n46 a_n7636_8799.n45 0.189894
R751 a_n7636_8799.n47 a_n7636_8799.n46 0.189894
R752 a_n7636_8799.n47 a_n7636_8799.n20 0.189894
R753 a_n7636_8799.n51 a_n7636_8799.n20 0.189894
R754 a_n7636_8799.n52 a_n7636_8799.n51 0.189894
R755 a_n7636_8799.n53 a_n7636_8799.n52 0.189894
R756 a_n7636_8799.n53 a_n7636_8799.n18 0.189894
R757 a_n7636_8799.n57 a_n7636_8799.n18 0.189894
R758 a_n7636_8799.n58 a_n7636_8799.n57 0.189894
R759 a_n7636_8799.n59 a_n7636_8799.n58 0.189894
R760 a_n7636_8799.n59 a_n7636_8799.n16 0.189894
R761 a_n7636_8799.n63 a_n7636_8799.n16 0.189894
R762 a_n7636_8799.n77 a_n7636_8799.n74 0.189894
R763 a_n7636_8799.n81 a_n7636_8799.n74 0.189894
R764 a_n7636_8799.n82 a_n7636_8799.n81 0.189894
R765 a_n7636_8799.n83 a_n7636_8799.n82 0.189894
R766 a_n7636_8799.n83 a_n7636_8799.n72 0.189894
R767 a_n7636_8799.n87 a_n7636_8799.n72 0.189894
R768 a_n7636_8799.n88 a_n7636_8799.n87 0.189894
R769 a_n7636_8799.n89 a_n7636_8799.n88 0.189894
R770 a_n7636_8799.n89 a_n7636_8799.n70 0.189894
R771 a_n7636_8799.n93 a_n7636_8799.n70 0.189894
R772 a_n7636_8799.n94 a_n7636_8799.n93 0.189894
R773 a_n7636_8799.n95 a_n7636_8799.n94 0.189894
R774 a_n7636_8799.n95 a_n7636_8799.n68 0.189894
R775 a_n7636_8799.n99 a_n7636_8799.n68 0.189894
R776 a_n7636_8799.n100 a_n7636_8799.n99 0.189894
R777 a_n7636_8799.n101 a_n7636_8799.n100 0.189894
R778 a_n7636_8799.n101 a_n7636_8799.n66 0.189894
R779 a_n7636_8799.n105 a_n7636_8799.n66 0.189894
R780 a_n7636_8799.n106 a_n7636_8799.n105 0.189894
R781 a_n7636_8799.n107 a_n7636_8799.n106 0.189894
R782 a_n7636_8799.n107 a_n7636_8799.n64 0.189894
R783 a_n7636_8799.n111 a_n7636_8799.n64 0.189894
R784 a_n7636_8799.n126 a_n7636_8799.n123 0.189894
R785 a_n7636_8799.n130 a_n7636_8799.n123 0.189894
R786 a_n7636_8799.n131 a_n7636_8799.n130 0.189894
R787 a_n7636_8799.n132 a_n7636_8799.n131 0.189894
R788 a_n7636_8799.n132 a_n7636_8799.n121 0.189894
R789 a_n7636_8799.n136 a_n7636_8799.n121 0.189894
R790 a_n7636_8799.n137 a_n7636_8799.n136 0.189894
R791 a_n7636_8799.n138 a_n7636_8799.n137 0.189894
R792 a_n7636_8799.n138 a_n7636_8799.n119 0.189894
R793 a_n7636_8799.n142 a_n7636_8799.n119 0.189894
R794 a_n7636_8799.n143 a_n7636_8799.n142 0.189894
R795 a_n7636_8799.n144 a_n7636_8799.n143 0.189894
R796 a_n7636_8799.n144 a_n7636_8799.n117 0.189894
R797 a_n7636_8799.n148 a_n7636_8799.n117 0.189894
R798 a_n7636_8799.n149 a_n7636_8799.n148 0.189894
R799 a_n7636_8799.n150 a_n7636_8799.n149 0.189894
R800 a_n7636_8799.n150 a_n7636_8799.n115 0.189894
R801 a_n7636_8799.n154 a_n7636_8799.n115 0.189894
R802 a_n7636_8799.n155 a_n7636_8799.n154 0.189894
R803 a_n7636_8799.n156 a_n7636_8799.n155 0.189894
R804 a_n7636_8799.n156 a_n7636_8799.n113 0.189894
R805 a_n7636_8799.n160 a_n7636_8799.n113 0.189894
R806 gnd.n7003 gnd.n546 965.481
R807 gnd.n3813 gnd.n3812 939.716
R808 gnd.n3720 gnd.n2339 766.379
R809 gnd.n3723 gnd.n3722 766.379
R810 gnd.n2962 gnd.n2865 766.379
R811 gnd.n2958 gnd.n2863 766.379
R812 gnd.n3811 gnd.n2361 756.769
R813 gnd.n3714 gnd.n3713 756.769
R814 gnd.n3055 gnd.n2772 756.769
R815 gnd.n3053 gnd.n2775 756.769
R816 gnd.n6581 gnd.n798 756.769
R817 gnd.n7002 gnd.n547 756.769
R818 gnd.n7214 gnd.n7213 756.769
R819 gnd.n6404 gnd.n963 756.769
R820 gnd.n7509 gnd.n129 751.963
R821 gnd.n7667 gnd.n7666 751.963
R822 gnd.n1337 gnd.n1284 751.963
R823 gnd.n6078 gnd.n1339 751.963
R824 gnd.n6323 gnd.n1113 751.963
R825 gnd.n4849 gnd.n1111 751.963
R826 gnd.n3880 gnd.n3815 751.963
R827 gnd.n4200 gnd.n2338 751.963
R828 gnd.n7664 gnd.n131 732.745
R829 gnd.n199 gnd.n127 732.745
R830 gnd.n6081 gnd.n6080 732.745
R831 gnd.n6153 gnd.n1288 732.745
R832 gnd.n6325 gnd.n1108 732.745
R833 gnd.n2123 gnd.n1110 732.745
R834 gnd.n4119 gnd.n3814 732.745
R835 gnd.n4198 gnd.n3978 732.745
R836 gnd.n4895 gnd.n1118 711.122
R837 gnd.n6165 gnd.n1244 711.122
R838 gnd.n4905 gnd.n1975 711.122
R839 gnd.n5883 gnd.n1247 711.122
R840 gnd.n6577 gnd.n798 585
R841 gnd.n798 gnd.n797 585
R842 gnd.n6576 gnd.n6575 585
R843 gnd.n6575 gnd.n6574 585
R844 gnd.n801 gnd.n800 585
R845 gnd.n6573 gnd.n801 585
R846 gnd.n6571 gnd.n6570 585
R847 gnd.n6572 gnd.n6571 585
R848 gnd.n6569 gnd.n803 585
R849 gnd.n803 gnd.n802 585
R850 gnd.n6568 gnd.n6567 585
R851 gnd.n6567 gnd.n6566 585
R852 gnd.n809 gnd.n808 585
R853 gnd.n6565 gnd.n809 585
R854 gnd.n6563 gnd.n6562 585
R855 gnd.n6564 gnd.n6563 585
R856 gnd.n6561 gnd.n811 585
R857 gnd.n811 gnd.n810 585
R858 gnd.n6560 gnd.n6559 585
R859 gnd.n6559 gnd.n6558 585
R860 gnd.n817 gnd.n816 585
R861 gnd.n6557 gnd.n817 585
R862 gnd.n6555 gnd.n6554 585
R863 gnd.n6556 gnd.n6555 585
R864 gnd.n6553 gnd.n819 585
R865 gnd.n819 gnd.n818 585
R866 gnd.n6552 gnd.n6551 585
R867 gnd.n6551 gnd.n6550 585
R868 gnd.n825 gnd.n824 585
R869 gnd.n6549 gnd.n825 585
R870 gnd.n6547 gnd.n6546 585
R871 gnd.n6548 gnd.n6547 585
R872 gnd.n6545 gnd.n827 585
R873 gnd.n827 gnd.n826 585
R874 gnd.n6544 gnd.n6543 585
R875 gnd.n6543 gnd.n6542 585
R876 gnd.n833 gnd.n832 585
R877 gnd.n6541 gnd.n833 585
R878 gnd.n6539 gnd.n6538 585
R879 gnd.n6540 gnd.n6539 585
R880 gnd.n6537 gnd.n835 585
R881 gnd.n835 gnd.n834 585
R882 gnd.n6536 gnd.n6535 585
R883 gnd.n6535 gnd.n6534 585
R884 gnd.n841 gnd.n840 585
R885 gnd.n6533 gnd.n841 585
R886 gnd.n6531 gnd.n6530 585
R887 gnd.n6532 gnd.n6531 585
R888 gnd.n6529 gnd.n843 585
R889 gnd.n843 gnd.n842 585
R890 gnd.n6528 gnd.n6527 585
R891 gnd.n6527 gnd.n6526 585
R892 gnd.n849 gnd.n848 585
R893 gnd.n6525 gnd.n849 585
R894 gnd.n6523 gnd.n6522 585
R895 gnd.n6524 gnd.n6523 585
R896 gnd.n6521 gnd.n851 585
R897 gnd.n851 gnd.n850 585
R898 gnd.n6520 gnd.n6519 585
R899 gnd.n6519 gnd.n6518 585
R900 gnd.n857 gnd.n856 585
R901 gnd.n6517 gnd.n857 585
R902 gnd.n6515 gnd.n6514 585
R903 gnd.n6516 gnd.n6515 585
R904 gnd.n6513 gnd.n859 585
R905 gnd.n859 gnd.n858 585
R906 gnd.n6512 gnd.n6511 585
R907 gnd.n6511 gnd.n6510 585
R908 gnd.n865 gnd.n864 585
R909 gnd.n6509 gnd.n865 585
R910 gnd.n6507 gnd.n6506 585
R911 gnd.n6508 gnd.n6507 585
R912 gnd.n6505 gnd.n867 585
R913 gnd.n867 gnd.n866 585
R914 gnd.n6504 gnd.n6503 585
R915 gnd.n6503 gnd.n6502 585
R916 gnd.n873 gnd.n872 585
R917 gnd.n6501 gnd.n873 585
R918 gnd.n6499 gnd.n6498 585
R919 gnd.n6500 gnd.n6499 585
R920 gnd.n6497 gnd.n875 585
R921 gnd.n875 gnd.n874 585
R922 gnd.n6496 gnd.n6495 585
R923 gnd.n6495 gnd.n6494 585
R924 gnd.n881 gnd.n880 585
R925 gnd.n6493 gnd.n881 585
R926 gnd.n6491 gnd.n6490 585
R927 gnd.n6492 gnd.n6491 585
R928 gnd.n6489 gnd.n883 585
R929 gnd.n883 gnd.n882 585
R930 gnd.n6488 gnd.n6487 585
R931 gnd.n6487 gnd.n6486 585
R932 gnd.n889 gnd.n888 585
R933 gnd.n6485 gnd.n889 585
R934 gnd.n6483 gnd.n6482 585
R935 gnd.n6484 gnd.n6483 585
R936 gnd.n6481 gnd.n891 585
R937 gnd.n891 gnd.n890 585
R938 gnd.n6480 gnd.n6479 585
R939 gnd.n6479 gnd.n6478 585
R940 gnd.n897 gnd.n896 585
R941 gnd.n6477 gnd.n897 585
R942 gnd.n6475 gnd.n6474 585
R943 gnd.n6476 gnd.n6475 585
R944 gnd.n6473 gnd.n899 585
R945 gnd.n899 gnd.n898 585
R946 gnd.n6472 gnd.n6471 585
R947 gnd.n6471 gnd.n6470 585
R948 gnd.n905 gnd.n904 585
R949 gnd.n6469 gnd.n905 585
R950 gnd.n6467 gnd.n6466 585
R951 gnd.n6468 gnd.n6467 585
R952 gnd.n6465 gnd.n907 585
R953 gnd.n907 gnd.n906 585
R954 gnd.n6464 gnd.n6463 585
R955 gnd.n6463 gnd.n6462 585
R956 gnd.n913 gnd.n912 585
R957 gnd.n6461 gnd.n913 585
R958 gnd.n6459 gnd.n6458 585
R959 gnd.n6460 gnd.n6459 585
R960 gnd.n6457 gnd.n915 585
R961 gnd.n915 gnd.n914 585
R962 gnd.n6456 gnd.n6455 585
R963 gnd.n6455 gnd.n6454 585
R964 gnd.n921 gnd.n920 585
R965 gnd.n6453 gnd.n921 585
R966 gnd.n6451 gnd.n6450 585
R967 gnd.n6452 gnd.n6451 585
R968 gnd.n6449 gnd.n923 585
R969 gnd.n923 gnd.n922 585
R970 gnd.n6448 gnd.n6447 585
R971 gnd.n6447 gnd.n6446 585
R972 gnd.n929 gnd.n928 585
R973 gnd.n6445 gnd.n929 585
R974 gnd.n6443 gnd.n6442 585
R975 gnd.n6444 gnd.n6443 585
R976 gnd.n6441 gnd.n931 585
R977 gnd.n931 gnd.n930 585
R978 gnd.n6440 gnd.n6439 585
R979 gnd.n6439 gnd.n6438 585
R980 gnd.n937 gnd.n936 585
R981 gnd.n6437 gnd.n937 585
R982 gnd.n6435 gnd.n6434 585
R983 gnd.n6436 gnd.n6435 585
R984 gnd.n6433 gnd.n939 585
R985 gnd.n939 gnd.n938 585
R986 gnd.n6432 gnd.n6431 585
R987 gnd.n6431 gnd.n6430 585
R988 gnd.n945 gnd.n944 585
R989 gnd.n6429 gnd.n945 585
R990 gnd.n6427 gnd.n6426 585
R991 gnd.n6428 gnd.n6427 585
R992 gnd.n6425 gnd.n947 585
R993 gnd.n947 gnd.n946 585
R994 gnd.n6424 gnd.n6423 585
R995 gnd.n6423 gnd.n6422 585
R996 gnd.n953 gnd.n952 585
R997 gnd.n6421 gnd.n953 585
R998 gnd.n6419 gnd.n6418 585
R999 gnd.n6420 gnd.n6419 585
R1000 gnd.n6417 gnd.n955 585
R1001 gnd.n955 gnd.n954 585
R1002 gnd.n6416 gnd.n6415 585
R1003 gnd.n6415 gnd.n6414 585
R1004 gnd.n961 gnd.n960 585
R1005 gnd.n6413 gnd.n961 585
R1006 gnd.n6411 gnd.n6410 585
R1007 gnd.n6412 gnd.n6411 585
R1008 gnd.n6581 gnd.n6580 585
R1009 gnd.n6582 gnd.n6581 585
R1010 gnd.n796 gnd.n795 585
R1011 gnd.n6583 gnd.n796 585
R1012 gnd.n6586 gnd.n6585 585
R1013 gnd.n6585 gnd.n6584 585
R1014 gnd.n793 gnd.n792 585
R1015 gnd.n792 gnd.n791 585
R1016 gnd.n6591 gnd.n6590 585
R1017 gnd.n6592 gnd.n6591 585
R1018 gnd.n790 gnd.n789 585
R1019 gnd.n6593 gnd.n790 585
R1020 gnd.n6596 gnd.n6595 585
R1021 gnd.n6595 gnd.n6594 585
R1022 gnd.n787 gnd.n786 585
R1023 gnd.n786 gnd.n785 585
R1024 gnd.n6601 gnd.n6600 585
R1025 gnd.n6602 gnd.n6601 585
R1026 gnd.n784 gnd.n783 585
R1027 gnd.n6603 gnd.n784 585
R1028 gnd.n6606 gnd.n6605 585
R1029 gnd.n6605 gnd.n6604 585
R1030 gnd.n781 gnd.n780 585
R1031 gnd.n780 gnd.n779 585
R1032 gnd.n6611 gnd.n6610 585
R1033 gnd.n6612 gnd.n6611 585
R1034 gnd.n778 gnd.n777 585
R1035 gnd.n6613 gnd.n778 585
R1036 gnd.n6616 gnd.n6615 585
R1037 gnd.n6615 gnd.n6614 585
R1038 gnd.n775 gnd.n774 585
R1039 gnd.n774 gnd.n773 585
R1040 gnd.n6621 gnd.n6620 585
R1041 gnd.n6622 gnd.n6621 585
R1042 gnd.n772 gnd.n771 585
R1043 gnd.n6623 gnd.n772 585
R1044 gnd.n6626 gnd.n6625 585
R1045 gnd.n6625 gnd.n6624 585
R1046 gnd.n769 gnd.n768 585
R1047 gnd.n768 gnd.n767 585
R1048 gnd.n6631 gnd.n6630 585
R1049 gnd.n6632 gnd.n6631 585
R1050 gnd.n766 gnd.n765 585
R1051 gnd.n6633 gnd.n766 585
R1052 gnd.n6636 gnd.n6635 585
R1053 gnd.n6635 gnd.n6634 585
R1054 gnd.n763 gnd.n762 585
R1055 gnd.n762 gnd.n761 585
R1056 gnd.n6641 gnd.n6640 585
R1057 gnd.n6642 gnd.n6641 585
R1058 gnd.n760 gnd.n759 585
R1059 gnd.n6643 gnd.n760 585
R1060 gnd.n6646 gnd.n6645 585
R1061 gnd.n6645 gnd.n6644 585
R1062 gnd.n757 gnd.n756 585
R1063 gnd.n756 gnd.n755 585
R1064 gnd.n6651 gnd.n6650 585
R1065 gnd.n6652 gnd.n6651 585
R1066 gnd.n754 gnd.n753 585
R1067 gnd.n6653 gnd.n754 585
R1068 gnd.n6656 gnd.n6655 585
R1069 gnd.n6655 gnd.n6654 585
R1070 gnd.n751 gnd.n750 585
R1071 gnd.n750 gnd.n749 585
R1072 gnd.n6661 gnd.n6660 585
R1073 gnd.n6662 gnd.n6661 585
R1074 gnd.n748 gnd.n747 585
R1075 gnd.n6663 gnd.n748 585
R1076 gnd.n6666 gnd.n6665 585
R1077 gnd.n6665 gnd.n6664 585
R1078 gnd.n745 gnd.n744 585
R1079 gnd.n744 gnd.n743 585
R1080 gnd.n6671 gnd.n6670 585
R1081 gnd.n6672 gnd.n6671 585
R1082 gnd.n742 gnd.n741 585
R1083 gnd.n6673 gnd.n742 585
R1084 gnd.n6676 gnd.n6675 585
R1085 gnd.n6675 gnd.n6674 585
R1086 gnd.n739 gnd.n738 585
R1087 gnd.n738 gnd.n737 585
R1088 gnd.n6681 gnd.n6680 585
R1089 gnd.n6682 gnd.n6681 585
R1090 gnd.n736 gnd.n735 585
R1091 gnd.n6683 gnd.n736 585
R1092 gnd.n6686 gnd.n6685 585
R1093 gnd.n6685 gnd.n6684 585
R1094 gnd.n733 gnd.n732 585
R1095 gnd.n732 gnd.n731 585
R1096 gnd.n6691 gnd.n6690 585
R1097 gnd.n6692 gnd.n6691 585
R1098 gnd.n730 gnd.n729 585
R1099 gnd.n6693 gnd.n730 585
R1100 gnd.n6696 gnd.n6695 585
R1101 gnd.n6695 gnd.n6694 585
R1102 gnd.n727 gnd.n726 585
R1103 gnd.n726 gnd.n725 585
R1104 gnd.n6701 gnd.n6700 585
R1105 gnd.n6702 gnd.n6701 585
R1106 gnd.n724 gnd.n723 585
R1107 gnd.n6703 gnd.n724 585
R1108 gnd.n6706 gnd.n6705 585
R1109 gnd.n6705 gnd.n6704 585
R1110 gnd.n721 gnd.n720 585
R1111 gnd.n720 gnd.n719 585
R1112 gnd.n6711 gnd.n6710 585
R1113 gnd.n6712 gnd.n6711 585
R1114 gnd.n718 gnd.n717 585
R1115 gnd.n6713 gnd.n718 585
R1116 gnd.n6716 gnd.n6715 585
R1117 gnd.n6715 gnd.n6714 585
R1118 gnd.n715 gnd.n714 585
R1119 gnd.n714 gnd.n713 585
R1120 gnd.n6721 gnd.n6720 585
R1121 gnd.n6722 gnd.n6721 585
R1122 gnd.n712 gnd.n711 585
R1123 gnd.n6723 gnd.n712 585
R1124 gnd.n6726 gnd.n6725 585
R1125 gnd.n6725 gnd.n6724 585
R1126 gnd.n709 gnd.n708 585
R1127 gnd.n708 gnd.n707 585
R1128 gnd.n6731 gnd.n6730 585
R1129 gnd.n6732 gnd.n6731 585
R1130 gnd.n706 gnd.n705 585
R1131 gnd.n6733 gnd.n706 585
R1132 gnd.n6736 gnd.n6735 585
R1133 gnd.n6735 gnd.n6734 585
R1134 gnd.n703 gnd.n702 585
R1135 gnd.n702 gnd.n701 585
R1136 gnd.n6741 gnd.n6740 585
R1137 gnd.n6742 gnd.n6741 585
R1138 gnd.n700 gnd.n699 585
R1139 gnd.n6743 gnd.n700 585
R1140 gnd.n6746 gnd.n6745 585
R1141 gnd.n6745 gnd.n6744 585
R1142 gnd.n697 gnd.n696 585
R1143 gnd.n696 gnd.n695 585
R1144 gnd.n6751 gnd.n6750 585
R1145 gnd.n6752 gnd.n6751 585
R1146 gnd.n694 gnd.n693 585
R1147 gnd.n6753 gnd.n694 585
R1148 gnd.n6756 gnd.n6755 585
R1149 gnd.n6755 gnd.n6754 585
R1150 gnd.n691 gnd.n690 585
R1151 gnd.n690 gnd.n689 585
R1152 gnd.n6761 gnd.n6760 585
R1153 gnd.n6762 gnd.n6761 585
R1154 gnd.n688 gnd.n687 585
R1155 gnd.n6763 gnd.n688 585
R1156 gnd.n6766 gnd.n6765 585
R1157 gnd.n6765 gnd.n6764 585
R1158 gnd.n685 gnd.n684 585
R1159 gnd.n684 gnd.n683 585
R1160 gnd.n6771 gnd.n6770 585
R1161 gnd.n6772 gnd.n6771 585
R1162 gnd.n682 gnd.n681 585
R1163 gnd.n6773 gnd.n682 585
R1164 gnd.n6776 gnd.n6775 585
R1165 gnd.n6775 gnd.n6774 585
R1166 gnd.n679 gnd.n678 585
R1167 gnd.n678 gnd.n677 585
R1168 gnd.n6781 gnd.n6780 585
R1169 gnd.n6782 gnd.n6781 585
R1170 gnd.n676 gnd.n675 585
R1171 gnd.n6783 gnd.n676 585
R1172 gnd.n6786 gnd.n6785 585
R1173 gnd.n6785 gnd.n6784 585
R1174 gnd.n673 gnd.n672 585
R1175 gnd.n672 gnd.n671 585
R1176 gnd.n6791 gnd.n6790 585
R1177 gnd.n6792 gnd.n6791 585
R1178 gnd.n670 gnd.n669 585
R1179 gnd.n6793 gnd.n670 585
R1180 gnd.n6796 gnd.n6795 585
R1181 gnd.n6795 gnd.n6794 585
R1182 gnd.n667 gnd.n666 585
R1183 gnd.n666 gnd.n665 585
R1184 gnd.n6801 gnd.n6800 585
R1185 gnd.n6802 gnd.n6801 585
R1186 gnd.n664 gnd.n663 585
R1187 gnd.n6803 gnd.n664 585
R1188 gnd.n6806 gnd.n6805 585
R1189 gnd.n6805 gnd.n6804 585
R1190 gnd.n661 gnd.n660 585
R1191 gnd.n660 gnd.n659 585
R1192 gnd.n6811 gnd.n6810 585
R1193 gnd.n6812 gnd.n6811 585
R1194 gnd.n658 gnd.n657 585
R1195 gnd.n6813 gnd.n658 585
R1196 gnd.n6816 gnd.n6815 585
R1197 gnd.n6815 gnd.n6814 585
R1198 gnd.n655 gnd.n654 585
R1199 gnd.n654 gnd.n653 585
R1200 gnd.n6821 gnd.n6820 585
R1201 gnd.n6822 gnd.n6821 585
R1202 gnd.n652 gnd.n651 585
R1203 gnd.n6823 gnd.n652 585
R1204 gnd.n6826 gnd.n6825 585
R1205 gnd.n6825 gnd.n6824 585
R1206 gnd.n649 gnd.n648 585
R1207 gnd.n648 gnd.n647 585
R1208 gnd.n6831 gnd.n6830 585
R1209 gnd.n6832 gnd.n6831 585
R1210 gnd.n646 gnd.n645 585
R1211 gnd.n6833 gnd.n646 585
R1212 gnd.n6836 gnd.n6835 585
R1213 gnd.n6835 gnd.n6834 585
R1214 gnd.n643 gnd.n642 585
R1215 gnd.n642 gnd.n641 585
R1216 gnd.n6841 gnd.n6840 585
R1217 gnd.n6842 gnd.n6841 585
R1218 gnd.n640 gnd.n639 585
R1219 gnd.n6843 gnd.n640 585
R1220 gnd.n6846 gnd.n6845 585
R1221 gnd.n6845 gnd.n6844 585
R1222 gnd.n637 gnd.n636 585
R1223 gnd.n636 gnd.n635 585
R1224 gnd.n6851 gnd.n6850 585
R1225 gnd.n6852 gnd.n6851 585
R1226 gnd.n634 gnd.n633 585
R1227 gnd.n6853 gnd.n634 585
R1228 gnd.n6856 gnd.n6855 585
R1229 gnd.n6855 gnd.n6854 585
R1230 gnd.n631 gnd.n630 585
R1231 gnd.n630 gnd.n629 585
R1232 gnd.n6861 gnd.n6860 585
R1233 gnd.n6862 gnd.n6861 585
R1234 gnd.n628 gnd.n627 585
R1235 gnd.n6863 gnd.n628 585
R1236 gnd.n6866 gnd.n6865 585
R1237 gnd.n6865 gnd.n6864 585
R1238 gnd.n625 gnd.n624 585
R1239 gnd.n624 gnd.n623 585
R1240 gnd.n6871 gnd.n6870 585
R1241 gnd.n6872 gnd.n6871 585
R1242 gnd.n622 gnd.n621 585
R1243 gnd.n6873 gnd.n622 585
R1244 gnd.n6876 gnd.n6875 585
R1245 gnd.n6875 gnd.n6874 585
R1246 gnd.n619 gnd.n618 585
R1247 gnd.n618 gnd.n617 585
R1248 gnd.n6881 gnd.n6880 585
R1249 gnd.n6882 gnd.n6881 585
R1250 gnd.n616 gnd.n615 585
R1251 gnd.n6883 gnd.n616 585
R1252 gnd.n6886 gnd.n6885 585
R1253 gnd.n6885 gnd.n6884 585
R1254 gnd.n613 gnd.n612 585
R1255 gnd.n612 gnd.n611 585
R1256 gnd.n6891 gnd.n6890 585
R1257 gnd.n6892 gnd.n6891 585
R1258 gnd.n610 gnd.n609 585
R1259 gnd.n6893 gnd.n610 585
R1260 gnd.n6896 gnd.n6895 585
R1261 gnd.n6895 gnd.n6894 585
R1262 gnd.n607 gnd.n606 585
R1263 gnd.n606 gnd.n605 585
R1264 gnd.n6901 gnd.n6900 585
R1265 gnd.n6902 gnd.n6901 585
R1266 gnd.n604 gnd.n603 585
R1267 gnd.n6903 gnd.n604 585
R1268 gnd.n6906 gnd.n6905 585
R1269 gnd.n6905 gnd.n6904 585
R1270 gnd.n601 gnd.n600 585
R1271 gnd.n600 gnd.n599 585
R1272 gnd.n6911 gnd.n6910 585
R1273 gnd.n6912 gnd.n6911 585
R1274 gnd.n598 gnd.n597 585
R1275 gnd.n6913 gnd.n598 585
R1276 gnd.n6916 gnd.n6915 585
R1277 gnd.n6915 gnd.n6914 585
R1278 gnd.n595 gnd.n594 585
R1279 gnd.n594 gnd.n593 585
R1280 gnd.n6921 gnd.n6920 585
R1281 gnd.n6922 gnd.n6921 585
R1282 gnd.n592 gnd.n591 585
R1283 gnd.n6923 gnd.n592 585
R1284 gnd.n6926 gnd.n6925 585
R1285 gnd.n6925 gnd.n6924 585
R1286 gnd.n589 gnd.n588 585
R1287 gnd.n588 gnd.n587 585
R1288 gnd.n6931 gnd.n6930 585
R1289 gnd.n6932 gnd.n6931 585
R1290 gnd.n586 gnd.n585 585
R1291 gnd.n6933 gnd.n586 585
R1292 gnd.n6936 gnd.n6935 585
R1293 gnd.n6935 gnd.n6934 585
R1294 gnd.n583 gnd.n582 585
R1295 gnd.n582 gnd.n581 585
R1296 gnd.n6941 gnd.n6940 585
R1297 gnd.n6942 gnd.n6941 585
R1298 gnd.n580 gnd.n579 585
R1299 gnd.n6943 gnd.n580 585
R1300 gnd.n6946 gnd.n6945 585
R1301 gnd.n6945 gnd.n6944 585
R1302 gnd.n577 gnd.n576 585
R1303 gnd.n576 gnd.n575 585
R1304 gnd.n6951 gnd.n6950 585
R1305 gnd.n6952 gnd.n6951 585
R1306 gnd.n574 gnd.n573 585
R1307 gnd.n6953 gnd.n574 585
R1308 gnd.n6956 gnd.n6955 585
R1309 gnd.n6955 gnd.n6954 585
R1310 gnd.n571 gnd.n570 585
R1311 gnd.n570 gnd.n569 585
R1312 gnd.n6961 gnd.n6960 585
R1313 gnd.n6962 gnd.n6961 585
R1314 gnd.n568 gnd.n567 585
R1315 gnd.n6963 gnd.n568 585
R1316 gnd.n6966 gnd.n6965 585
R1317 gnd.n6965 gnd.n6964 585
R1318 gnd.n565 gnd.n564 585
R1319 gnd.n564 gnd.n563 585
R1320 gnd.n6971 gnd.n6970 585
R1321 gnd.n6972 gnd.n6971 585
R1322 gnd.n562 gnd.n561 585
R1323 gnd.n6973 gnd.n562 585
R1324 gnd.n6976 gnd.n6975 585
R1325 gnd.n6975 gnd.n6974 585
R1326 gnd.n559 gnd.n558 585
R1327 gnd.n558 gnd.n557 585
R1328 gnd.n6981 gnd.n6980 585
R1329 gnd.n6982 gnd.n6981 585
R1330 gnd.n556 gnd.n555 585
R1331 gnd.n6983 gnd.n556 585
R1332 gnd.n6986 gnd.n6985 585
R1333 gnd.n6985 gnd.n6984 585
R1334 gnd.n553 gnd.n552 585
R1335 gnd.n552 gnd.n551 585
R1336 gnd.n6992 gnd.n6991 585
R1337 gnd.n6993 gnd.n6992 585
R1338 gnd.n550 gnd.n549 585
R1339 gnd.n6994 gnd.n550 585
R1340 gnd.n6997 gnd.n6996 585
R1341 gnd.n6996 gnd.n6995 585
R1342 gnd.n6998 gnd.n547 585
R1343 gnd.n547 gnd.n546 585
R1344 gnd.n422 gnd.n421 585
R1345 gnd.n7205 gnd.n421 585
R1346 gnd.n7208 gnd.n7207 585
R1347 gnd.n7207 gnd.n7206 585
R1348 gnd.n425 gnd.n424 585
R1349 gnd.n7204 gnd.n425 585
R1350 gnd.n7202 gnd.n7201 585
R1351 gnd.n7203 gnd.n7202 585
R1352 gnd.n428 gnd.n427 585
R1353 gnd.n427 gnd.n426 585
R1354 gnd.n7197 gnd.n7196 585
R1355 gnd.n7196 gnd.n7195 585
R1356 gnd.n431 gnd.n430 585
R1357 gnd.n7194 gnd.n431 585
R1358 gnd.n7192 gnd.n7191 585
R1359 gnd.n7193 gnd.n7192 585
R1360 gnd.n434 gnd.n433 585
R1361 gnd.n433 gnd.n432 585
R1362 gnd.n7187 gnd.n7186 585
R1363 gnd.n7186 gnd.n7185 585
R1364 gnd.n437 gnd.n436 585
R1365 gnd.n7184 gnd.n437 585
R1366 gnd.n7182 gnd.n7181 585
R1367 gnd.n7183 gnd.n7182 585
R1368 gnd.n440 gnd.n439 585
R1369 gnd.n439 gnd.n438 585
R1370 gnd.n7177 gnd.n7176 585
R1371 gnd.n7176 gnd.n7175 585
R1372 gnd.n443 gnd.n442 585
R1373 gnd.n7174 gnd.n443 585
R1374 gnd.n7172 gnd.n7171 585
R1375 gnd.n7173 gnd.n7172 585
R1376 gnd.n446 gnd.n445 585
R1377 gnd.n445 gnd.n444 585
R1378 gnd.n7167 gnd.n7166 585
R1379 gnd.n7166 gnd.n7165 585
R1380 gnd.n449 gnd.n448 585
R1381 gnd.n7164 gnd.n449 585
R1382 gnd.n7162 gnd.n7161 585
R1383 gnd.n7163 gnd.n7162 585
R1384 gnd.n452 gnd.n451 585
R1385 gnd.n451 gnd.n450 585
R1386 gnd.n7157 gnd.n7156 585
R1387 gnd.n7156 gnd.n7155 585
R1388 gnd.n455 gnd.n454 585
R1389 gnd.n7154 gnd.n455 585
R1390 gnd.n7152 gnd.n7151 585
R1391 gnd.n7153 gnd.n7152 585
R1392 gnd.n458 gnd.n457 585
R1393 gnd.n457 gnd.n456 585
R1394 gnd.n7147 gnd.n7146 585
R1395 gnd.n7146 gnd.n7145 585
R1396 gnd.n461 gnd.n460 585
R1397 gnd.n7144 gnd.n461 585
R1398 gnd.n7142 gnd.n7141 585
R1399 gnd.n7143 gnd.n7142 585
R1400 gnd.n464 gnd.n463 585
R1401 gnd.n463 gnd.n462 585
R1402 gnd.n7137 gnd.n7136 585
R1403 gnd.n7136 gnd.n7135 585
R1404 gnd.n467 gnd.n466 585
R1405 gnd.n7134 gnd.n467 585
R1406 gnd.n7132 gnd.n7131 585
R1407 gnd.n7133 gnd.n7132 585
R1408 gnd.n470 gnd.n469 585
R1409 gnd.n469 gnd.n468 585
R1410 gnd.n7127 gnd.n7126 585
R1411 gnd.n7126 gnd.n7125 585
R1412 gnd.n473 gnd.n472 585
R1413 gnd.n7124 gnd.n473 585
R1414 gnd.n7122 gnd.n7121 585
R1415 gnd.n7123 gnd.n7122 585
R1416 gnd.n476 gnd.n475 585
R1417 gnd.n475 gnd.n474 585
R1418 gnd.n7117 gnd.n7116 585
R1419 gnd.n7116 gnd.n7115 585
R1420 gnd.n479 gnd.n478 585
R1421 gnd.n7114 gnd.n479 585
R1422 gnd.n7112 gnd.n7111 585
R1423 gnd.n7113 gnd.n7112 585
R1424 gnd.n482 gnd.n481 585
R1425 gnd.n481 gnd.n480 585
R1426 gnd.n7107 gnd.n7106 585
R1427 gnd.n7106 gnd.n7105 585
R1428 gnd.n485 gnd.n484 585
R1429 gnd.n7104 gnd.n485 585
R1430 gnd.n7102 gnd.n7101 585
R1431 gnd.n7103 gnd.n7102 585
R1432 gnd.n488 gnd.n487 585
R1433 gnd.n487 gnd.n486 585
R1434 gnd.n7097 gnd.n7096 585
R1435 gnd.n7096 gnd.n7095 585
R1436 gnd.n491 gnd.n490 585
R1437 gnd.n7094 gnd.n491 585
R1438 gnd.n7092 gnd.n7091 585
R1439 gnd.n7093 gnd.n7092 585
R1440 gnd.n494 gnd.n493 585
R1441 gnd.n493 gnd.n492 585
R1442 gnd.n7087 gnd.n7086 585
R1443 gnd.n7086 gnd.n7085 585
R1444 gnd.n497 gnd.n496 585
R1445 gnd.n7084 gnd.n497 585
R1446 gnd.n7082 gnd.n7081 585
R1447 gnd.n7083 gnd.n7082 585
R1448 gnd.n500 gnd.n499 585
R1449 gnd.n499 gnd.n498 585
R1450 gnd.n7077 gnd.n7076 585
R1451 gnd.n7076 gnd.n7075 585
R1452 gnd.n503 gnd.n502 585
R1453 gnd.n7074 gnd.n503 585
R1454 gnd.n7072 gnd.n7071 585
R1455 gnd.n7073 gnd.n7072 585
R1456 gnd.n506 gnd.n505 585
R1457 gnd.n505 gnd.n504 585
R1458 gnd.n7067 gnd.n7066 585
R1459 gnd.n7066 gnd.n7065 585
R1460 gnd.n509 gnd.n508 585
R1461 gnd.n7064 gnd.n509 585
R1462 gnd.n7062 gnd.n7061 585
R1463 gnd.n7063 gnd.n7062 585
R1464 gnd.n512 gnd.n511 585
R1465 gnd.n511 gnd.n510 585
R1466 gnd.n7057 gnd.n7056 585
R1467 gnd.n7056 gnd.n7055 585
R1468 gnd.n515 gnd.n514 585
R1469 gnd.n7054 gnd.n515 585
R1470 gnd.n7052 gnd.n7051 585
R1471 gnd.n7053 gnd.n7052 585
R1472 gnd.n518 gnd.n517 585
R1473 gnd.n517 gnd.n516 585
R1474 gnd.n7047 gnd.n7046 585
R1475 gnd.n7046 gnd.n7045 585
R1476 gnd.n521 gnd.n520 585
R1477 gnd.n7044 gnd.n521 585
R1478 gnd.n7042 gnd.n7041 585
R1479 gnd.n7043 gnd.n7042 585
R1480 gnd.n524 gnd.n523 585
R1481 gnd.n523 gnd.n522 585
R1482 gnd.n7037 gnd.n7036 585
R1483 gnd.n7036 gnd.n7035 585
R1484 gnd.n527 gnd.n526 585
R1485 gnd.n7034 gnd.n527 585
R1486 gnd.n7032 gnd.n7031 585
R1487 gnd.n7033 gnd.n7032 585
R1488 gnd.n530 gnd.n529 585
R1489 gnd.n529 gnd.n528 585
R1490 gnd.n7027 gnd.n7026 585
R1491 gnd.n7026 gnd.n7025 585
R1492 gnd.n533 gnd.n532 585
R1493 gnd.n7024 gnd.n533 585
R1494 gnd.n7022 gnd.n7021 585
R1495 gnd.n7023 gnd.n7022 585
R1496 gnd.n536 gnd.n535 585
R1497 gnd.n535 gnd.n534 585
R1498 gnd.n7017 gnd.n7016 585
R1499 gnd.n7016 gnd.n7015 585
R1500 gnd.n539 gnd.n538 585
R1501 gnd.n7014 gnd.n539 585
R1502 gnd.n7012 gnd.n7011 585
R1503 gnd.n7013 gnd.n7012 585
R1504 gnd.n542 gnd.n541 585
R1505 gnd.n541 gnd.n540 585
R1506 gnd.n7007 gnd.n7006 585
R1507 gnd.n7006 gnd.n7005 585
R1508 gnd.n545 gnd.n544 585
R1509 gnd.n7004 gnd.n545 585
R1510 gnd.n7002 gnd.n7001 585
R1511 gnd.n7003 gnd.n7002 585
R1512 gnd.n6323 gnd.n6322 585
R1513 gnd.n6324 gnd.n6323 585
R1514 gnd.n1099 gnd.n1098 585
R1515 gnd.n4568 gnd.n1099 585
R1516 gnd.n6332 gnd.n6331 585
R1517 gnd.n6331 gnd.n6330 585
R1518 gnd.n6333 gnd.n1093 585
R1519 gnd.n4530 gnd.n1093 585
R1520 gnd.n6335 gnd.n6334 585
R1521 gnd.n6336 gnd.n6335 585
R1522 gnd.n1078 gnd.n1077 585
R1523 gnd.n4521 gnd.n1078 585
R1524 gnd.n6344 gnd.n6343 585
R1525 gnd.n6343 gnd.n6342 585
R1526 gnd.n6345 gnd.n1072 585
R1527 gnd.n4513 gnd.n1072 585
R1528 gnd.n6347 gnd.n6346 585
R1529 gnd.n6348 gnd.n6347 585
R1530 gnd.n1056 gnd.n1055 585
R1531 gnd.n4451 gnd.n1056 585
R1532 gnd.n6356 gnd.n6355 585
R1533 gnd.n6355 gnd.n6354 585
R1534 gnd.n6357 gnd.n1050 585
R1535 gnd.n4439 gnd.n1050 585
R1536 gnd.n6359 gnd.n6358 585
R1537 gnd.n6360 gnd.n6359 585
R1538 gnd.n1036 gnd.n1035 585
R1539 gnd.n4462 gnd.n1036 585
R1540 gnd.n6368 gnd.n6367 585
R1541 gnd.n6367 gnd.n6366 585
R1542 gnd.n6369 gnd.n1030 585
R1543 gnd.n4431 gnd.n1030 585
R1544 gnd.n6371 gnd.n6370 585
R1545 gnd.n6372 gnd.n6371 585
R1546 gnd.n1014 gnd.n1013 585
R1547 gnd.n4398 gnd.n1014 585
R1548 gnd.n6380 gnd.n6379 585
R1549 gnd.n6379 gnd.n6378 585
R1550 gnd.n6381 gnd.n1008 585
R1551 gnd.n4390 gnd.n1008 585
R1552 gnd.n6383 gnd.n6382 585
R1553 gnd.n6384 gnd.n6383 585
R1554 gnd.n994 gnd.n993 585
R1555 gnd.n4413 gnd.n994 585
R1556 gnd.n6392 gnd.n6391 585
R1557 gnd.n6391 gnd.n6390 585
R1558 gnd.n6393 gnd.n988 585
R1559 gnd.n4382 gnd.n988 585
R1560 gnd.n6395 gnd.n6394 585
R1561 gnd.n6396 gnd.n6395 585
R1562 gnd.n989 gnd.n987 585
R1563 gnd.n4364 gnd.n987 585
R1564 gnd.n4341 gnd.n974 585
R1565 gnd.n6402 gnd.n974 585
R1566 gnd.n4343 gnd.n4342 585
R1567 gnd.n4342 gnd.n970 585
R1568 gnd.n4344 gnd.n2191 585
R1569 gnd.n4355 gnd.n2191 585
R1570 gnd.n4345 gnd.n2200 585
R1571 gnd.n2200 gnd.n2198 585
R1572 gnd.n4347 gnd.n4346 585
R1573 gnd.n4348 gnd.n4347 585
R1574 gnd.n2201 gnd.n2199 585
R1575 gnd.n2216 gnd.n2199 585
R1576 gnd.n2217 gnd.n2203 585
R1577 gnd.n4329 gnd.n2217 585
R1578 gnd.n4318 gnd.n2225 585
R1579 gnd.n2225 gnd.n2214 585
R1580 gnd.n4320 gnd.n4319 585
R1581 gnd.n4321 gnd.n4320 585
R1582 gnd.n2226 gnd.n2224 585
R1583 gnd.n2224 gnd.n2221 585
R1584 gnd.n4314 gnd.n4313 585
R1585 gnd.n4313 gnd.n4312 585
R1586 gnd.n2229 gnd.n2228 585
R1587 gnd.n2230 gnd.n2229 585
R1588 gnd.n4303 gnd.n4302 585
R1589 gnd.n4304 gnd.n4303 585
R1590 gnd.n2240 gnd.n2239 585
R1591 gnd.n2247 gnd.n2239 585
R1592 gnd.n4298 gnd.n4297 585
R1593 gnd.n4297 gnd.n4296 585
R1594 gnd.n2243 gnd.n2242 585
R1595 gnd.n2244 gnd.n2243 585
R1596 gnd.n4286 gnd.n4285 585
R1597 gnd.n4287 gnd.n4286 585
R1598 gnd.n2257 gnd.n2256 585
R1599 gnd.n2256 gnd.n2253 585
R1600 gnd.n4281 gnd.n4280 585
R1601 gnd.n4280 gnd.n4279 585
R1602 gnd.n2260 gnd.n2259 585
R1603 gnd.n2261 gnd.n2260 585
R1604 gnd.n4270 gnd.n4269 585
R1605 gnd.n4271 gnd.n4270 585
R1606 gnd.n2272 gnd.n2271 585
R1607 gnd.n2279 gnd.n2271 585
R1608 gnd.n4265 gnd.n4264 585
R1609 gnd.n4264 gnd.n4263 585
R1610 gnd.n2275 gnd.n2274 585
R1611 gnd.n2276 gnd.n2275 585
R1612 gnd.n4254 gnd.n4253 585
R1613 gnd.n4255 gnd.n4254 585
R1614 gnd.n2289 gnd.n2288 585
R1615 gnd.n2288 gnd.n2285 585
R1616 gnd.n4249 gnd.n4248 585
R1617 gnd.n4248 gnd.n4247 585
R1618 gnd.n2292 gnd.n2291 585
R1619 gnd.n2293 gnd.n2292 585
R1620 gnd.n4238 gnd.n4237 585
R1621 gnd.n4239 gnd.n4238 585
R1622 gnd.n2304 gnd.n2303 585
R1623 gnd.n2311 gnd.n2303 585
R1624 gnd.n4233 gnd.n4232 585
R1625 gnd.n4232 gnd.n4231 585
R1626 gnd.n2307 gnd.n2306 585
R1627 gnd.n2308 gnd.n2307 585
R1628 gnd.n4222 gnd.n4221 585
R1629 gnd.n4223 gnd.n4222 585
R1630 gnd.n2321 gnd.n2320 585
R1631 gnd.n2320 gnd.n2317 585
R1632 gnd.n4217 gnd.n4216 585
R1633 gnd.n4216 gnd.n4215 585
R1634 gnd.n2324 gnd.n2323 585
R1635 gnd.n2325 gnd.n2324 585
R1636 gnd.n4206 gnd.n4205 585
R1637 gnd.n4207 gnd.n4206 585
R1638 gnd.n2336 gnd.n2335 585
R1639 gnd.n3977 gnd.n2335 585
R1640 gnd.n4201 gnd.n4200 585
R1641 gnd.n4200 gnd.n4199 585
R1642 gnd.n3836 gnd.n2338 585
R1643 gnd.n3839 gnd.n3837 585
R1644 gnd.n3842 gnd.n3841 585
R1645 gnd.n3834 gnd.n3833 585
R1646 gnd.n3847 gnd.n3846 585
R1647 gnd.n3849 gnd.n3832 585
R1648 gnd.n3852 gnd.n3851 585
R1649 gnd.n3830 gnd.n3829 585
R1650 gnd.n3857 gnd.n3856 585
R1651 gnd.n3859 gnd.n3828 585
R1652 gnd.n3862 gnd.n3861 585
R1653 gnd.n3826 gnd.n3825 585
R1654 gnd.n3867 gnd.n3866 585
R1655 gnd.n3869 gnd.n3824 585
R1656 gnd.n3872 gnd.n3871 585
R1657 gnd.n3822 gnd.n3821 585
R1658 gnd.n3877 gnd.n3876 585
R1659 gnd.n3879 gnd.n3820 585
R1660 gnd.n3881 gnd.n3880 585
R1661 gnd.n3880 gnd.n3813 585
R1662 gnd.n4850 gnd.n4849 585
R1663 gnd.n2046 gnd.n2038 585
R1664 gnd.n4857 gnd.n2035 585
R1665 gnd.n4858 gnd.n2034 585
R1666 gnd.n2060 gnd.n2028 585
R1667 gnd.n4865 gnd.n2027 585
R1668 gnd.n4866 gnd.n2026 585
R1669 gnd.n2058 gnd.n2018 585
R1670 gnd.n4873 gnd.n2017 585
R1671 gnd.n4874 gnd.n2016 585
R1672 gnd.n2055 gnd.n2010 585
R1673 gnd.n4881 gnd.n2009 585
R1674 gnd.n4882 gnd.n2008 585
R1675 gnd.n2053 gnd.n2001 585
R1676 gnd.n4889 gnd.n2000 585
R1677 gnd.n4890 gnd.n1999 585
R1678 gnd.n2050 gnd.n1998 585
R1679 gnd.n2049 gnd.n2048 585
R1680 gnd.n1115 gnd.n1113 585
R1681 gnd.n4847 gnd.n1113 585
R1682 gnd.n2131 gnd.n1111 585
R1683 gnd.n6324 gnd.n1111 585
R1684 gnd.n4567 gnd.n4566 585
R1685 gnd.n4568 gnd.n4567 585
R1686 gnd.n2130 gnd.n1102 585
R1687 gnd.n6330 gnd.n1102 585
R1688 gnd.n4532 gnd.n4531 585
R1689 gnd.n4531 gnd.n4530 585
R1690 gnd.n2133 gnd.n1091 585
R1691 gnd.n6336 gnd.n1091 585
R1692 gnd.n4520 gnd.n4519 585
R1693 gnd.n4521 gnd.n4520 585
R1694 gnd.n2137 gnd.n1080 585
R1695 gnd.n6342 gnd.n1080 585
R1696 gnd.n4515 gnd.n4514 585
R1697 gnd.n4514 gnd.n4513 585
R1698 gnd.n2139 gnd.n1070 585
R1699 gnd.n6348 gnd.n1070 585
R1700 gnd.n4454 gnd.n4452 585
R1701 gnd.n4452 gnd.n4451 585
R1702 gnd.n4455 gnd.n1059 585
R1703 gnd.n6354 gnd.n1059 585
R1704 gnd.n4456 gnd.n2156 585
R1705 gnd.n4439 gnd.n2156 585
R1706 gnd.n2153 gnd.n1048 585
R1707 gnd.n6360 gnd.n1048 585
R1708 gnd.n4461 gnd.n4460 585
R1709 gnd.n4462 gnd.n4461 585
R1710 gnd.n2152 gnd.n1038 585
R1711 gnd.n6366 gnd.n1038 585
R1712 gnd.n4401 gnd.n2162 585
R1713 gnd.n4431 gnd.n2162 585
R1714 gnd.n4400 gnd.n1028 585
R1715 gnd.n6372 gnd.n1028 585
R1716 gnd.n4405 gnd.n4399 585
R1717 gnd.n4399 gnd.n4398 585
R1718 gnd.n4406 gnd.n1017 585
R1719 gnd.n6378 gnd.n1017 585
R1720 gnd.n4407 gnd.n2177 585
R1721 gnd.n4390 gnd.n2177 585
R1722 gnd.n2174 gnd.n1006 585
R1723 gnd.n6384 gnd.n1006 585
R1724 gnd.n4412 gnd.n4411 585
R1725 gnd.n4413 gnd.n4412 585
R1726 gnd.n2173 gnd.n996 585
R1727 gnd.n6390 gnd.n996 585
R1728 gnd.n4371 gnd.n4370 585
R1729 gnd.n4382 gnd.n4371 585
R1730 gnd.n2183 gnd.n985 585
R1731 gnd.n6396 gnd.n985 585
R1732 gnd.n4366 gnd.n4365 585
R1733 gnd.n4365 gnd.n4364 585
R1734 gnd.n2185 gnd.n972 585
R1735 gnd.n6402 gnd.n972 585
R1736 gnd.n3920 gnd.n3919 585
R1737 gnd.n3919 gnd.n970 585
R1738 gnd.n3923 gnd.n2190 585
R1739 gnd.n4355 gnd.n2190 585
R1740 gnd.n3924 gnd.n3918 585
R1741 gnd.n3918 gnd.n2198 585
R1742 gnd.n3925 gnd.n2196 585
R1743 gnd.n4348 gnd.n2196 585
R1744 gnd.n3916 gnd.n3915 585
R1745 gnd.n3915 gnd.n2216 585
R1746 gnd.n3929 gnd.n2215 585
R1747 gnd.n4329 gnd.n2215 585
R1748 gnd.n3931 gnd.n3930 585
R1749 gnd.n3930 gnd.n2214 585
R1750 gnd.n3932 gnd.n2223 585
R1751 gnd.n4321 gnd.n2223 585
R1752 gnd.n3934 gnd.n3933 585
R1753 gnd.n3933 gnd.n2221 585
R1754 gnd.n3935 gnd.n2232 585
R1755 gnd.n4312 gnd.n2232 585
R1756 gnd.n3937 gnd.n3936 585
R1757 gnd.n3936 gnd.n2230 585
R1758 gnd.n3938 gnd.n2238 585
R1759 gnd.n4304 gnd.n2238 585
R1760 gnd.n3940 gnd.n3939 585
R1761 gnd.n3939 gnd.n2247 585
R1762 gnd.n3941 gnd.n2246 585
R1763 gnd.n4296 gnd.n2246 585
R1764 gnd.n3943 gnd.n3942 585
R1765 gnd.n3942 gnd.n2244 585
R1766 gnd.n3944 gnd.n2255 585
R1767 gnd.n4287 gnd.n2255 585
R1768 gnd.n3946 gnd.n3945 585
R1769 gnd.n3945 gnd.n2253 585
R1770 gnd.n3947 gnd.n2263 585
R1771 gnd.n4279 gnd.n2263 585
R1772 gnd.n3949 gnd.n3948 585
R1773 gnd.n3948 gnd.n2261 585
R1774 gnd.n3950 gnd.n2270 585
R1775 gnd.n4271 gnd.n2270 585
R1776 gnd.n3952 gnd.n3951 585
R1777 gnd.n3951 gnd.n2279 585
R1778 gnd.n3953 gnd.n2278 585
R1779 gnd.n4263 gnd.n2278 585
R1780 gnd.n3955 gnd.n3954 585
R1781 gnd.n3954 gnd.n2276 585
R1782 gnd.n3956 gnd.n2287 585
R1783 gnd.n4255 gnd.n2287 585
R1784 gnd.n3958 gnd.n3957 585
R1785 gnd.n3957 gnd.n2285 585
R1786 gnd.n3959 gnd.n2295 585
R1787 gnd.n4247 gnd.n2295 585
R1788 gnd.n3961 gnd.n3960 585
R1789 gnd.n3960 gnd.n2293 585
R1790 gnd.n3962 gnd.n2302 585
R1791 gnd.n4239 gnd.n2302 585
R1792 gnd.n3964 gnd.n3963 585
R1793 gnd.n3963 gnd.n2311 585
R1794 gnd.n3965 gnd.n2310 585
R1795 gnd.n4231 gnd.n2310 585
R1796 gnd.n3967 gnd.n3966 585
R1797 gnd.n3966 gnd.n2308 585
R1798 gnd.n3968 gnd.n2319 585
R1799 gnd.n4223 gnd.n2319 585
R1800 gnd.n3970 gnd.n3969 585
R1801 gnd.n3969 gnd.n2317 585
R1802 gnd.n3971 gnd.n2327 585
R1803 gnd.n4215 gnd.n2327 585
R1804 gnd.n3973 gnd.n3972 585
R1805 gnd.n3972 gnd.n2325 585
R1806 gnd.n3974 gnd.n2334 585
R1807 gnd.n4207 gnd.n2334 585
R1808 gnd.n3976 gnd.n3975 585
R1809 gnd.n3977 gnd.n3976 585
R1810 gnd.n3816 gnd.n3815 585
R1811 gnd.n4199 gnd.n3815 585
R1812 gnd.n7569 gnd.n129 585
R1813 gnd.n7665 gnd.n129 585
R1814 gnd.n7570 gnd.n7507 585
R1815 gnd.n7507 gnd.n126 585
R1816 gnd.n7571 gnd.n207 585
R1817 gnd.n7585 gnd.n207 585
R1818 gnd.n219 gnd.n217 585
R1819 gnd.n217 gnd.n206 585
R1820 gnd.n7576 gnd.n7575 585
R1821 gnd.n7577 gnd.n7576 585
R1822 gnd.n218 gnd.n216 585
R1823 gnd.n216 gnd.n213 585
R1824 gnd.n7503 gnd.n7502 585
R1825 gnd.n7502 gnd.n7501 585
R1826 gnd.n222 gnd.n221 585
R1827 gnd.n232 gnd.n222 585
R1828 gnd.n7492 gnd.n7491 585
R1829 gnd.n7493 gnd.n7492 585
R1830 gnd.n234 gnd.n233 585
R1831 gnd.n233 gnd.n229 585
R1832 gnd.n7487 gnd.n7486 585
R1833 gnd.n7486 gnd.n7485 585
R1834 gnd.n237 gnd.n236 585
R1835 gnd.n247 gnd.n237 585
R1836 gnd.n7476 gnd.n7475 585
R1837 gnd.n7477 gnd.n7476 585
R1838 gnd.n249 gnd.n248 585
R1839 gnd.n254 gnd.n248 585
R1840 gnd.n7471 gnd.n7470 585
R1841 gnd.n7470 gnd.n7469 585
R1842 gnd.n252 gnd.n251 585
R1843 gnd.n263 gnd.n252 585
R1844 gnd.n7460 gnd.n7459 585
R1845 gnd.n7461 gnd.n7460 585
R1846 gnd.n265 gnd.n264 585
R1847 gnd.n264 gnd.n260 585
R1848 gnd.n7455 gnd.n7454 585
R1849 gnd.n7454 gnd.n7453 585
R1850 gnd.n268 gnd.n267 585
R1851 gnd.n269 gnd.n268 585
R1852 gnd.n7444 gnd.n7443 585
R1853 gnd.n7445 gnd.n7444 585
R1854 gnd.n279 gnd.n278 585
R1855 gnd.n284 gnd.n278 585
R1856 gnd.n7439 gnd.n7438 585
R1857 gnd.n7438 gnd.n7437 585
R1858 gnd.n282 gnd.n281 585
R1859 gnd.n293 gnd.n282 585
R1860 gnd.n7428 gnd.n7427 585
R1861 gnd.n7429 gnd.n7428 585
R1862 gnd.n295 gnd.n294 585
R1863 gnd.n294 gnd.n290 585
R1864 gnd.n7423 gnd.n7422 585
R1865 gnd.n7422 gnd.n7421 585
R1866 gnd.n298 gnd.n297 585
R1867 gnd.n299 gnd.n298 585
R1868 gnd.n7399 gnd.n7398 585
R1869 gnd.n7398 gnd.n7397 585
R1870 gnd.n7400 gnd.n327 585
R1871 gnd.n7393 gnd.n327 585
R1872 gnd.n333 gnd.n325 585
R1873 gnd.n334 gnd.n333 585
R1874 gnd.n7404 gnd.n324 585
R1875 gnd.n7320 gnd.n324 585
R1876 gnd.n7405 gnd.n323 585
R1877 gnd.n340 gnd.n323 585
R1878 gnd.n7406 gnd.n322 585
R1879 gnd.n7314 gnd.n322 585
R1880 gnd.n319 gnd.n317 585
R1881 gnd.n317 gnd.n315 585
R1882 gnd.n7411 gnd.n7410 585
R1883 gnd.n7412 gnd.n7411 585
R1884 gnd.n318 gnd.n316 585
R1885 gnd.n7305 gnd.n316 585
R1886 gnd.n7273 gnd.n7271 585
R1887 gnd.n7271 gnd.n350 585
R1888 gnd.n7274 gnd.n359 585
R1889 gnd.n7290 gnd.n359 585
R1890 gnd.n7275 gnd.n7270 585
R1891 gnd.n7270 gnd.n7269 585
R1892 gnd.n374 gnd.n372 585
R1893 gnd.n7253 gnd.n372 585
R1894 gnd.n7280 gnd.n7279 585
R1895 gnd.n7281 gnd.n7280 585
R1896 gnd.n373 gnd.n371 585
R1897 gnd.n7259 gnd.n371 585
R1898 gnd.n7228 gnd.n7227 585
R1899 gnd.n7227 gnd.n7226 585
R1900 gnd.n7229 gnd.n392 585
R1901 gnd.n7245 gnd.n392 585
R1902 gnd.n406 gnd.n404 585
R1903 gnd.n6004 gnd.n404 585
R1904 gnd.n7234 gnd.n7233 585
R1905 gnd.n7235 gnd.n7234 585
R1906 gnd.n405 gnd.n403 585
R1907 gnd.n5999 gnd.n403 585
R1908 gnd.n6053 gnd.n6051 585
R1909 gnd.n6051 gnd.n6050 585
R1910 gnd.n6054 gnd.n1360 585
R1911 gnd.n1373 gnd.n1360 585
R1912 gnd.n6055 gnd.n1359 585
R1913 gnd.n6042 gnd.n1359 585
R1914 gnd.n6019 gnd.n1357 585
R1915 gnd.n6020 gnd.n6019 585
R1916 gnd.n6059 gnd.n1356 585
R1917 gnd.n1398 gnd.n1356 585
R1918 gnd.n6060 gnd.n1355 585
R1919 gnd.n5982 gnd.n1355 585
R1920 gnd.n6061 gnd.n1354 585
R1921 gnd.n1407 gnd.n1354 585
R1922 gnd.n5971 gnd.n1352 585
R1923 gnd.n5972 gnd.n5971 585
R1924 gnd.n6065 gnd.n1351 585
R1925 gnd.n5959 gnd.n1351 585
R1926 gnd.n6066 gnd.n1350 585
R1927 gnd.n1414 gnd.n1350 585
R1928 gnd.n6067 gnd.n1349 585
R1929 gnd.n5945 gnd.n1349 585
R1930 gnd.n1434 gnd.n1347 585
R1931 gnd.n1435 gnd.n1434 585
R1932 gnd.n6071 gnd.n1346 585
R1933 gnd.n5935 gnd.n1346 585
R1934 gnd.n6072 gnd.n1345 585
R1935 gnd.n5923 gnd.n1345 585
R1936 gnd.n6073 gnd.n1344 585
R1937 gnd.n1452 gnd.n1344 585
R1938 gnd.n1341 gnd.n1340 585
R1939 gnd.n5914 gnd.n1340 585
R1940 gnd.n6078 gnd.n6077 585
R1941 gnd.n6079 gnd.n6078 585
R1942 gnd.n1517 gnd.n1339 585
R1943 gnd.n1522 gnd.n1521 585
R1944 gnd.n1524 gnd.n1523 585
R1945 gnd.n1527 gnd.n1526 585
R1946 gnd.n1525 gnd.n1510 585
R1947 gnd.n1541 gnd.n1540 585
R1948 gnd.n1543 gnd.n1542 585
R1949 gnd.n1546 gnd.n1545 585
R1950 gnd.n1544 gnd.n1503 585
R1951 gnd.n1560 gnd.n1559 585
R1952 gnd.n1562 gnd.n1561 585
R1953 gnd.n1565 gnd.n1564 585
R1954 gnd.n1563 gnd.n1496 585
R1955 gnd.n1578 gnd.n1577 585
R1956 gnd.n1580 gnd.n1579 585
R1957 gnd.n1489 gnd.n1488 585
R1958 gnd.n1593 gnd.n1490 585
R1959 gnd.n1594 gnd.n1485 585
R1960 gnd.n1595 gnd.n1284 585
R1961 gnd.n6155 gnd.n1284 585
R1962 gnd.n7668 gnd.n7667 585
R1963 gnd.n7540 gnd.n124 585
R1964 gnd.n7542 gnd.n7541 585
R1965 gnd.n7538 gnd.n7537 585
R1966 gnd.n7546 gnd.n7536 585
R1967 gnd.n7547 gnd.n7534 585
R1968 gnd.n7548 gnd.n7533 585
R1969 gnd.n7531 gnd.n7529 585
R1970 gnd.n7552 gnd.n7528 585
R1971 gnd.n7553 gnd.n7526 585
R1972 gnd.n7554 gnd.n7525 585
R1973 gnd.n7523 gnd.n7521 585
R1974 gnd.n7558 gnd.n7520 585
R1975 gnd.n7559 gnd.n7518 585
R1976 gnd.n7560 gnd.n7517 585
R1977 gnd.n7515 gnd.n7513 585
R1978 gnd.n7564 gnd.n7512 585
R1979 gnd.n7565 gnd.n7510 585
R1980 gnd.n7566 gnd.n7509 585
R1981 gnd.n7509 gnd.n128 585
R1982 gnd.n7666 gnd.n120 585
R1983 gnd.n7666 gnd.n7665 585
R1984 gnd.n7672 gnd.n119 585
R1985 gnd.n126 gnd.n119 585
R1986 gnd.n7673 gnd.n118 585
R1987 gnd.n7585 gnd.n118 585
R1988 gnd.n7674 gnd.n117 585
R1989 gnd.n206 gnd.n117 585
R1990 gnd.n215 gnd.n115 585
R1991 gnd.n7577 gnd.n215 585
R1992 gnd.n7678 gnd.n114 585
R1993 gnd.n213 gnd.n114 585
R1994 gnd.n7679 gnd.n113 585
R1995 gnd.n7501 gnd.n113 585
R1996 gnd.n7680 gnd.n112 585
R1997 gnd.n232 gnd.n112 585
R1998 gnd.n231 gnd.n110 585
R1999 gnd.n7493 gnd.n231 585
R2000 gnd.n7684 gnd.n109 585
R2001 gnd.n229 gnd.n109 585
R2002 gnd.n7685 gnd.n108 585
R2003 gnd.n7485 gnd.n108 585
R2004 gnd.n7686 gnd.n107 585
R2005 gnd.n247 gnd.n107 585
R2006 gnd.n246 gnd.n105 585
R2007 gnd.n7477 gnd.n246 585
R2008 gnd.n7690 gnd.n104 585
R2009 gnd.n254 gnd.n104 585
R2010 gnd.n7691 gnd.n103 585
R2011 gnd.n7469 gnd.n103 585
R2012 gnd.n7692 gnd.n102 585
R2013 gnd.n263 gnd.n102 585
R2014 gnd.n262 gnd.n100 585
R2015 gnd.n7461 gnd.n262 585
R2016 gnd.n7696 gnd.n99 585
R2017 gnd.n260 gnd.n99 585
R2018 gnd.n7697 gnd.n98 585
R2019 gnd.n7453 gnd.n98 585
R2020 gnd.n7698 gnd.n97 585
R2021 gnd.n269 gnd.n97 585
R2022 gnd.n277 gnd.n95 585
R2023 gnd.n7445 gnd.n277 585
R2024 gnd.n7702 gnd.n94 585
R2025 gnd.n284 gnd.n94 585
R2026 gnd.n7703 gnd.n93 585
R2027 gnd.n7437 gnd.n93 585
R2028 gnd.n7704 gnd.n92 585
R2029 gnd.n293 gnd.n92 585
R2030 gnd.n292 gnd.n90 585
R2031 gnd.n7429 gnd.n292 585
R2032 gnd.n7708 gnd.n89 585
R2033 gnd.n290 gnd.n89 585
R2034 gnd.n7709 gnd.n88 585
R2035 gnd.n7421 gnd.n88 585
R2036 gnd.n7710 gnd.n87 585
R2037 gnd.n299 gnd.n87 585
R2038 gnd.n329 gnd.n85 585
R2039 gnd.n7397 gnd.n329 585
R2040 gnd.n7714 gnd.n84 585
R2041 gnd.n7393 gnd.n84 585
R2042 gnd.n7715 gnd.n83 585
R2043 gnd.n334 gnd.n83 585
R2044 gnd.n7716 gnd.n82 585
R2045 gnd.n7320 gnd.n82 585
R2046 gnd.n345 gnd.n80 585
R2047 gnd.n345 gnd.n340 585
R2048 gnd.n7313 gnd.n7312 585
R2049 gnd.n7314 gnd.n7313 585
R2050 gnd.n7311 gnd.n344 585
R2051 gnd.n344 gnd.n315 585
R2052 gnd.n346 gnd.n314 585
R2053 gnd.n7412 gnd.n314 585
R2054 gnd.n7307 gnd.n7306 585
R2055 gnd.n7306 gnd.n7305 585
R2056 gnd.n349 gnd.n348 585
R2057 gnd.n350 gnd.n349 585
R2058 gnd.n380 gnd.n357 585
R2059 gnd.n7290 gnd.n357 585
R2060 gnd.n7268 gnd.n7267 585
R2061 gnd.n7269 gnd.n7268 585
R2062 gnd.n379 gnd.n378 585
R2063 gnd.n7253 gnd.n378 585
R2064 gnd.n7262 gnd.n369 585
R2065 gnd.n7281 gnd.n369 585
R2066 gnd.n7261 gnd.n7260 585
R2067 gnd.n7260 gnd.n7259 585
R2068 gnd.n383 gnd.n382 585
R2069 gnd.n7226 gnd.n383 585
R2070 gnd.n6006 gnd.n391 585
R2071 gnd.n7245 gnd.n391 585
R2072 gnd.n6007 gnd.n6005 585
R2073 gnd.n6005 gnd.n6004 585
R2074 gnd.n6001 gnd.n401 585
R2075 gnd.n7235 gnd.n401 585
R2076 gnd.n6011 gnd.n6000 585
R2077 gnd.n6000 gnd.n5999 585
R2078 gnd.n6012 gnd.n1363 585
R2079 gnd.n6050 gnd.n1363 585
R2080 gnd.n6013 gnd.n1386 585
R2081 gnd.n1386 gnd.n1373 585
R2082 gnd.n1383 gnd.n1372 585
R2083 gnd.n6042 gnd.n1372 585
R2084 gnd.n6018 gnd.n6017 585
R2085 gnd.n6020 gnd.n6018 585
R2086 gnd.n1382 gnd.n1381 585
R2087 gnd.n1398 gnd.n1381 585
R2088 gnd.n5952 gnd.n1395 585
R2089 gnd.n5982 gnd.n1395 585
R2090 gnd.n5953 gnd.n5951 585
R2091 gnd.n5951 gnd.n1407 585
R2092 gnd.n1418 gnd.n1406 585
R2093 gnd.n5972 gnd.n1406 585
R2094 gnd.n5958 gnd.n5957 585
R2095 gnd.n5959 gnd.n5958 585
R2096 gnd.n1417 gnd.n1416 585
R2097 gnd.n1416 gnd.n1414 585
R2098 gnd.n5947 gnd.n5946 585
R2099 gnd.n5946 gnd.n5945 585
R2100 gnd.n1421 gnd.n1420 585
R2101 gnd.n1435 gnd.n1421 585
R2102 gnd.n1477 gnd.n1433 585
R2103 gnd.n5935 gnd.n1433 585
R2104 gnd.n5922 gnd.n5921 585
R2105 gnd.n5923 gnd.n5922 585
R2106 gnd.n1476 gnd.n1475 585
R2107 gnd.n1475 gnd.n1452 585
R2108 gnd.n5916 gnd.n5915 585
R2109 gnd.n5915 gnd.n5914 585
R2110 gnd.n5904 gnd.n1337 585
R2111 gnd.n6079 gnd.n1337 585
R2112 gnd.n3720 gnd.n3719 585
R2113 gnd.n3721 gnd.n3720 585
R2114 gnd.n2415 gnd.n2414 585
R2115 gnd.n2421 gnd.n2414 585
R2116 gnd.n3695 gnd.n2433 585
R2117 gnd.n2433 gnd.n2420 585
R2118 gnd.n3697 gnd.n3696 585
R2119 gnd.n3698 gnd.n3697 585
R2120 gnd.n2434 gnd.n2432 585
R2121 gnd.n2432 gnd.n2428 585
R2122 gnd.n3429 gnd.n3428 585
R2123 gnd.n3428 gnd.n3427 585
R2124 gnd.n2439 gnd.n2438 585
R2125 gnd.n3398 gnd.n2439 585
R2126 gnd.n3418 gnd.n3417 585
R2127 gnd.n3417 gnd.n3416 585
R2128 gnd.n2446 gnd.n2445 585
R2129 gnd.n3404 gnd.n2446 585
R2130 gnd.n3374 gnd.n2466 585
R2131 gnd.n2466 gnd.n2465 585
R2132 gnd.n3376 gnd.n3375 585
R2133 gnd.n3377 gnd.n3376 585
R2134 gnd.n2467 gnd.n2464 585
R2135 gnd.n2475 gnd.n2464 585
R2136 gnd.n3352 gnd.n2487 585
R2137 gnd.n2487 gnd.n2474 585
R2138 gnd.n3354 gnd.n3353 585
R2139 gnd.n3355 gnd.n3354 585
R2140 gnd.n2488 gnd.n2486 585
R2141 gnd.n2486 gnd.n2482 585
R2142 gnd.n3340 gnd.n3339 585
R2143 gnd.n3339 gnd.n3338 585
R2144 gnd.n2493 gnd.n2492 585
R2145 gnd.n2503 gnd.n2493 585
R2146 gnd.n3329 gnd.n3328 585
R2147 gnd.n3328 gnd.n3327 585
R2148 gnd.n2500 gnd.n2499 585
R2149 gnd.n3315 gnd.n2500 585
R2150 gnd.n3289 gnd.n2521 585
R2151 gnd.n2521 gnd.n2510 585
R2152 gnd.n3291 gnd.n3290 585
R2153 gnd.n3292 gnd.n3291 585
R2154 gnd.n2522 gnd.n2520 585
R2155 gnd.n2530 gnd.n2520 585
R2156 gnd.n3267 gnd.n2542 585
R2157 gnd.n2542 gnd.n2529 585
R2158 gnd.n3269 gnd.n3268 585
R2159 gnd.n3270 gnd.n3269 585
R2160 gnd.n2543 gnd.n2541 585
R2161 gnd.n2541 gnd.n2537 585
R2162 gnd.n3255 gnd.n3254 585
R2163 gnd.n3254 gnd.n3253 585
R2164 gnd.n2548 gnd.n2547 585
R2165 gnd.n2557 gnd.n2548 585
R2166 gnd.n3244 gnd.n3243 585
R2167 gnd.n3243 gnd.n3242 585
R2168 gnd.n2555 gnd.n2554 585
R2169 gnd.n3230 gnd.n2555 585
R2170 gnd.n2668 gnd.n2667 585
R2171 gnd.n2668 gnd.n2564 585
R2172 gnd.n3187 gnd.n3186 585
R2173 gnd.n3186 gnd.n3185 585
R2174 gnd.n3188 gnd.n2662 585
R2175 gnd.n2673 gnd.n2662 585
R2176 gnd.n3190 gnd.n3189 585
R2177 gnd.n3191 gnd.n3190 585
R2178 gnd.n2663 gnd.n2661 585
R2179 gnd.n2686 gnd.n2661 585
R2180 gnd.n2646 gnd.n2645 585
R2181 gnd.n2649 gnd.n2646 585
R2182 gnd.n3201 gnd.n3200 585
R2183 gnd.n3200 gnd.n3199 585
R2184 gnd.n3202 gnd.n2640 585
R2185 gnd.n3161 gnd.n2640 585
R2186 gnd.n3204 gnd.n3203 585
R2187 gnd.n3205 gnd.n3204 585
R2188 gnd.n2641 gnd.n2639 585
R2189 gnd.n2700 gnd.n2639 585
R2190 gnd.n3153 gnd.n3152 585
R2191 gnd.n3152 gnd.n3151 585
R2192 gnd.n2697 gnd.n2696 585
R2193 gnd.n3135 gnd.n2697 585
R2194 gnd.n3122 gnd.n2716 585
R2195 gnd.n2716 gnd.n2715 585
R2196 gnd.n3124 gnd.n3123 585
R2197 gnd.n3125 gnd.n3124 585
R2198 gnd.n2717 gnd.n2714 585
R2199 gnd.n2723 gnd.n2714 585
R2200 gnd.n3103 gnd.n3102 585
R2201 gnd.n3104 gnd.n3103 585
R2202 gnd.n2734 gnd.n2733 585
R2203 gnd.n2733 gnd.n2729 585
R2204 gnd.n3093 gnd.n3092 585
R2205 gnd.n3094 gnd.n3093 585
R2206 gnd.n2744 gnd.n2743 585
R2207 gnd.n2749 gnd.n2743 585
R2208 gnd.n3071 gnd.n2762 585
R2209 gnd.n2762 gnd.n2748 585
R2210 gnd.n3073 gnd.n3072 585
R2211 gnd.n3074 gnd.n3073 585
R2212 gnd.n2763 gnd.n2761 585
R2213 gnd.n2761 gnd.n2757 585
R2214 gnd.n3062 gnd.n3061 585
R2215 gnd.n3063 gnd.n3062 585
R2216 gnd.n2770 gnd.n2769 585
R2217 gnd.n2774 gnd.n2769 585
R2218 gnd.n3039 gnd.n2791 585
R2219 gnd.n2791 gnd.n2773 585
R2220 gnd.n3041 gnd.n3040 585
R2221 gnd.n3042 gnd.n3041 585
R2222 gnd.n2792 gnd.n2790 585
R2223 gnd.n2790 gnd.n2781 585
R2224 gnd.n3034 gnd.n3033 585
R2225 gnd.n3033 gnd.n3032 585
R2226 gnd.n2839 gnd.n2838 585
R2227 gnd.n2840 gnd.n2839 585
R2228 gnd.n2993 gnd.n2992 585
R2229 gnd.n2994 gnd.n2993 585
R2230 gnd.n2849 gnd.n2848 585
R2231 gnd.n2848 gnd.n2847 585
R2232 gnd.n2988 gnd.n2987 585
R2233 gnd.n2987 gnd.n2986 585
R2234 gnd.n2852 gnd.n2851 585
R2235 gnd.n2853 gnd.n2852 585
R2236 gnd.n2977 gnd.n2976 585
R2237 gnd.n2978 gnd.n2977 585
R2238 gnd.n2860 gnd.n2859 585
R2239 gnd.n2969 gnd.n2859 585
R2240 gnd.n2972 gnd.n2971 585
R2241 gnd.n2971 gnd.n2970 585
R2242 gnd.n2863 gnd.n2862 585
R2243 gnd.n2864 gnd.n2863 585
R2244 gnd.n2958 gnd.n2957 585
R2245 gnd.n2956 gnd.n2882 585
R2246 gnd.n2955 gnd.n2881 585
R2247 gnd.n2960 gnd.n2881 585
R2248 gnd.n2954 gnd.n2953 585
R2249 gnd.n2952 gnd.n2951 585
R2250 gnd.n2950 gnd.n2949 585
R2251 gnd.n2948 gnd.n2947 585
R2252 gnd.n2946 gnd.n2945 585
R2253 gnd.n2944 gnd.n2943 585
R2254 gnd.n2942 gnd.n2941 585
R2255 gnd.n2940 gnd.n2939 585
R2256 gnd.n2938 gnd.n2937 585
R2257 gnd.n2936 gnd.n2935 585
R2258 gnd.n2934 gnd.n2933 585
R2259 gnd.n2932 gnd.n2931 585
R2260 gnd.n2930 gnd.n2929 585
R2261 gnd.n2928 gnd.n2927 585
R2262 gnd.n2926 gnd.n2925 585
R2263 gnd.n2924 gnd.n2923 585
R2264 gnd.n2922 gnd.n2921 585
R2265 gnd.n2920 gnd.n2919 585
R2266 gnd.n2918 gnd.n2917 585
R2267 gnd.n2916 gnd.n2915 585
R2268 gnd.n2914 gnd.n2913 585
R2269 gnd.n2912 gnd.n2911 585
R2270 gnd.n2869 gnd.n2868 585
R2271 gnd.n2963 gnd.n2962 585
R2272 gnd.n3724 gnd.n3723 585
R2273 gnd.n3726 gnd.n3725 585
R2274 gnd.n3728 gnd.n3727 585
R2275 gnd.n3730 gnd.n3729 585
R2276 gnd.n3732 gnd.n3731 585
R2277 gnd.n3734 gnd.n3733 585
R2278 gnd.n3736 gnd.n3735 585
R2279 gnd.n3738 gnd.n3737 585
R2280 gnd.n3740 gnd.n3739 585
R2281 gnd.n3742 gnd.n3741 585
R2282 gnd.n3744 gnd.n3743 585
R2283 gnd.n3746 gnd.n3745 585
R2284 gnd.n3748 gnd.n3747 585
R2285 gnd.n3750 gnd.n3749 585
R2286 gnd.n3752 gnd.n3751 585
R2287 gnd.n3754 gnd.n3753 585
R2288 gnd.n3756 gnd.n3755 585
R2289 gnd.n3758 gnd.n3757 585
R2290 gnd.n3760 gnd.n3759 585
R2291 gnd.n3762 gnd.n3761 585
R2292 gnd.n3764 gnd.n3763 585
R2293 gnd.n3766 gnd.n3765 585
R2294 gnd.n3768 gnd.n3767 585
R2295 gnd.n3770 gnd.n3769 585
R2296 gnd.n3772 gnd.n3771 585
R2297 gnd.n3773 gnd.n2381 585
R2298 gnd.n3774 gnd.n2339 585
R2299 gnd.n3812 gnd.n2339 585
R2300 gnd.n3722 gnd.n2411 585
R2301 gnd.n3722 gnd.n3721 585
R2302 gnd.n3391 gnd.n2410 585
R2303 gnd.n2421 gnd.n2410 585
R2304 gnd.n3393 gnd.n3392 585
R2305 gnd.n3392 gnd.n2420 585
R2306 gnd.n3394 gnd.n2430 585
R2307 gnd.n3698 gnd.n2430 585
R2308 gnd.n3396 gnd.n3395 585
R2309 gnd.n3395 gnd.n2428 585
R2310 gnd.n3397 gnd.n2441 585
R2311 gnd.n3427 gnd.n2441 585
R2312 gnd.n3400 gnd.n3399 585
R2313 gnd.n3399 gnd.n3398 585
R2314 gnd.n3401 gnd.n2448 585
R2315 gnd.n3416 gnd.n2448 585
R2316 gnd.n3403 gnd.n3402 585
R2317 gnd.n3404 gnd.n3403 585
R2318 gnd.n2458 gnd.n2457 585
R2319 gnd.n2465 gnd.n2457 585
R2320 gnd.n3379 gnd.n3378 585
R2321 gnd.n3378 gnd.n3377 585
R2322 gnd.n2461 gnd.n2460 585
R2323 gnd.n2475 gnd.n2461 585
R2324 gnd.n3305 gnd.n3304 585
R2325 gnd.n3304 gnd.n2474 585
R2326 gnd.n3306 gnd.n2484 585
R2327 gnd.n3355 gnd.n2484 585
R2328 gnd.n3308 gnd.n3307 585
R2329 gnd.n3307 gnd.n2482 585
R2330 gnd.n3309 gnd.n2495 585
R2331 gnd.n3338 gnd.n2495 585
R2332 gnd.n3311 gnd.n3310 585
R2333 gnd.n3310 gnd.n2503 585
R2334 gnd.n3312 gnd.n2502 585
R2335 gnd.n3327 gnd.n2502 585
R2336 gnd.n3314 gnd.n3313 585
R2337 gnd.n3315 gnd.n3314 585
R2338 gnd.n2514 gnd.n2513 585
R2339 gnd.n2513 gnd.n2510 585
R2340 gnd.n3294 gnd.n3293 585
R2341 gnd.n3293 gnd.n3292 585
R2342 gnd.n2517 gnd.n2516 585
R2343 gnd.n2530 gnd.n2517 585
R2344 gnd.n3218 gnd.n3217 585
R2345 gnd.n3217 gnd.n2529 585
R2346 gnd.n3219 gnd.n2539 585
R2347 gnd.n3270 gnd.n2539 585
R2348 gnd.n3221 gnd.n3220 585
R2349 gnd.n3220 gnd.n2537 585
R2350 gnd.n3222 gnd.n2550 585
R2351 gnd.n3253 gnd.n2550 585
R2352 gnd.n3224 gnd.n3223 585
R2353 gnd.n3223 gnd.n2557 585
R2354 gnd.n3225 gnd.n2556 585
R2355 gnd.n3242 gnd.n2556 585
R2356 gnd.n3227 gnd.n3226 585
R2357 gnd.n3230 gnd.n3227 585
R2358 gnd.n2567 gnd.n2566 585
R2359 gnd.n2566 gnd.n2564 585
R2360 gnd.n2670 gnd.n2669 585
R2361 gnd.n3185 gnd.n2669 585
R2362 gnd.n2672 gnd.n2671 585
R2363 gnd.n2673 gnd.n2672 585
R2364 gnd.n2683 gnd.n2659 585
R2365 gnd.n3191 gnd.n2659 585
R2366 gnd.n2685 gnd.n2684 585
R2367 gnd.n2686 gnd.n2685 585
R2368 gnd.n2682 gnd.n2681 585
R2369 gnd.n2682 gnd.n2649 585
R2370 gnd.n2680 gnd.n2647 585
R2371 gnd.n3199 gnd.n2647 585
R2372 gnd.n2636 gnd.n2634 585
R2373 gnd.n3161 gnd.n2636 585
R2374 gnd.n3207 gnd.n3206 585
R2375 gnd.n3206 gnd.n3205 585
R2376 gnd.n2635 gnd.n2633 585
R2377 gnd.n2700 gnd.n2635 585
R2378 gnd.n3132 gnd.n2699 585
R2379 gnd.n3151 gnd.n2699 585
R2380 gnd.n3134 gnd.n3133 585
R2381 gnd.n3135 gnd.n3134 585
R2382 gnd.n2709 gnd.n2708 585
R2383 gnd.n2715 gnd.n2708 585
R2384 gnd.n3127 gnd.n3126 585
R2385 gnd.n3126 gnd.n3125 585
R2386 gnd.n2712 gnd.n2711 585
R2387 gnd.n2723 gnd.n2712 585
R2388 gnd.n3012 gnd.n2731 585
R2389 gnd.n3104 gnd.n2731 585
R2390 gnd.n3014 gnd.n3013 585
R2391 gnd.n3013 gnd.n2729 585
R2392 gnd.n3015 gnd.n2742 585
R2393 gnd.n3094 gnd.n2742 585
R2394 gnd.n3017 gnd.n3016 585
R2395 gnd.n3017 gnd.n2749 585
R2396 gnd.n3019 gnd.n3018 585
R2397 gnd.n3018 gnd.n2748 585
R2398 gnd.n3020 gnd.n2759 585
R2399 gnd.n3074 gnd.n2759 585
R2400 gnd.n3022 gnd.n3021 585
R2401 gnd.n3021 gnd.n2757 585
R2402 gnd.n3023 gnd.n2768 585
R2403 gnd.n3063 gnd.n2768 585
R2404 gnd.n3025 gnd.n3024 585
R2405 gnd.n3025 gnd.n2774 585
R2406 gnd.n3027 gnd.n3026 585
R2407 gnd.n3026 gnd.n2773 585
R2408 gnd.n3028 gnd.n2789 585
R2409 gnd.n3042 gnd.n2789 585
R2410 gnd.n3029 gnd.n2842 585
R2411 gnd.n2842 gnd.n2781 585
R2412 gnd.n3031 gnd.n3030 585
R2413 gnd.n3032 gnd.n3031 585
R2414 gnd.n2843 gnd.n2841 585
R2415 gnd.n2841 gnd.n2840 585
R2416 gnd.n2996 gnd.n2995 585
R2417 gnd.n2995 gnd.n2994 585
R2418 gnd.n2846 gnd.n2845 585
R2419 gnd.n2847 gnd.n2846 585
R2420 gnd.n2985 gnd.n2984 585
R2421 gnd.n2986 gnd.n2985 585
R2422 gnd.n2855 gnd.n2854 585
R2423 gnd.n2854 gnd.n2853 585
R2424 gnd.n2980 gnd.n2979 585
R2425 gnd.n2979 gnd.n2978 585
R2426 gnd.n2858 gnd.n2857 585
R2427 gnd.n2969 gnd.n2858 585
R2428 gnd.n2968 gnd.n2967 585
R2429 gnd.n2970 gnd.n2968 585
R2430 gnd.n2866 gnd.n2865 585
R2431 gnd.n2865 gnd.n2864 585
R2432 gnd.n3707 gnd.n2361 585
R2433 gnd.n2413 gnd.n2361 585
R2434 gnd.n3708 gnd.n2423 585
R2435 gnd.n2423 gnd.n2412 585
R2436 gnd.n3710 gnd.n3709 585
R2437 gnd.n3711 gnd.n3710 585
R2438 gnd.n2424 gnd.n2422 585
R2439 gnd.n2431 gnd.n2422 585
R2440 gnd.n3701 gnd.n3700 585
R2441 gnd.n3700 gnd.n3699 585
R2442 gnd.n2427 gnd.n2426 585
R2443 gnd.n3426 gnd.n2427 585
R2444 gnd.n3412 gnd.n2450 585
R2445 gnd.n2450 gnd.n2440 585
R2446 gnd.n3414 gnd.n3413 585
R2447 gnd.n3415 gnd.n3414 585
R2448 gnd.n2451 gnd.n2449 585
R2449 gnd.n2449 gnd.n2447 585
R2450 gnd.n3407 gnd.n3406 585
R2451 gnd.n3406 gnd.n3405 585
R2452 gnd.n2454 gnd.n2453 585
R2453 gnd.n2463 gnd.n2454 585
R2454 gnd.n3363 gnd.n2477 585
R2455 gnd.n2477 gnd.n2462 585
R2456 gnd.n3365 gnd.n3364 585
R2457 gnd.n3366 gnd.n3365 585
R2458 gnd.n2478 gnd.n2476 585
R2459 gnd.n2485 gnd.n2476 585
R2460 gnd.n3358 gnd.n3357 585
R2461 gnd.n3357 gnd.n3356 585
R2462 gnd.n2481 gnd.n2480 585
R2463 gnd.n3337 gnd.n2481 585
R2464 gnd.n3323 gnd.n2505 585
R2465 gnd.n2505 gnd.n2494 585
R2466 gnd.n3325 gnd.n3324 585
R2467 gnd.n3326 gnd.n3325 585
R2468 gnd.n2506 gnd.n2504 585
R2469 gnd.n2504 gnd.n2501 585
R2470 gnd.n3318 gnd.n3317 585
R2471 gnd.n3317 gnd.n3316 585
R2472 gnd.n2509 gnd.n2508 585
R2473 gnd.n2519 gnd.n2509 585
R2474 gnd.n3278 gnd.n2532 585
R2475 gnd.n2532 gnd.n2518 585
R2476 gnd.n3280 gnd.n3279 585
R2477 gnd.n3281 gnd.n3280 585
R2478 gnd.n2533 gnd.n2531 585
R2479 gnd.n2540 gnd.n2531 585
R2480 gnd.n3273 gnd.n3272 585
R2481 gnd.n3272 gnd.n3271 585
R2482 gnd.n2536 gnd.n2535 585
R2483 gnd.n3252 gnd.n2536 585
R2484 gnd.n3238 gnd.n2559 585
R2485 gnd.n2559 gnd.n2549 585
R2486 gnd.n3240 gnd.n3239 585
R2487 gnd.n3241 gnd.n3240 585
R2488 gnd.n2560 gnd.n2558 585
R2489 gnd.n3229 gnd.n2558 585
R2490 gnd.n3233 gnd.n3232 585
R2491 gnd.n3232 gnd.n3231 585
R2492 gnd.n2563 gnd.n2562 585
R2493 gnd.n3184 gnd.n2563 585
R2494 gnd.n2677 gnd.n2676 585
R2495 gnd.n2678 gnd.n2677 585
R2496 gnd.n2657 gnd.n2656 585
R2497 gnd.n2660 gnd.n2657 585
R2498 gnd.n3194 gnd.n3193 585
R2499 gnd.n3193 gnd.n3192 585
R2500 gnd.n3195 gnd.n2651 585
R2501 gnd.n2687 gnd.n2651 585
R2502 gnd.n3197 gnd.n3196 585
R2503 gnd.n3198 gnd.n3197 585
R2504 gnd.n2652 gnd.n2650 585
R2505 gnd.n3162 gnd.n2650 585
R2506 gnd.n3146 gnd.n3145 585
R2507 gnd.n3145 gnd.n2638 585
R2508 gnd.n3147 gnd.n2702 585
R2509 gnd.n2702 gnd.n2637 585
R2510 gnd.n3149 gnd.n3148 585
R2511 gnd.n3150 gnd.n3149 585
R2512 gnd.n2703 gnd.n2701 585
R2513 gnd.n2701 gnd.n2698 585
R2514 gnd.n3138 gnd.n3137 585
R2515 gnd.n3137 gnd.n3136 585
R2516 gnd.n2706 gnd.n2705 585
R2517 gnd.n2713 gnd.n2706 585
R2518 gnd.n3112 gnd.n3111 585
R2519 gnd.n3113 gnd.n3112 585
R2520 gnd.n2725 gnd.n2724 585
R2521 gnd.n2732 gnd.n2724 585
R2522 gnd.n3107 gnd.n3106 585
R2523 gnd.n3106 gnd.n3105 585
R2524 gnd.n2728 gnd.n2727 585
R2525 gnd.n3095 gnd.n2728 585
R2526 gnd.n3082 gnd.n2752 585
R2527 gnd.n2752 gnd.n2751 585
R2528 gnd.n3084 gnd.n3083 585
R2529 gnd.n3085 gnd.n3084 585
R2530 gnd.n2753 gnd.n2750 585
R2531 gnd.n2760 gnd.n2750 585
R2532 gnd.n3077 gnd.n3076 585
R2533 gnd.n3076 gnd.n3075 585
R2534 gnd.n2756 gnd.n2755 585
R2535 gnd.n3064 gnd.n2756 585
R2536 gnd.n3051 gnd.n2777 585
R2537 gnd.n2777 gnd.n2776 585
R2538 gnd.n3053 gnd.n3052 585
R2539 gnd.n3054 gnd.n3053 585
R2540 gnd.n3047 gnd.n2775 585
R2541 gnd.n3046 gnd.n3045 585
R2542 gnd.n2780 gnd.n2779 585
R2543 gnd.n3043 gnd.n2780 585
R2544 gnd.n2802 gnd.n2801 585
R2545 gnd.n2805 gnd.n2804 585
R2546 gnd.n2803 gnd.n2798 585
R2547 gnd.n2810 gnd.n2809 585
R2548 gnd.n2812 gnd.n2811 585
R2549 gnd.n2815 gnd.n2814 585
R2550 gnd.n2813 gnd.n2796 585
R2551 gnd.n2820 gnd.n2819 585
R2552 gnd.n2822 gnd.n2821 585
R2553 gnd.n2825 gnd.n2824 585
R2554 gnd.n2823 gnd.n2794 585
R2555 gnd.n2830 gnd.n2829 585
R2556 gnd.n2834 gnd.n2831 585
R2557 gnd.n2835 gnd.n2772 585
R2558 gnd.n3713 gnd.n2376 585
R2559 gnd.n3780 gnd.n3779 585
R2560 gnd.n3782 gnd.n3781 585
R2561 gnd.n3784 gnd.n3783 585
R2562 gnd.n3786 gnd.n3785 585
R2563 gnd.n3788 gnd.n3787 585
R2564 gnd.n3790 gnd.n3789 585
R2565 gnd.n3792 gnd.n3791 585
R2566 gnd.n3794 gnd.n3793 585
R2567 gnd.n3796 gnd.n3795 585
R2568 gnd.n3798 gnd.n3797 585
R2569 gnd.n3800 gnd.n3799 585
R2570 gnd.n3802 gnd.n3801 585
R2571 gnd.n3805 gnd.n3804 585
R2572 gnd.n3803 gnd.n2364 585
R2573 gnd.n3809 gnd.n2362 585
R2574 gnd.n3811 gnd.n3810 585
R2575 gnd.n3812 gnd.n3811 585
R2576 gnd.n3714 gnd.n2418 585
R2577 gnd.n3714 gnd.n2413 585
R2578 gnd.n3716 gnd.n3715 585
R2579 gnd.n3715 gnd.n2412 585
R2580 gnd.n3712 gnd.n2417 585
R2581 gnd.n3712 gnd.n3711 585
R2582 gnd.n3691 gnd.n2419 585
R2583 gnd.n2431 gnd.n2419 585
R2584 gnd.n3690 gnd.n2429 585
R2585 gnd.n3699 gnd.n2429 585
R2586 gnd.n3425 gnd.n2436 585
R2587 gnd.n3426 gnd.n3425 585
R2588 gnd.n3424 gnd.n3423 585
R2589 gnd.n3424 gnd.n2440 585
R2590 gnd.n3422 gnd.n2442 585
R2591 gnd.n3415 gnd.n2442 585
R2592 gnd.n2455 gnd.n2443 585
R2593 gnd.n2455 gnd.n2447 585
R2594 gnd.n3371 gnd.n2456 585
R2595 gnd.n3405 gnd.n2456 585
R2596 gnd.n3370 gnd.n3369 585
R2597 gnd.n3369 gnd.n2463 585
R2598 gnd.n3368 gnd.n2471 585
R2599 gnd.n3368 gnd.n2462 585
R2600 gnd.n3367 gnd.n2473 585
R2601 gnd.n3367 gnd.n3366 585
R2602 gnd.n3346 gnd.n2472 585
R2603 gnd.n2485 gnd.n2472 585
R2604 gnd.n3345 gnd.n2483 585
R2605 gnd.n3356 gnd.n2483 585
R2606 gnd.n3336 gnd.n2490 585
R2607 gnd.n3337 gnd.n3336 585
R2608 gnd.n3335 gnd.n3334 585
R2609 gnd.n3335 gnd.n2494 585
R2610 gnd.n3333 gnd.n2496 585
R2611 gnd.n3326 gnd.n2496 585
R2612 gnd.n2511 gnd.n2497 585
R2613 gnd.n2511 gnd.n2501 585
R2614 gnd.n3286 gnd.n2512 585
R2615 gnd.n3316 gnd.n2512 585
R2616 gnd.n3285 gnd.n3284 585
R2617 gnd.n3284 gnd.n2519 585
R2618 gnd.n3283 gnd.n2526 585
R2619 gnd.n3283 gnd.n2518 585
R2620 gnd.n3282 gnd.n2528 585
R2621 gnd.n3282 gnd.n3281 585
R2622 gnd.n3261 gnd.n2527 585
R2623 gnd.n2540 gnd.n2527 585
R2624 gnd.n3260 gnd.n2538 585
R2625 gnd.n3271 gnd.n2538 585
R2626 gnd.n3251 gnd.n2545 585
R2627 gnd.n3252 gnd.n3251 585
R2628 gnd.n3250 gnd.n3249 585
R2629 gnd.n3250 gnd.n2549 585
R2630 gnd.n3248 gnd.n2551 585
R2631 gnd.n3241 gnd.n2551 585
R2632 gnd.n3228 gnd.n2552 585
R2633 gnd.n3229 gnd.n3228 585
R2634 gnd.n3181 gnd.n2565 585
R2635 gnd.n3231 gnd.n2565 585
R2636 gnd.n3183 gnd.n3182 585
R2637 gnd.n3184 gnd.n3183 585
R2638 gnd.n3176 gnd.n2679 585
R2639 gnd.n2679 gnd.n2678 585
R2640 gnd.n3174 gnd.n3173 585
R2641 gnd.n3173 gnd.n2660 585
R2642 gnd.n3171 gnd.n2658 585
R2643 gnd.n3192 gnd.n2658 585
R2644 gnd.n2689 gnd.n2688 585
R2645 gnd.n2688 gnd.n2687 585
R2646 gnd.n3165 gnd.n2648 585
R2647 gnd.n3198 gnd.n2648 585
R2648 gnd.n3164 gnd.n3163 585
R2649 gnd.n3163 gnd.n3162 585
R2650 gnd.n3160 gnd.n2691 585
R2651 gnd.n3160 gnd.n2638 585
R2652 gnd.n3159 gnd.n3158 585
R2653 gnd.n3159 gnd.n2637 585
R2654 gnd.n2694 gnd.n2693 585
R2655 gnd.n3150 gnd.n2693 585
R2656 gnd.n3118 gnd.n3117 585
R2657 gnd.n3117 gnd.n2698 585
R2658 gnd.n3119 gnd.n2707 585
R2659 gnd.n3136 gnd.n2707 585
R2660 gnd.n3116 gnd.n3115 585
R2661 gnd.n3115 gnd.n2713 585
R2662 gnd.n3114 gnd.n2721 585
R2663 gnd.n3114 gnd.n3113 585
R2664 gnd.n3099 gnd.n2722 585
R2665 gnd.n2732 gnd.n2722 585
R2666 gnd.n3098 gnd.n2730 585
R2667 gnd.n3105 gnd.n2730 585
R2668 gnd.n3097 gnd.n3096 585
R2669 gnd.n3096 gnd.n3095 585
R2670 gnd.n2741 gnd.n2738 585
R2671 gnd.n2751 gnd.n2741 585
R2672 gnd.n3087 gnd.n3086 585
R2673 gnd.n3086 gnd.n3085 585
R2674 gnd.n2747 gnd.n2746 585
R2675 gnd.n2760 gnd.n2747 585
R2676 gnd.n3067 gnd.n2758 585
R2677 gnd.n3075 gnd.n2758 585
R2678 gnd.n3066 gnd.n3065 585
R2679 gnd.n3065 gnd.n3064 585
R2680 gnd.n2767 gnd.n2765 585
R2681 gnd.n2776 gnd.n2767 585
R2682 gnd.n3056 gnd.n3055 585
R2683 gnd.n3055 gnd.n3054 585
R2684 gnd.n6326 gnd.n6325 585
R2685 gnd.n6325 gnd.n6324 585
R2686 gnd.n6327 gnd.n1103 585
R2687 gnd.n4568 gnd.n1103 585
R2688 gnd.n6329 gnd.n6328 585
R2689 gnd.n6330 gnd.n6329 585
R2690 gnd.n1088 gnd.n1087 585
R2691 gnd.n4530 gnd.n1088 585
R2692 gnd.n6338 gnd.n6337 585
R2693 gnd.n6337 gnd.n6336 585
R2694 gnd.n6339 gnd.n1082 585
R2695 gnd.n4521 gnd.n1082 585
R2696 gnd.n6341 gnd.n6340 585
R2697 gnd.n6342 gnd.n6341 585
R2698 gnd.n1067 gnd.n1066 585
R2699 gnd.n4513 gnd.n1067 585
R2700 gnd.n6350 gnd.n6349 585
R2701 gnd.n6349 gnd.n6348 585
R2702 gnd.n6351 gnd.n1061 585
R2703 gnd.n4451 gnd.n1061 585
R2704 gnd.n6353 gnd.n6352 585
R2705 gnd.n6354 gnd.n6353 585
R2706 gnd.n1046 gnd.n1045 585
R2707 gnd.n4439 gnd.n1046 585
R2708 gnd.n6362 gnd.n6361 585
R2709 gnd.n6361 gnd.n6360 585
R2710 gnd.n6363 gnd.n1040 585
R2711 gnd.n4462 gnd.n1040 585
R2712 gnd.n6365 gnd.n6364 585
R2713 gnd.n6366 gnd.n6365 585
R2714 gnd.n1025 gnd.n1024 585
R2715 gnd.n4431 gnd.n1025 585
R2716 gnd.n6374 gnd.n6373 585
R2717 gnd.n6373 gnd.n6372 585
R2718 gnd.n6375 gnd.n1019 585
R2719 gnd.n4398 gnd.n1019 585
R2720 gnd.n6377 gnd.n6376 585
R2721 gnd.n6378 gnd.n6377 585
R2722 gnd.n1004 gnd.n1003 585
R2723 gnd.n4390 gnd.n1004 585
R2724 gnd.n6386 gnd.n6385 585
R2725 gnd.n6385 gnd.n6384 585
R2726 gnd.n6387 gnd.n998 585
R2727 gnd.n4413 gnd.n998 585
R2728 gnd.n6389 gnd.n6388 585
R2729 gnd.n6390 gnd.n6389 585
R2730 gnd.n982 gnd.n981 585
R2731 gnd.n4382 gnd.n982 585
R2732 gnd.n6398 gnd.n6397 585
R2733 gnd.n6397 gnd.n6396 585
R2734 gnd.n6399 gnd.n976 585
R2735 gnd.n4364 gnd.n976 585
R2736 gnd.n6401 gnd.n6400 585
R2737 gnd.n6402 gnd.n6401 585
R2738 gnd.n977 gnd.n975 585
R2739 gnd.n975 gnd.n970 585
R2740 gnd.n4354 gnd.n4353 585
R2741 gnd.n4355 gnd.n4354 585
R2742 gnd.n4351 gnd.n2192 585
R2743 gnd.n2198 gnd.n2192 585
R2744 gnd.n4350 gnd.n4349 585
R2745 gnd.n4349 gnd.n4348 585
R2746 gnd.n4326 gnd.n2194 585
R2747 gnd.n2216 gnd.n2194 585
R2748 gnd.n4328 gnd.n4327 585
R2749 gnd.n4329 gnd.n4328 585
R2750 gnd.n4324 gnd.n2218 585
R2751 gnd.n2218 gnd.n2214 585
R2752 gnd.n4323 gnd.n4322 585
R2753 gnd.n4322 gnd.n4321 585
R2754 gnd.n4309 gnd.n2220 585
R2755 gnd.n2221 gnd.n2220 585
R2756 gnd.n4311 gnd.n4310 585
R2757 gnd.n4312 gnd.n4311 585
R2758 gnd.n4307 gnd.n2233 585
R2759 gnd.n2233 gnd.n2230 585
R2760 gnd.n4306 gnd.n4305 585
R2761 gnd.n4305 gnd.n4304 585
R2762 gnd.n2236 gnd.n2234 585
R2763 gnd.n2247 gnd.n2236 585
R2764 gnd.n4295 gnd.n4294 585
R2765 gnd.n4296 gnd.n4295 585
R2766 gnd.n2249 gnd.n2248 585
R2767 gnd.n2248 gnd.n2244 585
R2768 gnd.n4289 gnd.n4288 585
R2769 gnd.n4288 gnd.n4287 585
R2770 gnd.n2252 gnd.n2251 585
R2771 gnd.n2253 gnd.n2252 585
R2772 gnd.n4278 gnd.n4277 585
R2773 gnd.n4279 gnd.n4278 585
R2774 gnd.n2265 gnd.n2264 585
R2775 gnd.n2264 gnd.n2261 585
R2776 gnd.n4273 gnd.n4272 585
R2777 gnd.n4272 gnd.n4271 585
R2778 gnd.n2268 gnd.n2267 585
R2779 gnd.n2279 gnd.n2268 585
R2780 gnd.n4262 gnd.n4261 585
R2781 gnd.n4263 gnd.n4262 585
R2782 gnd.n2281 gnd.n2280 585
R2783 gnd.n2280 gnd.n2276 585
R2784 gnd.n4257 gnd.n4256 585
R2785 gnd.n4256 gnd.n4255 585
R2786 gnd.n2284 gnd.n2283 585
R2787 gnd.n2285 gnd.n2284 585
R2788 gnd.n4246 gnd.n4245 585
R2789 gnd.n4247 gnd.n4246 585
R2790 gnd.n2297 gnd.n2296 585
R2791 gnd.n2296 gnd.n2293 585
R2792 gnd.n4241 gnd.n4240 585
R2793 gnd.n4240 gnd.n4239 585
R2794 gnd.n2300 gnd.n2299 585
R2795 gnd.n2311 gnd.n2300 585
R2796 gnd.n4230 gnd.n4229 585
R2797 gnd.n4231 gnd.n4230 585
R2798 gnd.n2313 gnd.n2312 585
R2799 gnd.n2312 gnd.n2308 585
R2800 gnd.n4225 gnd.n4224 585
R2801 gnd.n4224 gnd.n4223 585
R2802 gnd.n2316 gnd.n2315 585
R2803 gnd.n2317 gnd.n2316 585
R2804 gnd.n4214 gnd.n4213 585
R2805 gnd.n4215 gnd.n4214 585
R2806 gnd.n2329 gnd.n2328 585
R2807 gnd.n2328 gnd.n2325 585
R2808 gnd.n4209 gnd.n4208 585
R2809 gnd.n4208 gnd.n4207 585
R2810 gnd.n2332 gnd.n2331 585
R2811 gnd.n3977 gnd.n2332 585
R2812 gnd.n4198 gnd.n4197 585
R2813 gnd.n4199 gnd.n4198 585
R2814 gnd.n4194 gnd.n3978 585
R2815 gnd.n4193 gnd.n4192 585
R2816 gnd.n4190 gnd.n3980 585
R2817 gnd.n4190 gnd.n3813 585
R2818 gnd.n4189 gnd.n4188 585
R2819 gnd.n4187 gnd.n4186 585
R2820 gnd.n4185 gnd.n3985 585
R2821 gnd.n4183 gnd.n4182 585
R2822 gnd.n4181 gnd.n3986 585
R2823 gnd.n4180 gnd.n4179 585
R2824 gnd.n4177 gnd.n3991 585
R2825 gnd.n4175 gnd.n4174 585
R2826 gnd.n4173 gnd.n3992 585
R2827 gnd.n4172 gnd.n4171 585
R2828 gnd.n4169 gnd.n3997 585
R2829 gnd.n4167 gnd.n4166 585
R2830 gnd.n4165 gnd.n3998 585
R2831 gnd.n4164 gnd.n4163 585
R2832 gnd.n4161 gnd.n4003 585
R2833 gnd.n4159 gnd.n4158 585
R2834 gnd.n4157 gnd.n4004 585
R2835 gnd.n4156 gnd.n4155 585
R2836 gnd.n4153 gnd.n4012 585
R2837 gnd.n4151 gnd.n4150 585
R2838 gnd.n4149 gnd.n4013 585
R2839 gnd.n4148 gnd.n4147 585
R2840 gnd.n4145 gnd.n4018 585
R2841 gnd.n4143 gnd.n4142 585
R2842 gnd.n4141 gnd.n4019 585
R2843 gnd.n4140 gnd.n4139 585
R2844 gnd.n4137 gnd.n4024 585
R2845 gnd.n4135 gnd.n4134 585
R2846 gnd.n4133 gnd.n4025 585
R2847 gnd.n4132 gnd.n4131 585
R2848 gnd.n4129 gnd.n4030 585
R2849 gnd.n4127 gnd.n4126 585
R2850 gnd.n4125 gnd.n4031 585
R2851 gnd.n4124 gnd.n4036 585
R2852 gnd.n4117 gnd.n4039 585
R2853 gnd.n4120 gnd.n4119 585
R2854 gnd.n2124 gnd.n2123 585
R2855 gnd.n4576 gnd.n4575 585
R2856 gnd.n4578 gnd.n4577 585
R2857 gnd.n4580 gnd.n4579 585
R2858 gnd.n4582 gnd.n4581 585
R2859 gnd.n4584 gnd.n4583 585
R2860 gnd.n4586 gnd.n4585 585
R2861 gnd.n4588 gnd.n4587 585
R2862 gnd.n4590 gnd.n4589 585
R2863 gnd.n4592 gnd.n4591 585
R2864 gnd.n4594 gnd.n4593 585
R2865 gnd.n4596 gnd.n4595 585
R2866 gnd.n4598 gnd.n4597 585
R2867 gnd.n4600 gnd.n4599 585
R2868 gnd.n4602 gnd.n4601 585
R2869 gnd.n4604 gnd.n4603 585
R2870 gnd.n4606 gnd.n4605 585
R2871 gnd.n4608 gnd.n4607 585
R2872 gnd.n4610 gnd.n4609 585
R2873 gnd.n4613 gnd.n4612 585
R2874 gnd.n4611 gnd.n2102 585
R2875 gnd.n4820 gnd.n4819 585
R2876 gnd.n4822 gnd.n4821 585
R2877 gnd.n4824 gnd.n4823 585
R2878 gnd.n4826 gnd.n4825 585
R2879 gnd.n4828 gnd.n4827 585
R2880 gnd.n4830 gnd.n4829 585
R2881 gnd.n4832 gnd.n4831 585
R2882 gnd.n4834 gnd.n4833 585
R2883 gnd.n4836 gnd.n4835 585
R2884 gnd.n4838 gnd.n4837 585
R2885 gnd.n4840 gnd.n4839 585
R2886 gnd.n4842 gnd.n4841 585
R2887 gnd.n4843 gnd.n2083 585
R2888 gnd.n4845 gnd.n4844 585
R2889 gnd.n2084 gnd.n2082 585
R2890 gnd.n2085 gnd.n1108 585
R2891 gnd.n4847 gnd.n1108 585
R2892 gnd.n4571 gnd.n1110 585
R2893 gnd.n6324 gnd.n1110 585
R2894 gnd.n4570 gnd.n4569 585
R2895 gnd.n4569 gnd.n4568 585
R2896 gnd.n2128 gnd.n1101 585
R2897 gnd.n6330 gnd.n1101 585
R2898 gnd.n4529 gnd.n4528 585
R2899 gnd.n4530 gnd.n4529 585
R2900 gnd.n2134 gnd.n1090 585
R2901 gnd.n6336 gnd.n1090 585
R2902 gnd.n4523 gnd.n4522 585
R2903 gnd.n4522 gnd.n4521 585
R2904 gnd.n2136 gnd.n1079 585
R2905 gnd.n6342 gnd.n1079 585
R2906 gnd.n4447 gnd.n2140 585
R2907 gnd.n4513 gnd.n2140 585
R2908 gnd.n4448 gnd.n1069 585
R2909 gnd.n6348 gnd.n1069 585
R2910 gnd.n4450 gnd.n4449 585
R2911 gnd.n4451 gnd.n4450 585
R2912 gnd.n2157 gnd.n1058 585
R2913 gnd.n6354 gnd.n1058 585
R2914 gnd.n4441 gnd.n4440 585
R2915 gnd.n4440 gnd.n4439 585
R2916 gnd.n4438 gnd.n1047 585
R2917 gnd.n6360 gnd.n1047 585
R2918 gnd.n4437 gnd.n2151 585
R2919 gnd.n4462 gnd.n2151 585
R2920 gnd.n2159 gnd.n1037 585
R2921 gnd.n6366 gnd.n1037 585
R2922 gnd.n4433 gnd.n4432 585
R2923 gnd.n4432 gnd.n4431 585
R2924 gnd.n2161 gnd.n1027 585
R2925 gnd.n6372 gnd.n1027 585
R2926 gnd.n4397 gnd.n4396 585
R2927 gnd.n4398 gnd.n4397 585
R2928 gnd.n2178 gnd.n1016 585
R2929 gnd.n6378 gnd.n1016 585
R2930 gnd.n4392 gnd.n4391 585
R2931 gnd.n4391 gnd.n4390 585
R2932 gnd.n4389 gnd.n1005 585
R2933 gnd.n6384 gnd.n1005 585
R2934 gnd.n4388 gnd.n2172 585
R2935 gnd.n4413 gnd.n2172 585
R2936 gnd.n2180 gnd.n995 585
R2937 gnd.n6390 gnd.n995 585
R2938 gnd.n4384 gnd.n4383 585
R2939 gnd.n4383 gnd.n4382 585
R2940 gnd.n2182 gnd.n984 585
R2941 gnd.n6396 gnd.n984 585
R2942 gnd.n4363 gnd.n4362 585
R2943 gnd.n4364 gnd.n4363 585
R2944 gnd.n2186 gnd.n971 585
R2945 gnd.n6402 gnd.n971 585
R2946 gnd.n4358 gnd.n4357 585
R2947 gnd.n4357 gnd.n970 585
R2948 gnd.n4356 gnd.n2188 585
R2949 gnd.n4356 gnd.n4355 585
R2950 gnd.n2209 gnd.n2189 585
R2951 gnd.n2198 gnd.n2189 585
R2952 gnd.n2210 gnd.n2195 585
R2953 gnd.n4348 gnd.n2195 585
R2954 gnd.n2213 gnd.n2211 585
R2955 gnd.n2216 gnd.n2213 585
R2956 gnd.n4331 gnd.n4330 585
R2957 gnd.n4330 gnd.n4329 585
R2958 gnd.n2212 gnd.n2206 585
R2959 gnd.n2214 gnd.n2212 585
R2960 gnd.n4071 gnd.n2222 585
R2961 gnd.n4321 gnd.n2222 585
R2962 gnd.n4073 gnd.n4072 585
R2963 gnd.n4072 gnd.n2221 585
R2964 gnd.n4074 gnd.n2231 585
R2965 gnd.n4312 gnd.n2231 585
R2966 gnd.n4076 gnd.n4075 585
R2967 gnd.n4075 gnd.n2230 585
R2968 gnd.n4077 gnd.n2237 585
R2969 gnd.n4304 gnd.n2237 585
R2970 gnd.n4079 gnd.n4078 585
R2971 gnd.n4078 gnd.n2247 585
R2972 gnd.n4080 gnd.n2245 585
R2973 gnd.n4296 gnd.n2245 585
R2974 gnd.n4082 gnd.n4081 585
R2975 gnd.n4081 gnd.n2244 585
R2976 gnd.n4083 gnd.n2254 585
R2977 gnd.n4287 gnd.n2254 585
R2978 gnd.n4085 gnd.n4084 585
R2979 gnd.n4084 gnd.n2253 585
R2980 gnd.n4086 gnd.n2262 585
R2981 gnd.n4279 gnd.n2262 585
R2982 gnd.n4088 gnd.n4087 585
R2983 gnd.n4087 gnd.n2261 585
R2984 gnd.n4089 gnd.n2269 585
R2985 gnd.n4271 gnd.n2269 585
R2986 gnd.n4091 gnd.n4090 585
R2987 gnd.n4090 gnd.n2279 585
R2988 gnd.n4092 gnd.n2277 585
R2989 gnd.n4263 gnd.n2277 585
R2990 gnd.n4094 gnd.n4093 585
R2991 gnd.n4093 gnd.n2276 585
R2992 gnd.n4095 gnd.n2286 585
R2993 gnd.n4255 gnd.n2286 585
R2994 gnd.n4097 gnd.n4096 585
R2995 gnd.n4096 gnd.n2285 585
R2996 gnd.n4098 gnd.n2294 585
R2997 gnd.n4247 gnd.n2294 585
R2998 gnd.n4100 gnd.n4099 585
R2999 gnd.n4099 gnd.n2293 585
R3000 gnd.n4101 gnd.n2301 585
R3001 gnd.n4239 gnd.n2301 585
R3002 gnd.n4103 gnd.n4102 585
R3003 gnd.n4102 gnd.n2311 585
R3004 gnd.n4104 gnd.n2309 585
R3005 gnd.n4231 gnd.n2309 585
R3006 gnd.n4106 gnd.n4105 585
R3007 gnd.n4105 gnd.n2308 585
R3008 gnd.n4107 gnd.n2318 585
R3009 gnd.n4223 gnd.n2318 585
R3010 gnd.n4109 gnd.n4108 585
R3011 gnd.n4108 gnd.n2317 585
R3012 gnd.n4110 gnd.n2326 585
R3013 gnd.n4215 gnd.n2326 585
R3014 gnd.n4112 gnd.n4111 585
R3015 gnd.n4111 gnd.n2325 585
R3016 gnd.n4113 gnd.n2333 585
R3017 gnd.n4207 gnd.n2333 585
R3018 gnd.n4114 gnd.n4041 585
R3019 gnd.n4041 gnd.n3977 585
R3020 gnd.n4115 gnd.n3814 585
R3021 gnd.n4199 gnd.n3814 585
R3022 gnd.n7664 gnd.n7663 585
R3023 gnd.n7665 gnd.n7664 585
R3024 gnd.n132 gnd.n130 585
R3025 gnd.n130 gnd.n126 585
R3026 gnd.n7584 gnd.n7583 585
R3027 gnd.n7585 gnd.n7584 585
R3028 gnd.n209 gnd.n208 585
R3029 gnd.n208 gnd.n206 585
R3030 gnd.n7579 gnd.n7578 585
R3031 gnd.n7578 gnd.n7577 585
R3032 gnd.n212 gnd.n211 585
R3033 gnd.n213 gnd.n212 585
R3034 gnd.n7500 gnd.n7499 585
R3035 gnd.n7501 gnd.n7500 585
R3036 gnd.n225 gnd.n224 585
R3037 gnd.n232 gnd.n224 585
R3038 gnd.n7495 gnd.n7494 585
R3039 gnd.n7494 gnd.n7493 585
R3040 gnd.n228 gnd.n227 585
R3041 gnd.n229 gnd.n228 585
R3042 gnd.n7484 gnd.n7483 585
R3043 gnd.n7485 gnd.n7484 585
R3044 gnd.n241 gnd.n240 585
R3045 gnd.n247 gnd.n240 585
R3046 gnd.n7479 gnd.n7478 585
R3047 gnd.n7478 gnd.n7477 585
R3048 gnd.n244 gnd.n243 585
R3049 gnd.n254 gnd.n244 585
R3050 gnd.n7468 gnd.n7467 585
R3051 gnd.n7469 gnd.n7468 585
R3052 gnd.n256 gnd.n255 585
R3053 gnd.n263 gnd.n255 585
R3054 gnd.n7463 gnd.n7462 585
R3055 gnd.n7462 gnd.n7461 585
R3056 gnd.n259 gnd.n258 585
R3057 gnd.n260 gnd.n259 585
R3058 gnd.n7452 gnd.n7451 585
R3059 gnd.n7453 gnd.n7452 585
R3060 gnd.n272 gnd.n271 585
R3061 gnd.n271 gnd.n269 585
R3062 gnd.n7447 gnd.n7446 585
R3063 gnd.n7446 gnd.n7445 585
R3064 gnd.n275 gnd.n274 585
R3065 gnd.n284 gnd.n275 585
R3066 gnd.n7436 gnd.n7435 585
R3067 gnd.n7437 gnd.n7436 585
R3068 gnd.n286 gnd.n285 585
R3069 gnd.n293 gnd.n285 585
R3070 gnd.n7431 gnd.n7430 585
R3071 gnd.n7430 gnd.n7429 585
R3072 gnd.n289 gnd.n288 585
R3073 gnd.n290 gnd.n289 585
R3074 gnd.n7420 gnd.n7419 585
R3075 gnd.n7421 gnd.n7420 585
R3076 gnd.n302 gnd.n301 585
R3077 gnd.n301 gnd.n299 585
R3078 gnd.n7396 gnd.n7395 585
R3079 gnd.n7397 gnd.n7396 585
R3080 gnd.n7394 gnd.n332 585
R3081 gnd.n7394 gnd.n7393 585
R3082 gnd.n331 gnd.n330 585
R3083 gnd.n334 gnd.n330 585
R3084 gnd.n7319 gnd.n7318 585
R3085 gnd.n7320 gnd.n7319 585
R3086 gnd.n7317 gnd.n7316 585
R3087 gnd.n7316 gnd.n340 585
R3088 gnd.n7315 gnd.n342 585
R3089 gnd.n7315 gnd.n7314 585
R3090 gnd.n341 gnd.n311 585
R3091 gnd.n315 gnd.n311 585
R3092 gnd.n7414 gnd.n7413 585
R3093 gnd.n7413 gnd.n7412 585
R3094 gnd.n7415 gnd.n310 585
R3095 gnd.n7305 gnd.n310 585
R3096 gnd.n361 gnd.n309 585
R3097 gnd.n361 gnd.n350 585
R3098 gnd.n7289 gnd.n7288 585
R3099 gnd.n7290 gnd.n7289 585
R3100 gnd.n7287 gnd.n360 585
R3101 gnd.n7269 gnd.n360 585
R3102 gnd.n366 gnd.n362 585
R3103 gnd.n7253 gnd.n366 585
R3104 gnd.n7283 gnd.n7282 585
R3105 gnd.n7282 gnd.n7281 585
R3106 gnd.n365 gnd.n364 585
R3107 gnd.n7259 gnd.n365 585
R3108 gnd.n7242 gnd.n394 585
R3109 gnd.n7226 gnd.n394 585
R3110 gnd.n7244 gnd.n7243 585
R3111 gnd.n7245 gnd.n7244 585
R3112 gnd.n395 gnd.n393 585
R3113 gnd.n6004 gnd.n393 585
R3114 gnd.n7237 gnd.n7236 585
R3115 gnd.n7236 gnd.n7235 585
R3116 gnd.n398 gnd.n397 585
R3117 gnd.n5999 gnd.n398 585
R3118 gnd.n6049 gnd.n6048 585
R3119 gnd.n6050 gnd.n6049 585
R3120 gnd.n1366 gnd.n1365 585
R3121 gnd.n1373 gnd.n1365 585
R3122 gnd.n6044 gnd.n6043 585
R3123 gnd.n6043 gnd.n6042 585
R3124 gnd.n1369 gnd.n1368 585
R3125 gnd.n6020 gnd.n1369 585
R3126 gnd.n5979 gnd.n1399 585
R3127 gnd.n1399 gnd.n1398 585
R3128 gnd.n5981 gnd.n5980 585
R3129 gnd.n5982 gnd.n5981 585
R3130 gnd.n1400 gnd.n1397 585
R3131 gnd.n1407 gnd.n1397 585
R3132 gnd.n5974 gnd.n5973 585
R3133 gnd.n5973 gnd.n5972 585
R3134 gnd.n1403 gnd.n1402 585
R3135 gnd.n5959 gnd.n1403 585
R3136 gnd.n5942 gnd.n1426 585
R3137 gnd.n1426 gnd.n1414 585
R3138 gnd.n5944 gnd.n5943 585
R3139 gnd.n5945 gnd.n5944 585
R3140 gnd.n1427 gnd.n1425 585
R3141 gnd.n1435 gnd.n1425 585
R3142 gnd.n5937 gnd.n5936 585
R3143 gnd.n5936 gnd.n5935 585
R3144 gnd.n1430 gnd.n1429 585
R3145 gnd.n5923 gnd.n1430 585
R3146 gnd.n5911 gnd.n5906 585
R3147 gnd.n5906 gnd.n1452 585
R3148 gnd.n5913 gnd.n5912 585
R3149 gnd.n5914 gnd.n5913 585
R3150 gnd.n5907 gnd.n1288 585
R3151 gnd.n6079 gnd.n1288 585
R3152 gnd.n6153 gnd.n6152 585
R3153 gnd.n6151 gnd.n1287 585
R3154 gnd.n6150 gnd.n1286 585
R3155 gnd.n6155 gnd.n1286 585
R3156 gnd.n6149 gnd.n6148 585
R3157 gnd.n6147 gnd.n6146 585
R3158 gnd.n6145 gnd.n6144 585
R3159 gnd.n6143 gnd.n6142 585
R3160 gnd.n6141 gnd.n6140 585
R3161 gnd.n6139 gnd.n6138 585
R3162 gnd.n6137 gnd.n6136 585
R3163 gnd.n6135 gnd.n6134 585
R3164 gnd.n6133 gnd.n6132 585
R3165 gnd.n6131 gnd.n6130 585
R3166 gnd.n6129 gnd.n6128 585
R3167 gnd.n6127 gnd.n6126 585
R3168 gnd.n6125 gnd.n6124 585
R3169 gnd.n6122 gnd.n6121 585
R3170 gnd.n6120 gnd.n6119 585
R3171 gnd.n6118 gnd.n6117 585
R3172 gnd.n6116 gnd.n6115 585
R3173 gnd.n6114 gnd.n6113 585
R3174 gnd.n6112 gnd.n6111 585
R3175 gnd.n6110 gnd.n6109 585
R3176 gnd.n6108 gnd.n6107 585
R3177 gnd.n6106 gnd.n6105 585
R3178 gnd.n6104 gnd.n6103 585
R3179 gnd.n6102 gnd.n6101 585
R3180 gnd.n6100 gnd.n6099 585
R3181 gnd.n6098 gnd.n6097 585
R3182 gnd.n6096 gnd.n6095 585
R3183 gnd.n6094 gnd.n6093 585
R3184 gnd.n6092 gnd.n6091 585
R3185 gnd.n6090 gnd.n6089 585
R3186 gnd.n6088 gnd.n6087 585
R3187 gnd.n6086 gnd.n1328 585
R3188 gnd.n1332 gnd.n1329 585
R3189 gnd.n6082 gnd.n6081 585
R3190 gnd.n200 gnd.n199 585
R3191 gnd.n7593 gnd.n195 585
R3192 gnd.n7595 gnd.n7594 585
R3193 gnd.n7597 gnd.n193 585
R3194 gnd.n7599 gnd.n7598 585
R3195 gnd.n7600 gnd.n188 585
R3196 gnd.n7602 gnd.n7601 585
R3197 gnd.n7604 gnd.n186 585
R3198 gnd.n7606 gnd.n7605 585
R3199 gnd.n7607 gnd.n181 585
R3200 gnd.n7609 gnd.n7608 585
R3201 gnd.n7611 gnd.n179 585
R3202 gnd.n7613 gnd.n7612 585
R3203 gnd.n7614 gnd.n174 585
R3204 gnd.n7616 gnd.n7615 585
R3205 gnd.n7618 gnd.n172 585
R3206 gnd.n7620 gnd.n7619 585
R3207 gnd.n7621 gnd.n167 585
R3208 gnd.n7623 gnd.n7622 585
R3209 gnd.n7625 gnd.n165 585
R3210 gnd.n7627 gnd.n7626 585
R3211 gnd.n7631 gnd.n160 585
R3212 gnd.n7633 gnd.n7632 585
R3213 gnd.n7635 gnd.n158 585
R3214 gnd.n7637 gnd.n7636 585
R3215 gnd.n7638 gnd.n153 585
R3216 gnd.n7640 gnd.n7639 585
R3217 gnd.n7642 gnd.n151 585
R3218 gnd.n7644 gnd.n7643 585
R3219 gnd.n7645 gnd.n146 585
R3220 gnd.n7647 gnd.n7646 585
R3221 gnd.n7649 gnd.n144 585
R3222 gnd.n7651 gnd.n7650 585
R3223 gnd.n7652 gnd.n139 585
R3224 gnd.n7654 gnd.n7653 585
R3225 gnd.n7656 gnd.n137 585
R3226 gnd.n7658 gnd.n7657 585
R3227 gnd.n7659 gnd.n135 585
R3228 gnd.n7660 gnd.n131 585
R3229 gnd.n131 gnd.n128 585
R3230 gnd.n7589 gnd.n127 585
R3231 gnd.n7665 gnd.n127 585
R3232 gnd.n7588 gnd.n7587 585
R3233 gnd.n7587 gnd.n126 585
R3234 gnd.n7586 gnd.n204 585
R3235 gnd.n7586 gnd.n7585 585
R3236 gnd.n7353 gnd.n205 585
R3237 gnd.n206 gnd.n205 585
R3238 gnd.n7354 gnd.n214 585
R3239 gnd.n7577 gnd.n214 585
R3240 gnd.n7356 gnd.n7355 585
R3241 gnd.n7355 gnd.n213 585
R3242 gnd.n7357 gnd.n223 585
R3243 gnd.n7501 gnd.n223 585
R3244 gnd.n7359 gnd.n7358 585
R3245 gnd.n7358 gnd.n232 585
R3246 gnd.n7360 gnd.n230 585
R3247 gnd.n7493 gnd.n230 585
R3248 gnd.n7362 gnd.n7361 585
R3249 gnd.n7361 gnd.n229 585
R3250 gnd.n7363 gnd.n239 585
R3251 gnd.n7485 gnd.n239 585
R3252 gnd.n7365 gnd.n7364 585
R3253 gnd.n7364 gnd.n247 585
R3254 gnd.n7366 gnd.n245 585
R3255 gnd.n7477 gnd.n245 585
R3256 gnd.n7368 gnd.n7367 585
R3257 gnd.n7367 gnd.n254 585
R3258 gnd.n7369 gnd.n253 585
R3259 gnd.n7469 gnd.n253 585
R3260 gnd.n7371 gnd.n7370 585
R3261 gnd.n7370 gnd.n263 585
R3262 gnd.n7372 gnd.n261 585
R3263 gnd.n7461 gnd.n261 585
R3264 gnd.n7374 gnd.n7373 585
R3265 gnd.n7373 gnd.n260 585
R3266 gnd.n7375 gnd.n270 585
R3267 gnd.n7453 gnd.n270 585
R3268 gnd.n7377 gnd.n7376 585
R3269 gnd.n7376 gnd.n269 585
R3270 gnd.n7378 gnd.n276 585
R3271 gnd.n7445 gnd.n276 585
R3272 gnd.n7380 gnd.n7379 585
R3273 gnd.n7379 gnd.n284 585
R3274 gnd.n7381 gnd.n283 585
R3275 gnd.n7437 gnd.n283 585
R3276 gnd.n7383 gnd.n7382 585
R3277 gnd.n7382 gnd.n293 585
R3278 gnd.n7384 gnd.n291 585
R3279 gnd.n7429 gnd.n291 585
R3280 gnd.n7386 gnd.n7385 585
R3281 gnd.n7385 gnd.n290 585
R3282 gnd.n7387 gnd.n300 585
R3283 gnd.n7421 gnd.n300 585
R3284 gnd.n7389 gnd.n7388 585
R3285 gnd.n7388 gnd.n299 585
R3286 gnd.n7390 gnd.n328 585
R3287 gnd.n7397 gnd.n328 585
R3288 gnd.n7392 gnd.n7391 585
R3289 gnd.n7393 gnd.n7392 585
R3290 gnd.n336 gnd.n335 585
R3291 gnd.n335 gnd.n334 585
R3292 gnd.n7322 gnd.n7321 585
R3293 gnd.n7321 gnd.n7320 585
R3294 gnd.n339 gnd.n338 585
R3295 gnd.n340 gnd.n339 585
R3296 gnd.n7299 gnd.n343 585
R3297 gnd.n7314 gnd.n343 585
R3298 gnd.n7301 gnd.n7300 585
R3299 gnd.n7300 gnd.n315 585
R3300 gnd.n7302 gnd.n313 585
R3301 gnd.n7412 gnd.n313 585
R3302 gnd.n7304 gnd.n7303 585
R3303 gnd.n7305 gnd.n7304 585
R3304 gnd.n352 gnd.n351 585
R3305 gnd.n351 gnd.n350 585
R3306 gnd.n7292 gnd.n7291 585
R3307 gnd.n7291 gnd.n7290 585
R3308 gnd.n355 gnd.n354 585
R3309 gnd.n7269 gnd.n355 585
R3310 gnd.n7255 gnd.n7254 585
R3311 gnd.n7254 gnd.n7253 585
R3312 gnd.n7256 gnd.n368 585
R3313 gnd.n7281 gnd.n368 585
R3314 gnd.n7258 gnd.n7257 585
R3315 gnd.n7259 gnd.n7258 585
R3316 gnd.n386 gnd.n385 585
R3317 gnd.n7226 gnd.n385 585
R3318 gnd.n7247 gnd.n7246 585
R3319 gnd.n7246 gnd.n7245 585
R3320 gnd.n389 gnd.n388 585
R3321 gnd.n6004 gnd.n389 585
R3322 gnd.n5996 gnd.n400 585
R3323 gnd.n7235 gnd.n400 585
R3324 gnd.n5998 gnd.n5997 585
R3325 gnd.n5999 gnd.n5998 585
R3326 gnd.n1387 gnd.n1362 585
R3327 gnd.n6050 gnd.n1362 585
R3328 gnd.n5991 gnd.n5990 585
R3329 gnd.n5990 gnd.n1373 585
R3330 gnd.n5989 gnd.n1371 585
R3331 gnd.n6042 gnd.n1371 585
R3332 gnd.n5988 gnd.n1380 585
R3333 gnd.n6020 gnd.n1380 585
R3334 gnd.n1393 gnd.n1389 585
R3335 gnd.n1398 gnd.n1393 585
R3336 gnd.n5984 gnd.n5983 585
R3337 gnd.n5983 gnd.n5982 585
R3338 gnd.n1392 gnd.n1391 585
R3339 gnd.n1407 gnd.n1392 585
R3340 gnd.n1465 gnd.n1405 585
R3341 gnd.n5972 gnd.n1405 585
R3342 gnd.n1466 gnd.n1415 585
R3343 gnd.n5959 gnd.n1415 585
R3344 gnd.n1468 gnd.n1467 585
R3345 gnd.n1467 gnd.n1414 585
R3346 gnd.n1469 gnd.n1423 585
R3347 gnd.n5945 gnd.n1423 585
R3348 gnd.n1471 gnd.n1470 585
R3349 gnd.n1470 gnd.n1435 585
R3350 gnd.n1472 gnd.n1432 585
R3351 gnd.n5935 gnd.n1432 585
R3352 gnd.n1474 gnd.n1473 585
R3353 gnd.n5923 gnd.n1474 585
R3354 gnd.n1454 gnd.n1453 585
R3355 gnd.n1453 gnd.n1452 585
R3356 gnd.n1455 gnd.n1334 585
R3357 gnd.n5914 gnd.n1334 585
R3358 gnd.n6080 gnd.n1335 585
R3359 gnd.n6080 gnd.n6079 585
R3360 gnd.n5375 gnd.n5184 585
R3361 gnd.n5184 gnd.n1684 585
R3362 gnd.n5377 gnd.n5376 585
R3363 gnd.n5378 gnd.n5377 585
R3364 gnd.n5178 gnd.n5177 585
R3365 gnd.n5178 gnd.n1693 585
R3366 gnd.n5386 gnd.n5385 585
R3367 gnd.n5385 gnd.n5384 585
R3368 gnd.n5387 gnd.n5175 585
R3369 gnd.n5179 gnd.n5175 585
R3370 gnd.n5389 gnd.n5388 585
R3371 gnd.n5390 gnd.n5389 585
R3372 gnd.n5176 gnd.n5166 585
R3373 gnd.n5166 gnd.n1699 585
R3374 gnd.n5398 gnd.n5167 585
R3375 gnd.n5398 gnd.n5397 585
R3376 gnd.n5399 gnd.n5165 585
R3377 gnd.n5399 gnd.n1707 585
R3378 gnd.n5401 gnd.n5400 585
R3379 gnd.n5400 gnd.n1706 585
R3380 gnd.n5402 gnd.n5163 585
R3381 gnd.n5163 gnd.n5162 585
R3382 gnd.n5404 gnd.n5403 585
R3383 gnd.n5405 gnd.n5404 585
R3384 gnd.n5164 gnd.n5160 585
R3385 gnd.n5160 gnd.n1713 585
R3386 gnd.n5154 gnd.n5153 585
R3387 gnd.n5412 gnd.n5154 585
R3388 gnd.n5415 gnd.n5414 585
R3389 gnd.n5414 gnd.n5413 585
R3390 gnd.n5416 gnd.n5150 585
R3391 gnd.n5150 gnd.n1720 585
R3392 gnd.n5418 gnd.n5417 585
R3393 gnd.n5419 gnd.n5418 585
R3394 gnd.n5152 gnd.n5149 585
R3395 gnd.n5149 gnd.n5147 585
R3396 gnd.n5151 gnd.n5139 585
R3397 gnd.n5425 gnd.n5139 585
R3398 gnd.n5428 gnd.n5138 585
R3399 gnd.n5428 gnd.n5427 585
R3400 gnd.n5430 gnd.n5429 585
R3401 gnd.n5429 gnd.n1732 585
R3402 gnd.n5431 gnd.n5136 585
R3403 gnd.n5136 gnd.n5135 585
R3404 gnd.n5433 gnd.n5432 585
R3405 gnd.n5434 gnd.n5433 585
R3406 gnd.n5137 gnd.n5134 585
R3407 gnd.n5134 gnd.n1739 585
R3408 gnd.n5126 gnd.n5125 585
R3409 gnd.n5440 gnd.n5126 585
R3410 gnd.n5444 gnd.n5443 585
R3411 gnd.n5443 gnd.n5442 585
R3412 gnd.n5445 gnd.n5122 585
R3413 gnd.n5122 gnd.n1745 585
R3414 gnd.n5447 gnd.n5446 585
R3415 gnd.n5448 gnd.n5447 585
R3416 gnd.n5124 gnd.n5121 585
R3417 gnd.n5121 gnd.n1753 585
R3418 gnd.n5123 gnd.n1751 585
R3419 gnd.n5708 gnd.n1751 585
R3420 gnd.n5114 gnd.n5113 585
R3421 gnd.n5455 gnd.n5114 585
R3422 gnd.n5459 gnd.n5458 585
R3423 gnd.n5458 gnd.n5457 585
R3424 gnd.n5460 gnd.n5110 585
R3425 gnd.n5110 gnd.n1760 585
R3426 gnd.n5462 gnd.n5461 585
R3427 gnd.n5463 gnd.n5462 585
R3428 gnd.n5112 gnd.n5109 585
R3429 gnd.n5109 gnd.n1768 585
R3430 gnd.n5111 gnd.n5100 585
R3431 gnd.n5100 gnd.n1766 585
R3432 gnd.n5471 gnd.n5099 585
R3433 gnd.n5471 gnd.n5470 585
R3434 gnd.n5473 gnd.n5472 585
R3435 gnd.n5472 gnd.n1775 585
R3436 gnd.n5474 gnd.n5096 585
R3437 gnd.n5096 gnd.n1774 585
R3438 gnd.n5476 gnd.n5475 585
R3439 gnd.n5477 gnd.n5476 585
R3440 gnd.n5098 gnd.n5095 585
R3441 gnd.n5095 gnd.n1783 585
R3442 gnd.n5097 gnd.n5086 585
R3443 gnd.n5086 gnd.n1781 585
R3444 gnd.n5485 gnd.n5085 585
R3445 gnd.n5485 gnd.n5484 585
R3446 gnd.n5487 gnd.n5486 585
R3447 gnd.n5486 gnd.n1790 585
R3448 gnd.n5488 gnd.n5082 585
R3449 gnd.n5082 gnd.n1789 585
R3450 gnd.n5490 gnd.n5489 585
R3451 gnd.n5491 gnd.n5490 585
R3452 gnd.n5084 gnd.n5081 585
R3453 gnd.n5081 gnd.n1798 585
R3454 gnd.n5083 gnd.n5072 585
R3455 gnd.n5072 gnd.n1796 585
R3456 gnd.n5499 gnd.n5071 585
R3457 gnd.n5499 gnd.n5498 585
R3458 gnd.n5501 gnd.n5500 585
R3459 gnd.n5500 gnd.n1805 585
R3460 gnd.n5502 gnd.n5068 585
R3461 gnd.n5068 gnd.n1804 585
R3462 gnd.n5504 gnd.n5503 585
R3463 gnd.n5505 gnd.n5504 585
R3464 gnd.n5070 gnd.n5067 585
R3465 gnd.n5067 gnd.n1813 585
R3466 gnd.n5069 gnd.n5060 585
R3467 gnd.n5060 gnd.n1811 585
R3468 gnd.n5513 gnd.n5059 585
R3469 gnd.n5513 gnd.n5512 585
R3470 gnd.n5515 gnd.n5514 585
R3471 gnd.n5514 gnd.n1820 585
R3472 gnd.n5516 gnd.n5056 585
R3473 gnd.n5056 gnd.n1819 585
R3474 gnd.n5518 gnd.n5517 585
R3475 gnd.n5519 gnd.n5518 585
R3476 gnd.n5058 gnd.n5055 585
R3477 gnd.n5055 gnd.n1827 585
R3478 gnd.n5057 gnd.n5045 585
R3479 gnd.n5525 gnd.n5045 585
R3480 gnd.n5528 gnd.n5044 585
R3481 gnd.n5528 gnd.n5527 585
R3482 gnd.n5530 gnd.n5529 585
R3483 gnd.n5529 gnd.n1834 585
R3484 gnd.n5531 gnd.n5041 585
R3485 gnd.n5041 gnd.n1833 585
R3486 gnd.n5533 gnd.n5532 585
R3487 gnd.n5534 gnd.n5533 585
R3488 gnd.n5043 gnd.n5040 585
R3489 gnd.n5040 gnd.n1842 585
R3490 gnd.n5042 gnd.n5032 585
R3491 gnd.n5032 gnd.n1840 585
R3492 gnd.n5543 gnd.n5031 585
R3493 gnd.n5543 gnd.n5542 585
R3494 gnd.n5545 gnd.n5544 585
R3495 gnd.n5544 gnd.n1849 585
R3496 gnd.n5546 gnd.n5028 585
R3497 gnd.n5028 gnd.n1848 585
R3498 gnd.n5548 gnd.n5547 585
R3499 gnd.n5549 gnd.n5548 585
R3500 gnd.n5030 gnd.n5027 585
R3501 gnd.n5027 gnd.n1857 585
R3502 gnd.n5029 gnd.n5019 585
R3503 gnd.n5019 gnd.n1855 585
R3504 gnd.n5558 gnd.n5018 585
R3505 gnd.n5558 gnd.n5557 585
R3506 gnd.n5560 gnd.n5559 585
R3507 gnd.n5559 gnd.n1863 585
R3508 gnd.n5561 gnd.n1889 585
R3509 gnd.n1889 gnd.n1888 585
R3510 gnd.n5563 gnd.n5562 585
R3511 gnd.n5564 gnd.n5563 585
R3512 gnd.n5017 gnd.n1887 585
R3513 gnd.n1887 gnd.n1871 585
R3514 gnd.n5016 gnd.n5015 585
R3515 gnd.n5015 gnd.n1869 585
R3516 gnd.n5014 gnd.n5011 585
R3517 gnd.n5014 gnd.n5013 585
R3518 gnd.n5010 gnd.n1878 585
R3519 gnd.n5572 gnd.n1878 585
R3520 gnd.n5009 gnd.n5008 585
R3521 gnd.n5008 gnd.n1877 585
R3522 gnd.n5007 gnd.n1890 585
R3523 gnd.n5007 gnd.n5006 585
R3524 gnd.n4745 gnd.n1891 585
R3525 gnd.n4641 gnd.n1891 585
R3526 gnd.n4747 gnd.n4746 585
R3527 gnd.n4748 gnd.n4747 585
R3528 gnd.n4743 gnd.n4642 585
R3529 gnd.n4742 gnd.n4741 585
R3530 gnd.n4739 gnd.n4663 585
R3531 gnd.n4739 gnd.n1901 585
R3532 gnd.n4738 gnd.n4737 585
R3533 gnd.n4736 gnd.n4735 585
R3534 gnd.n4734 gnd.n4665 585
R3535 gnd.n4732 gnd.n4731 585
R3536 gnd.n4730 gnd.n4666 585
R3537 gnd.n4729 gnd.n4728 585
R3538 gnd.n4726 gnd.n4667 585
R3539 gnd.n4724 gnd.n4723 585
R3540 gnd.n4722 gnd.n4668 585
R3541 gnd.n4721 gnd.n4720 585
R3542 gnd.n4718 gnd.n4669 585
R3543 gnd.n4716 gnd.n4715 585
R3544 gnd.n4714 gnd.n4670 585
R3545 gnd.n4713 gnd.n4712 585
R3546 gnd.n4710 gnd.n4671 585
R3547 gnd.n4708 gnd.n4707 585
R3548 gnd.n4706 gnd.n4672 585
R3549 gnd.n4705 gnd.n4704 585
R3550 gnd.n4702 gnd.n4673 585
R3551 gnd.n4700 gnd.n4699 585
R3552 gnd.n4698 gnd.n4674 585
R3553 gnd.n4697 gnd.n4696 585
R3554 gnd.n4694 gnd.n4675 585
R3555 gnd.n4692 gnd.n4691 585
R3556 gnd.n4690 gnd.n4676 585
R3557 gnd.n4689 gnd.n4688 585
R3558 gnd.n4686 gnd.n4685 585
R3559 gnd.n4684 gnd.n4683 585
R3560 gnd.n4682 gnd.n4618 585
R3561 gnd.n4817 gnd.n4816 585
R3562 gnd.n4814 gnd.n4617 585
R3563 gnd.n4812 gnd.n4811 585
R3564 gnd.n4810 gnd.n4620 585
R3565 gnd.n4808 gnd.n4807 585
R3566 gnd.n4805 gnd.n4623 585
R3567 gnd.n4803 gnd.n4802 585
R3568 gnd.n4801 gnd.n4624 585
R3569 gnd.n4800 gnd.n4799 585
R3570 gnd.n4797 gnd.n4625 585
R3571 gnd.n4795 gnd.n4794 585
R3572 gnd.n4793 gnd.n4626 585
R3573 gnd.n4792 gnd.n4791 585
R3574 gnd.n4789 gnd.n4627 585
R3575 gnd.n4787 gnd.n4786 585
R3576 gnd.n4785 gnd.n4628 585
R3577 gnd.n4784 gnd.n4783 585
R3578 gnd.n4781 gnd.n4629 585
R3579 gnd.n4779 gnd.n4778 585
R3580 gnd.n4777 gnd.n4630 585
R3581 gnd.n4776 gnd.n4775 585
R3582 gnd.n4773 gnd.n4631 585
R3583 gnd.n4771 gnd.n4770 585
R3584 gnd.n4769 gnd.n4632 585
R3585 gnd.n4768 gnd.n4767 585
R3586 gnd.n4765 gnd.n4633 585
R3587 gnd.n4763 gnd.n4762 585
R3588 gnd.n4761 gnd.n4634 585
R3589 gnd.n4760 gnd.n4759 585
R3590 gnd.n4757 gnd.n4635 585
R3591 gnd.n4755 gnd.n4754 585
R3592 gnd.n4753 gnd.n4636 585
R3593 gnd.n4752 gnd.n4751 585
R3594 gnd.n5256 gnd.n5255 585
R3595 gnd.n5257 gnd.n5253 585
R3596 gnd.n5259 gnd.n5258 585
R3597 gnd.n5261 gnd.n5251 585
R3598 gnd.n5263 gnd.n5262 585
R3599 gnd.n5264 gnd.n5250 585
R3600 gnd.n5266 gnd.n5265 585
R3601 gnd.n5268 gnd.n5248 585
R3602 gnd.n5270 gnd.n5269 585
R3603 gnd.n5271 gnd.n5247 585
R3604 gnd.n5273 gnd.n5272 585
R3605 gnd.n5275 gnd.n5245 585
R3606 gnd.n5277 gnd.n5276 585
R3607 gnd.n5278 gnd.n5244 585
R3608 gnd.n5280 gnd.n5279 585
R3609 gnd.n5282 gnd.n5242 585
R3610 gnd.n5284 gnd.n5283 585
R3611 gnd.n5285 gnd.n5241 585
R3612 gnd.n5287 gnd.n5286 585
R3613 gnd.n5289 gnd.n5239 585
R3614 gnd.n5291 gnd.n5290 585
R3615 gnd.n5292 gnd.n5238 585
R3616 gnd.n5294 gnd.n5293 585
R3617 gnd.n5296 gnd.n5236 585
R3618 gnd.n5298 gnd.n5297 585
R3619 gnd.n5299 gnd.n5235 585
R3620 gnd.n5301 gnd.n5300 585
R3621 gnd.n5303 gnd.n5233 585
R3622 gnd.n5305 gnd.n5304 585
R3623 gnd.n5307 gnd.n5230 585
R3624 gnd.n5309 gnd.n5308 585
R3625 gnd.n5311 gnd.n5229 585
R3626 gnd.n5312 gnd.n1687 585
R3627 gnd.n5315 gnd.n1305 585
R3628 gnd.n5317 gnd.n5316 585
R3629 gnd.n5319 gnd.n5227 585
R3630 gnd.n5321 gnd.n5320 585
R3631 gnd.n5323 gnd.n5224 585
R3632 gnd.n5325 gnd.n5324 585
R3633 gnd.n5327 gnd.n5222 585
R3634 gnd.n5329 gnd.n5328 585
R3635 gnd.n5330 gnd.n5221 585
R3636 gnd.n5332 gnd.n5331 585
R3637 gnd.n5334 gnd.n5219 585
R3638 gnd.n5336 gnd.n5335 585
R3639 gnd.n5337 gnd.n5218 585
R3640 gnd.n5339 gnd.n5338 585
R3641 gnd.n5341 gnd.n5216 585
R3642 gnd.n5343 gnd.n5342 585
R3643 gnd.n5344 gnd.n5215 585
R3644 gnd.n5346 gnd.n5345 585
R3645 gnd.n5348 gnd.n5213 585
R3646 gnd.n5350 gnd.n5349 585
R3647 gnd.n5351 gnd.n5212 585
R3648 gnd.n5353 gnd.n5352 585
R3649 gnd.n5355 gnd.n5210 585
R3650 gnd.n5357 gnd.n5356 585
R3651 gnd.n5358 gnd.n5209 585
R3652 gnd.n5360 gnd.n5359 585
R3653 gnd.n5362 gnd.n5207 585
R3654 gnd.n5364 gnd.n5363 585
R3655 gnd.n5365 gnd.n5206 585
R3656 gnd.n5367 gnd.n5366 585
R3657 gnd.n5369 gnd.n5205 585
R3658 gnd.n5370 gnd.n5204 585
R3659 gnd.n5373 gnd.n5372 585
R3660 gnd.n5182 gnd.n5181 585
R3661 gnd.n5182 gnd.n1684 585
R3662 gnd.n5380 gnd.n5379 585
R3663 gnd.n5379 gnd.n5378 585
R3664 gnd.n5381 gnd.n5180 585
R3665 gnd.n5180 gnd.n1693 585
R3666 gnd.n5383 gnd.n5382 585
R3667 gnd.n5384 gnd.n5383 585
R3668 gnd.n5174 gnd.n5173 585
R3669 gnd.n5179 gnd.n5174 585
R3670 gnd.n5392 gnd.n5391 585
R3671 gnd.n5391 gnd.n5390 585
R3672 gnd.n5393 gnd.n5169 585
R3673 gnd.n5169 gnd.n1699 585
R3674 gnd.n5395 gnd.n5394 585
R3675 gnd.n5397 gnd.n5395 585
R3676 gnd.n5172 gnd.n5168 585
R3677 gnd.n5168 gnd.n1707 585
R3678 gnd.n5171 gnd.n5170 585
R3679 gnd.n5170 gnd.n1706 585
R3680 gnd.n5159 gnd.n5158 585
R3681 gnd.n5162 gnd.n5159 585
R3682 gnd.n5407 gnd.n5406 585
R3683 gnd.n5406 gnd.n5405 585
R3684 gnd.n5408 gnd.n5156 585
R3685 gnd.n5156 gnd.n1713 585
R3686 gnd.n5410 gnd.n5409 585
R3687 gnd.n5412 gnd.n5410 585
R3688 gnd.n5157 gnd.n5155 585
R3689 gnd.n5413 gnd.n5155 585
R3690 gnd.n5146 gnd.n5145 585
R3691 gnd.n5146 gnd.n1720 585
R3692 gnd.n5421 gnd.n5420 585
R3693 gnd.n5420 gnd.n5419 585
R3694 gnd.n5422 gnd.n5141 585
R3695 gnd.n5147 gnd.n5141 585
R3696 gnd.n5424 gnd.n5423 585
R3697 gnd.n5425 gnd.n5424 585
R3698 gnd.n5144 gnd.n5140 585
R3699 gnd.n5427 gnd.n5140 585
R3700 gnd.n5143 gnd.n5142 585
R3701 gnd.n5142 gnd.n1732 585
R3702 gnd.n5132 gnd.n5131 585
R3703 gnd.n5135 gnd.n5132 585
R3704 gnd.n5436 gnd.n5435 585
R3705 gnd.n5435 gnd.n5434 585
R3706 gnd.n5437 gnd.n5128 585
R3707 gnd.n5128 gnd.n1739 585
R3708 gnd.n5439 gnd.n5438 585
R3709 gnd.n5440 gnd.n5439 585
R3710 gnd.n5130 gnd.n5127 585
R3711 gnd.n5442 gnd.n5127 585
R3712 gnd.n5129 gnd.n5119 585
R3713 gnd.n5119 gnd.n1745 585
R3714 gnd.n5449 gnd.n5118 585
R3715 gnd.n5449 gnd.n5448 585
R3716 gnd.n5451 gnd.n5450 585
R3717 gnd.n5450 gnd.n1753 585
R3718 gnd.n5452 gnd.n1754 585
R3719 gnd.n5708 gnd.n1754 585
R3720 gnd.n5454 gnd.n5453 585
R3721 gnd.n5455 gnd.n5454 585
R3722 gnd.n5117 gnd.n5115 585
R3723 gnd.n5457 gnd.n5115 585
R3724 gnd.n5116 gnd.n5107 585
R3725 gnd.n5107 gnd.n1760 585
R3726 gnd.n5464 gnd.n5106 585
R3727 gnd.n5464 gnd.n5463 585
R3728 gnd.n5466 gnd.n5465 585
R3729 gnd.n5465 gnd.n1768 585
R3730 gnd.n5467 gnd.n5103 585
R3731 gnd.n5103 gnd.n1766 585
R3732 gnd.n5469 gnd.n5468 585
R3733 gnd.n5470 gnd.n5469 585
R3734 gnd.n5105 gnd.n5102 585
R3735 gnd.n5102 gnd.n1775 585
R3736 gnd.n5104 gnd.n5093 585
R3737 gnd.n5093 gnd.n1774 585
R3738 gnd.n5478 gnd.n5092 585
R3739 gnd.n5478 gnd.n5477 585
R3740 gnd.n5480 gnd.n5479 585
R3741 gnd.n5479 gnd.n1783 585
R3742 gnd.n5481 gnd.n5089 585
R3743 gnd.n5089 gnd.n1781 585
R3744 gnd.n5483 gnd.n5482 585
R3745 gnd.n5484 gnd.n5483 585
R3746 gnd.n5091 gnd.n5088 585
R3747 gnd.n5088 gnd.n1790 585
R3748 gnd.n5090 gnd.n5079 585
R3749 gnd.n5079 gnd.n1789 585
R3750 gnd.n5492 gnd.n5078 585
R3751 gnd.n5492 gnd.n5491 585
R3752 gnd.n5494 gnd.n5493 585
R3753 gnd.n5493 gnd.n1798 585
R3754 gnd.n5495 gnd.n5075 585
R3755 gnd.n5075 gnd.n1796 585
R3756 gnd.n5497 gnd.n5496 585
R3757 gnd.n5498 gnd.n5497 585
R3758 gnd.n5077 gnd.n5074 585
R3759 gnd.n5074 gnd.n1805 585
R3760 gnd.n5076 gnd.n5065 585
R3761 gnd.n5065 gnd.n1804 585
R3762 gnd.n5506 gnd.n5064 585
R3763 gnd.n5506 gnd.n5505 585
R3764 gnd.n5508 gnd.n5507 585
R3765 gnd.n5507 gnd.n1813 585
R3766 gnd.n5509 gnd.n5062 585
R3767 gnd.n5062 gnd.n1811 585
R3768 gnd.n5511 gnd.n5510 585
R3769 gnd.n5512 gnd.n5511 585
R3770 gnd.n5063 gnd.n5061 585
R3771 gnd.n5061 gnd.n1820 585
R3772 gnd.n5053 gnd.n5052 585
R3773 gnd.n5053 gnd.n1819 585
R3774 gnd.n5521 gnd.n5520 585
R3775 gnd.n5520 gnd.n5519 585
R3776 gnd.n5522 gnd.n5047 585
R3777 gnd.n5047 gnd.n1827 585
R3778 gnd.n5524 gnd.n5523 585
R3779 gnd.n5525 gnd.n5524 585
R3780 gnd.n5051 gnd.n5046 585
R3781 gnd.n5527 gnd.n5046 585
R3782 gnd.n5050 gnd.n5049 585
R3783 gnd.n5049 gnd.n1834 585
R3784 gnd.n5048 gnd.n5038 585
R3785 gnd.n5038 gnd.n1833 585
R3786 gnd.n5535 gnd.n5037 585
R3787 gnd.n5535 gnd.n5534 585
R3788 gnd.n5537 gnd.n5536 585
R3789 gnd.n5536 gnd.n1842 585
R3790 gnd.n5538 gnd.n5034 585
R3791 gnd.n5034 gnd.n1840 585
R3792 gnd.n5540 gnd.n5539 585
R3793 gnd.n5542 gnd.n5540 585
R3794 gnd.n5036 gnd.n5033 585
R3795 gnd.n5033 gnd.n1849 585
R3796 gnd.n5035 gnd.n5025 585
R3797 gnd.n5025 gnd.n1848 585
R3798 gnd.n5550 gnd.n5024 585
R3799 gnd.n5550 gnd.n5549 585
R3800 gnd.n5552 gnd.n5551 585
R3801 gnd.n5551 gnd.n1857 585
R3802 gnd.n5553 gnd.n5021 585
R3803 gnd.n5021 gnd.n1855 585
R3804 gnd.n5555 gnd.n5554 585
R3805 gnd.n5557 gnd.n5555 585
R3806 gnd.n5023 gnd.n5020 585
R3807 gnd.n5020 gnd.n1863 585
R3808 gnd.n5022 gnd.n1884 585
R3809 gnd.n1888 gnd.n1884 585
R3810 gnd.n5565 gnd.n1885 585
R3811 gnd.n5565 gnd.n5564 585
R3812 gnd.n5566 gnd.n1883 585
R3813 gnd.n5566 gnd.n1871 585
R3814 gnd.n5568 gnd.n5567 585
R3815 gnd.n5567 gnd.n1869 585
R3816 gnd.n5569 gnd.n1881 585
R3817 gnd.n5013 gnd.n1881 585
R3818 gnd.n5571 gnd.n5570 585
R3819 gnd.n5572 gnd.n5571 585
R3820 gnd.n1882 gnd.n1880 585
R3821 gnd.n1880 gnd.n1877 585
R3822 gnd.n4638 gnd.n1894 585
R3823 gnd.n5006 gnd.n1894 585
R3824 gnd.n4640 gnd.n4639 585
R3825 gnd.n4641 gnd.n4640 585
R3826 gnd.n4749 gnd.n4637 585
R3827 gnd.n4749 gnd.n4748 585
R3828 gnd.n6409 gnd.n963 585
R3829 gnd.n2197 gnd.n963 585
R3830 gnd.n7213 gnd.n7212 585
R3831 gnd.n7213 gnd.n312 585
R3832 gnd.n7215 gnd.n7214 585
R3833 gnd.n7214 gnd.n358 585
R3834 gnd.n7216 gnd.n416 585
R3835 gnd.n416 gnd.n356 585
R3836 gnd.n7218 gnd.n7217 585
R3837 gnd.n7218 gnd.n377 585
R3838 gnd.n7219 gnd.n415 585
R3839 gnd.n7219 gnd.n370 585
R3840 gnd.n7221 gnd.n7220 585
R3841 gnd.n7220 gnd.n367 585
R3842 gnd.n7222 gnd.n410 585
R3843 gnd.n410 gnd.n384 585
R3844 gnd.n7224 gnd.n7223 585
R3845 gnd.n7225 gnd.n7224 585
R3846 gnd.n411 gnd.n409 585
R3847 gnd.n409 gnd.n390 585
R3848 gnd.n6034 gnd.n6033 585
R3849 gnd.n6034 gnd.n402 585
R3850 gnd.n6035 gnd.n6029 585
R3851 gnd.n6035 gnd.n399 585
R3852 gnd.n6037 gnd.n6036 585
R3853 gnd.n6036 gnd.n1364 585
R3854 gnd.n6038 gnd.n1375 585
R3855 gnd.n1375 gnd.n1361 585
R3856 gnd.n6040 gnd.n6039 585
R3857 gnd.n6041 gnd.n6040 585
R3858 gnd.n1376 gnd.n1374 585
R3859 gnd.n1374 gnd.n1370 585
R3860 gnd.n6023 gnd.n6022 585
R3861 gnd.n6022 gnd.n6021 585
R3862 gnd.n1379 gnd.n1378 585
R3863 gnd.n1396 gnd.n1379 585
R3864 gnd.n5967 gnd.n1409 585
R3865 gnd.n1409 gnd.n1394 585
R3866 gnd.n5969 gnd.n5968 585
R3867 gnd.n5970 gnd.n5969 585
R3868 gnd.n1410 gnd.n1408 585
R3869 gnd.n1408 gnd.n1404 585
R3870 gnd.n5962 gnd.n5961 585
R3871 gnd.n5961 gnd.n5960 585
R3872 gnd.n1413 gnd.n1412 585
R3873 gnd.n1424 gnd.n1413 585
R3874 gnd.n5931 gnd.n1437 585
R3875 gnd.n1437 gnd.n1422 585
R3876 gnd.n5933 gnd.n5932 585
R3877 gnd.n5934 gnd.n5933 585
R3878 gnd.n1438 gnd.n1436 585
R3879 gnd.n1436 gnd.n1431 585
R3880 gnd.n5926 gnd.n5925 585
R3881 gnd.n5925 gnd.n5924 585
R3882 gnd.n1451 gnd.n1440 585
R3883 gnd.n5905 gnd.n1451 585
R3884 gnd.n1450 gnd.n1449 585
R3885 gnd.n1450 gnd.n1338 585
R3886 gnd.n1442 gnd.n1441 585
R3887 gnd.n1441 gnd.n1336 585
R3888 gnd.n1445 gnd.n1444 585
R3889 gnd.n1444 gnd.n1285 585
R3890 gnd.n1255 gnd.n1254 585
R3891 gnd.n6156 gnd.n1255 585
R3892 gnd.n6159 gnd.n6158 585
R3893 gnd.n6158 gnd.n6157 585
R3894 gnd.n6160 gnd.n1249 585
R3895 gnd.n1256 gnd.n1249 585
R3896 gnd.n6162 gnd.n6161 585
R3897 gnd.n6163 gnd.n6162 585
R3898 gnd.n1250 gnd.n1246 585
R3899 gnd.n6164 gnd.n1246 585
R3900 gnd.n5870 gnd.n1621 585
R3901 gnd.n1621 gnd.n1245 585
R3902 gnd.n5872 gnd.n5871 585
R3903 gnd.n5873 gnd.n5872 585
R3904 gnd.n1622 gnd.n1620 585
R3905 gnd.n1620 gnd.n1618 585
R3906 gnd.n5864 gnd.n5863 585
R3907 gnd.n5863 gnd.n5862 585
R3908 gnd.n1625 gnd.n1624 585
R3909 gnd.n1626 gnd.n1625 585
R3910 gnd.n5851 gnd.n5850 585
R3911 gnd.n5852 gnd.n5851 585
R3912 gnd.n1635 gnd.n1634 585
R3913 gnd.n1640 gnd.n1634 585
R3914 gnd.n5846 gnd.n5845 585
R3915 gnd.n5845 gnd.n5844 585
R3916 gnd.n1638 gnd.n1637 585
R3917 gnd.n1639 gnd.n1638 585
R3918 gnd.n5835 gnd.n5834 585
R3919 gnd.n5836 gnd.n5835 585
R3920 gnd.n1649 gnd.n1648 585
R3921 gnd.n1648 gnd.n1646 585
R3922 gnd.n5830 gnd.n5829 585
R3923 gnd.n5829 gnd.n5828 585
R3924 gnd.n1652 gnd.n1651 585
R3925 gnd.n1653 gnd.n1652 585
R3926 gnd.n5819 gnd.n5818 585
R3927 gnd.n5820 gnd.n5819 585
R3928 gnd.n1662 gnd.n1661 585
R3929 gnd.n1661 gnd.n1659 585
R3930 gnd.n5814 gnd.n5813 585
R3931 gnd.n5813 gnd.n5812 585
R3932 gnd.n1665 gnd.n1664 585
R3933 gnd.n1666 gnd.n1665 585
R3934 gnd.n5803 gnd.n5802 585
R3935 gnd.n5804 gnd.n5803 585
R3936 gnd.n1675 gnd.n1674 585
R3937 gnd.n1674 gnd.n1672 585
R3938 gnd.n5798 gnd.n5797 585
R3939 gnd.n5797 gnd.n5796 585
R3940 gnd.n1678 gnd.n1677 585
R3941 gnd.n1686 gnd.n1678 585
R3942 gnd.n5787 gnd.n5786 585
R3943 gnd.n5788 gnd.n5787 585
R3944 gnd.n1689 gnd.n1688 585
R3945 gnd.n5183 gnd.n1688 585
R3946 gnd.n5782 gnd.n5781 585
R3947 gnd.n5781 gnd.n5780 585
R3948 gnd.n1692 gnd.n1691 585
R3949 gnd.n5179 gnd.n1692 585
R3950 gnd.n5771 gnd.n5770 585
R3951 gnd.n5772 gnd.n5771 585
R3952 gnd.n1702 gnd.n1701 585
R3953 gnd.n5396 gnd.n1701 585
R3954 gnd.n5766 gnd.n5765 585
R3955 gnd.n5765 gnd.n5764 585
R3956 gnd.n1705 gnd.n1704 585
R3957 gnd.n5161 gnd.n1705 585
R3958 gnd.n5755 gnd.n5754 585
R3959 gnd.n5756 gnd.n5755 585
R3960 gnd.n1716 gnd.n1715 585
R3961 gnd.n5411 gnd.n1715 585
R3962 gnd.n5750 gnd.n5749 585
R3963 gnd.n5749 gnd.n5748 585
R3964 gnd.n1719 gnd.n1718 585
R3965 gnd.n5148 gnd.n1719 585
R3966 gnd.n5739 gnd.n5738 585
R3967 gnd.n5740 gnd.n5739 585
R3968 gnd.n1728 gnd.n1727 585
R3969 gnd.n5426 gnd.n1727 585
R3970 gnd.n5734 gnd.n5733 585
R3971 gnd.n5733 gnd.n5732 585
R3972 gnd.n1731 gnd.n1730 585
R3973 gnd.n5133 gnd.n1731 585
R3974 gnd.n5723 gnd.n5722 585
R3975 gnd.n5724 gnd.n5723 585
R3976 gnd.n1741 gnd.n1740 585
R3977 gnd.n5441 gnd.n1740 585
R3978 gnd.n5718 gnd.n5717 585
R3979 gnd.n5717 gnd.n5716 585
R3980 gnd.n1744 gnd.n1743 585
R3981 gnd.n5120 gnd.n1744 585
R3982 gnd.n5707 gnd.n5706 585
R3983 gnd.n5708 gnd.n5707 585
R3984 gnd.n1756 gnd.n1755 585
R3985 gnd.n5456 gnd.n1755 585
R3986 gnd.n5702 gnd.n5701 585
R3987 gnd.n5701 gnd.n5700 585
R3988 gnd.n1759 gnd.n1758 585
R3989 gnd.n5108 gnd.n1759 585
R3990 gnd.n5691 gnd.n5690 585
R3991 gnd.n5692 gnd.n5691 585
R3992 gnd.n1770 gnd.n1769 585
R3993 gnd.n5101 gnd.n1769 585
R3994 gnd.n5686 gnd.n5685 585
R3995 gnd.n5685 gnd.n5684 585
R3996 gnd.n1773 gnd.n1772 585
R3997 gnd.n5094 gnd.n1773 585
R3998 gnd.n5675 gnd.n5674 585
R3999 gnd.n5676 gnd.n5675 585
R4000 gnd.n1785 gnd.n1784 585
R4001 gnd.n5087 gnd.n1784 585
R4002 gnd.n5670 gnd.n5669 585
R4003 gnd.n5669 gnd.n5668 585
R4004 gnd.n1788 gnd.n1787 585
R4005 gnd.n5080 gnd.n1788 585
R4006 gnd.n5659 gnd.n5658 585
R4007 gnd.n5660 gnd.n5659 585
R4008 gnd.n1800 gnd.n1799 585
R4009 gnd.n5073 gnd.n1799 585
R4010 gnd.n5654 gnd.n5653 585
R4011 gnd.n5653 gnd.n5652 585
R4012 gnd.n1803 gnd.n1802 585
R4013 gnd.n5066 gnd.n1803 585
R4014 gnd.n5643 gnd.n5642 585
R4015 gnd.n5644 gnd.n5643 585
R4016 gnd.n1815 gnd.n1814 585
R4017 gnd.n5512 gnd.n1814 585
R4018 gnd.n5638 gnd.n5637 585
R4019 gnd.n5637 gnd.n5636 585
R4020 gnd.n1818 gnd.n1817 585
R4021 gnd.n5054 gnd.n1818 585
R4022 gnd.n5627 gnd.n5626 585
R4023 gnd.n5628 gnd.n5627 585
R4024 gnd.n1829 gnd.n1828 585
R4025 gnd.n5526 gnd.n1828 585
R4026 gnd.n5622 gnd.n5621 585
R4027 gnd.n5621 gnd.n5620 585
R4028 gnd.n1832 gnd.n1831 585
R4029 gnd.n5039 gnd.n1832 585
R4030 gnd.n5611 gnd.n5610 585
R4031 gnd.n5612 gnd.n5611 585
R4032 gnd.n1844 gnd.n1843 585
R4033 gnd.n5541 gnd.n1843 585
R4034 gnd.n5606 gnd.n5605 585
R4035 gnd.n5605 gnd.n5604 585
R4036 gnd.n1847 gnd.n1846 585
R4037 gnd.n5026 gnd.n1847 585
R4038 gnd.n5595 gnd.n5594 585
R4039 gnd.n5596 gnd.n5595 585
R4040 gnd.n1859 gnd.n1858 585
R4041 gnd.n5556 gnd.n1858 585
R4042 gnd.n5590 gnd.n5589 585
R4043 gnd.n5589 gnd.n5588 585
R4044 gnd.n1862 gnd.n1861 585
R4045 gnd.n1886 gnd.n1862 585
R4046 gnd.n5579 gnd.n5578 585
R4047 gnd.n5580 gnd.n5579 585
R4048 gnd.n1873 gnd.n1872 585
R4049 gnd.n5012 gnd.n1872 585
R4050 gnd.n5574 gnd.n5573 585
R4051 gnd.n5573 gnd.n5572 585
R4052 gnd.n1876 gnd.n1875 585
R4053 gnd.n5005 gnd.n1876 585
R4054 gnd.n4993 gnd.n1903 585
R4055 gnd.n1903 gnd.n1893 585
R4056 gnd.n4995 gnd.n4994 585
R4057 gnd.n4996 gnd.n4995 585
R4058 gnd.n1904 gnd.n1902 585
R4059 gnd.n1910 gnd.n1902 585
R4060 gnd.n4988 gnd.n4987 585
R4061 gnd.n4987 gnd.n4986 585
R4062 gnd.n1907 gnd.n1906 585
R4063 gnd.n1909 gnd.n1907 585
R4064 gnd.n4977 gnd.n4976 585
R4065 gnd.n4978 gnd.n4977 585
R4066 gnd.n1918 gnd.n1917 585
R4067 gnd.n1917 gnd.n1916 585
R4068 gnd.n4972 gnd.n4971 585
R4069 gnd.n4971 gnd.n4970 585
R4070 gnd.n1921 gnd.n1920 585
R4071 gnd.n1929 gnd.n1921 585
R4072 gnd.n4961 gnd.n4960 585
R4073 gnd.n4962 gnd.n4961 585
R4074 gnd.n1931 gnd.n1930 585
R4075 gnd.n1930 gnd.n1927 585
R4076 gnd.n4956 gnd.n4955 585
R4077 gnd.n4955 gnd.n4954 585
R4078 gnd.n1934 gnd.n1933 585
R4079 gnd.n1942 gnd.n1934 585
R4080 gnd.n4945 gnd.n4944 585
R4081 gnd.n4946 gnd.n4945 585
R4082 gnd.n1944 gnd.n1943 585
R4083 gnd.n1943 gnd.n1940 585
R4084 gnd.n4940 gnd.n4939 585
R4085 gnd.n4939 gnd.n4938 585
R4086 gnd.n1947 gnd.n1946 585
R4087 gnd.n1949 gnd.n1947 585
R4088 gnd.n4929 gnd.n4928 585
R4089 gnd.n4930 gnd.n4929 585
R4090 gnd.n1957 gnd.n1956 585
R4091 gnd.n1956 gnd.n1955 585
R4092 gnd.n4924 gnd.n4923 585
R4093 gnd.n4923 gnd.n4922 585
R4094 gnd.n1960 gnd.n1959 585
R4095 gnd.n1962 gnd.n1960 585
R4096 gnd.n4913 gnd.n4912 585
R4097 gnd.n4914 gnd.n4913 585
R4098 gnd.n1969 gnd.n1968 585
R4099 gnd.n1974 gnd.n1968 585
R4100 gnd.n4908 gnd.n4907 585
R4101 gnd.n4907 gnd.n4906 585
R4102 gnd.n1972 gnd.n1971 585
R4103 gnd.n1973 gnd.n1972 585
R4104 gnd.n4493 gnd.n4492 585
R4105 gnd.n4493 gnd.n1979 585
R4106 gnd.n4496 gnd.n4495 585
R4107 gnd.n4495 gnd.n4494 585
R4108 gnd.n4497 gnd.n4486 585
R4109 gnd.n4486 gnd.n2063 585
R4110 gnd.n4499 gnd.n4498 585
R4111 gnd.n4499 gnd.n2047 585
R4112 gnd.n4500 gnd.n4485 585
R4113 gnd.n4500 gnd.n1112 585
R4114 gnd.n4502 gnd.n4501 585
R4115 gnd.n4501 gnd.n1109 585
R4116 gnd.n4503 gnd.n4480 585
R4117 gnd.n4480 gnd.n2129 585
R4118 gnd.n4505 gnd.n4504 585
R4119 gnd.n4505 gnd.n1100 585
R4120 gnd.n4506 gnd.n4479 585
R4121 gnd.n4506 gnd.n1092 585
R4122 gnd.n4508 gnd.n4507 585
R4123 gnd.n4507 gnd.n1089 585
R4124 gnd.n4509 gnd.n2142 585
R4125 gnd.n2142 gnd.n1081 585
R4126 gnd.n4511 gnd.n4510 585
R4127 gnd.n4512 gnd.n4511 585
R4128 gnd.n2143 gnd.n2141 585
R4129 gnd.n2141 gnd.n1071 585
R4130 gnd.n4473 gnd.n4472 585
R4131 gnd.n4472 gnd.n1068 585
R4132 gnd.n4471 gnd.n2145 585
R4133 gnd.n4471 gnd.n1060 585
R4134 gnd.n4470 gnd.n4469 585
R4135 gnd.n4470 gnd.n1057 585
R4136 gnd.n2147 gnd.n2146 585
R4137 gnd.n2146 gnd.n1049 585
R4138 gnd.n4465 gnd.n4464 585
R4139 gnd.n4464 gnd.n4463 585
R4140 gnd.n2150 gnd.n2149 585
R4141 gnd.n2150 gnd.n1039 585
R4142 gnd.n4429 gnd.n4428 585
R4143 gnd.n4430 gnd.n4429 585
R4144 gnd.n2164 gnd.n2163 585
R4145 gnd.n2163 gnd.n1029 585
R4146 gnd.n4424 gnd.n4423 585
R4147 gnd.n4423 gnd.n1026 585
R4148 gnd.n4422 gnd.n2166 585
R4149 gnd.n4422 gnd.n1018 585
R4150 gnd.n4421 gnd.n4420 585
R4151 gnd.n4421 gnd.n1015 585
R4152 gnd.n2168 gnd.n2167 585
R4153 gnd.n2167 gnd.n1007 585
R4154 gnd.n4416 gnd.n4415 585
R4155 gnd.n4415 gnd.n4414 585
R4156 gnd.n2171 gnd.n2170 585
R4157 gnd.n2171 gnd.n997 585
R4158 gnd.n4380 gnd.n4379 585
R4159 gnd.n4381 gnd.n4380 585
R4160 gnd.n4373 gnd.n4372 585
R4161 gnd.n4372 gnd.n986 585
R4162 gnd.n4375 gnd.n4374 585
R4163 gnd.n4374 gnd.n983 585
R4164 gnd.n969 gnd.n968 585
R4165 gnd.n973 gnd.n969 585
R4166 gnd.n6405 gnd.n6404 585
R4167 gnd.n6404 gnd.n6403 585
R4168 gnd.n6166 gnd.n6165 585
R4169 gnd.n6165 gnd.n6164 585
R4170 gnd.n6167 gnd.n1243 585
R4171 gnd.n1245 gnd.n1243 585
R4172 gnd.n1619 gnd.n1241 585
R4173 gnd.n5873 gnd.n1619 585
R4174 gnd.n6171 gnd.n1240 585
R4175 gnd.n1618 gnd.n1240 585
R4176 gnd.n6172 gnd.n1239 585
R4177 gnd.n5862 gnd.n1239 585
R4178 gnd.n6173 gnd.n1238 585
R4179 gnd.n1626 gnd.n1238 585
R4180 gnd.n1633 gnd.n1236 585
R4181 gnd.n5852 gnd.n1633 585
R4182 gnd.n6177 gnd.n1235 585
R4183 gnd.n1640 gnd.n1235 585
R4184 gnd.n6178 gnd.n1234 585
R4185 gnd.n5844 gnd.n1234 585
R4186 gnd.n6179 gnd.n1233 585
R4187 gnd.n1639 gnd.n1233 585
R4188 gnd.n1647 gnd.n1231 585
R4189 gnd.n5836 gnd.n1647 585
R4190 gnd.n6183 gnd.n1230 585
R4191 gnd.n1646 gnd.n1230 585
R4192 gnd.n6184 gnd.n1229 585
R4193 gnd.n5828 gnd.n1229 585
R4194 gnd.n6185 gnd.n1228 585
R4195 gnd.n1653 gnd.n1228 585
R4196 gnd.n1660 gnd.n1226 585
R4197 gnd.n5820 gnd.n1660 585
R4198 gnd.n6189 gnd.n1225 585
R4199 gnd.n1659 gnd.n1225 585
R4200 gnd.n6190 gnd.n1224 585
R4201 gnd.n5812 gnd.n1224 585
R4202 gnd.n6191 gnd.n1223 585
R4203 gnd.n1666 gnd.n1223 585
R4204 gnd.n1673 gnd.n1221 585
R4205 gnd.n5804 gnd.n1673 585
R4206 gnd.n6195 gnd.n1220 585
R4207 gnd.n1672 gnd.n1220 585
R4208 gnd.n6196 gnd.n1219 585
R4209 gnd.n5796 gnd.n1219 585
R4210 gnd.n6197 gnd.n1218 585
R4211 gnd.n1686 gnd.n1218 585
R4212 gnd.n1685 gnd.n1216 585
R4213 gnd.n5788 gnd.n1685 585
R4214 gnd.n6201 gnd.n1215 585
R4215 gnd.n5183 gnd.n1215 585
R4216 gnd.n6202 gnd.n1214 585
R4217 gnd.n5780 gnd.n1214 585
R4218 gnd.n6203 gnd.n1213 585
R4219 gnd.n5179 gnd.n1213 585
R4220 gnd.n1700 gnd.n1211 585
R4221 gnd.n5772 gnd.n1700 585
R4222 gnd.n6207 gnd.n1210 585
R4223 gnd.n5396 gnd.n1210 585
R4224 gnd.n6208 gnd.n1209 585
R4225 gnd.n5764 gnd.n1209 585
R4226 gnd.n6209 gnd.n1208 585
R4227 gnd.n5161 gnd.n1208 585
R4228 gnd.n1714 gnd.n1206 585
R4229 gnd.n5756 gnd.n1714 585
R4230 gnd.n6213 gnd.n1205 585
R4231 gnd.n5411 gnd.n1205 585
R4232 gnd.n6214 gnd.n1204 585
R4233 gnd.n5748 gnd.n1204 585
R4234 gnd.n6215 gnd.n1203 585
R4235 gnd.n5148 gnd.n1203 585
R4236 gnd.n1726 gnd.n1201 585
R4237 gnd.n5740 gnd.n1726 585
R4238 gnd.n6219 gnd.n1200 585
R4239 gnd.n5426 gnd.n1200 585
R4240 gnd.n6220 gnd.n1199 585
R4241 gnd.n5732 gnd.n1199 585
R4242 gnd.n6221 gnd.n1198 585
R4243 gnd.n5133 gnd.n1198 585
R4244 gnd.n1738 gnd.n1196 585
R4245 gnd.n5724 gnd.n1738 585
R4246 gnd.n6225 gnd.n1195 585
R4247 gnd.n5441 gnd.n1195 585
R4248 gnd.n6226 gnd.n1194 585
R4249 gnd.n5716 gnd.n1194 585
R4250 gnd.n6227 gnd.n1193 585
R4251 gnd.n5120 gnd.n1193 585
R4252 gnd.n1752 gnd.n1191 585
R4253 gnd.n5708 gnd.n1752 585
R4254 gnd.n6231 gnd.n1190 585
R4255 gnd.n5456 gnd.n1190 585
R4256 gnd.n6232 gnd.n1189 585
R4257 gnd.n5700 gnd.n1189 585
R4258 gnd.n6233 gnd.n1188 585
R4259 gnd.n5108 gnd.n1188 585
R4260 gnd.n1767 gnd.n1186 585
R4261 gnd.n5692 gnd.n1767 585
R4262 gnd.n6237 gnd.n1185 585
R4263 gnd.n5101 gnd.n1185 585
R4264 gnd.n6238 gnd.n1184 585
R4265 gnd.n5684 gnd.n1184 585
R4266 gnd.n6239 gnd.n1183 585
R4267 gnd.n5094 gnd.n1183 585
R4268 gnd.n1782 gnd.n1181 585
R4269 gnd.n5676 gnd.n1782 585
R4270 gnd.n6243 gnd.n1180 585
R4271 gnd.n5087 gnd.n1180 585
R4272 gnd.n6244 gnd.n1179 585
R4273 gnd.n5668 gnd.n1179 585
R4274 gnd.n6245 gnd.n1178 585
R4275 gnd.n5080 gnd.n1178 585
R4276 gnd.n1797 gnd.n1176 585
R4277 gnd.n5660 gnd.n1797 585
R4278 gnd.n6249 gnd.n1175 585
R4279 gnd.n5073 gnd.n1175 585
R4280 gnd.n6250 gnd.n1174 585
R4281 gnd.n5652 gnd.n1174 585
R4282 gnd.n6251 gnd.n1173 585
R4283 gnd.n5066 gnd.n1173 585
R4284 gnd.n1812 gnd.n1171 585
R4285 gnd.n5644 gnd.n1812 585
R4286 gnd.n6255 gnd.n1170 585
R4287 gnd.n5512 gnd.n1170 585
R4288 gnd.n6256 gnd.n1169 585
R4289 gnd.n5636 gnd.n1169 585
R4290 gnd.n6257 gnd.n1168 585
R4291 gnd.n5054 gnd.n1168 585
R4292 gnd.n1826 gnd.n1166 585
R4293 gnd.n5628 gnd.n1826 585
R4294 gnd.n6261 gnd.n1165 585
R4295 gnd.n5526 gnd.n1165 585
R4296 gnd.n6262 gnd.n1164 585
R4297 gnd.n5620 gnd.n1164 585
R4298 gnd.n6263 gnd.n1163 585
R4299 gnd.n5039 gnd.n1163 585
R4300 gnd.n1841 gnd.n1161 585
R4301 gnd.n5612 gnd.n1841 585
R4302 gnd.n6267 gnd.n1160 585
R4303 gnd.n5541 gnd.n1160 585
R4304 gnd.n6268 gnd.n1159 585
R4305 gnd.n5604 gnd.n1159 585
R4306 gnd.n6269 gnd.n1158 585
R4307 gnd.n5026 gnd.n1158 585
R4308 gnd.n1856 gnd.n1156 585
R4309 gnd.n5596 gnd.n1856 585
R4310 gnd.n6273 gnd.n1155 585
R4311 gnd.n5556 gnd.n1155 585
R4312 gnd.n6274 gnd.n1154 585
R4313 gnd.n5588 gnd.n1154 585
R4314 gnd.n6275 gnd.n1153 585
R4315 gnd.n1886 gnd.n1153 585
R4316 gnd.n1870 gnd.n1151 585
R4317 gnd.n5580 gnd.n1870 585
R4318 gnd.n6279 gnd.n1150 585
R4319 gnd.n5012 gnd.n1150 585
R4320 gnd.n6280 gnd.n1149 585
R4321 gnd.n5572 gnd.n1149 585
R4322 gnd.n6281 gnd.n1148 585
R4323 gnd.n5005 gnd.n1148 585
R4324 gnd.n1892 gnd.n1146 585
R4325 gnd.n1893 gnd.n1892 585
R4326 gnd.n6285 gnd.n1145 585
R4327 gnd.n4996 gnd.n1145 585
R4328 gnd.n6286 gnd.n1144 585
R4329 gnd.n1910 gnd.n1144 585
R4330 gnd.n6287 gnd.n1143 585
R4331 gnd.n4986 gnd.n1143 585
R4332 gnd.n1908 gnd.n1141 585
R4333 gnd.n1909 gnd.n1908 585
R4334 gnd.n6291 gnd.n1140 585
R4335 gnd.n4978 gnd.n1140 585
R4336 gnd.n6292 gnd.n1139 585
R4337 gnd.n1916 gnd.n1139 585
R4338 gnd.n6293 gnd.n1138 585
R4339 gnd.n4970 gnd.n1138 585
R4340 gnd.n1928 gnd.n1136 585
R4341 gnd.n1929 gnd.n1928 585
R4342 gnd.n6297 gnd.n1135 585
R4343 gnd.n4962 gnd.n1135 585
R4344 gnd.n6298 gnd.n1134 585
R4345 gnd.n1927 gnd.n1134 585
R4346 gnd.n6299 gnd.n1133 585
R4347 gnd.n4954 gnd.n1133 585
R4348 gnd.n1941 gnd.n1131 585
R4349 gnd.n1942 gnd.n1941 585
R4350 gnd.n6303 gnd.n1130 585
R4351 gnd.n4946 gnd.n1130 585
R4352 gnd.n6304 gnd.n1129 585
R4353 gnd.n1940 gnd.n1129 585
R4354 gnd.n6305 gnd.n1128 585
R4355 gnd.n4938 gnd.n1128 585
R4356 gnd.n1948 gnd.n1126 585
R4357 gnd.n1949 gnd.n1948 585
R4358 gnd.n6309 gnd.n1125 585
R4359 gnd.n4930 gnd.n1125 585
R4360 gnd.n6310 gnd.n1124 585
R4361 gnd.n1955 gnd.n1124 585
R4362 gnd.n6311 gnd.n1123 585
R4363 gnd.n4922 gnd.n1123 585
R4364 gnd.n1961 gnd.n1121 585
R4365 gnd.n1962 gnd.n1961 585
R4366 gnd.n6315 gnd.n1120 585
R4367 gnd.n4914 gnd.n1120 585
R4368 gnd.n6316 gnd.n1119 585
R4369 gnd.n1974 gnd.n1119 585
R4370 gnd.n6317 gnd.n1118 585
R4371 gnd.n4906 gnd.n1118 585
R4372 gnd.n4895 gnd.n4894 585
R4373 gnd.n4893 gnd.n1993 585
R4374 gnd.n1995 gnd.n1992 585
R4375 gnd.n4897 gnd.n1992 585
R4376 gnd.n4886 gnd.n2003 585
R4377 gnd.n4885 gnd.n2004 585
R4378 gnd.n2006 gnd.n2005 585
R4379 gnd.n4878 gnd.n2012 585
R4380 gnd.n4877 gnd.n2013 585
R4381 gnd.n2020 gnd.n2014 585
R4382 gnd.n4870 gnd.n2021 585
R4383 gnd.n4869 gnd.n2022 585
R4384 gnd.n2024 gnd.n2023 585
R4385 gnd.n4862 gnd.n2030 585
R4386 gnd.n4861 gnd.n2031 585
R4387 gnd.n2040 gnd.n2032 585
R4388 gnd.n4854 gnd.n2041 585
R4389 gnd.n4853 gnd.n2042 585
R4390 gnd.n2044 gnd.n2043 585
R4391 gnd.n4561 gnd.n4536 585
R4392 gnd.n4560 gnd.n4537 585
R4393 gnd.n4559 gnd.n4538 585
R4394 gnd.n4540 gnd.n4539 585
R4395 gnd.n4555 gnd.n4542 585
R4396 gnd.n4554 gnd.n4543 585
R4397 gnd.n4553 gnd.n4544 585
R4398 gnd.n4550 gnd.n4549 585
R4399 gnd.n1978 gnd.n1977 585
R4400 gnd.n4900 gnd.n4899 585
R4401 gnd.n4901 gnd.n1975 585
R4402 gnd.n5877 gnd.n1247 585
R4403 gnd.n6164 gnd.n1247 585
R4404 gnd.n5876 gnd.n5875 585
R4405 gnd.n5875 gnd.n1245 585
R4406 gnd.n5874 gnd.n1616 585
R4407 gnd.n5874 gnd.n5873 585
R4408 gnd.n1629 gnd.n1617 585
R4409 gnd.n1618 gnd.n1617 585
R4410 gnd.n5861 gnd.n5860 585
R4411 gnd.n5862 gnd.n5861 585
R4412 gnd.n1628 gnd.n1627 585
R4413 gnd.n1627 gnd.n1626 585
R4414 gnd.n5854 gnd.n5853 585
R4415 gnd.n5853 gnd.n5852 585
R4416 gnd.n1632 gnd.n1631 585
R4417 gnd.n1640 gnd.n1632 585
R4418 gnd.n5843 gnd.n5842 585
R4419 gnd.n5844 gnd.n5843 585
R4420 gnd.n1642 gnd.n1641 585
R4421 gnd.n1641 gnd.n1639 585
R4422 gnd.n5838 gnd.n5837 585
R4423 gnd.n5837 gnd.n5836 585
R4424 gnd.n1645 gnd.n1644 585
R4425 gnd.n1646 gnd.n1645 585
R4426 gnd.n5827 gnd.n5826 585
R4427 gnd.n5828 gnd.n5827 585
R4428 gnd.n1655 gnd.n1654 585
R4429 gnd.n1654 gnd.n1653 585
R4430 gnd.n5822 gnd.n5821 585
R4431 gnd.n5821 gnd.n5820 585
R4432 gnd.n1658 gnd.n1657 585
R4433 gnd.n1659 gnd.n1658 585
R4434 gnd.n5811 gnd.n5810 585
R4435 gnd.n5812 gnd.n5811 585
R4436 gnd.n1668 gnd.n1667 585
R4437 gnd.n1667 gnd.n1666 585
R4438 gnd.n5806 gnd.n5805 585
R4439 gnd.n5805 gnd.n5804 585
R4440 gnd.n1671 gnd.n1670 585
R4441 gnd.n1672 gnd.n1671 585
R4442 gnd.n5795 gnd.n5794 585
R4443 gnd.n5796 gnd.n5795 585
R4444 gnd.n1680 gnd.n1679 585
R4445 gnd.n1686 gnd.n1679 585
R4446 gnd.n5790 gnd.n5789 585
R4447 gnd.n5789 gnd.n5788 585
R4448 gnd.n1683 gnd.n1682 585
R4449 gnd.n5183 gnd.n1683 585
R4450 gnd.n5779 gnd.n5778 585
R4451 gnd.n5780 gnd.n5779 585
R4452 gnd.n1695 gnd.n1694 585
R4453 gnd.n5179 gnd.n1694 585
R4454 gnd.n5774 gnd.n5773 585
R4455 gnd.n5773 gnd.n5772 585
R4456 gnd.n1698 gnd.n1697 585
R4457 gnd.n5396 gnd.n1698 585
R4458 gnd.n5763 gnd.n5762 585
R4459 gnd.n5764 gnd.n5763 585
R4460 gnd.n1709 gnd.n1708 585
R4461 gnd.n5161 gnd.n1708 585
R4462 gnd.n5758 gnd.n5757 585
R4463 gnd.n5757 gnd.n5756 585
R4464 gnd.n1712 gnd.n1711 585
R4465 gnd.n5411 gnd.n1712 585
R4466 gnd.n5747 gnd.n5746 585
R4467 gnd.n5748 gnd.n5747 585
R4468 gnd.n1722 gnd.n1721 585
R4469 gnd.n5148 gnd.n1721 585
R4470 gnd.n5742 gnd.n5741 585
R4471 gnd.n5741 gnd.n5740 585
R4472 gnd.n1725 gnd.n1724 585
R4473 gnd.n5426 gnd.n1725 585
R4474 gnd.n5731 gnd.n5730 585
R4475 gnd.n5732 gnd.n5731 585
R4476 gnd.n1734 gnd.n1733 585
R4477 gnd.n5133 gnd.n1733 585
R4478 gnd.n5726 gnd.n5725 585
R4479 gnd.n5725 gnd.n5724 585
R4480 gnd.n1737 gnd.n1736 585
R4481 gnd.n5441 gnd.n1737 585
R4482 gnd.n5715 gnd.n5714 585
R4483 gnd.n5716 gnd.n5715 585
R4484 gnd.n1747 gnd.n1746 585
R4485 gnd.n5120 gnd.n1746 585
R4486 gnd.n5710 gnd.n5709 585
R4487 gnd.n5709 gnd.n5708 585
R4488 gnd.n1750 gnd.n1749 585
R4489 gnd.n5456 gnd.n1750 585
R4490 gnd.n5699 gnd.n5698 585
R4491 gnd.n5700 gnd.n5699 585
R4492 gnd.n1762 gnd.n1761 585
R4493 gnd.n5108 gnd.n1761 585
R4494 gnd.n5694 gnd.n5693 585
R4495 gnd.n5693 gnd.n5692 585
R4496 gnd.n1765 gnd.n1764 585
R4497 gnd.n5101 gnd.n1765 585
R4498 gnd.n5683 gnd.n5682 585
R4499 gnd.n5684 gnd.n5683 585
R4500 gnd.n1777 gnd.n1776 585
R4501 gnd.n5094 gnd.n1776 585
R4502 gnd.n5678 gnd.n5677 585
R4503 gnd.n5677 gnd.n5676 585
R4504 gnd.n1780 gnd.n1779 585
R4505 gnd.n5087 gnd.n1780 585
R4506 gnd.n5667 gnd.n5666 585
R4507 gnd.n5668 gnd.n5667 585
R4508 gnd.n1792 gnd.n1791 585
R4509 gnd.n5080 gnd.n1791 585
R4510 gnd.n5662 gnd.n5661 585
R4511 gnd.n5661 gnd.n5660 585
R4512 gnd.n1795 gnd.n1794 585
R4513 gnd.n5073 gnd.n1795 585
R4514 gnd.n5651 gnd.n5650 585
R4515 gnd.n5652 gnd.n5651 585
R4516 gnd.n1807 gnd.n1806 585
R4517 gnd.n5066 gnd.n1806 585
R4518 gnd.n5646 gnd.n5645 585
R4519 gnd.n5645 gnd.n5644 585
R4520 gnd.n1810 gnd.n1809 585
R4521 gnd.n5512 gnd.n1810 585
R4522 gnd.n5635 gnd.n5634 585
R4523 gnd.n5636 gnd.n5635 585
R4524 gnd.n1822 gnd.n1821 585
R4525 gnd.n5054 gnd.n1821 585
R4526 gnd.n5630 gnd.n5629 585
R4527 gnd.n5629 gnd.n5628 585
R4528 gnd.n1825 gnd.n1824 585
R4529 gnd.n5526 gnd.n1825 585
R4530 gnd.n5619 gnd.n5618 585
R4531 gnd.n5620 gnd.n5619 585
R4532 gnd.n1836 gnd.n1835 585
R4533 gnd.n5039 gnd.n1835 585
R4534 gnd.n5614 gnd.n5613 585
R4535 gnd.n5613 gnd.n5612 585
R4536 gnd.n1839 gnd.n1838 585
R4537 gnd.n5541 gnd.n1839 585
R4538 gnd.n5603 gnd.n5602 585
R4539 gnd.n5604 gnd.n5603 585
R4540 gnd.n1851 gnd.n1850 585
R4541 gnd.n5026 gnd.n1850 585
R4542 gnd.n5598 gnd.n5597 585
R4543 gnd.n5597 gnd.n5596 585
R4544 gnd.n1854 gnd.n1853 585
R4545 gnd.n5556 gnd.n1854 585
R4546 gnd.n5587 gnd.n5586 585
R4547 gnd.n5588 gnd.n5587 585
R4548 gnd.n1865 gnd.n1864 585
R4549 gnd.n1886 gnd.n1864 585
R4550 gnd.n5582 gnd.n5581 585
R4551 gnd.n5581 gnd.n5580 585
R4552 gnd.n1868 gnd.n1867 585
R4553 gnd.n5012 gnd.n1868 585
R4554 gnd.n1897 gnd.n1879 585
R4555 gnd.n5572 gnd.n1879 585
R4556 gnd.n5004 gnd.n5003 585
R4557 gnd.n5005 gnd.n5004 585
R4558 gnd.n1896 gnd.n1895 585
R4559 gnd.n1895 gnd.n1893 585
R4560 gnd.n4998 gnd.n4997 585
R4561 gnd.n4997 gnd.n4996 585
R4562 gnd.n1900 gnd.n1899 585
R4563 gnd.n1910 gnd.n1900 585
R4564 gnd.n4985 gnd.n4984 585
R4565 gnd.n4986 gnd.n4985 585
R4566 gnd.n1912 gnd.n1911 585
R4567 gnd.n1911 gnd.n1909 585
R4568 gnd.n4980 gnd.n4979 585
R4569 gnd.n4979 gnd.n4978 585
R4570 gnd.n1915 gnd.n1914 585
R4571 gnd.n1916 gnd.n1915 585
R4572 gnd.n4969 gnd.n4968 585
R4573 gnd.n4970 gnd.n4969 585
R4574 gnd.n1923 gnd.n1922 585
R4575 gnd.n1929 gnd.n1922 585
R4576 gnd.n4964 gnd.n4963 585
R4577 gnd.n4963 gnd.n4962 585
R4578 gnd.n1926 gnd.n1925 585
R4579 gnd.n1927 gnd.n1926 585
R4580 gnd.n4953 gnd.n4952 585
R4581 gnd.n4954 gnd.n4953 585
R4582 gnd.n1936 gnd.n1935 585
R4583 gnd.n1942 gnd.n1935 585
R4584 gnd.n4948 gnd.n4947 585
R4585 gnd.n4947 gnd.n4946 585
R4586 gnd.n1939 gnd.n1938 585
R4587 gnd.n1940 gnd.n1939 585
R4588 gnd.n4937 gnd.n4936 585
R4589 gnd.n4938 gnd.n4937 585
R4590 gnd.n1951 gnd.n1950 585
R4591 gnd.n1950 gnd.n1949 585
R4592 gnd.n4932 gnd.n4931 585
R4593 gnd.n4931 gnd.n4930 585
R4594 gnd.n1954 gnd.n1953 585
R4595 gnd.n1955 gnd.n1954 585
R4596 gnd.n4921 gnd.n4920 585
R4597 gnd.n4922 gnd.n4921 585
R4598 gnd.n1964 gnd.n1963 585
R4599 gnd.n1963 gnd.n1962 585
R4600 gnd.n4916 gnd.n4915 585
R4601 gnd.n4915 gnd.n4914 585
R4602 gnd.n1967 gnd.n1966 585
R4603 gnd.n1974 gnd.n1967 585
R4604 gnd.n4905 gnd.n4904 585
R4605 gnd.n4906 gnd.n4905 585
R4606 gnd.n5884 gnd.n5883 585
R4607 gnd.n5883 gnd.n1248 585
R4608 gnd.n5885 gnd.n5882 585
R4609 gnd.n5880 gnd.n1614 585
R4610 gnd.n5889 gnd.n1613 585
R4611 gnd.n5893 gnd.n1611 585
R4612 gnd.n5894 gnd.n1610 585
R4613 gnd.n1608 gnd.n1606 585
R4614 gnd.n5898 gnd.n1605 585
R4615 gnd.n5899 gnd.n1603 585
R4616 gnd.n5900 gnd.n1602 585
R4617 gnd.n1600 gnd.n1480 585
R4618 gnd.n1599 gnd.n1598 585
R4619 gnd.n1588 gnd.n1482 585
R4620 gnd.n1590 gnd.n1589 585
R4621 gnd.n1586 gnd.n1492 585
R4622 gnd.n1585 gnd.n1584 585
R4623 gnd.n1572 gnd.n1494 585
R4624 gnd.n1574 gnd.n1573 585
R4625 gnd.n1570 gnd.n1498 585
R4626 gnd.n1569 gnd.n1568 585
R4627 gnd.n1553 gnd.n1500 585
R4628 gnd.n1555 gnd.n1554 585
R4629 gnd.n1551 gnd.n1505 585
R4630 gnd.n1550 gnd.n1549 585
R4631 gnd.n1534 gnd.n1507 585
R4632 gnd.n1536 gnd.n1535 585
R4633 gnd.n1532 gnd.n1512 585
R4634 gnd.n1531 gnd.n1530 585
R4635 gnd.n1514 gnd.n1244 585
R4636 gnd.n5372 gnd.n5184 473.281
R4637 gnd.n5255 gnd.n5182 473.281
R4638 gnd.n4751 gnd.n4749 473.281
R4639 gnd.n4747 gnd.n4642 473.281
R4640 gnd.n4621 gnd.t298 443.966
R4641 gnd.n5231 gnd.t251 443.966
R4642 gnd.n4677 gnd.t244 443.966
R4643 gnd.n5225 gnd.t288 443.966
R4644 gnd.n6582 gnd.n797 440.005
R4645 gnd.n4545 gnd.t265 371.625
R4646 gnd.n122 gnd.t279 371.625
R4647 gnd.n1486 gnd.t291 371.625
R4648 gnd.n2036 gnd.t315 371.625
R4649 gnd.n1308 gnd.t262 371.625
R4650 gnd.n1330 gnd.t240 371.625
R4651 gnd.n201 gnd.t308 371.625
R4652 gnd.n7628 gnd.t222 371.625
R4653 gnd.n4005 gnd.t324 371.625
R4654 gnd.n4037 gnd.t304 371.625
R4655 gnd.n3818 gnd.t321 371.625
R4656 gnd.n2125 gnd.t318 371.625
R4657 gnd.n2103 gnd.t236 371.625
R4658 gnd.n5890 gnd.t232 371.625
R4659 gnd.n2832 gnd.t311 323.425
R4660 gnd.n2377 gnd.t255 323.425
R4661 gnd.n3680 gnd.n3654 289.615
R4662 gnd.n3648 gnd.n3622 289.615
R4663 gnd.n3616 gnd.n3590 289.615
R4664 gnd.n3585 gnd.n3559 289.615
R4665 gnd.n3553 gnd.n3527 289.615
R4666 gnd.n3521 gnd.n3495 289.615
R4667 gnd.n3489 gnd.n3463 289.615
R4668 gnd.n3458 gnd.n3432 289.615
R4669 gnd.n2906 gnd.t294 279.217
R4670 gnd.n2403 gnd.t272 279.217
R4671 gnd.n4649 gnd.t231 260.649
R4672 gnd.n5196 gnd.t271 260.649
R4673 gnd.n4740 gnd.n1901 256.663
R4674 gnd.n4664 gnd.n1901 256.663
R4675 gnd.n4733 gnd.n1901 256.663
R4676 gnd.n4727 gnd.n1901 256.663
R4677 gnd.n4725 gnd.n1901 256.663
R4678 gnd.n4719 gnd.n1901 256.663
R4679 gnd.n4717 gnd.n1901 256.663
R4680 gnd.n4711 gnd.n1901 256.663
R4681 gnd.n4709 gnd.n1901 256.663
R4682 gnd.n4703 gnd.n1901 256.663
R4683 gnd.n4701 gnd.n1901 256.663
R4684 gnd.n4695 gnd.n1901 256.663
R4685 gnd.n4693 gnd.n1901 256.663
R4686 gnd.n4687 gnd.n1901 256.663
R4687 gnd.n4680 gnd.n1901 256.663
R4688 gnd.n4681 gnd.n1901 256.663
R4689 gnd.n4817 gnd.n4619 256.663
R4690 gnd.n4815 gnd.n1901 256.663
R4691 gnd.n4813 gnd.n1901 256.663
R4692 gnd.n4806 gnd.n1901 256.663
R4693 gnd.n4804 gnd.n1901 256.663
R4694 gnd.n4798 gnd.n1901 256.663
R4695 gnd.n4796 gnd.n1901 256.663
R4696 gnd.n4790 gnd.n1901 256.663
R4697 gnd.n4788 gnd.n1901 256.663
R4698 gnd.n4782 gnd.n1901 256.663
R4699 gnd.n4780 gnd.n1901 256.663
R4700 gnd.n4774 gnd.n1901 256.663
R4701 gnd.n4772 gnd.n1901 256.663
R4702 gnd.n4766 gnd.n1901 256.663
R4703 gnd.n4764 gnd.n1901 256.663
R4704 gnd.n4758 gnd.n1901 256.663
R4705 gnd.n4756 gnd.n1901 256.663
R4706 gnd.n4750 gnd.n1901 256.663
R4707 gnd.n5254 gnd.n1687 256.663
R4708 gnd.n5260 gnd.n1687 256.663
R4709 gnd.n5252 gnd.n1687 256.663
R4710 gnd.n5267 gnd.n1687 256.663
R4711 gnd.n5249 gnd.n1687 256.663
R4712 gnd.n5274 gnd.n1687 256.663
R4713 gnd.n5246 gnd.n1687 256.663
R4714 gnd.n5281 gnd.n1687 256.663
R4715 gnd.n5243 gnd.n1687 256.663
R4716 gnd.n5288 gnd.n1687 256.663
R4717 gnd.n5240 gnd.n1687 256.663
R4718 gnd.n5295 gnd.n1687 256.663
R4719 gnd.n5237 gnd.n1687 256.663
R4720 gnd.n5302 gnd.n1687 256.663
R4721 gnd.n5234 gnd.n1687 256.663
R4722 gnd.n5310 gnd.n1687 256.663
R4723 gnd.n5313 gnd.n1305 256.663
R4724 gnd.n5314 gnd.n1687 256.663
R4725 gnd.n5318 gnd.n1687 256.663
R4726 gnd.n5228 gnd.n1687 256.663
R4727 gnd.n5326 gnd.n1687 256.663
R4728 gnd.n5223 gnd.n1687 256.663
R4729 gnd.n5333 gnd.n1687 256.663
R4730 gnd.n5220 gnd.n1687 256.663
R4731 gnd.n5340 gnd.n1687 256.663
R4732 gnd.n5217 gnd.n1687 256.663
R4733 gnd.n5347 gnd.n1687 256.663
R4734 gnd.n5214 gnd.n1687 256.663
R4735 gnd.n5354 gnd.n1687 256.663
R4736 gnd.n5211 gnd.n1687 256.663
R4737 gnd.n5361 gnd.n1687 256.663
R4738 gnd.n5208 gnd.n1687 256.663
R4739 gnd.n5368 gnd.n1687 256.663
R4740 gnd.n5371 gnd.n1687 256.663
R4741 gnd.n3838 gnd.n3813 242.672
R4742 gnd.n3840 gnd.n3813 242.672
R4743 gnd.n3848 gnd.n3813 242.672
R4744 gnd.n3850 gnd.n3813 242.672
R4745 gnd.n3858 gnd.n3813 242.672
R4746 gnd.n3860 gnd.n3813 242.672
R4747 gnd.n3868 gnd.n3813 242.672
R4748 gnd.n3870 gnd.n3813 242.672
R4749 gnd.n3878 gnd.n3813 242.672
R4750 gnd.n4848 gnd.n4847 242.672
R4751 gnd.n4847 gnd.n2062 242.672
R4752 gnd.n4847 gnd.n2061 242.672
R4753 gnd.n4847 gnd.n2059 242.672
R4754 gnd.n4847 gnd.n2057 242.672
R4755 gnd.n4847 gnd.n2056 242.672
R4756 gnd.n4847 gnd.n2054 242.672
R4757 gnd.n4847 gnd.n2052 242.672
R4758 gnd.n4847 gnd.n2051 242.672
R4759 gnd.n6155 gnd.n1275 242.672
R4760 gnd.n6155 gnd.n1276 242.672
R4761 gnd.n6155 gnd.n1277 242.672
R4762 gnd.n6155 gnd.n1278 242.672
R4763 gnd.n6155 gnd.n1279 242.672
R4764 gnd.n6155 gnd.n1280 242.672
R4765 gnd.n6155 gnd.n1281 242.672
R4766 gnd.n6155 gnd.n1282 242.672
R4767 gnd.n6155 gnd.n1283 242.672
R4768 gnd.n128 gnd.n125 242.672
R4769 gnd.n7539 gnd.n128 242.672
R4770 gnd.n7535 gnd.n128 242.672
R4771 gnd.n7532 gnd.n128 242.672
R4772 gnd.n7527 gnd.n128 242.672
R4773 gnd.n7524 gnd.n128 242.672
R4774 gnd.n7519 gnd.n128 242.672
R4775 gnd.n7516 gnd.n128 242.672
R4776 gnd.n7511 gnd.n128 242.672
R4777 gnd.n2960 gnd.n2959 242.672
R4778 gnd.n2960 gnd.n2870 242.672
R4779 gnd.n2960 gnd.n2871 242.672
R4780 gnd.n2960 gnd.n2872 242.672
R4781 gnd.n2960 gnd.n2873 242.672
R4782 gnd.n2960 gnd.n2874 242.672
R4783 gnd.n2960 gnd.n2875 242.672
R4784 gnd.n2960 gnd.n2876 242.672
R4785 gnd.n2960 gnd.n2877 242.672
R4786 gnd.n2960 gnd.n2878 242.672
R4787 gnd.n2960 gnd.n2879 242.672
R4788 gnd.n2960 gnd.n2880 242.672
R4789 gnd.n2961 gnd.n2960 242.672
R4790 gnd.n3812 gnd.n2352 242.672
R4791 gnd.n3812 gnd.n2351 242.672
R4792 gnd.n3812 gnd.n2350 242.672
R4793 gnd.n3812 gnd.n2349 242.672
R4794 gnd.n3812 gnd.n2348 242.672
R4795 gnd.n3812 gnd.n2347 242.672
R4796 gnd.n3812 gnd.n2346 242.672
R4797 gnd.n3812 gnd.n2345 242.672
R4798 gnd.n3812 gnd.n2344 242.672
R4799 gnd.n3812 gnd.n2343 242.672
R4800 gnd.n3812 gnd.n2342 242.672
R4801 gnd.n3812 gnd.n2341 242.672
R4802 gnd.n3812 gnd.n2340 242.672
R4803 gnd.n3044 gnd.n3043 242.672
R4804 gnd.n3043 gnd.n2782 242.672
R4805 gnd.n3043 gnd.n2783 242.672
R4806 gnd.n3043 gnd.n2784 242.672
R4807 gnd.n3043 gnd.n2785 242.672
R4808 gnd.n3043 gnd.n2786 242.672
R4809 gnd.n3043 gnd.n2787 242.672
R4810 gnd.n3043 gnd.n2788 242.672
R4811 gnd.n3812 gnd.n2353 242.672
R4812 gnd.n3812 gnd.n2354 242.672
R4813 gnd.n3812 gnd.n2355 242.672
R4814 gnd.n3812 gnd.n2356 242.672
R4815 gnd.n3812 gnd.n2357 242.672
R4816 gnd.n3812 gnd.n2358 242.672
R4817 gnd.n3812 gnd.n2359 242.672
R4818 gnd.n3812 gnd.n2360 242.672
R4819 gnd.n4191 gnd.n3813 242.672
R4820 gnd.n3981 gnd.n3813 242.672
R4821 gnd.n4184 gnd.n3813 242.672
R4822 gnd.n4178 gnd.n3813 242.672
R4823 gnd.n4176 gnd.n3813 242.672
R4824 gnd.n4170 gnd.n3813 242.672
R4825 gnd.n4168 gnd.n3813 242.672
R4826 gnd.n4162 gnd.n3813 242.672
R4827 gnd.n4160 gnd.n3813 242.672
R4828 gnd.n4154 gnd.n3813 242.672
R4829 gnd.n4152 gnd.n3813 242.672
R4830 gnd.n4146 gnd.n3813 242.672
R4831 gnd.n4144 gnd.n3813 242.672
R4832 gnd.n4138 gnd.n3813 242.672
R4833 gnd.n4136 gnd.n3813 242.672
R4834 gnd.n4130 gnd.n3813 242.672
R4835 gnd.n4128 gnd.n3813 242.672
R4836 gnd.n4035 gnd.n3813 242.672
R4837 gnd.n4118 gnd.n3813 242.672
R4838 gnd.n4847 gnd.n2064 242.672
R4839 gnd.n4847 gnd.n2065 242.672
R4840 gnd.n4847 gnd.n2066 242.672
R4841 gnd.n4847 gnd.n2067 242.672
R4842 gnd.n4847 gnd.n2068 242.672
R4843 gnd.n4847 gnd.n2069 242.672
R4844 gnd.n4847 gnd.n2070 242.672
R4845 gnd.n4847 gnd.n2071 242.672
R4846 gnd.n4847 gnd.n2072 242.672
R4847 gnd.n4847 gnd.n2073 242.672
R4848 gnd.n4847 gnd.n2074 242.672
R4849 gnd.n4818 gnd.n2105 242.672
R4850 gnd.n4847 gnd.n2075 242.672
R4851 gnd.n4847 gnd.n2076 242.672
R4852 gnd.n4847 gnd.n2077 242.672
R4853 gnd.n4847 gnd.n2078 242.672
R4854 gnd.n4847 gnd.n2079 242.672
R4855 gnd.n4847 gnd.n2080 242.672
R4856 gnd.n4847 gnd.n2081 242.672
R4857 gnd.n4847 gnd.n4846 242.672
R4858 gnd.n6155 gnd.n6154 242.672
R4859 gnd.n6155 gnd.n1257 242.672
R4860 gnd.n6155 gnd.n1258 242.672
R4861 gnd.n6155 gnd.n1259 242.672
R4862 gnd.n6155 gnd.n1260 242.672
R4863 gnd.n6155 gnd.n1261 242.672
R4864 gnd.n6155 gnd.n1262 242.672
R4865 gnd.n6155 gnd.n1263 242.672
R4866 gnd.n6123 gnd.n1306 242.672
R4867 gnd.n6155 gnd.n1264 242.672
R4868 gnd.n6155 gnd.n1265 242.672
R4869 gnd.n6155 gnd.n1266 242.672
R4870 gnd.n6155 gnd.n1267 242.672
R4871 gnd.n6155 gnd.n1268 242.672
R4872 gnd.n6155 gnd.n1269 242.672
R4873 gnd.n6155 gnd.n1270 242.672
R4874 gnd.n6155 gnd.n1271 242.672
R4875 gnd.n6155 gnd.n1272 242.672
R4876 gnd.n6155 gnd.n1273 242.672
R4877 gnd.n6155 gnd.n1274 242.672
R4878 gnd.n198 gnd.n128 242.672
R4879 gnd.n7596 gnd.n128 242.672
R4880 gnd.n194 gnd.n128 242.672
R4881 gnd.n7603 gnd.n128 242.672
R4882 gnd.n187 gnd.n128 242.672
R4883 gnd.n7610 gnd.n128 242.672
R4884 gnd.n180 gnd.n128 242.672
R4885 gnd.n7617 gnd.n128 242.672
R4886 gnd.n173 gnd.n128 242.672
R4887 gnd.n7624 gnd.n128 242.672
R4888 gnd.n166 gnd.n128 242.672
R4889 gnd.n7634 gnd.n128 242.672
R4890 gnd.n159 gnd.n128 242.672
R4891 gnd.n7641 gnd.n128 242.672
R4892 gnd.n152 gnd.n128 242.672
R4893 gnd.n7648 gnd.n128 242.672
R4894 gnd.n145 gnd.n128 242.672
R4895 gnd.n7655 gnd.n128 242.672
R4896 gnd.n138 gnd.n128 242.672
R4897 gnd.n4897 gnd.n4896 242.672
R4898 gnd.n4897 gnd.n1980 242.672
R4899 gnd.n4897 gnd.n1981 242.672
R4900 gnd.n4897 gnd.n1982 242.672
R4901 gnd.n4897 gnd.n1983 242.672
R4902 gnd.n4897 gnd.n1984 242.672
R4903 gnd.n4897 gnd.n1985 242.672
R4904 gnd.n4897 gnd.n1986 242.672
R4905 gnd.n4897 gnd.n1987 242.672
R4906 gnd.n4897 gnd.n1988 242.672
R4907 gnd.n4897 gnd.n1989 242.672
R4908 gnd.n4897 gnd.n1990 242.672
R4909 gnd.n4897 gnd.n1991 242.672
R4910 gnd.n4898 gnd.n4897 242.672
R4911 gnd.n5881 gnd.n1248 242.672
R4912 gnd.n1612 gnd.n1248 242.672
R4913 gnd.n1609 gnd.n1248 242.672
R4914 gnd.n1604 gnd.n1248 242.672
R4915 gnd.n1601 gnd.n1248 242.672
R4916 gnd.n1481 gnd.n1248 242.672
R4917 gnd.n1587 gnd.n1248 242.672
R4918 gnd.n1493 gnd.n1248 242.672
R4919 gnd.n1571 gnd.n1248 242.672
R4920 gnd.n1499 gnd.n1248 242.672
R4921 gnd.n1552 gnd.n1248 242.672
R4922 gnd.n1506 gnd.n1248 242.672
R4923 gnd.n1533 gnd.n1248 242.672
R4924 gnd.n1513 gnd.n1248 242.672
R4925 gnd.n135 gnd.n131 240.244
R4926 gnd.n7657 gnd.n7656 240.244
R4927 gnd.n7654 gnd.n139 240.244
R4928 gnd.n7650 gnd.n7649 240.244
R4929 gnd.n7647 gnd.n146 240.244
R4930 gnd.n7643 gnd.n7642 240.244
R4931 gnd.n7640 gnd.n153 240.244
R4932 gnd.n7636 gnd.n7635 240.244
R4933 gnd.n7633 gnd.n160 240.244
R4934 gnd.n7626 gnd.n7625 240.244
R4935 gnd.n7623 gnd.n167 240.244
R4936 gnd.n7619 gnd.n7618 240.244
R4937 gnd.n7616 gnd.n174 240.244
R4938 gnd.n7612 gnd.n7611 240.244
R4939 gnd.n7609 gnd.n181 240.244
R4940 gnd.n7605 gnd.n7604 240.244
R4941 gnd.n7602 gnd.n188 240.244
R4942 gnd.n7598 gnd.n7597 240.244
R4943 gnd.n7595 gnd.n195 240.244
R4944 gnd.n6080 gnd.n1334 240.244
R4945 gnd.n1453 gnd.n1334 240.244
R4946 gnd.n1474 gnd.n1453 240.244
R4947 gnd.n1474 gnd.n1432 240.244
R4948 gnd.n1470 gnd.n1432 240.244
R4949 gnd.n1470 gnd.n1423 240.244
R4950 gnd.n1467 gnd.n1423 240.244
R4951 gnd.n1467 gnd.n1415 240.244
R4952 gnd.n1415 gnd.n1405 240.244
R4953 gnd.n1405 gnd.n1392 240.244
R4954 gnd.n5983 gnd.n1392 240.244
R4955 gnd.n5983 gnd.n1393 240.244
R4956 gnd.n1393 gnd.n1380 240.244
R4957 gnd.n1380 gnd.n1371 240.244
R4958 gnd.n5990 gnd.n1371 240.244
R4959 gnd.n5990 gnd.n1362 240.244
R4960 gnd.n5998 gnd.n1362 240.244
R4961 gnd.n5998 gnd.n400 240.244
R4962 gnd.n400 gnd.n389 240.244
R4963 gnd.n7246 gnd.n389 240.244
R4964 gnd.n7246 gnd.n385 240.244
R4965 gnd.n7258 gnd.n385 240.244
R4966 gnd.n7258 gnd.n368 240.244
R4967 gnd.n7254 gnd.n368 240.244
R4968 gnd.n7254 gnd.n355 240.244
R4969 gnd.n7291 gnd.n355 240.244
R4970 gnd.n7291 gnd.n351 240.244
R4971 gnd.n7304 gnd.n351 240.244
R4972 gnd.n7304 gnd.n313 240.244
R4973 gnd.n7300 gnd.n313 240.244
R4974 gnd.n7300 gnd.n343 240.244
R4975 gnd.n343 gnd.n339 240.244
R4976 gnd.n7321 gnd.n339 240.244
R4977 gnd.n7321 gnd.n335 240.244
R4978 gnd.n7392 gnd.n335 240.244
R4979 gnd.n7392 gnd.n328 240.244
R4980 gnd.n7388 gnd.n328 240.244
R4981 gnd.n7388 gnd.n300 240.244
R4982 gnd.n7385 gnd.n300 240.244
R4983 gnd.n7385 gnd.n291 240.244
R4984 gnd.n7382 gnd.n291 240.244
R4985 gnd.n7382 gnd.n283 240.244
R4986 gnd.n7379 gnd.n283 240.244
R4987 gnd.n7379 gnd.n276 240.244
R4988 gnd.n7376 gnd.n276 240.244
R4989 gnd.n7376 gnd.n270 240.244
R4990 gnd.n7373 gnd.n270 240.244
R4991 gnd.n7373 gnd.n261 240.244
R4992 gnd.n7370 gnd.n261 240.244
R4993 gnd.n7370 gnd.n253 240.244
R4994 gnd.n7367 gnd.n253 240.244
R4995 gnd.n7367 gnd.n245 240.244
R4996 gnd.n7364 gnd.n245 240.244
R4997 gnd.n7364 gnd.n239 240.244
R4998 gnd.n7361 gnd.n239 240.244
R4999 gnd.n7361 gnd.n230 240.244
R5000 gnd.n7358 gnd.n230 240.244
R5001 gnd.n7358 gnd.n223 240.244
R5002 gnd.n7355 gnd.n223 240.244
R5003 gnd.n7355 gnd.n214 240.244
R5004 gnd.n214 gnd.n205 240.244
R5005 gnd.n7586 gnd.n205 240.244
R5006 gnd.n7587 gnd.n7586 240.244
R5007 gnd.n7587 gnd.n127 240.244
R5008 gnd.n1287 gnd.n1286 240.244
R5009 gnd.n6148 gnd.n1286 240.244
R5010 gnd.n6146 gnd.n6145 240.244
R5011 gnd.n6142 gnd.n6141 240.244
R5012 gnd.n6138 gnd.n6137 240.244
R5013 gnd.n6134 gnd.n6133 240.244
R5014 gnd.n6130 gnd.n6129 240.244
R5015 gnd.n6126 gnd.n6125 240.244
R5016 gnd.n6121 gnd.n6120 240.244
R5017 gnd.n6117 gnd.n6116 240.244
R5018 gnd.n6113 gnd.n6112 240.244
R5019 gnd.n6109 gnd.n6108 240.244
R5020 gnd.n6105 gnd.n6104 240.244
R5021 gnd.n6101 gnd.n6100 240.244
R5022 gnd.n6097 gnd.n6096 240.244
R5023 gnd.n6093 gnd.n6092 240.244
R5024 gnd.n6089 gnd.n6088 240.244
R5025 gnd.n1329 gnd.n1328 240.244
R5026 gnd.n5913 gnd.n1288 240.244
R5027 gnd.n5913 gnd.n5906 240.244
R5028 gnd.n5906 gnd.n1430 240.244
R5029 gnd.n5936 gnd.n1430 240.244
R5030 gnd.n5936 gnd.n1425 240.244
R5031 gnd.n5944 gnd.n1425 240.244
R5032 gnd.n5944 gnd.n1426 240.244
R5033 gnd.n1426 gnd.n1403 240.244
R5034 gnd.n5973 gnd.n1403 240.244
R5035 gnd.n5973 gnd.n1397 240.244
R5036 gnd.n5981 gnd.n1397 240.244
R5037 gnd.n5981 gnd.n1399 240.244
R5038 gnd.n1399 gnd.n1369 240.244
R5039 gnd.n6043 gnd.n1369 240.244
R5040 gnd.n6043 gnd.n1365 240.244
R5041 gnd.n6049 gnd.n1365 240.244
R5042 gnd.n6049 gnd.n398 240.244
R5043 gnd.n7236 gnd.n398 240.244
R5044 gnd.n7236 gnd.n393 240.244
R5045 gnd.n7244 gnd.n393 240.244
R5046 gnd.n7244 gnd.n394 240.244
R5047 gnd.n394 gnd.n365 240.244
R5048 gnd.n7282 gnd.n365 240.244
R5049 gnd.n7282 gnd.n366 240.244
R5050 gnd.n366 gnd.n360 240.244
R5051 gnd.n7289 gnd.n360 240.244
R5052 gnd.n7289 gnd.n361 240.244
R5053 gnd.n361 gnd.n310 240.244
R5054 gnd.n7413 gnd.n310 240.244
R5055 gnd.n7413 gnd.n311 240.244
R5056 gnd.n7315 gnd.n311 240.244
R5057 gnd.n7316 gnd.n7315 240.244
R5058 gnd.n7319 gnd.n7316 240.244
R5059 gnd.n7319 gnd.n330 240.244
R5060 gnd.n7394 gnd.n330 240.244
R5061 gnd.n7396 gnd.n7394 240.244
R5062 gnd.n7396 gnd.n301 240.244
R5063 gnd.n7420 gnd.n301 240.244
R5064 gnd.n7420 gnd.n289 240.244
R5065 gnd.n7430 gnd.n289 240.244
R5066 gnd.n7430 gnd.n285 240.244
R5067 gnd.n7436 gnd.n285 240.244
R5068 gnd.n7436 gnd.n275 240.244
R5069 gnd.n7446 gnd.n275 240.244
R5070 gnd.n7446 gnd.n271 240.244
R5071 gnd.n7452 gnd.n271 240.244
R5072 gnd.n7452 gnd.n259 240.244
R5073 gnd.n7462 gnd.n259 240.244
R5074 gnd.n7462 gnd.n255 240.244
R5075 gnd.n7468 gnd.n255 240.244
R5076 gnd.n7468 gnd.n244 240.244
R5077 gnd.n7478 gnd.n244 240.244
R5078 gnd.n7478 gnd.n240 240.244
R5079 gnd.n7484 gnd.n240 240.244
R5080 gnd.n7484 gnd.n228 240.244
R5081 gnd.n7494 gnd.n228 240.244
R5082 gnd.n7494 gnd.n224 240.244
R5083 gnd.n7500 gnd.n224 240.244
R5084 gnd.n7500 gnd.n212 240.244
R5085 gnd.n7578 gnd.n212 240.244
R5086 gnd.n7578 gnd.n208 240.244
R5087 gnd.n7584 gnd.n208 240.244
R5088 gnd.n7584 gnd.n130 240.244
R5089 gnd.n7664 gnd.n130 240.244
R5090 gnd.n2082 gnd.n1108 240.244
R5091 gnd.n4845 gnd.n2083 240.244
R5092 gnd.n4841 gnd.n4840 240.244
R5093 gnd.n4837 gnd.n4836 240.244
R5094 gnd.n4833 gnd.n4832 240.244
R5095 gnd.n4829 gnd.n4828 240.244
R5096 gnd.n4825 gnd.n4824 240.244
R5097 gnd.n4821 gnd.n4820 240.244
R5098 gnd.n4612 gnd.n4611 240.244
R5099 gnd.n4609 gnd.n4608 240.244
R5100 gnd.n4605 gnd.n4604 240.244
R5101 gnd.n4601 gnd.n4600 240.244
R5102 gnd.n4597 gnd.n4596 240.244
R5103 gnd.n4593 gnd.n4592 240.244
R5104 gnd.n4589 gnd.n4588 240.244
R5105 gnd.n4585 gnd.n4584 240.244
R5106 gnd.n4581 gnd.n4580 240.244
R5107 gnd.n4577 gnd.n4576 240.244
R5108 gnd.n4041 gnd.n3814 240.244
R5109 gnd.n4041 gnd.n2333 240.244
R5110 gnd.n4111 gnd.n2333 240.244
R5111 gnd.n4111 gnd.n2326 240.244
R5112 gnd.n4108 gnd.n2326 240.244
R5113 gnd.n4108 gnd.n2318 240.244
R5114 gnd.n4105 gnd.n2318 240.244
R5115 gnd.n4105 gnd.n2309 240.244
R5116 gnd.n4102 gnd.n2309 240.244
R5117 gnd.n4102 gnd.n2301 240.244
R5118 gnd.n4099 gnd.n2301 240.244
R5119 gnd.n4099 gnd.n2294 240.244
R5120 gnd.n4096 gnd.n2294 240.244
R5121 gnd.n4096 gnd.n2286 240.244
R5122 gnd.n4093 gnd.n2286 240.244
R5123 gnd.n4093 gnd.n2277 240.244
R5124 gnd.n4090 gnd.n2277 240.244
R5125 gnd.n4090 gnd.n2269 240.244
R5126 gnd.n4087 gnd.n2269 240.244
R5127 gnd.n4087 gnd.n2262 240.244
R5128 gnd.n4084 gnd.n2262 240.244
R5129 gnd.n4084 gnd.n2254 240.244
R5130 gnd.n4081 gnd.n2254 240.244
R5131 gnd.n4081 gnd.n2245 240.244
R5132 gnd.n4078 gnd.n2245 240.244
R5133 gnd.n4078 gnd.n2237 240.244
R5134 gnd.n4075 gnd.n2237 240.244
R5135 gnd.n4075 gnd.n2231 240.244
R5136 gnd.n4072 gnd.n2231 240.244
R5137 gnd.n4072 gnd.n2222 240.244
R5138 gnd.n2222 gnd.n2212 240.244
R5139 gnd.n4330 gnd.n2212 240.244
R5140 gnd.n4330 gnd.n2213 240.244
R5141 gnd.n2213 gnd.n2195 240.244
R5142 gnd.n2195 gnd.n2189 240.244
R5143 gnd.n4356 gnd.n2189 240.244
R5144 gnd.n4357 gnd.n4356 240.244
R5145 gnd.n4357 gnd.n971 240.244
R5146 gnd.n4363 gnd.n971 240.244
R5147 gnd.n4363 gnd.n984 240.244
R5148 gnd.n4383 gnd.n984 240.244
R5149 gnd.n4383 gnd.n995 240.244
R5150 gnd.n2172 gnd.n995 240.244
R5151 gnd.n2172 gnd.n1005 240.244
R5152 gnd.n4391 gnd.n1005 240.244
R5153 gnd.n4391 gnd.n1016 240.244
R5154 gnd.n4397 gnd.n1016 240.244
R5155 gnd.n4397 gnd.n1027 240.244
R5156 gnd.n4432 gnd.n1027 240.244
R5157 gnd.n4432 gnd.n1037 240.244
R5158 gnd.n2151 gnd.n1037 240.244
R5159 gnd.n2151 gnd.n1047 240.244
R5160 gnd.n4440 gnd.n1047 240.244
R5161 gnd.n4440 gnd.n1058 240.244
R5162 gnd.n4450 gnd.n1058 240.244
R5163 gnd.n4450 gnd.n1069 240.244
R5164 gnd.n2140 gnd.n1069 240.244
R5165 gnd.n2140 gnd.n1079 240.244
R5166 gnd.n4522 gnd.n1079 240.244
R5167 gnd.n4522 gnd.n1090 240.244
R5168 gnd.n4529 gnd.n1090 240.244
R5169 gnd.n4529 gnd.n1101 240.244
R5170 gnd.n4569 gnd.n1101 240.244
R5171 gnd.n4569 gnd.n1110 240.244
R5172 gnd.n4192 gnd.n4190 240.244
R5173 gnd.n4190 gnd.n4189 240.244
R5174 gnd.n4186 gnd.n4185 240.244
R5175 gnd.n4183 gnd.n3986 240.244
R5176 gnd.n4179 gnd.n4177 240.244
R5177 gnd.n4175 gnd.n3992 240.244
R5178 gnd.n4171 gnd.n4169 240.244
R5179 gnd.n4167 gnd.n3998 240.244
R5180 gnd.n4163 gnd.n4161 240.244
R5181 gnd.n4159 gnd.n4004 240.244
R5182 gnd.n4155 gnd.n4153 240.244
R5183 gnd.n4151 gnd.n4013 240.244
R5184 gnd.n4147 gnd.n4145 240.244
R5185 gnd.n4143 gnd.n4019 240.244
R5186 gnd.n4139 gnd.n4137 240.244
R5187 gnd.n4135 gnd.n4025 240.244
R5188 gnd.n4131 gnd.n4129 240.244
R5189 gnd.n4127 gnd.n4031 240.244
R5190 gnd.n4117 gnd.n4036 240.244
R5191 gnd.n4198 gnd.n2332 240.244
R5192 gnd.n4208 gnd.n2332 240.244
R5193 gnd.n4208 gnd.n2328 240.244
R5194 gnd.n4214 gnd.n2328 240.244
R5195 gnd.n4214 gnd.n2316 240.244
R5196 gnd.n4224 gnd.n2316 240.244
R5197 gnd.n4224 gnd.n2312 240.244
R5198 gnd.n4230 gnd.n2312 240.244
R5199 gnd.n4230 gnd.n2300 240.244
R5200 gnd.n4240 gnd.n2300 240.244
R5201 gnd.n4240 gnd.n2296 240.244
R5202 gnd.n4246 gnd.n2296 240.244
R5203 gnd.n4246 gnd.n2284 240.244
R5204 gnd.n4256 gnd.n2284 240.244
R5205 gnd.n4256 gnd.n2280 240.244
R5206 gnd.n4262 gnd.n2280 240.244
R5207 gnd.n4262 gnd.n2268 240.244
R5208 gnd.n4272 gnd.n2268 240.244
R5209 gnd.n4272 gnd.n2264 240.244
R5210 gnd.n4278 gnd.n2264 240.244
R5211 gnd.n4278 gnd.n2252 240.244
R5212 gnd.n4288 gnd.n2252 240.244
R5213 gnd.n4288 gnd.n2248 240.244
R5214 gnd.n4295 gnd.n2248 240.244
R5215 gnd.n4295 gnd.n2236 240.244
R5216 gnd.n4305 gnd.n2236 240.244
R5217 gnd.n4305 gnd.n2233 240.244
R5218 gnd.n4311 gnd.n2233 240.244
R5219 gnd.n4311 gnd.n2220 240.244
R5220 gnd.n4322 gnd.n2220 240.244
R5221 gnd.n4322 gnd.n2218 240.244
R5222 gnd.n4328 gnd.n2218 240.244
R5223 gnd.n4328 gnd.n2194 240.244
R5224 gnd.n4349 gnd.n2194 240.244
R5225 gnd.n4349 gnd.n2192 240.244
R5226 gnd.n4354 gnd.n2192 240.244
R5227 gnd.n4354 gnd.n975 240.244
R5228 gnd.n6401 gnd.n975 240.244
R5229 gnd.n6401 gnd.n976 240.244
R5230 gnd.n6397 gnd.n976 240.244
R5231 gnd.n6397 gnd.n982 240.244
R5232 gnd.n6389 gnd.n982 240.244
R5233 gnd.n6389 gnd.n998 240.244
R5234 gnd.n6385 gnd.n998 240.244
R5235 gnd.n6385 gnd.n1004 240.244
R5236 gnd.n6377 gnd.n1004 240.244
R5237 gnd.n6377 gnd.n1019 240.244
R5238 gnd.n6373 gnd.n1019 240.244
R5239 gnd.n6373 gnd.n1025 240.244
R5240 gnd.n6365 gnd.n1025 240.244
R5241 gnd.n6365 gnd.n1040 240.244
R5242 gnd.n6361 gnd.n1040 240.244
R5243 gnd.n6361 gnd.n1046 240.244
R5244 gnd.n6353 gnd.n1046 240.244
R5245 gnd.n6353 gnd.n1061 240.244
R5246 gnd.n6349 gnd.n1061 240.244
R5247 gnd.n6349 gnd.n1067 240.244
R5248 gnd.n6341 gnd.n1067 240.244
R5249 gnd.n6341 gnd.n1082 240.244
R5250 gnd.n6337 gnd.n1082 240.244
R5251 gnd.n6337 gnd.n1088 240.244
R5252 gnd.n6329 gnd.n1088 240.244
R5253 gnd.n6329 gnd.n1103 240.244
R5254 gnd.n6325 gnd.n1103 240.244
R5255 gnd.n3811 gnd.n2362 240.244
R5256 gnd.n3804 gnd.n3803 240.244
R5257 gnd.n3801 gnd.n3800 240.244
R5258 gnd.n3797 gnd.n3796 240.244
R5259 gnd.n3793 gnd.n3792 240.244
R5260 gnd.n3789 gnd.n3788 240.244
R5261 gnd.n3785 gnd.n3784 240.244
R5262 gnd.n3781 gnd.n3780 240.244
R5263 gnd.n3055 gnd.n2767 240.244
R5264 gnd.n3065 gnd.n2767 240.244
R5265 gnd.n3065 gnd.n2758 240.244
R5266 gnd.n2758 gnd.n2747 240.244
R5267 gnd.n3086 gnd.n2747 240.244
R5268 gnd.n3086 gnd.n2741 240.244
R5269 gnd.n3096 gnd.n2741 240.244
R5270 gnd.n3096 gnd.n2730 240.244
R5271 gnd.n2730 gnd.n2722 240.244
R5272 gnd.n3114 gnd.n2722 240.244
R5273 gnd.n3115 gnd.n3114 240.244
R5274 gnd.n3115 gnd.n2707 240.244
R5275 gnd.n3117 gnd.n2707 240.244
R5276 gnd.n3117 gnd.n2693 240.244
R5277 gnd.n3159 gnd.n2693 240.244
R5278 gnd.n3160 gnd.n3159 240.244
R5279 gnd.n3163 gnd.n3160 240.244
R5280 gnd.n3163 gnd.n2648 240.244
R5281 gnd.n2688 gnd.n2648 240.244
R5282 gnd.n2688 gnd.n2658 240.244
R5283 gnd.n3173 gnd.n2658 240.244
R5284 gnd.n3173 gnd.n2679 240.244
R5285 gnd.n3183 gnd.n2679 240.244
R5286 gnd.n3183 gnd.n2565 240.244
R5287 gnd.n3228 gnd.n2565 240.244
R5288 gnd.n3228 gnd.n2551 240.244
R5289 gnd.n3250 gnd.n2551 240.244
R5290 gnd.n3251 gnd.n3250 240.244
R5291 gnd.n3251 gnd.n2538 240.244
R5292 gnd.n2538 gnd.n2527 240.244
R5293 gnd.n3282 gnd.n2527 240.244
R5294 gnd.n3283 gnd.n3282 240.244
R5295 gnd.n3284 gnd.n3283 240.244
R5296 gnd.n3284 gnd.n2512 240.244
R5297 gnd.n2512 gnd.n2511 240.244
R5298 gnd.n2511 gnd.n2496 240.244
R5299 gnd.n3335 gnd.n2496 240.244
R5300 gnd.n3336 gnd.n3335 240.244
R5301 gnd.n3336 gnd.n2483 240.244
R5302 gnd.n2483 gnd.n2472 240.244
R5303 gnd.n3367 gnd.n2472 240.244
R5304 gnd.n3368 gnd.n3367 240.244
R5305 gnd.n3369 gnd.n3368 240.244
R5306 gnd.n3369 gnd.n2456 240.244
R5307 gnd.n2456 gnd.n2455 240.244
R5308 gnd.n2455 gnd.n2442 240.244
R5309 gnd.n3424 gnd.n2442 240.244
R5310 gnd.n3425 gnd.n3424 240.244
R5311 gnd.n3425 gnd.n2429 240.244
R5312 gnd.n2429 gnd.n2419 240.244
R5313 gnd.n3712 gnd.n2419 240.244
R5314 gnd.n3715 gnd.n3712 240.244
R5315 gnd.n3715 gnd.n3714 240.244
R5316 gnd.n3045 gnd.n2780 240.244
R5317 gnd.n2801 gnd.n2780 240.244
R5318 gnd.n2804 gnd.n2803 240.244
R5319 gnd.n2811 gnd.n2810 240.244
R5320 gnd.n2814 gnd.n2813 240.244
R5321 gnd.n2821 gnd.n2820 240.244
R5322 gnd.n2824 gnd.n2823 240.244
R5323 gnd.n2831 gnd.n2830 240.244
R5324 gnd.n3053 gnd.n2777 240.244
R5325 gnd.n2777 gnd.n2756 240.244
R5326 gnd.n3076 gnd.n2756 240.244
R5327 gnd.n3076 gnd.n2750 240.244
R5328 gnd.n3084 gnd.n2750 240.244
R5329 gnd.n3084 gnd.n2752 240.244
R5330 gnd.n2752 gnd.n2728 240.244
R5331 gnd.n3106 gnd.n2728 240.244
R5332 gnd.n3106 gnd.n2724 240.244
R5333 gnd.n3112 gnd.n2724 240.244
R5334 gnd.n3112 gnd.n2706 240.244
R5335 gnd.n3137 gnd.n2706 240.244
R5336 gnd.n3137 gnd.n2701 240.244
R5337 gnd.n3149 gnd.n2701 240.244
R5338 gnd.n3149 gnd.n2702 240.244
R5339 gnd.n3145 gnd.n2702 240.244
R5340 gnd.n3145 gnd.n2650 240.244
R5341 gnd.n3197 gnd.n2650 240.244
R5342 gnd.n3197 gnd.n2651 240.244
R5343 gnd.n3193 gnd.n2651 240.244
R5344 gnd.n3193 gnd.n2657 240.244
R5345 gnd.n2677 gnd.n2657 240.244
R5346 gnd.n2677 gnd.n2563 240.244
R5347 gnd.n3232 gnd.n2563 240.244
R5348 gnd.n3232 gnd.n2558 240.244
R5349 gnd.n3240 gnd.n2558 240.244
R5350 gnd.n3240 gnd.n2559 240.244
R5351 gnd.n2559 gnd.n2536 240.244
R5352 gnd.n3272 gnd.n2536 240.244
R5353 gnd.n3272 gnd.n2531 240.244
R5354 gnd.n3280 gnd.n2531 240.244
R5355 gnd.n3280 gnd.n2532 240.244
R5356 gnd.n2532 gnd.n2509 240.244
R5357 gnd.n3317 gnd.n2509 240.244
R5358 gnd.n3317 gnd.n2504 240.244
R5359 gnd.n3325 gnd.n2504 240.244
R5360 gnd.n3325 gnd.n2505 240.244
R5361 gnd.n2505 gnd.n2481 240.244
R5362 gnd.n3357 gnd.n2481 240.244
R5363 gnd.n3357 gnd.n2476 240.244
R5364 gnd.n3365 gnd.n2476 240.244
R5365 gnd.n3365 gnd.n2477 240.244
R5366 gnd.n2477 gnd.n2454 240.244
R5367 gnd.n3406 gnd.n2454 240.244
R5368 gnd.n3406 gnd.n2449 240.244
R5369 gnd.n3414 gnd.n2449 240.244
R5370 gnd.n3414 gnd.n2450 240.244
R5371 gnd.n2450 gnd.n2427 240.244
R5372 gnd.n3700 gnd.n2427 240.244
R5373 gnd.n3700 gnd.n2422 240.244
R5374 gnd.n3710 gnd.n2422 240.244
R5375 gnd.n3710 gnd.n2423 240.244
R5376 gnd.n2423 gnd.n2361 240.244
R5377 gnd.n2381 gnd.n2339 240.244
R5378 gnd.n3771 gnd.n3770 240.244
R5379 gnd.n3767 gnd.n3766 240.244
R5380 gnd.n3763 gnd.n3762 240.244
R5381 gnd.n3759 gnd.n3758 240.244
R5382 gnd.n3755 gnd.n3754 240.244
R5383 gnd.n3751 gnd.n3750 240.244
R5384 gnd.n3747 gnd.n3746 240.244
R5385 gnd.n3743 gnd.n3742 240.244
R5386 gnd.n3739 gnd.n3738 240.244
R5387 gnd.n3735 gnd.n3734 240.244
R5388 gnd.n3731 gnd.n3730 240.244
R5389 gnd.n3727 gnd.n3726 240.244
R5390 gnd.n2968 gnd.n2865 240.244
R5391 gnd.n2968 gnd.n2858 240.244
R5392 gnd.n2979 gnd.n2858 240.244
R5393 gnd.n2979 gnd.n2854 240.244
R5394 gnd.n2985 gnd.n2854 240.244
R5395 gnd.n2985 gnd.n2846 240.244
R5396 gnd.n2995 gnd.n2846 240.244
R5397 gnd.n2995 gnd.n2841 240.244
R5398 gnd.n3031 gnd.n2841 240.244
R5399 gnd.n3031 gnd.n2842 240.244
R5400 gnd.n2842 gnd.n2789 240.244
R5401 gnd.n3026 gnd.n2789 240.244
R5402 gnd.n3026 gnd.n3025 240.244
R5403 gnd.n3025 gnd.n2768 240.244
R5404 gnd.n3021 gnd.n2768 240.244
R5405 gnd.n3021 gnd.n2759 240.244
R5406 gnd.n3018 gnd.n2759 240.244
R5407 gnd.n3018 gnd.n3017 240.244
R5408 gnd.n3017 gnd.n2742 240.244
R5409 gnd.n3013 gnd.n2742 240.244
R5410 gnd.n3013 gnd.n2731 240.244
R5411 gnd.n2731 gnd.n2712 240.244
R5412 gnd.n3126 gnd.n2712 240.244
R5413 gnd.n3126 gnd.n2708 240.244
R5414 gnd.n3134 gnd.n2708 240.244
R5415 gnd.n3134 gnd.n2699 240.244
R5416 gnd.n2699 gnd.n2635 240.244
R5417 gnd.n3206 gnd.n2635 240.244
R5418 gnd.n3206 gnd.n2636 240.244
R5419 gnd.n2647 gnd.n2636 240.244
R5420 gnd.n2682 gnd.n2647 240.244
R5421 gnd.n2685 gnd.n2682 240.244
R5422 gnd.n2685 gnd.n2659 240.244
R5423 gnd.n2672 gnd.n2659 240.244
R5424 gnd.n2672 gnd.n2669 240.244
R5425 gnd.n2669 gnd.n2566 240.244
R5426 gnd.n3227 gnd.n2566 240.244
R5427 gnd.n3227 gnd.n2556 240.244
R5428 gnd.n3223 gnd.n2556 240.244
R5429 gnd.n3223 gnd.n2550 240.244
R5430 gnd.n3220 gnd.n2550 240.244
R5431 gnd.n3220 gnd.n2539 240.244
R5432 gnd.n3217 gnd.n2539 240.244
R5433 gnd.n3217 gnd.n2517 240.244
R5434 gnd.n3293 gnd.n2517 240.244
R5435 gnd.n3293 gnd.n2513 240.244
R5436 gnd.n3314 gnd.n2513 240.244
R5437 gnd.n3314 gnd.n2502 240.244
R5438 gnd.n3310 gnd.n2502 240.244
R5439 gnd.n3310 gnd.n2495 240.244
R5440 gnd.n3307 gnd.n2495 240.244
R5441 gnd.n3307 gnd.n2484 240.244
R5442 gnd.n3304 gnd.n2484 240.244
R5443 gnd.n3304 gnd.n2461 240.244
R5444 gnd.n3378 gnd.n2461 240.244
R5445 gnd.n3378 gnd.n2457 240.244
R5446 gnd.n3403 gnd.n2457 240.244
R5447 gnd.n3403 gnd.n2448 240.244
R5448 gnd.n3399 gnd.n2448 240.244
R5449 gnd.n3399 gnd.n2441 240.244
R5450 gnd.n3395 gnd.n2441 240.244
R5451 gnd.n3395 gnd.n2430 240.244
R5452 gnd.n3392 gnd.n2430 240.244
R5453 gnd.n3392 gnd.n2410 240.244
R5454 gnd.n3722 gnd.n2410 240.244
R5455 gnd.n2882 gnd.n2881 240.244
R5456 gnd.n2953 gnd.n2881 240.244
R5457 gnd.n2951 gnd.n2950 240.244
R5458 gnd.n2947 gnd.n2946 240.244
R5459 gnd.n2943 gnd.n2942 240.244
R5460 gnd.n2939 gnd.n2938 240.244
R5461 gnd.n2935 gnd.n2934 240.244
R5462 gnd.n2931 gnd.n2930 240.244
R5463 gnd.n2927 gnd.n2926 240.244
R5464 gnd.n2923 gnd.n2922 240.244
R5465 gnd.n2919 gnd.n2918 240.244
R5466 gnd.n2915 gnd.n2914 240.244
R5467 gnd.n2911 gnd.n2869 240.244
R5468 gnd.n2971 gnd.n2863 240.244
R5469 gnd.n2971 gnd.n2859 240.244
R5470 gnd.n2977 gnd.n2859 240.244
R5471 gnd.n2977 gnd.n2852 240.244
R5472 gnd.n2987 gnd.n2852 240.244
R5473 gnd.n2987 gnd.n2848 240.244
R5474 gnd.n2993 gnd.n2848 240.244
R5475 gnd.n2993 gnd.n2839 240.244
R5476 gnd.n3033 gnd.n2839 240.244
R5477 gnd.n3033 gnd.n2790 240.244
R5478 gnd.n3041 gnd.n2790 240.244
R5479 gnd.n3041 gnd.n2791 240.244
R5480 gnd.n2791 gnd.n2769 240.244
R5481 gnd.n3062 gnd.n2769 240.244
R5482 gnd.n3062 gnd.n2761 240.244
R5483 gnd.n3073 gnd.n2761 240.244
R5484 gnd.n3073 gnd.n2762 240.244
R5485 gnd.n2762 gnd.n2743 240.244
R5486 gnd.n3093 gnd.n2743 240.244
R5487 gnd.n3093 gnd.n2733 240.244
R5488 gnd.n3103 gnd.n2733 240.244
R5489 gnd.n3103 gnd.n2714 240.244
R5490 gnd.n3124 gnd.n2714 240.244
R5491 gnd.n3124 gnd.n2716 240.244
R5492 gnd.n2716 gnd.n2697 240.244
R5493 gnd.n3152 gnd.n2697 240.244
R5494 gnd.n3152 gnd.n2639 240.244
R5495 gnd.n3204 gnd.n2639 240.244
R5496 gnd.n3204 gnd.n2640 240.244
R5497 gnd.n3200 gnd.n2640 240.244
R5498 gnd.n3200 gnd.n2646 240.244
R5499 gnd.n2661 gnd.n2646 240.244
R5500 gnd.n3190 gnd.n2661 240.244
R5501 gnd.n3190 gnd.n2662 240.244
R5502 gnd.n3186 gnd.n2662 240.244
R5503 gnd.n3186 gnd.n2668 240.244
R5504 gnd.n2668 gnd.n2555 240.244
R5505 gnd.n3243 gnd.n2555 240.244
R5506 gnd.n3243 gnd.n2548 240.244
R5507 gnd.n3254 gnd.n2548 240.244
R5508 gnd.n3254 gnd.n2541 240.244
R5509 gnd.n3269 gnd.n2541 240.244
R5510 gnd.n3269 gnd.n2542 240.244
R5511 gnd.n2542 gnd.n2520 240.244
R5512 gnd.n3291 gnd.n2520 240.244
R5513 gnd.n3291 gnd.n2521 240.244
R5514 gnd.n2521 gnd.n2500 240.244
R5515 gnd.n3328 gnd.n2500 240.244
R5516 gnd.n3328 gnd.n2493 240.244
R5517 gnd.n3339 gnd.n2493 240.244
R5518 gnd.n3339 gnd.n2486 240.244
R5519 gnd.n3354 gnd.n2486 240.244
R5520 gnd.n3354 gnd.n2487 240.244
R5521 gnd.n2487 gnd.n2464 240.244
R5522 gnd.n3376 gnd.n2464 240.244
R5523 gnd.n3376 gnd.n2466 240.244
R5524 gnd.n2466 gnd.n2446 240.244
R5525 gnd.n3417 gnd.n2446 240.244
R5526 gnd.n3417 gnd.n2439 240.244
R5527 gnd.n3428 gnd.n2439 240.244
R5528 gnd.n3428 gnd.n2432 240.244
R5529 gnd.n3697 gnd.n2432 240.244
R5530 gnd.n3697 gnd.n2433 240.244
R5531 gnd.n2433 gnd.n2414 240.244
R5532 gnd.n3720 gnd.n2414 240.244
R5533 gnd.n7510 gnd.n7509 240.244
R5534 gnd.n7515 gnd.n7512 240.244
R5535 gnd.n7518 gnd.n7517 240.244
R5536 gnd.n7523 gnd.n7520 240.244
R5537 gnd.n7526 gnd.n7525 240.244
R5538 gnd.n7531 gnd.n7528 240.244
R5539 gnd.n7534 gnd.n7533 240.244
R5540 gnd.n7538 gnd.n7536 240.244
R5541 gnd.n7541 gnd.n7540 240.244
R5542 gnd.n5915 gnd.n1337 240.244
R5543 gnd.n5915 gnd.n1475 240.244
R5544 gnd.n5922 gnd.n1475 240.244
R5545 gnd.n5922 gnd.n1433 240.244
R5546 gnd.n1433 gnd.n1421 240.244
R5547 gnd.n5946 gnd.n1421 240.244
R5548 gnd.n5946 gnd.n1416 240.244
R5549 gnd.n5958 gnd.n1416 240.244
R5550 gnd.n5958 gnd.n1406 240.244
R5551 gnd.n5951 gnd.n1406 240.244
R5552 gnd.n5951 gnd.n1395 240.244
R5553 gnd.n1395 gnd.n1381 240.244
R5554 gnd.n6018 gnd.n1381 240.244
R5555 gnd.n6018 gnd.n1372 240.244
R5556 gnd.n1386 gnd.n1372 240.244
R5557 gnd.n1386 gnd.n1363 240.244
R5558 gnd.n6000 gnd.n1363 240.244
R5559 gnd.n6000 gnd.n401 240.244
R5560 gnd.n6005 gnd.n401 240.244
R5561 gnd.n6005 gnd.n391 240.244
R5562 gnd.n391 gnd.n383 240.244
R5563 gnd.n7260 gnd.n383 240.244
R5564 gnd.n7260 gnd.n369 240.244
R5565 gnd.n378 gnd.n369 240.244
R5566 gnd.n7268 gnd.n378 240.244
R5567 gnd.n7268 gnd.n357 240.244
R5568 gnd.n357 gnd.n349 240.244
R5569 gnd.n7306 gnd.n349 240.244
R5570 gnd.n7306 gnd.n314 240.244
R5571 gnd.n344 gnd.n314 240.244
R5572 gnd.n7313 gnd.n344 240.244
R5573 gnd.n7313 gnd.n345 240.244
R5574 gnd.n345 gnd.n82 240.244
R5575 gnd.n83 gnd.n82 240.244
R5576 gnd.n84 gnd.n83 240.244
R5577 gnd.n329 gnd.n84 240.244
R5578 gnd.n329 gnd.n87 240.244
R5579 gnd.n88 gnd.n87 240.244
R5580 gnd.n89 gnd.n88 240.244
R5581 gnd.n292 gnd.n89 240.244
R5582 gnd.n292 gnd.n92 240.244
R5583 gnd.n93 gnd.n92 240.244
R5584 gnd.n94 gnd.n93 240.244
R5585 gnd.n277 gnd.n94 240.244
R5586 gnd.n277 gnd.n97 240.244
R5587 gnd.n98 gnd.n97 240.244
R5588 gnd.n99 gnd.n98 240.244
R5589 gnd.n262 gnd.n99 240.244
R5590 gnd.n262 gnd.n102 240.244
R5591 gnd.n103 gnd.n102 240.244
R5592 gnd.n104 gnd.n103 240.244
R5593 gnd.n246 gnd.n104 240.244
R5594 gnd.n246 gnd.n107 240.244
R5595 gnd.n108 gnd.n107 240.244
R5596 gnd.n109 gnd.n108 240.244
R5597 gnd.n231 gnd.n109 240.244
R5598 gnd.n231 gnd.n112 240.244
R5599 gnd.n113 gnd.n112 240.244
R5600 gnd.n114 gnd.n113 240.244
R5601 gnd.n215 gnd.n114 240.244
R5602 gnd.n215 gnd.n117 240.244
R5603 gnd.n118 gnd.n117 240.244
R5604 gnd.n119 gnd.n118 240.244
R5605 gnd.n7666 gnd.n119 240.244
R5606 gnd.n1523 gnd.n1522 240.244
R5607 gnd.n1526 gnd.n1525 240.244
R5608 gnd.n1542 gnd.n1541 240.244
R5609 gnd.n1545 gnd.n1544 240.244
R5610 gnd.n1561 gnd.n1560 240.244
R5611 gnd.n1564 gnd.n1563 240.244
R5612 gnd.n1579 gnd.n1578 240.244
R5613 gnd.n1490 gnd.n1489 240.244
R5614 gnd.n1485 gnd.n1284 240.244
R5615 gnd.n6078 gnd.n1340 240.244
R5616 gnd.n1344 gnd.n1340 240.244
R5617 gnd.n1345 gnd.n1344 240.244
R5618 gnd.n1346 gnd.n1345 240.244
R5619 gnd.n1434 gnd.n1346 240.244
R5620 gnd.n1434 gnd.n1349 240.244
R5621 gnd.n1350 gnd.n1349 240.244
R5622 gnd.n1351 gnd.n1350 240.244
R5623 gnd.n5971 gnd.n1351 240.244
R5624 gnd.n5971 gnd.n1354 240.244
R5625 gnd.n1355 gnd.n1354 240.244
R5626 gnd.n1356 gnd.n1355 240.244
R5627 gnd.n6019 gnd.n1356 240.244
R5628 gnd.n6019 gnd.n1359 240.244
R5629 gnd.n1360 gnd.n1359 240.244
R5630 gnd.n6051 gnd.n1360 240.244
R5631 gnd.n6051 gnd.n403 240.244
R5632 gnd.n7234 gnd.n403 240.244
R5633 gnd.n7234 gnd.n404 240.244
R5634 gnd.n404 gnd.n392 240.244
R5635 gnd.n7227 gnd.n392 240.244
R5636 gnd.n7227 gnd.n371 240.244
R5637 gnd.n7280 gnd.n371 240.244
R5638 gnd.n7280 gnd.n372 240.244
R5639 gnd.n7270 gnd.n372 240.244
R5640 gnd.n7270 gnd.n359 240.244
R5641 gnd.n7271 gnd.n359 240.244
R5642 gnd.n7271 gnd.n316 240.244
R5643 gnd.n7411 gnd.n316 240.244
R5644 gnd.n7411 gnd.n317 240.244
R5645 gnd.n322 gnd.n317 240.244
R5646 gnd.n323 gnd.n322 240.244
R5647 gnd.n324 gnd.n323 240.244
R5648 gnd.n333 gnd.n324 240.244
R5649 gnd.n333 gnd.n327 240.244
R5650 gnd.n7398 gnd.n327 240.244
R5651 gnd.n7398 gnd.n298 240.244
R5652 gnd.n7422 gnd.n298 240.244
R5653 gnd.n7422 gnd.n294 240.244
R5654 gnd.n7428 gnd.n294 240.244
R5655 gnd.n7428 gnd.n282 240.244
R5656 gnd.n7438 gnd.n282 240.244
R5657 gnd.n7438 gnd.n278 240.244
R5658 gnd.n7444 gnd.n278 240.244
R5659 gnd.n7444 gnd.n268 240.244
R5660 gnd.n7454 gnd.n268 240.244
R5661 gnd.n7454 gnd.n264 240.244
R5662 gnd.n7460 gnd.n264 240.244
R5663 gnd.n7460 gnd.n252 240.244
R5664 gnd.n7470 gnd.n252 240.244
R5665 gnd.n7470 gnd.n248 240.244
R5666 gnd.n7476 gnd.n248 240.244
R5667 gnd.n7476 gnd.n237 240.244
R5668 gnd.n7486 gnd.n237 240.244
R5669 gnd.n7486 gnd.n233 240.244
R5670 gnd.n7492 gnd.n233 240.244
R5671 gnd.n7492 gnd.n222 240.244
R5672 gnd.n7502 gnd.n222 240.244
R5673 gnd.n7502 gnd.n216 240.244
R5674 gnd.n7576 gnd.n216 240.244
R5675 gnd.n7576 gnd.n217 240.244
R5676 gnd.n217 gnd.n207 240.244
R5677 gnd.n7507 gnd.n207 240.244
R5678 gnd.n7507 gnd.n129 240.244
R5679 gnd.n2049 gnd.n1113 240.244
R5680 gnd.n2050 gnd.n1999 240.244
R5681 gnd.n2053 gnd.n2000 240.244
R5682 gnd.n2009 gnd.n2008 240.244
R5683 gnd.n2055 gnd.n2016 240.244
R5684 gnd.n2058 gnd.n2017 240.244
R5685 gnd.n2027 gnd.n2026 240.244
R5686 gnd.n2060 gnd.n2034 240.244
R5687 gnd.n2046 gnd.n2035 240.244
R5688 gnd.n3976 gnd.n3815 240.244
R5689 gnd.n3976 gnd.n2334 240.244
R5690 gnd.n3972 gnd.n2334 240.244
R5691 gnd.n3972 gnd.n2327 240.244
R5692 gnd.n3969 gnd.n2327 240.244
R5693 gnd.n3969 gnd.n2319 240.244
R5694 gnd.n3966 gnd.n2319 240.244
R5695 gnd.n3966 gnd.n2310 240.244
R5696 gnd.n3963 gnd.n2310 240.244
R5697 gnd.n3963 gnd.n2302 240.244
R5698 gnd.n3960 gnd.n2302 240.244
R5699 gnd.n3960 gnd.n2295 240.244
R5700 gnd.n3957 gnd.n2295 240.244
R5701 gnd.n3957 gnd.n2287 240.244
R5702 gnd.n3954 gnd.n2287 240.244
R5703 gnd.n3954 gnd.n2278 240.244
R5704 gnd.n3951 gnd.n2278 240.244
R5705 gnd.n3951 gnd.n2270 240.244
R5706 gnd.n3948 gnd.n2270 240.244
R5707 gnd.n3948 gnd.n2263 240.244
R5708 gnd.n3945 gnd.n2263 240.244
R5709 gnd.n3945 gnd.n2255 240.244
R5710 gnd.n3942 gnd.n2255 240.244
R5711 gnd.n3942 gnd.n2246 240.244
R5712 gnd.n3939 gnd.n2246 240.244
R5713 gnd.n3939 gnd.n2238 240.244
R5714 gnd.n3936 gnd.n2238 240.244
R5715 gnd.n3936 gnd.n2232 240.244
R5716 gnd.n3933 gnd.n2232 240.244
R5717 gnd.n3933 gnd.n2223 240.244
R5718 gnd.n3930 gnd.n2223 240.244
R5719 gnd.n3930 gnd.n2215 240.244
R5720 gnd.n3915 gnd.n2215 240.244
R5721 gnd.n3915 gnd.n2196 240.244
R5722 gnd.n3918 gnd.n2196 240.244
R5723 gnd.n3918 gnd.n2190 240.244
R5724 gnd.n3919 gnd.n2190 240.244
R5725 gnd.n3919 gnd.n972 240.244
R5726 gnd.n4365 gnd.n972 240.244
R5727 gnd.n4365 gnd.n985 240.244
R5728 gnd.n4371 gnd.n985 240.244
R5729 gnd.n4371 gnd.n996 240.244
R5730 gnd.n4412 gnd.n996 240.244
R5731 gnd.n4412 gnd.n1006 240.244
R5732 gnd.n2177 gnd.n1006 240.244
R5733 gnd.n2177 gnd.n1017 240.244
R5734 gnd.n4399 gnd.n1017 240.244
R5735 gnd.n4399 gnd.n1028 240.244
R5736 gnd.n2162 gnd.n1028 240.244
R5737 gnd.n2162 gnd.n1038 240.244
R5738 gnd.n4461 gnd.n1038 240.244
R5739 gnd.n4461 gnd.n1048 240.244
R5740 gnd.n2156 gnd.n1048 240.244
R5741 gnd.n2156 gnd.n1059 240.244
R5742 gnd.n4452 gnd.n1059 240.244
R5743 gnd.n4452 gnd.n1070 240.244
R5744 gnd.n4514 gnd.n1070 240.244
R5745 gnd.n4514 gnd.n1080 240.244
R5746 gnd.n4520 gnd.n1080 240.244
R5747 gnd.n4520 gnd.n1091 240.244
R5748 gnd.n4531 gnd.n1091 240.244
R5749 gnd.n4531 gnd.n1102 240.244
R5750 gnd.n4567 gnd.n1102 240.244
R5751 gnd.n4567 gnd.n1111 240.244
R5752 gnd.n3841 gnd.n3839 240.244
R5753 gnd.n3847 gnd.n3833 240.244
R5754 gnd.n3851 gnd.n3849 240.244
R5755 gnd.n3857 gnd.n3829 240.244
R5756 gnd.n3861 gnd.n3859 240.244
R5757 gnd.n3867 gnd.n3825 240.244
R5758 gnd.n3871 gnd.n3869 240.244
R5759 gnd.n3877 gnd.n3821 240.244
R5760 gnd.n3880 gnd.n3879 240.244
R5761 gnd.n4200 gnd.n2335 240.244
R5762 gnd.n4206 gnd.n2335 240.244
R5763 gnd.n4206 gnd.n2324 240.244
R5764 gnd.n4216 gnd.n2324 240.244
R5765 gnd.n4216 gnd.n2320 240.244
R5766 gnd.n4222 gnd.n2320 240.244
R5767 gnd.n4222 gnd.n2307 240.244
R5768 gnd.n4232 gnd.n2307 240.244
R5769 gnd.n4232 gnd.n2303 240.244
R5770 gnd.n4238 gnd.n2303 240.244
R5771 gnd.n4238 gnd.n2292 240.244
R5772 gnd.n4248 gnd.n2292 240.244
R5773 gnd.n4248 gnd.n2288 240.244
R5774 gnd.n4254 gnd.n2288 240.244
R5775 gnd.n4254 gnd.n2275 240.244
R5776 gnd.n4264 gnd.n2275 240.244
R5777 gnd.n4264 gnd.n2271 240.244
R5778 gnd.n4270 gnd.n2271 240.244
R5779 gnd.n4270 gnd.n2260 240.244
R5780 gnd.n4280 gnd.n2260 240.244
R5781 gnd.n4280 gnd.n2256 240.244
R5782 gnd.n4286 gnd.n2256 240.244
R5783 gnd.n4286 gnd.n2243 240.244
R5784 gnd.n4297 gnd.n2243 240.244
R5785 gnd.n4297 gnd.n2239 240.244
R5786 gnd.n4303 gnd.n2239 240.244
R5787 gnd.n4303 gnd.n2229 240.244
R5788 gnd.n4313 gnd.n2229 240.244
R5789 gnd.n4313 gnd.n2224 240.244
R5790 gnd.n4320 gnd.n2224 240.244
R5791 gnd.n4320 gnd.n2225 240.244
R5792 gnd.n2225 gnd.n2217 240.244
R5793 gnd.n2217 gnd.n2199 240.244
R5794 gnd.n4347 gnd.n2199 240.244
R5795 gnd.n4347 gnd.n2200 240.244
R5796 gnd.n2200 gnd.n2191 240.244
R5797 gnd.n4342 gnd.n2191 240.244
R5798 gnd.n4342 gnd.n974 240.244
R5799 gnd.n987 gnd.n974 240.244
R5800 gnd.n6395 gnd.n987 240.244
R5801 gnd.n6395 gnd.n988 240.244
R5802 gnd.n6391 gnd.n988 240.244
R5803 gnd.n6391 gnd.n994 240.244
R5804 gnd.n6383 gnd.n994 240.244
R5805 gnd.n6383 gnd.n1008 240.244
R5806 gnd.n6379 gnd.n1008 240.244
R5807 gnd.n6379 gnd.n1014 240.244
R5808 gnd.n6371 gnd.n1014 240.244
R5809 gnd.n6371 gnd.n1030 240.244
R5810 gnd.n6367 gnd.n1030 240.244
R5811 gnd.n6367 gnd.n1036 240.244
R5812 gnd.n6359 gnd.n1036 240.244
R5813 gnd.n6359 gnd.n1050 240.244
R5814 gnd.n6355 gnd.n1050 240.244
R5815 gnd.n6355 gnd.n1056 240.244
R5816 gnd.n6347 gnd.n1056 240.244
R5817 gnd.n6347 gnd.n1072 240.244
R5818 gnd.n6343 gnd.n1072 240.244
R5819 gnd.n6343 gnd.n1078 240.244
R5820 gnd.n6335 gnd.n1078 240.244
R5821 gnd.n6335 gnd.n1093 240.244
R5822 gnd.n6331 gnd.n1093 240.244
R5823 gnd.n6331 gnd.n1099 240.244
R5824 gnd.n6323 gnd.n1099 240.244
R5825 gnd.n6581 gnd.n796 240.244
R5826 gnd.n6585 gnd.n796 240.244
R5827 gnd.n6585 gnd.n792 240.244
R5828 gnd.n6591 gnd.n792 240.244
R5829 gnd.n6591 gnd.n790 240.244
R5830 gnd.n6595 gnd.n790 240.244
R5831 gnd.n6595 gnd.n786 240.244
R5832 gnd.n6601 gnd.n786 240.244
R5833 gnd.n6601 gnd.n784 240.244
R5834 gnd.n6605 gnd.n784 240.244
R5835 gnd.n6605 gnd.n780 240.244
R5836 gnd.n6611 gnd.n780 240.244
R5837 gnd.n6611 gnd.n778 240.244
R5838 gnd.n6615 gnd.n778 240.244
R5839 gnd.n6615 gnd.n774 240.244
R5840 gnd.n6621 gnd.n774 240.244
R5841 gnd.n6621 gnd.n772 240.244
R5842 gnd.n6625 gnd.n772 240.244
R5843 gnd.n6625 gnd.n768 240.244
R5844 gnd.n6631 gnd.n768 240.244
R5845 gnd.n6631 gnd.n766 240.244
R5846 gnd.n6635 gnd.n766 240.244
R5847 gnd.n6635 gnd.n762 240.244
R5848 gnd.n6641 gnd.n762 240.244
R5849 gnd.n6641 gnd.n760 240.244
R5850 gnd.n6645 gnd.n760 240.244
R5851 gnd.n6645 gnd.n756 240.244
R5852 gnd.n6651 gnd.n756 240.244
R5853 gnd.n6651 gnd.n754 240.244
R5854 gnd.n6655 gnd.n754 240.244
R5855 gnd.n6655 gnd.n750 240.244
R5856 gnd.n6661 gnd.n750 240.244
R5857 gnd.n6661 gnd.n748 240.244
R5858 gnd.n6665 gnd.n748 240.244
R5859 gnd.n6665 gnd.n744 240.244
R5860 gnd.n6671 gnd.n744 240.244
R5861 gnd.n6671 gnd.n742 240.244
R5862 gnd.n6675 gnd.n742 240.244
R5863 gnd.n6675 gnd.n738 240.244
R5864 gnd.n6681 gnd.n738 240.244
R5865 gnd.n6681 gnd.n736 240.244
R5866 gnd.n6685 gnd.n736 240.244
R5867 gnd.n6685 gnd.n732 240.244
R5868 gnd.n6691 gnd.n732 240.244
R5869 gnd.n6691 gnd.n730 240.244
R5870 gnd.n6695 gnd.n730 240.244
R5871 gnd.n6695 gnd.n726 240.244
R5872 gnd.n6701 gnd.n726 240.244
R5873 gnd.n6701 gnd.n724 240.244
R5874 gnd.n6705 gnd.n724 240.244
R5875 gnd.n6705 gnd.n720 240.244
R5876 gnd.n6711 gnd.n720 240.244
R5877 gnd.n6711 gnd.n718 240.244
R5878 gnd.n6715 gnd.n718 240.244
R5879 gnd.n6715 gnd.n714 240.244
R5880 gnd.n6721 gnd.n714 240.244
R5881 gnd.n6721 gnd.n712 240.244
R5882 gnd.n6725 gnd.n712 240.244
R5883 gnd.n6725 gnd.n708 240.244
R5884 gnd.n6731 gnd.n708 240.244
R5885 gnd.n6731 gnd.n706 240.244
R5886 gnd.n6735 gnd.n706 240.244
R5887 gnd.n6735 gnd.n702 240.244
R5888 gnd.n6741 gnd.n702 240.244
R5889 gnd.n6741 gnd.n700 240.244
R5890 gnd.n6745 gnd.n700 240.244
R5891 gnd.n6745 gnd.n696 240.244
R5892 gnd.n6751 gnd.n696 240.244
R5893 gnd.n6751 gnd.n694 240.244
R5894 gnd.n6755 gnd.n694 240.244
R5895 gnd.n6755 gnd.n690 240.244
R5896 gnd.n6761 gnd.n690 240.244
R5897 gnd.n6761 gnd.n688 240.244
R5898 gnd.n6765 gnd.n688 240.244
R5899 gnd.n6765 gnd.n684 240.244
R5900 gnd.n6771 gnd.n684 240.244
R5901 gnd.n6771 gnd.n682 240.244
R5902 gnd.n6775 gnd.n682 240.244
R5903 gnd.n6775 gnd.n678 240.244
R5904 gnd.n6781 gnd.n678 240.244
R5905 gnd.n6781 gnd.n676 240.244
R5906 gnd.n6785 gnd.n676 240.244
R5907 gnd.n6785 gnd.n672 240.244
R5908 gnd.n6791 gnd.n672 240.244
R5909 gnd.n6791 gnd.n670 240.244
R5910 gnd.n6795 gnd.n670 240.244
R5911 gnd.n6795 gnd.n666 240.244
R5912 gnd.n6801 gnd.n666 240.244
R5913 gnd.n6801 gnd.n664 240.244
R5914 gnd.n6805 gnd.n664 240.244
R5915 gnd.n6805 gnd.n660 240.244
R5916 gnd.n6811 gnd.n660 240.244
R5917 gnd.n6811 gnd.n658 240.244
R5918 gnd.n6815 gnd.n658 240.244
R5919 gnd.n6815 gnd.n654 240.244
R5920 gnd.n6821 gnd.n654 240.244
R5921 gnd.n6821 gnd.n652 240.244
R5922 gnd.n6825 gnd.n652 240.244
R5923 gnd.n6825 gnd.n648 240.244
R5924 gnd.n6831 gnd.n648 240.244
R5925 gnd.n6831 gnd.n646 240.244
R5926 gnd.n6835 gnd.n646 240.244
R5927 gnd.n6835 gnd.n642 240.244
R5928 gnd.n6841 gnd.n642 240.244
R5929 gnd.n6841 gnd.n640 240.244
R5930 gnd.n6845 gnd.n640 240.244
R5931 gnd.n6845 gnd.n636 240.244
R5932 gnd.n6851 gnd.n636 240.244
R5933 gnd.n6851 gnd.n634 240.244
R5934 gnd.n6855 gnd.n634 240.244
R5935 gnd.n6855 gnd.n630 240.244
R5936 gnd.n6861 gnd.n630 240.244
R5937 gnd.n6861 gnd.n628 240.244
R5938 gnd.n6865 gnd.n628 240.244
R5939 gnd.n6865 gnd.n624 240.244
R5940 gnd.n6871 gnd.n624 240.244
R5941 gnd.n6871 gnd.n622 240.244
R5942 gnd.n6875 gnd.n622 240.244
R5943 gnd.n6875 gnd.n618 240.244
R5944 gnd.n6881 gnd.n618 240.244
R5945 gnd.n6881 gnd.n616 240.244
R5946 gnd.n6885 gnd.n616 240.244
R5947 gnd.n6885 gnd.n612 240.244
R5948 gnd.n6891 gnd.n612 240.244
R5949 gnd.n6891 gnd.n610 240.244
R5950 gnd.n6895 gnd.n610 240.244
R5951 gnd.n6895 gnd.n606 240.244
R5952 gnd.n6901 gnd.n606 240.244
R5953 gnd.n6901 gnd.n604 240.244
R5954 gnd.n6905 gnd.n604 240.244
R5955 gnd.n6905 gnd.n600 240.244
R5956 gnd.n6911 gnd.n600 240.244
R5957 gnd.n6911 gnd.n598 240.244
R5958 gnd.n6915 gnd.n598 240.244
R5959 gnd.n6915 gnd.n594 240.244
R5960 gnd.n6921 gnd.n594 240.244
R5961 gnd.n6921 gnd.n592 240.244
R5962 gnd.n6925 gnd.n592 240.244
R5963 gnd.n6925 gnd.n588 240.244
R5964 gnd.n6931 gnd.n588 240.244
R5965 gnd.n6931 gnd.n586 240.244
R5966 gnd.n6935 gnd.n586 240.244
R5967 gnd.n6935 gnd.n582 240.244
R5968 gnd.n6941 gnd.n582 240.244
R5969 gnd.n6941 gnd.n580 240.244
R5970 gnd.n6945 gnd.n580 240.244
R5971 gnd.n6945 gnd.n576 240.244
R5972 gnd.n6951 gnd.n576 240.244
R5973 gnd.n6951 gnd.n574 240.244
R5974 gnd.n6955 gnd.n574 240.244
R5975 gnd.n6955 gnd.n570 240.244
R5976 gnd.n6961 gnd.n570 240.244
R5977 gnd.n6961 gnd.n568 240.244
R5978 gnd.n6965 gnd.n568 240.244
R5979 gnd.n6965 gnd.n564 240.244
R5980 gnd.n6971 gnd.n564 240.244
R5981 gnd.n6971 gnd.n562 240.244
R5982 gnd.n6975 gnd.n562 240.244
R5983 gnd.n6975 gnd.n558 240.244
R5984 gnd.n6981 gnd.n558 240.244
R5985 gnd.n6981 gnd.n556 240.244
R5986 gnd.n6985 gnd.n556 240.244
R5987 gnd.n6985 gnd.n552 240.244
R5988 gnd.n6992 gnd.n552 240.244
R5989 gnd.n6992 gnd.n550 240.244
R5990 gnd.n6996 gnd.n550 240.244
R5991 gnd.n6996 gnd.n547 240.244
R5992 gnd.n7002 gnd.n545 240.244
R5993 gnd.n7006 gnd.n545 240.244
R5994 gnd.n7006 gnd.n541 240.244
R5995 gnd.n7012 gnd.n541 240.244
R5996 gnd.n7012 gnd.n539 240.244
R5997 gnd.n7016 gnd.n539 240.244
R5998 gnd.n7016 gnd.n535 240.244
R5999 gnd.n7022 gnd.n535 240.244
R6000 gnd.n7022 gnd.n533 240.244
R6001 gnd.n7026 gnd.n533 240.244
R6002 gnd.n7026 gnd.n529 240.244
R6003 gnd.n7032 gnd.n529 240.244
R6004 gnd.n7032 gnd.n527 240.244
R6005 gnd.n7036 gnd.n527 240.244
R6006 gnd.n7036 gnd.n523 240.244
R6007 gnd.n7042 gnd.n523 240.244
R6008 gnd.n7042 gnd.n521 240.244
R6009 gnd.n7046 gnd.n521 240.244
R6010 gnd.n7046 gnd.n517 240.244
R6011 gnd.n7052 gnd.n517 240.244
R6012 gnd.n7052 gnd.n515 240.244
R6013 gnd.n7056 gnd.n515 240.244
R6014 gnd.n7056 gnd.n511 240.244
R6015 gnd.n7062 gnd.n511 240.244
R6016 gnd.n7062 gnd.n509 240.244
R6017 gnd.n7066 gnd.n509 240.244
R6018 gnd.n7066 gnd.n505 240.244
R6019 gnd.n7072 gnd.n505 240.244
R6020 gnd.n7072 gnd.n503 240.244
R6021 gnd.n7076 gnd.n503 240.244
R6022 gnd.n7076 gnd.n499 240.244
R6023 gnd.n7082 gnd.n499 240.244
R6024 gnd.n7082 gnd.n497 240.244
R6025 gnd.n7086 gnd.n497 240.244
R6026 gnd.n7086 gnd.n493 240.244
R6027 gnd.n7092 gnd.n493 240.244
R6028 gnd.n7092 gnd.n491 240.244
R6029 gnd.n7096 gnd.n491 240.244
R6030 gnd.n7096 gnd.n487 240.244
R6031 gnd.n7102 gnd.n487 240.244
R6032 gnd.n7102 gnd.n485 240.244
R6033 gnd.n7106 gnd.n485 240.244
R6034 gnd.n7106 gnd.n481 240.244
R6035 gnd.n7112 gnd.n481 240.244
R6036 gnd.n7112 gnd.n479 240.244
R6037 gnd.n7116 gnd.n479 240.244
R6038 gnd.n7116 gnd.n475 240.244
R6039 gnd.n7122 gnd.n475 240.244
R6040 gnd.n7122 gnd.n473 240.244
R6041 gnd.n7126 gnd.n473 240.244
R6042 gnd.n7126 gnd.n469 240.244
R6043 gnd.n7132 gnd.n469 240.244
R6044 gnd.n7132 gnd.n467 240.244
R6045 gnd.n7136 gnd.n467 240.244
R6046 gnd.n7136 gnd.n463 240.244
R6047 gnd.n7142 gnd.n463 240.244
R6048 gnd.n7142 gnd.n461 240.244
R6049 gnd.n7146 gnd.n461 240.244
R6050 gnd.n7146 gnd.n457 240.244
R6051 gnd.n7152 gnd.n457 240.244
R6052 gnd.n7152 gnd.n455 240.244
R6053 gnd.n7156 gnd.n455 240.244
R6054 gnd.n7156 gnd.n451 240.244
R6055 gnd.n7162 gnd.n451 240.244
R6056 gnd.n7162 gnd.n449 240.244
R6057 gnd.n7166 gnd.n449 240.244
R6058 gnd.n7166 gnd.n445 240.244
R6059 gnd.n7172 gnd.n445 240.244
R6060 gnd.n7172 gnd.n443 240.244
R6061 gnd.n7176 gnd.n443 240.244
R6062 gnd.n7176 gnd.n439 240.244
R6063 gnd.n7182 gnd.n439 240.244
R6064 gnd.n7182 gnd.n437 240.244
R6065 gnd.n7186 gnd.n437 240.244
R6066 gnd.n7186 gnd.n433 240.244
R6067 gnd.n7192 gnd.n433 240.244
R6068 gnd.n7192 gnd.n431 240.244
R6069 gnd.n7196 gnd.n431 240.244
R6070 gnd.n7196 gnd.n427 240.244
R6071 gnd.n7202 gnd.n427 240.244
R6072 gnd.n7202 gnd.n425 240.244
R6073 gnd.n7207 gnd.n425 240.244
R6074 gnd.n7207 gnd.n421 240.244
R6075 gnd.n7213 gnd.n421 240.244
R6076 gnd.n6404 gnd.n969 240.244
R6077 gnd.n4374 gnd.n969 240.244
R6078 gnd.n4374 gnd.n4372 240.244
R6079 gnd.n4380 gnd.n4372 240.244
R6080 gnd.n4380 gnd.n2171 240.244
R6081 gnd.n4415 gnd.n2171 240.244
R6082 gnd.n4415 gnd.n2167 240.244
R6083 gnd.n4421 gnd.n2167 240.244
R6084 gnd.n4422 gnd.n4421 240.244
R6085 gnd.n4423 gnd.n4422 240.244
R6086 gnd.n4423 gnd.n2163 240.244
R6087 gnd.n4429 gnd.n2163 240.244
R6088 gnd.n4429 gnd.n2150 240.244
R6089 gnd.n4464 gnd.n2150 240.244
R6090 gnd.n4464 gnd.n2146 240.244
R6091 gnd.n4470 gnd.n2146 240.244
R6092 gnd.n4471 gnd.n4470 240.244
R6093 gnd.n4472 gnd.n4471 240.244
R6094 gnd.n4472 gnd.n2141 240.244
R6095 gnd.n4511 gnd.n2141 240.244
R6096 gnd.n4511 gnd.n2142 240.244
R6097 gnd.n4507 gnd.n2142 240.244
R6098 gnd.n4507 gnd.n4506 240.244
R6099 gnd.n4506 gnd.n4505 240.244
R6100 gnd.n4505 gnd.n4480 240.244
R6101 gnd.n4501 gnd.n4480 240.244
R6102 gnd.n4501 gnd.n4500 240.244
R6103 gnd.n4500 gnd.n4499 240.244
R6104 gnd.n4499 gnd.n4486 240.244
R6105 gnd.n4495 gnd.n4486 240.244
R6106 gnd.n4495 gnd.n4493 240.244
R6107 gnd.n4493 gnd.n1972 240.244
R6108 gnd.n4907 gnd.n1972 240.244
R6109 gnd.n4907 gnd.n1968 240.244
R6110 gnd.n4913 gnd.n1968 240.244
R6111 gnd.n4913 gnd.n1960 240.244
R6112 gnd.n4923 gnd.n1960 240.244
R6113 gnd.n4923 gnd.n1956 240.244
R6114 gnd.n4929 gnd.n1956 240.244
R6115 gnd.n4929 gnd.n1947 240.244
R6116 gnd.n4939 gnd.n1947 240.244
R6117 gnd.n4939 gnd.n1943 240.244
R6118 gnd.n4945 gnd.n1943 240.244
R6119 gnd.n4945 gnd.n1934 240.244
R6120 gnd.n4955 gnd.n1934 240.244
R6121 gnd.n4955 gnd.n1930 240.244
R6122 gnd.n4961 gnd.n1930 240.244
R6123 gnd.n4961 gnd.n1921 240.244
R6124 gnd.n4971 gnd.n1921 240.244
R6125 gnd.n4971 gnd.n1917 240.244
R6126 gnd.n4977 gnd.n1917 240.244
R6127 gnd.n4977 gnd.n1907 240.244
R6128 gnd.n4987 gnd.n1907 240.244
R6129 gnd.n4987 gnd.n1902 240.244
R6130 gnd.n4995 gnd.n1902 240.244
R6131 gnd.n4995 gnd.n1903 240.244
R6132 gnd.n1903 gnd.n1876 240.244
R6133 gnd.n5573 gnd.n1876 240.244
R6134 gnd.n5573 gnd.n1872 240.244
R6135 gnd.n5579 gnd.n1872 240.244
R6136 gnd.n5579 gnd.n1862 240.244
R6137 gnd.n5589 gnd.n1862 240.244
R6138 gnd.n5589 gnd.n1858 240.244
R6139 gnd.n5595 gnd.n1858 240.244
R6140 gnd.n5595 gnd.n1847 240.244
R6141 gnd.n5605 gnd.n1847 240.244
R6142 gnd.n5605 gnd.n1843 240.244
R6143 gnd.n5611 gnd.n1843 240.244
R6144 gnd.n5611 gnd.n1832 240.244
R6145 gnd.n5621 gnd.n1832 240.244
R6146 gnd.n5621 gnd.n1828 240.244
R6147 gnd.n5627 gnd.n1828 240.244
R6148 gnd.n5627 gnd.n1818 240.244
R6149 gnd.n5637 gnd.n1818 240.244
R6150 gnd.n5637 gnd.n1814 240.244
R6151 gnd.n5643 gnd.n1814 240.244
R6152 gnd.n5643 gnd.n1803 240.244
R6153 gnd.n5653 gnd.n1803 240.244
R6154 gnd.n5653 gnd.n1799 240.244
R6155 gnd.n5659 gnd.n1799 240.244
R6156 gnd.n5659 gnd.n1788 240.244
R6157 gnd.n5669 gnd.n1788 240.244
R6158 gnd.n5669 gnd.n1784 240.244
R6159 gnd.n5675 gnd.n1784 240.244
R6160 gnd.n5675 gnd.n1773 240.244
R6161 gnd.n5685 gnd.n1773 240.244
R6162 gnd.n5685 gnd.n1769 240.244
R6163 gnd.n5691 gnd.n1769 240.244
R6164 gnd.n5691 gnd.n1759 240.244
R6165 gnd.n5701 gnd.n1759 240.244
R6166 gnd.n5701 gnd.n1755 240.244
R6167 gnd.n5707 gnd.n1755 240.244
R6168 gnd.n5707 gnd.n1744 240.244
R6169 gnd.n5717 gnd.n1744 240.244
R6170 gnd.n5717 gnd.n1740 240.244
R6171 gnd.n5723 gnd.n1740 240.244
R6172 gnd.n5723 gnd.n1731 240.244
R6173 gnd.n5733 gnd.n1731 240.244
R6174 gnd.n5733 gnd.n1727 240.244
R6175 gnd.n5739 gnd.n1727 240.244
R6176 gnd.n5739 gnd.n1719 240.244
R6177 gnd.n5749 gnd.n1719 240.244
R6178 gnd.n5749 gnd.n1715 240.244
R6179 gnd.n5755 gnd.n1715 240.244
R6180 gnd.n5755 gnd.n1705 240.244
R6181 gnd.n5765 gnd.n1705 240.244
R6182 gnd.n5765 gnd.n1701 240.244
R6183 gnd.n5771 gnd.n1701 240.244
R6184 gnd.n5771 gnd.n1692 240.244
R6185 gnd.n5781 gnd.n1692 240.244
R6186 gnd.n5781 gnd.n1688 240.244
R6187 gnd.n5787 gnd.n1688 240.244
R6188 gnd.n5787 gnd.n1678 240.244
R6189 gnd.n5797 gnd.n1678 240.244
R6190 gnd.n5797 gnd.n1674 240.244
R6191 gnd.n5803 gnd.n1674 240.244
R6192 gnd.n5803 gnd.n1665 240.244
R6193 gnd.n5813 gnd.n1665 240.244
R6194 gnd.n5813 gnd.n1661 240.244
R6195 gnd.n5819 gnd.n1661 240.244
R6196 gnd.n5819 gnd.n1652 240.244
R6197 gnd.n5829 gnd.n1652 240.244
R6198 gnd.n5829 gnd.n1648 240.244
R6199 gnd.n5835 gnd.n1648 240.244
R6200 gnd.n5835 gnd.n1638 240.244
R6201 gnd.n5845 gnd.n1638 240.244
R6202 gnd.n5845 gnd.n1634 240.244
R6203 gnd.n5851 gnd.n1634 240.244
R6204 gnd.n5851 gnd.n1625 240.244
R6205 gnd.n5863 gnd.n1625 240.244
R6206 gnd.n5863 gnd.n1620 240.244
R6207 gnd.n5872 gnd.n1620 240.244
R6208 gnd.n5872 gnd.n1621 240.244
R6209 gnd.n1621 gnd.n1246 240.244
R6210 gnd.n6162 gnd.n1246 240.244
R6211 gnd.n6162 gnd.n1249 240.244
R6212 gnd.n6158 gnd.n1249 240.244
R6213 gnd.n6158 gnd.n1255 240.244
R6214 gnd.n1444 gnd.n1255 240.244
R6215 gnd.n1444 gnd.n1441 240.244
R6216 gnd.n1450 gnd.n1441 240.244
R6217 gnd.n1451 gnd.n1450 240.244
R6218 gnd.n5925 gnd.n1451 240.244
R6219 gnd.n5925 gnd.n1436 240.244
R6220 gnd.n5933 gnd.n1436 240.244
R6221 gnd.n5933 gnd.n1437 240.244
R6222 gnd.n1437 gnd.n1413 240.244
R6223 gnd.n5961 gnd.n1413 240.244
R6224 gnd.n5961 gnd.n1408 240.244
R6225 gnd.n5969 gnd.n1408 240.244
R6226 gnd.n5969 gnd.n1409 240.244
R6227 gnd.n1409 gnd.n1379 240.244
R6228 gnd.n6022 gnd.n1379 240.244
R6229 gnd.n6022 gnd.n1374 240.244
R6230 gnd.n6040 gnd.n1374 240.244
R6231 gnd.n6040 gnd.n1375 240.244
R6232 gnd.n6036 gnd.n1375 240.244
R6233 gnd.n6036 gnd.n6035 240.244
R6234 gnd.n6035 gnd.n6034 240.244
R6235 gnd.n6034 gnd.n409 240.244
R6236 gnd.n7224 gnd.n409 240.244
R6237 gnd.n7224 gnd.n410 240.244
R6238 gnd.n7220 gnd.n410 240.244
R6239 gnd.n7220 gnd.n7219 240.244
R6240 gnd.n7219 gnd.n7218 240.244
R6241 gnd.n7218 gnd.n416 240.244
R6242 gnd.n7214 gnd.n416 240.244
R6243 gnd.n6575 gnd.n798 240.244
R6244 gnd.n6575 gnd.n801 240.244
R6245 gnd.n6571 gnd.n801 240.244
R6246 gnd.n6571 gnd.n803 240.244
R6247 gnd.n6567 gnd.n803 240.244
R6248 gnd.n6567 gnd.n809 240.244
R6249 gnd.n6563 gnd.n809 240.244
R6250 gnd.n6563 gnd.n811 240.244
R6251 gnd.n6559 gnd.n811 240.244
R6252 gnd.n6559 gnd.n817 240.244
R6253 gnd.n6555 gnd.n817 240.244
R6254 gnd.n6555 gnd.n819 240.244
R6255 gnd.n6551 gnd.n819 240.244
R6256 gnd.n6551 gnd.n825 240.244
R6257 gnd.n6547 gnd.n825 240.244
R6258 gnd.n6547 gnd.n827 240.244
R6259 gnd.n6543 gnd.n827 240.244
R6260 gnd.n6543 gnd.n833 240.244
R6261 gnd.n6539 gnd.n833 240.244
R6262 gnd.n6539 gnd.n835 240.244
R6263 gnd.n6535 gnd.n835 240.244
R6264 gnd.n6535 gnd.n841 240.244
R6265 gnd.n6531 gnd.n841 240.244
R6266 gnd.n6531 gnd.n843 240.244
R6267 gnd.n6527 gnd.n843 240.244
R6268 gnd.n6527 gnd.n849 240.244
R6269 gnd.n6523 gnd.n849 240.244
R6270 gnd.n6523 gnd.n851 240.244
R6271 gnd.n6519 gnd.n851 240.244
R6272 gnd.n6519 gnd.n857 240.244
R6273 gnd.n6515 gnd.n857 240.244
R6274 gnd.n6515 gnd.n859 240.244
R6275 gnd.n6511 gnd.n859 240.244
R6276 gnd.n6511 gnd.n865 240.244
R6277 gnd.n6507 gnd.n865 240.244
R6278 gnd.n6507 gnd.n867 240.244
R6279 gnd.n6503 gnd.n867 240.244
R6280 gnd.n6503 gnd.n873 240.244
R6281 gnd.n6499 gnd.n873 240.244
R6282 gnd.n6499 gnd.n875 240.244
R6283 gnd.n6495 gnd.n875 240.244
R6284 gnd.n6495 gnd.n881 240.244
R6285 gnd.n6491 gnd.n881 240.244
R6286 gnd.n6491 gnd.n883 240.244
R6287 gnd.n6487 gnd.n883 240.244
R6288 gnd.n6487 gnd.n889 240.244
R6289 gnd.n6483 gnd.n889 240.244
R6290 gnd.n6483 gnd.n891 240.244
R6291 gnd.n6479 gnd.n891 240.244
R6292 gnd.n6479 gnd.n897 240.244
R6293 gnd.n6475 gnd.n897 240.244
R6294 gnd.n6475 gnd.n899 240.244
R6295 gnd.n6471 gnd.n899 240.244
R6296 gnd.n6471 gnd.n905 240.244
R6297 gnd.n6467 gnd.n905 240.244
R6298 gnd.n6467 gnd.n907 240.244
R6299 gnd.n6463 gnd.n907 240.244
R6300 gnd.n6463 gnd.n913 240.244
R6301 gnd.n6459 gnd.n913 240.244
R6302 gnd.n6459 gnd.n915 240.244
R6303 gnd.n6455 gnd.n915 240.244
R6304 gnd.n6455 gnd.n921 240.244
R6305 gnd.n6451 gnd.n921 240.244
R6306 gnd.n6451 gnd.n923 240.244
R6307 gnd.n6447 gnd.n923 240.244
R6308 gnd.n6447 gnd.n929 240.244
R6309 gnd.n6443 gnd.n929 240.244
R6310 gnd.n6443 gnd.n931 240.244
R6311 gnd.n6439 gnd.n931 240.244
R6312 gnd.n6439 gnd.n937 240.244
R6313 gnd.n6435 gnd.n937 240.244
R6314 gnd.n6435 gnd.n939 240.244
R6315 gnd.n6431 gnd.n939 240.244
R6316 gnd.n6431 gnd.n945 240.244
R6317 gnd.n6427 gnd.n945 240.244
R6318 gnd.n6427 gnd.n947 240.244
R6319 gnd.n6423 gnd.n947 240.244
R6320 gnd.n6423 gnd.n953 240.244
R6321 gnd.n6419 gnd.n953 240.244
R6322 gnd.n6419 gnd.n955 240.244
R6323 gnd.n6415 gnd.n955 240.244
R6324 gnd.n6415 gnd.n961 240.244
R6325 gnd.n6411 gnd.n961 240.244
R6326 gnd.n6411 gnd.n963 240.244
R6327 gnd.n1119 gnd.n1118 240.244
R6328 gnd.n1120 gnd.n1119 240.244
R6329 gnd.n1961 gnd.n1120 240.244
R6330 gnd.n1961 gnd.n1123 240.244
R6331 gnd.n1124 gnd.n1123 240.244
R6332 gnd.n1125 gnd.n1124 240.244
R6333 gnd.n1948 gnd.n1125 240.244
R6334 gnd.n1948 gnd.n1128 240.244
R6335 gnd.n1129 gnd.n1128 240.244
R6336 gnd.n1130 gnd.n1129 240.244
R6337 gnd.n1941 gnd.n1130 240.244
R6338 gnd.n1941 gnd.n1133 240.244
R6339 gnd.n1134 gnd.n1133 240.244
R6340 gnd.n1135 gnd.n1134 240.244
R6341 gnd.n1928 gnd.n1135 240.244
R6342 gnd.n1928 gnd.n1138 240.244
R6343 gnd.n1139 gnd.n1138 240.244
R6344 gnd.n1140 gnd.n1139 240.244
R6345 gnd.n1908 gnd.n1140 240.244
R6346 gnd.n1908 gnd.n1143 240.244
R6347 gnd.n1144 gnd.n1143 240.244
R6348 gnd.n1145 gnd.n1144 240.244
R6349 gnd.n1892 gnd.n1145 240.244
R6350 gnd.n1892 gnd.n1148 240.244
R6351 gnd.n1149 gnd.n1148 240.244
R6352 gnd.n1150 gnd.n1149 240.244
R6353 gnd.n1870 gnd.n1150 240.244
R6354 gnd.n1870 gnd.n1153 240.244
R6355 gnd.n1154 gnd.n1153 240.244
R6356 gnd.n1155 gnd.n1154 240.244
R6357 gnd.n1856 gnd.n1155 240.244
R6358 gnd.n1856 gnd.n1158 240.244
R6359 gnd.n1159 gnd.n1158 240.244
R6360 gnd.n1160 gnd.n1159 240.244
R6361 gnd.n1841 gnd.n1160 240.244
R6362 gnd.n1841 gnd.n1163 240.244
R6363 gnd.n1164 gnd.n1163 240.244
R6364 gnd.n1165 gnd.n1164 240.244
R6365 gnd.n1826 gnd.n1165 240.244
R6366 gnd.n1826 gnd.n1168 240.244
R6367 gnd.n1169 gnd.n1168 240.244
R6368 gnd.n1170 gnd.n1169 240.244
R6369 gnd.n1812 gnd.n1170 240.244
R6370 gnd.n1812 gnd.n1173 240.244
R6371 gnd.n1174 gnd.n1173 240.244
R6372 gnd.n1175 gnd.n1174 240.244
R6373 gnd.n1797 gnd.n1175 240.244
R6374 gnd.n1797 gnd.n1178 240.244
R6375 gnd.n1179 gnd.n1178 240.244
R6376 gnd.n1180 gnd.n1179 240.244
R6377 gnd.n1782 gnd.n1180 240.244
R6378 gnd.n1782 gnd.n1183 240.244
R6379 gnd.n1184 gnd.n1183 240.244
R6380 gnd.n1185 gnd.n1184 240.244
R6381 gnd.n1767 gnd.n1185 240.244
R6382 gnd.n1767 gnd.n1188 240.244
R6383 gnd.n1189 gnd.n1188 240.244
R6384 gnd.n1190 gnd.n1189 240.244
R6385 gnd.n1752 gnd.n1190 240.244
R6386 gnd.n1752 gnd.n1193 240.244
R6387 gnd.n1194 gnd.n1193 240.244
R6388 gnd.n1195 gnd.n1194 240.244
R6389 gnd.n1738 gnd.n1195 240.244
R6390 gnd.n1738 gnd.n1198 240.244
R6391 gnd.n1199 gnd.n1198 240.244
R6392 gnd.n1200 gnd.n1199 240.244
R6393 gnd.n1726 gnd.n1200 240.244
R6394 gnd.n1726 gnd.n1203 240.244
R6395 gnd.n1204 gnd.n1203 240.244
R6396 gnd.n1205 gnd.n1204 240.244
R6397 gnd.n1714 gnd.n1205 240.244
R6398 gnd.n1714 gnd.n1208 240.244
R6399 gnd.n1209 gnd.n1208 240.244
R6400 gnd.n1210 gnd.n1209 240.244
R6401 gnd.n1700 gnd.n1210 240.244
R6402 gnd.n1700 gnd.n1213 240.244
R6403 gnd.n1214 gnd.n1213 240.244
R6404 gnd.n1215 gnd.n1214 240.244
R6405 gnd.n1685 gnd.n1215 240.244
R6406 gnd.n1685 gnd.n1218 240.244
R6407 gnd.n1219 gnd.n1218 240.244
R6408 gnd.n1220 gnd.n1219 240.244
R6409 gnd.n1673 gnd.n1220 240.244
R6410 gnd.n1673 gnd.n1223 240.244
R6411 gnd.n1224 gnd.n1223 240.244
R6412 gnd.n1225 gnd.n1224 240.244
R6413 gnd.n1660 gnd.n1225 240.244
R6414 gnd.n1660 gnd.n1228 240.244
R6415 gnd.n1229 gnd.n1228 240.244
R6416 gnd.n1230 gnd.n1229 240.244
R6417 gnd.n1647 gnd.n1230 240.244
R6418 gnd.n1647 gnd.n1233 240.244
R6419 gnd.n1234 gnd.n1233 240.244
R6420 gnd.n1235 gnd.n1234 240.244
R6421 gnd.n1633 gnd.n1235 240.244
R6422 gnd.n1633 gnd.n1238 240.244
R6423 gnd.n1239 gnd.n1238 240.244
R6424 gnd.n1240 gnd.n1239 240.244
R6425 gnd.n1619 gnd.n1240 240.244
R6426 gnd.n1619 gnd.n1243 240.244
R6427 gnd.n6165 gnd.n1243 240.244
R6428 gnd.n1993 gnd.n1992 240.244
R6429 gnd.n2003 gnd.n1992 240.244
R6430 gnd.n2005 gnd.n2004 240.244
R6431 gnd.n2013 gnd.n2012 240.244
R6432 gnd.n2021 gnd.n2020 240.244
R6433 gnd.n2023 gnd.n2022 240.244
R6434 gnd.n2031 gnd.n2030 240.244
R6435 gnd.n2041 gnd.n2040 240.244
R6436 gnd.n2043 gnd.n2042 240.244
R6437 gnd.n4537 gnd.n4536 240.244
R6438 gnd.n4539 gnd.n4538 240.244
R6439 gnd.n4543 gnd.n4542 240.244
R6440 gnd.n4549 gnd.n4544 240.244
R6441 gnd.n4899 gnd.n1978 240.244
R6442 gnd.n4905 gnd.n1967 240.244
R6443 gnd.n4915 gnd.n1967 240.244
R6444 gnd.n4915 gnd.n1963 240.244
R6445 gnd.n4921 gnd.n1963 240.244
R6446 gnd.n4921 gnd.n1954 240.244
R6447 gnd.n4931 gnd.n1954 240.244
R6448 gnd.n4931 gnd.n1950 240.244
R6449 gnd.n4937 gnd.n1950 240.244
R6450 gnd.n4937 gnd.n1939 240.244
R6451 gnd.n4947 gnd.n1939 240.244
R6452 gnd.n4947 gnd.n1935 240.244
R6453 gnd.n4953 gnd.n1935 240.244
R6454 gnd.n4953 gnd.n1926 240.244
R6455 gnd.n4963 gnd.n1926 240.244
R6456 gnd.n4963 gnd.n1922 240.244
R6457 gnd.n4969 gnd.n1922 240.244
R6458 gnd.n4969 gnd.n1915 240.244
R6459 gnd.n4979 gnd.n1915 240.244
R6460 gnd.n4979 gnd.n1911 240.244
R6461 gnd.n4985 gnd.n1911 240.244
R6462 gnd.n4985 gnd.n1900 240.244
R6463 gnd.n4997 gnd.n1900 240.244
R6464 gnd.n4997 gnd.n1895 240.244
R6465 gnd.n5004 gnd.n1895 240.244
R6466 gnd.n5004 gnd.n1879 240.244
R6467 gnd.n1879 gnd.n1868 240.244
R6468 gnd.n5581 gnd.n1868 240.244
R6469 gnd.n5581 gnd.n1864 240.244
R6470 gnd.n5587 gnd.n1864 240.244
R6471 gnd.n5587 gnd.n1854 240.244
R6472 gnd.n5597 gnd.n1854 240.244
R6473 gnd.n5597 gnd.n1850 240.244
R6474 gnd.n5603 gnd.n1850 240.244
R6475 gnd.n5603 gnd.n1839 240.244
R6476 gnd.n5613 gnd.n1839 240.244
R6477 gnd.n5613 gnd.n1835 240.244
R6478 gnd.n5619 gnd.n1835 240.244
R6479 gnd.n5619 gnd.n1825 240.244
R6480 gnd.n5629 gnd.n1825 240.244
R6481 gnd.n5629 gnd.n1821 240.244
R6482 gnd.n5635 gnd.n1821 240.244
R6483 gnd.n5635 gnd.n1810 240.244
R6484 gnd.n5645 gnd.n1810 240.244
R6485 gnd.n5645 gnd.n1806 240.244
R6486 gnd.n5651 gnd.n1806 240.244
R6487 gnd.n5651 gnd.n1795 240.244
R6488 gnd.n5661 gnd.n1795 240.244
R6489 gnd.n5661 gnd.n1791 240.244
R6490 gnd.n5667 gnd.n1791 240.244
R6491 gnd.n5667 gnd.n1780 240.244
R6492 gnd.n5677 gnd.n1780 240.244
R6493 gnd.n5677 gnd.n1776 240.244
R6494 gnd.n5683 gnd.n1776 240.244
R6495 gnd.n5683 gnd.n1765 240.244
R6496 gnd.n5693 gnd.n1765 240.244
R6497 gnd.n5693 gnd.n1761 240.244
R6498 gnd.n5699 gnd.n1761 240.244
R6499 gnd.n5699 gnd.n1750 240.244
R6500 gnd.n5709 gnd.n1750 240.244
R6501 gnd.n5709 gnd.n1746 240.244
R6502 gnd.n5715 gnd.n1746 240.244
R6503 gnd.n5715 gnd.n1737 240.244
R6504 gnd.n5725 gnd.n1737 240.244
R6505 gnd.n5725 gnd.n1733 240.244
R6506 gnd.n5731 gnd.n1733 240.244
R6507 gnd.n5731 gnd.n1725 240.244
R6508 gnd.n5741 gnd.n1725 240.244
R6509 gnd.n5741 gnd.n1721 240.244
R6510 gnd.n5747 gnd.n1721 240.244
R6511 gnd.n5747 gnd.n1712 240.244
R6512 gnd.n5757 gnd.n1712 240.244
R6513 gnd.n5757 gnd.n1708 240.244
R6514 gnd.n5763 gnd.n1708 240.244
R6515 gnd.n5763 gnd.n1698 240.244
R6516 gnd.n5773 gnd.n1698 240.244
R6517 gnd.n5773 gnd.n1694 240.244
R6518 gnd.n5779 gnd.n1694 240.244
R6519 gnd.n5779 gnd.n1683 240.244
R6520 gnd.n5789 gnd.n1683 240.244
R6521 gnd.n5789 gnd.n1679 240.244
R6522 gnd.n5795 gnd.n1679 240.244
R6523 gnd.n5795 gnd.n1671 240.244
R6524 gnd.n5805 gnd.n1671 240.244
R6525 gnd.n5805 gnd.n1667 240.244
R6526 gnd.n5811 gnd.n1667 240.244
R6527 gnd.n5811 gnd.n1658 240.244
R6528 gnd.n5821 gnd.n1658 240.244
R6529 gnd.n5821 gnd.n1654 240.244
R6530 gnd.n5827 gnd.n1654 240.244
R6531 gnd.n5827 gnd.n1645 240.244
R6532 gnd.n5837 gnd.n1645 240.244
R6533 gnd.n5837 gnd.n1641 240.244
R6534 gnd.n5843 gnd.n1641 240.244
R6535 gnd.n5843 gnd.n1632 240.244
R6536 gnd.n5853 gnd.n1632 240.244
R6537 gnd.n5853 gnd.n1627 240.244
R6538 gnd.n5861 gnd.n1627 240.244
R6539 gnd.n5861 gnd.n1617 240.244
R6540 gnd.n5874 gnd.n1617 240.244
R6541 gnd.n5875 gnd.n5874 240.244
R6542 gnd.n5875 gnd.n1247 240.244
R6543 gnd.n1532 gnd.n1531 240.244
R6544 gnd.n1535 gnd.n1534 240.244
R6545 gnd.n1551 gnd.n1550 240.244
R6546 gnd.n1554 gnd.n1553 240.244
R6547 gnd.n1570 gnd.n1569 240.244
R6548 gnd.n1573 gnd.n1572 240.244
R6549 gnd.n1586 gnd.n1585 240.244
R6550 gnd.n1589 gnd.n1588 240.244
R6551 gnd.n1600 gnd.n1599 240.244
R6552 gnd.n1603 gnd.n1602 240.244
R6553 gnd.n1608 gnd.n1605 240.244
R6554 gnd.n1611 gnd.n1610 240.244
R6555 gnd.n5880 gnd.n1613 240.244
R6556 gnd.n5883 gnd.n5882 240.244
R6557 gnd.n4649 gnd.n4648 240.132
R6558 gnd.n5196 gnd.n5195 240.132
R6559 gnd.n6583 gnd.n6582 225.874
R6560 gnd.n6584 gnd.n6583 225.874
R6561 gnd.n6584 gnd.n791 225.874
R6562 gnd.n6592 gnd.n791 225.874
R6563 gnd.n6593 gnd.n6592 225.874
R6564 gnd.n6594 gnd.n6593 225.874
R6565 gnd.n6594 gnd.n785 225.874
R6566 gnd.n6602 gnd.n785 225.874
R6567 gnd.n6603 gnd.n6602 225.874
R6568 gnd.n6604 gnd.n6603 225.874
R6569 gnd.n6604 gnd.n779 225.874
R6570 gnd.n6612 gnd.n779 225.874
R6571 gnd.n6613 gnd.n6612 225.874
R6572 gnd.n6614 gnd.n6613 225.874
R6573 gnd.n6614 gnd.n773 225.874
R6574 gnd.n6622 gnd.n773 225.874
R6575 gnd.n6623 gnd.n6622 225.874
R6576 gnd.n6624 gnd.n6623 225.874
R6577 gnd.n6624 gnd.n767 225.874
R6578 gnd.n6632 gnd.n767 225.874
R6579 gnd.n6633 gnd.n6632 225.874
R6580 gnd.n6634 gnd.n6633 225.874
R6581 gnd.n6634 gnd.n761 225.874
R6582 gnd.n6642 gnd.n761 225.874
R6583 gnd.n6643 gnd.n6642 225.874
R6584 gnd.n6644 gnd.n6643 225.874
R6585 gnd.n6644 gnd.n755 225.874
R6586 gnd.n6652 gnd.n755 225.874
R6587 gnd.n6653 gnd.n6652 225.874
R6588 gnd.n6654 gnd.n6653 225.874
R6589 gnd.n6654 gnd.n749 225.874
R6590 gnd.n6662 gnd.n749 225.874
R6591 gnd.n6663 gnd.n6662 225.874
R6592 gnd.n6664 gnd.n6663 225.874
R6593 gnd.n6664 gnd.n743 225.874
R6594 gnd.n6672 gnd.n743 225.874
R6595 gnd.n6673 gnd.n6672 225.874
R6596 gnd.n6674 gnd.n6673 225.874
R6597 gnd.n6674 gnd.n737 225.874
R6598 gnd.n6682 gnd.n737 225.874
R6599 gnd.n6683 gnd.n6682 225.874
R6600 gnd.n6684 gnd.n6683 225.874
R6601 gnd.n6684 gnd.n731 225.874
R6602 gnd.n6692 gnd.n731 225.874
R6603 gnd.n6693 gnd.n6692 225.874
R6604 gnd.n6694 gnd.n6693 225.874
R6605 gnd.n6694 gnd.n725 225.874
R6606 gnd.n6702 gnd.n725 225.874
R6607 gnd.n6703 gnd.n6702 225.874
R6608 gnd.n6704 gnd.n6703 225.874
R6609 gnd.n6704 gnd.n719 225.874
R6610 gnd.n6712 gnd.n719 225.874
R6611 gnd.n6713 gnd.n6712 225.874
R6612 gnd.n6714 gnd.n6713 225.874
R6613 gnd.n6714 gnd.n713 225.874
R6614 gnd.n6722 gnd.n713 225.874
R6615 gnd.n6723 gnd.n6722 225.874
R6616 gnd.n6724 gnd.n6723 225.874
R6617 gnd.n6724 gnd.n707 225.874
R6618 gnd.n6732 gnd.n707 225.874
R6619 gnd.n6733 gnd.n6732 225.874
R6620 gnd.n6734 gnd.n6733 225.874
R6621 gnd.n6734 gnd.n701 225.874
R6622 gnd.n6742 gnd.n701 225.874
R6623 gnd.n6743 gnd.n6742 225.874
R6624 gnd.n6744 gnd.n6743 225.874
R6625 gnd.n6744 gnd.n695 225.874
R6626 gnd.n6752 gnd.n695 225.874
R6627 gnd.n6753 gnd.n6752 225.874
R6628 gnd.n6754 gnd.n6753 225.874
R6629 gnd.n6754 gnd.n689 225.874
R6630 gnd.n6762 gnd.n689 225.874
R6631 gnd.n6763 gnd.n6762 225.874
R6632 gnd.n6764 gnd.n6763 225.874
R6633 gnd.n6764 gnd.n683 225.874
R6634 gnd.n6772 gnd.n683 225.874
R6635 gnd.n6773 gnd.n6772 225.874
R6636 gnd.n6774 gnd.n6773 225.874
R6637 gnd.n6774 gnd.n677 225.874
R6638 gnd.n6782 gnd.n677 225.874
R6639 gnd.n6783 gnd.n6782 225.874
R6640 gnd.n6784 gnd.n6783 225.874
R6641 gnd.n6784 gnd.n671 225.874
R6642 gnd.n6792 gnd.n671 225.874
R6643 gnd.n6793 gnd.n6792 225.874
R6644 gnd.n6794 gnd.n6793 225.874
R6645 gnd.n6794 gnd.n665 225.874
R6646 gnd.n6802 gnd.n665 225.874
R6647 gnd.n6803 gnd.n6802 225.874
R6648 gnd.n6804 gnd.n6803 225.874
R6649 gnd.n6804 gnd.n659 225.874
R6650 gnd.n6812 gnd.n659 225.874
R6651 gnd.n6813 gnd.n6812 225.874
R6652 gnd.n6814 gnd.n6813 225.874
R6653 gnd.n6814 gnd.n653 225.874
R6654 gnd.n6822 gnd.n653 225.874
R6655 gnd.n6823 gnd.n6822 225.874
R6656 gnd.n6824 gnd.n6823 225.874
R6657 gnd.n6824 gnd.n647 225.874
R6658 gnd.n6832 gnd.n647 225.874
R6659 gnd.n6833 gnd.n6832 225.874
R6660 gnd.n6834 gnd.n6833 225.874
R6661 gnd.n6834 gnd.n641 225.874
R6662 gnd.n6842 gnd.n641 225.874
R6663 gnd.n6843 gnd.n6842 225.874
R6664 gnd.n6844 gnd.n6843 225.874
R6665 gnd.n6844 gnd.n635 225.874
R6666 gnd.n6852 gnd.n635 225.874
R6667 gnd.n6853 gnd.n6852 225.874
R6668 gnd.n6854 gnd.n6853 225.874
R6669 gnd.n6854 gnd.n629 225.874
R6670 gnd.n6862 gnd.n629 225.874
R6671 gnd.n6863 gnd.n6862 225.874
R6672 gnd.n6864 gnd.n6863 225.874
R6673 gnd.n6864 gnd.n623 225.874
R6674 gnd.n6872 gnd.n623 225.874
R6675 gnd.n6873 gnd.n6872 225.874
R6676 gnd.n6874 gnd.n6873 225.874
R6677 gnd.n6874 gnd.n617 225.874
R6678 gnd.n6882 gnd.n617 225.874
R6679 gnd.n6883 gnd.n6882 225.874
R6680 gnd.n6884 gnd.n6883 225.874
R6681 gnd.n6884 gnd.n611 225.874
R6682 gnd.n6892 gnd.n611 225.874
R6683 gnd.n6893 gnd.n6892 225.874
R6684 gnd.n6894 gnd.n6893 225.874
R6685 gnd.n6894 gnd.n605 225.874
R6686 gnd.n6902 gnd.n605 225.874
R6687 gnd.n6903 gnd.n6902 225.874
R6688 gnd.n6904 gnd.n6903 225.874
R6689 gnd.n6904 gnd.n599 225.874
R6690 gnd.n6912 gnd.n599 225.874
R6691 gnd.n6913 gnd.n6912 225.874
R6692 gnd.n6914 gnd.n6913 225.874
R6693 gnd.n6914 gnd.n593 225.874
R6694 gnd.n6922 gnd.n593 225.874
R6695 gnd.n6923 gnd.n6922 225.874
R6696 gnd.n6924 gnd.n6923 225.874
R6697 gnd.n6924 gnd.n587 225.874
R6698 gnd.n6932 gnd.n587 225.874
R6699 gnd.n6933 gnd.n6932 225.874
R6700 gnd.n6934 gnd.n6933 225.874
R6701 gnd.n6934 gnd.n581 225.874
R6702 gnd.n6942 gnd.n581 225.874
R6703 gnd.n6943 gnd.n6942 225.874
R6704 gnd.n6944 gnd.n6943 225.874
R6705 gnd.n6944 gnd.n575 225.874
R6706 gnd.n6952 gnd.n575 225.874
R6707 gnd.n6953 gnd.n6952 225.874
R6708 gnd.n6954 gnd.n6953 225.874
R6709 gnd.n6954 gnd.n569 225.874
R6710 gnd.n6962 gnd.n569 225.874
R6711 gnd.n6963 gnd.n6962 225.874
R6712 gnd.n6964 gnd.n6963 225.874
R6713 gnd.n6964 gnd.n563 225.874
R6714 gnd.n6972 gnd.n563 225.874
R6715 gnd.n6973 gnd.n6972 225.874
R6716 gnd.n6974 gnd.n6973 225.874
R6717 gnd.n6974 gnd.n557 225.874
R6718 gnd.n6982 gnd.n557 225.874
R6719 gnd.n6983 gnd.n6982 225.874
R6720 gnd.n6984 gnd.n6983 225.874
R6721 gnd.n6984 gnd.n551 225.874
R6722 gnd.n6993 gnd.n551 225.874
R6723 gnd.n6994 gnd.n6993 225.874
R6724 gnd.n6995 gnd.n6994 225.874
R6725 gnd.n6995 gnd.n546 225.874
R6726 gnd.n2906 gnd.t297 224.174
R6727 gnd.n2403 gnd.t274 224.174
R6728 gnd.n1306 gnd.n1263 199.319
R6729 gnd.n1306 gnd.n1264 199.319
R6730 gnd.n2105 gnd.n2075 199.319
R6731 gnd.n2105 gnd.n2074 199.319
R6732 gnd.n4650 gnd.n4647 186.49
R6733 gnd.n5197 gnd.n5194 186.49
R6734 gnd.n3681 gnd.n3680 185
R6735 gnd.n3679 gnd.n3678 185
R6736 gnd.n3658 gnd.n3657 185
R6737 gnd.n3673 gnd.n3672 185
R6738 gnd.n3671 gnd.n3670 185
R6739 gnd.n3662 gnd.n3661 185
R6740 gnd.n3665 gnd.n3664 185
R6741 gnd.n3649 gnd.n3648 185
R6742 gnd.n3647 gnd.n3646 185
R6743 gnd.n3626 gnd.n3625 185
R6744 gnd.n3641 gnd.n3640 185
R6745 gnd.n3639 gnd.n3638 185
R6746 gnd.n3630 gnd.n3629 185
R6747 gnd.n3633 gnd.n3632 185
R6748 gnd.n3617 gnd.n3616 185
R6749 gnd.n3615 gnd.n3614 185
R6750 gnd.n3594 gnd.n3593 185
R6751 gnd.n3609 gnd.n3608 185
R6752 gnd.n3607 gnd.n3606 185
R6753 gnd.n3598 gnd.n3597 185
R6754 gnd.n3601 gnd.n3600 185
R6755 gnd.n3586 gnd.n3585 185
R6756 gnd.n3584 gnd.n3583 185
R6757 gnd.n3563 gnd.n3562 185
R6758 gnd.n3578 gnd.n3577 185
R6759 gnd.n3576 gnd.n3575 185
R6760 gnd.n3567 gnd.n3566 185
R6761 gnd.n3570 gnd.n3569 185
R6762 gnd.n3554 gnd.n3553 185
R6763 gnd.n3552 gnd.n3551 185
R6764 gnd.n3531 gnd.n3530 185
R6765 gnd.n3546 gnd.n3545 185
R6766 gnd.n3544 gnd.n3543 185
R6767 gnd.n3535 gnd.n3534 185
R6768 gnd.n3538 gnd.n3537 185
R6769 gnd.n3522 gnd.n3521 185
R6770 gnd.n3520 gnd.n3519 185
R6771 gnd.n3499 gnd.n3498 185
R6772 gnd.n3514 gnd.n3513 185
R6773 gnd.n3512 gnd.n3511 185
R6774 gnd.n3503 gnd.n3502 185
R6775 gnd.n3506 gnd.n3505 185
R6776 gnd.n3490 gnd.n3489 185
R6777 gnd.n3488 gnd.n3487 185
R6778 gnd.n3467 gnd.n3466 185
R6779 gnd.n3482 gnd.n3481 185
R6780 gnd.n3480 gnd.n3479 185
R6781 gnd.n3471 gnd.n3470 185
R6782 gnd.n3474 gnd.n3473 185
R6783 gnd.n3459 gnd.n3458 185
R6784 gnd.n3457 gnd.n3456 185
R6785 gnd.n3436 gnd.n3435 185
R6786 gnd.n3451 gnd.n3450 185
R6787 gnd.n3449 gnd.n3448 185
R6788 gnd.n3440 gnd.n3439 185
R6789 gnd.n3443 gnd.n3442 185
R6790 gnd.n2907 gnd.t296 178.987
R6791 gnd.n2404 gnd.t275 178.987
R6792 gnd.n1 gnd.t154 170.774
R6793 gnd.n9 gnd.t355 170.103
R6794 gnd.n8 gnd.t6 170.103
R6795 gnd.n7 gnd.t351 170.103
R6796 gnd.n6 gnd.t152 170.103
R6797 gnd.n5 gnd.t343 170.103
R6798 gnd.n4 gnd.t45 170.103
R6799 gnd.n3 gnd.t187 170.103
R6800 gnd.n2 gnd.t60 170.103
R6801 gnd.n1 gnd.t150 170.103
R6802 gnd.n6123 gnd.n1305 164.544
R6803 gnd.n4818 gnd.n4817 164.544
R6804 gnd.n5370 gnd.n5369 163.367
R6805 gnd.n5367 gnd.n5206 163.367
R6806 gnd.n5363 gnd.n5362 163.367
R6807 gnd.n5360 gnd.n5209 163.367
R6808 gnd.n5356 gnd.n5355 163.367
R6809 gnd.n5353 gnd.n5212 163.367
R6810 gnd.n5349 gnd.n5348 163.367
R6811 gnd.n5346 gnd.n5215 163.367
R6812 gnd.n5342 gnd.n5341 163.367
R6813 gnd.n5339 gnd.n5218 163.367
R6814 gnd.n5335 gnd.n5334 163.367
R6815 gnd.n5332 gnd.n5221 163.367
R6816 gnd.n5328 gnd.n5327 163.367
R6817 gnd.n5325 gnd.n5224 163.367
R6818 gnd.n5320 gnd.n5319 163.367
R6819 gnd.n5317 gnd.n5315 163.367
R6820 gnd.n5312 gnd.n5311 163.367
R6821 gnd.n5309 gnd.n5230 163.367
R6822 gnd.n5304 gnd.n5303 163.367
R6823 gnd.n5301 gnd.n5235 163.367
R6824 gnd.n5297 gnd.n5296 163.367
R6825 gnd.n5294 gnd.n5238 163.367
R6826 gnd.n5290 gnd.n5289 163.367
R6827 gnd.n5287 gnd.n5241 163.367
R6828 gnd.n5283 gnd.n5282 163.367
R6829 gnd.n5280 gnd.n5244 163.367
R6830 gnd.n5276 gnd.n5275 163.367
R6831 gnd.n5273 gnd.n5247 163.367
R6832 gnd.n5269 gnd.n5268 163.367
R6833 gnd.n5266 gnd.n5250 163.367
R6834 gnd.n5262 gnd.n5261 163.367
R6835 gnd.n5259 gnd.n5253 163.367
R6836 gnd.n4749 gnd.n4640 163.367
R6837 gnd.n4640 gnd.n1894 163.367
R6838 gnd.n1894 gnd.n1880 163.367
R6839 gnd.n5571 gnd.n1880 163.367
R6840 gnd.n5571 gnd.n1881 163.367
R6841 gnd.n5567 gnd.n1881 163.367
R6842 gnd.n5567 gnd.n5566 163.367
R6843 gnd.n5566 gnd.n5565 163.367
R6844 gnd.n5565 gnd.n1884 163.367
R6845 gnd.n5020 gnd.n1884 163.367
R6846 gnd.n5555 gnd.n5020 163.367
R6847 gnd.n5555 gnd.n5021 163.367
R6848 gnd.n5551 gnd.n5021 163.367
R6849 gnd.n5551 gnd.n5550 163.367
R6850 gnd.n5550 gnd.n5025 163.367
R6851 gnd.n5033 gnd.n5025 163.367
R6852 gnd.n5540 gnd.n5033 163.367
R6853 gnd.n5540 gnd.n5034 163.367
R6854 gnd.n5536 gnd.n5034 163.367
R6855 gnd.n5536 gnd.n5535 163.367
R6856 gnd.n5535 gnd.n5038 163.367
R6857 gnd.n5049 gnd.n5038 163.367
R6858 gnd.n5049 gnd.n5046 163.367
R6859 gnd.n5524 gnd.n5046 163.367
R6860 gnd.n5524 gnd.n5047 163.367
R6861 gnd.n5520 gnd.n5047 163.367
R6862 gnd.n5520 gnd.n5053 163.367
R6863 gnd.n5061 gnd.n5053 163.367
R6864 gnd.n5511 gnd.n5061 163.367
R6865 gnd.n5511 gnd.n5062 163.367
R6866 gnd.n5507 gnd.n5062 163.367
R6867 gnd.n5507 gnd.n5506 163.367
R6868 gnd.n5506 gnd.n5065 163.367
R6869 gnd.n5074 gnd.n5065 163.367
R6870 gnd.n5497 gnd.n5074 163.367
R6871 gnd.n5497 gnd.n5075 163.367
R6872 gnd.n5493 gnd.n5075 163.367
R6873 gnd.n5493 gnd.n5492 163.367
R6874 gnd.n5492 gnd.n5079 163.367
R6875 gnd.n5088 gnd.n5079 163.367
R6876 gnd.n5483 gnd.n5088 163.367
R6877 gnd.n5483 gnd.n5089 163.367
R6878 gnd.n5479 gnd.n5089 163.367
R6879 gnd.n5479 gnd.n5478 163.367
R6880 gnd.n5478 gnd.n5093 163.367
R6881 gnd.n5102 gnd.n5093 163.367
R6882 gnd.n5469 gnd.n5102 163.367
R6883 gnd.n5469 gnd.n5103 163.367
R6884 gnd.n5465 gnd.n5103 163.367
R6885 gnd.n5465 gnd.n5464 163.367
R6886 gnd.n5464 gnd.n5107 163.367
R6887 gnd.n5115 gnd.n5107 163.367
R6888 gnd.n5454 gnd.n5115 163.367
R6889 gnd.n5454 gnd.n1754 163.367
R6890 gnd.n5450 gnd.n1754 163.367
R6891 gnd.n5450 gnd.n5449 163.367
R6892 gnd.n5449 gnd.n5119 163.367
R6893 gnd.n5127 gnd.n5119 163.367
R6894 gnd.n5439 gnd.n5127 163.367
R6895 gnd.n5439 gnd.n5128 163.367
R6896 gnd.n5435 gnd.n5128 163.367
R6897 gnd.n5435 gnd.n5132 163.367
R6898 gnd.n5142 gnd.n5132 163.367
R6899 gnd.n5142 gnd.n5140 163.367
R6900 gnd.n5424 gnd.n5140 163.367
R6901 gnd.n5424 gnd.n5141 163.367
R6902 gnd.n5420 gnd.n5141 163.367
R6903 gnd.n5420 gnd.n5146 163.367
R6904 gnd.n5155 gnd.n5146 163.367
R6905 gnd.n5410 gnd.n5155 163.367
R6906 gnd.n5410 gnd.n5156 163.367
R6907 gnd.n5406 gnd.n5156 163.367
R6908 gnd.n5406 gnd.n5159 163.367
R6909 gnd.n5170 gnd.n5159 163.367
R6910 gnd.n5170 gnd.n5168 163.367
R6911 gnd.n5395 gnd.n5168 163.367
R6912 gnd.n5395 gnd.n5169 163.367
R6913 gnd.n5391 gnd.n5169 163.367
R6914 gnd.n5391 gnd.n5174 163.367
R6915 gnd.n5383 gnd.n5174 163.367
R6916 gnd.n5383 gnd.n5180 163.367
R6917 gnd.n5379 gnd.n5180 163.367
R6918 gnd.n5379 gnd.n5182 163.367
R6919 gnd.n4741 gnd.n4739 163.367
R6920 gnd.n4739 gnd.n4738 163.367
R6921 gnd.n4735 gnd.n4734 163.367
R6922 gnd.n4732 gnd.n4666 163.367
R6923 gnd.n4728 gnd.n4726 163.367
R6924 gnd.n4724 gnd.n4668 163.367
R6925 gnd.n4720 gnd.n4718 163.367
R6926 gnd.n4716 gnd.n4670 163.367
R6927 gnd.n4712 gnd.n4710 163.367
R6928 gnd.n4708 gnd.n4672 163.367
R6929 gnd.n4704 gnd.n4702 163.367
R6930 gnd.n4700 gnd.n4674 163.367
R6931 gnd.n4696 gnd.n4694 163.367
R6932 gnd.n4692 gnd.n4676 163.367
R6933 gnd.n4688 gnd.n4686 163.367
R6934 gnd.n4683 gnd.n4682 163.367
R6935 gnd.n4816 gnd.n4814 163.367
R6936 gnd.n4812 gnd.n4620 163.367
R6937 gnd.n4807 gnd.n4805 163.367
R6938 gnd.n4803 gnd.n4624 163.367
R6939 gnd.n4799 gnd.n4797 163.367
R6940 gnd.n4795 gnd.n4626 163.367
R6941 gnd.n4791 gnd.n4789 163.367
R6942 gnd.n4787 gnd.n4628 163.367
R6943 gnd.n4783 gnd.n4781 163.367
R6944 gnd.n4779 gnd.n4630 163.367
R6945 gnd.n4775 gnd.n4773 163.367
R6946 gnd.n4771 gnd.n4632 163.367
R6947 gnd.n4767 gnd.n4765 163.367
R6948 gnd.n4763 gnd.n4634 163.367
R6949 gnd.n4759 gnd.n4757 163.367
R6950 gnd.n4755 gnd.n4636 163.367
R6951 gnd.n4747 gnd.n1891 163.367
R6952 gnd.n5007 gnd.n1891 163.367
R6953 gnd.n5008 gnd.n5007 163.367
R6954 gnd.n5008 gnd.n1878 163.367
R6955 gnd.n5014 gnd.n1878 163.367
R6956 gnd.n5015 gnd.n5014 163.367
R6957 gnd.n5015 gnd.n1887 163.367
R6958 gnd.n5563 gnd.n1887 163.367
R6959 gnd.n5563 gnd.n1889 163.367
R6960 gnd.n5559 gnd.n1889 163.367
R6961 gnd.n5559 gnd.n5558 163.367
R6962 gnd.n5558 gnd.n5019 163.367
R6963 gnd.n5027 gnd.n5019 163.367
R6964 gnd.n5548 gnd.n5027 163.367
R6965 gnd.n5548 gnd.n5028 163.367
R6966 gnd.n5544 gnd.n5028 163.367
R6967 gnd.n5544 gnd.n5543 163.367
R6968 gnd.n5543 gnd.n5032 163.367
R6969 gnd.n5040 gnd.n5032 163.367
R6970 gnd.n5533 gnd.n5040 163.367
R6971 gnd.n5533 gnd.n5041 163.367
R6972 gnd.n5529 gnd.n5041 163.367
R6973 gnd.n5529 gnd.n5528 163.367
R6974 gnd.n5528 gnd.n5045 163.367
R6975 gnd.n5055 gnd.n5045 163.367
R6976 gnd.n5518 gnd.n5055 163.367
R6977 gnd.n5518 gnd.n5056 163.367
R6978 gnd.n5514 gnd.n5056 163.367
R6979 gnd.n5514 gnd.n5513 163.367
R6980 gnd.n5513 gnd.n5060 163.367
R6981 gnd.n5067 gnd.n5060 163.367
R6982 gnd.n5504 gnd.n5067 163.367
R6983 gnd.n5504 gnd.n5068 163.367
R6984 gnd.n5500 gnd.n5068 163.367
R6985 gnd.n5500 gnd.n5499 163.367
R6986 gnd.n5499 gnd.n5072 163.367
R6987 gnd.n5081 gnd.n5072 163.367
R6988 gnd.n5490 gnd.n5081 163.367
R6989 gnd.n5490 gnd.n5082 163.367
R6990 gnd.n5486 gnd.n5082 163.367
R6991 gnd.n5486 gnd.n5485 163.367
R6992 gnd.n5485 gnd.n5086 163.367
R6993 gnd.n5095 gnd.n5086 163.367
R6994 gnd.n5476 gnd.n5095 163.367
R6995 gnd.n5476 gnd.n5096 163.367
R6996 gnd.n5472 gnd.n5096 163.367
R6997 gnd.n5472 gnd.n5471 163.367
R6998 gnd.n5471 gnd.n5100 163.367
R6999 gnd.n5109 gnd.n5100 163.367
R7000 gnd.n5462 gnd.n5109 163.367
R7001 gnd.n5462 gnd.n5110 163.367
R7002 gnd.n5458 gnd.n5110 163.367
R7003 gnd.n5458 gnd.n5114 163.367
R7004 gnd.n5114 gnd.n1751 163.367
R7005 gnd.n5121 gnd.n1751 163.367
R7006 gnd.n5447 gnd.n5121 163.367
R7007 gnd.n5447 gnd.n5122 163.367
R7008 gnd.n5443 gnd.n5122 163.367
R7009 gnd.n5443 gnd.n5126 163.367
R7010 gnd.n5134 gnd.n5126 163.367
R7011 gnd.n5433 gnd.n5134 163.367
R7012 gnd.n5433 gnd.n5136 163.367
R7013 gnd.n5429 gnd.n5136 163.367
R7014 gnd.n5429 gnd.n5428 163.367
R7015 gnd.n5428 gnd.n5139 163.367
R7016 gnd.n5149 gnd.n5139 163.367
R7017 gnd.n5418 gnd.n5149 163.367
R7018 gnd.n5418 gnd.n5150 163.367
R7019 gnd.n5414 gnd.n5150 163.367
R7020 gnd.n5414 gnd.n5154 163.367
R7021 gnd.n5160 gnd.n5154 163.367
R7022 gnd.n5404 gnd.n5160 163.367
R7023 gnd.n5404 gnd.n5163 163.367
R7024 gnd.n5400 gnd.n5163 163.367
R7025 gnd.n5400 gnd.n5399 163.367
R7026 gnd.n5399 gnd.n5398 163.367
R7027 gnd.n5398 gnd.n5166 163.367
R7028 gnd.n5389 gnd.n5166 163.367
R7029 gnd.n5389 gnd.n5175 163.367
R7030 gnd.n5385 gnd.n5175 163.367
R7031 gnd.n5385 gnd.n5178 163.367
R7032 gnd.n5377 gnd.n5178 163.367
R7033 gnd.n5377 gnd.n5184 163.367
R7034 gnd.n5203 gnd.n5202 156.462
R7035 gnd.n3621 gnd.n3589 153.042
R7036 gnd.n3685 gnd.n3684 152.079
R7037 gnd.n3653 gnd.n3652 152.079
R7038 gnd.n3621 gnd.n3620 152.079
R7039 gnd.n4655 gnd.n4654 152
R7040 gnd.n4656 gnd.n4645 152
R7041 gnd.n4658 gnd.n4657 152
R7042 gnd.n4660 gnd.n4643 152
R7043 gnd.n4662 gnd.n4661 152
R7044 gnd.n5201 gnd.n5185 152
R7045 gnd.n5193 gnd.n5186 152
R7046 gnd.n5192 gnd.n5191 152
R7047 gnd.n5190 gnd.n5187 152
R7048 gnd.n5188 gnd.t269 150.546
R7049 gnd.t117 gnd.n3663 147.661
R7050 gnd.t40 gnd.n3631 147.661
R7051 gnd.t168 gnd.n3599 147.661
R7052 gnd.t4 gnd.n3568 147.661
R7053 gnd.t341 gnd.n3536 147.661
R7054 gnd.t331 gnd.n3504 147.661
R7055 gnd.t158 gnd.n3472 147.661
R7056 gnd.t170 gnd.n3441 147.661
R7057 gnd.n5314 gnd.n5313 143.351
R7058 gnd.n4681 gnd.n4619 143.351
R7059 gnd.n4815 gnd.n4619 143.351
R7060 gnd.n4652 gnd.t226 130.484
R7061 gnd.n4661 gnd.t229 126.766
R7062 gnd.n4659 gnd.t301 126.766
R7063 gnd.n4645 gnd.t327 126.766
R7064 gnd.n4653 gnd.t276 126.766
R7065 gnd.n5189 gnd.t248 126.766
R7066 gnd.n5191 gnd.t282 126.766
R7067 gnd.n5200 gnd.t259 126.766
R7068 gnd.n5202 gnd.t285 126.766
R7069 gnd.n3680 gnd.n3679 104.615
R7070 gnd.n3679 gnd.n3657 104.615
R7071 gnd.n3672 gnd.n3657 104.615
R7072 gnd.n3672 gnd.n3671 104.615
R7073 gnd.n3671 gnd.n3661 104.615
R7074 gnd.n3664 gnd.n3661 104.615
R7075 gnd.n3648 gnd.n3647 104.615
R7076 gnd.n3647 gnd.n3625 104.615
R7077 gnd.n3640 gnd.n3625 104.615
R7078 gnd.n3640 gnd.n3639 104.615
R7079 gnd.n3639 gnd.n3629 104.615
R7080 gnd.n3632 gnd.n3629 104.615
R7081 gnd.n3616 gnd.n3615 104.615
R7082 gnd.n3615 gnd.n3593 104.615
R7083 gnd.n3608 gnd.n3593 104.615
R7084 gnd.n3608 gnd.n3607 104.615
R7085 gnd.n3607 gnd.n3597 104.615
R7086 gnd.n3600 gnd.n3597 104.615
R7087 gnd.n3585 gnd.n3584 104.615
R7088 gnd.n3584 gnd.n3562 104.615
R7089 gnd.n3577 gnd.n3562 104.615
R7090 gnd.n3577 gnd.n3576 104.615
R7091 gnd.n3576 gnd.n3566 104.615
R7092 gnd.n3569 gnd.n3566 104.615
R7093 gnd.n3553 gnd.n3552 104.615
R7094 gnd.n3552 gnd.n3530 104.615
R7095 gnd.n3545 gnd.n3530 104.615
R7096 gnd.n3545 gnd.n3544 104.615
R7097 gnd.n3544 gnd.n3534 104.615
R7098 gnd.n3537 gnd.n3534 104.615
R7099 gnd.n3521 gnd.n3520 104.615
R7100 gnd.n3520 gnd.n3498 104.615
R7101 gnd.n3513 gnd.n3498 104.615
R7102 gnd.n3513 gnd.n3512 104.615
R7103 gnd.n3512 gnd.n3502 104.615
R7104 gnd.n3505 gnd.n3502 104.615
R7105 gnd.n3489 gnd.n3488 104.615
R7106 gnd.n3488 gnd.n3466 104.615
R7107 gnd.n3481 gnd.n3466 104.615
R7108 gnd.n3481 gnd.n3480 104.615
R7109 gnd.n3480 gnd.n3470 104.615
R7110 gnd.n3473 gnd.n3470 104.615
R7111 gnd.n3458 gnd.n3457 104.615
R7112 gnd.n3457 gnd.n3435 104.615
R7113 gnd.n3450 gnd.n3435 104.615
R7114 gnd.n3450 gnd.n3449 104.615
R7115 gnd.n3449 gnd.n3439 104.615
R7116 gnd.n3442 gnd.n3439 104.615
R7117 gnd.n2832 gnd.t314 100.632
R7118 gnd.n2377 gnd.t257 100.632
R7119 gnd.n7657 gnd.n138 99.6594
R7120 gnd.n7655 gnd.n7654 99.6594
R7121 gnd.n7650 gnd.n145 99.6594
R7122 gnd.n7648 gnd.n7647 99.6594
R7123 gnd.n7643 gnd.n152 99.6594
R7124 gnd.n7641 gnd.n7640 99.6594
R7125 gnd.n7636 gnd.n159 99.6594
R7126 gnd.n7634 gnd.n7633 99.6594
R7127 gnd.n7626 gnd.n166 99.6594
R7128 gnd.n7624 gnd.n7623 99.6594
R7129 gnd.n7619 gnd.n173 99.6594
R7130 gnd.n7617 gnd.n7616 99.6594
R7131 gnd.n7612 gnd.n180 99.6594
R7132 gnd.n7610 gnd.n7609 99.6594
R7133 gnd.n7605 gnd.n187 99.6594
R7134 gnd.n7603 gnd.n7602 99.6594
R7135 gnd.n7598 gnd.n194 99.6594
R7136 gnd.n7596 gnd.n7595 99.6594
R7137 gnd.n199 gnd.n198 99.6594
R7138 gnd.n6154 gnd.n6153 99.6594
R7139 gnd.n6148 gnd.n1257 99.6594
R7140 gnd.n6145 gnd.n1258 99.6594
R7141 gnd.n6141 gnd.n1259 99.6594
R7142 gnd.n6137 gnd.n1260 99.6594
R7143 gnd.n6133 gnd.n1261 99.6594
R7144 gnd.n6129 gnd.n1262 99.6594
R7145 gnd.n6125 gnd.n1263 99.6594
R7146 gnd.n6120 gnd.n1265 99.6594
R7147 gnd.n6116 gnd.n1266 99.6594
R7148 gnd.n6112 gnd.n1267 99.6594
R7149 gnd.n6108 gnd.n1268 99.6594
R7150 gnd.n6104 gnd.n1269 99.6594
R7151 gnd.n6100 gnd.n1270 99.6594
R7152 gnd.n6096 gnd.n1271 99.6594
R7153 gnd.n6092 gnd.n1272 99.6594
R7154 gnd.n6088 gnd.n1273 99.6594
R7155 gnd.n1329 gnd.n1274 99.6594
R7156 gnd.n4846 gnd.n4845 99.6594
R7157 gnd.n4841 gnd.n2081 99.6594
R7158 gnd.n4837 gnd.n2080 99.6594
R7159 gnd.n4833 gnd.n2079 99.6594
R7160 gnd.n4829 gnd.n2078 99.6594
R7161 gnd.n4825 gnd.n2077 99.6594
R7162 gnd.n4821 gnd.n2076 99.6594
R7163 gnd.n4611 gnd.n2074 99.6594
R7164 gnd.n4609 gnd.n2073 99.6594
R7165 gnd.n4605 gnd.n2072 99.6594
R7166 gnd.n4601 gnd.n2071 99.6594
R7167 gnd.n4597 gnd.n2070 99.6594
R7168 gnd.n4593 gnd.n2069 99.6594
R7169 gnd.n4589 gnd.n2068 99.6594
R7170 gnd.n4585 gnd.n2067 99.6594
R7171 gnd.n4581 gnd.n2066 99.6594
R7172 gnd.n4577 gnd.n2065 99.6594
R7173 gnd.n2123 gnd.n2064 99.6594
R7174 gnd.n4191 gnd.n3978 99.6594
R7175 gnd.n4189 gnd.n3981 99.6594
R7176 gnd.n4185 gnd.n4184 99.6594
R7177 gnd.n4178 gnd.n3986 99.6594
R7178 gnd.n4177 gnd.n4176 99.6594
R7179 gnd.n4170 gnd.n3992 99.6594
R7180 gnd.n4169 gnd.n4168 99.6594
R7181 gnd.n4162 gnd.n3998 99.6594
R7182 gnd.n4161 gnd.n4160 99.6594
R7183 gnd.n4154 gnd.n4004 99.6594
R7184 gnd.n4153 gnd.n4152 99.6594
R7185 gnd.n4146 gnd.n4013 99.6594
R7186 gnd.n4145 gnd.n4144 99.6594
R7187 gnd.n4138 gnd.n4019 99.6594
R7188 gnd.n4137 gnd.n4136 99.6594
R7189 gnd.n4130 gnd.n4025 99.6594
R7190 gnd.n4129 gnd.n4128 99.6594
R7191 gnd.n4035 gnd.n4031 99.6594
R7192 gnd.n4118 gnd.n4117 99.6594
R7193 gnd.n3803 gnd.n2360 99.6594
R7194 gnd.n3801 gnd.n2359 99.6594
R7195 gnd.n3797 gnd.n2358 99.6594
R7196 gnd.n3793 gnd.n2357 99.6594
R7197 gnd.n3789 gnd.n2356 99.6594
R7198 gnd.n3785 gnd.n2355 99.6594
R7199 gnd.n3781 gnd.n2354 99.6594
R7200 gnd.n3713 gnd.n2353 99.6594
R7201 gnd.n3044 gnd.n2775 99.6594
R7202 gnd.n2801 gnd.n2782 99.6594
R7203 gnd.n2803 gnd.n2783 99.6594
R7204 gnd.n2811 gnd.n2784 99.6594
R7205 gnd.n2813 gnd.n2785 99.6594
R7206 gnd.n2821 gnd.n2786 99.6594
R7207 gnd.n2823 gnd.n2787 99.6594
R7208 gnd.n2831 gnd.n2788 99.6594
R7209 gnd.n3771 gnd.n2340 99.6594
R7210 gnd.n3767 gnd.n2341 99.6594
R7211 gnd.n3763 gnd.n2342 99.6594
R7212 gnd.n3759 gnd.n2343 99.6594
R7213 gnd.n3755 gnd.n2344 99.6594
R7214 gnd.n3751 gnd.n2345 99.6594
R7215 gnd.n3747 gnd.n2346 99.6594
R7216 gnd.n3743 gnd.n2347 99.6594
R7217 gnd.n3739 gnd.n2348 99.6594
R7218 gnd.n3735 gnd.n2349 99.6594
R7219 gnd.n3731 gnd.n2350 99.6594
R7220 gnd.n3727 gnd.n2351 99.6594
R7221 gnd.n3723 gnd.n2352 99.6594
R7222 gnd.n2959 gnd.n2958 99.6594
R7223 gnd.n2953 gnd.n2870 99.6594
R7224 gnd.n2950 gnd.n2871 99.6594
R7225 gnd.n2946 gnd.n2872 99.6594
R7226 gnd.n2942 gnd.n2873 99.6594
R7227 gnd.n2938 gnd.n2874 99.6594
R7228 gnd.n2934 gnd.n2875 99.6594
R7229 gnd.n2930 gnd.n2876 99.6594
R7230 gnd.n2926 gnd.n2877 99.6594
R7231 gnd.n2922 gnd.n2878 99.6594
R7232 gnd.n2918 gnd.n2879 99.6594
R7233 gnd.n2914 gnd.n2880 99.6594
R7234 gnd.n2961 gnd.n2869 99.6594
R7235 gnd.n7512 gnd.n7511 99.6594
R7236 gnd.n7517 gnd.n7516 99.6594
R7237 gnd.n7520 gnd.n7519 99.6594
R7238 gnd.n7525 gnd.n7524 99.6594
R7239 gnd.n7528 gnd.n7527 99.6594
R7240 gnd.n7533 gnd.n7532 99.6594
R7241 gnd.n7536 gnd.n7535 99.6594
R7242 gnd.n7541 gnd.n7539 99.6594
R7243 gnd.n7667 gnd.n125 99.6594
R7244 gnd.n1339 gnd.n1275 99.6594
R7245 gnd.n1523 gnd.n1276 99.6594
R7246 gnd.n1525 gnd.n1277 99.6594
R7247 gnd.n1542 gnd.n1278 99.6594
R7248 gnd.n1544 gnd.n1279 99.6594
R7249 gnd.n1561 gnd.n1280 99.6594
R7250 gnd.n1563 gnd.n1281 99.6594
R7251 gnd.n1579 gnd.n1282 99.6594
R7252 gnd.n1490 gnd.n1283 99.6594
R7253 gnd.n2051 gnd.n2050 99.6594
R7254 gnd.n2052 gnd.n2000 99.6594
R7255 gnd.n2054 gnd.n2008 99.6594
R7256 gnd.n2056 gnd.n2055 99.6594
R7257 gnd.n2057 gnd.n2017 99.6594
R7258 gnd.n2059 gnd.n2026 99.6594
R7259 gnd.n2061 gnd.n2060 99.6594
R7260 gnd.n2062 gnd.n2035 99.6594
R7261 gnd.n4849 gnd.n4848 99.6594
R7262 gnd.n3838 gnd.n2338 99.6594
R7263 gnd.n3841 gnd.n3840 99.6594
R7264 gnd.n3848 gnd.n3847 99.6594
R7265 gnd.n3851 gnd.n3850 99.6594
R7266 gnd.n3858 gnd.n3857 99.6594
R7267 gnd.n3861 gnd.n3860 99.6594
R7268 gnd.n3868 gnd.n3867 99.6594
R7269 gnd.n3871 gnd.n3870 99.6594
R7270 gnd.n3878 gnd.n3877 99.6594
R7271 gnd.n3839 gnd.n3838 99.6594
R7272 gnd.n3840 gnd.n3833 99.6594
R7273 gnd.n3849 gnd.n3848 99.6594
R7274 gnd.n3850 gnd.n3829 99.6594
R7275 gnd.n3859 gnd.n3858 99.6594
R7276 gnd.n3860 gnd.n3825 99.6594
R7277 gnd.n3869 gnd.n3868 99.6594
R7278 gnd.n3870 gnd.n3821 99.6594
R7279 gnd.n3879 gnd.n3878 99.6594
R7280 gnd.n4848 gnd.n2046 99.6594
R7281 gnd.n2062 gnd.n2034 99.6594
R7282 gnd.n2061 gnd.n2027 99.6594
R7283 gnd.n2059 gnd.n2058 99.6594
R7284 gnd.n2057 gnd.n2016 99.6594
R7285 gnd.n2056 gnd.n2009 99.6594
R7286 gnd.n2054 gnd.n2053 99.6594
R7287 gnd.n2052 gnd.n1999 99.6594
R7288 gnd.n2051 gnd.n2049 99.6594
R7289 gnd.n1522 gnd.n1275 99.6594
R7290 gnd.n1526 gnd.n1276 99.6594
R7291 gnd.n1541 gnd.n1277 99.6594
R7292 gnd.n1545 gnd.n1278 99.6594
R7293 gnd.n1560 gnd.n1279 99.6594
R7294 gnd.n1564 gnd.n1280 99.6594
R7295 gnd.n1578 gnd.n1281 99.6594
R7296 gnd.n1489 gnd.n1282 99.6594
R7297 gnd.n1485 gnd.n1283 99.6594
R7298 gnd.n7540 gnd.n125 99.6594
R7299 gnd.n7539 gnd.n7538 99.6594
R7300 gnd.n7535 gnd.n7534 99.6594
R7301 gnd.n7532 gnd.n7531 99.6594
R7302 gnd.n7527 gnd.n7526 99.6594
R7303 gnd.n7524 gnd.n7523 99.6594
R7304 gnd.n7519 gnd.n7518 99.6594
R7305 gnd.n7516 gnd.n7515 99.6594
R7306 gnd.n7511 gnd.n7510 99.6594
R7307 gnd.n2959 gnd.n2882 99.6594
R7308 gnd.n2951 gnd.n2870 99.6594
R7309 gnd.n2947 gnd.n2871 99.6594
R7310 gnd.n2943 gnd.n2872 99.6594
R7311 gnd.n2939 gnd.n2873 99.6594
R7312 gnd.n2935 gnd.n2874 99.6594
R7313 gnd.n2931 gnd.n2875 99.6594
R7314 gnd.n2927 gnd.n2876 99.6594
R7315 gnd.n2923 gnd.n2877 99.6594
R7316 gnd.n2919 gnd.n2878 99.6594
R7317 gnd.n2915 gnd.n2879 99.6594
R7318 gnd.n2911 gnd.n2880 99.6594
R7319 gnd.n2962 gnd.n2961 99.6594
R7320 gnd.n3726 gnd.n2352 99.6594
R7321 gnd.n3730 gnd.n2351 99.6594
R7322 gnd.n3734 gnd.n2350 99.6594
R7323 gnd.n3738 gnd.n2349 99.6594
R7324 gnd.n3742 gnd.n2348 99.6594
R7325 gnd.n3746 gnd.n2347 99.6594
R7326 gnd.n3750 gnd.n2346 99.6594
R7327 gnd.n3754 gnd.n2345 99.6594
R7328 gnd.n3758 gnd.n2344 99.6594
R7329 gnd.n3762 gnd.n2343 99.6594
R7330 gnd.n3766 gnd.n2342 99.6594
R7331 gnd.n3770 gnd.n2341 99.6594
R7332 gnd.n2381 gnd.n2340 99.6594
R7333 gnd.n3045 gnd.n3044 99.6594
R7334 gnd.n2804 gnd.n2782 99.6594
R7335 gnd.n2810 gnd.n2783 99.6594
R7336 gnd.n2814 gnd.n2784 99.6594
R7337 gnd.n2820 gnd.n2785 99.6594
R7338 gnd.n2824 gnd.n2786 99.6594
R7339 gnd.n2830 gnd.n2787 99.6594
R7340 gnd.n2788 gnd.n2772 99.6594
R7341 gnd.n3780 gnd.n2353 99.6594
R7342 gnd.n3784 gnd.n2354 99.6594
R7343 gnd.n3788 gnd.n2355 99.6594
R7344 gnd.n3792 gnd.n2356 99.6594
R7345 gnd.n3796 gnd.n2357 99.6594
R7346 gnd.n3800 gnd.n2358 99.6594
R7347 gnd.n3804 gnd.n2359 99.6594
R7348 gnd.n2362 gnd.n2360 99.6594
R7349 gnd.n4192 gnd.n4191 99.6594
R7350 gnd.n4186 gnd.n3981 99.6594
R7351 gnd.n4184 gnd.n4183 99.6594
R7352 gnd.n4179 gnd.n4178 99.6594
R7353 gnd.n4176 gnd.n4175 99.6594
R7354 gnd.n4171 gnd.n4170 99.6594
R7355 gnd.n4168 gnd.n4167 99.6594
R7356 gnd.n4163 gnd.n4162 99.6594
R7357 gnd.n4160 gnd.n4159 99.6594
R7358 gnd.n4155 gnd.n4154 99.6594
R7359 gnd.n4152 gnd.n4151 99.6594
R7360 gnd.n4147 gnd.n4146 99.6594
R7361 gnd.n4144 gnd.n4143 99.6594
R7362 gnd.n4139 gnd.n4138 99.6594
R7363 gnd.n4136 gnd.n4135 99.6594
R7364 gnd.n4131 gnd.n4130 99.6594
R7365 gnd.n4128 gnd.n4127 99.6594
R7366 gnd.n4036 gnd.n4035 99.6594
R7367 gnd.n4119 gnd.n4118 99.6594
R7368 gnd.n4576 gnd.n2064 99.6594
R7369 gnd.n4580 gnd.n2065 99.6594
R7370 gnd.n4584 gnd.n2066 99.6594
R7371 gnd.n4588 gnd.n2067 99.6594
R7372 gnd.n4592 gnd.n2068 99.6594
R7373 gnd.n4596 gnd.n2069 99.6594
R7374 gnd.n4600 gnd.n2070 99.6594
R7375 gnd.n4604 gnd.n2071 99.6594
R7376 gnd.n4608 gnd.n2072 99.6594
R7377 gnd.n4612 gnd.n2073 99.6594
R7378 gnd.n4820 gnd.n2075 99.6594
R7379 gnd.n4824 gnd.n2076 99.6594
R7380 gnd.n4828 gnd.n2077 99.6594
R7381 gnd.n4832 gnd.n2078 99.6594
R7382 gnd.n4836 gnd.n2079 99.6594
R7383 gnd.n4840 gnd.n2080 99.6594
R7384 gnd.n2083 gnd.n2081 99.6594
R7385 gnd.n4846 gnd.n2082 99.6594
R7386 gnd.n6154 gnd.n1287 99.6594
R7387 gnd.n6146 gnd.n1257 99.6594
R7388 gnd.n6142 gnd.n1258 99.6594
R7389 gnd.n6138 gnd.n1259 99.6594
R7390 gnd.n6134 gnd.n1260 99.6594
R7391 gnd.n6130 gnd.n1261 99.6594
R7392 gnd.n6126 gnd.n1262 99.6594
R7393 gnd.n6121 gnd.n1264 99.6594
R7394 gnd.n6117 gnd.n1265 99.6594
R7395 gnd.n6113 gnd.n1266 99.6594
R7396 gnd.n6109 gnd.n1267 99.6594
R7397 gnd.n6105 gnd.n1268 99.6594
R7398 gnd.n6101 gnd.n1269 99.6594
R7399 gnd.n6097 gnd.n1270 99.6594
R7400 gnd.n6093 gnd.n1271 99.6594
R7401 gnd.n6089 gnd.n1272 99.6594
R7402 gnd.n1328 gnd.n1273 99.6594
R7403 gnd.n6081 gnd.n1274 99.6594
R7404 gnd.n198 gnd.n195 99.6594
R7405 gnd.n7597 gnd.n7596 99.6594
R7406 gnd.n194 gnd.n188 99.6594
R7407 gnd.n7604 gnd.n7603 99.6594
R7408 gnd.n187 gnd.n181 99.6594
R7409 gnd.n7611 gnd.n7610 99.6594
R7410 gnd.n180 gnd.n174 99.6594
R7411 gnd.n7618 gnd.n7617 99.6594
R7412 gnd.n173 gnd.n167 99.6594
R7413 gnd.n7625 gnd.n7624 99.6594
R7414 gnd.n166 gnd.n160 99.6594
R7415 gnd.n7635 gnd.n7634 99.6594
R7416 gnd.n159 gnd.n153 99.6594
R7417 gnd.n7642 gnd.n7641 99.6594
R7418 gnd.n152 gnd.n146 99.6594
R7419 gnd.n7649 gnd.n7648 99.6594
R7420 gnd.n145 gnd.n139 99.6594
R7421 gnd.n7656 gnd.n7655 99.6594
R7422 gnd.n138 gnd.n135 99.6594
R7423 gnd.n4896 gnd.n4895 99.6594
R7424 gnd.n2003 gnd.n1980 99.6594
R7425 gnd.n2005 gnd.n1981 99.6594
R7426 gnd.n2013 gnd.n1982 99.6594
R7427 gnd.n2021 gnd.n1983 99.6594
R7428 gnd.n2023 gnd.n1984 99.6594
R7429 gnd.n2031 gnd.n1985 99.6594
R7430 gnd.n2041 gnd.n1986 99.6594
R7431 gnd.n2043 gnd.n1987 99.6594
R7432 gnd.n4537 gnd.n1988 99.6594
R7433 gnd.n4539 gnd.n1989 99.6594
R7434 gnd.n4543 gnd.n1990 99.6594
R7435 gnd.n4549 gnd.n1991 99.6594
R7436 gnd.n4899 gnd.n4898 99.6594
R7437 gnd.n4896 gnd.n1993 99.6594
R7438 gnd.n2004 gnd.n1980 99.6594
R7439 gnd.n2012 gnd.n1981 99.6594
R7440 gnd.n2020 gnd.n1982 99.6594
R7441 gnd.n2022 gnd.n1983 99.6594
R7442 gnd.n2030 gnd.n1984 99.6594
R7443 gnd.n2040 gnd.n1985 99.6594
R7444 gnd.n2042 gnd.n1986 99.6594
R7445 gnd.n4536 gnd.n1987 99.6594
R7446 gnd.n4538 gnd.n1988 99.6594
R7447 gnd.n4542 gnd.n1989 99.6594
R7448 gnd.n4544 gnd.n1990 99.6594
R7449 gnd.n1991 gnd.n1978 99.6594
R7450 gnd.n4898 gnd.n1975 99.6594
R7451 gnd.n1531 gnd.n1513 99.6594
R7452 gnd.n1535 gnd.n1533 99.6594
R7453 gnd.n1550 gnd.n1506 99.6594
R7454 gnd.n1554 gnd.n1552 99.6594
R7455 gnd.n1569 gnd.n1499 99.6594
R7456 gnd.n1573 gnd.n1571 99.6594
R7457 gnd.n1585 gnd.n1493 99.6594
R7458 gnd.n1589 gnd.n1587 99.6594
R7459 gnd.n1599 gnd.n1481 99.6594
R7460 gnd.n1602 gnd.n1601 99.6594
R7461 gnd.n1605 gnd.n1604 99.6594
R7462 gnd.n1610 gnd.n1609 99.6594
R7463 gnd.n1613 gnd.n1612 99.6594
R7464 gnd.n5882 gnd.n5881 99.6594
R7465 gnd.n5881 gnd.n5880 99.6594
R7466 gnd.n1612 gnd.n1611 99.6594
R7467 gnd.n1609 gnd.n1608 99.6594
R7468 gnd.n1604 gnd.n1603 99.6594
R7469 gnd.n1601 gnd.n1600 99.6594
R7470 gnd.n1588 gnd.n1481 99.6594
R7471 gnd.n1587 gnd.n1586 99.6594
R7472 gnd.n1572 gnd.n1493 99.6594
R7473 gnd.n1571 gnd.n1570 99.6594
R7474 gnd.n1553 gnd.n1499 99.6594
R7475 gnd.n1552 gnd.n1551 99.6594
R7476 gnd.n1534 gnd.n1506 99.6594
R7477 gnd.n1533 gnd.n1532 99.6594
R7478 gnd.n1513 gnd.n1244 99.6594
R7479 gnd.n4545 gnd.t268 98.63
R7480 gnd.n122 gnd.t280 98.63
R7481 gnd.n1486 gnd.t293 98.63
R7482 gnd.n2036 gnd.t316 98.63
R7483 gnd.n1308 gnd.t264 98.63
R7484 gnd.n1330 gnd.t243 98.63
R7485 gnd.n201 gnd.t309 98.63
R7486 gnd.n7628 gnd.t224 98.63
R7487 gnd.n4005 gnd.t326 98.63
R7488 gnd.n4037 gnd.t307 98.63
R7489 gnd.n3818 gnd.t323 98.63
R7490 gnd.n2125 gnd.t319 98.63
R7491 gnd.n2103 gnd.t238 98.63
R7492 gnd.n5890 gnd.t234 98.63
R7493 gnd.n4621 gnd.t300 92.8196
R7494 gnd.n5231 gnd.t253 92.8196
R7495 gnd.n4677 gnd.t247 92.8118
R7496 gnd.n5225 gnd.t289 92.8118
R7497 gnd.n7004 gnd.n7003 84.8607
R7498 gnd.n7005 gnd.n7004 84.8607
R7499 gnd.n7005 gnd.n540 84.8607
R7500 gnd.n7013 gnd.n540 84.8607
R7501 gnd.n7014 gnd.n7013 84.8607
R7502 gnd.n7015 gnd.n7014 84.8607
R7503 gnd.n7015 gnd.n534 84.8607
R7504 gnd.n7023 gnd.n534 84.8607
R7505 gnd.n7024 gnd.n7023 84.8607
R7506 gnd.n7025 gnd.n7024 84.8607
R7507 gnd.n7025 gnd.n528 84.8607
R7508 gnd.n7033 gnd.n528 84.8607
R7509 gnd.n7034 gnd.n7033 84.8607
R7510 gnd.n7035 gnd.n7034 84.8607
R7511 gnd.n7035 gnd.n522 84.8607
R7512 gnd.n7043 gnd.n522 84.8607
R7513 gnd.n7044 gnd.n7043 84.8607
R7514 gnd.n7045 gnd.n7044 84.8607
R7515 gnd.n7045 gnd.n516 84.8607
R7516 gnd.n7053 gnd.n516 84.8607
R7517 gnd.n7054 gnd.n7053 84.8607
R7518 gnd.n7055 gnd.n7054 84.8607
R7519 gnd.n7055 gnd.n510 84.8607
R7520 gnd.n7063 gnd.n510 84.8607
R7521 gnd.n7064 gnd.n7063 84.8607
R7522 gnd.n7065 gnd.n7064 84.8607
R7523 gnd.n7065 gnd.n504 84.8607
R7524 gnd.n7073 gnd.n504 84.8607
R7525 gnd.n7074 gnd.n7073 84.8607
R7526 gnd.n7075 gnd.n7074 84.8607
R7527 gnd.n7075 gnd.n498 84.8607
R7528 gnd.n7083 gnd.n498 84.8607
R7529 gnd.n7084 gnd.n7083 84.8607
R7530 gnd.n7085 gnd.n7084 84.8607
R7531 gnd.n7085 gnd.n492 84.8607
R7532 gnd.n7093 gnd.n492 84.8607
R7533 gnd.n7094 gnd.n7093 84.8607
R7534 gnd.n7095 gnd.n7094 84.8607
R7535 gnd.n7095 gnd.n486 84.8607
R7536 gnd.n7103 gnd.n486 84.8607
R7537 gnd.n7104 gnd.n7103 84.8607
R7538 gnd.n7105 gnd.n7104 84.8607
R7539 gnd.n7105 gnd.n480 84.8607
R7540 gnd.n7113 gnd.n480 84.8607
R7541 gnd.n7114 gnd.n7113 84.8607
R7542 gnd.n7115 gnd.n7114 84.8607
R7543 gnd.n7115 gnd.n474 84.8607
R7544 gnd.n7123 gnd.n474 84.8607
R7545 gnd.n7124 gnd.n7123 84.8607
R7546 gnd.n7125 gnd.n7124 84.8607
R7547 gnd.n7125 gnd.n468 84.8607
R7548 gnd.n7133 gnd.n468 84.8607
R7549 gnd.n7134 gnd.n7133 84.8607
R7550 gnd.n7135 gnd.n7134 84.8607
R7551 gnd.n7135 gnd.n462 84.8607
R7552 gnd.n7143 gnd.n462 84.8607
R7553 gnd.n7144 gnd.n7143 84.8607
R7554 gnd.n7145 gnd.n7144 84.8607
R7555 gnd.n7145 gnd.n456 84.8607
R7556 gnd.n7153 gnd.n456 84.8607
R7557 gnd.n7154 gnd.n7153 84.8607
R7558 gnd.n7155 gnd.n7154 84.8607
R7559 gnd.n7155 gnd.n450 84.8607
R7560 gnd.n7163 gnd.n450 84.8607
R7561 gnd.n7164 gnd.n7163 84.8607
R7562 gnd.n7165 gnd.n7164 84.8607
R7563 gnd.n7165 gnd.n444 84.8607
R7564 gnd.n7173 gnd.n444 84.8607
R7565 gnd.n7174 gnd.n7173 84.8607
R7566 gnd.n7175 gnd.n7174 84.8607
R7567 gnd.n7175 gnd.n438 84.8607
R7568 gnd.n7183 gnd.n438 84.8607
R7569 gnd.n7184 gnd.n7183 84.8607
R7570 gnd.n7185 gnd.n7184 84.8607
R7571 gnd.n7185 gnd.n432 84.8607
R7572 gnd.n7193 gnd.n432 84.8607
R7573 gnd.n7194 gnd.n7193 84.8607
R7574 gnd.n7195 gnd.n7194 84.8607
R7575 gnd.n7195 gnd.n426 84.8607
R7576 gnd.n7203 gnd.n426 84.8607
R7577 gnd.n7204 gnd.n7203 84.8607
R7578 gnd.n7206 gnd.n7204 84.8607
R7579 gnd.n7206 gnd.n7205 84.8607
R7580 gnd.n4652 gnd.n4651 81.8399
R7581 gnd.n2833 gnd.t313 74.8376
R7582 gnd.n2378 gnd.t258 74.8376
R7583 gnd.n4622 gnd.t299 72.8438
R7584 gnd.n5232 gnd.t254 72.8438
R7585 gnd.n4653 gnd.n4646 72.8411
R7586 gnd.n4659 gnd.n4644 72.8411
R7587 gnd.n5200 gnd.n5199 72.8411
R7588 gnd.n4546 gnd.t267 72.836
R7589 gnd.n4678 gnd.t246 72.836
R7590 gnd.n5226 gnd.t290 72.836
R7591 gnd.n123 gnd.t281 72.836
R7592 gnd.n1487 gnd.t292 72.836
R7593 gnd.n2037 gnd.t317 72.836
R7594 gnd.n1309 gnd.t263 72.836
R7595 gnd.n1331 gnd.t242 72.836
R7596 gnd.n202 gnd.t310 72.836
R7597 gnd.n7629 gnd.t225 72.836
R7598 gnd.n4006 gnd.t325 72.836
R7599 gnd.n4038 gnd.t306 72.836
R7600 gnd.n3819 gnd.t322 72.836
R7601 gnd.n2126 gnd.t320 72.836
R7602 gnd.n2104 gnd.t239 72.836
R7603 gnd.n5891 gnd.t235 72.836
R7604 gnd.n5371 gnd.n5370 71.676
R7605 gnd.n5368 gnd.n5367 71.676
R7606 gnd.n5363 gnd.n5208 71.676
R7607 gnd.n5361 gnd.n5360 71.676
R7608 gnd.n5356 gnd.n5211 71.676
R7609 gnd.n5354 gnd.n5353 71.676
R7610 gnd.n5349 gnd.n5214 71.676
R7611 gnd.n5347 gnd.n5346 71.676
R7612 gnd.n5342 gnd.n5217 71.676
R7613 gnd.n5340 gnd.n5339 71.676
R7614 gnd.n5335 gnd.n5220 71.676
R7615 gnd.n5333 gnd.n5332 71.676
R7616 gnd.n5328 gnd.n5223 71.676
R7617 gnd.n5326 gnd.n5325 71.676
R7618 gnd.n5320 gnd.n5228 71.676
R7619 gnd.n5318 gnd.n5317 71.676
R7620 gnd.n5313 gnd.n5312 71.676
R7621 gnd.n5310 gnd.n5309 71.676
R7622 gnd.n5304 gnd.n5234 71.676
R7623 gnd.n5302 gnd.n5301 71.676
R7624 gnd.n5297 gnd.n5237 71.676
R7625 gnd.n5295 gnd.n5294 71.676
R7626 gnd.n5290 gnd.n5240 71.676
R7627 gnd.n5288 gnd.n5287 71.676
R7628 gnd.n5283 gnd.n5243 71.676
R7629 gnd.n5281 gnd.n5280 71.676
R7630 gnd.n5276 gnd.n5246 71.676
R7631 gnd.n5274 gnd.n5273 71.676
R7632 gnd.n5269 gnd.n5249 71.676
R7633 gnd.n5267 gnd.n5266 71.676
R7634 gnd.n5262 gnd.n5252 71.676
R7635 gnd.n5260 gnd.n5259 71.676
R7636 gnd.n5255 gnd.n5254 71.676
R7637 gnd.n4740 gnd.n4642 71.676
R7638 gnd.n4738 gnd.n4664 71.676
R7639 gnd.n4734 gnd.n4733 71.676
R7640 gnd.n4727 gnd.n4666 71.676
R7641 gnd.n4726 gnd.n4725 71.676
R7642 gnd.n4719 gnd.n4668 71.676
R7643 gnd.n4718 gnd.n4717 71.676
R7644 gnd.n4711 gnd.n4670 71.676
R7645 gnd.n4710 gnd.n4709 71.676
R7646 gnd.n4703 gnd.n4672 71.676
R7647 gnd.n4702 gnd.n4701 71.676
R7648 gnd.n4695 gnd.n4674 71.676
R7649 gnd.n4694 gnd.n4693 71.676
R7650 gnd.n4687 gnd.n4676 71.676
R7651 gnd.n4686 gnd.n4680 71.676
R7652 gnd.n4682 gnd.n4681 71.676
R7653 gnd.n4814 gnd.n4813 71.676
R7654 gnd.n4806 gnd.n4620 71.676
R7655 gnd.n4805 gnd.n4804 71.676
R7656 gnd.n4798 gnd.n4624 71.676
R7657 gnd.n4797 gnd.n4796 71.676
R7658 gnd.n4790 gnd.n4626 71.676
R7659 gnd.n4789 gnd.n4788 71.676
R7660 gnd.n4782 gnd.n4628 71.676
R7661 gnd.n4781 gnd.n4780 71.676
R7662 gnd.n4774 gnd.n4630 71.676
R7663 gnd.n4773 gnd.n4772 71.676
R7664 gnd.n4766 gnd.n4632 71.676
R7665 gnd.n4765 gnd.n4764 71.676
R7666 gnd.n4758 gnd.n4634 71.676
R7667 gnd.n4757 gnd.n4756 71.676
R7668 gnd.n4750 gnd.n4636 71.676
R7669 gnd.n4741 gnd.n4740 71.676
R7670 gnd.n4735 gnd.n4664 71.676
R7671 gnd.n4733 gnd.n4732 71.676
R7672 gnd.n4728 gnd.n4727 71.676
R7673 gnd.n4725 gnd.n4724 71.676
R7674 gnd.n4720 gnd.n4719 71.676
R7675 gnd.n4717 gnd.n4716 71.676
R7676 gnd.n4712 gnd.n4711 71.676
R7677 gnd.n4709 gnd.n4708 71.676
R7678 gnd.n4704 gnd.n4703 71.676
R7679 gnd.n4701 gnd.n4700 71.676
R7680 gnd.n4696 gnd.n4695 71.676
R7681 gnd.n4693 gnd.n4692 71.676
R7682 gnd.n4688 gnd.n4687 71.676
R7683 gnd.n4683 gnd.n4680 71.676
R7684 gnd.n4816 gnd.n4815 71.676
R7685 gnd.n4813 gnd.n4812 71.676
R7686 gnd.n4807 gnd.n4806 71.676
R7687 gnd.n4804 gnd.n4803 71.676
R7688 gnd.n4799 gnd.n4798 71.676
R7689 gnd.n4796 gnd.n4795 71.676
R7690 gnd.n4791 gnd.n4790 71.676
R7691 gnd.n4788 gnd.n4787 71.676
R7692 gnd.n4783 gnd.n4782 71.676
R7693 gnd.n4780 gnd.n4779 71.676
R7694 gnd.n4775 gnd.n4774 71.676
R7695 gnd.n4772 gnd.n4771 71.676
R7696 gnd.n4767 gnd.n4766 71.676
R7697 gnd.n4764 gnd.n4763 71.676
R7698 gnd.n4759 gnd.n4758 71.676
R7699 gnd.n4756 gnd.n4755 71.676
R7700 gnd.n4751 gnd.n4750 71.676
R7701 gnd.n5254 gnd.n5253 71.676
R7702 gnd.n5261 gnd.n5260 71.676
R7703 gnd.n5252 gnd.n5250 71.676
R7704 gnd.n5268 gnd.n5267 71.676
R7705 gnd.n5249 gnd.n5247 71.676
R7706 gnd.n5275 gnd.n5274 71.676
R7707 gnd.n5246 gnd.n5244 71.676
R7708 gnd.n5282 gnd.n5281 71.676
R7709 gnd.n5243 gnd.n5241 71.676
R7710 gnd.n5289 gnd.n5288 71.676
R7711 gnd.n5240 gnd.n5238 71.676
R7712 gnd.n5296 gnd.n5295 71.676
R7713 gnd.n5237 gnd.n5235 71.676
R7714 gnd.n5303 gnd.n5302 71.676
R7715 gnd.n5234 gnd.n5230 71.676
R7716 gnd.n5311 gnd.n5310 71.676
R7717 gnd.n5315 gnd.n5314 71.676
R7718 gnd.n5319 gnd.n5318 71.676
R7719 gnd.n5228 gnd.n5224 71.676
R7720 gnd.n5327 gnd.n5326 71.676
R7721 gnd.n5223 gnd.n5221 71.676
R7722 gnd.n5334 gnd.n5333 71.676
R7723 gnd.n5220 gnd.n5218 71.676
R7724 gnd.n5341 gnd.n5340 71.676
R7725 gnd.n5217 gnd.n5215 71.676
R7726 gnd.n5348 gnd.n5347 71.676
R7727 gnd.n5214 gnd.n5212 71.676
R7728 gnd.n5355 gnd.n5354 71.676
R7729 gnd.n5211 gnd.n5209 71.676
R7730 gnd.n5362 gnd.n5361 71.676
R7731 gnd.n5208 gnd.n5206 71.676
R7732 gnd.n5369 gnd.n5368 71.676
R7733 gnd.n5372 gnd.n5371 71.676
R7734 gnd.n10 gnd.t206 69.1507
R7735 gnd.n18 gnd.t217 68.4792
R7736 gnd.n17 gnd.t156 68.4792
R7737 gnd.n16 gnd.t219 68.4792
R7738 gnd.n15 gnd.t359 68.4792
R7739 gnd.n14 gnd.t111 68.4792
R7740 gnd.n13 gnd.t353 68.4792
R7741 gnd.n12 gnd.t109 68.4792
R7742 gnd.n11 gnd.t120 68.4792
R7743 gnd.n10 gnd.t123 68.4792
R7744 gnd.n2960 gnd.n2864 64.369
R7745 gnd.n4809 gnd.n4622 59.5399
R7746 gnd.n5306 gnd.n5232 59.5399
R7747 gnd.n4679 gnd.n4678 59.5399
R7748 gnd.n5322 gnd.n5226 59.5399
R7749 gnd.n4744 gnd.n4662 59.1804
R7750 gnd.n2611 gnd.t107 56.607
R7751 gnd.n60 gnd.t339 56.607
R7752 gnd.n2572 gnd.t335 56.407
R7753 gnd.n2591 gnd.t173 56.407
R7754 gnd.n21 gnd.t12 56.407
R7755 gnd.n40 gnd.t133 56.407
R7756 gnd.n2628 gnd.t144 55.8337
R7757 gnd.n2589 gnd.t346 55.8337
R7758 gnd.n2608 gnd.t334 55.8337
R7759 gnd.n77 gnd.t15 55.8337
R7760 gnd.n38 gnd.t14 55.8337
R7761 gnd.n57 gnd.t130 55.8337
R7762 gnd.n4650 gnd.n4649 54.358
R7763 gnd.n5197 gnd.n5196 54.358
R7764 gnd.n2611 gnd.n2610 53.0052
R7765 gnd.n2613 gnd.n2612 53.0052
R7766 gnd.n2615 gnd.n2614 53.0052
R7767 gnd.n2617 gnd.n2616 53.0052
R7768 gnd.n2619 gnd.n2618 53.0052
R7769 gnd.n2621 gnd.n2620 53.0052
R7770 gnd.n2623 gnd.n2622 53.0052
R7771 gnd.n2625 gnd.n2624 53.0052
R7772 gnd.n2627 gnd.n2626 53.0052
R7773 gnd.n2572 gnd.n2571 53.0052
R7774 gnd.n2574 gnd.n2573 53.0052
R7775 gnd.n2576 gnd.n2575 53.0052
R7776 gnd.n2578 gnd.n2577 53.0052
R7777 gnd.n2580 gnd.n2579 53.0052
R7778 gnd.n2582 gnd.n2581 53.0052
R7779 gnd.n2584 gnd.n2583 53.0052
R7780 gnd.n2586 gnd.n2585 53.0052
R7781 gnd.n2588 gnd.n2587 53.0052
R7782 gnd.n2591 gnd.n2590 53.0052
R7783 gnd.n2593 gnd.n2592 53.0052
R7784 gnd.n2595 gnd.n2594 53.0052
R7785 gnd.n2597 gnd.n2596 53.0052
R7786 gnd.n2599 gnd.n2598 53.0052
R7787 gnd.n2601 gnd.n2600 53.0052
R7788 gnd.n2603 gnd.n2602 53.0052
R7789 gnd.n2605 gnd.n2604 53.0052
R7790 gnd.n2607 gnd.n2606 53.0052
R7791 gnd.n76 gnd.n75 53.0052
R7792 gnd.n74 gnd.n73 53.0052
R7793 gnd.n72 gnd.n71 53.0052
R7794 gnd.n70 gnd.n69 53.0052
R7795 gnd.n68 gnd.n67 53.0052
R7796 gnd.n66 gnd.n65 53.0052
R7797 gnd.n64 gnd.n63 53.0052
R7798 gnd.n62 gnd.n61 53.0052
R7799 gnd.n60 gnd.n59 53.0052
R7800 gnd.n37 gnd.n36 53.0052
R7801 gnd.n35 gnd.n34 53.0052
R7802 gnd.n33 gnd.n32 53.0052
R7803 gnd.n31 gnd.n30 53.0052
R7804 gnd.n29 gnd.n28 53.0052
R7805 gnd.n27 gnd.n26 53.0052
R7806 gnd.n25 gnd.n24 53.0052
R7807 gnd.n23 gnd.n22 53.0052
R7808 gnd.n21 gnd.n20 53.0052
R7809 gnd.n56 gnd.n55 53.0052
R7810 gnd.n54 gnd.n53 53.0052
R7811 gnd.n52 gnd.n51 53.0052
R7812 gnd.n50 gnd.n49 53.0052
R7813 gnd.n48 gnd.n47 53.0052
R7814 gnd.n46 gnd.n45 53.0052
R7815 gnd.n44 gnd.n43 53.0052
R7816 gnd.n42 gnd.n41 53.0052
R7817 gnd.n40 gnd.n39 53.0052
R7818 gnd.n5188 gnd.n5187 52.4801
R7819 gnd.n3664 gnd.t117 52.3082
R7820 gnd.n3632 gnd.t40 52.3082
R7821 gnd.n3600 gnd.t168 52.3082
R7822 gnd.n3569 gnd.t4 52.3082
R7823 gnd.n3537 gnd.t341 52.3082
R7824 gnd.n3505 gnd.t331 52.3082
R7825 gnd.n3473 gnd.t158 52.3082
R7826 gnd.n3442 gnd.t170 52.3082
R7827 gnd.n4199 gnd.n3813 51.6227
R7828 gnd.n7665 gnd.n128 51.6227
R7829 gnd.n3494 gnd.n3462 51.4173
R7830 gnd.n7205 gnd.n238 50.9166
R7831 gnd.n3558 gnd.n3557 50.455
R7832 gnd.n3526 gnd.n3525 50.455
R7833 gnd.n3494 gnd.n3493 50.455
R7834 gnd.n2907 gnd.n2906 45.1884
R7835 gnd.n2404 gnd.n2403 45.1884
R7836 gnd.n5374 gnd.n5203 44.3322
R7837 gnd.n4653 gnd.n4652 44.3189
R7838 gnd.n4547 gnd.n4546 42.4732
R7839 gnd.n5892 gnd.n5891 42.4732
R7840 gnd.n2908 gnd.n2907 42.2793
R7841 gnd.n2405 gnd.n2404 42.2793
R7842 gnd.n2834 gnd.n2833 42.2793
R7843 gnd.n3779 gnd.n2378 42.2793
R7844 gnd.n124 gnd.n123 42.2793
R7845 gnd.n1594 gnd.n1487 42.2793
R7846 gnd.n2038 gnd.n2037 42.2793
R7847 gnd.n1332 gnd.n1331 42.2793
R7848 gnd.n7593 gnd.n202 42.2793
R7849 gnd.n7630 gnd.n7629 42.2793
R7850 gnd.n4007 gnd.n4006 42.2793
R7851 gnd.n4039 gnd.n4038 42.2793
R7852 gnd.n3820 gnd.n3819 42.2793
R7853 gnd.n4575 gnd.n2126 42.2793
R7854 gnd.n4651 gnd.n4650 41.6274
R7855 gnd.n5198 gnd.n5197 41.6274
R7856 gnd.n4660 gnd.n4659 40.8975
R7857 gnd.n5201 gnd.n5200 40.8975
R7858 gnd.n6123 gnd.n1309 36.9518
R7859 gnd.n4818 gnd.n2104 36.9518
R7860 gnd.n4659 gnd.n4658 35.055
R7861 gnd.n4654 gnd.n4653 35.055
R7862 gnd.n5190 gnd.n5189 35.055
R7863 gnd.n5200 gnd.n5186 35.055
R7864 gnd.n6574 gnd.n797 31.9958
R7865 gnd.n6574 gnd.n6573 31.9958
R7866 gnd.n6573 gnd.n6572 31.9958
R7867 gnd.n6572 gnd.n802 31.9958
R7868 gnd.n6566 gnd.n802 31.9958
R7869 gnd.n6566 gnd.n6565 31.9958
R7870 gnd.n6565 gnd.n6564 31.9958
R7871 gnd.n6564 gnd.n810 31.9958
R7872 gnd.n6558 gnd.n810 31.9958
R7873 gnd.n6558 gnd.n6557 31.9958
R7874 gnd.n6557 gnd.n6556 31.9958
R7875 gnd.n6556 gnd.n818 31.9958
R7876 gnd.n6550 gnd.n818 31.9958
R7877 gnd.n6550 gnd.n6549 31.9958
R7878 gnd.n6549 gnd.n6548 31.9958
R7879 gnd.n6548 gnd.n826 31.9958
R7880 gnd.n6542 gnd.n826 31.9958
R7881 gnd.n6542 gnd.n6541 31.9958
R7882 gnd.n6541 gnd.n6540 31.9958
R7883 gnd.n6540 gnd.n834 31.9958
R7884 gnd.n6534 gnd.n834 31.9958
R7885 gnd.n6534 gnd.n6533 31.9958
R7886 gnd.n6533 gnd.n6532 31.9958
R7887 gnd.n6532 gnd.n842 31.9958
R7888 gnd.n6526 gnd.n842 31.9958
R7889 gnd.n6526 gnd.n6525 31.9958
R7890 gnd.n6525 gnd.n6524 31.9958
R7891 gnd.n6524 gnd.n850 31.9958
R7892 gnd.n6518 gnd.n850 31.9958
R7893 gnd.n6518 gnd.n6517 31.9958
R7894 gnd.n6517 gnd.n6516 31.9958
R7895 gnd.n6516 gnd.n858 31.9958
R7896 gnd.n6510 gnd.n858 31.9958
R7897 gnd.n6510 gnd.n6509 31.9958
R7898 gnd.n6509 gnd.n6508 31.9958
R7899 gnd.n6508 gnd.n866 31.9958
R7900 gnd.n6502 gnd.n866 31.9958
R7901 gnd.n6502 gnd.n6501 31.9958
R7902 gnd.n6501 gnd.n6500 31.9958
R7903 gnd.n6500 gnd.n874 31.9958
R7904 gnd.n6494 gnd.n874 31.9958
R7905 gnd.n6494 gnd.n6493 31.9958
R7906 gnd.n6493 gnd.n6492 31.9958
R7907 gnd.n6492 gnd.n882 31.9958
R7908 gnd.n6486 gnd.n882 31.9958
R7909 gnd.n6486 gnd.n6485 31.9958
R7910 gnd.n6485 gnd.n6484 31.9958
R7911 gnd.n6484 gnd.n890 31.9958
R7912 gnd.n6478 gnd.n890 31.9958
R7913 gnd.n6478 gnd.n6477 31.9958
R7914 gnd.n6477 gnd.n6476 31.9958
R7915 gnd.n6476 gnd.n898 31.9958
R7916 gnd.n6470 gnd.n898 31.9958
R7917 gnd.n6470 gnd.n6469 31.9958
R7918 gnd.n6469 gnd.n6468 31.9958
R7919 gnd.n6468 gnd.n906 31.9958
R7920 gnd.n6462 gnd.n906 31.9958
R7921 gnd.n6462 gnd.n6461 31.9958
R7922 gnd.n6461 gnd.n6460 31.9958
R7923 gnd.n6460 gnd.n914 31.9958
R7924 gnd.n6454 gnd.n914 31.9958
R7925 gnd.n6454 gnd.n6453 31.9958
R7926 gnd.n6453 gnd.n6452 31.9958
R7927 gnd.n6452 gnd.n922 31.9958
R7928 gnd.n6446 gnd.n922 31.9958
R7929 gnd.n6446 gnd.n6445 31.9958
R7930 gnd.n6445 gnd.n6444 31.9958
R7931 gnd.n6444 gnd.n930 31.9958
R7932 gnd.n6438 gnd.n930 31.9958
R7933 gnd.n6438 gnd.n6437 31.9958
R7934 gnd.n6437 gnd.n6436 31.9958
R7935 gnd.n6436 gnd.n938 31.9958
R7936 gnd.n6430 gnd.n938 31.9958
R7937 gnd.n6430 gnd.n6429 31.9958
R7938 gnd.n6429 gnd.n6428 31.9958
R7939 gnd.n6428 gnd.n946 31.9958
R7940 gnd.n6422 gnd.n946 31.9958
R7941 gnd.n6422 gnd.n6421 31.9958
R7942 gnd.n6421 gnd.n6420 31.9958
R7943 gnd.n6420 gnd.n954 31.9958
R7944 gnd.n6414 gnd.n954 31.9958
R7945 gnd.n6414 gnd.n6413 31.9958
R7946 gnd.n6413 gnd.n6412 31.9958
R7947 gnd.n2970 gnd.n2864 31.8661
R7948 gnd.n2970 gnd.n2969 31.8661
R7949 gnd.n2978 gnd.n2853 31.8661
R7950 gnd.n2986 gnd.n2853 31.8661
R7951 gnd.n2986 gnd.n2847 31.8661
R7952 gnd.n2994 gnd.n2847 31.8661
R7953 gnd.n2994 gnd.n2840 31.8661
R7954 gnd.n3032 gnd.n2840 31.8661
R7955 gnd.n3042 gnd.n2773 31.8661
R7956 gnd.n4199 gnd.n3977 31.8661
R7957 gnd.n4207 gnd.n2325 31.8661
R7958 gnd.n4215 gnd.n2325 31.8661
R7959 gnd.n4215 gnd.n2317 31.8661
R7960 gnd.n4223 gnd.n2317 31.8661
R7961 gnd.n4231 gnd.n2308 31.8661
R7962 gnd.n4231 gnd.n2311 31.8661
R7963 gnd.n4239 gnd.n2293 31.8661
R7964 gnd.n4247 gnd.n2293 31.8661
R7965 gnd.n4255 gnd.n2285 31.8661
R7966 gnd.n4263 gnd.n2276 31.8661
R7967 gnd.n4263 gnd.n2279 31.8661
R7968 gnd.n4271 gnd.n2261 31.8661
R7969 gnd.n4279 gnd.n2261 31.8661
R7970 gnd.n4287 gnd.n2253 31.8661
R7971 gnd.n4296 gnd.n2244 31.8661
R7972 gnd.n4296 gnd.n2247 31.8661
R7973 gnd.n4304 gnd.n2230 31.8661
R7974 gnd.n4312 gnd.n2230 31.8661
R7975 gnd.n4321 gnd.n2221 31.8661
R7976 gnd.n4329 gnd.n2214 31.8661
R7977 gnd.n4329 gnd.n2216 31.8661
R7978 gnd.n4348 gnd.n2198 31.8661
R7979 gnd.n4355 gnd.n970 31.8661
R7980 gnd.n2047 gnd.n1112 31.8661
R7981 gnd.n4494 gnd.n2063 31.8661
R7982 gnd.n4494 gnd.n1979 31.8661
R7983 gnd.n4906 gnd.n1973 31.8661
R7984 gnd.n4906 gnd.n1974 31.8661
R7985 gnd.n4914 gnd.n1962 31.8661
R7986 gnd.n4922 gnd.n1962 31.8661
R7987 gnd.n4922 gnd.n1955 31.8661
R7988 gnd.n4930 gnd.n1955 31.8661
R7989 gnd.n4938 gnd.n1949 31.8661
R7990 gnd.n4938 gnd.n1940 31.8661
R7991 gnd.n4946 gnd.n1940 31.8661
R7992 gnd.n4946 gnd.n1942 31.8661
R7993 gnd.n4954 gnd.n1927 31.8661
R7994 gnd.n4962 gnd.n1927 31.8661
R7995 gnd.n4962 gnd.n1929 31.8661
R7996 gnd.n4970 gnd.n1916 31.8661
R7997 gnd.n4978 gnd.n1916 31.8661
R7998 gnd.n4978 gnd.n1909 31.8661
R7999 gnd.n4986 gnd.n1909 31.8661
R8000 gnd.n5796 gnd.n1672 31.8661
R8001 gnd.n5804 gnd.n1672 31.8661
R8002 gnd.n5804 gnd.n1666 31.8661
R8003 gnd.n5812 gnd.n1666 31.8661
R8004 gnd.n5820 gnd.n1659 31.8661
R8005 gnd.n5820 gnd.n1653 31.8661
R8006 gnd.n5828 gnd.n1653 31.8661
R8007 gnd.n5836 gnd.n1646 31.8661
R8008 gnd.n5836 gnd.n1639 31.8661
R8009 gnd.n5844 gnd.n1639 31.8661
R8010 gnd.n5844 gnd.n1640 31.8661
R8011 gnd.n5852 gnd.n1626 31.8661
R8012 gnd.n5862 gnd.n1626 31.8661
R8013 gnd.n5862 gnd.n1618 31.8661
R8014 gnd.n5873 gnd.n1618 31.8661
R8015 gnd.n6164 gnd.n1245 31.8661
R8016 gnd.n6164 gnd.n6163 31.8661
R8017 gnd.n6157 gnd.n1256 31.8661
R8018 gnd.n6157 gnd.n6156 31.8661
R8019 gnd.n1336 gnd.n1285 31.8661
R8020 gnd.n7305 gnd.n350 31.8661
R8021 gnd.n7412 gnd.n315 31.8661
R8022 gnd.n7314 gnd.n340 31.8661
R8023 gnd.n7320 gnd.n340 31.8661
R8024 gnd.n7393 gnd.n334 31.8661
R8025 gnd.n7397 gnd.n299 31.8661
R8026 gnd.n7421 gnd.n299 31.8661
R8027 gnd.n7429 gnd.n290 31.8661
R8028 gnd.n7429 gnd.n293 31.8661
R8029 gnd.n7437 gnd.n284 31.8661
R8030 gnd.n7445 gnd.n269 31.8661
R8031 gnd.n7453 gnd.n269 31.8661
R8032 gnd.n7461 gnd.n260 31.8661
R8033 gnd.n7461 gnd.n263 31.8661
R8034 gnd.n7469 gnd.n254 31.8661
R8035 gnd.n7477 gnd.n247 31.8661
R8036 gnd.n7493 gnd.n229 31.8661
R8037 gnd.n7493 gnd.n232 31.8661
R8038 gnd.n7501 gnd.n213 31.8661
R8039 gnd.n7577 gnd.n213 31.8661
R8040 gnd.n7577 gnd.n206 31.8661
R8041 gnd.n7585 gnd.n206 31.8661
R8042 gnd.n7665 gnd.n126 31.8661
R8043 gnd.t63 gnd.n2221 31.5474
R8044 gnd.n7393 gnd.t32 31.5474
R8045 gnd.t136 gnd.n2253 30.9101
R8046 gnd.n284 gnd.t25 30.9101
R8047 gnd.n5256 gnd.n5181 30.7517
R8048 gnd.n4752 gnd.n4637 30.7517
R8049 gnd.n3812 gnd.n962 30.2728
R8050 gnd.t75 gnd.n2285 30.2728
R8051 gnd.n254 gnd.t21 30.2728
R8052 gnd.n4996 gnd.n1901 28.9982
R8053 gnd.n5788 gnd.n1687 28.9982
R8054 gnd.n3977 gnd.t305 28.3609
R8055 gnd.t223 gnd.n126 28.3609
R8056 gnd.n2413 gnd.n962 27.0862
R8057 gnd.n1929 gnd.t149 27.0862
R8058 gnd.t155 gnd.n1659 27.0862
R8059 gnd.n4546 gnd.n4545 25.7944
R8060 gnd.n2833 gnd.n2832 25.7944
R8061 gnd.n2378 gnd.n2377 25.7944
R8062 gnd.n123 gnd.n122 25.7944
R8063 gnd.n1487 gnd.n1486 25.7944
R8064 gnd.n2037 gnd.n2036 25.7944
R8065 gnd.n1309 gnd.n1308 25.7944
R8066 gnd.n1331 gnd.n1330 25.7944
R8067 gnd.n202 gnd.n201 25.7944
R8068 gnd.n7629 gnd.n7628 25.7944
R8069 gnd.n4006 gnd.n4005 25.7944
R8070 gnd.n4038 gnd.n4037 25.7944
R8071 gnd.n3819 gnd.n3818 25.7944
R8072 gnd.n2126 gnd.n2125 25.7944
R8073 gnd.n2104 gnd.n2103 25.7944
R8074 gnd.n5891 gnd.n5890 25.7944
R8075 gnd.n3054 gnd.n2774 24.8557
R8076 gnd.n3064 gnd.n2757 24.8557
R8077 gnd.n2760 gnd.n2748 24.8557
R8078 gnd.n3085 gnd.n2749 24.8557
R8079 gnd.n3095 gnd.n2729 24.8557
R8080 gnd.n3105 gnd.n3104 24.8557
R8081 gnd.n2715 gnd.n2713 24.8557
R8082 gnd.n3136 gnd.n3135 24.8557
R8083 gnd.n3151 gnd.n2698 24.8557
R8084 gnd.n3205 gnd.n2637 24.8557
R8085 gnd.n3161 gnd.n2638 24.8557
R8086 gnd.n3198 gnd.n2649 24.8557
R8087 gnd.n2687 gnd.n2686 24.8557
R8088 gnd.n3192 gnd.n3191 24.8557
R8089 gnd.n2673 gnd.n2660 24.8557
R8090 gnd.n3231 gnd.n3230 24.8557
R8091 gnd.n3241 gnd.n2557 24.8557
R8092 gnd.n3253 gnd.n2549 24.8557
R8093 gnd.n3252 gnd.n2537 24.8557
R8094 gnd.n3271 gnd.n3270 24.8557
R8095 gnd.n3281 gnd.n2530 24.8557
R8096 gnd.n3292 gnd.n2518 24.8557
R8097 gnd.n3316 gnd.n3315 24.8557
R8098 gnd.n3327 gnd.n2501 24.8557
R8099 gnd.n3326 gnd.n2503 24.8557
R8100 gnd.n3338 gnd.n2494 24.8557
R8101 gnd.n3356 gnd.n3355 24.8557
R8102 gnd.n2485 gnd.n2474 24.8557
R8103 gnd.n3377 gnd.n2462 24.8557
R8104 gnd.n3405 gnd.n3404 24.8557
R8105 gnd.n3416 gnd.n2447 24.8557
R8106 gnd.n3427 gnd.n2440 24.8557
R8107 gnd.n3426 gnd.n2428 24.8557
R8108 gnd.n3699 gnd.n3698 24.8557
R8109 gnd.n3721 gnd.n2412 24.8557
R8110 gnd.n1974 gnd.t266 24.537
R8111 gnd.n4954 gnd.t205 24.537
R8112 gnd.n5828 gnd.t354 24.537
R8113 gnd.t233 gnd.n1245 24.537
R8114 gnd.n7485 gnd.n238 24.537
R8115 gnd.n6403 gnd.n6402 24.2183
R8116 gnd.n6396 gnd.n983 24.2183
R8117 gnd.n4382 gnd.n986 24.2183
R8118 gnd.n4413 gnd.n997 24.2183
R8119 gnd.n4390 gnd.n1007 24.2183
R8120 gnd.n6378 gnd.n1015 24.2183
R8121 gnd.n6372 gnd.n1026 24.2183
R8122 gnd.n4431 gnd.n1029 24.2183
R8123 gnd.n4462 gnd.n1039 24.2183
R8124 gnd.n4439 gnd.n1049 24.2183
R8125 gnd.n6354 gnd.n1057 24.2183
R8126 gnd.n6348 gnd.n1068 24.2183
R8127 gnd.n4513 gnd.n1071 24.2183
R8128 gnd.n4521 gnd.n1081 24.2183
R8129 gnd.n6336 gnd.n1089 24.2183
R8130 gnd.n4530 gnd.n1092 24.2183
R8131 gnd.n6330 gnd.n1100 24.2183
R8132 gnd.n4568 gnd.n2129 24.2183
R8133 gnd.n6324 gnd.n1109 24.2183
R8134 gnd.n6079 gnd.n1338 24.2183
R8135 gnd.n5914 gnd.n5905 24.2183
R8136 gnd.n5924 gnd.n1452 24.2183
R8137 gnd.n5923 gnd.n1431 24.2183
R8138 gnd.n5935 gnd.n5934 24.2183
R8139 gnd.n1435 gnd.n1422 24.2183
R8140 gnd.n5960 gnd.n1414 24.2183
R8141 gnd.n5959 gnd.n1404 24.2183
R8142 gnd.n1407 gnd.n1394 24.2183
R8143 gnd.n5982 gnd.n1396 24.2183
R8144 gnd.n6020 gnd.n1370 24.2183
R8145 gnd.n1373 gnd.n1361 24.2183
R8146 gnd.n6050 gnd.n1364 24.2183
R8147 gnd.n7235 gnd.n402 24.2183
R8148 gnd.n6004 gnd.n390 24.2183
R8149 gnd.n7226 gnd.n384 24.2183
R8150 gnd.n7281 gnd.n370 24.2183
R8151 gnd.n7253 gnd.n377 24.2183
R8152 gnd.n7290 gnd.n358 24.2183
R8153 gnd.n4897 gnd.n1973 23.8997
R8154 gnd.n6163 gnd.n1248 23.8997
R8155 gnd.n3075 gnd.t169 23.2624
R8156 gnd.n4223 gnd.t143 23.2624
R8157 gnd.n4414 gnd.t30 23.2624
R8158 gnd.n6342 gnd.t106 23.2624
R8159 gnd.n5945 gnd.t11 23.2624
R8160 gnd.n7225 gnd.t50 23.2624
R8161 gnd.n7501 gnd.t13 23.2624
R8162 gnd.n2776 gnd.t312 22.6251
R8163 gnd.n4255 gnd.t131 22.6251
R8164 gnd.n6366 gnd.t77 22.6251
R8165 gnd.n4463 gnd.t34 22.6251
R8166 gnd.n6021 gnd.t61 22.6251
R8167 gnd.n6042 gnd.t138 22.6251
R8168 gnd.n7469 gnd.t69 22.6251
R8169 gnd.n2197 gnd.t9 22.3064
R8170 gnd.t197 gnd.n312 22.3064
R8171 gnd.n4287 gnd.t97 21.9878
R8172 gnd.n6390 gnd.t83 21.9878
R8173 gnd.n7259 gnd.t46 21.9878
R8174 gnd.n7437 gnd.t183 21.9878
R8175 gnd.n4748 gnd.n4641 21.6691
R8176 gnd.n5572 gnd.n1877 21.6691
R8177 gnd.n5549 gnd.n1857 21.6691
R8178 gnd.n5542 gnd.n1849 21.6691
R8179 gnd.n5534 gnd.n1842 21.6691
R8180 gnd.n5527 gnd.n1834 21.6691
R8181 gnd.n5519 gnd.n1827 21.6691
R8182 gnd.n5512 gnd.n1820 21.6691
R8183 gnd.n5484 gnd.n1781 21.6691
R8184 gnd.n5708 gnd.n1753 21.6691
R8185 gnd.n5442 gnd.n1745 21.6691
R8186 gnd.n5434 gnd.n1739 21.6691
R8187 gnd.n5427 gnd.n1732 21.6691
R8188 gnd.n5419 gnd.n5147 21.6691
R8189 gnd.n5413 gnd.n5412 21.6691
R8190 gnd.n5384 gnd.n5179 21.6691
R8191 gnd.t3 gnd.n2781 21.3504
R8192 gnd.n4321 gnd.t19 21.3504
R8193 gnd.n4348 gnd.t36 21.3504
R8194 gnd.t86 gnd.n315 21.3504
R8195 gnd.t71 gnd.n334 21.3504
R8196 gnd.n5564 gnd.t277 21.0318
R8197 gnd.t57 gnd.n2475 20.7131
R8198 gnd.n4304 gnd.t65 20.7131
R8199 gnd.n7421 gnd.t73 20.7131
R8200 gnd.n5006 gnd.n1893 20.3945
R8201 gnd.n5580 gnd.n1869 20.3945
R8202 gnd.n5396 gnd.n1699 20.3945
R8203 gnd.n5183 gnd.n1693 20.3945
R8204 gnd.t55 gnd.n2510 20.0758
R8205 gnd.n4271 gnd.t90 20.0758
R8206 gnd.t119 gnd.n1863 20.0758
R8207 gnd.n5162 gnd.t350 20.0758
R8208 gnd.n7453 gnd.t104 20.0758
R8209 gnd.n4622 gnd.n4621 19.9763
R8210 gnd.n5232 gnd.n5231 19.9763
R8211 gnd.n4678 gnd.n4677 19.9763
R8212 gnd.n5226 gnd.n5225 19.9763
R8213 gnd.n4647 gnd.t278 19.8005
R8214 gnd.n4647 gnd.t228 19.8005
R8215 gnd.n4648 gnd.t303 19.8005
R8216 gnd.n4648 gnd.t329 19.8005
R8217 gnd.n5194 gnd.t261 19.8005
R8218 gnd.n5194 gnd.t287 19.8005
R8219 gnd.n5195 gnd.t250 19.8005
R8220 gnd.n5195 gnd.t284 19.8005
R8221 gnd.n4847 gnd.n2063 19.7572
R8222 gnd.n6156 gnd.n6155 19.7572
R8223 gnd.n4644 gnd.n4643 19.5087
R8224 gnd.n4657 gnd.n4644 19.5087
R8225 gnd.n4655 gnd.n4646 19.5087
R8226 gnd.n5199 gnd.n5193 19.5087
R8227 gnd.n3242 gnd.t214 19.4385
R8228 gnd.n4239 gnd.t162 19.4385
R8229 gnd.n4930 gnd.t153 19.4385
R8230 gnd.n5852 gnd.t216 19.4385
R8231 gnd.n7485 gnd.t48 19.4385
R8232 gnd.n4904 gnd.n1966 19.3944
R8233 gnd.n4916 gnd.n1966 19.3944
R8234 gnd.n4916 gnd.n1964 19.3944
R8235 gnd.n4920 gnd.n1964 19.3944
R8236 gnd.n4920 gnd.n1953 19.3944
R8237 gnd.n4932 gnd.n1953 19.3944
R8238 gnd.n4932 gnd.n1951 19.3944
R8239 gnd.n4936 gnd.n1951 19.3944
R8240 gnd.n4936 gnd.n1938 19.3944
R8241 gnd.n4948 gnd.n1938 19.3944
R8242 gnd.n4948 gnd.n1936 19.3944
R8243 gnd.n4952 gnd.n1936 19.3944
R8244 gnd.n4952 gnd.n1925 19.3944
R8245 gnd.n4964 gnd.n1925 19.3944
R8246 gnd.n4964 gnd.n1923 19.3944
R8247 gnd.n4968 gnd.n1923 19.3944
R8248 gnd.n4968 gnd.n1914 19.3944
R8249 gnd.n4980 gnd.n1914 19.3944
R8250 gnd.n4980 gnd.n1912 19.3944
R8251 gnd.n4984 gnd.n1912 19.3944
R8252 gnd.n4984 gnd.n1899 19.3944
R8253 gnd.n4998 gnd.n1899 19.3944
R8254 gnd.n4998 gnd.n1896 19.3944
R8255 gnd.n5003 gnd.n1896 19.3944
R8256 gnd.n5003 gnd.n1897 19.3944
R8257 gnd.n1897 gnd.n1867 19.3944
R8258 gnd.n5582 gnd.n1867 19.3944
R8259 gnd.n5582 gnd.n1865 19.3944
R8260 gnd.n5586 gnd.n1865 19.3944
R8261 gnd.n5586 gnd.n1853 19.3944
R8262 gnd.n5598 gnd.n1853 19.3944
R8263 gnd.n5598 gnd.n1851 19.3944
R8264 gnd.n5602 gnd.n1851 19.3944
R8265 gnd.n5602 gnd.n1838 19.3944
R8266 gnd.n5614 gnd.n1838 19.3944
R8267 gnd.n5614 gnd.n1836 19.3944
R8268 gnd.n5618 gnd.n1836 19.3944
R8269 gnd.n5618 gnd.n1824 19.3944
R8270 gnd.n5630 gnd.n1824 19.3944
R8271 gnd.n5630 gnd.n1822 19.3944
R8272 gnd.n5634 gnd.n1822 19.3944
R8273 gnd.n5634 gnd.n1809 19.3944
R8274 gnd.n5646 gnd.n1809 19.3944
R8275 gnd.n5646 gnd.n1807 19.3944
R8276 gnd.n5650 gnd.n1807 19.3944
R8277 gnd.n5650 gnd.n1794 19.3944
R8278 gnd.n5662 gnd.n1794 19.3944
R8279 gnd.n5662 gnd.n1792 19.3944
R8280 gnd.n5666 gnd.n1792 19.3944
R8281 gnd.n5666 gnd.n1779 19.3944
R8282 gnd.n5678 gnd.n1779 19.3944
R8283 gnd.n5678 gnd.n1777 19.3944
R8284 gnd.n5682 gnd.n1777 19.3944
R8285 gnd.n5682 gnd.n1764 19.3944
R8286 gnd.n5694 gnd.n1764 19.3944
R8287 gnd.n5694 gnd.n1762 19.3944
R8288 gnd.n5698 gnd.n1762 19.3944
R8289 gnd.n5698 gnd.n1749 19.3944
R8290 gnd.n5710 gnd.n1749 19.3944
R8291 gnd.n5710 gnd.n1747 19.3944
R8292 gnd.n5714 gnd.n1747 19.3944
R8293 gnd.n5714 gnd.n1736 19.3944
R8294 gnd.n5726 gnd.n1736 19.3944
R8295 gnd.n5726 gnd.n1734 19.3944
R8296 gnd.n5730 gnd.n1734 19.3944
R8297 gnd.n5730 gnd.n1724 19.3944
R8298 gnd.n5742 gnd.n1724 19.3944
R8299 gnd.n5742 gnd.n1722 19.3944
R8300 gnd.n5746 gnd.n1722 19.3944
R8301 gnd.n5746 gnd.n1711 19.3944
R8302 gnd.n5758 gnd.n1711 19.3944
R8303 gnd.n5758 gnd.n1709 19.3944
R8304 gnd.n5762 gnd.n1709 19.3944
R8305 gnd.n5762 gnd.n1697 19.3944
R8306 gnd.n5774 gnd.n1697 19.3944
R8307 gnd.n5774 gnd.n1695 19.3944
R8308 gnd.n5778 gnd.n1695 19.3944
R8309 gnd.n5778 gnd.n1682 19.3944
R8310 gnd.n5790 gnd.n1682 19.3944
R8311 gnd.n5790 gnd.n1680 19.3944
R8312 gnd.n5794 gnd.n1680 19.3944
R8313 gnd.n5794 gnd.n1670 19.3944
R8314 gnd.n5806 gnd.n1670 19.3944
R8315 gnd.n5806 gnd.n1668 19.3944
R8316 gnd.n5810 gnd.n1668 19.3944
R8317 gnd.n5810 gnd.n1657 19.3944
R8318 gnd.n5822 gnd.n1657 19.3944
R8319 gnd.n5822 gnd.n1655 19.3944
R8320 gnd.n5826 gnd.n1655 19.3944
R8321 gnd.n5826 gnd.n1644 19.3944
R8322 gnd.n5838 gnd.n1644 19.3944
R8323 gnd.n5838 gnd.n1642 19.3944
R8324 gnd.n5842 gnd.n1642 19.3944
R8325 gnd.n5842 gnd.n1631 19.3944
R8326 gnd.n5854 gnd.n1631 19.3944
R8327 gnd.n5854 gnd.n1628 19.3944
R8328 gnd.n5860 gnd.n1628 19.3944
R8329 gnd.n5860 gnd.n1629 19.3944
R8330 gnd.n1629 gnd.n1616 19.3944
R8331 gnd.n5876 gnd.n1616 19.3944
R8332 gnd.n5877 gnd.n5876 19.3944
R8333 gnd.n4550 gnd.n1977 19.3944
R8334 gnd.n4900 gnd.n1977 19.3944
R8335 gnd.n4901 gnd.n4900 19.3944
R8336 gnd.n4894 gnd.n4893 19.3944
R8337 gnd.n4893 gnd.n1995 19.3944
R8338 gnd.n4886 gnd.n1995 19.3944
R8339 gnd.n4886 gnd.n4885 19.3944
R8340 gnd.n4885 gnd.n2006 19.3944
R8341 gnd.n4878 gnd.n2006 19.3944
R8342 gnd.n4878 gnd.n4877 19.3944
R8343 gnd.n4877 gnd.n2014 19.3944
R8344 gnd.n4870 gnd.n2014 19.3944
R8345 gnd.n4870 gnd.n4869 19.3944
R8346 gnd.n4869 gnd.n2024 19.3944
R8347 gnd.n4862 gnd.n2024 19.3944
R8348 gnd.n4862 gnd.n4861 19.3944
R8349 gnd.n4861 gnd.n2032 19.3944
R8350 gnd.n4854 gnd.n2032 19.3944
R8351 gnd.n4854 gnd.n4853 19.3944
R8352 gnd.n4853 gnd.n2044 19.3944
R8353 gnd.n4561 gnd.n2044 19.3944
R8354 gnd.n4561 gnd.n4560 19.3944
R8355 gnd.n4560 gnd.n4559 19.3944
R8356 gnd.n4559 gnd.n4540 19.3944
R8357 gnd.n4555 gnd.n4540 19.3944
R8358 gnd.n4555 gnd.n4554 19.3944
R8359 gnd.n4554 gnd.n4553 19.3944
R8360 gnd.n2957 gnd.n2956 19.3944
R8361 gnd.n2956 gnd.n2955 19.3944
R8362 gnd.n2955 gnd.n2954 19.3944
R8363 gnd.n2954 gnd.n2952 19.3944
R8364 gnd.n2952 gnd.n2949 19.3944
R8365 gnd.n2949 gnd.n2948 19.3944
R8366 gnd.n2948 gnd.n2945 19.3944
R8367 gnd.n2945 gnd.n2944 19.3944
R8368 gnd.n2944 gnd.n2941 19.3944
R8369 gnd.n2941 gnd.n2940 19.3944
R8370 gnd.n2940 gnd.n2937 19.3944
R8371 gnd.n2937 gnd.n2936 19.3944
R8372 gnd.n2936 gnd.n2933 19.3944
R8373 gnd.n2933 gnd.n2932 19.3944
R8374 gnd.n2932 gnd.n2929 19.3944
R8375 gnd.n2929 gnd.n2928 19.3944
R8376 gnd.n2928 gnd.n2925 19.3944
R8377 gnd.n2925 gnd.n2924 19.3944
R8378 gnd.n2924 gnd.n2921 19.3944
R8379 gnd.n2921 gnd.n2920 19.3944
R8380 gnd.n2920 gnd.n2917 19.3944
R8381 gnd.n2917 gnd.n2916 19.3944
R8382 gnd.n2913 gnd.n2912 19.3944
R8383 gnd.n2912 gnd.n2868 19.3944
R8384 gnd.n2963 gnd.n2868 19.3944
R8385 gnd.n3729 gnd.n3728 19.3944
R8386 gnd.n3728 gnd.n3725 19.3944
R8387 gnd.n3725 gnd.n3724 19.3944
R8388 gnd.n3774 gnd.n3773 19.3944
R8389 gnd.n3773 gnd.n3772 19.3944
R8390 gnd.n3772 gnd.n3769 19.3944
R8391 gnd.n3769 gnd.n3768 19.3944
R8392 gnd.n3768 gnd.n3765 19.3944
R8393 gnd.n3765 gnd.n3764 19.3944
R8394 gnd.n3764 gnd.n3761 19.3944
R8395 gnd.n3761 gnd.n3760 19.3944
R8396 gnd.n3760 gnd.n3757 19.3944
R8397 gnd.n3757 gnd.n3756 19.3944
R8398 gnd.n3756 gnd.n3753 19.3944
R8399 gnd.n3753 gnd.n3752 19.3944
R8400 gnd.n3752 gnd.n3749 19.3944
R8401 gnd.n3749 gnd.n3748 19.3944
R8402 gnd.n3748 gnd.n3745 19.3944
R8403 gnd.n3745 gnd.n3744 19.3944
R8404 gnd.n3744 gnd.n3741 19.3944
R8405 gnd.n3741 gnd.n3740 19.3944
R8406 gnd.n3740 gnd.n3737 19.3944
R8407 gnd.n3737 gnd.n3736 19.3944
R8408 gnd.n3736 gnd.n3733 19.3944
R8409 gnd.n3733 gnd.n3732 19.3944
R8410 gnd.n3056 gnd.n2765 19.3944
R8411 gnd.n3066 gnd.n2765 19.3944
R8412 gnd.n3067 gnd.n3066 19.3944
R8413 gnd.n3067 gnd.n2746 19.3944
R8414 gnd.n3087 gnd.n2746 19.3944
R8415 gnd.n3087 gnd.n2738 19.3944
R8416 gnd.n3097 gnd.n2738 19.3944
R8417 gnd.n3098 gnd.n3097 19.3944
R8418 gnd.n3099 gnd.n3098 19.3944
R8419 gnd.n3099 gnd.n2721 19.3944
R8420 gnd.n3116 gnd.n2721 19.3944
R8421 gnd.n3119 gnd.n3116 19.3944
R8422 gnd.n3119 gnd.n3118 19.3944
R8423 gnd.n3118 gnd.n2694 19.3944
R8424 gnd.n3158 gnd.n2694 19.3944
R8425 gnd.n3158 gnd.n2691 19.3944
R8426 gnd.n3164 gnd.n2691 19.3944
R8427 gnd.n3165 gnd.n3164 19.3944
R8428 gnd.n3165 gnd.n2689 19.3944
R8429 gnd.n3171 gnd.n2689 19.3944
R8430 gnd.n3174 gnd.n3171 19.3944
R8431 gnd.n3176 gnd.n3174 19.3944
R8432 gnd.n3182 gnd.n3176 19.3944
R8433 gnd.n3182 gnd.n3181 19.3944
R8434 gnd.n3181 gnd.n2552 19.3944
R8435 gnd.n3248 gnd.n2552 19.3944
R8436 gnd.n3249 gnd.n3248 19.3944
R8437 gnd.n3249 gnd.n2545 19.3944
R8438 gnd.n3260 gnd.n2545 19.3944
R8439 gnd.n3261 gnd.n3260 19.3944
R8440 gnd.n3261 gnd.n2528 19.3944
R8441 gnd.n2528 gnd.n2526 19.3944
R8442 gnd.n3285 gnd.n2526 19.3944
R8443 gnd.n3286 gnd.n3285 19.3944
R8444 gnd.n3286 gnd.n2497 19.3944
R8445 gnd.n3333 gnd.n2497 19.3944
R8446 gnd.n3334 gnd.n3333 19.3944
R8447 gnd.n3334 gnd.n2490 19.3944
R8448 gnd.n3345 gnd.n2490 19.3944
R8449 gnd.n3346 gnd.n3345 19.3944
R8450 gnd.n3346 gnd.n2473 19.3944
R8451 gnd.n2473 gnd.n2471 19.3944
R8452 gnd.n3370 gnd.n2471 19.3944
R8453 gnd.n3371 gnd.n3370 19.3944
R8454 gnd.n3371 gnd.n2443 19.3944
R8455 gnd.n3422 gnd.n2443 19.3944
R8456 gnd.n3423 gnd.n3422 19.3944
R8457 gnd.n3423 gnd.n2436 19.3944
R8458 gnd.n3690 gnd.n2436 19.3944
R8459 gnd.n3691 gnd.n3690 19.3944
R8460 gnd.n3691 gnd.n2417 19.3944
R8461 gnd.n3716 gnd.n2417 19.3944
R8462 gnd.n3716 gnd.n2418 19.3944
R8463 gnd.n3047 gnd.n3046 19.3944
R8464 gnd.n3046 gnd.n2779 19.3944
R8465 gnd.n2802 gnd.n2779 19.3944
R8466 gnd.n2805 gnd.n2802 19.3944
R8467 gnd.n2805 gnd.n2798 19.3944
R8468 gnd.n2809 gnd.n2798 19.3944
R8469 gnd.n2812 gnd.n2809 19.3944
R8470 gnd.n2815 gnd.n2812 19.3944
R8471 gnd.n2815 gnd.n2796 19.3944
R8472 gnd.n2819 gnd.n2796 19.3944
R8473 gnd.n2822 gnd.n2819 19.3944
R8474 gnd.n2825 gnd.n2822 19.3944
R8475 gnd.n2825 gnd.n2794 19.3944
R8476 gnd.n2829 gnd.n2794 19.3944
R8477 gnd.n3052 gnd.n3051 19.3944
R8478 gnd.n3051 gnd.n2755 19.3944
R8479 gnd.n3077 gnd.n2755 19.3944
R8480 gnd.n3077 gnd.n2753 19.3944
R8481 gnd.n3083 gnd.n2753 19.3944
R8482 gnd.n3083 gnd.n3082 19.3944
R8483 gnd.n3082 gnd.n2727 19.3944
R8484 gnd.n3107 gnd.n2727 19.3944
R8485 gnd.n3107 gnd.n2725 19.3944
R8486 gnd.n3111 gnd.n2725 19.3944
R8487 gnd.n3111 gnd.n2705 19.3944
R8488 gnd.n3138 gnd.n2705 19.3944
R8489 gnd.n3138 gnd.n2703 19.3944
R8490 gnd.n3148 gnd.n2703 19.3944
R8491 gnd.n3148 gnd.n3147 19.3944
R8492 gnd.n3147 gnd.n3146 19.3944
R8493 gnd.n3146 gnd.n2652 19.3944
R8494 gnd.n3196 gnd.n2652 19.3944
R8495 gnd.n3196 gnd.n3195 19.3944
R8496 gnd.n3195 gnd.n3194 19.3944
R8497 gnd.n3194 gnd.n2656 19.3944
R8498 gnd.n2676 gnd.n2656 19.3944
R8499 gnd.n2676 gnd.n2562 19.3944
R8500 gnd.n3233 gnd.n2562 19.3944
R8501 gnd.n3233 gnd.n2560 19.3944
R8502 gnd.n3239 gnd.n2560 19.3944
R8503 gnd.n3239 gnd.n3238 19.3944
R8504 gnd.n3238 gnd.n2535 19.3944
R8505 gnd.n3273 gnd.n2535 19.3944
R8506 gnd.n3273 gnd.n2533 19.3944
R8507 gnd.n3279 gnd.n2533 19.3944
R8508 gnd.n3279 gnd.n3278 19.3944
R8509 gnd.n3278 gnd.n2508 19.3944
R8510 gnd.n3318 gnd.n2508 19.3944
R8511 gnd.n3318 gnd.n2506 19.3944
R8512 gnd.n3324 gnd.n2506 19.3944
R8513 gnd.n3324 gnd.n3323 19.3944
R8514 gnd.n3323 gnd.n2480 19.3944
R8515 gnd.n3358 gnd.n2480 19.3944
R8516 gnd.n3358 gnd.n2478 19.3944
R8517 gnd.n3364 gnd.n2478 19.3944
R8518 gnd.n3364 gnd.n3363 19.3944
R8519 gnd.n3363 gnd.n2453 19.3944
R8520 gnd.n3407 gnd.n2453 19.3944
R8521 gnd.n3407 gnd.n2451 19.3944
R8522 gnd.n3413 gnd.n2451 19.3944
R8523 gnd.n3413 gnd.n3412 19.3944
R8524 gnd.n3412 gnd.n2426 19.3944
R8525 gnd.n3701 gnd.n2426 19.3944
R8526 gnd.n3701 gnd.n2424 19.3944
R8527 gnd.n3709 gnd.n2424 19.3944
R8528 gnd.n3709 gnd.n3708 19.3944
R8529 gnd.n3708 gnd.n3707 19.3944
R8530 gnd.n3810 gnd.n3809 19.3944
R8531 gnd.n3809 gnd.n2364 19.3944
R8532 gnd.n3805 gnd.n2364 19.3944
R8533 gnd.n3805 gnd.n3802 19.3944
R8534 gnd.n3802 gnd.n3799 19.3944
R8535 gnd.n3799 gnd.n3798 19.3944
R8536 gnd.n3798 gnd.n3795 19.3944
R8537 gnd.n3795 gnd.n3794 19.3944
R8538 gnd.n3794 gnd.n3791 19.3944
R8539 gnd.n3791 gnd.n3790 19.3944
R8540 gnd.n3790 gnd.n3787 19.3944
R8541 gnd.n3787 gnd.n3786 19.3944
R8542 gnd.n3786 gnd.n3783 19.3944
R8543 gnd.n3783 gnd.n3782 19.3944
R8544 gnd.n2967 gnd.n2866 19.3944
R8545 gnd.n2967 gnd.n2857 19.3944
R8546 gnd.n2980 gnd.n2857 19.3944
R8547 gnd.n2980 gnd.n2855 19.3944
R8548 gnd.n2984 gnd.n2855 19.3944
R8549 gnd.n2984 gnd.n2845 19.3944
R8550 gnd.n2996 gnd.n2845 19.3944
R8551 gnd.n2996 gnd.n2843 19.3944
R8552 gnd.n3030 gnd.n2843 19.3944
R8553 gnd.n3030 gnd.n3029 19.3944
R8554 gnd.n3029 gnd.n3028 19.3944
R8555 gnd.n3028 gnd.n3027 19.3944
R8556 gnd.n3027 gnd.n3024 19.3944
R8557 gnd.n3024 gnd.n3023 19.3944
R8558 gnd.n3023 gnd.n3022 19.3944
R8559 gnd.n3022 gnd.n3020 19.3944
R8560 gnd.n3020 gnd.n3019 19.3944
R8561 gnd.n3019 gnd.n3016 19.3944
R8562 gnd.n3016 gnd.n3015 19.3944
R8563 gnd.n3015 gnd.n3014 19.3944
R8564 gnd.n3014 gnd.n3012 19.3944
R8565 gnd.n3012 gnd.n2711 19.3944
R8566 gnd.n3127 gnd.n2711 19.3944
R8567 gnd.n3127 gnd.n2709 19.3944
R8568 gnd.n3133 gnd.n2709 19.3944
R8569 gnd.n3133 gnd.n3132 19.3944
R8570 gnd.n3132 gnd.n2633 19.3944
R8571 gnd.n3207 gnd.n2633 19.3944
R8572 gnd.n3207 gnd.n2634 19.3944
R8573 gnd.n2681 gnd.n2680 19.3944
R8574 gnd.n2684 gnd.n2683 19.3944
R8575 gnd.n2671 gnd.n2670 19.3944
R8576 gnd.n3226 gnd.n2567 19.3944
R8577 gnd.n3226 gnd.n3225 19.3944
R8578 gnd.n3225 gnd.n3224 19.3944
R8579 gnd.n3224 gnd.n3222 19.3944
R8580 gnd.n3222 gnd.n3221 19.3944
R8581 gnd.n3221 gnd.n3219 19.3944
R8582 gnd.n3219 gnd.n3218 19.3944
R8583 gnd.n3218 gnd.n2516 19.3944
R8584 gnd.n3294 gnd.n2516 19.3944
R8585 gnd.n3294 gnd.n2514 19.3944
R8586 gnd.n3313 gnd.n2514 19.3944
R8587 gnd.n3313 gnd.n3312 19.3944
R8588 gnd.n3312 gnd.n3311 19.3944
R8589 gnd.n3311 gnd.n3309 19.3944
R8590 gnd.n3309 gnd.n3308 19.3944
R8591 gnd.n3308 gnd.n3306 19.3944
R8592 gnd.n3306 gnd.n3305 19.3944
R8593 gnd.n3305 gnd.n2460 19.3944
R8594 gnd.n3379 gnd.n2460 19.3944
R8595 gnd.n3379 gnd.n2458 19.3944
R8596 gnd.n3402 gnd.n2458 19.3944
R8597 gnd.n3402 gnd.n3401 19.3944
R8598 gnd.n3401 gnd.n3400 19.3944
R8599 gnd.n3400 gnd.n3397 19.3944
R8600 gnd.n3397 gnd.n3396 19.3944
R8601 gnd.n3396 gnd.n3394 19.3944
R8602 gnd.n3394 gnd.n3393 19.3944
R8603 gnd.n3393 gnd.n3391 19.3944
R8604 gnd.n3391 gnd.n2411 19.3944
R8605 gnd.n2972 gnd.n2862 19.3944
R8606 gnd.n2972 gnd.n2860 19.3944
R8607 gnd.n2976 gnd.n2860 19.3944
R8608 gnd.n2976 gnd.n2851 19.3944
R8609 gnd.n2988 gnd.n2851 19.3944
R8610 gnd.n2988 gnd.n2849 19.3944
R8611 gnd.n2992 gnd.n2849 19.3944
R8612 gnd.n2992 gnd.n2838 19.3944
R8613 gnd.n3034 gnd.n2838 19.3944
R8614 gnd.n3034 gnd.n2792 19.3944
R8615 gnd.n3040 gnd.n2792 19.3944
R8616 gnd.n3040 gnd.n3039 19.3944
R8617 gnd.n3039 gnd.n2770 19.3944
R8618 gnd.n3061 gnd.n2770 19.3944
R8619 gnd.n3061 gnd.n2763 19.3944
R8620 gnd.n3072 gnd.n2763 19.3944
R8621 gnd.n3072 gnd.n3071 19.3944
R8622 gnd.n3071 gnd.n2744 19.3944
R8623 gnd.n3092 gnd.n2744 19.3944
R8624 gnd.n3092 gnd.n2734 19.3944
R8625 gnd.n3102 gnd.n2734 19.3944
R8626 gnd.n3102 gnd.n2717 19.3944
R8627 gnd.n3123 gnd.n2717 19.3944
R8628 gnd.n3123 gnd.n3122 19.3944
R8629 gnd.n3122 gnd.n2696 19.3944
R8630 gnd.n3153 gnd.n2696 19.3944
R8631 gnd.n3153 gnd.n2641 19.3944
R8632 gnd.n3203 gnd.n2641 19.3944
R8633 gnd.n3203 gnd.n3202 19.3944
R8634 gnd.n3202 gnd.n3201 19.3944
R8635 gnd.n3201 gnd.n2645 19.3944
R8636 gnd.n2663 gnd.n2645 19.3944
R8637 gnd.n3189 gnd.n2663 19.3944
R8638 gnd.n3189 gnd.n3188 19.3944
R8639 gnd.n3188 gnd.n3187 19.3944
R8640 gnd.n3187 gnd.n2667 19.3944
R8641 gnd.n2667 gnd.n2554 19.3944
R8642 gnd.n3244 gnd.n2554 19.3944
R8643 gnd.n3244 gnd.n2547 19.3944
R8644 gnd.n3255 gnd.n2547 19.3944
R8645 gnd.n3255 gnd.n2543 19.3944
R8646 gnd.n3268 gnd.n2543 19.3944
R8647 gnd.n3268 gnd.n3267 19.3944
R8648 gnd.n3267 gnd.n2522 19.3944
R8649 gnd.n3290 gnd.n2522 19.3944
R8650 gnd.n3290 gnd.n3289 19.3944
R8651 gnd.n3289 gnd.n2499 19.3944
R8652 gnd.n3329 gnd.n2499 19.3944
R8653 gnd.n3329 gnd.n2492 19.3944
R8654 gnd.n3340 gnd.n2492 19.3944
R8655 gnd.n3340 gnd.n2488 19.3944
R8656 gnd.n3353 gnd.n2488 19.3944
R8657 gnd.n3353 gnd.n3352 19.3944
R8658 gnd.n3352 gnd.n2467 19.3944
R8659 gnd.n3375 gnd.n2467 19.3944
R8660 gnd.n3375 gnd.n3374 19.3944
R8661 gnd.n3374 gnd.n2445 19.3944
R8662 gnd.n3418 gnd.n2445 19.3944
R8663 gnd.n3418 gnd.n2438 19.3944
R8664 gnd.n3429 gnd.n2438 19.3944
R8665 gnd.n3429 gnd.n2434 19.3944
R8666 gnd.n3696 gnd.n2434 19.3944
R8667 gnd.n3696 gnd.n3695 19.3944
R8668 gnd.n3695 gnd.n2415 19.3944
R8669 gnd.n3719 gnd.n2415 19.3944
R8670 gnd.n5916 gnd.n5904 19.3944
R8671 gnd.n5916 gnd.n1476 19.3944
R8672 gnd.n5921 gnd.n1476 19.3944
R8673 gnd.n5921 gnd.n1477 19.3944
R8674 gnd.n1477 gnd.n1420 19.3944
R8675 gnd.n5947 gnd.n1420 19.3944
R8676 gnd.n5947 gnd.n1417 19.3944
R8677 gnd.n5957 gnd.n1417 19.3944
R8678 gnd.n5957 gnd.n1418 19.3944
R8679 gnd.n5953 gnd.n1418 19.3944
R8680 gnd.n5953 gnd.n5952 19.3944
R8681 gnd.n5952 gnd.n1382 19.3944
R8682 gnd.n6017 gnd.n1382 19.3944
R8683 gnd.n6017 gnd.n1383 19.3944
R8684 gnd.n6013 gnd.n1383 19.3944
R8685 gnd.n6013 gnd.n6012 19.3944
R8686 gnd.n6012 gnd.n6011 19.3944
R8687 gnd.n6011 gnd.n6001 19.3944
R8688 gnd.n6007 gnd.n6001 19.3944
R8689 gnd.n6007 gnd.n6006 19.3944
R8690 gnd.n6006 gnd.n382 19.3944
R8691 gnd.n7261 gnd.n382 19.3944
R8692 gnd.n7262 gnd.n7261 19.3944
R8693 gnd.n7262 gnd.n379 19.3944
R8694 gnd.n7267 gnd.n379 19.3944
R8695 gnd.n7267 gnd.n380 19.3944
R8696 gnd.n380 gnd.n348 19.3944
R8697 gnd.n7307 gnd.n348 19.3944
R8698 gnd.n7307 gnd.n346 19.3944
R8699 gnd.n7311 gnd.n346 19.3944
R8700 gnd.n7312 gnd.n7311 19.3944
R8701 gnd.n7312 gnd.n80 19.3944
R8702 gnd.n7716 gnd.n80 19.3944
R8703 gnd.n7716 gnd.n7715 19.3944
R8704 gnd.n7715 gnd.n7714 19.3944
R8705 gnd.n7714 gnd.n85 19.3944
R8706 gnd.n7710 gnd.n85 19.3944
R8707 gnd.n7710 gnd.n7709 19.3944
R8708 gnd.n7709 gnd.n7708 19.3944
R8709 gnd.n7708 gnd.n90 19.3944
R8710 gnd.n7704 gnd.n90 19.3944
R8711 gnd.n7704 gnd.n7703 19.3944
R8712 gnd.n7703 gnd.n7702 19.3944
R8713 gnd.n7702 gnd.n95 19.3944
R8714 gnd.n7698 gnd.n95 19.3944
R8715 gnd.n7698 gnd.n7697 19.3944
R8716 gnd.n7697 gnd.n7696 19.3944
R8717 gnd.n7696 gnd.n100 19.3944
R8718 gnd.n7692 gnd.n100 19.3944
R8719 gnd.n7692 gnd.n7691 19.3944
R8720 gnd.n7691 gnd.n7690 19.3944
R8721 gnd.n7690 gnd.n105 19.3944
R8722 gnd.n7686 gnd.n105 19.3944
R8723 gnd.n7686 gnd.n7685 19.3944
R8724 gnd.n7685 gnd.n7684 19.3944
R8725 gnd.n7684 gnd.n110 19.3944
R8726 gnd.n7680 gnd.n110 19.3944
R8727 gnd.n7680 gnd.n7679 19.3944
R8728 gnd.n7679 gnd.n7678 19.3944
R8729 gnd.n7678 gnd.n115 19.3944
R8730 gnd.n7674 gnd.n115 19.3944
R8731 gnd.n7674 gnd.n7673 19.3944
R8732 gnd.n7673 gnd.n7672 19.3944
R8733 gnd.n7672 gnd.n120 19.3944
R8734 gnd.n7566 gnd.n7565 19.3944
R8735 gnd.n7565 gnd.n7564 19.3944
R8736 gnd.n7564 gnd.n7513 19.3944
R8737 gnd.n7560 gnd.n7513 19.3944
R8738 gnd.n7560 gnd.n7559 19.3944
R8739 gnd.n7559 gnd.n7558 19.3944
R8740 gnd.n7558 gnd.n7521 19.3944
R8741 gnd.n7554 gnd.n7521 19.3944
R8742 gnd.n7554 gnd.n7553 19.3944
R8743 gnd.n7553 gnd.n7552 19.3944
R8744 gnd.n7552 gnd.n7529 19.3944
R8745 gnd.n7548 gnd.n7529 19.3944
R8746 gnd.n7548 gnd.n7547 19.3944
R8747 gnd.n7547 gnd.n7546 19.3944
R8748 gnd.n7546 gnd.n7537 19.3944
R8749 gnd.n7542 gnd.n7537 19.3944
R8750 gnd.n1521 gnd.n1517 19.3944
R8751 gnd.n1524 gnd.n1521 19.3944
R8752 gnd.n1527 gnd.n1524 19.3944
R8753 gnd.n1527 gnd.n1510 19.3944
R8754 gnd.n1540 gnd.n1510 19.3944
R8755 gnd.n1543 gnd.n1540 19.3944
R8756 gnd.n1546 gnd.n1543 19.3944
R8757 gnd.n1546 gnd.n1503 19.3944
R8758 gnd.n1559 gnd.n1503 19.3944
R8759 gnd.n1562 gnd.n1559 19.3944
R8760 gnd.n1565 gnd.n1562 19.3944
R8761 gnd.n1565 gnd.n1496 19.3944
R8762 gnd.n1577 gnd.n1496 19.3944
R8763 gnd.n1580 gnd.n1577 19.3944
R8764 gnd.n1580 gnd.n1488 19.3944
R8765 gnd.n1593 gnd.n1488 19.3944
R8766 gnd.n6077 gnd.n1341 19.3944
R8767 gnd.n6073 gnd.n1341 19.3944
R8768 gnd.n6073 gnd.n6072 19.3944
R8769 gnd.n6072 gnd.n6071 19.3944
R8770 gnd.n6071 gnd.n1347 19.3944
R8771 gnd.n6067 gnd.n1347 19.3944
R8772 gnd.n6067 gnd.n6066 19.3944
R8773 gnd.n6066 gnd.n6065 19.3944
R8774 gnd.n6065 gnd.n1352 19.3944
R8775 gnd.n6061 gnd.n1352 19.3944
R8776 gnd.n6061 gnd.n6060 19.3944
R8777 gnd.n6060 gnd.n6059 19.3944
R8778 gnd.n6059 gnd.n1357 19.3944
R8779 gnd.n6055 gnd.n1357 19.3944
R8780 gnd.n6055 gnd.n6054 19.3944
R8781 gnd.n6054 gnd.n6053 19.3944
R8782 gnd.n6053 gnd.n405 19.3944
R8783 gnd.n7233 gnd.n405 19.3944
R8784 gnd.n7233 gnd.n406 19.3944
R8785 gnd.n7229 gnd.n406 19.3944
R8786 gnd.n7229 gnd.n7228 19.3944
R8787 gnd.n7228 gnd.n373 19.3944
R8788 gnd.n7279 gnd.n373 19.3944
R8789 gnd.n7279 gnd.n374 19.3944
R8790 gnd.n7275 gnd.n374 19.3944
R8791 gnd.n7275 gnd.n7274 19.3944
R8792 gnd.n7274 gnd.n7273 19.3944
R8793 gnd.n7273 gnd.n318 19.3944
R8794 gnd.n7410 gnd.n318 19.3944
R8795 gnd.n7410 gnd.n319 19.3944
R8796 gnd.n7406 gnd.n319 19.3944
R8797 gnd.n7406 gnd.n7405 19.3944
R8798 gnd.n7405 gnd.n7404 19.3944
R8799 gnd.n7404 gnd.n325 19.3944
R8800 gnd.n7400 gnd.n325 19.3944
R8801 gnd.n7400 gnd.n7399 19.3944
R8802 gnd.n7399 gnd.n297 19.3944
R8803 gnd.n7423 gnd.n297 19.3944
R8804 gnd.n7423 gnd.n295 19.3944
R8805 gnd.n7427 gnd.n295 19.3944
R8806 gnd.n7427 gnd.n281 19.3944
R8807 gnd.n7439 gnd.n281 19.3944
R8808 gnd.n7439 gnd.n279 19.3944
R8809 gnd.n7443 gnd.n279 19.3944
R8810 gnd.n7443 gnd.n267 19.3944
R8811 gnd.n7455 gnd.n267 19.3944
R8812 gnd.n7455 gnd.n265 19.3944
R8813 gnd.n7459 gnd.n265 19.3944
R8814 gnd.n7459 gnd.n251 19.3944
R8815 gnd.n7471 gnd.n251 19.3944
R8816 gnd.n7471 gnd.n249 19.3944
R8817 gnd.n7475 gnd.n249 19.3944
R8818 gnd.n7475 gnd.n236 19.3944
R8819 gnd.n7487 gnd.n236 19.3944
R8820 gnd.n7487 gnd.n234 19.3944
R8821 gnd.n7491 gnd.n234 19.3944
R8822 gnd.n7491 gnd.n221 19.3944
R8823 gnd.n7503 gnd.n221 19.3944
R8824 gnd.n7503 gnd.n218 19.3944
R8825 gnd.n7575 gnd.n218 19.3944
R8826 gnd.n7575 gnd.n219 19.3944
R8827 gnd.n7571 gnd.n219 19.3944
R8828 gnd.n7571 gnd.n7570 19.3944
R8829 gnd.n7570 gnd.n7569 19.3944
R8830 gnd.n2048 gnd.n1115 19.3944
R8831 gnd.n2048 gnd.n1998 19.3944
R8832 gnd.n4890 gnd.n1998 19.3944
R8833 gnd.n4890 gnd.n4889 19.3944
R8834 gnd.n4889 gnd.n2001 19.3944
R8835 gnd.n4882 gnd.n2001 19.3944
R8836 gnd.n4882 gnd.n4881 19.3944
R8837 gnd.n4881 gnd.n2010 19.3944
R8838 gnd.n4874 gnd.n2010 19.3944
R8839 gnd.n4874 gnd.n4873 19.3944
R8840 gnd.n4873 gnd.n2018 19.3944
R8841 gnd.n4866 gnd.n2018 19.3944
R8842 gnd.n4866 gnd.n4865 19.3944
R8843 gnd.n4865 gnd.n2028 19.3944
R8844 gnd.n4858 gnd.n2028 19.3944
R8845 gnd.n4858 gnd.n4857 19.3944
R8846 gnd.n6405 gnd.n968 19.3944
R8847 gnd.n4375 gnd.n968 19.3944
R8848 gnd.n4375 gnd.n4373 19.3944
R8849 gnd.n4379 gnd.n4373 19.3944
R8850 gnd.n4379 gnd.n2170 19.3944
R8851 gnd.n4416 gnd.n2170 19.3944
R8852 gnd.n4416 gnd.n2168 19.3944
R8853 gnd.n4420 gnd.n2168 19.3944
R8854 gnd.n4420 gnd.n2166 19.3944
R8855 gnd.n4424 gnd.n2166 19.3944
R8856 gnd.n4424 gnd.n2164 19.3944
R8857 gnd.n4428 gnd.n2164 19.3944
R8858 gnd.n4428 gnd.n2149 19.3944
R8859 gnd.n4465 gnd.n2149 19.3944
R8860 gnd.n4465 gnd.n2147 19.3944
R8861 gnd.n4469 gnd.n2147 19.3944
R8862 gnd.n4469 gnd.n2145 19.3944
R8863 gnd.n4473 gnd.n2145 19.3944
R8864 gnd.n4473 gnd.n2143 19.3944
R8865 gnd.n4510 gnd.n2143 19.3944
R8866 gnd.n4510 gnd.n4509 19.3944
R8867 gnd.n4509 gnd.n4508 19.3944
R8868 gnd.n4508 gnd.n4479 19.3944
R8869 gnd.n4504 gnd.n4479 19.3944
R8870 gnd.n4504 gnd.n4503 19.3944
R8871 gnd.n4503 gnd.n4502 19.3944
R8872 gnd.n4502 gnd.n4485 19.3944
R8873 gnd.n4498 gnd.n4485 19.3944
R8874 gnd.n4498 gnd.n4497 19.3944
R8875 gnd.n4497 gnd.n4496 19.3944
R8876 gnd.n4496 gnd.n4492 19.3944
R8877 gnd.n4492 gnd.n1971 19.3944
R8878 gnd.n4908 gnd.n1971 19.3944
R8879 gnd.n4908 gnd.n1969 19.3944
R8880 gnd.n4912 gnd.n1969 19.3944
R8881 gnd.n4912 gnd.n1959 19.3944
R8882 gnd.n4924 gnd.n1959 19.3944
R8883 gnd.n4924 gnd.n1957 19.3944
R8884 gnd.n4928 gnd.n1957 19.3944
R8885 gnd.n4928 gnd.n1946 19.3944
R8886 gnd.n4940 gnd.n1946 19.3944
R8887 gnd.n4940 gnd.n1944 19.3944
R8888 gnd.n4944 gnd.n1944 19.3944
R8889 gnd.n4944 gnd.n1933 19.3944
R8890 gnd.n4956 gnd.n1933 19.3944
R8891 gnd.n4956 gnd.n1931 19.3944
R8892 gnd.n4960 gnd.n1931 19.3944
R8893 gnd.n4960 gnd.n1920 19.3944
R8894 gnd.n4972 gnd.n1920 19.3944
R8895 gnd.n4972 gnd.n1918 19.3944
R8896 gnd.n4976 gnd.n1918 19.3944
R8897 gnd.n4976 gnd.n1906 19.3944
R8898 gnd.n4988 gnd.n1906 19.3944
R8899 gnd.n4988 gnd.n1904 19.3944
R8900 gnd.n4994 gnd.n1904 19.3944
R8901 gnd.n4994 gnd.n4993 19.3944
R8902 gnd.n4993 gnd.n1875 19.3944
R8903 gnd.n5574 gnd.n1875 19.3944
R8904 gnd.n5574 gnd.n1873 19.3944
R8905 gnd.n5578 gnd.n1873 19.3944
R8906 gnd.n5578 gnd.n1861 19.3944
R8907 gnd.n5590 gnd.n1861 19.3944
R8908 gnd.n5590 gnd.n1859 19.3944
R8909 gnd.n5594 gnd.n1859 19.3944
R8910 gnd.n5594 gnd.n1846 19.3944
R8911 gnd.n5606 gnd.n1846 19.3944
R8912 gnd.n5606 gnd.n1844 19.3944
R8913 gnd.n5610 gnd.n1844 19.3944
R8914 gnd.n5610 gnd.n1831 19.3944
R8915 gnd.n5622 gnd.n1831 19.3944
R8916 gnd.n5622 gnd.n1829 19.3944
R8917 gnd.n5626 gnd.n1829 19.3944
R8918 gnd.n5626 gnd.n1817 19.3944
R8919 gnd.n5638 gnd.n1817 19.3944
R8920 gnd.n5638 gnd.n1815 19.3944
R8921 gnd.n5642 gnd.n1815 19.3944
R8922 gnd.n5642 gnd.n1802 19.3944
R8923 gnd.n5654 gnd.n1802 19.3944
R8924 gnd.n5654 gnd.n1800 19.3944
R8925 gnd.n5658 gnd.n1800 19.3944
R8926 gnd.n5658 gnd.n1787 19.3944
R8927 gnd.n5670 gnd.n1787 19.3944
R8928 gnd.n5670 gnd.n1785 19.3944
R8929 gnd.n5674 gnd.n1785 19.3944
R8930 gnd.n5674 gnd.n1772 19.3944
R8931 gnd.n5686 gnd.n1772 19.3944
R8932 gnd.n5686 gnd.n1770 19.3944
R8933 gnd.n5690 gnd.n1770 19.3944
R8934 gnd.n5690 gnd.n1758 19.3944
R8935 gnd.n5702 gnd.n1758 19.3944
R8936 gnd.n5702 gnd.n1756 19.3944
R8937 gnd.n5706 gnd.n1756 19.3944
R8938 gnd.n5706 gnd.n1743 19.3944
R8939 gnd.n5718 gnd.n1743 19.3944
R8940 gnd.n5718 gnd.n1741 19.3944
R8941 gnd.n5722 gnd.n1741 19.3944
R8942 gnd.n5722 gnd.n1730 19.3944
R8943 gnd.n5734 gnd.n1730 19.3944
R8944 gnd.n5734 gnd.n1728 19.3944
R8945 gnd.n5738 gnd.n1728 19.3944
R8946 gnd.n5738 gnd.n1718 19.3944
R8947 gnd.n5750 gnd.n1718 19.3944
R8948 gnd.n5750 gnd.n1716 19.3944
R8949 gnd.n5754 gnd.n1716 19.3944
R8950 gnd.n5754 gnd.n1704 19.3944
R8951 gnd.n5766 gnd.n1704 19.3944
R8952 gnd.n5766 gnd.n1702 19.3944
R8953 gnd.n5770 gnd.n1702 19.3944
R8954 gnd.n5770 gnd.n1691 19.3944
R8955 gnd.n5782 gnd.n1691 19.3944
R8956 gnd.n5782 gnd.n1689 19.3944
R8957 gnd.n5786 gnd.n1689 19.3944
R8958 gnd.n5786 gnd.n1677 19.3944
R8959 gnd.n5798 gnd.n1677 19.3944
R8960 gnd.n5798 gnd.n1675 19.3944
R8961 gnd.n5802 gnd.n1675 19.3944
R8962 gnd.n5802 gnd.n1664 19.3944
R8963 gnd.n5814 gnd.n1664 19.3944
R8964 gnd.n5814 gnd.n1662 19.3944
R8965 gnd.n5818 gnd.n1662 19.3944
R8966 gnd.n5818 gnd.n1651 19.3944
R8967 gnd.n5830 gnd.n1651 19.3944
R8968 gnd.n5830 gnd.n1649 19.3944
R8969 gnd.n5834 gnd.n1649 19.3944
R8970 gnd.n5834 gnd.n1637 19.3944
R8971 gnd.n5846 gnd.n1637 19.3944
R8972 gnd.n5846 gnd.n1635 19.3944
R8973 gnd.n5850 gnd.n1635 19.3944
R8974 gnd.n5850 gnd.n1624 19.3944
R8975 gnd.n5864 gnd.n1624 19.3944
R8976 gnd.n5864 gnd.n1622 19.3944
R8977 gnd.n5871 gnd.n1622 19.3944
R8978 gnd.n5871 gnd.n5870 19.3944
R8979 gnd.n5870 gnd.n1250 19.3944
R8980 gnd.n6161 gnd.n1250 19.3944
R8981 gnd.n6161 gnd.n6160 19.3944
R8982 gnd.n6160 gnd.n6159 19.3944
R8983 gnd.n6159 gnd.n1254 19.3944
R8984 gnd.n1445 gnd.n1254 19.3944
R8985 gnd.n1445 gnd.n1442 19.3944
R8986 gnd.n1449 gnd.n1442 19.3944
R8987 gnd.n1449 gnd.n1440 19.3944
R8988 gnd.n5926 gnd.n1440 19.3944
R8989 gnd.n5926 gnd.n1438 19.3944
R8990 gnd.n5932 gnd.n1438 19.3944
R8991 gnd.n5932 gnd.n5931 19.3944
R8992 gnd.n5931 gnd.n1412 19.3944
R8993 gnd.n5962 gnd.n1412 19.3944
R8994 gnd.n5962 gnd.n1410 19.3944
R8995 gnd.n5968 gnd.n1410 19.3944
R8996 gnd.n5968 gnd.n5967 19.3944
R8997 gnd.n5967 gnd.n1378 19.3944
R8998 gnd.n6023 gnd.n1378 19.3944
R8999 gnd.n6023 gnd.n1376 19.3944
R9000 gnd.n6039 gnd.n1376 19.3944
R9001 gnd.n6039 gnd.n6038 19.3944
R9002 gnd.n6038 gnd.n6037 19.3944
R9003 gnd.n6037 gnd.n6029 19.3944
R9004 gnd.n6033 gnd.n6029 19.3944
R9005 gnd.n6033 gnd.n411 19.3944
R9006 gnd.n7223 gnd.n411 19.3944
R9007 gnd.n7223 gnd.n7222 19.3944
R9008 gnd.n7222 gnd.n7221 19.3944
R9009 gnd.n7221 gnd.n415 19.3944
R9010 gnd.n7217 gnd.n415 19.3944
R9011 gnd.n7217 gnd.n7216 19.3944
R9012 gnd.n7216 gnd.n7215 19.3944
R9013 gnd.n7001 gnd.n544 19.3944
R9014 gnd.n7007 gnd.n544 19.3944
R9015 gnd.n7007 gnd.n542 19.3944
R9016 gnd.n7011 gnd.n542 19.3944
R9017 gnd.n7011 gnd.n538 19.3944
R9018 gnd.n7017 gnd.n538 19.3944
R9019 gnd.n7017 gnd.n536 19.3944
R9020 gnd.n7021 gnd.n536 19.3944
R9021 gnd.n7021 gnd.n532 19.3944
R9022 gnd.n7027 gnd.n532 19.3944
R9023 gnd.n7027 gnd.n530 19.3944
R9024 gnd.n7031 gnd.n530 19.3944
R9025 gnd.n7031 gnd.n526 19.3944
R9026 gnd.n7037 gnd.n526 19.3944
R9027 gnd.n7037 gnd.n524 19.3944
R9028 gnd.n7041 gnd.n524 19.3944
R9029 gnd.n7041 gnd.n520 19.3944
R9030 gnd.n7047 gnd.n520 19.3944
R9031 gnd.n7047 gnd.n518 19.3944
R9032 gnd.n7051 gnd.n518 19.3944
R9033 gnd.n7051 gnd.n514 19.3944
R9034 gnd.n7057 gnd.n514 19.3944
R9035 gnd.n7057 gnd.n512 19.3944
R9036 gnd.n7061 gnd.n512 19.3944
R9037 gnd.n7061 gnd.n508 19.3944
R9038 gnd.n7067 gnd.n508 19.3944
R9039 gnd.n7067 gnd.n506 19.3944
R9040 gnd.n7071 gnd.n506 19.3944
R9041 gnd.n7071 gnd.n502 19.3944
R9042 gnd.n7077 gnd.n502 19.3944
R9043 gnd.n7077 gnd.n500 19.3944
R9044 gnd.n7081 gnd.n500 19.3944
R9045 gnd.n7081 gnd.n496 19.3944
R9046 gnd.n7087 gnd.n496 19.3944
R9047 gnd.n7087 gnd.n494 19.3944
R9048 gnd.n7091 gnd.n494 19.3944
R9049 gnd.n7091 gnd.n490 19.3944
R9050 gnd.n7097 gnd.n490 19.3944
R9051 gnd.n7097 gnd.n488 19.3944
R9052 gnd.n7101 gnd.n488 19.3944
R9053 gnd.n7101 gnd.n484 19.3944
R9054 gnd.n7107 gnd.n484 19.3944
R9055 gnd.n7107 gnd.n482 19.3944
R9056 gnd.n7111 gnd.n482 19.3944
R9057 gnd.n7111 gnd.n478 19.3944
R9058 gnd.n7117 gnd.n478 19.3944
R9059 gnd.n7117 gnd.n476 19.3944
R9060 gnd.n7121 gnd.n476 19.3944
R9061 gnd.n7121 gnd.n472 19.3944
R9062 gnd.n7127 gnd.n472 19.3944
R9063 gnd.n7127 gnd.n470 19.3944
R9064 gnd.n7131 gnd.n470 19.3944
R9065 gnd.n7131 gnd.n466 19.3944
R9066 gnd.n7137 gnd.n466 19.3944
R9067 gnd.n7137 gnd.n464 19.3944
R9068 gnd.n7141 gnd.n464 19.3944
R9069 gnd.n7141 gnd.n460 19.3944
R9070 gnd.n7147 gnd.n460 19.3944
R9071 gnd.n7147 gnd.n458 19.3944
R9072 gnd.n7151 gnd.n458 19.3944
R9073 gnd.n7151 gnd.n454 19.3944
R9074 gnd.n7157 gnd.n454 19.3944
R9075 gnd.n7157 gnd.n452 19.3944
R9076 gnd.n7161 gnd.n452 19.3944
R9077 gnd.n7161 gnd.n448 19.3944
R9078 gnd.n7167 gnd.n448 19.3944
R9079 gnd.n7167 gnd.n446 19.3944
R9080 gnd.n7171 gnd.n446 19.3944
R9081 gnd.n7171 gnd.n442 19.3944
R9082 gnd.n7177 gnd.n442 19.3944
R9083 gnd.n7177 gnd.n440 19.3944
R9084 gnd.n7181 gnd.n440 19.3944
R9085 gnd.n7181 gnd.n436 19.3944
R9086 gnd.n7187 gnd.n436 19.3944
R9087 gnd.n7187 gnd.n434 19.3944
R9088 gnd.n7191 gnd.n434 19.3944
R9089 gnd.n7191 gnd.n430 19.3944
R9090 gnd.n7197 gnd.n430 19.3944
R9091 gnd.n7197 gnd.n428 19.3944
R9092 gnd.n7201 gnd.n428 19.3944
R9093 gnd.n7201 gnd.n424 19.3944
R9094 gnd.n7208 gnd.n424 19.3944
R9095 gnd.n7208 gnd.n422 19.3944
R9096 gnd.n7212 gnd.n422 19.3944
R9097 gnd.n6580 gnd.n795 19.3944
R9098 gnd.n6586 gnd.n795 19.3944
R9099 gnd.n6586 gnd.n793 19.3944
R9100 gnd.n6590 gnd.n793 19.3944
R9101 gnd.n6590 gnd.n789 19.3944
R9102 gnd.n6596 gnd.n789 19.3944
R9103 gnd.n6596 gnd.n787 19.3944
R9104 gnd.n6600 gnd.n787 19.3944
R9105 gnd.n6600 gnd.n783 19.3944
R9106 gnd.n6606 gnd.n783 19.3944
R9107 gnd.n6606 gnd.n781 19.3944
R9108 gnd.n6610 gnd.n781 19.3944
R9109 gnd.n6610 gnd.n777 19.3944
R9110 gnd.n6616 gnd.n777 19.3944
R9111 gnd.n6616 gnd.n775 19.3944
R9112 gnd.n6620 gnd.n775 19.3944
R9113 gnd.n6620 gnd.n771 19.3944
R9114 gnd.n6626 gnd.n771 19.3944
R9115 gnd.n6626 gnd.n769 19.3944
R9116 gnd.n6630 gnd.n769 19.3944
R9117 gnd.n6630 gnd.n765 19.3944
R9118 gnd.n6636 gnd.n765 19.3944
R9119 gnd.n6636 gnd.n763 19.3944
R9120 gnd.n6640 gnd.n763 19.3944
R9121 gnd.n6640 gnd.n759 19.3944
R9122 gnd.n6646 gnd.n759 19.3944
R9123 gnd.n6646 gnd.n757 19.3944
R9124 gnd.n6650 gnd.n757 19.3944
R9125 gnd.n6650 gnd.n753 19.3944
R9126 gnd.n6656 gnd.n753 19.3944
R9127 gnd.n6656 gnd.n751 19.3944
R9128 gnd.n6660 gnd.n751 19.3944
R9129 gnd.n6660 gnd.n747 19.3944
R9130 gnd.n6666 gnd.n747 19.3944
R9131 gnd.n6666 gnd.n745 19.3944
R9132 gnd.n6670 gnd.n745 19.3944
R9133 gnd.n6670 gnd.n741 19.3944
R9134 gnd.n6676 gnd.n741 19.3944
R9135 gnd.n6676 gnd.n739 19.3944
R9136 gnd.n6680 gnd.n739 19.3944
R9137 gnd.n6680 gnd.n735 19.3944
R9138 gnd.n6686 gnd.n735 19.3944
R9139 gnd.n6686 gnd.n733 19.3944
R9140 gnd.n6690 gnd.n733 19.3944
R9141 gnd.n6690 gnd.n729 19.3944
R9142 gnd.n6696 gnd.n729 19.3944
R9143 gnd.n6696 gnd.n727 19.3944
R9144 gnd.n6700 gnd.n727 19.3944
R9145 gnd.n6700 gnd.n723 19.3944
R9146 gnd.n6706 gnd.n723 19.3944
R9147 gnd.n6706 gnd.n721 19.3944
R9148 gnd.n6710 gnd.n721 19.3944
R9149 gnd.n6710 gnd.n717 19.3944
R9150 gnd.n6716 gnd.n717 19.3944
R9151 gnd.n6716 gnd.n715 19.3944
R9152 gnd.n6720 gnd.n715 19.3944
R9153 gnd.n6720 gnd.n711 19.3944
R9154 gnd.n6726 gnd.n711 19.3944
R9155 gnd.n6726 gnd.n709 19.3944
R9156 gnd.n6730 gnd.n709 19.3944
R9157 gnd.n6730 gnd.n705 19.3944
R9158 gnd.n6736 gnd.n705 19.3944
R9159 gnd.n6736 gnd.n703 19.3944
R9160 gnd.n6740 gnd.n703 19.3944
R9161 gnd.n6740 gnd.n699 19.3944
R9162 gnd.n6746 gnd.n699 19.3944
R9163 gnd.n6746 gnd.n697 19.3944
R9164 gnd.n6750 gnd.n697 19.3944
R9165 gnd.n6750 gnd.n693 19.3944
R9166 gnd.n6756 gnd.n693 19.3944
R9167 gnd.n6756 gnd.n691 19.3944
R9168 gnd.n6760 gnd.n691 19.3944
R9169 gnd.n6760 gnd.n687 19.3944
R9170 gnd.n6766 gnd.n687 19.3944
R9171 gnd.n6766 gnd.n685 19.3944
R9172 gnd.n6770 gnd.n685 19.3944
R9173 gnd.n6770 gnd.n681 19.3944
R9174 gnd.n6776 gnd.n681 19.3944
R9175 gnd.n6776 gnd.n679 19.3944
R9176 gnd.n6780 gnd.n679 19.3944
R9177 gnd.n6780 gnd.n675 19.3944
R9178 gnd.n6786 gnd.n675 19.3944
R9179 gnd.n6786 gnd.n673 19.3944
R9180 gnd.n6790 gnd.n673 19.3944
R9181 gnd.n6790 gnd.n669 19.3944
R9182 gnd.n6796 gnd.n669 19.3944
R9183 gnd.n6796 gnd.n667 19.3944
R9184 gnd.n6800 gnd.n667 19.3944
R9185 gnd.n6800 gnd.n663 19.3944
R9186 gnd.n6806 gnd.n663 19.3944
R9187 gnd.n6806 gnd.n661 19.3944
R9188 gnd.n6810 gnd.n661 19.3944
R9189 gnd.n6810 gnd.n657 19.3944
R9190 gnd.n6816 gnd.n657 19.3944
R9191 gnd.n6816 gnd.n655 19.3944
R9192 gnd.n6820 gnd.n655 19.3944
R9193 gnd.n6820 gnd.n651 19.3944
R9194 gnd.n6826 gnd.n651 19.3944
R9195 gnd.n6826 gnd.n649 19.3944
R9196 gnd.n6830 gnd.n649 19.3944
R9197 gnd.n6830 gnd.n645 19.3944
R9198 gnd.n6836 gnd.n645 19.3944
R9199 gnd.n6836 gnd.n643 19.3944
R9200 gnd.n6840 gnd.n643 19.3944
R9201 gnd.n6840 gnd.n639 19.3944
R9202 gnd.n6846 gnd.n639 19.3944
R9203 gnd.n6846 gnd.n637 19.3944
R9204 gnd.n6850 gnd.n637 19.3944
R9205 gnd.n6850 gnd.n633 19.3944
R9206 gnd.n6856 gnd.n633 19.3944
R9207 gnd.n6856 gnd.n631 19.3944
R9208 gnd.n6860 gnd.n631 19.3944
R9209 gnd.n6860 gnd.n627 19.3944
R9210 gnd.n6866 gnd.n627 19.3944
R9211 gnd.n6866 gnd.n625 19.3944
R9212 gnd.n6870 gnd.n625 19.3944
R9213 gnd.n6870 gnd.n621 19.3944
R9214 gnd.n6876 gnd.n621 19.3944
R9215 gnd.n6876 gnd.n619 19.3944
R9216 gnd.n6880 gnd.n619 19.3944
R9217 gnd.n6880 gnd.n615 19.3944
R9218 gnd.n6886 gnd.n615 19.3944
R9219 gnd.n6886 gnd.n613 19.3944
R9220 gnd.n6890 gnd.n613 19.3944
R9221 gnd.n6890 gnd.n609 19.3944
R9222 gnd.n6896 gnd.n609 19.3944
R9223 gnd.n6896 gnd.n607 19.3944
R9224 gnd.n6900 gnd.n607 19.3944
R9225 gnd.n6900 gnd.n603 19.3944
R9226 gnd.n6906 gnd.n603 19.3944
R9227 gnd.n6906 gnd.n601 19.3944
R9228 gnd.n6910 gnd.n601 19.3944
R9229 gnd.n6910 gnd.n597 19.3944
R9230 gnd.n6916 gnd.n597 19.3944
R9231 gnd.n6916 gnd.n595 19.3944
R9232 gnd.n6920 gnd.n595 19.3944
R9233 gnd.n6920 gnd.n591 19.3944
R9234 gnd.n6926 gnd.n591 19.3944
R9235 gnd.n6926 gnd.n589 19.3944
R9236 gnd.n6930 gnd.n589 19.3944
R9237 gnd.n6930 gnd.n585 19.3944
R9238 gnd.n6936 gnd.n585 19.3944
R9239 gnd.n6936 gnd.n583 19.3944
R9240 gnd.n6940 gnd.n583 19.3944
R9241 gnd.n6940 gnd.n579 19.3944
R9242 gnd.n6946 gnd.n579 19.3944
R9243 gnd.n6946 gnd.n577 19.3944
R9244 gnd.n6950 gnd.n577 19.3944
R9245 gnd.n6950 gnd.n573 19.3944
R9246 gnd.n6956 gnd.n573 19.3944
R9247 gnd.n6956 gnd.n571 19.3944
R9248 gnd.n6960 gnd.n571 19.3944
R9249 gnd.n6960 gnd.n567 19.3944
R9250 gnd.n6966 gnd.n567 19.3944
R9251 gnd.n6966 gnd.n565 19.3944
R9252 gnd.n6970 gnd.n565 19.3944
R9253 gnd.n6970 gnd.n561 19.3944
R9254 gnd.n6976 gnd.n561 19.3944
R9255 gnd.n6976 gnd.n559 19.3944
R9256 gnd.n6980 gnd.n559 19.3944
R9257 gnd.n6980 gnd.n555 19.3944
R9258 gnd.n6986 gnd.n555 19.3944
R9259 gnd.n6986 gnd.n553 19.3944
R9260 gnd.n6991 gnd.n553 19.3944
R9261 gnd.n6991 gnd.n549 19.3944
R9262 gnd.n6997 gnd.n549 19.3944
R9263 gnd.n6998 gnd.n6997 19.3944
R9264 gnd.n6152 gnd.n6151 19.3944
R9265 gnd.n6151 gnd.n6150 19.3944
R9266 gnd.n6150 gnd.n6149 19.3944
R9267 gnd.n6149 gnd.n6147 19.3944
R9268 gnd.n6147 gnd.n6144 19.3944
R9269 gnd.n6144 gnd.n6143 19.3944
R9270 gnd.n6143 gnd.n6140 19.3944
R9271 gnd.n6140 gnd.n6139 19.3944
R9272 gnd.n6139 gnd.n6136 19.3944
R9273 gnd.n6136 gnd.n6135 19.3944
R9274 gnd.n6135 gnd.n6132 19.3944
R9275 gnd.n6132 gnd.n6131 19.3944
R9276 gnd.n6131 gnd.n6128 19.3944
R9277 gnd.n6128 gnd.n6127 19.3944
R9278 gnd.n6127 gnd.n6124 19.3944
R9279 gnd.n6122 gnd.n6119 19.3944
R9280 gnd.n6119 gnd.n6118 19.3944
R9281 gnd.n6118 gnd.n6115 19.3944
R9282 gnd.n6115 gnd.n6114 19.3944
R9283 gnd.n6114 gnd.n6111 19.3944
R9284 gnd.n6111 gnd.n6110 19.3944
R9285 gnd.n6110 gnd.n6107 19.3944
R9286 gnd.n6107 gnd.n6106 19.3944
R9287 gnd.n6106 gnd.n6103 19.3944
R9288 gnd.n6103 gnd.n6102 19.3944
R9289 gnd.n6102 gnd.n6099 19.3944
R9290 gnd.n6099 gnd.n6098 19.3944
R9291 gnd.n6098 gnd.n6095 19.3944
R9292 gnd.n6095 gnd.n6094 19.3944
R9293 gnd.n6094 gnd.n6091 19.3944
R9294 gnd.n6091 gnd.n6090 19.3944
R9295 gnd.n6090 gnd.n6087 19.3944
R9296 gnd.n6087 gnd.n6086 19.3944
R9297 gnd.n1455 gnd.n1335 19.3944
R9298 gnd.n1455 gnd.n1454 19.3944
R9299 gnd.n1473 gnd.n1454 19.3944
R9300 gnd.n1473 gnd.n1472 19.3944
R9301 gnd.n1472 gnd.n1471 19.3944
R9302 gnd.n1471 gnd.n1469 19.3944
R9303 gnd.n1469 gnd.n1468 19.3944
R9304 gnd.n1468 gnd.n1466 19.3944
R9305 gnd.n1466 gnd.n1465 19.3944
R9306 gnd.n1465 gnd.n1391 19.3944
R9307 gnd.n5984 gnd.n1391 19.3944
R9308 gnd.n5984 gnd.n1389 19.3944
R9309 gnd.n5988 gnd.n1389 19.3944
R9310 gnd.n5989 gnd.n5988 19.3944
R9311 gnd.n5991 gnd.n5989 19.3944
R9312 gnd.n5991 gnd.n1387 19.3944
R9313 gnd.n5997 gnd.n1387 19.3944
R9314 gnd.n5997 gnd.n5996 19.3944
R9315 gnd.n5996 gnd.n388 19.3944
R9316 gnd.n7247 gnd.n388 19.3944
R9317 gnd.n7247 gnd.n386 19.3944
R9318 gnd.n7257 gnd.n386 19.3944
R9319 gnd.n7257 gnd.n7256 19.3944
R9320 gnd.n7256 gnd.n7255 19.3944
R9321 gnd.n7255 gnd.n354 19.3944
R9322 gnd.n7292 gnd.n354 19.3944
R9323 gnd.n7292 gnd.n352 19.3944
R9324 gnd.n7303 gnd.n352 19.3944
R9325 gnd.n7303 gnd.n7302 19.3944
R9326 gnd.n7302 gnd.n7301 19.3944
R9327 gnd.n7301 gnd.n7299 19.3944
R9328 gnd.n7299 gnd.n338 19.3944
R9329 gnd.n7322 gnd.n338 19.3944
R9330 gnd.n7322 gnd.n336 19.3944
R9331 gnd.n7391 gnd.n336 19.3944
R9332 gnd.n7391 gnd.n7390 19.3944
R9333 gnd.n7390 gnd.n7389 19.3944
R9334 gnd.n7389 gnd.n7387 19.3944
R9335 gnd.n7387 gnd.n7386 19.3944
R9336 gnd.n7386 gnd.n7384 19.3944
R9337 gnd.n7384 gnd.n7383 19.3944
R9338 gnd.n7383 gnd.n7381 19.3944
R9339 gnd.n7381 gnd.n7380 19.3944
R9340 gnd.n7380 gnd.n7378 19.3944
R9341 gnd.n7378 gnd.n7377 19.3944
R9342 gnd.n7377 gnd.n7375 19.3944
R9343 gnd.n7375 gnd.n7374 19.3944
R9344 gnd.n7374 gnd.n7372 19.3944
R9345 gnd.n7372 gnd.n7371 19.3944
R9346 gnd.n7371 gnd.n7369 19.3944
R9347 gnd.n7369 gnd.n7368 19.3944
R9348 gnd.n7368 gnd.n7366 19.3944
R9349 gnd.n7366 gnd.n7365 19.3944
R9350 gnd.n7365 gnd.n7363 19.3944
R9351 gnd.n7363 gnd.n7362 19.3944
R9352 gnd.n7362 gnd.n7360 19.3944
R9353 gnd.n7360 gnd.n7359 19.3944
R9354 gnd.n7359 gnd.n7357 19.3944
R9355 gnd.n7357 gnd.n7356 19.3944
R9356 gnd.n7356 gnd.n7354 19.3944
R9357 gnd.n7354 gnd.n7353 19.3944
R9358 gnd.n7353 gnd.n204 19.3944
R9359 gnd.n7588 gnd.n204 19.3944
R9360 gnd.n7589 gnd.n7588 19.3944
R9361 gnd.n7627 gnd.n165 19.3944
R9362 gnd.n7622 gnd.n165 19.3944
R9363 gnd.n7622 gnd.n7621 19.3944
R9364 gnd.n7621 gnd.n7620 19.3944
R9365 gnd.n7620 gnd.n172 19.3944
R9366 gnd.n7615 gnd.n172 19.3944
R9367 gnd.n7615 gnd.n7614 19.3944
R9368 gnd.n7614 gnd.n7613 19.3944
R9369 gnd.n7613 gnd.n179 19.3944
R9370 gnd.n7608 gnd.n179 19.3944
R9371 gnd.n7608 gnd.n7607 19.3944
R9372 gnd.n7607 gnd.n7606 19.3944
R9373 gnd.n7606 gnd.n186 19.3944
R9374 gnd.n7601 gnd.n186 19.3944
R9375 gnd.n7601 gnd.n7600 19.3944
R9376 gnd.n7600 gnd.n7599 19.3944
R9377 gnd.n7599 gnd.n193 19.3944
R9378 gnd.n7594 gnd.n193 19.3944
R9379 gnd.n7660 gnd.n7659 19.3944
R9380 gnd.n7659 gnd.n7658 19.3944
R9381 gnd.n7658 gnd.n137 19.3944
R9382 gnd.n7653 gnd.n137 19.3944
R9383 gnd.n7653 gnd.n7652 19.3944
R9384 gnd.n7652 gnd.n7651 19.3944
R9385 gnd.n7651 gnd.n144 19.3944
R9386 gnd.n7646 gnd.n144 19.3944
R9387 gnd.n7646 gnd.n7645 19.3944
R9388 gnd.n7645 gnd.n7644 19.3944
R9389 gnd.n7644 gnd.n151 19.3944
R9390 gnd.n7639 gnd.n151 19.3944
R9391 gnd.n7639 gnd.n7638 19.3944
R9392 gnd.n7638 gnd.n7637 19.3944
R9393 gnd.n7637 gnd.n158 19.3944
R9394 gnd.n7632 gnd.n158 19.3944
R9395 gnd.n7632 gnd.n7631 19.3944
R9396 gnd.n5912 gnd.n5907 19.3944
R9397 gnd.n5912 gnd.n5911 19.3944
R9398 gnd.n5911 gnd.n1429 19.3944
R9399 gnd.n5937 gnd.n1429 19.3944
R9400 gnd.n5937 gnd.n1427 19.3944
R9401 gnd.n5943 gnd.n1427 19.3944
R9402 gnd.n5943 gnd.n5942 19.3944
R9403 gnd.n5942 gnd.n1402 19.3944
R9404 gnd.n5974 gnd.n1402 19.3944
R9405 gnd.n5974 gnd.n1400 19.3944
R9406 gnd.n5980 gnd.n1400 19.3944
R9407 gnd.n5980 gnd.n5979 19.3944
R9408 gnd.n5979 gnd.n1368 19.3944
R9409 gnd.n6044 gnd.n1368 19.3944
R9410 gnd.n6044 gnd.n1366 19.3944
R9411 gnd.n6048 gnd.n1366 19.3944
R9412 gnd.n6048 gnd.n397 19.3944
R9413 gnd.n7237 gnd.n397 19.3944
R9414 gnd.n7237 gnd.n395 19.3944
R9415 gnd.n7243 gnd.n395 19.3944
R9416 gnd.n7243 gnd.n7242 19.3944
R9417 gnd.n7242 gnd.n364 19.3944
R9418 gnd.n7283 gnd.n364 19.3944
R9419 gnd.n7283 gnd.n362 19.3944
R9420 gnd.n7287 gnd.n362 19.3944
R9421 gnd.n7288 gnd.n7287 19.3944
R9422 gnd.n7288 gnd.n309 19.3944
R9423 gnd.n7415 gnd.n7414 19.3944
R9424 gnd.n342 gnd.n341 19.3944
R9425 gnd.n7318 gnd.n7317 19.3944
R9426 gnd.n332 gnd.n331 19.3944
R9427 gnd.n7395 gnd.n302 19.3944
R9428 gnd.n7419 gnd.n302 19.3944
R9429 gnd.n7419 gnd.n288 19.3944
R9430 gnd.n7431 gnd.n288 19.3944
R9431 gnd.n7431 gnd.n286 19.3944
R9432 gnd.n7435 gnd.n286 19.3944
R9433 gnd.n7435 gnd.n274 19.3944
R9434 gnd.n7447 gnd.n274 19.3944
R9435 gnd.n7447 gnd.n272 19.3944
R9436 gnd.n7451 gnd.n272 19.3944
R9437 gnd.n7451 gnd.n258 19.3944
R9438 gnd.n7463 gnd.n258 19.3944
R9439 gnd.n7463 gnd.n256 19.3944
R9440 gnd.n7467 gnd.n256 19.3944
R9441 gnd.n7467 gnd.n243 19.3944
R9442 gnd.n7479 gnd.n243 19.3944
R9443 gnd.n7479 gnd.n241 19.3944
R9444 gnd.n7483 gnd.n241 19.3944
R9445 gnd.n7483 gnd.n227 19.3944
R9446 gnd.n7495 gnd.n227 19.3944
R9447 gnd.n7495 gnd.n225 19.3944
R9448 gnd.n7499 gnd.n225 19.3944
R9449 gnd.n7499 gnd.n211 19.3944
R9450 gnd.n7579 gnd.n211 19.3944
R9451 gnd.n7579 gnd.n209 19.3944
R9452 gnd.n7583 gnd.n209 19.3944
R9453 gnd.n7583 gnd.n132 19.3944
R9454 gnd.n7663 gnd.n132 19.3944
R9455 gnd.n4194 gnd.n4193 19.3944
R9456 gnd.n4193 gnd.n3980 19.3944
R9457 gnd.n4188 gnd.n3980 19.3944
R9458 gnd.n4188 gnd.n4187 19.3944
R9459 gnd.n4187 gnd.n3985 19.3944
R9460 gnd.n4182 gnd.n3985 19.3944
R9461 gnd.n4182 gnd.n4181 19.3944
R9462 gnd.n4181 gnd.n4180 19.3944
R9463 gnd.n4180 gnd.n3991 19.3944
R9464 gnd.n4174 gnd.n3991 19.3944
R9465 gnd.n4174 gnd.n4173 19.3944
R9466 gnd.n4173 gnd.n4172 19.3944
R9467 gnd.n4172 gnd.n3997 19.3944
R9468 gnd.n4166 gnd.n3997 19.3944
R9469 gnd.n4166 gnd.n4165 19.3944
R9470 gnd.n4165 gnd.n4164 19.3944
R9471 gnd.n4164 gnd.n4003 19.3944
R9472 gnd.n4158 gnd.n4157 19.3944
R9473 gnd.n4157 gnd.n4156 19.3944
R9474 gnd.n4156 gnd.n4012 19.3944
R9475 gnd.n4150 gnd.n4012 19.3944
R9476 gnd.n4150 gnd.n4149 19.3944
R9477 gnd.n4149 gnd.n4148 19.3944
R9478 gnd.n4148 gnd.n4018 19.3944
R9479 gnd.n4142 gnd.n4018 19.3944
R9480 gnd.n4142 gnd.n4141 19.3944
R9481 gnd.n4141 gnd.n4140 19.3944
R9482 gnd.n4140 gnd.n4024 19.3944
R9483 gnd.n4134 gnd.n4024 19.3944
R9484 gnd.n4134 gnd.n4133 19.3944
R9485 gnd.n4133 gnd.n4132 19.3944
R9486 gnd.n4132 gnd.n4030 19.3944
R9487 gnd.n4126 gnd.n4030 19.3944
R9488 gnd.n4126 gnd.n4125 19.3944
R9489 gnd.n4125 gnd.n4124 19.3944
R9490 gnd.n4201 gnd.n2336 19.3944
R9491 gnd.n4205 gnd.n2336 19.3944
R9492 gnd.n4205 gnd.n2323 19.3944
R9493 gnd.n4217 gnd.n2323 19.3944
R9494 gnd.n4217 gnd.n2321 19.3944
R9495 gnd.n4221 gnd.n2321 19.3944
R9496 gnd.n4221 gnd.n2306 19.3944
R9497 gnd.n4233 gnd.n2306 19.3944
R9498 gnd.n4233 gnd.n2304 19.3944
R9499 gnd.n4237 gnd.n2304 19.3944
R9500 gnd.n4237 gnd.n2291 19.3944
R9501 gnd.n4249 gnd.n2291 19.3944
R9502 gnd.n4249 gnd.n2289 19.3944
R9503 gnd.n4253 gnd.n2289 19.3944
R9504 gnd.n4253 gnd.n2274 19.3944
R9505 gnd.n4265 gnd.n2274 19.3944
R9506 gnd.n4265 gnd.n2272 19.3944
R9507 gnd.n4269 gnd.n2272 19.3944
R9508 gnd.n4269 gnd.n2259 19.3944
R9509 gnd.n4281 gnd.n2259 19.3944
R9510 gnd.n4281 gnd.n2257 19.3944
R9511 gnd.n4285 gnd.n2257 19.3944
R9512 gnd.n4285 gnd.n2242 19.3944
R9513 gnd.n4298 gnd.n2242 19.3944
R9514 gnd.n4298 gnd.n2240 19.3944
R9515 gnd.n4302 gnd.n2240 19.3944
R9516 gnd.n4302 gnd.n2228 19.3944
R9517 gnd.n4314 gnd.n2228 19.3944
R9518 gnd.n4314 gnd.n2226 19.3944
R9519 gnd.n4319 gnd.n2226 19.3944
R9520 gnd.n4319 gnd.n4318 19.3944
R9521 gnd.n4318 gnd.n2203 19.3944
R9522 gnd.n2203 gnd.n2201 19.3944
R9523 gnd.n4346 gnd.n2201 19.3944
R9524 gnd.n4346 gnd.n4345 19.3944
R9525 gnd.n4345 gnd.n4344 19.3944
R9526 gnd.n4344 gnd.n4343 19.3944
R9527 gnd.n4343 gnd.n4341 19.3944
R9528 gnd.n4341 gnd.n989 19.3944
R9529 gnd.n6394 gnd.n989 19.3944
R9530 gnd.n6394 gnd.n6393 19.3944
R9531 gnd.n6393 gnd.n6392 19.3944
R9532 gnd.n6392 gnd.n993 19.3944
R9533 gnd.n6382 gnd.n993 19.3944
R9534 gnd.n6382 gnd.n6381 19.3944
R9535 gnd.n6381 gnd.n6380 19.3944
R9536 gnd.n6380 gnd.n1013 19.3944
R9537 gnd.n6370 gnd.n1013 19.3944
R9538 gnd.n6370 gnd.n6369 19.3944
R9539 gnd.n6369 gnd.n6368 19.3944
R9540 gnd.n6368 gnd.n1035 19.3944
R9541 gnd.n6358 gnd.n1035 19.3944
R9542 gnd.n6358 gnd.n6357 19.3944
R9543 gnd.n6357 gnd.n6356 19.3944
R9544 gnd.n6356 gnd.n1055 19.3944
R9545 gnd.n6346 gnd.n1055 19.3944
R9546 gnd.n6346 gnd.n6345 19.3944
R9547 gnd.n6345 gnd.n6344 19.3944
R9548 gnd.n6344 gnd.n1077 19.3944
R9549 gnd.n6334 gnd.n1077 19.3944
R9550 gnd.n6334 gnd.n6333 19.3944
R9551 gnd.n6333 gnd.n6332 19.3944
R9552 gnd.n6332 gnd.n1098 19.3944
R9553 gnd.n6322 gnd.n1098 19.3944
R9554 gnd.n3837 gnd.n3836 19.3944
R9555 gnd.n3842 gnd.n3837 19.3944
R9556 gnd.n3842 gnd.n3834 19.3944
R9557 gnd.n3846 gnd.n3834 19.3944
R9558 gnd.n3846 gnd.n3832 19.3944
R9559 gnd.n3852 gnd.n3832 19.3944
R9560 gnd.n3852 gnd.n3830 19.3944
R9561 gnd.n3856 gnd.n3830 19.3944
R9562 gnd.n3856 gnd.n3828 19.3944
R9563 gnd.n3862 gnd.n3828 19.3944
R9564 gnd.n3862 gnd.n3826 19.3944
R9565 gnd.n3866 gnd.n3826 19.3944
R9566 gnd.n3866 gnd.n3824 19.3944
R9567 gnd.n3872 gnd.n3824 19.3944
R9568 gnd.n3872 gnd.n3822 19.3944
R9569 gnd.n3876 gnd.n3822 19.3944
R9570 gnd.n3975 gnd.n3816 19.3944
R9571 gnd.n3975 gnd.n3974 19.3944
R9572 gnd.n3974 gnd.n3973 19.3944
R9573 gnd.n3973 gnd.n3971 19.3944
R9574 gnd.n3971 gnd.n3970 19.3944
R9575 gnd.n3970 gnd.n3968 19.3944
R9576 gnd.n3968 gnd.n3967 19.3944
R9577 gnd.n3967 gnd.n3965 19.3944
R9578 gnd.n3965 gnd.n3964 19.3944
R9579 gnd.n3964 gnd.n3962 19.3944
R9580 gnd.n3962 gnd.n3961 19.3944
R9581 gnd.n3961 gnd.n3959 19.3944
R9582 gnd.n3959 gnd.n3958 19.3944
R9583 gnd.n3958 gnd.n3956 19.3944
R9584 gnd.n3956 gnd.n3955 19.3944
R9585 gnd.n3955 gnd.n3953 19.3944
R9586 gnd.n3953 gnd.n3952 19.3944
R9587 gnd.n3952 gnd.n3950 19.3944
R9588 gnd.n3950 gnd.n3949 19.3944
R9589 gnd.n3949 gnd.n3947 19.3944
R9590 gnd.n3947 gnd.n3946 19.3944
R9591 gnd.n3946 gnd.n3944 19.3944
R9592 gnd.n3944 gnd.n3943 19.3944
R9593 gnd.n3943 gnd.n3941 19.3944
R9594 gnd.n3941 gnd.n3940 19.3944
R9595 gnd.n3940 gnd.n3938 19.3944
R9596 gnd.n3938 gnd.n3937 19.3944
R9597 gnd.n3937 gnd.n3935 19.3944
R9598 gnd.n3935 gnd.n3934 19.3944
R9599 gnd.n3934 gnd.n3932 19.3944
R9600 gnd.n3932 gnd.n3931 19.3944
R9601 gnd.n3931 gnd.n3929 19.3944
R9602 gnd.n3929 gnd.n3916 19.3944
R9603 gnd.n3925 gnd.n3916 19.3944
R9604 gnd.n3925 gnd.n3924 19.3944
R9605 gnd.n3924 gnd.n3923 19.3944
R9606 gnd.n3923 gnd.n3920 19.3944
R9607 gnd.n3920 gnd.n2185 19.3944
R9608 gnd.n4366 gnd.n2185 19.3944
R9609 gnd.n4366 gnd.n2183 19.3944
R9610 gnd.n4370 gnd.n2183 19.3944
R9611 gnd.n4370 gnd.n2173 19.3944
R9612 gnd.n4411 gnd.n2173 19.3944
R9613 gnd.n4411 gnd.n2174 19.3944
R9614 gnd.n4407 gnd.n2174 19.3944
R9615 gnd.n4407 gnd.n4406 19.3944
R9616 gnd.n4406 gnd.n4405 19.3944
R9617 gnd.n4405 gnd.n4400 19.3944
R9618 gnd.n4401 gnd.n4400 19.3944
R9619 gnd.n4401 gnd.n2152 19.3944
R9620 gnd.n4460 gnd.n2152 19.3944
R9621 gnd.n4460 gnd.n2153 19.3944
R9622 gnd.n4456 gnd.n2153 19.3944
R9623 gnd.n4456 gnd.n4455 19.3944
R9624 gnd.n4455 gnd.n4454 19.3944
R9625 gnd.n4454 gnd.n2139 19.3944
R9626 gnd.n4515 gnd.n2139 19.3944
R9627 gnd.n4515 gnd.n2137 19.3944
R9628 gnd.n4519 gnd.n2137 19.3944
R9629 gnd.n4519 gnd.n2133 19.3944
R9630 gnd.n4532 gnd.n2133 19.3944
R9631 gnd.n4532 gnd.n2130 19.3944
R9632 gnd.n4566 gnd.n2130 19.3944
R9633 gnd.n4566 gnd.n2131 19.3944
R9634 gnd.n4115 gnd.n4114 19.3944
R9635 gnd.n4114 gnd.n4113 19.3944
R9636 gnd.n4113 gnd.n4112 19.3944
R9637 gnd.n4112 gnd.n4110 19.3944
R9638 gnd.n4110 gnd.n4109 19.3944
R9639 gnd.n4109 gnd.n4107 19.3944
R9640 gnd.n4107 gnd.n4106 19.3944
R9641 gnd.n4106 gnd.n4104 19.3944
R9642 gnd.n4104 gnd.n4103 19.3944
R9643 gnd.n4103 gnd.n4101 19.3944
R9644 gnd.n4101 gnd.n4100 19.3944
R9645 gnd.n4100 gnd.n4098 19.3944
R9646 gnd.n4098 gnd.n4097 19.3944
R9647 gnd.n4097 gnd.n4095 19.3944
R9648 gnd.n4095 gnd.n4094 19.3944
R9649 gnd.n4094 gnd.n4092 19.3944
R9650 gnd.n4092 gnd.n4091 19.3944
R9651 gnd.n4091 gnd.n4089 19.3944
R9652 gnd.n4089 gnd.n4088 19.3944
R9653 gnd.n4088 gnd.n4086 19.3944
R9654 gnd.n4086 gnd.n4085 19.3944
R9655 gnd.n4085 gnd.n4083 19.3944
R9656 gnd.n4083 gnd.n4082 19.3944
R9657 gnd.n4082 gnd.n4080 19.3944
R9658 gnd.n4080 gnd.n4079 19.3944
R9659 gnd.n4079 gnd.n4077 19.3944
R9660 gnd.n4077 gnd.n4076 19.3944
R9661 gnd.n4076 gnd.n4074 19.3944
R9662 gnd.n4074 gnd.n4073 19.3944
R9663 gnd.n4073 gnd.n4071 19.3944
R9664 gnd.n4071 gnd.n2206 19.3944
R9665 gnd.n4331 gnd.n2206 19.3944
R9666 gnd.n4331 gnd.n2211 19.3944
R9667 gnd.n2211 gnd.n2210 19.3944
R9668 gnd.n2210 gnd.n2209 19.3944
R9669 gnd.n2209 gnd.n2188 19.3944
R9670 gnd.n4358 gnd.n2188 19.3944
R9671 gnd.n4358 gnd.n2186 19.3944
R9672 gnd.n4362 gnd.n2186 19.3944
R9673 gnd.n4362 gnd.n2182 19.3944
R9674 gnd.n4384 gnd.n2182 19.3944
R9675 gnd.n4384 gnd.n2180 19.3944
R9676 gnd.n4388 gnd.n2180 19.3944
R9677 gnd.n4389 gnd.n4388 19.3944
R9678 gnd.n4392 gnd.n4389 19.3944
R9679 gnd.n4392 gnd.n2178 19.3944
R9680 gnd.n4396 gnd.n2178 19.3944
R9681 gnd.n4396 gnd.n2161 19.3944
R9682 gnd.n4433 gnd.n2161 19.3944
R9683 gnd.n4433 gnd.n2159 19.3944
R9684 gnd.n4437 gnd.n2159 19.3944
R9685 gnd.n4438 gnd.n4437 19.3944
R9686 gnd.n4441 gnd.n4438 19.3944
R9687 gnd.n4441 gnd.n2157 19.3944
R9688 gnd.n4449 gnd.n2157 19.3944
R9689 gnd.n4449 gnd.n4448 19.3944
R9690 gnd.n4448 gnd.n4447 19.3944
R9691 gnd.n4447 gnd.n2136 19.3944
R9692 gnd.n4523 gnd.n2136 19.3944
R9693 gnd.n4523 gnd.n2134 19.3944
R9694 gnd.n4528 gnd.n2134 19.3944
R9695 gnd.n4528 gnd.n2128 19.3944
R9696 gnd.n4570 gnd.n2128 19.3944
R9697 gnd.n4571 gnd.n4570 19.3944
R9698 gnd.n4613 gnd.n2102 19.3944
R9699 gnd.n4613 gnd.n4610 19.3944
R9700 gnd.n4610 gnd.n4607 19.3944
R9701 gnd.n4607 gnd.n4606 19.3944
R9702 gnd.n4606 gnd.n4603 19.3944
R9703 gnd.n4603 gnd.n4602 19.3944
R9704 gnd.n4602 gnd.n4599 19.3944
R9705 gnd.n4599 gnd.n4598 19.3944
R9706 gnd.n4598 gnd.n4595 19.3944
R9707 gnd.n4595 gnd.n4594 19.3944
R9708 gnd.n4594 gnd.n4591 19.3944
R9709 gnd.n4591 gnd.n4590 19.3944
R9710 gnd.n4590 gnd.n4587 19.3944
R9711 gnd.n4587 gnd.n4586 19.3944
R9712 gnd.n4586 gnd.n4583 19.3944
R9713 gnd.n4583 gnd.n4582 19.3944
R9714 gnd.n4582 gnd.n4579 19.3944
R9715 gnd.n4579 gnd.n4578 19.3944
R9716 gnd.n2085 gnd.n2084 19.3944
R9717 gnd.n4844 gnd.n2084 19.3944
R9718 gnd.n4844 gnd.n4843 19.3944
R9719 gnd.n4843 gnd.n4842 19.3944
R9720 gnd.n4842 gnd.n4839 19.3944
R9721 gnd.n4839 gnd.n4838 19.3944
R9722 gnd.n4838 gnd.n4835 19.3944
R9723 gnd.n4835 gnd.n4834 19.3944
R9724 gnd.n4834 gnd.n4831 19.3944
R9725 gnd.n4831 gnd.n4830 19.3944
R9726 gnd.n4830 gnd.n4827 19.3944
R9727 gnd.n4827 gnd.n4826 19.3944
R9728 gnd.n4826 gnd.n4823 19.3944
R9729 gnd.n4823 gnd.n4822 19.3944
R9730 gnd.n4822 gnd.n4819 19.3944
R9731 gnd.n4197 gnd.n2331 19.3944
R9732 gnd.n4209 gnd.n2331 19.3944
R9733 gnd.n4209 gnd.n2329 19.3944
R9734 gnd.n4213 gnd.n2329 19.3944
R9735 gnd.n4213 gnd.n2315 19.3944
R9736 gnd.n4225 gnd.n2315 19.3944
R9737 gnd.n4225 gnd.n2313 19.3944
R9738 gnd.n4229 gnd.n2313 19.3944
R9739 gnd.n4229 gnd.n2299 19.3944
R9740 gnd.n4241 gnd.n2299 19.3944
R9741 gnd.n4241 gnd.n2297 19.3944
R9742 gnd.n4245 gnd.n2297 19.3944
R9743 gnd.n4245 gnd.n2283 19.3944
R9744 gnd.n4257 gnd.n2283 19.3944
R9745 gnd.n4257 gnd.n2281 19.3944
R9746 gnd.n4261 gnd.n2281 19.3944
R9747 gnd.n4261 gnd.n2267 19.3944
R9748 gnd.n4273 gnd.n2267 19.3944
R9749 gnd.n4273 gnd.n2265 19.3944
R9750 gnd.n4277 gnd.n2265 19.3944
R9751 gnd.n4277 gnd.n2251 19.3944
R9752 gnd.n4289 gnd.n2251 19.3944
R9753 gnd.n4289 gnd.n2249 19.3944
R9754 gnd.n4294 gnd.n2249 19.3944
R9755 gnd.n4294 gnd.n2234 19.3944
R9756 gnd.n4306 gnd.n2234 19.3944
R9757 gnd.n4307 gnd.n4306 19.3944
R9758 gnd.n4310 gnd.n4309 19.3944
R9759 gnd.n4324 gnd.n4323 19.3944
R9760 gnd.n4327 gnd.n4326 19.3944
R9761 gnd.n4351 gnd.n4350 19.3944
R9762 gnd.n4353 gnd.n977 19.3944
R9763 gnd.n6400 gnd.n977 19.3944
R9764 gnd.n6400 gnd.n6399 19.3944
R9765 gnd.n6399 gnd.n6398 19.3944
R9766 gnd.n6398 gnd.n981 19.3944
R9767 gnd.n6388 gnd.n981 19.3944
R9768 gnd.n6388 gnd.n6387 19.3944
R9769 gnd.n6387 gnd.n6386 19.3944
R9770 gnd.n6386 gnd.n1003 19.3944
R9771 gnd.n6376 gnd.n1003 19.3944
R9772 gnd.n6376 gnd.n6375 19.3944
R9773 gnd.n6375 gnd.n6374 19.3944
R9774 gnd.n6374 gnd.n1024 19.3944
R9775 gnd.n6364 gnd.n1024 19.3944
R9776 gnd.n6364 gnd.n6363 19.3944
R9777 gnd.n6363 gnd.n6362 19.3944
R9778 gnd.n6362 gnd.n1045 19.3944
R9779 gnd.n6352 gnd.n1045 19.3944
R9780 gnd.n6352 gnd.n6351 19.3944
R9781 gnd.n6351 gnd.n6350 19.3944
R9782 gnd.n6350 gnd.n1066 19.3944
R9783 gnd.n6340 gnd.n1066 19.3944
R9784 gnd.n6340 gnd.n6339 19.3944
R9785 gnd.n6339 gnd.n6338 19.3944
R9786 gnd.n6338 gnd.n1087 19.3944
R9787 gnd.n6328 gnd.n1087 19.3944
R9788 gnd.n6328 gnd.n6327 19.3944
R9789 gnd.n6327 gnd.n6326 19.3944
R9790 gnd.n6577 gnd.n6576 19.3944
R9791 gnd.n6576 gnd.n800 19.3944
R9792 gnd.n6570 gnd.n800 19.3944
R9793 gnd.n6570 gnd.n6569 19.3944
R9794 gnd.n6569 gnd.n6568 19.3944
R9795 gnd.n6568 gnd.n808 19.3944
R9796 gnd.n6562 gnd.n808 19.3944
R9797 gnd.n6562 gnd.n6561 19.3944
R9798 gnd.n6561 gnd.n6560 19.3944
R9799 gnd.n6560 gnd.n816 19.3944
R9800 gnd.n6554 gnd.n816 19.3944
R9801 gnd.n6554 gnd.n6553 19.3944
R9802 gnd.n6553 gnd.n6552 19.3944
R9803 gnd.n6552 gnd.n824 19.3944
R9804 gnd.n6546 gnd.n824 19.3944
R9805 gnd.n6546 gnd.n6545 19.3944
R9806 gnd.n6545 gnd.n6544 19.3944
R9807 gnd.n6544 gnd.n832 19.3944
R9808 gnd.n6538 gnd.n832 19.3944
R9809 gnd.n6538 gnd.n6537 19.3944
R9810 gnd.n6537 gnd.n6536 19.3944
R9811 gnd.n6536 gnd.n840 19.3944
R9812 gnd.n6530 gnd.n840 19.3944
R9813 gnd.n6530 gnd.n6529 19.3944
R9814 gnd.n6529 gnd.n6528 19.3944
R9815 gnd.n6528 gnd.n848 19.3944
R9816 gnd.n6522 gnd.n848 19.3944
R9817 gnd.n6522 gnd.n6521 19.3944
R9818 gnd.n6521 gnd.n6520 19.3944
R9819 gnd.n6520 gnd.n856 19.3944
R9820 gnd.n6514 gnd.n856 19.3944
R9821 gnd.n6514 gnd.n6513 19.3944
R9822 gnd.n6513 gnd.n6512 19.3944
R9823 gnd.n6512 gnd.n864 19.3944
R9824 gnd.n6506 gnd.n864 19.3944
R9825 gnd.n6506 gnd.n6505 19.3944
R9826 gnd.n6505 gnd.n6504 19.3944
R9827 gnd.n6504 gnd.n872 19.3944
R9828 gnd.n6498 gnd.n872 19.3944
R9829 gnd.n6498 gnd.n6497 19.3944
R9830 gnd.n6497 gnd.n6496 19.3944
R9831 gnd.n6496 gnd.n880 19.3944
R9832 gnd.n6490 gnd.n880 19.3944
R9833 gnd.n6490 gnd.n6489 19.3944
R9834 gnd.n6489 gnd.n6488 19.3944
R9835 gnd.n6488 gnd.n888 19.3944
R9836 gnd.n6482 gnd.n888 19.3944
R9837 gnd.n6482 gnd.n6481 19.3944
R9838 gnd.n6481 gnd.n6480 19.3944
R9839 gnd.n6480 gnd.n896 19.3944
R9840 gnd.n6474 gnd.n896 19.3944
R9841 gnd.n6474 gnd.n6473 19.3944
R9842 gnd.n6473 gnd.n6472 19.3944
R9843 gnd.n6472 gnd.n904 19.3944
R9844 gnd.n6466 gnd.n904 19.3944
R9845 gnd.n6466 gnd.n6465 19.3944
R9846 gnd.n6465 gnd.n6464 19.3944
R9847 gnd.n6464 gnd.n912 19.3944
R9848 gnd.n6458 gnd.n912 19.3944
R9849 gnd.n6458 gnd.n6457 19.3944
R9850 gnd.n6457 gnd.n6456 19.3944
R9851 gnd.n6456 gnd.n920 19.3944
R9852 gnd.n6450 gnd.n920 19.3944
R9853 gnd.n6450 gnd.n6449 19.3944
R9854 gnd.n6449 gnd.n6448 19.3944
R9855 gnd.n6448 gnd.n928 19.3944
R9856 gnd.n6442 gnd.n928 19.3944
R9857 gnd.n6442 gnd.n6441 19.3944
R9858 gnd.n6441 gnd.n6440 19.3944
R9859 gnd.n6440 gnd.n936 19.3944
R9860 gnd.n6434 gnd.n936 19.3944
R9861 gnd.n6434 gnd.n6433 19.3944
R9862 gnd.n6433 gnd.n6432 19.3944
R9863 gnd.n6432 gnd.n944 19.3944
R9864 gnd.n6426 gnd.n944 19.3944
R9865 gnd.n6426 gnd.n6425 19.3944
R9866 gnd.n6425 gnd.n6424 19.3944
R9867 gnd.n6424 gnd.n952 19.3944
R9868 gnd.n6418 gnd.n952 19.3944
R9869 gnd.n6418 gnd.n6417 19.3944
R9870 gnd.n6417 gnd.n6416 19.3944
R9871 gnd.n6416 gnd.n960 19.3944
R9872 gnd.n6410 gnd.n960 19.3944
R9873 gnd.n6410 gnd.n6409 19.3944
R9874 gnd.n6317 gnd.n6316 19.3944
R9875 gnd.n6316 gnd.n6315 19.3944
R9876 gnd.n6315 gnd.n1121 19.3944
R9877 gnd.n6311 gnd.n1121 19.3944
R9878 gnd.n6311 gnd.n6310 19.3944
R9879 gnd.n6310 gnd.n6309 19.3944
R9880 gnd.n6309 gnd.n1126 19.3944
R9881 gnd.n6305 gnd.n1126 19.3944
R9882 gnd.n6305 gnd.n6304 19.3944
R9883 gnd.n6304 gnd.n6303 19.3944
R9884 gnd.n6303 gnd.n1131 19.3944
R9885 gnd.n6299 gnd.n1131 19.3944
R9886 gnd.n6299 gnd.n6298 19.3944
R9887 gnd.n6298 gnd.n6297 19.3944
R9888 gnd.n6297 gnd.n1136 19.3944
R9889 gnd.n6293 gnd.n1136 19.3944
R9890 gnd.n6293 gnd.n6292 19.3944
R9891 gnd.n6292 gnd.n6291 19.3944
R9892 gnd.n6291 gnd.n1141 19.3944
R9893 gnd.n6287 gnd.n1141 19.3944
R9894 gnd.n6287 gnd.n6286 19.3944
R9895 gnd.n6286 gnd.n6285 19.3944
R9896 gnd.n6285 gnd.n1146 19.3944
R9897 gnd.n6281 gnd.n1146 19.3944
R9898 gnd.n6281 gnd.n6280 19.3944
R9899 gnd.n6280 gnd.n6279 19.3944
R9900 gnd.n6279 gnd.n1151 19.3944
R9901 gnd.n6275 gnd.n1151 19.3944
R9902 gnd.n6275 gnd.n6274 19.3944
R9903 gnd.n6274 gnd.n6273 19.3944
R9904 gnd.n6273 gnd.n1156 19.3944
R9905 gnd.n6269 gnd.n1156 19.3944
R9906 gnd.n6269 gnd.n6268 19.3944
R9907 gnd.n6268 gnd.n6267 19.3944
R9908 gnd.n6267 gnd.n1161 19.3944
R9909 gnd.n6263 gnd.n1161 19.3944
R9910 gnd.n6263 gnd.n6262 19.3944
R9911 gnd.n6262 gnd.n6261 19.3944
R9912 gnd.n6261 gnd.n1166 19.3944
R9913 gnd.n6257 gnd.n1166 19.3944
R9914 gnd.n6257 gnd.n6256 19.3944
R9915 gnd.n6256 gnd.n6255 19.3944
R9916 gnd.n6255 gnd.n1171 19.3944
R9917 gnd.n6251 gnd.n1171 19.3944
R9918 gnd.n6251 gnd.n6250 19.3944
R9919 gnd.n6250 gnd.n6249 19.3944
R9920 gnd.n6249 gnd.n1176 19.3944
R9921 gnd.n6245 gnd.n1176 19.3944
R9922 gnd.n6245 gnd.n6244 19.3944
R9923 gnd.n6244 gnd.n6243 19.3944
R9924 gnd.n6243 gnd.n1181 19.3944
R9925 gnd.n6239 gnd.n1181 19.3944
R9926 gnd.n6239 gnd.n6238 19.3944
R9927 gnd.n6238 gnd.n6237 19.3944
R9928 gnd.n6237 gnd.n1186 19.3944
R9929 gnd.n6233 gnd.n1186 19.3944
R9930 gnd.n6233 gnd.n6232 19.3944
R9931 gnd.n6232 gnd.n6231 19.3944
R9932 gnd.n6231 gnd.n1191 19.3944
R9933 gnd.n6227 gnd.n1191 19.3944
R9934 gnd.n6227 gnd.n6226 19.3944
R9935 gnd.n6226 gnd.n6225 19.3944
R9936 gnd.n6225 gnd.n1196 19.3944
R9937 gnd.n6221 gnd.n1196 19.3944
R9938 gnd.n6221 gnd.n6220 19.3944
R9939 gnd.n6220 gnd.n6219 19.3944
R9940 gnd.n6219 gnd.n1201 19.3944
R9941 gnd.n6215 gnd.n1201 19.3944
R9942 gnd.n6215 gnd.n6214 19.3944
R9943 gnd.n6214 gnd.n6213 19.3944
R9944 gnd.n6213 gnd.n1206 19.3944
R9945 gnd.n6209 gnd.n1206 19.3944
R9946 gnd.n6209 gnd.n6208 19.3944
R9947 gnd.n6208 gnd.n6207 19.3944
R9948 gnd.n6207 gnd.n1211 19.3944
R9949 gnd.n6203 gnd.n1211 19.3944
R9950 gnd.n6203 gnd.n6202 19.3944
R9951 gnd.n6202 gnd.n6201 19.3944
R9952 gnd.n6201 gnd.n1216 19.3944
R9953 gnd.n6197 gnd.n1216 19.3944
R9954 gnd.n6197 gnd.n6196 19.3944
R9955 gnd.n6196 gnd.n6195 19.3944
R9956 gnd.n6195 gnd.n1221 19.3944
R9957 gnd.n6191 gnd.n1221 19.3944
R9958 gnd.n6191 gnd.n6190 19.3944
R9959 gnd.n6190 gnd.n6189 19.3944
R9960 gnd.n6189 gnd.n1226 19.3944
R9961 gnd.n6185 gnd.n1226 19.3944
R9962 gnd.n6185 gnd.n6184 19.3944
R9963 gnd.n6184 gnd.n6183 19.3944
R9964 gnd.n6183 gnd.n1231 19.3944
R9965 gnd.n6179 gnd.n1231 19.3944
R9966 gnd.n6179 gnd.n6178 19.3944
R9967 gnd.n6178 gnd.n6177 19.3944
R9968 gnd.n6177 gnd.n1236 19.3944
R9969 gnd.n6173 gnd.n1236 19.3944
R9970 gnd.n6173 gnd.n6172 19.3944
R9971 gnd.n6172 gnd.n6171 19.3944
R9972 gnd.n6171 gnd.n1241 19.3944
R9973 gnd.n6167 gnd.n1241 19.3944
R9974 gnd.n6167 gnd.n6166 19.3944
R9975 gnd.n5889 gnd.n1614 19.3944
R9976 gnd.n5885 gnd.n1614 19.3944
R9977 gnd.n5885 gnd.n5884 19.3944
R9978 gnd.n1530 gnd.n1514 19.3944
R9979 gnd.n1530 gnd.n1512 19.3944
R9980 gnd.n1536 gnd.n1512 19.3944
R9981 gnd.n1536 gnd.n1507 19.3944
R9982 gnd.n1549 gnd.n1507 19.3944
R9983 gnd.n1549 gnd.n1505 19.3944
R9984 gnd.n1555 gnd.n1505 19.3944
R9985 gnd.n1555 gnd.n1500 19.3944
R9986 gnd.n1568 gnd.n1500 19.3944
R9987 gnd.n1568 gnd.n1498 19.3944
R9988 gnd.n1574 gnd.n1498 19.3944
R9989 gnd.n1574 gnd.n1494 19.3944
R9990 gnd.n1584 gnd.n1494 19.3944
R9991 gnd.n1584 gnd.n1492 19.3944
R9992 gnd.n1590 gnd.n1492 19.3944
R9993 gnd.n1590 gnd.n1482 19.3944
R9994 gnd.n1598 gnd.n1482 19.3944
R9995 gnd.n1598 gnd.n1480 19.3944
R9996 gnd.n5900 gnd.n1480 19.3944
R9997 gnd.n5900 gnd.n5899 19.3944
R9998 gnd.n5899 gnd.n5898 19.3944
R9999 gnd.n5898 gnd.n1606 19.3944
R10000 gnd.n5894 gnd.n1606 19.3944
R10001 gnd.n5894 gnd.n5893 19.3944
R10002 gnd.n6412 gnd.n962 19.1977
R10003 gnd.n5073 gnd.n1805 19.1199
R10004 gnd.n5692 gnd.n1768 19.1199
R10005 gnd.n5161 gnd.n1706 19.1199
R10006 gnd.n3199 gnd.t16 18.8012
R10007 gnd.n3184 gnd.t39 18.8012
R10008 gnd.n4746 gnd.n4744 18.5761
R10009 gnd.n5375 gnd.n5374 18.5761
R10010 gnd.n3043 gnd.n3042 18.4825
R10011 gnd.n6124 gnd.n6123 18.4247
R10012 gnd.n4819 gnd.n4818 18.4247
R10013 gnd.n7542 gnd.n124 18.2308
R10014 gnd.n1594 gnd.n1593 18.2308
R10015 gnd.n4857 gnd.n2038 18.2308
R10016 gnd.n3876 gnd.n3820 18.2308
R10017 gnd.t58 gnd.n2723 18.1639
R10018 gnd.n5596 gnd.n1855 17.8452
R10019 gnd.n5080 gnd.n1798 17.8452
R10020 gnd.n5684 gnd.n1775 17.8452
R10021 gnd.n5411 gnd.n1713 17.8452
R10022 gnd.n2751 gnd.t18 17.5266
R10023 gnd.t0 gnd.n1833 17.2079
R10024 gnd.n5135 gnd.t8 17.2079
R10025 gnd.n5397 gnd.t270 17.2079
R10026 gnd.n3150 gnd.t215 16.8893
R10027 gnd.t122 gnd.n1910 16.8893
R10028 gnd.n5604 gnd.n1848 16.5706
R10029 gnd.t208 gnd.n5525 16.5706
R10030 gnd.n5087 gnd.n1790 16.5706
R10031 gnd.n5676 gnd.n1783 16.5706
R10032 gnd.n5440 gnd.t27 16.5706
R10033 gnd.n5148 gnd.n1720 16.5706
R10034 gnd.n2978 gnd.t295 16.2519
R10035 gnd.n2678 gnd.t88 16.2519
R10036 gnd.t218 gnd.t252 16.2519
R10037 gnd.t209 gnd.n1819 15.9333
R10038 gnd.n5448 gnd.t28 15.9333
R10039 gnd.n3665 gnd.n3663 15.6674
R10040 gnd.n3633 gnd.n3631 15.6674
R10041 gnd.n3601 gnd.n3599 15.6674
R10042 gnd.n3570 gnd.n3568 15.6674
R10043 gnd.n3538 gnd.n3536 15.6674
R10044 gnd.n3506 gnd.n3504 15.6674
R10045 gnd.n3474 gnd.n3472 15.6674
R10046 gnd.n3443 gnd.n3441 15.6674
R10047 gnd.n2969 gnd.t295 15.6146
R10048 gnd.t273 gnd.n2420 15.6146
R10049 gnd.t256 gnd.n2421 15.6146
R10050 gnd.n5026 gnd.n1848 15.296
R10051 gnd.n5612 gnd.n1840 15.296
R10052 gnd.t207 gnd.n1811 15.296
R10053 gnd.n5668 gnd.n1790 15.296
R10054 gnd.n5094 gnd.n1783 15.296
R10055 gnd.n5455 gnd.t2 15.296
R10056 gnd.n5426 gnd.n5425 15.296
R10057 gnd.n5748 gnd.n1720 15.296
R10058 gnd.n5189 gnd.n5188 15.0827
R10059 gnd.n4651 gnd.n4646 15.0481
R10060 gnd.n5199 gnd.n5198 15.0481
R10061 gnd.n3337 gnd.t56 14.9773
R10062 gnd.n4986 gnd.t122 14.9773
R10063 gnd.t286 gnd.t5 14.9773
R10064 gnd.n5796 gnd.t5 14.9773
R10065 gnd.t171 gnd.n1804 14.6587
R10066 gnd.n5463 gnd.t112 14.6587
R10067 gnd.t340 gnd.n2463 14.34
R10068 gnd.n3415 gnd.t42 14.34
R10069 gnd.n5556 gnd.n1855 14.0214
R10070 gnd.n5620 gnd.n1833 14.0214
R10071 gnd.t7 gnd.n1796 14.0214
R10072 gnd.n5660 gnd.n1798 14.0214
R10073 gnd.n5101 gnd.n1775 14.0214
R10074 gnd.n5470 gnd.t210 14.0214
R10075 gnd.n5135 gnd.n5133 14.0214
R10076 gnd.n5756 gnd.n1713 14.0214
R10077 gnd.n3125 gnd.t167 13.7027
R10078 gnd.n5066 gnd.t44 13.7027
R10079 gnd.n5700 gnd.t110 13.7027
R10080 gnd.n2835 gnd.n2834 13.5763
R10081 gnd.n3779 gnd.n2376 13.5763
R10082 gnd.n6086 gnd.n1332 13.5763
R10083 gnd.n7594 gnd.n7593 13.5763
R10084 gnd.n4124 gnd.n4039 13.5763
R10085 gnd.n4578 gnd.n4575 13.5763
R10086 gnd.n3043 gnd.n2781 13.384
R10087 gnd.t121 gnd.n1789 13.384
R10088 gnd.n5477 gnd.t29 13.384
R10089 gnd.n4662 gnd.n4643 13.1884
R10090 gnd.n4657 gnd.n4656 13.1884
R10091 gnd.n4656 gnd.n4655 13.1884
R10092 gnd.n5192 gnd.n5187 13.1884
R10093 gnd.n5193 gnd.n5192 13.1884
R10094 gnd.n4658 gnd.n4645 13.146
R10095 gnd.n4654 gnd.n4645 13.146
R10096 gnd.n5191 gnd.n5190 13.146
R10097 gnd.n5191 gnd.n5186 13.146
R10098 gnd.t93 gnd.n973 13.0654
R10099 gnd.t23 gnd.n356 13.0654
R10100 gnd.n3666 gnd.n3662 12.8005
R10101 gnd.n3634 gnd.n3630 12.8005
R10102 gnd.n3602 gnd.n3598 12.8005
R10103 gnd.n3571 gnd.n3567 12.8005
R10104 gnd.n3539 gnd.n3535 12.8005
R10105 gnd.n3507 gnd.n3503 12.8005
R10106 gnd.n3475 gnd.n3471 12.8005
R10107 gnd.n3444 gnd.n3440 12.8005
R10108 gnd.n1888 gnd.n1886 12.7467
R10109 gnd.n5652 gnd.n1805 12.7467
R10110 gnd.n5108 gnd.n1768 12.7467
R10111 gnd.n5764 gnd.n1706 12.7467
R10112 gnd.n2311 gnd.t162 12.4281
R10113 gnd.t95 gnd.n1018 12.4281
R10114 gnd.n4451 gnd.t128 12.4281
R10115 gnd.t153 gnd.n1949 12.4281
R10116 gnd.n1640 gnd.t216 12.4281
R10117 gnd.n5972 gnd.t145 12.4281
R10118 gnd.t80 gnd.n399 12.4281
R10119 gnd.t48 gnd.n229 12.4281
R10120 gnd.n2834 gnd.n2829 12.4126
R10121 gnd.n3782 gnd.n3779 12.4126
R10122 gnd.n6082 gnd.n1332 12.4126
R10123 gnd.n7593 gnd.n200 12.4126
R10124 gnd.n4120 gnd.n4039 12.4126
R10125 gnd.n4575 gnd.n2124 12.4126
R10126 gnd.n4744 gnd.n4743 12.1761
R10127 gnd.n5374 gnd.n5373 12.1761
R10128 gnd.n4847 gnd.n2047 12.1094
R10129 gnd.n6155 gnd.n1285 12.1094
R10130 gnd.n3670 gnd.n3669 12.0247
R10131 gnd.n3638 gnd.n3637 12.0247
R10132 gnd.n3606 gnd.n3605 12.0247
R10133 gnd.n3575 gnd.n3574 12.0247
R10134 gnd.n3543 gnd.n3542 12.0247
R10135 gnd.n3511 gnd.n3510 12.0247
R10136 gnd.n3479 gnd.n3478 12.0247
R10137 gnd.n3448 gnd.n3447 12.0247
R10138 gnd.n2279 gnd.t90 11.7908
R10139 gnd.n4398 gnd.t95 11.7908
R10140 gnd.t128 gnd.n1060 11.7908
R10141 gnd.t145 gnd.n5970 11.7908
R10142 gnd.n5999 gnd.t80 11.7908
R10143 gnd.t104 gnd.n260 11.7908
R10144 gnd.n5012 gnd.n1869 11.4721
R10145 gnd.n5636 gnd.n1819 11.4721
R10146 gnd.n5644 gnd.n1813 11.4721
R10147 gnd.n5457 gnd.n5456 11.4721
R10148 gnd.n5448 gnd.n5120 11.4721
R10149 gnd.n5772 gnd.n1699 11.4721
R10150 gnd.n5780 gnd.n1693 11.4721
R10151 gnd.n5378 gnd.t260 11.4721
R10152 gnd.n3673 gnd.n3660 11.249
R10153 gnd.n3641 gnd.n3628 11.249
R10154 gnd.n3609 gnd.n3596 11.249
R10155 gnd.n3578 gnd.n3565 11.249
R10156 gnd.n3546 gnd.n3533 11.249
R10157 gnd.n3514 gnd.n3501 11.249
R10158 gnd.n3482 gnd.n3469 11.249
R10159 gnd.n3451 gnd.n3438 11.249
R10160 gnd.n3113 gnd.t167 11.1535
R10161 gnd.n2247 gnd.t65 11.1535
R10162 gnd.n4364 gnd.t93 11.1535
R10163 gnd.n5525 gnd.t108 11.1535
R10164 gnd.t151 gnd.n5440 11.1535
R10165 gnd.n7269 gnd.t23 11.1535
R10166 gnd.t73 gnd.n290 11.1535
R10167 gnd.n5308 gnd.n5229 10.6151
R10168 gnd.n5308 gnd.n5307 10.6151
R10169 gnd.n5305 gnd.n5233 10.6151
R10170 gnd.n5300 gnd.n5233 10.6151
R10171 gnd.n5300 gnd.n5299 10.6151
R10172 gnd.n5299 gnd.n5298 10.6151
R10173 gnd.n5298 gnd.n5236 10.6151
R10174 gnd.n5293 gnd.n5236 10.6151
R10175 gnd.n5293 gnd.n5292 10.6151
R10176 gnd.n5292 gnd.n5291 10.6151
R10177 gnd.n5291 gnd.n5239 10.6151
R10178 gnd.n5286 gnd.n5239 10.6151
R10179 gnd.n5286 gnd.n5285 10.6151
R10180 gnd.n5285 gnd.n5284 10.6151
R10181 gnd.n5284 gnd.n5242 10.6151
R10182 gnd.n5279 gnd.n5242 10.6151
R10183 gnd.n5279 gnd.n5278 10.6151
R10184 gnd.n5278 gnd.n5277 10.6151
R10185 gnd.n5277 gnd.n5245 10.6151
R10186 gnd.n5272 gnd.n5245 10.6151
R10187 gnd.n5272 gnd.n5271 10.6151
R10188 gnd.n5271 gnd.n5270 10.6151
R10189 gnd.n5270 gnd.n5248 10.6151
R10190 gnd.n5265 gnd.n5248 10.6151
R10191 gnd.n5265 gnd.n5264 10.6151
R10192 gnd.n5264 gnd.n5263 10.6151
R10193 gnd.n5263 gnd.n5251 10.6151
R10194 gnd.n5258 gnd.n5251 10.6151
R10195 gnd.n5258 gnd.n5257 10.6151
R10196 gnd.n5257 gnd.n5256 10.6151
R10197 gnd.n4639 gnd.n4637 10.6151
R10198 gnd.n4639 gnd.n4638 10.6151
R10199 gnd.n4638 gnd.n1882 10.6151
R10200 gnd.n5570 gnd.n1882 10.6151
R10201 gnd.n5570 gnd.n5569 10.6151
R10202 gnd.n5569 gnd.n5568 10.6151
R10203 gnd.n5568 gnd.n1883 10.6151
R10204 gnd.n1885 gnd.n1883 10.6151
R10205 gnd.n5022 gnd.n1885 10.6151
R10206 gnd.n5023 gnd.n5022 10.6151
R10207 gnd.n5554 gnd.n5023 10.6151
R10208 gnd.n5554 gnd.n5553 10.6151
R10209 gnd.n5553 gnd.n5552 10.6151
R10210 gnd.n5552 gnd.n5024 10.6151
R10211 gnd.n5035 gnd.n5024 10.6151
R10212 gnd.n5036 gnd.n5035 10.6151
R10213 gnd.n5539 gnd.n5036 10.6151
R10214 gnd.n5539 gnd.n5538 10.6151
R10215 gnd.n5538 gnd.n5537 10.6151
R10216 gnd.n5537 gnd.n5037 10.6151
R10217 gnd.n5048 gnd.n5037 10.6151
R10218 gnd.n5050 gnd.n5048 10.6151
R10219 gnd.n5051 gnd.n5050 10.6151
R10220 gnd.n5523 gnd.n5051 10.6151
R10221 gnd.n5523 gnd.n5522 10.6151
R10222 gnd.n5522 gnd.n5521 10.6151
R10223 gnd.n5521 gnd.n5052 10.6151
R10224 gnd.n5063 gnd.n5052 10.6151
R10225 gnd.n5510 gnd.n5063 10.6151
R10226 gnd.n5510 gnd.n5509 10.6151
R10227 gnd.n5509 gnd.n5508 10.6151
R10228 gnd.n5508 gnd.n5064 10.6151
R10229 gnd.n5076 gnd.n5064 10.6151
R10230 gnd.n5077 gnd.n5076 10.6151
R10231 gnd.n5496 gnd.n5077 10.6151
R10232 gnd.n5496 gnd.n5495 10.6151
R10233 gnd.n5495 gnd.n5494 10.6151
R10234 gnd.n5494 gnd.n5078 10.6151
R10235 gnd.n5090 gnd.n5078 10.6151
R10236 gnd.n5091 gnd.n5090 10.6151
R10237 gnd.n5482 gnd.n5091 10.6151
R10238 gnd.n5482 gnd.n5481 10.6151
R10239 gnd.n5481 gnd.n5480 10.6151
R10240 gnd.n5480 gnd.n5092 10.6151
R10241 gnd.n5104 gnd.n5092 10.6151
R10242 gnd.n5105 gnd.n5104 10.6151
R10243 gnd.n5468 gnd.n5105 10.6151
R10244 gnd.n5468 gnd.n5467 10.6151
R10245 gnd.n5467 gnd.n5466 10.6151
R10246 gnd.n5466 gnd.n5106 10.6151
R10247 gnd.n5116 gnd.n5106 10.6151
R10248 gnd.n5117 gnd.n5116 10.6151
R10249 gnd.n5453 gnd.n5117 10.6151
R10250 gnd.n5453 gnd.n5452 10.6151
R10251 gnd.n5452 gnd.n5451 10.6151
R10252 gnd.n5451 gnd.n5118 10.6151
R10253 gnd.n5129 gnd.n5118 10.6151
R10254 gnd.n5130 gnd.n5129 10.6151
R10255 gnd.n5438 gnd.n5130 10.6151
R10256 gnd.n5438 gnd.n5437 10.6151
R10257 gnd.n5437 gnd.n5436 10.6151
R10258 gnd.n5436 gnd.n5131 10.6151
R10259 gnd.n5143 gnd.n5131 10.6151
R10260 gnd.n5144 gnd.n5143 10.6151
R10261 gnd.n5423 gnd.n5144 10.6151
R10262 gnd.n5423 gnd.n5422 10.6151
R10263 gnd.n5422 gnd.n5421 10.6151
R10264 gnd.n5421 gnd.n5145 10.6151
R10265 gnd.n5157 gnd.n5145 10.6151
R10266 gnd.n5409 gnd.n5157 10.6151
R10267 gnd.n5409 gnd.n5408 10.6151
R10268 gnd.n5408 gnd.n5407 10.6151
R10269 gnd.n5407 gnd.n5158 10.6151
R10270 gnd.n5171 gnd.n5158 10.6151
R10271 gnd.n5172 gnd.n5171 10.6151
R10272 gnd.n5394 gnd.n5172 10.6151
R10273 gnd.n5394 gnd.n5393 10.6151
R10274 gnd.n5393 gnd.n5392 10.6151
R10275 gnd.n5392 gnd.n5173 10.6151
R10276 gnd.n5382 gnd.n5173 10.6151
R10277 gnd.n5382 gnd.n5381 10.6151
R10278 gnd.n5381 gnd.n5380 10.6151
R10279 gnd.n5380 gnd.n5181 10.6151
R10280 gnd.n4811 gnd.n4617 10.6151
R10281 gnd.n4811 gnd.n4810 10.6151
R10282 gnd.n4808 gnd.n4623 10.6151
R10283 gnd.n4802 gnd.n4623 10.6151
R10284 gnd.n4802 gnd.n4801 10.6151
R10285 gnd.n4801 gnd.n4800 10.6151
R10286 gnd.n4800 gnd.n4625 10.6151
R10287 gnd.n4794 gnd.n4625 10.6151
R10288 gnd.n4794 gnd.n4793 10.6151
R10289 gnd.n4793 gnd.n4792 10.6151
R10290 gnd.n4792 gnd.n4627 10.6151
R10291 gnd.n4786 gnd.n4627 10.6151
R10292 gnd.n4786 gnd.n4785 10.6151
R10293 gnd.n4785 gnd.n4784 10.6151
R10294 gnd.n4784 gnd.n4629 10.6151
R10295 gnd.n4778 gnd.n4629 10.6151
R10296 gnd.n4778 gnd.n4777 10.6151
R10297 gnd.n4777 gnd.n4776 10.6151
R10298 gnd.n4776 gnd.n4631 10.6151
R10299 gnd.n4770 gnd.n4631 10.6151
R10300 gnd.n4770 gnd.n4769 10.6151
R10301 gnd.n4769 gnd.n4768 10.6151
R10302 gnd.n4768 gnd.n4633 10.6151
R10303 gnd.n4762 gnd.n4633 10.6151
R10304 gnd.n4762 gnd.n4761 10.6151
R10305 gnd.n4761 gnd.n4760 10.6151
R10306 gnd.n4760 gnd.n4635 10.6151
R10307 gnd.n4754 gnd.n4635 10.6151
R10308 gnd.n4754 gnd.n4753 10.6151
R10309 gnd.n4753 gnd.n4752 10.6151
R10310 gnd.n4743 gnd.n4742 10.6151
R10311 gnd.n4742 gnd.n4663 10.6151
R10312 gnd.n4737 gnd.n4663 10.6151
R10313 gnd.n4737 gnd.n4736 10.6151
R10314 gnd.n4736 gnd.n4665 10.6151
R10315 gnd.n4731 gnd.n4665 10.6151
R10316 gnd.n4731 gnd.n4730 10.6151
R10317 gnd.n4730 gnd.n4729 10.6151
R10318 gnd.n4729 gnd.n4667 10.6151
R10319 gnd.n4723 gnd.n4667 10.6151
R10320 gnd.n4723 gnd.n4722 10.6151
R10321 gnd.n4722 gnd.n4721 10.6151
R10322 gnd.n4721 gnd.n4669 10.6151
R10323 gnd.n4715 gnd.n4669 10.6151
R10324 gnd.n4715 gnd.n4714 10.6151
R10325 gnd.n4714 gnd.n4713 10.6151
R10326 gnd.n4713 gnd.n4671 10.6151
R10327 gnd.n4707 gnd.n4671 10.6151
R10328 gnd.n4707 gnd.n4706 10.6151
R10329 gnd.n4706 gnd.n4705 10.6151
R10330 gnd.n4705 gnd.n4673 10.6151
R10331 gnd.n4699 gnd.n4673 10.6151
R10332 gnd.n4699 gnd.n4698 10.6151
R10333 gnd.n4698 gnd.n4697 10.6151
R10334 gnd.n4697 gnd.n4675 10.6151
R10335 gnd.n4691 gnd.n4675 10.6151
R10336 gnd.n4691 gnd.n4690 10.6151
R10337 gnd.n4690 gnd.n4689 10.6151
R10338 gnd.n4685 gnd.n4684 10.6151
R10339 gnd.n4684 gnd.n4618 10.6151
R10340 gnd.n5373 gnd.n5204 10.6151
R10341 gnd.n5205 gnd.n5204 10.6151
R10342 gnd.n5366 gnd.n5205 10.6151
R10343 gnd.n5366 gnd.n5365 10.6151
R10344 gnd.n5365 gnd.n5364 10.6151
R10345 gnd.n5364 gnd.n5207 10.6151
R10346 gnd.n5359 gnd.n5207 10.6151
R10347 gnd.n5359 gnd.n5358 10.6151
R10348 gnd.n5358 gnd.n5357 10.6151
R10349 gnd.n5357 gnd.n5210 10.6151
R10350 gnd.n5352 gnd.n5210 10.6151
R10351 gnd.n5352 gnd.n5351 10.6151
R10352 gnd.n5351 gnd.n5350 10.6151
R10353 gnd.n5350 gnd.n5213 10.6151
R10354 gnd.n5345 gnd.n5213 10.6151
R10355 gnd.n5345 gnd.n5344 10.6151
R10356 gnd.n5344 gnd.n5343 10.6151
R10357 gnd.n5343 gnd.n5216 10.6151
R10358 gnd.n5338 gnd.n5216 10.6151
R10359 gnd.n5338 gnd.n5337 10.6151
R10360 gnd.n5337 gnd.n5336 10.6151
R10361 gnd.n5336 gnd.n5219 10.6151
R10362 gnd.n5331 gnd.n5219 10.6151
R10363 gnd.n5331 gnd.n5330 10.6151
R10364 gnd.n5330 gnd.n5329 10.6151
R10365 gnd.n5329 gnd.n5222 10.6151
R10366 gnd.n5324 gnd.n5222 10.6151
R10367 gnd.n5324 gnd.n5323 10.6151
R10368 gnd.n5321 gnd.n5227 10.6151
R10369 gnd.n5316 gnd.n5227 10.6151
R10370 gnd.n4746 gnd.n4745 10.6151
R10371 gnd.n4745 gnd.n1890 10.6151
R10372 gnd.n5009 gnd.n1890 10.6151
R10373 gnd.n5010 gnd.n5009 10.6151
R10374 gnd.n5011 gnd.n5010 10.6151
R10375 gnd.n5016 gnd.n5011 10.6151
R10376 gnd.n5017 gnd.n5016 10.6151
R10377 gnd.n5562 gnd.n5017 10.6151
R10378 gnd.n5562 gnd.n5561 10.6151
R10379 gnd.n5561 gnd.n5560 10.6151
R10380 gnd.n5560 gnd.n5018 10.6151
R10381 gnd.n5029 gnd.n5018 10.6151
R10382 gnd.n5030 gnd.n5029 10.6151
R10383 gnd.n5547 gnd.n5030 10.6151
R10384 gnd.n5547 gnd.n5546 10.6151
R10385 gnd.n5546 gnd.n5545 10.6151
R10386 gnd.n5545 gnd.n5031 10.6151
R10387 gnd.n5042 gnd.n5031 10.6151
R10388 gnd.n5043 gnd.n5042 10.6151
R10389 gnd.n5532 gnd.n5043 10.6151
R10390 gnd.n5532 gnd.n5531 10.6151
R10391 gnd.n5531 gnd.n5530 10.6151
R10392 gnd.n5530 gnd.n5044 10.6151
R10393 gnd.n5057 gnd.n5044 10.6151
R10394 gnd.n5058 gnd.n5057 10.6151
R10395 gnd.n5517 gnd.n5058 10.6151
R10396 gnd.n5517 gnd.n5516 10.6151
R10397 gnd.n5516 gnd.n5515 10.6151
R10398 gnd.n5515 gnd.n5059 10.6151
R10399 gnd.n5069 gnd.n5059 10.6151
R10400 gnd.n5070 gnd.n5069 10.6151
R10401 gnd.n5503 gnd.n5070 10.6151
R10402 gnd.n5503 gnd.n5502 10.6151
R10403 gnd.n5502 gnd.n5501 10.6151
R10404 gnd.n5501 gnd.n5071 10.6151
R10405 gnd.n5083 gnd.n5071 10.6151
R10406 gnd.n5084 gnd.n5083 10.6151
R10407 gnd.n5489 gnd.n5084 10.6151
R10408 gnd.n5489 gnd.n5488 10.6151
R10409 gnd.n5488 gnd.n5487 10.6151
R10410 gnd.n5487 gnd.n5085 10.6151
R10411 gnd.n5097 gnd.n5085 10.6151
R10412 gnd.n5098 gnd.n5097 10.6151
R10413 gnd.n5475 gnd.n5098 10.6151
R10414 gnd.n5475 gnd.n5474 10.6151
R10415 gnd.n5474 gnd.n5473 10.6151
R10416 gnd.n5473 gnd.n5099 10.6151
R10417 gnd.n5111 gnd.n5099 10.6151
R10418 gnd.n5112 gnd.n5111 10.6151
R10419 gnd.n5461 gnd.n5112 10.6151
R10420 gnd.n5461 gnd.n5460 10.6151
R10421 gnd.n5460 gnd.n5459 10.6151
R10422 gnd.n5459 gnd.n5113 10.6151
R10423 gnd.n5123 gnd.n5113 10.6151
R10424 gnd.n5124 gnd.n5123 10.6151
R10425 gnd.n5446 gnd.n5124 10.6151
R10426 gnd.n5446 gnd.n5445 10.6151
R10427 gnd.n5445 gnd.n5444 10.6151
R10428 gnd.n5444 gnd.n5125 10.6151
R10429 gnd.n5137 gnd.n5125 10.6151
R10430 gnd.n5432 gnd.n5137 10.6151
R10431 gnd.n5432 gnd.n5431 10.6151
R10432 gnd.n5431 gnd.n5430 10.6151
R10433 gnd.n5430 gnd.n5138 10.6151
R10434 gnd.n5151 gnd.n5138 10.6151
R10435 gnd.n5152 gnd.n5151 10.6151
R10436 gnd.n5417 gnd.n5152 10.6151
R10437 gnd.n5417 gnd.n5416 10.6151
R10438 gnd.n5416 gnd.n5415 10.6151
R10439 gnd.n5415 gnd.n5153 10.6151
R10440 gnd.n5164 gnd.n5153 10.6151
R10441 gnd.n5403 gnd.n5164 10.6151
R10442 gnd.n5403 gnd.n5402 10.6151
R10443 gnd.n5402 gnd.n5401 10.6151
R10444 gnd.n5401 gnd.n5165 10.6151
R10445 gnd.n5167 gnd.n5165 10.6151
R10446 gnd.n5176 gnd.n5167 10.6151
R10447 gnd.n5388 gnd.n5176 10.6151
R10448 gnd.n5388 gnd.n5387 10.6151
R10449 gnd.n5387 gnd.n5386 10.6151
R10450 gnd.n5386 gnd.n5177 10.6151
R10451 gnd.n5376 gnd.n5177 10.6151
R10452 gnd.n5376 gnd.n5375 10.6151
R10453 gnd.n3032 gnd.t3 10.5161
R10454 gnd.n2465 gnd.t340 10.5161
R10455 gnd.n3398 gnd.t42 10.5161
R10456 gnd.t19 gnd.n2214 10.5161
R10457 gnd.n2216 gnd.t36 10.5161
R10458 gnd.n5541 gnd.t186 10.5161
R10459 gnd.n5740 gnd.t358 10.5161
R10460 gnd.n7314 gnd.t86 10.5161
R10461 gnd.n7320 gnd.t71 10.5161
R10462 gnd.n3674 gnd.n3658 10.4732
R10463 gnd.n3642 gnd.n3626 10.4732
R10464 gnd.n3610 gnd.n3594 10.4732
R10465 gnd.n3579 gnd.n3563 10.4732
R10466 gnd.n3547 gnd.n3531 10.4732
R10467 gnd.n3515 gnd.n3499 10.4732
R10468 gnd.n3483 gnd.n3467 10.4732
R10469 gnd.n3452 gnd.n3436 10.4732
R10470 gnd.n5005 gnd.n1877 10.1975
R10471 gnd.n5013 gnd.n5012 10.1975
R10472 gnd.n1888 gnd.t227 10.1975
R10473 gnd.n5636 gnd.n1820 10.1975
R10474 gnd.n5644 gnd.n1811 10.1975
R10475 gnd.n5456 gnd.n5455 10.1975
R10476 gnd.n5120 gnd.n1753 10.1975
R10477 gnd.t260 gnd.n1684 10.1975
R10478 gnd.t56 gnd.n2482 9.87883
R10479 gnd.t97 gnd.n2244 9.87883
R10480 gnd.t328 gnd.t59 9.87883
R10481 gnd.n293 gnd.t183 9.87883
R10482 gnd.n7719 gnd.n78 9.81789
R10483 gnd.n3678 gnd.n3677 9.69747
R10484 gnd.n3646 gnd.n3645 9.69747
R10485 gnd.n3614 gnd.n3613 9.69747
R10486 gnd.n3583 gnd.n3582 9.69747
R10487 gnd.n3551 gnd.n3550 9.69747
R10488 gnd.n3519 gnd.n3518 9.69747
R10489 gnd.n3487 gnd.n3486 9.69747
R10490 gnd.n3456 gnd.n3455 9.69747
R10491 gnd.n6320 gnd.n1115 9.45751
R10492 gnd.n1517 gnd.n1342 9.45599
R10493 gnd.n3684 gnd.n3683 9.45567
R10494 gnd.n3652 gnd.n3651 9.45567
R10495 gnd.n3620 gnd.n3619 9.45567
R10496 gnd.n3589 gnd.n3588 9.45567
R10497 gnd.n3557 gnd.n3556 9.45567
R10498 gnd.n3525 gnd.n3524 9.45567
R10499 gnd.n3493 gnd.n3492 9.45567
R10500 gnd.n3462 gnd.n3461 9.45567
R10501 gnd.n2630 gnd.n2629 9.39724
R10502 gnd.n3683 gnd.n3682 9.3005
R10503 gnd.n3656 gnd.n3655 9.3005
R10504 gnd.n3677 gnd.n3676 9.3005
R10505 gnd.n3675 gnd.n3674 9.3005
R10506 gnd.n3660 gnd.n3659 9.3005
R10507 gnd.n3669 gnd.n3668 9.3005
R10508 gnd.n3667 gnd.n3666 9.3005
R10509 gnd.n3651 gnd.n3650 9.3005
R10510 gnd.n3624 gnd.n3623 9.3005
R10511 gnd.n3645 gnd.n3644 9.3005
R10512 gnd.n3643 gnd.n3642 9.3005
R10513 gnd.n3628 gnd.n3627 9.3005
R10514 gnd.n3637 gnd.n3636 9.3005
R10515 gnd.n3635 gnd.n3634 9.3005
R10516 gnd.n3619 gnd.n3618 9.3005
R10517 gnd.n3592 gnd.n3591 9.3005
R10518 gnd.n3613 gnd.n3612 9.3005
R10519 gnd.n3611 gnd.n3610 9.3005
R10520 gnd.n3596 gnd.n3595 9.3005
R10521 gnd.n3605 gnd.n3604 9.3005
R10522 gnd.n3603 gnd.n3602 9.3005
R10523 gnd.n3588 gnd.n3587 9.3005
R10524 gnd.n3561 gnd.n3560 9.3005
R10525 gnd.n3582 gnd.n3581 9.3005
R10526 gnd.n3580 gnd.n3579 9.3005
R10527 gnd.n3565 gnd.n3564 9.3005
R10528 gnd.n3574 gnd.n3573 9.3005
R10529 gnd.n3572 gnd.n3571 9.3005
R10530 gnd.n3556 gnd.n3555 9.3005
R10531 gnd.n3529 gnd.n3528 9.3005
R10532 gnd.n3550 gnd.n3549 9.3005
R10533 gnd.n3548 gnd.n3547 9.3005
R10534 gnd.n3533 gnd.n3532 9.3005
R10535 gnd.n3542 gnd.n3541 9.3005
R10536 gnd.n3540 gnd.n3539 9.3005
R10537 gnd.n3524 gnd.n3523 9.3005
R10538 gnd.n3497 gnd.n3496 9.3005
R10539 gnd.n3518 gnd.n3517 9.3005
R10540 gnd.n3516 gnd.n3515 9.3005
R10541 gnd.n3501 gnd.n3500 9.3005
R10542 gnd.n3510 gnd.n3509 9.3005
R10543 gnd.n3508 gnd.n3507 9.3005
R10544 gnd.n3492 gnd.n3491 9.3005
R10545 gnd.n3465 gnd.n3464 9.3005
R10546 gnd.n3486 gnd.n3485 9.3005
R10547 gnd.n3484 gnd.n3483 9.3005
R10548 gnd.n3469 gnd.n3468 9.3005
R10549 gnd.n3478 gnd.n3477 9.3005
R10550 gnd.n3476 gnd.n3475 9.3005
R10551 gnd.n3461 gnd.n3460 9.3005
R10552 gnd.n3434 gnd.n3433 9.3005
R10553 gnd.n3455 gnd.n3454 9.3005
R10554 gnd.n3453 gnd.n3452 9.3005
R10555 gnd.n3438 gnd.n3437 9.3005
R10556 gnd.n3447 gnd.n3446 9.3005
R10557 gnd.n3445 gnd.n3444 9.3005
R10558 gnd.n3809 gnd.n3808 9.3005
R10559 gnd.n3807 gnd.n2364 9.3005
R10560 gnd.n3806 gnd.n3805 9.3005
R10561 gnd.n3802 gnd.n2365 9.3005
R10562 gnd.n3799 gnd.n2366 9.3005
R10563 gnd.n3798 gnd.n2367 9.3005
R10564 gnd.n3795 gnd.n2368 9.3005
R10565 gnd.n3794 gnd.n2369 9.3005
R10566 gnd.n3791 gnd.n2370 9.3005
R10567 gnd.n3790 gnd.n2371 9.3005
R10568 gnd.n3787 gnd.n2372 9.3005
R10569 gnd.n3786 gnd.n2373 9.3005
R10570 gnd.n3783 gnd.n2374 9.3005
R10571 gnd.n3782 gnd.n2375 9.3005
R10572 gnd.n3779 gnd.n3778 9.3005
R10573 gnd.n3777 gnd.n2376 9.3005
R10574 gnd.n3810 gnd.n2363 9.3005
R10575 gnd.n3051 gnd.n3050 9.3005
R10576 gnd.n2755 gnd.n2754 9.3005
R10577 gnd.n3078 gnd.n3077 9.3005
R10578 gnd.n3079 gnd.n2753 9.3005
R10579 gnd.n3083 gnd.n3080 9.3005
R10580 gnd.n3082 gnd.n3081 9.3005
R10581 gnd.n2727 gnd.n2726 9.3005
R10582 gnd.n3108 gnd.n3107 9.3005
R10583 gnd.n3109 gnd.n2725 9.3005
R10584 gnd.n3111 gnd.n3110 9.3005
R10585 gnd.n2705 gnd.n2704 9.3005
R10586 gnd.n3139 gnd.n3138 9.3005
R10587 gnd.n3140 gnd.n2703 9.3005
R10588 gnd.n3148 gnd.n3141 9.3005
R10589 gnd.n3147 gnd.n3142 9.3005
R10590 gnd.n3146 gnd.n3144 9.3005
R10591 gnd.n3143 gnd.n2652 9.3005
R10592 gnd.n3196 gnd.n2653 9.3005
R10593 gnd.n3195 gnd.n2654 9.3005
R10594 gnd.n3194 gnd.n2655 9.3005
R10595 gnd.n2674 gnd.n2656 9.3005
R10596 gnd.n2676 gnd.n2675 9.3005
R10597 gnd.n2562 gnd.n2561 9.3005
R10598 gnd.n3234 gnd.n3233 9.3005
R10599 gnd.n3235 gnd.n2560 9.3005
R10600 gnd.n3239 gnd.n3236 9.3005
R10601 gnd.n3238 gnd.n3237 9.3005
R10602 gnd.n2535 gnd.n2534 9.3005
R10603 gnd.n3274 gnd.n3273 9.3005
R10604 gnd.n3275 gnd.n2533 9.3005
R10605 gnd.n3279 gnd.n3276 9.3005
R10606 gnd.n3278 gnd.n3277 9.3005
R10607 gnd.n2508 gnd.n2507 9.3005
R10608 gnd.n3319 gnd.n3318 9.3005
R10609 gnd.n3320 gnd.n2506 9.3005
R10610 gnd.n3324 gnd.n3321 9.3005
R10611 gnd.n3323 gnd.n3322 9.3005
R10612 gnd.n2480 gnd.n2479 9.3005
R10613 gnd.n3359 gnd.n3358 9.3005
R10614 gnd.n3360 gnd.n2478 9.3005
R10615 gnd.n3364 gnd.n3361 9.3005
R10616 gnd.n3363 gnd.n3362 9.3005
R10617 gnd.n2453 gnd.n2452 9.3005
R10618 gnd.n3408 gnd.n3407 9.3005
R10619 gnd.n3409 gnd.n2451 9.3005
R10620 gnd.n3413 gnd.n3410 9.3005
R10621 gnd.n3412 gnd.n3411 9.3005
R10622 gnd.n2426 gnd.n2425 9.3005
R10623 gnd.n3702 gnd.n3701 9.3005
R10624 gnd.n3703 gnd.n2424 9.3005
R10625 gnd.n3709 gnd.n3704 9.3005
R10626 gnd.n3708 gnd.n3705 9.3005
R10627 gnd.n3707 gnd.n3706 9.3005
R10628 gnd.n3052 gnd.n3049 9.3005
R10629 gnd.n2834 gnd.n2793 9.3005
R10630 gnd.n2829 gnd.n2828 9.3005
R10631 gnd.n2827 gnd.n2794 9.3005
R10632 gnd.n2826 gnd.n2825 9.3005
R10633 gnd.n2822 gnd.n2795 9.3005
R10634 gnd.n2819 gnd.n2818 9.3005
R10635 gnd.n2817 gnd.n2796 9.3005
R10636 gnd.n2816 gnd.n2815 9.3005
R10637 gnd.n2812 gnd.n2797 9.3005
R10638 gnd.n2809 gnd.n2808 9.3005
R10639 gnd.n2807 gnd.n2798 9.3005
R10640 gnd.n2806 gnd.n2805 9.3005
R10641 gnd.n2802 gnd.n2800 9.3005
R10642 gnd.n2799 gnd.n2779 9.3005
R10643 gnd.n3046 gnd.n2778 9.3005
R10644 gnd.n3048 gnd.n3047 9.3005
R10645 gnd.n2836 gnd.n2835 9.3005
R10646 gnd.n3059 gnd.n2765 9.3005
R10647 gnd.n3066 gnd.n2766 9.3005
R10648 gnd.n3068 gnd.n3067 9.3005
R10649 gnd.n3069 gnd.n2746 9.3005
R10650 gnd.n3088 gnd.n3087 9.3005
R10651 gnd.n3090 gnd.n2738 9.3005
R10652 gnd.n3097 gnd.n2740 9.3005
R10653 gnd.n3098 gnd.n2735 9.3005
R10654 gnd.n3100 gnd.n3099 9.3005
R10655 gnd.n2736 gnd.n2721 9.3005
R10656 gnd.n3116 gnd.n2719 9.3005
R10657 gnd.n3120 gnd.n3119 9.3005
R10658 gnd.n3118 gnd.n2695 9.3005
R10659 gnd.n3155 gnd.n2694 9.3005
R10660 gnd.n3158 gnd.n3157 9.3005
R10661 gnd.n2691 gnd.n2690 9.3005
R10662 gnd.n3164 gnd.n2692 9.3005
R10663 gnd.n3166 gnd.n3165 9.3005
R10664 gnd.n3168 gnd.n2689 9.3005
R10665 gnd.n3171 gnd.n3170 9.3005
R10666 gnd.n3174 gnd.n3172 9.3005
R10667 gnd.n3176 gnd.n3175 9.3005
R10668 gnd.n3182 gnd.n3177 9.3005
R10669 gnd.n3181 gnd.n3180 9.3005
R10670 gnd.n2553 gnd.n2552 9.3005
R10671 gnd.n3248 gnd.n3247 9.3005
R10672 gnd.n3249 gnd.n2546 9.3005
R10673 gnd.n3257 gnd.n2545 9.3005
R10674 gnd.n3260 gnd.n3259 9.3005
R10675 gnd.n3262 gnd.n3261 9.3005
R10676 gnd.n3265 gnd.n2528 9.3005
R10677 gnd.n3263 gnd.n2526 9.3005
R10678 gnd.n3285 gnd.n2524 9.3005
R10679 gnd.n3287 gnd.n3286 9.3005
R10680 gnd.n2498 gnd.n2497 9.3005
R10681 gnd.n3333 gnd.n3332 9.3005
R10682 gnd.n3334 gnd.n2491 9.3005
R10683 gnd.n3342 gnd.n2490 9.3005
R10684 gnd.n3345 gnd.n3344 9.3005
R10685 gnd.n3347 gnd.n3346 9.3005
R10686 gnd.n3350 gnd.n2473 9.3005
R10687 gnd.n3348 gnd.n2471 9.3005
R10688 gnd.n3370 gnd.n2469 9.3005
R10689 gnd.n3372 gnd.n3371 9.3005
R10690 gnd.n2444 gnd.n2443 9.3005
R10691 gnd.n3422 gnd.n3421 9.3005
R10692 gnd.n3423 gnd.n2437 9.3005
R10693 gnd.n3431 gnd.n2436 9.3005
R10694 gnd.n3690 gnd.n3689 9.3005
R10695 gnd.n3692 gnd.n3691 9.3005
R10696 gnd.n3693 gnd.n2417 9.3005
R10697 gnd.n3717 gnd.n3716 9.3005
R10698 gnd.n2418 gnd.n2379 9.3005
R10699 gnd.n3057 gnd.n3056 9.3005
R10700 gnd.n3773 gnd.n2380 9.3005
R10701 gnd.n3772 gnd.n2382 9.3005
R10702 gnd.n3769 gnd.n2383 9.3005
R10703 gnd.n3768 gnd.n2384 9.3005
R10704 gnd.n3765 gnd.n2385 9.3005
R10705 gnd.n3764 gnd.n2386 9.3005
R10706 gnd.n3761 gnd.n2387 9.3005
R10707 gnd.n3760 gnd.n2388 9.3005
R10708 gnd.n3757 gnd.n2389 9.3005
R10709 gnd.n3756 gnd.n2390 9.3005
R10710 gnd.n3753 gnd.n2391 9.3005
R10711 gnd.n3752 gnd.n2392 9.3005
R10712 gnd.n3749 gnd.n2393 9.3005
R10713 gnd.n3748 gnd.n2394 9.3005
R10714 gnd.n3745 gnd.n2395 9.3005
R10715 gnd.n3744 gnd.n2396 9.3005
R10716 gnd.n3741 gnd.n2397 9.3005
R10717 gnd.n3740 gnd.n2398 9.3005
R10718 gnd.n3737 gnd.n2399 9.3005
R10719 gnd.n3736 gnd.n2400 9.3005
R10720 gnd.n3733 gnd.n2401 9.3005
R10721 gnd.n3732 gnd.n2402 9.3005
R10722 gnd.n3729 gnd.n2406 9.3005
R10723 gnd.n3728 gnd.n2407 9.3005
R10724 gnd.n3725 gnd.n2408 9.3005
R10725 gnd.n3724 gnd.n2409 9.3005
R10726 gnd.n3775 gnd.n3774 9.3005
R10727 gnd.n3226 gnd.n3210 9.3005
R10728 gnd.n3225 gnd.n3211 9.3005
R10729 gnd.n3224 gnd.n3212 9.3005
R10730 gnd.n3222 gnd.n3213 9.3005
R10731 gnd.n3221 gnd.n3214 9.3005
R10732 gnd.n3219 gnd.n3215 9.3005
R10733 gnd.n3218 gnd.n3216 9.3005
R10734 gnd.n2516 gnd.n2515 9.3005
R10735 gnd.n3295 gnd.n3294 9.3005
R10736 gnd.n3296 gnd.n2514 9.3005
R10737 gnd.n3313 gnd.n3297 9.3005
R10738 gnd.n3312 gnd.n3298 9.3005
R10739 gnd.n3311 gnd.n3299 9.3005
R10740 gnd.n3309 gnd.n3300 9.3005
R10741 gnd.n3308 gnd.n3301 9.3005
R10742 gnd.n3306 gnd.n3302 9.3005
R10743 gnd.n3305 gnd.n3303 9.3005
R10744 gnd.n2460 gnd.n2459 9.3005
R10745 gnd.n3380 gnd.n3379 9.3005
R10746 gnd.n3381 gnd.n2458 9.3005
R10747 gnd.n3402 gnd.n3382 9.3005
R10748 gnd.n3401 gnd.n3383 9.3005
R10749 gnd.n3400 gnd.n3384 9.3005
R10750 gnd.n3397 gnd.n3385 9.3005
R10751 gnd.n3396 gnd.n3386 9.3005
R10752 gnd.n3394 gnd.n3387 9.3005
R10753 gnd.n3393 gnd.n3388 9.3005
R10754 gnd.n3391 gnd.n3390 9.3005
R10755 gnd.n3389 gnd.n2411 9.3005
R10756 gnd.n2967 gnd.n2966 9.3005
R10757 gnd.n2857 gnd.n2856 9.3005
R10758 gnd.n2981 gnd.n2980 9.3005
R10759 gnd.n2982 gnd.n2855 9.3005
R10760 gnd.n2984 gnd.n2983 9.3005
R10761 gnd.n2845 gnd.n2844 9.3005
R10762 gnd.n2997 gnd.n2996 9.3005
R10763 gnd.n2998 gnd.n2843 9.3005
R10764 gnd.n3030 gnd.n2999 9.3005
R10765 gnd.n3029 gnd.n3000 9.3005
R10766 gnd.n3028 gnd.n3001 9.3005
R10767 gnd.n3027 gnd.n3002 9.3005
R10768 gnd.n3024 gnd.n3003 9.3005
R10769 gnd.n3023 gnd.n3004 9.3005
R10770 gnd.n3022 gnd.n3005 9.3005
R10771 gnd.n3020 gnd.n3006 9.3005
R10772 gnd.n3019 gnd.n3007 9.3005
R10773 gnd.n3016 gnd.n3008 9.3005
R10774 gnd.n3015 gnd.n3009 9.3005
R10775 gnd.n3014 gnd.n3010 9.3005
R10776 gnd.n3012 gnd.n3011 9.3005
R10777 gnd.n2711 gnd.n2710 9.3005
R10778 gnd.n3128 gnd.n3127 9.3005
R10779 gnd.n3129 gnd.n2709 9.3005
R10780 gnd.n3133 gnd.n3130 9.3005
R10781 gnd.n3132 gnd.n3131 9.3005
R10782 gnd.n2633 gnd.n2632 9.3005
R10783 gnd.n3208 gnd.n3207 9.3005
R10784 gnd.n2965 gnd.n2866 9.3005
R10785 gnd.n2868 gnd.n2867 9.3005
R10786 gnd.n2912 gnd.n2910 9.3005
R10787 gnd.n2913 gnd.n2909 9.3005
R10788 gnd.n2916 gnd.n2905 9.3005
R10789 gnd.n2917 gnd.n2904 9.3005
R10790 gnd.n2920 gnd.n2903 9.3005
R10791 gnd.n2921 gnd.n2902 9.3005
R10792 gnd.n2924 gnd.n2901 9.3005
R10793 gnd.n2925 gnd.n2900 9.3005
R10794 gnd.n2928 gnd.n2899 9.3005
R10795 gnd.n2929 gnd.n2898 9.3005
R10796 gnd.n2932 gnd.n2897 9.3005
R10797 gnd.n2933 gnd.n2896 9.3005
R10798 gnd.n2936 gnd.n2895 9.3005
R10799 gnd.n2937 gnd.n2894 9.3005
R10800 gnd.n2940 gnd.n2893 9.3005
R10801 gnd.n2941 gnd.n2892 9.3005
R10802 gnd.n2944 gnd.n2891 9.3005
R10803 gnd.n2945 gnd.n2890 9.3005
R10804 gnd.n2948 gnd.n2889 9.3005
R10805 gnd.n2949 gnd.n2888 9.3005
R10806 gnd.n2952 gnd.n2887 9.3005
R10807 gnd.n2954 gnd.n2886 9.3005
R10808 gnd.n2955 gnd.n2885 9.3005
R10809 gnd.n2956 gnd.n2884 9.3005
R10810 gnd.n2957 gnd.n2883 9.3005
R10811 gnd.n2964 gnd.n2963 9.3005
R10812 gnd.n2973 gnd.n2972 9.3005
R10813 gnd.n2974 gnd.n2860 9.3005
R10814 gnd.n2976 gnd.n2975 9.3005
R10815 gnd.n2851 gnd.n2850 9.3005
R10816 gnd.n2989 gnd.n2988 9.3005
R10817 gnd.n2990 gnd.n2849 9.3005
R10818 gnd.n2992 gnd.n2991 9.3005
R10819 gnd.n2838 gnd.n2837 9.3005
R10820 gnd.n3035 gnd.n3034 9.3005
R10821 gnd.n3036 gnd.n2792 9.3005
R10822 gnd.n3040 gnd.n3038 9.3005
R10823 gnd.n3039 gnd.n2771 9.3005
R10824 gnd.n3058 gnd.n2770 9.3005
R10825 gnd.n3061 gnd.n3060 9.3005
R10826 gnd.n2764 gnd.n2763 9.3005
R10827 gnd.n3072 gnd.n3070 9.3005
R10828 gnd.n3071 gnd.n2745 9.3005
R10829 gnd.n3089 gnd.n2744 9.3005
R10830 gnd.n3092 gnd.n3091 9.3005
R10831 gnd.n2739 gnd.n2734 9.3005
R10832 gnd.n3102 gnd.n3101 9.3005
R10833 gnd.n2737 gnd.n2717 9.3005
R10834 gnd.n3123 gnd.n2718 9.3005
R10835 gnd.n3122 gnd.n3121 9.3005
R10836 gnd.n2720 gnd.n2696 9.3005
R10837 gnd.n3154 gnd.n3153 9.3005
R10838 gnd.n3156 gnd.n2641 9.3005
R10839 gnd.n3203 gnd.n2642 9.3005
R10840 gnd.n3202 gnd.n2643 9.3005
R10841 gnd.n3201 gnd.n2644 9.3005
R10842 gnd.n3167 gnd.n2645 9.3005
R10843 gnd.n3169 gnd.n2663 9.3005
R10844 gnd.n3189 gnd.n2664 9.3005
R10845 gnd.n3188 gnd.n2665 9.3005
R10846 gnd.n3187 gnd.n2666 9.3005
R10847 gnd.n3178 gnd.n2667 9.3005
R10848 gnd.n3179 gnd.n2554 9.3005
R10849 gnd.n3245 gnd.n3244 9.3005
R10850 gnd.n3246 gnd.n2547 9.3005
R10851 gnd.n3256 gnd.n3255 9.3005
R10852 gnd.n3258 gnd.n2543 9.3005
R10853 gnd.n3268 gnd.n2544 9.3005
R10854 gnd.n3267 gnd.n3266 9.3005
R10855 gnd.n3264 gnd.n2522 9.3005
R10856 gnd.n3290 gnd.n2523 9.3005
R10857 gnd.n3289 gnd.n3288 9.3005
R10858 gnd.n2525 gnd.n2499 9.3005
R10859 gnd.n3330 gnd.n3329 9.3005
R10860 gnd.n3331 gnd.n2492 9.3005
R10861 gnd.n3341 gnd.n3340 9.3005
R10862 gnd.n3343 gnd.n2488 9.3005
R10863 gnd.n3353 gnd.n2489 9.3005
R10864 gnd.n3352 gnd.n3351 9.3005
R10865 gnd.n3349 gnd.n2467 9.3005
R10866 gnd.n3375 gnd.n2468 9.3005
R10867 gnd.n3374 gnd.n3373 9.3005
R10868 gnd.n2470 gnd.n2445 9.3005
R10869 gnd.n3419 gnd.n3418 9.3005
R10870 gnd.n3420 gnd.n2438 9.3005
R10871 gnd.n3430 gnd.n3429 9.3005
R10872 gnd.n3688 gnd.n2434 9.3005
R10873 gnd.n3696 gnd.n2435 9.3005
R10874 gnd.n3695 gnd.n3694 9.3005
R10875 gnd.n2416 gnd.n2415 9.3005
R10876 gnd.n3719 gnd.n3718 9.3005
R10877 gnd.n2862 gnd.n2861 9.3005
R10878 gnd.n6580 gnd.n6579 9.3005
R10879 gnd.n795 gnd.n794 9.3005
R10880 gnd.n6587 gnd.n6586 9.3005
R10881 gnd.n6588 gnd.n793 9.3005
R10882 gnd.n6590 gnd.n6589 9.3005
R10883 gnd.n789 gnd.n788 9.3005
R10884 gnd.n6597 gnd.n6596 9.3005
R10885 gnd.n6598 gnd.n787 9.3005
R10886 gnd.n6600 gnd.n6599 9.3005
R10887 gnd.n783 gnd.n782 9.3005
R10888 gnd.n6607 gnd.n6606 9.3005
R10889 gnd.n6608 gnd.n781 9.3005
R10890 gnd.n6610 gnd.n6609 9.3005
R10891 gnd.n777 gnd.n776 9.3005
R10892 gnd.n6617 gnd.n6616 9.3005
R10893 gnd.n6618 gnd.n775 9.3005
R10894 gnd.n6620 gnd.n6619 9.3005
R10895 gnd.n771 gnd.n770 9.3005
R10896 gnd.n6627 gnd.n6626 9.3005
R10897 gnd.n6628 gnd.n769 9.3005
R10898 gnd.n6630 gnd.n6629 9.3005
R10899 gnd.n765 gnd.n764 9.3005
R10900 gnd.n6637 gnd.n6636 9.3005
R10901 gnd.n6638 gnd.n763 9.3005
R10902 gnd.n6640 gnd.n6639 9.3005
R10903 gnd.n759 gnd.n758 9.3005
R10904 gnd.n6647 gnd.n6646 9.3005
R10905 gnd.n6648 gnd.n757 9.3005
R10906 gnd.n6650 gnd.n6649 9.3005
R10907 gnd.n753 gnd.n752 9.3005
R10908 gnd.n6657 gnd.n6656 9.3005
R10909 gnd.n6658 gnd.n751 9.3005
R10910 gnd.n6660 gnd.n6659 9.3005
R10911 gnd.n747 gnd.n746 9.3005
R10912 gnd.n6667 gnd.n6666 9.3005
R10913 gnd.n6668 gnd.n745 9.3005
R10914 gnd.n6670 gnd.n6669 9.3005
R10915 gnd.n741 gnd.n740 9.3005
R10916 gnd.n6677 gnd.n6676 9.3005
R10917 gnd.n6678 gnd.n739 9.3005
R10918 gnd.n6680 gnd.n6679 9.3005
R10919 gnd.n735 gnd.n734 9.3005
R10920 gnd.n6687 gnd.n6686 9.3005
R10921 gnd.n6688 gnd.n733 9.3005
R10922 gnd.n6690 gnd.n6689 9.3005
R10923 gnd.n729 gnd.n728 9.3005
R10924 gnd.n6697 gnd.n6696 9.3005
R10925 gnd.n6698 gnd.n727 9.3005
R10926 gnd.n6700 gnd.n6699 9.3005
R10927 gnd.n723 gnd.n722 9.3005
R10928 gnd.n6707 gnd.n6706 9.3005
R10929 gnd.n6708 gnd.n721 9.3005
R10930 gnd.n6710 gnd.n6709 9.3005
R10931 gnd.n717 gnd.n716 9.3005
R10932 gnd.n6717 gnd.n6716 9.3005
R10933 gnd.n6718 gnd.n715 9.3005
R10934 gnd.n6720 gnd.n6719 9.3005
R10935 gnd.n711 gnd.n710 9.3005
R10936 gnd.n6727 gnd.n6726 9.3005
R10937 gnd.n6728 gnd.n709 9.3005
R10938 gnd.n6730 gnd.n6729 9.3005
R10939 gnd.n705 gnd.n704 9.3005
R10940 gnd.n6737 gnd.n6736 9.3005
R10941 gnd.n6738 gnd.n703 9.3005
R10942 gnd.n6740 gnd.n6739 9.3005
R10943 gnd.n699 gnd.n698 9.3005
R10944 gnd.n6747 gnd.n6746 9.3005
R10945 gnd.n6748 gnd.n697 9.3005
R10946 gnd.n6750 gnd.n6749 9.3005
R10947 gnd.n693 gnd.n692 9.3005
R10948 gnd.n6757 gnd.n6756 9.3005
R10949 gnd.n6758 gnd.n691 9.3005
R10950 gnd.n6760 gnd.n6759 9.3005
R10951 gnd.n687 gnd.n686 9.3005
R10952 gnd.n6767 gnd.n6766 9.3005
R10953 gnd.n6768 gnd.n685 9.3005
R10954 gnd.n6770 gnd.n6769 9.3005
R10955 gnd.n681 gnd.n680 9.3005
R10956 gnd.n6777 gnd.n6776 9.3005
R10957 gnd.n6778 gnd.n679 9.3005
R10958 gnd.n6780 gnd.n6779 9.3005
R10959 gnd.n675 gnd.n674 9.3005
R10960 gnd.n6787 gnd.n6786 9.3005
R10961 gnd.n6788 gnd.n673 9.3005
R10962 gnd.n6790 gnd.n6789 9.3005
R10963 gnd.n669 gnd.n668 9.3005
R10964 gnd.n6797 gnd.n6796 9.3005
R10965 gnd.n6798 gnd.n667 9.3005
R10966 gnd.n6800 gnd.n6799 9.3005
R10967 gnd.n663 gnd.n662 9.3005
R10968 gnd.n6807 gnd.n6806 9.3005
R10969 gnd.n6808 gnd.n661 9.3005
R10970 gnd.n6810 gnd.n6809 9.3005
R10971 gnd.n657 gnd.n656 9.3005
R10972 gnd.n6817 gnd.n6816 9.3005
R10973 gnd.n6818 gnd.n655 9.3005
R10974 gnd.n6820 gnd.n6819 9.3005
R10975 gnd.n651 gnd.n650 9.3005
R10976 gnd.n6827 gnd.n6826 9.3005
R10977 gnd.n6828 gnd.n649 9.3005
R10978 gnd.n6830 gnd.n6829 9.3005
R10979 gnd.n645 gnd.n644 9.3005
R10980 gnd.n6837 gnd.n6836 9.3005
R10981 gnd.n6838 gnd.n643 9.3005
R10982 gnd.n6840 gnd.n6839 9.3005
R10983 gnd.n639 gnd.n638 9.3005
R10984 gnd.n6847 gnd.n6846 9.3005
R10985 gnd.n6848 gnd.n637 9.3005
R10986 gnd.n6850 gnd.n6849 9.3005
R10987 gnd.n633 gnd.n632 9.3005
R10988 gnd.n6857 gnd.n6856 9.3005
R10989 gnd.n6858 gnd.n631 9.3005
R10990 gnd.n6860 gnd.n6859 9.3005
R10991 gnd.n627 gnd.n626 9.3005
R10992 gnd.n6867 gnd.n6866 9.3005
R10993 gnd.n6868 gnd.n625 9.3005
R10994 gnd.n6870 gnd.n6869 9.3005
R10995 gnd.n621 gnd.n620 9.3005
R10996 gnd.n6877 gnd.n6876 9.3005
R10997 gnd.n6878 gnd.n619 9.3005
R10998 gnd.n6880 gnd.n6879 9.3005
R10999 gnd.n615 gnd.n614 9.3005
R11000 gnd.n6887 gnd.n6886 9.3005
R11001 gnd.n6888 gnd.n613 9.3005
R11002 gnd.n6890 gnd.n6889 9.3005
R11003 gnd.n609 gnd.n608 9.3005
R11004 gnd.n6897 gnd.n6896 9.3005
R11005 gnd.n6898 gnd.n607 9.3005
R11006 gnd.n6900 gnd.n6899 9.3005
R11007 gnd.n603 gnd.n602 9.3005
R11008 gnd.n6907 gnd.n6906 9.3005
R11009 gnd.n6908 gnd.n601 9.3005
R11010 gnd.n6910 gnd.n6909 9.3005
R11011 gnd.n597 gnd.n596 9.3005
R11012 gnd.n6917 gnd.n6916 9.3005
R11013 gnd.n6918 gnd.n595 9.3005
R11014 gnd.n6920 gnd.n6919 9.3005
R11015 gnd.n591 gnd.n590 9.3005
R11016 gnd.n6927 gnd.n6926 9.3005
R11017 gnd.n6928 gnd.n589 9.3005
R11018 gnd.n6930 gnd.n6929 9.3005
R11019 gnd.n585 gnd.n584 9.3005
R11020 gnd.n6937 gnd.n6936 9.3005
R11021 gnd.n6938 gnd.n583 9.3005
R11022 gnd.n6940 gnd.n6939 9.3005
R11023 gnd.n579 gnd.n578 9.3005
R11024 gnd.n6947 gnd.n6946 9.3005
R11025 gnd.n6948 gnd.n577 9.3005
R11026 gnd.n6950 gnd.n6949 9.3005
R11027 gnd.n573 gnd.n572 9.3005
R11028 gnd.n6957 gnd.n6956 9.3005
R11029 gnd.n6958 gnd.n571 9.3005
R11030 gnd.n6960 gnd.n6959 9.3005
R11031 gnd.n567 gnd.n566 9.3005
R11032 gnd.n6967 gnd.n6966 9.3005
R11033 gnd.n6968 gnd.n565 9.3005
R11034 gnd.n6970 gnd.n6969 9.3005
R11035 gnd.n561 gnd.n560 9.3005
R11036 gnd.n6977 gnd.n6976 9.3005
R11037 gnd.n6978 gnd.n559 9.3005
R11038 gnd.n6980 gnd.n6979 9.3005
R11039 gnd.n555 gnd.n554 9.3005
R11040 gnd.n6987 gnd.n6986 9.3005
R11041 gnd.n6988 gnd.n553 9.3005
R11042 gnd.n6991 gnd.n6990 9.3005
R11043 gnd.n6989 gnd.n549 9.3005
R11044 gnd.n6997 gnd.n548 9.3005
R11045 gnd.n6999 gnd.n6998 9.3005
R11046 gnd.n544 gnd.n543 9.3005
R11047 gnd.n7008 gnd.n7007 9.3005
R11048 gnd.n7009 gnd.n542 9.3005
R11049 gnd.n7011 gnd.n7010 9.3005
R11050 gnd.n538 gnd.n537 9.3005
R11051 gnd.n7018 gnd.n7017 9.3005
R11052 gnd.n7019 gnd.n536 9.3005
R11053 gnd.n7021 gnd.n7020 9.3005
R11054 gnd.n532 gnd.n531 9.3005
R11055 gnd.n7028 gnd.n7027 9.3005
R11056 gnd.n7029 gnd.n530 9.3005
R11057 gnd.n7031 gnd.n7030 9.3005
R11058 gnd.n526 gnd.n525 9.3005
R11059 gnd.n7038 gnd.n7037 9.3005
R11060 gnd.n7039 gnd.n524 9.3005
R11061 gnd.n7041 gnd.n7040 9.3005
R11062 gnd.n520 gnd.n519 9.3005
R11063 gnd.n7048 gnd.n7047 9.3005
R11064 gnd.n7049 gnd.n518 9.3005
R11065 gnd.n7051 gnd.n7050 9.3005
R11066 gnd.n514 gnd.n513 9.3005
R11067 gnd.n7058 gnd.n7057 9.3005
R11068 gnd.n7059 gnd.n512 9.3005
R11069 gnd.n7061 gnd.n7060 9.3005
R11070 gnd.n508 gnd.n507 9.3005
R11071 gnd.n7068 gnd.n7067 9.3005
R11072 gnd.n7069 gnd.n506 9.3005
R11073 gnd.n7071 gnd.n7070 9.3005
R11074 gnd.n502 gnd.n501 9.3005
R11075 gnd.n7078 gnd.n7077 9.3005
R11076 gnd.n7079 gnd.n500 9.3005
R11077 gnd.n7081 gnd.n7080 9.3005
R11078 gnd.n496 gnd.n495 9.3005
R11079 gnd.n7088 gnd.n7087 9.3005
R11080 gnd.n7089 gnd.n494 9.3005
R11081 gnd.n7091 gnd.n7090 9.3005
R11082 gnd.n490 gnd.n489 9.3005
R11083 gnd.n7098 gnd.n7097 9.3005
R11084 gnd.n7099 gnd.n488 9.3005
R11085 gnd.n7101 gnd.n7100 9.3005
R11086 gnd.n484 gnd.n483 9.3005
R11087 gnd.n7108 gnd.n7107 9.3005
R11088 gnd.n7109 gnd.n482 9.3005
R11089 gnd.n7111 gnd.n7110 9.3005
R11090 gnd.n478 gnd.n477 9.3005
R11091 gnd.n7118 gnd.n7117 9.3005
R11092 gnd.n7119 gnd.n476 9.3005
R11093 gnd.n7121 gnd.n7120 9.3005
R11094 gnd.n472 gnd.n471 9.3005
R11095 gnd.n7128 gnd.n7127 9.3005
R11096 gnd.n7129 gnd.n470 9.3005
R11097 gnd.n7131 gnd.n7130 9.3005
R11098 gnd.n466 gnd.n465 9.3005
R11099 gnd.n7138 gnd.n7137 9.3005
R11100 gnd.n7139 gnd.n464 9.3005
R11101 gnd.n7141 gnd.n7140 9.3005
R11102 gnd.n460 gnd.n459 9.3005
R11103 gnd.n7148 gnd.n7147 9.3005
R11104 gnd.n7149 gnd.n458 9.3005
R11105 gnd.n7151 gnd.n7150 9.3005
R11106 gnd.n454 gnd.n453 9.3005
R11107 gnd.n7158 gnd.n7157 9.3005
R11108 gnd.n7159 gnd.n452 9.3005
R11109 gnd.n7161 gnd.n7160 9.3005
R11110 gnd.n448 gnd.n447 9.3005
R11111 gnd.n7168 gnd.n7167 9.3005
R11112 gnd.n7169 gnd.n446 9.3005
R11113 gnd.n7171 gnd.n7170 9.3005
R11114 gnd.n442 gnd.n441 9.3005
R11115 gnd.n7178 gnd.n7177 9.3005
R11116 gnd.n7179 gnd.n440 9.3005
R11117 gnd.n7181 gnd.n7180 9.3005
R11118 gnd.n436 gnd.n435 9.3005
R11119 gnd.n7188 gnd.n7187 9.3005
R11120 gnd.n7189 gnd.n434 9.3005
R11121 gnd.n7191 gnd.n7190 9.3005
R11122 gnd.n430 gnd.n429 9.3005
R11123 gnd.n7198 gnd.n7197 9.3005
R11124 gnd.n7199 gnd.n428 9.3005
R11125 gnd.n7201 gnd.n7200 9.3005
R11126 gnd.n424 gnd.n423 9.3005
R11127 gnd.n7209 gnd.n7208 9.3005
R11128 gnd.n7210 gnd.n422 9.3005
R11129 gnd.n7212 gnd.n7211 9.3005
R11130 gnd.n7001 gnd.n7000 9.3005
R11131 gnd.n7659 gnd.n134 9.3005
R11132 gnd.n7658 gnd.n136 9.3005
R11133 gnd.n140 gnd.n137 9.3005
R11134 gnd.n7653 gnd.n141 9.3005
R11135 gnd.n7652 gnd.n142 9.3005
R11136 gnd.n7651 gnd.n143 9.3005
R11137 gnd.n147 gnd.n144 9.3005
R11138 gnd.n7646 gnd.n148 9.3005
R11139 gnd.n7645 gnd.n149 9.3005
R11140 gnd.n7644 gnd.n150 9.3005
R11141 gnd.n154 gnd.n151 9.3005
R11142 gnd.n7639 gnd.n155 9.3005
R11143 gnd.n7638 gnd.n156 9.3005
R11144 gnd.n7637 gnd.n157 9.3005
R11145 gnd.n161 gnd.n158 9.3005
R11146 gnd.n7632 gnd.n162 9.3005
R11147 gnd.n7631 gnd.n163 9.3005
R11148 gnd.n7627 gnd.n164 9.3005
R11149 gnd.n168 gnd.n165 9.3005
R11150 gnd.n7622 gnd.n169 9.3005
R11151 gnd.n7621 gnd.n170 9.3005
R11152 gnd.n7620 gnd.n171 9.3005
R11153 gnd.n175 gnd.n172 9.3005
R11154 gnd.n7615 gnd.n176 9.3005
R11155 gnd.n7614 gnd.n177 9.3005
R11156 gnd.n7613 gnd.n178 9.3005
R11157 gnd.n182 gnd.n179 9.3005
R11158 gnd.n7608 gnd.n183 9.3005
R11159 gnd.n7607 gnd.n184 9.3005
R11160 gnd.n7606 gnd.n185 9.3005
R11161 gnd.n189 gnd.n186 9.3005
R11162 gnd.n7601 gnd.n190 9.3005
R11163 gnd.n7600 gnd.n191 9.3005
R11164 gnd.n7599 gnd.n192 9.3005
R11165 gnd.n196 gnd.n193 9.3005
R11166 gnd.n7594 gnd.n197 9.3005
R11167 gnd.n7593 gnd.n7592 9.3005
R11168 gnd.n7591 gnd.n200 9.3005
R11169 gnd.n7661 gnd.n7660 9.3005
R11170 gnd.n1456 gnd.n1455 9.3005
R11171 gnd.n1457 gnd.n1454 9.3005
R11172 gnd.n1473 gnd.n1458 9.3005
R11173 gnd.n1472 gnd.n1459 9.3005
R11174 gnd.n1471 gnd.n1460 9.3005
R11175 gnd.n1469 gnd.n1461 9.3005
R11176 gnd.n1468 gnd.n1462 9.3005
R11177 gnd.n1466 gnd.n1463 9.3005
R11178 gnd.n1465 gnd.n1464 9.3005
R11179 gnd.n1391 gnd.n1390 9.3005
R11180 gnd.n5985 gnd.n5984 9.3005
R11181 gnd.n5986 gnd.n1389 9.3005
R11182 gnd.n5988 gnd.n5987 9.3005
R11183 gnd.n5989 gnd.n1388 9.3005
R11184 gnd.n5992 gnd.n5991 9.3005
R11185 gnd.n5993 gnd.n1387 9.3005
R11186 gnd.n5997 gnd.n5994 9.3005
R11187 gnd.n5996 gnd.n5995 9.3005
R11188 gnd.n388 gnd.n387 9.3005
R11189 gnd.n7248 gnd.n7247 9.3005
R11190 gnd.n7249 gnd.n386 9.3005
R11191 gnd.n7257 gnd.n7250 9.3005
R11192 gnd.n7256 gnd.n7251 9.3005
R11193 gnd.n7255 gnd.n7252 9.3005
R11194 gnd.n354 gnd.n353 9.3005
R11195 gnd.n7293 gnd.n7292 9.3005
R11196 gnd.n7294 gnd.n352 9.3005
R11197 gnd.n7303 gnd.n7295 9.3005
R11198 gnd.n7302 gnd.n7296 9.3005
R11199 gnd.n7301 gnd.n7297 9.3005
R11200 gnd.n7299 gnd.n7298 9.3005
R11201 gnd.n338 gnd.n337 9.3005
R11202 gnd.n7323 gnd.n7322 9.3005
R11203 gnd.n7324 gnd.n336 9.3005
R11204 gnd.n7391 gnd.n7325 9.3005
R11205 gnd.n7390 gnd.n7326 9.3005
R11206 gnd.n7389 gnd.n7327 9.3005
R11207 gnd.n7387 gnd.n7328 9.3005
R11208 gnd.n7386 gnd.n7329 9.3005
R11209 gnd.n7384 gnd.n7330 9.3005
R11210 gnd.n7383 gnd.n7331 9.3005
R11211 gnd.n7381 gnd.n7332 9.3005
R11212 gnd.n7380 gnd.n7333 9.3005
R11213 gnd.n7378 gnd.n7334 9.3005
R11214 gnd.n7377 gnd.n7335 9.3005
R11215 gnd.n7375 gnd.n7336 9.3005
R11216 gnd.n7374 gnd.n7337 9.3005
R11217 gnd.n7372 gnd.n7338 9.3005
R11218 gnd.n7371 gnd.n7339 9.3005
R11219 gnd.n7369 gnd.n7340 9.3005
R11220 gnd.n7368 gnd.n7341 9.3005
R11221 gnd.n7366 gnd.n7342 9.3005
R11222 gnd.n7365 gnd.n7343 9.3005
R11223 gnd.n7363 gnd.n7344 9.3005
R11224 gnd.n7362 gnd.n7345 9.3005
R11225 gnd.n7360 gnd.n7346 9.3005
R11226 gnd.n7359 gnd.n7347 9.3005
R11227 gnd.n7357 gnd.n7348 9.3005
R11228 gnd.n7356 gnd.n7349 9.3005
R11229 gnd.n7354 gnd.n7350 9.3005
R11230 gnd.n7353 gnd.n7352 9.3005
R11231 gnd.n7351 gnd.n204 9.3005
R11232 gnd.n7588 gnd.n203 9.3005
R11233 gnd.n7590 gnd.n7589 9.3005
R11234 gnd.n1335 gnd.n1333 9.3005
R11235 gnd.n6086 gnd.n6085 9.3005
R11236 gnd.n6087 gnd.n1327 9.3005
R11237 gnd.n6090 gnd.n1326 9.3005
R11238 gnd.n6091 gnd.n1325 9.3005
R11239 gnd.n6094 gnd.n1324 9.3005
R11240 gnd.n6095 gnd.n1323 9.3005
R11241 gnd.n6098 gnd.n1322 9.3005
R11242 gnd.n6099 gnd.n1321 9.3005
R11243 gnd.n6102 gnd.n1320 9.3005
R11244 gnd.n6103 gnd.n1319 9.3005
R11245 gnd.n6106 gnd.n1318 9.3005
R11246 gnd.n6107 gnd.n1317 9.3005
R11247 gnd.n6110 gnd.n1316 9.3005
R11248 gnd.n6111 gnd.n1315 9.3005
R11249 gnd.n6114 gnd.n1314 9.3005
R11250 gnd.n6115 gnd.n1313 9.3005
R11251 gnd.n6118 gnd.n1312 9.3005
R11252 gnd.n6119 gnd.n1311 9.3005
R11253 gnd.n6122 gnd.n1310 9.3005
R11254 gnd.n6124 gnd.n1304 9.3005
R11255 gnd.n6127 gnd.n1303 9.3005
R11256 gnd.n6128 gnd.n1302 9.3005
R11257 gnd.n6131 gnd.n1301 9.3005
R11258 gnd.n6132 gnd.n1300 9.3005
R11259 gnd.n6135 gnd.n1299 9.3005
R11260 gnd.n6136 gnd.n1298 9.3005
R11261 gnd.n6139 gnd.n1297 9.3005
R11262 gnd.n6140 gnd.n1296 9.3005
R11263 gnd.n6143 gnd.n1295 9.3005
R11264 gnd.n6144 gnd.n1294 9.3005
R11265 gnd.n6147 gnd.n1293 9.3005
R11266 gnd.n6149 gnd.n1292 9.3005
R11267 gnd.n6150 gnd.n1291 9.3005
R11268 gnd.n6151 gnd.n1290 9.3005
R11269 gnd.n6152 gnd.n1289 9.3005
R11270 gnd.n6084 gnd.n1332 9.3005
R11271 gnd.n6083 gnd.n6082 9.3005
R11272 gnd.n5912 gnd.n5909 9.3005
R11273 gnd.n5911 gnd.n5910 9.3005
R11274 gnd.n1429 gnd.n1428 9.3005
R11275 gnd.n5938 gnd.n5937 9.3005
R11276 gnd.n5939 gnd.n1427 9.3005
R11277 gnd.n5943 gnd.n5940 9.3005
R11278 gnd.n5942 gnd.n5941 9.3005
R11279 gnd.n1402 gnd.n1401 9.3005
R11280 gnd.n5975 gnd.n5974 9.3005
R11281 gnd.n5976 gnd.n1400 9.3005
R11282 gnd.n5980 gnd.n5977 9.3005
R11283 gnd.n5979 gnd.n5978 9.3005
R11284 gnd.n1368 gnd.n1367 9.3005
R11285 gnd.n6045 gnd.n6044 9.3005
R11286 gnd.n6046 gnd.n1366 9.3005
R11287 gnd.n6048 gnd.n6047 9.3005
R11288 gnd.n397 gnd.n396 9.3005
R11289 gnd.n7238 gnd.n7237 9.3005
R11290 gnd.n7239 gnd.n395 9.3005
R11291 gnd.n7243 gnd.n7240 9.3005
R11292 gnd.n7242 gnd.n7241 9.3005
R11293 gnd.n364 gnd.n363 9.3005
R11294 gnd.n7284 gnd.n7283 9.3005
R11295 gnd.n7285 gnd.n362 9.3005
R11296 gnd.n7287 gnd.n7286 9.3005
R11297 gnd.n7288 gnd.n303 9.3005
R11298 gnd.n7419 gnd.n7418 9.3005
R11299 gnd.n288 gnd.n287 9.3005
R11300 gnd.n7432 gnd.n7431 9.3005
R11301 gnd.n7433 gnd.n286 9.3005
R11302 gnd.n7435 gnd.n7434 9.3005
R11303 gnd.n274 gnd.n273 9.3005
R11304 gnd.n7448 gnd.n7447 9.3005
R11305 gnd.n7449 gnd.n272 9.3005
R11306 gnd.n7451 gnd.n7450 9.3005
R11307 gnd.n258 gnd.n257 9.3005
R11308 gnd.n7464 gnd.n7463 9.3005
R11309 gnd.n7465 gnd.n256 9.3005
R11310 gnd.n7467 gnd.n7466 9.3005
R11311 gnd.n243 gnd.n242 9.3005
R11312 gnd.n7480 gnd.n7479 9.3005
R11313 gnd.n7481 gnd.n241 9.3005
R11314 gnd.n7483 gnd.n7482 9.3005
R11315 gnd.n227 gnd.n226 9.3005
R11316 gnd.n7496 gnd.n7495 9.3005
R11317 gnd.n7497 gnd.n225 9.3005
R11318 gnd.n7499 gnd.n7498 9.3005
R11319 gnd.n211 gnd.n210 9.3005
R11320 gnd.n7580 gnd.n7579 9.3005
R11321 gnd.n7581 gnd.n209 9.3005
R11322 gnd.n7583 gnd.n7582 9.3005
R11323 gnd.n133 gnd.n132 9.3005
R11324 gnd.n7663 gnd.n7662 9.3005
R11325 gnd.n5908 gnd.n5907 9.3005
R11326 gnd.n7417 gnd.n302 9.3005
R11327 gnd.n968 gnd.n967 9.3005
R11328 gnd.n4376 gnd.n4375 9.3005
R11329 gnd.n4377 gnd.n4373 9.3005
R11330 gnd.n4379 gnd.n4378 9.3005
R11331 gnd.n2170 gnd.n2169 9.3005
R11332 gnd.n4417 gnd.n4416 9.3005
R11333 gnd.n4418 gnd.n2168 9.3005
R11334 gnd.n4420 gnd.n4419 9.3005
R11335 gnd.n2166 gnd.n2165 9.3005
R11336 gnd.n4425 gnd.n4424 9.3005
R11337 gnd.n4426 gnd.n2164 9.3005
R11338 gnd.n4428 gnd.n4427 9.3005
R11339 gnd.n2149 gnd.n2148 9.3005
R11340 gnd.n4466 gnd.n4465 9.3005
R11341 gnd.n4467 gnd.n2147 9.3005
R11342 gnd.n4469 gnd.n4468 9.3005
R11343 gnd.n2145 gnd.n2144 9.3005
R11344 gnd.n4474 gnd.n4473 9.3005
R11345 gnd.n4475 gnd.n2143 9.3005
R11346 gnd.n4510 gnd.n4476 9.3005
R11347 gnd.n4509 gnd.n4477 9.3005
R11348 gnd.n4508 gnd.n4478 9.3005
R11349 gnd.n4481 gnd.n4479 9.3005
R11350 gnd.n4504 gnd.n4482 9.3005
R11351 gnd.n4503 gnd.n4483 9.3005
R11352 gnd.n4502 gnd.n4484 9.3005
R11353 gnd.n4487 gnd.n4485 9.3005
R11354 gnd.n4498 gnd.n4488 9.3005
R11355 gnd.n4497 gnd.n4489 9.3005
R11356 gnd.n4496 gnd.n4490 9.3005
R11357 gnd.n4492 gnd.n4491 9.3005
R11358 gnd.n1971 gnd.n1970 9.3005
R11359 gnd.n4909 gnd.n4908 9.3005
R11360 gnd.n4910 gnd.n1969 9.3005
R11361 gnd.n4912 gnd.n4911 9.3005
R11362 gnd.n1959 gnd.n1958 9.3005
R11363 gnd.n4925 gnd.n4924 9.3005
R11364 gnd.n4926 gnd.n1957 9.3005
R11365 gnd.n4928 gnd.n4927 9.3005
R11366 gnd.n1946 gnd.n1945 9.3005
R11367 gnd.n4941 gnd.n4940 9.3005
R11368 gnd.n4942 gnd.n1944 9.3005
R11369 gnd.n4944 gnd.n4943 9.3005
R11370 gnd.n1933 gnd.n1932 9.3005
R11371 gnd.n4957 gnd.n4956 9.3005
R11372 gnd.n4958 gnd.n1931 9.3005
R11373 gnd.n4960 gnd.n4959 9.3005
R11374 gnd.n1920 gnd.n1919 9.3005
R11375 gnd.n4973 gnd.n4972 9.3005
R11376 gnd.n4974 gnd.n1918 9.3005
R11377 gnd.n4976 gnd.n4975 9.3005
R11378 gnd.n1906 gnd.n1905 9.3005
R11379 gnd.n4989 gnd.n4988 9.3005
R11380 gnd.n4990 gnd.n1904 9.3005
R11381 gnd.n4994 gnd.n4991 9.3005
R11382 gnd.n4993 gnd.n4992 9.3005
R11383 gnd.n1875 gnd.n1874 9.3005
R11384 gnd.n5575 gnd.n5574 9.3005
R11385 gnd.n5576 gnd.n1873 9.3005
R11386 gnd.n5578 gnd.n5577 9.3005
R11387 gnd.n1861 gnd.n1860 9.3005
R11388 gnd.n5591 gnd.n5590 9.3005
R11389 gnd.n5592 gnd.n1859 9.3005
R11390 gnd.n5594 gnd.n5593 9.3005
R11391 gnd.n1846 gnd.n1845 9.3005
R11392 gnd.n5607 gnd.n5606 9.3005
R11393 gnd.n5608 gnd.n1844 9.3005
R11394 gnd.n5610 gnd.n5609 9.3005
R11395 gnd.n1831 gnd.n1830 9.3005
R11396 gnd.n5623 gnd.n5622 9.3005
R11397 gnd.n5624 gnd.n1829 9.3005
R11398 gnd.n5626 gnd.n5625 9.3005
R11399 gnd.n1817 gnd.n1816 9.3005
R11400 gnd.n5639 gnd.n5638 9.3005
R11401 gnd.n5640 gnd.n1815 9.3005
R11402 gnd.n5642 gnd.n5641 9.3005
R11403 gnd.n1802 gnd.n1801 9.3005
R11404 gnd.n5655 gnd.n5654 9.3005
R11405 gnd.n5656 gnd.n1800 9.3005
R11406 gnd.n5658 gnd.n5657 9.3005
R11407 gnd.n1787 gnd.n1786 9.3005
R11408 gnd.n5671 gnd.n5670 9.3005
R11409 gnd.n5672 gnd.n1785 9.3005
R11410 gnd.n5674 gnd.n5673 9.3005
R11411 gnd.n1772 gnd.n1771 9.3005
R11412 gnd.n5687 gnd.n5686 9.3005
R11413 gnd.n5688 gnd.n1770 9.3005
R11414 gnd.n5690 gnd.n5689 9.3005
R11415 gnd.n1758 gnd.n1757 9.3005
R11416 gnd.n5703 gnd.n5702 9.3005
R11417 gnd.n5704 gnd.n1756 9.3005
R11418 gnd.n5706 gnd.n5705 9.3005
R11419 gnd.n1743 gnd.n1742 9.3005
R11420 gnd.n5719 gnd.n5718 9.3005
R11421 gnd.n5720 gnd.n1741 9.3005
R11422 gnd.n5722 gnd.n5721 9.3005
R11423 gnd.n1730 gnd.n1729 9.3005
R11424 gnd.n5735 gnd.n5734 9.3005
R11425 gnd.n5736 gnd.n1728 9.3005
R11426 gnd.n5738 gnd.n5737 9.3005
R11427 gnd.n1718 gnd.n1717 9.3005
R11428 gnd.n5751 gnd.n5750 9.3005
R11429 gnd.n5752 gnd.n1716 9.3005
R11430 gnd.n5754 gnd.n5753 9.3005
R11431 gnd.n1704 gnd.n1703 9.3005
R11432 gnd.n5767 gnd.n5766 9.3005
R11433 gnd.n5768 gnd.n1702 9.3005
R11434 gnd.n5770 gnd.n5769 9.3005
R11435 gnd.n1691 gnd.n1690 9.3005
R11436 gnd.n5783 gnd.n5782 9.3005
R11437 gnd.n5784 gnd.n1689 9.3005
R11438 gnd.n5786 gnd.n5785 9.3005
R11439 gnd.n1677 gnd.n1676 9.3005
R11440 gnd.n5799 gnd.n5798 9.3005
R11441 gnd.n5800 gnd.n1675 9.3005
R11442 gnd.n5802 gnd.n5801 9.3005
R11443 gnd.n1664 gnd.n1663 9.3005
R11444 gnd.n5815 gnd.n5814 9.3005
R11445 gnd.n5816 gnd.n1662 9.3005
R11446 gnd.n5818 gnd.n5817 9.3005
R11447 gnd.n1651 gnd.n1650 9.3005
R11448 gnd.n5831 gnd.n5830 9.3005
R11449 gnd.n5832 gnd.n1649 9.3005
R11450 gnd.n5834 gnd.n5833 9.3005
R11451 gnd.n1637 gnd.n1636 9.3005
R11452 gnd.n5847 gnd.n5846 9.3005
R11453 gnd.n5848 gnd.n1635 9.3005
R11454 gnd.n5850 gnd.n5849 9.3005
R11455 gnd.n1624 gnd.n1623 9.3005
R11456 gnd.n5865 gnd.n5864 9.3005
R11457 gnd.n5866 gnd.n1622 9.3005
R11458 gnd.n5871 gnd.n5867 9.3005
R11459 gnd.n5870 gnd.n5869 9.3005
R11460 gnd.n5868 gnd.n1250 9.3005
R11461 gnd.n6161 gnd.n1251 9.3005
R11462 gnd.n6160 gnd.n1252 9.3005
R11463 gnd.n6159 gnd.n1253 9.3005
R11464 gnd.n1443 gnd.n1254 9.3005
R11465 gnd.n1446 gnd.n1445 9.3005
R11466 gnd.n1447 gnd.n1442 9.3005
R11467 gnd.n1449 gnd.n1448 9.3005
R11468 gnd.n1440 gnd.n1439 9.3005
R11469 gnd.n5927 gnd.n5926 9.3005
R11470 gnd.n5928 gnd.n1438 9.3005
R11471 gnd.n5932 gnd.n5929 9.3005
R11472 gnd.n5931 gnd.n5930 9.3005
R11473 gnd.n1412 gnd.n1411 9.3005
R11474 gnd.n5963 gnd.n5962 9.3005
R11475 gnd.n5964 gnd.n1410 9.3005
R11476 gnd.n5968 gnd.n5965 9.3005
R11477 gnd.n5967 gnd.n5966 9.3005
R11478 gnd.n1378 gnd.n1377 9.3005
R11479 gnd.n6024 gnd.n6023 9.3005
R11480 gnd.n6025 gnd.n1376 9.3005
R11481 gnd.n6039 gnd.n6026 9.3005
R11482 gnd.n6038 gnd.n6027 9.3005
R11483 gnd.n6037 gnd.n6028 9.3005
R11484 gnd.n6030 gnd.n6029 9.3005
R11485 gnd.n6033 gnd.n6032 9.3005
R11486 gnd.n6031 gnd.n411 9.3005
R11487 gnd.n7223 gnd.n412 9.3005
R11488 gnd.n7222 gnd.n413 9.3005
R11489 gnd.n7221 gnd.n414 9.3005
R11490 gnd.n417 gnd.n415 9.3005
R11491 gnd.n7217 gnd.n418 9.3005
R11492 gnd.n7216 gnd.n419 9.3005
R11493 gnd.n7215 gnd.n420 9.3005
R11494 gnd.n6406 gnd.n6405 9.3005
R11495 gnd.n3929 gnd.n3928 9.3005
R11496 gnd.n3975 gnd.n3884 9.3005
R11497 gnd.n3974 gnd.n3885 9.3005
R11498 gnd.n3973 gnd.n3886 9.3005
R11499 gnd.n3971 gnd.n3887 9.3005
R11500 gnd.n3970 gnd.n3888 9.3005
R11501 gnd.n3968 gnd.n3889 9.3005
R11502 gnd.n3967 gnd.n3890 9.3005
R11503 gnd.n3965 gnd.n3891 9.3005
R11504 gnd.n3964 gnd.n3892 9.3005
R11505 gnd.n3962 gnd.n3893 9.3005
R11506 gnd.n3961 gnd.n3894 9.3005
R11507 gnd.n3959 gnd.n3895 9.3005
R11508 gnd.n3958 gnd.n3896 9.3005
R11509 gnd.n3956 gnd.n3897 9.3005
R11510 gnd.n3955 gnd.n3898 9.3005
R11511 gnd.n3953 gnd.n3899 9.3005
R11512 gnd.n3952 gnd.n3900 9.3005
R11513 gnd.n3950 gnd.n3901 9.3005
R11514 gnd.n3949 gnd.n3902 9.3005
R11515 gnd.n3947 gnd.n3903 9.3005
R11516 gnd.n3946 gnd.n3904 9.3005
R11517 gnd.n3944 gnd.n3905 9.3005
R11518 gnd.n3943 gnd.n3906 9.3005
R11519 gnd.n3941 gnd.n3907 9.3005
R11520 gnd.n3940 gnd.n3908 9.3005
R11521 gnd.n3938 gnd.n3909 9.3005
R11522 gnd.n3937 gnd.n3910 9.3005
R11523 gnd.n3935 gnd.n3911 9.3005
R11524 gnd.n3934 gnd.n3912 9.3005
R11525 gnd.n3932 gnd.n3913 9.3005
R11526 gnd.n3931 gnd.n3914 9.3005
R11527 gnd.n3883 gnd.n3816 9.3005
R11528 gnd.n3876 gnd.n3875 9.3005
R11529 gnd.n3874 gnd.n3822 9.3005
R11530 gnd.n3873 gnd.n3872 9.3005
R11531 gnd.n3824 gnd.n3823 9.3005
R11532 gnd.n3866 gnd.n3865 9.3005
R11533 gnd.n3864 gnd.n3826 9.3005
R11534 gnd.n3863 gnd.n3862 9.3005
R11535 gnd.n3828 gnd.n3827 9.3005
R11536 gnd.n3856 gnd.n3855 9.3005
R11537 gnd.n3854 gnd.n3830 9.3005
R11538 gnd.n3853 gnd.n3852 9.3005
R11539 gnd.n3832 gnd.n3831 9.3005
R11540 gnd.n3846 gnd.n3845 9.3005
R11541 gnd.n3844 gnd.n3834 9.3005
R11542 gnd.n3843 gnd.n3842 9.3005
R11543 gnd.n3837 gnd.n3835 9.3005
R11544 gnd.n3836 gnd.n2337 9.3005
R11545 gnd.n3820 gnd.n3817 9.3005
R11546 gnd.n3882 gnd.n3881 9.3005
R11547 gnd.n4203 gnd.n2336 9.3005
R11548 gnd.n4205 gnd.n4204 9.3005
R11549 gnd.n2323 gnd.n2322 9.3005
R11550 gnd.n4218 gnd.n4217 9.3005
R11551 gnd.n4219 gnd.n2321 9.3005
R11552 gnd.n4221 gnd.n4220 9.3005
R11553 gnd.n2306 gnd.n2305 9.3005
R11554 gnd.n4234 gnd.n4233 9.3005
R11555 gnd.n4235 gnd.n2304 9.3005
R11556 gnd.n4237 gnd.n4236 9.3005
R11557 gnd.n2291 gnd.n2290 9.3005
R11558 gnd.n4250 gnd.n4249 9.3005
R11559 gnd.n4251 gnd.n2289 9.3005
R11560 gnd.n4253 gnd.n4252 9.3005
R11561 gnd.n2274 gnd.n2273 9.3005
R11562 gnd.n4266 gnd.n4265 9.3005
R11563 gnd.n4267 gnd.n2272 9.3005
R11564 gnd.n4269 gnd.n4268 9.3005
R11565 gnd.n2259 gnd.n2258 9.3005
R11566 gnd.n4282 gnd.n4281 9.3005
R11567 gnd.n4283 gnd.n2257 9.3005
R11568 gnd.n4285 gnd.n4284 9.3005
R11569 gnd.n2242 gnd.n2241 9.3005
R11570 gnd.n4299 gnd.n4298 9.3005
R11571 gnd.n4300 gnd.n2240 9.3005
R11572 gnd.n4302 gnd.n4301 9.3005
R11573 gnd.n2228 gnd.n2227 9.3005
R11574 gnd.n4315 gnd.n4314 9.3005
R11575 gnd.n4316 gnd.n2226 9.3005
R11576 gnd.n4319 gnd.n4317 9.3005
R11577 gnd.n4318 gnd.n2202 9.3005
R11578 gnd.n4333 gnd.n2203 9.3005
R11579 gnd.n4334 gnd.n2201 9.3005
R11580 gnd.n4346 gnd.n4335 9.3005
R11581 gnd.n4345 gnd.n4336 9.3005
R11582 gnd.n4344 gnd.n4337 9.3005
R11583 gnd.n4343 gnd.n4338 9.3005
R11584 gnd.n4341 gnd.n4340 9.3005
R11585 gnd.n4339 gnd.n989 9.3005
R11586 gnd.n6394 gnd.n990 9.3005
R11587 gnd.n6393 gnd.n991 9.3005
R11588 gnd.n6392 gnd.n992 9.3005
R11589 gnd.n1009 gnd.n993 9.3005
R11590 gnd.n6382 gnd.n1010 9.3005
R11591 gnd.n6381 gnd.n1011 9.3005
R11592 gnd.n6380 gnd.n1012 9.3005
R11593 gnd.n1031 gnd.n1013 9.3005
R11594 gnd.n6370 gnd.n1032 9.3005
R11595 gnd.n6369 gnd.n1033 9.3005
R11596 gnd.n6368 gnd.n1034 9.3005
R11597 gnd.n1051 gnd.n1035 9.3005
R11598 gnd.n6358 gnd.n1052 9.3005
R11599 gnd.n6357 gnd.n1053 9.3005
R11600 gnd.n6356 gnd.n1054 9.3005
R11601 gnd.n1073 gnd.n1055 9.3005
R11602 gnd.n6346 gnd.n1074 9.3005
R11603 gnd.n6345 gnd.n1075 9.3005
R11604 gnd.n6344 gnd.n1076 9.3005
R11605 gnd.n1094 gnd.n1077 9.3005
R11606 gnd.n6334 gnd.n1095 9.3005
R11607 gnd.n6333 gnd.n1096 9.3005
R11608 gnd.n6332 gnd.n1097 9.3005
R11609 gnd.n1114 gnd.n1098 9.3005
R11610 gnd.n6322 gnd.n6321 9.3005
R11611 gnd.n4202 gnd.n4201 9.3005
R11612 gnd.n4819 gnd.n2101 9.3005
R11613 gnd.n4822 gnd.n2100 9.3005
R11614 gnd.n4823 gnd.n2099 9.3005
R11615 gnd.n4826 gnd.n2098 9.3005
R11616 gnd.n4827 gnd.n2097 9.3005
R11617 gnd.n4830 gnd.n2096 9.3005
R11618 gnd.n4831 gnd.n2095 9.3005
R11619 gnd.n4834 gnd.n2094 9.3005
R11620 gnd.n4835 gnd.n2093 9.3005
R11621 gnd.n4838 gnd.n2092 9.3005
R11622 gnd.n4839 gnd.n2091 9.3005
R11623 gnd.n4842 gnd.n2090 9.3005
R11624 gnd.n4843 gnd.n2089 9.3005
R11625 gnd.n4844 gnd.n2088 9.3005
R11626 gnd.n2087 gnd.n2084 9.3005
R11627 gnd.n2086 gnd.n2085 9.3005
R11628 gnd.n4614 gnd.n4613 9.3005
R11629 gnd.n4610 gnd.n2106 9.3005
R11630 gnd.n4607 gnd.n2107 9.3005
R11631 gnd.n4606 gnd.n2108 9.3005
R11632 gnd.n4603 gnd.n2109 9.3005
R11633 gnd.n4602 gnd.n2110 9.3005
R11634 gnd.n4599 gnd.n2111 9.3005
R11635 gnd.n4598 gnd.n2112 9.3005
R11636 gnd.n4595 gnd.n2113 9.3005
R11637 gnd.n4594 gnd.n2114 9.3005
R11638 gnd.n4591 gnd.n2115 9.3005
R11639 gnd.n4590 gnd.n2116 9.3005
R11640 gnd.n4587 gnd.n2117 9.3005
R11641 gnd.n4586 gnd.n2118 9.3005
R11642 gnd.n4583 gnd.n2119 9.3005
R11643 gnd.n4582 gnd.n2120 9.3005
R11644 gnd.n4579 gnd.n2121 9.3005
R11645 gnd.n4578 gnd.n2122 9.3005
R11646 gnd.n4575 gnd.n4574 9.3005
R11647 gnd.n4573 gnd.n2124 9.3005
R11648 gnd.n4615 gnd.n2102 9.3005
R11649 gnd.n4114 gnd.n4040 9.3005
R11650 gnd.n4113 gnd.n4042 9.3005
R11651 gnd.n4112 gnd.n4043 9.3005
R11652 gnd.n4110 gnd.n4044 9.3005
R11653 gnd.n4109 gnd.n4045 9.3005
R11654 gnd.n4107 gnd.n4046 9.3005
R11655 gnd.n4106 gnd.n4047 9.3005
R11656 gnd.n4104 gnd.n4048 9.3005
R11657 gnd.n4103 gnd.n4049 9.3005
R11658 gnd.n4101 gnd.n4050 9.3005
R11659 gnd.n4100 gnd.n4051 9.3005
R11660 gnd.n4098 gnd.n4052 9.3005
R11661 gnd.n4097 gnd.n4053 9.3005
R11662 gnd.n4095 gnd.n4054 9.3005
R11663 gnd.n4094 gnd.n4055 9.3005
R11664 gnd.n4092 gnd.n4056 9.3005
R11665 gnd.n4091 gnd.n4057 9.3005
R11666 gnd.n4089 gnd.n4058 9.3005
R11667 gnd.n4088 gnd.n4059 9.3005
R11668 gnd.n4086 gnd.n4060 9.3005
R11669 gnd.n4085 gnd.n4061 9.3005
R11670 gnd.n4083 gnd.n4062 9.3005
R11671 gnd.n4082 gnd.n4063 9.3005
R11672 gnd.n4080 gnd.n4064 9.3005
R11673 gnd.n4079 gnd.n4065 9.3005
R11674 gnd.n4077 gnd.n4066 9.3005
R11675 gnd.n4076 gnd.n4067 9.3005
R11676 gnd.n4074 gnd.n4068 9.3005
R11677 gnd.n4073 gnd.n4069 9.3005
R11678 gnd.n4071 gnd.n4070 9.3005
R11679 gnd.n2206 gnd.n2204 9.3005
R11680 gnd.n4332 gnd.n4331 9.3005
R11681 gnd.n2211 gnd.n2205 9.3005
R11682 gnd.n2210 gnd.n2207 9.3005
R11683 gnd.n2209 gnd.n2208 9.3005
R11684 gnd.n2188 gnd.n2187 9.3005
R11685 gnd.n4359 gnd.n4358 9.3005
R11686 gnd.n4360 gnd.n2186 9.3005
R11687 gnd.n4362 gnd.n4361 9.3005
R11688 gnd.n2182 gnd.n2181 9.3005
R11689 gnd.n4385 gnd.n4384 9.3005
R11690 gnd.n4386 gnd.n2180 9.3005
R11691 gnd.n4388 gnd.n4387 9.3005
R11692 gnd.n4389 gnd.n2179 9.3005
R11693 gnd.n4393 gnd.n4392 9.3005
R11694 gnd.n4394 gnd.n2178 9.3005
R11695 gnd.n4396 gnd.n4395 9.3005
R11696 gnd.n2161 gnd.n2160 9.3005
R11697 gnd.n4434 gnd.n4433 9.3005
R11698 gnd.n4435 gnd.n2159 9.3005
R11699 gnd.n4437 gnd.n4436 9.3005
R11700 gnd.n4438 gnd.n2158 9.3005
R11701 gnd.n4442 gnd.n4441 9.3005
R11702 gnd.n4443 gnd.n2157 9.3005
R11703 gnd.n4449 gnd.n4444 9.3005
R11704 gnd.n4448 gnd.n4445 9.3005
R11705 gnd.n4447 gnd.n4446 9.3005
R11706 gnd.n2136 gnd.n2135 9.3005
R11707 gnd.n4524 gnd.n4523 9.3005
R11708 gnd.n4525 gnd.n2134 9.3005
R11709 gnd.n4528 gnd.n4527 9.3005
R11710 gnd.n4526 gnd.n2128 9.3005
R11711 gnd.n4570 gnd.n2127 9.3005
R11712 gnd.n4572 gnd.n4571 9.3005
R11713 gnd.n4116 gnd.n4115 9.3005
R11714 gnd.n4124 gnd.n4123 9.3005
R11715 gnd.n4125 gnd.n4034 9.3005
R11716 gnd.n4126 gnd.n4033 9.3005
R11717 gnd.n4032 gnd.n4030 9.3005
R11718 gnd.n4132 gnd.n4029 9.3005
R11719 gnd.n4133 gnd.n4028 9.3005
R11720 gnd.n4134 gnd.n4027 9.3005
R11721 gnd.n4026 gnd.n4024 9.3005
R11722 gnd.n4140 gnd.n4023 9.3005
R11723 gnd.n4141 gnd.n4022 9.3005
R11724 gnd.n4142 gnd.n4021 9.3005
R11725 gnd.n4020 gnd.n4018 9.3005
R11726 gnd.n4148 gnd.n4017 9.3005
R11727 gnd.n4149 gnd.n4016 9.3005
R11728 gnd.n4150 gnd.n4015 9.3005
R11729 gnd.n4014 gnd.n4012 9.3005
R11730 gnd.n4156 gnd.n4011 9.3005
R11731 gnd.n4157 gnd.n4010 9.3005
R11732 gnd.n4158 gnd.n4009 9.3005
R11733 gnd.n4008 gnd.n4003 9.3005
R11734 gnd.n4164 gnd.n4002 9.3005
R11735 gnd.n4165 gnd.n4001 9.3005
R11736 gnd.n4166 gnd.n4000 9.3005
R11737 gnd.n3999 gnd.n3997 9.3005
R11738 gnd.n4172 gnd.n3996 9.3005
R11739 gnd.n4173 gnd.n3995 9.3005
R11740 gnd.n4174 gnd.n3994 9.3005
R11741 gnd.n3993 gnd.n3991 9.3005
R11742 gnd.n4180 gnd.n3990 9.3005
R11743 gnd.n4181 gnd.n3989 9.3005
R11744 gnd.n4182 gnd.n3988 9.3005
R11745 gnd.n3987 gnd.n3985 9.3005
R11746 gnd.n4187 gnd.n3984 9.3005
R11747 gnd.n4188 gnd.n3983 9.3005
R11748 gnd.n3982 gnd.n3980 9.3005
R11749 gnd.n4193 gnd.n3979 9.3005
R11750 gnd.n4195 gnd.n4194 9.3005
R11751 gnd.n4122 gnd.n4039 9.3005
R11752 gnd.n4121 gnd.n4120 9.3005
R11753 gnd.n2331 gnd.n2330 9.3005
R11754 gnd.n4210 gnd.n4209 9.3005
R11755 gnd.n4211 gnd.n2329 9.3005
R11756 gnd.n4213 gnd.n4212 9.3005
R11757 gnd.n2315 gnd.n2314 9.3005
R11758 gnd.n4226 gnd.n4225 9.3005
R11759 gnd.n4227 gnd.n2313 9.3005
R11760 gnd.n4229 gnd.n4228 9.3005
R11761 gnd.n2299 gnd.n2298 9.3005
R11762 gnd.n4242 gnd.n4241 9.3005
R11763 gnd.n4243 gnd.n2297 9.3005
R11764 gnd.n4245 gnd.n4244 9.3005
R11765 gnd.n2283 gnd.n2282 9.3005
R11766 gnd.n4258 gnd.n4257 9.3005
R11767 gnd.n4259 gnd.n2281 9.3005
R11768 gnd.n4261 gnd.n4260 9.3005
R11769 gnd.n2267 gnd.n2266 9.3005
R11770 gnd.n4274 gnd.n4273 9.3005
R11771 gnd.n4275 gnd.n2265 9.3005
R11772 gnd.n4277 gnd.n4276 9.3005
R11773 gnd.n2251 gnd.n2250 9.3005
R11774 gnd.n4290 gnd.n4289 9.3005
R11775 gnd.n4291 gnd.n2249 9.3005
R11776 gnd.n4294 gnd.n4293 9.3005
R11777 gnd.n4292 gnd.n2234 9.3005
R11778 gnd.n4306 gnd.n2235 9.3005
R11779 gnd.n6400 gnd.n978 9.3005
R11780 gnd.n6399 gnd.n979 9.3005
R11781 gnd.n6398 gnd.n980 9.3005
R11782 gnd.n999 gnd.n981 9.3005
R11783 gnd.n6388 gnd.n1000 9.3005
R11784 gnd.n6387 gnd.n1001 9.3005
R11785 gnd.n6386 gnd.n1002 9.3005
R11786 gnd.n1020 gnd.n1003 9.3005
R11787 gnd.n6376 gnd.n1021 9.3005
R11788 gnd.n6375 gnd.n1022 9.3005
R11789 gnd.n6374 gnd.n1023 9.3005
R11790 gnd.n1041 gnd.n1024 9.3005
R11791 gnd.n6364 gnd.n1042 9.3005
R11792 gnd.n6363 gnd.n1043 9.3005
R11793 gnd.n6362 gnd.n1044 9.3005
R11794 gnd.n1062 gnd.n1045 9.3005
R11795 gnd.n6352 gnd.n1063 9.3005
R11796 gnd.n6351 gnd.n1064 9.3005
R11797 gnd.n6350 gnd.n1065 9.3005
R11798 gnd.n1083 gnd.n1066 9.3005
R11799 gnd.n6340 gnd.n1084 9.3005
R11800 gnd.n6339 gnd.n1085 9.3005
R11801 gnd.n6338 gnd.n1086 9.3005
R11802 gnd.n1104 gnd.n1087 9.3005
R11803 gnd.n6328 gnd.n1105 9.3005
R11804 gnd.n6327 gnd.n1106 9.3005
R11805 gnd.n6326 gnd.n1107 9.3005
R11806 gnd.n4197 gnd.n4196 9.3005
R11807 gnd.n977 gnd.n966 9.3005
R11808 gnd.n6410 gnd.n965 9.3005
R11809 gnd.n964 gnd.n960 9.3005
R11810 gnd.n6416 gnd.n959 9.3005
R11811 gnd.n6417 gnd.n958 9.3005
R11812 gnd.n6418 gnd.n957 9.3005
R11813 gnd.n956 gnd.n952 9.3005
R11814 gnd.n6424 gnd.n951 9.3005
R11815 gnd.n6425 gnd.n950 9.3005
R11816 gnd.n6426 gnd.n949 9.3005
R11817 gnd.n948 gnd.n944 9.3005
R11818 gnd.n6432 gnd.n943 9.3005
R11819 gnd.n6433 gnd.n942 9.3005
R11820 gnd.n6434 gnd.n941 9.3005
R11821 gnd.n940 gnd.n936 9.3005
R11822 gnd.n6440 gnd.n935 9.3005
R11823 gnd.n6441 gnd.n934 9.3005
R11824 gnd.n6442 gnd.n933 9.3005
R11825 gnd.n932 gnd.n928 9.3005
R11826 gnd.n6448 gnd.n927 9.3005
R11827 gnd.n6449 gnd.n926 9.3005
R11828 gnd.n6450 gnd.n925 9.3005
R11829 gnd.n924 gnd.n920 9.3005
R11830 gnd.n6456 gnd.n919 9.3005
R11831 gnd.n6457 gnd.n918 9.3005
R11832 gnd.n6458 gnd.n917 9.3005
R11833 gnd.n916 gnd.n912 9.3005
R11834 gnd.n6464 gnd.n911 9.3005
R11835 gnd.n6465 gnd.n910 9.3005
R11836 gnd.n6466 gnd.n909 9.3005
R11837 gnd.n908 gnd.n904 9.3005
R11838 gnd.n6472 gnd.n903 9.3005
R11839 gnd.n6473 gnd.n902 9.3005
R11840 gnd.n6474 gnd.n901 9.3005
R11841 gnd.n900 gnd.n896 9.3005
R11842 gnd.n6480 gnd.n895 9.3005
R11843 gnd.n6481 gnd.n894 9.3005
R11844 gnd.n6482 gnd.n893 9.3005
R11845 gnd.n892 gnd.n888 9.3005
R11846 gnd.n6488 gnd.n887 9.3005
R11847 gnd.n6489 gnd.n886 9.3005
R11848 gnd.n6490 gnd.n885 9.3005
R11849 gnd.n884 gnd.n880 9.3005
R11850 gnd.n6496 gnd.n879 9.3005
R11851 gnd.n6497 gnd.n878 9.3005
R11852 gnd.n6498 gnd.n877 9.3005
R11853 gnd.n876 gnd.n872 9.3005
R11854 gnd.n6504 gnd.n871 9.3005
R11855 gnd.n6505 gnd.n870 9.3005
R11856 gnd.n6506 gnd.n869 9.3005
R11857 gnd.n868 gnd.n864 9.3005
R11858 gnd.n6512 gnd.n863 9.3005
R11859 gnd.n6513 gnd.n862 9.3005
R11860 gnd.n6514 gnd.n861 9.3005
R11861 gnd.n860 gnd.n856 9.3005
R11862 gnd.n6520 gnd.n855 9.3005
R11863 gnd.n6521 gnd.n854 9.3005
R11864 gnd.n6522 gnd.n853 9.3005
R11865 gnd.n852 gnd.n848 9.3005
R11866 gnd.n6528 gnd.n847 9.3005
R11867 gnd.n6529 gnd.n846 9.3005
R11868 gnd.n6530 gnd.n845 9.3005
R11869 gnd.n844 gnd.n840 9.3005
R11870 gnd.n6536 gnd.n839 9.3005
R11871 gnd.n6537 gnd.n838 9.3005
R11872 gnd.n6538 gnd.n837 9.3005
R11873 gnd.n836 gnd.n832 9.3005
R11874 gnd.n6544 gnd.n831 9.3005
R11875 gnd.n6545 gnd.n830 9.3005
R11876 gnd.n6546 gnd.n829 9.3005
R11877 gnd.n828 gnd.n824 9.3005
R11878 gnd.n6552 gnd.n823 9.3005
R11879 gnd.n6553 gnd.n822 9.3005
R11880 gnd.n6554 gnd.n821 9.3005
R11881 gnd.n820 gnd.n816 9.3005
R11882 gnd.n6560 gnd.n815 9.3005
R11883 gnd.n6561 gnd.n814 9.3005
R11884 gnd.n6562 gnd.n813 9.3005
R11885 gnd.n812 gnd.n808 9.3005
R11886 gnd.n6568 gnd.n807 9.3005
R11887 gnd.n6569 gnd.n806 9.3005
R11888 gnd.n6570 gnd.n805 9.3005
R11889 gnd.n804 gnd.n800 9.3005
R11890 gnd.n6576 gnd.n799 9.3005
R11891 gnd.n6578 gnd.n6577 9.3005
R11892 gnd.n6409 gnd.n6408 9.3005
R11893 gnd.n1530 gnd.n1529 9.3005
R11894 gnd.n1516 gnd.n1512 9.3005
R11895 gnd.n1537 gnd.n1536 9.3005
R11896 gnd.n1538 gnd.n1507 9.3005
R11897 gnd.n1549 gnd.n1548 9.3005
R11898 gnd.n1509 gnd.n1505 9.3005
R11899 gnd.n1556 gnd.n1555 9.3005
R11900 gnd.n1557 gnd.n1500 9.3005
R11901 gnd.n1568 gnd.n1567 9.3005
R11902 gnd.n1502 gnd.n1498 9.3005
R11903 gnd.n1575 gnd.n1574 9.3005
R11904 gnd.n1495 gnd.n1494 9.3005
R11905 gnd.n1584 gnd.n1583 9.3005
R11906 gnd.n1492 gnd.n1491 9.3005
R11907 gnd.n1591 gnd.n1590 9.3005
R11908 gnd.n1483 gnd.n1482 9.3005
R11909 gnd.n1598 gnd.n1597 9.3005
R11910 gnd.n1480 gnd.n1478 9.3005
R11911 gnd.n1519 gnd.n1514 9.3005
R11912 gnd.n1593 gnd.n1592 9.3005
R11913 gnd.n1582 gnd.n1488 9.3005
R11914 gnd.n1581 gnd.n1580 9.3005
R11915 gnd.n1577 gnd.n1576 9.3005
R11916 gnd.n1497 gnd.n1496 9.3005
R11917 gnd.n1566 gnd.n1565 9.3005
R11918 gnd.n1562 gnd.n1501 9.3005
R11919 gnd.n1559 gnd.n1558 9.3005
R11920 gnd.n1504 gnd.n1503 9.3005
R11921 gnd.n1547 gnd.n1546 9.3005
R11922 gnd.n1543 gnd.n1508 9.3005
R11923 gnd.n1540 gnd.n1539 9.3005
R11924 gnd.n1511 gnd.n1510 9.3005
R11925 gnd.n1528 gnd.n1527 9.3005
R11926 gnd.n1524 gnd.n1515 9.3005
R11927 gnd.n1521 gnd.n1520 9.3005
R11928 gnd.n1594 gnd.n1484 9.3005
R11929 gnd.n1596 gnd.n1595 9.3005
R11930 gnd.n5901 gnd.n5900 9.3005
R11931 gnd.n5899 gnd.n1479 9.3005
R11932 gnd.n5898 gnd.n5897 9.3005
R11933 gnd.n5896 gnd.n1606 9.3005
R11934 gnd.n5895 gnd.n5894 9.3005
R11935 gnd.n5893 gnd.n1607 9.3005
R11936 gnd.n5889 gnd.n5888 9.3005
R11937 gnd.n5887 gnd.n1614 9.3005
R11938 gnd.n5886 gnd.n5885 9.3005
R11939 gnd.n5884 gnd.n5879 9.3005
R11940 gnd.n1966 gnd.n1965 9.3005
R11941 gnd.n4917 gnd.n4916 9.3005
R11942 gnd.n4918 gnd.n1964 9.3005
R11943 gnd.n4920 gnd.n4919 9.3005
R11944 gnd.n1953 gnd.n1952 9.3005
R11945 gnd.n4933 gnd.n4932 9.3005
R11946 gnd.n4934 gnd.n1951 9.3005
R11947 gnd.n4936 gnd.n4935 9.3005
R11948 gnd.n1938 gnd.n1937 9.3005
R11949 gnd.n4949 gnd.n4948 9.3005
R11950 gnd.n4950 gnd.n1936 9.3005
R11951 gnd.n4952 gnd.n4951 9.3005
R11952 gnd.n1925 gnd.n1924 9.3005
R11953 gnd.n4965 gnd.n4964 9.3005
R11954 gnd.n4966 gnd.n1923 9.3005
R11955 gnd.n4968 gnd.n4967 9.3005
R11956 gnd.n1914 gnd.n1913 9.3005
R11957 gnd.n4981 gnd.n4980 9.3005
R11958 gnd.n4982 gnd.n1912 9.3005
R11959 gnd.n4984 gnd.n4983 9.3005
R11960 gnd.n1899 gnd.n1898 9.3005
R11961 gnd.n4999 gnd.n4998 9.3005
R11962 gnd.n5000 gnd.n1896 9.3005
R11963 gnd.n5003 gnd.n5002 9.3005
R11964 gnd.n5001 gnd.n1897 9.3005
R11965 gnd.n1867 gnd.n1866 9.3005
R11966 gnd.n5583 gnd.n5582 9.3005
R11967 gnd.n5584 gnd.n1865 9.3005
R11968 gnd.n5586 gnd.n5585 9.3005
R11969 gnd.n1853 gnd.n1852 9.3005
R11970 gnd.n5599 gnd.n5598 9.3005
R11971 gnd.n5600 gnd.n1851 9.3005
R11972 gnd.n5602 gnd.n5601 9.3005
R11973 gnd.n1838 gnd.n1837 9.3005
R11974 gnd.n5615 gnd.n5614 9.3005
R11975 gnd.n5616 gnd.n1836 9.3005
R11976 gnd.n5618 gnd.n5617 9.3005
R11977 gnd.n1824 gnd.n1823 9.3005
R11978 gnd.n5631 gnd.n5630 9.3005
R11979 gnd.n5632 gnd.n1822 9.3005
R11980 gnd.n5634 gnd.n5633 9.3005
R11981 gnd.n1809 gnd.n1808 9.3005
R11982 gnd.n5647 gnd.n5646 9.3005
R11983 gnd.n5648 gnd.n1807 9.3005
R11984 gnd.n5650 gnd.n5649 9.3005
R11985 gnd.n1794 gnd.n1793 9.3005
R11986 gnd.n5663 gnd.n5662 9.3005
R11987 gnd.n5664 gnd.n1792 9.3005
R11988 gnd.n5666 gnd.n5665 9.3005
R11989 gnd.n1779 gnd.n1778 9.3005
R11990 gnd.n5679 gnd.n5678 9.3005
R11991 gnd.n5680 gnd.n1777 9.3005
R11992 gnd.n5682 gnd.n5681 9.3005
R11993 gnd.n1764 gnd.n1763 9.3005
R11994 gnd.n5695 gnd.n5694 9.3005
R11995 gnd.n5696 gnd.n1762 9.3005
R11996 gnd.n5698 gnd.n5697 9.3005
R11997 gnd.n1749 gnd.n1748 9.3005
R11998 gnd.n5711 gnd.n5710 9.3005
R11999 gnd.n5712 gnd.n1747 9.3005
R12000 gnd.n5714 gnd.n5713 9.3005
R12001 gnd.n1736 gnd.n1735 9.3005
R12002 gnd.n5727 gnd.n5726 9.3005
R12003 gnd.n5728 gnd.n1734 9.3005
R12004 gnd.n5730 gnd.n5729 9.3005
R12005 gnd.n1724 gnd.n1723 9.3005
R12006 gnd.n5743 gnd.n5742 9.3005
R12007 gnd.n5744 gnd.n1722 9.3005
R12008 gnd.n5746 gnd.n5745 9.3005
R12009 gnd.n1711 gnd.n1710 9.3005
R12010 gnd.n5759 gnd.n5758 9.3005
R12011 gnd.n5760 gnd.n1709 9.3005
R12012 gnd.n5762 gnd.n5761 9.3005
R12013 gnd.n1697 gnd.n1696 9.3005
R12014 gnd.n5775 gnd.n5774 9.3005
R12015 gnd.n5776 gnd.n1695 9.3005
R12016 gnd.n5778 gnd.n5777 9.3005
R12017 gnd.n1682 gnd.n1681 9.3005
R12018 gnd.n5791 gnd.n5790 9.3005
R12019 gnd.n5792 gnd.n1680 9.3005
R12020 gnd.n5794 gnd.n5793 9.3005
R12021 gnd.n1670 gnd.n1669 9.3005
R12022 gnd.n5807 gnd.n5806 9.3005
R12023 gnd.n5808 gnd.n1668 9.3005
R12024 gnd.n5810 gnd.n5809 9.3005
R12025 gnd.n1657 gnd.n1656 9.3005
R12026 gnd.n5823 gnd.n5822 9.3005
R12027 gnd.n5824 gnd.n1655 9.3005
R12028 gnd.n5826 gnd.n5825 9.3005
R12029 gnd.n1644 gnd.n1643 9.3005
R12030 gnd.n5839 gnd.n5838 9.3005
R12031 gnd.n5840 gnd.n1642 9.3005
R12032 gnd.n5842 gnd.n5841 9.3005
R12033 gnd.n1631 gnd.n1630 9.3005
R12034 gnd.n5855 gnd.n5854 9.3005
R12035 gnd.n5856 gnd.n1628 9.3005
R12036 gnd.n5860 gnd.n5859 9.3005
R12037 gnd.n5858 gnd.n1629 9.3005
R12038 gnd.n5857 gnd.n1616 9.3005
R12039 gnd.n5876 gnd.n1615 9.3005
R12040 gnd.n5878 gnd.n5877 9.3005
R12041 gnd.n4904 gnd.n4903 9.3005
R12042 gnd.n4900 gnd.n1976 9.3005
R12043 gnd.n4548 gnd.n1977 9.3005
R12044 gnd.n4551 gnd.n4550 9.3005
R12045 gnd.n4553 gnd.n4552 9.3005
R12046 gnd.n4554 gnd.n4541 9.3005
R12047 gnd.n4556 gnd.n4555 9.3005
R12048 gnd.n4557 gnd.n4540 9.3005
R12049 gnd.n4559 gnd.n4558 9.3005
R12050 gnd.n4560 gnd.n4535 9.3005
R12051 gnd.n4902 gnd.n4901 9.3005
R12052 gnd.n3927 gnd.n3916 9.3005
R12053 gnd.n3926 gnd.n3925 9.3005
R12054 gnd.n3924 gnd.n3917 9.3005
R12055 gnd.n3923 gnd.n3922 9.3005
R12056 gnd.n3921 gnd.n3920 9.3005
R12057 gnd.n2185 gnd.n2184 9.3005
R12058 gnd.n4367 gnd.n4366 9.3005
R12059 gnd.n4368 gnd.n2183 9.3005
R12060 gnd.n4370 gnd.n4369 9.3005
R12061 gnd.n2175 gnd.n2173 9.3005
R12062 gnd.n4411 gnd.n4410 9.3005
R12063 gnd.n4409 gnd.n2174 9.3005
R12064 gnd.n4408 gnd.n4407 9.3005
R12065 gnd.n4406 gnd.n2176 9.3005
R12066 gnd.n4405 gnd.n4404 9.3005
R12067 gnd.n4403 gnd.n4400 9.3005
R12068 gnd.n4402 gnd.n4401 9.3005
R12069 gnd.n2154 gnd.n2152 9.3005
R12070 gnd.n4460 gnd.n4459 9.3005
R12071 gnd.n4458 gnd.n2153 9.3005
R12072 gnd.n4457 gnd.n4456 9.3005
R12073 gnd.n4455 gnd.n2155 9.3005
R12074 gnd.n4454 gnd.n4453 9.3005
R12075 gnd.n2139 gnd.n2138 9.3005
R12076 gnd.n4516 gnd.n4515 9.3005
R12077 gnd.n4517 gnd.n2137 9.3005
R12078 gnd.n4519 gnd.n4518 9.3005
R12079 gnd.n2133 gnd.n2132 9.3005
R12080 gnd.n4533 gnd.n4532 9.3005
R12081 gnd.n4534 gnd.n2130 9.3005
R12082 gnd.n4566 gnd.n4565 9.3005
R12083 gnd.n4564 gnd.n2131 9.3005
R12084 gnd.n4562 gnd.n4561 9.3005
R12085 gnd.n2045 gnd.n2044 9.3005
R12086 gnd.n4853 gnd.n4852 9.3005
R12087 gnd.n4855 gnd.n4854 9.3005
R12088 gnd.n2033 gnd.n2032 9.3005
R12089 gnd.n4861 gnd.n4860 9.3005
R12090 gnd.n4863 gnd.n4862 9.3005
R12091 gnd.n2025 gnd.n2024 9.3005
R12092 gnd.n4869 gnd.n4868 9.3005
R12093 gnd.n4871 gnd.n4870 9.3005
R12094 gnd.n2015 gnd.n2014 9.3005
R12095 gnd.n4877 gnd.n4876 9.3005
R12096 gnd.n4879 gnd.n4878 9.3005
R12097 gnd.n2007 gnd.n2006 9.3005
R12098 gnd.n4885 gnd.n4884 9.3005
R12099 gnd.n4887 gnd.n4886 9.3005
R12100 gnd.n1997 gnd.n1995 9.3005
R12101 gnd.n4893 gnd.n4892 9.3005
R12102 gnd.n4894 gnd.n1994 9.3005
R12103 gnd.n2048 gnd.n1116 9.3005
R12104 gnd.n1998 gnd.n1996 9.3005
R12105 gnd.n4891 gnd.n4890 9.3005
R12106 gnd.n4889 gnd.n4888 9.3005
R12107 gnd.n2002 gnd.n2001 9.3005
R12108 gnd.n4883 gnd.n4882 9.3005
R12109 gnd.n4881 gnd.n4880 9.3005
R12110 gnd.n2011 gnd.n2010 9.3005
R12111 gnd.n4875 gnd.n4874 9.3005
R12112 gnd.n4873 gnd.n4872 9.3005
R12113 gnd.n2019 gnd.n2018 9.3005
R12114 gnd.n4867 gnd.n4866 9.3005
R12115 gnd.n4865 gnd.n4864 9.3005
R12116 gnd.n2029 gnd.n2028 9.3005
R12117 gnd.n4859 gnd.n4858 9.3005
R12118 gnd.n4857 gnd.n4856 9.3005
R12119 gnd.n2039 gnd.n2038 9.3005
R12120 gnd.n4851 gnd.n4850 9.3005
R12121 gnd.n6316 gnd.n1117 9.3005
R12122 gnd.n6315 gnd.n6314 9.3005
R12123 gnd.n6313 gnd.n1121 9.3005
R12124 gnd.n6312 gnd.n6311 9.3005
R12125 gnd.n6310 gnd.n1122 9.3005
R12126 gnd.n6309 gnd.n6308 9.3005
R12127 gnd.n6307 gnd.n1126 9.3005
R12128 gnd.n6306 gnd.n6305 9.3005
R12129 gnd.n6304 gnd.n1127 9.3005
R12130 gnd.n6303 gnd.n6302 9.3005
R12131 gnd.n6301 gnd.n1131 9.3005
R12132 gnd.n6300 gnd.n6299 9.3005
R12133 gnd.n6298 gnd.n1132 9.3005
R12134 gnd.n6297 gnd.n6296 9.3005
R12135 gnd.n6295 gnd.n1136 9.3005
R12136 gnd.n6294 gnd.n6293 9.3005
R12137 gnd.n6292 gnd.n1137 9.3005
R12138 gnd.n6291 gnd.n6290 9.3005
R12139 gnd.n6289 gnd.n1141 9.3005
R12140 gnd.n6288 gnd.n6287 9.3005
R12141 gnd.n6286 gnd.n1142 9.3005
R12142 gnd.n6285 gnd.n6284 9.3005
R12143 gnd.n6283 gnd.n1146 9.3005
R12144 gnd.n6282 gnd.n6281 9.3005
R12145 gnd.n6280 gnd.n1147 9.3005
R12146 gnd.n6279 gnd.n6278 9.3005
R12147 gnd.n6277 gnd.n1151 9.3005
R12148 gnd.n6276 gnd.n6275 9.3005
R12149 gnd.n6274 gnd.n1152 9.3005
R12150 gnd.n6273 gnd.n6272 9.3005
R12151 gnd.n6271 gnd.n1156 9.3005
R12152 gnd.n6270 gnd.n6269 9.3005
R12153 gnd.n6268 gnd.n1157 9.3005
R12154 gnd.n6267 gnd.n6266 9.3005
R12155 gnd.n6265 gnd.n1161 9.3005
R12156 gnd.n6264 gnd.n6263 9.3005
R12157 gnd.n6262 gnd.n1162 9.3005
R12158 gnd.n6261 gnd.n6260 9.3005
R12159 gnd.n6259 gnd.n1166 9.3005
R12160 gnd.n6258 gnd.n6257 9.3005
R12161 gnd.n6256 gnd.n1167 9.3005
R12162 gnd.n6255 gnd.n6254 9.3005
R12163 gnd.n6253 gnd.n1171 9.3005
R12164 gnd.n6252 gnd.n6251 9.3005
R12165 gnd.n6250 gnd.n1172 9.3005
R12166 gnd.n6249 gnd.n6248 9.3005
R12167 gnd.n6247 gnd.n1176 9.3005
R12168 gnd.n6246 gnd.n6245 9.3005
R12169 gnd.n6244 gnd.n1177 9.3005
R12170 gnd.n6243 gnd.n6242 9.3005
R12171 gnd.n6241 gnd.n1181 9.3005
R12172 gnd.n6240 gnd.n6239 9.3005
R12173 gnd.n6238 gnd.n1182 9.3005
R12174 gnd.n6237 gnd.n6236 9.3005
R12175 gnd.n6235 gnd.n1186 9.3005
R12176 gnd.n6234 gnd.n6233 9.3005
R12177 gnd.n6232 gnd.n1187 9.3005
R12178 gnd.n6231 gnd.n6230 9.3005
R12179 gnd.n6229 gnd.n1191 9.3005
R12180 gnd.n6228 gnd.n6227 9.3005
R12181 gnd.n6226 gnd.n1192 9.3005
R12182 gnd.n6225 gnd.n6224 9.3005
R12183 gnd.n6223 gnd.n1196 9.3005
R12184 gnd.n6222 gnd.n6221 9.3005
R12185 gnd.n6220 gnd.n1197 9.3005
R12186 gnd.n6219 gnd.n6218 9.3005
R12187 gnd.n6217 gnd.n1201 9.3005
R12188 gnd.n6216 gnd.n6215 9.3005
R12189 gnd.n6214 gnd.n1202 9.3005
R12190 gnd.n6213 gnd.n6212 9.3005
R12191 gnd.n6211 gnd.n1206 9.3005
R12192 gnd.n6210 gnd.n6209 9.3005
R12193 gnd.n6208 gnd.n1207 9.3005
R12194 gnd.n6207 gnd.n6206 9.3005
R12195 gnd.n6205 gnd.n1211 9.3005
R12196 gnd.n6204 gnd.n6203 9.3005
R12197 gnd.n6202 gnd.n1212 9.3005
R12198 gnd.n6201 gnd.n6200 9.3005
R12199 gnd.n6199 gnd.n1216 9.3005
R12200 gnd.n6198 gnd.n6197 9.3005
R12201 gnd.n6196 gnd.n1217 9.3005
R12202 gnd.n6195 gnd.n6194 9.3005
R12203 gnd.n6193 gnd.n1221 9.3005
R12204 gnd.n6192 gnd.n6191 9.3005
R12205 gnd.n6190 gnd.n1222 9.3005
R12206 gnd.n6189 gnd.n6188 9.3005
R12207 gnd.n6187 gnd.n1226 9.3005
R12208 gnd.n6186 gnd.n6185 9.3005
R12209 gnd.n6184 gnd.n1227 9.3005
R12210 gnd.n6183 gnd.n6182 9.3005
R12211 gnd.n6181 gnd.n1231 9.3005
R12212 gnd.n6180 gnd.n6179 9.3005
R12213 gnd.n6178 gnd.n1232 9.3005
R12214 gnd.n6177 gnd.n6176 9.3005
R12215 gnd.n6175 gnd.n1236 9.3005
R12216 gnd.n6174 gnd.n6173 9.3005
R12217 gnd.n6172 gnd.n1237 9.3005
R12218 gnd.n6171 gnd.n6170 9.3005
R12219 gnd.n6169 gnd.n1241 9.3005
R12220 gnd.n6168 gnd.n6167 9.3005
R12221 gnd.n6166 gnd.n1242 9.3005
R12222 gnd.n6318 gnd.n6317 9.3005
R12223 gnd.n6075 gnd.n1341 9.3005
R12224 gnd.n6074 gnd.n6073 9.3005
R12225 gnd.n6072 gnd.n1343 9.3005
R12226 gnd.n6071 gnd.n6070 9.3005
R12227 gnd.n6069 gnd.n1347 9.3005
R12228 gnd.n6068 gnd.n6067 9.3005
R12229 gnd.n6066 gnd.n1348 9.3005
R12230 gnd.n6065 gnd.n6064 9.3005
R12231 gnd.n6063 gnd.n1352 9.3005
R12232 gnd.n6062 gnd.n6061 9.3005
R12233 gnd.n6060 gnd.n1353 9.3005
R12234 gnd.n6059 gnd.n6058 9.3005
R12235 gnd.n6057 gnd.n1357 9.3005
R12236 gnd.n6056 gnd.n6055 9.3005
R12237 gnd.n6054 gnd.n1358 9.3005
R12238 gnd.n6053 gnd.n6052 9.3005
R12239 gnd.n407 gnd.n405 9.3005
R12240 gnd.n7233 gnd.n7232 9.3005
R12241 gnd.n7231 gnd.n406 9.3005
R12242 gnd.n7230 gnd.n7229 9.3005
R12243 gnd.n7228 gnd.n408 9.3005
R12244 gnd.n375 gnd.n373 9.3005
R12245 gnd.n7279 gnd.n7278 9.3005
R12246 gnd.n7277 gnd.n374 9.3005
R12247 gnd.n7276 gnd.n7275 9.3005
R12248 gnd.n7274 gnd.n376 9.3005
R12249 gnd.n7273 gnd.n7272 9.3005
R12250 gnd.n320 gnd.n318 9.3005
R12251 gnd.n7410 gnd.n7409 9.3005
R12252 gnd.n7408 gnd.n319 9.3005
R12253 gnd.n7407 gnd.n7406 9.3005
R12254 gnd.n7405 gnd.n321 9.3005
R12255 gnd.n7404 gnd.n7403 9.3005
R12256 gnd.n7402 gnd.n325 9.3005
R12257 gnd.n7401 gnd.n7400 9.3005
R12258 gnd.n7399 gnd.n326 9.3005
R12259 gnd.n297 gnd.n296 9.3005
R12260 gnd.n7424 gnd.n7423 9.3005
R12261 gnd.n7425 gnd.n295 9.3005
R12262 gnd.n7427 gnd.n7426 9.3005
R12263 gnd.n281 gnd.n280 9.3005
R12264 gnd.n7440 gnd.n7439 9.3005
R12265 gnd.n7441 gnd.n279 9.3005
R12266 gnd.n7443 gnd.n7442 9.3005
R12267 gnd.n267 gnd.n266 9.3005
R12268 gnd.n7456 gnd.n7455 9.3005
R12269 gnd.n7457 gnd.n265 9.3005
R12270 gnd.n7459 gnd.n7458 9.3005
R12271 gnd.n251 gnd.n250 9.3005
R12272 gnd.n7472 gnd.n7471 9.3005
R12273 gnd.n7473 gnd.n249 9.3005
R12274 gnd.n7475 gnd.n7474 9.3005
R12275 gnd.n236 gnd.n235 9.3005
R12276 gnd.n7488 gnd.n7487 9.3005
R12277 gnd.n7489 gnd.n234 9.3005
R12278 gnd.n7491 gnd.n7490 9.3005
R12279 gnd.n221 gnd.n220 9.3005
R12280 gnd.n7504 gnd.n7503 9.3005
R12281 gnd.n7505 gnd.n218 9.3005
R12282 gnd.n7575 gnd.n7574 9.3005
R12283 gnd.n7573 gnd.n219 9.3005
R12284 gnd.n7572 gnd.n7571 9.3005
R12285 gnd.n7570 gnd.n7506 9.3005
R12286 gnd.n7569 gnd.n7568 9.3005
R12287 gnd.n6077 gnd.n6076 9.3005
R12288 gnd.n7565 gnd.n7508 9.3005
R12289 gnd.n7564 gnd.n7563 9.3005
R12290 gnd.n7562 gnd.n7513 9.3005
R12291 gnd.n7561 gnd.n7560 9.3005
R12292 gnd.n7559 gnd.n7514 9.3005
R12293 gnd.n7558 gnd.n7557 9.3005
R12294 gnd.n7556 gnd.n7521 9.3005
R12295 gnd.n7555 gnd.n7554 9.3005
R12296 gnd.n7553 gnd.n7522 9.3005
R12297 gnd.n7552 gnd.n7551 9.3005
R12298 gnd.n7550 gnd.n7529 9.3005
R12299 gnd.n7549 gnd.n7548 9.3005
R12300 gnd.n7547 gnd.n7530 9.3005
R12301 gnd.n7546 gnd.n7545 9.3005
R12302 gnd.n7544 gnd.n7537 9.3005
R12303 gnd.n7543 gnd.n7542 9.3005
R12304 gnd.n124 gnd.n121 9.3005
R12305 gnd.n7669 gnd.n7668 9.3005
R12306 gnd.n7567 gnd.n7566 9.3005
R12307 gnd.n5917 gnd.n5916 9.3005
R12308 gnd.n5918 gnd.n1476 9.3005
R12309 gnd.n5921 gnd.n5920 9.3005
R12310 gnd.n5919 gnd.n1477 9.3005
R12311 gnd.n1420 gnd.n1419 9.3005
R12312 gnd.n5948 gnd.n5947 9.3005
R12313 gnd.n5949 gnd.n1417 9.3005
R12314 gnd.n5957 gnd.n5956 9.3005
R12315 gnd.n5955 gnd.n1418 9.3005
R12316 gnd.n5954 gnd.n5953 9.3005
R12317 gnd.n5952 gnd.n5950 9.3005
R12318 gnd.n1384 gnd.n1382 9.3005
R12319 gnd.n6017 gnd.n6016 9.3005
R12320 gnd.n6015 gnd.n1383 9.3005
R12321 gnd.n6014 gnd.n6013 9.3005
R12322 gnd.n6012 gnd.n1385 9.3005
R12323 gnd.n6011 gnd.n6010 9.3005
R12324 gnd.n6009 gnd.n6001 9.3005
R12325 gnd.n6008 gnd.n6007 9.3005
R12326 gnd.n6006 gnd.n6003 9.3005
R12327 gnd.n6002 gnd.n382 9.3005
R12328 gnd.n7261 gnd.n381 9.3005
R12329 gnd.n7263 gnd.n7262 9.3005
R12330 gnd.n7264 gnd.n379 9.3005
R12331 gnd.n7267 gnd.n7266 9.3005
R12332 gnd.n7265 gnd.n380 9.3005
R12333 gnd.n348 gnd.n347 9.3005
R12334 gnd.n7308 gnd.n7307 9.3005
R12335 gnd.n7309 gnd.n346 9.3005
R12336 gnd.n7311 gnd.n7310 9.3005
R12337 gnd.n7312 gnd.n79 9.3005
R12338 gnd.n7718 gnd.n80 9.3005
R12339 gnd.n7717 gnd.n7716 9.3005
R12340 gnd.n7715 gnd.n81 9.3005
R12341 gnd.n7714 gnd.n7713 9.3005
R12342 gnd.n7712 gnd.n85 9.3005
R12343 gnd.n7711 gnd.n7710 9.3005
R12344 gnd.n7709 gnd.n86 9.3005
R12345 gnd.n7708 gnd.n7707 9.3005
R12346 gnd.n7706 gnd.n90 9.3005
R12347 gnd.n7705 gnd.n7704 9.3005
R12348 gnd.n7703 gnd.n91 9.3005
R12349 gnd.n7702 gnd.n7701 9.3005
R12350 gnd.n7700 gnd.n95 9.3005
R12351 gnd.n7699 gnd.n7698 9.3005
R12352 gnd.n7697 gnd.n96 9.3005
R12353 gnd.n7696 gnd.n7695 9.3005
R12354 gnd.n7694 gnd.n100 9.3005
R12355 gnd.n7693 gnd.n7692 9.3005
R12356 gnd.n7691 gnd.n101 9.3005
R12357 gnd.n7690 gnd.n7689 9.3005
R12358 gnd.n7688 gnd.n105 9.3005
R12359 gnd.n7687 gnd.n7686 9.3005
R12360 gnd.n7685 gnd.n106 9.3005
R12361 gnd.n7684 gnd.n7683 9.3005
R12362 gnd.n7682 gnd.n110 9.3005
R12363 gnd.n7681 gnd.n7680 9.3005
R12364 gnd.n7679 gnd.n111 9.3005
R12365 gnd.n7678 gnd.n7677 9.3005
R12366 gnd.n7676 gnd.n115 9.3005
R12367 gnd.n7675 gnd.n7674 9.3005
R12368 gnd.n7673 gnd.n116 9.3005
R12369 gnd.n7672 gnd.n7671 9.3005
R12370 gnd.n7670 gnd.n120 9.3005
R12371 gnd.n5904 gnd.n5903 9.3005
R12372 gnd.t54 gnd.n2529 9.24152
R12373 gnd.n2431 gnd.t273 9.24152
R12374 gnd.n3711 gnd.t256 9.24152
R12375 gnd.t131 gnd.n2276 9.24152
R12376 gnd.n2198 gnd.n2197 9.24152
R12377 gnd.n7412 gnd.n312 9.24152
R12378 gnd.n263 gnd.t69 9.24152
R12379 gnd.t330 gnd.t54 8.92286
R12380 gnd.n5564 gnd.n1886 8.92286
R12381 gnd.n5588 gnd.t227 8.92286
R12382 gnd.n5628 gnd.n1827 8.92286
R12383 gnd.n5652 gnd.n1804 8.92286
R12384 gnd.n5463 gnd.n5108 8.92286
R12385 gnd.n5442 gnd.n5441 8.92286
R12386 gnd.n5764 gnd.n1707 8.92286
R12387 gnd.n5788 gnd.n1684 8.92286
R12388 gnd.n3681 gnd.n3656 8.92171
R12389 gnd.n3649 gnd.n3624 8.92171
R12390 gnd.n3617 gnd.n3592 8.92171
R12391 gnd.n3586 gnd.n3561 8.92171
R12392 gnd.n3554 gnd.n3529 8.92171
R12393 gnd.n3522 gnd.n3497 8.92171
R12394 gnd.n3490 gnd.n3465 8.92171
R12395 gnd.n3459 gnd.n3434 8.92171
R12396 gnd.n5203 gnd.n5185 8.72777
R12397 gnd.n3185 gnd.t88 8.60421
R12398 gnd.t143 gnd.n2308 8.60421
R12399 gnd.n232 gnd.t13 8.60421
R12400 gnd.n2609 gnd.n2589 8.43467
R12401 gnd.n58 gnd.n38 8.43467
R12402 gnd.n3928 gnd.n0 8.41456
R12403 gnd.n7719 gnd.n7718 8.41456
R12404 gnd.t302 gnd.n5005 8.28555
R12405 gnd.n5780 gnd.t283 8.28555
R12406 gnd.n3682 gnd.n3654 8.14595
R12407 gnd.n3650 gnd.n3622 8.14595
R12408 gnd.n3618 gnd.n3590 8.14595
R12409 gnd.n3587 gnd.n3559 8.14595
R12410 gnd.n3555 gnd.n3527 8.14595
R12411 gnd.n3523 gnd.n3495 8.14595
R12412 gnd.n3491 gnd.n3463 8.14595
R12413 gnd.n3460 gnd.n3432 8.14595
R12414 gnd.n3687 gnd.n3686 7.97301
R12415 gnd.t215 gnd.n2700 7.9669
R12416 gnd.n4897 gnd.n1979 7.9669
R12417 gnd.n1256 gnd.n1248 7.9669
R12418 gnd.n7668 gnd.n124 7.75808
R12419 gnd.n1595 gnd.n1594 7.75808
R12420 gnd.n4850 gnd.n2038 7.75808
R12421 gnd.n3881 gnd.n3820 7.75808
R12422 gnd.n6403 gnd.n970 7.64824
R12423 gnd.n6402 gnd.n973 7.64824
R12424 gnd.n4364 gnd.n983 7.64824
R12425 gnd.n6396 gnd.n986 7.64824
R12426 gnd.n4382 gnd.n4381 7.64824
R12427 gnd.n6390 gnd.n997 7.64824
R12428 gnd.n4414 gnd.n4413 7.64824
R12429 gnd.n6384 gnd.n1007 7.64824
R12430 gnd.n4390 gnd.n1015 7.64824
R12431 gnd.n6378 gnd.n1018 7.64824
R12432 gnd.n4398 gnd.n1026 7.64824
R12433 gnd.n6372 gnd.n1029 7.64824
R12434 gnd.n4431 gnd.n4430 7.64824
R12435 gnd.n6366 gnd.n1039 7.64824
R12436 gnd.n4463 gnd.n4462 7.64824
R12437 gnd.n6360 gnd.n1049 7.64824
R12438 gnd.n4439 gnd.n1057 7.64824
R12439 gnd.n6354 gnd.n1060 7.64824
R12440 gnd.n4451 gnd.n1068 7.64824
R12441 gnd.n6348 gnd.n1071 7.64824
R12442 gnd.n4513 gnd.n4512 7.64824
R12443 gnd.n6342 gnd.n1081 7.64824
R12444 gnd.n4521 gnd.n1089 7.64824
R12445 gnd.n6336 gnd.n1092 7.64824
R12446 gnd.n4530 gnd.n1100 7.64824
R12447 gnd.n4568 gnd.n1109 7.64824
R12448 gnd.n6324 gnd.n1112 7.64824
R12449 gnd.n5620 gnd.n1834 7.64824
R12450 gnd.n5498 gnd.t7 7.64824
R12451 gnd.n5660 gnd.n1796 7.64824
R12452 gnd.n5470 gnd.n5101 7.64824
R12453 gnd.t210 gnd.n1766 7.64824
R12454 gnd.n5434 gnd.n5133 7.64824
R12455 gnd.n5390 gnd.t249 7.64824
R12456 gnd.n6079 gnd.n1336 7.64824
R12457 gnd.n5914 gnd.n1338 7.64824
R12458 gnd.n5924 gnd.n5923 7.64824
R12459 gnd.n5935 gnd.n1431 7.64824
R12460 gnd.n5934 gnd.n1435 7.64824
R12461 gnd.n5945 gnd.n1422 7.64824
R12462 gnd.n1424 gnd.n1414 7.64824
R12463 gnd.n5960 gnd.n5959 7.64824
R12464 gnd.n5972 gnd.n1404 7.64824
R12465 gnd.n5970 gnd.n1407 7.64824
R12466 gnd.n5982 gnd.n1394 7.64824
R12467 gnd.n1398 gnd.n1396 7.64824
R12468 gnd.n6021 gnd.n6020 7.64824
R12469 gnd.n6042 gnd.n1370 7.64824
R12470 gnd.n6041 gnd.n1373 7.64824
R12471 gnd.n6050 gnd.n1361 7.64824
R12472 gnd.n5999 gnd.n1364 7.64824
R12473 gnd.n7235 gnd.n399 7.64824
R12474 gnd.n6004 gnd.n402 7.64824
R12475 gnd.n7245 gnd.n390 7.64824
R12476 gnd.n7226 gnd.n7225 7.64824
R12477 gnd.n7259 gnd.n384 7.64824
R12478 gnd.n7281 gnd.n367 7.64824
R12479 gnd.n7253 gnd.n370 7.64824
R12480 gnd.n7269 gnd.n377 7.64824
R12481 gnd.n7290 gnd.n356 7.64824
R12482 gnd.n358 gnd.n350 7.64824
R12483 gnd.n3094 gnd.t18 7.32958
R12484 gnd.n4914 gnd.t266 7.32958
R12485 gnd.n1942 gnd.t205 7.32958
R12486 gnd.t354 gnd.n1646 7.32958
R12487 gnd.n5873 gnd.t233 7.32958
R12488 gnd.n247 gnd.n238 7.32958
R12489 gnd.n4661 gnd.n4660 7.30353
R12490 gnd.n5202 gnd.n5201 7.30353
R12491 gnd.n3054 gnd.n2773 7.01093
R12492 gnd.n2776 gnd.n2774 7.01093
R12493 gnd.n3064 gnd.n3063 7.01093
R12494 gnd.n3075 gnd.n2757 7.01093
R12495 gnd.n3074 gnd.n2760 7.01093
R12496 gnd.n3085 gnd.n2748 7.01093
R12497 gnd.n2751 gnd.n2749 7.01093
R12498 gnd.n3095 gnd.n3094 7.01093
R12499 gnd.n3105 gnd.n2729 7.01093
R12500 gnd.n3104 gnd.n2732 7.01093
R12501 gnd.n3113 gnd.n2723 7.01093
R12502 gnd.n3125 gnd.n2713 7.01093
R12503 gnd.n3135 gnd.n2698 7.01093
R12504 gnd.n3151 gnd.n3150 7.01093
R12505 gnd.n2700 gnd.n2637 7.01093
R12506 gnd.n3205 gnd.n2638 7.01093
R12507 gnd.n3199 gnd.n3198 7.01093
R12508 gnd.n2687 gnd.n2649 7.01093
R12509 gnd.n3191 gnd.n2660 7.01093
R12510 gnd.n2678 gnd.n2673 7.01093
R12511 gnd.n3185 gnd.n3184 7.01093
R12512 gnd.n3231 gnd.n2564 7.01093
R12513 gnd.n3230 gnd.n3229 7.01093
R12514 gnd.n3242 gnd.n3241 7.01093
R12515 gnd.n2557 gnd.n2549 7.01093
R12516 gnd.n3271 gnd.n2537 7.01093
R12517 gnd.n3270 gnd.n2540 7.01093
R12518 gnd.n3281 gnd.n2529 7.01093
R12519 gnd.n2530 gnd.n2518 7.01093
R12520 gnd.n3292 gnd.n2519 7.01093
R12521 gnd.n3316 gnd.n2510 7.01093
R12522 gnd.n3315 gnd.n2501 7.01093
R12523 gnd.n3338 gnd.n3337 7.01093
R12524 gnd.n3356 gnd.n2482 7.01093
R12525 gnd.n3355 gnd.n2485 7.01093
R12526 gnd.n3366 gnd.n2474 7.01093
R12527 gnd.n2475 gnd.n2462 7.01093
R12528 gnd.n3377 gnd.n2463 7.01093
R12529 gnd.n3404 gnd.n2447 7.01093
R12530 gnd.n3416 gnd.n3415 7.01093
R12531 gnd.n3398 gnd.n2440 7.01093
R12532 gnd.n3427 gnd.n3426 7.01093
R12533 gnd.n3699 gnd.n2428 7.01093
R12534 gnd.n3698 gnd.n2431 7.01093
R12535 gnd.n3711 gnd.n2420 7.01093
R12536 gnd.n2421 gnd.n2412 7.01093
R12537 gnd.n3721 gnd.n2413 7.01093
R12538 gnd.n5505 gnd.t171 7.01093
R12539 gnd.t112 gnd.n1760 7.01093
R12540 gnd.n2732 gnd.t58 6.69227
R12541 gnd.n2540 gnd.t330 6.69227
R12542 gnd.n3405 gnd.t89 6.69227
R12543 gnd.t44 gnd.n1813 6.69227
R12544 gnd.n5457 gnd.t110 6.69227
R12545 gnd.n5307 gnd.n5306 6.5566
R12546 gnd.n4810 gnd.n4809 6.5566
R12547 gnd.n4685 gnd.n4679 6.5566
R12548 gnd.n5322 gnd.n5321 6.5566
R12549 gnd.n4748 gnd.t230 6.37362
R12550 gnd.t245 gnd.t328 6.37362
R12551 gnd.n5612 gnd.n1842 6.37362
R12552 gnd.n5512 gnd.t207 6.37362
R12553 gnd.n5668 gnd.n1789 6.37362
R12554 gnd.n5477 gnd.n5094 6.37362
R12555 gnd.n5708 gnd.t2 6.37362
R12556 gnd.n5427 gnd.n5426 6.37362
R12557 gnd.n4550 gnd.n4547 6.20656
R12558 gnd.n7630 gnd.n7627 6.20656
R12559 gnd.n4158 gnd.n4007 6.20656
R12560 gnd.n5892 gnd.n5889 6.20656
R12561 gnd.t157 gnd.n3161 6.05496
R12562 gnd.n3162 gnd.t16 6.05496
R12563 gnd.t39 gnd.n2564 6.05496
R12564 gnd.t43 gnd.n3326 6.05496
R12565 gnd.t186 gnd.n1840 6.05496
R12566 gnd.t352 gnd.t121 6.05496
R12567 gnd.t29 gnd.t342 6.05496
R12568 gnd.n5425 gnd.t358 6.05496
R12569 gnd.n3684 gnd.n3654 5.81868
R12570 gnd.n3652 gnd.n3622 5.81868
R12571 gnd.n3620 gnd.n3590 5.81868
R12572 gnd.n3589 gnd.n3559 5.81868
R12573 gnd.n3557 gnd.n3527 5.81868
R12574 gnd.n3525 gnd.n3495 5.81868
R12575 gnd.n3493 gnd.n3463 5.81868
R12576 gnd.n3462 gnd.n3432 5.81868
R12577 gnd.n5229 gnd.n1305 5.62001
R12578 gnd.n4817 gnd.n4617 5.62001
R12579 gnd.n4817 gnd.n4618 5.62001
R12580 gnd.n5316 gnd.n1305 5.62001
R12581 gnd.n2913 gnd.n2908 5.4308
R12582 gnd.n3729 gnd.n2405 5.4308
R12583 gnd.n3229 gnd.t214 5.41765
R12584 gnd.t41 gnd.n3252 5.41765
R12585 gnd.t116 gnd.n2494 5.41765
R12586 gnd.t118 gnd.n5556 5.09899
R12587 gnd.n5604 gnd.n1849 5.09899
R12588 gnd.n5484 gnd.n5087 5.09899
R12589 gnd.n5676 gnd.n1781 5.09899
R12590 gnd.n5419 gnd.n5148 5.09899
R12591 gnd.n5756 gnd.t1 5.09899
R12592 gnd.n3682 gnd.n3681 5.04292
R12593 gnd.n3650 gnd.n3649 5.04292
R12594 gnd.n3618 gnd.n3617 5.04292
R12595 gnd.n3587 gnd.n3586 5.04292
R12596 gnd.n3555 gnd.n3554 5.04292
R12597 gnd.n3523 gnd.n3522 5.04292
R12598 gnd.n3491 gnd.n3490 5.04292
R12599 gnd.n3460 gnd.n3459 5.04292
R12600 gnd.n2629 gnd.n2628 4.82753
R12601 gnd.n78 gnd.n77 4.82753
R12602 gnd.n3192 gnd.t17 4.78034
R12603 gnd.n2519 gnd.t55 4.78034
R12604 gnd.n4970 gnd.t149 4.78034
R12605 gnd.n5812 gnd.t155 4.78034
R12606 gnd.n2634 gnd.n2631 4.74817
R12607 gnd.n2684 gnd.n2570 4.74817
R12608 gnd.n2671 gnd.n2569 4.74817
R12609 gnd.n2568 gnd.n2567 4.74817
R12610 gnd.n2680 gnd.n2631 4.74817
R12611 gnd.n2681 gnd.n2570 4.74817
R12612 gnd.n2683 gnd.n2569 4.74817
R12613 gnd.n2670 gnd.n2568 4.74817
R12614 gnd.n7416 gnd.n7415 4.74817
R12615 gnd.n341 gnd.n308 4.74817
R12616 gnd.n7317 gnd.n307 4.74817
R12617 gnd.n331 gnd.n306 4.74817
R12618 gnd.n7395 gnd.n305 4.74817
R12619 gnd.n7416 gnd.n309 4.74817
R12620 gnd.n7414 gnd.n308 4.74817
R12621 gnd.n342 gnd.n307 4.74817
R12622 gnd.n7318 gnd.n306 4.74817
R12623 gnd.n332 gnd.n305 4.74817
R12624 gnd.n4310 gnd.n4308 4.74817
R12625 gnd.n4323 gnd.n2219 4.74817
R12626 gnd.n4327 gnd.n4325 4.74817
R12627 gnd.n4350 gnd.n2193 4.74817
R12628 gnd.n4353 gnd.n4352 4.74817
R12629 gnd.n4308 gnd.n4307 4.74817
R12630 gnd.n4309 gnd.n2219 4.74817
R12631 gnd.n4325 gnd.n4324 4.74817
R12632 gnd.n4326 gnd.n2193 4.74817
R12633 gnd.n4352 gnd.n4351 4.74817
R12634 gnd.n2609 gnd.n2608 4.7074
R12635 gnd.n58 gnd.n57 4.7074
R12636 gnd.n2629 gnd.n2609 4.65959
R12637 gnd.n78 gnd.n58 4.65959
R12638 gnd.n6123 gnd.n1307 4.6132
R12639 gnd.n4818 gnd.n4616 4.6132
R12640 gnd.n5054 gnd.t209 4.46168
R12641 gnd.n5716 gnd.t28 4.46168
R12642 gnd.t270 gnd.n1707 4.46168
R12643 gnd.n5198 gnd.n5185 4.46111
R12644 gnd.n3667 gnd.n3663 4.38594
R12645 gnd.n3635 gnd.n3631 4.38594
R12646 gnd.n3603 gnd.n3599 4.38594
R12647 gnd.n3572 gnd.n3568 4.38594
R12648 gnd.n3540 gnd.n3536 4.38594
R12649 gnd.n3508 gnd.n3504 4.38594
R12650 gnd.n3476 gnd.n3472 4.38594
R12651 gnd.n3445 gnd.n3441 4.38594
R12652 gnd.n3678 gnd.n3656 4.26717
R12653 gnd.n3646 gnd.n3624 4.26717
R12654 gnd.n3614 gnd.n3592 4.26717
R12655 gnd.n3583 gnd.n3561 4.26717
R12656 gnd.n3551 gnd.n3529 4.26717
R12657 gnd.n3519 gnd.n3497 4.26717
R12658 gnd.n3487 gnd.n3465 4.26717
R12659 gnd.n3456 gnd.n3434 4.26717
R12660 gnd.n3136 gnd.t53 4.14303
R12661 gnd.n3366 gnd.t57 4.14303
R12662 gnd.n2129 gnd.t237 4.14303
R12663 gnd.n5905 gnd.t241 4.14303
R12664 gnd.n3686 gnd.n3685 4.08274
R12665 gnd.n5306 gnd.n5305 4.05904
R12666 gnd.n4809 gnd.n4808 4.05904
R12667 gnd.n4689 gnd.n4679 4.05904
R12668 gnd.n5323 gnd.n5322 4.05904
R12669 gnd.n19 gnd.n9 3.99943
R12670 gnd.n5596 gnd.n1857 3.82437
R12671 gnd.n5542 gnd.t124 3.82437
R12672 gnd.n5534 gnd.n5039 3.82437
R12673 gnd.n5491 gnd.n5080 3.82437
R12674 gnd.n5684 gnd.n1774 3.82437
R12675 gnd.n5732 gnd.n1732 3.82437
R12676 gnd.n5147 gnd.t188 3.82437
R12677 gnd.n5412 gnd.n5411 3.82437
R12678 gnd.n3686 gnd.n3558 3.70378
R12679 gnd.n3209 gnd.n2630 3.65935
R12680 gnd.n19 gnd.n18 3.60163
R12681 gnd.n4207 gnd.t305 3.50571
R12682 gnd.n6330 gnd.t237 3.50571
R12683 gnd.t241 gnd.n1452 3.50571
R12684 gnd.n7585 gnd.t223 3.50571
R12685 gnd.n3677 gnd.n3658 3.49141
R12686 gnd.n3645 gnd.n3626 3.49141
R12687 gnd.n3613 gnd.n3594 3.49141
R12688 gnd.n3582 gnd.n3563 3.49141
R12689 gnd.n3550 gnd.n3531 3.49141
R12690 gnd.n3518 gnd.n3499 3.49141
R12691 gnd.n3486 gnd.n3467 3.49141
R12692 gnd.n3455 gnd.n3436 3.49141
R12693 gnd.n5006 gnd.t302 3.18706
R12694 gnd.n5549 gnd.t85 3.18706
R12695 gnd.t85 gnd.n5026 3.18706
R12696 gnd.n5748 gnd.t189 3.18706
R12697 gnd.n5413 gnd.t189 3.18706
R12698 gnd.n2715 gnd.t53 2.8684
R12699 gnd.n1910 gnd.n1901 2.8684
R12700 gnd.n5572 gnd.t59 2.8684
R12701 gnd.n5179 gnd.t218 2.8684
R12702 gnd.n1687 gnd.n1686 2.8684
R12703 gnd.n2610 gnd.t161 2.82907
R12704 gnd.n2610 gnd.t192 2.82907
R12705 gnd.n2612 gnd.t204 2.82907
R12706 gnd.n2612 gnd.t194 2.82907
R12707 gnd.n2614 gnd.t191 2.82907
R12708 gnd.n2614 gnd.t196 2.82907
R12709 gnd.n2616 gnd.t142 2.82907
R12710 gnd.n2616 gnd.t94 2.82907
R12711 gnd.n2618 gnd.t202 2.82907
R12712 gnd.n2618 gnd.t185 2.82907
R12713 gnd.n2620 gnd.t92 2.82907
R12714 gnd.n2620 gnd.t99 2.82907
R12715 gnd.n2622 gnd.t203 2.82907
R12716 gnd.n2622 gnd.t213 2.82907
R12717 gnd.n2624 gnd.t147 2.82907
R12718 gnd.n2624 gnd.t91 2.82907
R12719 gnd.n2626 gnd.t163 2.82907
R12720 gnd.n2626 gnd.t100 2.82907
R12721 gnd.n2571 gnd.t356 2.82907
R12722 gnd.n2571 gnd.t129 2.82907
R12723 gnd.n2573 gnd.t165 2.82907
R12724 gnd.n2573 gnd.t135 2.82907
R12725 gnd.n2575 gnd.t84 2.82907
R12726 gnd.n2575 gnd.t31 2.82907
R12727 gnd.n2577 gnd.t160 2.82907
R12728 gnd.n2577 gnd.t180 2.82907
R12729 gnd.n2579 gnd.t20 2.82907
R12730 gnd.n2579 gnd.t172 2.82907
R12731 gnd.n2581 gnd.t164 2.82907
R12732 gnd.n2581 gnd.t67 2.82907
R12733 gnd.n2583 gnd.t221 2.82907
R12734 gnd.n2583 gnd.t98 2.82907
R12735 gnd.n2585 gnd.t132 2.82907
R12736 gnd.n2585 gnd.t179 2.82907
R12737 gnd.n2587 gnd.t220 2.82907
R12738 gnd.n2587 gnd.t159 2.82907
R12739 gnd.n2590 gnd.t35 2.82907
R12740 gnd.n2590 gnd.t344 2.82907
R12741 gnd.n2592 gnd.t96 2.82907
R12742 gnd.n2592 gnd.t78 2.82907
R12743 gnd.n2594 gnd.t115 2.82907
R12744 gnd.n2594 gnd.t82 2.82907
R12745 gnd.n2596 gnd.t10 2.82907
R12746 gnd.n2596 gnd.t177 2.82907
R12747 gnd.n2598 gnd.t348 2.82907
R12748 gnd.n2598 gnd.t37 2.82907
R12749 gnd.n2600 gnd.t66 2.82907
R12750 gnd.n2600 gnd.t64 2.82907
R12751 gnd.n2602 gnd.t137 2.82907
R12752 gnd.n2602 gnd.t126 2.82907
R12753 gnd.n2604 gnd.t166 2.82907
R12754 gnd.n2604 gnd.t134 2.82907
R12755 gnd.n2606 gnd.t212 2.82907
R12756 gnd.n2606 gnd.t76 2.82907
R12757 gnd.n75 gnd.t52 2.82907
R12758 gnd.n75 gnd.t141 2.82907
R12759 gnd.n73 gnd.t105 2.82907
R12760 gnd.n73 gnd.t190 2.82907
R12761 gnd.n71 gnd.t184 2.82907
R12762 gnd.n71 gnd.t195 2.82907
R12763 gnd.n69 gnd.t38 2.82907
R12764 gnd.n69 gnd.t74 2.82907
R12765 gnd.n67 gnd.t101 2.82907
R12766 gnd.n67 gnd.t72 2.82907
R12767 gnd.n65 gnd.t102 2.82907
R12768 gnd.n65 gnd.t198 2.82907
R12769 gnd.n63 gnd.t51 2.82907
R12770 gnd.n63 gnd.t103 2.82907
R12771 gnd.n61 gnd.t148 2.82907
R12772 gnd.n61 gnd.t193 2.82907
R12773 gnd.n59 gnd.t146 2.82907
R12774 gnd.n59 gnd.t140 2.82907
R12775 gnd.n36 gnd.t68 2.82907
R12776 gnd.n36 gnd.t176 2.82907
R12777 gnd.n34 gnd.t182 2.82907
R12778 gnd.n34 gnd.t113 2.82907
R12779 gnd.n32 gnd.t332 2.82907
R12780 gnd.n32 gnd.t26 2.82907
R12781 gnd.n30 gnd.t33 2.82907
R12782 gnd.n30 gnd.t211 2.82907
R12783 gnd.n28 gnd.t345 2.82907
R12784 gnd.n28 gnd.t125 2.82907
R12785 gnd.n26 gnd.t349 2.82907
R12786 gnd.n26 gnd.t338 2.82907
R12787 gnd.n24 gnd.t79 2.82907
R12788 gnd.n24 gnd.t175 2.82907
R12789 gnd.n22 gnd.t181 2.82907
R12790 gnd.n22 gnd.t174 2.82907
R12791 gnd.n20 gnd.t337 2.82907
R12792 gnd.n20 gnd.t199 2.82907
R12793 gnd.n55 gnd.t22 2.82907
R12794 gnd.n55 gnd.t49 2.82907
R12795 gnd.n53 gnd.t347 2.82907
R12796 gnd.n53 gnd.t70 2.82907
R12797 gnd.n51 gnd.t357 2.82907
R12798 gnd.n51 gnd.t178 2.82907
R12799 gnd.n49 gnd.t333 2.82907
R12800 gnd.n49 gnd.t336 2.82907
R12801 gnd.n47 gnd.t87 2.82907
R12802 gnd.n47 gnd.t114 2.82907
R12803 gnd.n45 gnd.t24 2.82907
R12804 gnd.n45 gnd.t201 2.82907
R12805 gnd.n43 gnd.t127 2.82907
R12806 gnd.n43 gnd.t47 2.82907
R12807 gnd.n41 gnd.t139 2.82907
R12808 gnd.n41 gnd.t81 2.82907
R12809 gnd.n39 gnd.t200 2.82907
R12810 gnd.n39 gnd.t62 2.82907
R12811 gnd.n3674 gnd.n3673 2.71565
R12812 gnd.n3642 gnd.n3641 2.71565
R12813 gnd.n3610 gnd.n3609 2.71565
R12814 gnd.n3579 gnd.n3578 2.71565
R12815 gnd.n3547 gnd.n3546 2.71565
R12816 gnd.n3515 gnd.n3514 2.71565
R12817 gnd.n3483 gnd.n3482 2.71565
R12818 gnd.n3452 gnd.n3451 2.71565
R12819 gnd.n4996 gnd.t230 2.54975
R12820 gnd.n5013 gnd.t245 2.54975
R12821 gnd.n5588 gnd.n1863 2.54975
R12822 gnd.n5557 gnd.t118 2.54975
R12823 gnd.n5527 gnd.n5526 2.54975
R12824 gnd.n5526 gnd.t208 2.54975
R12825 gnd.n5498 gnd.n5073 2.54975
R12826 gnd.n5692 gnd.n1766 2.54975
R12827 gnd.n5724 gnd.t27 2.54975
R12828 gnd.n5724 gnd.n1739 2.54975
R12829 gnd.n5405 gnd.t1 2.54975
R12830 gnd.n5162 gnd.n5161 2.54975
R12831 gnd.n5772 gnd.t249 2.54975
R12832 gnd.n5390 gnd.t252 2.54975
R12833 gnd.n3209 gnd.n2631 2.27742
R12834 gnd.n3209 gnd.n2570 2.27742
R12835 gnd.n3209 gnd.n2569 2.27742
R12836 gnd.n3209 gnd.n2568 2.27742
R12837 gnd.n7417 gnd.n7416 2.27742
R12838 gnd.n7417 gnd.n308 2.27742
R12839 gnd.n7417 gnd.n307 2.27742
R12840 gnd.n7417 gnd.n306 2.27742
R12841 gnd.n7417 gnd.n305 2.27742
R12842 gnd.n4308 gnd.n966 2.27742
R12843 gnd.n2219 gnd.n966 2.27742
R12844 gnd.n4325 gnd.n966 2.27742
R12845 gnd.n2193 gnd.n966 2.27742
R12846 gnd.n4352 gnd.n966 2.27742
R12847 gnd.n3063 gnd.t312 2.23109
R12848 gnd.n2686 gnd.t17 2.23109
R12849 gnd.n4381 gnd.t83 2.23109
R12850 gnd.n5491 gnd.t352 2.23109
R12851 gnd.t342 gnd.n1774 2.23109
R12852 gnd.t46 gnd.n367 2.23109
R12853 gnd.n3670 gnd.n3660 1.93989
R12854 gnd.n3638 gnd.n3628 1.93989
R12855 gnd.n3606 gnd.n3596 1.93989
R12856 gnd.n3575 gnd.n3565 1.93989
R12857 gnd.n3543 gnd.n3533 1.93989
R12858 gnd.n3511 gnd.n3501 1.93989
R12859 gnd.n3479 gnd.n3469 1.93989
R12860 gnd.n3448 gnd.n3438 1.93989
R12861 gnd.n5384 gnd.t283 1.91244
R12862 gnd.n1686 gnd.t286 1.91244
R12863 gnd.t169 gnd.n3074 1.59378
R12864 gnd.n3253 gnd.t41 1.59378
R12865 gnd.n2503 gnd.t116 1.59378
R12866 gnd.n4247 gnd.t75 1.59378
R12867 gnd.n4430 gnd.t77 1.59378
R12868 gnd.n6360 gnd.t34 1.59378
R12869 gnd.n5557 gnd.t119 1.59378
R12870 gnd.n5628 gnd.t108 1.59378
R12871 gnd.n5441 gnd.t151 1.59378
R12872 gnd.n5405 gnd.t350 1.59378
R12873 gnd.n1398 gnd.t61 1.59378
R12874 gnd.t138 gnd.n6041 1.59378
R12875 gnd.n7477 gnd.t21 1.59378
R12876 gnd.n4641 gnd.n1893 1.27512
R12877 gnd.n5580 gnd.n1871 1.27512
R12878 gnd.t124 gnd.n5541 1.27512
R12879 gnd.n5519 gnd.n5054 1.27512
R12880 gnd.n5505 gnd.n5066 1.27512
R12881 gnd.n5700 gnd.n1760 1.27512
R12882 gnd.n5716 gnd.n1745 1.27512
R12883 gnd.n5740 gnd.t188 1.27512
R12884 gnd.n5397 gnd.n5396 1.27512
R12885 gnd.n5378 gnd.n5183 1.27512
R12886 gnd.n2916 gnd.n2908 1.16414
R12887 gnd.n3732 gnd.n2405 1.16414
R12888 gnd.n3669 gnd.n3662 1.16414
R12889 gnd.n3637 gnd.n3630 1.16414
R12890 gnd.n3605 gnd.n3598 1.16414
R12891 gnd.n3574 gnd.n3567 1.16414
R12892 gnd.n3542 gnd.n3535 1.16414
R12893 gnd.n3510 gnd.n3503 1.16414
R12894 gnd.n3478 gnd.n3471 1.16414
R12895 gnd.n3447 gnd.n3440 1.16414
R12896 gnd.n6123 gnd.n6122 0.970197
R12897 gnd.n4818 gnd.n2102 0.970197
R12898 gnd.n3653 gnd.n3621 0.962709
R12899 gnd.n3685 gnd.n3653 0.962709
R12900 gnd.n3526 gnd.n3494 0.962709
R12901 gnd.n3558 gnd.n3526 0.962709
R12902 gnd.n3162 gnd.t157 0.956468
R12903 gnd.n3327 gnd.t43 0.956468
R12904 gnd.n4279 gnd.t136 0.956468
R12905 gnd.n6384 gnd.t30 0.956468
R12906 gnd.n4512 gnd.t106 0.956468
R12907 gnd.t11 gnd.n1424 0.956468
R12908 gnd.n7245 gnd.t50 0.956468
R12909 gnd.n7445 gnd.t25 0.956468
R12910 gnd.n2621 gnd.n2619 0.773756
R12911 gnd.n70 gnd.n68 0.773756
R12912 gnd.n2628 gnd.n2627 0.773756
R12913 gnd.n2627 gnd.n2625 0.773756
R12914 gnd.n2625 gnd.n2623 0.773756
R12915 gnd.n2623 gnd.n2621 0.773756
R12916 gnd.n2619 gnd.n2617 0.773756
R12917 gnd.n2617 gnd.n2615 0.773756
R12918 gnd.n2615 gnd.n2613 0.773756
R12919 gnd.n2613 gnd.n2611 0.773756
R12920 gnd.n62 gnd.n60 0.773756
R12921 gnd.n64 gnd.n62 0.773756
R12922 gnd.n66 gnd.n64 0.773756
R12923 gnd.n68 gnd.n66 0.773756
R12924 gnd.n72 gnd.n70 0.773756
R12925 gnd.n74 gnd.n72 0.773756
R12926 gnd.n76 gnd.n74 0.773756
R12927 gnd.n77 gnd.n76 0.773756
R12928 gnd gnd.n0 0.70738
R12929 gnd.n2 gnd.n1 0.672012
R12930 gnd.n3 gnd.n2 0.672012
R12931 gnd.n4 gnd.n3 0.672012
R12932 gnd.n5 gnd.n4 0.672012
R12933 gnd.n6 gnd.n5 0.672012
R12934 gnd.n7 gnd.n6 0.672012
R12935 gnd.n8 gnd.n7 0.672012
R12936 gnd.n9 gnd.n8 0.672012
R12937 gnd.n11 gnd.n10 0.672012
R12938 gnd.n12 gnd.n11 0.672012
R12939 gnd.n13 gnd.n12 0.672012
R12940 gnd.n14 gnd.n13 0.672012
R12941 gnd.n15 gnd.n14 0.672012
R12942 gnd.n16 gnd.n15 0.672012
R12943 gnd.n17 gnd.n16 0.672012
R12944 gnd.n18 gnd.n17 0.672012
R12945 gnd.t277 gnd.n1871 0.637812
R12946 gnd.n5039 gnd.t0 0.637812
R12947 gnd.n5732 gnd.t8 0.637812
R12948 gnd.n7720 gnd.n7719 0.637193
R12949 gnd.n2589 gnd.n2588 0.573776
R12950 gnd.n2588 gnd.n2586 0.573776
R12951 gnd.n2586 gnd.n2584 0.573776
R12952 gnd.n2584 gnd.n2582 0.573776
R12953 gnd.n2582 gnd.n2580 0.573776
R12954 gnd.n2580 gnd.n2578 0.573776
R12955 gnd.n2578 gnd.n2576 0.573776
R12956 gnd.n2576 gnd.n2574 0.573776
R12957 gnd.n2574 gnd.n2572 0.573776
R12958 gnd.n2608 gnd.n2607 0.573776
R12959 gnd.n2607 gnd.n2605 0.573776
R12960 gnd.n2605 gnd.n2603 0.573776
R12961 gnd.n2603 gnd.n2601 0.573776
R12962 gnd.n2601 gnd.n2599 0.573776
R12963 gnd.n2599 gnd.n2597 0.573776
R12964 gnd.n2597 gnd.n2595 0.573776
R12965 gnd.n2595 gnd.n2593 0.573776
R12966 gnd.n2593 gnd.n2591 0.573776
R12967 gnd.n23 gnd.n21 0.573776
R12968 gnd.n25 gnd.n23 0.573776
R12969 gnd.n27 gnd.n25 0.573776
R12970 gnd.n29 gnd.n27 0.573776
R12971 gnd.n31 gnd.n29 0.573776
R12972 gnd.n33 gnd.n31 0.573776
R12973 gnd.n35 gnd.n33 0.573776
R12974 gnd.n37 gnd.n35 0.573776
R12975 gnd.n38 gnd.n37 0.573776
R12976 gnd.n42 gnd.n40 0.573776
R12977 gnd.n44 gnd.n42 0.573776
R12978 gnd.n46 gnd.n44 0.573776
R12979 gnd.n48 gnd.n46 0.573776
R12980 gnd.n50 gnd.n48 0.573776
R12981 gnd.n52 gnd.n50 0.573776
R12982 gnd.n54 gnd.n52 0.573776
R12983 gnd.n56 gnd.n54 0.573776
R12984 gnd.n57 gnd.n56 0.573776
R12985 gnd.n7417 gnd.n304 0.5435
R12986 gnd.n6407 gnd.n966 0.5435
R12987 gnd.n3389 gnd.n2409 0.486781
R12988 gnd.n1518 gnd.n1242 0.486781
R12989 gnd.n2965 gnd.n2964 0.48678
R12990 gnd.n6319 gnd.n6318 0.485256
R12991 gnd.n3706 gnd.n2363 0.480683
R12992 gnd.n3049 gnd.n3048 0.480683
R12993 gnd.n6579 gnd.n6578 0.480683
R12994 gnd.n7000 gnd.n6999 0.480683
R12995 gnd.n3883 gnd.n3882 0.477634
R12996 gnd.n4202 gnd.n2337 0.477634
R12997 gnd.n7568 gnd.n7567 0.477634
R12998 gnd.n7670 gnd.n7669 0.477634
R12999 gnd.n7662 gnd.n7661 0.465439
R13000 gnd.n7591 gnd.n7590 0.465439
R13001 gnd.n6083 gnd.n1333 0.465439
R13002 gnd.n5908 gnd.n1289 0.465439
R13003 gnd.n2086 gnd.n1107 0.465439
R13004 gnd.n4573 gnd.n4572 0.465439
R13005 gnd.n4121 gnd.n4116 0.465439
R13006 gnd.n4196 gnd.n4195 0.465439
R13007 gnd.n5879 gnd.n5878 0.451719
R13008 gnd.n4903 gnd.n4902 0.451719
R13009 gnd.n4553 gnd.n4547 0.388379
R13010 gnd.n3666 gnd.n3665 0.388379
R13011 gnd.n3634 gnd.n3633 0.388379
R13012 gnd.n3602 gnd.n3601 0.388379
R13013 gnd.n3571 gnd.n3570 0.388379
R13014 gnd.n3539 gnd.n3538 0.388379
R13015 gnd.n3507 gnd.n3506 0.388379
R13016 gnd.n3475 gnd.n3474 0.388379
R13017 gnd.n3444 gnd.n3443 0.388379
R13018 gnd.n7631 gnd.n7630 0.388379
R13019 gnd.n4007 gnd.n4003 0.388379
R13020 gnd.n5893 gnd.n5892 0.388379
R13021 gnd.n6321 gnd.n6320 0.378829
R13022 gnd.n6076 gnd.n1342 0.377553
R13023 gnd.n7720 gnd.n19 0.374463
R13024 gnd gnd.n7720 0.367492
R13025 gnd.n2465 gnd.t89 0.319156
R13026 gnd.n4312 gnd.t63 0.319156
R13027 gnd.n4355 gnd.t9 0.319156
R13028 gnd.n7305 gnd.t197 0.319156
R13029 gnd.n7397 gnd.t32 0.319156
R13030 gnd.n2883 gnd.n2861 0.311721
R13031 gnd.n7211 gnd.n304 0.282512
R13032 gnd.n6408 gnd.n6407 0.282512
R13033 gnd.n3777 gnd.n3776 0.268793
R13034 gnd.n4564 gnd.n4563 0.247451
R13035 gnd.n5903 gnd.n5902 0.247451
R13036 gnd.n3776 gnd.n3775 0.241354
R13037 gnd.n1307 gnd.n1304 0.229039
R13038 gnd.n1310 gnd.n1307 0.229039
R13039 gnd.n4616 gnd.n2101 0.229039
R13040 gnd.n4616 gnd.n4615 0.229039
R13041 gnd.n2630 gnd.n0 0.210825
R13042 gnd.n3037 gnd.n2836 0.206293
R13043 gnd.n420 gnd.n304 0.198671
R13044 gnd.n6407 gnd.n6406 0.198671
R13045 gnd.n3683 gnd.n3655 0.155672
R13046 gnd.n3676 gnd.n3655 0.155672
R13047 gnd.n3676 gnd.n3675 0.155672
R13048 gnd.n3675 gnd.n3659 0.155672
R13049 gnd.n3668 gnd.n3659 0.155672
R13050 gnd.n3668 gnd.n3667 0.155672
R13051 gnd.n3651 gnd.n3623 0.155672
R13052 gnd.n3644 gnd.n3623 0.155672
R13053 gnd.n3644 gnd.n3643 0.155672
R13054 gnd.n3643 gnd.n3627 0.155672
R13055 gnd.n3636 gnd.n3627 0.155672
R13056 gnd.n3636 gnd.n3635 0.155672
R13057 gnd.n3619 gnd.n3591 0.155672
R13058 gnd.n3612 gnd.n3591 0.155672
R13059 gnd.n3612 gnd.n3611 0.155672
R13060 gnd.n3611 gnd.n3595 0.155672
R13061 gnd.n3604 gnd.n3595 0.155672
R13062 gnd.n3604 gnd.n3603 0.155672
R13063 gnd.n3588 gnd.n3560 0.155672
R13064 gnd.n3581 gnd.n3560 0.155672
R13065 gnd.n3581 gnd.n3580 0.155672
R13066 gnd.n3580 gnd.n3564 0.155672
R13067 gnd.n3573 gnd.n3564 0.155672
R13068 gnd.n3573 gnd.n3572 0.155672
R13069 gnd.n3556 gnd.n3528 0.155672
R13070 gnd.n3549 gnd.n3528 0.155672
R13071 gnd.n3549 gnd.n3548 0.155672
R13072 gnd.n3548 gnd.n3532 0.155672
R13073 gnd.n3541 gnd.n3532 0.155672
R13074 gnd.n3541 gnd.n3540 0.155672
R13075 gnd.n3524 gnd.n3496 0.155672
R13076 gnd.n3517 gnd.n3496 0.155672
R13077 gnd.n3517 gnd.n3516 0.155672
R13078 gnd.n3516 gnd.n3500 0.155672
R13079 gnd.n3509 gnd.n3500 0.155672
R13080 gnd.n3509 gnd.n3508 0.155672
R13081 gnd.n3492 gnd.n3464 0.155672
R13082 gnd.n3485 gnd.n3464 0.155672
R13083 gnd.n3485 gnd.n3484 0.155672
R13084 gnd.n3484 gnd.n3468 0.155672
R13085 gnd.n3477 gnd.n3468 0.155672
R13086 gnd.n3477 gnd.n3476 0.155672
R13087 gnd.n3461 gnd.n3433 0.155672
R13088 gnd.n3454 gnd.n3433 0.155672
R13089 gnd.n3454 gnd.n3453 0.155672
R13090 gnd.n3453 gnd.n3437 0.155672
R13091 gnd.n3446 gnd.n3437 0.155672
R13092 gnd.n3446 gnd.n3445 0.155672
R13093 gnd.n3808 gnd.n2363 0.152939
R13094 gnd.n3808 gnd.n3807 0.152939
R13095 gnd.n3807 gnd.n3806 0.152939
R13096 gnd.n3806 gnd.n2365 0.152939
R13097 gnd.n2366 gnd.n2365 0.152939
R13098 gnd.n2367 gnd.n2366 0.152939
R13099 gnd.n2368 gnd.n2367 0.152939
R13100 gnd.n2369 gnd.n2368 0.152939
R13101 gnd.n2370 gnd.n2369 0.152939
R13102 gnd.n2371 gnd.n2370 0.152939
R13103 gnd.n2372 gnd.n2371 0.152939
R13104 gnd.n2373 gnd.n2372 0.152939
R13105 gnd.n2374 gnd.n2373 0.152939
R13106 gnd.n2375 gnd.n2374 0.152939
R13107 gnd.n3778 gnd.n2375 0.152939
R13108 gnd.n3778 gnd.n3777 0.152939
R13109 gnd.n3050 gnd.n3049 0.152939
R13110 gnd.n3050 gnd.n2754 0.152939
R13111 gnd.n3078 gnd.n2754 0.152939
R13112 gnd.n3079 gnd.n3078 0.152939
R13113 gnd.n3080 gnd.n3079 0.152939
R13114 gnd.n3081 gnd.n3080 0.152939
R13115 gnd.n3081 gnd.n2726 0.152939
R13116 gnd.n3108 gnd.n2726 0.152939
R13117 gnd.n3109 gnd.n3108 0.152939
R13118 gnd.n3110 gnd.n3109 0.152939
R13119 gnd.n3110 gnd.n2704 0.152939
R13120 gnd.n3139 gnd.n2704 0.152939
R13121 gnd.n3140 gnd.n3139 0.152939
R13122 gnd.n3141 gnd.n3140 0.152939
R13123 gnd.n3142 gnd.n3141 0.152939
R13124 gnd.n3144 gnd.n3142 0.152939
R13125 gnd.n3144 gnd.n3143 0.152939
R13126 gnd.n3143 gnd.n2653 0.152939
R13127 gnd.n2654 gnd.n2653 0.152939
R13128 gnd.n2655 gnd.n2654 0.152939
R13129 gnd.n2674 gnd.n2655 0.152939
R13130 gnd.n2675 gnd.n2674 0.152939
R13131 gnd.n2675 gnd.n2561 0.152939
R13132 gnd.n3234 gnd.n2561 0.152939
R13133 gnd.n3235 gnd.n3234 0.152939
R13134 gnd.n3236 gnd.n3235 0.152939
R13135 gnd.n3237 gnd.n3236 0.152939
R13136 gnd.n3237 gnd.n2534 0.152939
R13137 gnd.n3274 gnd.n2534 0.152939
R13138 gnd.n3275 gnd.n3274 0.152939
R13139 gnd.n3276 gnd.n3275 0.152939
R13140 gnd.n3277 gnd.n3276 0.152939
R13141 gnd.n3277 gnd.n2507 0.152939
R13142 gnd.n3319 gnd.n2507 0.152939
R13143 gnd.n3320 gnd.n3319 0.152939
R13144 gnd.n3321 gnd.n3320 0.152939
R13145 gnd.n3322 gnd.n3321 0.152939
R13146 gnd.n3322 gnd.n2479 0.152939
R13147 gnd.n3359 gnd.n2479 0.152939
R13148 gnd.n3360 gnd.n3359 0.152939
R13149 gnd.n3361 gnd.n3360 0.152939
R13150 gnd.n3362 gnd.n3361 0.152939
R13151 gnd.n3362 gnd.n2452 0.152939
R13152 gnd.n3408 gnd.n2452 0.152939
R13153 gnd.n3409 gnd.n3408 0.152939
R13154 gnd.n3410 gnd.n3409 0.152939
R13155 gnd.n3411 gnd.n3410 0.152939
R13156 gnd.n3411 gnd.n2425 0.152939
R13157 gnd.n3702 gnd.n2425 0.152939
R13158 gnd.n3703 gnd.n3702 0.152939
R13159 gnd.n3704 gnd.n3703 0.152939
R13160 gnd.n3705 gnd.n3704 0.152939
R13161 gnd.n3706 gnd.n3705 0.152939
R13162 gnd.n3048 gnd.n2778 0.152939
R13163 gnd.n2799 gnd.n2778 0.152939
R13164 gnd.n2800 gnd.n2799 0.152939
R13165 gnd.n2806 gnd.n2800 0.152939
R13166 gnd.n2807 gnd.n2806 0.152939
R13167 gnd.n2808 gnd.n2807 0.152939
R13168 gnd.n2808 gnd.n2797 0.152939
R13169 gnd.n2816 gnd.n2797 0.152939
R13170 gnd.n2817 gnd.n2816 0.152939
R13171 gnd.n2818 gnd.n2817 0.152939
R13172 gnd.n2818 gnd.n2795 0.152939
R13173 gnd.n2826 gnd.n2795 0.152939
R13174 gnd.n2827 gnd.n2826 0.152939
R13175 gnd.n2828 gnd.n2827 0.152939
R13176 gnd.n2828 gnd.n2793 0.152939
R13177 gnd.n2836 gnd.n2793 0.152939
R13178 gnd.n3775 gnd.n2380 0.152939
R13179 gnd.n2382 gnd.n2380 0.152939
R13180 gnd.n2383 gnd.n2382 0.152939
R13181 gnd.n2384 gnd.n2383 0.152939
R13182 gnd.n2385 gnd.n2384 0.152939
R13183 gnd.n2386 gnd.n2385 0.152939
R13184 gnd.n2387 gnd.n2386 0.152939
R13185 gnd.n2388 gnd.n2387 0.152939
R13186 gnd.n2389 gnd.n2388 0.152939
R13187 gnd.n2390 gnd.n2389 0.152939
R13188 gnd.n2391 gnd.n2390 0.152939
R13189 gnd.n2392 gnd.n2391 0.152939
R13190 gnd.n2393 gnd.n2392 0.152939
R13191 gnd.n2394 gnd.n2393 0.152939
R13192 gnd.n2395 gnd.n2394 0.152939
R13193 gnd.n2396 gnd.n2395 0.152939
R13194 gnd.n2397 gnd.n2396 0.152939
R13195 gnd.n2398 gnd.n2397 0.152939
R13196 gnd.n2399 gnd.n2398 0.152939
R13197 gnd.n2400 gnd.n2399 0.152939
R13198 gnd.n2401 gnd.n2400 0.152939
R13199 gnd.n2402 gnd.n2401 0.152939
R13200 gnd.n2406 gnd.n2402 0.152939
R13201 gnd.n2407 gnd.n2406 0.152939
R13202 gnd.n2408 gnd.n2407 0.152939
R13203 gnd.n2409 gnd.n2408 0.152939
R13204 gnd.n3211 gnd.n3210 0.152939
R13205 gnd.n3212 gnd.n3211 0.152939
R13206 gnd.n3213 gnd.n3212 0.152939
R13207 gnd.n3214 gnd.n3213 0.152939
R13208 gnd.n3215 gnd.n3214 0.152939
R13209 gnd.n3216 gnd.n3215 0.152939
R13210 gnd.n3216 gnd.n2515 0.152939
R13211 gnd.n3295 gnd.n2515 0.152939
R13212 gnd.n3296 gnd.n3295 0.152939
R13213 gnd.n3297 gnd.n3296 0.152939
R13214 gnd.n3298 gnd.n3297 0.152939
R13215 gnd.n3299 gnd.n3298 0.152939
R13216 gnd.n3300 gnd.n3299 0.152939
R13217 gnd.n3301 gnd.n3300 0.152939
R13218 gnd.n3302 gnd.n3301 0.152939
R13219 gnd.n3303 gnd.n3302 0.152939
R13220 gnd.n3303 gnd.n2459 0.152939
R13221 gnd.n3380 gnd.n2459 0.152939
R13222 gnd.n3381 gnd.n3380 0.152939
R13223 gnd.n3382 gnd.n3381 0.152939
R13224 gnd.n3383 gnd.n3382 0.152939
R13225 gnd.n3384 gnd.n3383 0.152939
R13226 gnd.n3385 gnd.n3384 0.152939
R13227 gnd.n3386 gnd.n3385 0.152939
R13228 gnd.n3387 gnd.n3386 0.152939
R13229 gnd.n3388 gnd.n3387 0.152939
R13230 gnd.n3390 gnd.n3388 0.152939
R13231 gnd.n3390 gnd.n3389 0.152939
R13232 gnd.n2966 gnd.n2965 0.152939
R13233 gnd.n2966 gnd.n2856 0.152939
R13234 gnd.n2981 gnd.n2856 0.152939
R13235 gnd.n2982 gnd.n2981 0.152939
R13236 gnd.n2983 gnd.n2982 0.152939
R13237 gnd.n2983 gnd.n2844 0.152939
R13238 gnd.n2997 gnd.n2844 0.152939
R13239 gnd.n2998 gnd.n2997 0.152939
R13240 gnd.n2999 gnd.n2998 0.152939
R13241 gnd.n3000 gnd.n2999 0.152939
R13242 gnd.n3001 gnd.n3000 0.152939
R13243 gnd.n3002 gnd.n3001 0.152939
R13244 gnd.n3003 gnd.n3002 0.152939
R13245 gnd.n3004 gnd.n3003 0.152939
R13246 gnd.n3005 gnd.n3004 0.152939
R13247 gnd.n3006 gnd.n3005 0.152939
R13248 gnd.n3007 gnd.n3006 0.152939
R13249 gnd.n3008 gnd.n3007 0.152939
R13250 gnd.n3009 gnd.n3008 0.152939
R13251 gnd.n3010 gnd.n3009 0.152939
R13252 gnd.n3011 gnd.n3010 0.152939
R13253 gnd.n3011 gnd.n2710 0.152939
R13254 gnd.n3128 gnd.n2710 0.152939
R13255 gnd.n3129 gnd.n3128 0.152939
R13256 gnd.n3130 gnd.n3129 0.152939
R13257 gnd.n3131 gnd.n3130 0.152939
R13258 gnd.n3131 gnd.n2632 0.152939
R13259 gnd.n3208 gnd.n2632 0.152939
R13260 gnd.n2884 gnd.n2883 0.152939
R13261 gnd.n2885 gnd.n2884 0.152939
R13262 gnd.n2886 gnd.n2885 0.152939
R13263 gnd.n2887 gnd.n2886 0.152939
R13264 gnd.n2888 gnd.n2887 0.152939
R13265 gnd.n2889 gnd.n2888 0.152939
R13266 gnd.n2890 gnd.n2889 0.152939
R13267 gnd.n2891 gnd.n2890 0.152939
R13268 gnd.n2892 gnd.n2891 0.152939
R13269 gnd.n2893 gnd.n2892 0.152939
R13270 gnd.n2894 gnd.n2893 0.152939
R13271 gnd.n2895 gnd.n2894 0.152939
R13272 gnd.n2896 gnd.n2895 0.152939
R13273 gnd.n2897 gnd.n2896 0.152939
R13274 gnd.n2898 gnd.n2897 0.152939
R13275 gnd.n2899 gnd.n2898 0.152939
R13276 gnd.n2900 gnd.n2899 0.152939
R13277 gnd.n2901 gnd.n2900 0.152939
R13278 gnd.n2902 gnd.n2901 0.152939
R13279 gnd.n2903 gnd.n2902 0.152939
R13280 gnd.n2904 gnd.n2903 0.152939
R13281 gnd.n2905 gnd.n2904 0.152939
R13282 gnd.n2909 gnd.n2905 0.152939
R13283 gnd.n2910 gnd.n2909 0.152939
R13284 gnd.n2910 gnd.n2867 0.152939
R13285 gnd.n2964 gnd.n2867 0.152939
R13286 gnd.n6579 gnd.n794 0.152939
R13287 gnd.n6587 gnd.n794 0.152939
R13288 gnd.n6588 gnd.n6587 0.152939
R13289 gnd.n6589 gnd.n6588 0.152939
R13290 gnd.n6589 gnd.n788 0.152939
R13291 gnd.n6597 gnd.n788 0.152939
R13292 gnd.n6598 gnd.n6597 0.152939
R13293 gnd.n6599 gnd.n6598 0.152939
R13294 gnd.n6599 gnd.n782 0.152939
R13295 gnd.n6607 gnd.n782 0.152939
R13296 gnd.n6608 gnd.n6607 0.152939
R13297 gnd.n6609 gnd.n6608 0.152939
R13298 gnd.n6609 gnd.n776 0.152939
R13299 gnd.n6617 gnd.n776 0.152939
R13300 gnd.n6618 gnd.n6617 0.152939
R13301 gnd.n6619 gnd.n6618 0.152939
R13302 gnd.n6619 gnd.n770 0.152939
R13303 gnd.n6627 gnd.n770 0.152939
R13304 gnd.n6628 gnd.n6627 0.152939
R13305 gnd.n6629 gnd.n6628 0.152939
R13306 gnd.n6629 gnd.n764 0.152939
R13307 gnd.n6637 gnd.n764 0.152939
R13308 gnd.n6638 gnd.n6637 0.152939
R13309 gnd.n6639 gnd.n6638 0.152939
R13310 gnd.n6639 gnd.n758 0.152939
R13311 gnd.n6647 gnd.n758 0.152939
R13312 gnd.n6648 gnd.n6647 0.152939
R13313 gnd.n6649 gnd.n6648 0.152939
R13314 gnd.n6649 gnd.n752 0.152939
R13315 gnd.n6657 gnd.n752 0.152939
R13316 gnd.n6658 gnd.n6657 0.152939
R13317 gnd.n6659 gnd.n6658 0.152939
R13318 gnd.n6659 gnd.n746 0.152939
R13319 gnd.n6667 gnd.n746 0.152939
R13320 gnd.n6668 gnd.n6667 0.152939
R13321 gnd.n6669 gnd.n6668 0.152939
R13322 gnd.n6669 gnd.n740 0.152939
R13323 gnd.n6677 gnd.n740 0.152939
R13324 gnd.n6678 gnd.n6677 0.152939
R13325 gnd.n6679 gnd.n6678 0.152939
R13326 gnd.n6679 gnd.n734 0.152939
R13327 gnd.n6687 gnd.n734 0.152939
R13328 gnd.n6688 gnd.n6687 0.152939
R13329 gnd.n6689 gnd.n6688 0.152939
R13330 gnd.n6689 gnd.n728 0.152939
R13331 gnd.n6697 gnd.n728 0.152939
R13332 gnd.n6698 gnd.n6697 0.152939
R13333 gnd.n6699 gnd.n6698 0.152939
R13334 gnd.n6699 gnd.n722 0.152939
R13335 gnd.n6707 gnd.n722 0.152939
R13336 gnd.n6708 gnd.n6707 0.152939
R13337 gnd.n6709 gnd.n6708 0.152939
R13338 gnd.n6709 gnd.n716 0.152939
R13339 gnd.n6717 gnd.n716 0.152939
R13340 gnd.n6718 gnd.n6717 0.152939
R13341 gnd.n6719 gnd.n6718 0.152939
R13342 gnd.n6719 gnd.n710 0.152939
R13343 gnd.n6727 gnd.n710 0.152939
R13344 gnd.n6728 gnd.n6727 0.152939
R13345 gnd.n6729 gnd.n6728 0.152939
R13346 gnd.n6729 gnd.n704 0.152939
R13347 gnd.n6737 gnd.n704 0.152939
R13348 gnd.n6738 gnd.n6737 0.152939
R13349 gnd.n6739 gnd.n6738 0.152939
R13350 gnd.n6739 gnd.n698 0.152939
R13351 gnd.n6747 gnd.n698 0.152939
R13352 gnd.n6748 gnd.n6747 0.152939
R13353 gnd.n6749 gnd.n6748 0.152939
R13354 gnd.n6749 gnd.n692 0.152939
R13355 gnd.n6757 gnd.n692 0.152939
R13356 gnd.n6758 gnd.n6757 0.152939
R13357 gnd.n6759 gnd.n6758 0.152939
R13358 gnd.n6759 gnd.n686 0.152939
R13359 gnd.n6767 gnd.n686 0.152939
R13360 gnd.n6768 gnd.n6767 0.152939
R13361 gnd.n6769 gnd.n6768 0.152939
R13362 gnd.n6769 gnd.n680 0.152939
R13363 gnd.n6777 gnd.n680 0.152939
R13364 gnd.n6778 gnd.n6777 0.152939
R13365 gnd.n6779 gnd.n6778 0.152939
R13366 gnd.n6779 gnd.n674 0.152939
R13367 gnd.n6787 gnd.n674 0.152939
R13368 gnd.n6788 gnd.n6787 0.152939
R13369 gnd.n6789 gnd.n6788 0.152939
R13370 gnd.n6789 gnd.n668 0.152939
R13371 gnd.n6797 gnd.n668 0.152939
R13372 gnd.n6798 gnd.n6797 0.152939
R13373 gnd.n6799 gnd.n6798 0.152939
R13374 gnd.n6799 gnd.n662 0.152939
R13375 gnd.n6807 gnd.n662 0.152939
R13376 gnd.n6808 gnd.n6807 0.152939
R13377 gnd.n6809 gnd.n6808 0.152939
R13378 gnd.n6809 gnd.n656 0.152939
R13379 gnd.n6817 gnd.n656 0.152939
R13380 gnd.n6818 gnd.n6817 0.152939
R13381 gnd.n6819 gnd.n6818 0.152939
R13382 gnd.n6819 gnd.n650 0.152939
R13383 gnd.n6827 gnd.n650 0.152939
R13384 gnd.n6828 gnd.n6827 0.152939
R13385 gnd.n6829 gnd.n6828 0.152939
R13386 gnd.n6829 gnd.n644 0.152939
R13387 gnd.n6837 gnd.n644 0.152939
R13388 gnd.n6838 gnd.n6837 0.152939
R13389 gnd.n6839 gnd.n6838 0.152939
R13390 gnd.n6839 gnd.n638 0.152939
R13391 gnd.n6847 gnd.n638 0.152939
R13392 gnd.n6848 gnd.n6847 0.152939
R13393 gnd.n6849 gnd.n6848 0.152939
R13394 gnd.n6849 gnd.n632 0.152939
R13395 gnd.n6857 gnd.n632 0.152939
R13396 gnd.n6858 gnd.n6857 0.152939
R13397 gnd.n6859 gnd.n6858 0.152939
R13398 gnd.n6859 gnd.n626 0.152939
R13399 gnd.n6867 gnd.n626 0.152939
R13400 gnd.n6868 gnd.n6867 0.152939
R13401 gnd.n6869 gnd.n6868 0.152939
R13402 gnd.n6869 gnd.n620 0.152939
R13403 gnd.n6877 gnd.n620 0.152939
R13404 gnd.n6878 gnd.n6877 0.152939
R13405 gnd.n6879 gnd.n6878 0.152939
R13406 gnd.n6879 gnd.n614 0.152939
R13407 gnd.n6887 gnd.n614 0.152939
R13408 gnd.n6888 gnd.n6887 0.152939
R13409 gnd.n6889 gnd.n6888 0.152939
R13410 gnd.n6889 gnd.n608 0.152939
R13411 gnd.n6897 gnd.n608 0.152939
R13412 gnd.n6898 gnd.n6897 0.152939
R13413 gnd.n6899 gnd.n6898 0.152939
R13414 gnd.n6899 gnd.n602 0.152939
R13415 gnd.n6907 gnd.n602 0.152939
R13416 gnd.n6908 gnd.n6907 0.152939
R13417 gnd.n6909 gnd.n6908 0.152939
R13418 gnd.n6909 gnd.n596 0.152939
R13419 gnd.n6917 gnd.n596 0.152939
R13420 gnd.n6918 gnd.n6917 0.152939
R13421 gnd.n6919 gnd.n6918 0.152939
R13422 gnd.n6919 gnd.n590 0.152939
R13423 gnd.n6927 gnd.n590 0.152939
R13424 gnd.n6928 gnd.n6927 0.152939
R13425 gnd.n6929 gnd.n6928 0.152939
R13426 gnd.n6929 gnd.n584 0.152939
R13427 gnd.n6937 gnd.n584 0.152939
R13428 gnd.n6938 gnd.n6937 0.152939
R13429 gnd.n6939 gnd.n6938 0.152939
R13430 gnd.n6939 gnd.n578 0.152939
R13431 gnd.n6947 gnd.n578 0.152939
R13432 gnd.n6948 gnd.n6947 0.152939
R13433 gnd.n6949 gnd.n6948 0.152939
R13434 gnd.n6949 gnd.n572 0.152939
R13435 gnd.n6957 gnd.n572 0.152939
R13436 gnd.n6958 gnd.n6957 0.152939
R13437 gnd.n6959 gnd.n6958 0.152939
R13438 gnd.n6959 gnd.n566 0.152939
R13439 gnd.n6967 gnd.n566 0.152939
R13440 gnd.n6968 gnd.n6967 0.152939
R13441 gnd.n6969 gnd.n6968 0.152939
R13442 gnd.n6969 gnd.n560 0.152939
R13443 gnd.n6977 gnd.n560 0.152939
R13444 gnd.n6978 gnd.n6977 0.152939
R13445 gnd.n6979 gnd.n6978 0.152939
R13446 gnd.n6979 gnd.n554 0.152939
R13447 gnd.n6987 gnd.n554 0.152939
R13448 gnd.n6988 gnd.n6987 0.152939
R13449 gnd.n6990 gnd.n6988 0.152939
R13450 gnd.n6990 gnd.n6989 0.152939
R13451 gnd.n6989 gnd.n548 0.152939
R13452 gnd.n6999 gnd.n548 0.152939
R13453 gnd.n7000 gnd.n543 0.152939
R13454 gnd.n7008 gnd.n543 0.152939
R13455 gnd.n7009 gnd.n7008 0.152939
R13456 gnd.n7010 gnd.n7009 0.152939
R13457 gnd.n7010 gnd.n537 0.152939
R13458 gnd.n7018 gnd.n537 0.152939
R13459 gnd.n7019 gnd.n7018 0.152939
R13460 gnd.n7020 gnd.n7019 0.152939
R13461 gnd.n7020 gnd.n531 0.152939
R13462 gnd.n7028 gnd.n531 0.152939
R13463 gnd.n7029 gnd.n7028 0.152939
R13464 gnd.n7030 gnd.n7029 0.152939
R13465 gnd.n7030 gnd.n525 0.152939
R13466 gnd.n7038 gnd.n525 0.152939
R13467 gnd.n7039 gnd.n7038 0.152939
R13468 gnd.n7040 gnd.n7039 0.152939
R13469 gnd.n7040 gnd.n519 0.152939
R13470 gnd.n7048 gnd.n519 0.152939
R13471 gnd.n7049 gnd.n7048 0.152939
R13472 gnd.n7050 gnd.n7049 0.152939
R13473 gnd.n7050 gnd.n513 0.152939
R13474 gnd.n7058 gnd.n513 0.152939
R13475 gnd.n7059 gnd.n7058 0.152939
R13476 gnd.n7060 gnd.n7059 0.152939
R13477 gnd.n7060 gnd.n507 0.152939
R13478 gnd.n7068 gnd.n507 0.152939
R13479 gnd.n7069 gnd.n7068 0.152939
R13480 gnd.n7070 gnd.n7069 0.152939
R13481 gnd.n7070 gnd.n501 0.152939
R13482 gnd.n7078 gnd.n501 0.152939
R13483 gnd.n7079 gnd.n7078 0.152939
R13484 gnd.n7080 gnd.n7079 0.152939
R13485 gnd.n7080 gnd.n495 0.152939
R13486 gnd.n7088 gnd.n495 0.152939
R13487 gnd.n7089 gnd.n7088 0.152939
R13488 gnd.n7090 gnd.n7089 0.152939
R13489 gnd.n7090 gnd.n489 0.152939
R13490 gnd.n7098 gnd.n489 0.152939
R13491 gnd.n7099 gnd.n7098 0.152939
R13492 gnd.n7100 gnd.n7099 0.152939
R13493 gnd.n7100 gnd.n483 0.152939
R13494 gnd.n7108 gnd.n483 0.152939
R13495 gnd.n7109 gnd.n7108 0.152939
R13496 gnd.n7110 gnd.n7109 0.152939
R13497 gnd.n7110 gnd.n477 0.152939
R13498 gnd.n7118 gnd.n477 0.152939
R13499 gnd.n7119 gnd.n7118 0.152939
R13500 gnd.n7120 gnd.n7119 0.152939
R13501 gnd.n7120 gnd.n471 0.152939
R13502 gnd.n7128 gnd.n471 0.152939
R13503 gnd.n7129 gnd.n7128 0.152939
R13504 gnd.n7130 gnd.n7129 0.152939
R13505 gnd.n7130 gnd.n465 0.152939
R13506 gnd.n7138 gnd.n465 0.152939
R13507 gnd.n7139 gnd.n7138 0.152939
R13508 gnd.n7140 gnd.n7139 0.152939
R13509 gnd.n7140 gnd.n459 0.152939
R13510 gnd.n7148 gnd.n459 0.152939
R13511 gnd.n7149 gnd.n7148 0.152939
R13512 gnd.n7150 gnd.n7149 0.152939
R13513 gnd.n7150 gnd.n453 0.152939
R13514 gnd.n7158 gnd.n453 0.152939
R13515 gnd.n7159 gnd.n7158 0.152939
R13516 gnd.n7160 gnd.n7159 0.152939
R13517 gnd.n7160 gnd.n447 0.152939
R13518 gnd.n7168 gnd.n447 0.152939
R13519 gnd.n7169 gnd.n7168 0.152939
R13520 gnd.n7170 gnd.n7169 0.152939
R13521 gnd.n7170 gnd.n441 0.152939
R13522 gnd.n7178 gnd.n441 0.152939
R13523 gnd.n7179 gnd.n7178 0.152939
R13524 gnd.n7180 gnd.n7179 0.152939
R13525 gnd.n7180 gnd.n435 0.152939
R13526 gnd.n7188 gnd.n435 0.152939
R13527 gnd.n7189 gnd.n7188 0.152939
R13528 gnd.n7190 gnd.n7189 0.152939
R13529 gnd.n7190 gnd.n429 0.152939
R13530 gnd.n7198 gnd.n429 0.152939
R13531 gnd.n7199 gnd.n7198 0.152939
R13532 gnd.n7200 gnd.n7199 0.152939
R13533 gnd.n7200 gnd.n423 0.152939
R13534 gnd.n7209 gnd.n423 0.152939
R13535 gnd.n7210 gnd.n7209 0.152939
R13536 gnd.n7211 gnd.n7210 0.152939
R13537 gnd.n7418 gnd.n7417 0.152939
R13538 gnd.n7418 gnd.n287 0.152939
R13539 gnd.n7432 gnd.n287 0.152939
R13540 gnd.n7433 gnd.n7432 0.152939
R13541 gnd.n7434 gnd.n7433 0.152939
R13542 gnd.n7434 gnd.n273 0.152939
R13543 gnd.n7448 gnd.n273 0.152939
R13544 gnd.n7449 gnd.n7448 0.152939
R13545 gnd.n7450 gnd.n7449 0.152939
R13546 gnd.n7450 gnd.n257 0.152939
R13547 gnd.n7464 gnd.n257 0.152939
R13548 gnd.n7465 gnd.n7464 0.152939
R13549 gnd.n7466 gnd.n7465 0.152939
R13550 gnd.n7466 gnd.n242 0.152939
R13551 gnd.n7480 gnd.n242 0.152939
R13552 gnd.n7481 gnd.n7480 0.152939
R13553 gnd.n7482 gnd.n7481 0.152939
R13554 gnd.n7482 gnd.n226 0.152939
R13555 gnd.n7496 gnd.n226 0.152939
R13556 gnd.n7497 gnd.n7496 0.152939
R13557 gnd.n7498 gnd.n7497 0.152939
R13558 gnd.n7498 gnd.n210 0.152939
R13559 gnd.n7580 gnd.n210 0.152939
R13560 gnd.n7581 gnd.n7580 0.152939
R13561 gnd.n7582 gnd.n7581 0.152939
R13562 gnd.n7582 gnd.n133 0.152939
R13563 gnd.n7662 gnd.n133 0.152939
R13564 gnd.n7661 gnd.n134 0.152939
R13565 gnd.n136 gnd.n134 0.152939
R13566 gnd.n140 gnd.n136 0.152939
R13567 gnd.n141 gnd.n140 0.152939
R13568 gnd.n142 gnd.n141 0.152939
R13569 gnd.n143 gnd.n142 0.152939
R13570 gnd.n147 gnd.n143 0.152939
R13571 gnd.n148 gnd.n147 0.152939
R13572 gnd.n149 gnd.n148 0.152939
R13573 gnd.n150 gnd.n149 0.152939
R13574 gnd.n154 gnd.n150 0.152939
R13575 gnd.n155 gnd.n154 0.152939
R13576 gnd.n156 gnd.n155 0.152939
R13577 gnd.n157 gnd.n156 0.152939
R13578 gnd.n161 gnd.n157 0.152939
R13579 gnd.n162 gnd.n161 0.152939
R13580 gnd.n163 gnd.n162 0.152939
R13581 gnd.n164 gnd.n163 0.152939
R13582 gnd.n168 gnd.n164 0.152939
R13583 gnd.n169 gnd.n168 0.152939
R13584 gnd.n170 gnd.n169 0.152939
R13585 gnd.n171 gnd.n170 0.152939
R13586 gnd.n175 gnd.n171 0.152939
R13587 gnd.n176 gnd.n175 0.152939
R13588 gnd.n177 gnd.n176 0.152939
R13589 gnd.n178 gnd.n177 0.152939
R13590 gnd.n182 gnd.n178 0.152939
R13591 gnd.n183 gnd.n182 0.152939
R13592 gnd.n184 gnd.n183 0.152939
R13593 gnd.n185 gnd.n184 0.152939
R13594 gnd.n189 gnd.n185 0.152939
R13595 gnd.n190 gnd.n189 0.152939
R13596 gnd.n191 gnd.n190 0.152939
R13597 gnd.n192 gnd.n191 0.152939
R13598 gnd.n196 gnd.n192 0.152939
R13599 gnd.n197 gnd.n196 0.152939
R13600 gnd.n7592 gnd.n197 0.152939
R13601 gnd.n7592 gnd.n7591 0.152939
R13602 gnd.n1456 gnd.n1333 0.152939
R13603 gnd.n1457 gnd.n1456 0.152939
R13604 gnd.n1458 gnd.n1457 0.152939
R13605 gnd.n1459 gnd.n1458 0.152939
R13606 gnd.n1460 gnd.n1459 0.152939
R13607 gnd.n1461 gnd.n1460 0.152939
R13608 gnd.n1462 gnd.n1461 0.152939
R13609 gnd.n1463 gnd.n1462 0.152939
R13610 gnd.n1464 gnd.n1463 0.152939
R13611 gnd.n1464 gnd.n1390 0.152939
R13612 gnd.n5985 gnd.n1390 0.152939
R13613 gnd.n5986 gnd.n5985 0.152939
R13614 gnd.n5987 gnd.n5986 0.152939
R13615 gnd.n5987 gnd.n1388 0.152939
R13616 gnd.n5992 gnd.n1388 0.152939
R13617 gnd.n5993 gnd.n5992 0.152939
R13618 gnd.n5994 gnd.n5993 0.152939
R13619 gnd.n5995 gnd.n5994 0.152939
R13620 gnd.n5995 gnd.n387 0.152939
R13621 gnd.n7248 gnd.n387 0.152939
R13622 gnd.n7249 gnd.n7248 0.152939
R13623 gnd.n7250 gnd.n7249 0.152939
R13624 gnd.n7251 gnd.n7250 0.152939
R13625 gnd.n7252 gnd.n7251 0.152939
R13626 gnd.n7252 gnd.n353 0.152939
R13627 gnd.n7293 gnd.n353 0.152939
R13628 gnd.n7294 gnd.n7293 0.152939
R13629 gnd.n7295 gnd.n7294 0.152939
R13630 gnd.n7296 gnd.n7295 0.152939
R13631 gnd.n7297 gnd.n7296 0.152939
R13632 gnd.n7298 gnd.n7297 0.152939
R13633 gnd.n7298 gnd.n337 0.152939
R13634 gnd.n7323 gnd.n337 0.152939
R13635 gnd.n7324 gnd.n7323 0.152939
R13636 gnd.n7325 gnd.n7324 0.152939
R13637 gnd.n7326 gnd.n7325 0.152939
R13638 gnd.n7327 gnd.n7326 0.152939
R13639 gnd.n7328 gnd.n7327 0.152939
R13640 gnd.n7329 gnd.n7328 0.152939
R13641 gnd.n7330 gnd.n7329 0.152939
R13642 gnd.n7331 gnd.n7330 0.152939
R13643 gnd.n7332 gnd.n7331 0.152939
R13644 gnd.n7333 gnd.n7332 0.152939
R13645 gnd.n7334 gnd.n7333 0.152939
R13646 gnd.n7335 gnd.n7334 0.152939
R13647 gnd.n7336 gnd.n7335 0.152939
R13648 gnd.n7337 gnd.n7336 0.152939
R13649 gnd.n7338 gnd.n7337 0.152939
R13650 gnd.n7339 gnd.n7338 0.152939
R13651 gnd.n7340 gnd.n7339 0.152939
R13652 gnd.n7341 gnd.n7340 0.152939
R13653 gnd.n7342 gnd.n7341 0.152939
R13654 gnd.n7343 gnd.n7342 0.152939
R13655 gnd.n7344 gnd.n7343 0.152939
R13656 gnd.n7345 gnd.n7344 0.152939
R13657 gnd.n7346 gnd.n7345 0.152939
R13658 gnd.n7347 gnd.n7346 0.152939
R13659 gnd.n7348 gnd.n7347 0.152939
R13660 gnd.n7349 gnd.n7348 0.152939
R13661 gnd.n7350 gnd.n7349 0.152939
R13662 gnd.n7352 gnd.n7350 0.152939
R13663 gnd.n7352 gnd.n7351 0.152939
R13664 gnd.n7351 gnd.n203 0.152939
R13665 gnd.n7590 gnd.n203 0.152939
R13666 gnd.n1290 gnd.n1289 0.152939
R13667 gnd.n1291 gnd.n1290 0.152939
R13668 gnd.n1292 gnd.n1291 0.152939
R13669 gnd.n1293 gnd.n1292 0.152939
R13670 gnd.n1294 gnd.n1293 0.152939
R13671 gnd.n1295 gnd.n1294 0.152939
R13672 gnd.n1296 gnd.n1295 0.152939
R13673 gnd.n1297 gnd.n1296 0.152939
R13674 gnd.n1298 gnd.n1297 0.152939
R13675 gnd.n1299 gnd.n1298 0.152939
R13676 gnd.n1300 gnd.n1299 0.152939
R13677 gnd.n1301 gnd.n1300 0.152939
R13678 gnd.n1302 gnd.n1301 0.152939
R13679 gnd.n1303 gnd.n1302 0.152939
R13680 gnd.n1304 gnd.n1303 0.152939
R13681 gnd.n1311 gnd.n1310 0.152939
R13682 gnd.n1312 gnd.n1311 0.152939
R13683 gnd.n1313 gnd.n1312 0.152939
R13684 gnd.n1314 gnd.n1313 0.152939
R13685 gnd.n1315 gnd.n1314 0.152939
R13686 gnd.n1316 gnd.n1315 0.152939
R13687 gnd.n1317 gnd.n1316 0.152939
R13688 gnd.n1318 gnd.n1317 0.152939
R13689 gnd.n1319 gnd.n1318 0.152939
R13690 gnd.n1320 gnd.n1319 0.152939
R13691 gnd.n1321 gnd.n1320 0.152939
R13692 gnd.n1322 gnd.n1321 0.152939
R13693 gnd.n1323 gnd.n1322 0.152939
R13694 gnd.n1324 gnd.n1323 0.152939
R13695 gnd.n1325 gnd.n1324 0.152939
R13696 gnd.n1326 gnd.n1325 0.152939
R13697 gnd.n1327 gnd.n1326 0.152939
R13698 gnd.n6085 gnd.n1327 0.152939
R13699 gnd.n6085 gnd.n6084 0.152939
R13700 gnd.n6084 gnd.n6083 0.152939
R13701 gnd.n5909 gnd.n5908 0.152939
R13702 gnd.n5910 gnd.n5909 0.152939
R13703 gnd.n5910 gnd.n1428 0.152939
R13704 gnd.n5938 gnd.n1428 0.152939
R13705 gnd.n5939 gnd.n5938 0.152939
R13706 gnd.n5940 gnd.n5939 0.152939
R13707 gnd.n5941 gnd.n5940 0.152939
R13708 gnd.n5941 gnd.n1401 0.152939
R13709 gnd.n5975 gnd.n1401 0.152939
R13710 gnd.n5976 gnd.n5975 0.152939
R13711 gnd.n5977 gnd.n5976 0.152939
R13712 gnd.n5978 gnd.n5977 0.152939
R13713 gnd.n5978 gnd.n1367 0.152939
R13714 gnd.n6045 gnd.n1367 0.152939
R13715 gnd.n6046 gnd.n6045 0.152939
R13716 gnd.n6047 gnd.n6046 0.152939
R13717 gnd.n6047 gnd.n396 0.152939
R13718 gnd.n7238 gnd.n396 0.152939
R13719 gnd.n7239 gnd.n7238 0.152939
R13720 gnd.n7240 gnd.n7239 0.152939
R13721 gnd.n7241 gnd.n7240 0.152939
R13722 gnd.n7241 gnd.n363 0.152939
R13723 gnd.n7284 gnd.n363 0.152939
R13724 gnd.n7285 gnd.n7284 0.152939
R13725 gnd.n7286 gnd.n7285 0.152939
R13726 gnd.n7286 gnd.n303 0.152939
R13727 gnd.n7417 gnd.n303 0.152939
R13728 gnd.n6406 gnd.n967 0.152939
R13729 gnd.n4376 gnd.n967 0.152939
R13730 gnd.n4377 gnd.n4376 0.152939
R13731 gnd.n4378 gnd.n4377 0.152939
R13732 gnd.n4378 gnd.n2169 0.152939
R13733 gnd.n4417 gnd.n2169 0.152939
R13734 gnd.n4418 gnd.n4417 0.152939
R13735 gnd.n4419 gnd.n4418 0.152939
R13736 gnd.n4419 gnd.n2165 0.152939
R13737 gnd.n4425 gnd.n2165 0.152939
R13738 gnd.n4426 gnd.n4425 0.152939
R13739 gnd.n4427 gnd.n4426 0.152939
R13740 gnd.n4427 gnd.n2148 0.152939
R13741 gnd.n4466 gnd.n2148 0.152939
R13742 gnd.n4467 gnd.n4466 0.152939
R13743 gnd.n4468 gnd.n4467 0.152939
R13744 gnd.n4468 gnd.n2144 0.152939
R13745 gnd.n4474 gnd.n2144 0.152939
R13746 gnd.n4475 gnd.n4474 0.152939
R13747 gnd.n4476 gnd.n4475 0.152939
R13748 gnd.n4477 gnd.n4476 0.152939
R13749 gnd.n4478 gnd.n4477 0.152939
R13750 gnd.n4481 gnd.n4478 0.152939
R13751 gnd.n4482 gnd.n4481 0.152939
R13752 gnd.n4483 gnd.n4482 0.152939
R13753 gnd.n4484 gnd.n4483 0.152939
R13754 gnd.n4487 gnd.n4484 0.152939
R13755 gnd.n4488 gnd.n4487 0.152939
R13756 gnd.n4489 gnd.n4488 0.152939
R13757 gnd.n4490 gnd.n4489 0.152939
R13758 gnd.n4491 gnd.n4490 0.152939
R13759 gnd.n4491 gnd.n1970 0.152939
R13760 gnd.n4909 gnd.n1970 0.152939
R13761 gnd.n4910 gnd.n4909 0.152939
R13762 gnd.n4911 gnd.n4910 0.152939
R13763 gnd.n4911 gnd.n1958 0.152939
R13764 gnd.n4925 gnd.n1958 0.152939
R13765 gnd.n4926 gnd.n4925 0.152939
R13766 gnd.n4927 gnd.n4926 0.152939
R13767 gnd.n4927 gnd.n1945 0.152939
R13768 gnd.n4941 gnd.n1945 0.152939
R13769 gnd.n4942 gnd.n4941 0.152939
R13770 gnd.n4943 gnd.n4942 0.152939
R13771 gnd.n4943 gnd.n1932 0.152939
R13772 gnd.n4957 gnd.n1932 0.152939
R13773 gnd.n4958 gnd.n4957 0.152939
R13774 gnd.n4959 gnd.n4958 0.152939
R13775 gnd.n4959 gnd.n1919 0.152939
R13776 gnd.n4973 gnd.n1919 0.152939
R13777 gnd.n4974 gnd.n4973 0.152939
R13778 gnd.n4975 gnd.n4974 0.152939
R13779 gnd.n4975 gnd.n1905 0.152939
R13780 gnd.n4989 gnd.n1905 0.152939
R13781 gnd.n4990 gnd.n4989 0.152939
R13782 gnd.n4991 gnd.n4990 0.152939
R13783 gnd.n4992 gnd.n4991 0.152939
R13784 gnd.n4992 gnd.n1874 0.152939
R13785 gnd.n5575 gnd.n1874 0.152939
R13786 gnd.n5576 gnd.n5575 0.152939
R13787 gnd.n5577 gnd.n5576 0.152939
R13788 gnd.n5577 gnd.n1860 0.152939
R13789 gnd.n5591 gnd.n1860 0.152939
R13790 gnd.n5592 gnd.n5591 0.152939
R13791 gnd.n5593 gnd.n5592 0.152939
R13792 gnd.n5593 gnd.n1845 0.152939
R13793 gnd.n5607 gnd.n1845 0.152939
R13794 gnd.n5608 gnd.n5607 0.152939
R13795 gnd.n5609 gnd.n5608 0.152939
R13796 gnd.n5609 gnd.n1830 0.152939
R13797 gnd.n5623 gnd.n1830 0.152939
R13798 gnd.n5624 gnd.n5623 0.152939
R13799 gnd.n5625 gnd.n5624 0.152939
R13800 gnd.n5625 gnd.n1816 0.152939
R13801 gnd.n5639 gnd.n1816 0.152939
R13802 gnd.n5640 gnd.n5639 0.152939
R13803 gnd.n5641 gnd.n5640 0.152939
R13804 gnd.n5641 gnd.n1801 0.152939
R13805 gnd.n5655 gnd.n1801 0.152939
R13806 gnd.n5656 gnd.n5655 0.152939
R13807 gnd.n5657 gnd.n5656 0.152939
R13808 gnd.n5657 gnd.n1786 0.152939
R13809 gnd.n5671 gnd.n1786 0.152939
R13810 gnd.n5672 gnd.n5671 0.152939
R13811 gnd.n5673 gnd.n5672 0.152939
R13812 gnd.n5673 gnd.n1771 0.152939
R13813 gnd.n5687 gnd.n1771 0.152939
R13814 gnd.n5688 gnd.n5687 0.152939
R13815 gnd.n5689 gnd.n5688 0.152939
R13816 gnd.n5689 gnd.n1757 0.152939
R13817 gnd.n5703 gnd.n1757 0.152939
R13818 gnd.n5704 gnd.n5703 0.152939
R13819 gnd.n5705 gnd.n5704 0.152939
R13820 gnd.n5705 gnd.n1742 0.152939
R13821 gnd.n5719 gnd.n1742 0.152939
R13822 gnd.n5720 gnd.n5719 0.152939
R13823 gnd.n5721 gnd.n5720 0.152939
R13824 gnd.n5721 gnd.n1729 0.152939
R13825 gnd.n5735 gnd.n1729 0.152939
R13826 gnd.n5736 gnd.n5735 0.152939
R13827 gnd.n5737 gnd.n5736 0.152939
R13828 gnd.n5737 gnd.n1717 0.152939
R13829 gnd.n5751 gnd.n1717 0.152939
R13830 gnd.n5752 gnd.n5751 0.152939
R13831 gnd.n5753 gnd.n5752 0.152939
R13832 gnd.n5753 gnd.n1703 0.152939
R13833 gnd.n5767 gnd.n1703 0.152939
R13834 gnd.n5768 gnd.n5767 0.152939
R13835 gnd.n5769 gnd.n5768 0.152939
R13836 gnd.n5769 gnd.n1690 0.152939
R13837 gnd.n5783 gnd.n1690 0.152939
R13838 gnd.n5784 gnd.n5783 0.152939
R13839 gnd.n5785 gnd.n5784 0.152939
R13840 gnd.n5785 gnd.n1676 0.152939
R13841 gnd.n5799 gnd.n1676 0.152939
R13842 gnd.n5800 gnd.n5799 0.152939
R13843 gnd.n5801 gnd.n5800 0.152939
R13844 gnd.n5801 gnd.n1663 0.152939
R13845 gnd.n5815 gnd.n1663 0.152939
R13846 gnd.n5816 gnd.n5815 0.152939
R13847 gnd.n5817 gnd.n5816 0.152939
R13848 gnd.n5817 gnd.n1650 0.152939
R13849 gnd.n5831 gnd.n1650 0.152939
R13850 gnd.n5832 gnd.n5831 0.152939
R13851 gnd.n5833 gnd.n5832 0.152939
R13852 gnd.n5833 gnd.n1636 0.152939
R13853 gnd.n5847 gnd.n1636 0.152939
R13854 gnd.n5848 gnd.n5847 0.152939
R13855 gnd.n5849 gnd.n5848 0.152939
R13856 gnd.n5849 gnd.n1623 0.152939
R13857 gnd.n5865 gnd.n1623 0.152939
R13858 gnd.n5866 gnd.n5865 0.152939
R13859 gnd.n5867 gnd.n5866 0.152939
R13860 gnd.n5869 gnd.n5867 0.152939
R13861 gnd.n5869 gnd.n5868 0.152939
R13862 gnd.n5868 gnd.n1251 0.152939
R13863 gnd.n1252 gnd.n1251 0.152939
R13864 gnd.n1253 gnd.n1252 0.152939
R13865 gnd.n1443 gnd.n1253 0.152939
R13866 gnd.n1446 gnd.n1443 0.152939
R13867 gnd.n1447 gnd.n1446 0.152939
R13868 gnd.n1448 gnd.n1447 0.152939
R13869 gnd.n1448 gnd.n1439 0.152939
R13870 gnd.n5927 gnd.n1439 0.152939
R13871 gnd.n5928 gnd.n5927 0.152939
R13872 gnd.n5929 gnd.n5928 0.152939
R13873 gnd.n5930 gnd.n5929 0.152939
R13874 gnd.n5930 gnd.n1411 0.152939
R13875 gnd.n5963 gnd.n1411 0.152939
R13876 gnd.n5964 gnd.n5963 0.152939
R13877 gnd.n5965 gnd.n5964 0.152939
R13878 gnd.n5966 gnd.n5965 0.152939
R13879 gnd.n5966 gnd.n1377 0.152939
R13880 gnd.n6024 gnd.n1377 0.152939
R13881 gnd.n6025 gnd.n6024 0.152939
R13882 gnd.n6026 gnd.n6025 0.152939
R13883 gnd.n6027 gnd.n6026 0.152939
R13884 gnd.n6028 gnd.n6027 0.152939
R13885 gnd.n6030 gnd.n6028 0.152939
R13886 gnd.n6032 gnd.n6030 0.152939
R13887 gnd.n6032 gnd.n6031 0.152939
R13888 gnd.n6031 gnd.n412 0.152939
R13889 gnd.n413 gnd.n412 0.152939
R13890 gnd.n414 gnd.n413 0.152939
R13891 gnd.n417 gnd.n414 0.152939
R13892 gnd.n418 gnd.n417 0.152939
R13893 gnd.n419 gnd.n418 0.152939
R13894 gnd.n420 gnd.n419 0.152939
R13895 gnd.n3884 gnd.n3883 0.152939
R13896 gnd.n3885 gnd.n3884 0.152939
R13897 gnd.n3886 gnd.n3885 0.152939
R13898 gnd.n3887 gnd.n3886 0.152939
R13899 gnd.n3888 gnd.n3887 0.152939
R13900 gnd.n3889 gnd.n3888 0.152939
R13901 gnd.n3890 gnd.n3889 0.152939
R13902 gnd.n3891 gnd.n3890 0.152939
R13903 gnd.n3892 gnd.n3891 0.152939
R13904 gnd.n3893 gnd.n3892 0.152939
R13905 gnd.n3894 gnd.n3893 0.152939
R13906 gnd.n3895 gnd.n3894 0.152939
R13907 gnd.n3896 gnd.n3895 0.152939
R13908 gnd.n3897 gnd.n3896 0.152939
R13909 gnd.n3898 gnd.n3897 0.152939
R13910 gnd.n3899 gnd.n3898 0.152939
R13911 gnd.n3900 gnd.n3899 0.152939
R13912 gnd.n3901 gnd.n3900 0.152939
R13913 gnd.n3902 gnd.n3901 0.152939
R13914 gnd.n3903 gnd.n3902 0.152939
R13915 gnd.n3904 gnd.n3903 0.152939
R13916 gnd.n3905 gnd.n3904 0.152939
R13917 gnd.n3906 gnd.n3905 0.152939
R13918 gnd.n3907 gnd.n3906 0.152939
R13919 gnd.n3908 gnd.n3907 0.152939
R13920 gnd.n3909 gnd.n3908 0.152939
R13921 gnd.n3910 gnd.n3909 0.152939
R13922 gnd.n3911 gnd.n3910 0.152939
R13923 gnd.n3912 gnd.n3911 0.152939
R13924 gnd.n3913 gnd.n3912 0.152939
R13925 gnd.n3914 gnd.n3913 0.152939
R13926 gnd.n3835 gnd.n2337 0.152939
R13927 gnd.n3843 gnd.n3835 0.152939
R13928 gnd.n3844 gnd.n3843 0.152939
R13929 gnd.n3845 gnd.n3844 0.152939
R13930 gnd.n3845 gnd.n3831 0.152939
R13931 gnd.n3853 gnd.n3831 0.152939
R13932 gnd.n3854 gnd.n3853 0.152939
R13933 gnd.n3855 gnd.n3854 0.152939
R13934 gnd.n3855 gnd.n3827 0.152939
R13935 gnd.n3863 gnd.n3827 0.152939
R13936 gnd.n3864 gnd.n3863 0.152939
R13937 gnd.n3865 gnd.n3864 0.152939
R13938 gnd.n3865 gnd.n3823 0.152939
R13939 gnd.n3873 gnd.n3823 0.152939
R13940 gnd.n3874 gnd.n3873 0.152939
R13941 gnd.n3875 gnd.n3874 0.152939
R13942 gnd.n3875 gnd.n3817 0.152939
R13943 gnd.n3882 gnd.n3817 0.152939
R13944 gnd.n4203 gnd.n4202 0.152939
R13945 gnd.n4204 gnd.n4203 0.152939
R13946 gnd.n4204 gnd.n2322 0.152939
R13947 gnd.n4218 gnd.n2322 0.152939
R13948 gnd.n4219 gnd.n4218 0.152939
R13949 gnd.n4220 gnd.n4219 0.152939
R13950 gnd.n4220 gnd.n2305 0.152939
R13951 gnd.n4234 gnd.n2305 0.152939
R13952 gnd.n4235 gnd.n4234 0.152939
R13953 gnd.n4236 gnd.n4235 0.152939
R13954 gnd.n4236 gnd.n2290 0.152939
R13955 gnd.n4250 gnd.n2290 0.152939
R13956 gnd.n4251 gnd.n4250 0.152939
R13957 gnd.n4252 gnd.n4251 0.152939
R13958 gnd.n4252 gnd.n2273 0.152939
R13959 gnd.n4266 gnd.n2273 0.152939
R13960 gnd.n4267 gnd.n4266 0.152939
R13961 gnd.n4268 gnd.n4267 0.152939
R13962 gnd.n4268 gnd.n2258 0.152939
R13963 gnd.n4282 gnd.n2258 0.152939
R13964 gnd.n4283 gnd.n4282 0.152939
R13965 gnd.n4284 gnd.n4283 0.152939
R13966 gnd.n4284 gnd.n2241 0.152939
R13967 gnd.n4299 gnd.n2241 0.152939
R13968 gnd.n4300 gnd.n4299 0.152939
R13969 gnd.n4301 gnd.n4300 0.152939
R13970 gnd.n4301 gnd.n2227 0.152939
R13971 gnd.n4315 gnd.n2227 0.152939
R13972 gnd.n4316 gnd.n4315 0.152939
R13973 gnd.n4317 gnd.n4316 0.152939
R13974 gnd.n4317 gnd.n2202 0.152939
R13975 gnd.n4333 gnd.n2202 0.152939
R13976 gnd.n4334 gnd.n4333 0.152939
R13977 gnd.n4335 gnd.n4334 0.152939
R13978 gnd.n4336 gnd.n4335 0.152939
R13979 gnd.n4337 gnd.n4336 0.152939
R13980 gnd.n4338 gnd.n4337 0.152939
R13981 gnd.n4340 gnd.n4338 0.152939
R13982 gnd.n4340 gnd.n4339 0.152939
R13983 gnd.n4339 gnd.n990 0.152939
R13984 gnd.n991 gnd.n990 0.152939
R13985 gnd.n992 gnd.n991 0.152939
R13986 gnd.n1009 gnd.n992 0.152939
R13987 gnd.n1010 gnd.n1009 0.152939
R13988 gnd.n1011 gnd.n1010 0.152939
R13989 gnd.n1012 gnd.n1011 0.152939
R13990 gnd.n1031 gnd.n1012 0.152939
R13991 gnd.n1032 gnd.n1031 0.152939
R13992 gnd.n1033 gnd.n1032 0.152939
R13993 gnd.n1034 gnd.n1033 0.152939
R13994 gnd.n1051 gnd.n1034 0.152939
R13995 gnd.n1052 gnd.n1051 0.152939
R13996 gnd.n1053 gnd.n1052 0.152939
R13997 gnd.n1054 gnd.n1053 0.152939
R13998 gnd.n1073 gnd.n1054 0.152939
R13999 gnd.n1074 gnd.n1073 0.152939
R14000 gnd.n1075 gnd.n1074 0.152939
R14001 gnd.n1076 gnd.n1075 0.152939
R14002 gnd.n1094 gnd.n1076 0.152939
R14003 gnd.n1095 gnd.n1094 0.152939
R14004 gnd.n1096 gnd.n1095 0.152939
R14005 gnd.n1097 gnd.n1096 0.152939
R14006 gnd.n1114 gnd.n1097 0.152939
R14007 gnd.n6321 gnd.n1114 0.152939
R14008 gnd.n978 gnd.n966 0.152939
R14009 gnd.n979 gnd.n978 0.152939
R14010 gnd.n980 gnd.n979 0.152939
R14011 gnd.n999 gnd.n980 0.152939
R14012 gnd.n1000 gnd.n999 0.152939
R14013 gnd.n1001 gnd.n1000 0.152939
R14014 gnd.n1002 gnd.n1001 0.152939
R14015 gnd.n1020 gnd.n1002 0.152939
R14016 gnd.n1021 gnd.n1020 0.152939
R14017 gnd.n1022 gnd.n1021 0.152939
R14018 gnd.n1023 gnd.n1022 0.152939
R14019 gnd.n1041 gnd.n1023 0.152939
R14020 gnd.n1042 gnd.n1041 0.152939
R14021 gnd.n1043 gnd.n1042 0.152939
R14022 gnd.n1044 gnd.n1043 0.152939
R14023 gnd.n1062 gnd.n1044 0.152939
R14024 gnd.n1063 gnd.n1062 0.152939
R14025 gnd.n1064 gnd.n1063 0.152939
R14026 gnd.n1065 gnd.n1064 0.152939
R14027 gnd.n1083 gnd.n1065 0.152939
R14028 gnd.n1084 gnd.n1083 0.152939
R14029 gnd.n1085 gnd.n1084 0.152939
R14030 gnd.n1086 gnd.n1085 0.152939
R14031 gnd.n1104 gnd.n1086 0.152939
R14032 gnd.n1105 gnd.n1104 0.152939
R14033 gnd.n1106 gnd.n1105 0.152939
R14034 gnd.n1107 gnd.n1106 0.152939
R14035 gnd.n2087 gnd.n2086 0.152939
R14036 gnd.n2088 gnd.n2087 0.152939
R14037 gnd.n2089 gnd.n2088 0.152939
R14038 gnd.n2090 gnd.n2089 0.152939
R14039 gnd.n2091 gnd.n2090 0.152939
R14040 gnd.n2092 gnd.n2091 0.152939
R14041 gnd.n2093 gnd.n2092 0.152939
R14042 gnd.n2094 gnd.n2093 0.152939
R14043 gnd.n2095 gnd.n2094 0.152939
R14044 gnd.n2096 gnd.n2095 0.152939
R14045 gnd.n2097 gnd.n2096 0.152939
R14046 gnd.n2098 gnd.n2097 0.152939
R14047 gnd.n2099 gnd.n2098 0.152939
R14048 gnd.n2100 gnd.n2099 0.152939
R14049 gnd.n2101 gnd.n2100 0.152939
R14050 gnd.n4615 gnd.n4614 0.152939
R14051 gnd.n4614 gnd.n2106 0.152939
R14052 gnd.n2107 gnd.n2106 0.152939
R14053 gnd.n2108 gnd.n2107 0.152939
R14054 gnd.n2109 gnd.n2108 0.152939
R14055 gnd.n2110 gnd.n2109 0.152939
R14056 gnd.n2111 gnd.n2110 0.152939
R14057 gnd.n2112 gnd.n2111 0.152939
R14058 gnd.n2113 gnd.n2112 0.152939
R14059 gnd.n2114 gnd.n2113 0.152939
R14060 gnd.n2115 gnd.n2114 0.152939
R14061 gnd.n2116 gnd.n2115 0.152939
R14062 gnd.n2117 gnd.n2116 0.152939
R14063 gnd.n2118 gnd.n2117 0.152939
R14064 gnd.n2119 gnd.n2118 0.152939
R14065 gnd.n2120 gnd.n2119 0.152939
R14066 gnd.n2121 gnd.n2120 0.152939
R14067 gnd.n2122 gnd.n2121 0.152939
R14068 gnd.n4574 gnd.n2122 0.152939
R14069 gnd.n4574 gnd.n4573 0.152939
R14070 gnd.n4116 gnd.n4040 0.152939
R14071 gnd.n4042 gnd.n4040 0.152939
R14072 gnd.n4043 gnd.n4042 0.152939
R14073 gnd.n4044 gnd.n4043 0.152939
R14074 gnd.n4045 gnd.n4044 0.152939
R14075 gnd.n4046 gnd.n4045 0.152939
R14076 gnd.n4047 gnd.n4046 0.152939
R14077 gnd.n4048 gnd.n4047 0.152939
R14078 gnd.n4049 gnd.n4048 0.152939
R14079 gnd.n4050 gnd.n4049 0.152939
R14080 gnd.n4051 gnd.n4050 0.152939
R14081 gnd.n4052 gnd.n4051 0.152939
R14082 gnd.n4053 gnd.n4052 0.152939
R14083 gnd.n4054 gnd.n4053 0.152939
R14084 gnd.n4055 gnd.n4054 0.152939
R14085 gnd.n4056 gnd.n4055 0.152939
R14086 gnd.n4057 gnd.n4056 0.152939
R14087 gnd.n4058 gnd.n4057 0.152939
R14088 gnd.n4059 gnd.n4058 0.152939
R14089 gnd.n4060 gnd.n4059 0.152939
R14090 gnd.n4061 gnd.n4060 0.152939
R14091 gnd.n4062 gnd.n4061 0.152939
R14092 gnd.n4063 gnd.n4062 0.152939
R14093 gnd.n4064 gnd.n4063 0.152939
R14094 gnd.n4065 gnd.n4064 0.152939
R14095 gnd.n4066 gnd.n4065 0.152939
R14096 gnd.n4067 gnd.n4066 0.152939
R14097 gnd.n4068 gnd.n4067 0.152939
R14098 gnd.n4069 gnd.n4068 0.152939
R14099 gnd.n4070 gnd.n4069 0.152939
R14100 gnd.n4070 gnd.n2204 0.152939
R14101 gnd.n4332 gnd.n2204 0.152939
R14102 gnd.n4332 gnd.n2205 0.152939
R14103 gnd.n2207 gnd.n2205 0.152939
R14104 gnd.n2208 gnd.n2207 0.152939
R14105 gnd.n2208 gnd.n2187 0.152939
R14106 gnd.n4359 gnd.n2187 0.152939
R14107 gnd.n4360 gnd.n4359 0.152939
R14108 gnd.n4361 gnd.n4360 0.152939
R14109 gnd.n4361 gnd.n2181 0.152939
R14110 gnd.n4385 gnd.n2181 0.152939
R14111 gnd.n4386 gnd.n4385 0.152939
R14112 gnd.n4387 gnd.n4386 0.152939
R14113 gnd.n4387 gnd.n2179 0.152939
R14114 gnd.n4393 gnd.n2179 0.152939
R14115 gnd.n4394 gnd.n4393 0.152939
R14116 gnd.n4395 gnd.n4394 0.152939
R14117 gnd.n4395 gnd.n2160 0.152939
R14118 gnd.n4434 gnd.n2160 0.152939
R14119 gnd.n4435 gnd.n4434 0.152939
R14120 gnd.n4436 gnd.n4435 0.152939
R14121 gnd.n4436 gnd.n2158 0.152939
R14122 gnd.n4442 gnd.n2158 0.152939
R14123 gnd.n4443 gnd.n4442 0.152939
R14124 gnd.n4444 gnd.n4443 0.152939
R14125 gnd.n4445 gnd.n4444 0.152939
R14126 gnd.n4446 gnd.n4445 0.152939
R14127 gnd.n4446 gnd.n2135 0.152939
R14128 gnd.n4524 gnd.n2135 0.152939
R14129 gnd.n4525 gnd.n4524 0.152939
R14130 gnd.n4527 gnd.n4525 0.152939
R14131 gnd.n4527 gnd.n4526 0.152939
R14132 gnd.n4526 gnd.n2127 0.152939
R14133 gnd.n4572 gnd.n2127 0.152939
R14134 gnd.n4195 gnd.n3979 0.152939
R14135 gnd.n3982 gnd.n3979 0.152939
R14136 gnd.n3983 gnd.n3982 0.152939
R14137 gnd.n3984 gnd.n3983 0.152939
R14138 gnd.n3987 gnd.n3984 0.152939
R14139 gnd.n3988 gnd.n3987 0.152939
R14140 gnd.n3989 gnd.n3988 0.152939
R14141 gnd.n3990 gnd.n3989 0.152939
R14142 gnd.n3993 gnd.n3990 0.152939
R14143 gnd.n3994 gnd.n3993 0.152939
R14144 gnd.n3995 gnd.n3994 0.152939
R14145 gnd.n3996 gnd.n3995 0.152939
R14146 gnd.n3999 gnd.n3996 0.152939
R14147 gnd.n4000 gnd.n3999 0.152939
R14148 gnd.n4001 gnd.n4000 0.152939
R14149 gnd.n4002 gnd.n4001 0.152939
R14150 gnd.n4008 gnd.n4002 0.152939
R14151 gnd.n4009 gnd.n4008 0.152939
R14152 gnd.n4010 gnd.n4009 0.152939
R14153 gnd.n4011 gnd.n4010 0.152939
R14154 gnd.n4014 gnd.n4011 0.152939
R14155 gnd.n4015 gnd.n4014 0.152939
R14156 gnd.n4016 gnd.n4015 0.152939
R14157 gnd.n4017 gnd.n4016 0.152939
R14158 gnd.n4020 gnd.n4017 0.152939
R14159 gnd.n4021 gnd.n4020 0.152939
R14160 gnd.n4022 gnd.n4021 0.152939
R14161 gnd.n4023 gnd.n4022 0.152939
R14162 gnd.n4026 gnd.n4023 0.152939
R14163 gnd.n4027 gnd.n4026 0.152939
R14164 gnd.n4028 gnd.n4027 0.152939
R14165 gnd.n4029 gnd.n4028 0.152939
R14166 gnd.n4032 gnd.n4029 0.152939
R14167 gnd.n4033 gnd.n4032 0.152939
R14168 gnd.n4034 gnd.n4033 0.152939
R14169 gnd.n4123 gnd.n4034 0.152939
R14170 gnd.n4123 gnd.n4122 0.152939
R14171 gnd.n4122 gnd.n4121 0.152939
R14172 gnd.n4196 gnd.n2330 0.152939
R14173 gnd.n4210 gnd.n2330 0.152939
R14174 gnd.n4211 gnd.n4210 0.152939
R14175 gnd.n4212 gnd.n4211 0.152939
R14176 gnd.n4212 gnd.n2314 0.152939
R14177 gnd.n4226 gnd.n2314 0.152939
R14178 gnd.n4227 gnd.n4226 0.152939
R14179 gnd.n4228 gnd.n4227 0.152939
R14180 gnd.n4228 gnd.n2298 0.152939
R14181 gnd.n4242 gnd.n2298 0.152939
R14182 gnd.n4243 gnd.n4242 0.152939
R14183 gnd.n4244 gnd.n4243 0.152939
R14184 gnd.n4244 gnd.n2282 0.152939
R14185 gnd.n4258 gnd.n2282 0.152939
R14186 gnd.n4259 gnd.n4258 0.152939
R14187 gnd.n4260 gnd.n4259 0.152939
R14188 gnd.n4260 gnd.n2266 0.152939
R14189 gnd.n4274 gnd.n2266 0.152939
R14190 gnd.n4275 gnd.n4274 0.152939
R14191 gnd.n4276 gnd.n4275 0.152939
R14192 gnd.n4276 gnd.n2250 0.152939
R14193 gnd.n4290 gnd.n2250 0.152939
R14194 gnd.n4291 gnd.n4290 0.152939
R14195 gnd.n4293 gnd.n4291 0.152939
R14196 gnd.n4293 gnd.n4292 0.152939
R14197 gnd.n4292 gnd.n2235 0.152939
R14198 gnd.n2235 gnd.n966 0.152939
R14199 gnd.n6578 gnd.n799 0.152939
R14200 gnd.n804 gnd.n799 0.152939
R14201 gnd.n805 gnd.n804 0.152939
R14202 gnd.n806 gnd.n805 0.152939
R14203 gnd.n807 gnd.n806 0.152939
R14204 gnd.n812 gnd.n807 0.152939
R14205 gnd.n813 gnd.n812 0.152939
R14206 gnd.n814 gnd.n813 0.152939
R14207 gnd.n815 gnd.n814 0.152939
R14208 gnd.n820 gnd.n815 0.152939
R14209 gnd.n821 gnd.n820 0.152939
R14210 gnd.n822 gnd.n821 0.152939
R14211 gnd.n823 gnd.n822 0.152939
R14212 gnd.n828 gnd.n823 0.152939
R14213 gnd.n829 gnd.n828 0.152939
R14214 gnd.n830 gnd.n829 0.152939
R14215 gnd.n831 gnd.n830 0.152939
R14216 gnd.n836 gnd.n831 0.152939
R14217 gnd.n837 gnd.n836 0.152939
R14218 gnd.n838 gnd.n837 0.152939
R14219 gnd.n839 gnd.n838 0.152939
R14220 gnd.n844 gnd.n839 0.152939
R14221 gnd.n845 gnd.n844 0.152939
R14222 gnd.n846 gnd.n845 0.152939
R14223 gnd.n847 gnd.n846 0.152939
R14224 gnd.n852 gnd.n847 0.152939
R14225 gnd.n853 gnd.n852 0.152939
R14226 gnd.n854 gnd.n853 0.152939
R14227 gnd.n855 gnd.n854 0.152939
R14228 gnd.n860 gnd.n855 0.152939
R14229 gnd.n861 gnd.n860 0.152939
R14230 gnd.n862 gnd.n861 0.152939
R14231 gnd.n863 gnd.n862 0.152939
R14232 gnd.n868 gnd.n863 0.152939
R14233 gnd.n869 gnd.n868 0.152939
R14234 gnd.n870 gnd.n869 0.152939
R14235 gnd.n871 gnd.n870 0.152939
R14236 gnd.n876 gnd.n871 0.152939
R14237 gnd.n877 gnd.n876 0.152939
R14238 gnd.n878 gnd.n877 0.152939
R14239 gnd.n879 gnd.n878 0.152939
R14240 gnd.n884 gnd.n879 0.152939
R14241 gnd.n885 gnd.n884 0.152939
R14242 gnd.n886 gnd.n885 0.152939
R14243 gnd.n887 gnd.n886 0.152939
R14244 gnd.n892 gnd.n887 0.152939
R14245 gnd.n893 gnd.n892 0.152939
R14246 gnd.n894 gnd.n893 0.152939
R14247 gnd.n895 gnd.n894 0.152939
R14248 gnd.n900 gnd.n895 0.152939
R14249 gnd.n901 gnd.n900 0.152939
R14250 gnd.n902 gnd.n901 0.152939
R14251 gnd.n903 gnd.n902 0.152939
R14252 gnd.n908 gnd.n903 0.152939
R14253 gnd.n909 gnd.n908 0.152939
R14254 gnd.n910 gnd.n909 0.152939
R14255 gnd.n911 gnd.n910 0.152939
R14256 gnd.n916 gnd.n911 0.152939
R14257 gnd.n917 gnd.n916 0.152939
R14258 gnd.n918 gnd.n917 0.152939
R14259 gnd.n919 gnd.n918 0.152939
R14260 gnd.n924 gnd.n919 0.152939
R14261 gnd.n925 gnd.n924 0.152939
R14262 gnd.n926 gnd.n925 0.152939
R14263 gnd.n927 gnd.n926 0.152939
R14264 gnd.n932 gnd.n927 0.152939
R14265 gnd.n933 gnd.n932 0.152939
R14266 gnd.n934 gnd.n933 0.152939
R14267 gnd.n935 gnd.n934 0.152939
R14268 gnd.n940 gnd.n935 0.152939
R14269 gnd.n941 gnd.n940 0.152939
R14270 gnd.n942 gnd.n941 0.152939
R14271 gnd.n943 gnd.n942 0.152939
R14272 gnd.n948 gnd.n943 0.152939
R14273 gnd.n949 gnd.n948 0.152939
R14274 gnd.n950 gnd.n949 0.152939
R14275 gnd.n951 gnd.n950 0.152939
R14276 gnd.n956 gnd.n951 0.152939
R14277 gnd.n957 gnd.n956 0.152939
R14278 gnd.n958 gnd.n957 0.152939
R14279 gnd.n959 gnd.n958 0.152939
R14280 gnd.n964 gnd.n959 0.152939
R14281 gnd.n965 gnd.n964 0.152939
R14282 gnd.n6408 gnd.n965 0.152939
R14283 gnd.n5901 gnd.n1479 0.152939
R14284 gnd.n5897 gnd.n1479 0.152939
R14285 gnd.n5897 gnd.n5896 0.152939
R14286 gnd.n5896 gnd.n5895 0.152939
R14287 gnd.n5895 gnd.n1607 0.152939
R14288 gnd.n5888 gnd.n1607 0.152939
R14289 gnd.n5888 gnd.n5887 0.152939
R14290 gnd.n5887 gnd.n5886 0.152939
R14291 gnd.n5886 gnd.n5879 0.152939
R14292 gnd.n4903 gnd.n1965 0.152939
R14293 gnd.n4917 gnd.n1965 0.152939
R14294 gnd.n4918 gnd.n4917 0.152939
R14295 gnd.n4919 gnd.n4918 0.152939
R14296 gnd.n4919 gnd.n1952 0.152939
R14297 gnd.n4933 gnd.n1952 0.152939
R14298 gnd.n4934 gnd.n4933 0.152939
R14299 gnd.n4935 gnd.n4934 0.152939
R14300 gnd.n4935 gnd.n1937 0.152939
R14301 gnd.n4949 gnd.n1937 0.152939
R14302 gnd.n4950 gnd.n4949 0.152939
R14303 gnd.n4951 gnd.n4950 0.152939
R14304 gnd.n4951 gnd.n1924 0.152939
R14305 gnd.n4965 gnd.n1924 0.152939
R14306 gnd.n4966 gnd.n4965 0.152939
R14307 gnd.n4967 gnd.n4966 0.152939
R14308 gnd.n4967 gnd.n1913 0.152939
R14309 gnd.n4981 gnd.n1913 0.152939
R14310 gnd.n4982 gnd.n4981 0.152939
R14311 gnd.n4983 gnd.n4982 0.152939
R14312 gnd.n4983 gnd.n1898 0.152939
R14313 gnd.n4999 gnd.n1898 0.152939
R14314 gnd.n5000 gnd.n4999 0.152939
R14315 gnd.n5002 gnd.n5000 0.152939
R14316 gnd.n5002 gnd.n5001 0.152939
R14317 gnd.n5001 gnd.n1866 0.152939
R14318 gnd.n5583 gnd.n1866 0.152939
R14319 gnd.n5584 gnd.n5583 0.152939
R14320 gnd.n5585 gnd.n5584 0.152939
R14321 gnd.n5585 gnd.n1852 0.152939
R14322 gnd.n5599 gnd.n1852 0.152939
R14323 gnd.n5600 gnd.n5599 0.152939
R14324 gnd.n5601 gnd.n5600 0.152939
R14325 gnd.n5601 gnd.n1837 0.152939
R14326 gnd.n5615 gnd.n1837 0.152939
R14327 gnd.n5616 gnd.n5615 0.152939
R14328 gnd.n5617 gnd.n5616 0.152939
R14329 gnd.n5617 gnd.n1823 0.152939
R14330 gnd.n5631 gnd.n1823 0.152939
R14331 gnd.n5632 gnd.n5631 0.152939
R14332 gnd.n5633 gnd.n5632 0.152939
R14333 gnd.n5633 gnd.n1808 0.152939
R14334 gnd.n5647 gnd.n1808 0.152939
R14335 gnd.n5648 gnd.n5647 0.152939
R14336 gnd.n5649 gnd.n5648 0.152939
R14337 gnd.n5649 gnd.n1793 0.152939
R14338 gnd.n5663 gnd.n1793 0.152939
R14339 gnd.n5664 gnd.n5663 0.152939
R14340 gnd.n5665 gnd.n5664 0.152939
R14341 gnd.n5665 gnd.n1778 0.152939
R14342 gnd.n5679 gnd.n1778 0.152939
R14343 gnd.n5680 gnd.n5679 0.152939
R14344 gnd.n5681 gnd.n5680 0.152939
R14345 gnd.n5681 gnd.n1763 0.152939
R14346 gnd.n5695 gnd.n1763 0.152939
R14347 gnd.n5696 gnd.n5695 0.152939
R14348 gnd.n5697 gnd.n5696 0.152939
R14349 gnd.n5697 gnd.n1748 0.152939
R14350 gnd.n5711 gnd.n1748 0.152939
R14351 gnd.n5712 gnd.n5711 0.152939
R14352 gnd.n5713 gnd.n5712 0.152939
R14353 gnd.n5713 gnd.n1735 0.152939
R14354 gnd.n5727 gnd.n1735 0.152939
R14355 gnd.n5728 gnd.n5727 0.152939
R14356 gnd.n5729 gnd.n5728 0.152939
R14357 gnd.n5729 gnd.n1723 0.152939
R14358 gnd.n5743 gnd.n1723 0.152939
R14359 gnd.n5744 gnd.n5743 0.152939
R14360 gnd.n5745 gnd.n5744 0.152939
R14361 gnd.n5745 gnd.n1710 0.152939
R14362 gnd.n5759 gnd.n1710 0.152939
R14363 gnd.n5760 gnd.n5759 0.152939
R14364 gnd.n5761 gnd.n5760 0.152939
R14365 gnd.n5761 gnd.n1696 0.152939
R14366 gnd.n5775 gnd.n1696 0.152939
R14367 gnd.n5776 gnd.n5775 0.152939
R14368 gnd.n5777 gnd.n5776 0.152939
R14369 gnd.n5777 gnd.n1681 0.152939
R14370 gnd.n5791 gnd.n1681 0.152939
R14371 gnd.n5792 gnd.n5791 0.152939
R14372 gnd.n5793 gnd.n5792 0.152939
R14373 gnd.n5793 gnd.n1669 0.152939
R14374 gnd.n5807 gnd.n1669 0.152939
R14375 gnd.n5808 gnd.n5807 0.152939
R14376 gnd.n5809 gnd.n5808 0.152939
R14377 gnd.n5809 gnd.n1656 0.152939
R14378 gnd.n5823 gnd.n1656 0.152939
R14379 gnd.n5824 gnd.n5823 0.152939
R14380 gnd.n5825 gnd.n5824 0.152939
R14381 gnd.n5825 gnd.n1643 0.152939
R14382 gnd.n5839 gnd.n1643 0.152939
R14383 gnd.n5840 gnd.n5839 0.152939
R14384 gnd.n5841 gnd.n5840 0.152939
R14385 gnd.n5841 gnd.n1630 0.152939
R14386 gnd.n5855 gnd.n1630 0.152939
R14387 gnd.n5856 gnd.n5855 0.152939
R14388 gnd.n5859 gnd.n5856 0.152939
R14389 gnd.n5859 gnd.n5858 0.152939
R14390 gnd.n5858 gnd.n5857 0.152939
R14391 gnd.n5857 gnd.n1615 0.152939
R14392 gnd.n5878 gnd.n1615 0.152939
R14393 gnd.n4558 gnd.n4535 0.152939
R14394 gnd.n4558 gnd.n4557 0.152939
R14395 gnd.n4557 gnd.n4556 0.152939
R14396 gnd.n4556 gnd.n4541 0.152939
R14397 gnd.n4552 gnd.n4541 0.152939
R14398 gnd.n4552 gnd.n4551 0.152939
R14399 gnd.n4551 gnd.n4548 0.152939
R14400 gnd.n4548 gnd.n1976 0.152939
R14401 gnd.n4902 gnd.n1976 0.152939
R14402 gnd.n3927 gnd.n3926 0.152939
R14403 gnd.n3926 gnd.n3917 0.152939
R14404 gnd.n3922 gnd.n3917 0.152939
R14405 gnd.n3922 gnd.n3921 0.152939
R14406 gnd.n3921 gnd.n2184 0.152939
R14407 gnd.n4367 gnd.n2184 0.152939
R14408 gnd.n4368 gnd.n4367 0.152939
R14409 gnd.n4369 gnd.n4368 0.152939
R14410 gnd.n4369 gnd.n2175 0.152939
R14411 gnd.n4410 gnd.n2175 0.152939
R14412 gnd.n4410 gnd.n4409 0.152939
R14413 gnd.n4409 gnd.n4408 0.152939
R14414 gnd.n4408 gnd.n2176 0.152939
R14415 gnd.n4404 gnd.n2176 0.152939
R14416 gnd.n4404 gnd.n4403 0.152939
R14417 gnd.n4403 gnd.n4402 0.152939
R14418 gnd.n4402 gnd.n2154 0.152939
R14419 gnd.n4459 gnd.n2154 0.152939
R14420 gnd.n4459 gnd.n4458 0.152939
R14421 gnd.n4458 gnd.n4457 0.152939
R14422 gnd.n4457 gnd.n2155 0.152939
R14423 gnd.n4453 gnd.n2155 0.152939
R14424 gnd.n4453 gnd.n2138 0.152939
R14425 gnd.n4516 gnd.n2138 0.152939
R14426 gnd.n4517 gnd.n4516 0.152939
R14427 gnd.n4518 gnd.n4517 0.152939
R14428 gnd.n4518 gnd.n2132 0.152939
R14429 gnd.n4533 gnd.n2132 0.152939
R14430 gnd.n4534 gnd.n4533 0.152939
R14431 gnd.n4565 gnd.n4534 0.152939
R14432 gnd.n4565 gnd.n4564 0.152939
R14433 gnd.n6318 gnd.n1117 0.152939
R14434 gnd.n6314 gnd.n1117 0.152939
R14435 gnd.n6314 gnd.n6313 0.152939
R14436 gnd.n6313 gnd.n6312 0.152939
R14437 gnd.n6312 gnd.n1122 0.152939
R14438 gnd.n6308 gnd.n1122 0.152939
R14439 gnd.n6308 gnd.n6307 0.152939
R14440 gnd.n6307 gnd.n6306 0.152939
R14441 gnd.n6306 gnd.n1127 0.152939
R14442 gnd.n6302 gnd.n1127 0.152939
R14443 gnd.n6302 gnd.n6301 0.152939
R14444 gnd.n6301 gnd.n6300 0.152939
R14445 gnd.n6300 gnd.n1132 0.152939
R14446 gnd.n6296 gnd.n1132 0.152939
R14447 gnd.n6296 gnd.n6295 0.152939
R14448 gnd.n6295 gnd.n6294 0.152939
R14449 gnd.n6294 gnd.n1137 0.152939
R14450 gnd.n6290 gnd.n1137 0.152939
R14451 gnd.n6290 gnd.n6289 0.152939
R14452 gnd.n6289 gnd.n6288 0.152939
R14453 gnd.n6288 gnd.n1142 0.152939
R14454 gnd.n6284 gnd.n1142 0.152939
R14455 gnd.n6284 gnd.n6283 0.152939
R14456 gnd.n6283 gnd.n6282 0.152939
R14457 gnd.n6282 gnd.n1147 0.152939
R14458 gnd.n6278 gnd.n1147 0.152939
R14459 gnd.n6278 gnd.n6277 0.152939
R14460 gnd.n6277 gnd.n6276 0.152939
R14461 gnd.n6276 gnd.n1152 0.152939
R14462 gnd.n6272 gnd.n1152 0.152939
R14463 gnd.n6272 gnd.n6271 0.152939
R14464 gnd.n6271 gnd.n6270 0.152939
R14465 gnd.n6270 gnd.n1157 0.152939
R14466 gnd.n6266 gnd.n1157 0.152939
R14467 gnd.n6266 gnd.n6265 0.152939
R14468 gnd.n6265 gnd.n6264 0.152939
R14469 gnd.n6264 gnd.n1162 0.152939
R14470 gnd.n6260 gnd.n1162 0.152939
R14471 gnd.n6260 gnd.n6259 0.152939
R14472 gnd.n6259 gnd.n6258 0.152939
R14473 gnd.n6258 gnd.n1167 0.152939
R14474 gnd.n6254 gnd.n1167 0.152939
R14475 gnd.n6254 gnd.n6253 0.152939
R14476 gnd.n6253 gnd.n6252 0.152939
R14477 gnd.n6252 gnd.n1172 0.152939
R14478 gnd.n6248 gnd.n1172 0.152939
R14479 gnd.n6248 gnd.n6247 0.152939
R14480 gnd.n6247 gnd.n6246 0.152939
R14481 gnd.n6246 gnd.n1177 0.152939
R14482 gnd.n6242 gnd.n1177 0.152939
R14483 gnd.n6242 gnd.n6241 0.152939
R14484 gnd.n6241 gnd.n6240 0.152939
R14485 gnd.n6240 gnd.n1182 0.152939
R14486 gnd.n6236 gnd.n1182 0.152939
R14487 gnd.n6236 gnd.n6235 0.152939
R14488 gnd.n6235 gnd.n6234 0.152939
R14489 gnd.n6234 gnd.n1187 0.152939
R14490 gnd.n6230 gnd.n1187 0.152939
R14491 gnd.n6230 gnd.n6229 0.152939
R14492 gnd.n6229 gnd.n6228 0.152939
R14493 gnd.n6228 gnd.n1192 0.152939
R14494 gnd.n6224 gnd.n1192 0.152939
R14495 gnd.n6224 gnd.n6223 0.152939
R14496 gnd.n6223 gnd.n6222 0.152939
R14497 gnd.n6222 gnd.n1197 0.152939
R14498 gnd.n6218 gnd.n1197 0.152939
R14499 gnd.n6218 gnd.n6217 0.152939
R14500 gnd.n6217 gnd.n6216 0.152939
R14501 gnd.n6216 gnd.n1202 0.152939
R14502 gnd.n6212 gnd.n1202 0.152939
R14503 gnd.n6212 gnd.n6211 0.152939
R14504 gnd.n6211 gnd.n6210 0.152939
R14505 gnd.n6210 gnd.n1207 0.152939
R14506 gnd.n6206 gnd.n1207 0.152939
R14507 gnd.n6206 gnd.n6205 0.152939
R14508 gnd.n6205 gnd.n6204 0.152939
R14509 gnd.n6204 gnd.n1212 0.152939
R14510 gnd.n6200 gnd.n1212 0.152939
R14511 gnd.n6200 gnd.n6199 0.152939
R14512 gnd.n6199 gnd.n6198 0.152939
R14513 gnd.n6198 gnd.n1217 0.152939
R14514 gnd.n6194 gnd.n1217 0.152939
R14515 gnd.n6194 gnd.n6193 0.152939
R14516 gnd.n6193 gnd.n6192 0.152939
R14517 gnd.n6192 gnd.n1222 0.152939
R14518 gnd.n6188 gnd.n1222 0.152939
R14519 gnd.n6188 gnd.n6187 0.152939
R14520 gnd.n6187 gnd.n6186 0.152939
R14521 gnd.n6186 gnd.n1227 0.152939
R14522 gnd.n6182 gnd.n1227 0.152939
R14523 gnd.n6182 gnd.n6181 0.152939
R14524 gnd.n6181 gnd.n6180 0.152939
R14525 gnd.n6180 gnd.n1232 0.152939
R14526 gnd.n6176 gnd.n1232 0.152939
R14527 gnd.n6176 gnd.n6175 0.152939
R14528 gnd.n6175 gnd.n6174 0.152939
R14529 gnd.n6174 gnd.n1237 0.152939
R14530 gnd.n6170 gnd.n1237 0.152939
R14531 gnd.n6170 gnd.n6169 0.152939
R14532 gnd.n6169 gnd.n6168 0.152939
R14533 gnd.n6168 gnd.n1242 0.152939
R14534 gnd.n6076 gnd.n6075 0.152939
R14535 gnd.n6075 gnd.n6074 0.152939
R14536 gnd.n6074 gnd.n1343 0.152939
R14537 gnd.n6070 gnd.n1343 0.152939
R14538 gnd.n6070 gnd.n6069 0.152939
R14539 gnd.n6069 gnd.n6068 0.152939
R14540 gnd.n6068 gnd.n1348 0.152939
R14541 gnd.n6064 gnd.n1348 0.152939
R14542 gnd.n6064 gnd.n6063 0.152939
R14543 gnd.n6063 gnd.n6062 0.152939
R14544 gnd.n6062 gnd.n1353 0.152939
R14545 gnd.n6058 gnd.n1353 0.152939
R14546 gnd.n6058 gnd.n6057 0.152939
R14547 gnd.n6057 gnd.n6056 0.152939
R14548 gnd.n6056 gnd.n1358 0.152939
R14549 gnd.n6052 gnd.n1358 0.152939
R14550 gnd.n6052 gnd.n407 0.152939
R14551 gnd.n7232 gnd.n407 0.152939
R14552 gnd.n7232 gnd.n7231 0.152939
R14553 gnd.n7231 gnd.n7230 0.152939
R14554 gnd.n7230 gnd.n408 0.152939
R14555 gnd.n408 gnd.n375 0.152939
R14556 gnd.n7278 gnd.n375 0.152939
R14557 gnd.n7278 gnd.n7277 0.152939
R14558 gnd.n7277 gnd.n7276 0.152939
R14559 gnd.n7276 gnd.n376 0.152939
R14560 gnd.n7272 gnd.n376 0.152939
R14561 gnd.n7272 gnd.n320 0.152939
R14562 gnd.n7409 gnd.n320 0.152939
R14563 gnd.n7409 gnd.n7408 0.152939
R14564 gnd.n7408 gnd.n7407 0.152939
R14565 gnd.n7407 gnd.n321 0.152939
R14566 gnd.n7403 gnd.n321 0.152939
R14567 gnd.n7403 gnd.n7402 0.152939
R14568 gnd.n7402 gnd.n7401 0.152939
R14569 gnd.n7401 gnd.n326 0.152939
R14570 gnd.n326 gnd.n296 0.152939
R14571 gnd.n7424 gnd.n296 0.152939
R14572 gnd.n7425 gnd.n7424 0.152939
R14573 gnd.n7426 gnd.n7425 0.152939
R14574 gnd.n7426 gnd.n280 0.152939
R14575 gnd.n7440 gnd.n280 0.152939
R14576 gnd.n7441 gnd.n7440 0.152939
R14577 gnd.n7442 gnd.n7441 0.152939
R14578 gnd.n7442 gnd.n266 0.152939
R14579 gnd.n7456 gnd.n266 0.152939
R14580 gnd.n7457 gnd.n7456 0.152939
R14581 gnd.n7458 gnd.n7457 0.152939
R14582 gnd.n7458 gnd.n250 0.152939
R14583 gnd.n7472 gnd.n250 0.152939
R14584 gnd.n7473 gnd.n7472 0.152939
R14585 gnd.n7474 gnd.n7473 0.152939
R14586 gnd.n7474 gnd.n235 0.152939
R14587 gnd.n7488 gnd.n235 0.152939
R14588 gnd.n7489 gnd.n7488 0.152939
R14589 gnd.n7490 gnd.n7489 0.152939
R14590 gnd.n7490 gnd.n220 0.152939
R14591 gnd.n7504 gnd.n220 0.152939
R14592 gnd.n7505 gnd.n7504 0.152939
R14593 gnd.n7574 gnd.n7505 0.152939
R14594 gnd.n7574 gnd.n7573 0.152939
R14595 gnd.n7573 gnd.n7572 0.152939
R14596 gnd.n7572 gnd.n7506 0.152939
R14597 gnd.n7568 gnd.n7506 0.152939
R14598 gnd.n7567 gnd.n7508 0.152939
R14599 gnd.n7563 gnd.n7508 0.152939
R14600 gnd.n7563 gnd.n7562 0.152939
R14601 gnd.n7562 gnd.n7561 0.152939
R14602 gnd.n7561 gnd.n7514 0.152939
R14603 gnd.n7557 gnd.n7514 0.152939
R14604 gnd.n7557 gnd.n7556 0.152939
R14605 gnd.n7556 gnd.n7555 0.152939
R14606 gnd.n7555 gnd.n7522 0.152939
R14607 gnd.n7551 gnd.n7522 0.152939
R14608 gnd.n7551 gnd.n7550 0.152939
R14609 gnd.n7550 gnd.n7549 0.152939
R14610 gnd.n7549 gnd.n7530 0.152939
R14611 gnd.n7545 gnd.n7530 0.152939
R14612 gnd.n7545 gnd.n7544 0.152939
R14613 gnd.n7544 gnd.n7543 0.152939
R14614 gnd.n7543 gnd.n121 0.152939
R14615 gnd.n7669 gnd.n121 0.152939
R14616 gnd.n5917 gnd.n5903 0.152939
R14617 gnd.n5918 gnd.n5917 0.152939
R14618 gnd.n5920 gnd.n5918 0.152939
R14619 gnd.n5920 gnd.n5919 0.152939
R14620 gnd.n5919 gnd.n1419 0.152939
R14621 gnd.n5948 gnd.n1419 0.152939
R14622 gnd.n5949 gnd.n5948 0.152939
R14623 gnd.n5956 gnd.n5949 0.152939
R14624 gnd.n5956 gnd.n5955 0.152939
R14625 gnd.n5955 gnd.n5954 0.152939
R14626 gnd.n5954 gnd.n5950 0.152939
R14627 gnd.n5950 gnd.n1384 0.152939
R14628 gnd.n6016 gnd.n1384 0.152939
R14629 gnd.n6016 gnd.n6015 0.152939
R14630 gnd.n6015 gnd.n6014 0.152939
R14631 gnd.n6014 gnd.n1385 0.152939
R14632 gnd.n6010 gnd.n1385 0.152939
R14633 gnd.n6010 gnd.n6009 0.152939
R14634 gnd.n6009 gnd.n6008 0.152939
R14635 gnd.n6008 gnd.n6003 0.152939
R14636 gnd.n6003 gnd.n6002 0.152939
R14637 gnd.n6002 gnd.n381 0.152939
R14638 gnd.n7263 gnd.n381 0.152939
R14639 gnd.n7264 gnd.n7263 0.152939
R14640 gnd.n7266 gnd.n7264 0.152939
R14641 gnd.n7266 gnd.n7265 0.152939
R14642 gnd.n7265 gnd.n347 0.152939
R14643 gnd.n7308 gnd.n347 0.152939
R14644 gnd.n7309 gnd.n7308 0.152939
R14645 gnd.n7310 gnd.n7309 0.152939
R14646 gnd.n7310 gnd.n79 0.152939
R14647 gnd.n7718 gnd.n79 0.152939
R14648 gnd.n7718 gnd.n7717 0.152939
R14649 gnd.n7717 gnd.n81 0.152939
R14650 gnd.n7713 gnd.n81 0.152939
R14651 gnd.n7713 gnd.n7712 0.152939
R14652 gnd.n7712 gnd.n7711 0.152939
R14653 gnd.n7711 gnd.n86 0.152939
R14654 gnd.n7707 gnd.n86 0.152939
R14655 gnd.n7707 gnd.n7706 0.152939
R14656 gnd.n7706 gnd.n7705 0.152939
R14657 gnd.n7705 gnd.n91 0.152939
R14658 gnd.n7701 gnd.n91 0.152939
R14659 gnd.n7701 gnd.n7700 0.152939
R14660 gnd.n7700 gnd.n7699 0.152939
R14661 gnd.n7699 gnd.n96 0.152939
R14662 gnd.n7695 gnd.n96 0.152939
R14663 gnd.n7695 gnd.n7694 0.152939
R14664 gnd.n7694 gnd.n7693 0.152939
R14665 gnd.n7693 gnd.n101 0.152939
R14666 gnd.n7689 gnd.n101 0.152939
R14667 gnd.n7689 gnd.n7688 0.152939
R14668 gnd.n7688 gnd.n7687 0.152939
R14669 gnd.n7687 gnd.n106 0.152939
R14670 gnd.n7683 gnd.n106 0.152939
R14671 gnd.n7683 gnd.n7682 0.152939
R14672 gnd.n7682 gnd.n7681 0.152939
R14673 gnd.n7681 gnd.n111 0.152939
R14674 gnd.n7677 gnd.n111 0.152939
R14675 gnd.n7677 gnd.n7676 0.152939
R14676 gnd.n7676 gnd.n7675 0.152939
R14677 gnd.n7675 gnd.n116 0.152939
R14678 gnd.n7671 gnd.n116 0.152939
R14679 gnd.n7671 gnd.n7670 0.152939
R14680 gnd.n5902 gnd.n5901 0.151415
R14681 gnd.n4563 gnd.n4535 0.151415
R14682 gnd.n3928 gnd.n3914 0.145814
R14683 gnd.n3928 gnd.n3927 0.145814
R14684 gnd.n3210 gnd.n3209 0.0767195
R14685 gnd.n3209 gnd.n3208 0.0767195
R14686 gnd.n6320 gnd.n6319 0.063
R14687 gnd.n1518 gnd.n1342 0.063
R14688 gnd.n3776 gnd.n2379 0.0477147
R14689 gnd.n2973 gnd.n2861 0.0442063
R14690 gnd.n2974 gnd.n2973 0.0442063
R14691 gnd.n2975 gnd.n2974 0.0442063
R14692 gnd.n2975 gnd.n2850 0.0442063
R14693 gnd.n2989 gnd.n2850 0.0442063
R14694 gnd.n2990 gnd.n2989 0.0442063
R14695 gnd.n2991 gnd.n2990 0.0442063
R14696 gnd.n2991 gnd.n2837 0.0442063
R14697 gnd.n3035 gnd.n2837 0.0442063
R14698 gnd.n3036 gnd.n3035 0.0442063
R14699 gnd.n3038 gnd.n2771 0.0344674
R14700 gnd.n1597 gnd.n1478 0.0343753
R14701 gnd.n4562 gnd.n2045 0.0343753
R14702 gnd.n3058 gnd.n3057 0.0269946
R14703 gnd.n3060 gnd.n3059 0.0269946
R14704 gnd.n2766 gnd.n2764 0.0269946
R14705 gnd.n3070 gnd.n3068 0.0269946
R14706 gnd.n3069 gnd.n2745 0.0269946
R14707 gnd.n3089 gnd.n3088 0.0269946
R14708 gnd.n3091 gnd.n3090 0.0269946
R14709 gnd.n2740 gnd.n2739 0.0269946
R14710 gnd.n3101 gnd.n2735 0.0269946
R14711 gnd.n3100 gnd.n2737 0.0269946
R14712 gnd.n2736 gnd.n2718 0.0269946
R14713 gnd.n3121 gnd.n2719 0.0269946
R14714 gnd.n3120 gnd.n2720 0.0269946
R14715 gnd.n3154 gnd.n2695 0.0269946
R14716 gnd.n3156 gnd.n3155 0.0269946
R14717 gnd.n3157 gnd.n2642 0.0269946
R14718 gnd.n2690 gnd.n2643 0.0269946
R14719 gnd.n2692 gnd.n2644 0.0269946
R14720 gnd.n3167 gnd.n3166 0.0269946
R14721 gnd.n3169 gnd.n3168 0.0269946
R14722 gnd.n3170 gnd.n2664 0.0269946
R14723 gnd.n3172 gnd.n2665 0.0269946
R14724 gnd.n3175 gnd.n2666 0.0269946
R14725 gnd.n3178 gnd.n3177 0.0269946
R14726 gnd.n3180 gnd.n3179 0.0269946
R14727 gnd.n3245 gnd.n2553 0.0269946
R14728 gnd.n3247 gnd.n3246 0.0269946
R14729 gnd.n3256 gnd.n2546 0.0269946
R14730 gnd.n3258 gnd.n3257 0.0269946
R14731 gnd.n3259 gnd.n2544 0.0269946
R14732 gnd.n3266 gnd.n3262 0.0269946
R14733 gnd.n3265 gnd.n3264 0.0269946
R14734 gnd.n3263 gnd.n2523 0.0269946
R14735 gnd.n3288 gnd.n2524 0.0269946
R14736 gnd.n3287 gnd.n2525 0.0269946
R14737 gnd.n3330 gnd.n2498 0.0269946
R14738 gnd.n3332 gnd.n3331 0.0269946
R14739 gnd.n3341 gnd.n2491 0.0269946
R14740 gnd.n3343 gnd.n3342 0.0269946
R14741 gnd.n3344 gnd.n2489 0.0269946
R14742 gnd.n3351 gnd.n3347 0.0269946
R14743 gnd.n3350 gnd.n3349 0.0269946
R14744 gnd.n3348 gnd.n2468 0.0269946
R14745 gnd.n3373 gnd.n2469 0.0269946
R14746 gnd.n3372 gnd.n2470 0.0269946
R14747 gnd.n3419 gnd.n2444 0.0269946
R14748 gnd.n3421 gnd.n3420 0.0269946
R14749 gnd.n3430 gnd.n2437 0.0269946
R14750 gnd.n3689 gnd.n2435 0.0269946
R14751 gnd.n3694 gnd.n3692 0.0269946
R14752 gnd.n3693 gnd.n2416 0.0269946
R14753 gnd.n3718 gnd.n3717 0.0269946
R14754 gnd.n1520 gnd.n1518 0.0245515
R14755 gnd.n6319 gnd.n1116 0.0245515
R14756 gnd.n3038 gnd.n3037 0.0202011
R14757 gnd.n1520 gnd.n1519 0.0174377
R14758 gnd.n1519 gnd.n1515 0.0174377
R14759 gnd.n1529 gnd.n1515 0.0174377
R14760 gnd.n1529 gnd.n1528 0.0174377
R14761 gnd.n1528 gnd.n1516 0.0174377
R14762 gnd.n1516 gnd.n1511 0.0174377
R14763 gnd.n1537 gnd.n1511 0.0174377
R14764 gnd.n1539 gnd.n1537 0.0174377
R14765 gnd.n1539 gnd.n1538 0.0174377
R14766 gnd.n1538 gnd.n1508 0.0174377
R14767 gnd.n1548 gnd.n1508 0.0174377
R14768 gnd.n1548 gnd.n1547 0.0174377
R14769 gnd.n1547 gnd.n1509 0.0174377
R14770 gnd.n1509 gnd.n1504 0.0174377
R14771 gnd.n1556 gnd.n1504 0.0174377
R14772 gnd.n1558 gnd.n1556 0.0174377
R14773 gnd.n1558 gnd.n1557 0.0174377
R14774 gnd.n1557 gnd.n1501 0.0174377
R14775 gnd.n1567 gnd.n1501 0.0174377
R14776 gnd.n1567 gnd.n1566 0.0174377
R14777 gnd.n1566 gnd.n1502 0.0174377
R14778 gnd.n1502 gnd.n1497 0.0174377
R14779 gnd.n1575 gnd.n1497 0.0174377
R14780 gnd.n1576 gnd.n1575 0.0174377
R14781 gnd.n1576 gnd.n1495 0.0174377
R14782 gnd.n1581 gnd.n1495 0.0174377
R14783 gnd.n1583 gnd.n1581 0.0174377
R14784 gnd.n1583 gnd.n1582 0.0174377
R14785 gnd.n1582 gnd.n1491 0.0174377
R14786 gnd.n1592 gnd.n1491 0.0174377
R14787 gnd.n1592 gnd.n1591 0.0174377
R14788 gnd.n1591 gnd.n1484 0.0174377
R14789 gnd.n1484 gnd.n1483 0.0174377
R14790 gnd.n1596 gnd.n1483 0.0174377
R14791 gnd.n1597 gnd.n1596 0.0174377
R14792 gnd.n1994 gnd.n1116 0.0174377
R14793 gnd.n1996 gnd.n1994 0.0174377
R14794 gnd.n4892 gnd.n1996 0.0174377
R14795 gnd.n4892 gnd.n4891 0.0174377
R14796 gnd.n4891 gnd.n1997 0.0174377
R14797 gnd.n4888 gnd.n1997 0.0174377
R14798 gnd.n4888 gnd.n4887 0.0174377
R14799 gnd.n4887 gnd.n2002 0.0174377
R14800 gnd.n4884 gnd.n2002 0.0174377
R14801 gnd.n4884 gnd.n4883 0.0174377
R14802 gnd.n4883 gnd.n2007 0.0174377
R14803 gnd.n4880 gnd.n2007 0.0174377
R14804 gnd.n4880 gnd.n4879 0.0174377
R14805 gnd.n4879 gnd.n2011 0.0174377
R14806 gnd.n4876 gnd.n2011 0.0174377
R14807 gnd.n4876 gnd.n4875 0.0174377
R14808 gnd.n4875 gnd.n2015 0.0174377
R14809 gnd.n4872 gnd.n2015 0.0174377
R14810 gnd.n4872 gnd.n4871 0.0174377
R14811 gnd.n4871 gnd.n2019 0.0174377
R14812 gnd.n4868 gnd.n2019 0.0174377
R14813 gnd.n4868 gnd.n4867 0.0174377
R14814 gnd.n4867 gnd.n2025 0.0174377
R14815 gnd.n4864 gnd.n2025 0.0174377
R14816 gnd.n4864 gnd.n4863 0.0174377
R14817 gnd.n4863 gnd.n2029 0.0174377
R14818 gnd.n4860 gnd.n2029 0.0174377
R14819 gnd.n4860 gnd.n4859 0.0174377
R14820 gnd.n4859 gnd.n2033 0.0174377
R14821 gnd.n4856 gnd.n2033 0.0174377
R14822 gnd.n4856 gnd.n4855 0.0174377
R14823 gnd.n4855 gnd.n2039 0.0174377
R14824 gnd.n4852 gnd.n2039 0.0174377
R14825 gnd.n4852 gnd.n4851 0.0174377
R14826 gnd.n4851 gnd.n2045 0.0174377
R14827 gnd.n3037 gnd.n3036 0.0148637
R14828 gnd.n3687 gnd.n3431 0.0144266
R14829 gnd.n3688 gnd.n3687 0.0130679
R14830 gnd.n3057 gnd.n2771 0.00797283
R14831 gnd.n3059 gnd.n3058 0.00797283
R14832 gnd.n3060 gnd.n2766 0.00797283
R14833 gnd.n3068 gnd.n2764 0.00797283
R14834 gnd.n3070 gnd.n3069 0.00797283
R14835 gnd.n3088 gnd.n2745 0.00797283
R14836 gnd.n3090 gnd.n3089 0.00797283
R14837 gnd.n3091 gnd.n2740 0.00797283
R14838 gnd.n2739 gnd.n2735 0.00797283
R14839 gnd.n3101 gnd.n3100 0.00797283
R14840 gnd.n2737 gnd.n2736 0.00797283
R14841 gnd.n2719 gnd.n2718 0.00797283
R14842 gnd.n3121 gnd.n3120 0.00797283
R14843 gnd.n2720 gnd.n2695 0.00797283
R14844 gnd.n3155 gnd.n3154 0.00797283
R14845 gnd.n3157 gnd.n3156 0.00797283
R14846 gnd.n2690 gnd.n2642 0.00797283
R14847 gnd.n2692 gnd.n2643 0.00797283
R14848 gnd.n3166 gnd.n2644 0.00797283
R14849 gnd.n3168 gnd.n3167 0.00797283
R14850 gnd.n3170 gnd.n3169 0.00797283
R14851 gnd.n3172 gnd.n2664 0.00797283
R14852 gnd.n3175 gnd.n2665 0.00797283
R14853 gnd.n3177 gnd.n2666 0.00797283
R14854 gnd.n3180 gnd.n3178 0.00797283
R14855 gnd.n3179 gnd.n2553 0.00797283
R14856 gnd.n3247 gnd.n3245 0.00797283
R14857 gnd.n3246 gnd.n2546 0.00797283
R14858 gnd.n3257 gnd.n3256 0.00797283
R14859 gnd.n3259 gnd.n3258 0.00797283
R14860 gnd.n3262 gnd.n2544 0.00797283
R14861 gnd.n3266 gnd.n3265 0.00797283
R14862 gnd.n3264 gnd.n3263 0.00797283
R14863 gnd.n2524 gnd.n2523 0.00797283
R14864 gnd.n3288 gnd.n3287 0.00797283
R14865 gnd.n2525 gnd.n2498 0.00797283
R14866 gnd.n3332 gnd.n3330 0.00797283
R14867 gnd.n3331 gnd.n2491 0.00797283
R14868 gnd.n3342 gnd.n3341 0.00797283
R14869 gnd.n3344 gnd.n3343 0.00797283
R14870 gnd.n3347 gnd.n2489 0.00797283
R14871 gnd.n3351 gnd.n3350 0.00797283
R14872 gnd.n3349 gnd.n3348 0.00797283
R14873 gnd.n2469 gnd.n2468 0.00797283
R14874 gnd.n3373 gnd.n3372 0.00797283
R14875 gnd.n2470 gnd.n2444 0.00797283
R14876 gnd.n3421 gnd.n3419 0.00797283
R14877 gnd.n3420 gnd.n2437 0.00797283
R14878 gnd.n3431 gnd.n3430 0.00797283
R14879 gnd.n3689 gnd.n3688 0.00797283
R14880 gnd.n3692 gnd.n2435 0.00797283
R14881 gnd.n3694 gnd.n3693 0.00797283
R14882 gnd.n3717 gnd.n2416 0.00797283
R14883 gnd.n3718 gnd.n2379 0.00797283
R14884 gnd.n337 gnd.n321 0.00433921
R14885 gnd.n4333 gnd.n4332 0.00433921
R14886 gnd.n5902 gnd.n1478 0.000838753
R14887 gnd.n4563 gnd.n4562 0.000838753
R14888 vdd.n315 vdd.n279 756.745
R14889 vdd.n260 vdd.n224 756.745
R14890 vdd.n217 vdd.n181 756.745
R14891 vdd.n162 vdd.n126 756.745
R14892 vdd.n120 vdd.n84 756.745
R14893 vdd.n65 vdd.n29 756.745
R14894 vdd.n2046 vdd.n2010 756.745
R14895 vdd.n2101 vdd.n2065 756.745
R14896 vdd.n1948 vdd.n1912 756.745
R14897 vdd.n2003 vdd.n1967 756.745
R14898 vdd.n1851 vdd.n1815 756.745
R14899 vdd.n1906 vdd.n1870 756.745
R14900 vdd.n1224 vdd.t16 640.208
R14901 vdd.n952 vdd.t58 640.208
R14902 vdd.n1244 vdd.t31 640.208
R14903 vdd.n943 vdd.t76 640.208
R14904 vdd.n843 vdd.t34 640.208
R14905 vdd.n2621 vdd.t73 640.208
R14906 vdd.n804 vdd.t82 640.208
R14907 vdd.n2618 vdd.t62 640.208
R14908 vdd.n768 vdd.t12 640.208
R14909 vdd.n1014 vdd.t66 640.208
R14910 vdd.n1510 vdd.t49 592.009
R14911 vdd.n1666 vdd.t41 592.009
R14912 vdd.n1702 vdd.t52 592.009
R14913 vdd.n2186 vdd.t24 592.009
R14914 vdd.n1161 vdd.t55 592.009
R14915 vdd.n1121 vdd.t70 592.009
R14916 vdd.n405 vdd.t45 592.009
R14917 vdd.n419 vdd.t79 592.009
R14918 vdd.n431 vdd.t85 592.009
R14919 vdd.n723 vdd.t28 592.009
R14920 vdd.n686 vdd.t38 592.009
R14921 vdd.n3105 vdd.t20 592.009
R14922 vdd.n316 vdd.n315 585
R14923 vdd.n314 vdd.n281 585
R14924 vdd.n313 vdd.n312 585
R14925 vdd.n284 vdd.n282 585
R14926 vdd.n307 vdd.n306 585
R14927 vdd.n305 vdd.n304 585
R14928 vdd.n288 vdd.n287 585
R14929 vdd.n299 vdd.n298 585
R14930 vdd.n297 vdd.n296 585
R14931 vdd.n292 vdd.n291 585
R14932 vdd.n261 vdd.n260 585
R14933 vdd.n259 vdd.n226 585
R14934 vdd.n258 vdd.n257 585
R14935 vdd.n229 vdd.n227 585
R14936 vdd.n252 vdd.n251 585
R14937 vdd.n250 vdd.n249 585
R14938 vdd.n233 vdd.n232 585
R14939 vdd.n244 vdd.n243 585
R14940 vdd.n242 vdd.n241 585
R14941 vdd.n237 vdd.n236 585
R14942 vdd.n218 vdd.n217 585
R14943 vdd.n216 vdd.n183 585
R14944 vdd.n215 vdd.n214 585
R14945 vdd.n186 vdd.n184 585
R14946 vdd.n209 vdd.n208 585
R14947 vdd.n207 vdd.n206 585
R14948 vdd.n190 vdd.n189 585
R14949 vdd.n201 vdd.n200 585
R14950 vdd.n199 vdd.n198 585
R14951 vdd.n194 vdd.n193 585
R14952 vdd.n163 vdd.n162 585
R14953 vdd.n161 vdd.n128 585
R14954 vdd.n160 vdd.n159 585
R14955 vdd.n131 vdd.n129 585
R14956 vdd.n154 vdd.n153 585
R14957 vdd.n152 vdd.n151 585
R14958 vdd.n135 vdd.n134 585
R14959 vdd.n146 vdd.n145 585
R14960 vdd.n144 vdd.n143 585
R14961 vdd.n139 vdd.n138 585
R14962 vdd.n121 vdd.n120 585
R14963 vdd.n119 vdd.n86 585
R14964 vdd.n118 vdd.n117 585
R14965 vdd.n89 vdd.n87 585
R14966 vdd.n112 vdd.n111 585
R14967 vdd.n110 vdd.n109 585
R14968 vdd.n93 vdd.n92 585
R14969 vdd.n104 vdd.n103 585
R14970 vdd.n102 vdd.n101 585
R14971 vdd.n97 vdd.n96 585
R14972 vdd.n66 vdd.n65 585
R14973 vdd.n64 vdd.n31 585
R14974 vdd.n63 vdd.n62 585
R14975 vdd.n34 vdd.n32 585
R14976 vdd.n57 vdd.n56 585
R14977 vdd.n55 vdd.n54 585
R14978 vdd.n38 vdd.n37 585
R14979 vdd.n49 vdd.n48 585
R14980 vdd.n47 vdd.n46 585
R14981 vdd.n42 vdd.n41 585
R14982 vdd.n2047 vdd.n2046 585
R14983 vdd.n2045 vdd.n2012 585
R14984 vdd.n2044 vdd.n2043 585
R14985 vdd.n2015 vdd.n2013 585
R14986 vdd.n2038 vdd.n2037 585
R14987 vdd.n2036 vdd.n2035 585
R14988 vdd.n2019 vdd.n2018 585
R14989 vdd.n2030 vdd.n2029 585
R14990 vdd.n2028 vdd.n2027 585
R14991 vdd.n2023 vdd.n2022 585
R14992 vdd.n2102 vdd.n2101 585
R14993 vdd.n2100 vdd.n2067 585
R14994 vdd.n2099 vdd.n2098 585
R14995 vdd.n2070 vdd.n2068 585
R14996 vdd.n2093 vdd.n2092 585
R14997 vdd.n2091 vdd.n2090 585
R14998 vdd.n2074 vdd.n2073 585
R14999 vdd.n2085 vdd.n2084 585
R15000 vdd.n2083 vdd.n2082 585
R15001 vdd.n2078 vdd.n2077 585
R15002 vdd.n1949 vdd.n1948 585
R15003 vdd.n1947 vdd.n1914 585
R15004 vdd.n1946 vdd.n1945 585
R15005 vdd.n1917 vdd.n1915 585
R15006 vdd.n1940 vdd.n1939 585
R15007 vdd.n1938 vdd.n1937 585
R15008 vdd.n1921 vdd.n1920 585
R15009 vdd.n1932 vdd.n1931 585
R15010 vdd.n1930 vdd.n1929 585
R15011 vdd.n1925 vdd.n1924 585
R15012 vdd.n2004 vdd.n2003 585
R15013 vdd.n2002 vdd.n1969 585
R15014 vdd.n2001 vdd.n2000 585
R15015 vdd.n1972 vdd.n1970 585
R15016 vdd.n1995 vdd.n1994 585
R15017 vdd.n1993 vdd.n1992 585
R15018 vdd.n1976 vdd.n1975 585
R15019 vdd.n1987 vdd.n1986 585
R15020 vdd.n1985 vdd.n1984 585
R15021 vdd.n1980 vdd.n1979 585
R15022 vdd.n1852 vdd.n1851 585
R15023 vdd.n1850 vdd.n1817 585
R15024 vdd.n1849 vdd.n1848 585
R15025 vdd.n1820 vdd.n1818 585
R15026 vdd.n1843 vdd.n1842 585
R15027 vdd.n1841 vdd.n1840 585
R15028 vdd.n1824 vdd.n1823 585
R15029 vdd.n1835 vdd.n1834 585
R15030 vdd.n1833 vdd.n1832 585
R15031 vdd.n1828 vdd.n1827 585
R15032 vdd.n1907 vdd.n1906 585
R15033 vdd.n1905 vdd.n1872 585
R15034 vdd.n1904 vdd.n1903 585
R15035 vdd.n1875 vdd.n1873 585
R15036 vdd.n1898 vdd.n1897 585
R15037 vdd.n1896 vdd.n1895 585
R15038 vdd.n1879 vdd.n1878 585
R15039 vdd.n1890 vdd.n1889 585
R15040 vdd.n1888 vdd.n1887 585
R15041 vdd.n1883 vdd.n1882 585
R15042 vdd.n445 vdd.n370 462.44
R15043 vdd.n3343 vdd.n372 462.44
R15044 vdd.n3238 vdd.n657 462.44
R15045 vdd.n3236 vdd.n660 462.44
R15046 vdd.n2181 vdd.n1409 462.44
R15047 vdd.n2184 vdd.n2183 462.44
R15048 vdd.n1737 vdd.n1507 462.44
R15049 vdd.n1734 vdd.n1505 462.44
R15050 vdd.n293 vdd.t220 329.043
R15051 vdd.n238 vdd.t198 329.043
R15052 vdd.n195 vdd.t210 329.043
R15053 vdd.n140 vdd.t185 329.043
R15054 vdd.n98 vdd.t172 329.043
R15055 vdd.n43 vdd.t153 329.043
R15056 vdd.n2024 vdd.t231 329.043
R15057 vdd.n2079 vdd.t141 329.043
R15058 vdd.n1926 vdd.t221 329.043
R15059 vdd.n1981 vdd.t120 329.043
R15060 vdd.n1829 vdd.t155 329.043
R15061 vdd.n1884 vdd.t173 329.043
R15062 vdd.n1510 vdd.t51 319.788
R15063 vdd.n1666 vdd.t44 319.788
R15064 vdd.n1702 vdd.t54 319.788
R15065 vdd.n2186 vdd.t26 319.788
R15066 vdd.n1161 vdd.t56 319.788
R15067 vdd.n1121 vdd.t71 319.788
R15068 vdd.n405 vdd.t47 319.788
R15069 vdd.n419 vdd.t80 319.788
R15070 vdd.n431 vdd.t86 319.788
R15071 vdd.n723 vdd.t30 319.788
R15072 vdd.n686 vdd.t40 319.788
R15073 vdd.n3105 vdd.t23 319.788
R15074 vdd.n1511 vdd.t50 303.69
R15075 vdd.n1667 vdd.t43 303.69
R15076 vdd.n1703 vdd.t53 303.69
R15077 vdd.n2187 vdd.t27 303.69
R15078 vdd.n1162 vdd.t57 303.69
R15079 vdd.n1122 vdd.t72 303.69
R15080 vdd.n406 vdd.t48 303.69
R15081 vdd.n420 vdd.t81 303.69
R15082 vdd.n432 vdd.t87 303.69
R15083 vdd.n724 vdd.t29 303.69
R15084 vdd.n687 vdd.t39 303.69
R15085 vdd.n3106 vdd.t22 303.69
R15086 vdd.n2853 vdd.n898 291.221
R15087 vdd.n3067 vdd.n778 291.221
R15088 vdd.n3004 vdd.n775 291.221
R15089 vdd.n2785 vdd.n2784 291.221
R15090 vdd.n2581 vdd.n940 291.221
R15091 vdd.n2512 vdd.n2511 291.221
R15092 vdd.n1280 vdd.n1279 291.221
R15093 vdd.n2332 vdd.n1046 291.221
R15094 vdd.n2983 vdd.n776 291.221
R15095 vdd.n3070 vdd.n3069 291.221
R15096 vdd.n2689 vdd.n2615 291.221
R15097 vdd.n2857 vdd.n902 291.221
R15098 vdd.n2509 vdd.n950 291.221
R15099 vdd.n948 vdd.n922 291.221
R15100 vdd.n1358 vdd.n1087 291.221
R15101 vdd.n2336 vdd.n1051 291.221
R15102 vdd.n2985 vdd.n776 185
R15103 vdd.n3068 vdd.n776 185
R15104 vdd.n2987 vdd.n2986 185
R15105 vdd.n2986 vdd.n774 185
R15106 vdd.n2988 vdd.n810 185
R15107 vdd.n2998 vdd.n810 185
R15108 vdd.n2989 vdd.n819 185
R15109 vdd.n819 vdd.n817 185
R15110 vdd.n2991 vdd.n2990 185
R15111 vdd.n2992 vdd.n2991 185
R15112 vdd.n2944 vdd.n818 185
R15113 vdd.n818 vdd.n814 185
R15114 vdd.n2943 vdd.n2942 185
R15115 vdd.n2942 vdd.n2941 185
R15116 vdd.n821 vdd.n820 185
R15117 vdd.n822 vdd.n821 185
R15118 vdd.n2934 vdd.n2933 185
R15119 vdd.n2935 vdd.n2934 185
R15120 vdd.n2932 vdd.n831 185
R15121 vdd.n831 vdd.n828 185
R15122 vdd.n2931 vdd.n2930 185
R15123 vdd.n2930 vdd.n2929 185
R15124 vdd.n833 vdd.n832 185
R15125 vdd.n841 vdd.n833 185
R15126 vdd.n2922 vdd.n2921 185
R15127 vdd.n2923 vdd.n2922 185
R15128 vdd.n2919 vdd.n842 185
R15129 vdd.n849 vdd.n842 185
R15130 vdd.n2918 vdd.n2917 185
R15131 vdd.n2917 vdd.n2916 185
R15132 vdd.n845 vdd.n844 185
R15133 vdd.n846 vdd.n845 185
R15134 vdd.n2909 vdd.n2908 185
R15135 vdd.n2910 vdd.n2909 185
R15136 vdd.n2907 vdd.n856 185
R15137 vdd.n856 vdd.n853 185
R15138 vdd.n2906 vdd.n2905 185
R15139 vdd.n2905 vdd.n2904 185
R15140 vdd.n858 vdd.n857 185
R15141 vdd.n866 vdd.n858 185
R15142 vdd.n2897 vdd.n2896 185
R15143 vdd.n2898 vdd.n2897 185
R15144 vdd.n2895 vdd.n867 185
R15145 vdd.n872 vdd.n867 185
R15146 vdd.n2894 vdd.n2893 185
R15147 vdd.n2893 vdd.n2892 185
R15148 vdd.n869 vdd.n868 185
R15149 vdd.n2764 vdd.n869 185
R15150 vdd.n2885 vdd.n2884 185
R15151 vdd.n2886 vdd.n2885 185
R15152 vdd.n2883 vdd.n879 185
R15153 vdd.n879 vdd.n876 185
R15154 vdd.n2882 vdd.n2881 185
R15155 vdd.n2881 vdd.n2880 185
R15156 vdd.n881 vdd.n880 185
R15157 vdd.n882 vdd.n881 185
R15158 vdd.n2873 vdd.n2872 185
R15159 vdd.n2874 vdd.n2873 185
R15160 vdd.n2871 vdd.n891 185
R15161 vdd.n891 vdd.n888 185
R15162 vdd.n2870 vdd.n2869 185
R15163 vdd.n2869 vdd.n2868 185
R15164 vdd.n893 vdd.n892 185
R15165 vdd.n2779 vdd.n893 185
R15166 vdd.n2861 vdd.n2860 185
R15167 vdd.n2862 vdd.n2861 185
R15168 vdd.n2859 vdd.n902 185
R15169 vdd.n902 vdd.n899 185
R15170 vdd.n2858 vdd.n2857 185
R15171 vdd.n904 vdd.n903 185
R15172 vdd.n2625 vdd.n2624 185
R15173 vdd.n2627 vdd.n2626 185
R15174 vdd.n2629 vdd.n2628 185
R15175 vdd.n2631 vdd.n2630 185
R15176 vdd.n2633 vdd.n2632 185
R15177 vdd.n2635 vdd.n2634 185
R15178 vdd.n2637 vdd.n2636 185
R15179 vdd.n2639 vdd.n2638 185
R15180 vdd.n2641 vdd.n2640 185
R15181 vdd.n2643 vdd.n2642 185
R15182 vdd.n2645 vdd.n2644 185
R15183 vdd.n2647 vdd.n2646 185
R15184 vdd.n2649 vdd.n2648 185
R15185 vdd.n2651 vdd.n2650 185
R15186 vdd.n2653 vdd.n2652 185
R15187 vdd.n2655 vdd.n2654 185
R15188 vdd.n2657 vdd.n2656 185
R15189 vdd.n2659 vdd.n2658 185
R15190 vdd.n2661 vdd.n2660 185
R15191 vdd.n2663 vdd.n2662 185
R15192 vdd.n2665 vdd.n2664 185
R15193 vdd.n2667 vdd.n2666 185
R15194 vdd.n2669 vdd.n2668 185
R15195 vdd.n2671 vdd.n2670 185
R15196 vdd.n2673 vdd.n2672 185
R15197 vdd.n2675 vdd.n2674 185
R15198 vdd.n2677 vdd.n2676 185
R15199 vdd.n2679 vdd.n2678 185
R15200 vdd.n2681 vdd.n2680 185
R15201 vdd.n2683 vdd.n2682 185
R15202 vdd.n2685 vdd.n2684 185
R15203 vdd.n2687 vdd.n2686 185
R15204 vdd.n2688 vdd.n2615 185
R15205 vdd.n2855 vdd.n2615 185
R15206 vdd.n3071 vdd.n3070 185
R15207 vdd.n3072 vdd.n767 185
R15208 vdd.n3074 vdd.n3073 185
R15209 vdd.n3076 vdd.n765 185
R15210 vdd.n3078 vdd.n3077 185
R15211 vdd.n3079 vdd.n764 185
R15212 vdd.n3081 vdd.n3080 185
R15213 vdd.n3083 vdd.n762 185
R15214 vdd.n3085 vdd.n3084 185
R15215 vdd.n3086 vdd.n761 185
R15216 vdd.n3088 vdd.n3087 185
R15217 vdd.n3090 vdd.n759 185
R15218 vdd.n3092 vdd.n3091 185
R15219 vdd.n3093 vdd.n758 185
R15220 vdd.n3095 vdd.n3094 185
R15221 vdd.n3097 vdd.n757 185
R15222 vdd.n3098 vdd.n754 185
R15223 vdd.n3101 vdd.n3100 185
R15224 vdd.n755 vdd.n753 185
R15225 vdd.n2957 vdd.n2956 185
R15226 vdd.n2959 vdd.n2958 185
R15227 vdd.n2961 vdd.n2953 185
R15228 vdd.n2963 vdd.n2962 185
R15229 vdd.n2964 vdd.n2952 185
R15230 vdd.n2966 vdd.n2965 185
R15231 vdd.n2968 vdd.n2950 185
R15232 vdd.n2970 vdd.n2969 185
R15233 vdd.n2971 vdd.n2949 185
R15234 vdd.n2973 vdd.n2972 185
R15235 vdd.n2975 vdd.n2947 185
R15236 vdd.n2977 vdd.n2976 185
R15237 vdd.n2978 vdd.n2946 185
R15238 vdd.n2980 vdd.n2979 185
R15239 vdd.n2982 vdd.n2945 185
R15240 vdd.n2984 vdd.n2983 185
R15241 vdd.n2983 vdd.n756 185
R15242 vdd.n3069 vdd.n771 185
R15243 vdd.n3069 vdd.n3068 185
R15244 vdd.n2692 vdd.n773 185
R15245 vdd.n774 vdd.n773 185
R15246 vdd.n2693 vdd.n809 185
R15247 vdd.n2998 vdd.n809 185
R15248 vdd.n2695 vdd.n2694 185
R15249 vdd.n2694 vdd.n817 185
R15250 vdd.n2696 vdd.n816 185
R15251 vdd.n2992 vdd.n816 185
R15252 vdd.n2698 vdd.n2697 185
R15253 vdd.n2697 vdd.n814 185
R15254 vdd.n2699 vdd.n824 185
R15255 vdd.n2941 vdd.n824 185
R15256 vdd.n2701 vdd.n2700 185
R15257 vdd.n2700 vdd.n822 185
R15258 vdd.n2702 vdd.n830 185
R15259 vdd.n2935 vdd.n830 185
R15260 vdd.n2704 vdd.n2703 185
R15261 vdd.n2703 vdd.n828 185
R15262 vdd.n2705 vdd.n835 185
R15263 vdd.n2929 vdd.n835 185
R15264 vdd.n2707 vdd.n2706 185
R15265 vdd.n2706 vdd.n841 185
R15266 vdd.n2708 vdd.n840 185
R15267 vdd.n2923 vdd.n840 185
R15268 vdd.n2710 vdd.n2709 185
R15269 vdd.n2709 vdd.n849 185
R15270 vdd.n2711 vdd.n848 185
R15271 vdd.n2916 vdd.n848 185
R15272 vdd.n2713 vdd.n2712 185
R15273 vdd.n2712 vdd.n846 185
R15274 vdd.n2714 vdd.n855 185
R15275 vdd.n2910 vdd.n855 185
R15276 vdd.n2716 vdd.n2715 185
R15277 vdd.n2715 vdd.n853 185
R15278 vdd.n2717 vdd.n860 185
R15279 vdd.n2904 vdd.n860 185
R15280 vdd.n2719 vdd.n2718 185
R15281 vdd.n2718 vdd.n866 185
R15282 vdd.n2720 vdd.n865 185
R15283 vdd.n2898 vdd.n865 185
R15284 vdd.n2722 vdd.n2721 185
R15285 vdd.n2721 vdd.n872 185
R15286 vdd.n2723 vdd.n871 185
R15287 vdd.n2892 vdd.n871 185
R15288 vdd.n2766 vdd.n2765 185
R15289 vdd.n2765 vdd.n2764 185
R15290 vdd.n2767 vdd.n878 185
R15291 vdd.n2886 vdd.n878 185
R15292 vdd.n2769 vdd.n2768 185
R15293 vdd.n2768 vdd.n876 185
R15294 vdd.n2770 vdd.n884 185
R15295 vdd.n2880 vdd.n884 185
R15296 vdd.n2772 vdd.n2771 185
R15297 vdd.n2771 vdd.n882 185
R15298 vdd.n2773 vdd.n890 185
R15299 vdd.n2874 vdd.n890 185
R15300 vdd.n2775 vdd.n2774 185
R15301 vdd.n2774 vdd.n888 185
R15302 vdd.n2776 vdd.n895 185
R15303 vdd.n2868 vdd.n895 185
R15304 vdd.n2778 vdd.n2777 185
R15305 vdd.n2779 vdd.n2778 185
R15306 vdd.n2691 vdd.n901 185
R15307 vdd.n2862 vdd.n901 185
R15308 vdd.n2690 vdd.n2689 185
R15309 vdd.n2689 vdd.n899 185
R15310 vdd.n2181 vdd.n2180 185
R15311 vdd.n2182 vdd.n2181 185
R15312 vdd.n1410 vdd.n1408 185
R15313 vdd.n1408 vdd.n1407 185
R15314 vdd.n2176 vdd.n2175 185
R15315 vdd.n2175 vdd.n2174 185
R15316 vdd.n1413 vdd.n1412 185
R15317 vdd.n1414 vdd.n1413 185
R15318 vdd.n2163 vdd.n2162 185
R15319 vdd.n2164 vdd.n2163 185
R15320 vdd.n1422 vdd.n1421 185
R15321 vdd.n2155 vdd.n1421 185
R15322 vdd.n2158 vdd.n2157 185
R15323 vdd.n2157 vdd.n2156 185
R15324 vdd.n1425 vdd.n1424 185
R15325 vdd.n1431 vdd.n1425 185
R15326 vdd.n2146 vdd.n2145 185
R15327 vdd.n2147 vdd.n2146 185
R15328 vdd.n1433 vdd.n1432 185
R15329 vdd.n2138 vdd.n1432 185
R15330 vdd.n2141 vdd.n2140 185
R15331 vdd.n2140 vdd.n2139 185
R15332 vdd.n1436 vdd.n1435 185
R15333 vdd.n1437 vdd.n1436 185
R15334 vdd.n2129 vdd.n2128 185
R15335 vdd.n2130 vdd.n2129 185
R15336 vdd.n1445 vdd.n1444 185
R15337 vdd.n1444 vdd.n1443 185
R15338 vdd.n2124 vdd.n2123 185
R15339 vdd.n2123 vdd.n2122 185
R15340 vdd.n1448 vdd.n1447 185
R15341 vdd.n1454 vdd.n1448 185
R15342 vdd.n2113 vdd.n2112 185
R15343 vdd.n2114 vdd.n2113 185
R15344 vdd.n1456 vdd.n1455 185
R15345 vdd.n1810 vdd.n1455 185
R15346 vdd.n1813 vdd.n1812 185
R15347 vdd.n1812 vdd.n1811 185
R15348 vdd.n1459 vdd.n1458 185
R15349 vdd.n1466 vdd.n1459 185
R15350 vdd.n1801 vdd.n1800 185
R15351 vdd.n1802 vdd.n1801 185
R15352 vdd.n1468 vdd.n1467 185
R15353 vdd.n1467 vdd.n1465 185
R15354 vdd.n1796 vdd.n1795 185
R15355 vdd.n1795 vdd.n1794 185
R15356 vdd.n1471 vdd.n1470 185
R15357 vdd.n1472 vdd.n1471 185
R15358 vdd.n1785 vdd.n1784 185
R15359 vdd.n1786 vdd.n1785 185
R15360 vdd.n1479 vdd.n1478 185
R15361 vdd.n1777 vdd.n1478 185
R15362 vdd.n1780 vdd.n1779 185
R15363 vdd.n1779 vdd.n1778 185
R15364 vdd.n1482 vdd.n1481 185
R15365 vdd.n1488 vdd.n1482 185
R15366 vdd.n1768 vdd.n1767 185
R15367 vdd.n1769 vdd.n1768 185
R15368 vdd.n1490 vdd.n1489 185
R15369 vdd.n1760 vdd.n1489 185
R15370 vdd.n1763 vdd.n1762 185
R15371 vdd.n1762 vdd.n1761 185
R15372 vdd.n1493 vdd.n1492 185
R15373 vdd.n1494 vdd.n1493 185
R15374 vdd.n1751 vdd.n1750 185
R15375 vdd.n1752 vdd.n1751 185
R15376 vdd.n1502 vdd.n1501 185
R15377 vdd.n1501 vdd.n1500 185
R15378 vdd.n1746 vdd.n1745 185
R15379 vdd.n1745 vdd.n1744 185
R15380 vdd.n1505 vdd.n1504 185
R15381 vdd.n1506 vdd.n1505 185
R15382 vdd.n1734 vdd.n1733 185
R15383 vdd.n1732 vdd.n1545 185
R15384 vdd.n1547 vdd.n1544 185
R15385 vdd.n1736 vdd.n1544 185
R15386 vdd.n1728 vdd.n1549 185
R15387 vdd.n1727 vdd.n1550 185
R15388 vdd.n1726 vdd.n1551 185
R15389 vdd.n1554 vdd.n1552 185
R15390 vdd.n1722 vdd.n1555 185
R15391 vdd.n1721 vdd.n1556 185
R15392 vdd.n1720 vdd.n1557 185
R15393 vdd.n1560 vdd.n1558 185
R15394 vdd.n1716 vdd.n1561 185
R15395 vdd.n1715 vdd.n1562 185
R15396 vdd.n1714 vdd.n1563 185
R15397 vdd.n1566 vdd.n1564 185
R15398 vdd.n1710 vdd.n1567 185
R15399 vdd.n1709 vdd.n1568 185
R15400 vdd.n1708 vdd.n1569 185
R15401 vdd.n1700 vdd.n1570 185
R15402 vdd.n1704 vdd.n1701 185
R15403 vdd.n1699 vdd.n1572 185
R15404 vdd.n1698 vdd.n1573 185
R15405 vdd.n1576 vdd.n1574 185
R15406 vdd.n1694 vdd.n1577 185
R15407 vdd.n1693 vdd.n1578 185
R15408 vdd.n1692 vdd.n1579 185
R15409 vdd.n1582 vdd.n1580 185
R15410 vdd.n1688 vdd.n1583 185
R15411 vdd.n1687 vdd.n1584 185
R15412 vdd.n1686 vdd.n1585 185
R15413 vdd.n1588 vdd.n1586 185
R15414 vdd.n1682 vdd.n1589 185
R15415 vdd.n1681 vdd.n1590 185
R15416 vdd.n1680 vdd.n1591 185
R15417 vdd.n1594 vdd.n1592 185
R15418 vdd.n1676 vdd.n1595 185
R15419 vdd.n1675 vdd.n1596 185
R15420 vdd.n1674 vdd.n1597 185
R15421 vdd.n1600 vdd.n1598 185
R15422 vdd.n1670 vdd.n1601 185
R15423 vdd.n1669 vdd.n1602 185
R15424 vdd.n1668 vdd.n1665 185
R15425 vdd.n1605 vdd.n1603 185
R15426 vdd.n1661 vdd.n1606 185
R15427 vdd.n1660 vdd.n1607 185
R15428 vdd.n1659 vdd.n1608 185
R15429 vdd.n1611 vdd.n1609 185
R15430 vdd.n1655 vdd.n1612 185
R15431 vdd.n1654 vdd.n1613 185
R15432 vdd.n1653 vdd.n1614 185
R15433 vdd.n1617 vdd.n1615 185
R15434 vdd.n1649 vdd.n1618 185
R15435 vdd.n1648 vdd.n1619 185
R15436 vdd.n1647 vdd.n1620 185
R15437 vdd.n1623 vdd.n1621 185
R15438 vdd.n1643 vdd.n1624 185
R15439 vdd.n1642 vdd.n1625 185
R15440 vdd.n1641 vdd.n1626 185
R15441 vdd.n1629 vdd.n1627 185
R15442 vdd.n1637 vdd.n1630 185
R15443 vdd.n1636 vdd.n1631 185
R15444 vdd.n1635 vdd.n1632 185
R15445 vdd.n1633 vdd.n1513 185
R15446 vdd.n1738 vdd.n1737 185
R15447 vdd.n1737 vdd.n1736 185
R15448 vdd.n2185 vdd.n2184 185
R15449 vdd.n2189 vdd.n1403 185
R15450 vdd.n1402 vdd.n1396 185
R15451 vdd.n1400 vdd.n1399 185
R15452 vdd.n1398 vdd.n1192 185
R15453 vdd.n2193 vdd.n1189 185
R15454 vdd.n2195 vdd.n2194 185
R15455 vdd.n2197 vdd.n1187 185
R15456 vdd.n2199 vdd.n2198 185
R15457 vdd.n2200 vdd.n1182 185
R15458 vdd.n2202 vdd.n2201 185
R15459 vdd.n2204 vdd.n1180 185
R15460 vdd.n2206 vdd.n2205 185
R15461 vdd.n2207 vdd.n1175 185
R15462 vdd.n2209 vdd.n2208 185
R15463 vdd.n2211 vdd.n1173 185
R15464 vdd.n2213 vdd.n2212 185
R15465 vdd.n2214 vdd.n1169 185
R15466 vdd.n2216 vdd.n2215 185
R15467 vdd.n2218 vdd.n1166 185
R15468 vdd.n2220 vdd.n2219 185
R15469 vdd.n1167 vdd.n1160 185
R15470 vdd.n2224 vdd.n1164 185
R15471 vdd.n2225 vdd.n1156 185
R15472 vdd.n2227 vdd.n2226 185
R15473 vdd.n2229 vdd.n1154 185
R15474 vdd.n2231 vdd.n2230 185
R15475 vdd.n2232 vdd.n1149 185
R15476 vdd.n2234 vdd.n2233 185
R15477 vdd.n2236 vdd.n1147 185
R15478 vdd.n2238 vdd.n2237 185
R15479 vdd.n2239 vdd.n1142 185
R15480 vdd.n2241 vdd.n2240 185
R15481 vdd.n2243 vdd.n1140 185
R15482 vdd.n2245 vdd.n2244 185
R15483 vdd.n2246 vdd.n1135 185
R15484 vdd.n2248 vdd.n2247 185
R15485 vdd.n2250 vdd.n1133 185
R15486 vdd.n2252 vdd.n2251 185
R15487 vdd.n2253 vdd.n1129 185
R15488 vdd.n2255 vdd.n2254 185
R15489 vdd.n2257 vdd.n1126 185
R15490 vdd.n2259 vdd.n2258 185
R15491 vdd.n1127 vdd.n1120 185
R15492 vdd.n2263 vdd.n1124 185
R15493 vdd.n2264 vdd.n1116 185
R15494 vdd.n2266 vdd.n2265 185
R15495 vdd.n2268 vdd.n1114 185
R15496 vdd.n2270 vdd.n2269 185
R15497 vdd.n2271 vdd.n1109 185
R15498 vdd.n2273 vdd.n2272 185
R15499 vdd.n2275 vdd.n1107 185
R15500 vdd.n2277 vdd.n2276 185
R15501 vdd.n2278 vdd.n1102 185
R15502 vdd.n2280 vdd.n2279 185
R15503 vdd.n2282 vdd.n1100 185
R15504 vdd.n2284 vdd.n2283 185
R15505 vdd.n2285 vdd.n1098 185
R15506 vdd.n2287 vdd.n2286 185
R15507 vdd.n2290 vdd.n2289 185
R15508 vdd.n2292 vdd.n2291 185
R15509 vdd.n2294 vdd.n1096 185
R15510 vdd.n2296 vdd.n2295 185
R15511 vdd.n1409 vdd.n1095 185
R15512 vdd.n2183 vdd.n1406 185
R15513 vdd.n2183 vdd.n2182 185
R15514 vdd.n1417 vdd.n1405 185
R15515 vdd.n1407 vdd.n1405 185
R15516 vdd.n2173 vdd.n2172 185
R15517 vdd.n2174 vdd.n2173 185
R15518 vdd.n1416 vdd.n1415 185
R15519 vdd.n1415 vdd.n1414 185
R15520 vdd.n2166 vdd.n2165 185
R15521 vdd.n2165 vdd.n2164 185
R15522 vdd.n1420 vdd.n1419 185
R15523 vdd.n2155 vdd.n1420 185
R15524 vdd.n2154 vdd.n2153 185
R15525 vdd.n2156 vdd.n2154 185
R15526 vdd.n1427 vdd.n1426 185
R15527 vdd.n1431 vdd.n1426 185
R15528 vdd.n2149 vdd.n2148 185
R15529 vdd.n2148 vdd.n2147 185
R15530 vdd.n1430 vdd.n1429 185
R15531 vdd.n2138 vdd.n1430 185
R15532 vdd.n2137 vdd.n2136 185
R15533 vdd.n2139 vdd.n2137 185
R15534 vdd.n1439 vdd.n1438 185
R15535 vdd.n1438 vdd.n1437 185
R15536 vdd.n2132 vdd.n2131 185
R15537 vdd.n2131 vdd.n2130 185
R15538 vdd.n1442 vdd.n1441 185
R15539 vdd.n1443 vdd.n1442 185
R15540 vdd.n2121 vdd.n2120 185
R15541 vdd.n2122 vdd.n2121 185
R15542 vdd.n1450 vdd.n1449 185
R15543 vdd.n1454 vdd.n1449 185
R15544 vdd.n2116 vdd.n2115 185
R15545 vdd.n2115 vdd.n2114 185
R15546 vdd.n1453 vdd.n1452 185
R15547 vdd.n1810 vdd.n1453 185
R15548 vdd.n1809 vdd.n1808 185
R15549 vdd.n1811 vdd.n1809 185
R15550 vdd.n1461 vdd.n1460 185
R15551 vdd.n1466 vdd.n1460 185
R15552 vdd.n1804 vdd.n1803 185
R15553 vdd.n1803 vdd.n1802 185
R15554 vdd.n1464 vdd.n1463 185
R15555 vdd.n1465 vdd.n1464 185
R15556 vdd.n1793 vdd.n1792 185
R15557 vdd.n1794 vdd.n1793 185
R15558 vdd.n1474 vdd.n1473 185
R15559 vdd.n1473 vdd.n1472 185
R15560 vdd.n1788 vdd.n1787 185
R15561 vdd.n1787 vdd.n1786 185
R15562 vdd.n1477 vdd.n1476 185
R15563 vdd.n1777 vdd.n1477 185
R15564 vdd.n1776 vdd.n1775 185
R15565 vdd.n1778 vdd.n1776 185
R15566 vdd.n1484 vdd.n1483 185
R15567 vdd.n1488 vdd.n1483 185
R15568 vdd.n1771 vdd.n1770 185
R15569 vdd.n1770 vdd.n1769 185
R15570 vdd.n1487 vdd.n1486 185
R15571 vdd.n1760 vdd.n1487 185
R15572 vdd.n1759 vdd.n1758 185
R15573 vdd.n1761 vdd.n1759 185
R15574 vdd.n1496 vdd.n1495 185
R15575 vdd.n1495 vdd.n1494 185
R15576 vdd.n1754 vdd.n1753 185
R15577 vdd.n1753 vdd.n1752 185
R15578 vdd.n1499 vdd.n1498 185
R15579 vdd.n1500 vdd.n1499 185
R15580 vdd.n1743 vdd.n1742 185
R15581 vdd.n1744 vdd.n1743 185
R15582 vdd.n1508 vdd.n1507 185
R15583 vdd.n1507 vdd.n1506 185
R15584 vdd.n942 vdd.n940 185
R15585 vdd.n2510 vdd.n940 185
R15586 vdd.n2432 vdd.n960 185
R15587 vdd.n960 vdd.n947 185
R15588 vdd.n2434 vdd.n2433 185
R15589 vdd.n2435 vdd.n2434 185
R15590 vdd.n2431 vdd.n959 185
R15591 vdd.n1309 vdd.n959 185
R15592 vdd.n2430 vdd.n2429 185
R15593 vdd.n2429 vdd.n2428 185
R15594 vdd.n962 vdd.n961 185
R15595 vdd.n963 vdd.n962 185
R15596 vdd.n2419 vdd.n2418 185
R15597 vdd.n2420 vdd.n2419 185
R15598 vdd.n2417 vdd.n973 185
R15599 vdd.n973 vdd.n970 185
R15600 vdd.n2416 vdd.n2415 185
R15601 vdd.n2415 vdd.n2414 185
R15602 vdd.n975 vdd.n974 185
R15603 vdd.n976 vdd.n975 185
R15604 vdd.n2407 vdd.n2406 185
R15605 vdd.n2408 vdd.n2407 185
R15606 vdd.n2405 vdd.n984 185
R15607 vdd.n989 vdd.n984 185
R15608 vdd.n2404 vdd.n2403 185
R15609 vdd.n2403 vdd.n2402 185
R15610 vdd.n986 vdd.n985 185
R15611 vdd.n995 vdd.n986 185
R15612 vdd.n2395 vdd.n2394 185
R15613 vdd.n2396 vdd.n2395 185
R15614 vdd.n2393 vdd.n996 185
R15615 vdd.n1330 vdd.n996 185
R15616 vdd.n2392 vdd.n2391 185
R15617 vdd.n2391 vdd.n2390 185
R15618 vdd.n998 vdd.n997 185
R15619 vdd.n999 vdd.n998 185
R15620 vdd.n2383 vdd.n2382 185
R15621 vdd.n2384 vdd.n2383 185
R15622 vdd.n2381 vdd.n1008 185
R15623 vdd.n1008 vdd.n1005 185
R15624 vdd.n2380 vdd.n2379 185
R15625 vdd.n2379 vdd.n2378 185
R15626 vdd.n1010 vdd.n1009 185
R15627 vdd.n1019 vdd.n1010 185
R15628 vdd.n2370 vdd.n2369 185
R15629 vdd.n2371 vdd.n2370 185
R15630 vdd.n2368 vdd.n1020 185
R15631 vdd.n1026 vdd.n1020 185
R15632 vdd.n2367 vdd.n2366 185
R15633 vdd.n2366 vdd.n2365 185
R15634 vdd.n1022 vdd.n1021 185
R15635 vdd.n1023 vdd.n1022 185
R15636 vdd.n2358 vdd.n2357 185
R15637 vdd.n2359 vdd.n2358 185
R15638 vdd.n2356 vdd.n1033 185
R15639 vdd.n1033 vdd.n1030 185
R15640 vdd.n2355 vdd.n2354 185
R15641 vdd.n2354 vdd.n2353 185
R15642 vdd.n1035 vdd.n1034 185
R15643 vdd.n1036 vdd.n1035 185
R15644 vdd.n2346 vdd.n2345 185
R15645 vdd.n2347 vdd.n2346 185
R15646 vdd.n2344 vdd.n1044 185
R15647 vdd.n1050 vdd.n1044 185
R15648 vdd.n2343 vdd.n2342 185
R15649 vdd.n2342 vdd.n2341 185
R15650 vdd.n1046 vdd.n1045 185
R15651 vdd.n1047 vdd.n1046 185
R15652 vdd.n2332 vdd.n2331 185
R15653 vdd.n2330 vdd.n1089 185
R15654 vdd.n2329 vdd.n1088 185
R15655 vdd.n2334 vdd.n1088 185
R15656 vdd.n2328 vdd.n2327 185
R15657 vdd.n2326 vdd.n2325 185
R15658 vdd.n2324 vdd.n2323 185
R15659 vdd.n2322 vdd.n2321 185
R15660 vdd.n2320 vdd.n2319 185
R15661 vdd.n2318 vdd.n2317 185
R15662 vdd.n2316 vdd.n2315 185
R15663 vdd.n2314 vdd.n2313 185
R15664 vdd.n2312 vdd.n2311 185
R15665 vdd.n2310 vdd.n2309 185
R15666 vdd.n2308 vdd.n2307 185
R15667 vdd.n2306 vdd.n2305 185
R15668 vdd.n2304 vdd.n2303 185
R15669 vdd.n2302 vdd.n2301 185
R15670 vdd.n2300 vdd.n2299 185
R15671 vdd.n1246 vdd.n1090 185
R15672 vdd.n1248 vdd.n1247 185
R15673 vdd.n1250 vdd.n1249 185
R15674 vdd.n1252 vdd.n1251 185
R15675 vdd.n1254 vdd.n1253 185
R15676 vdd.n1256 vdd.n1255 185
R15677 vdd.n1258 vdd.n1257 185
R15678 vdd.n1260 vdd.n1259 185
R15679 vdd.n1262 vdd.n1261 185
R15680 vdd.n1264 vdd.n1263 185
R15681 vdd.n1266 vdd.n1265 185
R15682 vdd.n1268 vdd.n1267 185
R15683 vdd.n1270 vdd.n1269 185
R15684 vdd.n1272 vdd.n1271 185
R15685 vdd.n1275 vdd.n1274 185
R15686 vdd.n1277 vdd.n1276 185
R15687 vdd.n1279 vdd.n1278 185
R15688 vdd.n2513 vdd.n2512 185
R15689 vdd.n2515 vdd.n2514 185
R15690 vdd.n2517 vdd.n2516 185
R15691 vdd.n2520 vdd.n2519 185
R15692 vdd.n2522 vdd.n2521 185
R15693 vdd.n2524 vdd.n2523 185
R15694 vdd.n2526 vdd.n2525 185
R15695 vdd.n2528 vdd.n2527 185
R15696 vdd.n2530 vdd.n2529 185
R15697 vdd.n2532 vdd.n2531 185
R15698 vdd.n2534 vdd.n2533 185
R15699 vdd.n2536 vdd.n2535 185
R15700 vdd.n2538 vdd.n2537 185
R15701 vdd.n2540 vdd.n2539 185
R15702 vdd.n2542 vdd.n2541 185
R15703 vdd.n2544 vdd.n2543 185
R15704 vdd.n2546 vdd.n2545 185
R15705 vdd.n2548 vdd.n2547 185
R15706 vdd.n2550 vdd.n2549 185
R15707 vdd.n2552 vdd.n2551 185
R15708 vdd.n2554 vdd.n2553 185
R15709 vdd.n2556 vdd.n2555 185
R15710 vdd.n2558 vdd.n2557 185
R15711 vdd.n2560 vdd.n2559 185
R15712 vdd.n2562 vdd.n2561 185
R15713 vdd.n2564 vdd.n2563 185
R15714 vdd.n2566 vdd.n2565 185
R15715 vdd.n2568 vdd.n2567 185
R15716 vdd.n2570 vdd.n2569 185
R15717 vdd.n2572 vdd.n2571 185
R15718 vdd.n2574 vdd.n2573 185
R15719 vdd.n2576 vdd.n2575 185
R15720 vdd.n2578 vdd.n2577 185
R15721 vdd.n2579 vdd.n941 185
R15722 vdd.n2581 vdd.n2580 185
R15723 vdd.n2582 vdd.n2581 185
R15724 vdd.n2511 vdd.n945 185
R15725 vdd.n2511 vdd.n2510 185
R15726 vdd.n1307 vdd.n946 185
R15727 vdd.n947 vdd.n946 185
R15728 vdd.n1308 vdd.n957 185
R15729 vdd.n2435 vdd.n957 185
R15730 vdd.n1311 vdd.n1310 185
R15731 vdd.n1310 vdd.n1309 185
R15732 vdd.n1312 vdd.n964 185
R15733 vdd.n2428 vdd.n964 185
R15734 vdd.n1314 vdd.n1313 185
R15735 vdd.n1313 vdd.n963 185
R15736 vdd.n1315 vdd.n971 185
R15737 vdd.n2420 vdd.n971 185
R15738 vdd.n1317 vdd.n1316 185
R15739 vdd.n1316 vdd.n970 185
R15740 vdd.n1318 vdd.n977 185
R15741 vdd.n2414 vdd.n977 185
R15742 vdd.n1320 vdd.n1319 185
R15743 vdd.n1319 vdd.n976 185
R15744 vdd.n1321 vdd.n982 185
R15745 vdd.n2408 vdd.n982 185
R15746 vdd.n1323 vdd.n1322 185
R15747 vdd.n1322 vdd.n989 185
R15748 vdd.n1324 vdd.n987 185
R15749 vdd.n2402 vdd.n987 185
R15750 vdd.n1326 vdd.n1325 185
R15751 vdd.n1325 vdd.n995 185
R15752 vdd.n1327 vdd.n993 185
R15753 vdd.n2396 vdd.n993 185
R15754 vdd.n1329 vdd.n1328 185
R15755 vdd.n1330 vdd.n1329 185
R15756 vdd.n1306 vdd.n1000 185
R15757 vdd.n2390 vdd.n1000 185
R15758 vdd.n1305 vdd.n1304 185
R15759 vdd.n1304 vdd.n999 185
R15760 vdd.n1303 vdd.n1006 185
R15761 vdd.n2384 vdd.n1006 185
R15762 vdd.n1302 vdd.n1301 185
R15763 vdd.n1301 vdd.n1005 185
R15764 vdd.n1300 vdd.n1011 185
R15765 vdd.n2378 vdd.n1011 185
R15766 vdd.n1299 vdd.n1298 185
R15767 vdd.n1298 vdd.n1019 185
R15768 vdd.n1297 vdd.n1017 185
R15769 vdd.n2371 vdd.n1017 185
R15770 vdd.n1296 vdd.n1295 185
R15771 vdd.n1295 vdd.n1026 185
R15772 vdd.n1294 vdd.n1024 185
R15773 vdd.n2365 vdd.n1024 185
R15774 vdd.n1293 vdd.n1292 185
R15775 vdd.n1292 vdd.n1023 185
R15776 vdd.n1291 vdd.n1031 185
R15777 vdd.n2359 vdd.n1031 185
R15778 vdd.n1290 vdd.n1289 185
R15779 vdd.n1289 vdd.n1030 185
R15780 vdd.n1288 vdd.n1037 185
R15781 vdd.n2353 vdd.n1037 185
R15782 vdd.n1287 vdd.n1286 185
R15783 vdd.n1286 vdd.n1036 185
R15784 vdd.n1285 vdd.n1042 185
R15785 vdd.n2347 vdd.n1042 185
R15786 vdd.n1284 vdd.n1283 185
R15787 vdd.n1283 vdd.n1050 185
R15788 vdd.n1282 vdd.n1048 185
R15789 vdd.n2341 vdd.n1048 185
R15790 vdd.n1281 vdd.n1280 185
R15791 vdd.n1280 vdd.n1047 185
R15792 vdd.n370 vdd.n369 185
R15793 vdd.n3346 vdd.n370 185
R15794 vdd.n3349 vdd.n3348 185
R15795 vdd.n3348 vdd.n3347 185
R15796 vdd.n3350 vdd.n364 185
R15797 vdd.n364 vdd.n363 185
R15798 vdd.n3352 vdd.n3351 185
R15799 vdd.n3353 vdd.n3352 185
R15800 vdd.n359 vdd.n358 185
R15801 vdd.n3354 vdd.n359 185
R15802 vdd.n3357 vdd.n3356 185
R15803 vdd.n3356 vdd.n3355 185
R15804 vdd.n3358 vdd.n353 185
R15805 vdd.n3328 vdd.n353 185
R15806 vdd.n3360 vdd.n3359 185
R15807 vdd.n3361 vdd.n3360 185
R15808 vdd.n348 vdd.n347 185
R15809 vdd.n3362 vdd.n348 185
R15810 vdd.n3365 vdd.n3364 185
R15811 vdd.n3364 vdd.n3363 185
R15812 vdd.n3366 vdd.n342 185
R15813 vdd.n349 vdd.n342 185
R15814 vdd.n3368 vdd.n3367 185
R15815 vdd.n3369 vdd.n3368 185
R15816 vdd.n338 vdd.n337 185
R15817 vdd.n3370 vdd.n338 185
R15818 vdd.n3373 vdd.n3372 185
R15819 vdd.n3372 vdd.n3371 185
R15820 vdd.n3374 vdd.n333 185
R15821 vdd.n333 vdd.n332 185
R15822 vdd.n3376 vdd.n3375 185
R15823 vdd.n3377 vdd.n3376 185
R15824 vdd.n327 vdd.n325 185
R15825 vdd.n3378 vdd.n327 185
R15826 vdd.n3381 vdd.n3380 185
R15827 vdd.n3380 vdd.n3379 185
R15828 vdd.n326 vdd.n324 185
R15829 vdd.n328 vdd.n326 185
R15830 vdd.n3304 vdd.n3303 185
R15831 vdd.n3305 vdd.n3304 185
R15832 vdd.n615 vdd.n614 185
R15833 vdd.n614 vdd.n613 185
R15834 vdd.n3299 vdd.n3298 185
R15835 vdd.n3298 vdd.n3297 185
R15836 vdd.n618 vdd.n617 185
R15837 vdd.n624 vdd.n618 185
R15838 vdd.n3285 vdd.n3284 185
R15839 vdd.n3286 vdd.n3285 185
R15840 vdd.n626 vdd.n625 185
R15841 vdd.n3277 vdd.n625 185
R15842 vdd.n3280 vdd.n3279 185
R15843 vdd.n3279 vdd.n3278 185
R15844 vdd.n629 vdd.n628 185
R15845 vdd.n636 vdd.n629 185
R15846 vdd.n3268 vdd.n3267 185
R15847 vdd.n3269 vdd.n3268 185
R15848 vdd.n638 vdd.n637 185
R15849 vdd.n637 vdd.n635 185
R15850 vdd.n3263 vdd.n3262 185
R15851 vdd.n3262 vdd.n3261 185
R15852 vdd.n641 vdd.n640 185
R15853 vdd.n642 vdd.n641 185
R15854 vdd.n3252 vdd.n3251 185
R15855 vdd.n3253 vdd.n3252 185
R15856 vdd.n650 vdd.n649 185
R15857 vdd.n649 vdd.n648 185
R15858 vdd.n3247 vdd.n3246 185
R15859 vdd.n3246 vdd.n3245 185
R15860 vdd.n653 vdd.n652 185
R15861 vdd.n659 vdd.n653 185
R15862 vdd.n3236 vdd.n3235 185
R15863 vdd.n3237 vdd.n3236 185
R15864 vdd.n3232 vdd.n660 185
R15865 vdd.n3231 vdd.n3230 185
R15866 vdd.n3228 vdd.n662 185
R15867 vdd.n3228 vdd.n658 185
R15868 vdd.n3227 vdd.n3226 185
R15869 vdd.n3225 vdd.n3224 185
R15870 vdd.n3223 vdd.n3222 185
R15871 vdd.n3221 vdd.n3220 185
R15872 vdd.n3219 vdd.n668 185
R15873 vdd.n3217 vdd.n3216 185
R15874 vdd.n3215 vdd.n669 185
R15875 vdd.n3214 vdd.n3213 185
R15876 vdd.n3211 vdd.n674 185
R15877 vdd.n3209 vdd.n3208 185
R15878 vdd.n3207 vdd.n675 185
R15879 vdd.n3206 vdd.n3205 185
R15880 vdd.n3203 vdd.n680 185
R15881 vdd.n3201 vdd.n3200 185
R15882 vdd.n3199 vdd.n681 185
R15883 vdd.n3198 vdd.n3197 185
R15884 vdd.n3195 vdd.n688 185
R15885 vdd.n3193 vdd.n3192 185
R15886 vdd.n3191 vdd.n689 185
R15887 vdd.n3190 vdd.n3189 185
R15888 vdd.n3187 vdd.n694 185
R15889 vdd.n3185 vdd.n3184 185
R15890 vdd.n3183 vdd.n695 185
R15891 vdd.n3182 vdd.n3181 185
R15892 vdd.n3179 vdd.n700 185
R15893 vdd.n3177 vdd.n3176 185
R15894 vdd.n3175 vdd.n701 185
R15895 vdd.n3174 vdd.n3173 185
R15896 vdd.n3171 vdd.n706 185
R15897 vdd.n3169 vdd.n3168 185
R15898 vdd.n3167 vdd.n707 185
R15899 vdd.n3166 vdd.n3165 185
R15900 vdd.n3163 vdd.n712 185
R15901 vdd.n3161 vdd.n3160 185
R15902 vdd.n3159 vdd.n713 185
R15903 vdd.n3158 vdd.n3157 185
R15904 vdd.n3155 vdd.n718 185
R15905 vdd.n3153 vdd.n3152 185
R15906 vdd.n3151 vdd.n719 185
R15907 vdd.n728 vdd.n722 185
R15908 vdd.n3147 vdd.n3146 185
R15909 vdd.n3144 vdd.n726 185
R15910 vdd.n3143 vdd.n3142 185
R15911 vdd.n3141 vdd.n3140 185
R15912 vdd.n3139 vdd.n732 185
R15913 vdd.n3137 vdd.n3136 185
R15914 vdd.n3135 vdd.n733 185
R15915 vdd.n3134 vdd.n3133 185
R15916 vdd.n3131 vdd.n738 185
R15917 vdd.n3129 vdd.n3128 185
R15918 vdd.n3127 vdd.n739 185
R15919 vdd.n3126 vdd.n3125 185
R15920 vdd.n3123 vdd.n744 185
R15921 vdd.n3121 vdd.n3120 185
R15922 vdd.n3119 vdd.n745 185
R15923 vdd.n3118 vdd.n3117 185
R15924 vdd.n3115 vdd.n3114 185
R15925 vdd.n3113 vdd.n3112 185
R15926 vdd.n3111 vdd.n3110 185
R15927 vdd.n3109 vdd.n3108 185
R15928 vdd.n3104 vdd.n657 185
R15929 vdd.n658 vdd.n657 185
R15930 vdd.n3343 vdd.n3342 185
R15931 vdd.n599 vdd.n404 185
R15932 vdd.n598 vdd.n597 185
R15933 vdd.n596 vdd.n595 185
R15934 vdd.n594 vdd.n409 185
R15935 vdd.n590 vdd.n589 185
R15936 vdd.n588 vdd.n587 185
R15937 vdd.n586 vdd.n585 185
R15938 vdd.n584 vdd.n411 185
R15939 vdd.n580 vdd.n579 185
R15940 vdd.n578 vdd.n577 185
R15941 vdd.n576 vdd.n575 185
R15942 vdd.n574 vdd.n413 185
R15943 vdd.n570 vdd.n569 185
R15944 vdd.n568 vdd.n567 185
R15945 vdd.n566 vdd.n565 185
R15946 vdd.n564 vdd.n415 185
R15947 vdd.n560 vdd.n559 185
R15948 vdd.n558 vdd.n557 185
R15949 vdd.n556 vdd.n555 185
R15950 vdd.n554 vdd.n417 185
R15951 vdd.n550 vdd.n549 185
R15952 vdd.n548 vdd.n547 185
R15953 vdd.n546 vdd.n545 185
R15954 vdd.n544 vdd.n421 185
R15955 vdd.n540 vdd.n539 185
R15956 vdd.n538 vdd.n537 185
R15957 vdd.n536 vdd.n535 185
R15958 vdd.n534 vdd.n423 185
R15959 vdd.n530 vdd.n529 185
R15960 vdd.n528 vdd.n527 185
R15961 vdd.n526 vdd.n525 185
R15962 vdd.n524 vdd.n425 185
R15963 vdd.n520 vdd.n519 185
R15964 vdd.n518 vdd.n517 185
R15965 vdd.n516 vdd.n515 185
R15966 vdd.n514 vdd.n427 185
R15967 vdd.n510 vdd.n509 185
R15968 vdd.n508 vdd.n507 185
R15969 vdd.n506 vdd.n505 185
R15970 vdd.n504 vdd.n429 185
R15971 vdd.n500 vdd.n499 185
R15972 vdd.n498 vdd.n497 185
R15973 vdd.n496 vdd.n495 185
R15974 vdd.n494 vdd.n433 185
R15975 vdd.n490 vdd.n489 185
R15976 vdd.n488 vdd.n487 185
R15977 vdd.n486 vdd.n485 185
R15978 vdd.n484 vdd.n435 185
R15979 vdd.n480 vdd.n479 185
R15980 vdd.n478 vdd.n477 185
R15981 vdd.n476 vdd.n475 185
R15982 vdd.n474 vdd.n437 185
R15983 vdd.n470 vdd.n469 185
R15984 vdd.n468 vdd.n467 185
R15985 vdd.n466 vdd.n465 185
R15986 vdd.n464 vdd.n439 185
R15987 vdd.n460 vdd.n459 185
R15988 vdd.n458 vdd.n457 185
R15989 vdd.n456 vdd.n455 185
R15990 vdd.n454 vdd.n441 185
R15991 vdd.n450 vdd.n449 185
R15992 vdd.n448 vdd.n447 185
R15993 vdd.n446 vdd.n445 185
R15994 vdd.n3339 vdd.n372 185
R15995 vdd.n3346 vdd.n372 185
R15996 vdd.n3338 vdd.n371 185
R15997 vdd.n3347 vdd.n371 185
R15998 vdd.n3337 vdd.n3336 185
R15999 vdd.n3336 vdd.n363 185
R16000 vdd.n602 vdd.n362 185
R16001 vdd.n3353 vdd.n362 185
R16002 vdd.n3332 vdd.n361 185
R16003 vdd.n3354 vdd.n361 185
R16004 vdd.n3331 vdd.n360 185
R16005 vdd.n3355 vdd.n360 185
R16006 vdd.n3330 vdd.n3329 185
R16007 vdd.n3329 vdd.n3328 185
R16008 vdd.n604 vdd.n352 185
R16009 vdd.n3361 vdd.n352 185
R16010 vdd.n3324 vdd.n351 185
R16011 vdd.n3362 vdd.n351 185
R16012 vdd.n3323 vdd.n350 185
R16013 vdd.n3363 vdd.n350 185
R16014 vdd.n3322 vdd.n3321 185
R16015 vdd.n3321 vdd.n349 185
R16016 vdd.n606 vdd.n341 185
R16017 vdd.n3369 vdd.n341 185
R16018 vdd.n3317 vdd.n340 185
R16019 vdd.n3370 vdd.n340 185
R16020 vdd.n3316 vdd.n339 185
R16021 vdd.n3371 vdd.n339 185
R16022 vdd.n3315 vdd.n3314 185
R16023 vdd.n3314 vdd.n332 185
R16024 vdd.n608 vdd.n331 185
R16025 vdd.n3377 vdd.n331 185
R16026 vdd.n3310 vdd.n330 185
R16027 vdd.n3378 vdd.n330 185
R16028 vdd.n3309 vdd.n329 185
R16029 vdd.n3379 vdd.n329 185
R16030 vdd.n3308 vdd.n3307 185
R16031 vdd.n3307 vdd.n328 185
R16032 vdd.n3306 vdd.n610 185
R16033 vdd.n3306 vdd.n3305 185
R16034 vdd.n3294 vdd.n612 185
R16035 vdd.n613 vdd.n612 185
R16036 vdd.n3296 vdd.n3295 185
R16037 vdd.n3297 vdd.n3296 185
R16038 vdd.n620 vdd.n619 185
R16039 vdd.n624 vdd.n619 185
R16040 vdd.n3288 vdd.n3287 185
R16041 vdd.n3287 vdd.n3286 185
R16042 vdd.n623 vdd.n622 185
R16043 vdd.n3277 vdd.n623 185
R16044 vdd.n3276 vdd.n3275 185
R16045 vdd.n3278 vdd.n3276 185
R16046 vdd.n631 vdd.n630 185
R16047 vdd.n636 vdd.n630 185
R16048 vdd.n3271 vdd.n3270 185
R16049 vdd.n3270 vdd.n3269 185
R16050 vdd.n634 vdd.n633 185
R16051 vdd.n635 vdd.n634 185
R16052 vdd.n3260 vdd.n3259 185
R16053 vdd.n3261 vdd.n3260 185
R16054 vdd.n644 vdd.n643 185
R16055 vdd.n643 vdd.n642 185
R16056 vdd.n3255 vdd.n3254 185
R16057 vdd.n3254 vdd.n3253 185
R16058 vdd.n647 vdd.n646 185
R16059 vdd.n648 vdd.n647 185
R16060 vdd.n3244 vdd.n3243 185
R16061 vdd.n3245 vdd.n3244 185
R16062 vdd.n655 vdd.n654 185
R16063 vdd.n659 vdd.n654 185
R16064 vdd.n3239 vdd.n3238 185
R16065 vdd.n3238 vdd.n3237 185
R16066 vdd.n2853 vdd.n2852 185
R16067 vdd.n2851 vdd.n2617 185
R16068 vdd.n2850 vdd.n2616 185
R16069 vdd.n2855 vdd.n2616 185
R16070 vdd.n2849 vdd.n2848 185
R16071 vdd.n2847 vdd.n2846 185
R16072 vdd.n2845 vdd.n2844 185
R16073 vdd.n2843 vdd.n2842 185
R16074 vdd.n2841 vdd.n2840 185
R16075 vdd.n2839 vdd.n2838 185
R16076 vdd.n2837 vdd.n2836 185
R16077 vdd.n2835 vdd.n2834 185
R16078 vdd.n2833 vdd.n2832 185
R16079 vdd.n2831 vdd.n2830 185
R16080 vdd.n2829 vdd.n2828 185
R16081 vdd.n2827 vdd.n2826 185
R16082 vdd.n2825 vdd.n2824 185
R16083 vdd.n2823 vdd.n2822 185
R16084 vdd.n2821 vdd.n2820 185
R16085 vdd.n2819 vdd.n2818 185
R16086 vdd.n2817 vdd.n2816 185
R16087 vdd.n2815 vdd.n2814 185
R16088 vdd.n2813 vdd.n2812 185
R16089 vdd.n2811 vdd.n2810 185
R16090 vdd.n2809 vdd.n2808 185
R16091 vdd.n2807 vdd.n2806 185
R16092 vdd.n2805 vdd.n2804 185
R16093 vdd.n2803 vdd.n2802 185
R16094 vdd.n2801 vdd.n2800 185
R16095 vdd.n2799 vdd.n2798 185
R16096 vdd.n2797 vdd.n2796 185
R16097 vdd.n2795 vdd.n2794 185
R16098 vdd.n2793 vdd.n2792 185
R16099 vdd.n2790 vdd.n2789 185
R16100 vdd.n2788 vdd.n2787 185
R16101 vdd.n2786 vdd.n2785 185
R16102 vdd.n3005 vdd.n3004 185
R16103 vdd.n3006 vdd.n803 185
R16104 vdd.n3008 vdd.n3007 185
R16105 vdd.n3010 vdd.n801 185
R16106 vdd.n3012 vdd.n3011 185
R16107 vdd.n3013 vdd.n800 185
R16108 vdd.n3015 vdd.n3014 185
R16109 vdd.n3017 vdd.n798 185
R16110 vdd.n3019 vdd.n3018 185
R16111 vdd.n3020 vdd.n797 185
R16112 vdd.n3022 vdd.n3021 185
R16113 vdd.n3024 vdd.n795 185
R16114 vdd.n3026 vdd.n3025 185
R16115 vdd.n3027 vdd.n794 185
R16116 vdd.n3029 vdd.n3028 185
R16117 vdd.n3031 vdd.n792 185
R16118 vdd.n3033 vdd.n3032 185
R16119 vdd.n3035 vdd.n791 185
R16120 vdd.n3037 vdd.n3036 185
R16121 vdd.n3039 vdd.n789 185
R16122 vdd.n3041 vdd.n3040 185
R16123 vdd.n3042 vdd.n788 185
R16124 vdd.n3044 vdd.n3043 185
R16125 vdd.n3046 vdd.n786 185
R16126 vdd.n3048 vdd.n3047 185
R16127 vdd.n3049 vdd.n785 185
R16128 vdd.n3051 vdd.n3050 185
R16129 vdd.n3053 vdd.n783 185
R16130 vdd.n3055 vdd.n3054 185
R16131 vdd.n3056 vdd.n782 185
R16132 vdd.n3058 vdd.n3057 185
R16133 vdd.n3060 vdd.n781 185
R16134 vdd.n3061 vdd.n780 185
R16135 vdd.n3064 vdd.n3063 185
R16136 vdd.n3065 vdd.n778 185
R16137 vdd.n778 vdd.n756 185
R16138 vdd.n3002 vdd.n775 185
R16139 vdd.n3068 vdd.n775 185
R16140 vdd.n3001 vdd.n3000 185
R16141 vdd.n3000 vdd.n774 185
R16142 vdd.n2999 vdd.n807 185
R16143 vdd.n2999 vdd.n2998 185
R16144 vdd.n2733 vdd.n808 185
R16145 vdd.n817 vdd.n808 185
R16146 vdd.n2734 vdd.n815 185
R16147 vdd.n2992 vdd.n815 185
R16148 vdd.n2736 vdd.n2735 185
R16149 vdd.n2735 vdd.n814 185
R16150 vdd.n2737 vdd.n823 185
R16151 vdd.n2941 vdd.n823 185
R16152 vdd.n2739 vdd.n2738 185
R16153 vdd.n2738 vdd.n822 185
R16154 vdd.n2740 vdd.n829 185
R16155 vdd.n2935 vdd.n829 185
R16156 vdd.n2742 vdd.n2741 185
R16157 vdd.n2741 vdd.n828 185
R16158 vdd.n2743 vdd.n834 185
R16159 vdd.n2929 vdd.n834 185
R16160 vdd.n2745 vdd.n2744 185
R16161 vdd.n2744 vdd.n841 185
R16162 vdd.n2746 vdd.n839 185
R16163 vdd.n2923 vdd.n839 185
R16164 vdd.n2748 vdd.n2747 185
R16165 vdd.n2747 vdd.n849 185
R16166 vdd.n2749 vdd.n847 185
R16167 vdd.n2916 vdd.n847 185
R16168 vdd.n2751 vdd.n2750 185
R16169 vdd.n2750 vdd.n846 185
R16170 vdd.n2752 vdd.n854 185
R16171 vdd.n2910 vdd.n854 185
R16172 vdd.n2754 vdd.n2753 185
R16173 vdd.n2753 vdd.n853 185
R16174 vdd.n2755 vdd.n859 185
R16175 vdd.n2904 vdd.n859 185
R16176 vdd.n2757 vdd.n2756 185
R16177 vdd.n2756 vdd.n866 185
R16178 vdd.n2758 vdd.n864 185
R16179 vdd.n2898 vdd.n864 185
R16180 vdd.n2760 vdd.n2759 185
R16181 vdd.n2759 vdd.n872 185
R16182 vdd.n2761 vdd.n870 185
R16183 vdd.n2892 vdd.n870 185
R16184 vdd.n2763 vdd.n2762 185
R16185 vdd.n2764 vdd.n2763 185
R16186 vdd.n2732 vdd.n877 185
R16187 vdd.n2886 vdd.n877 185
R16188 vdd.n2731 vdd.n2730 185
R16189 vdd.n2730 vdd.n876 185
R16190 vdd.n2729 vdd.n883 185
R16191 vdd.n2880 vdd.n883 185
R16192 vdd.n2728 vdd.n2727 185
R16193 vdd.n2727 vdd.n882 185
R16194 vdd.n2726 vdd.n889 185
R16195 vdd.n2874 vdd.n889 185
R16196 vdd.n2725 vdd.n2724 185
R16197 vdd.n2724 vdd.n888 185
R16198 vdd.n2620 vdd.n894 185
R16199 vdd.n2868 vdd.n894 185
R16200 vdd.n2781 vdd.n2780 185
R16201 vdd.n2780 vdd.n2779 185
R16202 vdd.n2782 vdd.n900 185
R16203 vdd.n2862 vdd.n900 185
R16204 vdd.n2784 vdd.n2783 185
R16205 vdd.n2784 vdd.n899 185
R16206 vdd.n898 vdd.n897 185
R16207 vdd.n899 vdd.n898 185
R16208 vdd.n2864 vdd.n2863 185
R16209 vdd.n2863 vdd.n2862 185
R16210 vdd.n2865 vdd.n896 185
R16211 vdd.n2779 vdd.n896 185
R16212 vdd.n2867 vdd.n2866 185
R16213 vdd.n2868 vdd.n2867 185
R16214 vdd.n887 vdd.n886 185
R16215 vdd.n888 vdd.n887 185
R16216 vdd.n2876 vdd.n2875 185
R16217 vdd.n2875 vdd.n2874 185
R16218 vdd.n2877 vdd.n885 185
R16219 vdd.n885 vdd.n882 185
R16220 vdd.n2879 vdd.n2878 185
R16221 vdd.n2880 vdd.n2879 185
R16222 vdd.n875 vdd.n874 185
R16223 vdd.n876 vdd.n875 185
R16224 vdd.n2888 vdd.n2887 185
R16225 vdd.n2887 vdd.n2886 185
R16226 vdd.n2889 vdd.n873 185
R16227 vdd.n2764 vdd.n873 185
R16228 vdd.n2891 vdd.n2890 185
R16229 vdd.n2892 vdd.n2891 185
R16230 vdd.n863 vdd.n862 185
R16231 vdd.n872 vdd.n863 185
R16232 vdd.n2900 vdd.n2899 185
R16233 vdd.n2899 vdd.n2898 185
R16234 vdd.n2901 vdd.n861 185
R16235 vdd.n866 vdd.n861 185
R16236 vdd.n2903 vdd.n2902 185
R16237 vdd.n2904 vdd.n2903 185
R16238 vdd.n852 vdd.n851 185
R16239 vdd.n853 vdd.n852 185
R16240 vdd.n2912 vdd.n2911 185
R16241 vdd.n2911 vdd.n2910 185
R16242 vdd.n2913 vdd.n850 185
R16243 vdd.n850 vdd.n846 185
R16244 vdd.n2915 vdd.n2914 185
R16245 vdd.n2916 vdd.n2915 185
R16246 vdd.n838 vdd.n837 185
R16247 vdd.n849 vdd.n838 185
R16248 vdd.n2925 vdd.n2924 185
R16249 vdd.n2924 vdd.n2923 185
R16250 vdd.n2926 vdd.n836 185
R16251 vdd.n841 vdd.n836 185
R16252 vdd.n2928 vdd.n2927 185
R16253 vdd.n2929 vdd.n2928 185
R16254 vdd.n827 vdd.n826 185
R16255 vdd.n828 vdd.n827 185
R16256 vdd.n2937 vdd.n2936 185
R16257 vdd.n2936 vdd.n2935 185
R16258 vdd.n2938 vdd.n825 185
R16259 vdd.n825 vdd.n822 185
R16260 vdd.n2940 vdd.n2939 185
R16261 vdd.n2941 vdd.n2940 185
R16262 vdd.n813 vdd.n812 185
R16263 vdd.n814 vdd.n813 185
R16264 vdd.n2994 vdd.n2993 185
R16265 vdd.n2993 vdd.n2992 185
R16266 vdd.n2995 vdd.n811 185
R16267 vdd.n817 vdd.n811 185
R16268 vdd.n2997 vdd.n2996 185
R16269 vdd.n2998 vdd.n2997 185
R16270 vdd.n779 vdd.n777 185
R16271 vdd.n777 vdd.n774 185
R16272 vdd.n3067 vdd.n3066 185
R16273 vdd.n3068 vdd.n3067 185
R16274 vdd.n2509 vdd.n2508 185
R16275 vdd.n2510 vdd.n2509 185
R16276 vdd.n951 vdd.n949 185
R16277 vdd.n949 vdd.n947 185
R16278 vdd.n2424 vdd.n958 185
R16279 vdd.n2435 vdd.n958 185
R16280 vdd.n2425 vdd.n967 185
R16281 vdd.n1309 vdd.n967 185
R16282 vdd.n2427 vdd.n2426 185
R16283 vdd.n2428 vdd.n2427 185
R16284 vdd.n2423 vdd.n966 185
R16285 vdd.n966 vdd.n963 185
R16286 vdd.n2422 vdd.n2421 185
R16287 vdd.n2421 vdd.n2420 185
R16288 vdd.n969 vdd.n968 185
R16289 vdd.n970 vdd.n969 185
R16290 vdd.n2413 vdd.n2412 185
R16291 vdd.n2414 vdd.n2413 185
R16292 vdd.n2411 vdd.n979 185
R16293 vdd.n979 vdd.n976 185
R16294 vdd.n2410 vdd.n2409 185
R16295 vdd.n2409 vdd.n2408 185
R16296 vdd.n981 vdd.n980 185
R16297 vdd.n989 vdd.n981 185
R16298 vdd.n2401 vdd.n2400 185
R16299 vdd.n2402 vdd.n2401 185
R16300 vdd.n2399 vdd.n990 185
R16301 vdd.n995 vdd.n990 185
R16302 vdd.n2398 vdd.n2397 185
R16303 vdd.n2397 vdd.n2396 185
R16304 vdd.n992 vdd.n991 185
R16305 vdd.n1330 vdd.n992 185
R16306 vdd.n2389 vdd.n2388 185
R16307 vdd.n2390 vdd.n2389 185
R16308 vdd.n2387 vdd.n1002 185
R16309 vdd.n1002 vdd.n999 185
R16310 vdd.n2386 vdd.n2385 185
R16311 vdd.n2385 vdd.n2384 185
R16312 vdd.n1004 vdd.n1003 185
R16313 vdd.n1005 vdd.n1004 185
R16314 vdd.n2377 vdd.n2376 185
R16315 vdd.n2378 vdd.n2377 185
R16316 vdd.n2374 vdd.n1013 185
R16317 vdd.n1019 vdd.n1013 185
R16318 vdd.n2373 vdd.n2372 185
R16319 vdd.n2372 vdd.n2371 185
R16320 vdd.n1016 vdd.n1015 185
R16321 vdd.n1026 vdd.n1016 185
R16322 vdd.n2364 vdd.n2363 185
R16323 vdd.n2365 vdd.n2364 185
R16324 vdd.n2362 vdd.n1027 185
R16325 vdd.n1027 vdd.n1023 185
R16326 vdd.n2361 vdd.n2360 185
R16327 vdd.n2360 vdd.n2359 185
R16328 vdd.n1029 vdd.n1028 185
R16329 vdd.n1030 vdd.n1029 185
R16330 vdd.n2352 vdd.n2351 185
R16331 vdd.n2353 vdd.n2352 185
R16332 vdd.n2350 vdd.n1039 185
R16333 vdd.n1039 vdd.n1036 185
R16334 vdd.n2349 vdd.n2348 185
R16335 vdd.n2348 vdd.n2347 185
R16336 vdd.n1041 vdd.n1040 185
R16337 vdd.n1050 vdd.n1041 185
R16338 vdd.n2340 vdd.n2339 185
R16339 vdd.n2341 vdd.n2340 185
R16340 vdd.n2338 vdd.n1051 185
R16341 vdd.n1051 vdd.n1047 185
R16342 vdd.n2440 vdd.n922 185
R16343 vdd.n2582 vdd.n922 185
R16344 vdd.n2442 vdd.n2441 185
R16345 vdd.n2444 vdd.n2443 185
R16346 vdd.n2446 vdd.n2445 185
R16347 vdd.n2448 vdd.n2447 185
R16348 vdd.n2450 vdd.n2449 185
R16349 vdd.n2452 vdd.n2451 185
R16350 vdd.n2454 vdd.n2453 185
R16351 vdd.n2456 vdd.n2455 185
R16352 vdd.n2458 vdd.n2457 185
R16353 vdd.n2460 vdd.n2459 185
R16354 vdd.n2462 vdd.n2461 185
R16355 vdd.n2464 vdd.n2463 185
R16356 vdd.n2466 vdd.n2465 185
R16357 vdd.n2468 vdd.n2467 185
R16358 vdd.n2470 vdd.n2469 185
R16359 vdd.n2472 vdd.n2471 185
R16360 vdd.n2474 vdd.n2473 185
R16361 vdd.n2476 vdd.n2475 185
R16362 vdd.n2478 vdd.n2477 185
R16363 vdd.n2480 vdd.n2479 185
R16364 vdd.n2482 vdd.n2481 185
R16365 vdd.n2484 vdd.n2483 185
R16366 vdd.n2486 vdd.n2485 185
R16367 vdd.n2488 vdd.n2487 185
R16368 vdd.n2490 vdd.n2489 185
R16369 vdd.n2492 vdd.n2491 185
R16370 vdd.n2494 vdd.n2493 185
R16371 vdd.n2496 vdd.n2495 185
R16372 vdd.n2498 vdd.n2497 185
R16373 vdd.n2500 vdd.n2499 185
R16374 vdd.n2502 vdd.n2501 185
R16375 vdd.n2504 vdd.n2503 185
R16376 vdd.n2506 vdd.n2505 185
R16377 vdd.n2507 vdd.n950 185
R16378 vdd.n2439 vdd.n948 185
R16379 vdd.n2510 vdd.n948 185
R16380 vdd.n2438 vdd.n2437 185
R16381 vdd.n2437 vdd.n947 185
R16382 vdd.n2436 vdd.n955 185
R16383 vdd.n2436 vdd.n2435 185
R16384 vdd.n1227 vdd.n956 185
R16385 vdd.n1309 vdd.n956 185
R16386 vdd.n1228 vdd.n965 185
R16387 vdd.n2428 vdd.n965 185
R16388 vdd.n1230 vdd.n1229 185
R16389 vdd.n1229 vdd.n963 185
R16390 vdd.n1231 vdd.n972 185
R16391 vdd.n2420 vdd.n972 185
R16392 vdd.n1233 vdd.n1232 185
R16393 vdd.n1232 vdd.n970 185
R16394 vdd.n1234 vdd.n978 185
R16395 vdd.n2414 vdd.n978 185
R16396 vdd.n1236 vdd.n1235 185
R16397 vdd.n1235 vdd.n976 185
R16398 vdd.n1237 vdd.n983 185
R16399 vdd.n2408 vdd.n983 185
R16400 vdd.n1239 vdd.n1238 185
R16401 vdd.n1238 vdd.n989 185
R16402 vdd.n1240 vdd.n988 185
R16403 vdd.n2402 vdd.n988 185
R16404 vdd.n1242 vdd.n1241 185
R16405 vdd.n1241 vdd.n995 185
R16406 vdd.n1243 vdd.n994 185
R16407 vdd.n2396 vdd.n994 185
R16408 vdd.n1332 vdd.n1331 185
R16409 vdd.n1331 vdd.n1330 185
R16410 vdd.n1333 vdd.n1001 185
R16411 vdd.n2390 vdd.n1001 185
R16412 vdd.n1335 vdd.n1334 185
R16413 vdd.n1334 vdd.n999 185
R16414 vdd.n1336 vdd.n1007 185
R16415 vdd.n2384 vdd.n1007 185
R16416 vdd.n1338 vdd.n1337 185
R16417 vdd.n1337 vdd.n1005 185
R16418 vdd.n1339 vdd.n1012 185
R16419 vdd.n2378 vdd.n1012 185
R16420 vdd.n1341 vdd.n1340 185
R16421 vdd.n1340 vdd.n1019 185
R16422 vdd.n1342 vdd.n1018 185
R16423 vdd.n2371 vdd.n1018 185
R16424 vdd.n1344 vdd.n1343 185
R16425 vdd.n1343 vdd.n1026 185
R16426 vdd.n1345 vdd.n1025 185
R16427 vdd.n2365 vdd.n1025 185
R16428 vdd.n1347 vdd.n1346 185
R16429 vdd.n1346 vdd.n1023 185
R16430 vdd.n1348 vdd.n1032 185
R16431 vdd.n2359 vdd.n1032 185
R16432 vdd.n1350 vdd.n1349 185
R16433 vdd.n1349 vdd.n1030 185
R16434 vdd.n1351 vdd.n1038 185
R16435 vdd.n2353 vdd.n1038 185
R16436 vdd.n1353 vdd.n1352 185
R16437 vdd.n1352 vdd.n1036 185
R16438 vdd.n1354 vdd.n1043 185
R16439 vdd.n2347 vdd.n1043 185
R16440 vdd.n1356 vdd.n1355 185
R16441 vdd.n1355 vdd.n1050 185
R16442 vdd.n1357 vdd.n1049 185
R16443 vdd.n2341 vdd.n1049 185
R16444 vdd.n1359 vdd.n1358 185
R16445 vdd.n1358 vdd.n1047 185
R16446 vdd.n2337 vdd.n2336 185
R16447 vdd.n1053 vdd.n1052 185
R16448 vdd.n1194 vdd.n1193 185
R16449 vdd.n1196 vdd.n1195 185
R16450 vdd.n1198 vdd.n1197 185
R16451 vdd.n1200 vdd.n1199 185
R16452 vdd.n1202 vdd.n1201 185
R16453 vdd.n1204 vdd.n1203 185
R16454 vdd.n1206 vdd.n1205 185
R16455 vdd.n1208 vdd.n1207 185
R16456 vdd.n1210 vdd.n1209 185
R16457 vdd.n1212 vdd.n1211 185
R16458 vdd.n1214 vdd.n1213 185
R16459 vdd.n1216 vdd.n1215 185
R16460 vdd.n1218 vdd.n1217 185
R16461 vdd.n1220 vdd.n1219 185
R16462 vdd.n1222 vdd.n1221 185
R16463 vdd.n1393 vdd.n1223 185
R16464 vdd.n1392 vdd.n1391 185
R16465 vdd.n1390 vdd.n1389 185
R16466 vdd.n1388 vdd.n1387 185
R16467 vdd.n1386 vdd.n1385 185
R16468 vdd.n1384 vdd.n1383 185
R16469 vdd.n1382 vdd.n1381 185
R16470 vdd.n1380 vdd.n1379 185
R16471 vdd.n1378 vdd.n1377 185
R16472 vdd.n1376 vdd.n1375 185
R16473 vdd.n1374 vdd.n1373 185
R16474 vdd.n1372 vdd.n1371 185
R16475 vdd.n1370 vdd.n1369 185
R16476 vdd.n1368 vdd.n1367 185
R16477 vdd.n1366 vdd.n1365 185
R16478 vdd.n1364 vdd.n1363 185
R16479 vdd.n1362 vdd.n1361 185
R16480 vdd.n1360 vdd.n1087 185
R16481 vdd.n2334 vdd.n1087 185
R16482 vdd.n2334 vdd.n1054 179.345
R16483 vdd.n756 vdd.n658 179.345
R16484 vdd.n315 vdd.n314 171.744
R16485 vdd.n314 vdd.n313 171.744
R16486 vdd.n313 vdd.n282 171.744
R16487 vdd.n306 vdd.n282 171.744
R16488 vdd.n306 vdd.n305 171.744
R16489 vdd.n305 vdd.n287 171.744
R16490 vdd.n298 vdd.n287 171.744
R16491 vdd.n298 vdd.n297 171.744
R16492 vdd.n297 vdd.n291 171.744
R16493 vdd.n260 vdd.n259 171.744
R16494 vdd.n259 vdd.n258 171.744
R16495 vdd.n258 vdd.n227 171.744
R16496 vdd.n251 vdd.n227 171.744
R16497 vdd.n251 vdd.n250 171.744
R16498 vdd.n250 vdd.n232 171.744
R16499 vdd.n243 vdd.n232 171.744
R16500 vdd.n243 vdd.n242 171.744
R16501 vdd.n242 vdd.n236 171.744
R16502 vdd.n217 vdd.n216 171.744
R16503 vdd.n216 vdd.n215 171.744
R16504 vdd.n215 vdd.n184 171.744
R16505 vdd.n208 vdd.n184 171.744
R16506 vdd.n208 vdd.n207 171.744
R16507 vdd.n207 vdd.n189 171.744
R16508 vdd.n200 vdd.n189 171.744
R16509 vdd.n200 vdd.n199 171.744
R16510 vdd.n199 vdd.n193 171.744
R16511 vdd.n162 vdd.n161 171.744
R16512 vdd.n161 vdd.n160 171.744
R16513 vdd.n160 vdd.n129 171.744
R16514 vdd.n153 vdd.n129 171.744
R16515 vdd.n153 vdd.n152 171.744
R16516 vdd.n152 vdd.n134 171.744
R16517 vdd.n145 vdd.n134 171.744
R16518 vdd.n145 vdd.n144 171.744
R16519 vdd.n144 vdd.n138 171.744
R16520 vdd.n120 vdd.n119 171.744
R16521 vdd.n119 vdd.n118 171.744
R16522 vdd.n118 vdd.n87 171.744
R16523 vdd.n111 vdd.n87 171.744
R16524 vdd.n111 vdd.n110 171.744
R16525 vdd.n110 vdd.n92 171.744
R16526 vdd.n103 vdd.n92 171.744
R16527 vdd.n103 vdd.n102 171.744
R16528 vdd.n102 vdd.n96 171.744
R16529 vdd.n65 vdd.n64 171.744
R16530 vdd.n64 vdd.n63 171.744
R16531 vdd.n63 vdd.n32 171.744
R16532 vdd.n56 vdd.n32 171.744
R16533 vdd.n56 vdd.n55 171.744
R16534 vdd.n55 vdd.n37 171.744
R16535 vdd.n48 vdd.n37 171.744
R16536 vdd.n48 vdd.n47 171.744
R16537 vdd.n47 vdd.n41 171.744
R16538 vdd.n2046 vdd.n2045 171.744
R16539 vdd.n2045 vdd.n2044 171.744
R16540 vdd.n2044 vdd.n2013 171.744
R16541 vdd.n2037 vdd.n2013 171.744
R16542 vdd.n2037 vdd.n2036 171.744
R16543 vdd.n2036 vdd.n2018 171.744
R16544 vdd.n2029 vdd.n2018 171.744
R16545 vdd.n2029 vdd.n2028 171.744
R16546 vdd.n2028 vdd.n2022 171.744
R16547 vdd.n2101 vdd.n2100 171.744
R16548 vdd.n2100 vdd.n2099 171.744
R16549 vdd.n2099 vdd.n2068 171.744
R16550 vdd.n2092 vdd.n2068 171.744
R16551 vdd.n2092 vdd.n2091 171.744
R16552 vdd.n2091 vdd.n2073 171.744
R16553 vdd.n2084 vdd.n2073 171.744
R16554 vdd.n2084 vdd.n2083 171.744
R16555 vdd.n2083 vdd.n2077 171.744
R16556 vdd.n1948 vdd.n1947 171.744
R16557 vdd.n1947 vdd.n1946 171.744
R16558 vdd.n1946 vdd.n1915 171.744
R16559 vdd.n1939 vdd.n1915 171.744
R16560 vdd.n1939 vdd.n1938 171.744
R16561 vdd.n1938 vdd.n1920 171.744
R16562 vdd.n1931 vdd.n1920 171.744
R16563 vdd.n1931 vdd.n1930 171.744
R16564 vdd.n1930 vdd.n1924 171.744
R16565 vdd.n2003 vdd.n2002 171.744
R16566 vdd.n2002 vdd.n2001 171.744
R16567 vdd.n2001 vdd.n1970 171.744
R16568 vdd.n1994 vdd.n1970 171.744
R16569 vdd.n1994 vdd.n1993 171.744
R16570 vdd.n1993 vdd.n1975 171.744
R16571 vdd.n1986 vdd.n1975 171.744
R16572 vdd.n1986 vdd.n1985 171.744
R16573 vdd.n1985 vdd.n1979 171.744
R16574 vdd.n1851 vdd.n1850 171.744
R16575 vdd.n1850 vdd.n1849 171.744
R16576 vdd.n1849 vdd.n1818 171.744
R16577 vdd.n1842 vdd.n1818 171.744
R16578 vdd.n1842 vdd.n1841 171.744
R16579 vdd.n1841 vdd.n1823 171.744
R16580 vdd.n1834 vdd.n1823 171.744
R16581 vdd.n1834 vdd.n1833 171.744
R16582 vdd.n1833 vdd.n1827 171.744
R16583 vdd.n1906 vdd.n1905 171.744
R16584 vdd.n1905 vdd.n1904 171.744
R16585 vdd.n1904 vdd.n1873 171.744
R16586 vdd.n1897 vdd.n1873 171.744
R16587 vdd.n1897 vdd.n1896 171.744
R16588 vdd.n1896 vdd.n1878 171.744
R16589 vdd.n1889 vdd.n1878 171.744
R16590 vdd.n1889 vdd.n1888 171.744
R16591 vdd.n1888 vdd.n1882 171.744
R16592 vdd.n449 vdd.n448 146.341
R16593 vdd.n455 vdd.n454 146.341
R16594 vdd.n459 vdd.n458 146.341
R16595 vdd.n465 vdd.n464 146.341
R16596 vdd.n469 vdd.n468 146.341
R16597 vdd.n475 vdd.n474 146.341
R16598 vdd.n479 vdd.n478 146.341
R16599 vdd.n485 vdd.n484 146.341
R16600 vdd.n489 vdd.n488 146.341
R16601 vdd.n495 vdd.n494 146.341
R16602 vdd.n499 vdd.n498 146.341
R16603 vdd.n505 vdd.n504 146.341
R16604 vdd.n509 vdd.n508 146.341
R16605 vdd.n515 vdd.n514 146.341
R16606 vdd.n519 vdd.n518 146.341
R16607 vdd.n525 vdd.n524 146.341
R16608 vdd.n529 vdd.n528 146.341
R16609 vdd.n535 vdd.n534 146.341
R16610 vdd.n539 vdd.n538 146.341
R16611 vdd.n545 vdd.n544 146.341
R16612 vdd.n549 vdd.n548 146.341
R16613 vdd.n555 vdd.n554 146.341
R16614 vdd.n559 vdd.n558 146.341
R16615 vdd.n565 vdd.n564 146.341
R16616 vdd.n569 vdd.n568 146.341
R16617 vdd.n575 vdd.n574 146.341
R16618 vdd.n579 vdd.n578 146.341
R16619 vdd.n585 vdd.n584 146.341
R16620 vdd.n589 vdd.n588 146.341
R16621 vdd.n595 vdd.n594 146.341
R16622 vdd.n597 vdd.n404 146.341
R16623 vdd.n3238 vdd.n654 146.341
R16624 vdd.n3244 vdd.n654 146.341
R16625 vdd.n3244 vdd.n647 146.341
R16626 vdd.n3254 vdd.n647 146.341
R16627 vdd.n3254 vdd.n643 146.341
R16628 vdd.n3260 vdd.n643 146.341
R16629 vdd.n3260 vdd.n634 146.341
R16630 vdd.n3270 vdd.n634 146.341
R16631 vdd.n3270 vdd.n630 146.341
R16632 vdd.n3276 vdd.n630 146.341
R16633 vdd.n3276 vdd.n623 146.341
R16634 vdd.n3287 vdd.n623 146.341
R16635 vdd.n3287 vdd.n619 146.341
R16636 vdd.n3296 vdd.n619 146.341
R16637 vdd.n3296 vdd.n612 146.341
R16638 vdd.n3306 vdd.n612 146.341
R16639 vdd.n3307 vdd.n3306 146.341
R16640 vdd.n3307 vdd.n329 146.341
R16641 vdd.n330 vdd.n329 146.341
R16642 vdd.n331 vdd.n330 146.341
R16643 vdd.n3314 vdd.n331 146.341
R16644 vdd.n3314 vdd.n339 146.341
R16645 vdd.n340 vdd.n339 146.341
R16646 vdd.n341 vdd.n340 146.341
R16647 vdd.n3321 vdd.n341 146.341
R16648 vdd.n3321 vdd.n350 146.341
R16649 vdd.n351 vdd.n350 146.341
R16650 vdd.n352 vdd.n351 146.341
R16651 vdd.n3329 vdd.n352 146.341
R16652 vdd.n3329 vdd.n360 146.341
R16653 vdd.n361 vdd.n360 146.341
R16654 vdd.n362 vdd.n361 146.341
R16655 vdd.n3336 vdd.n362 146.341
R16656 vdd.n3336 vdd.n371 146.341
R16657 vdd.n372 vdd.n371 146.341
R16658 vdd.n3230 vdd.n3228 146.341
R16659 vdd.n3228 vdd.n3227 146.341
R16660 vdd.n3224 vdd.n3223 146.341
R16661 vdd.n3220 vdd.n3219 146.341
R16662 vdd.n3217 vdd.n669 146.341
R16663 vdd.n3213 vdd.n3211 146.341
R16664 vdd.n3209 vdd.n675 146.341
R16665 vdd.n3205 vdd.n3203 146.341
R16666 vdd.n3201 vdd.n681 146.341
R16667 vdd.n3197 vdd.n3195 146.341
R16668 vdd.n3193 vdd.n689 146.341
R16669 vdd.n3189 vdd.n3187 146.341
R16670 vdd.n3185 vdd.n695 146.341
R16671 vdd.n3181 vdd.n3179 146.341
R16672 vdd.n3177 vdd.n701 146.341
R16673 vdd.n3173 vdd.n3171 146.341
R16674 vdd.n3169 vdd.n707 146.341
R16675 vdd.n3165 vdd.n3163 146.341
R16676 vdd.n3161 vdd.n713 146.341
R16677 vdd.n3157 vdd.n3155 146.341
R16678 vdd.n3153 vdd.n719 146.341
R16679 vdd.n3146 vdd.n728 146.341
R16680 vdd.n3144 vdd.n3143 146.341
R16681 vdd.n3140 vdd.n3139 146.341
R16682 vdd.n3137 vdd.n733 146.341
R16683 vdd.n3133 vdd.n3131 146.341
R16684 vdd.n3129 vdd.n739 146.341
R16685 vdd.n3125 vdd.n3123 146.341
R16686 vdd.n3121 vdd.n745 146.341
R16687 vdd.n3117 vdd.n3115 146.341
R16688 vdd.n3112 vdd.n3111 146.341
R16689 vdd.n3108 vdd.n657 146.341
R16690 vdd.n3236 vdd.n653 146.341
R16691 vdd.n3246 vdd.n653 146.341
R16692 vdd.n3246 vdd.n649 146.341
R16693 vdd.n3252 vdd.n649 146.341
R16694 vdd.n3252 vdd.n641 146.341
R16695 vdd.n3262 vdd.n641 146.341
R16696 vdd.n3262 vdd.n637 146.341
R16697 vdd.n3268 vdd.n637 146.341
R16698 vdd.n3268 vdd.n629 146.341
R16699 vdd.n3279 vdd.n629 146.341
R16700 vdd.n3279 vdd.n625 146.341
R16701 vdd.n3285 vdd.n625 146.341
R16702 vdd.n3285 vdd.n618 146.341
R16703 vdd.n3298 vdd.n618 146.341
R16704 vdd.n3298 vdd.n614 146.341
R16705 vdd.n3304 vdd.n614 146.341
R16706 vdd.n3304 vdd.n326 146.341
R16707 vdd.n3380 vdd.n326 146.341
R16708 vdd.n3380 vdd.n327 146.341
R16709 vdd.n3376 vdd.n327 146.341
R16710 vdd.n3376 vdd.n333 146.341
R16711 vdd.n3372 vdd.n333 146.341
R16712 vdd.n3372 vdd.n338 146.341
R16713 vdd.n3368 vdd.n338 146.341
R16714 vdd.n3368 vdd.n342 146.341
R16715 vdd.n3364 vdd.n342 146.341
R16716 vdd.n3364 vdd.n348 146.341
R16717 vdd.n3360 vdd.n348 146.341
R16718 vdd.n3360 vdd.n353 146.341
R16719 vdd.n3356 vdd.n353 146.341
R16720 vdd.n3356 vdd.n359 146.341
R16721 vdd.n3352 vdd.n359 146.341
R16722 vdd.n3352 vdd.n364 146.341
R16723 vdd.n3348 vdd.n364 146.341
R16724 vdd.n3348 vdd.n370 146.341
R16725 vdd.n2295 vdd.n2294 146.341
R16726 vdd.n2292 vdd.n2289 146.341
R16727 vdd.n2287 vdd.n1098 146.341
R16728 vdd.n2283 vdd.n2282 146.341
R16729 vdd.n2280 vdd.n1102 146.341
R16730 vdd.n2276 vdd.n2275 146.341
R16731 vdd.n2273 vdd.n1109 146.341
R16732 vdd.n2269 vdd.n2268 146.341
R16733 vdd.n2266 vdd.n1116 146.341
R16734 vdd.n1127 vdd.n1124 146.341
R16735 vdd.n2258 vdd.n2257 146.341
R16736 vdd.n2255 vdd.n1129 146.341
R16737 vdd.n2251 vdd.n2250 146.341
R16738 vdd.n2248 vdd.n1135 146.341
R16739 vdd.n2244 vdd.n2243 146.341
R16740 vdd.n2241 vdd.n1142 146.341
R16741 vdd.n2237 vdd.n2236 146.341
R16742 vdd.n2234 vdd.n1149 146.341
R16743 vdd.n2230 vdd.n2229 146.341
R16744 vdd.n2227 vdd.n1156 146.341
R16745 vdd.n1167 vdd.n1164 146.341
R16746 vdd.n2219 vdd.n2218 146.341
R16747 vdd.n2216 vdd.n1169 146.341
R16748 vdd.n2212 vdd.n2211 146.341
R16749 vdd.n2209 vdd.n1175 146.341
R16750 vdd.n2205 vdd.n2204 146.341
R16751 vdd.n2202 vdd.n1182 146.341
R16752 vdd.n2198 vdd.n2197 146.341
R16753 vdd.n2195 vdd.n1189 146.341
R16754 vdd.n1400 vdd.n1398 146.341
R16755 vdd.n1403 vdd.n1402 146.341
R16756 vdd.n1743 vdd.n1507 146.341
R16757 vdd.n1743 vdd.n1499 146.341
R16758 vdd.n1753 vdd.n1499 146.341
R16759 vdd.n1753 vdd.n1495 146.341
R16760 vdd.n1759 vdd.n1495 146.341
R16761 vdd.n1759 vdd.n1487 146.341
R16762 vdd.n1770 vdd.n1487 146.341
R16763 vdd.n1770 vdd.n1483 146.341
R16764 vdd.n1776 vdd.n1483 146.341
R16765 vdd.n1776 vdd.n1477 146.341
R16766 vdd.n1787 vdd.n1477 146.341
R16767 vdd.n1787 vdd.n1473 146.341
R16768 vdd.n1793 vdd.n1473 146.341
R16769 vdd.n1793 vdd.n1464 146.341
R16770 vdd.n1803 vdd.n1464 146.341
R16771 vdd.n1803 vdd.n1460 146.341
R16772 vdd.n1809 vdd.n1460 146.341
R16773 vdd.n1809 vdd.n1453 146.341
R16774 vdd.n2115 vdd.n1453 146.341
R16775 vdd.n2115 vdd.n1449 146.341
R16776 vdd.n2121 vdd.n1449 146.341
R16777 vdd.n2121 vdd.n1442 146.341
R16778 vdd.n2131 vdd.n1442 146.341
R16779 vdd.n2131 vdd.n1438 146.341
R16780 vdd.n2137 vdd.n1438 146.341
R16781 vdd.n2137 vdd.n1430 146.341
R16782 vdd.n2148 vdd.n1430 146.341
R16783 vdd.n2148 vdd.n1426 146.341
R16784 vdd.n2154 vdd.n1426 146.341
R16785 vdd.n2154 vdd.n1420 146.341
R16786 vdd.n2165 vdd.n1420 146.341
R16787 vdd.n2165 vdd.n1415 146.341
R16788 vdd.n2173 vdd.n1415 146.341
R16789 vdd.n2173 vdd.n1405 146.341
R16790 vdd.n2183 vdd.n1405 146.341
R16791 vdd.n1545 vdd.n1544 146.341
R16792 vdd.n1549 vdd.n1544 146.341
R16793 vdd.n1551 vdd.n1550 146.341
R16794 vdd.n1555 vdd.n1554 146.341
R16795 vdd.n1557 vdd.n1556 146.341
R16796 vdd.n1561 vdd.n1560 146.341
R16797 vdd.n1563 vdd.n1562 146.341
R16798 vdd.n1567 vdd.n1566 146.341
R16799 vdd.n1569 vdd.n1568 146.341
R16800 vdd.n1701 vdd.n1700 146.341
R16801 vdd.n1573 vdd.n1572 146.341
R16802 vdd.n1577 vdd.n1576 146.341
R16803 vdd.n1579 vdd.n1578 146.341
R16804 vdd.n1583 vdd.n1582 146.341
R16805 vdd.n1585 vdd.n1584 146.341
R16806 vdd.n1589 vdd.n1588 146.341
R16807 vdd.n1591 vdd.n1590 146.341
R16808 vdd.n1595 vdd.n1594 146.341
R16809 vdd.n1597 vdd.n1596 146.341
R16810 vdd.n1601 vdd.n1600 146.341
R16811 vdd.n1665 vdd.n1602 146.341
R16812 vdd.n1606 vdd.n1605 146.341
R16813 vdd.n1608 vdd.n1607 146.341
R16814 vdd.n1612 vdd.n1611 146.341
R16815 vdd.n1614 vdd.n1613 146.341
R16816 vdd.n1618 vdd.n1617 146.341
R16817 vdd.n1620 vdd.n1619 146.341
R16818 vdd.n1624 vdd.n1623 146.341
R16819 vdd.n1626 vdd.n1625 146.341
R16820 vdd.n1630 vdd.n1629 146.341
R16821 vdd.n1632 vdd.n1631 146.341
R16822 vdd.n1737 vdd.n1513 146.341
R16823 vdd.n1745 vdd.n1505 146.341
R16824 vdd.n1745 vdd.n1501 146.341
R16825 vdd.n1751 vdd.n1501 146.341
R16826 vdd.n1751 vdd.n1493 146.341
R16827 vdd.n1762 vdd.n1493 146.341
R16828 vdd.n1762 vdd.n1489 146.341
R16829 vdd.n1768 vdd.n1489 146.341
R16830 vdd.n1768 vdd.n1482 146.341
R16831 vdd.n1779 vdd.n1482 146.341
R16832 vdd.n1779 vdd.n1478 146.341
R16833 vdd.n1785 vdd.n1478 146.341
R16834 vdd.n1785 vdd.n1471 146.341
R16835 vdd.n1795 vdd.n1471 146.341
R16836 vdd.n1795 vdd.n1467 146.341
R16837 vdd.n1801 vdd.n1467 146.341
R16838 vdd.n1801 vdd.n1459 146.341
R16839 vdd.n1812 vdd.n1459 146.341
R16840 vdd.n1812 vdd.n1455 146.341
R16841 vdd.n2113 vdd.n1455 146.341
R16842 vdd.n2113 vdd.n1448 146.341
R16843 vdd.n2123 vdd.n1448 146.341
R16844 vdd.n2123 vdd.n1444 146.341
R16845 vdd.n2129 vdd.n1444 146.341
R16846 vdd.n2129 vdd.n1436 146.341
R16847 vdd.n2140 vdd.n1436 146.341
R16848 vdd.n2140 vdd.n1432 146.341
R16849 vdd.n2146 vdd.n1432 146.341
R16850 vdd.n2146 vdd.n1425 146.341
R16851 vdd.n2157 vdd.n1425 146.341
R16852 vdd.n2157 vdd.n1421 146.341
R16853 vdd.n2163 vdd.n1421 146.341
R16854 vdd.n2163 vdd.n1413 146.341
R16855 vdd.n2175 vdd.n1413 146.341
R16856 vdd.n2175 vdd.n1408 146.341
R16857 vdd.n2181 vdd.n1408 146.341
R16858 vdd.n1224 vdd.t19 127.284
R16859 vdd.n952 vdd.t60 127.284
R16860 vdd.n1244 vdd.t33 127.284
R16861 vdd.n943 vdd.t77 127.284
R16862 vdd.n843 vdd.t36 127.284
R16863 vdd.n843 vdd.t37 127.284
R16864 vdd.n2621 vdd.t75 127.284
R16865 vdd.n804 vdd.t83 127.284
R16866 vdd.n2618 vdd.t65 127.284
R16867 vdd.n768 vdd.t14 127.284
R16868 vdd.n1014 vdd.t68 127.284
R16869 vdd.n1014 vdd.t69 127.284
R16870 vdd.n22 vdd.n20 117.314
R16871 vdd.n17 vdd.n15 117.314
R16872 vdd.n27 vdd.n26 116.927
R16873 vdd.n24 vdd.n23 116.927
R16874 vdd.n22 vdd.n21 116.927
R16875 vdd.n17 vdd.n16 116.927
R16876 vdd.n19 vdd.n18 116.927
R16877 vdd.n27 vdd.n25 116.927
R16878 vdd.n1225 vdd.t18 111.188
R16879 vdd.n953 vdd.t61 111.188
R16880 vdd.n1245 vdd.t32 111.188
R16881 vdd.n944 vdd.t78 111.188
R16882 vdd.n2622 vdd.t74 111.188
R16883 vdd.n805 vdd.t84 111.188
R16884 vdd.n2619 vdd.t64 111.188
R16885 vdd.n769 vdd.t15 111.188
R16886 vdd.n2863 vdd.n898 99.5127
R16887 vdd.n2863 vdd.n896 99.5127
R16888 vdd.n2867 vdd.n896 99.5127
R16889 vdd.n2867 vdd.n887 99.5127
R16890 vdd.n2875 vdd.n887 99.5127
R16891 vdd.n2875 vdd.n885 99.5127
R16892 vdd.n2879 vdd.n885 99.5127
R16893 vdd.n2879 vdd.n875 99.5127
R16894 vdd.n2887 vdd.n875 99.5127
R16895 vdd.n2887 vdd.n873 99.5127
R16896 vdd.n2891 vdd.n873 99.5127
R16897 vdd.n2891 vdd.n863 99.5127
R16898 vdd.n2899 vdd.n863 99.5127
R16899 vdd.n2899 vdd.n861 99.5127
R16900 vdd.n2903 vdd.n861 99.5127
R16901 vdd.n2903 vdd.n852 99.5127
R16902 vdd.n2911 vdd.n852 99.5127
R16903 vdd.n2911 vdd.n850 99.5127
R16904 vdd.n2915 vdd.n850 99.5127
R16905 vdd.n2915 vdd.n838 99.5127
R16906 vdd.n2924 vdd.n838 99.5127
R16907 vdd.n2924 vdd.n836 99.5127
R16908 vdd.n2928 vdd.n836 99.5127
R16909 vdd.n2928 vdd.n827 99.5127
R16910 vdd.n2936 vdd.n827 99.5127
R16911 vdd.n2936 vdd.n825 99.5127
R16912 vdd.n2940 vdd.n825 99.5127
R16913 vdd.n2940 vdd.n813 99.5127
R16914 vdd.n2993 vdd.n813 99.5127
R16915 vdd.n2993 vdd.n811 99.5127
R16916 vdd.n2997 vdd.n811 99.5127
R16917 vdd.n2997 vdd.n777 99.5127
R16918 vdd.n3067 vdd.n777 99.5127
R16919 vdd.n3063 vdd.n778 99.5127
R16920 vdd.n3061 vdd.n3060 99.5127
R16921 vdd.n3058 vdd.n782 99.5127
R16922 vdd.n3054 vdd.n3053 99.5127
R16923 vdd.n3051 vdd.n785 99.5127
R16924 vdd.n3047 vdd.n3046 99.5127
R16925 vdd.n3044 vdd.n788 99.5127
R16926 vdd.n3040 vdd.n3039 99.5127
R16927 vdd.n3037 vdd.n791 99.5127
R16928 vdd.n3032 vdd.n3031 99.5127
R16929 vdd.n3029 vdd.n794 99.5127
R16930 vdd.n3025 vdd.n3024 99.5127
R16931 vdd.n3022 vdd.n797 99.5127
R16932 vdd.n3018 vdd.n3017 99.5127
R16933 vdd.n3015 vdd.n800 99.5127
R16934 vdd.n3011 vdd.n3010 99.5127
R16935 vdd.n3008 vdd.n803 99.5127
R16936 vdd.n2784 vdd.n900 99.5127
R16937 vdd.n2780 vdd.n900 99.5127
R16938 vdd.n2780 vdd.n894 99.5127
R16939 vdd.n2724 vdd.n894 99.5127
R16940 vdd.n2724 vdd.n889 99.5127
R16941 vdd.n2727 vdd.n889 99.5127
R16942 vdd.n2727 vdd.n883 99.5127
R16943 vdd.n2730 vdd.n883 99.5127
R16944 vdd.n2730 vdd.n877 99.5127
R16945 vdd.n2763 vdd.n877 99.5127
R16946 vdd.n2763 vdd.n870 99.5127
R16947 vdd.n2759 vdd.n870 99.5127
R16948 vdd.n2759 vdd.n864 99.5127
R16949 vdd.n2756 vdd.n864 99.5127
R16950 vdd.n2756 vdd.n859 99.5127
R16951 vdd.n2753 vdd.n859 99.5127
R16952 vdd.n2753 vdd.n854 99.5127
R16953 vdd.n2750 vdd.n854 99.5127
R16954 vdd.n2750 vdd.n847 99.5127
R16955 vdd.n2747 vdd.n847 99.5127
R16956 vdd.n2747 vdd.n839 99.5127
R16957 vdd.n2744 vdd.n839 99.5127
R16958 vdd.n2744 vdd.n834 99.5127
R16959 vdd.n2741 vdd.n834 99.5127
R16960 vdd.n2741 vdd.n829 99.5127
R16961 vdd.n2738 vdd.n829 99.5127
R16962 vdd.n2738 vdd.n823 99.5127
R16963 vdd.n2735 vdd.n823 99.5127
R16964 vdd.n2735 vdd.n815 99.5127
R16965 vdd.n815 vdd.n808 99.5127
R16966 vdd.n2999 vdd.n808 99.5127
R16967 vdd.n3000 vdd.n2999 99.5127
R16968 vdd.n3000 vdd.n775 99.5127
R16969 vdd.n2617 vdd.n2616 99.5127
R16970 vdd.n2848 vdd.n2616 99.5127
R16971 vdd.n2846 vdd.n2845 99.5127
R16972 vdd.n2842 vdd.n2841 99.5127
R16973 vdd.n2838 vdd.n2837 99.5127
R16974 vdd.n2834 vdd.n2833 99.5127
R16975 vdd.n2830 vdd.n2829 99.5127
R16976 vdd.n2826 vdd.n2825 99.5127
R16977 vdd.n2822 vdd.n2821 99.5127
R16978 vdd.n2818 vdd.n2817 99.5127
R16979 vdd.n2814 vdd.n2813 99.5127
R16980 vdd.n2810 vdd.n2809 99.5127
R16981 vdd.n2806 vdd.n2805 99.5127
R16982 vdd.n2802 vdd.n2801 99.5127
R16983 vdd.n2798 vdd.n2797 99.5127
R16984 vdd.n2794 vdd.n2793 99.5127
R16985 vdd.n2789 vdd.n2788 99.5127
R16986 vdd.n2581 vdd.n941 99.5127
R16987 vdd.n2577 vdd.n2576 99.5127
R16988 vdd.n2573 vdd.n2572 99.5127
R16989 vdd.n2569 vdd.n2568 99.5127
R16990 vdd.n2565 vdd.n2564 99.5127
R16991 vdd.n2561 vdd.n2560 99.5127
R16992 vdd.n2557 vdd.n2556 99.5127
R16993 vdd.n2553 vdd.n2552 99.5127
R16994 vdd.n2549 vdd.n2548 99.5127
R16995 vdd.n2545 vdd.n2544 99.5127
R16996 vdd.n2541 vdd.n2540 99.5127
R16997 vdd.n2537 vdd.n2536 99.5127
R16998 vdd.n2533 vdd.n2532 99.5127
R16999 vdd.n2529 vdd.n2528 99.5127
R17000 vdd.n2525 vdd.n2524 99.5127
R17001 vdd.n2521 vdd.n2520 99.5127
R17002 vdd.n2516 vdd.n2515 99.5127
R17003 vdd.n1280 vdd.n1048 99.5127
R17004 vdd.n1283 vdd.n1048 99.5127
R17005 vdd.n1283 vdd.n1042 99.5127
R17006 vdd.n1286 vdd.n1042 99.5127
R17007 vdd.n1286 vdd.n1037 99.5127
R17008 vdd.n1289 vdd.n1037 99.5127
R17009 vdd.n1289 vdd.n1031 99.5127
R17010 vdd.n1292 vdd.n1031 99.5127
R17011 vdd.n1292 vdd.n1024 99.5127
R17012 vdd.n1295 vdd.n1024 99.5127
R17013 vdd.n1295 vdd.n1017 99.5127
R17014 vdd.n1298 vdd.n1017 99.5127
R17015 vdd.n1298 vdd.n1011 99.5127
R17016 vdd.n1301 vdd.n1011 99.5127
R17017 vdd.n1301 vdd.n1006 99.5127
R17018 vdd.n1304 vdd.n1006 99.5127
R17019 vdd.n1304 vdd.n1000 99.5127
R17020 vdd.n1329 vdd.n1000 99.5127
R17021 vdd.n1329 vdd.n993 99.5127
R17022 vdd.n1325 vdd.n993 99.5127
R17023 vdd.n1325 vdd.n987 99.5127
R17024 vdd.n1322 vdd.n987 99.5127
R17025 vdd.n1322 vdd.n982 99.5127
R17026 vdd.n1319 vdd.n982 99.5127
R17027 vdd.n1319 vdd.n977 99.5127
R17028 vdd.n1316 vdd.n977 99.5127
R17029 vdd.n1316 vdd.n971 99.5127
R17030 vdd.n1313 vdd.n971 99.5127
R17031 vdd.n1313 vdd.n964 99.5127
R17032 vdd.n1310 vdd.n964 99.5127
R17033 vdd.n1310 vdd.n957 99.5127
R17034 vdd.n957 vdd.n946 99.5127
R17035 vdd.n2511 vdd.n946 99.5127
R17036 vdd.n1089 vdd.n1088 99.5127
R17037 vdd.n2327 vdd.n1088 99.5127
R17038 vdd.n2325 vdd.n2324 99.5127
R17039 vdd.n2321 vdd.n2320 99.5127
R17040 vdd.n2317 vdd.n2316 99.5127
R17041 vdd.n2313 vdd.n2312 99.5127
R17042 vdd.n2309 vdd.n2308 99.5127
R17043 vdd.n2305 vdd.n2304 99.5127
R17044 vdd.n2301 vdd.n2300 99.5127
R17045 vdd.n1247 vdd.n1246 99.5127
R17046 vdd.n1251 vdd.n1250 99.5127
R17047 vdd.n1255 vdd.n1254 99.5127
R17048 vdd.n1259 vdd.n1258 99.5127
R17049 vdd.n1263 vdd.n1262 99.5127
R17050 vdd.n1267 vdd.n1266 99.5127
R17051 vdd.n1271 vdd.n1270 99.5127
R17052 vdd.n1276 vdd.n1275 99.5127
R17053 vdd.n2342 vdd.n1046 99.5127
R17054 vdd.n2342 vdd.n1044 99.5127
R17055 vdd.n2346 vdd.n1044 99.5127
R17056 vdd.n2346 vdd.n1035 99.5127
R17057 vdd.n2354 vdd.n1035 99.5127
R17058 vdd.n2354 vdd.n1033 99.5127
R17059 vdd.n2358 vdd.n1033 99.5127
R17060 vdd.n2358 vdd.n1022 99.5127
R17061 vdd.n2366 vdd.n1022 99.5127
R17062 vdd.n2366 vdd.n1020 99.5127
R17063 vdd.n2370 vdd.n1020 99.5127
R17064 vdd.n2370 vdd.n1010 99.5127
R17065 vdd.n2379 vdd.n1010 99.5127
R17066 vdd.n2379 vdd.n1008 99.5127
R17067 vdd.n2383 vdd.n1008 99.5127
R17068 vdd.n2383 vdd.n998 99.5127
R17069 vdd.n2391 vdd.n998 99.5127
R17070 vdd.n2391 vdd.n996 99.5127
R17071 vdd.n2395 vdd.n996 99.5127
R17072 vdd.n2395 vdd.n986 99.5127
R17073 vdd.n2403 vdd.n986 99.5127
R17074 vdd.n2403 vdd.n984 99.5127
R17075 vdd.n2407 vdd.n984 99.5127
R17076 vdd.n2407 vdd.n975 99.5127
R17077 vdd.n2415 vdd.n975 99.5127
R17078 vdd.n2415 vdd.n973 99.5127
R17079 vdd.n2419 vdd.n973 99.5127
R17080 vdd.n2419 vdd.n962 99.5127
R17081 vdd.n2429 vdd.n962 99.5127
R17082 vdd.n2429 vdd.n959 99.5127
R17083 vdd.n2434 vdd.n959 99.5127
R17084 vdd.n2434 vdd.n960 99.5127
R17085 vdd.n960 vdd.n940 99.5127
R17086 vdd.n2983 vdd.n2982 99.5127
R17087 vdd.n2980 vdd.n2946 99.5127
R17088 vdd.n2976 vdd.n2975 99.5127
R17089 vdd.n2973 vdd.n2949 99.5127
R17090 vdd.n2969 vdd.n2968 99.5127
R17091 vdd.n2966 vdd.n2952 99.5127
R17092 vdd.n2962 vdd.n2961 99.5127
R17093 vdd.n2959 vdd.n2956 99.5127
R17094 vdd.n3100 vdd.n755 99.5127
R17095 vdd.n3098 vdd.n3097 99.5127
R17096 vdd.n3095 vdd.n758 99.5127
R17097 vdd.n3091 vdd.n3090 99.5127
R17098 vdd.n3088 vdd.n761 99.5127
R17099 vdd.n3084 vdd.n3083 99.5127
R17100 vdd.n3081 vdd.n764 99.5127
R17101 vdd.n3077 vdd.n3076 99.5127
R17102 vdd.n3074 vdd.n767 99.5127
R17103 vdd.n2689 vdd.n901 99.5127
R17104 vdd.n2778 vdd.n901 99.5127
R17105 vdd.n2778 vdd.n895 99.5127
R17106 vdd.n2774 vdd.n895 99.5127
R17107 vdd.n2774 vdd.n890 99.5127
R17108 vdd.n2771 vdd.n890 99.5127
R17109 vdd.n2771 vdd.n884 99.5127
R17110 vdd.n2768 vdd.n884 99.5127
R17111 vdd.n2768 vdd.n878 99.5127
R17112 vdd.n2765 vdd.n878 99.5127
R17113 vdd.n2765 vdd.n871 99.5127
R17114 vdd.n2721 vdd.n871 99.5127
R17115 vdd.n2721 vdd.n865 99.5127
R17116 vdd.n2718 vdd.n865 99.5127
R17117 vdd.n2718 vdd.n860 99.5127
R17118 vdd.n2715 vdd.n860 99.5127
R17119 vdd.n2715 vdd.n855 99.5127
R17120 vdd.n2712 vdd.n855 99.5127
R17121 vdd.n2712 vdd.n848 99.5127
R17122 vdd.n2709 vdd.n848 99.5127
R17123 vdd.n2709 vdd.n840 99.5127
R17124 vdd.n2706 vdd.n840 99.5127
R17125 vdd.n2706 vdd.n835 99.5127
R17126 vdd.n2703 vdd.n835 99.5127
R17127 vdd.n2703 vdd.n830 99.5127
R17128 vdd.n2700 vdd.n830 99.5127
R17129 vdd.n2700 vdd.n824 99.5127
R17130 vdd.n2697 vdd.n824 99.5127
R17131 vdd.n2697 vdd.n816 99.5127
R17132 vdd.n2694 vdd.n816 99.5127
R17133 vdd.n2694 vdd.n809 99.5127
R17134 vdd.n809 vdd.n773 99.5127
R17135 vdd.n3069 vdd.n773 99.5127
R17136 vdd.n2624 vdd.n904 99.5127
R17137 vdd.n2628 vdd.n2627 99.5127
R17138 vdd.n2632 vdd.n2631 99.5127
R17139 vdd.n2636 vdd.n2635 99.5127
R17140 vdd.n2640 vdd.n2639 99.5127
R17141 vdd.n2644 vdd.n2643 99.5127
R17142 vdd.n2648 vdd.n2647 99.5127
R17143 vdd.n2652 vdd.n2651 99.5127
R17144 vdd.n2656 vdd.n2655 99.5127
R17145 vdd.n2660 vdd.n2659 99.5127
R17146 vdd.n2664 vdd.n2663 99.5127
R17147 vdd.n2668 vdd.n2667 99.5127
R17148 vdd.n2672 vdd.n2671 99.5127
R17149 vdd.n2676 vdd.n2675 99.5127
R17150 vdd.n2680 vdd.n2679 99.5127
R17151 vdd.n2684 vdd.n2683 99.5127
R17152 vdd.n2686 vdd.n2615 99.5127
R17153 vdd.n2861 vdd.n902 99.5127
R17154 vdd.n2861 vdd.n893 99.5127
R17155 vdd.n2869 vdd.n893 99.5127
R17156 vdd.n2869 vdd.n891 99.5127
R17157 vdd.n2873 vdd.n891 99.5127
R17158 vdd.n2873 vdd.n881 99.5127
R17159 vdd.n2881 vdd.n881 99.5127
R17160 vdd.n2881 vdd.n879 99.5127
R17161 vdd.n2885 vdd.n879 99.5127
R17162 vdd.n2885 vdd.n869 99.5127
R17163 vdd.n2893 vdd.n869 99.5127
R17164 vdd.n2893 vdd.n867 99.5127
R17165 vdd.n2897 vdd.n867 99.5127
R17166 vdd.n2897 vdd.n858 99.5127
R17167 vdd.n2905 vdd.n858 99.5127
R17168 vdd.n2905 vdd.n856 99.5127
R17169 vdd.n2909 vdd.n856 99.5127
R17170 vdd.n2909 vdd.n845 99.5127
R17171 vdd.n2917 vdd.n845 99.5127
R17172 vdd.n2917 vdd.n842 99.5127
R17173 vdd.n2922 vdd.n842 99.5127
R17174 vdd.n2922 vdd.n833 99.5127
R17175 vdd.n2930 vdd.n833 99.5127
R17176 vdd.n2930 vdd.n831 99.5127
R17177 vdd.n2934 vdd.n831 99.5127
R17178 vdd.n2934 vdd.n821 99.5127
R17179 vdd.n2942 vdd.n821 99.5127
R17180 vdd.n2942 vdd.n818 99.5127
R17181 vdd.n2991 vdd.n818 99.5127
R17182 vdd.n2991 vdd.n819 99.5127
R17183 vdd.n819 vdd.n810 99.5127
R17184 vdd.n2986 vdd.n810 99.5127
R17185 vdd.n2986 vdd.n776 99.5127
R17186 vdd.n2505 vdd.n2504 99.5127
R17187 vdd.n2501 vdd.n2500 99.5127
R17188 vdd.n2497 vdd.n2496 99.5127
R17189 vdd.n2493 vdd.n2492 99.5127
R17190 vdd.n2489 vdd.n2488 99.5127
R17191 vdd.n2485 vdd.n2484 99.5127
R17192 vdd.n2481 vdd.n2480 99.5127
R17193 vdd.n2477 vdd.n2476 99.5127
R17194 vdd.n2473 vdd.n2472 99.5127
R17195 vdd.n2469 vdd.n2468 99.5127
R17196 vdd.n2465 vdd.n2464 99.5127
R17197 vdd.n2461 vdd.n2460 99.5127
R17198 vdd.n2457 vdd.n2456 99.5127
R17199 vdd.n2453 vdd.n2452 99.5127
R17200 vdd.n2449 vdd.n2448 99.5127
R17201 vdd.n2445 vdd.n2444 99.5127
R17202 vdd.n2441 vdd.n922 99.5127
R17203 vdd.n1358 vdd.n1049 99.5127
R17204 vdd.n1355 vdd.n1049 99.5127
R17205 vdd.n1355 vdd.n1043 99.5127
R17206 vdd.n1352 vdd.n1043 99.5127
R17207 vdd.n1352 vdd.n1038 99.5127
R17208 vdd.n1349 vdd.n1038 99.5127
R17209 vdd.n1349 vdd.n1032 99.5127
R17210 vdd.n1346 vdd.n1032 99.5127
R17211 vdd.n1346 vdd.n1025 99.5127
R17212 vdd.n1343 vdd.n1025 99.5127
R17213 vdd.n1343 vdd.n1018 99.5127
R17214 vdd.n1340 vdd.n1018 99.5127
R17215 vdd.n1340 vdd.n1012 99.5127
R17216 vdd.n1337 vdd.n1012 99.5127
R17217 vdd.n1337 vdd.n1007 99.5127
R17218 vdd.n1334 vdd.n1007 99.5127
R17219 vdd.n1334 vdd.n1001 99.5127
R17220 vdd.n1331 vdd.n1001 99.5127
R17221 vdd.n1331 vdd.n994 99.5127
R17222 vdd.n1241 vdd.n994 99.5127
R17223 vdd.n1241 vdd.n988 99.5127
R17224 vdd.n1238 vdd.n988 99.5127
R17225 vdd.n1238 vdd.n983 99.5127
R17226 vdd.n1235 vdd.n983 99.5127
R17227 vdd.n1235 vdd.n978 99.5127
R17228 vdd.n1232 vdd.n978 99.5127
R17229 vdd.n1232 vdd.n972 99.5127
R17230 vdd.n1229 vdd.n972 99.5127
R17231 vdd.n1229 vdd.n965 99.5127
R17232 vdd.n965 vdd.n956 99.5127
R17233 vdd.n2436 vdd.n956 99.5127
R17234 vdd.n2437 vdd.n2436 99.5127
R17235 vdd.n2437 vdd.n948 99.5127
R17236 vdd.n1193 vdd.n1053 99.5127
R17237 vdd.n1197 vdd.n1196 99.5127
R17238 vdd.n1201 vdd.n1200 99.5127
R17239 vdd.n1205 vdd.n1204 99.5127
R17240 vdd.n1209 vdd.n1208 99.5127
R17241 vdd.n1213 vdd.n1212 99.5127
R17242 vdd.n1217 vdd.n1216 99.5127
R17243 vdd.n1221 vdd.n1220 99.5127
R17244 vdd.n1391 vdd.n1223 99.5127
R17245 vdd.n1389 vdd.n1388 99.5127
R17246 vdd.n1385 vdd.n1384 99.5127
R17247 vdd.n1381 vdd.n1380 99.5127
R17248 vdd.n1377 vdd.n1376 99.5127
R17249 vdd.n1373 vdd.n1372 99.5127
R17250 vdd.n1369 vdd.n1368 99.5127
R17251 vdd.n1365 vdd.n1364 99.5127
R17252 vdd.n1361 vdd.n1087 99.5127
R17253 vdd.n2340 vdd.n1051 99.5127
R17254 vdd.n2340 vdd.n1041 99.5127
R17255 vdd.n2348 vdd.n1041 99.5127
R17256 vdd.n2348 vdd.n1039 99.5127
R17257 vdd.n2352 vdd.n1039 99.5127
R17258 vdd.n2352 vdd.n1029 99.5127
R17259 vdd.n2360 vdd.n1029 99.5127
R17260 vdd.n2360 vdd.n1027 99.5127
R17261 vdd.n2364 vdd.n1027 99.5127
R17262 vdd.n2364 vdd.n1016 99.5127
R17263 vdd.n2372 vdd.n1016 99.5127
R17264 vdd.n2372 vdd.n1013 99.5127
R17265 vdd.n2377 vdd.n1013 99.5127
R17266 vdd.n2377 vdd.n1004 99.5127
R17267 vdd.n2385 vdd.n1004 99.5127
R17268 vdd.n2385 vdd.n1002 99.5127
R17269 vdd.n2389 vdd.n1002 99.5127
R17270 vdd.n2389 vdd.n992 99.5127
R17271 vdd.n2397 vdd.n992 99.5127
R17272 vdd.n2397 vdd.n990 99.5127
R17273 vdd.n2401 vdd.n990 99.5127
R17274 vdd.n2401 vdd.n981 99.5127
R17275 vdd.n2409 vdd.n981 99.5127
R17276 vdd.n2409 vdd.n979 99.5127
R17277 vdd.n2413 vdd.n979 99.5127
R17278 vdd.n2413 vdd.n969 99.5127
R17279 vdd.n2421 vdd.n969 99.5127
R17280 vdd.n2421 vdd.n966 99.5127
R17281 vdd.n2427 vdd.n966 99.5127
R17282 vdd.n2427 vdd.n967 99.5127
R17283 vdd.n967 vdd.n958 99.5127
R17284 vdd.n958 vdd.n949 99.5127
R17285 vdd.n2509 vdd.n949 99.5127
R17286 vdd.n9 vdd.n7 98.9633
R17287 vdd.n2 vdd.n0 98.9633
R17288 vdd.n9 vdd.n8 98.6055
R17289 vdd.n11 vdd.n10 98.6055
R17290 vdd.n13 vdd.n12 98.6055
R17291 vdd.n6 vdd.n5 98.6055
R17292 vdd.n4 vdd.n3 98.6055
R17293 vdd.n2 vdd.n1 98.6055
R17294 vdd.t220 vdd.n291 85.8723
R17295 vdd.t198 vdd.n236 85.8723
R17296 vdd.t210 vdd.n193 85.8723
R17297 vdd.t185 vdd.n138 85.8723
R17298 vdd.t172 vdd.n96 85.8723
R17299 vdd.t153 vdd.n41 85.8723
R17300 vdd.t231 vdd.n2022 85.8723
R17301 vdd.t141 vdd.n2077 85.8723
R17302 vdd.t221 vdd.n1924 85.8723
R17303 vdd.t120 vdd.n1979 85.8723
R17304 vdd.t155 vdd.n1827 85.8723
R17305 vdd.t173 vdd.n1882 85.8723
R17306 vdd.n2920 vdd.n843 78.546
R17307 vdd.n2375 vdd.n1014 78.546
R17308 vdd.n278 vdd.n277 75.1835
R17309 vdd.n276 vdd.n275 75.1835
R17310 vdd.n274 vdd.n273 75.1835
R17311 vdd.n272 vdd.n271 75.1835
R17312 vdd.n270 vdd.n269 75.1835
R17313 vdd.n268 vdd.n267 75.1835
R17314 vdd.n266 vdd.n265 75.1835
R17315 vdd.n180 vdd.n179 75.1835
R17316 vdd.n178 vdd.n177 75.1835
R17317 vdd.n176 vdd.n175 75.1835
R17318 vdd.n174 vdd.n173 75.1835
R17319 vdd.n172 vdd.n171 75.1835
R17320 vdd.n170 vdd.n169 75.1835
R17321 vdd.n168 vdd.n167 75.1835
R17322 vdd.n83 vdd.n82 75.1835
R17323 vdd.n81 vdd.n80 75.1835
R17324 vdd.n79 vdd.n78 75.1835
R17325 vdd.n77 vdd.n76 75.1835
R17326 vdd.n75 vdd.n74 75.1835
R17327 vdd.n73 vdd.n72 75.1835
R17328 vdd.n71 vdd.n70 75.1835
R17329 vdd.n2052 vdd.n2051 75.1835
R17330 vdd.n2054 vdd.n2053 75.1835
R17331 vdd.n2056 vdd.n2055 75.1835
R17332 vdd.n2058 vdd.n2057 75.1835
R17333 vdd.n2060 vdd.n2059 75.1835
R17334 vdd.n2062 vdd.n2061 75.1835
R17335 vdd.n2064 vdd.n2063 75.1835
R17336 vdd.n1954 vdd.n1953 75.1835
R17337 vdd.n1956 vdd.n1955 75.1835
R17338 vdd.n1958 vdd.n1957 75.1835
R17339 vdd.n1960 vdd.n1959 75.1835
R17340 vdd.n1962 vdd.n1961 75.1835
R17341 vdd.n1964 vdd.n1963 75.1835
R17342 vdd.n1966 vdd.n1965 75.1835
R17343 vdd.n1857 vdd.n1856 75.1835
R17344 vdd.n1859 vdd.n1858 75.1835
R17345 vdd.n1861 vdd.n1860 75.1835
R17346 vdd.n1863 vdd.n1862 75.1835
R17347 vdd.n1865 vdd.n1864 75.1835
R17348 vdd.n1867 vdd.n1866 75.1835
R17349 vdd.n1869 vdd.n1868 75.1835
R17350 vdd.n2856 vdd.n2855 72.8958
R17351 vdd.n2855 vdd.n2599 72.8958
R17352 vdd.n2855 vdd.n2600 72.8958
R17353 vdd.n2855 vdd.n2601 72.8958
R17354 vdd.n2855 vdd.n2602 72.8958
R17355 vdd.n2855 vdd.n2603 72.8958
R17356 vdd.n2855 vdd.n2604 72.8958
R17357 vdd.n2855 vdd.n2605 72.8958
R17358 vdd.n2855 vdd.n2606 72.8958
R17359 vdd.n2855 vdd.n2607 72.8958
R17360 vdd.n2855 vdd.n2608 72.8958
R17361 vdd.n2855 vdd.n2609 72.8958
R17362 vdd.n2855 vdd.n2610 72.8958
R17363 vdd.n2855 vdd.n2611 72.8958
R17364 vdd.n2855 vdd.n2612 72.8958
R17365 vdd.n2855 vdd.n2613 72.8958
R17366 vdd.n2855 vdd.n2614 72.8958
R17367 vdd.n772 vdd.n756 72.8958
R17368 vdd.n3075 vdd.n756 72.8958
R17369 vdd.n766 vdd.n756 72.8958
R17370 vdd.n3082 vdd.n756 72.8958
R17371 vdd.n763 vdd.n756 72.8958
R17372 vdd.n3089 vdd.n756 72.8958
R17373 vdd.n760 vdd.n756 72.8958
R17374 vdd.n3096 vdd.n756 72.8958
R17375 vdd.n3099 vdd.n756 72.8958
R17376 vdd.n2955 vdd.n756 72.8958
R17377 vdd.n2960 vdd.n756 72.8958
R17378 vdd.n2954 vdd.n756 72.8958
R17379 vdd.n2967 vdd.n756 72.8958
R17380 vdd.n2951 vdd.n756 72.8958
R17381 vdd.n2974 vdd.n756 72.8958
R17382 vdd.n2948 vdd.n756 72.8958
R17383 vdd.n2981 vdd.n756 72.8958
R17384 vdd.n2334 vdd.n2333 72.8958
R17385 vdd.n2334 vdd.n1055 72.8958
R17386 vdd.n2334 vdd.n1056 72.8958
R17387 vdd.n2334 vdd.n1057 72.8958
R17388 vdd.n2334 vdd.n1058 72.8958
R17389 vdd.n2334 vdd.n1059 72.8958
R17390 vdd.n2334 vdd.n1060 72.8958
R17391 vdd.n2334 vdd.n1061 72.8958
R17392 vdd.n2334 vdd.n1062 72.8958
R17393 vdd.n2334 vdd.n1063 72.8958
R17394 vdd.n2334 vdd.n1064 72.8958
R17395 vdd.n2334 vdd.n1065 72.8958
R17396 vdd.n2334 vdd.n1066 72.8958
R17397 vdd.n2334 vdd.n1067 72.8958
R17398 vdd.n2334 vdd.n1068 72.8958
R17399 vdd.n2334 vdd.n1069 72.8958
R17400 vdd.n2334 vdd.n1070 72.8958
R17401 vdd.n2582 vdd.n923 72.8958
R17402 vdd.n2582 vdd.n924 72.8958
R17403 vdd.n2582 vdd.n925 72.8958
R17404 vdd.n2582 vdd.n926 72.8958
R17405 vdd.n2582 vdd.n927 72.8958
R17406 vdd.n2582 vdd.n928 72.8958
R17407 vdd.n2582 vdd.n929 72.8958
R17408 vdd.n2582 vdd.n930 72.8958
R17409 vdd.n2582 vdd.n931 72.8958
R17410 vdd.n2582 vdd.n932 72.8958
R17411 vdd.n2582 vdd.n933 72.8958
R17412 vdd.n2582 vdd.n934 72.8958
R17413 vdd.n2582 vdd.n935 72.8958
R17414 vdd.n2582 vdd.n936 72.8958
R17415 vdd.n2582 vdd.n937 72.8958
R17416 vdd.n2582 vdd.n938 72.8958
R17417 vdd.n2582 vdd.n939 72.8958
R17418 vdd.n2855 vdd.n2854 72.8958
R17419 vdd.n2855 vdd.n2583 72.8958
R17420 vdd.n2855 vdd.n2584 72.8958
R17421 vdd.n2855 vdd.n2585 72.8958
R17422 vdd.n2855 vdd.n2586 72.8958
R17423 vdd.n2855 vdd.n2587 72.8958
R17424 vdd.n2855 vdd.n2588 72.8958
R17425 vdd.n2855 vdd.n2589 72.8958
R17426 vdd.n2855 vdd.n2590 72.8958
R17427 vdd.n2855 vdd.n2591 72.8958
R17428 vdd.n2855 vdd.n2592 72.8958
R17429 vdd.n2855 vdd.n2593 72.8958
R17430 vdd.n2855 vdd.n2594 72.8958
R17431 vdd.n2855 vdd.n2595 72.8958
R17432 vdd.n2855 vdd.n2596 72.8958
R17433 vdd.n2855 vdd.n2597 72.8958
R17434 vdd.n2855 vdd.n2598 72.8958
R17435 vdd.n3003 vdd.n756 72.8958
R17436 vdd.n3009 vdd.n756 72.8958
R17437 vdd.n802 vdd.n756 72.8958
R17438 vdd.n3016 vdd.n756 72.8958
R17439 vdd.n799 vdd.n756 72.8958
R17440 vdd.n3023 vdd.n756 72.8958
R17441 vdd.n796 vdd.n756 72.8958
R17442 vdd.n3030 vdd.n756 72.8958
R17443 vdd.n793 vdd.n756 72.8958
R17444 vdd.n3038 vdd.n756 72.8958
R17445 vdd.n790 vdd.n756 72.8958
R17446 vdd.n3045 vdd.n756 72.8958
R17447 vdd.n787 vdd.n756 72.8958
R17448 vdd.n3052 vdd.n756 72.8958
R17449 vdd.n784 vdd.n756 72.8958
R17450 vdd.n3059 vdd.n756 72.8958
R17451 vdd.n3062 vdd.n756 72.8958
R17452 vdd.n2582 vdd.n921 72.8958
R17453 vdd.n2582 vdd.n920 72.8958
R17454 vdd.n2582 vdd.n919 72.8958
R17455 vdd.n2582 vdd.n918 72.8958
R17456 vdd.n2582 vdd.n917 72.8958
R17457 vdd.n2582 vdd.n916 72.8958
R17458 vdd.n2582 vdd.n915 72.8958
R17459 vdd.n2582 vdd.n914 72.8958
R17460 vdd.n2582 vdd.n913 72.8958
R17461 vdd.n2582 vdd.n912 72.8958
R17462 vdd.n2582 vdd.n911 72.8958
R17463 vdd.n2582 vdd.n910 72.8958
R17464 vdd.n2582 vdd.n909 72.8958
R17465 vdd.n2582 vdd.n908 72.8958
R17466 vdd.n2582 vdd.n907 72.8958
R17467 vdd.n2582 vdd.n906 72.8958
R17468 vdd.n2582 vdd.n905 72.8958
R17469 vdd.n2335 vdd.n2334 72.8958
R17470 vdd.n2334 vdd.n1071 72.8958
R17471 vdd.n2334 vdd.n1072 72.8958
R17472 vdd.n2334 vdd.n1073 72.8958
R17473 vdd.n2334 vdd.n1074 72.8958
R17474 vdd.n2334 vdd.n1075 72.8958
R17475 vdd.n2334 vdd.n1076 72.8958
R17476 vdd.n2334 vdd.n1077 72.8958
R17477 vdd.n2334 vdd.n1078 72.8958
R17478 vdd.n2334 vdd.n1079 72.8958
R17479 vdd.n2334 vdd.n1080 72.8958
R17480 vdd.n2334 vdd.n1081 72.8958
R17481 vdd.n2334 vdd.n1082 72.8958
R17482 vdd.n2334 vdd.n1083 72.8958
R17483 vdd.n2334 vdd.n1084 72.8958
R17484 vdd.n2334 vdd.n1085 72.8958
R17485 vdd.n2334 vdd.n1086 72.8958
R17486 vdd.n1736 vdd.n1735 66.2847
R17487 vdd.n1736 vdd.n1514 66.2847
R17488 vdd.n1736 vdd.n1515 66.2847
R17489 vdd.n1736 vdd.n1516 66.2847
R17490 vdd.n1736 vdd.n1517 66.2847
R17491 vdd.n1736 vdd.n1518 66.2847
R17492 vdd.n1736 vdd.n1519 66.2847
R17493 vdd.n1736 vdd.n1520 66.2847
R17494 vdd.n1736 vdd.n1521 66.2847
R17495 vdd.n1736 vdd.n1522 66.2847
R17496 vdd.n1736 vdd.n1523 66.2847
R17497 vdd.n1736 vdd.n1524 66.2847
R17498 vdd.n1736 vdd.n1525 66.2847
R17499 vdd.n1736 vdd.n1526 66.2847
R17500 vdd.n1736 vdd.n1527 66.2847
R17501 vdd.n1736 vdd.n1528 66.2847
R17502 vdd.n1736 vdd.n1529 66.2847
R17503 vdd.n1736 vdd.n1530 66.2847
R17504 vdd.n1736 vdd.n1531 66.2847
R17505 vdd.n1736 vdd.n1532 66.2847
R17506 vdd.n1736 vdd.n1533 66.2847
R17507 vdd.n1736 vdd.n1534 66.2847
R17508 vdd.n1736 vdd.n1535 66.2847
R17509 vdd.n1736 vdd.n1536 66.2847
R17510 vdd.n1736 vdd.n1537 66.2847
R17511 vdd.n1736 vdd.n1538 66.2847
R17512 vdd.n1736 vdd.n1539 66.2847
R17513 vdd.n1736 vdd.n1540 66.2847
R17514 vdd.n1736 vdd.n1541 66.2847
R17515 vdd.n1736 vdd.n1542 66.2847
R17516 vdd.n1736 vdd.n1543 66.2847
R17517 vdd.n1404 vdd.n1054 66.2847
R17518 vdd.n1401 vdd.n1054 66.2847
R17519 vdd.n1397 vdd.n1054 66.2847
R17520 vdd.n2196 vdd.n1054 66.2847
R17521 vdd.n1188 vdd.n1054 66.2847
R17522 vdd.n2203 vdd.n1054 66.2847
R17523 vdd.n1181 vdd.n1054 66.2847
R17524 vdd.n2210 vdd.n1054 66.2847
R17525 vdd.n1174 vdd.n1054 66.2847
R17526 vdd.n2217 vdd.n1054 66.2847
R17527 vdd.n1168 vdd.n1054 66.2847
R17528 vdd.n1163 vdd.n1054 66.2847
R17529 vdd.n2228 vdd.n1054 66.2847
R17530 vdd.n1155 vdd.n1054 66.2847
R17531 vdd.n2235 vdd.n1054 66.2847
R17532 vdd.n1148 vdd.n1054 66.2847
R17533 vdd.n2242 vdd.n1054 66.2847
R17534 vdd.n1141 vdd.n1054 66.2847
R17535 vdd.n2249 vdd.n1054 66.2847
R17536 vdd.n1134 vdd.n1054 66.2847
R17537 vdd.n2256 vdd.n1054 66.2847
R17538 vdd.n1128 vdd.n1054 66.2847
R17539 vdd.n1123 vdd.n1054 66.2847
R17540 vdd.n2267 vdd.n1054 66.2847
R17541 vdd.n1115 vdd.n1054 66.2847
R17542 vdd.n2274 vdd.n1054 66.2847
R17543 vdd.n1108 vdd.n1054 66.2847
R17544 vdd.n2281 vdd.n1054 66.2847
R17545 vdd.n1101 vdd.n1054 66.2847
R17546 vdd.n2288 vdd.n1054 66.2847
R17547 vdd.n2293 vdd.n1054 66.2847
R17548 vdd.n1097 vdd.n1054 66.2847
R17549 vdd.n3229 vdd.n658 66.2847
R17550 vdd.n663 vdd.n658 66.2847
R17551 vdd.n666 vdd.n658 66.2847
R17552 vdd.n3218 vdd.n658 66.2847
R17553 vdd.n3212 vdd.n658 66.2847
R17554 vdd.n3210 vdd.n658 66.2847
R17555 vdd.n3204 vdd.n658 66.2847
R17556 vdd.n3202 vdd.n658 66.2847
R17557 vdd.n3196 vdd.n658 66.2847
R17558 vdd.n3194 vdd.n658 66.2847
R17559 vdd.n3188 vdd.n658 66.2847
R17560 vdd.n3186 vdd.n658 66.2847
R17561 vdd.n3180 vdd.n658 66.2847
R17562 vdd.n3178 vdd.n658 66.2847
R17563 vdd.n3172 vdd.n658 66.2847
R17564 vdd.n3170 vdd.n658 66.2847
R17565 vdd.n3164 vdd.n658 66.2847
R17566 vdd.n3162 vdd.n658 66.2847
R17567 vdd.n3156 vdd.n658 66.2847
R17568 vdd.n3154 vdd.n658 66.2847
R17569 vdd.n727 vdd.n658 66.2847
R17570 vdd.n3145 vdd.n658 66.2847
R17571 vdd.n729 vdd.n658 66.2847
R17572 vdd.n3138 vdd.n658 66.2847
R17573 vdd.n3132 vdd.n658 66.2847
R17574 vdd.n3130 vdd.n658 66.2847
R17575 vdd.n3124 vdd.n658 66.2847
R17576 vdd.n3122 vdd.n658 66.2847
R17577 vdd.n3116 vdd.n658 66.2847
R17578 vdd.n750 vdd.n658 66.2847
R17579 vdd.n752 vdd.n658 66.2847
R17580 vdd.n3345 vdd.n3344 66.2847
R17581 vdd.n3345 vdd.n403 66.2847
R17582 vdd.n3345 vdd.n402 66.2847
R17583 vdd.n3345 vdd.n401 66.2847
R17584 vdd.n3345 vdd.n400 66.2847
R17585 vdd.n3345 vdd.n399 66.2847
R17586 vdd.n3345 vdd.n398 66.2847
R17587 vdd.n3345 vdd.n397 66.2847
R17588 vdd.n3345 vdd.n396 66.2847
R17589 vdd.n3345 vdd.n395 66.2847
R17590 vdd.n3345 vdd.n394 66.2847
R17591 vdd.n3345 vdd.n393 66.2847
R17592 vdd.n3345 vdd.n392 66.2847
R17593 vdd.n3345 vdd.n391 66.2847
R17594 vdd.n3345 vdd.n390 66.2847
R17595 vdd.n3345 vdd.n389 66.2847
R17596 vdd.n3345 vdd.n388 66.2847
R17597 vdd.n3345 vdd.n387 66.2847
R17598 vdd.n3345 vdd.n386 66.2847
R17599 vdd.n3345 vdd.n385 66.2847
R17600 vdd.n3345 vdd.n384 66.2847
R17601 vdd.n3345 vdd.n383 66.2847
R17602 vdd.n3345 vdd.n382 66.2847
R17603 vdd.n3345 vdd.n381 66.2847
R17604 vdd.n3345 vdd.n380 66.2847
R17605 vdd.n3345 vdd.n379 66.2847
R17606 vdd.n3345 vdd.n378 66.2847
R17607 vdd.n3345 vdd.n377 66.2847
R17608 vdd.n3345 vdd.n376 66.2847
R17609 vdd.n3345 vdd.n375 66.2847
R17610 vdd.n3345 vdd.n374 66.2847
R17611 vdd.n3345 vdd.n373 66.2847
R17612 vdd.n448 vdd.n373 52.4337
R17613 vdd.n454 vdd.n374 52.4337
R17614 vdd.n458 vdd.n375 52.4337
R17615 vdd.n464 vdd.n376 52.4337
R17616 vdd.n468 vdd.n377 52.4337
R17617 vdd.n474 vdd.n378 52.4337
R17618 vdd.n478 vdd.n379 52.4337
R17619 vdd.n484 vdd.n380 52.4337
R17620 vdd.n488 vdd.n381 52.4337
R17621 vdd.n494 vdd.n382 52.4337
R17622 vdd.n498 vdd.n383 52.4337
R17623 vdd.n504 vdd.n384 52.4337
R17624 vdd.n508 vdd.n385 52.4337
R17625 vdd.n514 vdd.n386 52.4337
R17626 vdd.n518 vdd.n387 52.4337
R17627 vdd.n524 vdd.n388 52.4337
R17628 vdd.n528 vdd.n389 52.4337
R17629 vdd.n534 vdd.n390 52.4337
R17630 vdd.n538 vdd.n391 52.4337
R17631 vdd.n544 vdd.n392 52.4337
R17632 vdd.n548 vdd.n393 52.4337
R17633 vdd.n554 vdd.n394 52.4337
R17634 vdd.n558 vdd.n395 52.4337
R17635 vdd.n564 vdd.n396 52.4337
R17636 vdd.n568 vdd.n397 52.4337
R17637 vdd.n574 vdd.n398 52.4337
R17638 vdd.n578 vdd.n399 52.4337
R17639 vdd.n584 vdd.n400 52.4337
R17640 vdd.n588 vdd.n401 52.4337
R17641 vdd.n594 vdd.n402 52.4337
R17642 vdd.n597 vdd.n403 52.4337
R17643 vdd.n3344 vdd.n3343 52.4337
R17644 vdd.n3229 vdd.n660 52.4337
R17645 vdd.n3227 vdd.n663 52.4337
R17646 vdd.n3223 vdd.n666 52.4337
R17647 vdd.n3219 vdd.n3218 52.4337
R17648 vdd.n3212 vdd.n669 52.4337
R17649 vdd.n3211 vdd.n3210 52.4337
R17650 vdd.n3204 vdd.n675 52.4337
R17651 vdd.n3203 vdd.n3202 52.4337
R17652 vdd.n3196 vdd.n681 52.4337
R17653 vdd.n3195 vdd.n3194 52.4337
R17654 vdd.n3188 vdd.n689 52.4337
R17655 vdd.n3187 vdd.n3186 52.4337
R17656 vdd.n3180 vdd.n695 52.4337
R17657 vdd.n3179 vdd.n3178 52.4337
R17658 vdd.n3172 vdd.n701 52.4337
R17659 vdd.n3171 vdd.n3170 52.4337
R17660 vdd.n3164 vdd.n707 52.4337
R17661 vdd.n3163 vdd.n3162 52.4337
R17662 vdd.n3156 vdd.n713 52.4337
R17663 vdd.n3155 vdd.n3154 52.4337
R17664 vdd.n727 vdd.n719 52.4337
R17665 vdd.n3146 vdd.n3145 52.4337
R17666 vdd.n3143 vdd.n729 52.4337
R17667 vdd.n3139 vdd.n3138 52.4337
R17668 vdd.n3132 vdd.n733 52.4337
R17669 vdd.n3131 vdd.n3130 52.4337
R17670 vdd.n3124 vdd.n739 52.4337
R17671 vdd.n3123 vdd.n3122 52.4337
R17672 vdd.n3116 vdd.n745 52.4337
R17673 vdd.n3115 vdd.n750 52.4337
R17674 vdd.n3111 vdd.n752 52.4337
R17675 vdd.n2295 vdd.n1097 52.4337
R17676 vdd.n2293 vdd.n2292 52.4337
R17677 vdd.n2288 vdd.n2287 52.4337
R17678 vdd.n2283 vdd.n1101 52.4337
R17679 vdd.n2281 vdd.n2280 52.4337
R17680 vdd.n2276 vdd.n1108 52.4337
R17681 vdd.n2274 vdd.n2273 52.4337
R17682 vdd.n2269 vdd.n1115 52.4337
R17683 vdd.n2267 vdd.n2266 52.4337
R17684 vdd.n1124 vdd.n1123 52.4337
R17685 vdd.n2258 vdd.n1128 52.4337
R17686 vdd.n2256 vdd.n2255 52.4337
R17687 vdd.n2251 vdd.n1134 52.4337
R17688 vdd.n2249 vdd.n2248 52.4337
R17689 vdd.n2244 vdd.n1141 52.4337
R17690 vdd.n2242 vdd.n2241 52.4337
R17691 vdd.n2237 vdd.n1148 52.4337
R17692 vdd.n2235 vdd.n2234 52.4337
R17693 vdd.n2230 vdd.n1155 52.4337
R17694 vdd.n2228 vdd.n2227 52.4337
R17695 vdd.n1164 vdd.n1163 52.4337
R17696 vdd.n2219 vdd.n1168 52.4337
R17697 vdd.n2217 vdd.n2216 52.4337
R17698 vdd.n2212 vdd.n1174 52.4337
R17699 vdd.n2210 vdd.n2209 52.4337
R17700 vdd.n2205 vdd.n1181 52.4337
R17701 vdd.n2203 vdd.n2202 52.4337
R17702 vdd.n2198 vdd.n1188 52.4337
R17703 vdd.n2196 vdd.n2195 52.4337
R17704 vdd.n1398 vdd.n1397 52.4337
R17705 vdd.n1402 vdd.n1401 52.4337
R17706 vdd.n2184 vdd.n1404 52.4337
R17707 vdd.n1735 vdd.n1734 52.4337
R17708 vdd.n1549 vdd.n1514 52.4337
R17709 vdd.n1551 vdd.n1515 52.4337
R17710 vdd.n1555 vdd.n1516 52.4337
R17711 vdd.n1557 vdd.n1517 52.4337
R17712 vdd.n1561 vdd.n1518 52.4337
R17713 vdd.n1563 vdd.n1519 52.4337
R17714 vdd.n1567 vdd.n1520 52.4337
R17715 vdd.n1569 vdd.n1521 52.4337
R17716 vdd.n1701 vdd.n1522 52.4337
R17717 vdd.n1573 vdd.n1523 52.4337
R17718 vdd.n1577 vdd.n1524 52.4337
R17719 vdd.n1579 vdd.n1525 52.4337
R17720 vdd.n1583 vdd.n1526 52.4337
R17721 vdd.n1585 vdd.n1527 52.4337
R17722 vdd.n1589 vdd.n1528 52.4337
R17723 vdd.n1591 vdd.n1529 52.4337
R17724 vdd.n1595 vdd.n1530 52.4337
R17725 vdd.n1597 vdd.n1531 52.4337
R17726 vdd.n1601 vdd.n1532 52.4337
R17727 vdd.n1665 vdd.n1533 52.4337
R17728 vdd.n1606 vdd.n1534 52.4337
R17729 vdd.n1608 vdd.n1535 52.4337
R17730 vdd.n1612 vdd.n1536 52.4337
R17731 vdd.n1614 vdd.n1537 52.4337
R17732 vdd.n1618 vdd.n1538 52.4337
R17733 vdd.n1620 vdd.n1539 52.4337
R17734 vdd.n1624 vdd.n1540 52.4337
R17735 vdd.n1626 vdd.n1541 52.4337
R17736 vdd.n1630 vdd.n1542 52.4337
R17737 vdd.n1632 vdd.n1543 52.4337
R17738 vdd.n1735 vdd.n1545 52.4337
R17739 vdd.n1550 vdd.n1514 52.4337
R17740 vdd.n1554 vdd.n1515 52.4337
R17741 vdd.n1556 vdd.n1516 52.4337
R17742 vdd.n1560 vdd.n1517 52.4337
R17743 vdd.n1562 vdd.n1518 52.4337
R17744 vdd.n1566 vdd.n1519 52.4337
R17745 vdd.n1568 vdd.n1520 52.4337
R17746 vdd.n1700 vdd.n1521 52.4337
R17747 vdd.n1572 vdd.n1522 52.4337
R17748 vdd.n1576 vdd.n1523 52.4337
R17749 vdd.n1578 vdd.n1524 52.4337
R17750 vdd.n1582 vdd.n1525 52.4337
R17751 vdd.n1584 vdd.n1526 52.4337
R17752 vdd.n1588 vdd.n1527 52.4337
R17753 vdd.n1590 vdd.n1528 52.4337
R17754 vdd.n1594 vdd.n1529 52.4337
R17755 vdd.n1596 vdd.n1530 52.4337
R17756 vdd.n1600 vdd.n1531 52.4337
R17757 vdd.n1602 vdd.n1532 52.4337
R17758 vdd.n1605 vdd.n1533 52.4337
R17759 vdd.n1607 vdd.n1534 52.4337
R17760 vdd.n1611 vdd.n1535 52.4337
R17761 vdd.n1613 vdd.n1536 52.4337
R17762 vdd.n1617 vdd.n1537 52.4337
R17763 vdd.n1619 vdd.n1538 52.4337
R17764 vdd.n1623 vdd.n1539 52.4337
R17765 vdd.n1625 vdd.n1540 52.4337
R17766 vdd.n1629 vdd.n1541 52.4337
R17767 vdd.n1631 vdd.n1542 52.4337
R17768 vdd.n1543 vdd.n1513 52.4337
R17769 vdd.n1404 vdd.n1403 52.4337
R17770 vdd.n1401 vdd.n1400 52.4337
R17771 vdd.n1397 vdd.n1189 52.4337
R17772 vdd.n2197 vdd.n2196 52.4337
R17773 vdd.n1188 vdd.n1182 52.4337
R17774 vdd.n2204 vdd.n2203 52.4337
R17775 vdd.n1181 vdd.n1175 52.4337
R17776 vdd.n2211 vdd.n2210 52.4337
R17777 vdd.n1174 vdd.n1169 52.4337
R17778 vdd.n2218 vdd.n2217 52.4337
R17779 vdd.n1168 vdd.n1167 52.4337
R17780 vdd.n1163 vdd.n1156 52.4337
R17781 vdd.n2229 vdd.n2228 52.4337
R17782 vdd.n1155 vdd.n1149 52.4337
R17783 vdd.n2236 vdd.n2235 52.4337
R17784 vdd.n1148 vdd.n1142 52.4337
R17785 vdd.n2243 vdd.n2242 52.4337
R17786 vdd.n1141 vdd.n1135 52.4337
R17787 vdd.n2250 vdd.n2249 52.4337
R17788 vdd.n1134 vdd.n1129 52.4337
R17789 vdd.n2257 vdd.n2256 52.4337
R17790 vdd.n1128 vdd.n1127 52.4337
R17791 vdd.n1123 vdd.n1116 52.4337
R17792 vdd.n2268 vdd.n2267 52.4337
R17793 vdd.n1115 vdd.n1109 52.4337
R17794 vdd.n2275 vdd.n2274 52.4337
R17795 vdd.n1108 vdd.n1102 52.4337
R17796 vdd.n2282 vdd.n2281 52.4337
R17797 vdd.n1101 vdd.n1098 52.4337
R17798 vdd.n2289 vdd.n2288 52.4337
R17799 vdd.n2294 vdd.n2293 52.4337
R17800 vdd.n1409 vdd.n1097 52.4337
R17801 vdd.n3230 vdd.n3229 52.4337
R17802 vdd.n3224 vdd.n663 52.4337
R17803 vdd.n3220 vdd.n666 52.4337
R17804 vdd.n3218 vdd.n3217 52.4337
R17805 vdd.n3213 vdd.n3212 52.4337
R17806 vdd.n3210 vdd.n3209 52.4337
R17807 vdd.n3205 vdd.n3204 52.4337
R17808 vdd.n3202 vdd.n3201 52.4337
R17809 vdd.n3197 vdd.n3196 52.4337
R17810 vdd.n3194 vdd.n3193 52.4337
R17811 vdd.n3189 vdd.n3188 52.4337
R17812 vdd.n3186 vdd.n3185 52.4337
R17813 vdd.n3181 vdd.n3180 52.4337
R17814 vdd.n3178 vdd.n3177 52.4337
R17815 vdd.n3173 vdd.n3172 52.4337
R17816 vdd.n3170 vdd.n3169 52.4337
R17817 vdd.n3165 vdd.n3164 52.4337
R17818 vdd.n3162 vdd.n3161 52.4337
R17819 vdd.n3157 vdd.n3156 52.4337
R17820 vdd.n3154 vdd.n3153 52.4337
R17821 vdd.n728 vdd.n727 52.4337
R17822 vdd.n3145 vdd.n3144 52.4337
R17823 vdd.n3140 vdd.n729 52.4337
R17824 vdd.n3138 vdd.n3137 52.4337
R17825 vdd.n3133 vdd.n3132 52.4337
R17826 vdd.n3130 vdd.n3129 52.4337
R17827 vdd.n3125 vdd.n3124 52.4337
R17828 vdd.n3122 vdd.n3121 52.4337
R17829 vdd.n3117 vdd.n3116 52.4337
R17830 vdd.n3112 vdd.n750 52.4337
R17831 vdd.n3108 vdd.n752 52.4337
R17832 vdd.n3344 vdd.n404 52.4337
R17833 vdd.n595 vdd.n403 52.4337
R17834 vdd.n589 vdd.n402 52.4337
R17835 vdd.n585 vdd.n401 52.4337
R17836 vdd.n579 vdd.n400 52.4337
R17837 vdd.n575 vdd.n399 52.4337
R17838 vdd.n569 vdd.n398 52.4337
R17839 vdd.n565 vdd.n397 52.4337
R17840 vdd.n559 vdd.n396 52.4337
R17841 vdd.n555 vdd.n395 52.4337
R17842 vdd.n549 vdd.n394 52.4337
R17843 vdd.n545 vdd.n393 52.4337
R17844 vdd.n539 vdd.n392 52.4337
R17845 vdd.n535 vdd.n391 52.4337
R17846 vdd.n529 vdd.n390 52.4337
R17847 vdd.n525 vdd.n389 52.4337
R17848 vdd.n519 vdd.n388 52.4337
R17849 vdd.n515 vdd.n387 52.4337
R17850 vdd.n509 vdd.n386 52.4337
R17851 vdd.n505 vdd.n385 52.4337
R17852 vdd.n499 vdd.n384 52.4337
R17853 vdd.n495 vdd.n383 52.4337
R17854 vdd.n489 vdd.n382 52.4337
R17855 vdd.n485 vdd.n381 52.4337
R17856 vdd.n479 vdd.n380 52.4337
R17857 vdd.n475 vdd.n379 52.4337
R17858 vdd.n469 vdd.n378 52.4337
R17859 vdd.n465 vdd.n377 52.4337
R17860 vdd.n459 vdd.n376 52.4337
R17861 vdd.n455 vdd.n375 52.4337
R17862 vdd.n449 vdd.n374 52.4337
R17863 vdd.n445 vdd.n373 52.4337
R17864 vdd.t101 vdd.t258 51.4683
R17865 vdd.n266 vdd.n264 42.0461
R17866 vdd.n168 vdd.n166 42.0461
R17867 vdd.n71 vdd.n69 42.0461
R17868 vdd.n2052 vdd.n2050 42.0461
R17869 vdd.n1954 vdd.n1952 42.0461
R17870 vdd.n1857 vdd.n1855 42.0461
R17871 vdd.n320 vdd.n319 41.6884
R17872 vdd.n222 vdd.n221 41.6884
R17873 vdd.n125 vdd.n124 41.6884
R17874 vdd.n2106 vdd.n2105 41.6884
R17875 vdd.n2008 vdd.n2007 41.6884
R17876 vdd.n1911 vdd.n1910 41.6884
R17877 vdd.n1512 vdd.n1511 41.1157
R17878 vdd.n1668 vdd.n1667 41.1157
R17879 vdd.n1704 vdd.n1703 41.1157
R17880 vdd.n407 vdd.n406 41.1157
R17881 vdd.n547 vdd.n420 41.1157
R17882 vdd.n433 vdd.n432 41.1157
R17883 vdd.n3062 vdd.n3061 39.2114
R17884 vdd.n3059 vdd.n3058 39.2114
R17885 vdd.n3054 vdd.n784 39.2114
R17886 vdd.n3052 vdd.n3051 39.2114
R17887 vdd.n3047 vdd.n787 39.2114
R17888 vdd.n3045 vdd.n3044 39.2114
R17889 vdd.n3040 vdd.n790 39.2114
R17890 vdd.n3038 vdd.n3037 39.2114
R17891 vdd.n3032 vdd.n793 39.2114
R17892 vdd.n3030 vdd.n3029 39.2114
R17893 vdd.n3025 vdd.n796 39.2114
R17894 vdd.n3023 vdd.n3022 39.2114
R17895 vdd.n3018 vdd.n799 39.2114
R17896 vdd.n3016 vdd.n3015 39.2114
R17897 vdd.n3011 vdd.n802 39.2114
R17898 vdd.n3009 vdd.n3008 39.2114
R17899 vdd.n3004 vdd.n3003 39.2114
R17900 vdd.n2854 vdd.n2853 39.2114
R17901 vdd.n2848 vdd.n2583 39.2114
R17902 vdd.n2845 vdd.n2584 39.2114
R17903 vdd.n2841 vdd.n2585 39.2114
R17904 vdd.n2837 vdd.n2586 39.2114
R17905 vdd.n2833 vdd.n2587 39.2114
R17906 vdd.n2829 vdd.n2588 39.2114
R17907 vdd.n2825 vdd.n2589 39.2114
R17908 vdd.n2821 vdd.n2590 39.2114
R17909 vdd.n2817 vdd.n2591 39.2114
R17910 vdd.n2813 vdd.n2592 39.2114
R17911 vdd.n2809 vdd.n2593 39.2114
R17912 vdd.n2805 vdd.n2594 39.2114
R17913 vdd.n2801 vdd.n2595 39.2114
R17914 vdd.n2797 vdd.n2596 39.2114
R17915 vdd.n2793 vdd.n2597 39.2114
R17916 vdd.n2788 vdd.n2598 39.2114
R17917 vdd.n2577 vdd.n939 39.2114
R17918 vdd.n2573 vdd.n938 39.2114
R17919 vdd.n2569 vdd.n937 39.2114
R17920 vdd.n2565 vdd.n936 39.2114
R17921 vdd.n2561 vdd.n935 39.2114
R17922 vdd.n2557 vdd.n934 39.2114
R17923 vdd.n2553 vdd.n933 39.2114
R17924 vdd.n2549 vdd.n932 39.2114
R17925 vdd.n2545 vdd.n931 39.2114
R17926 vdd.n2541 vdd.n930 39.2114
R17927 vdd.n2537 vdd.n929 39.2114
R17928 vdd.n2533 vdd.n928 39.2114
R17929 vdd.n2529 vdd.n927 39.2114
R17930 vdd.n2525 vdd.n926 39.2114
R17931 vdd.n2521 vdd.n925 39.2114
R17932 vdd.n2516 vdd.n924 39.2114
R17933 vdd.n2512 vdd.n923 39.2114
R17934 vdd.n2333 vdd.n2332 39.2114
R17935 vdd.n2327 vdd.n1055 39.2114
R17936 vdd.n2324 vdd.n1056 39.2114
R17937 vdd.n2320 vdd.n1057 39.2114
R17938 vdd.n2316 vdd.n1058 39.2114
R17939 vdd.n2312 vdd.n1059 39.2114
R17940 vdd.n2308 vdd.n1060 39.2114
R17941 vdd.n2304 vdd.n1061 39.2114
R17942 vdd.n2300 vdd.n1062 39.2114
R17943 vdd.n1247 vdd.n1063 39.2114
R17944 vdd.n1251 vdd.n1064 39.2114
R17945 vdd.n1255 vdd.n1065 39.2114
R17946 vdd.n1259 vdd.n1066 39.2114
R17947 vdd.n1263 vdd.n1067 39.2114
R17948 vdd.n1267 vdd.n1068 39.2114
R17949 vdd.n1271 vdd.n1069 39.2114
R17950 vdd.n1276 vdd.n1070 39.2114
R17951 vdd.n2981 vdd.n2980 39.2114
R17952 vdd.n2976 vdd.n2948 39.2114
R17953 vdd.n2974 vdd.n2973 39.2114
R17954 vdd.n2969 vdd.n2951 39.2114
R17955 vdd.n2967 vdd.n2966 39.2114
R17956 vdd.n2962 vdd.n2954 39.2114
R17957 vdd.n2960 vdd.n2959 39.2114
R17958 vdd.n2955 vdd.n755 39.2114
R17959 vdd.n3099 vdd.n3098 39.2114
R17960 vdd.n3096 vdd.n3095 39.2114
R17961 vdd.n3091 vdd.n760 39.2114
R17962 vdd.n3089 vdd.n3088 39.2114
R17963 vdd.n3084 vdd.n763 39.2114
R17964 vdd.n3082 vdd.n3081 39.2114
R17965 vdd.n3077 vdd.n766 39.2114
R17966 vdd.n3075 vdd.n3074 39.2114
R17967 vdd.n3070 vdd.n772 39.2114
R17968 vdd.n2857 vdd.n2856 39.2114
R17969 vdd.n2624 vdd.n2599 39.2114
R17970 vdd.n2628 vdd.n2600 39.2114
R17971 vdd.n2632 vdd.n2601 39.2114
R17972 vdd.n2636 vdd.n2602 39.2114
R17973 vdd.n2640 vdd.n2603 39.2114
R17974 vdd.n2644 vdd.n2604 39.2114
R17975 vdd.n2648 vdd.n2605 39.2114
R17976 vdd.n2652 vdd.n2606 39.2114
R17977 vdd.n2656 vdd.n2607 39.2114
R17978 vdd.n2660 vdd.n2608 39.2114
R17979 vdd.n2664 vdd.n2609 39.2114
R17980 vdd.n2668 vdd.n2610 39.2114
R17981 vdd.n2672 vdd.n2611 39.2114
R17982 vdd.n2676 vdd.n2612 39.2114
R17983 vdd.n2680 vdd.n2613 39.2114
R17984 vdd.n2684 vdd.n2614 39.2114
R17985 vdd.n2856 vdd.n904 39.2114
R17986 vdd.n2627 vdd.n2599 39.2114
R17987 vdd.n2631 vdd.n2600 39.2114
R17988 vdd.n2635 vdd.n2601 39.2114
R17989 vdd.n2639 vdd.n2602 39.2114
R17990 vdd.n2643 vdd.n2603 39.2114
R17991 vdd.n2647 vdd.n2604 39.2114
R17992 vdd.n2651 vdd.n2605 39.2114
R17993 vdd.n2655 vdd.n2606 39.2114
R17994 vdd.n2659 vdd.n2607 39.2114
R17995 vdd.n2663 vdd.n2608 39.2114
R17996 vdd.n2667 vdd.n2609 39.2114
R17997 vdd.n2671 vdd.n2610 39.2114
R17998 vdd.n2675 vdd.n2611 39.2114
R17999 vdd.n2679 vdd.n2612 39.2114
R18000 vdd.n2683 vdd.n2613 39.2114
R18001 vdd.n2686 vdd.n2614 39.2114
R18002 vdd.n772 vdd.n767 39.2114
R18003 vdd.n3076 vdd.n3075 39.2114
R18004 vdd.n766 vdd.n764 39.2114
R18005 vdd.n3083 vdd.n3082 39.2114
R18006 vdd.n763 vdd.n761 39.2114
R18007 vdd.n3090 vdd.n3089 39.2114
R18008 vdd.n760 vdd.n758 39.2114
R18009 vdd.n3097 vdd.n3096 39.2114
R18010 vdd.n3100 vdd.n3099 39.2114
R18011 vdd.n2956 vdd.n2955 39.2114
R18012 vdd.n2961 vdd.n2960 39.2114
R18013 vdd.n2954 vdd.n2952 39.2114
R18014 vdd.n2968 vdd.n2967 39.2114
R18015 vdd.n2951 vdd.n2949 39.2114
R18016 vdd.n2975 vdd.n2974 39.2114
R18017 vdd.n2948 vdd.n2946 39.2114
R18018 vdd.n2982 vdd.n2981 39.2114
R18019 vdd.n2333 vdd.n1089 39.2114
R18020 vdd.n2325 vdd.n1055 39.2114
R18021 vdd.n2321 vdd.n1056 39.2114
R18022 vdd.n2317 vdd.n1057 39.2114
R18023 vdd.n2313 vdd.n1058 39.2114
R18024 vdd.n2309 vdd.n1059 39.2114
R18025 vdd.n2305 vdd.n1060 39.2114
R18026 vdd.n2301 vdd.n1061 39.2114
R18027 vdd.n1246 vdd.n1062 39.2114
R18028 vdd.n1250 vdd.n1063 39.2114
R18029 vdd.n1254 vdd.n1064 39.2114
R18030 vdd.n1258 vdd.n1065 39.2114
R18031 vdd.n1262 vdd.n1066 39.2114
R18032 vdd.n1266 vdd.n1067 39.2114
R18033 vdd.n1270 vdd.n1068 39.2114
R18034 vdd.n1275 vdd.n1069 39.2114
R18035 vdd.n1279 vdd.n1070 39.2114
R18036 vdd.n2515 vdd.n923 39.2114
R18037 vdd.n2520 vdd.n924 39.2114
R18038 vdd.n2524 vdd.n925 39.2114
R18039 vdd.n2528 vdd.n926 39.2114
R18040 vdd.n2532 vdd.n927 39.2114
R18041 vdd.n2536 vdd.n928 39.2114
R18042 vdd.n2540 vdd.n929 39.2114
R18043 vdd.n2544 vdd.n930 39.2114
R18044 vdd.n2548 vdd.n931 39.2114
R18045 vdd.n2552 vdd.n932 39.2114
R18046 vdd.n2556 vdd.n933 39.2114
R18047 vdd.n2560 vdd.n934 39.2114
R18048 vdd.n2564 vdd.n935 39.2114
R18049 vdd.n2568 vdd.n936 39.2114
R18050 vdd.n2572 vdd.n937 39.2114
R18051 vdd.n2576 vdd.n938 39.2114
R18052 vdd.n941 vdd.n939 39.2114
R18053 vdd.n2854 vdd.n2617 39.2114
R18054 vdd.n2846 vdd.n2583 39.2114
R18055 vdd.n2842 vdd.n2584 39.2114
R18056 vdd.n2838 vdd.n2585 39.2114
R18057 vdd.n2834 vdd.n2586 39.2114
R18058 vdd.n2830 vdd.n2587 39.2114
R18059 vdd.n2826 vdd.n2588 39.2114
R18060 vdd.n2822 vdd.n2589 39.2114
R18061 vdd.n2818 vdd.n2590 39.2114
R18062 vdd.n2814 vdd.n2591 39.2114
R18063 vdd.n2810 vdd.n2592 39.2114
R18064 vdd.n2806 vdd.n2593 39.2114
R18065 vdd.n2802 vdd.n2594 39.2114
R18066 vdd.n2798 vdd.n2595 39.2114
R18067 vdd.n2794 vdd.n2596 39.2114
R18068 vdd.n2789 vdd.n2597 39.2114
R18069 vdd.n2785 vdd.n2598 39.2114
R18070 vdd.n3003 vdd.n803 39.2114
R18071 vdd.n3010 vdd.n3009 39.2114
R18072 vdd.n802 vdd.n800 39.2114
R18073 vdd.n3017 vdd.n3016 39.2114
R18074 vdd.n799 vdd.n797 39.2114
R18075 vdd.n3024 vdd.n3023 39.2114
R18076 vdd.n796 vdd.n794 39.2114
R18077 vdd.n3031 vdd.n3030 39.2114
R18078 vdd.n793 vdd.n791 39.2114
R18079 vdd.n3039 vdd.n3038 39.2114
R18080 vdd.n790 vdd.n788 39.2114
R18081 vdd.n3046 vdd.n3045 39.2114
R18082 vdd.n787 vdd.n785 39.2114
R18083 vdd.n3053 vdd.n3052 39.2114
R18084 vdd.n784 vdd.n782 39.2114
R18085 vdd.n3060 vdd.n3059 39.2114
R18086 vdd.n3063 vdd.n3062 39.2114
R18087 vdd.n950 vdd.n905 39.2114
R18088 vdd.n2504 vdd.n906 39.2114
R18089 vdd.n2500 vdd.n907 39.2114
R18090 vdd.n2496 vdd.n908 39.2114
R18091 vdd.n2492 vdd.n909 39.2114
R18092 vdd.n2488 vdd.n910 39.2114
R18093 vdd.n2484 vdd.n911 39.2114
R18094 vdd.n2480 vdd.n912 39.2114
R18095 vdd.n2476 vdd.n913 39.2114
R18096 vdd.n2472 vdd.n914 39.2114
R18097 vdd.n2468 vdd.n915 39.2114
R18098 vdd.n2464 vdd.n916 39.2114
R18099 vdd.n2460 vdd.n917 39.2114
R18100 vdd.n2456 vdd.n918 39.2114
R18101 vdd.n2452 vdd.n919 39.2114
R18102 vdd.n2448 vdd.n920 39.2114
R18103 vdd.n2444 vdd.n921 39.2114
R18104 vdd.n2336 vdd.n2335 39.2114
R18105 vdd.n1193 vdd.n1071 39.2114
R18106 vdd.n1197 vdd.n1072 39.2114
R18107 vdd.n1201 vdd.n1073 39.2114
R18108 vdd.n1205 vdd.n1074 39.2114
R18109 vdd.n1209 vdd.n1075 39.2114
R18110 vdd.n1213 vdd.n1076 39.2114
R18111 vdd.n1217 vdd.n1077 39.2114
R18112 vdd.n1221 vdd.n1078 39.2114
R18113 vdd.n1391 vdd.n1079 39.2114
R18114 vdd.n1388 vdd.n1080 39.2114
R18115 vdd.n1384 vdd.n1081 39.2114
R18116 vdd.n1380 vdd.n1082 39.2114
R18117 vdd.n1376 vdd.n1083 39.2114
R18118 vdd.n1372 vdd.n1084 39.2114
R18119 vdd.n1368 vdd.n1085 39.2114
R18120 vdd.n1364 vdd.n1086 39.2114
R18121 vdd.n2441 vdd.n921 39.2114
R18122 vdd.n2445 vdd.n920 39.2114
R18123 vdd.n2449 vdd.n919 39.2114
R18124 vdd.n2453 vdd.n918 39.2114
R18125 vdd.n2457 vdd.n917 39.2114
R18126 vdd.n2461 vdd.n916 39.2114
R18127 vdd.n2465 vdd.n915 39.2114
R18128 vdd.n2469 vdd.n914 39.2114
R18129 vdd.n2473 vdd.n913 39.2114
R18130 vdd.n2477 vdd.n912 39.2114
R18131 vdd.n2481 vdd.n911 39.2114
R18132 vdd.n2485 vdd.n910 39.2114
R18133 vdd.n2489 vdd.n909 39.2114
R18134 vdd.n2493 vdd.n908 39.2114
R18135 vdd.n2497 vdd.n907 39.2114
R18136 vdd.n2501 vdd.n906 39.2114
R18137 vdd.n2505 vdd.n905 39.2114
R18138 vdd.n2335 vdd.n1053 39.2114
R18139 vdd.n1196 vdd.n1071 39.2114
R18140 vdd.n1200 vdd.n1072 39.2114
R18141 vdd.n1204 vdd.n1073 39.2114
R18142 vdd.n1208 vdd.n1074 39.2114
R18143 vdd.n1212 vdd.n1075 39.2114
R18144 vdd.n1216 vdd.n1076 39.2114
R18145 vdd.n1220 vdd.n1077 39.2114
R18146 vdd.n1223 vdd.n1078 39.2114
R18147 vdd.n1389 vdd.n1079 39.2114
R18148 vdd.n1385 vdd.n1080 39.2114
R18149 vdd.n1381 vdd.n1081 39.2114
R18150 vdd.n1377 vdd.n1082 39.2114
R18151 vdd.n1373 vdd.n1083 39.2114
R18152 vdd.n1369 vdd.n1084 39.2114
R18153 vdd.n1365 vdd.n1085 39.2114
R18154 vdd.n1361 vdd.n1086 39.2114
R18155 vdd.n2188 vdd.n2187 37.2369
R18156 vdd.n2224 vdd.n1162 37.2369
R18157 vdd.n2263 vdd.n1122 37.2369
R18158 vdd.n3151 vdd.n724 37.2369
R18159 vdd.n688 vdd.n687 37.2369
R18160 vdd.n3107 vdd.n3106 37.2369
R18161 vdd.n2331 vdd.n1045 31.0639
R18162 vdd.n2580 vdd.n942 31.0639
R18163 vdd.n2513 vdd.n945 31.0639
R18164 vdd.n1281 vdd.n1278 31.0639
R18165 vdd.n2786 vdd.n2783 31.0639
R18166 vdd.n3005 vdd.n3002 31.0639
R18167 vdd.n2852 vdd.n897 31.0639
R18168 vdd.n3066 vdd.n3065 31.0639
R18169 vdd.n2985 vdd.n2984 31.0639
R18170 vdd.n3071 vdd.n771 31.0639
R18171 vdd.n2690 vdd.n2688 31.0639
R18172 vdd.n2859 vdd.n2858 31.0639
R18173 vdd.n2338 vdd.n2337 31.0639
R18174 vdd.n2508 vdd.n2507 31.0639
R18175 vdd.n2440 vdd.n2439 31.0639
R18176 vdd.n1360 vdd.n1359 31.0639
R18177 vdd.n1226 vdd.n1225 30.449
R18178 vdd.n954 vdd.n953 30.449
R18179 vdd.n1273 vdd.n1245 30.449
R18180 vdd.n2518 vdd.n944 30.449
R18181 vdd.n2623 vdd.n2622 30.449
R18182 vdd.n806 vdd.n805 30.449
R18183 vdd.n2791 vdd.n2619 30.449
R18184 vdd.n770 vdd.n769 30.449
R18185 vdd.n1742 vdd.n1508 19.3944
R18186 vdd.n1742 vdd.n1498 19.3944
R18187 vdd.n1754 vdd.n1498 19.3944
R18188 vdd.n1754 vdd.n1496 19.3944
R18189 vdd.n1758 vdd.n1496 19.3944
R18190 vdd.n1758 vdd.n1486 19.3944
R18191 vdd.n1771 vdd.n1486 19.3944
R18192 vdd.n1771 vdd.n1484 19.3944
R18193 vdd.n1775 vdd.n1484 19.3944
R18194 vdd.n1775 vdd.n1476 19.3944
R18195 vdd.n1788 vdd.n1476 19.3944
R18196 vdd.n1788 vdd.n1474 19.3944
R18197 vdd.n1792 vdd.n1474 19.3944
R18198 vdd.n1792 vdd.n1463 19.3944
R18199 vdd.n1804 vdd.n1463 19.3944
R18200 vdd.n1804 vdd.n1461 19.3944
R18201 vdd.n1808 vdd.n1461 19.3944
R18202 vdd.n1808 vdd.n1452 19.3944
R18203 vdd.n2116 vdd.n1452 19.3944
R18204 vdd.n2116 vdd.n1450 19.3944
R18205 vdd.n2120 vdd.n1450 19.3944
R18206 vdd.n2120 vdd.n1441 19.3944
R18207 vdd.n2132 vdd.n1441 19.3944
R18208 vdd.n2132 vdd.n1439 19.3944
R18209 vdd.n2136 vdd.n1439 19.3944
R18210 vdd.n2136 vdd.n1429 19.3944
R18211 vdd.n2149 vdd.n1429 19.3944
R18212 vdd.n2149 vdd.n1427 19.3944
R18213 vdd.n2153 vdd.n1427 19.3944
R18214 vdd.n2153 vdd.n1419 19.3944
R18215 vdd.n2166 vdd.n1419 19.3944
R18216 vdd.n2166 vdd.n1416 19.3944
R18217 vdd.n2172 vdd.n1416 19.3944
R18218 vdd.n2172 vdd.n1417 19.3944
R18219 vdd.n1417 vdd.n1406 19.3944
R18220 vdd.n1661 vdd.n1603 19.3944
R18221 vdd.n1661 vdd.n1660 19.3944
R18222 vdd.n1660 vdd.n1659 19.3944
R18223 vdd.n1659 vdd.n1609 19.3944
R18224 vdd.n1655 vdd.n1609 19.3944
R18225 vdd.n1655 vdd.n1654 19.3944
R18226 vdd.n1654 vdd.n1653 19.3944
R18227 vdd.n1653 vdd.n1615 19.3944
R18228 vdd.n1649 vdd.n1615 19.3944
R18229 vdd.n1649 vdd.n1648 19.3944
R18230 vdd.n1648 vdd.n1647 19.3944
R18231 vdd.n1647 vdd.n1621 19.3944
R18232 vdd.n1643 vdd.n1621 19.3944
R18233 vdd.n1643 vdd.n1642 19.3944
R18234 vdd.n1642 vdd.n1641 19.3944
R18235 vdd.n1641 vdd.n1627 19.3944
R18236 vdd.n1637 vdd.n1627 19.3944
R18237 vdd.n1637 vdd.n1636 19.3944
R18238 vdd.n1636 vdd.n1635 19.3944
R18239 vdd.n1635 vdd.n1633 19.3944
R18240 vdd.n1699 vdd.n1698 19.3944
R18241 vdd.n1698 vdd.n1574 19.3944
R18242 vdd.n1694 vdd.n1574 19.3944
R18243 vdd.n1694 vdd.n1693 19.3944
R18244 vdd.n1693 vdd.n1692 19.3944
R18245 vdd.n1692 vdd.n1580 19.3944
R18246 vdd.n1688 vdd.n1580 19.3944
R18247 vdd.n1688 vdd.n1687 19.3944
R18248 vdd.n1687 vdd.n1686 19.3944
R18249 vdd.n1686 vdd.n1586 19.3944
R18250 vdd.n1682 vdd.n1586 19.3944
R18251 vdd.n1682 vdd.n1681 19.3944
R18252 vdd.n1681 vdd.n1680 19.3944
R18253 vdd.n1680 vdd.n1592 19.3944
R18254 vdd.n1676 vdd.n1592 19.3944
R18255 vdd.n1676 vdd.n1675 19.3944
R18256 vdd.n1675 vdd.n1674 19.3944
R18257 vdd.n1674 vdd.n1598 19.3944
R18258 vdd.n1670 vdd.n1598 19.3944
R18259 vdd.n1670 vdd.n1669 19.3944
R18260 vdd.n1733 vdd.n1732 19.3944
R18261 vdd.n1732 vdd.n1547 19.3944
R18262 vdd.n1728 vdd.n1547 19.3944
R18263 vdd.n1728 vdd.n1727 19.3944
R18264 vdd.n1727 vdd.n1726 19.3944
R18265 vdd.n1726 vdd.n1552 19.3944
R18266 vdd.n1722 vdd.n1552 19.3944
R18267 vdd.n1722 vdd.n1721 19.3944
R18268 vdd.n1721 vdd.n1720 19.3944
R18269 vdd.n1720 vdd.n1558 19.3944
R18270 vdd.n1716 vdd.n1558 19.3944
R18271 vdd.n1716 vdd.n1715 19.3944
R18272 vdd.n1715 vdd.n1714 19.3944
R18273 vdd.n1714 vdd.n1564 19.3944
R18274 vdd.n1710 vdd.n1564 19.3944
R18275 vdd.n1710 vdd.n1709 19.3944
R18276 vdd.n1709 vdd.n1708 19.3944
R18277 vdd.n1708 vdd.n1570 19.3944
R18278 vdd.n2220 vdd.n1160 19.3944
R18279 vdd.n2220 vdd.n1166 19.3944
R18280 vdd.n2215 vdd.n1166 19.3944
R18281 vdd.n2215 vdd.n2214 19.3944
R18282 vdd.n2214 vdd.n2213 19.3944
R18283 vdd.n2213 vdd.n1173 19.3944
R18284 vdd.n2208 vdd.n1173 19.3944
R18285 vdd.n2208 vdd.n2207 19.3944
R18286 vdd.n2207 vdd.n2206 19.3944
R18287 vdd.n2206 vdd.n1180 19.3944
R18288 vdd.n2201 vdd.n1180 19.3944
R18289 vdd.n2201 vdd.n2200 19.3944
R18290 vdd.n2200 vdd.n2199 19.3944
R18291 vdd.n2199 vdd.n1187 19.3944
R18292 vdd.n2194 vdd.n1187 19.3944
R18293 vdd.n2194 vdd.n2193 19.3944
R18294 vdd.n1399 vdd.n1192 19.3944
R18295 vdd.n2189 vdd.n1396 19.3944
R18296 vdd.n2259 vdd.n1120 19.3944
R18297 vdd.n2259 vdd.n1126 19.3944
R18298 vdd.n2254 vdd.n1126 19.3944
R18299 vdd.n2254 vdd.n2253 19.3944
R18300 vdd.n2253 vdd.n2252 19.3944
R18301 vdd.n2252 vdd.n1133 19.3944
R18302 vdd.n2247 vdd.n1133 19.3944
R18303 vdd.n2247 vdd.n2246 19.3944
R18304 vdd.n2246 vdd.n2245 19.3944
R18305 vdd.n2245 vdd.n1140 19.3944
R18306 vdd.n2240 vdd.n1140 19.3944
R18307 vdd.n2240 vdd.n2239 19.3944
R18308 vdd.n2239 vdd.n2238 19.3944
R18309 vdd.n2238 vdd.n1147 19.3944
R18310 vdd.n2233 vdd.n1147 19.3944
R18311 vdd.n2233 vdd.n2232 19.3944
R18312 vdd.n2232 vdd.n2231 19.3944
R18313 vdd.n2231 vdd.n1154 19.3944
R18314 vdd.n2226 vdd.n1154 19.3944
R18315 vdd.n2226 vdd.n2225 19.3944
R18316 vdd.n2296 vdd.n1095 19.3944
R18317 vdd.n2296 vdd.n1096 19.3944
R18318 vdd.n2291 vdd.n2290 19.3944
R18319 vdd.n2286 vdd.n2285 19.3944
R18320 vdd.n2285 vdd.n2284 19.3944
R18321 vdd.n2284 vdd.n1100 19.3944
R18322 vdd.n2279 vdd.n1100 19.3944
R18323 vdd.n2279 vdd.n2278 19.3944
R18324 vdd.n2278 vdd.n2277 19.3944
R18325 vdd.n2277 vdd.n1107 19.3944
R18326 vdd.n2272 vdd.n1107 19.3944
R18327 vdd.n2272 vdd.n2271 19.3944
R18328 vdd.n2271 vdd.n2270 19.3944
R18329 vdd.n2270 vdd.n1114 19.3944
R18330 vdd.n2265 vdd.n1114 19.3944
R18331 vdd.n2265 vdd.n2264 19.3944
R18332 vdd.n1746 vdd.n1504 19.3944
R18333 vdd.n1746 vdd.n1502 19.3944
R18334 vdd.n1750 vdd.n1502 19.3944
R18335 vdd.n1750 vdd.n1492 19.3944
R18336 vdd.n1763 vdd.n1492 19.3944
R18337 vdd.n1763 vdd.n1490 19.3944
R18338 vdd.n1767 vdd.n1490 19.3944
R18339 vdd.n1767 vdd.n1481 19.3944
R18340 vdd.n1780 vdd.n1481 19.3944
R18341 vdd.n1780 vdd.n1479 19.3944
R18342 vdd.n1784 vdd.n1479 19.3944
R18343 vdd.n1784 vdd.n1470 19.3944
R18344 vdd.n1796 vdd.n1470 19.3944
R18345 vdd.n1796 vdd.n1468 19.3944
R18346 vdd.n1800 vdd.n1468 19.3944
R18347 vdd.n1800 vdd.n1458 19.3944
R18348 vdd.n1813 vdd.n1458 19.3944
R18349 vdd.n1813 vdd.n1456 19.3944
R18350 vdd.n2112 vdd.n1456 19.3944
R18351 vdd.n2112 vdd.n1447 19.3944
R18352 vdd.n2124 vdd.n1447 19.3944
R18353 vdd.n2124 vdd.n1445 19.3944
R18354 vdd.n2128 vdd.n1445 19.3944
R18355 vdd.n2128 vdd.n1435 19.3944
R18356 vdd.n2141 vdd.n1435 19.3944
R18357 vdd.n2141 vdd.n1433 19.3944
R18358 vdd.n2145 vdd.n1433 19.3944
R18359 vdd.n2145 vdd.n1424 19.3944
R18360 vdd.n2158 vdd.n1424 19.3944
R18361 vdd.n2158 vdd.n1422 19.3944
R18362 vdd.n2162 vdd.n1422 19.3944
R18363 vdd.n2162 vdd.n1412 19.3944
R18364 vdd.n2176 vdd.n1412 19.3944
R18365 vdd.n2176 vdd.n1410 19.3944
R18366 vdd.n2180 vdd.n1410 19.3944
R18367 vdd.n3239 vdd.n655 19.3944
R18368 vdd.n3243 vdd.n655 19.3944
R18369 vdd.n3243 vdd.n646 19.3944
R18370 vdd.n3255 vdd.n646 19.3944
R18371 vdd.n3255 vdd.n644 19.3944
R18372 vdd.n3259 vdd.n644 19.3944
R18373 vdd.n3259 vdd.n633 19.3944
R18374 vdd.n3271 vdd.n633 19.3944
R18375 vdd.n3271 vdd.n631 19.3944
R18376 vdd.n3275 vdd.n631 19.3944
R18377 vdd.n3275 vdd.n622 19.3944
R18378 vdd.n3288 vdd.n622 19.3944
R18379 vdd.n3288 vdd.n620 19.3944
R18380 vdd.n3295 vdd.n620 19.3944
R18381 vdd.n3295 vdd.n3294 19.3944
R18382 vdd.n3294 vdd.n610 19.3944
R18383 vdd.n3308 vdd.n610 19.3944
R18384 vdd.n3309 vdd.n3308 19.3944
R18385 vdd.n3310 vdd.n3309 19.3944
R18386 vdd.n3310 vdd.n608 19.3944
R18387 vdd.n3315 vdd.n608 19.3944
R18388 vdd.n3316 vdd.n3315 19.3944
R18389 vdd.n3317 vdd.n3316 19.3944
R18390 vdd.n3317 vdd.n606 19.3944
R18391 vdd.n3322 vdd.n606 19.3944
R18392 vdd.n3323 vdd.n3322 19.3944
R18393 vdd.n3324 vdd.n3323 19.3944
R18394 vdd.n3324 vdd.n604 19.3944
R18395 vdd.n3330 vdd.n604 19.3944
R18396 vdd.n3331 vdd.n3330 19.3944
R18397 vdd.n3332 vdd.n3331 19.3944
R18398 vdd.n3332 vdd.n602 19.3944
R18399 vdd.n3337 vdd.n602 19.3944
R18400 vdd.n3338 vdd.n3337 19.3944
R18401 vdd.n3339 vdd.n3338 19.3944
R18402 vdd.n550 vdd.n417 19.3944
R18403 vdd.n556 vdd.n417 19.3944
R18404 vdd.n557 vdd.n556 19.3944
R18405 vdd.n560 vdd.n557 19.3944
R18406 vdd.n560 vdd.n415 19.3944
R18407 vdd.n566 vdd.n415 19.3944
R18408 vdd.n567 vdd.n566 19.3944
R18409 vdd.n570 vdd.n567 19.3944
R18410 vdd.n570 vdd.n413 19.3944
R18411 vdd.n576 vdd.n413 19.3944
R18412 vdd.n577 vdd.n576 19.3944
R18413 vdd.n580 vdd.n577 19.3944
R18414 vdd.n580 vdd.n411 19.3944
R18415 vdd.n586 vdd.n411 19.3944
R18416 vdd.n587 vdd.n586 19.3944
R18417 vdd.n590 vdd.n587 19.3944
R18418 vdd.n590 vdd.n409 19.3944
R18419 vdd.n596 vdd.n409 19.3944
R18420 vdd.n598 vdd.n596 19.3944
R18421 vdd.n599 vdd.n598 19.3944
R18422 vdd.n497 vdd.n496 19.3944
R18423 vdd.n500 vdd.n497 19.3944
R18424 vdd.n500 vdd.n429 19.3944
R18425 vdd.n506 vdd.n429 19.3944
R18426 vdd.n507 vdd.n506 19.3944
R18427 vdd.n510 vdd.n507 19.3944
R18428 vdd.n510 vdd.n427 19.3944
R18429 vdd.n516 vdd.n427 19.3944
R18430 vdd.n517 vdd.n516 19.3944
R18431 vdd.n520 vdd.n517 19.3944
R18432 vdd.n520 vdd.n425 19.3944
R18433 vdd.n526 vdd.n425 19.3944
R18434 vdd.n527 vdd.n526 19.3944
R18435 vdd.n530 vdd.n527 19.3944
R18436 vdd.n530 vdd.n423 19.3944
R18437 vdd.n536 vdd.n423 19.3944
R18438 vdd.n537 vdd.n536 19.3944
R18439 vdd.n540 vdd.n537 19.3944
R18440 vdd.n540 vdd.n421 19.3944
R18441 vdd.n546 vdd.n421 19.3944
R18442 vdd.n447 vdd.n446 19.3944
R18443 vdd.n450 vdd.n447 19.3944
R18444 vdd.n450 vdd.n441 19.3944
R18445 vdd.n456 vdd.n441 19.3944
R18446 vdd.n457 vdd.n456 19.3944
R18447 vdd.n460 vdd.n457 19.3944
R18448 vdd.n460 vdd.n439 19.3944
R18449 vdd.n466 vdd.n439 19.3944
R18450 vdd.n467 vdd.n466 19.3944
R18451 vdd.n470 vdd.n467 19.3944
R18452 vdd.n470 vdd.n437 19.3944
R18453 vdd.n476 vdd.n437 19.3944
R18454 vdd.n477 vdd.n476 19.3944
R18455 vdd.n480 vdd.n477 19.3944
R18456 vdd.n480 vdd.n435 19.3944
R18457 vdd.n486 vdd.n435 19.3944
R18458 vdd.n487 vdd.n486 19.3944
R18459 vdd.n490 vdd.n487 19.3944
R18460 vdd.n3235 vdd.n652 19.3944
R18461 vdd.n3247 vdd.n652 19.3944
R18462 vdd.n3247 vdd.n650 19.3944
R18463 vdd.n3251 vdd.n650 19.3944
R18464 vdd.n3251 vdd.n640 19.3944
R18465 vdd.n3263 vdd.n640 19.3944
R18466 vdd.n3263 vdd.n638 19.3944
R18467 vdd.n3267 vdd.n638 19.3944
R18468 vdd.n3267 vdd.n628 19.3944
R18469 vdd.n3280 vdd.n628 19.3944
R18470 vdd.n3280 vdd.n626 19.3944
R18471 vdd.n3284 vdd.n626 19.3944
R18472 vdd.n3284 vdd.n617 19.3944
R18473 vdd.n3299 vdd.n617 19.3944
R18474 vdd.n3299 vdd.n615 19.3944
R18475 vdd.n3303 vdd.n615 19.3944
R18476 vdd.n3303 vdd.n324 19.3944
R18477 vdd.n3381 vdd.n324 19.3944
R18478 vdd.n3381 vdd.n325 19.3944
R18479 vdd.n3375 vdd.n325 19.3944
R18480 vdd.n3375 vdd.n3374 19.3944
R18481 vdd.n3374 vdd.n3373 19.3944
R18482 vdd.n3373 vdd.n337 19.3944
R18483 vdd.n3367 vdd.n337 19.3944
R18484 vdd.n3367 vdd.n3366 19.3944
R18485 vdd.n3366 vdd.n3365 19.3944
R18486 vdd.n3365 vdd.n347 19.3944
R18487 vdd.n3359 vdd.n347 19.3944
R18488 vdd.n3359 vdd.n3358 19.3944
R18489 vdd.n3358 vdd.n3357 19.3944
R18490 vdd.n3357 vdd.n358 19.3944
R18491 vdd.n3351 vdd.n358 19.3944
R18492 vdd.n3351 vdd.n3350 19.3944
R18493 vdd.n3350 vdd.n3349 19.3944
R18494 vdd.n3349 vdd.n369 19.3944
R18495 vdd.n3192 vdd.n3191 19.3944
R18496 vdd.n3191 vdd.n3190 19.3944
R18497 vdd.n3190 vdd.n694 19.3944
R18498 vdd.n3184 vdd.n694 19.3944
R18499 vdd.n3184 vdd.n3183 19.3944
R18500 vdd.n3183 vdd.n3182 19.3944
R18501 vdd.n3182 vdd.n700 19.3944
R18502 vdd.n3176 vdd.n700 19.3944
R18503 vdd.n3176 vdd.n3175 19.3944
R18504 vdd.n3175 vdd.n3174 19.3944
R18505 vdd.n3174 vdd.n706 19.3944
R18506 vdd.n3168 vdd.n706 19.3944
R18507 vdd.n3168 vdd.n3167 19.3944
R18508 vdd.n3167 vdd.n3166 19.3944
R18509 vdd.n3166 vdd.n712 19.3944
R18510 vdd.n3160 vdd.n712 19.3944
R18511 vdd.n3160 vdd.n3159 19.3944
R18512 vdd.n3159 vdd.n3158 19.3944
R18513 vdd.n3158 vdd.n718 19.3944
R18514 vdd.n3152 vdd.n718 19.3944
R18515 vdd.n3232 vdd.n3231 19.3944
R18516 vdd.n3231 vdd.n662 19.3944
R18517 vdd.n3226 vdd.n3225 19.3944
R18518 vdd.n3222 vdd.n3221 19.3944
R18519 vdd.n3221 vdd.n668 19.3944
R18520 vdd.n3216 vdd.n668 19.3944
R18521 vdd.n3216 vdd.n3215 19.3944
R18522 vdd.n3215 vdd.n3214 19.3944
R18523 vdd.n3214 vdd.n674 19.3944
R18524 vdd.n3208 vdd.n674 19.3944
R18525 vdd.n3208 vdd.n3207 19.3944
R18526 vdd.n3207 vdd.n3206 19.3944
R18527 vdd.n3206 vdd.n680 19.3944
R18528 vdd.n3200 vdd.n680 19.3944
R18529 vdd.n3200 vdd.n3199 19.3944
R18530 vdd.n3199 vdd.n3198 19.3944
R18531 vdd.n3147 vdd.n722 19.3944
R18532 vdd.n3147 vdd.n726 19.3944
R18533 vdd.n3142 vdd.n726 19.3944
R18534 vdd.n3142 vdd.n3141 19.3944
R18535 vdd.n3141 vdd.n732 19.3944
R18536 vdd.n3136 vdd.n732 19.3944
R18537 vdd.n3136 vdd.n3135 19.3944
R18538 vdd.n3135 vdd.n3134 19.3944
R18539 vdd.n3134 vdd.n738 19.3944
R18540 vdd.n3128 vdd.n738 19.3944
R18541 vdd.n3128 vdd.n3127 19.3944
R18542 vdd.n3127 vdd.n3126 19.3944
R18543 vdd.n3126 vdd.n744 19.3944
R18544 vdd.n3120 vdd.n744 19.3944
R18545 vdd.n3120 vdd.n3119 19.3944
R18546 vdd.n3119 vdd.n3118 19.3944
R18547 vdd.n3114 vdd.n3113 19.3944
R18548 vdd.n3110 vdd.n3109 19.3944
R18549 vdd.n1668 vdd.n1603 19.0066
R18550 vdd.n2224 vdd.n1160 19.0066
R18551 vdd.n550 vdd.n547 19.0066
R18552 vdd.n3151 vdd.n722 19.0066
R18553 vdd.n1736 vdd.n1506 18.5924
R18554 vdd.n2182 vdd.n1054 18.5924
R18555 vdd.n3237 vdd.n658 18.5924
R18556 vdd.n3346 vdd.n3345 18.5924
R18557 vdd.n1225 vdd.n1224 16.0975
R18558 vdd.n953 vdd.n952 16.0975
R18559 vdd.n1511 vdd.n1510 16.0975
R18560 vdd.n1667 vdd.n1666 16.0975
R18561 vdd.n1703 vdd.n1702 16.0975
R18562 vdd.n2187 vdd.n2186 16.0975
R18563 vdd.n1162 vdd.n1161 16.0975
R18564 vdd.n1122 vdd.n1121 16.0975
R18565 vdd.n1245 vdd.n1244 16.0975
R18566 vdd.n944 vdd.n943 16.0975
R18567 vdd.n2622 vdd.n2621 16.0975
R18568 vdd.n406 vdd.n405 16.0975
R18569 vdd.n420 vdd.n419 16.0975
R18570 vdd.n432 vdd.n431 16.0975
R18571 vdd.n724 vdd.n723 16.0975
R18572 vdd.n687 vdd.n686 16.0975
R18573 vdd.n805 vdd.n804 16.0975
R18574 vdd.n2619 vdd.n2618 16.0975
R18575 vdd.n3106 vdd.n3105 16.0975
R18576 vdd.n769 vdd.n768 16.0975
R18577 vdd.t258 vdd.n2582 15.4182
R18578 vdd.n2855 vdd.t101 15.4182
R18579 vdd.n28 vdd.n27 15.0023
R18580 vdd.n2334 vdd.n1047 14.0578
R18581 vdd.n3068 vdd.n756 14.0578
R18582 vdd.n316 vdd.n281 13.1884
R18583 vdd.n261 vdd.n226 13.1884
R18584 vdd.n218 vdd.n183 13.1884
R18585 vdd.n163 vdd.n128 13.1884
R18586 vdd.n121 vdd.n86 13.1884
R18587 vdd.n66 vdd.n31 13.1884
R18588 vdd.n2047 vdd.n2012 13.1884
R18589 vdd.n2102 vdd.n2067 13.1884
R18590 vdd.n1949 vdd.n1914 13.1884
R18591 vdd.n2004 vdd.n1969 13.1884
R18592 vdd.n1852 vdd.n1817 13.1884
R18593 vdd.n1907 vdd.n1872 13.1884
R18594 vdd.n1704 vdd.n1699 12.9944
R18595 vdd.n1704 vdd.n1570 12.9944
R18596 vdd.n2263 vdd.n1120 12.9944
R18597 vdd.n2264 vdd.n2263 12.9944
R18598 vdd.n496 vdd.n433 12.9944
R18599 vdd.n490 vdd.n433 12.9944
R18600 vdd.n3192 vdd.n688 12.9944
R18601 vdd.n3198 vdd.n688 12.9944
R18602 vdd.n317 vdd.n279 12.8005
R18603 vdd.n312 vdd.n283 12.8005
R18604 vdd.n262 vdd.n224 12.8005
R18605 vdd.n257 vdd.n228 12.8005
R18606 vdd.n219 vdd.n181 12.8005
R18607 vdd.n214 vdd.n185 12.8005
R18608 vdd.n164 vdd.n126 12.8005
R18609 vdd.n159 vdd.n130 12.8005
R18610 vdd.n122 vdd.n84 12.8005
R18611 vdd.n117 vdd.n88 12.8005
R18612 vdd.n67 vdd.n29 12.8005
R18613 vdd.n62 vdd.n33 12.8005
R18614 vdd.n2048 vdd.n2010 12.8005
R18615 vdd.n2043 vdd.n2014 12.8005
R18616 vdd.n2103 vdd.n2065 12.8005
R18617 vdd.n2098 vdd.n2069 12.8005
R18618 vdd.n1950 vdd.n1912 12.8005
R18619 vdd.n1945 vdd.n1916 12.8005
R18620 vdd.n2005 vdd.n1967 12.8005
R18621 vdd.n2000 vdd.n1971 12.8005
R18622 vdd.n1853 vdd.n1815 12.8005
R18623 vdd.n1848 vdd.n1819 12.8005
R18624 vdd.n1908 vdd.n1870 12.8005
R18625 vdd.n1903 vdd.n1874 12.8005
R18626 vdd.n311 vdd.n284 12.0247
R18627 vdd.n256 vdd.n229 12.0247
R18628 vdd.n213 vdd.n186 12.0247
R18629 vdd.n158 vdd.n131 12.0247
R18630 vdd.n116 vdd.n89 12.0247
R18631 vdd.n61 vdd.n34 12.0247
R18632 vdd.n2042 vdd.n2015 12.0247
R18633 vdd.n2097 vdd.n2070 12.0247
R18634 vdd.n1944 vdd.n1917 12.0247
R18635 vdd.n1999 vdd.n1972 12.0247
R18636 vdd.n1847 vdd.n1820 12.0247
R18637 vdd.n1902 vdd.n1875 12.0247
R18638 vdd.n1744 vdd.n1506 11.337
R18639 vdd.n1752 vdd.n1500 11.337
R18640 vdd.n1752 vdd.n1494 11.337
R18641 vdd.n1761 vdd.n1494 11.337
R18642 vdd.n1769 vdd.n1488 11.337
R18643 vdd.n1778 vdd.n1777 11.337
R18644 vdd.n1794 vdd.n1472 11.337
R18645 vdd.n1802 vdd.n1465 11.337
R18646 vdd.n1811 vdd.n1810 11.337
R18647 vdd.n2114 vdd.n1454 11.337
R18648 vdd.n2130 vdd.n1443 11.337
R18649 vdd.n2139 vdd.n1437 11.337
R18650 vdd.n2147 vdd.n1431 11.337
R18651 vdd.n2156 vdd.n2155 11.337
R18652 vdd.n2164 vdd.n1414 11.337
R18653 vdd.n2174 vdd.n1414 11.337
R18654 vdd.n2182 vdd.n1407 11.337
R18655 vdd.n3237 vdd.n659 11.337
R18656 vdd.n3245 vdd.n648 11.337
R18657 vdd.n3253 vdd.n648 11.337
R18658 vdd.n3261 vdd.n642 11.337
R18659 vdd.n3269 vdd.n635 11.337
R18660 vdd.n3278 vdd.n3277 11.337
R18661 vdd.n3286 vdd.n624 11.337
R18662 vdd.n3305 vdd.n613 11.337
R18663 vdd.n3379 vdd.n328 11.337
R18664 vdd.n3377 vdd.n332 11.337
R18665 vdd.n3371 vdd.n3370 11.337
R18666 vdd.n3363 vdd.n349 11.337
R18667 vdd.n3362 vdd.n3361 11.337
R18668 vdd.n3355 vdd.n3354 11.337
R18669 vdd.n3354 vdd.n3353 11.337
R18670 vdd.n3353 vdd.n363 11.337
R18671 vdd.n3347 vdd.n3346 11.337
R18672 vdd.n308 vdd.n307 11.249
R18673 vdd.n253 vdd.n252 11.249
R18674 vdd.n210 vdd.n209 11.249
R18675 vdd.n155 vdd.n154 11.249
R18676 vdd.n113 vdd.n112 11.249
R18677 vdd.n58 vdd.n57 11.249
R18678 vdd.n2039 vdd.n2038 11.249
R18679 vdd.n2094 vdd.n2093 11.249
R18680 vdd.n1941 vdd.n1940 11.249
R18681 vdd.n1996 vdd.n1995 11.249
R18682 vdd.n1844 vdd.n1843 11.249
R18683 vdd.n1899 vdd.n1898 11.249
R18684 vdd.n2164 vdd.t154 10.7702
R18685 vdd.n3253 vdd.t152 10.7702
R18686 vdd.n293 vdd.n292 10.7238
R18687 vdd.n238 vdd.n237 10.7238
R18688 vdd.n195 vdd.n194 10.7238
R18689 vdd.n140 vdd.n139 10.7238
R18690 vdd.n98 vdd.n97 10.7238
R18691 vdd.n43 vdd.n42 10.7238
R18692 vdd.n2024 vdd.n2023 10.7238
R18693 vdd.n2079 vdd.n2078 10.7238
R18694 vdd.n1926 vdd.n1925 10.7238
R18695 vdd.n1981 vdd.n1980 10.7238
R18696 vdd.n1829 vdd.n1828 10.7238
R18697 vdd.n1884 vdd.n1883 10.7238
R18698 vdd.n2510 vdd.t245 10.6568
R18699 vdd.t247 vdd.n899 10.6568
R18700 vdd.n2343 vdd.n1045 10.6151
R18701 vdd.n2344 vdd.n2343 10.6151
R18702 vdd.n2345 vdd.n2344 10.6151
R18703 vdd.n2345 vdd.n1034 10.6151
R18704 vdd.n2355 vdd.n1034 10.6151
R18705 vdd.n2356 vdd.n2355 10.6151
R18706 vdd.n2357 vdd.n2356 10.6151
R18707 vdd.n2357 vdd.n1021 10.6151
R18708 vdd.n2367 vdd.n1021 10.6151
R18709 vdd.n2368 vdd.n2367 10.6151
R18710 vdd.n2369 vdd.n2368 10.6151
R18711 vdd.n2369 vdd.n1009 10.6151
R18712 vdd.n2380 vdd.n1009 10.6151
R18713 vdd.n2381 vdd.n2380 10.6151
R18714 vdd.n2382 vdd.n2381 10.6151
R18715 vdd.n2382 vdd.n997 10.6151
R18716 vdd.n2392 vdd.n997 10.6151
R18717 vdd.n2393 vdd.n2392 10.6151
R18718 vdd.n2394 vdd.n2393 10.6151
R18719 vdd.n2394 vdd.n985 10.6151
R18720 vdd.n2404 vdd.n985 10.6151
R18721 vdd.n2405 vdd.n2404 10.6151
R18722 vdd.n2406 vdd.n2405 10.6151
R18723 vdd.n2406 vdd.n974 10.6151
R18724 vdd.n2416 vdd.n974 10.6151
R18725 vdd.n2417 vdd.n2416 10.6151
R18726 vdd.n2418 vdd.n2417 10.6151
R18727 vdd.n2418 vdd.n961 10.6151
R18728 vdd.n2430 vdd.n961 10.6151
R18729 vdd.n2431 vdd.n2430 10.6151
R18730 vdd.n2433 vdd.n2431 10.6151
R18731 vdd.n2433 vdd.n2432 10.6151
R18732 vdd.n2432 vdd.n942 10.6151
R18733 vdd.n2580 vdd.n2579 10.6151
R18734 vdd.n2579 vdd.n2578 10.6151
R18735 vdd.n2578 vdd.n2575 10.6151
R18736 vdd.n2575 vdd.n2574 10.6151
R18737 vdd.n2574 vdd.n2571 10.6151
R18738 vdd.n2571 vdd.n2570 10.6151
R18739 vdd.n2570 vdd.n2567 10.6151
R18740 vdd.n2567 vdd.n2566 10.6151
R18741 vdd.n2566 vdd.n2563 10.6151
R18742 vdd.n2563 vdd.n2562 10.6151
R18743 vdd.n2562 vdd.n2559 10.6151
R18744 vdd.n2559 vdd.n2558 10.6151
R18745 vdd.n2558 vdd.n2555 10.6151
R18746 vdd.n2555 vdd.n2554 10.6151
R18747 vdd.n2554 vdd.n2551 10.6151
R18748 vdd.n2551 vdd.n2550 10.6151
R18749 vdd.n2550 vdd.n2547 10.6151
R18750 vdd.n2547 vdd.n2546 10.6151
R18751 vdd.n2546 vdd.n2543 10.6151
R18752 vdd.n2543 vdd.n2542 10.6151
R18753 vdd.n2542 vdd.n2539 10.6151
R18754 vdd.n2539 vdd.n2538 10.6151
R18755 vdd.n2538 vdd.n2535 10.6151
R18756 vdd.n2535 vdd.n2534 10.6151
R18757 vdd.n2534 vdd.n2531 10.6151
R18758 vdd.n2531 vdd.n2530 10.6151
R18759 vdd.n2530 vdd.n2527 10.6151
R18760 vdd.n2527 vdd.n2526 10.6151
R18761 vdd.n2526 vdd.n2523 10.6151
R18762 vdd.n2523 vdd.n2522 10.6151
R18763 vdd.n2522 vdd.n2519 10.6151
R18764 vdd.n2517 vdd.n2514 10.6151
R18765 vdd.n2514 vdd.n2513 10.6151
R18766 vdd.n1282 vdd.n1281 10.6151
R18767 vdd.n1284 vdd.n1282 10.6151
R18768 vdd.n1285 vdd.n1284 10.6151
R18769 vdd.n1287 vdd.n1285 10.6151
R18770 vdd.n1288 vdd.n1287 10.6151
R18771 vdd.n1290 vdd.n1288 10.6151
R18772 vdd.n1291 vdd.n1290 10.6151
R18773 vdd.n1293 vdd.n1291 10.6151
R18774 vdd.n1294 vdd.n1293 10.6151
R18775 vdd.n1296 vdd.n1294 10.6151
R18776 vdd.n1297 vdd.n1296 10.6151
R18777 vdd.n1299 vdd.n1297 10.6151
R18778 vdd.n1300 vdd.n1299 10.6151
R18779 vdd.n1302 vdd.n1300 10.6151
R18780 vdd.n1303 vdd.n1302 10.6151
R18781 vdd.n1305 vdd.n1303 10.6151
R18782 vdd.n1306 vdd.n1305 10.6151
R18783 vdd.n1328 vdd.n1306 10.6151
R18784 vdd.n1328 vdd.n1327 10.6151
R18785 vdd.n1327 vdd.n1326 10.6151
R18786 vdd.n1326 vdd.n1324 10.6151
R18787 vdd.n1324 vdd.n1323 10.6151
R18788 vdd.n1323 vdd.n1321 10.6151
R18789 vdd.n1321 vdd.n1320 10.6151
R18790 vdd.n1320 vdd.n1318 10.6151
R18791 vdd.n1318 vdd.n1317 10.6151
R18792 vdd.n1317 vdd.n1315 10.6151
R18793 vdd.n1315 vdd.n1314 10.6151
R18794 vdd.n1314 vdd.n1312 10.6151
R18795 vdd.n1312 vdd.n1311 10.6151
R18796 vdd.n1311 vdd.n1308 10.6151
R18797 vdd.n1308 vdd.n1307 10.6151
R18798 vdd.n1307 vdd.n945 10.6151
R18799 vdd.n2331 vdd.n2330 10.6151
R18800 vdd.n2330 vdd.n2329 10.6151
R18801 vdd.n2329 vdd.n2328 10.6151
R18802 vdd.n2328 vdd.n2326 10.6151
R18803 vdd.n2326 vdd.n2323 10.6151
R18804 vdd.n2323 vdd.n2322 10.6151
R18805 vdd.n2322 vdd.n2319 10.6151
R18806 vdd.n2319 vdd.n2318 10.6151
R18807 vdd.n2318 vdd.n2315 10.6151
R18808 vdd.n2315 vdd.n2314 10.6151
R18809 vdd.n2314 vdd.n2311 10.6151
R18810 vdd.n2311 vdd.n2310 10.6151
R18811 vdd.n2310 vdd.n2307 10.6151
R18812 vdd.n2307 vdd.n2306 10.6151
R18813 vdd.n2306 vdd.n2303 10.6151
R18814 vdd.n2303 vdd.n2302 10.6151
R18815 vdd.n2302 vdd.n2299 10.6151
R18816 vdd.n2299 vdd.n1090 10.6151
R18817 vdd.n1248 vdd.n1090 10.6151
R18818 vdd.n1249 vdd.n1248 10.6151
R18819 vdd.n1252 vdd.n1249 10.6151
R18820 vdd.n1253 vdd.n1252 10.6151
R18821 vdd.n1256 vdd.n1253 10.6151
R18822 vdd.n1257 vdd.n1256 10.6151
R18823 vdd.n1260 vdd.n1257 10.6151
R18824 vdd.n1261 vdd.n1260 10.6151
R18825 vdd.n1264 vdd.n1261 10.6151
R18826 vdd.n1265 vdd.n1264 10.6151
R18827 vdd.n1268 vdd.n1265 10.6151
R18828 vdd.n1269 vdd.n1268 10.6151
R18829 vdd.n1272 vdd.n1269 10.6151
R18830 vdd.n1277 vdd.n1274 10.6151
R18831 vdd.n1278 vdd.n1277 10.6151
R18832 vdd.n2783 vdd.n2782 10.6151
R18833 vdd.n2782 vdd.n2781 10.6151
R18834 vdd.n2781 vdd.n2620 10.6151
R18835 vdd.n2725 vdd.n2620 10.6151
R18836 vdd.n2726 vdd.n2725 10.6151
R18837 vdd.n2728 vdd.n2726 10.6151
R18838 vdd.n2729 vdd.n2728 10.6151
R18839 vdd.n2731 vdd.n2729 10.6151
R18840 vdd.n2732 vdd.n2731 10.6151
R18841 vdd.n2762 vdd.n2732 10.6151
R18842 vdd.n2762 vdd.n2761 10.6151
R18843 vdd.n2761 vdd.n2760 10.6151
R18844 vdd.n2760 vdd.n2758 10.6151
R18845 vdd.n2758 vdd.n2757 10.6151
R18846 vdd.n2757 vdd.n2755 10.6151
R18847 vdd.n2755 vdd.n2754 10.6151
R18848 vdd.n2754 vdd.n2752 10.6151
R18849 vdd.n2752 vdd.n2751 10.6151
R18850 vdd.n2751 vdd.n2749 10.6151
R18851 vdd.n2749 vdd.n2748 10.6151
R18852 vdd.n2748 vdd.n2746 10.6151
R18853 vdd.n2746 vdd.n2745 10.6151
R18854 vdd.n2745 vdd.n2743 10.6151
R18855 vdd.n2743 vdd.n2742 10.6151
R18856 vdd.n2742 vdd.n2740 10.6151
R18857 vdd.n2740 vdd.n2739 10.6151
R18858 vdd.n2739 vdd.n2737 10.6151
R18859 vdd.n2737 vdd.n2736 10.6151
R18860 vdd.n2736 vdd.n2734 10.6151
R18861 vdd.n2734 vdd.n2733 10.6151
R18862 vdd.n2733 vdd.n807 10.6151
R18863 vdd.n3001 vdd.n807 10.6151
R18864 vdd.n3002 vdd.n3001 10.6151
R18865 vdd.n2852 vdd.n2851 10.6151
R18866 vdd.n2851 vdd.n2850 10.6151
R18867 vdd.n2850 vdd.n2849 10.6151
R18868 vdd.n2849 vdd.n2847 10.6151
R18869 vdd.n2847 vdd.n2844 10.6151
R18870 vdd.n2844 vdd.n2843 10.6151
R18871 vdd.n2843 vdd.n2840 10.6151
R18872 vdd.n2840 vdd.n2839 10.6151
R18873 vdd.n2839 vdd.n2836 10.6151
R18874 vdd.n2836 vdd.n2835 10.6151
R18875 vdd.n2835 vdd.n2832 10.6151
R18876 vdd.n2832 vdd.n2831 10.6151
R18877 vdd.n2831 vdd.n2828 10.6151
R18878 vdd.n2828 vdd.n2827 10.6151
R18879 vdd.n2827 vdd.n2824 10.6151
R18880 vdd.n2824 vdd.n2823 10.6151
R18881 vdd.n2823 vdd.n2820 10.6151
R18882 vdd.n2820 vdd.n2819 10.6151
R18883 vdd.n2819 vdd.n2816 10.6151
R18884 vdd.n2816 vdd.n2815 10.6151
R18885 vdd.n2815 vdd.n2812 10.6151
R18886 vdd.n2812 vdd.n2811 10.6151
R18887 vdd.n2811 vdd.n2808 10.6151
R18888 vdd.n2808 vdd.n2807 10.6151
R18889 vdd.n2807 vdd.n2804 10.6151
R18890 vdd.n2804 vdd.n2803 10.6151
R18891 vdd.n2803 vdd.n2800 10.6151
R18892 vdd.n2800 vdd.n2799 10.6151
R18893 vdd.n2799 vdd.n2796 10.6151
R18894 vdd.n2796 vdd.n2795 10.6151
R18895 vdd.n2795 vdd.n2792 10.6151
R18896 vdd.n2790 vdd.n2787 10.6151
R18897 vdd.n2787 vdd.n2786 10.6151
R18898 vdd.n2864 vdd.n897 10.6151
R18899 vdd.n2865 vdd.n2864 10.6151
R18900 vdd.n2866 vdd.n2865 10.6151
R18901 vdd.n2866 vdd.n886 10.6151
R18902 vdd.n2876 vdd.n886 10.6151
R18903 vdd.n2877 vdd.n2876 10.6151
R18904 vdd.n2878 vdd.n2877 10.6151
R18905 vdd.n2878 vdd.n874 10.6151
R18906 vdd.n2888 vdd.n874 10.6151
R18907 vdd.n2889 vdd.n2888 10.6151
R18908 vdd.n2890 vdd.n2889 10.6151
R18909 vdd.n2890 vdd.n862 10.6151
R18910 vdd.n2900 vdd.n862 10.6151
R18911 vdd.n2901 vdd.n2900 10.6151
R18912 vdd.n2902 vdd.n2901 10.6151
R18913 vdd.n2902 vdd.n851 10.6151
R18914 vdd.n2912 vdd.n851 10.6151
R18915 vdd.n2913 vdd.n2912 10.6151
R18916 vdd.n2914 vdd.n2913 10.6151
R18917 vdd.n2914 vdd.n837 10.6151
R18918 vdd.n2925 vdd.n837 10.6151
R18919 vdd.n2926 vdd.n2925 10.6151
R18920 vdd.n2927 vdd.n2926 10.6151
R18921 vdd.n2927 vdd.n826 10.6151
R18922 vdd.n2937 vdd.n826 10.6151
R18923 vdd.n2938 vdd.n2937 10.6151
R18924 vdd.n2939 vdd.n2938 10.6151
R18925 vdd.n2939 vdd.n812 10.6151
R18926 vdd.n2994 vdd.n812 10.6151
R18927 vdd.n2995 vdd.n2994 10.6151
R18928 vdd.n2996 vdd.n2995 10.6151
R18929 vdd.n2996 vdd.n779 10.6151
R18930 vdd.n3066 vdd.n779 10.6151
R18931 vdd.n3065 vdd.n3064 10.6151
R18932 vdd.n3064 vdd.n780 10.6151
R18933 vdd.n781 vdd.n780 10.6151
R18934 vdd.n3057 vdd.n781 10.6151
R18935 vdd.n3057 vdd.n3056 10.6151
R18936 vdd.n3056 vdd.n3055 10.6151
R18937 vdd.n3055 vdd.n783 10.6151
R18938 vdd.n3050 vdd.n783 10.6151
R18939 vdd.n3050 vdd.n3049 10.6151
R18940 vdd.n3049 vdd.n3048 10.6151
R18941 vdd.n3048 vdd.n786 10.6151
R18942 vdd.n3043 vdd.n786 10.6151
R18943 vdd.n3043 vdd.n3042 10.6151
R18944 vdd.n3042 vdd.n3041 10.6151
R18945 vdd.n3041 vdd.n789 10.6151
R18946 vdd.n3036 vdd.n789 10.6151
R18947 vdd.n3036 vdd.n3035 10.6151
R18948 vdd.n3035 vdd.n3033 10.6151
R18949 vdd.n3033 vdd.n792 10.6151
R18950 vdd.n3028 vdd.n792 10.6151
R18951 vdd.n3028 vdd.n3027 10.6151
R18952 vdd.n3027 vdd.n3026 10.6151
R18953 vdd.n3026 vdd.n795 10.6151
R18954 vdd.n3021 vdd.n795 10.6151
R18955 vdd.n3021 vdd.n3020 10.6151
R18956 vdd.n3020 vdd.n3019 10.6151
R18957 vdd.n3019 vdd.n798 10.6151
R18958 vdd.n3014 vdd.n798 10.6151
R18959 vdd.n3014 vdd.n3013 10.6151
R18960 vdd.n3013 vdd.n3012 10.6151
R18961 vdd.n3012 vdd.n801 10.6151
R18962 vdd.n3007 vdd.n3006 10.6151
R18963 vdd.n3006 vdd.n3005 10.6151
R18964 vdd.n2984 vdd.n2945 10.6151
R18965 vdd.n2979 vdd.n2945 10.6151
R18966 vdd.n2979 vdd.n2978 10.6151
R18967 vdd.n2978 vdd.n2977 10.6151
R18968 vdd.n2977 vdd.n2947 10.6151
R18969 vdd.n2972 vdd.n2947 10.6151
R18970 vdd.n2972 vdd.n2971 10.6151
R18971 vdd.n2971 vdd.n2970 10.6151
R18972 vdd.n2970 vdd.n2950 10.6151
R18973 vdd.n2965 vdd.n2950 10.6151
R18974 vdd.n2965 vdd.n2964 10.6151
R18975 vdd.n2964 vdd.n2963 10.6151
R18976 vdd.n2963 vdd.n2953 10.6151
R18977 vdd.n2958 vdd.n2953 10.6151
R18978 vdd.n2958 vdd.n2957 10.6151
R18979 vdd.n2957 vdd.n753 10.6151
R18980 vdd.n3101 vdd.n753 10.6151
R18981 vdd.n3101 vdd.n754 10.6151
R18982 vdd.n757 vdd.n754 10.6151
R18983 vdd.n3094 vdd.n757 10.6151
R18984 vdd.n3094 vdd.n3093 10.6151
R18985 vdd.n3093 vdd.n3092 10.6151
R18986 vdd.n3092 vdd.n759 10.6151
R18987 vdd.n3087 vdd.n759 10.6151
R18988 vdd.n3087 vdd.n3086 10.6151
R18989 vdd.n3086 vdd.n3085 10.6151
R18990 vdd.n3085 vdd.n762 10.6151
R18991 vdd.n3080 vdd.n762 10.6151
R18992 vdd.n3080 vdd.n3079 10.6151
R18993 vdd.n3079 vdd.n3078 10.6151
R18994 vdd.n3078 vdd.n765 10.6151
R18995 vdd.n3073 vdd.n3072 10.6151
R18996 vdd.n3072 vdd.n3071 10.6151
R18997 vdd.n2691 vdd.n2690 10.6151
R18998 vdd.n2777 vdd.n2691 10.6151
R18999 vdd.n2777 vdd.n2776 10.6151
R19000 vdd.n2776 vdd.n2775 10.6151
R19001 vdd.n2775 vdd.n2773 10.6151
R19002 vdd.n2773 vdd.n2772 10.6151
R19003 vdd.n2772 vdd.n2770 10.6151
R19004 vdd.n2770 vdd.n2769 10.6151
R19005 vdd.n2769 vdd.n2767 10.6151
R19006 vdd.n2767 vdd.n2766 10.6151
R19007 vdd.n2766 vdd.n2723 10.6151
R19008 vdd.n2723 vdd.n2722 10.6151
R19009 vdd.n2722 vdd.n2720 10.6151
R19010 vdd.n2720 vdd.n2719 10.6151
R19011 vdd.n2719 vdd.n2717 10.6151
R19012 vdd.n2717 vdd.n2716 10.6151
R19013 vdd.n2716 vdd.n2714 10.6151
R19014 vdd.n2714 vdd.n2713 10.6151
R19015 vdd.n2713 vdd.n2711 10.6151
R19016 vdd.n2711 vdd.n2710 10.6151
R19017 vdd.n2710 vdd.n2708 10.6151
R19018 vdd.n2708 vdd.n2707 10.6151
R19019 vdd.n2707 vdd.n2705 10.6151
R19020 vdd.n2705 vdd.n2704 10.6151
R19021 vdd.n2704 vdd.n2702 10.6151
R19022 vdd.n2702 vdd.n2701 10.6151
R19023 vdd.n2701 vdd.n2699 10.6151
R19024 vdd.n2699 vdd.n2698 10.6151
R19025 vdd.n2698 vdd.n2696 10.6151
R19026 vdd.n2696 vdd.n2695 10.6151
R19027 vdd.n2695 vdd.n2693 10.6151
R19028 vdd.n2693 vdd.n2692 10.6151
R19029 vdd.n2692 vdd.n771 10.6151
R19030 vdd.n2858 vdd.n903 10.6151
R19031 vdd.n2625 vdd.n903 10.6151
R19032 vdd.n2626 vdd.n2625 10.6151
R19033 vdd.n2629 vdd.n2626 10.6151
R19034 vdd.n2630 vdd.n2629 10.6151
R19035 vdd.n2633 vdd.n2630 10.6151
R19036 vdd.n2634 vdd.n2633 10.6151
R19037 vdd.n2637 vdd.n2634 10.6151
R19038 vdd.n2638 vdd.n2637 10.6151
R19039 vdd.n2641 vdd.n2638 10.6151
R19040 vdd.n2642 vdd.n2641 10.6151
R19041 vdd.n2645 vdd.n2642 10.6151
R19042 vdd.n2646 vdd.n2645 10.6151
R19043 vdd.n2649 vdd.n2646 10.6151
R19044 vdd.n2650 vdd.n2649 10.6151
R19045 vdd.n2653 vdd.n2650 10.6151
R19046 vdd.n2654 vdd.n2653 10.6151
R19047 vdd.n2657 vdd.n2654 10.6151
R19048 vdd.n2658 vdd.n2657 10.6151
R19049 vdd.n2661 vdd.n2658 10.6151
R19050 vdd.n2662 vdd.n2661 10.6151
R19051 vdd.n2665 vdd.n2662 10.6151
R19052 vdd.n2666 vdd.n2665 10.6151
R19053 vdd.n2669 vdd.n2666 10.6151
R19054 vdd.n2670 vdd.n2669 10.6151
R19055 vdd.n2673 vdd.n2670 10.6151
R19056 vdd.n2674 vdd.n2673 10.6151
R19057 vdd.n2677 vdd.n2674 10.6151
R19058 vdd.n2678 vdd.n2677 10.6151
R19059 vdd.n2681 vdd.n2678 10.6151
R19060 vdd.n2682 vdd.n2681 10.6151
R19061 vdd.n2687 vdd.n2685 10.6151
R19062 vdd.n2688 vdd.n2687 10.6151
R19063 vdd.n2860 vdd.n2859 10.6151
R19064 vdd.n2860 vdd.n892 10.6151
R19065 vdd.n2870 vdd.n892 10.6151
R19066 vdd.n2871 vdd.n2870 10.6151
R19067 vdd.n2872 vdd.n2871 10.6151
R19068 vdd.n2872 vdd.n880 10.6151
R19069 vdd.n2882 vdd.n880 10.6151
R19070 vdd.n2883 vdd.n2882 10.6151
R19071 vdd.n2884 vdd.n2883 10.6151
R19072 vdd.n2884 vdd.n868 10.6151
R19073 vdd.n2894 vdd.n868 10.6151
R19074 vdd.n2895 vdd.n2894 10.6151
R19075 vdd.n2896 vdd.n2895 10.6151
R19076 vdd.n2896 vdd.n857 10.6151
R19077 vdd.n2906 vdd.n857 10.6151
R19078 vdd.n2907 vdd.n2906 10.6151
R19079 vdd.n2908 vdd.n2907 10.6151
R19080 vdd.n2908 vdd.n844 10.6151
R19081 vdd.n2918 vdd.n844 10.6151
R19082 vdd.n2919 vdd.n2918 10.6151
R19083 vdd.n2921 vdd.n832 10.6151
R19084 vdd.n2931 vdd.n832 10.6151
R19085 vdd.n2932 vdd.n2931 10.6151
R19086 vdd.n2933 vdd.n2932 10.6151
R19087 vdd.n2933 vdd.n820 10.6151
R19088 vdd.n2943 vdd.n820 10.6151
R19089 vdd.n2944 vdd.n2943 10.6151
R19090 vdd.n2990 vdd.n2944 10.6151
R19091 vdd.n2990 vdd.n2989 10.6151
R19092 vdd.n2989 vdd.n2988 10.6151
R19093 vdd.n2988 vdd.n2987 10.6151
R19094 vdd.n2987 vdd.n2985 10.6151
R19095 vdd.n2339 vdd.n2338 10.6151
R19096 vdd.n2339 vdd.n1040 10.6151
R19097 vdd.n2349 vdd.n1040 10.6151
R19098 vdd.n2350 vdd.n2349 10.6151
R19099 vdd.n2351 vdd.n2350 10.6151
R19100 vdd.n2351 vdd.n1028 10.6151
R19101 vdd.n2361 vdd.n1028 10.6151
R19102 vdd.n2362 vdd.n2361 10.6151
R19103 vdd.n2363 vdd.n2362 10.6151
R19104 vdd.n2363 vdd.n1015 10.6151
R19105 vdd.n2373 vdd.n1015 10.6151
R19106 vdd.n2374 vdd.n2373 10.6151
R19107 vdd.n2376 vdd.n1003 10.6151
R19108 vdd.n2386 vdd.n1003 10.6151
R19109 vdd.n2387 vdd.n2386 10.6151
R19110 vdd.n2388 vdd.n2387 10.6151
R19111 vdd.n2388 vdd.n991 10.6151
R19112 vdd.n2398 vdd.n991 10.6151
R19113 vdd.n2399 vdd.n2398 10.6151
R19114 vdd.n2400 vdd.n2399 10.6151
R19115 vdd.n2400 vdd.n980 10.6151
R19116 vdd.n2410 vdd.n980 10.6151
R19117 vdd.n2411 vdd.n2410 10.6151
R19118 vdd.n2412 vdd.n2411 10.6151
R19119 vdd.n2412 vdd.n968 10.6151
R19120 vdd.n2422 vdd.n968 10.6151
R19121 vdd.n2423 vdd.n2422 10.6151
R19122 vdd.n2426 vdd.n2423 10.6151
R19123 vdd.n2426 vdd.n2425 10.6151
R19124 vdd.n2425 vdd.n2424 10.6151
R19125 vdd.n2424 vdd.n951 10.6151
R19126 vdd.n2508 vdd.n951 10.6151
R19127 vdd.n2507 vdd.n2506 10.6151
R19128 vdd.n2506 vdd.n2503 10.6151
R19129 vdd.n2503 vdd.n2502 10.6151
R19130 vdd.n2502 vdd.n2499 10.6151
R19131 vdd.n2499 vdd.n2498 10.6151
R19132 vdd.n2498 vdd.n2495 10.6151
R19133 vdd.n2495 vdd.n2494 10.6151
R19134 vdd.n2494 vdd.n2491 10.6151
R19135 vdd.n2491 vdd.n2490 10.6151
R19136 vdd.n2490 vdd.n2487 10.6151
R19137 vdd.n2487 vdd.n2486 10.6151
R19138 vdd.n2486 vdd.n2483 10.6151
R19139 vdd.n2483 vdd.n2482 10.6151
R19140 vdd.n2482 vdd.n2479 10.6151
R19141 vdd.n2479 vdd.n2478 10.6151
R19142 vdd.n2478 vdd.n2475 10.6151
R19143 vdd.n2475 vdd.n2474 10.6151
R19144 vdd.n2474 vdd.n2471 10.6151
R19145 vdd.n2471 vdd.n2470 10.6151
R19146 vdd.n2470 vdd.n2467 10.6151
R19147 vdd.n2467 vdd.n2466 10.6151
R19148 vdd.n2466 vdd.n2463 10.6151
R19149 vdd.n2463 vdd.n2462 10.6151
R19150 vdd.n2462 vdd.n2459 10.6151
R19151 vdd.n2459 vdd.n2458 10.6151
R19152 vdd.n2458 vdd.n2455 10.6151
R19153 vdd.n2455 vdd.n2454 10.6151
R19154 vdd.n2454 vdd.n2451 10.6151
R19155 vdd.n2451 vdd.n2450 10.6151
R19156 vdd.n2450 vdd.n2447 10.6151
R19157 vdd.n2447 vdd.n2446 10.6151
R19158 vdd.n2443 vdd.n2442 10.6151
R19159 vdd.n2442 vdd.n2440 10.6151
R19160 vdd.n1359 vdd.n1357 10.6151
R19161 vdd.n1357 vdd.n1356 10.6151
R19162 vdd.n1356 vdd.n1354 10.6151
R19163 vdd.n1354 vdd.n1353 10.6151
R19164 vdd.n1353 vdd.n1351 10.6151
R19165 vdd.n1351 vdd.n1350 10.6151
R19166 vdd.n1350 vdd.n1348 10.6151
R19167 vdd.n1348 vdd.n1347 10.6151
R19168 vdd.n1347 vdd.n1345 10.6151
R19169 vdd.n1345 vdd.n1344 10.6151
R19170 vdd.n1344 vdd.n1342 10.6151
R19171 vdd.n1342 vdd.n1341 10.6151
R19172 vdd.n1341 vdd.n1339 10.6151
R19173 vdd.n1339 vdd.n1338 10.6151
R19174 vdd.n1338 vdd.n1336 10.6151
R19175 vdd.n1336 vdd.n1335 10.6151
R19176 vdd.n1335 vdd.n1333 10.6151
R19177 vdd.n1333 vdd.n1332 10.6151
R19178 vdd.n1332 vdd.n1243 10.6151
R19179 vdd.n1243 vdd.n1242 10.6151
R19180 vdd.n1242 vdd.n1240 10.6151
R19181 vdd.n1240 vdd.n1239 10.6151
R19182 vdd.n1239 vdd.n1237 10.6151
R19183 vdd.n1237 vdd.n1236 10.6151
R19184 vdd.n1236 vdd.n1234 10.6151
R19185 vdd.n1234 vdd.n1233 10.6151
R19186 vdd.n1233 vdd.n1231 10.6151
R19187 vdd.n1231 vdd.n1230 10.6151
R19188 vdd.n1230 vdd.n1228 10.6151
R19189 vdd.n1228 vdd.n1227 10.6151
R19190 vdd.n1227 vdd.n955 10.6151
R19191 vdd.n2438 vdd.n955 10.6151
R19192 vdd.n2439 vdd.n2438 10.6151
R19193 vdd.n2337 vdd.n1052 10.6151
R19194 vdd.n1194 vdd.n1052 10.6151
R19195 vdd.n1195 vdd.n1194 10.6151
R19196 vdd.n1198 vdd.n1195 10.6151
R19197 vdd.n1199 vdd.n1198 10.6151
R19198 vdd.n1202 vdd.n1199 10.6151
R19199 vdd.n1203 vdd.n1202 10.6151
R19200 vdd.n1206 vdd.n1203 10.6151
R19201 vdd.n1207 vdd.n1206 10.6151
R19202 vdd.n1210 vdd.n1207 10.6151
R19203 vdd.n1211 vdd.n1210 10.6151
R19204 vdd.n1214 vdd.n1211 10.6151
R19205 vdd.n1215 vdd.n1214 10.6151
R19206 vdd.n1218 vdd.n1215 10.6151
R19207 vdd.n1219 vdd.n1218 10.6151
R19208 vdd.n1222 vdd.n1219 10.6151
R19209 vdd.n1393 vdd.n1222 10.6151
R19210 vdd.n1393 vdd.n1392 10.6151
R19211 vdd.n1392 vdd.n1390 10.6151
R19212 vdd.n1390 vdd.n1387 10.6151
R19213 vdd.n1387 vdd.n1386 10.6151
R19214 vdd.n1386 vdd.n1383 10.6151
R19215 vdd.n1383 vdd.n1382 10.6151
R19216 vdd.n1382 vdd.n1379 10.6151
R19217 vdd.n1379 vdd.n1378 10.6151
R19218 vdd.n1378 vdd.n1375 10.6151
R19219 vdd.n1375 vdd.n1374 10.6151
R19220 vdd.n1374 vdd.n1371 10.6151
R19221 vdd.n1371 vdd.n1370 10.6151
R19222 vdd.n1370 vdd.n1367 10.6151
R19223 vdd.n1367 vdd.n1366 10.6151
R19224 vdd.n1363 vdd.n1362 10.6151
R19225 vdd.n1362 vdd.n1360 10.6151
R19226 vdd.t208 vdd.n2138 10.5435
R19227 vdd.n636 vdd.t162 10.5435
R19228 vdd.n304 vdd.n286 10.4732
R19229 vdd.n249 vdd.n231 10.4732
R19230 vdd.n206 vdd.n188 10.4732
R19231 vdd.n151 vdd.n133 10.4732
R19232 vdd.n109 vdd.n91 10.4732
R19233 vdd.n54 vdd.n36 10.4732
R19234 vdd.n2035 vdd.n2017 10.4732
R19235 vdd.n2090 vdd.n2072 10.4732
R19236 vdd.n1937 vdd.n1919 10.4732
R19237 vdd.n1992 vdd.n1974 10.4732
R19238 vdd.n1840 vdd.n1822 10.4732
R19239 vdd.n1895 vdd.n1877 10.4732
R19240 vdd.n2122 vdd.t169 10.3167
R19241 vdd.n3297 vdd.t157 10.3167
R19242 vdd.t190 vdd.n1466 10.09
R19243 vdd.n2174 vdd.t25 10.09
R19244 vdd.n3245 vdd.t21 10.09
R19245 vdd.n3378 vdd.t160 10.09
R19246 vdd.n1786 vdd.t147 9.86327
R19247 vdd.n3369 vdd.t205 9.86327
R19248 vdd.n2299 vdd.n2298 9.78206
R19249 vdd.n3035 vdd.n3034 9.78206
R19250 vdd.n3102 vdd.n3101 9.78206
R19251 vdd.n2191 vdd.n1393 9.78206
R19252 vdd.n303 vdd.n288 9.69747
R19253 vdd.n248 vdd.n233 9.69747
R19254 vdd.n205 vdd.n190 9.69747
R19255 vdd.n150 vdd.n135 9.69747
R19256 vdd.n108 vdd.n93 9.69747
R19257 vdd.n53 vdd.n38 9.69747
R19258 vdd.n2034 vdd.n2019 9.69747
R19259 vdd.n2089 vdd.n2074 9.69747
R19260 vdd.n1936 vdd.n1921 9.69747
R19261 vdd.n1991 vdd.n1976 9.69747
R19262 vdd.n1839 vdd.n1824 9.69747
R19263 vdd.n1894 vdd.n1879 9.69747
R19264 vdd.t119 vdd.n1760 9.63654
R19265 vdd.n3328 vdd.t171 9.63654
R19266 vdd.n319 vdd.n318 9.45567
R19267 vdd.n264 vdd.n263 9.45567
R19268 vdd.n221 vdd.n220 9.45567
R19269 vdd.n166 vdd.n165 9.45567
R19270 vdd.n124 vdd.n123 9.45567
R19271 vdd.n69 vdd.n68 9.45567
R19272 vdd.n2050 vdd.n2049 9.45567
R19273 vdd.n2105 vdd.n2104 9.45567
R19274 vdd.n1952 vdd.n1951 9.45567
R19275 vdd.n2007 vdd.n2006 9.45567
R19276 vdd.n1855 vdd.n1854 9.45567
R19277 vdd.n1910 vdd.n1909 9.45567
R19278 vdd.n2261 vdd.n1120 9.3005
R19279 vdd.n2260 vdd.n2259 9.3005
R19280 vdd.n1126 vdd.n1125 9.3005
R19281 vdd.n2254 vdd.n1130 9.3005
R19282 vdd.n2253 vdd.n1131 9.3005
R19283 vdd.n2252 vdd.n1132 9.3005
R19284 vdd.n1136 vdd.n1133 9.3005
R19285 vdd.n2247 vdd.n1137 9.3005
R19286 vdd.n2246 vdd.n1138 9.3005
R19287 vdd.n2245 vdd.n1139 9.3005
R19288 vdd.n1143 vdd.n1140 9.3005
R19289 vdd.n2240 vdd.n1144 9.3005
R19290 vdd.n2239 vdd.n1145 9.3005
R19291 vdd.n2238 vdd.n1146 9.3005
R19292 vdd.n1150 vdd.n1147 9.3005
R19293 vdd.n2233 vdd.n1151 9.3005
R19294 vdd.n2232 vdd.n1152 9.3005
R19295 vdd.n2231 vdd.n1153 9.3005
R19296 vdd.n1157 vdd.n1154 9.3005
R19297 vdd.n2226 vdd.n1158 9.3005
R19298 vdd.n2225 vdd.n1159 9.3005
R19299 vdd.n2224 vdd.n2223 9.3005
R19300 vdd.n2222 vdd.n1160 9.3005
R19301 vdd.n2221 vdd.n2220 9.3005
R19302 vdd.n1166 vdd.n1165 9.3005
R19303 vdd.n2215 vdd.n1170 9.3005
R19304 vdd.n2214 vdd.n1171 9.3005
R19305 vdd.n2213 vdd.n1172 9.3005
R19306 vdd.n1176 vdd.n1173 9.3005
R19307 vdd.n2208 vdd.n1177 9.3005
R19308 vdd.n2207 vdd.n1178 9.3005
R19309 vdd.n2206 vdd.n1179 9.3005
R19310 vdd.n1183 vdd.n1180 9.3005
R19311 vdd.n2201 vdd.n1184 9.3005
R19312 vdd.n2200 vdd.n1185 9.3005
R19313 vdd.n2199 vdd.n1186 9.3005
R19314 vdd.n1190 vdd.n1187 9.3005
R19315 vdd.n2194 vdd.n1191 9.3005
R19316 vdd.n2263 vdd.n2262 9.3005
R19317 vdd.n2285 vdd.n1091 9.3005
R19318 vdd.n2284 vdd.n1099 9.3005
R19319 vdd.n1103 vdd.n1100 9.3005
R19320 vdd.n2279 vdd.n1104 9.3005
R19321 vdd.n2278 vdd.n1105 9.3005
R19322 vdd.n2277 vdd.n1106 9.3005
R19323 vdd.n1110 vdd.n1107 9.3005
R19324 vdd.n2272 vdd.n1111 9.3005
R19325 vdd.n2271 vdd.n1112 9.3005
R19326 vdd.n2270 vdd.n1113 9.3005
R19327 vdd.n1117 vdd.n1114 9.3005
R19328 vdd.n2265 vdd.n1118 9.3005
R19329 vdd.n2264 vdd.n1119 9.3005
R19330 vdd.n2297 vdd.n2296 9.3005
R19331 vdd.n1095 vdd.n1094 9.3005
R19332 vdd.n2110 vdd.n1456 9.3005
R19333 vdd.n2112 vdd.n2111 9.3005
R19334 vdd.n1447 vdd.n1446 9.3005
R19335 vdd.n2125 vdd.n2124 9.3005
R19336 vdd.n2126 vdd.n1445 9.3005
R19337 vdd.n2128 vdd.n2127 9.3005
R19338 vdd.n1435 vdd.n1434 9.3005
R19339 vdd.n2142 vdd.n2141 9.3005
R19340 vdd.n2143 vdd.n1433 9.3005
R19341 vdd.n2145 vdd.n2144 9.3005
R19342 vdd.n1424 vdd.n1423 9.3005
R19343 vdd.n2159 vdd.n2158 9.3005
R19344 vdd.n2160 vdd.n1422 9.3005
R19345 vdd.n2162 vdd.n2161 9.3005
R19346 vdd.n1412 vdd.n1411 9.3005
R19347 vdd.n2177 vdd.n2176 9.3005
R19348 vdd.n2178 vdd.n1410 9.3005
R19349 vdd.n2180 vdd.n2179 9.3005
R19350 vdd.n295 vdd.n294 9.3005
R19351 vdd.n290 vdd.n289 9.3005
R19352 vdd.n301 vdd.n300 9.3005
R19353 vdd.n303 vdd.n302 9.3005
R19354 vdd.n286 vdd.n285 9.3005
R19355 vdd.n309 vdd.n308 9.3005
R19356 vdd.n311 vdd.n310 9.3005
R19357 vdd.n283 vdd.n280 9.3005
R19358 vdd.n318 vdd.n317 9.3005
R19359 vdd.n240 vdd.n239 9.3005
R19360 vdd.n235 vdd.n234 9.3005
R19361 vdd.n246 vdd.n245 9.3005
R19362 vdd.n248 vdd.n247 9.3005
R19363 vdd.n231 vdd.n230 9.3005
R19364 vdd.n254 vdd.n253 9.3005
R19365 vdd.n256 vdd.n255 9.3005
R19366 vdd.n228 vdd.n225 9.3005
R19367 vdd.n263 vdd.n262 9.3005
R19368 vdd.n197 vdd.n196 9.3005
R19369 vdd.n192 vdd.n191 9.3005
R19370 vdd.n203 vdd.n202 9.3005
R19371 vdd.n205 vdd.n204 9.3005
R19372 vdd.n188 vdd.n187 9.3005
R19373 vdd.n211 vdd.n210 9.3005
R19374 vdd.n213 vdd.n212 9.3005
R19375 vdd.n185 vdd.n182 9.3005
R19376 vdd.n220 vdd.n219 9.3005
R19377 vdd.n142 vdd.n141 9.3005
R19378 vdd.n137 vdd.n136 9.3005
R19379 vdd.n148 vdd.n147 9.3005
R19380 vdd.n150 vdd.n149 9.3005
R19381 vdd.n133 vdd.n132 9.3005
R19382 vdd.n156 vdd.n155 9.3005
R19383 vdd.n158 vdd.n157 9.3005
R19384 vdd.n130 vdd.n127 9.3005
R19385 vdd.n165 vdd.n164 9.3005
R19386 vdd.n100 vdd.n99 9.3005
R19387 vdd.n95 vdd.n94 9.3005
R19388 vdd.n106 vdd.n105 9.3005
R19389 vdd.n108 vdd.n107 9.3005
R19390 vdd.n91 vdd.n90 9.3005
R19391 vdd.n114 vdd.n113 9.3005
R19392 vdd.n116 vdd.n115 9.3005
R19393 vdd.n88 vdd.n85 9.3005
R19394 vdd.n123 vdd.n122 9.3005
R19395 vdd.n45 vdd.n44 9.3005
R19396 vdd.n40 vdd.n39 9.3005
R19397 vdd.n51 vdd.n50 9.3005
R19398 vdd.n53 vdd.n52 9.3005
R19399 vdd.n36 vdd.n35 9.3005
R19400 vdd.n59 vdd.n58 9.3005
R19401 vdd.n61 vdd.n60 9.3005
R19402 vdd.n33 vdd.n30 9.3005
R19403 vdd.n68 vdd.n67 9.3005
R19404 vdd.n3151 vdd.n3150 9.3005
R19405 vdd.n3152 vdd.n721 9.3005
R19406 vdd.n720 vdd.n718 9.3005
R19407 vdd.n3158 vdd.n717 9.3005
R19408 vdd.n3159 vdd.n716 9.3005
R19409 vdd.n3160 vdd.n715 9.3005
R19410 vdd.n714 vdd.n712 9.3005
R19411 vdd.n3166 vdd.n711 9.3005
R19412 vdd.n3167 vdd.n710 9.3005
R19413 vdd.n3168 vdd.n709 9.3005
R19414 vdd.n708 vdd.n706 9.3005
R19415 vdd.n3174 vdd.n705 9.3005
R19416 vdd.n3175 vdd.n704 9.3005
R19417 vdd.n3176 vdd.n703 9.3005
R19418 vdd.n702 vdd.n700 9.3005
R19419 vdd.n3182 vdd.n699 9.3005
R19420 vdd.n3183 vdd.n698 9.3005
R19421 vdd.n3184 vdd.n697 9.3005
R19422 vdd.n696 vdd.n694 9.3005
R19423 vdd.n3190 vdd.n693 9.3005
R19424 vdd.n3191 vdd.n692 9.3005
R19425 vdd.n3192 vdd.n691 9.3005
R19426 vdd.n690 vdd.n688 9.3005
R19427 vdd.n3198 vdd.n685 9.3005
R19428 vdd.n3199 vdd.n684 9.3005
R19429 vdd.n3200 vdd.n683 9.3005
R19430 vdd.n682 vdd.n680 9.3005
R19431 vdd.n3206 vdd.n679 9.3005
R19432 vdd.n3207 vdd.n678 9.3005
R19433 vdd.n3208 vdd.n677 9.3005
R19434 vdd.n676 vdd.n674 9.3005
R19435 vdd.n3214 vdd.n673 9.3005
R19436 vdd.n3215 vdd.n672 9.3005
R19437 vdd.n3216 vdd.n671 9.3005
R19438 vdd.n670 vdd.n668 9.3005
R19439 vdd.n3221 vdd.n667 9.3005
R19440 vdd.n3231 vdd.n661 9.3005
R19441 vdd.n3233 vdd.n3232 9.3005
R19442 vdd.n652 vdd.n651 9.3005
R19443 vdd.n3248 vdd.n3247 9.3005
R19444 vdd.n3249 vdd.n650 9.3005
R19445 vdd.n3251 vdd.n3250 9.3005
R19446 vdd.n640 vdd.n639 9.3005
R19447 vdd.n3264 vdd.n3263 9.3005
R19448 vdd.n3265 vdd.n638 9.3005
R19449 vdd.n3267 vdd.n3266 9.3005
R19450 vdd.n628 vdd.n627 9.3005
R19451 vdd.n3281 vdd.n3280 9.3005
R19452 vdd.n3282 vdd.n626 9.3005
R19453 vdd.n3284 vdd.n3283 9.3005
R19454 vdd.n617 vdd.n616 9.3005
R19455 vdd.n3300 vdd.n3299 9.3005
R19456 vdd.n3301 vdd.n615 9.3005
R19457 vdd.n3303 vdd.n3302 9.3005
R19458 vdd.n324 vdd.n322 9.3005
R19459 vdd.n3235 vdd.n3234 9.3005
R19460 vdd.n3382 vdd.n3381 9.3005
R19461 vdd.n325 vdd.n323 9.3005
R19462 vdd.n3375 vdd.n334 9.3005
R19463 vdd.n3374 vdd.n335 9.3005
R19464 vdd.n3373 vdd.n336 9.3005
R19465 vdd.n343 vdd.n337 9.3005
R19466 vdd.n3367 vdd.n344 9.3005
R19467 vdd.n3366 vdd.n345 9.3005
R19468 vdd.n3365 vdd.n346 9.3005
R19469 vdd.n354 vdd.n347 9.3005
R19470 vdd.n3359 vdd.n355 9.3005
R19471 vdd.n3358 vdd.n356 9.3005
R19472 vdd.n3357 vdd.n357 9.3005
R19473 vdd.n365 vdd.n358 9.3005
R19474 vdd.n3351 vdd.n366 9.3005
R19475 vdd.n3350 vdd.n367 9.3005
R19476 vdd.n3349 vdd.n368 9.3005
R19477 vdd.n443 vdd.n369 9.3005
R19478 vdd.n447 vdd.n442 9.3005
R19479 vdd.n451 vdd.n450 9.3005
R19480 vdd.n452 vdd.n441 9.3005
R19481 vdd.n456 vdd.n453 9.3005
R19482 vdd.n457 vdd.n440 9.3005
R19483 vdd.n461 vdd.n460 9.3005
R19484 vdd.n462 vdd.n439 9.3005
R19485 vdd.n466 vdd.n463 9.3005
R19486 vdd.n467 vdd.n438 9.3005
R19487 vdd.n471 vdd.n470 9.3005
R19488 vdd.n472 vdd.n437 9.3005
R19489 vdd.n476 vdd.n473 9.3005
R19490 vdd.n477 vdd.n436 9.3005
R19491 vdd.n481 vdd.n480 9.3005
R19492 vdd.n482 vdd.n435 9.3005
R19493 vdd.n486 vdd.n483 9.3005
R19494 vdd.n487 vdd.n434 9.3005
R19495 vdd.n491 vdd.n490 9.3005
R19496 vdd.n492 vdd.n433 9.3005
R19497 vdd.n496 vdd.n493 9.3005
R19498 vdd.n497 vdd.n430 9.3005
R19499 vdd.n501 vdd.n500 9.3005
R19500 vdd.n502 vdd.n429 9.3005
R19501 vdd.n506 vdd.n503 9.3005
R19502 vdd.n507 vdd.n428 9.3005
R19503 vdd.n511 vdd.n510 9.3005
R19504 vdd.n512 vdd.n427 9.3005
R19505 vdd.n516 vdd.n513 9.3005
R19506 vdd.n517 vdd.n426 9.3005
R19507 vdd.n521 vdd.n520 9.3005
R19508 vdd.n522 vdd.n425 9.3005
R19509 vdd.n526 vdd.n523 9.3005
R19510 vdd.n527 vdd.n424 9.3005
R19511 vdd.n531 vdd.n530 9.3005
R19512 vdd.n532 vdd.n423 9.3005
R19513 vdd.n536 vdd.n533 9.3005
R19514 vdd.n537 vdd.n422 9.3005
R19515 vdd.n541 vdd.n540 9.3005
R19516 vdd.n542 vdd.n421 9.3005
R19517 vdd.n546 vdd.n543 9.3005
R19518 vdd.n547 vdd.n418 9.3005
R19519 vdd.n551 vdd.n550 9.3005
R19520 vdd.n552 vdd.n417 9.3005
R19521 vdd.n556 vdd.n553 9.3005
R19522 vdd.n557 vdd.n416 9.3005
R19523 vdd.n561 vdd.n560 9.3005
R19524 vdd.n562 vdd.n415 9.3005
R19525 vdd.n566 vdd.n563 9.3005
R19526 vdd.n567 vdd.n414 9.3005
R19527 vdd.n571 vdd.n570 9.3005
R19528 vdd.n572 vdd.n413 9.3005
R19529 vdd.n576 vdd.n573 9.3005
R19530 vdd.n577 vdd.n412 9.3005
R19531 vdd.n581 vdd.n580 9.3005
R19532 vdd.n582 vdd.n411 9.3005
R19533 vdd.n586 vdd.n583 9.3005
R19534 vdd.n587 vdd.n410 9.3005
R19535 vdd.n591 vdd.n590 9.3005
R19536 vdd.n592 vdd.n409 9.3005
R19537 vdd.n596 vdd.n593 9.3005
R19538 vdd.n598 vdd.n408 9.3005
R19539 vdd.n600 vdd.n599 9.3005
R19540 vdd.n3342 vdd.n3341 9.3005
R19541 vdd.n446 vdd.n444 9.3005
R19542 vdd.n3241 vdd.n655 9.3005
R19543 vdd.n3243 vdd.n3242 9.3005
R19544 vdd.n646 vdd.n645 9.3005
R19545 vdd.n3256 vdd.n3255 9.3005
R19546 vdd.n3257 vdd.n644 9.3005
R19547 vdd.n3259 vdd.n3258 9.3005
R19548 vdd.n633 vdd.n632 9.3005
R19549 vdd.n3272 vdd.n3271 9.3005
R19550 vdd.n3273 vdd.n631 9.3005
R19551 vdd.n3275 vdd.n3274 9.3005
R19552 vdd.n622 vdd.n621 9.3005
R19553 vdd.n3289 vdd.n3288 9.3005
R19554 vdd.n3290 vdd.n620 9.3005
R19555 vdd.n3295 vdd.n3291 9.3005
R19556 vdd.n3294 vdd.n3293 9.3005
R19557 vdd.n3292 vdd.n610 9.3005
R19558 vdd.n3308 vdd.n611 9.3005
R19559 vdd.n3309 vdd.n609 9.3005
R19560 vdd.n3311 vdd.n3310 9.3005
R19561 vdd.n3312 vdd.n608 9.3005
R19562 vdd.n3315 vdd.n3313 9.3005
R19563 vdd.n3316 vdd.n607 9.3005
R19564 vdd.n3318 vdd.n3317 9.3005
R19565 vdd.n3319 vdd.n606 9.3005
R19566 vdd.n3322 vdd.n3320 9.3005
R19567 vdd.n3323 vdd.n605 9.3005
R19568 vdd.n3325 vdd.n3324 9.3005
R19569 vdd.n3326 vdd.n604 9.3005
R19570 vdd.n3330 vdd.n3327 9.3005
R19571 vdd.n3331 vdd.n603 9.3005
R19572 vdd.n3333 vdd.n3332 9.3005
R19573 vdd.n3334 vdd.n602 9.3005
R19574 vdd.n3337 vdd.n3335 9.3005
R19575 vdd.n3338 vdd.n601 9.3005
R19576 vdd.n3340 vdd.n3339 9.3005
R19577 vdd.n3240 vdd.n3239 9.3005
R19578 vdd.n3104 vdd.n656 9.3005
R19579 vdd.n3109 vdd.n3103 9.3005
R19580 vdd.n3119 vdd.n748 9.3005
R19581 vdd.n3120 vdd.n747 9.3005
R19582 vdd.n746 vdd.n744 9.3005
R19583 vdd.n3126 vdd.n743 9.3005
R19584 vdd.n3127 vdd.n742 9.3005
R19585 vdd.n3128 vdd.n741 9.3005
R19586 vdd.n740 vdd.n738 9.3005
R19587 vdd.n3134 vdd.n737 9.3005
R19588 vdd.n3135 vdd.n736 9.3005
R19589 vdd.n3136 vdd.n735 9.3005
R19590 vdd.n734 vdd.n732 9.3005
R19591 vdd.n3141 vdd.n731 9.3005
R19592 vdd.n3142 vdd.n730 9.3005
R19593 vdd.n726 vdd.n725 9.3005
R19594 vdd.n3148 vdd.n3147 9.3005
R19595 vdd.n3149 vdd.n722 9.3005
R19596 vdd.n2190 vdd.n2189 9.3005
R19597 vdd.n2185 vdd.n1395 9.3005
R19598 vdd.n1742 vdd.n1741 9.3005
R19599 vdd.n1498 vdd.n1497 9.3005
R19600 vdd.n1755 vdd.n1754 9.3005
R19601 vdd.n1756 vdd.n1496 9.3005
R19602 vdd.n1758 vdd.n1757 9.3005
R19603 vdd.n1486 vdd.n1485 9.3005
R19604 vdd.n1772 vdd.n1771 9.3005
R19605 vdd.n1773 vdd.n1484 9.3005
R19606 vdd.n1775 vdd.n1774 9.3005
R19607 vdd.n1476 vdd.n1475 9.3005
R19608 vdd.n1789 vdd.n1788 9.3005
R19609 vdd.n1790 vdd.n1474 9.3005
R19610 vdd.n1792 vdd.n1791 9.3005
R19611 vdd.n1463 vdd.n1462 9.3005
R19612 vdd.n1805 vdd.n1804 9.3005
R19613 vdd.n1806 vdd.n1461 9.3005
R19614 vdd.n1808 vdd.n1807 9.3005
R19615 vdd.n1452 vdd.n1451 9.3005
R19616 vdd.n2117 vdd.n2116 9.3005
R19617 vdd.n2118 vdd.n1450 9.3005
R19618 vdd.n2120 vdd.n2119 9.3005
R19619 vdd.n1441 vdd.n1440 9.3005
R19620 vdd.n2133 vdd.n2132 9.3005
R19621 vdd.n2134 vdd.n1439 9.3005
R19622 vdd.n2136 vdd.n2135 9.3005
R19623 vdd.n1429 vdd.n1428 9.3005
R19624 vdd.n2150 vdd.n2149 9.3005
R19625 vdd.n2151 vdd.n1427 9.3005
R19626 vdd.n2153 vdd.n2152 9.3005
R19627 vdd.n1419 vdd.n1418 9.3005
R19628 vdd.n2167 vdd.n2166 9.3005
R19629 vdd.n2168 vdd.n1416 9.3005
R19630 vdd.n2172 vdd.n2171 9.3005
R19631 vdd.n2170 vdd.n1417 9.3005
R19632 vdd.n2169 vdd.n1406 9.3005
R19633 vdd.n1740 vdd.n1508 9.3005
R19634 vdd.n1633 vdd.n1509 9.3005
R19635 vdd.n1635 vdd.n1634 9.3005
R19636 vdd.n1636 vdd.n1628 9.3005
R19637 vdd.n1638 vdd.n1637 9.3005
R19638 vdd.n1639 vdd.n1627 9.3005
R19639 vdd.n1641 vdd.n1640 9.3005
R19640 vdd.n1642 vdd.n1622 9.3005
R19641 vdd.n1644 vdd.n1643 9.3005
R19642 vdd.n1645 vdd.n1621 9.3005
R19643 vdd.n1647 vdd.n1646 9.3005
R19644 vdd.n1648 vdd.n1616 9.3005
R19645 vdd.n1650 vdd.n1649 9.3005
R19646 vdd.n1651 vdd.n1615 9.3005
R19647 vdd.n1653 vdd.n1652 9.3005
R19648 vdd.n1654 vdd.n1610 9.3005
R19649 vdd.n1656 vdd.n1655 9.3005
R19650 vdd.n1657 vdd.n1609 9.3005
R19651 vdd.n1659 vdd.n1658 9.3005
R19652 vdd.n1660 vdd.n1604 9.3005
R19653 vdd.n1662 vdd.n1661 9.3005
R19654 vdd.n1663 vdd.n1603 9.3005
R19655 vdd.n1668 vdd.n1664 9.3005
R19656 vdd.n1669 vdd.n1599 9.3005
R19657 vdd.n1671 vdd.n1670 9.3005
R19658 vdd.n1672 vdd.n1598 9.3005
R19659 vdd.n1674 vdd.n1673 9.3005
R19660 vdd.n1675 vdd.n1593 9.3005
R19661 vdd.n1677 vdd.n1676 9.3005
R19662 vdd.n1678 vdd.n1592 9.3005
R19663 vdd.n1680 vdd.n1679 9.3005
R19664 vdd.n1681 vdd.n1587 9.3005
R19665 vdd.n1683 vdd.n1682 9.3005
R19666 vdd.n1684 vdd.n1586 9.3005
R19667 vdd.n1686 vdd.n1685 9.3005
R19668 vdd.n1687 vdd.n1581 9.3005
R19669 vdd.n1689 vdd.n1688 9.3005
R19670 vdd.n1690 vdd.n1580 9.3005
R19671 vdd.n1692 vdd.n1691 9.3005
R19672 vdd.n1693 vdd.n1575 9.3005
R19673 vdd.n1695 vdd.n1694 9.3005
R19674 vdd.n1696 vdd.n1574 9.3005
R19675 vdd.n1698 vdd.n1697 9.3005
R19676 vdd.n1699 vdd.n1571 9.3005
R19677 vdd.n1705 vdd.n1704 9.3005
R19678 vdd.n1706 vdd.n1570 9.3005
R19679 vdd.n1708 vdd.n1707 9.3005
R19680 vdd.n1709 vdd.n1565 9.3005
R19681 vdd.n1711 vdd.n1710 9.3005
R19682 vdd.n1712 vdd.n1564 9.3005
R19683 vdd.n1714 vdd.n1713 9.3005
R19684 vdd.n1715 vdd.n1559 9.3005
R19685 vdd.n1717 vdd.n1716 9.3005
R19686 vdd.n1718 vdd.n1558 9.3005
R19687 vdd.n1720 vdd.n1719 9.3005
R19688 vdd.n1721 vdd.n1553 9.3005
R19689 vdd.n1723 vdd.n1722 9.3005
R19690 vdd.n1724 vdd.n1552 9.3005
R19691 vdd.n1726 vdd.n1725 9.3005
R19692 vdd.n1727 vdd.n1548 9.3005
R19693 vdd.n1729 vdd.n1728 9.3005
R19694 vdd.n1730 vdd.n1547 9.3005
R19695 vdd.n1732 vdd.n1731 9.3005
R19696 vdd.n1733 vdd.n1546 9.3005
R19697 vdd.n1739 vdd.n1738 9.3005
R19698 vdd.n1747 vdd.n1746 9.3005
R19699 vdd.n1748 vdd.n1502 9.3005
R19700 vdd.n1750 vdd.n1749 9.3005
R19701 vdd.n1492 vdd.n1491 9.3005
R19702 vdd.n1764 vdd.n1763 9.3005
R19703 vdd.n1765 vdd.n1490 9.3005
R19704 vdd.n1767 vdd.n1766 9.3005
R19705 vdd.n1481 vdd.n1480 9.3005
R19706 vdd.n1781 vdd.n1780 9.3005
R19707 vdd.n1782 vdd.n1479 9.3005
R19708 vdd.n1784 vdd.n1783 9.3005
R19709 vdd.n1470 vdd.n1469 9.3005
R19710 vdd.n1797 vdd.n1796 9.3005
R19711 vdd.n1798 vdd.n1468 9.3005
R19712 vdd.n1800 vdd.n1799 9.3005
R19713 vdd.n1458 vdd.n1457 9.3005
R19714 vdd.n1814 vdd.n1813 9.3005
R19715 vdd.n1504 vdd.n1503 9.3005
R19716 vdd.n2026 vdd.n2025 9.3005
R19717 vdd.n2021 vdd.n2020 9.3005
R19718 vdd.n2032 vdd.n2031 9.3005
R19719 vdd.n2034 vdd.n2033 9.3005
R19720 vdd.n2017 vdd.n2016 9.3005
R19721 vdd.n2040 vdd.n2039 9.3005
R19722 vdd.n2042 vdd.n2041 9.3005
R19723 vdd.n2014 vdd.n2011 9.3005
R19724 vdd.n2049 vdd.n2048 9.3005
R19725 vdd.n2081 vdd.n2080 9.3005
R19726 vdd.n2076 vdd.n2075 9.3005
R19727 vdd.n2087 vdd.n2086 9.3005
R19728 vdd.n2089 vdd.n2088 9.3005
R19729 vdd.n2072 vdd.n2071 9.3005
R19730 vdd.n2095 vdd.n2094 9.3005
R19731 vdd.n2097 vdd.n2096 9.3005
R19732 vdd.n2069 vdd.n2066 9.3005
R19733 vdd.n2104 vdd.n2103 9.3005
R19734 vdd.n1928 vdd.n1927 9.3005
R19735 vdd.n1923 vdd.n1922 9.3005
R19736 vdd.n1934 vdd.n1933 9.3005
R19737 vdd.n1936 vdd.n1935 9.3005
R19738 vdd.n1919 vdd.n1918 9.3005
R19739 vdd.n1942 vdd.n1941 9.3005
R19740 vdd.n1944 vdd.n1943 9.3005
R19741 vdd.n1916 vdd.n1913 9.3005
R19742 vdd.n1951 vdd.n1950 9.3005
R19743 vdd.n1983 vdd.n1982 9.3005
R19744 vdd.n1978 vdd.n1977 9.3005
R19745 vdd.n1989 vdd.n1988 9.3005
R19746 vdd.n1991 vdd.n1990 9.3005
R19747 vdd.n1974 vdd.n1973 9.3005
R19748 vdd.n1997 vdd.n1996 9.3005
R19749 vdd.n1999 vdd.n1998 9.3005
R19750 vdd.n1971 vdd.n1968 9.3005
R19751 vdd.n2006 vdd.n2005 9.3005
R19752 vdd.n1831 vdd.n1830 9.3005
R19753 vdd.n1826 vdd.n1825 9.3005
R19754 vdd.n1837 vdd.n1836 9.3005
R19755 vdd.n1839 vdd.n1838 9.3005
R19756 vdd.n1822 vdd.n1821 9.3005
R19757 vdd.n1845 vdd.n1844 9.3005
R19758 vdd.n1847 vdd.n1846 9.3005
R19759 vdd.n1819 vdd.n1816 9.3005
R19760 vdd.n1854 vdd.n1853 9.3005
R19761 vdd.n1886 vdd.n1885 9.3005
R19762 vdd.n1881 vdd.n1880 9.3005
R19763 vdd.n1892 vdd.n1891 9.3005
R19764 vdd.n1894 vdd.n1893 9.3005
R19765 vdd.n1877 vdd.n1876 9.3005
R19766 vdd.n1900 vdd.n1899 9.3005
R19767 vdd.n1902 vdd.n1901 9.3005
R19768 vdd.n1874 vdd.n1871 9.3005
R19769 vdd.n1909 vdd.n1908 9.3005
R19770 vdd.n1760 vdd.t115 9.18308
R19771 vdd.n3328 vdd.t181 9.18308
R19772 vdd.n1786 vdd.t123 8.95635
R19773 vdd.t136 vdd.n3369 8.95635
R19774 vdd.n300 vdd.n299 8.92171
R19775 vdd.n245 vdd.n244 8.92171
R19776 vdd.n202 vdd.n201 8.92171
R19777 vdd.n147 vdd.n146 8.92171
R19778 vdd.n105 vdd.n104 8.92171
R19779 vdd.n50 vdd.n49 8.92171
R19780 vdd.n2031 vdd.n2030 8.92171
R19781 vdd.n2086 vdd.n2085 8.92171
R19782 vdd.n1933 vdd.n1932 8.92171
R19783 vdd.n1988 vdd.n1987 8.92171
R19784 vdd.n1836 vdd.n1835 8.92171
R19785 vdd.n1891 vdd.n1890 8.92171
R19786 vdd.n223 vdd.n125 8.81535
R19787 vdd.n2009 vdd.n1911 8.81535
R19788 vdd.n1466 vdd.t144 8.72962
R19789 vdd.t186 vdd.n3378 8.72962
R19790 vdd.n2122 vdd.t125 8.50289
R19791 vdd.n3297 vdd.t121 8.50289
R19792 vdd.n28 vdd.n14 8.42249
R19793 vdd.n2138 vdd.t178 8.27616
R19794 vdd.t113 vdd.n636 8.27616
R19795 vdd.n3384 vdd.n3383 8.16225
R19796 vdd.n2109 vdd.n2108 8.16225
R19797 vdd.n296 vdd.n290 8.14595
R19798 vdd.n241 vdd.n235 8.14595
R19799 vdd.n198 vdd.n192 8.14595
R19800 vdd.n143 vdd.n137 8.14595
R19801 vdd.n101 vdd.n95 8.14595
R19802 vdd.n46 vdd.n40 8.14595
R19803 vdd.n2027 vdd.n2021 8.14595
R19804 vdd.n2082 vdd.n2076 8.14595
R19805 vdd.n1929 vdd.n1923 8.14595
R19806 vdd.n1984 vdd.n1978 8.14595
R19807 vdd.n1832 vdd.n1826 8.14595
R19808 vdd.n1887 vdd.n1881 8.14595
R19809 vdd.t42 vdd.n1500 7.8227
R19810 vdd.t46 vdd.n363 7.8227
R19811 vdd.n2341 vdd.n1047 7.70933
R19812 vdd.n2341 vdd.n1050 7.70933
R19813 vdd.n2347 vdd.n1036 7.70933
R19814 vdd.n2353 vdd.n1036 7.70933
R19815 vdd.n2353 vdd.n1030 7.70933
R19816 vdd.n2359 vdd.n1030 7.70933
R19817 vdd.n2365 vdd.n1023 7.70933
R19818 vdd.n2365 vdd.n1026 7.70933
R19819 vdd.n2371 vdd.n1019 7.70933
R19820 vdd.n2378 vdd.n1005 7.70933
R19821 vdd.n2384 vdd.n1005 7.70933
R19822 vdd.n2390 vdd.n999 7.70933
R19823 vdd.n2396 vdd.n995 7.70933
R19824 vdd.n2402 vdd.n989 7.70933
R19825 vdd.n2414 vdd.n976 7.70933
R19826 vdd.n2420 vdd.n970 7.70933
R19827 vdd.n2420 vdd.n963 7.70933
R19828 vdd.n2428 vdd.n963 7.70933
R19829 vdd.n2510 vdd.n947 7.70933
R19830 vdd.n2862 vdd.n899 7.70933
R19831 vdd.n2874 vdd.n888 7.70933
R19832 vdd.n2874 vdd.n882 7.70933
R19833 vdd.n2880 vdd.n882 7.70933
R19834 vdd.n2886 vdd.n876 7.70933
R19835 vdd.n2892 vdd.n872 7.70933
R19836 vdd.n2898 vdd.n866 7.70933
R19837 vdd.n2910 vdd.n853 7.70933
R19838 vdd.n2916 vdd.n846 7.70933
R19839 vdd.n2916 vdd.n849 7.70933
R19840 vdd.n2923 vdd.n841 7.70933
R19841 vdd.n2929 vdd.n828 7.70933
R19842 vdd.n2935 vdd.n828 7.70933
R19843 vdd.n2941 vdd.n822 7.70933
R19844 vdd.n2941 vdd.n814 7.70933
R19845 vdd.n2992 vdd.n814 7.70933
R19846 vdd.n2992 vdd.n817 7.70933
R19847 vdd.n2998 vdd.n774 7.70933
R19848 vdd.n3068 vdd.n774 7.70933
R19849 vdd.n2921 vdd.n2920 7.49318
R19850 vdd.n2375 vdd.n2374 7.49318
R19851 vdd.n295 vdd.n292 7.3702
R19852 vdd.n240 vdd.n237 7.3702
R19853 vdd.n197 vdd.n194 7.3702
R19854 vdd.n142 vdd.n139 7.3702
R19855 vdd.n100 vdd.n97 7.3702
R19856 vdd.n45 vdd.n42 7.3702
R19857 vdd.n2026 vdd.n2023 7.3702
R19858 vdd.n2081 vdd.n2078 7.3702
R19859 vdd.n1928 vdd.n1925 7.3702
R19860 vdd.n1983 vdd.n1980 7.3702
R19861 vdd.n1831 vdd.n1828 7.3702
R19862 vdd.n1886 vdd.n1883 7.3702
R19863 vdd.n2359 vdd.t94 7.36923
R19864 vdd.t104 vdd.n822 7.36923
R19865 vdd.n2435 vdd.t243 7.25587
R19866 vdd.n2779 vdd.t252 7.25587
R19867 vdd.n1669 vdd.n1668 6.98232
R19868 vdd.n2225 vdd.n2224 6.98232
R19869 vdd.n547 vdd.n546 6.98232
R19870 vdd.n3152 vdd.n3151 6.98232
R19871 vdd.n2156 vdd.t117 6.91577
R19872 vdd.n3261 vdd.t211 6.91577
R19873 vdd.t196 vdd.n1437 6.68904
R19874 vdd.n3277 vdd.t164 6.68904
R19875 vdd.n2114 vdd.t131 6.46231
R19876 vdd.n3305 vdd.t133 6.46231
R19877 vdd.n3384 vdd.n321 6.32949
R19878 vdd.n2108 vdd.n2107 6.32949
R19879 vdd.t193 vdd.n1465 6.23558
R19880 vdd.t129 vdd.n332 6.23558
R19881 vdd.n1778 vdd.t149 6.00885
R19882 vdd.n3363 vdd.t127 6.00885
R19883 vdd.t108 vdd.n976 5.89549
R19884 vdd.n2886 vdd.t254 5.89549
R19885 vdd.n296 vdd.n295 5.81868
R19886 vdd.n241 vdd.n240 5.81868
R19887 vdd.n198 vdd.n197 5.81868
R19888 vdd.n143 vdd.n142 5.81868
R19889 vdd.n101 vdd.n100 5.81868
R19890 vdd.n46 vdd.n45 5.81868
R19891 vdd.n2027 vdd.n2026 5.81868
R19892 vdd.n2082 vdd.n2081 5.81868
R19893 vdd.n1929 vdd.n1928 5.81868
R19894 vdd.n1984 vdd.n1983 5.81868
R19895 vdd.n1832 vdd.n1831 5.81868
R19896 vdd.n1887 vdd.n1886 5.81868
R19897 vdd.n2518 vdd.n2517 5.77611
R19898 vdd.n1274 vdd.n1273 5.77611
R19899 vdd.n2791 vdd.n2790 5.77611
R19900 vdd.n3007 vdd.n806 5.77611
R19901 vdd.n3073 vdd.n770 5.77611
R19902 vdd.n2685 vdd.n2623 5.77611
R19903 vdd.n2443 vdd.n954 5.77611
R19904 vdd.n1363 vdd.n1226 5.77611
R19905 vdd.n1738 vdd.n1512 5.62474
R19906 vdd.n2188 vdd.n2185 5.62474
R19907 vdd.n3342 vdd.n407 5.62474
R19908 vdd.n3107 vdd.n3104 5.62474
R19909 vdd.t100 vdd.n999 5.55539
R19910 vdd.n2390 vdd.t103 5.55539
R19911 vdd.t249 vdd.n853 5.55539
R19912 vdd.n2910 vdd.t111 5.55539
R19913 vdd.n1019 vdd.t67 5.44203
R19914 vdd.n2923 vdd.t35 5.44203
R19915 vdd.n1488 vdd.t149 5.32866
R19916 vdd.n2347 vdd.t17 5.32866
R19917 vdd.n1309 vdd.t59 5.32866
R19918 vdd.n2868 vdd.t63 5.32866
R19919 vdd.n817 vdd.t13 5.32866
R19920 vdd.t127 vdd.n3362 5.32866
R19921 vdd.n1794 vdd.t193 5.10193
R19922 vdd.n3371 vdd.t129 5.10193
R19923 vdd.n299 vdd.n290 5.04292
R19924 vdd.n244 vdd.n235 5.04292
R19925 vdd.n201 vdd.n192 5.04292
R19926 vdd.n146 vdd.n137 5.04292
R19927 vdd.n104 vdd.n95 5.04292
R19928 vdd.n49 vdd.n40 5.04292
R19929 vdd.n2030 vdd.n2021 5.04292
R19930 vdd.n2085 vdd.n2076 5.04292
R19931 vdd.n1932 vdd.n1923 5.04292
R19932 vdd.n1987 vdd.n1978 5.04292
R19933 vdd.n1835 vdd.n1826 5.04292
R19934 vdd.n1890 vdd.n1881 5.04292
R19935 vdd.n2396 vdd.t256 4.98857
R19936 vdd.n866 vdd.t266 4.98857
R19937 vdd.n1810 vdd.t131 4.8752
R19938 vdd.t88 vdd.t262 4.8752
R19939 vdd.t112 vdd.t250 4.8752
R19940 vdd.t260 vdd.t107 4.8752
R19941 vdd.t105 vdd.t97 4.8752
R19942 vdd.t133 vdd.n328 4.8752
R19943 vdd.n2519 vdd.n2518 4.83952
R19944 vdd.n1273 vdd.n1272 4.83952
R19945 vdd.n2792 vdd.n2791 4.83952
R19946 vdd.n806 vdd.n801 4.83952
R19947 vdd.n770 vdd.n765 4.83952
R19948 vdd.n2682 vdd.n2623 4.83952
R19949 vdd.n2446 vdd.n954 4.83952
R19950 vdd.n1366 vdd.n1226 4.83952
R19951 vdd.n2193 vdd.n2192 4.74817
R19952 vdd.n1399 vdd.n1394 4.74817
R19953 vdd.n1096 vdd.n1093 4.74817
R19954 vdd.n2286 vdd.n1092 4.74817
R19955 vdd.n2291 vdd.n1093 4.74817
R19956 vdd.n2290 vdd.n1092 4.74817
R19957 vdd.n664 vdd.n662 4.74817
R19958 vdd.n3222 vdd.n665 4.74817
R19959 vdd.n3225 vdd.n665 4.74817
R19960 vdd.n3226 vdd.n664 4.74817
R19961 vdd.n3114 vdd.n749 4.74817
R19962 vdd.n3110 vdd.n751 4.74817
R19963 vdd.n3113 vdd.n751 4.74817
R19964 vdd.n3118 vdd.n749 4.74817
R19965 vdd.n2192 vdd.n1192 4.74817
R19966 vdd.n1396 vdd.n1394 4.74817
R19967 vdd.n321 vdd.n320 4.7074
R19968 vdd.n223 vdd.n222 4.7074
R19969 vdd.n2107 vdd.n2106 4.7074
R19970 vdd.n2009 vdd.n2008 4.7074
R19971 vdd.n2130 vdd.t196 4.64847
R19972 vdd.n2371 vdd.t95 4.64847
R19973 vdd.n989 vdd.t110 4.64847
R19974 vdd.n2892 vdd.t96 4.64847
R19975 vdd.n841 vdd.t89 4.64847
R19976 vdd.n3286 vdd.t164 4.64847
R19977 vdd.n1431 vdd.t117 4.42174
R19978 vdd.t211 vdd.n635 4.42174
R19979 vdd.n300 vdd.n288 4.26717
R19980 vdd.n245 vdd.n233 4.26717
R19981 vdd.n202 vdd.n190 4.26717
R19982 vdd.n147 vdd.n135 4.26717
R19983 vdd.n105 vdd.n93 4.26717
R19984 vdd.n50 vdd.n38 4.26717
R19985 vdd.n2031 vdd.n2019 4.26717
R19986 vdd.n2086 vdd.n2074 4.26717
R19987 vdd.n1933 vdd.n1921 4.26717
R19988 vdd.n1988 vdd.n1976 4.26717
R19989 vdd.n1836 vdd.n1824 4.26717
R19990 vdd.n1891 vdd.n1879 4.26717
R19991 vdd.n321 vdd.n223 4.10845
R19992 vdd.n2107 vdd.n2009 4.10845
R19993 vdd.n277 vdd.t146 4.06363
R19994 vdd.n277 vdd.t199 4.06363
R19995 vdd.n275 vdd.t226 4.06363
R19996 vdd.n275 vdd.t233 4.06363
R19997 vdd.n273 vdd.t237 4.06363
R19998 vdd.n273 vdd.t151 4.06363
R19999 vdd.n271 vdd.t176 4.06363
R20000 vdd.n271 vdd.t236 4.06363
R20001 vdd.n269 vdd.t238 4.06363
R20002 vdd.n269 vdd.t175 4.06363
R20003 vdd.n267 vdd.t180 4.06363
R20004 vdd.n267 vdd.t184 4.06363
R20005 vdd.n265 vdd.t219 4.06363
R20006 vdd.n265 vdd.t135 4.06363
R20007 vdd.n179 vdd.t128 4.06363
R20008 vdd.n179 vdd.t182 4.06363
R20009 vdd.n177 vdd.t213 4.06363
R20010 vdd.n177 vdd.t227 4.06363
R20011 vdd.n175 vdd.t224 4.06363
R20012 vdd.n175 vdd.t130 4.06363
R20013 vdd.n173 vdd.t159 4.06363
R20014 vdd.n173 vdd.t229 4.06363
R20015 vdd.n171 vdd.t230 4.06363
R20016 vdd.n171 vdd.t158 4.06363
R20017 vdd.n169 vdd.t163 4.06363
R20018 vdd.n169 vdd.t165 4.06363
R20019 vdd.n167 vdd.t212 4.06363
R20020 vdd.n167 vdd.t114 4.06363
R20021 vdd.n82 vdd.t143 4.06363
R20022 vdd.n82 vdd.t218 4.06363
R20023 vdd.n80 vdd.t137 4.06363
R20024 vdd.n80 vdd.t206 4.06363
R20025 vdd.n78 vdd.t161 4.06363
R20026 vdd.n78 vdd.t223 4.06363
R20027 vdd.n76 vdd.t134 4.06363
R20028 vdd.n76 vdd.t187 4.06363
R20029 vdd.n74 vdd.t122 4.06363
R20030 vdd.n74 vdd.t168 4.06363
R20031 vdd.n72 vdd.t234 4.06363
R20032 vdd.n72 vdd.t217 4.06363
R20033 vdd.n70 vdd.t222 4.06363
R20034 vdd.n70 vdd.t177 4.06363
R20035 vdd.n2051 vdd.t195 4.06363
R20036 vdd.n2051 vdd.t140 4.06363
R20037 vdd.n2053 vdd.t240 4.06363
R20038 vdd.n2053 vdd.t216 4.06363
R20039 vdd.n2055 vdd.t214 4.06363
R20040 vdd.n2055 vdd.t174 4.06363
R20041 vdd.n2057 vdd.t167 4.06363
R20042 vdd.n2057 vdd.t215 4.06363
R20043 vdd.n2059 vdd.t202 4.06363
R20044 vdd.n2059 vdd.t201 4.06363
R20045 vdd.n2061 vdd.t166 4.06363
R20046 vdd.n2061 vdd.t142 4.06363
R20047 vdd.n2063 vdd.t139 4.06363
R20048 vdd.n2063 vdd.t200 4.06363
R20049 vdd.n1953 vdd.t183 4.06363
R20050 vdd.n1953 vdd.t118 4.06363
R20051 vdd.n1955 vdd.t232 4.06363
R20052 vdd.n1955 vdd.t209 4.06363
R20053 vdd.n1957 vdd.t203 4.06363
R20054 vdd.n1957 vdd.t156 4.06363
R20055 vdd.n1959 vdd.t145 4.06363
R20056 vdd.n1959 vdd.t204 4.06363
R20057 vdd.n1961 vdd.t194 4.06363
R20058 vdd.n1961 vdd.t191 4.06363
R20059 vdd.n1963 vdd.t148 4.06363
R20060 vdd.n1963 vdd.t124 4.06363
R20061 vdd.n1965 vdd.t116 4.06363
R20062 vdd.n1965 vdd.t189 4.06363
R20063 vdd.n1856 vdd.t179 4.06363
R20064 vdd.n1856 vdd.t225 4.06363
R20065 vdd.n1858 vdd.t197 4.06363
R20066 vdd.n1858 vdd.t235 4.06363
R20067 vdd.n1860 vdd.t170 4.06363
R20068 vdd.n1860 vdd.t126 4.06363
R20069 vdd.n1862 vdd.t188 4.06363
R20070 vdd.n1862 vdd.t132 4.06363
R20071 vdd.n1864 vdd.t228 4.06363
R20072 vdd.n1864 vdd.t239 4.06363
R20073 vdd.n1866 vdd.t207 4.06363
R20074 vdd.n1866 vdd.t138 4.06363
R20075 vdd.n1868 vdd.t192 4.06363
R20076 vdd.n1868 vdd.t150 4.06363
R20077 vdd.n26 vdd.t3 3.9605
R20078 vdd.n26 vdd.t7 3.9605
R20079 vdd.n23 vdd.t0 3.9605
R20080 vdd.n23 vdd.t1 3.9605
R20081 vdd.n21 vdd.t6 3.9605
R20082 vdd.n21 vdd.t242 3.9605
R20083 vdd.n20 vdd.t2 3.9605
R20084 vdd.n20 vdd.t11 3.9605
R20085 vdd.n15 vdd.t91 3.9605
R20086 vdd.n15 vdd.t4 3.9605
R20087 vdd.n16 vdd.t9 3.9605
R20088 vdd.n16 vdd.t10 3.9605
R20089 vdd.n18 vdd.t8 3.9605
R20090 vdd.n18 vdd.t5 3.9605
R20091 vdd.n25 vdd.t90 3.9605
R20092 vdd.n25 vdd.t241 3.9605
R20093 vdd.n2428 vdd.t264 3.85492
R20094 vdd.n1309 vdd.t264 3.85492
R20095 vdd.n2868 vdd.t98 3.85492
R20096 vdd.t98 vdd.n888 3.85492
R20097 vdd.n7 vdd.t106 3.61217
R20098 vdd.n7 vdd.t267 3.61217
R20099 vdd.n8 vdd.t261 3.61217
R20100 vdd.n8 vdd.t255 3.61217
R20101 vdd.n10 vdd.t253 3.61217
R20102 vdd.n10 vdd.t99 3.61217
R20103 vdd.n12 vdd.t102 3.61217
R20104 vdd.n12 vdd.t248 3.61217
R20105 vdd.n5 vdd.t246 3.61217
R20106 vdd.n5 vdd.t259 3.61217
R20107 vdd.n3 vdd.t265 3.61217
R20108 vdd.n3 vdd.t244 3.61217
R20109 vdd.n1 vdd.t109 3.61217
R20110 vdd.n1 vdd.t251 3.61217
R20111 vdd.n0 vdd.t257 3.61217
R20112 vdd.n0 vdd.t263 3.61217
R20113 vdd.n1744 vdd.t42 3.51482
R20114 vdd.n3347 vdd.t46 3.51482
R20115 vdd.n304 vdd.n303 3.49141
R20116 vdd.n249 vdd.n248 3.49141
R20117 vdd.n206 vdd.n205 3.49141
R20118 vdd.n151 vdd.n150 3.49141
R20119 vdd.n109 vdd.n108 3.49141
R20120 vdd.n54 vdd.n53 3.49141
R20121 vdd.n2035 vdd.n2034 3.49141
R20122 vdd.n2090 vdd.n2089 3.49141
R20123 vdd.n1937 vdd.n1936 3.49141
R20124 vdd.n1992 vdd.n1991 3.49141
R20125 vdd.n1840 vdd.n1839 3.49141
R20126 vdd.n1895 vdd.n1894 3.49141
R20127 vdd.n2582 vdd.t245 3.40145
R20128 vdd.n2855 vdd.t247 3.40145
R20129 vdd.n2920 vdd.n2919 3.12245
R20130 vdd.n2376 vdd.n2375 3.12245
R20131 vdd.n2147 vdd.t178 3.06136
R20132 vdd.n1026 vdd.t95 3.06136
R20133 vdd.n2408 vdd.t110 3.06136
R20134 vdd.n2764 vdd.t96 3.06136
R20135 vdd.n2929 vdd.t89 3.06136
R20136 vdd.n3269 vdd.t113 3.06136
R20137 vdd.t125 vdd.n1443 2.83463
R20138 vdd.n624 vdd.t121 2.83463
R20139 vdd.n1330 vdd.t256 2.72126
R20140 vdd.n2904 vdd.t266 2.72126
R20141 vdd.n307 vdd.n286 2.71565
R20142 vdd.n252 vdd.n231 2.71565
R20143 vdd.n209 vdd.n188 2.71565
R20144 vdd.n154 vdd.n133 2.71565
R20145 vdd.n112 vdd.n91 2.71565
R20146 vdd.n57 vdd.n36 2.71565
R20147 vdd.n2038 vdd.n2017 2.71565
R20148 vdd.n2093 vdd.n2072 2.71565
R20149 vdd.n1940 vdd.n1919 2.71565
R20150 vdd.n1995 vdd.n1974 2.71565
R20151 vdd.n1843 vdd.n1822 2.71565
R20152 vdd.n1898 vdd.n1877 2.71565
R20153 vdd.n1811 vdd.t144 2.6079
R20154 vdd.n3379 vdd.t186 2.6079
R20155 vdd.t250 vdd.n970 2.49453
R20156 vdd.n2880 vdd.t260 2.49453
R20157 vdd.n294 vdd.n293 2.4129
R20158 vdd.n239 vdd.n238 2.4129
R20159 vdd.n196 vdd.n195 2.4129
R20160 vdd.n141 vdd.n140 2.4129
R20161 vdd.n99 vdd.n98 2.4129
R20162 vdd.n44 vdd.n43 2.4129
R20163 vdd.n2025 vdd.n2024 2.4129
R20164 vdd.n2080 vdd.n2079 2.4129
R20165 vdd.n1927 vdd.n1926 2.4129
R20166 vdd.n1982 vdd.n1981 2.4129
R20167 vdd.n1830 vdd.n1829 2.4129
R20168 vdd.n1885 vdd.n1884 2.4129
R20169 vdd.t123 vdd.n1472 2.38117
R20170 vdd.n1050 vdd.t17 2.38117
R20171 vdd.n2435 vdd.t59 2.38117
R20172 vdd.n2779 vdd.t63 2.38117
R20173 vdd.n2998 vdd.t13 2.38117
R20174 vdd.n3370 vdd.t136 2.38117
R20175 vdd.n2298 vdd.n1093 2.27742
R20176 vdd.n2298 vdd.n1092 2.27742
R20177 vdd.n3034 vdd.n665 2.27742
R20178 vdd.n3034 vdd.n664 2.27742
R20179 vdd.n3102 vdd.n751 2.27742
R20180 vdd.n3102 vdd.n749 2.27742
R20181 vdd.n2192 vdd.n2191 2.27742
R20182 vdd.n2191 vdd.n1394 2.27742
R20183 vdd.n1769 vdd.t115 2.15444
R20184 vdd.n2384 vdd.t100 2.15444
R20185 vdd.n1330 vdd.t103 2.15444
R20186 vdd.n2904 vdd.t249 2.15444
R20187 vdd.t111 vdd.n846 2.15444
R20188 vdd.n3361 vdd.t181 2.15444
R20189 vdd.n308 vdd.n284 1.93989
R20190 vdd.n253 vdd.n229 1.93989
R20191 vdd.n210 vdd.n186 1.93989
R20192 vdd.n155 vdd.n131 1.93989
R20193 vdd.n113 vdd.n89 1.93989
R20194 vdd.n58 vdd.n34 1.93989
R20195 vdd.n2039 vdd.n2015 1.93989
R20196 vdd.n2094 vdd.n2070 1.93989
R20197 vdd.n1941 vdd.n1917 1.93989
R20198 vdd.n1996 vdd.n1972 1.93989
R20199 vdd.n1844 vdd.n1820 1.93989
R20200 vdd.n1899 vdd.n1875 1.93989
R20201 vdd.n2408 vdd.t108 1.81434
R20202 vdd.n2764 vdd.t254 1.81434
R20203 vdd.n1761 vdd.t119 1.70098
R20204 vdd.n3355 vdd.t171 1.70098
R20205 vdd.n2402 vdd.t262 1.58761
R20206 vdd.n872 vdd.t105 1.58761
R20207 vdd.n1777 vdd.t147 1.47425
R20208 vdd.n349 vdd.t205 1.47425
R20209 vdd.n1802 vdd.t190 1.24752
R20210 vdd.t25 vdd.n1407 1.24752
R20211 vdd.n2378 vdd.t93 1.24752
R20212 vdd.n995 vdd.t88 1.24752
R20213 vdd.n2898 vdd.t97 1.24752
R20214 vdd.n849 vdd.t92 1.24752
R20215 vdd.n659 vdd.t21 1.24752
R20216 vdd.t160 vdd.n3377 1.24752
R20217 vdd.n319 vdd.n279 1.16414
R20218 vdd.n312 vdd.n311 1.16414
R20219 vdd.n264 vdd.n224 1.16414
R20220 vdd.n257 vdd.n256 1.16414
R20221 vdd.n221 vdd.n181 1.16414
R20222 vdd.n214 vdd.n213 1.16414
R20223 vdd.n166 vdd.n126 1.16414
R20224 vdd.n159 vdd.n158 1.16414
R20225 vdd.n124 vdd.n84 1.16414
R20226 vdd.n117 vdd.n116 1.16414
R20227 vdd.n69 vdd.n29 1.16414
R20228 vdd.n62 vdd.n61 1.16414
R20229 vdd.n2050 vdd.n2010 1.16414
R20230 vdd.n2043 vdd.n2042 1.16414
R20231 vdd.n2105 vdd.n2065 1.16414
R20232 vdd.n2098 vdd.n2097 1.16414
R20233 vdd.n1952 vdd.n1912 1.16414
R20234 vdd.n1945 vdd.n1944 1.16414
R20235 vdd.n2007 vdd.n1967 1.16414
R20236 vdd.n2000 vdd.n1999 1.16414
R20237 vdd.n1855 vdd.n1815 1.16414
R20238 vdd.n1848 vdd.n1847 1.16414
R20239 vdd.n1910 vdd.n1870 1.16414
R20240 vdd.n1903 vdd.n1902 1.16414
R20241 vdd.n1454 vdd.t169 1.02079
R20242 vdd.t67 vdd.t93 1.02079
R20243 vdd.t92 vdd.t35 1.02079
R20244 vdd.t157 vdd.n613 1.02079
R20245 vdd.n1633 vdd.n1512 0.970197
R20246 vdd.n2189 vdd.n2188 0.970197
R20247 vdd.n599 vdd.n407 0.970197
R20248 vdd.n3109 vdd.n3107 0.970197
R20249 vdd.n2108 vdd.n28 0.956323
R20250 vdd vdd.n3384 0.94849
R20251 vdd.n2139 vdd.t208 0.794056
R20252 vdd.n3278 vdd.t162 0.794056
R20253 vdd.n2155 vdd.t154 0.567326
R20254 vdd.t152 vdd.n642 0.567326
R20255 vdd.n2179 vdd.n1094 0.482207
R20256 vdd.n3234 vdd.n3233 0.482207
R20257 vdd.n444 vdd.n443 0.482207
R20258 vdd.n3341 vdd.n3340 0.482207
R20259 vdd.n3240 vdd.n656 0.482207
R20260 vdd.n2169 vdd.n1395 0.482207
R20261 vdd.n1740 vdd.n1739 0.482207
R20262 vdd.n1546 vdd.n1503 0.482207
R20263 vdd.n4 vdd.n2 0.459552
R20264 vdd.n11 vdd.n9 0.459552
R20265 vdd.t243 vdd.n947 0.453961
R20266 vdd.n2862 vdd.t252 0.453961
R20267 vdd.n317 vdd.n316 0.388379
R20268 vdd.n283 vdd.n281 0.388379
R20269 vdd.n262 vdd.n261 0.388379
R20270 vdd.n228 vdd.n226 0.388379
R20271 vdd.n219 vdd.n218 0.388379
R20272 vdd.n185 vdd.n183 0.388379
R20273 vdd.n164 vdd.n163 0.388379
R20274 vdd.n130 vdd.n128 0.388379
R20275 vdd.n122 vdd.n121 0.388379
R20276 vdd.n88 vdd.n86 0.388379
R20277 vdd.n67 vdd.n66 0.388379
R20278 vdd.n33 vdd.n31 0.388379
R20279 vdd.n2048 vdd.n2047 0.388379
R20280 vdd.n2014 vdd.n2012 0.388379
R20281 vdd.n2103 vdd.n2102 0.388379
R20282 vdd.n2069 vdd.n2067 0.388379
R20283 vdd.n1950 vdd.n1949 0.388379
R20284 vdd.n1916 vdd.n1914 0.388379
R20285 vdd.n2005 vdd.n2004 0.388379
R20286 vdd.n1971 vdd.n1969 0.388379
R20287 vdd.n1853 vdd.n1852 0.388379
R20288 vdd.n1819 vdd.n1817 0.388379
R20289 vdd.n1908 vdd.n1907 0.388379
R20290 vdd.n1874 vdd.n1872 0.388379
R20291 vdd.n19 vdd.n17 0.387128
R20292 vdd.n24 vdd.n22 0.387128
R20293 vdd.n6 vdd.n4 0.358259
R20294 vdd.n13 vdd.n11 0.358259
R20295 vdd.n268 vdd.n266 0.358259
R20296 vdd.n270 vdd.n268 0.358259
R20297 vdd.n272 vdd.n270 0.358259
R20298 vdd.n274 vdd.n272 0.358259
R20299 vdd.n276 vdd.n274 0.358259
R20300 vdd.n278 vdd.n276 0.358259
R20301 vdd.n320 vdd.n278 0.358259
R20302 vdd.n170 vdd.n168 0.358259
R20303 vdd.n172 vdd.n170 0.358259
R20304 vdd.n174 vdd.n172 0.358259
R20305 vdd.n176 vdd.n174 0.358259
R20306 vdd.n178 vdd.n176 0.358259
R20307 vdd.n180 vdd.n178 0.358259
R20308 vdd.n222 vdd.n180 0.358259
R20309 vdd.n73 vdd.n71 0.358259
R20310 vdd.n75 vdd.n73 0.358259
R20311 vdd.n77 vdd.n75 0.358259
R20312 vdd.n79 vdd.n77 0.358259
R20313 vdd.n81 vdd.n79 0.358259
R20314 vdd.n83 vdd.n81 0.358259
R20315 vdd.n125 vdd.n83 0.358259
R20316 vdd.n2106 vdd.n2064 0.358259
R20317 vdd.n2064 vdd.n2062 0.358259
R20318 vdd.n2062 vdd.n2060 0.358259
R20319 vdd.n2060 vdd.n2058 0.358259
R20320 vdd.n2058 vdd.n2056 0.358259
R20321 vdd.n2056 vdd.n2054 0.358259
R20322 vdd.n2054 vdd.n2052 0.358259
R20323 vdd.n2008 vdd.n1966 0.358259
R20324 vdd.n1966 vdd.n1964 0.358259
R20325 vdd.n1964 vdd.n1962 0.358259
R20326 vdd.n1962 vdd.n1960 0.358259
R20327 vdd.n1960 vdd.n1958 0.358259
R20328 vdd.n1958 vdd.n1956 0.358259
R20329 vdd.n1956 vdd.n1954 0.358259
R20330 vdd.n1911 vdd.n1869 0.358259
R20331 vdd.n1869 vdd.n1867 0.358259
R20332 vdd.n1867 vdd.n1865 0.358259
R20333 vdd.n1865 vdd.n1863 0.358259
R20334 vdd.n1863 vdd.n1861 0.358259
R20335 vdd.n1861 vdd.n1859 0.358259
R20336 vdd.n1859 vdd.n1857 0.358259
R20337 vdd.t94 vdd.n1023 0.340595
R20338 vdd.n2414 vdd.t112 0.340595
R20339 vdd.t107 vdd.n876 0.340595
R20340 vdd.n2935 vdd.t104 0.340595
R20341 vdd.n14 vdd.n6 0.334552
R20342 vdd.n14 vdd.n13 0.334552
R20343 vdd.n27 vdd.n19 0.21707
R20344 vdd.n27 vdd.n24 0.21707
R20345 vdd.n318 vdd.n280 0.155672
R20346 vdd.n310 vdd.n280 0.155672
R20347 vdd.n310 vdd.n309 0.155672
R20348 vdd.n309 vdd.n285 0.155672
R20349 vdd.n302 vdd.n285 0.155672
R20350 vdd.n302 vdd.n301 0.155672
R20351 vdd.n301 vdd.n289 0.155672
R20352 vdd.n294 vdd.n289 0.155672
R20353 vdd.n263 vdd.n225 0.155672
R20354 vdd.n255 vdd.n225 0.155672
R20355 vdd.n255 vdd.n254 0.155672
R20356 vdd.n254 vdd.n230 0.155672
R20357 vdd.n247 vdd.n230 0.155672
R20358 vdd.n247 vdd.n246 0.155672
R20359 vdd.n246 vdd.n234 0.155672
R20360 vdd.n239 vdd.n234 0.155672
R20361 vdd.n220 vdd.n182 0.155672
R20362 vdd.n212 vdd.n182 0.155672
R20363 vdd.n212 vdd.n211 0.155672
R20364 vdd.n211 vdd.n187 0.155672
R20365 vdd.n204 vdd.n187 0.155672
R20366 vdd.n204 vdd.n203 0.155672
R20367 vdd.n203 vdd.n191 0.155672
R20368 vdd.n196 vdd.n191 0.155672
R20369 vdd.n165 vdd.n127 0.155672
R20370 vdd.n157 vdd.n127 0.155672
R20371 vdd.n157 vdd.n156 0.155672
R20372 vdd.n156 vdd.n132 0.155672
R20373 vdd.n149 vdd.n132 0.155672
R20374 vdd.n149 vdd.n148 0.155672
R20375 vdd.n148 vdd.n136 0.155672
R20376 vdd.n141 vdd.n136 0.155672
R20377 vdd.n123 vdd.n85 0.155672
R20378 vdd.n115 vdd.n85 0.155672
R20379 vdd.n115 vdd.n114 0.155672
R20380 vdd.n114 vdd.n90 0.155672
R20381 vdd.n107 vdd.n90 0.155672
R20382 vdd.n107 vdd.n106 0.155672
R20383 vdd.n106 vdd.n94 0.155672
R20384 vdd.n99 vdd.n94 0.155672
R20385 vdd.n68 vdd.n30 0.155672
R20386 vdd.n60 vdd.n30 0.155672
R20387 vdd.n60 vdd.n59 0.155672
R20388 vdd.n59 vdd.n35 0.155672
R20389 vdd.n52 vdd.n35 0.155672
R20390 vdd.n52 vdd.n51 0.155672
R20391 vdd.n51 vdd.n39 0.155672
R20392 vdd.n44 vdd.n39 0.155672
R20393 vdd.n2049 vdd.n2011 0.155672
R20394 vdd.n2041 vdd.n2011 0.155672
R20395 vdd.n2041 vdd.n2040 0.155672
R20396 vdd.n2040 vdd.n2016 0.155672
R20397 vdd.n2033 vdd.n2016 0.155672
R20398 vdd.n2033 vdd.n2032 0.155672
R20399 vdd.n2032 vdd.n2020 0.155672
R20400 vdd.n2025 vdd.n2020 0.155672
R20401 vdd.n2104 vdd.n2066 0.155672
R20402 vdd.n2096 vdd.n2066 0.155672
R20403 vdd.n2096 vdd.n2095 0.155672
R20404 vdd.n2095 vdd.n2071 0.155672
R20405 vdd.n2088 vdd.n2071 0.155672
R20406 vdd.n2088 vdd.n2087 0.155672
R20407 vdd.n2087 vdd.n2075 0.155672
R20408 vdd.n2080 vdd.n2075 0.155672
R20409 vdd.n1951 vdd.n1913 0.155672
R20410 vdd.n1943 vdd.n1913 0.155672
R20411 vdd.n1943 vdd.n1942 0.155672
R20412 vdd.n1942 vdd.n1918 0.155672
R20413 vdd.n1935 vdd.n1918 0.155672
R20414 vdd.n1935 vdd.n1934 0.155672
R20415 vdd.n1934 vdd.n1922 0.155672
R20416 vdd.n1927 vdd.n1922 0.155672
R20417 vdd.n2006 vdd.n1968 0.155672
R20418 vdd.n1998 vdd.n1968 0.155672
R20419 vdd.n1998 vdd.n1997 0.155672
R20420 vdd.n1997 vdd.n1973 0.155672
R20421 vdd.n1990 vdd.n1973 0.155672
R20422 vdd.n1990 vdd.n1989 0.155672
R20423 vdd.n1989 vdd.n1977 0.155672
R20424 vdd.n1982 vdd.n1977 0.155672
R20425 vdd.n1854 vdd.n1816 0.155672
R20426 vdd.n1846 vdd.n1816 0.155672
R20427 vdd.n1846 vdd.n1845 0.155672
R20428 vdd.n1845 vdd.n1821 0.155672
R20429 vdd.n1838 vdd.n1821 0.155672
R20430 vdd.n1838 vdd.n1837 0.155672
R20431 vdd.n1837 vdd.n1825 0.155672
R20432 vdd.n1830 vdd.n1825 0.155672
R20433 vdd.n1909 vdd.n1871 0.155672
R20434 vdd.n1901 vdd.n1871 0.155672
R20435 vdd.n1901 vdd.n1900 0.155672
R20436 vdd.n1900 vdd.n1876 0.155672
R20437 vdd.n1893 vdd.n1876 0.155672
R20438 vdd.n1893 vdd.n1892 0.155672
R20439 vdd.n1892 vdd.n1880 0.155672
R20440 vdd.n1885 vdd.n1880 0.155672
R20441 vdd.n1099 vdd.n1091 0.152939
R20442 vdd.n1103 vdd.n1099 0.152939
R20443 vdd.n1104 vdd.n1103 0.152939
R20444 vdd.n1105 vdd.n1104 0.152939
R20445 vdd.n1106 vdd.n1105 0.152939
R20446 vdd.n1110 vdd.n1106 0.152939
R20447 vdd.n1111 vdd.n1110 0.152939
R20448 vdd.n1112 vdd.n1111 0.152939
R20449 vdd.n1113 vdd.n1112 0.152939
R20450 vdd.n1117 vdd.n1113 0.152939
R20451 vdd.n1118 vdd.n1117 0.152939
R20452 vdd.n1119 vdd.n1118 0.152939
R20453 vdd.n2262 vdd.n1119 0.152939
R20454 vdd.n2262 vdd.n2261 0.152939
R20455 vdd.n2261 vdd.n2260 0.152939
R20456 vdd.n2260 vdd.n1125 0.152939
R20457 vdd.n1130 vdd.n1125 0.152939
R20458 vdd.n1131 vdd.n1130 0.152939
R20459 vdd.n1132 vdd.n1131 0.152939
R20460 vdd.n1136 vdd.n1132 0.152939
R20461 vdd.n1137 vdd.n1136 0.152939
R20462 vdd.n1138 vdd.n1137 0.152939
R20463 vdd.n1139 vdd.n1138 0.152939
R20464 vdd.n1143 vdd.n1139 0.152939
R20465 vdd.n1144 vdd.n1143 0.152939
R20466 vdd.n1145 vdd.n1144 0.152939
R20467 vdd.n1146 vdd.n1145 0.152939
R20468 vdd.n1150 vdd.n1146 0.152939
R20469 vdd.n1151 vdd.n1150 0.152939
R20470 vdd.n1152 vdd.n1151 0.152939
R20471 vdd.n1153 vdd.n1152 0.152939
R20472 vdd.n1157 vdd.n1153 0.152939
R20473 vdd.n1158 vdd.n1157 0.152939
R20474 vdd.n1159 vdd.n1158 0.152939
R20475 vdd.n2223 vdd.n1159 0.152939
R20476 vdd.n2223 vdd.n2222 0.152939
R20477 vdd.n2222 vdd.n2221 0.152939
R20478 vdd.n2221 vdd.n1165 0.152939
R20479 vdd.n1170 vdd.n1165 0.152939
R20480 vdd.n1171 vdd.n1170 0.152939
R20481 vdd.n1172 vdd.n1171 0.152939
R20482 vdd.n1176 vdd.n1172 0.152939
R20483 vdd.n1177 vdd.n1176 0.152939
R20484 vdd.n1178 vdd.n1177 0.152939
R20485 vdd.n1179 vdd.n1178 0.152939
R20486 vdd.n1183 vdd.n1179 0.152939
R20487 vdd.n1184 vdd.n1183 0.152939
R20488 vdd.n1185 vdd.n1184 0.152939
R20489 vdd.n1186 vdd.n1185 0.152939
R20490 vdd.n1190 vdd.n1186 0.152939
R20491 vdd.n1191 vdd.n1190 0.152939
R20492 vdd.n2297 vdd.n1094 0.152939
R20493 vdd.n2111 vdd.n2110 0.152939
R20494 vdd.n2111 vdd.n1446 0.152939
R20495 vdd.n2125 vdd.n1446 0.152939
R20496 vdd.n2126 vdd.n2125 0.152939
R20497 vdd.n2127 vdd.n2126 0.152939
R20498 vdd.n2127 vdd.n1434 0.152939
R20499 vdd.n2142 vdd.n1434 0.152939
R20500 vdd.n2143 vdd.n2142 0.152939
R20501 vdd.n2144 vdd.n2143 0.152939
R20502 vdd.n2144 vdd.n1423 0.152939
R20503 vdd.n2159 vdd.n1423 0.152939
R20504 vdd.n2160 vdd.n2159 0.152939
R20505 vdd.n2161 vdd.n2160 0.152939
R20506 vdd.n2161 vdd.n1411 0.152939
R20507 vdd.n2177 vdd.n1411 0.152939
R20508 vdd.n2178 vdd.n2177 0.152939
R20509 vdd.n2179 vdd.n2178 0.152939
R20510 vdd.n670 vdd.n667 0.152939
R20511 vdd.n671 vdd.n670 0.152939
R20512 vdd.n672 vdd.n671 0.152939
R20513 vdd.n673 vdd.n672 0.152939
R20514 vdd.n676 vdd.n673 0.152939
R20515 vdd.n677 vdd.n676 0.152939
R20516 vdd.n678 vdd.n677 0.152939
R20517 vdd.n679 vdd.n678 0.152939
R20518 vdd.n682 vdd.n679 0.152939
R20519 vdd.n683 vdd.n682 0.152939
R20520 vdd.n684 vdd.n683 0.152939
R20521 vdd.n685 vdd.n684 0.152939
R20522 vdd.n690 vdd.n685 0.152939
R20523 vdd.n691 vdd.n690 0.152939
R20524 vdd.n692 vdd.n691 0.152939
R20525 vdd.n693 vdd.n692 0.152939
R20526 vdd.n696 vdd.n693 0.152939
R20527 vdd.n697 vdd.n696 0.152939
R20528 vdd.n698 vdd.n697 0.152939
R20529 vdd.n699 vdd.n698 0.152939
R20530 vdd.n702 vdd.n699 0.152939
R20531 vdd.n703 vdd.n702 0.152939
R20532 vdd.n704 vdd.n703 0.152939
R20533 vdd.n705 vdd.n704 0.152939
R20534 vdd.n708 vdd.n705 0.152939
R20535 vdd.n709 vdd.n708 0.152939
R20536 vdd.n710 vdd.n709 0.152939
R20537 vdd.n711 vdd.n710 0.152939
R20538 vdd.n714 vdd.n711 0.152939
R20539 vdd.n715 vdd.n714 0.152939
R20540 vdd.n716 vdd.n715 0.152939
R20541 vdd.n717 vdd.n716 0.152939
R20542 vdd.n720 vdd.n717 0.152939
R20543 vdd.n721 vdd.n720 0.152939
R20544 vdd.n3150 vdd.n721 0.152939
R20545 vdd.n3150 vdd.n3149 0.152939
R20546 vdd.n3149 vdd.n3148 0.152939
R20547 vdd.n3148 vdd.n725 0.152939
R20548 vdd.n730 vdd.n725 0.152939
R20549 vdd.n731 vdd.n730 0.152939
R20550 vdd.n734 vdd.n731 0.152939
R20551 vdd.n735 vdd.n734 0.152939
R20552 vdd.n736 vdd.n735 0.152939
R20553 vdd.n737 vdd.n736 0.152939
R20554 vdd.n740 vdd.n737 0.152939
R20555 vdd.n741 vdd.n740 0.152939
R20556 vdd.n742 vdd.n741 0.152939
R20557 vdd.n743 vdd.n742 0.152939
R20558 vdd.n746 vdd.n743 0.152939
R20559 vdd.n747 vdd.n746 0.152939
R20560 vdd.n748 vdd.n747 0.152939
R20561 vdd.n3233 vdd.n661 0.152939
R20562 vdd.n3234 vdd.n651 0.152939
R20563 vdd.n3248 vdd.n651 0.152939
R20564 vdd.n3249 vdd.n3248 0.152939
R20565 vdd.n3250 vdd.n3249 0.152939
R20566 vdd.n3250 vdd.n639 0.152939
R20567 vdd.n3264 vdd.n639 0.152939
R20568 vdd.n3265 vdd.n3264 0.152939
R20569 vdd.n3266 vdd.n3265 0.152939
R20570 vdd.n3266 vdd.n627 0.152939
R20571 vdd.n3281 vdd.n627 0.152939
R20572 vdd.n3282 vdd.n3281 0.152939
R20573 vdd.n3283 vdd.n3282 0.152939
R20574 vdd.n3283 vdd.n616 0.152939
R20575 vdd.n3300 vdd.n616 0.152939
R20576 vdd.n3301 vdd.n3300 0.152939
R20577 vdd.n3302 vdd.n3301 0.152939
R20578 vdd.n3302 vdd.n322 0.152939
R20579 vdd.n3382 vdd.n323 0.152939
R20580 vdd.n334 vdd.n323 0.152939
R20581 vdd.n335 vdd.n334 0.152939
R20582 vdd.n336 vdd.n335 0.152939
R20583 vdd.n343 vdd.n336 0.152939
R20584 vdd.n344 vdd.n343 0.152939
R20585 vdd.n345 vdd.n344 0.152939
R20586 vdd.n346 vdd.n345 0.152939
R20587 vdd.n354 vdd.n346 0.152939
R20588 vdd.n355 vdd.n354 0.152939
R20589 vdd.n356 vdd.n355 0.152939
R20590 vdd.n357 vdd.n356 0.152939
R20591 vdd.n365 vdd.n357 0.152939
R20592 vdd.n366 vdd.n365 0.152939
R20593 vdd.n367 vdd.n366 0.152939
R20594 vdd.n368 vdd.n367 0.152939
R20595 vdd.n443 vdd.n368 0.152939
R20596 vdd.n444 vdd.n442 0.152939
R20597 vdd.n451 vdd.n442 0.152939
R20598 vdd.n452 vdd.n451 0.152939
R20599 vdd.n453 vdd.n452 0.152939
R20600 vdd.n453 vdd.n440 0.152939
R20601 vdd.n461 vdd.n440 0.152939
R20602 vdd.n462 vdd.n461 0.152939
R20603 vdd.n463 vdd.n462 0.152939
R20604 vdd.n463 vdd.n438 0.152939
R20605 vdd.n471 vdd.n438 0.152939
R20606 vdd.n472 vdd.n471 0.152939
R20607 vdd.n473 vdd.n472 0.152939
R20608 vdd.n473 vdd.n436 0.152939
R20609 vdd.n481 vdd.n436 0.152939
R20610 vdd.n482 vdd.n481 0.152939
R20611 vdd.n483 vdd.n482 0.152939
R20612 vdd.n483 vdd.n434 0.152939
R20613 vdd.n491 vdd.n434 0.152939
R20614 vdd.n492 vdd.n491 0.152939
R20615 vdd.n493 vdd.n492 0.152939
R20616 vdd.n493 vdd.n430 0.152939
R20617 vdd.n501 vdd.n430 0.152939
R20618 vdd.n502 vdd.n501 0.152939
R20619 vdd.n503 vdd.n502 0.152939
R20620 vdd.n503 vdd.n428 0.152939
R20621 vdd.n511 vdd.n428 0.152939
R20622 vdd.n512 vdd.n511 0.152939
R20623 vdd.n513 vdd.n512 0.152939
R20624 vdd.n513 vdd.n426 0.152939
R20625 vdd.n521 vdd.n426 0.152939
R20626 vdd.n522 vdd.n521 0.152939
R20627 vdd.n523 vdd.n522 0.152939
R20628 vdd.n523 vdd.n424 0.152939
R20629 vdd.n531 vdd.n424 0.152939
R20630 vdd.n532 vdd.n531 0.152939
R20631 vdd.n533 vdd.n532 0.152939
R20632 vdd.n533 vdd.n422 0.152939
R20633 vdd.n541 vdd.n422 0.152939
R20634 vdd.n542 vdd.n541 0.152939
R20635 vdd.n543 vdd.n542 0.152939
R20636 vdd.n543 vdd.n418 0.152939
R20637 vdd.n551 vdd.n418 0.152939
R20638 vdd.n552 vdd.n551 0.152939
R20639 vdd.n553 vdd.n552 0.152939
R20640 vdd.n553 vdd.n416 0.152939
R20641 vdd.n561 vdd.n416 0.152939
R20642 vdd.n562 vdd.n561 0.152939
R20643 vdd.n563 vdd.n562 0.152939
R20644 vdd.n563 vdd.n414 0.152939
R20645 vdd.n571 vdd.n414 0.152939
R20646 vdd.n572 vdd.n571 0.152939
R20647 vdd.n573 vdd.n572 0.152939
R20648 vdd.n573 vdd.n412 0.152939
R20649 vdd.n581 vdd.n412 0.152939
R20650 vdd.n582 vdd.n581 0.152939
R20651 vdd.n583 vdd.n582 0.152939
R20652 vdd.n583 vdd.n410 0.152939
R20653 vdd.n591 vdd.n410 0.152939
R20654 vdd.n592 vdd.n591 0.152939
R20655 vdd.n593 vdd.n592 0.152939
R20656 vdd.n593 vdd.n408 0.152939
R20657 vdd.n600 vdd.n408 0.152939
R20658 vdd.n3341 vdd.n600 0.152939
R20659 vdd.n3241 vdd.n3240 0.152939
R20660 vdd.n3242 vdd.n3241 0.152939
R20661 vdd.n3242 vdd.n645 0.152939
R20662 vdd.n3256 vdd.n645 0.152939
R20663 vdd.n3257 vdd.n3256 0.152939
R20664 vdd.n3258 vdd.n3257 0.152939
R20665 vdd.n3258 vdd.n632 0.152939
R20666 vdd.n3272 vdd.n632 0.152939
R20667 vdd.n3273 vdd.n3272 0.152939
R20668 vdd.n3274 vdd.n3273 0.152939
R20669 vdd.n3274 vdd.n621 0.152939
R20670 vdd.n3289 vdd.n621 0.152939
R20671 vdd.n3290 vdd.n3289 0.152939
R20672 vdd.n3291 vdd.n3290 0.152939
R20673 vdd.n3293 vdd.n3291 0.152939
R20674 vdd.n3293 vdd.n3292 0.152939
R20675 vdd.n3292 vdd.n611 0.152939
R20676 vdd.n611 vdd.n609 0.152939
R20677 vdd.n3311 vdd.n609 0.152939
R20678 vdd.n3312 vdd.n3311 0.152939
R20679 vdd.n3313 vdd.n3312 0.152939
R20680 vdd.n3313 vdd.n607 0.152939
R20681 vdd.n3318 vdd.n607 0.152939
R20682 vdd.n3319 vdd.n3318 0.152939
R20683 vdd.n3320 vdd.n3319 0.152939
R20684 vdd.n3320 vdd.n605 0.152939
R20685 vdd.n3325 vdd.n605 0.152939
R20686 vdd.n3326 vdd.n3325 0.152939
R20687 vdd.n3327 vdd.n3326 0.152939
R20688 vdd.n3327 vdd.n603 0.152939
R20689 vdd.n3333 vdd.n603 0.152939
R20690 vdd.n3334 vdd.n3333 0.152939
R20691 vdd.n3335 vdd.n3334 0.152939
R20692 vdd.n3335 vdd.n601 0.152939
R20693 vdd.n3340 vdd.n601 0.152939
R20694 vdd.n3103 vdd.n656 0.152939
R20695 vdd.n2190 vdd.n1395 0.152939
R20696 vdd.n1741 vdd.n1740 0.152939
R20697 vdd.n1741 vdd.n1497 0.152939
R20698 vdd.n1755 vdd.n1497 0.152939
R20699 vdd.n1756 vdd.n1755 0.152939
R20700 vdd.n1757 vdd.n1756 0.152939
R20701 vdd.n1757 vdd.n1485 0.152939
R20702 vdd.n1772 vdd.n1485 0.152939
R20703 vdd.n1773 vdd.n1772 0.152939
R20704 vdd.n1774 vdd.n1773 0.152939
R20705 vdd.n1774 vdd.n1475 0.152939
R20706 vdd.n1789 vdd.n1475 0.152939
R20707 vdd.n1790 vdd.n1789 0.152939
R20708 vdd.n1791 vdd.n1790 0.152939
R20709 vdd.n1791 vdd.n1462 0.152939
R20710 vdd.n1805 vdd.n1462 0.152939
R20711 vdd.n1806 vdd.n1805 0.152939
R20712 vdd.n1807 vdd.n1806 0.152939
R20713 vdd.n1807 vdd.n1451 0.152939
R20714 vdd.n2117 vdd.n1451 0.152939
R20715 vdd.n2118 vdd.n2117 0.152939
R20716 vdd.n2119 vdd.n2118 0.152939
R20717 vdd.n2119 vdd.n1440 0.152939
R20718 vdd.n2133 vdd.n1440 0.152939
R20719 vdd.n2134 vdd.n2133 0.152939
R20720 vdd.n2135 vdd.n2134 0.152939
R20721 vdd.n2135 vdd.n1428 0.152939
R20722 vdd.n2150 vdd.n1428 0.152939
R20723 vdd.n2151 vdd.n2150 0.152939
R20724 vdd.n2152 vdd.n2151 0.152939
R20725 vdd.n2152 vdd.n1418 0.152939
R20726 vdd.n2167 vdd.n1418 0.152939
R20727 vdd.n2168 vdd.n2167 0.152939
R20728 vdd.n2171 vdd.n2168 0.152939
R20729 vdd.n2171 vdd.n2170 0.152939
R20730 vdd.n2170 vdd.n2169 0.152939
R20731 vdd.n1731 vdd.n1546 0.152939
R20732 vdd.n1731 vdd.n1730 0.152939
R20733 vdd.n1730 vdd.n1729 0.152939
R20734 vdd.n1729 vdd.n1548 0.152939
R20735 vdd.n1725 vdd.n1548 0.152939
R20736 vdd.n1725 vdd.n1724 0.152939
R20737 vdd.n1724 vdd.n1723 0.152939
R20738 vdd.n1723 vdd.n1553 0.152939
R20739 vdd.n1719 vdd.n1553 0.152939
R20740 vdd.n1719 vdd.n1718 0.152939
R20741 vdd.n1718 vdd.n1717 0.152939
R20742 vdd.n1717 vdd.n1559 0.152939
R20743 vdd.n1713 vdd.n1559 0.152939
R20744 vdd.n1713 vdd.n1712 0.152939
R20745 vdd.n1712 vdd.n1711 0.152939
R20746 vdd.n1711 vdd.n1565 0.152939
R20747 vdd.n1707 vdd.n1565 0.152939
R20748 vdd.n1707 vdd.n1706 0.152939
R20749 vdd.n1706 vdd.n1705 0.152939
R20750 vdd.n1705 vdd.n1571 0.152939
R20751 vdd.n1697 vdd.n1571 0.152939
R20752 vdd.n1697 vdd.n1696 0.152939
R20753 vdd.n1696 vdd.n1695 0.152939
R20754 vdd.n1695 vdd.n1575 0.152939
R20755 vdd.n1691 vdd.n1575 0.152939
R20756 vdd.n1691 vdd.n1690 0.152939
R20757 vdd.n1690 vdd.n1689 0.152939
R20758 vdd.n1689 vdd.n1581 0.152939
R20759 vdd.n1685 vdd.n1581 0.152939
R20760 vdd.n1685 vdd.n1684 0.152939
R20761 vdd.n1684 vdd.n1683 0.152939
R20762 vdd.n1683 vdd.n1587 0.152939
R20763 vdd.n1679 vdd.n1587 0.152939
R20764 vdd.n1679 vdd.n1678 0.152939
R20765 vdd.n1678 vdd.n1677 0.152939
R20766 vdd.n1677 vdd.n1593 0.152939
R20767 vdd.n1673 vdd.n1593 0.152939
R20768 vdd.n1673 vdd.n1672 0.152939
R20769 vdd.n1672 vdd.n1671 0.152939
R20770 vdd.n1671 vdd.n1599 0.152939
R20771 vdd.n1664 vdd.n1599 0.152939
R20772 vdd.n1664 vdd.n1663 0.152939
R20773 vdd.n1663 vdd.n1662 0.152939
R20774 vdd.n1662 vdd.n1604 0.152939
R20775 vdd.n1658 vdd.n1604 0.152939
R20776 vdd.n1658 vdd.n1657 0.152939
R20777 vdd.n1657 vdd.n1656 0.152939
R20778 vdd.n1656 vdd.n1610 0.152939
R20779 vdd.n1652 vdd.n1610 0.152939
R20780 vdd.n1652 vdd.n1651 0.152939
R20781 vdd.n1651 vdd.n1650 0.152939
R20782 vdd.n1650 vdd.n1616 0.152939
R20783 vdd.n1646 vdd.n1616 0.152939
R20784 vdd.n1646 vdd.n1645 0.152939
R20785 vdd.n1645 vdd.n1644 0.152939
R20786 vdd.n1644 vdd.n1622 0.152939
R20787 vdd.n1640 vdd.n1622 0.152939
R20788 vdd.n1640 vdd.n1639 0.152939
R20789 vdd.n1639 vdd.n1638 0.152939
R20790 vdd.n1638 vdd.n1628 0.152939
R20791 vdd.n1634 vdd.n1628 0.152939
R20792 vdd.n1634 vdd.n1509 0.152939
R20793 vdd.n1739 vdd.n1509 0.152939
R20794 vdd.n1747 vdd.n1503 0.152939
R20795 vdd.n1748 vdd.n1747 0.152939
R20796 vdd.n1749 vdd.n1748 0.152939
R20797 vdd.n1749 vdd.n1491 0.152939
R20798 vdd.n1764 vdd.n1491 0.152939
R20799 vdd.n1765 vdd.n1764 0.152939
R20800 vdd.n1766 vdd.n1765 0.152939
R20801 vdd.n1766 vdd.n1480 0.152939
R20802 vdd.n1781 vdd.n1480 0.152939
R20803 vdd.n1782 vdd.n1781 0.152939
R20804 vdd.n1783 vdd.n1782 0.152939
R20805 vdd.n1783 vdd.n1469 0.152939
R20806 vdd.n1797 vdd.n1469 0.152939
R20807 vdd.n1798 vdd.n1797 0.152939
R20808 vdd.n1799 vdd.n1798 0.152939
R20809 vdd.n1799 vdd.n1457 0.152939
R20810 vdd.n1814 vdd.n1457 0.152939
R20811 vdd.n2298 vdd.n2297 0.110256
R20812 vdd.n3034 vdd.n661 0.110256
R20813 vdd.n3103 vdd.n3102 0.110256
R20814 vdd.n2191 vdd.n2190 0.110256
R20815 vdd.n2110 vdd.n2109 0.0695946
R20816 vdd.n3383 vdd.n322 0.0695946
R20817 vdd.n3383 vdd.n3382 0.0695946
R20818 vdd.n2109 vdd.n1814 0.0695946
R20819 vdd.n2298 vdd.n1091 0.0431829
R20820 vdd.n2191 vdd.n1191 0.0431829
R20821 vdd.n3034 vdd.n667 0.0431829
R20822 vdd.n3102 vdd.n748 0.0431829
R20823 vdd vdd.n28 0.00833333
R20824 CSoutput.n19 CSoutput.t180 184.661
R20825 CSoutput.n78 CSoutput.n77 165.8
R20826 CSoutput.n76 CSoutput.n0 165.8
R20827 CSoutput.n75 CSoutput.n74 165.8
R20828 CSoutput.n73 CSoutput.n72 165.8
R20829 CSoutput.n71 CSoutput.n2 165.8
R20830 CSoutput.n69 CSoutput.n68 165.8
R20831 CSoutput.n67 CSoutput.n3 165.8
R20832 CSoutput.n66 CSoutput.n65 165.8
R20833 CSoutput.n63 CSoutput.n4 165.8
R20834 CSoutput.n61 CSoutput.n60 165.8
R20835 CSoutput.n59 CSoutput.n5 165.8
R20836 CSoutput.n58 CSoutput.n57 165.8
R20837 CSoutput.n55 CSoutput.n6 165.8
R20838 CSoutput.n54 CSoutput.n53 165.8
R20839 CSoutput.n52 CSoutput.n51 165.8
R20840 CSoutput.n50 CSoutput.n8 165.8
R20841 CSoutput.n48 CSoutput.n47 165.8
R20842 CSoutput.n46 CSoutput.n9 165.8
R20843 CSoutput.n45 CSoutput.n44 165.8
R20844 CSoutput.n42 CSoutput.n10 165.8
R20845 CSoutput.n41 CSoutput.n40 165.8
R20846 CSoutput.n39 CSoutput.n38 165.8
R20847 CSoutput.n37 CSoutput.n12 165.8
R20848 CSoutput.n35 CSoutput.n34 165.8
R20849 CSoutput.n33 CSoutput.n13 165.8
R20850 CSoutput.n32 CSoutput.n31 165.8
R20851 CSoutput.n29 CSoutput.n14 165.8
R20852 CSoutput.n28 CSoutput.n27 165.8
R20853 CSoutput.n26 CSoutput.n25 165.8
R20854 CSoutput.n24 CSoutput.n16 165.8
R20855 CSoutput.n22 CSoutput.n21 165.8
R20856 CSoutput.n20 CSoutput.n17 165.8
R20857 CSoutput.n77 CSoutput.t183 162.194
R20858 CSoutput.n18 CSoutput.t177 120.501
R20859 CSoutput.n23 CSoutput.t194 120.501
R20860 CSoutput.n15 CSoutput.t189 120.501
R20861 CSoutput.n30 CSoutput.t178 120.501
R20862 CSoutput.n36 CSoutput.t179 120.501
R20863 CSoutput.n11 CSoutput.t191 120.501
R20864 CSoutput.n43 CSoutput.t188 120.501
R20865 CSoutput.n49 CSoutput.t182 120.501
R20866 CSoutput.n7 CSoutput.t195 120.501
R20867 CSoutput.n56 CSoutput.t196 120.501
R20868 CSoutput.n62 CSoutput.t185 120.501
R20869 CSoutput.n64 CSoutput.t197 120.501
R20870 CSoutput.n70 CSoutput.t176 120.501
R20871 CSoutput.n1 CSoutput.t193 120.501
R20872 CSoutput.n310 CSoutput.n308 103.469
R20873 CSoutput.n294 CSoutput.n292 103.469
R20874 CSoutput.n279 CSoutput.n277 103.469
R20875 CSoutput.n112 CSoutput.n110 103.469
R20876 CSoutput.n96 CSoutput.n94 103.469
R20877 CSoutput.n81 CSoutput.n79 103.469
R20878 CSoutput.n320 CSoutput.n319 103.111
R20879 CSoutput.n318 CSoutput.n317 103.111
R20880 CSoutput.n316 CSoutput.n315 103.111
R20881 CSoutput.n314 CSoutput.n313 103.111
R20882 CSoutput.n312 CSoutput.n311 103.111
R20883 CSoutput.n310 CSoutput.n309 103.111
R20884 CSoutput.n306 CSoutput.n305 103.111
R20885 CSoutput.n304 CSoutput.n303 103.111
R20886 CSoutput.n302 CSoutput.n301 103.111
R20887 CSoutput.n300 CSoutput.n299 103.111
R20888 CSoutput.n298 CSoutput.n297 103.111
R20889 CSoutput.n296 CSoutput.n295 103.111
R20890 CSoutput.n294 CSoutput.n293 103.111
R20891 CSoutput.n291 CSoutput.n290 103.111
R20892 CSoutput.n289 CSoutput.n288 103.111
R20893 CSoutput.n287 CSoutput.n286 103.111
R20894 CSoutput.n285 CSoutput.n284 103.111
R20895 CSoutput.n283 CSoutput.n282 103.111
R20896 CSoutput.n281 CSoutput.n280 103.111
R20897 CSoutput.n279 CSoutput.n278 103.111
R20898 CSoutput.n112 CSoutput.n111 103.111
R20899 CSoutput.n114 CSoutput.n113 103.111
R20900 CSoutput.n116 CSoutput.n115 103.111
R20901 CSoutput.n118 CSoutput.n117 103.111
R20902 CSoutput.n120 CSoutput.n119 103.111
R20903 CSoutput.n122 CSoutput.n121 103.111
R20904 CSoutput.n124 CSoutput.n123 103.111
R20905 CSoutput.n96 CSoutput.n95 103.111
R20906 CSoutput.n98 CSoutput.n97 103.111
R20907 CSoutput.n100 CSoutput.n99 103.111
R20908 CSoutput.n102 CSoutput.n101 103.111
R20909 CSoutput.n104 CSoutput.n103 103.111
R20910 CSoutput.n106 CSoutput.n105 103.111
R20911 CSoutput.n108 CSoutput.n107 103.111
R20912 CSoutput.n81 CSoutput.n80 103.111
R20913 CSoutput.n83 CSoutput.n82 103.111
R20914 CSoutput.n85 CSoutput.n84 103.111
R20915 CSoutput.n87 CSoutput.n86 103.111
R20916 CSoutput.n89 CSoutput.n88 103.111
R20917 CSoutput.n91 CSoutput.n90 103.111
R20918 CSoutput.n93 CSoutput.n92 103.111
R20919 CSoutput.n322 CSoutput.n321 103.111
R20920 CSoutput.n346 CSoutput.n344 81.5057
R20921 CSoutput.n327 CSoutput.n325 81.5057
R20922 CSoutput.n386 CSoutput.n384 81.5057
R20923 CSoutput.n367 CSoutput.n365 81.5057
R20924 CSoutput.n362 CSoutput.n361 80.9324
R20925 CSoutput.n360 CSoutput.n359 80.9324
R20926 CSoutput.n358 CSoutput.n357 80.9324
R20927 CSoutput.n356 CSoutput.n355 80.9324
R20928 CSoutput.n354 CSoutput.n353 80.9324
R20929 CSoutput.n352 CSoutput.n351 80.9324
R20930 CSoutput.n350 CSoutput.n349 80.9324
R20931 CSoutput.n348 CSoutput.n347 80.9324
R20932 CSoutput.n346 CSoutput.n345 80.9324
R20933 CSoutput.n343 CSoutput.n342 80.9324
R20934 CSoutput.n341 CSoutput.n340 80.9324
R20935 CSoutput.n339 CSoutput.n338 80.9324
R20936 CSoutput.n337 CSoutput.n336 80.9324
R20937 CSoutput.n335 CSoutput.n334 80.9324
R20938 CSoutput.n333 CSoutput.n332 80.9324
R20939 CSoutput.n331 CSoutput.n330 80.9324
R20940 CSoutput.n329 CSoutput.n328 80.9324
R20941 CSoutput.n327 CSoutput.n326 80.9324
R20942 CSoutput.n386 CSoutput.n385 80.9324
R20943 CSoutput.n388 CSoutput.n387 80.9324
R20944 CSoutput.n390 CSoutput.n389 80.9324
R20945 CSoutput.n392 CSoutput.n391 80.9324
R20946 CSoutput.n394 CSoutput.n393 80.9324
R20947 CSoutput.n396 CSoutput.n395 80.9324
R20948 CSoutput.n398 CSoutput.n397 80.9324
R20949 CSoutput.n400 CSoutput.n399 80.9324
R20950 CSoutput.n402 CSoutput.n401 80.9324
R20951 CSoutput.n367 CSoutput.n366 80.9324
R20952 CSoutput.n369 CSoutput.n368 80.9324
R20953 CSoutput.n371 CSoutput.n370 80.9324
R20954 CSoutput.n373 CSoutput.n372 80.9324
R20955 CSoutput.n375 CSoutput.n374 80.9324
R20956 CSoutput.n377 CSoutput.n376 80.9324
R20957 CSoutput.n379 CSoutput.n378 80.9324
R20958 CSoutput.n381 CSoutput.n380 80.9324
R20959 CSoutput.n383 CSoutput.n382 80.9324
R20960 CSoutput.n25 CSoutput.n24 48.1486
R20961 CSoutput.n69 CSoutput.n3 48.1486
R20962 CSoutput.n38 CSoutput.n37 48.1486
R20963 CSoutput.n42 CSoutput.n41 48.1486
R20964 CSoutput.n51 CSoutput.n50 48.1486
R20965 CSoutput.n55 CSoutput.n54 48.1486
R20966 CSoutput.n22 CSoutput.n17 46.462
R20967 CSoutput.n72 CSoutput.n71 46.462
R20968 CSoutput.n20 CSoutput.n19 44.9055
R20969 CSoutput.n29 CSoutput.n28 43.7635
R20970 CSoutput.n65 CSoutput.n63 43.7635
R20971 CSoutput.n35 CSoutput.n13 41.7396
R20972 CSoutput.n57 CSoutput.n5 41.7396
R20973 CSoutput.n44 CSoutput.n9 37.0171
R20974 CSoutput.n48 CSoutput.n9 37.0171
R20975 CSoutput.n76 CSoutput.n75 34.9932
R20976 CSoutput.n31 CSoutput.n13 32.2947
R20977 CSoutput.n61 CSoutput.n5 32.2947
R20978 CSoutput.n30 CSoutput.n29 29.6014
R20979 CSoutput.n63 CSoutput.n62 29.6014
R20980 CSoutput.n19 CSoutput.n18 28.4085
R20981 CSoutput.n18 CSoutput.n17 25.1176
R20982 CSoutput.n72 CSoutput.n1 25.1176
R20983 CSoutput.n43 CSoutput.n42 22.0922
R20984 CSoutput.n50 CSoutput.n49 22.0922
R20985 CSoutput.n77 CSoutput.n76 21.8586
R20986 CSoutput.n37 CSoutput.n36 18.9681
R20987 CSoutput.n56 CSoutput.n55 18.9681
R20988 CSoutput.n25 CSoutput.n15 17.6292
R20989 CSoutput.n64 CSoutput.n3 17.6292
R20990 CSoutput.n24 CSoutput.n23 15.844
R20991 CSoutput.n70 CSoutput.n69 15.844
R20992 CSoutput.n38 CSoutput.n11 14.5051
R20993 CSoutput.n54 CSoutput.n7 14.5051
R20994 CSoutput.n405 CSoutput.n78 11.6139
R20995 CSoutput.n41 CSoutput.n11 11.3811
R20996 CSoutput.n51 CSoutput.n7 11.3811
R20997 CSoutput.n23 CSoutput.n22 10.0422
R20998 CSoutput.n71 CSoutput.n70 10.0422
R20999 CSoutput.n307 CSoutput.n291 9.25285
R21000 CSoutput.n109 CSoutput.n93 9.25285
R21001 CSoutput.n364 CSoutput.n324 9.09467
R21002 CSoutput.n363 CSoutput.n343 8.97993
R21003 CSoutput.n403 CSoutput.n383 8.97993
R21004 CSoutput.n28 CSoutput.n15 8.25698
R21005 CSoutput.n65 CSoutput.n64 8.25698
R21006 CSoutput.n364 CSoutput.n363 7.89345
R21007 CSoutput.n404 CSoutput.n403 7.89345
R21008 CSoutput.n324 CSoutput.n323 7.12641
R21009 CSoutput.n126 CSoutput.n125 7.12641
R21010 CSoutput.n36 CSoutput.n35 6.91809
R21011 CSoutput.n57 CSoutput.n56 6.91809
R21012 CSoutput.n405 CSoutput.n126 5.50223
R21013 CSoutput.n363 CSoutput.n362 5.25266
R21014 CSoutput.n403 CSoutput.n402 5.25266
R21015 CSoutput.n323 CSoutput.n322 5.1449
R21016 CSoutput.n307 CSoutput.n306 5.1449
R21017 CSoutput.n125 CSoutput.n124 5.1449
R21018 CSoutput.n109 CSoutput.n108 5.1449
R21019 CSoutput.n217 CSoutput.n170 4.5005
R21020 CSoutput.n186 CSoutput.n170 4.5005
R21021 CSoutput.n181 CSoutput.n165 4.5005
R21022 CSoutput.n181 CSoutput.n167 4.5005
R21023 CSoutput.n181 CSoutput.n164 4.5005
R21024 CSoutput.n181 CSoutput.n168 4.5005
R21025 CSoutput.n181 CSoutput.n163 4.5005
R21026 CSoutput.n181 CSoutput.t184 4.5005
R21027 CSoutput.n181 CSoutput.n162 4.5005
R21028 CSoutput.n181 CSoutput.n169 4.5005
R21029 CSoutput.n181 CSoutput.n170 4.5005
R21030 CSoutput.n179 CSoutput.n165 4.5005
R21031 CSoutput.n179 CSoutput.n167 4.5005
R21032 CSoutput.n179 CSoutput.n164 4.5005
R21033 CSoutput.n179 CSoutput.n168 4.5005
R21034 CSoutput.n179 CSoutput.n163 4.5005
R21035 CSoutput.n179 CSoutput.t184 4.5005
R21036 CSoutput.n179 CSoutput.n162 4.5005
R21037 CSoutput.n179 CSoutput.n169 4.5005
R21038 CSoutput.n179 CSoutput.n170 4.5005
R21039 CSoutput.n178 CSoutput.n165 4.5005
R21040 CSoutput.n178 CSoutput.n167 4.5005
R21041 CSoutput.n178 CSoutput.n164 4.5005
R21042 CSoutput.n178 CSoutput.n168 4.5005
R21043 CSoutput.n178 CSoutput.n163 4.5005
R21044 CSoutput.n178 CSoutput.t184 4.5005
R21045 CSoutput.n178 CSoutput.n162 4.5005
R21046 CSoutput.n178 CSoutput.n169 4.5005
R21047 CSoutput.n178 CSoutput.n170 4.5005
R21048 CSoutput.n263 CSoutput.n165 4.5005
R21049 CSoutput.n263 CSoutput.n167 4.5005
R21050 CSoutput.n263 CSoutput.n164 4.5005
R21051 CSoutput.n263 CSoutput.n168 4.5005
R21052 CSoutput.n263 CSoutput.n163 4.5005
R21053 CSoutput.n263 CSoutput.t184 4.5005
R21054 CSoutput.n263 CSoutput.n162 4.5005
R21055 CSoutput.n263 CSoutput.n169 4.5005
R21056 CSoutput.n263 CSoutput.n170 4.5005
R21057 CSoutput.n261 CSoutput.n165 4.5005
R21058 CSoutput.n261 CSoutput.n167 4.5005
R21059 CSoutput.n261 CSoutput.n164 4.5005
R21060 CSoutput.n261 CSoutput.n168 4.5005
R21061 CSoutput.n261 CSoutput.n163 4.5005
R21062 CSoutput.n261 CSoutput.t184 4.5005
R21063 CSoutput.n261 CSoutput.n162 4.5005
R21064 CSoutput.n261 CSoutput.n169 4.5005
R21065 CSoutput.n259 CSoutput.n165 4.5005
R21066 CSoutput.n259 CSoutput.n167 4.5005
R21067 CSoutput.n259 CSoutput.n164 4.5005
R21068 CSoutput.n259 CSoutput.n168 4.5005
R21069 CSoutput.n259 CSoutput.n163 4.5005
R21070 CSoutput.n259 CSoutput.t184 4.5005
R21071 CSoutput.n259 CSoutput.n162 4.5005
R21072 CSoutput.n259 CSoutput.n169 4.5005
R21073 CSoutput.n189 CSoutput.n165 4.5005
R21074 CSoutput.n189 CSoutput.n167 4.5005
R21075 CSoutput.n189 CSoutput.n164 4.5005
R21076 CSoutput.n189 CSoutput.n168 4.5005
R21077 CSoutput.n189 CSoutput.n163 4.5005
R21078 CSoutput.n189 CSoutput.t184 4.5005
R21079 CSoutput.n189 CSoutput.n162 4.5005
R21080 CSoutput.n189 CSoutput.n169 4.5005
R21081 CSoutput.n189 CSoutput.n170 4.5005
R21082 CSoutput.n188 CSoutput.n165 4.5005
R21083 CSoutput.n188 CSoutput.n167 4.5005
R21084 CSoutput.n188 CSoutput.n164 4.5005
R21085 CSoutput.n188 CSoutput.n168 4.5005
R21086 CSoutput.n188 CSoutput.n163 4.5005
R21087 CSoutput.n188 CSoutput.t184 4.5005
R21088 CSoutput.n188 CSoutput.n162 4.5005
R21089 CSoutput.n188 CSoutput.n169 4.5005
R21090 CSoutput.n188 CSoutput.n170 4.5005
R21091 CSoutput.n192 CSoutput.n165 4.5005
R21092 CSoutput.n192 CSoutput.n167 4.5005
R21093 CSoutput.n192 CSoutput.n164 4.5005
R21094 CSoutput.n192 CSoutput.n168 4.5005
R21095 CSoutput.n192 CSoutput.n163 4.5005
R21096 CSoutput.n192 CSoutput.t184 4.5005
R21097 CSoutput.n192 CSoutput.n162 4.5005
R21098 CSoutput.n192 CSoutput.n169 4.5005
R21099 CSoutput.n192 CSoutput.n170 4.5005
R21100 CSoutput.n191 CSoutput.n165 4.5005
R21101 CSoutput.n191 CSoutput.n167 4.5005
R21102 CSoutput.n191 CSoutput.n164 4.5005
R21103 CSoutput.n191 CSoutput.n168 4.5005
R21104 CSoutput.n191 CSoutput.n163 4.5005
R21105 CSoutput.n191 CSoutput.t184 4.5005
R21106 CSoutput.n191 CSoutput.n162 4.5005
R21107 CSoutput.n191 CSoutput.n169 4.5005
R21108 CSoutput.n191 CSoutput.n170 4.5005
R21109 CSoutput.n174 CSoutput.n165 4.5005
R21110 CSoutput.n174 CSoutput.n167 4.5005
R21111 CSoutput.n174 CSoutput.n164 4.5005
R21112 CSoutput.n174 CSoutput.n168 4.5005
R21113 CSoutput.n174 CSoutput.n163 4.5005
R21114 CSoutput.n174 CSoutput.t184 4.5005
R21115 CSoutput.n174 CSoutput.n162 4.5005
R21116 CSoutput.n174 CSoutput.n169 4.5005
R21117 CSoutput.n174 CSoutput.n170 4.5005
R21118 CSoutput.n266 CSoutput.n165 4.5005
R21119 CSoutput.n266 CSoutput.n167 4.5005
R21120 CSoutput.n266 CSoutput.n164 4.5005
R21121 CSoutput.n266 CSoutput.n168 4.5005
R21122 CSoutput.n266 CSoutput.n163 4.5005
R21123 CSoutput.n266 CSoutput.t184 4.5005
R21124 CSoutput.n266 CSoutput.n162 4.5005
R21125 CSoutput.n266 CSoutput.n169 4.5005
R21126 CSoutput.n266 CSoutput.n170 4.5005
R21127 CSoutput.n253 CSoutput.n224 4.5005
R21128 CSoutput.n253 CSoutput.n230 4.5005
R21129 CSoutput.n211 CSoutput.n200 4.5005
R21130 CSoutput.n211 CSoutput.n202 4.5005
R21131 CSoutput.n211 CSoutput.n199 4.5005
R21132 CSoutput.n211 CSoutput.n203 4.5005
R21133 CSoutput.n211 CSoutput.n198 4.5005
R21134 CSoutput.n211 CSoutput.t186 4.5005
R21135 CSoutput.n211 CSoutput.n197 4.5005
R21136 CSoutput.n211 CSoutput.n204 4.5005
R21137 CSoutput.n253 CSoutput.n211 4.5005
R21138 CSoutput.n232 CSoutput.n200 4.5005
R21139 CSoutput.n232 CSoutput.n202 4.5005
R21140 CSoutput.n232 CSoutput.n199 4.5005
R21141 CSoutput.n232 CSoutput.n203 4.5005
R21142 CSoutput.n232 CSoutput.n198 4.5005
R21143 CSoutput.n232 CSoutput.t186 4.5005
R21144 CSoutput.n232 CSoutput.n197 4.5005
R21145 CSoutput.n232 CSoutput.n204 4.5005
R21146 CSoutput.n253 CSoutput.n232 4.5005
R21147 CSoutput.n210 CSoutput.n200 4.5005
R21148 CSoutput.n210 CSoutput.n202 4.5005
R21149 CSoutput.n210 CSoutput.n199 4.5005
R21150 CSoutput.n210 CSoutput.n203 4.5005
R21151 CSoutput.n210 CSoutput.n198 4.5005
R21152 CSoutput.n210 CSoutput.t186 4.5005
R21153 CSoutput.n210 CSoutput.n197 4.5005
R21154 CSoutput.n210 CSoutput.n204 4.5005
R21155 CSoutput.n253 CSoutput.n210 4.5005
R21156 CSoutput.n234 CSoutput.n200 4.5005
R21157 CSoutput.n234 CSoutput.n202 4.5005
R21158 CSoutput.n234 CSoutput.n199 4.5005
R21159 CSoutput.n234 CSoutput.n203 4.5005
R21160 CSoutput.n234 CSoutput.n198 4.5005
R21161 CSoutput.n234 CSoutput.t186 4.5005
R21162 CSoutput.n234 CSoutput.n197 4.5005
R21163 CSoutput.n234 CSoutput.n204 4.5005
R21164 CSoutput.n253 CSoutput.n234 4.5005
R21165 CSoutput.n200 CSoutput.n195 4.5005
R21166 CSoutput.n202 CSoutput.n195 4.5005
R21167 CSoutput.n199 CSoutput.n195 4.5005
R21168 CSoutput.n203 CSoutput.n195 4.5005
R21169 CSoutput.n198 CSoutput.n195 4.5005
R21170 CSoutput.t186 CSoutput.n195 4.5005
R21171 CSoutput.n197 CSoutput.n195 4.5005
R21172 CSoutput.n204 CSoutput.n195 4.5005
R21173 CSoutput.n256 CSoutput.n200 4.5005
R21174 CSoutput.n256 CSoutput.n202 4.5005
R21175 CSoutput.n256 CSoutput.n199 4.5005
R21176 CSoutput.n256 CSoutput.n203 4.5005
R21177 CSoutput.n256 CSoutput.n198 4.5005
R21178 CSoutput.n256 CSoutput.t186 4.5005
R21179 CSoutput.n256 CSoutput.n197 4.5005
R21180 CSoutput.n256 CSoutput.n204 4.5005
R21181 CSoutput.n254 CSoutput.n200 4.5005
R21182 CSoutput.n254 CSoutput.n202 4.5005
R21183 CSoutput.n254 CSoutput.n199 4.5005
R21184 CSoutput.n254 CSoutput.n203 4.5005
R21185 CSoutput.n254 CSoutput.n198 4.5005
R21186 CSoutput.n254 CSoutput.t186 4.5005
R21187 CSoutput.n254 CSoutput.n197 4.5005
R21188 CSoutput.n254 CSoutput.n204 4.5005
R21189 CSoutput.n254 CSoutput.n253 4.5005
R21190 CSoutput.n236 CSoutput.n200 4.5005
R21191 CSoutput.n236 CSoutput.n202 4.5005
R21192 CSoutput.n236 CSoutput.n199 4.5005
R21193 CSoutput.n236 CSoutput.n203 4.5005
R21194 CSoutput.n236 CSoutput.n198 4.5005
R21195 CSoutput.n236 CSoutput.t186 4.5005
R21196 CSoutput.n236 CSoutput.n197 4.5005
R21197 CSoutput.n236 CSoutput.n204 4.5005
R21198 CSoutput.n253 CSoutput.n236 4.5005
R21199 CSoutput.n208 CSoutput.n200 4.5005
R21200 CSoutput.n208 CSoutput.n202 4.5005
R21201 CSoutput.n208 CSoutput.n199 4.5005
R21202 CSoutput.n208 CSoutput.n203 4.5005
R21203 CSoutput.n208 CSoutput.n198 4.5005
R21204 CSoutput.n208 CSoutput.t186 4.5005
R21205 CSoutput.n208 CSoutput.n197 4.5005
R21206 CSoutput.n208 CSoutput.n204 4.5005
R21207 CSoutput.n253 CSoutput.n208 4.5005
R21208 CSoutput.n238 CSoutput.n200 4.5005
R21209 CSoutput.n238 CSoutput.n202 4.5005
R21210 CSoutput.n238 CSoutput.n199 4.5005
R21211 CSoutput.n238 CSoutput.n203 4.5005
R21212 CSoutput.n238 CSoutput.n198 4.5005
R21213 CSoutput.n238 CSoutput.t186 4.5005
R21214 CSoutput.n238 CSoutput.n197 4.5005
R21215 CSoutput.n238 CSoutput.n204 4.5005
R21216 CSoutput.n253 CSoutput.n238 4.5005
R21217 CSoutput.n207 CSoutput.n200 4.5005
R21218 CSoutput.n207 CSoutput.n202 4.5005
R21219 CSoutput.n207 CSoutput.n199 4.5005
R21220 CSoutput.n207 CSoutput.n203 4.5005
R21221 CSoutput.n207 CSoutput.n198 4.5005
R21222 CSoutput.n207 CSoutput.t186 4.5005
R21223 CSoutput.n207 CSoutput.n197 4.5005
R21224 CSoutput.n207 CSoutput.n204 4.5005
R21225 CSoutput.n253 CSoutput.n207 4.5005
R21226 CSoutput.n252 CSoutput.n200 4.5005
R21227 CSoutput.n252 CSoutput.n202 4.5005
R21228 CSoutput.n252 CSoutput.n199 4.5005
R21229 CSoutput.n252 CSoutput.n203 4.5005
R21230 CSoutput.n252 CSoutput.n198 4.5005
R21231 CSoutput.n252 CSoutput.t186 4.5005
R21232 CSoutput.n252 CSoutput.n197 4.5005
R21233 CSoutput.n252 CSoutput.n204 4.5005
R21234 CSoutput.n253 CSoutput.n252 4.5005
R21235 CSoutput.n251 CSoutput.n136 4.5005
R21236 CSoutput.n152 CSoutput.n136 4.5005
R21237 CSoutput.n147 CSoutput.n131 4.5005
R21238 CSoutput.n147 CSoutput.n133 4.5005
R21239 CSoutput.n147 CSoutput.n130 4.5005
R21240 CSoutput.n147 CSoutput.n134 4.5005
R21241 CSoutput.n147 CSoutput.n129 4.5005
R21242 CSoutput.n147 CSoutput.t187 4.5005
R21243 CSoutput.n147 CSoutput.n128 4.5005
R21244 CSoutput.n147 CSoutput.n135 4.5005
R21245 CSoutput.n147 CSoutput.n136 4.5005
R21246 CSoutput.n145 CSoutput.n131 4.5005
R21247 CSoutput.n145 CSoutput.n133 4.5005
R21248 CSoutput.n145 CSoutput.n130 4.5005
R21249 CSoutput.n145 CSoutput.n134 4.5005
R21250 CSoutput.n145 CSoutput.n129 4.5005
R21251 CSoutput.n145 CSoutput.t187 4.5005
R21252 CSoutput.n145 CSoutput.n128 4.5005
R21253 CSoutput.n145 CSoutput.n135 4.5005
R21254 CSoutput.n145 CSoutput.n136 4.5005
R21255 CSoutput.n144 CSoutput.n131 4.5005
R21256 CSoutput.n144 CSoutput.n133 4.5005
R21257 CSoutput.n144 CSoutput.n130 4.5005
R21258 CSoutput.n144 CSoutput.n134 4.5005
R21259 CSoutput.n144 CSoutput.n129 4.5005
R21260 CSoutput.n144 CSoutput.t187 4.5005
R21261 CSoutput.n144 CSoutput.n128 4.5005
R21262 CSoutput.n144 CSoutput.n135 4.5005
R21263 CSoutput.n144 CSoutput.n136 4.5005
R21264 CSoutput.n273 CSoutput.n131 4.5005
R21265 CSoutput.n273 CSoutput.n133 4.5005
R21266 CSoutput.n273 CSoutput.n130 4.5005
R21267 CSoutput.n273 CSoutput.n134 4.5005
R21268 CSoutput.n273 CSoutput.n129 4.5005
R21269 CSoutput.n273 CSoutput.t187 4.5005
R21270 CSoutput.n273 CSoutput.n128 4.5005
R21271 CSoutput.n273 CSoutput.n135 4.5005
R21272 CSoutput.n273 CSoutput.n136 4.5005
R21273 CSoutput.n271 CSoutput.n131 4.5005
R21274 CSoutput.n271 CSoutput.n133 4.5005
R21275 CSoutput.n271 CSoutput.n130 4.5005
R21276 CSoutput.n271 CSoutput.n134 4.5005
R21277 CSoutput.n271 CSoutput.n129 4.5005
R21278 CSoutput.n271 CSoutput.t187 4.5005
R21279 CSoutput.n271 CSoutput.n128 4.5005
R21280 CSoutput.n271 CSoutput.n135 4.5005
R21281 CSoutput.n269 CSoutput.n131 4.5005
R21282 CSoutput.n269 CSoutput.n133 4.5005
R21283 CSoutput.n269 CSoutput.n130 4.5005
R21284 CSoutput.n269 CSoutput.n134 4.5005
R21285 CSoutput.n269 CSoutput.n129 4.5005
R21286 CSoutput.n269 CSoutput.t187 4.5005
R21287 CSoutput.n269 CSoutput.n128 4.5005
R21288 CSoutput.n269 CSoutput.n135 4.5005
R21289 CSoutput.n155 CSoutput.n131 4.5005
R21290 CSoutput.n155 CSoutput.n133 4.5005
R21291 CSoutput.n155 CSoutput.n130 4.5005
R21292 CSoutput.n155 CSoutput.n134 4.5005
R21293 CSoutput.n155 CSoutput.n129 4.5005
R21294 CSoutput.n155 CSoutput.t187 4.5005
R21295 CSoutput.n155 CSoutput.n128 4.5005
R21296 CSoutput.n155 CSoutput.n135 4.5005
R21297 CSoutput.n155 CSoutput.n136 4.5005
R21298 CSoutput.n154 CSoutput.n131 4.5005
R21299 CSoutput.n154 CSoutput.n133 4.5005
R21300 CSoutput.n154 CSoutput.n130 4.5005
R21301 CSoutput.n154 CSoutput.n134 4.5005
R21302 CSoutput.n154 CSoutput.n129 4.5005
R21303 CSoutput.n154 CSoutput.t187 4.5005
R21304 CSoutput.n154 CSoutput.n128 4.5005
R21305 CSoutput.n154 CSoutput.n135 4.5005
R21306 CSoutput.n154 CSoutput.n136 4.5005
R21307 CSoutput.n158 CSoutput.n131 4.5005
R21308 CSoutput.n158 CSoutput.n133 4.5005
R21309 CSoutput.n158 CSoutput.n130 4.5005
R21310 CSoutput.n158 CSoutput.n134 4.5005
R21311 CSoutput.n158 CSoutput.n129 4.5005
R21312 CSoutput.n158 CSoutput.t187 4.5005
R21313 CSoutput.n158 CSoutput.n128 4.5005
R21314 CSoutput.n158 CSoutput.n135 4.5005
R21315 CSoutput.n158 CSoutput.n136 4.5005
R21316 CSoutput.n157 CSoutput.n131 4.5005
R21317 CSoutput.n157 CSoutput.n133 4.5005
R21318 CSoutput.n157 CSoutput.n130 4.5005
R21319 CSoutput.n157 CSoutput.n134 4.5005
R21320 CSoutput.n157 CSoutput.n129 4.5005
R21321 CSoutput.n157 CSoutput.t187 4.5005
R21322 CSoutput.n157 CSoutput.n128 4.5005
R21323 CSoutput.n157 CSoutput.n135 4.5005
R21324 CSoutput.n157 CSoutput.n136 4.5005
R21325 CSoutput.n140 CSoutput.n131 4.5005
R21326 CSoutput.n140 CSoutput.n133 4.5005
R21327 CSoutput.n140 CSoutput.n130 4.5005
R21328 CSoutput.n140 CSoutput.n134 4.5005
R21329 CSoutput.n140 CSoutput.n129 4.5005
R21330 CSoutput.n140 CSoutput.t187 4.5005
R21331 CSoutput.n140 CSoutput.n128 4.5005
R21332 CSoutput.n140 CSoutput.n135 4.5005
R21333 CSoutput.n140 CSoutput.n136 4.5005
R21334 CSoutput.n276 CSoutput.n131 4.5005
R21335 CSoutput.n276 CSoutput.n133 4.5005
R21336 CSoutput.n276 CSoutput.n130 4.5005
R21337 CSoutput.n276 CSoutput.n134 4.5005
R21338 CSoutput.n276 CSoutput.n129 4.5005
R21339 CSoutput.n276 CSoutput.t187 4.5005
R21340 CSoutput.n276 CSoutput.n128 4.5005
R21341 CSoutput.n276 CSoutput.n135 4.5005
R21342 CSoutput.n276 CSoutput.n136 4.5005
R21343 CSoutput.n323 CSoutput.n307 4.10845
R21344 CSoutput.n125 CSoutput.n109 4.10845
R21345 CSoutput.n321 CSoutput.t118 4.06363
R21346 CSoutput.n321 CSoutput.t136 4.06363
R21347 CSoutput.n319 CSoutput.t149 4.06363
R21348 CSoutput.n319 CSoutput.t80 4.06363
R21349 CSoutput.n317 CSoutput.t84 4.06363
R21350 CSoutput.n317 CSoutput.t140 4.06363
R21351 CSoutput.n315 CSoutput.t152 4.06363
R21352 CSoutput.n315 CSoutput.t153 4.06363
R21353 CSoutput.n313 CSoutput.t100 4.06363
R21354 CSoutput.n313 CSoutput.t101 4.06363
R21355 CSoutput.n311 CSoutput.t106 4.06363
R21356 CSoutput.n311 CSoutput.t154 4.06363
R21357 CSoutput.n309 CSoutput.t72 4.06363
R21358 CSoutput.n309 CSoutput.t104 4.06363
R21359 CSoutput.n308 CSoutput.t117 4.06363
R21360 CSoutput.n308 CSoutput.t135 4.06363
R21361 CSoutput.n305 CSoutput.t107 4.06363
R21362 CSoutput.n305 CSoutput.t127 4.06363
R21363 CSoutput.n303 CSoutput.t141 4.06363
R21364 CSoutput.n303 CSoutput.t68 4.06363
R21365 CSoutput.n301 CSoutput.t69 4.06363
R21366 CSoutput.n301 CSoutput.t129 4.06363
R21367 CSoutput.n299 CSoutput.t144 4.06363
R21368 CSoutput.n299 CSoutput.t145 4.06363
R21369 CSoutput.n297 CSoutput.t88 4.06363
R21370 CSoutput.n297 CSoutput.t89 4.06363
R21371 CSoutput.n295 CSoutput.t92 4.06363
R21372 CSoutput.n295 CSoutput.t146 4.06363
R21373 CSoutput.n293 CSoutput.t61 4.06363
R21374 CSoutput.n293 CSoutput.t91 4.06363
R21375 CSoutput.n292 CSoutput.t108 4.06363
R21376 CSoutput.n292 CSoutput.t128 4.06363
R21377 CSoutput.n290 CSoutput.t134 4.06363
R21378 CSoutput.n290 CSoutput.t97 4.06363
R21379 CSoutput.n288 CSoutput.t124 4.06363
R21380 CSoutput.n288 CSoutput.t79 4.06363
R21381 CSoutput.n286 CSoutput.t142 4.06363
R21382 CSoutput.n286 CSoutput.t73 4.06363
R21383 CSoutput.n284 CSoutput.t109 4.06363
R21384 CSoutput.n284 CSoutput.t90 4.06363
R21385 CSoutput.n282 CSoutput.t93 4.06363
R21386 CSoutput.n282 CSoutput.t70 4.06363
R21387 CSoutput.n280 CSoutput.t133 4.06363
R21388 CSoutput.n280 CSoutput.t65 4.06363
R21389 CSoutput.n278 CSoutput.t102 4.06363
R21390 CSoutput.n278 CSoutput.t150 4.06363
R21391 CSoutput.n277 CSoutput.t85 4.06363
R21392 CSoutput.n277 CSoutput.t138 4.06363
R21393 CSoutput.n110 CSoutput.t76 4.06363
R21394 CSoutput.n110 CSoutput.t147 4.06363
R21395 CSoutput.n111 CSoutput.t132 4.06363
R21396 CSoutput.n111 CSoutput.t114 4.06363
R21397 CSoutput.n113 CSoutput.t99 4.06363
R21398 CSoutput.n113 CSoutput.t156 4.06363
R21399 CSoutput.n115 CSoutput.t131 4.06363
R21400 CSoutput.n115 CSoutput.t130 4.06363
R21401 CSoutput.n117 CSoutput.t120 4.06363
R21402 CSoutput.n117 CSoutput.t96 4.06363
R21403 CSoutput.n119 CSoutput.t78 4.06363
R21404 CSoutput.n119 CSoutput.t121 4.06363
R21405 CSoutput.n121 CSoutput.t119 4.06363
R21406 CSoutput.n121 CSoutput.t94 4.06363
R21407 CSoutput.n123 CSoutput.t77 4.06363
R21408 CSoutput.n123 CSoutput.t75 4.06363
R21409 CSoutput.n94 CSoutput.t63 4.06363
R21410 CSoutput.n94 CSoutput.t137 4.06363
R21411 CSoutput.n95 CSoutput.t126 4.06363
R21412 CSoutput.n95 CSoutput.t105 4.06363
R21413 CSoutput.n97 CSoutput.t87 4.06363
R21414 CSoutput.n97 CSoutput.t148 4.06363
R21415 CSoutput.n99 CSoutput.t123 4.06363
R21416 CSoutput.n99 CSoutput.t122 4.06363
R21417 CSoutput.n101 CSoutput.t112 4.06363
R21418 CSoutput.n101 CSoutput.t83 4.06363
R21419 CSoutput.n103 CSoutput.t66 4.06363
R21420 CSoutput.n103 CSoutput.t113 4.06363
R21421 CSoutput.n105 CSoutput.t111 4.06363
R21422 CSoutput.n105 CSoutput.t81 4.06363
R21423 CSoutput.n107 CSoutput.t64 4.06363
R21424 CSoutput.n107 CSoutput.t62 4.06363
R21425 CSoutput.n79 CSoutput.t139 4.06363
R21426 CSoutput.n79 CSoutput.t86 4.06363
R21427 CSoutput.n80 CSoutput.t151 4.06363
R21428 CSoutput.n80 CSoutput.t103 4.06363
R21429 CSoutput.n82 CSoutput.t67 4.06363
R21430 CSoutput.n82 CSoutput.t115 4.06363
R21431 CSoutput.n84 CSoutput.t71 4.06363
R21432 CSoutput.n84 CSoutput.t95 4.06363
R21433 CSoutput.n86 CSoutput.t155 4.06363
R21434 CSoutput.n86 CSoutput.t110 4.06363
R21435 CSoutput.n88 CSoutput.t74 4.06363
R21436 CSoutput.n88 CSoutput.t143 4.06363
R21437 CSoutput.n90 CSoutput.t82 4.06363
R21438 CSoutput.n90 CSoutput.t125 4.06363
R21439 CSoutput.n92 CSoutput.t98 4.06363
R21440 CSoutput.n92 CSoutput.t116 4.06363
R21441 CSoutput.n44 CSoutput.n43 3.79402
R21442 CSoutput.n49 CSoutput.n48 3.79402
R21443 CSoutput.n404 CSoutput.n364 3.71319
R21444 CSoutput.n405 CSoutput.n404 3.57343
R21445 CSoutput.n361 CSoutput.t51 2.82907
R21446 CSoutput.n361 CSoutput.t2 2.82907
R21447 CSoutput.n359 CSoutput.t28 2.82907
R21448 CSoutput.n359 CSoutput.t17 2.82907
R21449 CSoutput.n357 CSoutput.t6 2.82907
R21450 CSoutput.n357 CSoutput.t57 2.82907
R21451 CSoutput.n355 CSoutput.t157 2.82907
R21452 CSoutput.n355 CSoutput.t161 2.82907
R21453 CSoutput.n353 CSoutput.t31 2.82907
R21454 CSoutput.n353 CSoutput.t8 2.82907
R21455 CSoutput.n351 CSoutput.t167 2.82907
R21456 CSoutput.n351 CSoutput.t169 2.82907
R21457 CSoutput.n349 CSoutput.t50 2.82907
R21458 CSoutput.n349 CSoutput.t173 2.82907
R21459 CSoutput.n347 CSoutput.t49 2.82907
R21460 CSoutput.n347 CSoutput.t21 2.82907
R21461 CSoutput.n345 CSoutput.t58 2.82907
R21462 CSoutput.n345 CSoutput.t56 2.82907
R21463 CSoutput.n344 CSoutput.t1 2.82907
R21464 CSoutput.n344 CSoutput.t166 2.82907
R21465 CSoutput.n342 CSoutput.t12 2.82907
R21466 CSoutput.n342 CSoutput.t35 2.82907
R21467 CSoutput.n340 CSoutput.t18 2.82907
R21468 CSoutput.n340 CSoutput.t4 2.82907
R21469 CSoutput.n338 CSoutput.t53 2.82907
R21470 CSoutput.n338 CSoutput.t171 2.82907
R21471 CSoutput.n336 CSoutput.t165 2.82907
R21472 CSoutput.n336 CSoutput.t175 2.82907
R21473 CSoutput.n334 CSoutput.t29 2.82907
R21474 CSoutput.n334 CSoutput.t162 2.82907
R21475 CSoutput.n332 CSoutput.t60 2.82907
R21476 CSoutput.n332 CSoutput.t25 2.82907
R21477 CSoutput.n330 CSoutput.t11 2.82907
R21478 CSoutput.n330 CSoutput.t5 2.82907
R21479 CSoutput.n328 CSoutput.t22 2.82907
R21480 CSoutput.n328 CSoutput.t33 2.82907
R21481 CSoutput.n326 CSoutput.t13 2.82907
R21482 CSoutput.n326 CSoutput.t41 2.82907
R21483 CSoutput.n325 CSoutput.t37 2.82907
R21484 CSoutput.n325 CSoutput.t59 2.82907
R21485 CSoutput.n384 CSoutput.t34 2.82907
R21486 CSoutput.n384 CSoutput.t164 2.82907
R21487 CSoutput.n385 CSoutput.t39 2.82907
R21488 CSoutput.n385 CSoutput.t174 2.82907
R21489 CSoutput.n387 CSoutput.t7 2.82907
R21490 CSoutput.n387 CSoutput.t45 2.82907
R21491 CSoutput.n389 CSoutput.t55 2.82907
R21492 CSoutput.n389 CSoutput.t24 2.82907
R21493 CSoutput.n391 CSoutput.t47 2.82907
R21494 CSoutput.n391 CSoutput.t43 2.82907
R21495 CSoutput.n393 CSoutput.t16 2.82907
R21496 CSoutput.n393 CSoutput.t3 2.82907
R21497 CSoutput.n395 CSoutput.t27 2.82907
R21498 CSoutput.n395 CSoutput.t44 2.82907
R21499 CSoutput.n397 CSoutput.t54 2.82907
R21500 CSoutput.n397 CSoutput.t160 2.82907
R21501 CSoutput.n399 CSoutput.t42 2.82907
R21502 CSoutput.n399 CSoutput.t36 2.82907
R21503 CSoutput.n401 CSoutput.t170 2.82907
R21504 CSoutput.n401 CSoutput.t159 2.82907
R21505 CSoutput.n365 CSoutput.t168 2.82907
R21506 CSoutput.n365 CSoutput.t48 2.82907
R21507 CSoutput.n366 CSoutput.t20 2.82907
R21508 CSoutput.n366 CSoutput.t9 2.82907
R21509 CSoutput.n368 CSoutput.t23 2.82907
R21510 CSoutput.n368 CSoutput.t26 2.82907
R21511 CSoutput.n370 CSoutput.t52 2.82907
R21512 CSoutput.n370 CSoutput.t30 2.82907
R21513 CSoutput.n372 CSoutput.t10 2.82907
R21514 CSoutput.n372 CSoutput.t0 2.82907
R21515 CSoutput.n374 CSoutput.t14 2.82907
R21516 CSoutput.n374 CSoutput.t172 2.82907
R21517 CSoutput.n376 CSoutput.t32 2.82907
R21518 CSoutput.n376 CSoutput.t15 2.82907
R21519 CSoutput.n378 CSoutput.t38 2.82907
R21520 CSoutput.n378 CSoutput.t40 2.82907
R21521 CSoutput.n380 CSoutput.t19 2.82907
R21522 CSoutput.n380 CSoutput.t46 2.82907
R21523 CSoutput.n382 CSoutput.t163 2.82907
R21524 CSoutput.n382 CSoutput.t158 2.82907
R21525 CSoutput.n324 CSoutput.n126 2.57547
R21526 CSoutput.n75 CSoutput.n1 2.45513
R21527 CSoutput.n217 CSoutput.n215 2.251
R21528 CSoutput.n217 CSoutput.n214 2.251
R21529 CSoutput.n217 CSoutput.n213 2.251
R21530 CSoutput.n217 CSoutput.n212 2.251
R21531 CSoutput.n186 CSoutput.n185 2.251
R21532 CSoutput.n186 CSoutput.n184 2.251
R21533 CSoutput.n186 CSoutput.n183 2.251
R21534 CSoutput.n186 CSoutput.n182 2.251
R21535 CSoutput.n259 CSoutput.n258 2.251
R21536 CSoutput.n224 CSoutput.n222 2.251
R21537 CSoutput.n224 CSoutput.n221 2.251
R21538 CSoutput.n224 CSoutput.n220 2.251
R21539 CSoutput.n242 CSoutput.n224 2.251
R21540 CSoutput.n230 CSoutput.n229 2.251
R21541 CSoutput.n230 CSoutput.n228 2.251
R21542 CSoutput.n230 CSoutput.n227 2.251
R21543 CSoutput.n230 CSoutput.n226 2.251
R21544 CSoutput.n256 CSoutput.n196 2.251
R21545 CSoutput.n251 CSoutput.n249 2.251
R21546 CSoutput.n251 CSoutput.n248 2.251
R21547 CSoutput.n251 CSoutput.n247 2.251
R21548 CSoutput.n251 CSoutput.n246 2.251
R21549 CSoutput.n152 CSoutput.n151 2.251
R21550 CSoutput.n152 CSoutput.n150 2.251
R21551 CSoutput.n152 CSoutput.n149 2.251
R21552 CSoutput.n152 CSoutput.n148 2.251
R21553 CSoutput.n269 CSoutput.n268 2.251
R21554 CSoutput.n186 CSoutput.n166 2.2505
R21555 CSoutput.n181 CSoutput.n166 2.2505
R21556 CSoutput.n179 CSoutput.n166 2.2505
R21557 CSoutput.n178 CSoutput.n166 2.2505
R21558 CSoutput.n263 CSoutput.n166 2.2505
R21559 CSoutput.n261 CSoutput.n166 2.2505
R21560 CSoutput.n259 CSoutput.n166 2.2505
R21561 CSoutput.n189 CSoutput.n166 2.2505
R21562 CSoutput.n188 CSoutput.n166 2.2505
R21563 CSoutput.n192 CSoutput.n166 2.2505
R21564 CSoutput.n191 CSoutput.n166 2.2505
R21565 CSoutput.n174 CSoutput.n166 2.2505
R21566 CSoutput.n266 CSoutput.n166 2.2505
R21567 CSoutput.n266 CSoutput.n265 2.2505
R21568 CSoutput.n230 CSoutput.n201 2.2505
R21569 CSoutput.n211 CSoutput.n201 2.2505
R21570 CSoutput.n232 CSoutput.n201 2.2505
R21571 CSoutput.n210 CSoutput.n201 2.2505
R21572 CSoutput.n234 CSoutput.n201 2.2505
R21573 CSoutput.n201 CSoutput.n195 2.2505
R21574 CSoutput.n256 CSoutput.n201 2.2505
R21575 CSoutput.n254 CSoutput.n201 2.2505
R21576 CSoutput.n236 CSoutput.n201 2.2505
R21577 CSoutput.n208 CSoutput.n201 2.2505
R21578 CSoutput.n238 CSoutput.n201 2.2505
R21579 CSoutput.n207 CSoutput.n201 2.2505
R21580 CSoutput.n252 CSoutput.n201 2.2505
R21581 CSoutput.n252 CSoutput.n205 2.2505
R21582 CSoutput.n152 CSoutput.n132 2.2505
R21583 CSoutput.n147 CSoutput.n132 2.2505
R21584 CSoutput.n145 CSoutput.n132 2.2505
R21585 CSoutput.n144 CSoutput.n132 2.2505
R21586 CSoutput.n273 CSoutput.n132 2.2505
R21587 CSoutput.n271 CSoutput.n132 2.2505
R21588 CSoutput.n269 CSoutput.n132 2.2505
R21589 CSoutput.n155 CSoutput.n132 2.2505
R21590 CSoutput.n154 CSoutput.n132 2.2505
R21591 CSoutput.n158 CSoutput.n132 2.2505
R21592 CSoutput.n157 CSoutput.n132 2.2505
R21593 CSoutput.n140 CSoutput.n132 2.2505
R21594 CSoutput.n276 CSoutput.n132 2.2505
R21595 CSoutput.n276 CSoutput.n275 2.2505
R21596 CSoutput.n194 CSoutput.n187 2.25024
R21597 CSoutput.n194 CSoutput.n180 2.25024
R21598 CSoutput.n262 CSoutput.n194 2.25024
R21599 CSoutput.n194 CSoutput.n190 2.25024
R21600 CSoutput.n194 CSoutput.n193 2.25024
R21601 CSoutput.n194 CSoutput.n161 2.25024
R21602 CSoutput.n244 CSoutput.n241 2.25024
R21603 CSoutput.n244 CSoutput.n240 2.25024
R21604 CSoutput.n244 CSoutput.n239 2.25024
R21605 CSoutput.n244 CSoutput.n206 2.25024
R21606 CSoutput.n244 CSoutput.n243 2.25024
R21607 CSoutput.n245 CSoutput.n244 2.25024
R21608 CSoutput.n160 CSoutput.n153 2.25024
R21609 CSoutput.n160 CSoutput.n146 2.25024
R21610 CSoutput.n272 CSoutput.n160 2.25024
R21611 CSoutput.n160 CSoutput.n156 2.25024
R21612 CSoutput.n160 CSoutput.n159 2.25024
R21613 CSoutput.n160 CSoutput.n127 2.25024
R21614 CSoutput.n261 CSoutput.n171 1.50111
R21615 CSoutput.n209 CSoutput.n195 1.50111
R21616 CSoutput.n271 CSoutput.n137 1.50111
R21617 CSoutput.n217 CSoutput.n216 1.501
R21618 CSoutput.n224 CSoutput.n223 1.501
R21619 CSoutput.n251 CSoutput.n250 1.501
R21620 CSoutput.n265 CSoutput.n176 1.12536
R21621 CSoutput.n265 CSoutput.n177 1.12536
R21622 CSoutput.n265 CSoutput.n264 1.12536
R21623 CSoutput.n225 CSoutput.n205 1.12536
R21624 CSoutput.n231 CSoutput.n205 1.12536
R21625 CSoutput.n233 CSoutput.n205 1.12536
R21626 CSoutput.n275 CSoutput.n142 1.12536
R21627 CSoutput.n275 CSoutput.n143 1.12536
R21628 CSoutput.n275 CSoutput.n274 1.12536
R21629 CSoutput.n265 CSoutput.n172 1.12536
R21630 CSoutput.n265 CSoutput.n173 1.12536
R21631 CSoutput.n265 CSoutput.n175 1.12536
R21632 CSoutput.n255 CSoutput.n205 1.12536
R21633 CSoutput.n235 CSoutput.n205 1.12536
R21634 CSoutput.n237 CSoutput.n205 1.12536
R21635 CSoutput.n275 CSoutput.n138 1.12536
R21636 CSoutput.n275 CSoutput.n139 1.12536
R21637 CSoutput.n275 CSoutput.n141 1.12536
R21638 CSoutput.n31 CSoutput.n30 0.669944
R21639 CSoutput.n62 CSoutput.n61 0.669944
R21640 CSoutput.n348 CSoutput.n346 0.573776
R21641 CSoutput.n350 CSoutput.n348 0.573776
R21642 CSoutput.n352 CSoutput.n350 0.573776
R21643 CSoutput.n354 CSoutput.n352 0.573776
R21644 CSoutput.n356 CSoutput.n354 0.573776
R21645 CSoutput.n358 CSoutput.n356 0.573776
R21646 CSoutput.n360 CSoutput.n358 0.573776
R21647 CSoutput.n362 CSoutput.n360 0.573776
R21648 CSoutput.n329 CSoutput.n327 0.573776
R21649 CSoutput.n331 CSoutput.n329 0.573776
R21650 CSoutput.n333 CSoutput.n331 0.573776
R21651 CSoutput.n335 CSoutput.n333 0.573776
R21652 CSoutput.n337 CSoutput.n335 0.573776
R21653 CSoutput.n339 CSoutput.n337 0.573776
R21654 CSoutput.n341 CSoutput.n339 0.573776
R21655 CSoutput.n343 CSoutput.n341 0.573776
R21656 CSoutput.n402 CSoutput.n400 0.573776
R21657 CSoutput.n400 CSoutput.n398 0.573776
R21658 CSoutput.n398 CSoutput.n396 0.573776
R21659 CSoutput.n396 CSoutput.n394 0.573776
R21660 CSoutput.n394 CSoutput.n392 0.573776
R21661 CSoutput.n392 CSoutput.n390 0.573776
R21662 CSoutput.n390 CSoutput.n388 0.573776
R21663 CSoutput.n388 CSoutput.n386 0.573776
R21664 CSoutput.n383 CSoutput.n381 0.573776
R21665 CSoutput.n381 CSoutput.n379 0.573776
R21666 CSoutput.n379 CSoutput.n377 0.573776
R21667 CSoutput.n377 CSoutput.n375 0.573776
R21668 CSoutput.n375 CSoutput.n373 0.573776
R21669 CSoutput.n373 CSoutput.n371 0.573776
R21670 CSoutput.n371 CSoutput.n369 0.573776
R21671 CSoutput.n369 CSoutput.n367 0.573776
R21672 CSoutput.n405 CSoutput.n276 0.53442
R21673 CSoutput.n312 CSoutput.n310 0.358259
R21674 CSoutput.n314 CSoutput.n312 0.358259
R21675 CSoutput.n316 CSoutput.n314 0.358259
R21676 CSoutput.n318 CSoutput.n316 0.358259
R21677 CSoutput.n320 CSoutput.n318 0.358259
R21678 CSoutput.n322 CSoutput.n320 0.358259
R21679 CSoutput.n296 CSoutput.n294 0.358259
R21680 CSoutput.n298 CSoutput.n296 0.358259
R21681 CSoutput.n300 CSoutput.n298 0.358259
R21682 CSoutput.n302 CSoutput.n300 0.358259
R21683 CSoutput.n304 CSoutput.n302 0.358259
R21684 CSoutput.n306 CSoutput.n304 0.358259
R21685 CSoutput.n281 CSoutput.n279 0.358259
R21686 CSoutput.n283 CSoutput.n281 0.358259
R21687 CSoutput.n285 CSoutput.n283 0.358259
R21688 CSoutput.n287 CSoutput.n285 0.358259
R21689 CSoutput.n289 CSoutput.n287 0.358259
R21690 CSoutput.n291 CSoutput.n289 0.358259
R21691 CSoutput.n124 CSoutput.n122 0.358259
R21692 CSoutput.n122 CSoutput.n120 0.358259
R21693 CSoutput.n120 CSoutput.n118 0.358259
R21694 CSoutput.n118 CSoutput.n116 0.358259
R21695 CSoutput.n116 CSoutput.n114 0.358259
R21696 CSoutput.n114 CSoutput.n112 0.358259
R21697 CSoutput.n108 CSoutput.n106 0.358259
R21698 CSoutput.n106 CSoutput.n104 0.358259
R21699 CSoutput.n104 CSoutput.n102 0.358259
R21700 CSoutput.n102 CSoutput.n100 0.358259
R21701 CSoutput.n100 CSoutput.n98 0.358259
R21702 CSoutput.n98 CSoutput.n96 0.358259
R21703 CSoutput.n93 CSoutput.n91 0.358259
R21704 CSoutput.n91 CSoutput.n89 0.358259
R21705 CSoutput.n89 CSoutput.n87 0.358259
R21706 CSoutput.n87 CSoutput.n85 0.358259
R21707 CSoutput.n85 CSoutput.n83 0.358259
R21708 CSoutput.n83 CSoutput.n81 0.358259
R21709 CSoutput.n21 CSoutput.n20 0.169105
R21710 CSoutput.n21 CSoutput.n16 0.169105
R21711 CSoutput.n26 CSoutput.n16 0.169105
R21712 CSoutput.n27 CSoutput.n26 0.169105
R21713 CSoutput.n27 CSoutput.n14 0.169105
R21714 CSoutput.n32 CSoutput.n14 0.169105
R21715 CSoutput.n33 CSoutput.n32 0.169105
R21716 CSoutput.n34 CSoutput.n33 0.169105
R21717 CSoutput.n34 CSoutput.n12 0.169105
R21718 CSoutput.n39 CSoutput.n12 0.169105
R21719 CSoutput.n40 CSoutput.n39 0.169105
R21720 CSoutput.n40 CSoutput.n10 0.169105
R21721 CSoutput.n45 CSoutput.n10 0.169105
R21722 CSoutput.n46 CSoutput.n45 0.169105
R21723 CSoutput.n47 CSoutput.n46 0.169105
R21724 CSoutput.n47 CSoutput.n8 0.169105
R21725 CSoutput.n52 CSoutput.n8 0.169105
R21726 CSoutput.n53 CSoutput.n52 0.169105
R21727 CSoutput.n53 CSoutput.n6 0.169105
R21728 CSoutput.n58 CSoutput.n6 0.169105
R21729 CSoutput.n59 CSoutput.n58 0.169105
R21730 CSoutput.n60 CSoutput.n59 0.169105
R21731 CSoutput.n60 CSoutput.n4 0.169105
R21732 CSoutput.n66 CSoutput.n4 0.169105
R21733 CSoutput.n67 CSoutput.n66 0.169105
R21734 CSoutput.n68 CSoutput.n67 0.169105
R21735 CSoutput.n68 CSoutput.n2 0.169105
R21736 CSoutput.n73 CSoutput.n2 0.169105
R21737 CSoutput.n74 CSoutput.n73 0.169105
R21738 CSoutput.n74 CSoutput.n0 0.169105
R21739 CSoutput.n78 CSoutput.n0 0.169105
R21740 CSoutput.n219 CSoutput.n218 0.0910737
R21741 CSoutput.n270 CSoutput.n267 0.0723685
R21742 CSoutput.n224 CSoutput.n219 0.0522944
R21743 CSoutput.n267 CSoutput.n266 0.0499135
R21744 CSoutput.n218 CSoutput.n217 0.0499135
R21745 CSoutput.n252 CSoutput.n251 0.0464294
R21746 CSoutput.n260 CSoutput.n257 0.0391444
R21747 CSoutput.n219 CSoutput.t192 0.023435
R21748 CSoutput.n267 CSoutput.t181 0.02262
R21749 CSoutput.n218 CSoutput.t190 0.02262
R21750 CSoutput CSoutput.n405 0.0052
R21751 CSoutput.n189 CSoutput.n172 0.00365111
R21752 CSoutput.n192 CSoutput.n173 0.00365111
R21753 CSoutput.n175 CSoutput.n174 0.00365111
R21754 CSoutput.n217 CSoutput.n176 0.00365111
R21755 CSoutput.n181 CSoutput.n177 0.00365111
R21756 CSoutput.n264 CSoutput.n178 0.00365111
R21757 CSoutput.n255 CSoutput.n254 0.00365111
R21758 CSoutput.n235 CSoutput.n208 0.00365111
R21759 CSoutput.n237 CSoutput.n207 0.00365111
R21760 CSoutput.n225 CSoutput.n224 0.00365111
R21761 CSoutput.n231 CSoutput.n211 0.00365111
R21762 CSoutput.n233 CSoutput.n210 0.00365111
R21763 CSoutput.n155 CSoutput.n138 0.00365111
R21764 CSoutput.n158 CSoutput.n139 0.00365111
R21765 CSoutput.n141 CSoutput.n140 0.00365111
R21766 CSoutput.n251 CSoutput.n142 0.00365111
R21767 CSoutput.n147 CSoutput.n143 0.00365111
R21768 CSoutput.n274 CSoutput.n144 0.00365111
R21769 CSoutput.n186 CSoutput.n176 0.00340054
R21770 CSoutput.n179 CSoutput.n177 0.00340054
R21771 CSoutput.n264 CSoutput.n263 0.00340054
R21772 CSoutput.n259 CSoutput.n172 0.00340054
R21773 CSoutput.n188 CSoutput.n173 0.00340054
R21774 CSoutput.n191 CSoutput.n175 0.00340054
R21775 CSoutput.n230 CSoutput.n225 0.00340054
R21776 CSoutput.n232 CSoutput.n231 0.00340054
R21777 CSoutput.n234 CSoutput.n233 0.00340054
R21778 CSoutput.n256 CSoutput.n255 0.00340054
R21779 CSoutput.n236 CSoutput.n235 0.00340054
R21780 CSoutput.n238 CSoutput.n237 0.00340054
R21781 CSoutput.n152 CSoutput.n142 0.00340054
R21782 CSoutput.n145 CSoutput.n143 0.00340054
R21783 CSoutput.n274 CSoutput.n273 0.00340054
R21784 CSoutput.n269 CSoutput.n138 0.00340054
R21785 CSoutput.n154 CSoutput.n139 0.00340054
R21786 CSoutput.n157 CSoutput.n141 0.00340054
R21787 CSoutput.n187 CSoutput.n181 0.00252698
R21788 CSoutput.n180 CSoutput.n178 0.00252698
R21789 CSoutput.n262 CSoutput.n261 0.00252698
R21790 CSoutput.n190 CSoutput.n188 0.00252698
R21791 CSoutput.n193 CSoutput.n191 0.00252698
R21792 CSoutput.n266 CSoutput.n161 0.00252698
R21793 CSoutput.n187 CSoutput.n186 0.00252698
R21794 CSoutput.n180 CSoutput.n179 0.00252698
R21795 CSoutput.n263 CSoutput.n262 0.00252698
R21796 CSoutput.n190 CSoutput.n189 0.00252698
R21797 CSoutput.n193 CSoutput.n192 0.00252698
R21798 CSoutput.n174 CSoutput.n161 0.00252698
R21799 CSoutput.n241 CSoutput.n211 0.00252698
R21800 CSoutput.n240 CSoutput.n210 0.00252698
R21801 CSoutput.n239 CSoutput.n195 0.00252698
R21802 CSoutput.n236 CSoutput.n206 0.00252698
R21803 CSoutput.n243 CSoutput.n238 0.00252698
R21804 CSoutput.n252 CSoutput.n245 0.00252698
R21805 CSoutput.n241 CSoutput.n230 0.00252698
R21806 CSoutput.n240 CSoutput.n232 0.00252698
R21807 CSoutput.n239 CSoutput.n234 0.00252698
R21808 CSoutput.n254 CSoutput.n206 0.00252698
R21809 CSoutput.n243 CSoutput.n208 0.00252698
R21810 CSoutput.n245 CSoutput.n207 0.00252698
R21811 CSoutput.n153 CSoutput.n147 0.00252698
R21812 CSoutput.n146 CSoutput.n144 0.00252698
R21813 CSoutput.n272 CSoutput.n271 0.00252698
R21814 CSoutput.n156 CSoutput.n154 0.00252698
R21815 CSoutput.n159 CSoutput.n157 0.00252698
R21816 CSoutput.n276 CSoutput.n127 0.00252698
R21817 CSoutput.n153 CSoutput.n152 0.00252698
R21818 CSoutput.n146 CSoutput.n145 0.00252698
R21819 CSoutput.n273 CSoutput.n272 0.00252698
R21820 CSoutput.n156 CSoutput.n155 0.00252698
R21821 CSoutput.n159 CSoutput.n158 0.00252698
R21822 CSoutput.n140 CSoutput.n127 0.00252698
R21823 CSoutput.n261 CSoutput.n260 0.0020275
R21824 CSoutput.n260 CSoutput.n259 0.0020275
R21825 CSoutput.n257 CSoutput.n195 0.0020275
R21826 CSoutput.n257 CSoutput.n256 0.0020275
R21827 CSoutput.n271 CSoutput.n270 0.0020275
R21828 CSoutput.n270 CSoutput.n269 0.0020275
R21829 CSoutput.n171 CSoutput.n170 0.00166668
R21830 CSoutput.n253 CSoutput.n209 0.00166668
R21831 CSoutput.n137 CSoutput.n136 0.00166668
R21832 CSoutput.n275 CSoutput.n137 0.00133328
R21833 CSoutput.n209 CSoutput.n205 0.00133328
R21834 CSoutput.n265 CSoutput.n171 0.00133328
R21835 CSoutput.n268 CSoutput.n160 0.001
R21836 CSoutput.n246 CSoutput.n160 0.001
R21837 CSoutput.n148 CSoutput.n128 0.001
R21838 CSoutput.n247 CSoutput.n128 0.001
R21839 CSoutput.n149 CSoutput.n129 0.001
R21840 CSoutput.n248 CSoutput.n129 0.001
R21841 CSoutput.n150 CSoutput.n130 0.001
R21842 CSoutput.n249 CSoutput.n130 0.001
R21843 CSoutput.n151 CSoutput.n131 0.001
R21844 CSoutput.n250 CSoutput.n131 0.001
R21845 CSoutput.n244 CSoutput.n196 0.001
R21846 CSoutput.n244 CSoutput.n242 0.001
R21847 CSoutput.n226 CSoutput.n197 0.001
R21848 CSoutput.n220 CSoutput.n197 0.001
R21849 CSoutput.n227 CSoutput.n198 0.001
R21850 CSoutput.n221 CSoutput.n198 0.001
R21851 CSoutput.n228 CSoutput.n199 0.001
R21852 CSoutput.n222 CSoutput.n199 0.001
R21853 CSoutput.n229 CSoutput.n200 0.001
R21854 CSoutput.n223 CSoutput.n200 0.001
R21855 CSoutput.n258 CSoutput.n194 0.001
R21856 CSoutput.n212 CSoutput.n194 0.001
R21857 CSoutput.n182 CSoutput.n162 0.001
R21858 CSoutput.n213 CSoutput.n162 0.001
R21859 CSoutput.n183 CSoutput.n163 0.001
R21860 CSoutput.n214 CSoutput.n163 0.001
R21861 CSoutput.n184 CSoutput.n164 0.001
R21862 CSoutput.n215 CSoutput.n164 0.001
R21863 CSoutput.n185 CSoutput.n165 0.001
R21864 CSoutput.n216 CSoutput.n165 0.001
R21865 CSoutput.n216 CSoutput.n166 0.001
R21866 CSoutput.n215 CSoutput.n167 0.001
R21867 CSoutput.n214 CSoutput.n168 0.001
R21868 CSoutput.n213 CSoutput.t184 0.001
R21869 CSoutput.n212 CSoutput.n169 0.001
R21870 CSoutput.n185 CSoutput.n167 0.001
R21871 CSoutput.n184 CSoutput.n168 0.001
R21872 CSoutput.n183 CSoutput.t184 0.001
R21873 CSoutput.n182 CSoutput.n169 0.001
R21874 CSoutput.n258 CSoutput.n170 0.001
R21875 CSoutput.n223 CSoutput.n201 0.001
R21876 CSoutput.n222 CSoutput.n202 0.001
R21877 CSoutput.n221 CSoutput.n203 0.001
R21878 CSoutput.n220 CSoutput.t186 0.001
R21879 CSoutput.n242 CSoutput.n204 0.001
R21880 CSoutput.n229 CSoutput.n202 0.001
R21881 CSoutput.n228 CSoutput.n203 0.001
R21882 CSoutput.n227 CSoutput.t186 0.001
R21883 CSoutput.n226 CSoutput.n204 0.001
R21884 CSoutput.n253 CSoutput.n196 0.001
R21885 CSoutput.n250 CSoutput.n132 0.001
R21886 CSoutput.n249 CSoutput.n133 0.001
R21887 CSoutput.n248 CSoutput.n134 0.001
R21888 CSoutput.n247 CSoutput.t187 0.001
R21889 CSoutput.n246 CSoutput.n135 0.001
R21890 CSoutput.n151 CSoutput.n133 0.001
R21891 CSoutput.n150 CSoutput.n134 0.001
R21892 CSoutput.n149 CSoutput.t187 0.001
R21893 CSoutput.n148 CSoutput.n135 0.001
R21894 CSoutput.n268 CSoutput.n136 0.001
R21895 a_n2318_13878.n101 a_n2318_13878.t69 512.366
R21896 a_n2318_13878.n100 a_n2318_13878.t60 512.366
R21897 a_n2318_13878.n99 a_n2318_13878.t52 512.366
R21898 a_n2318_13878.n103 a_n2318_13878.t77 512.366
R21899 a_n2318_13878.n102 a_n2318_13878.t66 512.366
R21900 a_n2318_13878.n98 a_n2318_13878.t65 512.366
R21901 a_n2318_13878.n105 a_n2318_13878.t73 512.366
R21902 a_n2318_13878.n104 a_n2318_13878.t58 512.366
R21903 a_n2318_13878.n97 a_n2318_13878.t59 512.366
R21904 a_n2318_13878.n107 a_n2318_13878.t61 512.366
R21905 a_n2318_13878.n106 a_n2318_13878.t70 512.366
R21906 a_n2318_13878.n96 a_n2318_13878.t83 512.366
R21907 a_n2318_13878.n29 a_n2318_13878.t82 533.335
R21908 a_n2318_13878.n87 a_n2318_13878.t63 512.366
R21909 a_n2318_13878.n82 a_n2318_13878.t67 512.366
R21910 a_n2318_13878.n86 a_n2318_13878.t57 512.366
R21911 a_n2318_13878.n85 a_n2318_13878.t72 512.366
R21912 a_n2318_13878.n83 a_n2318_13878.t79 512.366
R21913 a_n2318_13878.n84 a_n2318_13878.t80 512.366
R21914 a_n2318_13878.n36 a_n2318_13878.t18 533.335
R21915 a_n2318_13878.n91 a_n2318_13878.t38 512.366
R21916 a_n2318_13878.n70 a_n2318_13878.t20 512.366
R21917 a_n2318_13878.n90 a_n2318_13878.t34 512.366
R21918 a_n2318_13878.n89 a_n2318_13878.t10 512.366
R21919 a_n2318_13878.n71 a_n2318_13878.t30 512.366
R21920 a_n2318_13878.n88 a_n2318_13878.t22 512.366
R21921 a_n2318_13878.n49 a_n2318_13878.t36 533.335
R21922 a_n2318_13878.n114 a_n2318_13878.t14 512.366
R21923 a_n2318_13878.n115 a_n2318_13878.t24 512.366
R21924 a_n2318_13878.n116 a_n2318_13878.t16 512.366
R21925 a_n2318_13878.n117 a_n2318_13878.t26 512.366
R21926 a_n2318_13878.n68 a_n2318_13878.t12 512.366
R21927 a_n2318_13878.n118 a_n2318_13878.t32 512.366
R21928 a_n2318_13878.n42 a_n2318_13878.t78 533.335
R21929 a_n2318_13878.n109 a_n2318_13878.t56 512.366
R21930 a_n2318_13878.n110 a_n2318_13878.t75 512.366
R21931 a_n2318_13878.n111 a_n2318_13878.t76 512.366
R21932 a_n2318_13878.n112 a_n2318_13878.t53 512.366
R21933 a_n2318_13878.n69 a_n2318_13878.t62 512.366
R21934 a_n2318_13878.n113 a_n2318_13878.t71 512.366
R21935 a_n2318_13878.n4 a_n2318_13878.n63 70.1674
R21936 a_n2318_13878.n6 a_n2318_13878.n61 70.1674
R21937 a_n2318_13878.n8 a_n2318_13878.n59 70.1674
R21938 a_n2318_13878.n10 a_n2318_13878.n57 70.1674
R21939 a_n2318_13878.n35 a_n2318_13878.n21 70.1674
R21940 a_n2318_13878.n64 a_n2318_13878.n28 70.1674
R21941 a_n2318_13878.n84 a_n2318_13878.n35 20.9683
R21942 a_n2318_13878.n22 a_n2318_13878.n33 72.3034
R21943 a_n2318_13878.n33 a_n2318_13878.n83 16.6962
R21944 a_n2318_13878.n32 a_n2318_13878.n22 77.6622
R21945 a_n2318_13878.n85 a_n2318_13878.n32 5.97853
R21946 a_n2318_13878.n31 a_n2318_13878.n20 77.6622
R21947 a_n2318_13878.n20 a_n2318_13878.n30 72.3034
R21948 a_n2318_13878.n87 a_n2318_13878.n29 20.9683
R21949 a_n2318_13878.n23 a_n2318_13878.n29 70.1674
R21950 a_n2318_13878.n88 a_n2318_13878.n64 20.9683
R21951 a_n2318_13878.n28 a_n2318_13878.n41 72.3034
R21952 a_n2318_13878.n41 a_n2318_13878.n71 16.6962
R21953 a_n2318_13878.n40 a_n2318_13878.n39 77.6622
R21954 a_n2318_13878.n89 a_n2318_13878.n40 5.97853
R21955 a_n2318_13878.n38 a_n2318_13878.n19 77.6622
R21956 a_n2318_13878.n19 a_n2318_13878.n37 72.3034
R21957 a_n2318_13878.n91 a_n2318_13878.n36 20.9683
R21958 a_n2318_13878.n18 a_n2318_13878.n36 70.1674
R21959 a_n2318_13878.n12 a_n2318_13878.n55 70.1674
R21960 a_n2318_13878.n15 a_n2318_13878.n48 70.1674
R21961 a_n2318_13878.n113 a_n2318_13878.n48 20.9683
R21962 a_n2318_13878.n47 a_n2318_13878.n16 72.3034
R21963 a_n2318_13878.n47 a_n2318_13878.n69 16.6962
R21964 a_n2318_13878.n16 a_n2318_13878.n46 77.6622
R21965 a_n2318_13878.n112 a_n2318_13878.n46 5.97853
R21966 a_n2318_13878.n45 a_n2318_13878.n17 77.6622
R21967 a_n2318_13878.n17 a_n2318_13878.n44 72.3034
R21968 a_n2318_13878.n109 a_n2318_13878.n42 20.9683
R21969 a_n2318_13878.n43 a_n2318_13878.n42 70.1674
R21970 a_n2318_13878.n118 a_n2318_13878.n55 20.9683
R21971 a_n2318_13878.n54 a_n2318_13878.n13 72.3034
R21972 a_n2318_13878.n54 a_n2318_13878.n68 16.6962
R21973 a_n2318_13878.n13 a_n2318_13878.n53 77.6622
R21974 a_n2318_13878.n117 a_n2318_13878.n53 5.97853
R21975 a_n2318_13878.n52 a_n2318_13878.n14 77.6622
R21976 a_n2318_13878.n14 a_n2318_13878.n51 72.3034
R21977 a_n2318_13878.n114 a_n2318_13878.n49 20.9683
R21978 a_n2318_13878.n50 a_n2318_13878.n49 70.1674
R21979 a_n2318_13878.n57 a_n2318_13878.n96 20.9683
R21980 a_n2318_13878.n56 a_n2318_13878.n11 75.0448
R21981 a_n2318_13878.n106 a_n2318_13878.n56 11.2134
R21982 a_n2318_13878.n11 a_n2318_13878.n107 161.3
R21983 a_n2318_13878.n59 a_n2318_13878.n97 20.9683
R21984 a_n2318_13878.n58 a_n2318_13878.n9 75.0448
R21985 a_n2318_13878.n104 a_n2318_13878.n58 11.2134
R21986 a_n2318_13878.n9 a_n2318_13878.n105 161.3
R21987 a_n2318_13878.n61 a_n2318_13878.n98 20.9683
R21988 a_n2318_13878.n60 a_n2318_13878.n7 75.0448
R21989 a_n2318_13878.n102 a_n2318_13878.n60 11.2134
R21990 a_n2318_13878.n7 a_n2318_13878.n103 161.3
R21991 a_n2318_13878.n63 a_n2318_13878.n99 20.9683
R21992 a_n2318_13878.n62 a_n2318_13878.n5 75.0448
R21993 a_n2318_13878.n100 a_n2318_13878.n62 11.2134
R21994 a_n2318_13878.n5 a_n2318_13878.n101 161.3
R21995 a_n2318_13878.n3 a_n2318_13878.n80 81.3764
R21996 a_n2318_13878.n1 a_n2318_13878.n75 81.3764
R21997 a_n2318_13878.n0 a_n2318_13878.n72 81.3764
R21998 a_n2318_13878.n3 a_n2318_13878.n81 80.9324
R21999 a_n2318_13878.n3 a_n2318_13878.n79 80.9324
R22000 a_n2318_13878.n2 a_n2318_13878.n78 80.9324
R22001 a_n2318_13878.n2 a_n2318_13878.n77 80.9324
R22002 a_n2318_13878.n1 a_n2318_13878.n76 80.9324
R22003 a_n2318_13878.n1 a_n2318_13878.n74 80.9324
R22004 a_n2318_13878.n0 a_n2318_13878.n73 80.9324
R22005 a_n2318_13878.n26 a_n2318_13878.t37 74.6477
R22006 a_n2318_13878.n24 a_n2318_13878.t29 74.6477
R22007 a_n2318_13878.n25 a_n2318_13878.t19 74.2899
R22008 a_n2318_13878.t9 a_n2318_13878.n27 74.2898
R22009 a_n2318_13878.n27 a_n2318_13878.n67 70.6783
R22010 a_n2318_13878.n26 a_n2318_13878.n66 70.6783
R22011 a_n2318_13878.n26 a_n2318_13878.n65 70.6783
R22012 a_n2318_13878.n24 a_n2318_13878.n92 70.6783
R22013 a_n2318_13878.n24 a_n2318_13878.n93 70.6783
R22014 a_n2318_13878.n25 a_n2318_13878.n94 70.6783
R22015 a_n2318_13878.n101 a_n2318_13878.n100 48.2005
R22016 a_n2318_13878.t74 a_n2318_13878.n63 533.335
R22017 a_n2318_13878.n103 a_n2318_13878.n102 48.2005
R22018 a_n2318_13878.t81 a_n2318_13878.n61 533.335
R22019 a_n2318_13878.n105 a_n2318_13878.n104 48.2005
R22020 a_n2318_13878.t68 a_n2318_13878.n59 533.335
R22021 a_n2318_13878.n107 a_n2318_13878.n106 48.2005
R22022 a_n2318_13878.t64 a_n2318_13878.n57 533.335
R22023 a_n2318_13878.n86 a_n2318_13878.n85 48.2005
R22024 a_n2318_13878.n35 a_n2318_13878.t54 533.335
R22025 a_n2318_13878.n90 a_n2318_13878.n89 48.2005
R22026 a_n2318_13878.n64 a_n2318_13878.t28 533.335
R22027 a_n2318_13878.n117 a_n2318_13878.n116 48.2005
R22028 a_n2318_13878.t8 a_n2318_13878.n55 533.335
R22029 a_n2318_13878.n112 a_n2318_13878.n111 48.2005
R22030 a_n2318_13878.t55 a_n2318_13878.n48 533.335
R22031 a_n2318_13878.n30 a_n2318_13878.n82 16.6962
R22032 a_n2318_13878.n84 a_n2318_13878.n33 27.6507
R22033 a_n2318_13878.n37 a_n2318_13878.n70 16.6962
R22034 a_n2318_13878.n88 a_n2318_13878.n41 27.6507
R22035 a_n2318_13878.n115 a_n2318_13878.n51 16.6962
R22036 a_n2318_13878.n118 a_n2318_13878.n54 27.6507
R22037 a_n2318_13878.n110 a_n2318_13878.n44 16.6962
R22038 a_n2318_13878.n113 a_n2318_13878.n47 27.6507
R22039 a_n2318_13878.n31 a_n2318_13878.n82 41.7634
R22040 a_n2318_13878.n38 a_n2318_13878.n70 41.7634
R22041 a_n2318_13878.n115 a_n2318_13878.n52 41.7634
R22042 a_n2318_13878.n110 a_n2318_13878.n45 41.7634
R22043 a_n2318_13878.n2 a_n2318_13878.n1 32.0139
R22044 a_n2318_13878.n62 a_n2318_13878.n99 35.3134
R22045 a_n2318_13878.n60 a_n2318_13878.n98 35.3134
R22046 a_n2318_13878.n58 a_n2318_13878.n97 35.3134
R22047 a_n2318_13878.n56 a_n2318_13878.n96 35.3134
R22048 a_n2318_13878.n28 a_n2318_13878.n3 23.891
R22049 a_n2318_13878.n43 a_n2318_13878.n108 12.705
R22050 a_n2318_13878.n21 a_n2318_13878.n34 12.5005
R22051 a_n2318_13878.n31 a_n2318_13878.n86 5.97853
R22052 a_n2318_13878.n32 a_n2318_13878.n83 41.7634
R22053 a_n2318_13878.n38 a_n2318_13878.n90 5.97853
R22054 a_n2318_13878.n40 a_n2318_13878.n71 41.7634
R22055 a_n2318_13878.n116 a_n2318_13878.n52 5.97853
R22056 a_n2318_13878.n68 a_n2318_13878.n53 41.7634
R22057 a_n2318_13878.n111 a_n2318_13878.n45 5.97853
R22058 a_n2318_13878.n69 a_n2318_13878.n46 41.7634
R22059 a_n2318_13878.n95 a_n2318_13878.n18 11.1956
R22060 a_n2318_13878.n87 a_n2318_13878.n30 27.6507
R22061 a_n2318_13878.n91 a_n2318_13878.n37 27.6507
R22062 a_n2318_13878.n51 a_n2318_13878.n114 27.6507
R22063 a_n2318_13878.n44 a_n2318_13878.n109 27.6507
R22064 a_n2318_13878.n27 a_n2318_13878.n119 9.85898
R22065 a_n2318_13878.n108 a_n2318_13878.n11 8.73345
R22066 a_n2318_13878.n4 a_n2318_13878.n34 8.73345
R22067 a_n2318_13878.n119 a_n2318_13878.n12 7.36035
R22068 a_n2318_13878.n95 a_n2318_13878.n25 6.01559
R22069 a_n2318_13878.n119 a_n2318_13878.n34 5.3452
R22070 a_n2318_13878.n28 a_n2318_13878.n23 4.01186
R22071 a_n2318_13878.n50 a_n2318_13878.n15 4.01186
R22072 a_n2318_13878.n67 a_n2318_13878.t13 3.61217
R22073 a_n2318_13878.n67 a_n2318_13878.t33 3.61217
R22074 a_n2318_13878.n66 a_n2318_13878.t17 3.61217
R22075 a_n2318_13878.n66 a_n2318_13878.t27 3.61217
R22076 a_n2318_13878.n65 a_n2318_13878.t15 3.61217
R22077 a_n2318_13878.n65 a_n2318_13878.t25 3.61217
R22078 a_n2318_13878.n92 a_n2318_13878.t31 3.61217
R22079 a_n2318_13878.n92 a_n2318_13878.t23 3.61217
R22080 a_n2318_13878.n93 a_n2318_13878.t35 3.61217
R22081 a_n2318_13878.n93 a_n2318_13878.t11 3.61217
R22082 a_n2318_13878.n94 a_n2318_13878.t39 3.61217
R22083 a_n2318_13878.n94 a_n2318_13878.t21 3.61217
R22084 a_n2318_13878.n80 a_n2318_13878.t3 2.82907
R22085 a_n2318_13878.n80 a_n2318_13878.t43 2.82907
R22086 a_n2318_13878.n81 a_n2318_13878.t48 2.82907
R22087 a_n2318_13878.n81 a_n2318_13878.t45 2.82907
R22088 a_n2318_13878.n79 a_n2318_13878.t49 2.82907
R22089 a_n2318_13878.n79 a_n2318_13878.t50 2.82907
R22090 a_n2318_13878.n78 a_n2318_13878.t44 2.82907
R22091 a_n2318_13878.n78 a_n2318_13878.t0 2.82907
R22092 a_n2318_13878.n77 a_n2318_13878.t42 2.82907
R22093 a_n2318_13878.n77 a_n2318_13878.t40 2.82907
R22094 a_n2318_13878.n75 a_n2318_13878.t47 2.82907
R22095 a_n2318_13878.n75 a_n2318_13878.t1 2.82907
R22096 a_n2318_13878.n76 a_n2318_13878.t4 2.82907
R22097 a_n2318_13878.n76 a_n2318_13878.t46 2.82907
R22098 a_n2318_13878.n74 a_n2318_13878.t6 2.82907
R22099 a_n2318_13878.n74 a_n2318_13878.t5 2.82907
R22100 a_n2318_13878.n73 a_n2318_13878.t41 2.82907
R22101 a_n2318_13878.n73 a_n2318_13878.t2 2.82907
R22102 a_n2318_13878.n72 a_n2318_13878.t7 2.82907
R22103 a_n2318_13878.n72 a_n2318_13878.t51 2.82907
R22104 a_n2318_13878.n3 a_n2318_13878.n2 1.3324
R22105 a_n2318_13878.n108 a_n2318_13878.n95 1.30542
R22106 a_n2318_13878.n27 a_n2318_13878.n26 1.07378
R22107 a_n2318_13878.n25 a_n2318_13878.n24 1.07378
R22108 a_n2318_13878.n8 a_n2318_13878.n7 1.04595
R22109 a_n2318_13878.n1 a_n2318_13878.n0 0.888431
R22110 a_n2318_13878.n22 a_n2318_13878.n20 0.758076
R22111 a_n2318_13878.n22 a_n2318_13878.n21 0.758076
R22112 a_n2318_13878.n39 a_n2318_13878.n19 0.758076
R22113 a_n2318_13878.n17 a_n2318_13878.n16 0.758076
R22114 a_n2318_13878.n16 a_n2318_13878.n15 0.758076
R22115 a_n2318_13878.n14 a_n2318_13878.n13 0.758076
R22116 a_n2318_13878.n13 a_n2318_13878.n12 0.758076
R22117 a_n2318_13878.n11 a_n2318_13878.n10 0.758076
R22118 a_n2318_13878.n9 a_n2318_13878.n8 0.758076
R22119 a_n2318_13878.n7 a_n2318_13878.n6 0.758076
R22120 a_n2318_13878.n5 a_n2318_13878.n4 0.758076
R22121 a_n2318_13878.n39 a_n2318_13878.n28 0.720197
R22122 a_n2318_13878.n10 a_n2318_13878.n9 0.67853
R22123 a_n2318_13878.n6 a_n2318_13878.n5 0.67853
R22124 a_n2318_13878.n50 a_n2318_13878.n14 0.568682
R22125 a_n2318_13878.n43 a_n2318_13878.n17 0.568682
R22126 a_n2318_13878.n19 a_n2318_13878.n18 0.568682
R22127 a_n2318_13878.n20 a_n2318_13878.n23 0.568682
R22128 a_n2140_13878.n21 a_n2140_13878.n20 98.9632
R22129 a_n2140_13878.n2 a_n2140_13878.n0 98.7517
R22130 a_n2140_13878.n18 a_n2140_13878.n17 98.6055
R22131 a_n2140_13878.n20 a_n2140_13878.n19 98.6055
R22132 a_n2140_13878.n6 a_n2140_13878.n5 98.6055
R22133 a_n2140_13878.n4 a_n2140_13878.n3 98.6055
R22134 a_n2140_13878.n2 a_n2140_13878.n1 98.6055
R22135 a_n2140_13878.n16 a_n2140_13878.n15 98.6054
R22136 a_n2140_13878.n8 a_n2140_13878.t17 74.6477
R22137 a_n2140_13878.n13 a_n2140_13878.t18 74.2899
R22138 a_n2140_13878.n10 a_n2140_13878.t19 74.2899
R22139 a_n2140_13878.n9 a_n2140_13878.t16 74.2899
R22140 a_n2140_13878.n12 a_n2140_13878.n11 70.6783
R22141 a_n2140_13878.n8 a_n2140_13878.n7 70.6783
R22142 a_n2140_13878.n14 a_n2140_13878.n6 14.2849
R22143 a_n2140_13878.n16 a_n2140_13878.n14 11.9339
R22144 a_n2140_13878.n14 a_n2140_13878.n13 6.95632
R22145 a_n2140_13878.n15 a_n2140_13878.t6 3.61217
R22146 a_n2140_13878.n15 a_n2140_13878.t7 3.61217
R22147 a_n2140_13878.n17 a_n2140_13878.t13 3.61217
R22148 a_n2140_13878.n17 a_n2140_13878.t14 3.61217
R22149 a_n2140_13878.n19 a_n2140_13878.t0 3.61217
R22150 a_n2140_13878.n19 a_n2140_13878.t8 3.61217
R22151 a_n2140_13878.n11 a_n2140_13878.t22 3.61217
R22152 a_n2140_13878.n11 a_n2140_13878.t23 3.61217
R22153 a_n2140_13878.n7 a_n2140_13878.t20 3.61217
R22154 a_n2140_13878.n7 a_n2140_13878.t21 3.61217
R22155 a_n2140_13878.n5 a_n2140_13878.t9 3.61217
R22156 a_n2140_13878.n5 a_n2140_13878.t1 3.61217
R22157 a_n2140_13878.n3 a_n2140_13878.t12 3.61217
R22158 a_n2140_13878.n3 a_n2140_13878.t3 3.61217
R22159 a_n2140_13878.n1 a_n2140_13878.t2 3.61217
R22160 a_n2140_13878.n1 a_n2140_13878.t4 3.61217
R22161 a_n2140_13878.n0 a_n2140_13878.t10 3.61217
R22162 a_n2140_13878.n0 a_n2140_13878.t5 3.61217
R22163 a_n2140_13878.n21 a_n2140_13878.t11 3.61217
R22164 a_n2140_13878.t15 a_n2140_13878.n21 3.61217
R22165 a_n2140_13878.n9 a_n2140_13878.n8 0.358259
R22166 a_n2140_13878.n12 a_n2140_13878.n10 0.358259
R22167 a_n2140_13878.n13 a_n2140_13878.n12 0.358259
R22168 a_n2140_13878.n20 a_n2140_13878.n18 0.358259
R22169 a_n2140_13878.n18 a_n2140_13878.n16 0.358259
R22170 a_n2140_13878.n4 a_n2140_13878.n2 0.146627
R22171 a_n2140_13878.n6 a_n2140_13878.n4 0.146627
R22172 a_n2140_13878.n10 a_n2140_13878.n9 0.101793
R22173 outputibias.n27 outputibias.n1 289.615
R22174 outputibias.n58 outputibias.n32 289.615
R22175 outputibias.n90 outputibias.n64 289.615
R22176 outputibias.n122 outputibias.n96 289.615
R22177 outputibias.n28 outputibias.n27 185
R22178 outputibias.n26 outputibias.n25 185
R22179 outputibias.n5 outputibias.n4 185
R22180 outputibias.n20 outputibias.n19 185
R22181 outputibias.n18 outputibias.n17 185
R22182 outputibias.n9 outputibias.n8 185
R22183 outputibias.n12 outputibias.n11 185
R22184 outputibias.n59 outputibias.n58 185
R22185 outputibias.n57 outputibias.n56 185
R22186 outputibias.n36 outputibias.n35 185
R22187 outputibias.n51 outputibias.n50 185
R22188 outputibias.n49 outputibias.n48 185
R22189 outputibias.n40 outputibias.n39 185
R22190 outputibias.n43 outputibias.n42 185
R22191 outputibias.n91 outputibias.n90 185
R22192 outputibias.n89 outputibias.n88 185
R22193 outputibias.n68 outputibias.n67 185
R22194 outputibias.n83 outputibias.n82 185
R22195 outputibias.n81 outputibias.n80 185
R22196 outputibias.n72 outputibias.n71 185
R22197 outputibias.n75 outputibias.n74 185
R22198 outputibias.n123 outputibias.n122 185
R22199 outputibias.n121 outputibias.n120 185
R22200 outputibias.n100 outputibias.n99 185
R22201 outputibias.n115 outputibias.n114 185
R22202 outputibias.n113 outputibias.n112 185
R22203 outputibias.n104 outputibias.n103 185
R22204 outputibias.n107 outputibias.n106 185
R22205 outputibias.n0 outputibias.t8 178.945
R22206 outputibias.n133 outputibias.t9 177.018
R22207 outputibias.n132 outputibias.t11 177.018
R22208 outputibias.n0 outputibias.t10 177.018
R22209 outputibias.t5 outputibias.n10 147.661
R22210 outputibias.t3 outputibias.n41 147.661
R22211 outputibias.t1 outputibias.n73 147.661
R22212 outputibias.t7 outputibias.n105 147.661
R22213 outputibias.n128 outputibias.t4 132.363
R22214 outputibias.n128 outputibias.t2 130.436
R22215 outputibias.n129 outputibias.t0 130.436
R22216 outputibias.n130 outputibias.t6 130.436
R22217 outputibias.n27 outputibias.n26 104.615
R22218 outputibias.n26 outputibias.n4 104.615
R22219 outputibias.n19 outputibias.n4 104.615
R22220 outputibias.n19 outputibias.n18 104.615
R22221 outputibias.n18 outputibias.n8 104.615
R22222 outputibias.n11 outputibias.n8 104.615
R22223 outputibias.n58 outputibias.n57 104.615
R22224 outputibias.n57 outputibias.n35 104.615
R22225 outputibias.n50 outputibias.n35 104.615
R22226 outputibias.n50 outputibias.n49 104.615
R22227 outputibias.n49 outputibias.n39 104.615
R22228 outputibias.n42 outputibias.n39 104.615
R22229 outputibias.n90 outputibias.n89 104.615
R22230 outputibias.n89 outputibias.n67 104.615
R22231 outputibias.n82 outputibias.n67 104.615
R22232 outputibias.n82 outputibias.n81 104.615
R22233 outputibias.n81 outputibias.n71 104.615
R22234 outputibias.n74 outputibias.n71 104.615
R22235 outputibias.n122 outputibias.n121 104.615
R22236 outputibias.n121 outputibias.n99 104.615
R22237 outputibias.n114 outputibias.n99 104.615
R22238 outputibias.n114 outputibias.n113 104.615
R22239 outputibias.n113 outputibias.n103 104.615
R22240 outputibias.n106 outputibias.n103 104.615
R22241 outputibias.n63 outputibias.n31 95.6354
R22242 outputibias.n63 outputibias.n62 94.6732
R22243 outputibias.n95 outputibias.n94 94.6732
R22244 outputibias.n127 outputibias.n126 94.6732
R22245 outputibias.n11 outputibias.t5 52.3082
R22246 outputibias.n42 outputibias.t3 52.3082
R22247 outputibias.n74 outputibias.t1 52.3082
R22248 outputibias.n106 outputibias.t7 52.3082
R22249 outputibias.n12 outputibias.n10 15.6674
R22250 outputibias.n43 outputibias.n41 15.6674
R22251 outputibias.n75 outputibias.n73 15.6674
R22252 outputibias.n107 outputibias.n105 15.6674
R22253 outputibias.n13 outputibias.n9 12.8005
R22254 outputibias.n44 outputibias.n40 12.8005
R22255 outputibias.n76 outputibias.n72 12.8005
R22256 outputibias.n108 outputibias.n104 12.8005
R22257 outputibias.n17 outputibias.n16 12.0247
R22258 outputibias.n48 outputibias.n47 12.0247
R22259 outputibias.n80 outputibias.n79 12.0247
R22260 outputibias.n112 outputibias.n111 12.0247
R22261 outputibias.n20 outputibias.n7 11.249
R22262 outputibias.n51 outputibias.n38 11.249
R22263 outputibias.n83 outputibias.n70 11.249
R22264 outputibias.n115 outputibias.n102 11.249
R22265 outputibias.n21 outputibias.n5 10.4732
R22266 outputibias.n52 outputibias.n36 10.4732
R22267 outputibias.n84 outputibias.n68 10.4732
R22268 outputibias.n116 outputibias.n100 10.4732
R22269 outputibias.n25 outputibias.n24 9.69747
R22270 outputibias.n56 outputibias.n55 9.69747
R22271 outputibias.n88 outputibias.n87 9.69747
R22272 outputibias.n120 outputibias.n119 9.69747
R22273 outputibias.n31 outputibias.n30 9.45567
R22274 outputibias.n62 outputibias.n61 9.45567
R22275 outputibias.n94 outputibias.n93 9.45567
R22276 outputibias.n126 outputibias.n125 9.45567
R22277 outputibias.n30 outputibias.n29 9.3005
R22278 outputibias.n3 outputibias.n2 9.3005
R22279 outputibias.n24 outputibias.n23 9.3005
R22280 outputibias.n22 outputibias.n21 9.3005
R22281 outputibias.n7 outputibias.n6 9.3005
R22282 outputibias.n16 outputibias.n15 9.3005
R22283 outputibias.n14 outputibias.n13 9.3005
R22284 outputibias.n61 outputibias.n60 9.3005
R22285 outputibias.n34 outputibias.n33 9.3005
R22286 outputibias.n55 outputibias.n54 9.3005
R22287 outputibias.n53 outputibias.n52 9.3005
R22288 outputibias.n38 outputibias.n37 9.3005
R22289 outputibias.n47 outputibias.n46 9.3005
R22290 outputibias.n45 outputibias.n44 9.3005
R22291 outputibias.n93 outputibias.n92 9.3005
R22292 outputibias.n66 outputibias.n65 9.3005
R22293 outputibias.n87 outputibias.n86 9.3005
R22294 outputibias.n85 outputibias.n84 9.3005
R22295 outputibias.n70 outputibias.n69 9.3005
R22296 outputibias.n79 outputibias.n78 9.3005
R22297 outputibias.n77 outputibias.n76 9.3005
R22298 outputibias.n125 outputibias.n124 9.3005
R22299 outputibias.n98 outputibias.n97 9.3005
R22300 outputibias.n119 outputibias.n118 9.3005
R22301 outputibias.n117 outputibias.n116 9.3005
R22302 outputibias.n102 outputibias.n101 9.3005
R22303 outputibias.n111 outputibias.n110 9.3005
R22304 outputibias.n109 outputibias.n108 9.3005
R22305 outputibias.n28 outputibias.n3 8.92171
R22306 outputibias.n59 outputibias.n34 8.92171
R22307 outputibias.n91 outputibias.n66 8.92171
R22308 outputibias.n123 outputibias.n98 8.92171
R22309 outputibias.n29 outputibias.n1 8.14595
R22310 outputibias.n60 outputibias.n32 8.14595
R22311 outputibias.n92 outputibias.n64 8.14595
R22312 outputibias.n124 outputibias.n96 8.14595
R22313 outputibias.n31 outputibias.n1 5.81868
R22314 outputibias.n62 outputibias.n32 5.81868
R22315 outputibias.n94 outputibias.n64 5.81868
R22316 outputibias.n126 outputibias.n96 5.81868
R22317 outputibias.n131 outputibias.n130 5.20947
R22318 outputibias.n29 outputibias.n28 5.04292
R22319 outputibias.n60 outputibias.n59 5.04292
R22320 outputibias.n92 outputibias.n91 5.04292
R22321 outputibias.n124 outputibias.n123 5.04292
R22322 outputibias.n131 outputibias.n127 4.42209
R22323 outputibias.n14 outputibias.n10 4.38594
R22324 outputibias.n45 outputibias.n41 4.38594
R22325 outputibias.n77 outputibias.n73 4.38594
R22326 outputibias.n109 outputibias.n105 4.38594
R22327 outputibias.n132 outputibias.n131 4.28454
R22328 outputibias.n25 outputibias.n3 4.26717
R22329 outputibias.n56 outputibias.n34 4.26717
R22330 outputibias.n88 outputibias.n66 4.26717
R22331 outputibias.n120 outputibias.n98 4.26717
R22332 outputibias.n24 outputibias.n5 3.49141
R22333 outputibias.n55 outputibias.n36 3.49141
R22334 outputibias.n87 outputibias.n68 3.49141
R22335 outputibias.n119 outputibias.n100 3.49141
R22336 outputibias.n21 outputibias.n20 2.71565
R22337 outputibias.n52 outputibias.n51 2.71565
R22338 outputibias.n84 outputibias.n83 2.71565
R22339 outputibias.n116 outputibias.n115 2.71565
R22340 outputibias.n17 outputibias.n7 1.93989
R22341 outputibias.n48 outputibias.n38 1.93989
R22342 outputibias.n80 outputibias.n70 1.93989
R22343 outputibias.n112 outputibias.n102 1.93989
R22344 outputibias.n130 outputibias.n129 1.9266
R22345 outputibias.n129 outputibias.n128 1.9266
R22346 outputibias.n133 outputibias.n132 1.92658
R22347 outputibias.n134 outputibias.n133 1.29913
R22348 outputibias.n16 outputibias.n9 1.16414
R22349 outputibias.n47 outputibias.n40 1.16414
R22350 outputibias.n79 outputibias.n72 1.16414
R22351 outputibias.n111 outputibias.n104 1.16414
R22352 outputibias.n127 outputibias.n95 0.962709
R22353 outputibias.n95 outputibias.n63 0.962709
R22354 outputibias.n13 outputibias.n12 0.388379
R22355 outputibias.n44 outputibias.n43 0.388379
R22356 outputibias.n76 outputibias.n75 0.388379
R22357 outputibias.n108 outputibias.n107 0.388379
R22358 outputibias.n134 outputibias.n0 0.337251
R22359 outputibias outputibias.n134 0.302375
R22360 outputibias.n30 outputibias.n2 0.155672
R22361 outputibias.n23 outputibias.n2 0.155672
R22362 outputibias.n23 outputibias.n22 0.155672
R22363 outputibias.n22 outputibias.n6 0.155672
R22364 outputibias.n15 outputibias.n6 0.155672
R22365 outputibias.n15 outputibias.n14 0.155672
R22366 outputibias.n61 outputibias.n33 0.155672
R22367 outputibias.n54 outputibias.n33 0.155672
R22368 outputibias.n54 outputibias.n53 0.155672
R22369 outputibias.n53 outputibias.n37 0.155672
R22370 outputibias.n46 outputibias.n37 0.155672
R22371 outputibias.n46 outputibias.n45 0.155672
R22372 outputibias.n93 outputibias.n65 0.155672
R22373 outputibias.n86 outputibias.n65 0.155672
R22374 outputibias.n86 outputibias.n85 0.155672
R22375 outputibias.n85 outputibias.n69 0.155672
R22376 outputibias.n78 outputibias.n69 0.155672
R22377 outputibias.n78 outputibias.n77 0.155672
R22378 outputibias.n125 outputibias.n97 0.155672
R22379 outputibias.n118 outputibias.n97 0.155672
R22380 outputibias.n118 outputibias.n117 0.155672
R22381 outputibias.n117 outputibias.n101 0.155672
R22382 outputibias.n110 outputibias.n101 0.155672
R22383 outputibias.n110 outputibias.n109 0.155672
R22384 diffpairibias.n0 diffpairibias.t27 436.822
R22385 diffpairibias.n27 diffpairibias.t24 435.479
R22386 diffpairibias.n26 diffpairibias.t21 435.479
R22387 diffpairibias.n25 diffpairibias.t22 435.479
R22388 diffpairibias.n24 diffpairibias.t26 435.479
R22389 diffpairibias.n23 diffpairibias.t20 435.479
R22390 diffpairibias.n0 diffpairibias.t23 435.479
R22391 diffpairibias.n1 diffpairibias.t28 435.479
R22392 diffpairibias.n2 diffpairibias.t25 435.479
R22393 diffpairibias.n3 diffpairibias.t29 435.479
R22394 diffpairibias.n13 diffpairibias.t14 377.536
R22395 diffpairibias.n13 diffpairibias.t0 376.193
R22396 diffpairibias.n14 diffpairibias.t10 376.193
R22397 diffpairibias.n15 diffpairibias.t12 376.193
R22398 diffpairibias.n16 diffpairibias.t6 376.193
R22399 diffpairibias.n17 diffpairibias.t2 376.193
R22400 diffpairibias.n18 diffpairibias.t16 376.193
R22401 diffpairibias.n19 diffpairibias.t4 376.193
R22402 diffpairibias.n20 diffpairibias.t18 376.193
R22403 diffpairibias.n21 diffpairibias.t8 376.193
R22404 diffpairibias.n4 diffpairibias.t15 113.368
R22405 diffpairibias.n4 diffpairibias.t1 112.698
R22406 diffpairibias.n5 diffpairibias.t11 112.698
R22407 diffpairibias.n6 diffpairibias.t13 112.698
R22408 diffpairibias.n7 diffpairibias.t7 112.698
R22409 diffpairibias.n8 diffpairibias.t3 112.698
R22410 diffpairibias.n9 diffpairibias.t17 112.698
R22411 diffpairibias.n10 diffpairibias.t5 112.698
R22412 diffpairibias.n11 diffpairibias.t19 112.698
R22413 diffpairibias.n12 diffpairibias.t9 112.698
R22414 diffpairibias.n22 diffpairibias.n21 4.77242
R22415 diffpairibias.n22 diffpairibias.n12 4.30807
R22416 diffpairibias.n23 diffpairibias.n22 4.13945
R22417 diffpairibias.n21 diffpairibias.n20 1.34352
R22418 diffpairibias.n20 diffpairibias.n19 1.34352
R22419 diffpairibias.n19 diffpairibias.n18 1.34352
R22420 diffpairibias.n18 diffpairibias.n17 1.34352
R22421 diffpairibias.n17 diffpairibias.n16 1.34352
R22422 diffpairibias.n16 diffpairibias.n15 1.34352
R22423 diffpairibias.n15 diffpairibias.n14 1.34352
R22424 diffpairibias.n14 diffpairibias.n13 1.34352
R22425 diffpairibias.n3 diffpairibias.n2 1.34352
R22426 diffpairibias.n2 diffpairibias.n1 1.34352
R22427 diffpairibias.n1 diffpairibias.n0 1.34352
R22428 diffpairibias.n24 diffpairibias.n23 1.34352
R22429 diffpairibias.n25 diffpairibias.n24 1.34352
R22430 diffpairibias.n26 diffpairibias.n25 1.34352
R22431 diffpairibias.n27 diffpairibias.n26 1.34352
R22432 diffpairibias.n28 diffpairibias.n27 0.862419
R22433 diffpairibias diffpairibias.n28 0.684875
R22434 diffpairibias.n12 diffpairibias.n11 0.672012
R22435 diffpairibias.n11 diffpairibias.n10 0.672012
R22436 diffpairibias.n10 diffpairibias.n9 0.672012
R22437 diffpairibias.n9 diffpairibias.n8 0.672012
R22438 diffpairibias.n8 diffpairibias.n7 0.672012
R22439 diffpairibias.n7 diffpairibias.n6 0.672012
R22440 diffpairibias.n6 diffpairibias.n5 0.672012
R22441 diffpairibias.n5 diffpairibias.n4 0.672012
R22442 diffpairibias.n28 diffpairibias.n3 0.190907
R22443 commonsourceibias.n281 commonsourceibias.t101 222.032
R22444 commonsourceibias.n44 commonsourceibias.t78 222.032
R22445 commonsourceibias.n166 commonsourceibias.t117 222.032
R22446 commonsourceibias.n643 commonsourceibias.t106 222.032
R22447 commonsourceibias.n413 commonsourceibias.t28 222.032
R22448 commonsourceibias.n529 commonsourceibias.t123 222.032
R22449 commonsourceibias.n364 commonsourceibias.t100 207.983
R22450 commonsourceibias.n127 commonsourceibias.t74 207.983
R22451 commonsourceibias.n249 commonsourceibias.t115 207.983
R22452 commonsourceibias.n731 commonsourceibias.t122 207.983
R22453 commonsourceibias.n501 commonsourceibias.t14 207.983
R22454 commonsourceibias.n616 commonsourceibias.t140 207.983
R22455 commonsourceibias.n280 commonsourceibias.t87 168.701
R22456 commonsourceibias.n286 commonsourceibias.t129 168.701
R22457 commonsourceibias.n292 commonsourceibias.t110 168.701
R22458 commonsourceibias.n276 commonsourceibias.t93 168.701
R22459 commonsourceibias.n300 commonsourceibias.t95 168.701
R22460 commonsourceibias.n306 commonsourceibias.t121 168.701
R22461 commonsourceibias.n271 commonsourceibias.t102 168.701
R22462 commonsourceibias.n314 commonsourceibias.t108 168.701
R22463 commonsourceibias.n320 commonsourceibias.t159 168.701
R22464 commonsourceibias.n266 commonsourceibias.t138 168.701
R22465 commonsourceibias.n328 commonsourceibias.t118 168.701
R22466 commonsourceibias.n334 commonsourceibias.t83 168.701
R22467 commonsourceibias.n261 commonsourceibias.t86 168.701
R22468 commonsourceibias.n342 commonsourceibias.t128 168.701
R22469 commonsourceibias.n348 commonsourceibias.t109 168.701
R22470 commonsourceibias.n256 commonsourceibias.t92 168.701
R22471 commonsourceibias.n356 commonsourceibias.t137 168.701
R22472 commonsourceibias.n362 commonsourceibias.t119 168.701
R22473 commonsourceibias.n125 commonsourceibias.t20 168.701
R22474 commonsourceibias.n119 commonsourceibias.t50 168.701
R22475 commonsourceibias.n19 commonsourceibias.t8 168.701
R22476 commonsourceibias.n111 commonsourceibias.t36 168.701
R22477 commonsourceibias.n105 commonsourceibias.t76 168.701
R22478 commonsourceibias.n24 commonsourceibias.t24 168.701
R22479 commonsourceibias.n97 commonsourceibias.t34 168.701
R22480 commonsourceibias.n91 commonsourceibias.t10 168.701
R22481 commonsourceibias.n29 commonsourceibias.t40 168.701
R22482 commonsourceibias.n83 commonsourceibias.t56 168.701
R22483 commonsourceibias.n77 commonsourceibias.t26 168.701
R22484 commonsourceibias.n34 commonsourceibias.t38 168.701
R22485 commonsourceibias.n69 commonsourceibias.t70 168.701
R22486 commonsourceibias.n63 commonsourceibias.t18 168.701
R22487 commonsourceibias.n39 commonsourceibias.t22 168.701
R22488 commonsourceibias.n55 commonsourceibias.t54 168.701
R22489 commonsourceibias.n49 commonsourceibias.t4 168.701
R22490 commonsourceibias.n43 commonsourceibias.t46 168.701
R22491 commonsourceibias.n247 commonsourceibias.t136 168.701
R22492 commonsourceibias.n241 commonsourceibias.t151 168.701
R22493 commonsourceibias.n5 commonsourceibias.t105 168.701
R22494 commonsourceibias.n233 commonsourceibias.t126 168.701
R22495 commonsourceibias.n227 commonsourceibias.t144 168.701
R22496 commonsourceibias.n10 commonsourceibias.t98 168.701
R22497 commonsourceibias.n219 commonsourceibias.t94 168.701
R22498 commonsourceibias.n213 commonsourceibias.t135 168.701
R22499 commonsourceibias.n150 commonsourceibias.t153 168.701
R22500 commonsourceibias.n151 commonsourceibias.t88 168.701
R22501 commonsourceibias.n153 commonsourceibias.t125 168.701
R22502 commonsourceibias.n155 commonsourceibias.t120 168.701
R22503 commonsourceibias.n191 commonsourceibias.t139 168.701
R22504 commonsourceibias.n185 commonsourceibias.t112 168.701
R22505 commonsourceibias.n161 commonsourceibias.t107 168.701
R22506 commonsourceibias.n177 commonsourceibias.t127 168.701
R22507 commonsourceibias.n171 commonsourceibias.t146 168.701
R22508 commonsourceibias.n165 commonsourceibias.t99 168.701
R22509 commonsourceibias.n642 commonsourceibias.t90 168.701
R22510 commonsourceibias.n648 commonsourceibias.t134 168.701
R22511 commonsourceibias.n654 commonsourceibias.t116 168.701
R22512 commonsourceibias.n656 commonsourceibias.t96 168.701
R22513 commonsourceibias.n663 commonsourceibias.t91 168.701
R22514 commonsourceibias.n669 commonsourceibias.t145 168.701
R22515 commonsourceibias.n671 commonsourceibias.t124 168.701
R22516 commonsourceibias.n678 commonsourceibias.t131 168.701
R22517 commonsourceibias.n684 commonsourceibias.t152 168.701
R22518 commonsourceibias.n686 commonsourceibias.t157 168.701
R22519 commonsourceibias.n693 commonsourceibias.t141 168.701
R22520 commonsourceibias.n699 commonsourceibias.t97 168.701
R22521 commonsourceibias.n701 commonsourceibias.t81 168.701
R22522 commonsourceibias.n708 commonsourceibias.t149 168.701
R22523 commonsourceibias.n714 commonsourceibias.t132 168.701
R22524 commonsourceibias.n716 commonsourceibias.t111 168.701
R22525 commonsourceibias.n723 commonsourceibias.t156 168.701
R22526 commonsourceibias.n729 commonsourceibias.t142 168.701
R22527 commonsourceibias.n412 commonsourceibias.t2 168.701
R22528 commonsourceibias.n418 commonsourceibias.t48 168.701
R22529 commonsourceibias.n424 commonsourceibias.t12 168.701
R22530 commonsourceibias.n426 commonsourceibias.t68 168.701
R22531 commonsourceibias.n433 commonsourceibias.t66 168.701
R22532 commonsourceibias.n439 commonsourceibias.t6 168.701
R22533 commonsourceibias.n441 commonsourceibias.t62 168.701
R22534 commonsourceibias.n448 commonsourceibias.t52 168.701
R22535 commonsourceibias.n454 commonsourceibias.t72 168.701
R22536 commonsourceibias.n456 commonsourceibias.t64 168.701
R22537 commonsourceibias.n463 commonsourceibias.t32 168.701
R22538 commonsourceibias.n469 commonsourceibias.t58 168.701
R22539 commonsourceibias.n471 commonsourceibias.t44 168.701
R22540 commonsourceibias.n478 commonsourceibias.t16 168.701
R22541 commonsourceibias.n484 commonsourceibias.t60 168.701
R22542 commonsourceibias.n486 commonsourceibias.t30 168.701
R22543 commonsourceibias.n493 commonsourceibias.t0 168.701
R22544 commonsourceibias.n499 commonsourceibias.t42 168.701
R22545 commonsourceibias.n614 commonsourceibias.t155 168.701
R22546 commonsourceibias.n608 commonsourceibias.t84 168.701
R22547 commonsourceibias.n601 commonsourceibias.t130 168.701
R22548 commonsourceibias.n599 commonsourceibias.t148 168.701
R22549 commonsourceibias.n593 commonsourceibias.t80 168.701
R22550 commonsourceibias.n586 commonsourceibias.t89 168.701
R22551 commonsourceibias.n584 commonsourceibias.t113 168.701
R22552 commonsourceibias.n578 commonsourceibias.t154 168.701
R22553 commonsourceibias.n571 commonsourceibias.t85 168.701
R22554 commonsourceibias.n528 commonsourceibias.t103 168.701
R22555 commonsourceibias.n534 commonsourceibias.t150 168.701
R22556 commonsourceibias.n540 commonsourceibias.t133 168.701
R22557 commonsourceibias.n542 commonsourceibias.t114 168.701
R22558 commonsourceibias.n549 commonsourceibias.t104 168.701
R22559 commonsourceibias.n555 commonsourceibias.t158 168.701
R22560 commonsourceibias.n519 commonsourceibias.t143 168.701
R22561 commonsourceibias.n517 commonsourceibias.t147 168.701
R22562 commonsourceibias.n515 commonsourceibias.t82 168.701
R22563 commonsourceibias.n363 commonsourceibias.n251 161.3
R22564 commonsourceibias.n361 commonsourceibias.n360 161.3
R22565 commonsourceibias.n359 commonsourceibias.n252 161.3
R22566 commonsourceibias.n358 commonsourceibias.n357 161.3
R22567 commonsourceibias.n355 commonsourceibias.n253 161.3
R22568 commonsourceibias.n354 commonsourceibias.n353 161.3
R22569 commonsourceibias.n352 commonsourceibias.n254 161.3
R22570 commonsourceibias.n351 commonsourceibias.n350 161.3
R22571 commonsourceibias.n349 commonsourceibias.n255 161.3
R22572 commonsourceibias.n347 commonsourceibias.n346 161.3
R22573 commonsourceibias.n345 commonsourceibias.n257 161.3
R22574 commonsourceibias.n344 commonsourceibias.n343 161.3
R22575 commonsourceibias.n341 commonsourceibias.n258 161.3
R22576 commonsourceibias.n340 commonsourceibias.n339 161.3
R22577 commonsourceibias.n338 commonsourceibias.n259 161.3
R22578 commonsourceibias.n337 commonsourceibias.n336 161.3
R22579 commonsourceibias.n335 commonsourceibias.n260 161.3
R22580 commonsourceibias.n333 commonsourceibias.n332 161.3
R22581 commonsourceibias.n331 commonsourceibias.n262 161.3
R22582 commonsourceibias.n330 commonsourceibias.n329 161.3
R22583 commonsourceibias.n327 commonsourceibias.n263 161.3
R22584 commonsourceibias.n326 commonsourceibias.n325 161.3
R22585 commonsourceibias.n324 commonsourceibias.n264 161.3
R22586 commonsourceibias.n323 commonsourceibias.n322 161.3
R22587 commonsourceibias.n321 commonsourceibias.n265 161.3
R22588 commonsourceibias.n319 commonsourceibias.n318 161.3
R22589 commonsourceibias.n317 commonsourceibias.n267 161.3
R22590 commonsourceibias.n316 commonsourceibias.n315 161.3
R22591 commonsourceibias.n313 commonsourceibias.n268 161.3
R22592 commonsourceibias.n312 commonsourceibias.n311 161.3
R22593 commonsourceibias.n310 commonsourceibias.n269 161.3
R22594 commonsourceibias.n309 commonsourceibias.n308 161.3
R22595 commonsourceibias.n307 commonsourceibias.n270 161.3
R22596 commonsourceibias.n305 commonsourceibias.n304 161.3
R22597 commonsourceibias.n303 commonsourceibias.n272 161.3
R22598 commonsourceibias.n302 commonsourceibias.n301 161.3
R22599 commonsourceibias.n299 commonsourceibias.n273 161.3
R22600 commonsourceibias.n298 commonsourceibias.n297 161.3
R22601 commonsourceibias.n296 commonsourceibias.n274 161.3
R22602 commonsourceibias.n295 commonsourceibias.n294 161.3
R22603 commonsourceibias.n293 commonsourceibias.n275 161.3
R22604 commonsourceibias.n291 commonsourceibias.n290 161.3
R22605 commonsourceibias.n289 commonsourceibias.n277 161.3
R22606 commonsourceibias.n288 commonsourceibias.n287 161.3
R22607 commonsourceibias.n285 commonsourceibias.n278 161.3
R22608 commonsourceibias.n284 commonsourceibias.n283 161.3
R22609 commonsourceibias.n282 commonsourceibias.n279 161.3
R22610 commonsourceibias.n45 commonsourceibias.n42 161.3
R22611 commonsourceibias.n47 commonsourceibias.n46 161.3
R22612 commonsourceibias.n48 commonsourceibias.n41 161.3
R22613 commonsourceibias.n51 commonsourceibias.n50 161.3
R22614 commonsourceibias.n52 commonsourceibias.n40 161.3
R22615 commonsourceibias.n54 commonsourceibias.n53 161.3
R22616 commonsourceibias.n56 commonsourceibias.n38 161.3
R22617 commonsourceibias.n58 commonsourceibias.n57 161.3
R22618 commonsourceibias.n59 commonsourceibias.n37 161.3
R22619 commonsourceibias.n61 commonsourceibias.n60 161.3
R22620 commonsourceibias.n62 commonsourceibias.n36 161.3
R22621 commonsourceibias.n65 commonsourceibias.n64 161.3
R22622 commonsourceibias.n66 commonsourceibias.n35 161.3
R22623 commonsourceibias.n68 commonsourceibias.n67 161.3
R22624 commonsourceibias.n70 commonsourceibias.n33 161.3
R22625 commonsourceibias.n72 commonsourceibias.n71 161.3
R22626 commonsourceibias.n73 commonsourceibias.n32 161.3
R22627 commonsourceibias.n75 commonsourceibias.n74 161.3
R22628 commonsourceibias.n76 commonsourceibias.n31 161.3
R22629 commonsourceibias.n79 commonsourceibias.n78 161.3
R22630 commonsourceibias.n80 commonsourceibias.n30 161.3
R22631 commonsourceibias.n82 commonsourceibias.n81 161.3
R22632 commonsourceibias.n84 commonsourceibias.n28 161.3
R22633 commonsourceibias.n86 commonsourceibias.n85 161.3
R22634 commonsourceibias.n87 commonsourceibias.n27 161.3
R22635 commonsourceibias.n89 commonsourceibias.n88 161.3
R22636 commonsourceibias.n90 commonsourceibias.n26 161.3
R22637 commonsourceibias.n93 commonsourceibias.n92 161.3
R22638 commonsourceibias.n94 commonsourceibias.n25 161.3
R22639 commonsourceibias.n96 commonsourceibias.n95 161.3
R22640 commonsourceibias.n98 commonsourceibias.n23 161.3
R22641 commonsourceibias.n100 commonsourceibias.n99 161.3
R22642 commonsourceibias.n101 commonsourceibias.n22 161.3
R22643 commonsourceibias.n103 commonsourceibias.n102 161.3
R22644 commonsourceibias.n104 commonsourceibias.n21 161.3
R22645 commonsourceibias.n107 commonsourceibias.n106 161.3
R22646 commonsourceibias.n108 commonsourceibias.n20 161.3
R22647 commonsourceibias.n110 commonsourceibias.n109 161.3
R22648 commonsourceibias.n112 commonsourceibias.n18 161.3
R22649 commonsourceibias.n114 commonsourceibias.n113 161.3
R22650 commonsourceibias.n115 commonsourceibias.n17 161.3
R22651 commonsourceibias.n117 commonsourceibias.n116 161.3
R22652 commonsourceibias.n118 commonsourceibias.n16 161.3
R22653 commonsourceibias.n121 commonsourceibias.n120 161.3
R22654 commonsourceibias.n122 commonsourceibias.n15 161.3
R22655 commonsourceibias.n124 commonsourceibias.n123 161.3
R22656 commonsourceibias.n126 commonsourceibias.n14 161.3
R22657 commonsourceibias.n167 commonsourceibias.n164 161.3
R22658 commonsourceibias.n169 commonsourceibias.n168 161.3
R22659 commonsourceibias.n170 commonsourceibias.n163 161.3
R22660 commonsourceibias.n173 commonsourceibias.n172 161.3
R22661 commonsourceibias.n174 commonsourceibias.n162 161.3
R22662 commonsourceibias.n176 commonsourceibias.n175 161.3
R22663 commonsourceibias.n178 commonsourceibias.n160 161.3
R22664 commonsourceibias.n180 commonsourceibias.n179 161.3
R22665 commonsourceibias.n181 commonsourceibias.n159 161.3
R22666 commonsourceibias.n183 commonsourceibias.n182 161.3
R22667 commonsourceibias.n184 commonsourceibias.n158 161.3
R22668 commonsourceibias.n187 commonsourceibias.n186 161.3
R22669 commonsourceibias.n188 commonsourceibias.n157 161.3
R22670 commonsourceibias.n190 commonsourceibias.n189 161.3
R22671 commonsourceibias.n192 commonsourceibias.n156 161.3
R22672 commonsourceibias.n194 commonsourceibias.n193 161.3
R22673 commonsourceibias.n196 commonsourceibias.n195 161.3
R22674 commonsourceibias.n197 commonsourceibias.n154 161.3
R22675 commonsourceibias.n199 commonsourceibias.n198 161.3
R22676 commonsourceibias.n201 commonsourceibias.n200 161.3
R22677 commonsourceibias.n202 commonsourceibias.n152 161.3
R22678 commonsourceibias.n204 commonsourceibias.n203 161.3
R22679 commonsourceibias.n206 commonsourceibias.n205 161.3
R22680 commonsourceibias.n208 commonsourceibias.n207 161.3
R22681 commonsourceibias.n209 commonsourceibias.n13 161.3
R22682 commonsourceibias.n211 commonsourceibias.n210 161.3
R22683 commonsourceibias.n212 commonsourceibias.n12 161.3
R22684 commonsourceibias.n215 commonsourceibias.n214 161.3
R22685 commonsourceibias.n216 commonsourceibias.n11 161.3
R22686 commonsourceibias.n218 commonsourceibias.n217 161.3
R22687 commonsourceibias.n220 commonsourceibias.n9 161.3
R22688 commonsourceibias.n222 commonsourceibias.n221 161.3
R22689 commonsourceibias.n223 commonsourceibias.n8 161.3
R22690 commonsourceibias.n225 commonsourceibias.n224 161.3
R22691 commonsourceibias.n226 commonsourceibias.n7 161.3
R22692 commonsourceibias.n229 commonsourceibias.n228 161.3
R22693 commonsourceibias.n230 commonsourceibias.n6 161.3
R22694 commonsourceibias.n232 commonsourceibias.n231 161.3
R22695 commonsourceibias.n234 commonsourceibias.n4 161.3
R22696 commonsourceibias.n236 commonsourceibias.n235 161.3
R22697 commonsourceibias.n237 commonsourceibias.n3 161.3
R22698 commonsourceibias.n239 commonsourceibias.n238 161.3
R22699 commonsourceibias.n240 commonsourceibias.n2 161.3
R22700 commonsourceibias.n243 commonsourceibias.n242 161.3
R22701 commonsourceibias.n244 commonsourceibias.n1 161.3
R22702 commonsourceibias.n246 commonsourceibias.n245 161.3
R22703 commonsourceibias.n248 commonsourceibias.n0 161.3
R22704 commonsourceibias.n730 commonsourceibias.n618 161.3
R22705 commonsourceibias.n728 commonsourceibias.n727 161.3
R22706 commonsourceibias.n726 commonsourceibias.n619 161.3
R22707 commonsourceibias.n725 commonsourceibias.n724 161.3
R22708 commonsourceibias.n722 commonsourceibias.n620 161.3
R22709 commonsourceibias.n721 commonsourceibias.n720 161.3
R22710 commonsourceibias.n719 commonsourceibias.n621 161.3
R22711 commonsourceibias.n718 commonsourceibias.n717 161.3
R22712 commonsourceibias.n715 commonsourceibias.n622 161.3
R22713 commonsourceibias.n713 commonsourceibias.n712 161.3
R22714 commonsourceibias.n711 commonsourceibias.n623 161.3
R22715 commonsourceibias.n710 commonsourceibias.n709 161.3
R22716 commonsourceibias.n707 commonsourceibias.n624 161.3
R22717 commonsourceibias.n706 commonsourceibias.n705 161.3
R22718 commonsourceibias.n704 commonsourceibias.n625 161.3
R22719 commonsourceibias.n703 commonsourceibias.n702 161.3
R22720 commonsourceibias.n700 commonsourceibias.n626 161.3
R22721 commonsourceibias.n698 commonsourceibias.n697 161.3
R22722 commonsourceibias.n696 commonsourceibias.n627 161.3
R22723 commonsourceibias.n695 commonsourceibias.n694 161.3
R22724 commonsourceibias.n692 commonsourceibias.n628 161.3
R22725 commonsourceibias.n691 commonsourceibias.n690 161.3
R22726 commonsourceibias.n689 commonsourceibias.n629 161.3
R22727 commonsourceibias.n688 commonsourceibias.n687 161.3
R22728 commonsourceibias.n685 commonsourceibias.n630 161.3
R22729 commonsourceibias.n683 commonsourceibias.n682 161.3
R22730 commonsourceibias.n681 commonsourceibias.n631 161.3
R22731 commonsourceibias.n680 commonsourceibias.n679 161.3
R22732 commonsourceibias.n677 commonsourceibias.n632 161.3
R22733 commonsourceibias.n676 commonsourceibias.n675 161.3
R22734 commonsourceibias.n674 commonsourceibias.n633 161.3
R22735 commonsourceibias.n673 commonsourceibias.n672 161.3
R22736 commonsourceibias.n670 commonsourceibias.n634 161.3
R22737 commonsourceibias.n668 commonsourceibias.n667 161.3
R22738 commonsourceibias.n666 commonsourceibias.n635 161.3
R22739 commonsourceibias.n665 commonsourceibias.n664 161.3
R22740 commonsourceibias.n662 commonsourceibias.n636 161.3
R22741 commonsourceibias.n661 commonsourceibias.n660 161.3
R22742 commonsourceibias.n659 commonsourceibias.n637 161.3
R22743 commonsourceibias.n658 commonsourceibias.n657 161.3
R22744 commonsourceibias.n655 commonsourceibias.n638 161.3
R22745 commonsourceibias.n653 commonsourceibias.n652 161.3
R22746 commonsourceibias.n651 commonsourceibias.n639 161.3
R22747 commonsourceibias.n650 commonsourceibias.n649 161.3
R22748 commonsourceibias.n647 commonsourceibias.n640 161.3
R22749 commonsourceibias.n646 commonsourceibias.n645 161.3
R22750 commonsourceibias.n644 commonsourceibias.n641 161.3
R22751 commonsourceibias.n500 commonsourceibias.n388 161.3
R22752 commonsourceibias.n498 commonsourceibias.n497 161.3
R22753 commonsourceibias.n496 commonsourceibias.n389 161.3
R22754 commonsourceibias.n495 commonsourceibias.n494 161.3
R22755 commonsourceibias.n492 commonsourceibias.n390 161.3
R22756 commonsourceibias.n491 commonsourceibias.n490 161.3
R22757 commonsourceibias.n489 commonsourceibias.n391 161.3
R22758 commonsourceibias.n488 commonsourceibias.n487 161.3
R22759 commonsourceibias.n485 commonsourceibias.n392 161.3
R22760 commonsourceibias.n483 commonsourceibias.n482 161.3
R22761 commonsourceibias.n481 commonsourceibias.n393 161.3
R22762 commonsourceibias.n480 commonsourceibias.n479 161.3
R22763 commonsourceibias.n477 commonsourceibias.n394 161.3
R22764 commonsourceibias.n476 commonsourceibias.n475 161.3
R22765 commonsourceibias.n474 commonsourceibias.n395 161.3
R22766 commonsourceibias.n473 commonsourceibias.n472 161.3
R22767 commonsourceibias.n470 commonsourceibias.n396 161.3
R22768 commonsourceibias.n468 commonsourceibias.n467 161.3
R22769 commonsourceibias.n466 commonsourceibias.n397 161.3
R22770 commonsourceibias.n465 commonsourceibias.n464 161.3
R22771 commonsourceibias.n462 commonsourceibias.n398 161.3
R22772 commonsourceibias.n461 commonsourceibias.n460 161.3
R22773 commonsourceibias.n459 commonsourceibias.n399 161.3
R22774 commonsourceibias.n458 commonsourceibias.n457 161.3
R22775 commonsourceibias.n455 commonsourceibias.n400 161.3
R22776 commonsourceibias.n453 commonsourceibias.n452 161.3
R22777 commonsourceibias.n451 commonsourceibias.n401 161.3
R22778 commonsourceibias.n450 commonsourceibias.n449 161.3
R22779 commonsourceibias.n447 commonsourceibias.n402 161.3
R22780 commonsourceibias.n446 commonsourceibias.n445 161.3
R22781 commonsourceibias.n444 commonsourceibias.n403 161.3
R22782 commonsourceibias.n443 commonsourceibias.n442 161.3
R22783 commonsourceibias.n440 commonsourceibias.n404 161.3
R22784 commonsourceibias.n438 commonsourceibias.n437 161.3
R22785 commonsourceibias.n436 commonsourceibias.n405 161.3
R22786 commonsourceibias.n435 commonsourceibias.n434 161.3
R22787 commonsourceibias.n432 commonsourceibias.n406 161.3
R22788 commonsourceibias.n431 commonsourceibias.n430 161.3
R22789 commonsourceibias.n429 commonsourceibias.n407 161.3
R22790 commonsourceibias.n428 commonsourceibias.n427 161.3
R22791 commonsourceibias.n425 commonsourceibias.n408 161.3
R22792 commonsourceibias.n423 commonsourceibias.n422 161.3
R22793 commonsourceibias.n421 commonsourceibias.n409 161.3
R22794 commonsourceibias.n420 commonsourceibias.n419 161.3
R22795 commonsourceibias.n417 commonsourceibias.n410 161.3
R22796 commonsourceibias.n416 commonsourceibias.n415 161.3
R22797 commonsourceibias.n414 commonsourceibias.n411 161.3
R22798 commonsourceibias.n570 commonsourceibias.n569 161.3
R22799 commonsourceibias.n568 commonsourceibias.n567 161.3
R22800 commonsourceibias.n566 commonsourceibias.n516 161.3
R22801 commonsourceibias.n565 commonsourceibias.n564 161.3
R22802 commonsourceibias.n563 commonsourceibias.n562 161.3
R22803 commonsourceibias.n561 commonsourceibias.n518 161.3
R22804 commonsourceibias.n560 commonsourceibias.n559 161.3
R22805 commonsourceibias.n558 commonsourceibias.n557 161.3
R22806 commonsourceibias.n556 commonsourceibias.n520 161.3
R22807 commonsourceibias.n554 commonsourceibias.n553 161.3
R22808 commonsourceibias.n552 commonsourceibias.n521 161.3
R22809 commonsourceibias.n551 commonsourceibias.n550 161.3
R22810 commonsourceibias.n548 commonsourceibias.n522 161.3
R22811 commonsourceibias.n547 commonsourceibias.n546 161.3
R22812 commonsourceibias.n545 commonsourceibias.n523 161.3
R22813 commonsourceibias.n544 commonsourceibias.n543 161.3
R22814 commonsourceibias.n541 commonsourceibias.n524 161.3
R22815 commonsourceibias.n539 commonsourceibias.n538 161.3
R22816 commonsourceibias.n537 commonsourceibias.n525 161.3
R22817 commonsourceibias.n536 commonsourceibias.n535 161.3
R22818 commonsourceibias.n533 commonsourceibias.n526 161.3
R22819 commonsourceibias.n532 commonsourceibias.n531 161.3
R22820 commonsourceibias.n530 commonsourceibias.n527 161.3
R22821 commonsourceibias.n615 commonsourceibias.n367 161.3
R22822 commonsourceibias.n613 commonsourceibias.n612 161.3
R22823 commonsourceibias.n611 commonsourceibias.n368 161.3
R22824 commonsourceibias.n610 commonsourceibias.n609 161.3
R22825 commonsourceibias.n607 commonsourceibias.n369 161.3
R22826 commonsourceibias.n606 commonsourceibias.n605 161.3
R22827 commonsourceibias.n604 commonsourceibias.n370 161.3
R22828 commonsourceibias.n603 commonsourceibias.n602 161.3
R22829 commonsourceibias.n600 commonsourceibias.n371 161.3
R22830 commonsourceibias.n598 commonsourceibias.n597 161.3
R22831 commonsourceibias.n596 commonsourceibias.n372 161.3
R22832 commonsourceibias.n595 commonsourceibias.n594 161.3
R22833 commonsourceibias.n592 commonsourceibias.n373 161.3
R22834 commonsourceibias.n591 commonsourceibias.n590 161.3
R22835 commonsourceibias.n589 commonsourceibias.n374 161.3
R22836 commonsourceibias.n588 commonsourceibias.n587 161.3
R22837 commonsourceibias.n585 commonsourceibias.n375 161.3
R22838 commonsourceibias.n583 commonsourceibias.n582 161.3
R22839 commonsourceibias.n581 commonsourceibias.n376 161.3
R22840 commonsourceibias.n580 commonsourceibias.n579 161.3
R22841 commonsourceibias.n577 commonsourceibias.n377 161.3
R22842 commonsourceibias.n576 commonsourceibias.n575 161.3
R22843 commonsourceibias.n574 commonsourceibias.n378 161.3
R22844 commonsourceibias.n573 commonsourceibias.n572 161.3
R22845 commonsourceibias.n141 commonsourceibias.n139 81.5057
R22846 commonsourceibias.n381 commonsourceibias.n379 81.5057
R22847 commonsourceibias.n141 commonsourceibias.n140 80.9324
R22848 commonsourceibias.n143 commonsourceibias.n142 80.9324
R22849 commonsourceibias.n145 commonsourceibias.n144 80.9324
R22850 commonsourceibias.n147 commonsourceibias.n146 80.9324
R22851 commonsourceibias.n138 commonsourceibias.n137 80.9324
R22852 commonsourceibias.n136 commonsourceibias.n135 80.9324
R22853 commonsourceibias.n134 commonsourceibias.n133 80.9324
R22854 commonsourceibias.n132 commonsourceibias.n131 80.9324
R22855 commonsourceibias.n130 commonsourceibias.n129 80.9324
R22856 commonsourceibias.n504 commonsourceibias.n503 80.9324
R22857 commonsourceibias.n506 commonsourceibias.n505 80.9324
R22858 commonsourceibias.n508 commonsourceibias.n507 80.9324
R22859 commonsourceibias.n510 commonsourceibias.n509 80.9324
R22860 commonsourceibias.n512 commonsourceibias.n511 80.9324
R22861 commonsourceibias.n387 commonsourceibias.n386 80.9324
R22862 commonsourceibias.n385 commonsourceibias.n384 80.9324
R22863 commonsourceibias.n383 commonsourceibias.n382 80.9324
R22864 commonsourceibias.n381 commonsourceibias.n380 80.9324
R22865 commonsourceibias.n365 commonsourceibias.n364 80.6037
R22866 commonsourceibias.n128 commonsourceibias.n127 80.6037
R22867 commonsourceibias.n250 commonsourceibias.n249 80.6037
R22868 commonsourceibias.n732 commonsourceibias.n731 80.6037
R22869 commonsourceibias.n502 commonsourceibias.n501 80.6037
R22870 commonsourceibias.n617 commonsourceibias.n616 80.6037
R22871 commonsourceibias.n322 commonsourceibias.n321 56.5617
R22872 commonsourceibias.n336 commonsourceibias.n335 56.5617
R22873 commonsourceibias.n85 commonsourceibias.n84 56.5617
R22874 commonsourceibias.n71 commonsourceibias.n70 56.5617
R22875 commonsourceibias.n207 commonsourceibias.n206 56.5617
R22876 commonsourceibias.n193 commonsourceibias.n192 56.5617
R22877 commonsourceibias.n687 commonsourceibias.n685 56.5617
R22878 commonsourceibias.n702 commonsourceibias.n700 56.5617
R22879 commonsourceibias.n457 commonsourceibias.n455 56.5617
R22880 commonsourceibias.n472 commonsourceibias.n470 56.5617
R22881 commonsourceibias.n572 commonsourceibias.n570 56.5617
R22882 commonsourceibias.n294 commonsourceibias.n293 56.5617
R22883 commonsourceibias.n308 commonsourceibias.n307 56.5617
R22884 commonsourceibias.n350 commonsourceibias.n349 56.5617
R22885 commonsourceibias.n113 commonsourceibias.n112 56.5617
R22886 commonsourceibias.n99 commonsourceibias.n98 56.5617
R22887 commonsourceibias.n57 commonsourceibias.n56 56.5617
R22888 commonsourceibias.n235 commonsourceibias.n234 56.5617
R22889 commonsourceibias.n221 commonsourceibias.n220 56.5617
R22890 commonsourceibias.n179 commonsourceibias.n178 56.5617
R22891 commonsourceibias.n657 commonsourceibias.n655 56.5617
R22892 commonsourceibias.n672 commonsourceibias.n670 56.5617
R22893 commonsourceibias.n717 commonsourceibias.n715 56.5617
R22894 commonsourceibias.n427 commonsourceibias.n425 56.5617
R22895 commonsourceibias.n442 commonsourceibias.n440 56.5617
R22896 commonsourceibias.n487 commonsourceibias.n485 56.5617
R22897 commonsourceibias.n602 commonsourceibias.n600 56.5617
R22898 commonsourceibias.n587 commonsourceibias.n585 56.5617
R22899 commonsourceibias.n543 commonsourceibias.n541 56.5617
R22900 commonsourceibias.n557 commonsourceibias.n556 56.5617
R22901 commonsourceibias.n285 commonsourceibias.n284 51.2335
R22902 commonsourceibias.n357 commonsourceibias.n252 51.2335
R22903 commonsourceibias.n120 commonsourceibias.n15 51.2335
R22904 commonsourceibias.n48 commonsourceibias.n47 51.2335
R22905 commonsourceibias.n242 commonsourceibias.n1 51.2335
R22906 commonsourceibias.n170 commonsourceibias.n169 51.2335
R22907 commonsourceibias.n647 commonsourceibias.n646 51.2335
R22908 commonsourceibias.n724 commonsourceibias.n619 51.2335
R22909 commonsourceibias.n417 commonsourceibias.n416 51.2335
R22910 commonsourceibias.n494 commonsourceibias.n389 51.2335
R22911 commonsourceibias.n609 commonsourceibias.n368 51.2335
R22912 commonsourceibias.n533 commonsourceibias.n532 51.2335
R22913 commonsourceibias.n364 commonsourceibias.n363 50.9056
R22914 commonsourceibias.n127 commonsourceibias.n126 50.9056
R22915 commonsourceibias.n249 commonsourceibias.n248 50.9056
R22916 commonsourceibias.n731 commonsourceibias.n730 50.9056
R22917 commonsourceibias.n501 commonsourceibias.n500 50.9056
R22918 commonsourceibias.n616 commonsourceibias.n615 50.9056
R22919 commonsourceibias.n299 commonsourceibias.n298 50.2647
R22920 commonsourceibias.n343 commonsourceibias.n257 50.2647
R22921 commonsourceibias.n106 commonsourceibias.n20 50.2647
R22922 commonsourceibias.n62 commonsourceibias.n61 50.2647
R22923 commonsourceibias.n228 commonsourceibias.n6 50.2647
R22924 commonsourceibias.n184 commonsourceibias.n183 50.2647
R22925 commonsourceibias.n662 commonsourceibias.n661 50.2647
R22926 commonsourceibias.n709 commonsourceibias.n623 50.2647
R22927 commonsourceibias.n432 commonsourceibias.n431 50.2647
R22928 commonsourceibias.n479 commonsourceibias.n393 50.2647
R22929 commonsourceibias.n594 commonsourceibias.n372 50.2647
R22930 commonsourceibias.n548 commonsourceibias.n547 50.2647
R22931 commonsourceibias.n281 commonsourceibias.n280 49.9027
R22932 commonsourceibias.n44 commonsourceibias.n43 49.9027
R22933 commonsourceibias.n166 commonsourceibias.n165 49.9027
R22934 commonsourceibias.n643 commonsourceibias.n642 49.9027
R22935 commonsourceibias.n413 commonsourceibias.n412 49.9027
R22936 commonsourceibias.n529 commonsourceibias.n528 49.9027
R22937 commonsourceibias.n313 commonsourceibias.n312 49.296
R22938 commonsourceibias.n329 commonsourceibias.n262 49.296
R22939 commonsourceibias.n92 commonsourceibias.n25 49.296
R22940 commonsourceibias.n76 commonsourceibias.n75 49.296
R22941 commonsourceibias.n214 commonsourceibias.n11 49.296
R22942 commonsourceibias.n198 commonsourceibias.n197 49.296
R22943 commonsourceibias.n677 commonsourceibias.n676 49.296
R22944 commonsourceibias.n694 commonsourceibias.n627 49.296
R22945 commonsourceibias.n447 commonsourceibias.n446 49.296
R22946 commonsourceibias.n464 commonsourceibias.n397 49.296
R22947 commonsourceibias.n579 commonsourceibias.n376 49.296
R22948 commonsourceibias.n562 commonsourceibias.n561 49.296
R22949 commonsourceibias.n315 commonsourceibias.n267 48.3272
R22950 commonsourceibias.n327 commonsourceibias.n326 48.3272
R22951 commonsourceibias.n90 commonsourceibias.n89 48.3272
R22952 commonsourceibias.n78 commonsourceibias.n30 48.3272
R22953 commonsourceibias.n212 commonsourceibias.n211 48.3272
R22954 commonsourceibias.n202 commonsourceibias.n201 48.3272
R22955 commonsourceibias.n679 commonsourceibias.n631 48.3272
R22956 commonsourceibias.n692 commonsourceibias.n691 48.3272
R22957 commonsourceibias.n449 commonsourceibias.n401 48.3272
R22958 commonsourceibias.n462 commonsourceibias.n461 48.3272
R22959 commonsourceibias.n577 commonsourceibias.n576 48.3272
R22960 commonsourceibias.n566 commonsourceibias.n565 48.3272
R22961 commonsourceibias.n301 commonsourceibias.n272 47.3584
R22962 commonsourceibias.n341 commonsourceibias.n340 47.3584
R22963 commonsourceibias.n104 commonsourceibias.n103 47.3584
R22964 commonsourceibias.n64 commonsourceibias.n35 47.3584
R22965 commonsourceibias.n226 commonsourceibias.n225 47.3584
R22966 commonsourceibias.n186 commonsourceibias.n157 47.3584
R22967 commonsourceibias.n664 commonsourceibias.n635 47.3584
R22968 commonsourceibias.n707 commonsourceibias.n706 47.3584
R22969 commonsourceibias.n434 commonsourceibias.n405 47.3584
R22970 commonsourceibias.n477 commonsourceibias.n476 47.3584
R22971 commonsourceibias.n592 commonsourceibias.n591 47.3584
R22972 commonsourceibias.n550 commonsourceibias.n521 47.3584
R22973 commonsourceibias.n287 commonsourceibias.n277 46.3896
R22974 commonsourceibias.n355 commonsourceibias.n354 46.3896
R22975 commonsourceibias.n118 commonsourceibias.n117 46.3896
R22976 commonsourceibias.n50 commonsourceibias.n40 46.3896
R22977 commonsourceibias.n240 commonsourceibias.n239 46.3896
R22978 commonsourceibias.n172 commonsourceibias.n162 46.3896
R22979 commonsourceibias.n649 commonsourceibias.n639 46.3896
R22980 commonsourceibias.n722 commonsourceibias.n721 46.3896
R22981 commonsourceibias.n419 commonsourceibias.n409 46.3896
R22982 commonsourceibias.n492 commonsourceibias.n491 46.3896
R22983 commonsourceibias.n607 commonsourceibias.n606 46.3896
R22984 commonsourceibias.n535 commonsourceibias.n525 46.3896
R22985 commonsourceibias.n282 commonsourceibias.n281 44.7059
R22986 commonsourceibias.n644 commonsourceibias.n643 44.7059
R22987 commonsourceibias.n414 commonsourceibias.n413 44.7059
R22988 commonsourceibias.n530 commonsourceibias.n529 44.7059
R22989 commonsourceibias.n45 commonsourceibias.n44 44.7059
R22990 commonsourceibias.n167 commonsourceibias.n166 44.7059
R22991 commonsourceibias.n291 commonsourceibias.n277 34.7644
R22992 commonsourceibias.n354 commonsourceibias.n254 34.7644
R22993 commonsourceibias.n117 commonsourceibias.n17 34.7644
R22994 commonsourceibias.n54 commonsourceibias.n40 34.7644
R22995 commonsourceibias.n239 commonsourceibias.n3 34.7644
R22996 commonsourceibias.n176 commonsourceibias.n162 34.7644
R22997 commonsourceibias.n653 commonsourceibias.n639 34.7644
R22998 commonsourceibias.n721 commonsourceibias.n621 34.7644
R22999 commonsourceibias.n423 commonsourceibias.n409 34.7644
R23000 commonsourceibias.n491 commonsourceibias.n391 34.7644
R23001 commonsourceibias.n606 commonsourceibias.n370 34.7644
R23002 commonsourceibias.n539 commonsourceibias.n525 34.7644
R23003 commonsourceibias.n305 commonsourceibias.n272 33.7956
R23004 commonsourceibias.n340 commonsourceibias.n259 33.7956
R23005 commonsourceibias.n103 commonsourceibias.n22 33.7956
R23006 commonsourceibias.n68 commonsourceibias.n35 33.7956
R23007 commonsourceibias.n225 commonsourceibias.n8 33.7956
R23008 commonsourceibias.n190 commonsourceibias.n157 33.7956
R23009 commonsourceibias.n668 commonsourceibias.n635 33.7956
R23010 commonsourceibias.n706 commonsourceibias.n625 33.7956
R23011 commonsourceibias.n438 commonsourceibias.n405 33.7956
R23012 commonsourceibias.n476 commonsourceibias.n395 33.7956
R23013 commonsourceibias.n591 commonsourceibias.n374 33.7956
R23014 commonsourceibias.n554 commonsourceibias.n521 33.7956
R23015 commonsourceibias.n319 commonsourceibias.n267 32.8269
R23016 commonsourceibias.n326 commonsourceibias.n264 32.8269
R23017 commonsourceibias.n89 commonsourceibias.n27 32.8269
R23018 commonsourceibias.n82 commonsourceibias.n30 32.8269
R23019 commonsourceibias.n211 commonsourceibias.n13 32.8269
R23020 commonsourceibias.n203 commonsourceibias.n202 32.8269
R23021 commonsourceibias.n683 commonsourceibias.n631 32.8269
R23022 commonsourceibias.n691 commonsourceibias.n629 32.8269
R23023 commonsourceibias.n453 commonsourceibias.n401 32.8269
R23024 commonsourceibias.n461 commonsourceibias.n399 32.8269
R23025 commonsourceibias.n576 commonsourceibias.n378 32.8269
R23026 commonsourceibias.n567 commonsourceibias.n566 32.8269
R23027 commonsourceibias.n312 commonsourceibias.n269 31.8581
R23028 commonsourceibias.n333 commonsourceibias.n262 31.8581
R23029 commonsourceibias.n96 commonsourceibias.n25 31.8581
R23030 commonsourceibias.n75 commonsourceibias.n32 31.8581
R23031 commonsourceibias.n218 commonsourceibias.n11 31.8581
R23032 commonsourceibias.n197 commonsourceibias.n196 31.8581
R23033 commonsourceibias.n676 commonsourceibias.n633 31.8581
R23034 commonsourceibias.n698 commonsourceibias.n627 31.8581
R23035 commonsourceibias.n446 commonsourceibias.n403 31.8581
R23036 commonsourceibias.n468 commonsourceibias.n397 31.8581
R23037 commonsourceibias.n583 commonsourceibias.n376 31.8581
R23038 commonsourceibias.n561 commonsourceibias.n560 31.8581
R23039 commonsourceibias.n298 commonsourceibias.n274 30.8893
R23040 commonsourceibias.n347 commonsourceibias.n257 30.8893
R23041 commonsourceibias.n110 commonsourceibias.n20 30.8893
R23042 commonsourceibias.n61 commonsourceibias.n37 30.8893
R23043 commonsourceibias.n232 commonsourceibias.n6 30.8893
R23044 commonsourceibias.n183 commonsourceibias.n159 30.8893
R23045 commonsourceibias.n661 commonsourceibias.n637 30.8893
R23046 commonsourceibias.n713 commonsourceibias.n623 30.8893
R23047 commonsourceibias.n431 commonsourceibias.n407 30.8893
R23048 commonsourceibias.n483 commonsourceibias.n393 30.8893
R23049 commonsourceibias.n598 commonsourceibias.n372 30.8893
R23050 commonsourceibias.n547 commonsourceibias.n523 30.8893
R23051 commonsourceibias.n284 commonsourceibias.n279 29.9206
R23052 commonsourceibias.n361 commonsourceibias.n252 29.9206
R23053 commonsourceibias.n124 commonsourceibias.n15 29.9206
R23054 commonsourceibias.n47 commonsourceibias.n42 29.9206
R23055 commonsourceibias.n246 commonsourceibias.n1 29.9206
R23056 commonsourceibias.n169 commonsourceibias.n164 29.9206
R23057 commonsourceibias.n646 commonsourceibias.n641 29.9206
R23058 commonsourceibias.n728 commonsourceibias.n619 29.9206
R23059 commonsourceibias.n416 commonsourceibias.n411 29.9206
R23060 commonsourceibias.n498 commonsourceibias.n389 29.9206
R23061 commonsourceibias.n613 commonsourceibias.n368 29.9206
R23062 commonsourceibias.n532 commonsourceibias.n527 29.9206
R23063 commonsourceibias.n363 commonsourceibias.n362 21.8872
R23064 commonsourceibias.n126 commonsourceibias.n125 21.8872
R23065 commonsourceibias.n248 commonsourceibias.n247 21.8872
R23066 commonsourceibias.n730 commonsourceibias.n729 21.8872
R23067 commonsourceibias.n500 commonsourceibias.n499 21.8872
R23068 commonsourceibias.n615 commonsourceibias.n614 21.8872
R23069 commonsourceibias.n294 commonsourceibias.n276 21.3954
R23070 commonsourceibias.n349 commonsourceibias.n348 21.3954
R23071 commonsourceibias.n112 commonsourceibias.n111 21.3954
R23072 commonsourceibias.n57 commonsourceibias.n39 21.3954
R23073 commonsourceibias.n234 commonsourceibias.n233 21.3954
R23074 commonsourceibias.n179 commonsourceibias.n161 21.3954
R23075 commonsourceibias.n657 commonsourceibias.n656 21.3954
R23076 commonsourceibias.n715 commonsourceibias.n714 21.3954
R23077 commonsourceibias.n427 commonsourceibias.n426 21.3954
R23078 commonsourceibias.n485 commonsourceibias.n484 21.3954
R23079 commonsourceibias.n600 commonsourceibias.n599 21.3954
R23080 commonsourceibias.n543 commonsourceibias.n542 21.3954
R23081 commonsourceibias.n308 commonsourceibias.n271 20.9036
R23082 commonsourceibias.n335 commonsourceibias.n334 20.9036
R23083 commonsourceibias.n98 commonsourceibias.n97 20.9036
R23084 commonsourceibias.n71 commonsourceibias.n34 20.9036
R23085 commonsourceibias.n220 commonsourceibias.n219 20.9036
R23086 commonsourceibias.n193 commonsourceibias.n155 20.9036
R23087 commonsourceibias.n672 commonsourceibias.n671 20.9036
R23088 commonsourceibias.n700 commonsourceibias.n699 20.9036
R23089 commonsourceibias.n442 commonsourceibias.n441 20.9036
R23090 commonsourceibias.n470 commonsourceibias.n469 20.9036
R23091 commonsourceibias.n585 commonsourceibias.n584 20.9036
R23092 commonsourceibias.n557 commonsourceibias.n519 20.9036
R23093 commonsourceibias.n321 commonsourceibias.n320 20.4117
R23094 commonsourceibias.n322 commonsourceibias.n266 20.4117
R23095 commonsourceibias.n85 commonsourceibias.n29 20.4117
R23096 commonsourceibias.n84 commonsourceibias.n83 20.4117
R23097 commonsourceibias.n207 commonsourceibias.n150 20.4117
R23098 commonsourceibias.n206 commonsourceibias.n151 20.4117
R23099 commonsourceibias.n685 commonsourceibias.n684 20.4117
R23100 commonsourceibias.n687 commonsourceibias.n686 20.4117
R23101 commonsourceibias.n455 commonsourceibias.n454 20.4117
R23102 commonsourceibias.n457 commonsourceibias.n456 20.4117
R23103 commonsourceibias.n572 commonsourceibias.n571 20.4117
R23104 commonsourceibias.n570 commonsourceibias.n515 20.4117
R23105 commonsourceibias.n307 commonsourceibias.n306 19.9199
R23106 commonsourceibias.n336 commonsourceibias.n261 19.9199
R23107 commonsourceibias.n99 commonsourceibias.n24 19.9199
R23108 commonsourceibias.n70 commonsourceibias.n69 19.9199
R23109 commonsourceibias.n221 commonsourceibias.n10 19.9199
R23110 commonsourceibias.n192 commonsourceibias.n191 19.9199
R23111 commonsourceibias.n670 commonsourceibias.n669 19.9199
R23112 commonsourceibias.n702 commonsourceibias.n701 19.9199
R23113 commonsourceibias.n440 commonsourceibias.n439 19.9199
R23114 commonsourceibias.n472 commonsourceibias.n471 19.9199
R23115 commonsourceibias.n587 commonsourceibias.n586 19.9199
R23116 commonsourceibias.n556 commonsourceibias.n555 19.9199
R23117 commonsourceibias.n293 commonsourceibias.n292 19.4281
R23118 commonsourceibias.n350 commonsourceibias.n256 19.4281
R23119 commonsourceibias.n113 commonsourceibias.n19 19.4281
R23120 commonsourceibias.n56 commonsourceibias.n55 19.4281
R23121 commonsourceibias.n235 commonsourceibias.n5 19.4281
R23122 commonsourceibias.n178 commonsourceibias.n177 19.4281
R23123 commonsourceibias.n655 commonsourceibias.n654 19.4281
R23124 commonsourceibias.n717 commonsourceibias.n716 19.4281
R23125 commonsourceibias.n425 commonsourceibias.n424 19.4281
R23126 commonsourceibias.n487 commonsourceibias.n486 19.4281
R23127 commonsourceibias.n602 commonsourceibias.n601 19.4281
R23128 commonsourceibias.n541 commonsourceibias.n540 19.4281
R23129 commonsourceibias.n286 commonsourceibias.n285 13.526
R23130 commonsourceibias.n357 commonsourceibias.n356 13.526
R23131 commonsourceibias.n120 commonsourceibias.n119 13.526
R23132 commonsourceibias.n49 commonsourceibias.n48 13.526
R23133 commonsourceibias.n242 commonsourceibias.n241 13.526
R23134 commonsourceibias.n171 commonsourceibias.n170 13.526
R23135 commonsourceibias.n648 commonsourceibias.n647 13.526
R23136 commonsourceibias.n724 commonsourceibias.n723 13.526
R23137 commonsourceibias.n418 commonsourceibias.n417 13.526
R23138 commonsourceibias.n494 commonsourceibias.n493 13.526
R23139 commonsourceibias.n609 commonsourceibias.n608 13.526
R23140 commonsourceibias.n534 commonsourceibias.n533 13.526
R23141 commonsourceibias.n130 commonsourceibias.n128 13.2322
R23142 commonsourceibias.n504 commonsourceibias.n502 13.2322
R23143 commonsourceibias.n300 commonsourceibias.n299 13.0342
R23144 commonsourceibias.n343 commonsourceibias.n342 13.0342
R23145 commonsourceibias.n106 commonsourceibias.n105 13.0342
R23146 commonsourceibias.n63 commonsourceibias.n62 13.0342
R23147 commonsourceibias.n228 commonsourceibias.n227 13.0342
R23148 commonsourceibias.n185 commonsourceibias.n184 13.0342
R23149 commonsourceibias.n663 commonsourceibias.n662 13.0342
R23150 commonsourceibias.n709 commonsourceibias.n708 13.0342
R23151 commonsourceibias.n433 commonsourceibias.n432 13.0342
R23152 commonsourceibias.n479 commonsourceibias.n478 13.0342
R23153 commonsourceibias.n594 commonsourceibias.n593 13.0342
R23154 commonsourceibias.n549 commonsourceibias.n548 13.0342
R23155 commonsourceibias.n314 commonsourceibias.n313 12.5423
R23156 commonsourceibias.n329 commonsourceibias.n328 12.5423
R23157 commonsourceibias.n92 commonsourceibias.n91 12.5423
R23158 commonsourceibias.n77 commonsourceibias.n76 12.5423
R23159 commonsourceibias.n214 commonsourceibias.n213 12.5423
R23160 commonsourceibias.n198 commonsourceibias.n153 12.5423
R23161 commonsourceibias.n678 commonsourceibias.n677 12.5423
R23162 commonsourceibias.n694 commonsourceibias.n693 12.5423
R23163 commonsourceibias.n448 commonsourceibias.n447 12.5423
R23164 commonsourceibias.n464 commonsourceibias.n463 12.5423
R23165 commonsourceibias.n579 commonsourceibias.n578 12.5423
R23166 commonsourceibias.n562 commonsourceibias.n517 12.5423
R23167 commonsourceibias.n734 commonsourceibias.n366 12.2777
R23168 commonsourceibias.n315 commonsourceibias.n314 12.0505
R23169 commonsourceibias.n328 commonsourceibias.n327 12.0505
R23170 commonsourceibias.n91 commonsourceibias.n90 12.0505
R23171 commonsourceibias.n78 commonsourceibias.n77 12.0505
R23172 commonsourceibias.n213 commonsourceibias.n212 12.0505
R23173 commonsourceibias.n201 commonsourceibias.n153 12.0505
R23174 commonsourceibias.n679 commonsourceibias.n678 12.0505
R23175 commonsourceibias.n693 commonsourceibias.n692 12.0505
R23176 commonsourceibias.n449 commonsourceibias.n448 12.0505
R23177 commonsourceibias.n463 commonsourceibias.n462 12.0505
R23178 commonsourceibias.n578 commonsourceibias.n577 12.0505
R23179 commonsourceibias.n565 commonsourceibias.n517 12.0505
R23180 commonsourceibias.n301 commonsourceibias.n300 11.5587
R23181 commonsourceibias.n342 commonsourceibias.n341 11.5587
R23182 commonsourceibias.n105 commonsourceibias.n104 11.5587
R23183 commonsourceibias.n64 commonsourceibias.n63 11.5587
R23184 commonsourceibias.n227 commonsourceibias.n226 11.5587
R23185 commonsourceibias.n186 commonsourceibias.n185 11.5587
R23186 commonsourceibias.n664 commonsourceibias.n663 11.5587
R23187 commonsourceibias.n708 commonsourceibias.n707 11.5587
R23188 commonsourceibias.n434 commonsourceibias.n433 11.5587
R23189 commonsourceibias.n478 commonsourceibias.n477 11.5587
R23190 commonsourceibias.n593 commonsourceibias.n592 11.5587
R23191 commonsourceibias.n550 commonsourceibias.n549 11.5587
R23192 commonsourceibias.n287 commonsourceibias.n286 11.0668
R23193 commonsourceibias.n356 commonsourceibias.n355 11.0668
R23194 commonsourceibias.n119 commonsourceibias.n118 11.0668
R23195 commonsourceibias.n50 commonsourceibias.n49 11.0668
R23196 commonsourceibias.n241 commonsourceibias.n240 11.0668
R23197 commonsourceibias.n172 commonsourceibias.n171 11.0668
R23198 commonsourceibias.n649 commonsourceibias.n648 11.0668
R23199 commonsourceibias.n723 commonsourceibias.n722 11.0668
R23200 commonsourceibias.n419 commonsourceibias.n418 11.0668
R23201 commonsourceibias.n493 commonsourceibias.n492 11.0668
R23202 commonsourceibias.n608 commonsourceibias.n607 11.0668
R23203 commonsourceibias.n535 commonsourceibias.n534 11.0668
R23204 commonsourceibias.n734 commonsourceibias.n733 10.3347
R23205 commonsourceibias.n149 commonsourceibias.n148 9.50363
R23206 commonsourceibias.n514 commonsourceibias.n513 9.50363
R23207 commonsourceibias.n366 commonsourceibias.n250 8.75852
R23208 commonsourceibias.n733 commonsourceibias.n617 8.75852
R23209 commonsourceibias.n292 commonsourceibias.n291 5.16479
R23210 commonsourceibias.n256 commonsourceibias.n254 5.16479
R23211 commonsourceibias.n19 commonsourceibias.n17 5.16479
R23212 commonsourceibias.n55 commonsourceibias.n54 5.16479
R23213 commonsourceibias.n5 commonsourceibias.n3 5.16479
R23214 commonsourceibias.n177 commonsourceibias.n176 5.16479
R23215 commonsourceibias.n654 commonsourceibias.n653 5.16479
R23216 commonsourceibias.n716 commonsourceibias.n621 5.16479
R23217 commonsourceibias.n424 commonsourceibias.n423 5.16479
R23218 commonsourceibias.n486 commonsourceibias.n391 5.16479
R23219 commonsourceibias.n601 commonsourceibias.n370 5.16479
R23220 commonsourceibias.n540 commonsourceibias.n539 5.16479
R23221 commonsourceibias.n366 commonsourceibias.n365 5.03125
R23222 commonsourceibias.n733 commonsourceibias.n732 5.03125
R23223 commonsourceibias.n306 commonsourceibias.n305 4.67295
R23224 commonsourceibias.n261 commonsourceibias.n259 4.67295
R23225 commonsourceibias.n24 commonsourceibias.n22 4.67295
R23226 commonsourceibias.n69 commonsourceibias.n68 4.67295
R23227 commonsourceibias.n10 commonsourceibias.n8 4.67295
R23228 commonsourceibias.n191 commonsourceibias.n190 4.67295
R23229 commonsourceibias.n669 commonsourceibias.n668 4.67295
R23230 commonsourceibias.n701 commonsourceibias.n625 4.67295
R23231 commonsourceibias.n439 commonsourceibias.n438 4.67295
R23232 commonsourceibias.n471 commonsourceibias.n395 4.67295
R23233 commonsourceibias.n586 commonsourceibias.n374 4.67295
R23234 commonsourceibias.n555 commonsourceibias.n554 4.67295
R23235 commonsourceibias commonsourceibias.n734 4.20978
R23236 commonsourceibias.n320 commonsourceibias.n319 4.18111
R23237 commonsourceibias.n266 commonsourceibias.n264 4.18111
R23238 commonsourceibias.n29 commonsourceibias.n27 4.18111
R23239 commonsourceibias.n83 commonsourceibias.n82 4.18111
R23240 commonsourceibias.n150 commonsourceibias.n13 4.18111
R23241 commonsourceibias.n203 commonsourceibias.n151 4.18111
R23242 commonsourceibias.n684 commonsourceibias.n683 4.18111
R23243 commonsourceibias.n686 commonsourceibias.n629 4.18111
R23244 commonsourceibias.n454 commonsourceibias.n453 4.18111
R23245 commonsourceibias.n456 commonsourceibias.n399 4.18111
R23246 commonsourceibias.n571 commonsourceibias.n378 4.18111
R23247 commonsourceibias.n567 commonsourceibias.n515 4.18111
R23248 commonsourceibias.n271 commonsourceibias.n269 3.68928
R23249 commonsourceibias.n334 commonsourceibias.n333 3.68928
R23250 commonsourceibias.n97 commonsourceibias.n96 3.68928
R23251 commonsourceibias.n34 commonsourceibias.n32 3.68928
R23252 commonsourceibias.n219 commonsourceibias.n218 3.68928
R23253 commonsourceibias.n196 commonsourceibias.n155 3.68928
R23254 commonsourceibias.n671 commonsourceibias.n633 3.68928
R23255 commonsourceibias.n699 commonsourceibias.n698 3.68928
R23256 commonsourceibias.n441 commonsourceibias.n403 3.68928
R23257 commonsourceibias.n469 commonsourceibias.n468 3.68928
R23258 commonsourceibias.n584 commonsourceibias.n583 3.68928
R23259 commonsourceibias.n560 commonsourceibias.n519 3.68928
R23260 commonsourceibias.n276 commonsourceibias.n274 3.19744
R23261 commonsourceibias.n348 commonsourceibias.n347 3.19744
R23262 commonsourceibias.n111 commonsourceibias.n110 3.19744
R23263 commonsourceibias.n39 commonsourceibias.n37 3.19744
R23264 commonsourceibias.n233 commonsourceibias.n232 3.19744
R23265 commonsourceibias.n161 commonsourceibias.n159 3.19744
R23266 commonsourceibias.n656 commonsourceibias.n637 3.19744
R23267 commonsourceibias.n714 commonsourceibias.n713 3.19744
R23268 commonsourceibias.n426 commonsourceibias.n407 3.19744
R23269 commonsourceibias.n484 commonsourceibias.n483 3.19744
R23270 commonsourceibias.n599 commonsourceibias.n598 3.19744
R23271 commonsourceibias.n542 commonsourceibias.n523 3.19744
R23272 commonsourceibias.n139 commonsourceibias.t47 2.82907
R23273 commonsourceibias.n139 commonsourceibias.t79 2.82907
R23274 commonsourceibias.n140 commonsourceibias.t55 2.82907
R23275 commonsourceibias.n140 commonsourceibias.t5 2.82907
R23276 commonsourceibias.n142 commonsourceibias.t19 2.82907
R23277 commonsourceibias.n142 commonsourceibias.t23 2.82907
R23278 commonsourceibias.n144 commonsourceibias.t39 2.82907
R23279 commonsourceibias.n144 commonsourceibias.t71 2.82907
R23280 commonsourceibias.n146 commonsourceibias.t57 2.82907
R23281 commonsourceibias.n146 commonsourceibias.t27 2.82907
R23282 commonsourceibias.n137 commonsourceibias.t11 2.82907
R23283 commonsourceibias.n137 commonsourceibias.t41 2.82907
R23284 commonsourceibias.n135 commonsourceibias.t25 2.82907
R23285 commonsourceibias.n135 commonsourceibias.t35 2.82907
R23286 commonsourceibias.n133 commonsourceibias.t37 2.82907
R23287 commonsourceibias.n133 commonsourceibias.t77 2.82907
R23288 commonsourceibias.n131 commonsourceibias.t51 2.82907
R23289 commonsourceibias.n131 commonsourceibias.t9 2.82907
R23290 commonsourceibias.n129 commonsourceibias.t75 2.82907
R23291 commonsourceibias.n129 commonsourceibias.t21 2.82907
R23292 commonsourceibias.n503 commonsourceibias.t43 2.82907
R23293 commonsourceibias.n503 commonsourceibias.t15 2.82907
R23294 commonsourceibias.n505 commonsourceibias.t31 2.82907
R23295 commonsourceibias.n505 commonsourceibias.t1 2.82907
R23296 commonsourceibias.n507 commonsourceibias.t17 2.82907
R23297 commonsourceibias.n507 commonsourceibias.t61 2.82907
R23298 commonsourceibias.n509 commonsourceibias.t59 2.82907
R23299 commonsourceibias.n509 commonsourceibias.t45 2.82907
R23300 commonsourceibias.n511 commonsourceibias.t65 2.82907
R23301 commonsourceibias.n511 commonsourceibias.t33 2.82907
R23302 commonsourceibias.n386 commonsourceibias.t53 2.82907
R23303 commonsourceibias.n386 commonsourceibias.t73 2.82907
R23304 commonsourceibias.n384 commonsourceibias.t7 2.82907
R23305 commonsourceibias.n384 commonsourceibias.t63 2.82907
R23306 commonsourceibias.n382 commonsourceibias.t69 2.82907
R23307 commonsourceibias.n382 commonsourceibias.t67 2.82907
R23308 commonsourceibias.n380 commonsourceibias.t49 2.82907
R23309 commonsourceibias.n380 commonsourceibias.t13 2.82907
R23310 commonsourceibias.n379 commonsourceibias.t29 2.82907
R23311 commonsourceibias.n379 commonsourceibias.t3 2.82907
R23312 commonsourceibias.n280 commonsourceibias.n279 2.7056
R23313 commonsourceibias.n362 commonsourceibias.n361 2.7056
R23314 commonsourceibias.n125 commonsourceibias.n124 2.7056
R23315 commonsourceibias.n43 commonsourceibias.n42 2.7056
R23316 commonsourceibias.n247 commonsourceibias.n246 2.7056
R23317 commonsourceibias.n165 commonsourceibias.n164 2.7056
R23318 commonsourceibias.n642 commonsourceibias.n641 2.7056
R23319 commonsourceibias.n729 commonsourceibias.n728 2.7056
R23320 commonsourceibias.n412 commonsourceibias.n411 2.7056
R23321 commonsourceibias.n499 commonsourceibias.n498 2.7056
R23322 commonsourceibias.n614 commonsourceibias.n613 2.7056
R23323 commonsourceibias.n528 commonsourceibias.n527 2.7056
R23324 commonsourceibias.n132 commonsourceibias.n130 0.573776
R23325 commonsourceibias.n134 commonsourceibias.n132 0.573776
R23326 commonsourceibias.n136 commonsourceibias.n134 0.573776
R23327 commonsourceibias.n138 commonsourceibias.n136 0.573776
R23328 commonsourceibias.n147 commonsourceibias.n145 0.573776
R23329 commonsourceibias.n145 commonsourceibias.n143 0.573776
R23330 commonsourceibias.n143 commonsourceibias.n141 0.573776
R23331 commonsourceibias.n383 commonsourceibias.n381 0.573776
R23332 commonsourceibias.n385 commonsourceibias.n383 0.573776
R23333 commonsourceibias.n387 commonsourceibias.n385 0.573776
R23334 commonsourceibias.n512 commonsourceibias.n510 0.573776
R23335 commonsourceibias.n510 commonsourceibias.n508 0.573776
R23336 commonsourceibias.n508 commonsourceibias.n506 0.573776
R23337 commonsourceibias.n506 commonsourceibias.n504 0.573776
R23338 commonsourceibias.n148 commonsourceibias.n138 0.287138
R23339 commonsourceibias.n148 commonsourceibias.n147 0.287138
R23340 commonsourceibias.n513 commonsourceibias.n387 0.287138
R23341 commonsourceibias.n513 commonsourceibias.n512 0.287138
R23342 commonsourceibias.n365 commonsourceibias.n251 0.285035
R23343 commonsourceibias.n128 commonsourceibias.n14 0.285035
R23344 commonsourceibias.n250 commonsourceibias.n0 0.285035
R23345 commonsourceibias.n732 commonsourceibias.n618 0.285035
R23346 commonsourceibias.n502 commonsourceibias.n388 0.285035
R23347 commonsourceibias.n617 commonsourceibias.n367 0.285035
R23348 commonsourceibias.n360 commonsourceibias.n251 0.189894
R23349 commonsourceibias.n360 commonsourceibias.n359 0.189894
R23350 commonsourceibias.n359 commonsourceibias.n358 0.189894
R23351 commonsourceibias.n358 commonsourceibias.n253 0.189894
R23352 commonsourceibias.n353 commonsourceibias.n253 0.189894
R23353 commonsourceibias.n353 commonsourceibias.n352 0.189894
R23354 commonsourceibias.n352 commonsourceibias.n351 0.189894
R23355 commonsourceibias.n351 commonsourceibias.n255 0.189894
R23356 commonsourceibias.n346 commonsourceibias.n255 0.189894
R23357 commonsourceibias.n346 commonsourceibias.n345 0.189894
R23358 commonsourceibias.n345 commonsourceibias.n344 0.189894
R23359 commonsourceibias.n344 commonsourceibias.n258 0.189894
R23360 commonsourceibias.n339 commonsourceibias.n258 0.189894
R23361 commonsourceibias.n339 commonsourceibias.n338 0.189894
R23362 commonsourceibias.n338 commonsourceibias.n337 0.189894
R23363 commonsourceibias.n337 commonsourceibias.n260 0.189894
R23364 commonsourceibias.n332 commonsourceibias.n260 0.189894
R23365 commonsourceibias.n332 commonsourceibias.n331 0.189894
R23366 commonsourceibias.n331 commonsourceibias.n330 0.189894
R23367 commonsourceibias.n330 commonsourceibias.n263 0.189894
R23368 commonsourceibias.n325 commonsourceibias.n263 0.189894
R23369 commonsourceibias.n325 commonsourceibias.n324 0.189894
R23370 commonsourceibias.n324 commonsourceibias.n323 0.189894
R23371 commonsourceibias.n323 commonsourceibias.n265 0.189894
R23372 commonsourceibias.n318 commonsourceibias.n265 0.189894
R23373 commonsourceibias.n318 commonsourceibias.n317 0.189894
R23374 commonsourceibias.n317 commonsourceibias.n316 0.189894
R23375 commonsourceibias.n316 commonsourceibias.n268 0.189894
R23376 commonsourceibias.n311 commonsourceibias.n268 0.189894
R23377 commonsourceibias.n311 commonsourceibias.n310 0.189894
R23378 commonsourceibias.n310 commonsourceibias.n309 0.189894
R23379 commonsourceibias.n309 commonsourceibias.n270 0.189894
R23380 commonsourceibias.n304 commonsourceibias.n270 0.189894
R23381 commonsourceibias.n304 commonsourceibias.n303 0.189894
R23382 commonsourceibias.n303 commonsourceibias.n302 0.189894
R23383 commonsourceibias.n302 commonsourceibias.n273 0.189894
R23384 commonsourceibias.n297 commonsourceibias.n273 0.189894
R23385 commonsourceibias.n297 commonsourceibias.n296 0.189894
R23386 commonsourceibias.n296 commonsourceibias.n295 0.189894
R23387 commonsourceibias.n295 commonsourceibias.n275 0.189894
R23388 commonsourceibias.n290 commonsourceibias.n275 0.189894
R23389 commonsourceibias.n290 commonsourceibias.n289 0.189894
R23390 commonsourceibias.n289 commonsourceibias.n288 0.189894
R23391 commonsourceibias.n288 commonsourceibias.n278 0.189894
R23392 commonsourceibias.n283 commonsourceibias.n278 0.189894
R23393 commonsourceibias.n283 commonsourceibias.n282 0.189894
R23394 commonsourceibias.n123 commonsourceibias.n14 0.189894
R23395 commonsourceibias.n123 commonsourceibias.n122 0.189894
R23396 commonsourceibias.n122 commonsourceibias.n121 0.189894
R23397 commonsourceibias.n121 commonsourceibias.n16 0.189894
R23398 commonsourceibias.n116 commonsourceibias.n16 0.189894
R23399 commonsourceibias.n116 commonsourceibias.n115 0.189894
R23400 commonsourceibias.n115 commonsourceibias.n114 0.189894
R23401 commonsourceibias.n114 commonsourceibias.n18 0.189894
R23402 commonsourceibias.n109 commonsourceibias.n18 0.189894
R23403 commonsourceibias.n109 commonsourceibias.n108 0.189894
R23404 commonsourceibias.n108 commonsourceibias.n107 0.189894
R23405 commonsourceibias.n107 commonsourceibias.n21 0.189894
R23406 commonsourceibias.n102 commonsourceibias.n21 0.189894
R23407 commonsourceibias.n102 commonsourceibias.n101 0.189894
R23408 commonsourceibias.n101 commonsourceibias.n100 0.189894
R23409 commonsourceibias.n100 commonsourceibias.n23 0.189894
R23410 commonsourceibias.n95 commonsourceibias.n23 0.189894
R23411 commonsourceibias.n95 commonsourceibias.n94 0.189894
R23412 commonsourceibias.n94 commonsourceibias.n93 0.189894
R23413 commonsourceibias.n93 commonsourceibias.n26 0.189894
R23414 commonsourceibias.n88 commonsourceibias.n26 0.189894
R23415 commonsourceibias.n88 commonsourceibias.n87 0.189894
R23416 commonsourceibias.n87 commonsourceibias.n86 0.189894
R23417 commonsourceibias.n86 commonsourceibias.n28 0.189894
R23418 commonsourceibias.n81 commonsourceibias.n28 0.189894
R23419 commonsourceibias.n81 commonsourceibias.n80 0.189894
R23420 commonsourceibias.n80 commonsourceibias.n79 0.189894
R23421 commonsourceibias.n79 commonsourceibias.n31 0.189894
R23422 commonsourceibias.n74 commonsourceibias.n31 0.189894
R23423 commonsourceibias.n74 commonsourceibias.n73 0.189894
R23424 commonsourceibias.n73 commonsourceibias.n72 0.189894
R23425 commonsourceibias.n72 commonsourceibias.n33 0.189894
R23426 commonsourceibias.n67 commonsourceibias.n33 0.189894
R23427 commonsourceibias.n67 commonsourceibias.n66 0.189894
R23428 commonsourceibias.n66 commonsourceibias.n65 0.189894
R23429 commonsourceibias.n65 commonsourceibias.n36 0.189894
R23430 commonsourceibias.n60 commonsourceibias.n36 0.189894
R23431 commonsourceibias.n60 commonsourceibias.n59 0.189894
R23432 commonsourceibias.n59 commonsourceibias.n58 0.189894
R23433 commonsourceibias.n58 commonsourceibias.n38 0.189894
R23434 commonsourceibias.n53 commonsourceibias.n38 0.189894
R23435 commonsourceibias.n53 commonsourceibias.n52 0.189894
R23436 commonsourceibias.n52 commonsourceibias.n51 0.189894
R23437 commonsourceibias.n51 commonsourceibias.n41 0.189894
R23438 commonsourceibias.n46 commonsourceibias.n41 0.189894
R23439 commonsourceibias.n46 commonsourceibias.n45 0.189894
R23440 commonsourceibias.n205 commonsourceibias.n204 0.189894
R23441 commonsourceibias.n204 commonsourceibias.n152 0.189894
R23442 commonsourceibias.n200 commonsourceibias.n152 0.189894
R23443 commonsourceibias.n200 commonsourceibias.n199 0.189894
R23444 commonsourceibias.n199 commonsourceibias.n154 0.189894
R23445 commonsourceibias.n195 commonsourceibias.n154 0.189894
R23446 commonsourceibias.n195 commonsourceibias.n194 0.189894
R23447 commonsourceibias.n194 commonsourceibias.n156 0.189894
R23448 commonsourceibias.n189 commonsourceibias.n156 0.189894
R23449 commonsourceibias.n189 commonsourceibias.n188 0.189894
R23450 commonsourceibias.n188 commonsourceibias.n187 0.189894
R23451 commonsourceibias.n187 commonsourceibias.n158 0.189894
R23452 commonsourceibias.n182 commonsourceibias.n158 0.189894
R23453 commonsourceibias.n182 commonsourceibias.n181 0.189894
R23454 commonsourceibias.n181 commonsourceibias.n180 0.189894
R23455 commonsourceibias.n180 commonsourceibias.n160 0.189894
R23456 commonsourceibias.n175 commonsourceibias.n160 0.189894
R23457 commonsourceibias.n175 commonsourceibias.n174 0.189894
R23458 commonsourceibias.n174 commonsourceibias.n173 0.189894
R23459 commonsourceibias.n173 commonsourceibias.n163 0.189894
R23460 commonsourceibias.n168 commonsourceibias.n163 0.189894
R23461 commonsourceibias.n168 commonsourceibias.n167 0.189894
R23462 commonsourceibias.n245 commonsourceibias.n0 0.189894
R23463 commonsourceibias.n245 commonsourceibias.n244 0.189894
R23464 commonsourceibias.n244 commonsourceibias.n243 0.189894
R23465 commonsourceibias.n243 commonsourceibias.n2 0.189894
R23466 commonsourceibias.n238 commonsourceibias.n2 0.189894
R23467 commonsourceibias.n238 commonsourceibias.n237 0.189894
R23468 commonsourceibias.n237 commonsourceibias.n236 0.189894
R23469 commonsourceibias.n236 commonsourceibias.n4 0.189894
R23470 commonsourceibias.n231 commonsourceibias.n4 0.189894
R23471 commonsourceibias.n231 commonsourceibias.n230 0.189894
R23472 commonsourceibias.n230 commonsourceibias.n229 0.189894
R23473 commonsourceibias.n229 commonsourceibias.n7 0.189894
R23474 commonsourceibias.n224 commonsourceibias.n7 0.189894
R23475 commonsourceibias.n224 commonsourceibias.n223 0.189894
R23476 commonsourceibias.n223 commonsourceibias.n222 0.189894
R23477 commonsourceibias.n222 commonsourceibias.n9 0.189894
R23478 commonsourceibias.n217 commonsourceibias.n9 0.189894
R23479 commonsourceibias.n217 commonsourceibias.n216 0.189894
R23480 commonsourceibias.n216 commonsourceibias.n215 0.189894
R23481 commonsourceibias.n215 commonsourceibias.n12 0.189894
R23482 commonsourceibias.n210 commonsourceibias.n12 0.189894
R23483 commonsourceibias.n210 commonsourceibias.n209 0.189894
R23484 commonsourceibias.n209 commonsourceibias.n208 0.189894
R23485 commonsourceibias.n645 commonsourceibias.n644 0.189894
R23486 commonsourceibias.n645 commonsourceibias.n640 0.189894
R23487 commonsourceibias.n650 commonsourceibias.n640 0.189894
R23488 commonsourceibias.n651 commonsourceibias.n650 0.189894
R23489 commonsourceibias.n652 commonsourceibias.n651 0.189894
R23490 commonsourceibias.n652 commonsourceibias.n638 0.189894
R23491 commonsourceibias.n658 commonsourceibias.n638 0.189894
R23492 commonsourceibias.n659 commonsourceibias.n658 0.189894
R23493 commonsourceibias.n660 commonsourceibias.n659 0.189894
R23494 commonsourceibias.n660 commonsourceibias.n636 0.189894
R23495 commonsourceibias.n665 commonsourceibias.n636 0.189894
R23496 commonsourceibias.n666 commonsourceibias.n665 0.189894
R23497 commonsourceibias.n667 commonsourceibias.n666 0.189894
R23498 commonsourceibias.n667 commonsourceibias.n634 0.189894
R23499 commonsourceibias.n673 commonsourceibias.n634 0.189894
R23500 commonsourceibias.n674 commonsourceibias.n673 0.189894
R23501 commonsourceibias.n675 commonsourceibias.n674 0.189894
R23502 commonsourceibias.n675 commonsourceibias.n632 0.189894
R23503 commonsourceibias.n680 commonsourceibias.n632 0.189894
R23504 commonsourceibias.n681 commonsourceibias.n680 0.189894
R23505 commonsourceibias.n682 commonsourceibias.n681 0.189894
R23506 commonsourceibias.n682 commonsourceibias.n630 0.189894
R23507 commonsourceibias.n688 commonsourceibias.n630 0.189894
R23508 commonsourceibias.n689 commonsourceibias.n688 0.189894
R23509 commonsourceibias.n690 commonsourceibias.n689 0.189894
R23510 commonsourceibias.n690 commonsourceibias.n628 0.189894
R23511 commonsourceibias.n695 commonsourceibias.n628 0.189894
R23512 commonsourceibias.n696 commonsourceibias.n695 0.189894
R23513 commonsourceibias.n697 commonsourceibias.n696 0.189894
R23514 commonsourceibias.n697 commonsourceibias.n626 0.189894
R23515 commonsourceibias.n703 commonsourceibias.n626 0.189894
R23516 commonsourceibias.n704 commonsourceibias.n703 0.189894
R23517 commonsourceibias.n705 commonsourceibias.n704 0.189894
R23518 commonsourceibias.n705 commonsourceibias.n624 0.189894
R23519 commonsourceibias.n710 commonsourceibias.n624 0.189894
R23520 commonsourceibias.n711 commonsourceibias.n710 0.189894
R23521 commonsourceibias.n712 commonsourceibias.n711 0.189894
R23522 commonsourceibias.n712 commonsourceibias.n622 0.189894
R23523 commonsourceibias.n718 commonsourceibias.n622 0.189894
R23524 commonsourceibias.n719 commonsourceibias.n718 0.189894
R23525 commonsourceibias.n720 commonsourceibias.n719 0.189894
R23526 commonsourceibias.n720 commonsourceibias.n620 0.189894
R23527 commonsourceibias.n725 commonsourceibias.n620 0.189894
R23528 commonsourceibias.n726 commonsourceibias.n725 0.189894
R23529 commonsourceibias.n727 commonsourceibias.n726 0.189894
R23530 commonsourceibias.n727 commonsourceibias.n618 0.189894
R23531 commonsourceibias.n415 commonsourceibias.n414 0.189894
R23532 commonsourceibias.n415 commonsourceibias.n410 0.189894
R23533 commonsourceibias.n420 commonsourceibias.n410 0.189894
R23534 commonsourceibias.n421 commonsourceibias.n420 0.189894
R23535 commonsourceibias.n422 commonsourceibias.n421 0.189894
R23536 commonsourceibias.n422 commonsourceibias.n408 0.189894
R23537 commonsourceibias.n428 commonsourceibias.n408 0.189894
R23538 commonsourceibias.n429 commonsourceibias.n428 0.189894
R23539 commonsourceibias.n430 commonsourceibias.n429 0.189894
R23540 commonsourceibias.n430 commonsourceibias.n406 0.189894
R23541 commonsourceibias.n435 commonsourceibias.n406 0.189894
R23542 commonsourceibias.n436 commonsourceibias.n435 0.189894
R23543 commonsourceibias.n437 commonsourceibias.n436 0.189894
R23544 commonsourceibias.n437 commonsourceibias.n404 0.189894
R23545 commonsourceibias.n443 commonsourceibias.n404 0.189894
R23546 commonsourceibias.n444 commonsourceibias.n443 0.189894
R23547 commonsourceibias.n445 commonsourceibias.n444 0.189894
R23548 commonsourceibias.n445 commonsourceibias.n402 0.189894
R23549 commonsourceibias.n450 commonsourceibias.n402 0.189894
R23550 commonsourceibias.n451 commonsourceibias.n450 0.189894
R23551 commonsourceibias.n452 commonsourceibias.n451 0.189894
R23552 commonsourceibias.n452 commonsourceibias.n400 0.189894
R23553 commonsourceibias.n458 commonsourceibias.n400 0.189894
R23554 commonsourceibias.n459 commonsourceibias.n458 0.189894
R23555 commonsourceibias.n460 commonsourceibias.n459 0.189894
R23556 commonsourceibias.n460 commonsourceibias.n398 0.189894
R23557 commonsourceibias.n465 commonsourceibias.n398 0.189894
R23558 commonsourceibias.n466 commonsourceibias.n465 0.189894
R23559 commonsourceibias.n467 commonsourceibias.n466 0.189894
R23560 commonsourceibias.n467 commonsourceibias.n396 0.189894
R23561 commonsourceibias.n473 commonsourceibias.n396 0.189894
R23562 commonsourceibias.n474 commonsourceibias.n473 0.189894
R23563 commonsourceibias.n475 commonsourceibias.n474 0.189894
R23564 commonsourceibias.n475 commonsourceibias.n394 0.189894
R23565 commonsourceibias.n480 commonsourceibias.n394 0.189894
R23566 commonsourceibias.n481 commonsourceibias.n480 0.189894
R23567 commonsourceibias.n482 commonsourceibias.n481 0.189894
R23568 commonsourceibias.n482 commonsourceibias.n392 0.189894
R23569 commonsourceibias.n488 commonsourceibias.n392 0.189894
R23570 commonsourceibias.n489 commonsourceibias.n488 0.189894
R23571 commonsourceibias.n490 commonsourceibias.n489 0.189894
R23572 commonsourceibias.n490 commonsourceibias.n390 0.189894
R23573 commonsourceibias.n495 commonsourceibias.n390 0.189894
R23574 commonsourceibias.n496 commonsourceibias.n495 0.189894
R23575 commonsourceibias.n497 commonsourceibias.n496 0.189894
R23576 commonsourceibias.n497 commonsourceibias.n388 0.189894
R23577 commonsourceibias.n531 commonsourceibias.n530 0.189894
R23578 commonsourceibias.n531 commonsourceibias.n526 0.189894
R23579 commonsourceibias.n536 commonsourceibias.n526 0.189894
R23580 commonsourceibias.n537 commonsourceibias.n536 0.189894
R23581 commonsourceibias.n538 commonsourceibias.n537 0.189894
R23582 commonsourceibias.n538 commonsourceibias.n524 0.189894
R23583 commonsourceibias.n544 commonsourceibias.n524 0.189894
R23584 commonsourceibias.n545 commonsourceibias.n544 0.189894
R23585 commonsourceibias.n546 commonsourceibias.n545 0.189894
R23586 commonsourceibias.n546 commonsourceibias.n522 0.189894
R23587 commonsourceibias.n551 commonsourceibias.n522 0.189894
R23588 commonsourceibias.n552 commonsourceibias.n551 0.189894
R23589 commonsourceibias.n553 commonsourceibias.n552 0.189894
R23590 commonsourceibias.n553 commonsourceibias.n520 0.189894
R23591 commonsourceibias.n558 commonsourceibias.n520 0.189894
R23592 commonsourceibias.n559 commonsourceibias.n558 0.189894
R23593 commonsourceibias.n559 commonsourceibias.n518 0.189894
R23594 commonsourceibias.n563 commonsourceibias.n518 0.189894
R23595 commonsourceibias.n564 commonsourceibias.n563 0.189894
R23596 commonsourceibias.n564 commonsourceibias.n516 0.189894
R23597 commonsourceibias.n568 commonsourceibias.n516 0.189894
R23598 commonsourceibias.n569 commonsourceibias.n568 0.189894
R23599 commonsourceibias.n574 commonsourceibias.n573 0.189894
R23600 commonsourceibias.n575 commonsourceibias.n574 0.189894
R23601 commonsourceibias.n575 commonsourceibias.n377 0.189894
R23602 commonsourceibias.n580 commonsourceibias.n377 0.189894
R23603 commonsourceibias.n581 commonsourceibias.n580 0.189894
R23604 commonsourceibias.n582 commonsourceibias.n581 0.189894
R23605 commonsourceibias.n582 commonsourceibias.n375 0.189894
R23606 commonsourceibias.n588 commonsourceibias.n375 0.189894
R23607 commonsourceibias.n589 commonsourceibias.n588 0.189894
R23608 commonsourceibias.n590 commonsourceibias.n589 0.189894
R23609 commonsourceibias.n590 commonsourceibias.n373 0.189894
R23610 commonsourceibias.n595 commonsourceibias.n373 0.189894
R23611 commonsourceibias.n596 commonsourceibias.n595 0.189894
R23612 commonsourceibias.n597 commonsourceibias.n596 0.189894
R23613 commonsourceibias.n597 commonsourceibias.n371 0.189894
R23614 commonsourceibias.n603 commonsourceibias.n371 0.189894
R23615 commonsourceibias.n604 commonsourceibias.n603 0.189894
R23616 commonsourceibias.n605 commonsourceibias.n604 0.189894
R23617 commonsourceibias.n605 commonsourceibias.n369 0.189894
R23618 commonsourceibias.n610 commonsourceibias.n369 0.189894
R23619 commonsourceibias.n611 commonsourceibias.n610 0.189894
R23620 commonsourceibias.n612 commonsourceibias.n611 0.189894
R23621 commonsourceibias.n612 commonsourceibias.n367 0.189894
R23622 commonsourceibias.n205 commonsourceibias.n149 0.0762576
R23623 commonsourceibias.n208 commonsourceibias.n149 0.0762576
R23624 commonsourceibias.n569 commonsourceibias.n514 0.0762576
R23625 commonsourceibias.n573 commonsourceibias.n514 0.0762576
R23626 minus.n43 minus.t24 322.512
R23627 minus.n9 minus.t8 322.512
R23628 minus.n66 minus.t5 297.12
R23629 minus.n64 minus.t6 297.12
R23630 minus.n36 minus.t22 297.12
R23631 minus.n58 minus.t18 297.12
R23632 minus.n38 minus.t19 297.12
R23633 minus.n52 minus.t14 297.12
R23634 minus.n40 minus.t15 297.12
R23635 minus.n46 minus.t9 297.12
R23636 minus.n42 minus.t23 297.12
R23637 minus.n8 minus.t7 297.12
R23638 minus.n12 minus.t11 297.12
R23639 minus.n14 minus.t10 297.12
R23640 minus.n18 minus.t12 297.12
R23641 minus.n20 minus.t17 297.12
R23642 minus.n24 minus.t16 297.12
R23643 minus.n26 minus.t21 297.12
R23644 minus.n30 minus.t20 297.12
R23645 minus.n32 minus.t13 297.12
R23646 minus.n72 minus.t4 243.255
R23647 minus.n71 minus.n69 224.169
R23648 minus.n71 minus.n70 223.454
R23649 minus.n45 minus.n44 161.3
R23650 minus.n46 minus.n41 161.3
R23651 minus.n48 minus.n47 161.3
R23652 minus.n49 minus.n40 161.3
R23653 minus.n51 minus.n50 161.3
R23654 minus.n52 minus.n39 161.3
R23655 minus.n54 minus.n53 161.3
R23656 minus.n55 minus.n38 161.3
R23657 minus.n57 minus.n56 161.3
R23658 minus.n58 minus.n37 161.3
R23659 minus.n60 minus.n59 161.3
R23660 minus.n61 minus.n36 161.3
R23661 minus.n63 minus.n62 161.3
R23662 minus.n64 minus.n35 161.3
R23663 minus.n65 minus.n34 161.3
R23664 minus.n67 minus.n66 161.3
R23665 minus.n33 minus.n32 161.3
R23666 minus.n31 minus.n0 161.3
R23667 minus.n30 minus.n29 161.3
R23668 minus.n28 minus.n1 161.3
R23669 minus.n27 minus.n26 161.3
R23670 minus.n25 minus.n2 161.3
R23671 minus.n24 minus.n23 161.3
R23672 minus.n22 minus.n3 161.3
R23673 minus.n21 minus.n20 161.3
R23674 minus.n19 minus.n4 161.3
R23675 minus.n18 minus.n17 161.3
R23676 minus.n16 minus.n5 161.3
R23677 minus.n15 minus.n14 161.3
R23678 minus.n13 minus.n6 161.3
R23679 minus.n12 minus.n11 161.3
R23680 minus.n10 minus.n7 161.3
R23681 minus.n44 minus.n43 45.0031
R23682 minus.n10 minus.n9 45.0031
R23683 minus.n66 minus.n65 41.6278
R23684 minus.n32 minus.n31 41.6278
R23685 minus.n64 minus.n63 37.246
R23686 minus.n45 minus.n42 37.246
R23687 minus.n8 minus.n7 37.246
R23688 minus.n30 minus.n1 37.246
R23689 minus.n59 minus.n36 32.8641
R23690 minus.n47 minus.n46 32.8641
R23691 minus.n13 minus.n12 32.8641
R23692 minus.n26 minus.n25 32.8641
R23693 minus.n68 minus.n67 31.8206
R23694 minus.n58 minus.n57 28.4823
R23695 minus.n51 minus.n40 28.4823
R23696 minus.n14 minus.n5 28.4823
R23697 minus.n24 minus.n3 28.4823
R23698 minus.n53 minus.n38 24.1005
R23699 minus.n53 minus.n52 24.1005
R23700 minus.n19 minus.n18 24.1005
R23701 minus.n20 minus.n19 24.1005
R23702 minus.n70 minus.t3 19.8005
R23703 minus.n70 minus.t1 19.8005
R23704 minus.n69 minus.t2 19.8005
R23705 minus.n69 minus.t0 19.8005
R23706 minus.n57 minus.n38 19.7187
R23707 minus.n52 minus.n51 19.7187
R23708 minus.n18 minus.n5 19.7187
R23709 minus.n20 minus.n3 19.7187
R23710 minus.n43 minus.n42 15.6319
R23711 minus.n9 minus.n8 15.6319
R23712 minus.n59 minus.n58 15.3369
R23713 minus.n47 minus.n40 15.3369
R23714 minus.n14 minus.n13 15.3369
R23715 minus.n25 minus.n24 15.3369
R23716 minus minus.n73 12.1618
R23717 minus.n68 minus.n33 12.0819
R23718 minus.n63 minus.n36 10.955
R23719 minus.n46 minus.n45 10.955
R23720 minus.n12 minus.n7 10.955
R23721 minus.n26 minus.n1 10.955
R23722 minus.n65 minus.n64 6.57323
R23723 minus.n31 minus.n30 6.57323
R23724 minus.n73 minus.n72 4.80222
R23725 minus.n73 minus.n68 0.972091
R23726 minus.n72 minus.n71 0.716017
R23727 minus.n67 minus.n34 0.189894
R23728 minus.n35 minus.n34 0.189894
R23729 minus.n62 minus.n35 0.189894
R23730 minus.n62 minus.n61 0.189894
R23731 minus.n61 minus.n60 0.189894
R23732 minus.n60 minus.n37 0.189894
R23733 minus.n56 minus.n37 0.189894
R23734 minus.n56 minus.n55 0.189894
R23735 minus.n55 minus.n54 0.189894
R23736 minus.n54 minus.n39 0.189894
R23737 minus.n50 minus.n39 0.189894
R23738 minus.n50 minus.n49 0.189894
R23739 minus.n49 minus.n48 0.189894
R23740 minus.n48 minus.n41 0.189894
R23741 minus.n44 minus.n41 0.189894
R23742 minus.n11 minus.n10 0.189894
R23743 minus.n11 minus.n6 0.189894
R23744 minus.n15 minus.n6 0.189894
R23745 minus.n16 minus.n15 0.189894
R23746 minus.n17 minus.n16 0.189894
R23747 minus.n17 minus.n4 0.189894
R23748 minus.n21 minus.n4 0.189894
R23749 minus.n22 minus.n21 0.189894
R23750 minus.n23 minus.n22 0.189894
R23751 minus.n23 minus.n2 0.189894
R23752 minus.n27 minus.n2 0.189894
R23753 minus.n28 minus.n27 0.189894
R23754 minus.n29 minus.n28 0.189894
R23755 minus.n29 minus.n0 0.189894
R23756 minus.n33 minus.n0 0.189894
R23757 output.n41 output.n15 289.615
R23758 output.n72 output.n46 289.615
R23759 output.n104 output.n78 289.615
R23760 output.n136 output.n110 289.615
R23761 output.n77 output.n45 197.26
R23762 output.n77 output.n76 196.298
R23763 output.n109 output.n108 196.298
R23764 output.n141 output.n140 196.298
R23765 output.n42 output.n41 185
R23766 output.n40 output.n39 185
R23767 output.n19 output.n18 185
R23768 output.n34 output.n33 185
R23769 output.n32 output.n31 185
R23770 output.n23 output.n22 185
R23771 output.n26 output.n25 185
R23772 output.n73 output.n72 185
R23773 output.n71 output.n70 185
R23774 output.n50 output.n49 185
R23775 output.n65 output.n64 185
R23776 output.n63 output.n62 185
R23777 output.n54 output.n53 185
R23778 output.n57 output.n56 185
R23779 output.n105 output.n104 185
R23780 output.n103 output.n102 185
R23781 output.n82 output.n81 185
R23782 output.n97 output.n96 185
R23783 output.n95 output.n94 185
R23784 output.n86 output.n85 185
R23785 output.n89 output.n88 185
R23786 output.n137 output.n136 185
R23787 output.n135 output.n134 185
R23788 output.n114 output.n113 185
R23789 output.n129 output.n128 185
R23790 output.n127 output.n126 185
R23791 output.n118 output.n117 185
R23792 output.n121 output.n120 185
R23793 output.t3 output.n24 147.661
R23794 output.t1 output.n55 147.661
R23795 output.t2 output.n87 147.661
R23796 output.t0 output.n119 147.661
R23797 output.n41 output.n40 104.615
R23798 output.n40 output.n18 104.615
R23799 output.n33 output.n18 104.615
R23800 output.n33 output.n32 104.615
R23801 output.n32 output.n22 104.615
R23802 output.n25 output.n22 104.615
R23803 output.n72 output.n71 104.615
R23804 output.n71 output.n49 104.615
R23805 output.n64 output.n49 104.615
R23806 output.n64 output.n63 104.615
R23807 output.n63 output.n53 104.615
R23808 output.n56 output.n53 104.615
R23809 output.n104 output.n103 104.615
R23810 output.n103 output.n81 104.615
R23811 output.n96 output.n81 104.615
R23812 output.n96 output.n95 104.615
R23813 output.n95 output.n85 104.615
R23814 output.n88 output.n85 104.615
R23815 output.n136 output.n135 104.615
R23816 output.n135 output.n113 104.615
R23817 output.n128 output.n113 104.615
R23818 output.n128 output.n127 104.615
R23819 output.n127 output.n117 104.615
R23820 output.n120 output.n117 104.615
R23821 output.n1 output.t13 77.056
R23822 output.n14 output.t15 76.6694
R23823 output.n1 output.n0 72.7095
R23824 output.n3 output.n2 72.7095
R23825 output.n5 output.n4 72.7095
R23826 output.n7 output.n6 72.7095
R23827 output.n9 output.n8 72.7095
R23828 output.n11 output.n10 72.7095
R23829 output.n13 output.n12 72.7095
R23830 output.n25 output.t3 52.3082
R23831 output.n56 output.t1 52.3082
R23832 output.n88 output.t2 52.3082
R23833 output.n120 output.t0 52.3082
R23834 output.n26 output.n24 15.6674
R23835 output.n57 output.n55 15.6674
R23836 output.n89 output.n87 15.6674
R23837 output.n121 output.n119 15.6674
R23838 output.n27 output.n23 12.8005
R23839 output.n58 output.n54 12.8005
R23840 output.n90 output.n86 12.8005
R23841 output.n122 output.n118 12.8005
R23842 output.n31 output.n30 12.0247
R23843 output.n62 output.n61 12.0247
R23844 output.n94 output.n93 12.0247
R23845 output.n126 output.n125 12.0247
R23846 output.n34 output.n21 11.249
R23847 output.n65 output.n52 11.249
R23848 output.n97 output.n84 11.249
R23849 output.n129 output.n116 11.249
R23850 output.n35 output.n19 10.4732
R23851 output.n66 output.n50 10.4732
R23852 output.n98 output.n82 10.4732
R23853 output.n130 output.n114 10.4732
R23854 output.n39 output.n38 9.69747
R23855 output.n70 output.n69 9.69747
R23856 output.n102 output.n101 9.69747
R23857 output.n134 output.n133 9.69747
R23858 output.n45 output.n44 9.45567
R23859 output.n76 output.n75 9.45567
R23860 output.n108 output.n107 9.45567
R23861 output.n140 output.n139 9.45567
R23862 output.n44 output.n43 9.3005
R23863 output.n17 output.n16 9.3005
R23864 output.n38 output.n37 9.3005
R23865 output.n36 output.n35 9.3005
R23866 output.n21 output.n20 9.3005
R23867 output.n30 output.n29 9.3005
R23868 output.n28 output.n27 9.3005
R23869 output.n75 output.n74 9.3005
R23870 output.n48 output.n47 9.3005
R23871 output.n69 output.n68 9.3005
R23872 output.n67 output.n66 9.3005
R23873 output.n52 output.n51 9.3005
R23874 output.n61 output.n60 9.3005
R23875 output.n59 output.n58 9.3005
R23876 output.n107 output.n106 9.3005
R23877 output.n80 output.n79 9.3005
R23878 output.n101 output.n100 9.3005
R23879 output.n99 output.n98 9.3005
R23880 output.n84 output.n83 9.3005
R23881 output.n93 output.n92 9.3005
R23882 output.n91 output.n90 9.3005
R23883 output.n139 output.n138 9.3005
R23884 output.n112 output.n111 9.3005
R23885 output.n133 output.n132 9.3005
R23886 output.n131 output.n130 9.3005
R23887 output.n116 output.n115 9.3005
R23888 output.n125 output.n124 9.3005
R23889 output.n123 output.n122 9.3005
R23890 output.n42 output.n17 8.92171
R23891 output.n73 output.n48 8.92171
R23892 output.n105 output.n80 8.92171
R23893 output.n137 output.n112 8.92171
R23894 output output.n141 8.15037
R23895 output.n43 output.n15 8.14595
R23896 output.n74 output.n46 8.14595
R23897 output.n106 output.n78 8.14595
R23898 output.n138 output.n110 8.14595
R23899 output.n45 output.n15 5.81868
R23900 output.n76 output.n46 5.81868
R23901 output.n108 output.n78 5.81868
R23902 output.n140 output.n110 5.81868
R23903 output.n43 output.n42 5.04292
R23904 output.n74 output.n73 5.04292
R23905 output.n106 output.n105 5.04292
R23906 output.n138 output.n137 5.04292
R23907 output.n28 output.n24 4.38594
R23908 output.n59 output.n55 4.38594
R23909 output.n91 output.n87 4.38594
R23910 output.n123 output.n119 4.38594
R23911 output.n39 output.n17 4.26717
R23912 output.n70 output.n48 4.26717
R23913 output.n102 output.n80 4.26717
R23914 output.n134 output.n112 4.26717
R23915 output.n0 output.t19 3.9605
R23916 output.n0 output.t8 3.9605
R23917 output.n2 output.t12 3.9605
R23918 output.n2 output.t4 3.9605
R23919 output.n4 output.t6 3.9605
R23920 output.n4 output.t5 3.9605
R23921 output.n6 output.t11 3.9605
R23922 output.n6 output.t14 3.9605
R23923 output.n8 output.t16 3.9605
R23924 output.n8 output.t9 3.9605
R23925 output.n10 output.t10 3.9605
R23926 output.n10 output.t17 3.9605
R23927 output.n12 output.t18 3.9605
R23928 output.n12 output.t7 3.9605
R23929 output.n38 output.n19 3.49141
R23930 output.n69 output.n50 3.49141
R23931 output.n101 output.n82 3.49141
R23932 output.n133 output.n114 3.49141
R23933 output.n35 output.n34 2.71565
R23934 output.n66 output.n65 2.71565
R23935 output.n98 output.n97 2.71565
R23936 output.n130 output.n129 2.71565
R23937 output.n31 output.n21 1.93989
R23938 output.n62 output.n52 1.93989
R23939 output.n94 output.n84 1.93989
R23940 output.n126 output.n116 1.93989
R23941 output.n30 output.n23 1.16414
R23942 output.n61 output.n54 1.16414
R23943 output.n93 output.n86 1.16414
R23944 output.n125 output.n118 1.16414
R23945 output.n141 output.n109 0.962709
R23946 output.n109 output.n77 0.962709
R23947 output.n27 output.n26 0.388379
R23948 output.n58 output.n57 0.388379
R23949 output.n90 output.n89 0.388379
R23950 output.n122 output.n121 0.388379
R23951 output.n14 output.n13 0.387128
R23952 output.n13 output.n11 0.387128
R23953 output.n11 output.n9 0.387128
R23954 output.n9 output.n7 0.387128
R23955 output.n7 output.n5 0.387128
R23956 output.n5 output.n3 0.387128
R23957 output.n3 output.n1 0.387128
R23958 output.n44 output.n16 0.155672
R23959 output.n37 output.n16 0.155672
R23960 output.n37 output.n36 0.155672
R23961 output.n36 output.n20 0.155672
R23962 output.n29 output.n20 0.155672
R23963 output.n29 output.n28 0.155672
R23964 output.n75 output.n47 0.155672
R23965 output.n68 output.n47 0.155672
R23966 output.n68 output.n67 0.155672
R23967 output.n67 output.n51 0.155672
R23968 output.n60 output.n51 0.155672
R23969 output.n60 output.n59 0.155672
R23970 output.n107 output.n79 0.155672
R23971 output.n100 output.n79 0.155672
R23972 output.n100 output.n99 0.155672
R23973 output.n99 output.n83 0.155672
R23974 output.n92 output.n83 0.155672
R23975 output.n92 output.n91 0.155672
R23976 output.n139 output.n111 0.155672
R23977 output.n132 output.n111 0.155672
R23978 output.n132 output.n131 0.155672
R23979 output.n131 output.n115 0.155672
R23980 output.n124 output.n115 0.155672
R23981 output.n124 output.n123 0.155672
R23982 output output.n14 0.126227
R23983 a_n2318_8322.n8 a_n2318_8322.t3 74.6477
R23984 a_n2318_8322.n1 a_n2318_8322.t22 74.6477
R23985 a_n2318_8322.n20 a_n2318_8322.t21 74.6474
R23986 a_n2318_8322.n16 a_n2318_8322.t11 74.2899
R23987 a_n2318_8322.n9 a_n2318_8322.t1 74.2899
R23988 a_n2318_8322.n10 a_n2318_8322.t4 74.2899
R23989 a_n2318_8322.n13 a_n2318_8322.t5 74.2899
R23990 a_n2318_8322.n6 a_n2318_8322.t8 74.2899
R23991 a_n2318_8322.n20 a_n2318_8322.n19 70.6783
R23992 a_n2318_8322.n18 a_n2318_8322.n17 70.6783
R23993 a_n2318_8322.n8 a_n2318_8322.n7 70.6783
R23994 a_n2318_8322.n12 a_n2318_8322.n11 70.6783
R23995 a_n2318_8322.n1 a_n2318_8322.n0 70.6783
R23996 a_n2318_8322.n3 a_n2318_8322.n2 70.6783
R23997 a_n2318_8322.n5 a_n2318_8322.n4 70.6783
R23998 a_n2318_8322.n22 a_n2318_8322.n21 70.6782
R23999 a_n2318_8322.n14 a_n2318_8322.n6 23.4712
R24000 a_n2318_8322.n15 a_n2318_8322.t24 10.1716
R24001 a_n2318_8322.n14 a_n2318_8322.n13 6.95632
R24002 a_n2318_8322.n16 a_n2318_8322.n15 6.19447
R24003 a_n2318_8322.n15 a_n2318_8322.n14 5.3452
R24004 a_n2318_8322.n19 a_n2318_8322.t18 3.61217
R24005 a_n2318_8322.n19 a_n2318_8322.t15 3.61217
R24006 a_n2318_8322.n17 a_n2318_8322.t20 3.61217
R24007 a_n2318_8322.n17 a_n2318_8322.t13 3.61217
R24008 a_n2318_8322.n7 a_n2318_8322.t7 3.61217
R24009 a_n2318_8322.n7 a_n2318_8322.t6 3.61217
R24010 a_n2318_8322.n11 a_n2318_8322.t2 3.61217
R24011 a_n2318_8322.n11 a_n2318_8322.t0 3.61217
R24012 a_n2318_8322.n0 a_n2318_8322.t10 3.61217
R24013 a_n2318_8322.n0 a_n2318_8322.t9 3.61217
R24014 a_n2318_8322.n2 a_n2318_8322.t19 3.61217
R24015 a_n2318_8322.n2 a_n2318_8322.t14 3.61217
R24016 a_n2318_8322.n4 a_n2318_8322.t17 3.61217
R24017 a_n2318_8322.n4 a_n2318_8322.t16 3.61217
R24018 a_n2318_8322.n22 a_n2318_8322.t12 3.61217
R24019 a_n2318_8322.t23 a_n2318_8322.n22 3.61217
R24020 a_n2318_8322.n13 a_n2318_8322.n12 0.358259
R24021 a_n2318_8322.n12 a_n2318_8322.n10 0.358259
R24022 a_n2318_8322.n9 a_n2318_8322.n8 0.358259
R24023 a_n2318_8322.n6 a_n2318_8322.n5 0.358259
R24024 a_n2318_8322.n5 a_n2318_8322.n3 0.358259
R24025 a_n2318_8322.n3 a_n2318_8322.n1 0.358259
R24026 a_n2318_8322.n18 a_n2318_8322.n16 0.358259
R24027 a_n2318_8322.n21 a_n2318_8322.n18 0.358259
R24028 a_n2318_8322.n21 a_n2318_8322.n20 0.358259
R24029 a_n2318_8322.n10 a_n2318_8322.n9 0.101793
R24030 a_n2318_8322.t27 a_n2318_8322.t26 0.0788333
R24031 a_n2318_8322.t25 a_n2318_8322.t27 0.0631667
R24032 a_n2318_8322.t24 a_n2318_8322.t25 0.0471944
R24033 a_n2318_8322.t24 a_n2318_8322.t26 0.0453889
C0 minus diffpairibias 3.4e-19
C1 commonsourceibias output 0.006808f
C2 vdd plus 0.085467f
C3 CSoutput minus 3.2739f
C4 plus diffpairibias 3.42e-19
C5 commonsourceibias outputibias 0.003832f
C6 vdd commonsourceibias 0.004218f
C7 CSoutput plus 0.896085f
C8 commonsourceibias diffpairibias 0.052527f
C9 CSoutput commonsourceibias 45.462303f
C10 minus plus 9.93573f
C11 minus commonsourceibias 0.332601f
C12 plus commonsourceibias 0.278362f
C13 output outputibias 2.34152f
C14 vdd output 7.23429f
C15 CSoutput output 6.13571f
C16 CSoutput outputibias 0.032386f
C17 vdd CSoutput 0.116614p
C18 diffpairibias gnd 59.99123f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.182005p
C22 plus gnd 35.1617f
C23 minus gnd 29.882719f
C24 CSoutput gnd 0.115669p
C25 vdd gnd 0.443441p
C26 a_n2318_8322.t26 gnd 39.5788f
C27 a_n2318_8322.t24 gnd 29.8018f
C28 a_n2318_8322.t27 gnd 19.7198f
C29 a_n2318_8322.t25 gnd 39.5788f
C30 a_n2318_8322.t12 gnd 0.095725f
C31 a_n2318_8322.t22 gnd 0.89632f
C32 a_n2318_8322.t10 gnd 0.095725f
C33 a_n2318_8322.t9 gnd 0.095725f
C34 a_n2318_8322.n0 gnd 0.674286f
C35 a_n2318_8322.n1 gnd 0.753416f
C36 a_n2318_8322.t19 gnd 0.095725f
C37 a_n2318_8322.t14 gnd 0.095725f
C38 a_n2318_8322.n2 gnd 0.674286f
C39 a_n2318_8322.n3 gnd 0.382801f
C40 a_n2318_8322.t17 gnd 0.095725f
C41 a_n2318_8322.t16 gnd 0.095725f
C42 a_n2318_8322.n4 gnd 0.674286f
C43 a_n2318_8322.n5 gnd 0.382801f
C44 a_n2318_8322.t8 gnd 0.894535f
C45 a_n2318_8322.n6 gnd 1.55036f
C46 a_n2318_8322.t3 gnd 0.89632f
C47 a_n2318_8322.t7 gnd 0.095725f
C48 a_n2318_8322.t6 gnd 0.095725f
C49 a_n2318_8322.n7 gnd 0.674286f
C50 a_n2318_8322.n8 gnd 0.753416f
C51 a_n2318_8322.t1 gnd 0.894535f
C52 a_n2318_8322.n9 gnd 0.379129f
C53 a_n2318_8322.t4 gnd 0.894535f
C54 a_n2318_8322.n10 gnd 0.379129f
C55 a_n2318_8322.t2 gnd 0.095725f
C56 a_n2318_8322.t0 gnd 0.095725f
C57 a_n2318_8322.n11 gnd 0.674286f
C58 a_n2318_8322.n12 gnd 0.382801f
C59 a_n2318_8322.t5 gnd 0.894535f
C60 a_n2318_8322.n13 gnd 1.07361f
C61 a_n2318_8322.n14 gnd 1.82505f
C62 a_n2318_8322.n15 gnd 3.97113f
C63 a_n2318_8322.t11 gnd 0.894535f
C64 a_n2318_8322.n16 gnd 0.880601f
C65 a_n2318_8322.t20 gnd 0.095725f
C66 a_n2318_8322.t13 gnd 0.095725f
C67 a_n2318_8322.n17 gnd 0.674286f
C68 a_n2318_8322.n18 gnd 0.382801f
C69 a_n2318_8322.t21 gnd 0.896317f
C70 a_n2318_8322.t18 gnd 0.095725f
C71 a_n2318_8322.t15 gnd 0.095725f
C72 a_n2318_8322.n19 gnd 0.674286f
C73 a_n2318_8322.n20 gnd 0.753418f
C74 a_n2318_8322.n21 gnd 0.382799f
C75 a_n2318_8322.n22 gnd 0.674288f
C76 a_n2318_8322.t23 gnd 0.095725f
C77 output.t13 gnd 0.464308f
C78 output.t19 gnd 0.044422f
C79 output.t8 gnd 0.044422f
C80 output.n0 gnd 0.364624f
C81 output.n1 gnd 0.614102f
C82 output.t12 gnd 0.044422f
C83 output.t4 gnd 0.044422f
C84 output.n2 gnd 0.364624f
C85 output.n3 gnd 0.350265f
C86 output.t6 gnd 0.044422f
C87 output.t5 gnd 0.044422f
C88 output.n4 gnd 0.364624f
C89 output.n5 gnd 0.350265f
C90 output.t11 gnd 0.044422f
C91 output.t14 gnd 0.044422f
C92 output.n6 gnd 0.364624f
C93 output.n7 gnd 0.350265f
C94 output.t16 gnd 0.044422f
C95 output.t9 gnd 0.044422f
C96 output.n8 gnd 0.364624f
C97 output.n9 gnd 0.350265f
C98 output.t10 gnd 0.044422f
C99 output.t17 gnd 0.044422f
C100 output.n10 gnd 0.364624f
C101 output.n11 gnd 0.350265f
C102 output.t18 gnd 0.044422f
C103 output.t7 gnd 0.044422f
C104 output.n12 gnd 0.364624f
C105 output.n13 gnd 0.350265f
C106 output.t15 gnd 0.462979f
C107 output.n14 gnd 0.28994f
C108 output.n15 gnd 0.015803f
C109 output.n16 gnd 0.011243f
C110 output.n17 gnd 0.006041f
C111 output.n18 gnd 0.01428f
C112 output.n19 gnd 0.006397f
C113 output.n20 gnd 0.011243f
C114 output.n21 gnd 0.006041f
C115 output.n22 gnd 0.01428f
C116 output.n23 gnd 0.006397f
C117 output.n24 gnd 0.048111f
C118 output.t3 gnd 0.023274f
C119 output.n25 gnd 0.01071f
C120 output.n26 gnd 0.008435f
C121 output.n27 gnd 0.006041f
C122 output.n28 gnd 0.267512f
C123 output.n29 gnd 0.011243f
C124 output.n30 gnd 0.006041f
C125 output.n31 gnd 0.006397f
C126 output.n32 gnd 0.01428f
C127 output.n33 gnd 0.01428f
C128 output.n34 gnd 0.006397f
C129 output.n35 gnd 0.006041f
C130 output.n36 gnd 0.011243f
C131 output.n37 gnd 0.011243f
C132 output.n38 gnd 0.006041f
C133 output.n39 gnd 0.006397f
C134 output.n40 gnd 0.01428f
C135 output.n41 gnd 0.030913f
C136 output.n42 gnd 0.006397f
C137 output.n43 gnd 0.006041f
C138 output.n44 gnd 0.025987f
C139 output.n45 gnd 0.097665f
C140 output.n46 gnd 0.015803f
C141 output.n47 gnd 0.011243f
C142 output.n48 gnd 0.006041f
C143 output.n49 gnd 0.01428f
C144 output.n50 gnd 0.006397f
C145 output.n51 gnd 0.011243f
C146 output.n52 gnd 0.006041f
C147 output.n53 gnd 0.01428f
C148 output.n54 gnd 0.006397f
C149 output.n55 gnd 0.048111f
C150 output.t1 gnd 0.023274f
C151 output.n56 gnd 0.01071f
C152 output.n57 gnd 0.008435f
C153 output.n58 gnd 0.006041f
C154 output.n59 gnd 0.267512f
C155 output.n60 gnd 0.011243f
C156 output.n61 gnd 0.006041f
C157 output.n62 gnd 0.006397f
C158 output.n63 gnd 0.01428f
C159 output.n64 gnd 0.01428f
C160 output.n65 gnd 0.006397f
C161 output.n66 gnd 0.006041f
C162 output.n67 gnd 0.011243f
C163 output.n68 gnd 0.011243f
C164 output.n69 gnd 0.006041f
C165 output.n70 gnd 0.006397f
C166 output.n71 gnd 0.01428f
C167 output.n72 gnd 0.030913f
C168 output.n73 gnd 0.006397f
C169 output.n74 gnd 0.006041f
C170 output.n75 gnd 0.025987f
C171 output.n76 gnd 0.09306f
C172 output.n77 gnd 1.65264f
C173 output.n78 gnd 0.015803f
C174 output.n79 gnd 0.011243f
C175 output.n80 gnd 0.006041f
C176 output.n81 gnd 0.01428f
C177 output.n82 gnd 0.006397f
C178 output.n83 gnd 0.011243f
C179 output.n84 gnd 0.006041f
C180 output.n85 gnd 0.01428f
C181 output.n86 gnd 0.006397f
C182 output.n87 gnd 0.048111f
C183 output.t2 gnd 0.023274f
C184 output.n88 gnd 0.01071f
C185 output.n89 gnd 0.008435f
C186 output.n90 gnd 0.006041f
C187 output.n91 gnd 0.267512f
C188 output.n92 gnd 0.011243f
C189 output.n93 gnd 0.006041f
C190 output.n94 gnd 0.006397f
C191 output.n95 gnd 0.01428f
C192 output.n96 gnd 0.01428f
C193 output.n97 gnd 0.006397f
C194 output.n98 gnd 0.006041f
C195 output.n99 gnd 0.011243f
C196 output.n100 gnd 0.011243f
C197 output.n101 gnd 0.006041f
C198 output.n102 gnd 0.006397f
C199 output.n103 gnd 0.01428f
C200 output.n104 gnd 0.030913f
C201 output.n105 gnd 0.006397f
C202 output.n106 gnd 0.006041f
C203 output.n107 gnd 0.025987f
C204 output.n108 gnd 0.09306f
C205 output.n109 gnd 0.713089f
C206 output.n110 gnd 0.015803f
C207 output.n111 gnd 0.011243f
C208 output.n112 gnd 0.006041f
C209 output.n113 gnd 0.01428f
C210 output.n114 gnd 0.006397f
C211 output.n115 gnd 0.011243f
C212 output.n116 gnd 0.006041f
C213 output.n117 gnd 0.01428f
C214 output.n118 gnd 0.006397f
C215 output.n119 gnd 0.048111f
C216 output.t0 gnd 0.023274f
C217 output.n120 gnd 0.01071f
C218 output.n121 gnd 0.008435f
C219 output.n122 gnd 0.006041f
C220 output.n123 gnd 0.267512f
C221 output.n124 gnd 0.011243f
C222 output.n125 gnd 0.006041f
C223 output.n126 gnd 0.006397f
C224 output.n127 gnd 0.01428f
C225 output.n128 gnd 0.01428f
C226 output.n129 gnd 0.006397f
C227 output.n130 gnd 0.006041f
C228 output.n131 gnd 0.011243f
C229 output.n132 gnd 0.011243f
C230 output.n133 gnd 0.006041f
C231 output.n134 gnd 0.006397f
C232 output.n135 gnd 0.01428f
C233 output.n136 gnd 0.030913f
C234 output.n137 gnd 0.006397f
C235 output.n138 gnd 0.006041f
C236 output.n139 gnd 0.025987f
C237 output.n140 gnd 0.09306f
C238 output.n141 gnd 1.67353f
C239 minus.n0 gnd 0.030538f
C240 minus.n1 gnd 0.00693f
C241 minus.n2 gnd 0.030538f
C242 minus.n3 gnd 0.00693f
C243 minus.n4 gnd 0.030538f
C244 minus.n5 gnd 0.00693f
C245 minus.n6 gnd 0.030538f
C246 minus.n7 gnd 0.00693f
C247 minus.t8 gnd 0.447069f
C248 minus.t7 gnd 0.431937f
C249 minus.n8 gnd 0.196988f
C250 minus.n9 gnd 0.17894f
C251 minus.n10 gnd 0.13035f
C252 minus.n11 gnd 0.030538f
C253 minus.t11 gnd 0.431937f
C254 minus.n12 gnd 0.19188f
C255 minus.n13 gnd 0.00693f
C256 minus.t10 gnd 0.431937f
C257 minus.n14 gnd 0.19188f
C258 minus.n15 gnd 0.030538f
C259 minus.n16 gnd 0.030538f
C260 minus.n17 gnd 0.030538f
C261 minus.t12 gnd 0.431937f
C262 minus.n18 gnd 0.19188f
C263 minus.n19 gnd 0.00693f
C264 minus.t17 gnd 0.431937f
C265 minus.n20 gnd 0.19188f
C266 minus.n21 gnd 0.030538f
C267 minus.n22 gnd 0.030538f
C268 minus.n23 gnd 0.030538f
C269 minus.t16 gnd 0.431937f
C270 minus.n24 gnd 0.19188f
C271 minus.n25 gnd 0.00693f
C272 minus.t21 gnd 0.431937f
C273 minus.n26 gnd 0.19188f
C274 minus.n27 gnd 0.030538f
C275 minus.n28 gnd 0.030538f
C276 minus.n29 gnd 0.030538f
C277 minus.t20 gnd 0.431937f
C278 minus.n30 gnd 0.19188f
C279 minus.n31 gnd 0.00693f
C280 minus.t13 gnd 0.431937f
C281 minus.n32 gnd 0.191598f
C282 minus.n33 gnd 0.352847f
C283 minus.n34 gnd 0.030538f
C284 minus.t5 gnd 0.431937f
C285 minus.t6 gnd 0.431937f
C286 minus.n35 gnd 0.030538f
C287 minus.t22 gnd 0.431937f
C288 minus.n36 gnd 0.19188f
C289 minus.n37 gnd 0.030538f
C290 minus.t18 gnd 0.431937f
C291 minus.t19 gnd 0.431937f
C292 minus.n38 gnd 0.19188f
C293 minus.n39 gnd 0.030538f
C294 minus.t14 gnd 0.431937f
C295 minus.t15 gnd 0.431937f
C296 minus.n40 gnd 0.19188f
C297 minus.n41 gnd 0.030538f
C298 minus.t9 gnd 0.431937f
C299 minus.t23 gnd 0.431937f
C300 minus.n42 gnd 0.196988f
C301 minus.t24 gnd 0.447069f
C302 minus.n43 gnd 0.17894f
C303 minus.n44 gnd 0.13035f
C304 minus.n45 gnd 0.00693f
C305 minus.n46 gnd 0.19188f
C306 minus.n47 gnd 0.00693f
C307 minus.n48 gnd 0.030538f
C308 minus.n49 gnd 0.030538f
C309 minus.n50 gnd 0.030538f
C310 minus.n51 gnd 0.00693f
C311 minus.n52 gnd 0.19188f
C312 minus.n53 gnd 0.00693f
C313 minus.n54 gnd 0.030538f
C314 minus.n55 gnd 0.030538f
C315 minus.n56 gnd 0.030538f
C316 minus.n57 gnd 0.00693f
C317 minus.n58 gnd 0.19188f
C318 minus.n59 gnd 0.00693f
C319 minus.n60 gnd 0.030538f
C320 minus.n61 gnd 0.030538f
C321 minus.n62 gnd 0.030538f
C322 minus.n63 gnd 0.00693f
C323 minus.n64 gnd 0.19188f
C324 minus.n65 gnd 0.00693f
C325 minus.n66 gnd 0.191598f
C326 minus.n67 gnd 0.954237f
C327 minus.n68 gnd 1.43659f
C328 minus.t2 gnd 0.009414f
C329 minus.t0 gnd 0.009414f
C330 minus.n69 gnd 0.030956f
C331 minus.t3 gnd 0.009414f
C332 minus.t1 gnd 0.009414f
C333 minus.n70 gnd 0.030532f
C334 minus.n71 gnd 0.260573f
C335 minus.t4 gnd 0.052398f
C336 minus.n72 gnd 0.142192f
C337 minus.n73 gnd 2.36188f
C338 commonsourceibias.n0 gnd 0.010724f
C339 commonsourceibias.t115 gnd 0.162395f
C340 commonsourceibias.t136 gnd 0.150157f
C341 commonsourceibias.n1 gnd 0.007823f
C342 commonsourceibias.n2 gnd 0.008037f
C343 commonsourceibias.t151 gnd 0.150157f
C344 commonsourceibias.n3 gnd 0.01034f
C345 commonsourceibias.n4 gnd 0.008037f
C346 commonsourceibias.t105 gnd 0.150157f
C347 commonsourceibias.n5 gnd 0.059912f
C348 commonsourceibias.t126 gnd 0.150157f
C349 commonsourceibias.n6 gnd 0.007578f
C350 commonsourceibias.n7 gnd 0.008037f
C351 commonsourceibias.t144 gnd 0.150157f
C352 commonsourceibias.n8 gnd 0.010186f
C353 commonsourceibias.n9 gnd 0.008037f
C354 commonsourceibias.t98 gnd 0.150157f
C355 commonsourceibias.n10 gnd 0.059912f
C356 commonsourceibias.t94 gnd 0.150157f
C357 commonsourceibias.n11 gnd 0.007361f
C358 commonsourceibias.n12 gnd 0.008037f
C359 commonsourceibias.t135 gnd 0.150157f
C360 commonsourceibias.n13 gnd 0.010015f
C361 commonsourceibias.n14 gnd 0.010724f
C362 commonsourceibias.t74 gnd 0.162395f
C363 commonsourceibias.t20 gnd 0.150157f
C364 commonsourceibias.n15 gnd 0.007823f
C365 commonsourceibias.n16 gnd 0.008037f
C366 commonsourceibias.t50 gnd 0.150157f
C367 commonsourceibias.n17 gnd 0.01034f
C368 commonsourceibias.n18 gnd 0.008037f
C369 commonsourceibias.t8 gnd 0.150157f
C370 commonsourceibias.n19 gnd 0.059912f
C371 commonsourceibias.t36 gnd 0.150157f
C372 commonsourceibias.n20 gnd 0.007578f
C373 commonsourceibias.n21 gnd 0.008037f
C374 commonsourceibias.t76 gnd 0.150157f
C375 commonsourceibias.n22 gnd 0.010186f
C376 commonsourceibias.n23 gnd 0.008037f
C377 commonsourceibias.t24 gnd 0.150157f
C378 commonsourceibias.n24 gnd 0.059912f
C379 commonsourceibias.t34 gnd 0.150157f
C380 commonsourceibias.n25 gnd 0.007361f
C381 commonsourceibias.n26 gnd 0.008037f
C382 commonsourceibias.t10 gnd 0.150157f
C383 commonsourceibias.n27 gnd 0.010015f
C384 commonsourceibias.n28 gnd 0.008037f
C385 commonsourceibias.t40 gnd 0.150157f
C386 commonsourceibias.n29 gnd 0.059912f
C387 commonsourceibias.t56 gnd 0.150157f
C388 commonsourceibias.n30 gnd 0.007172f
C389 commonsourceibias.n31 gnd 0.008037f
C390 commonsourceibias.t26 gnd 0.150157f
C391 commonsourceibias.n32 gnd 0.009825f
C392 commonsourceibias.n33 gnd 0.008037f
C393 commonsourceibias.t38 gnd 0.150157f
C394 commonsourceibias.n34 gnd 0.059912f
C395 commonsourceibias.t70 gnd 0.150157f
C396 commonsourceibias.n35 gnd 0.007008f
C397 commonsourceibias.n36 gnd 0.008037f
C398 commonsourceibias.t18 gnd 0.150157f
C399 commonsourceibias.n37 gnd 0.009613f
C400 commonsourceibias.n38 gnd 0.008037f
C401 commonsourceibias.t22 gnd 0.150157f
C402 commonsourceibias.n39 gnd 0.059912f
C403 commonsourceibias.t54 gnd 0.150157f
C404 commonsourceibias.n40 gnd 0.006868f
C405 commonsourceibias.n41 gnd 0.008037f
C406 commonsourceibias.t4 gnd 0.150157f
C407 commonsourceibias.n42 gnd 0.009378f
C408 commonsourceibias.t78 gnd 0.166947f
C409 commonsourceibias.t46 gnd 0.150157f
C410 commonsourceibias.n43 gnd 0.065449f
C411 commonsourceibias.n44 gnd 0.071822f
C412 commonsourceibias.n45 gnd 0.033327f
C413 commonsourceibias.n46 gnd 0.008037f
C414 commonsourceibias.n47 gnd 0.007823f
C415 commonsourceibias.n48 gnd 0.01121f
C416 commonsourceibias.n49 gnd 0.059912f
C417 commonsourceibias.n50 gnd 0.011203f
C418 commonsourceibias.n51 gnd 0.008037f
C419 commonsourceibias.n52 gnd 0.008037f
C420 commonsourceibias.n53 gnd 0.008037f
C421 commonsourceibias.n54 gnd 0.01034f
C422 commonsourceibias.n55 gnd 0.059912f
C423 commonsourceibias.n56 gnd 0.010583f
C424 commonsourceibias.n57 gnd 0.010282f
C425 commonsourceibias.n58 gnd 0.008037f
C426 commonsourceibias.n59 gnd 0.008037f
C427 commonsourceibias.n60 gnd 0.008037f
C428 commonsourceibias.n61 gnd 0.007578f
C429 commonsourceibias.n62 gnd 0.01122f
C430 commonsourceibias.n63 gnd 0.059912f
C431 commonsourceibias.n64 gnd 0.011217f
C432 commonsourceibias.n65 gnd 0.008037f
C433 commonsourceibias.n66 gnd 0.008037f
C434 commonsourceibias.n67 gnd 0.008037f
C435 commonsourceibias.n68 gnd 0.010186f
C436 commonsourceibias.n69 gnd 0.059912f
C437 commonsourceibias.n70 gnd 0.010507f
C438 commonsourceibias.n71 gnd 0.010357f
C439 commonsourceibias.n72 gnd 0.008037f
C440 commonsourceibias.n73 gnd 0.008037f
C441 commonsourceibias.n74 gnd 0.008037f
C442 commonsourceibias.n75 gnd 0.007361f
C443 commonsourceibias.n76 gnd 0.011225f
C444 commonsourceibias.n77 gnd 0.059912f
C445 commonsourceibias.n78 gnd 0.011224f
C446 commonsourceibias.n79 gnd 0.008037f
C447 commonsourceibias.n80 gnd 0.008037f
C448 commonsourceibias.n81 gnd 0.008037f
C449 commonsourceibias.n82 gnd 0.010015f
C450 commonsourceibias.n83 gnd 0.059912f
C451 commonsourceibias.n84 gnd 0.010432f
C452 commonsourceibias.n85 gnd 0.010432f
C453 commonsourceibias.n86 gnd 0.008037f
C454 commonsourceibias.n87 gnd 0.008037f
C455 commonsourceibias.n88 gnd 0.008037f
C456 commonsourceibias.n89 gnd 0.007172f
C457 commonsourceibias.n90 gnd 0.011224f
C458 commonsourceibias.n91 gnd 0.059912f
C459 commonsourceibias.n92 gnd 0.011225f
C460 commonsourceibias.n93 gnd 0.008037f
C461 commonsourceibias.n94 gnd 0.008037f
C462 commonsourceibias.n95 gnd 0.008037f
C463 commonsourceibias.n96 gnd 0.009825f
C464 commonsourceibias.n97 gnd 0.059912f
C465 commonsourceibias.n98 gnd 0.010357f
C466 commonsourceibias.n99 gnd 0.010507f
C467 commonsourceibias.n100 gnd 0.008037f
C468 commonsourceibias.n101 gnd 0.008037f
C469 commonsourceibias.n102 gnd 0.008037f
C470 commonsourceibias.n103 gnd 0.007008f
C471 commonsourceibias.n104 gnd 0.011217f
C472 commonsourceibias.n105 gnd 0.059912f
C473 commonsourceibias.n106 gnd 0.01122f
C474 commonsourceibias.n107 gnd 0.008037f
C475 commonsourceibias.n108 gnd 0.008037f
C476 commonsourceibias.n109 gnd 0.008037f
C477 commonsourceibias.n110 gnd 0.009613f
C478 commonsourceibias.n111 gnd 0.059912f
C479 commonsourceibias.n112 gnd 0.010282f
C480 commonsourceibias.n113 gnd 0.010583f
C481 commonsourceibias.n114 gnd 0.008037f
C482 commonsourceibias.n115 gnd 0.008037f
C483 commonsourceibias.n116 gnd 0.008037f
C484 commonsourceibias.n117 gnd 0.006868f
C485 commonsourceibias.n118 gnd 0.011203f
C486 commonsourceibias.n119 gnd 0.059912f
C487 commonsourceibias.n120 gnd 0.01121f
C488 commonsourceibias.n121 gnd 0.008037f
C489 commonsourceibias.n122 gnd 0.008037f
C490 commonsourceibias.n123 gnd 0.008037f
C491 commonsourceibias.n124 gnd 0.009378f
C492 commonsourceibias.n125 gnd 0.059912f
C493 commonsourceibias.n126 gnd 0.009861f
C494 commonsourceibias.n127 gnd 0.07189f
C495 commonsourceibias.n128 gnd 0.080075f
C496 commonsourceibias.t75 gnd 0.017343f
C497 commonsourceibias.t21 gnd 0.017343f
C498 commonsourceibias.n129 gnd 0.15325f
C499 commonsourceibias.n130 gnd 0.132562f
C500 commonsourceibias.t51 gnd 0.017343f
C501 commonsourceibias.t9 gnd 0.017343f
C502 commonsourceibias.n131 gnd 0.15325f
C503 commonsourceibias.n132 gnd 0.070394f
C504 commonsourceibias.t37 gnd 0.017343f
C505 commonsourceibias.t77 gnd 0.017343f
C506 commonsourceibias.n133 gnd 0.15325f
C507 commonsourceibias.n134 gnd 0.070394f
C508 commonsourceibias.t25 gnd 0.017343f
C509 commonsourceibias.t35 gnd 0.017343f
C510 commonsourceibias.n135 gnd 0.15325f
C511 commonsourceibias.n136 gnd 0.070394f
C512 commonsourceibias.t11 gnd 0.017343f
C513 commonsourceibias.t41 gnd 0.017343f
C514 commonsourceibias.n137 gnd 0.15325f
C515 commonsourceibias.n138 gnd 0.058811f
C516 commonsourceibias.t47 gnd 0.017343f
C517 commonsourceibias.t79 gnd 0.017343f
C518 commonsourceibias.n139 gnd 0.153763f
C519 commonsourceibias.t55 gnd 0.017343f
C520 commonsourceibias.t5 gnd 0.017343f
C521 commonsourceibias.n140 gnd 0.15325f
C522 commonsourceibias.n141 gnd 0.1428f
C523 commonsourceibias.t19 gnd 0.017343f
C524 commonsourceibias.t23 gnd 0.017343f
C525 commonsourceibias.n142 gnd 0.15325f
C526 commonsourceibias.n143 gnd 0.070394f
C527 commonsourceibias.t39 gnd 0.017343f
C528 commonsourceibias.t71 gnd 0.017343f
C529 commonsourceibias.n144 gnd 0.15325f
C530 commonsourceibias.n145 gnd 0.070394f
C531 commonsourceibias.t57 gnd 0.017343f
C532 commonsourceibias.t27 gnd 0.017343f
C533 commonsourceibias.n146 gnd 0.15325f
C534 commonsourceibias.n147 gnd 0.058811f
C535 commonsourceibias.n148 gnd 0.071213f
C536 commonsourceibias.n149 gnd 0.052016f
C537 commonsourceibias.t153 gnd 0.150157f
C538 commonsourceibias.n150 gnd 0.059912f
C539 commonsourceibias.t88 gnd 0.150157f
C540 commonsourceibias.n151 gnd 0.059912f
C541 commonsourceibias.n152 gnd 0.008037f
C542 commonsourceibias.t125 gnd 0.150157f
C543 commonsourceibias.n153 gnd 0.059912f
C544 commonsourceibias.n154 gnd 0.008037f
C545 commonsourceibias.t120 gnd 0.150157f
C546 commonsourceibias.n155 gnd 0.059912f
C547 commonsourceibias.n156 gnd 0.008037f
C548 commonsourceibias.t139 gnd 0.150157f
C549 commonsourceibias.n157 gnd 0.007008f
C550 commonsourceibias.n158 gnd 0.008037f
C551 commonsourceibias.t112 gnd 0.150157f
C552 commonsourceibias.n159 gnd 0.009613f
C553 commonsourceibias.n160 gnd 0.008037f
C554 commonsourceibias.t107 gnd 0.150157f
C555 commonsourceibias.n161 gnd 0.059912f
C556 commonsourceibias.t127 gnd 0.150157f
C557 commonsourceibias.n162 gnd 0.006868f
C558 commonsourceibias.n163 gnd 0.008037f
C559 commonsourceibias.t146 gnd 0.150157f
C560 commonsourceibias.n164 gnd 0.009378f
C561 commonsourceibias.t117 gnd 0.166947f
C562 commonsourceibias.t99 gnd 0.150157f
C563 commonsourceibias.n165 gnd 0.065449f
C564 commonsourceibias.n166 gnd 0.071822f
C565 commonsourceibias.n167 gnd 0.033327f
C566 commonsourceibias.n168 gnd 0.008037f
C567 commonsourceibias.n169 gnd 0.007823f
C568 commonsourceibias.n170 gnd 0.01121f
C569 commonsourceibias.n171 gnd 0.059912f
C570 commonsourceibias.n172 gnd 0.011203f
C571 commonsourceibias.n173 gnd 0.008037f
C572 commonsourceibias.n174 gnd 0.008037f
C573 commonsourceibias.n175 gnd 0.008037f
C574 commonsourceibias.n176 gnd 0.01034f
C575 commonsourceibias.n177 gnd 0.059912f
C576 commonsourceibias.n178 gnd 0.010583f
C577 commonsourceibias.n179 gnd 0.010282f
C578 commonsourceibias.n180 gnd 0.008037f
C579 commonsourceibias.n181 gnd 0.008037f
C580 commonsourceibias.n182 gnd 0.008037f
C581 commonsourceibias.n183 gnd 0.007578f
C582 commonsourceibias.n184 gnd 0.01122f
C583 commonsourceibias.n185 gnd 0.059912f
C584 commonsourceibias.n186 gnd 0.011217f
C585 commonsourceibias.n187 gnd 0.008037f
C586 commonsourceibias.n188 gnd 0.008037f
C587 commonsourceibias.n189 gnd 0.008037f
C588 commonsourceibias.n190 gnd 0.010186f
C589 commonsourceibias.n191 gnd 0.059912f
C590 commonsourceibias.n192 gnd 0.010507f
C591 commonsourceibias.n193 gnd 0.010357f
C592 commonsourceibias.n194 gnd 0.008037f
C593 commonsourceibias.n195 gnd 0.008037f
C594 commonsourceibias.n196 gnd 0.009825f
C595 commonsourceibias.n197 gnd 0.007361f
C596 commonsourceibias.n198 gnd 0.011225f
C597 commonsourceibias.n199 gnd 0.008037f
C598 commonsourceibias.n200 gnd 0.008037f
C599 commonsourceibias.n201 gnd 0.011224f
C600 commonsourceibias.n202 gnd 0.007172f
C601 commonsourceibias.n203 gnd 0.010015f
C602 commonsourceibias.n204 gnd 0.008037f
C603 commonsourceibias.n205 gnd 0.007021f
C604 commonsourceibias.n206 gnd 0.010432f
C605 commonsourceibias.n207 gnd 0.010432f
C606 commonsourceibias.n208 gnd 0.007021f
C607 commonsourceibias.n209 gnd 0.008037f
C608 commonsourceibias.n210 gnd 0.008037f
C609 commonsourceibias.n211 gnd 0.007172f
C610 commonsourceibias.n212 gnd 0.011224f
C611 commonsourceibias.n213 gnd 0.059912f
C612 commonsourceibias.n214 gnd 0.011225f
C613 commonsourceibias.n215 gnd 0.008037f
C614 commonsourceibias.n216 gnd 0.008037f
C615 commonsourceibias.n217 gnd 0.008037f
C616 commonsourceibias.n218 gnd 0.009825f
C617 commonsourceibias.n219 gnd 0.059912f
C618 commonsourceibias.n220 gnd 0.010357f
C619 commonsourceibias.n221 gnd 0.010507f
C620 commonsourceibias.n222 gnd 0.008037f
C621 commonsourceibias.n223 gnd 0.008037f
C622 commonsourceibias.n224 gnd 0.008037f
C623 commonsourceibias.n225 gnd 0.007008f
C624 commonsourceibias.n226 gnd 0.011217f
C625 commonsourceibias.n227 gnd 0.059912f
C626 commonsourceibias.n228 gnd 0.01122f
C627 commonsourceibias.n229 gnd 0.008037f
C628 commonsourceibias.n230 gnd 0.008037f
C629 commonsourceibias.n231 gnd 0.008037f
C630 commonsourceibias.n232 gnd 0.009613f
C631 commonsourceibias.n233 gnd 0.059912f
C632 commonsourceibias.n234 gnd 0.010282f
C633 commonsourceibias.n235 gnd 0.010583f
C634 commonsourceibias.n236 gnd 0.008037f
C635 commonsourceibias.n237 gnd 0.008037f
C636 commonsourceibias.n238 gnd 0.008037f
C637 commonsourceibias.n239 gnd 0.006868f
C638 commonsourceibias.n240 gnd 0.011203f
C639 commonsourceibias.n241 gnd 0.059912f
C640 commonsourceibias.n242 gnd 0.01121f
C641 commonsourceibias.n243 gnd 0.008037f
C642 commonsourceibias.n244 gnd 0.008037f
C643 commonsourceibias.n245 gnd 0.008037f
C644 commonsourceibias.n246 gnd 0.009378f
C645 commonsourceibias.n247 gnd 0.059912f
C646 commonsourceibias.n248 gnd 0.009861f
C647 commonsourceibias.n249 gnd 0.07189f
C648 commonsourceibias.n250 gnd 0.04697f
C649 commonsourceibias.n251 gnd 0.010724f
C650 commonsourceibias.t119 gnd 0.150157f
C651 commonsourceibias.n252 gnd 0.007823f
C652 commonsourceibias.n253 gnd 0.008037f
C653 commonsourceibias.t137 gnd 0.150157f
C654 commonsourceibias.n254 gnd 0.01034f
C655 commonsourceibias.n255 gnd 0.008037f
C656 commonsourceibias.t92 gnd 0.150157f
C657 commonsourceibias.n256 gnd 0.059912f
C658 commonsourceibias.t109 gnd 0.150157f
C659 commonsourceibias.n257 gnd 0.007578f
C660 commonsourceibias.n258 gnd 0.008037f
C661 commonsourceibias.t128 gnd 0.150157f
C662 commonsourceibias.n259 gnd 0.010186f
C663 commonsourceibias.n260 gnd 0.008037f
C664 commonsourceibias.t86 gnd 0.150157f
C665 commonsourceibias.n261 gnd 0.059912f
C666 commonsourceibias.t83 gnd 0.150157f
C667 commonsourceibias.n262 gnd 0.007361f
C668 commonsourceibias.n263 gnd 0.008037f
C669 commonsourceibias.t118 gnd 0.150157f
C670 commonsourceibias.n264 gnd 0.010015f
C671 commonsourceibias.n265 gnd 0.008037f
C672 commonsourceibias.t138 gnd 0.150157f
C673 commonsourceibias.n266 gnd 0.059912f
C674 commonsourceibias.t159 gnd 0.150157f
C675 commonsourceibias.n267 gnd 0.007172f
C676 commonsourceibias.n268 gnd 0.008037f
C677 commonsourceibias.t108 gnd 0.150157f
C678 commonsourceibias.n269 gnd 0.009825f
C679 commonsourceibias.n270 gnd 0.008037f
C680 commonsourceibias.t102 gnd 0.150157f
C681 commonsourceibias.n271 gnd 0.059912f
C682 commonsourceibias.t121 gnd 0.150157f
C683 commonsourceibias.n272 gnd 0.007008f
C684 commonsourceibias.n273 gnd 0.008037f
C685 commonsourceibias.t95 gnd 0.150157f
C686 commonsourceibias.n274 gnd 0.009613f
C687 commonsourceibias.n275 gnd 0.008037f
C688 commonsourceibias.t93 gnd 0.150157f
C689 commonsourceibias.n276 gnd 0.059912f
C690 commonsourceibias.t110 gnd 0.150157f
C691 commonsourceibias.n277 gnd 0.006868f
C692 commonsourceibias.n278 gnd 0.008037f
C693 commonsourceibias.t129 gnd 0.150157f
C694 commonsourceibias.n279 gnd 0.009378f
C695 commonsourceibias.t101 gnd 0.166947f
C696 commonsourceibias.t87 gnd 0.150157f
C697 commonsourceibias.n280 gnd 0.065449f
C698 commonsourceibias.n281 gnd 0.071822f
C699 commonsourceibias.n282 gnd 0.033327f
C700 commonsourceibias.n283 gnd 0.008037f
C701 commonsourceibias.n284 gnd 0.007823f
C702 commonsourceibias.n285 gnd 0.01121f
C703 commonsourceibias.n286 gnd 0.059912f
C704 commonsourceibias.n287 gnd 0.011203f
C705 commonsourceibias.n288 gnd 0.008037f
C706 commonsourceibias.n289 gnd 0.008037f
C707 commonsourceibias.n290 gnd 0.008037f
C708 commonsourceibias.n291 gnd 0.01034f
C709 commonsourceibias.n292 gnd 0.059912f
C710 commonsourceibias.n293 gnd 0.010583f
C711 commonsourceibias.n294 gnd 0.010282f
C712 commonsourceibias.n295 gnd 0.008037f
C713 commonsourceibias.n296 gnd 0.008037f
C714 commonsourceibias.n297 gnd 0.008037f
C715 commonsourceibias.n298 gnd 0.007578f
C716 commonsourceibias.n299 gnd 0.01122f
C717 commonsourceibias.n300 gnd 0.059912f
C718 commonsourceibias.n301 gnd 0.011217f
C719 commonsourceibias.n302 gnd 0.008037f
C720 commonsourceibias.n303 gnd 0.008037f
C721 commonsourceibias.n304 gnd 0.008037f
C722 commonsourceibias.n305 gnd 0.010186f
C723 commonsourceibias.n306 gnd 0.059912f
C724 commonsourceibias.n307 gnd 0.010507f
C725 commonsourceibias.n308 gnd 0.010357f
C726 commonsourceibias.n309 gnd 0.008037f
C727 commonsourceibias.n310 gnd 0.008037f
C728 commonsourceibias.n311 gnd 0.008037f
C729 commonsourceibias.n312 gnd 0.007361f
C730 commonsourceibias.n313 gnd 0.011225f
C731 commonsourceibias.n314 gnd 0.059912f
C732 commonsourceibias.n315 gnd 0.011224f
C733 commonsourceibias.n316 gnd 0.008037f
C734 commonsourceibias.n317 gnd 0.008037f
C735 commonsourceibias.n318 gnd 0.008037f
C736 commonsourceibias.n319 gnd 0.010015f
C737 commonsourceibias.n320 gnd 0.059912f
C738 commonsourceibias.n321 gnd 0.010432f
C739 commonsourceibias.n322 gnd 0.010432f
C740 commonsourceibias.n323 gnd 0.008037f
C741 commonsourceibias.n324 gnd 0.008037f
C742 commonsourceibias.n325 gnd 0.008037f
C743 commonsourceibias.n326 gnd 0.007172f
C744 commonsourceibias.n327 gnd 0.011224f
C745 commonsourceibias.n328 gnd 0.059912f
C746 commonsourceibias.n329 gnd 0.011225f
C747 commonsourceibias.n330 gnd 0.008037f
C748 commonsourceibias.n331 gnd 0.008037f
C749 commonsourceibias.n332 gnd 0.008037f
C750 commonsourceibias.n333 gnd 0.009825f
C751 commonsourceibias.n334 gnd 0.059912f
C752 commonsourceibias.n335 gnd 0.010357f
C753 commonsourceibias.n336 gnd 0.010507f
C754 commonsourceibias.n337 gnd 0.008037f
C755 commonsourceibias.n338 gnd 0.008037f
C756 commonsourceibias.n339 gnd 0.008037f
C757 commonsourceibias.n340 gnd 0.007008f
C758 commonsourceibias.n341 gnd 0.011217f
C759 commonsourceibias.n342 gnd 0.059912f
C760 commonsourceibias.n343 gnd 0.01122f
C761 commonsourceibias.n344 gnd 0.008037f
C762 commonsourceibias.n345 gnd 0.008037f
C763 commonsourceibias.n346 gnd 0.008037f
C764 commonsourceibias.n347 gnd 0.009613f
C765 commonsourceibias.n348 gnd 0.059912f
C766 commonsourceibias.n349 gnd 0.010282f
C767 commonsourceibias.n350 gnd 0.010583f
C768 commonsourceibias.n351 gnd 0.008037f
C769 commonsourceibias.n352 gnd 0.008037f
C770 commonsourceibias.n353 gnd 0.008037f
C771 commonsourceibias.n354 gnd 0.006868f
C772 commonsourceibias.n355 gnd 0.011203f
C773 commonsourceibias.n356 gnd 0.059912f
C774 commonsourceibias.n357 gnd 0.01121f
C775 commonsourceibias.n358 gnd 0.008037f
C776 commonsourceibias.n359 gnd 0.008037f
C777 commonsourceibias.n360 gnd 0.008037f
C778 commonsourceibias.n361 gnd 0.009378f
C779 commonsourceibias.n362 gnd 0.059912f
C780 commonsourceibias.n363 gnd 0.009861f
C781 commonsourceibias.t100 gnd 0.162395f
C782 commonsourceibias.n364 gnd 0.07189f
C783 commonsourceibias.n365 gnd 0.025003f
C784 commonsourceibias.n366 gnd 0.464917f
C785 commonsourceibias.n367 gnd 0.010724f
C786 commonsourceibias.t140 gnd 0.162395f
C787 commonsourceibias.t155 gnd 0.150157f
C788 commonsourceibias.n368 gnd 0.007823f
C789 commonsourceibias.n369 gnd 0.008037f
C790 commonsourceibias.t84 gnd 0.150157f
C791 commonsourceibias.n370 gnd 0.01034f
C792 commonsourceibias.n371 gnd 0.008037f
C793 commonsourceibias.t148 gnd 0.150157f
C794 commonsourceibias.n372 gnd 0.007578f
C795 commonsourceibias.n373 gnd 0.008037f
C796 commonsourceibias.t80 gnd 0.150157f
C797 commonsourceibias.n374 gnd 0.010186f
C798 commonsourceibias.n375 gnd 0.008037f
C799 commonsourceibias.t113 gnd 0.150157f
C800 commonsourceibias.n376 gnd 0.007361f
C801 commonsourceibias.n377 gnd 0.008037f
C802 commonsourceibias.t154 gnd 0.150157f
C803 commonsourceibias.n378 gnd 0.010015f
C804 commonsourceibias.t29 gnd 0.017343f
C805 commonsourceibias.t3 gnd 0.017343f
C806 commonsourceibias.n379 gnd 0.153763f
C807 commonsourceibias.t49 gnd 0.017343f
C808 commonsourceibias.t13 gnd 0.017343f
C809 commonsourceibias.n380 gnd 0.15325f
C810 commonsourceibias.n381 gnd 0.1428f
C811 commonsourceibias.t69 gnd 0.017343f
C812 commonsourceibias.t67 gnd 0.017343f
C813 commonsourceibias.n382 gnd 0.15325f
C814 commonsourceibias.n383 gnd 0.070394f
C815 commonsourceibias.t7 gnd 0.017343f
C816 commonsourceibias.t63 gnd 0.017343f
C817 commonsourceibias.n384 gnd 0.15325f
C818 commonsourceibias.n385 gnd 0.070394f
C819 commonsourceibias.t53 gnd 0.017343f
C820 commonsourceibias.t73 gnd 0.017343f
C821 commonsourceibias.n386 gnd 0.15325f
C822 commonsourceibias.n387 gnd 0.058811f
C823 commonsourceibias.n388 gnd 0.010724f
C824 commonsourceibias.t42 gnd 0.150157f
C825 commonsourceibias.n389 gnd 0.007823f
C826 commonsourceibias.n390 gnd 0.008037f
C827 commonsourceibias.t0 gnd 0.150157f
C828 commonsourceibias.n391 gnd 0.01034f
C829 commonsourceibias.n392 gnd 0.008037f
C830 commonsourceibias.t60 gnd 0.150157f
C831 commonsourceibias.n393 gnd 0.007578f
C832 commonsourceibias.n394 gnd 0.008037f
C833 commonsourceibias.t16 gnd 0.150157f
C834 commonsourceibias.n395 gnd 0.010186f
C835 commonsourceibias.n396 gnd 0.008037f
C836 commonsourceibias.t58 gnd 0.150157f
C837 commonsourceibias.n397 gnd 0.007361f
C838 commonsourceibias.n398 gnd 0.008037f
C839 commonsourceibias.t32 gnd 0.150157f
C840 commonsourceibias.n399 gnd 0.010015f
C841 commonsourceibias.n400 gnd 0.008037f
C842 commonsourceibias.t72 gnd 0.150157f
C843 commonsourceibias.n401 gnd 0.007172f
C844 commonsourceibias.n402 gnd 0.008037f
C845 commonsourceibias.t52 gnd 0.150157f
C846 commonsourceibias.n403 gnd 0.009825f
C847 commonsourceibias.n404 gnd 0.008037f
C848 commonsourceibias.t6 gnd 0.150157f
C849 commonsourceibias.n405 gnd 0.007008f
C850 commonsourceibias.n406 gnd 0.008037f
C851 commonsourceibias.t66 gnd 0.150157f
C852 commonsourceibias.n407 gnd 0.009613f
C853 commonsourceibias.n408 gnd 0.008037f
C854 commonsourceibias.t12 gnd 0.150157f
C855 commonsourceibias.n409 gnd 0.006868f
C856 commonsourceibias.n410 gnd 0.008037f
C857 commonsourceibias.t48 gnd 0.150157f
C858 commonsourceibias.n411 gnd 0.009378f
C859 commonsourceibias.t28 gnd 0.166947f
C860 commonsourceibias.t2 gnd 0.150157f
C861 commonsourceibias.n412 gnd 0.065449f
C862 commonsourceibias.n413 gnd 0.071822f
C863 commonsourceibias.n414 gnd 0.033327f
C864 commonsourceibias.n415 gnd 0.008037f
C865 commonsourceibias.n416 gnd 0.007823f
C866 commonsourceibias.n417 gnd 0.01121f
C867 commonsourceibias.n418 gnd 0.059912f
C868 commonsourceibias.n419 gnd 0.011203f
C869 commonsourceibias.n420 gnd 0.008037f
C870 commonsourceibias.n421 gnd 0.008037f
C871 commonsourceibias.n422 gnd 0.008037f
C872 commonsourceibias.n423 gnd 0.01034f
C873 commonsourceibias.n424 gnd 0.059912f
C874 commonsourceibias.n425 gnd 0.010583f
C875 commonsourceibias.t68 gnd 0.150157f
C876 commonsourceibias.n426 gnd 0.059912f
C877 commonsourceibias.n427 gnd 0.010282f
C878 commonsourceibias.n428 gnd 0.008037f
C879 commonsourceibias.n429 gnd 0.008037f
C880 commonsourceibias.n430 gnd 0.008037f
C881 commonsourceibias.n431 gnd 0.007578f
C882 commonsourceibias.n432 gnd 0.01122f
C883 commonsourceibias.n433 gnd 0.059912f
C884 commonsourceibias.n434 gnd 0.011217f
C885 commonsourceibias.n435 gnd 0.008037f
C886 commonsourceibias.n436 gnd 0.008037f
C887 commonsourceibias.n437 gnd 0.008037f
C888 commonsourceibias.n438 gnd 0.010186f
C889 commonsourceibias.n439 gnd 0.059912f
C890 commonsourceibias.n440 gnd 0.010507f
C891 commonsourceibias.t62 gnd 0.150157f
C892 commonsourceibias.n441 gnd 0.059912f
C893 commonsourceibias.n442 gnd 0.010357f
C894 commonsourceibias.n443 gnd 0.008037f
C895 commonsourceibias.n444 gnd 0.008037f
C896 commonsourceibias.n445 gnd 0.008037f
C897 commonsourceibias.n446 gnd 0.007361f
C898 commonsourceibias.n447 gnd 0.011225f
C899 commonsourceibias.n448 gnd 0.059912f
C900 commonsourceibias.n449 gnd 0.011224f
C901 commonsourceibias.n450 gnd 0.008037f
C902 commonsourceibias.n451 gnd 0.008037f
C903 commonsourceibias.n452 gnd 0.008037f
C904 commonsourceibias.n453 gnd 0.010015f
C905 commonsourceibias.n454 gnd 0.059912f
C906 commonsourceibias.n455 gnd 0.010432f
C907 commonsourceibias.t64 gnd 0.150157f
C908 commonsourceibias.n456 gnd 0.059912f
C909 commonsourceibias.n457 gnd 0.010432f
C910 commonsourceibias.n458 gnd 0.008037f
C911 commonsourceibias.n459 gnd 0.008037f
C912 commonsourceibias.n460 gnd 0.008037f
C913 commonsourceibias.n461 gnd 0.007172f
C914 commonsourceibias.n462 gnd 0.011224f
C915 commonsourceibias.n463 gnd 0.059912f
C916 commonsourceibias.n464 gnd 0.011225f
C917 commonsourceibias.n465 gnd 0.008037f
C918 commonsourceibias.n466 gnd 0.008037f
C919 commonsourceibias.n467 gnd 0.008037f
C920 commonsourceibias.n468 gnd 0.009825f
C921 commonsourceibias.n469 gnd 0.059912f
C922 commonsourceibias.n470 gnd 0.010357f
C923 commonsourceibias.t44 gnd 0.150157f
C924 commonsourceibias.n471 gnd 0.059912f
C925 commonsourceibias.n472 gnd 0.010507f
C926 commonsourceibias.n473 gnd 0.008037f
C927 commonsourceibias.n474 gnd 0.008037f
C928 commonsourceibias.n475 gnd 0.008037f
C929 commonsourceibias.n476 gnd 0.007008f
C930 commonsourceibias.n477 gnd 0.011217f
C931 commonsourceibias.n478 gnd 0.059912f
C932 commonsourceibias.n479 gnd 0.01122f
C933 commonsourceibias.n480 gnd 0.008037f
C934 commonsourceibias.n481 gnd 0.008037f
C935 commonsourceibias.n482 gnd 0.008037f
C936 commonsourceibias.n483 gnd 0.009613f
C937 commonsourceibias.n484 gnd 0.059912f
C938 commonsourceibias.n485 gnd 0.010282f
C939 commonsourceibias.t30 gnd 0.150157f
C940 commonsourceibias.n486 gnd 0.059912f
C941 commonsourceibias.n487 gnd 0.010583f
C942 commonsourceibias.n488 gnd 0.008037f
C943 commonsourceibias.n489 gnd 0.008037f
C944 commonsourceibias.n490 gnd 0.008037f
C945 commonsourceibias.n491 gnd 0.006868f
C946 commonsourceibias.n492 gnd 0.011203f
C947 commonsourceibias.n493 gnd 0.059912f
C948 commonsourceibias.n494 gnd 0.01121f
C949 commonsourceibias.n495 gnd 0.008037f
C950 commonsourceibias.n496 gnd 0.008037f
C951 commonsourceibias.n497 gnd 0.008037f
C952 commonsourceibias.n498 gnd 0.009378f
C953 commonsourceibias.n499 gnd 0.059912f
C954 commonsourceibias.n500 gnd 0.009861f
C955 commonsourceibias.t14 gnd 0.162395f
C956 commonsourceibias.n501 gnd 0.07189f
C957 commonsourceibias.n502 gnd 0.080075f
C958 commonsourceibias.t43 gnd 0.017343f
C959 commonsourceibias.t15 gnd 0.017343f
C960 commonsourceibias.n503 gnd 0.15325f
C961 commonsourceibias.n504 gnd 0.132562f
C962 commonsourceibias.t31 gnd 0.017343f
C963 commonsourceibias.t1 gnd 0.017343f
C964 commonsourceibias.n505 gnd 0.15325f
C965 commonsourceibias.n506 gnd 0.070394f
C966 commonsourceibias.t17 gnd 0.017343f
C967 commonsourceibias.t61 gnd 0.017343f
C968 commonsourceibias.n507 gnd 0.15325f
C969 commonsourceibias.n508 gnd 0.070394f
C970 commonsourceibias.t59 gnd 0.017343f
C971 commonsourceibias.t45 gnd 0.017343f
C972 commonsourceibias.n509 gnd 0.15325f
C973 commonsourceibias.n510 gnd 0.070394f
C974 commonsourceibias.t65 gnd 0.017343f
C975 commonsourceibias.t33 gnd 0.017343f
C976 commonsourceibias.n511 gnd 0.15325f
C977 commonsourceibias.n512 gnd 0.058811f
C978 commonsourceibias.n513 gnd 0.071213f
C979 commonsourceibias.n514 gnd 0.052016f
C980 commonsourceibias.t82 gnd 0.150157f
C981 commonsourceibias.n515 gnd 0.059912f
C982 commonsourceibias.n516 gnd 0.008037f
C983 commonsourceibias.t147 gnd 0.150157f
C984 commonsourceibias.n517 gnd 0.059912f
C985 commonsourceibias.n518 gnd 0.008037f
C986 commonsourceibias.t143 gnd 0.150157f
C987 commonsourceibias.n519 gnd 0.059912f
C988 commonsourceibias.n520 gnd 0.008037f
C989 commonsourceibias.t158 gnd 0.150157f
C990 commonsourceibias.n521 gnd 0.007008f
C991 commonsourceibias.n522 gnd 0.008037f
C992 commonsourceibias.t104 gnd 0.150157f
C993 commonsourceibias.n523 gnd 0.009613f
C994 commonsourceibias.n524 gnd 0.008037f
C995 commonsourceibias.t133 gnd 0.150157f
C996 commonsourceibias.n525 gnd 0.006868f
C997 commonsourceibias.n526 gnd 0.008037f
C998 commonsourceibias.t150 gnd 0.150157f
C999 commonsourceibias.n527 gnd 0.009378f
C1000 commonsourceibias.t123 gnd 0.166947f
C1001 commonsourceibias.t103 gnd 0.150157f
C1002 commonsourceibias.n528 gnd 0.065449f
C1003 commonsourceibias.n529 gnd 0.071822f
C1004 commonsourceibias.n530 gnd 0.033327f
C1005 commonsourceibias.n531 gnd 0.008037f
C1006 commonsourceibias.n532 gnd 0.007823f
C1007 commonsourceibias.n533 gnd 0.01121f
C1008 commonsourceibias.n534 gnd 0.059912f
C1009 commonsourceibias.n535 gnd 0.011203f
C1010 commonsourceibias.n536 gnd 0.008037f
C1011 commonsourceibias.n537 gnd 0.008037f
C1012 commonsourceibias.n538 gnd 0.008037f
C1013 commonsourceibias.n539 gnd 0.01034f
C1014 commonsourceibias.n540 gnd 0.059912f
C1015 commonsourceibias.n541 gnd 0.010583f
C1016 commonsourceibias.t114 gnd 0.150157f
C1017 commonsourceibias.n542 gnd 0.059912f
C1018 commonsourceibias.n543 gnd 0.010282f
C1019 commonsourceibias.n544 gnd 0.008037f
C1020 commonsourceibias.n545 gnd 0.008037f
C1021 commonsourceibias.n546 gnd 0.008037f
C1022 commonsourceibias.n547 gnd 0.007578f
C1023 commonsourceibias.n548 gnd 0.01122f
C1024 commonsourceibias.n549 gnd 0.059912f
C1025 commonsourceibias.n550 gnd 0.011217f
C1026 commonsourceibias.n551 gnd 0.008037f
C1027 commonsourceibias.n552 gnd 0.008037f
C1028 commonsourceibias.n553 gnd 0.008037f
C1029 commonsourceibias.n554 gnd 0.010186f
C1030 commonsourceibias.n555 gnd 0.059912f
C1031 commonsourceibias.n556 gnd 0.010507f
C1032 commonsourceibias.n557 gnd 0.010357f
C1033 commonsourceibias.n558 gnd 0.008037f
C1034 commonsourceibias.n559 gnd 0.008037f
C1035 commonsourceibias.n560 gnd 0.009825f
C1036 commonsourceibias.n561 gnd 0.007361f
C1037 commonsourceibias.n562 gnd 0.011225f
C1038 commonsourceibias.n563 gnd 0.008037f
C1039 commonsourceibias.n564 gnd 0.008037f
C1040 commonsourceibias.n565 gnd 0.011224f
C1041 commonsourceibias.n566 gnd 0.007172f
C1042 commonsourceibias.n567 gnd 0.010015f
C1043 commonsourceibias.n568 gnd 0.008037f
C1044 commonsourceibias.n569 gnd 0.007021f
C1045 commonsourceibias.n570 gnd 0.010432f
C1046 commonsourceibias.t85 gnd 0.150157f
C1047 commonsourceibias.n571 gnd 0.059912f
C1048 commonsourceibias.n572 gnd 0.010432f
C1049 commonsourceibias.n573 gnd 0.007021f
C1050 commonsourceibias.n574 gnd 0.008037f
C1051 commonsourceibias.n575 gnd 0.008037f
C1052 commonsourceibias.n576 gnd 0.007172f
C1053 commonsourceibias.n577 gnd 0.011224f
C1054 commonsourceibias.n578 gnd 0.059912f
C1055 commonsourceibias.n579 gnd 0.011225f
C1056 commonsourceibias.n580 gnd 0.008037f
C1057 commonsourceibias.n581 gnd 0.008037f
C1058 commonsourceibias.n582 gnd 0.008037f
C1059 commonsourceibias.n583 gnd 0.009825f
C1060 commonsourceibias.n584 gnd 0.059912f
C1061 commonsourceibias.n585 gnd 0.010357f
C1062 commonsourceibias.t89 gnd 0.150157f
C1063 commonsourceibias.n586 gnd 0.059912f
C1064 commonsourceibias.n587 gnd 0.010507f
C1065 commonsourceibias.n588 gnd 0.008037f
C1066 commonsourceibias.n589 gnd 0.008037f
C1067 commonsourceibias.n590 gnd 0.008037f
C1068 commonsourceibias.n591 gnd 0.007008f
C1069 commonsourceibias.n592 gnd 0.011217f
C1070 commonsourceibias.n593 gnd 0.059912f
C1071 commonsourceibias.n594 gnd 0.01122f
C1072 commonsourceibias.n595 gnd 0.008037f
C1073 commonsourceibias.n596 gnd 0.008037f
C1074 commonsourceibias.n597 gnd 0.008037f
C1075 commonsourceibias.n598 gnd 0.009613f
C1076 commonsourceibias.n599 gnd 0.059912f
C1077 commonsourceibias.n600 gnd 0.010282f
C1078 commonsourceibias.t130 gnd 0.150157f
C1079 commonsourceibias.n601 gnd 0.059912f
C1080 commonsourceibias.n602 gnd 0.010583f
C1081 commonsourceibias.n603 gnd 0.008037f
C1082 commonsourceibias.n604 gnd 0.008037f
C1083 commonsourceibias.n605 gnd 0.008037f
C1084 commonsourceibias.n606 gnd 0.006868f
C1085 commonsourceibias.n607 gnd 0.011203f
C1086 commonsourceibias.n608 gnd 0.059912f
C1087 commonsourceibias.n609 gnd 0.01121f
C1088 commonsourceibias.n610 gnd 0.008037f
C1089 commonsourceibias.n611 gnd 0.008037f
C1090 commonsourceibias.n612 gnd 0.008037f
C1091 commonsourceibias.n613 gnd 0.009378f
C1092 commonsourceibias.n614 gnd 0.059912f
C1093 commonsourceibias.n615 gnd 0.009861f
C1094 commonsourceibias.n616 gnd 0.07189f
C1095 commonsourceibias.n617 gnd 0.04697f
C1096 commonsourceibias.n618 gnd 0.010724f
C1097 commonsourceibias.t142 gnd 0.150157f
C1098 commonsourceibias.n619 gnd 0.007823f
C1099 commonsourceibias.n620 gnd 0.008037f
C1100 commonsourceibias.t156 gnd 0.150157f
C1101 commonsourceibias.n621 gnd 0.01034f
C1102 commonsourceibias.n622 gnd 0.008037f
C1103 commonsourceibias.t132 gnd 0.150157f
C1104 commonsourceibias.n623 gnd 0.007578f
C1105 commonsourceibias.n624 gnd 0.008037f
C1106 commonsourceibias.t149 gnd 0.150157f
C1107 commonsourceibias.n625 gnd 0.010186f
C1108 commonsourceibias.n626 gnd 0.008037f
C1109 commonsourceibias.t97 gnd 0.150157f
C1110 commonsourceibias.n627 gnd 0.007361f
C1111 commonsourceibias.n628 gnd 0.008037f
C1112 commonsourceibias.t141 gnd 0.150157f
C1113 commonsourceibias.n629 gnd 0.010015f
C1114 commonsourceibias.n630 gnd 0.008037f
C1115 commonsourceibias.t152 gnd 0.150157f
C1116 commonsourceibias.n631 gnd 0.007172f
C1117 commonsourceibias.n632 gnd 0.008037f
C1118 commonsourceibias.t131 gnd 0.150157f
C1119 commonsourceibias.n633 gnd 0.009825f
C1120 commonsourceibias.n634 gnd 0.008037f
C1121 commonsourceibias.t145 gnd 0.150157f
C1122 commonsourceibias.n635 gnd 0.007008f
C1123 commonsourceibias.n636 gnd 0.008037f
C1124 commonsourceibias.t91 gnd 0.150157f
C1125 commonsourceibias.n637 gnd 0.009613f
C1126 commonsourceibias.n638 gnd 0.008037f
C1127 commonsourceibias.t116 gnd 0.150157f
C1128 commonsourceibias.n639 gnd 0.006868f
C1129 commonsourceibias.n640 gnd 0.008037f
C1130 commonsourceibias.t134 gnd 0.150157f
C1131 commonsourceibias.n641 gnd 0.009378f
C1132 commonsourceibias.t106 gnd 0.166947f
C1133 commonsourceibias.t90 gnd 0.150157f
C1134 commonsourceibias.n642 gnd 0.065449f
C1135 commonsourceibias.n643 gnd 0.071822f
C1136 commonsourceibias.n644 gnd 0.033327f
C1137 commonsourceibias.n645 gnd 0.008037f
C1138 commonsourceibias.n646 gnd 0.007823f
C1139 commonsourceibias.n647 gnd 0.01121f
C1140 commonsourceibias.n648 gnd 0.059912f
C1141 commonsourceibias.n649 gnd 0.011203f
C1142 commonsourceibias.n650 gnd 0.008037f
C1143 commonsourceibias.n651 gnd 0.008037f
C1144 commonsourceibias.n652 gnd 0.008037f
C1145 commonsourceibias.n653 gnd 0.01034f
C1146 commonsourceibias.n654 gnd 0.059912f
C1147 commonsourceibias.n655 gnd 0.010583f
C1148 commonsourceibias.t96 gnd 0.150157f
C1149 commonsourceibias.n656 gnd 0.059912f
C1150 commonsourceibias.n657 gnd 0.010282f
C1151 commonsourceibias.n658 gnd 0.008037f
C1152 commonsourceibias.n659 gnd 0.008037f
C1153 commonsourceibias.n660 gnd 0.008037f
C1154 commonsourceibias.n661 gnd 0.007578f
C1155 commonsourceibias.n662 gnd 0.01122f
C1156 commonsourceibias.n663 gnd 0.059912f
C1157 commonsourceibias.n664 gnd 0.011217f
C1158 commonsourceibias.n665 gnd 0.008037f
C1159 commonsourceibias.n666 gnd 0.008037f
C1160 commonsourceibias.n667 gnd 0.008037f
C1161 commonsourceibias.n668 gnd 0.010186f
C1162 commonsourceibias.n669 gnd 0.059912f
C1163 commonsourceibias.n670 gnd 0.010507f
C1164 commonsourceibias.t124 gnd 0.150157f
C1165 commonsourceibias.n671 gnd 0.059912f
C1166 commonsourceibias.n672 gnd 0.010357f
C1167 commonsourceibias.n673 gnd 0.008037f
C1168 commonsourceibias.n674 gnd 0.008037f
C1169 commonsourceibias.n675 gnd 0.008037f
C1170 commonsourceibias.n676 gnd 0.007361f
C1171 commonsourceibias.n677 gnd 0.011225f
C1172 commonsourceibias.n678 gnd 0.059912f
C1173 commonsourceibias.n679 gnd 0.011224f
C1174 commonsourceibias.n680 gnd 0.008037f
C1175 commonsourceibias.n681 gnd 0.008037f
C1176 commonsourceibias.n682 gnd 0.008037f
C1177 commonsourceibias.n683 gnd 0.010015f
C1178 commonsourceibias.n684 gnd 0.059912f
C1179 commonsourceibias.n685 gnd 0.010432f
C1180 commonsourceibias.t157 gnd 0.150157f
C1181 commonsourceibias.n686 gnd 0.059912f
C1182 commonsourceibias.n687 gnd 0.010432f
C1183 commonsourceibias.n688 gnd 0.008037f
C1184 commonsourceibias.n689 gnd 0.008037f
C1185 commonsourceibias.n690 gnd 0.008037f
C1186 commonsourceibias.n691 gnd 0.007172f
C1187 commonsourceibias.n692 gnd 0.011224f
C1188 commonsourceibias.n693 gnd 0.059912f
C1189 commonsourceibias.n694 gnd 0.011225f
C1190 commonsourceibias.n695 gnd 0.008037f
C1191 commonsourceibias.n696 gnd 0.008037f
C1192 commonsourceibias.n697 gnd 0.008037f
C1193 commonsourceibias.n698 gnd 0.009825f
C1194 commonsourceibias.n699 gnd 0.059912f
C1195 commonsourceibias.n700 gnd 0.010357f
C1196 commonsourceibias.t81 gnd 0.150157f
C1197 commonsourceibias.n701 gnd 0.059912f
C1198 commonsourceibias.n702 gnd 0.010507f
C1199 commonsourceibias.n703 gnd 0.008037f
C1200 commonsourceibias.n704 gnd 0.008037f
C1201 commonsourceibias.n705 gnd 0.008037f
C1202 commonsourceibias.n706 gnd 0.007008f
C1203 commonsourceibias.n707 gnd 0.011217f
C1204 commonsourceibias.n708 gnd 0.059912f
C1205 commonsourceibias.n709 gnd 0.01122f
C1206 commonsourceibias.n710 gnd 0.008037f
C1207 commonsourceibias.n711 gnd 0.008037f
C1208 commonsourceibias.n712 gnd 0.008037f
C1209 commonsourceibias.n713 gnd 0.009613f
C1210 commonsourceibias.n714 gnd 0.059912f
C1211 commonsourceibias.n715 gnd 0.010282f
C1212 commonsourceibias.t111 gnd 0.150157f
C1213 commonsourceibias.n716 gnd 0.059912f
C1214 commonsourceibias.n717 gnd 0.010583f
C1215 commonsourceibias.n718 gnd 0.008037f
C1216 commonsourceibias.n719 gnd 0.008037f
C1217 commonsourceibias.n720 gnd 0.008037f
C1218 commonsourceibias.n721 gnd 0.006868f
C1219 commonsourceibias.n722 gnd 0.011203f
C1220 commonsourceibias.n723 gnd 0.059912f
C1221 commonsourceibias.n724 gnd 0.01121f
C1222 commonsourceibias.n725 gnd 0.008037f
C1223 commonsourceibias.n726 gnd 0.008037f
C1224 commonsourceibias.n727 gnd 0.008037f
C1225 commonsourceibias.n728 gnd 0.009378f
C1226 commonsourceibias.n729 gnd 0.059912f
C1227 commonsourceibias.n730 gnd 0.009861f
C1228 commonsourceibias.t122 gnd 0.162395f
C1229 commonsourceibias.n731 gnd 0.07189f
C1230 commonsourceibias.n732 gnd 0.025003f
C1231 commonsourceibias.n733 gnd 0.221951f
C1232 commonsourceibias.n734 gnd 4.85761f
C1233 diffpairibias.t27 gnd 0.090128f
C1234 diffpairibias.t23 gnd 0.08996f
C1235 diffpairibias.n0 gnd 0.105991f
C1236 diffpairibias.t28 gnd 0.08996f
C1237 diffpairibias.n1 gnd 0.051736f
C1238 diffpairibias.t25 gnd 0.08996f
C1239 diffpairibias.n2 gnd 0.051736f
C1240 diffpairibias.t29 gnd 0.08996f
C1241 diffpairibias.n3 gnd 0.041084f
C1242 diffpairibias.t15 gnd 0.086371f
C1243 diffpairibias.t1 gnd 0.085993f
C1244 diffpairibias.n4 gnd 0.13579f
C1245 diffpairibias.t11 gnd 0.085993f
C1246 diffpairibias.n5 gnd 0.072463f
C1247 diffpairibias.t13 gnd 0.085993f
C1248 diffpairibias.n6 gnd 0.072463f
C1249 diffpairibias.t7 gnd 0.085993f
C1250 diffpairibias.n7 gnd 0.072463f
C1251 diffpairibias.t3 gnd 0.085993f
C1252 diffpairibias.n8 gnd 0.072463f
C1253 diffpairibias.t17 gnd 0.085993f
C1254 diffpairibias.n9 gnd 0.072463f
C1255 diffpairibias.t5 gnd 0.085993f
C1256 diffpairibias.n10 gnd 0.072463f
C1257 diffpairibias.t19 gnd 0.085993f
C1258 diffpairibias.n11 gnd 0.072463f
C1259 diffpairibias.t9 gnd 0.085993f
C1260 diffpairibias.n12 gnd 0.102883f
C1261 diffpairibias.t14 gnd 0.086899f
C1262 diffpairibias.t0 gnd 0.086748f
C1263 diffpairibias.n13 gnd 0.094648f
C1264 diffpairibias.t10 gnd 0.086748f
C1265 diffpairibias.n14 gnd 0.052262f
C1266 diffpairibias.t12 gnd 0.086748f
C1267 diffpairibias.n15 gnd 0.052262f
C1268 diffpairibias.t6 gnd 0.086748f
C1269 diffpairibias.n16 gnd 0.052262f
C1270 diffpairibias.t2 gnd 0.086748f
C1271 diffpairibias.n17 gnd 0.052262f
C1272 diffpairibias.t16 gnd 0.086748f
C1273 diffpairibias.n18 gnd 0.052262f
C1274 diffpairibias.t4 gnd 0.086748f
C1275 diffpairibias.n19 gnd 0.052262f
C1276 diffpairibias.t18 gnd 0.086748f
C1277 diffpairibias.n20 gnd 0.052262f
C1278 diffpairibias.t8 gnd 0.086748f
C1279 diffpairibias.n21 gnd 0.061849f
C1280 diffpairibias.n22 gnd 0.233513f
C1281 diffpairibias.t20 gnd 0.08996f
C1282 diffpairibias.n23 gnd 0.051747f
C1283 diffpairibias.t26 gnd 0.08996f
C1284 diffpairibias.n24 gnd 0.051736f
C1285 diffpairibias.t22 gnd 0.08996f
C1286 diffpairibias.n25 gnd 0.051736f
C1287 diffpairibias.t21 gnd 0.08996f
C1288 diffpairibias.n26 gnd 0.051736f
C1289 diffpairibias.t24 gnd 0.08996f
C1290 diffpairibias.n27 gnd 0.04729f
C1291 diffpairibias.n28 gnd 0.047711f
C1292 outputibias.t10 gnd 0.11477f
C1293 outputibias.t8 gnd 0.115567f
C1294 outputibias.n0 gnd 0.130108f
C1295 outputibias.n1 gnd 0.001372f
C1296 outputibias.n2 gnd 9.76e-19
C1297 outputibias.n3 gnd 5.24e-19
C1298 outputibias.n4 gnd 0.001239f
C1299 outputibias.n5 gnd 5.55e-19
C1300 outputibias.n6 gnd 9.76e-19
C1301 outputibias.n7 gnd 5.24e-19
C1302 outputibias.n8 gnd 0.001239f
C1303 outputibias.n9 gnd 5.55e-19
C1304 outputibias.n10 gnd 0.004176f
C1305 outputibias.t5 gnd 0.00202f
C1306 outputibias.n11 gnd 9.3e-19
C1307 outputibias.n12 gnd 7.32e-19
C1308 outputibias.n13 gnd 5.24e-19
C1309 outputibias.n14 gnd 0.02322f
C1310 outputibias.n15 gnd 9.76e-19
C1311 outputibias.n16 gnd 5.24e-19
C1312 outputibias.n17 gnd 5.55e-19
C1313 outputibias.n18 gnd 0.001239f
C1314 outputibias.n19 gnd 0.001239f
C1315 outputibias.n20 gnd 5.55e-19
C1316 outputibias.n21 gnd 5.24e-19
C1317 outputibias.n22 gnd 9.76e-19
C1318 outputibias.n23 gnd 9.76e-19
C1319 outputibias.n24 gnd 5.24e-19
C1320 outputibias.n25 gnd 5.55e-19
C1321 outputibias.n26 gnd 0.001239f
C1322 outputibias.n27 gnd 0.002683f
C1323 outputibias.n28 gnd 5.55e-19
C1324 outputibias.n29 gnd 5.24e-19
C1325 outputibias.n30 gnd 0.002256f
C1326 outputibias.n31 gnd 0.005781f
C1327 outputibias.n32 gnd 0.001372f
C1328 outputibias.n33 gnd 9.76e-19
C1329 outputibias.n34 gnd 5.24e-19
C1330 outputibias.n35 gnd 0.001239f
C1331 outputibias.n36 gnd 5.55e-19
C1332 outputibias.n37 gnd 9.76e-19
C1333 outputibias.n38 gnd 5.24e-19
C1334 outputibias.n39 gnd 0.001239f
C1335 outputibias.n40 gnd 5.55e-19
C1336 outputibias.n41 gnd 0.004176f
C1337 outputibias.t3 gnd 0.00202f
C1338 outputibias.n42 gnd 9.3e-19
C1339 outputibias.n43 gnd 7.32e-19
C1340 outputibias.n44 gnd 5.24e-19
C1341 outputibias.n45 gnd 0.02322f
C1342 outputibias.n46 gnd 9.76e-19
C1343 outputibias.n47 gnd 5.24e-19
C1344 outputibias.n48 gnd 5.55e-19
C1345 outputibias.n49 gnd 0.001239f
C1346 outputibias.n50 gnd 0.001239f
C1347 outputibias.n51 gnd 5.55e-19
C1348 outputibias.n52 gnd 5.24e-19
C1349 outputibias.n53 gnd 9.76e-19
C1350 outputibias.n54 gnd 9.76e-19
C1351 outputibias.n55 gnd 5.24e-19
C1352 outputibias.n56 gnd 5.55e-19
C1353 outputibias.n57 gnd 0.001239f
C1354 outputibias.n58 gnd 0.002683f
C1355 outputibias.n59 gnd 5.55e-19
C1356 outputibias.n60 gnd 5.24e-19
C1357 outputibias.n61 gnd 0.002256f
C1358 outputibias.n62 gnd 0.005197f
C1359 outputibias.n63 gnd 0.121892f
C1360 outputibias.n64 gnd 0.001372f
C1361 outputibias.n65 gnd 9.76e-19
C1362 outputibias.n66 gnd 5.24e-19
C1363 outputibias.n67 gnd 0.001239f
C1364 outputibias.n68 gnd 5.55e-19
C1365 outputibias.n69 gnd 9.76e-19
C1366 outputibias.n70 gnd 5.24e-19
C1367 outputibias.n71 gnd 0.001239f
C1368 outputibias.n72 gnd 5.55e-19
C1369 outputibias.n73 gnd 0.004176f
C1370 outputibias.t1 gnd 0.00202f
C1371 outputibias.n74 gnd 9.3e-19
C1372 outputibias.n75 gnd 7.32e-19
C1373 outputibias.n76 gnd 5.24e-19
C1374 outputibias.n77 gnd 0.02322f
C1375 outputibias.n78 gnd 9.76e-19
C1376 outputibias.n79 gnd 5.24e-19
C1377 outputibias.n80 gnd 5.55e-19
C1378 outputibias.n81 gnd 0.001239f
C1379 outputibias.n82 gnd 0.001239f
C1380 outputibias.n83 gnd 5.55e-19
C1381 outputibias.n84 gnd 5.24e-19
C1382 outputibias.n85 gnd 9.76e-19
C1383 outputibias.n86 gnd 9.76e-19
C1384 outputibias.n87 gnd 5.24e-19
C1385 outputibias.n88 gnd 5.55e-19
C1386 outputibias.n89 gnd 0.001239f
C1387 outputibias.n90 gnd 0.002683f
C1388 outputibias.n91 gnd 5.55e-19
C1389 outputibias.n92 gnd 5.24e-19
C1390 outputibias.n93 gnd 0.002256f
C1391 outputibias.n94 gnd 0.005197f
C1392 outputibias.n95 gnd 0.064513f
C1393 outputibias.n96 gnd 0.001372f
C1394 outputibias.n97 gnd 9.76e-19
C1395 outputibias.n98 gnd 5.24e-19
C1396 outputibias.n99 gnd 0.001239f
C1397 outputibias.n100 gnd 5.55e-19
C1398 outputibias.n101 gnd 9.76e-19
C1399 outputibias.n102 gnd 5.24e-19
C1400 outputibias.n103 gnd 0.001239f
C1401 outputibias.n104 gnd 5.55e-19
C1402 outputibias.n105 gnd 0.004176f
C1403 outputibias.t7 gnd 0.00202f
C1404 outputibias.n106 gnd 9.3e-19
C1405 outputibias.n107 gnd 7.32e-19
C1406 outputibias.n108 gnd 5.24e-19
C1407 outputibias.n109 gnd 0.02322f
C1408 outputibias.n110 gnd 9.76e-19
C1409 outputibias.n111 gnd 5.24e-19
C1410 outputibias.n112 gnd 5.55e-19
C1411 outputibias.n113 gnd 0.001239f
C1412 outputibias.n114 gnd 0.001239f
C1413 outputibias.n115 gnd 5.55e-19
C1414 outputibias.n116 gnd 5.24e-19
C1415 outputibias.n117 gnd 9.76e-19
C1416 outputibias.n118 gnd 9.76e-19
C1417 outputibias.n119 gnd 5.24e-19
C1418 outputibias.n120 gnd 5.55e-19
C1419 outputibias.n121 gnd 0.001239f
C1420 outputibias.n122 gnd 0.002683f
C1421 outputibias.n123 gnd 5.55e-19
C1422 outputibias.n124 gnd 5.24e-19
C1423 outputibias.n125 gnd 0.002256f
C1424 outputibias.n126 gnd 0.005197f
C1425 outputibias.n127 gnd 0.084814f
C1426 outputibias.t6 gnd 0.108319f
C1427 outputibias.t0 gnd 0.108319f
C1428 outputibias.t2 gnd 0.108319f
C1429 outputibias.t4 gnd 0.109238f
C1430 outputibias.n128 gnd 0.134674f
C1431 outputibias.n129 gnd 0.07244f
C1432 outputibias.n130 gnd 0.079818f
C1433 outputibias.n131 gnd 0.164901f
C1434 outputibias.t11 gnd 0.11477f
C1435 outputibias.n132 gnd 0.067481f
C1436 outputibias.t9 gnd 0.11477f
C1437 outputibias.n133 gnd 0.065115f
C1438 outputibias.n134 gnd 0.029159f
C1439 a_n2140_13878.t11 gnd 0.186868f
C1440 a_n2140_13878.t10 gnd 0.186868f
C1441 a_n2140_13878.t5 gnd 0.186868f
C1442 a_n2140_13878.n0 gnd 1.47299f
C1443 a_n2140_13878.t2 gnd 0.186868f
C1444 a_n2140_13878.t4 gnd 0.186868f
C1445 a_n2140_13878.n1 gnd 1.47143f
C1446 a_n2140_13878.n2 gnd 2.05603f
C1447 a_n2140_13878.t12 gnd 0.186868f
C1448 a_n2140_13878.t3 gnd 0.186868f
C1449 a_n2140_13878.n3 gnd 1.47143f
C1450 a_n2140_13878.n4 gnd 1.00289f
C1451 a_n2140_13878.t9 gnd 0.186868f
C1452 a_n2140_13878.t1 gnd 0.186868f
C1453 a_n2140_13878.n5 gnd 1.47143f
C1454 a_n2140_13878.n6 gnd 4.06212f
C1455 a_n2140_13878.t17 gnd 1.74974f
C1456 a_n2140_13878.t20 gnd 0.186868f
C1457 a_n2140_13878.t21 gnd 0.186868f
C1458 a_n2140_13878.n7 gnd 1.3163f
C1459 a_n2140_13878.n8 gnd 1.47077f
C1460 a_n2140_13878.t16 gnd 1.74626f
C1461 a_n2140_13878.n9 gnd 0.740113f
C1462 a_n2140_13878.t19 gnd 1.74626f
C1463 a_n2140_13878.n10 gnd 0.740113f
C1464 a_n2140_13878.t22 gnd 0.186868f
C1465 a_n2140_13878.t23 gnd 0.186868f
C1466 a_n2140_13878.n11 gnd 1.3163f
C1467 a_n2140_13878.n12 gnd 0.74728f
C1468 a_n2140_13878.t18 gnd 1.74626f
C1469 a_n2140_13878.n13 gnd 2.09583f
C1470 a_n2140_13878.n14 gnd 2.85974f
C1471 a_n2140_13878.t6 gnd 0.186868f
C1472 a_n2140_13878.t7 gnd 0.186868f
C1473 a_n2140_13878.n15 gnd 1.47142f
C1474 a_n2140_13878.n16 gnd 2.01665f
C1475 a_n2140_13878.t13 gnd 0.186868f
C1476 a_n2140_13878.t14 gnd 0.186868f
C1477 a_n2140_13878.n17 gnd 1.47143f
C1478 a_n2140_13878.n18 gnd 0.651951f
C1479 a_n2140_13878.t0 gnd 0.186868f
C1480 a_n2140_13878.t8 gnd 0.186868f
C1481 a_n2140_13878.n19 gnd 1.47143f
C1482 a_n2140_13878.n20 gnd 1.32263f
C1483 a_n2140_13878.n21 gnd 1.47386f
C1484 a_n2140_13878.t15 gnd 0.186868f
C1485 a_n2318_13878.n0 gnd 0.814024f
C1486 a_n2318_13878.n1 gnd 3.30896f
C1487 a_n2318_13878.n2 gnd 3.13757f
C1488 a_n2318_13878.n3 gnd 3.87452f
C1489 a_n2318_13878.n4 gnd 0.663692f
C1490 a_n2318_13878.n5 gnd 0.20341f
C1491 a_n2318_13878.n6 gnd 0.149815f
C1492 a_n2318_13878.n7 gnd 0.235462f
C1493 a_n2318_13878.n8 gnd 0.181867f
C1494 a_n2318_13878.n9 gnd 0.20341f
C1495 a_n2318_13878.n10 gnd 0.149815f
C1496 a_n2318_13878.n11 gnd 0.717286f
C1497 a_n2318_13878.n12 gnd 0.508687f
C1498 a_n2318_13878.n13 gnd 0.214378f
C1499 a_n2318_13878.n14 gnd 0.214378f
C1500 a_n2318_13878.n15 gnd 0.440597f
C1501 a_n2318_13878.n16 gnd 0.214378f
C1502 a_n2318_13878.n17 gnd 0.214378f
C1503 a_n2318_13878.n18 gnd 0.663715f
C1504 a_n2318_13878.n19 gnd 0.214378f
C1505 a_n2318_13878.n20 gnd 0.214378f
C1506 a_n2318_13878.n21 gnd 0.741582f
C1507 a_n2318_13878.n22 gnd 0.214378f
C1508 a_n2318_13878.n23 gnd 0.440597f
C1509 a_n2318_13878.n24 gnd 1.76495f
C1510 a_n2318_13878.n25 gnd 1.88382f
C1511 a_n2318_13878.n26 gnd 1.76495f
C1512 a_n2318_13878.n27 gnd 2.06406f
C1513 a_n2318_13878.n28 gnd 3.19629f
C1514 a_n2318_13878.n29 gnd 0.283193f
C1515 a_n2318_13878.n30 gnd 0.004818f
C1516 a_n2318_13878.n31 gnd 0.010421f
C1517 a_n2318_13878.n32 gnd 0.010421f
C1518 a_n2318_13878.n33 gnd 0.004818f
C1519 a_n2318_13878.n34 gnd 1.43973f
C1520 a_n2318_13878.n35 gnd 0.283193f
C1521 a_n2318_13878.n36 gnd 0.283193f
C1522 a_n2318_13878.n37 gnd 0.004818f
C1523 a_n2318_13878.n38 gnd 0.010421f
C1524 a_n2318_13878.n39 gnd 0.107189f
C1525 a_n2318_13878.n40 gnd 0.010421f
C1526 a_n2318_13878.n41 gnd 0.004818f
C1527 a_n2318_13878.n42 gnd 0.283193f
C1528 a_n2318_13878.n43 gnd 0.754458f
C1529 a_n2318_13878.n44 gnd 0.004818f
C1530 a_n2318_13878.n45 gnd 0.010421f
C1531 a_n2318_13878.n46 gnd 0.010421f
C1532 a_n2318_13878.n47 gnd 0.004818f
C1533 a_n2318_13878.n48 gnd 0.283193f
C1534 a_n2318_13878.n49 gnd 0.283193f
C1535 a_n2318_13878.n50 gnd 0.440597f
C1536 a_n2318_13878.n51 gnd 0.004818f
C1537 a_n2318_13878.n52 gnd 0.010421f
C1538 a_n2318_13878.n53 gnd 0.010421f
C1539 a_n2318_13878.n54 gnd 0.004818f
C1540 a_n2318_13878.n55 gnd 0.283193f
C1541 a_n2318_13878.n56 gnd 0.0083f
C1542 a_n2318_13878.n57 gnd 0.283193f
C1543 a_n2318_13878.n58 gnd 0.0083f
C1544 a_n2318_13878.n59 gnd 0.283193f
C1545 a_n2318_13878.n60 gnd 0.0083f
C1546 a_n2318_13878.n61 gnd 0.283193f
C1547 a_n2318_13878.n62 gnd 0.0083f
C1548 a_n2318_13878.n63 gnd 0.283193f
C1549 a_n2318_13878.n64 gnd 0.283193f
C1550 a_n2318_13878.t37 gnd 1.39231f
C1551 a_n2318_13878.t15 gnd 0.148695f
C1552 a_n2318_13878.t25 gnd 0.148695f
C1553 a_n2318_13878.n65 gnd 1.04741f
C1554 a_n2318_13878.t17 gnd 0.148695f
C1555 a_n2318_13878.t27 gnd 0.148695f
C1556 a_n2318_13878.n66 gnd 1.04741f
C1557 a_n2318_13878.t13 gnd 0.148695f
C1558 a_n2318_13878.t33 gnd 0.148695f
C1559 a_n2318_13878.n67 gnd 1.04741f
C1560 a_n2318_13878.t12 gnd 0.691658f
C1561 a_n2318_13878.n68 gnd 0.302141f
C1562 a_n2318_13878.t16 gnd 0.691658f
C1563 a_n2318_13878.t36 gnd 0.703247f
C1564 a_n2318_13878.t14 gnd 0.691658f
C1565 a_n2318_13878.t62 gnd 0.691658f
C1566 a_n2318_13878.n69 gnd 0.302141f
C1567 a_n2318_13878.t76 gnd 0.691658f
C1568 a_n2318_13878.t78 gnd 0.703247f
C1569 a_n2318_13878.t56 gnd 0.691658f
C1570 a_n2318_13878.t18 gnd 0.703247f
C1571 a_n2318_13878.t38 gnd 0.691658f
C1572 a_n2318_13878.t20 gnd 0.691658f
C1573 a_n2318_13878.n70 gnd 0.302141f
C1574 a_n2318_13878.t34 gnd 0.691658f
C1575 a_n2318_13878.t10 gnd 0.691658f
C1576 a_n2318_13878.t30 gnd 0.691658f
C1577 a_n2318_13878.n71 gnd 0.302141f
C1578 a_n2318_13878.t22 gnd 0.691658f
C1579 a_n2318_13878.t28 gnd 0.703247f
C1580 a_n2318_13878.t7 gnd 0.115652f
C1581 a_n2318_13878.t51 gnd 0.115652f
C1582 a_n2318_13878.n72 gnd 1.02421f
C1583 a_n2318_13878.t41 gnd 0.115652f
C1584 a_n2318_13878.t2 gnd 0.115652f
C1585 a_n2318_13878.n73 gnd 1.02194f
C1586 a_n2318_13878.t6 gnd 0.115652f
C1587 a_n2318_13878.t5 gnd 0.115652f
C1588 a_n2318_13878.n74 gnd 1.02194f
C1589 a_n2318_13878.t47 gnd 0.115652f
C1590 a_n2318_13878.t1 gnd 0.115652f
C1591 a_n2318_13878.n75 gnd 1.02421f
C1592 a_n2318_13878.t4 gnd 0.115652f
C1593 a_n2318_13878.t46 gnd 0.115652f
C1594 a_n2318_13878.n76 gnd 1.02194f
C1595 a_n2318_13878.t42 gnd 0.115652f
C1596 a_n2318_13878.t40 gnd 0.115652f
C1597 a_n2318_13878.n77 gnd 1.02194f
C1598 a_n2318_13878.t44 gnd 0.115652f
C1599 a_n2318_13878.t0 gnd 0.115652f
C1600 a_n2318_13878.n78 gnd 1.02194f
C1601 a_n2318_13878.t49 gnd 0.115652f
C1602 a_n2318_13878.t50 gnd 0.115652f
C1603 a_n2318_13878.n79 gnd 1.02194f
C1604 a_n2318_13878.t3 gnd 0.115652f
C1605 a_n2318_13878.t43 gnd 0.115652f
C1606 a_n2318_13878.n80 gnd 1.02421f
C1607 a_n2318_13878.t48 gnd 0.115652f
C1608 a_n2318_13878.t45 gnd 0.115652f
C1609 a_n2318_13878.n81 gnd 1.02194f
C1610 a_n2318_13878.t82 gnd 0.703247f
C1611 a_n2318_13878.t63 gnd 0.691658f
C1612 a_n2318_13878.t67 gnd 0.691658f
C1613 a_n2318_13878.n82 gnd 0.302141f
C1614 a_n2318_13878.t57 gnd 0.691658f
C1615 a_n2318_13878.t72 gnd 0.691658f
C1616 a_n2318_13878.t79 gnd 0.691658f
C1617 a_n2318_13878.n83 gnd 0.302141f
C1618 a_n2318_13878.t80 gnd 0.691658f
C1619 a_n2318_13878.t54 gnd 0.703247f
C1620 a_n2318_13878.n84 gnd 0.304604f
C1621 a_n2318_13878.n85 gnd 0.297591f
C1622 a_n2318_13878.n86 gnd 0.297591f
C1623 a_n2318_13878.n87 gnd 0.304604f
C1624 a_n2318_13878.n88 gnd 0.304604f
C1625 a_n2318_13878.n89 gnd 0.297591f
C1626 a_n2318_13878.n90 gnd 0.297591f
C1627 a_n2318_13878.n91 gnd 0.304604f
C1628 a_n2318_13878.t29 gnd 1.39231f
C1629 a_n2318_13878.t31 gnd 0.148695f
C1630 a_n2318_13878.t23 gnd 0.148695f
C1631 a_n2318_13878.n92 gnd 1.04741f
C1632 a_n2318_13878.t35 gnd 0.148695f
C1633 a_n2318_13878.t11 gnd 0.148695f
C1634 a_n2318_13878.n93 gnd 1.04741f
C1635 a_n2318_13878.t39 gnd 0.148695f
C1636 a_n2318_13878.t21 gnd 0.148695f
C1637 a_n2318_13878.n94 gnd 1.04741f
C1638 a_n2318_13878.t19 gnd 1.38953f
C1639 a_n2318_13878.n95 gnd 0.853399f
C1640 a_n2318_13878.t61 gnd 0.691658f
C1641 a_n2318_13878.t70 gnd 0.691658f
C1642 a_n2318_13878.t83 gnd 0.691658f
C1643 a_n2318_13878.n96 gnd 0.304097f
C1644 a_n2318_13878.t73 gnd 0.691658f
C1645 a_n2318_13878.t58 gnd 0.691658f
C1646 a_n2318_13878.t59 gnd 0.691658f
C1647 a_n2318_13878.n97 gnd 0.304097f
C1648 a_n2318_13878.t77 gnd 0.691658f
C1649 a_n2318_13878.t66 gnd 0.691658f
C1650 a_n2318_13878.t65 gnd 0.691658f
C1651 a_n2318_13878.n98 gnd 0.304097f
C1652 a_n2318_13878.t69 gnd 0.691658f
C1653 a_n2318_13878.t60 gnd 0.691658f
C1654 a_n2318_13878.t52 gnd 0.691658f
C1655 a_n2318_13878.n99 gnd 0.304097f
C1656 a_n2318_13878.t74 gnd 0.703247f
C1657 a_n2318_13878.n100 gnd 0.300235f
C1658 a_n2318_13878.n101 gnd 0.294783f
C1659 a_n2318_13878.t81 gnd 0.703247f
C1660 a_n2318_13878.n102 gnd 0.300235f
C1661 a_n2318_13878.n103 gnd 0.294783f
C1662 a_n2318_13878.t68 gnd 0.703247f
C1663 a_n2318_13878.n104 gnd 0.300235f
C1664 a_n2318_13878.n105 gnd 0.294783f
C1665 a_n2318_13878.t64 gnd 0.703247f
C1666 a_n2318_13878.n106 gnd 0.300235f
C1667 a_n2318_13878.n107 gnd 0.294783f
C1668 a_n2318_13878.n108 gnd 1.11013f
C1669 a_n2318_13878.n109 gnd 0.304604f
C1670 a_n2318_13878.t75 gnd 0.691658f
C1671 a_n2318_13878.n110 gnd 0.302141f
C1672 a_n2318_13878.n111 gnd 0.297591f
C1673 a_n2318_13878.t53 gnd 0.691658f
C1674 a_n2318_13878.n112 gnd 0.297591f
C1675 a_n2318_13878.t71 gnd 0.691658f
C1676 a_n2318_13878.n113 gnd 0.304604f
C1677 a_n2318_13878.t55 gnd 0.703247f
C1678 a_n2318_13878.n114 gnd 0.304604f
C1679 a_n2318_13878.t24 gnd 0.691658f
C1680 a_n2318_13878.n115 gnd 0.302141f
C1681 a_n2318_13878.n116 gnd 0.297591f
C1682 a_n2318_13878.t26 gnd 0.691658f
C1683 a_n2318_13878.n117 gnd 0.297591f
C1684 a_n2318_13878.t32 gnd 0.691658f
C1685 a_n2318_13878.n118 gnd 0.304604f
C1686 a_n2318_13878.t8 gnd 0.703247f
C1687 a_n2318_13878.n119 gnd 1.18985f
C1688 a_n2318_13878.t9 gnd 1.38954f
C1689 CSoutput.n0 gnd 0.044633f
C1690 CSoutput.t193 gnd 0.295236f
C1691 CSoutput.n1 gnd 0.133314f
C1692 CSoutput.n2 gnd 0.044633f
C1693 CSoutput.t176 gnd 0.295236f
C1694 CSoutput.n3 gnd 0.035375f
C1695 CSoutput.n4 gnd 0.044633f
C1696 CSoutput.t185 gnd 0.295236f
C1697 CSoutput.n5 gnd 0.030504f
C1698 CSoutput.n6 gnd 0.044633f
C1699 CSoutput.t196 gnd 0.295236f
C1700 CSoutput.t195 gnd 0.295236f
C1701 CSoutput.n7 gnd 0.131861f
C1702 CSoutput.n8 gnd 0.044633f
C1703 CSoutput.t182 gnd 0.295236f
C1704 CSoutput.n9 gnd 0.029084f
C1705 CSoutput.n10 gnd 0.044633f
C1706 CSoutput.t188 gnd 0.295236f
C1707 CSoutput.t191 gnd 0.295236f
C1708 CSoutput.n11 gnd 0.131861f
C1709 CSoutput.n12 gnd 0.044633f
C1710 CSoutput.t179 gnd 0.295236f
C1711 CSoutput.n13 gnd 0.030504f
C1712 CSoutput.n14 gnd 0.044633f
C1713 CSoutput.t178 gnd 0.295236f
C1714 CSoutput.t189 gnd 0.295236f
C1715 CSoutput.n15 gnd 0.131861f
C1716 CSoutput.n16 gnd 0.044633f
C1717 CSoutput.t194 gnd 0.295236f
C1718 CSoutput.n17 gnd 0.03258f
C1719 CSoutput.t180 gnd 0.352814f
C1720 CSoutput.t177 gnd 0.295236f
C1721 CSoutput.n18 gnd 0.168335f
C1722 CSoutput.n19 gnd 0.163343f
C1723 CSoutput.n20 gnd 0.189497f
C1724 CSoutput.n21 gnd 0.044633f
C1725 CSoutput.n22 gnd 0.037251f
C1726 CSoutput.n23 gnd 0.131861f
C1727 CSoutput.n24 gnd 0.035909f
C1728 CSoutput.n25 gnd 0.035375f
C1729 CSoutput.n26 gnd 0.044633f
C1730 CSoutput.n27 gnd 0.044633f
C1731 CSoutput.n28 gnd 0.036965f
C1732 CSoutput.n29 gnd 0.031384f
C1733 CSoutput.n30 gnd 0.134796f
C1734 CSoutput.n31 gnd 0.031816f
C1735 CSoutput.n32 gnd 0.044633f
C1736 CSoutput.n33 gnd 0.044633f
C1737 CSoutput.n34 gnd 0.044633f
C1738 CSoutput.n35 gnd 0.036571f
C1739 CSoutput.n36 gnd 0.131861f
C1740 CSoutput.n37 gnd 0.034975f
C1741 CSoutput.n38 gnd 0.036309f
C1742 CSoutput.n39 gnd 0.044633f
C1743 CSoutput.n40 gnd 0.044633f
C1744 CSoutput.n41 gnd 0.037243f
C1745 CSoutput.n42 gnd 0.03404f
C1746 CSoutput.n43 gnd 0.131861f
C1747 CSoutput.n44 gnd 0.034903f
C1748 CSoutput.n45 gnd 0.044633f
C1749 CSoutput.n46 gnd 0.044633f
C1750 CSoutput.n47 gnd 0.044633f
C1751 CSoutput.n48 gnd 0.034903f
C1752 CSoutput.n49 gnd 0.131861f
C1753 CSoutput.n50 gnd 0.03404f
C1754 CSoutput.n51 gnd 0.037243f
C1755 CSoutput.n52 gnd 0.044633f
C1756 CSoutput.n53 gnd 0.044633f
C1757 CSoutput.n54 gnd 0.036309f
C1758 CSoutput.n55 gnd 0.034975f
C1759 CSoutput.n56 gnd 0.131861f
C1760 CSoutput.n57 gnd 0.036571f
C1761 CSoutput.n58 gnd 0.044633f
C1762 CSoutput.n59 gnd 0.044633f
C1763 CSoutput.n60 gnd 0.044633f
C1764 CSoutput.n61 gnd 0.031816f
C1765 CSoutput.n62 gnd 0.134796f
C1766 CSoutput.n63 gnd 0.031384f
C1767 CSoutput.t197 gnd 0.295236f
C1768 CSoutput.n64 gnd 0.131861f
C1769 CSoutput.n65 gnd 0.036965f
C1770 CSoutput.n66 gnd 0.044633f
C1771 CSoutput.n67 gnd 0.044633f
C1772 CSoutput.n68 gnd 0.044633f
C1773 CSoutput.n69 gnd 0.035909f
C1774 CSoutput.n70 gnd 0.131861f
C1775 CSoutput.n71 gnd 0.037251f
C1776 CSoutput.n72 gnd 0.03258f
C1777 CSoutput.n73 gnd 0.044633f
C1778 CSoutput.n74 gnd 0.044633f
C1779 CSoutput.n75 gnd 0.033788f
C1780 CSoutput.n76 gnd 0.020067f
C1781 CSoutput.t183 gnd 0.331718f
C1782 CSoutput.n77 gnd 0.164784f
C1783 CSoutput.n78 gnd 0.705097f
C1784 CSoutput.t139 gnd 0.055673f
C1785 CSoutput.t86 gnd 0.055673f
C1786 CSoutput.n79 gnd 0.431039f
C1787 CSoutput.t151 gnd 0.055673f
C1788 CSoutput.t103 gnd 0.055673f
C1789 CSoutput.n80 gnd 0.43027f
C1790 CSoutput.n81 gnd 0.436724f
C1791 CSoutput.t67 gnd 0.055673f
C1792 CSoutput.t115 gnd 0.055673f
C1793 CSoutput.n82 gnd 0.43027f
C1794 CSoutput.n83 gnd 0.215199f
C1795 CSoutput.t71 gnd 0.055673f
C1796 CSoutput.t95 gnd 0.055673f
C1797 CSoutput.n84 gnd 0.43027f
C1798 CSoutput.n85 gnd 0.215199f
C1799 CSoutput.t155 gnd 0.055673f
C1800 CSoutput.t110 gnd 0.055673f
C1801 CSoutput.n86 gnd 0.43027f
C1802 CSoutput.n87 gnd 0.215199f
C1803 CSoutput.t74 gnd 0.055673f
C1804 CSoutput.t143 gnd 0.055673f
C1805 CSoutput.n88 gnd 0.43027f
C1806 CSoutput.n89 gnd 0.215199f
C1807 CSoutput.t82 gnd 0.055673f
C1808 CSoutput.t125 gnd 0.055673f
C1809 CSoutput.n90 gnd 0.43027f
C1810 CSoutput.n91 gnd 0.215199f
C1811 CSoutput.t98 gnd 0.055673f
C1812 CSoutput.t116 gnd 0.055673f
C1813 CSoutput.n92 gnd 0.43027f
C1814 CSoutput.n93 gnd 0.394625f
C1815 CSoutput.t63 gnd 0.055673f
C1816 CSoutput.t137 gnd 0.055673f
C1817 CSoutput.n94 gnd 0.431039f
C1818 CSoutput.t126 gnd 0.055673f
C1819 CSoutput.t105 gnd 0.055673f
C1820 CSoutput.n95 gnd 0.43027f
C1821 CSoutput.n96 gnd 0.436724f
C1822 CSoutput.t87 gnd 0.055673f
C1823 CSoutput.t148 gnd 0.055673f
C1824 CSoutput.n97 gnd 0.43027f
C1825 CSoutput.n98 gnd 0.215199f
C1826 CSoutput.t123 gnd 0.055673f
C1827 CSoutput.t122 gnd 0.055673f
C1828 CSoutput.n99 gnd 0.43027f
C1829 CSoutput.n100 gnd 0.215199f
C1830 CSoutput.t112 gnd 0.055673f
C1831 CSoutput.t83 gnd 0.055673f
C1832 CSoutput.n101 gnd 0.43027f
C1833 CSoutput.n102 gnd 0.215199f
C1834 CSoutput.t66 gnd 0.055673f
C1835 CSoutput.t113 gnd 0.055673f
C1836 CSoutput.n103 gnd 0.43027f
C1837 CSoutput.n104 gnd 0.215199f
C1838 CSoutput.t111 gnd 0.055673f
C1839 CSoutput.t81 gnd 0.055673f
C1840 CSoutput.n105 gnd 0.43027f
C1841 CSoutput.n106 gnd 0.215199f
C1842 CSoutput.t64 gnd 0.055673f
C1843 CSoutput.t62 gnd 0.055673f
C1844 CSoutput.n107 gnd 0.43027f
C1845 CSoutput.n108 gnd 0.320916f
C1846 CSoutput.n109 gnd 0.404673f
C1847 CSoutput.t76 gnd 0.055673f
C1848 CSoutput.t147 gnd 0.055673f
C1849 CSoutput.n110 gnd 0.431039f
C1850 CSoutput.t132 gnd 0.055673f
C1851 CSoutput.t114 gnd 0.055673f
C1852 CSoutput.n111 gnd 0.43027f
C1853 CSoutput.n112 gnd 0.436724f
C1854 CSoutput.t99 gnd 0.055673f
C1855 CSoutput.t156 gnd 0.055673f
C1856 CSoutput.n113 gnd 0.43027f
C1857 CSoutput.n114 gnd 0.215199f
C1858 CSoutput.t131 gnd 0.055673f
C1859 CSoutput.t130 gnd 0.055673f
C1860 CSoutput.n115 gnd 0.43027f
C1861 CSoutput.n116 gnd 0.215199f
C1862 CSoutput.t120 gnd 0.055673f
C1863 CSoutput.t96 gnd 0.055673f
C1864 CSoutput.n117 gnd 0.43027f
C1865 CSoutput.n118 gnd 0.215199f
C1866 CSoutput.t78 gnd 0.055673f
C1867 CSoutput.t121 gnd 0.055673f
C1868 CSoutput.n119 gnd 0.43027f
C1869 CSoutput.n120 gnd 0.215199f
C1870 CSoutput.t119 gnd 0.055673f
C1871 CSoutput.t94 gnd 0.055673f
C1872 CSoutput.n121 gnd 0.43027f
C1873 CSoutput.n122 gnd 0.215199f
C1874 CSoutput.t77 gnd 0.055673f
C1875 CSoutput.t75 gnd 0.055673f
C1876 CSoutput.n123 gnd 0.43027f
C1877 CSoutput.n124 gnd 0.320916f
C1878 CSoutput.n125 gnd 0.452321f
C1879 CSoutput.n126 gnd 9.421049f
C1880 CSoutput.n128 gnd 0.789544f
C1881 CSoutput.n129 gnd 0.592158f
C1882 CSoutput.n130 gnd 0.789544f
C1883 CSoutput.n131 gnd 0.789544f
C1884 CSoutput.n132 gnd 2.1257f
C1885 CSoutput.n133 gnd 0.789544f
C1886 CSoutput.n134 gnd 0.789544f
C1887 CSoutput.t187 gnd 0.986931f
C1888 CSoutput.n135 gnd 0.789544f
C1889 CSoutput.n136 gnd 0.789544f
C1890 CSoutput.n140 gnd 0.789544f
C1891 CSoutput.n144 gnd 0.789544f
C1892 CSoutput.n145 gnd 0.789544f
C1893 CSoutput.n147 gnd 0.789544f
C1894 CSoutput.n152 gnd 0.789544f
C1895 CSoutput.n154 gnd 0.789544f
C1896 CSoutput.n155 gnd 0.789544f
C1897 CSoutput.n157 gnd 0.789544f
C1898 CSoutput.n158 gnd 0.789544f
C1899 CSoutput.n160 gnd 0.789544f
C1900 CSoutput.t181 gnd 13.1932f
C1901 CSoutput.n162 gnd 0.789544f
C1902 CSoutput.n163 gnd 0.592158f
C1903 CSoutput.n164 gnd 0.789544f
C1904 CSoutput.n165 gnd 0.789544f
C1905 CSoutput.n166 gnd 2.1257f
C1906 CSoutput.n167 gnd 0.789544f
C1907 CSoutput.n168 gnd 0.789544f
C1908 CSoutput.t184 gnd 0.986931f
C1909 CSoutput.n169 gnd 0.789544f
C1910 CSoutput.n170 gnd 0.789544f
C1911 CSoutput.n174 gnd 0.789544f
C1912 CSoutput.n178 gnd 0.789544f
C1913 CSoutput.n179 gnd 0.789544f
C1914 CSoutput.n181 gnd 0.789544f
C1915 CSoutput.n186 gnd 0.789544f
C1916 CSoutput.n188 gnd 0.789544f
C1917 CSoutput.n189 gnd 0.789544f
C1918 CSoutput.n191 gnd 0.789544f
C1919 CSoutput.n192 gnd 0.789544f
C1920 CSoutput.n194 gnd 0.789544f
C1921 CSoutput.n195 gnd 0.592158f
C1922 CSoutput.n197 gnd 0.789544f
C1923 CSoutput.n198 gnd 0.592158f
C1924 CSoutput.n199 gnd 0.789544f
C1925 CSoutput.n200 gnd 0.789544f
C1926 CSoutput.n201 gnd 2.1257f
C1927 CSoutput.n202 gnd 0.789544f
C1928 CSoutput.n203 gnd 0.789544f
C1929 CSoutput.t186 gnd 0.986931f
C1930 CSoutput.n204 gnd 0.789544f
C1931 CSoutput.n205 gnd 2.1257f
C1932 CSoutput.n207 gnd 0.789544f
C1933 CSoutput.n208 gnd 0.789544f
C1934 CSoutput.n210 gnd 0.789544f
C1935 CSoutput.n211 gnd 0.789544f
C1936 CSoutput.t192 gnd 12.9782f
C1937 CSoutput.t190 gnd 13.1932f
C1938 CSoutput.n217 gnd 2.47692f
C1939 CSoutput.n218 gnd 10.090099f
C1940 CSoutput.n219 gnd 10.5123f
C1941 CSoutput.n224 gnd 2.68317f
C1942 CSoutput.n230 gnd 0.789544f
C1943 CSoutput.n232 gnd 0.789544f
C1944 CSoutput.n234 gnd 0.789544f
C1945 CSoutput.n236 gnd 0.789544f
C1946 CSoutput.n238 gnd 0.789544f
C1947 CSoutput.n244 gnd 0.789544f
C1948 CSoutput.n251 gnd 1.44851f
C1949 CSoutput.n252 gnd 1.44851f
C1950 CSoutput.n253 gnd 0.789544f
C1951 CSoutput.n254 gnd 0.789544f
C1952 CSoutput.n256 gnd 0.592158f
C1953 CSoutput.n257 gnd 0.50713f
C1954 CSoutput.n259 gnd 0.592158f
C1955 CSoutput.n260 gnd 0.50713f
C1956 CSoutput.n261 gnd 0.592158f
C1957 CSoutput.n263 gnd 0.789544f
C1958 CSoutput.n265 gnd 2.1257f
C1959 CSoutput.n266 gnd 2.47692f
C1960 CSoutput.n267 gnd 9.28026f
C1961 CSoutput.n269 gnd 0.592158f
C1962 CSoutput.n270 gnd 1.52366f
C1963 CSoutput.n271 gnd 0.592158f
C1964 CSoutput.n273 gnd 0.789544f
C1965 CSoutput.n275 gnd 2.1257f
C1966 CSoutput.n276 gnd 4.63011f
C1967 CSoutput.t85 gnd 0.055673f
C1968 CSoutput.t138 gnd 0.055673f
C1969 CSoutput.n277 gnd 0.431039f
C1970 CSoutput.t102 gnd 0.055673f
C1971 CSoutput.t150 gnd 0.055673f
C1972 CSoutput.n278 gnd 0.43027f
C1973 CSoutput.n279 gnd 0.436724f
C1974 CSoutput.t133 gnd 0.055673f
C1975 CSoutput.t65 gnd 0.055673f
C1976 CSoutput.n280 gnd 0.43027f
C1977 CSoutput.n281 gnd 0.215199f
C1978 CSoutput.t93 gnd 0.055673f
C1979 CSoutput.t70 gnd 0.055673f
C1980 CSoutput.n282 gnd 0.43027f
C1981 CSoutput.n283 gnd 0.215199f
C1982 CSoutput.t109 gnd 0.055673f
C1983 CSoutput.t90 gnd 0.055673f
C1984 CSoutput.n284 gnd 0.43027f
C1985 CSoutput.n285 gnd 0.215199f
C1986 CSoutput.t142 gnd 0.055673f
C1987 CSoutput.t73 gnd 0.055673f
C1988 CSoutput.n286 gnd 0.43027f
C1989 CSoutput.n287 gnd 0.215199f
C1990 CSoutput.t124 gnd 0.055673f
C1991 CSoutput.t79 gnd 0.055673f
C1992 CSoutput.n288 gnd 0.43027f
C1993 CSoutput.n289 gnd 0.215199f
C1994 CSoutput.t134 gnd 0.055673f
C1995 CSoutput.t97 gnd 0.055673f
C1996 CSoutput.n290 gnd 0.43027f
C1997 CSoutput.n291 gnd 0.394625f
C1998 CSoutput.t108 gnd 0.055673f
C1999 CSoutput.t128 gnd 0.055673f
C2000 CSoutput.n292 gnd 0.431039f
C2001 CSoutput.t61 gnd 0.055673f
C2002 CSoutput.t91 gnd 0.055673f
C2003 CSoutput.n293 gnd 0.43027f
C2004 CSoutput.n294 gnd 0.436724f
C2005 CSoutput.t92 gnd 0.055673f
C2006 CSoutput.t146 gnd 0.055673f
C2007 CSoutput.n295 gnd 0.43027f
C2008 CSoutput.n296 gnd 0.215199f
C2009 CSoutput.t88 gnd 0.055673f
C2010 CSoutput.t89 gnd 0.055673f
C2011 CSoutput.n297 gnd 0.43027f
C2012 CSoutput.n298 gnd 0.215199f
C2013 CSoutput.t144 gnd 0.055673f
C2014 CSoutput.t145 gnd 0.055673f
C2015 CSoutput.n299 gnd 0.43027f
C2016 CSoutput.n300 gnd 0.215199f
C2017 CSoutput.t69 gnd 0.055673f
C2018 CSoutput.t129 gnd 0.055673f
C2019 CSoutput.n301 gnd 0.43027f
C2020 CSoutput.n302 gnd 0.215199f
C2021 CSoutput.t141 gnd 0.055673f
C2022 CSoutput.t68 gnd 0.055673f
C2023 CSoutput.n303 gnd 0.43027f
C2024 CSoutput.n304 gnd 0.215199f
C2025 CSoutput.t107 gnd 0.055673f
C2026 CSoutput.t127 gnd 0.055673f
C2027 CSoutput.n305 gnd 0.43027f
C2028 CSoutput.n306 gnd 0.320916f
C2029 CSoutput.n307 gnd 0.404673f
C2030 CSoutput.t117 gnd 0.055673f
C2031 CSoutput.t135 gnd 0.055673f
C2032 CSoutput.n308 gnd 0.431039f
C2033 CSoutput.t72 gnd 0.055673f
C2034 CSoutput.t104 gnd 0.055673f
C2035 CSoutput.n309 gnd 0.43027f
C2036 CSoutput.n310 gnd 0.436724f
C2037 CSoutput.t106 gnd 0.055673f
C2038 CSoutput.t154 gnd 0.055673f
C2039 CSoutput.n311 gnd 0.43027f
C2040 CSoutput.n312 gnd 0.215199f
C2041 CSoutput.t100 gnd 0.055673f
C2042 CSoutput.t101 gnd 0.055673f
C2043 CSoutput.n313 gnd 0.43027f
C2044 CSoutput.n314 gnd 0.215199f
C2045 CSoutput.t152 gnd 0.055673f
C2046 CSoutput.t153 gnd 0.055673f
C2047 CSoutput.n315 gnd 0.43027f
C2048 CSoutput.n316 gnd 0.215199f
C2049 CSoutput.t84 gnd 0.055673f
C2050 CSoutput.t140 gnd 0.055673f
C2051 CSoutput.n317 gnd 0.43027f
C2052 CSoutput.n318 gnd 0.215199f
C2053 CSoutput.t149 gnd 0.055673f
C2054 CSoutput.t80 gnd 0.055673f
C2055 CSoutput.n319 gnd 0.43027f
C2056 CSoutput.n320 gnd 0.215199f
C2057 CSoutput.t118 gnd 0.055673f
C2058 CSoutput.t136 gnd 0.055673f
C2059 CSoutput.n321 gnd 0.430269f
C2060 CSoutput.n322 gnd 0.320917f
C2061 CSoutput.n323 gnd 0.452321f
C2062 CSoutput.n324 gnd 12.9662f
C2063 CSoutput.t37 gnd 0.048714f
C2064 CSoutput.t59 gnd 0.048714f
C2065 CSoutput.n325 gnd 0.431894f
C2066 CSoutput.t13 gnd 0.048714f
C2067 CSoutput.t41 gnd 0.048714f
C2068 CSoutput.n326 gnd 0.430453f
C2069 CSoutput.n327 gnd 0.401102f
C2070 CSoutput.t22 gnd 0.048714f
C2071 CSoutput.t33 gnd 0.048714f
C2072 CSoutput.n328 gnd 0.430453f
C2073 CSoutput.n329 gnd 0.197724f
C2074 CSoutput.t11 gnd 0.048714f
C2075 CSoutput.t5 gnd 0.048714f
C2076 CSoutput.n330 gnd 0.430453f
C2077 CSoutput.n331 gnd 0.197724f
C2078 CSoutput.t60 gnd 0.048714f
C2079 CSoutput.t25 gnd 0.048714f
C2080 CSoutput.n332 gnd 0.430453f
C2081 CSoutput.n333 gnd 0.197724f
C2082 CSoutput.t29 gnd 0.048714f
C2083 CSoutput.t162 gnd 0.048714f
C2084 CSoutput.n334 gnd 0.430453f
C2085 CSoutput.n335 gnd 0.197724f
C2086 CSoutput.t165 gnd 0.048714f
C2087 CSoutput.t175 gnd 0.048714f
C2088 CSoutput.n336 gnd 0.430453f
C2089 CSoutput.n337 gnd 0.197724f
C2090 CSoutput.t53 gnd 0.048714f
C2091 CSoutput.t171 gnd 0.048714f
C2092 CSoutput.n338 gnd 0.430453f
C2093 CSoutput.n339 gnd 0.197724f
C2094 CSoutput.t18 gnd 0.048714f
C2095 CSoutput.t4 gnd 0.048714f
C2096 CSoutput.n340 gnd 0.430453f
C2097 CSoutput.n341 gnd 0.197724f
C2098 CSoutput.t12 gnd 0.048714f
C2099 CSoutput.t35 gnd 0.048714f
C2100 CSoutput.n342 gnd 0.430453f
C2101 CSoutput.n343 gnd 0.364644f
C2102 CSoutput.t1 gnd 0.048714f
C2103 CSoutput.t166 gnd 0.048714f
C2104 CSoutput.n344 gnd 0.431894f
C2105 CSoutput.t58 gnd 0.048714f
C2106 CSoutput.t56 gnd 0.048714f
C2107 CSoutput.n345 gnd 0.430453f
C2108 CSoutput.n346 gnd 0.401102f
C2109 CSoutput.t49 gnd 0.048714f
C2110 CSoutput.t21 gnd 0.048714f
C2111 CSoutput.n347 gnd 0.430453f
C2112 CSoutput.n348 gnd 0.197724f
C2113 CSoutput.t50 gnd 0.048714f
C2114 CSoutput.t173 gnd 0.048714f
C2115 CSoutput.n349 gnd 0.430453f
C2116 CSoutput.n350 gnd 0.197724f
C2117 CSoutput.t167 gnd 0.048714f
C2118 CSoutput.t169 gnd 0.048714f
C2119 CSoutput.n351 gnd 0.430453f
C2120 CSoutput.n352 gnd 0.197724f
C2121 CSoutput.t31 gnd 0.048714f
C2122 CSoutput.t8 gnd 0.048714f
C2123 CSoutput.n353 gnd 0.430453f
C2124 CSoutput.n354 gnd 0.197724f
C2125 CSoutput.t157 gnd 0.048714f
C2126 CSoutput.t161 gnd 0.048714f
C2127 CSoutput.n355 gnd 0.430453f
C2128 CSoutput.n356 gnd 0.197724f
C2129 CSoutput.t6 gnd 0.048714f
C2130 CSoutput.t57 gnd 0.048714f
C2131 CSoutput.n357 gnd 0.430453f
C2132 CSoutput.n358 gnd 0.197724f
C2133 CSoutput.t28 gnd 0.048714f
C2134 CSoutput.t17 gnd 0.048714f
C2135 CSoutput.n359 gnd 0.430453f
C2136 CSoutput.n360 gnd 0.197724f
C2137 CSoutput.t51 gnd 0.048714f
C2138 CSoutput.t2 gnd 0.048714f
C2139 CSoutput.n361 gnd 0.430453f
C2140 CSoutput.n362 gnd 0.300188f
C2141 CSoutput.n363 gnd 0.557772f
C2142 CSoutput.n364 gnd 13.858099f
C2143 CSoutput.t168 gnd 0.048714f
C2144 CSoutput.t48 gnd 0.048714f
C2145 CSoutput.n365 gnd 0.431894f
C2146 CSoutput.t20 gnd 0.048714f
C2147 CSoutput.t9 gnd 0.048714f
C2148 CSoutput.n366 gnd 0.430453f
C2149 CSoutput.n367 gnd 0.401102f
C2150 CSoutput.t23 gnd 0.048714f
C2151 CSoutput.t26 gnd 0.048714f
C2152 CSoutput.n368 gnd 0.430453f
C2153 CSoutput.n369 gnd 0.197724f
C2154 CSoutput.t52 gnd 0.048714f
C2155 CSoutput.t30 gnd 0.048714f
C2156 CSoutput.n370 gnd 0.430453f
C2157 CSoutput.n371 gnd 0.197724f
C2158 CSoutput.t10 gnd 0.048714f
C2159 CSoutput.t0 gnd 0.048714f
C2160 CSoutput.n372 gnd 0.430453f
C2161 CSoutput.n373 gnd 0.197724f
C2162 CSoutput.t14 gnd 0.048714f
C2163 CSoutput.t172 gnd 0.048714f
C2164 CSoutput.n374 gnd 0.430453f
C2165 CSoutput.n375 gnd 0.197724f
C2166 CSoutput.t32 gnd 0.048714f
C2167 CSoutput.t15 gnd 0.048714f
C2168 CSoutput.n376 gnd 0.430453f
C2169 CSoutput.n377 gnd 0.197724f
C2170 CSoutput.t38 gnd 0.048714f
C2171 CSoutput.t40 gnd 0.048714f
C2172 CSoutput.n378 gnd 0.430453f
C2173 CSoutput.n379 gnd 0.197724f
C2174 CSoutput.t19 gnd 0.048714f
C2175 CSoutput.t46 gnd 0.048714f
C2176 CSoutput.n380 gnd 0.430453f
C2177 CSoutput.n381 gnd 0.197724f
C2178 CSoutput.t163 gnd 0.048714f
C2179 CSoutput.t158 gnd 0.048714f
C2180 CSoutput.n382 gnd 0.430453f
C2181 CSoutput.n383 gnd 0.364644f
C2182 CSoutput.t34 gnd 0.048714f
C2183 CSoutput.t164 gnd 0.048714f
C2184 CSoutput.n384 gnd 0.431894f
C2185 CSoutput.t39 gnd 0.048714f
C2186 CSoutput.t174 gnd 0.048714f
C2187 CSoutput.n385 gnd 0.430453f
C2188 CSoutput.n386 gnd 0.401102f
C2189 CSoutput.t7 gnd 0.048714f
C2190 CSoutput.t45 gnd 0.048714f
C2191 CSoutput.n387 gnd 0.430453f
C2192 CSoutput.n388 gnd 0.197724f
C2193 CSoutput.t55 gnd 0.048714f
C2194 CSoutput.t24 gnd 0.048714f
C2195 CSoutput.n389 gnd 0.430453f
C2196 CSoutput.n390 gnd 0.197724f
C2197 CSoutput.t47 gnd 0.048714f
C2198 CSoutput.t43 gnd 0.048714f
C2199 CSoutput.n391 gnd 0.430453f
C2200 CSoutput.n392 gnd 0.197724f
C2201 CSoutput.t16 gnd 0.048714f
C2202 CSoutput.t3 gnd 0.048714f
C2203 CSoutput.n393 gnd 0.430453f
C2204 CSoutput.n394 gnd 0.197724f
C2205 CSoutput.t27 gnd 0.048714f
C2206 CSoutput.t44 gnd 0.048714f
C2207 CSoutput.n395 gnd 0.430453f
C2208 CSoutput.n396 gnd 0.197724f
C2209 CSoutput.t54 gnd 0.048714f
C2210 CSoutput.t160 gnd 0.048714f
C2211 CSoutput.n397 gnd 0.430453f
C2212 CSoutput.n398 gnd 0.197724f
C2213 CSoutput.t42 gnd 0.048714f
C2214 CSoutput.t36 gnd 0.048714f
C2215 CSoutput.n399 gnd 0.430453f
C2216 CSoutput.n400 gnd 0.197724f
C2217 CSoutput.t170 gnd 0.048714f
C2218 CSoutput.t159 gnd 0.048714f
C2219 CSoutput.n401 gnd 0.430453f
C2220 CSoutput.n402 gnd 0.300188f
C2221 CSoutput.n403 gnd 0.557772f
C2222 CSoutput.n404 gnd 8.42815f
C2223 CSoutput.n405 gnd 14.5494f
C2224 vdd.t257 gnd 0.037026f
C2225 vdd.t263 gnd 0.037026f
C2226 vdd.n0 gnd 0.292027f
C2227 vdd.t109 gnd 0.037026f
C2228 vdd.t251 gnd 0.037026f
C2229 vdd.n1 gnd 0.291545f
C2230 vdd.n2 gnd 0.26886f
C2231 vdd.t265 gnd 0.037026f
C2232 vdd.t244 gnd 0.037026f
C2233 vdd.n3 gnd 0.291545f
C2234 vdd.n4 gnd 0.135973f
C2235 vdd.t246 gnd 0.037026f
C2236 vdd.t259 gnd 0.037026f
C2237 vdd.n5 gnd 0.291545f
C2238 vdd.n6 gnd 0.127585f
C2239 vdd.t106 gnd 0.037026f
C2240 vdd.t267 gnd 0.037026f
C2241 vdd.n7 gnd 0.292027f
C2242 vdd.t261 gnd 0.037026f
C2243 vdd.t255 gnd 0.037026f
C2244 vdd.n8 gnd 0.291545f
C2245 vdd.n9 gnd 0.26886f
C2246 vdd.t253 gnd 0.037026f
C2247 vdd.t99 gnd 0.037026f
C2248 vdd.n10 gnd 0.291545f
C2249 vdd.n11 gnd 0.135973f
C2250 vdd.t102 gnd 0.037026f
C2251 vdd.t248 gnd 0.037026f
C2252 vdd.n12 gnd 0.291545f
C2253 vdd.n13 gnd 0.127585f
C2254 vdd.n14 gnd 0.0902f
C2255 vdd.t91 gnd 0.02057f
C2256 vdd.t4 gnd 0.02057f
C2257 vdd.n15 gnd 0.189336f
C2258 vdd.t9 gnd 0.02057f
C2259 vdd.t10 gnd 0.02057f
C2260 vdd.n16 gnd 0.188782f
C2261 vdd.n17 gnd 0.32854f
C2262 vdd.t8 gnd 0.02057f
C2263 vdd.t5 gnd 0.02057f
C2264 vdd.n18 gnd 0.188782f
C2265 vdd.n19 gnd 0.135921f
C2266 vdd.t2 gnd 0.02057f
C2267 vdd.t11 gnd 0.02057f
C2268 vdd.n20 gnd 0.189336f
C2269 vdd.t6 gnd 0.02057f
C2270 vdd.t242 gnd 0.02057f
C2271 vdd.n21 gnd 0.188782f
C2272 vdd.n22 gnd 0.32854f
C2273 vdd.t0 gnd 0.02057f
C2274 vdd.t1 gnd 0.02057f
C2275 vdd.n23 gnd 0.188782f
C2276 vdd.n24 gnd 0.135921f
C2277 vdd.t90 gnd 0.02057f
C2278 vdd.t241 gnd 0.02057f
C2279 vdd.n25 gnd 0.188782f
C2280 vdd.t3 gnd 0.02057f
C2281 vdd.t7 gnd 0.02057f
C2282 vdd.n26 gnd 0.188782f
C2283 vdd.n27 gnd 22.171501f
C2284 vdd.n28 gnd 8.47832f
C2285 vdd.n29 gnd 0.00561f
C2286 vdd.n30 gnd 0.005206f
C2287 vdd.n31 gnd 0.00288f
C2288 vdd.n32 gnd 0.006612f
C2289 vdd.n33 gnd 0.002797f
C2290 vdd.n34 gnd 0.002962f
C2291 vdd.n35 gnd 0.005206f
C2292 vdd.n36 gnd 0.002797f
C2293 vdd.n37 gnd 0.006612f
C2294 vdd.n38 gnd 0.002962f
C2295 vdd.n39 gnd 0.005206f
C2296 vdd.n40 gnd 0.002797f
C2297 vdd.n41 gnd 0.004959f
C2298 vdd.n42 gnd 0.004974f
C2299 vdd.t153 gnd 0.014206f
C2300 vdd.n43 gnd 0.031608f
C2301 vdd.n44 gnd 0.164495f
C2302 vdd.n45 gnd 0.002797f
C2303 vdd.n46 gnd 0.002962f
C2304 vdd.n47 gnd 0.006612f
C2305 vdd.n48 gnd 0.006612f
C2306 vdd.n49 gnd 0.002962f
C2307 vdd.n50 gnd 0.002797f
C2308 vdd.n51 gnd 0.005206f
C2309 vdd.n52 gnd 0.005206f
C2310 vdd.n53 gnd 0.002797f
C2311 vdd.n54 gnd 0.002962f
C2312 vdd.n55 gnd 0.006612f
C2313 vdd.n56 gnd 0.006612f
C2314 vdd.n57 gnd 0.002962f
C2315 vdd.n58 gnd 0.002797f
C2316 vdd.n59 gnd 0.005206f
C2317 vdd.n60 gnd 0.005206f
C2318 vdd.n61 gnd 0.002797f
C2319 vdd.n62 gnd 0.002962f
C2320 vdd.n63 gnd 0.006612f
C2321 vdd.n64 gnd 0.006612f
C2322 vdd.n65 gnd 0.015633f
C2323 vdd.n66 gnd 0.00288f
C2324 vdd.n67 gnd 0.002797f
C2325 vdd.n68 gnd 0.013456f
C2326 vdd.n69 gnd 0.009394f
C2327 vdd.t222 gnd 0.032912f
C2328 vdd.t177 gnd 0.032912f
C2329 vdd.n70 gnd 0.226192f
C2330 vdd.n71 gnd 0.177865f
C2331 vdd.t234 gnd 0.032912f
C2332 vdd.t217 gnd 0.032912f
C2333 vdd.n72 gnd 0.226192f
C2334 vdd.n73 gnd 0.143536f
C2335 vdd.t122 gnd 0.032912f
C2336 vdd.t168 gnd 0.032912f
C2337 vdd.n74 gnd 0.226192f
C2338 vdd.n75 gnd 0.143536f
C2339 vdd.t134 gnd 0.032912f
C2340 vdd.t187 gnd 0.032912f
C2341 vdd.n76 gnd 0.226192f
C2342 vdd.n77 gnd 0.143536f
C2343 vdd.t161 gnd 0.032912f
C2344 vdd.t223 gnd 0.032912f
C2345 vdd.n78 gnd 0.226192f
C2346 vdd.n79 gnd 0.143536f
C2347 vdd.t137 gnd 0.032912f
C2348 vdd.t206 gnd 0.032912f
C2349 vdd.n80 gnd 0.226192f
C2350 vdd.n81 gnd 0.143536f
C2351 vdd.t143 gnd 0.032912f
C2352 vdd.t218 gnd 0.032912f
C2353 vdd.n82 gnd 0.226192f
C2354 vdd.n83 gnd 0.143536f
C2355 vdd.n84 gnd 0.00561f
C2356 vdd.n85 gnd 0.005206f
C2357 vdd.n86 gnd 0.00288f
C2358 vdd.n87 gnd 0.006612f
C2359 vdd.n88 gnd 0.002797f
C2360 vdd.n89 gnd 0.002962f
C2361 vdd.n90 gnd 0.005206f
C2362 vdd.n91 gnd 0.002797f
C2363 vdd.n92 gnd 0.006612f
C2364 vdd.n93 gnd 0.002962f
C2365 vdd.n94 gnd 0.005206f
C2366 vdd.n95 gnd 0.002797f
C2367 vdd.n96 gnd 0.004959f
C2368 vdd.n97 gnd 0.004974f
C2369 vdd.t172 gnd 0.014206f
C2370 vdd.n98 gnd 0.031608f
C2371 vdd.n99 gnd 0.164495f
C2372 vdd.n100 gnd 0.002797f
C2373 vdd.n101 gnd 0.002962f
C2374 vdd.n102 gnd 0.006612f
C2375 vdd.n103 gnd 0.006612f
C2376 vdd.n104 gnd 0.002962f
C2377 vdd.n105 gnd 0.002797f
C2378 vdd.n106 gnd 0.005206f
C2379 vdd.n107 gnd 0.005206f
C2380 vdd.n108 gnd 0.002797f
C2381 vdd.n109 gnd 0.002962f
C2382 vdd.n110 gnd 0.006612f
C2383 vdd.n111 gnd 0.006612f
C2384 vdd.n112 gnd 0.002962f
C2385 vdd.n113 gnd 0.002797f
C2386 vdd.n114 gnd 0.005206f
C2387 vdd.n115 gnd 0.005206f
C2388 vdd.n116 gnd 0.002797f
C2389 vdd.n117 gnd 0.002962f
C2390 vdd.n118 gnd 0.006612f
C2391 vdd.n119 gnd 0.006612f
C2392 vdd.n120 gnd 0.015633f
C2393 vdd.n121 gnd 0.00288f
C2394 vdd.n122 gnd 0.002797f
C2395 vdd.n123 gnd 0.013456f
C2396 vdd.n124 gnd 0.0091f
C2397 vdd.n125 gnd 0.106792f
C2398 vdd.n126 gnd 0.00561f
C2399 vdd.n127 gnd 0.005206f
C2400 vdd.n128 gnd 0.00288f
C2401 vdd.n129 gnd 0.006612f
C2402 vdd.n130 gnd 0.002797f
C2403 vdd.n131 gnd 0.002962f
C2404 vdd.n132 gnd 0.005206f
C2405 vdd.n133 gnd 0.002797f
C2406 vdd.n134 gnd 0.006612f
C2407 vdd.n135 gnd 0.002962f
C2408 vdd.n136 gnd 0.005206f
C2409 vdd.n137 gnd 0.002797f
C2410 vdd.n138 gnd 0.004959f
C2411 vdd.n139 gnd 0.004974f
C2412 vdd.t185 gnd 0.014206f
C2413 vdd.n140 gnd 0.031608f
C2414 vdd.n141 gnd 0.164495f
C2415 vdd.n142 gnd 0.002797f
C2416 vdd.n143 gnd 0.002962f
C2417 vdd.n144 gnd 0.006612f
C2418 vdd.n145 gnd 0.006612f
C2419 vdd.n146 gnd 0.002962f
C2420 vdd.n147 gnd 0.002797f
C2421 vdd.n148 gnd 0.005206f
C2422 vdd.n149 gnd 0.005206f
C2423 vdd.n150 gnd 0.002797f
C2424 vdd.n151 gnd 0.002962f
C2425 vdd.n152 gnd 0.006612f
C2426 vdd.n153 gnd 0.006612f
C2427 vdd.n154 gnd 0.002962f
C2428 vdd.n155 gnd 0.002797f
C2429 vdd.n156 gnd 0.005206f
C2430 vdd.n157 gnd 0.005206f
C2431 vdd.n158 gnd 0.002797f
C2432 vdd.n159 gnd 0.002962f
C2433 vdd.n160 gnd 0.006612f
C2434 vdd.n161 gnd 0.006612f
C2435 vdd.n162 gnd 0.015633f
C2436 vdd.n163 gnd 0.00288f
C2437 vdd.n164 gnd 0.002797f
C2438 vdd.n165 gnd 0.013456f
C2439 vdd.n166 gnd 0.009394f
C2440 vdd.t212 gnd 0.032912f
C2441 vdd.t114 gnd 0.032912f
C2442 vdd.n167 gnd 0.226192f
C2443 vdd.n168 gnd 0.177865f
C2444 vdd.t163 gnd 0.032912f
C2445 vdd.t165 gnd 0.032912f
C2446 vdd.n169 gnd 0.226192f
C2447 vdd.n170 gnd 0.143536f
C2448 vdd.t230 gnd 0.032912f
C2449 vdd.t158 gnd 0.032912f
C2450 vdd.n171 gnd 0.226192f
C2451 vdd.n172 gnd 0.143536f
C2452 vdd.t159 gnd 0.032912f
C2453 vdd.t229 gnd 0.032912f
C2454 vdd.n173 gnd 0.226192f
C2455 vdd.n174 gnd 0.143536f
C2456 vdd.t224 gnd 0.032912f
C2457 vdd.t130 gnd 0.032912f
C2458 vdd.n175 gnd 0.226192f
C2459 vdd.n176 gnd 0.143536f
C2460 vdd.t213 gnd 0.032912f
C2461 vdd.t227 gnd 0.032912f
C2462 vdd.n177 gnd 0.226192f
C2463 vdd.n178 gnd 0.143536f
C2464 vdd.t128 gnd 0.032912f
C2465 vdd.t182 gnd 0.032912f
C2466 vdd.n179 gnd 0.226192f
C2467 vdd.n180 gnd 0.143536f
C2468 vdd.n181 gnd 0.00561f
C2469 vdd.n182 gnd 0.005206f
C2470 vdd.n183 gnd 0.00288f
C2471 vdd.n184 gnd 0.006612f
C2472 vdd.n185 gnd 0.002797f
C2473 vdd.n186 gnd 0.002962f
C2474 vdd.n187 gnd 0.005206f
C2475 vdd.n188 gnd 0.002797f
C2476 vdd.n189 gnd 0.006612f
C2477 vdd.n190 gnd 0.002962f
C2478 vdd.n191 gnd 0.005206f
C2479 vdd.n192 gnd 0.002797f
C2480 vdd.n193 gnd 0.004959f
C2481 vdd.n194 gnd 0.004974f
C2482 vdd.t210 gnd 0.014206f
C2483 vdd.n195 gnd 0.031608f
C2484 vdd.n196 gnd 0.164495f
C2485 vdd.n197 gnd 0.002797f
C2486 vdd.n198 gnd 0.002962f
C2487 vdd.n199 gnd 0.006612f
C2488 vdd.n200 gnd 0.006612f
C2489 vdd.n201 gnd 0.002962f
C2490 vdd.n202 gnd 0.002797f
C2491 vdd.n203 gnd 0.005206f
C2492 vdd.n204 gnd 0.005206f
C2493 vdd.n205 gnd 0.002797f
C2494 vdd.n206 gnd 0.002962f
C2495 vdd.n207 gnd 0.006612f
C2496 vdd.n208 gnd 0.006612f
C2497 vdd.n209 gnd 0.002962f
C2498 vdd.n210 gnd 0.002797f
C2499 vdd.n211 gnd 0.005206f
C2500 vdd.n212 gnd 0.005206f
C2501 vdd.n213 gnd 0.002797f
C2502 vdd.n214 gnd 0.002962f
C2503 vdd.n215 gnd 0.006612f
C2504 vdd.n216 gnd 0.006612f
C2505 vdd.n217 gnd 0.015633f
C2506 vdd.n218 gnd 0.00288f
C2507 vdd.n219 gnd 0.002797f
C2508 vdd.n220 gnd 0.013456f
C2509 vdd.n221 gnd 0.0091f
C2510 vdd.n222 gnd 0.06353f
C2511 vdd.n223 gnd 0.228916f
C2512 vdd.n224 gnd 0.00561f
C2513 vdd.n225 gnd 0.005206f
C2514 vdd.n226 gnd 0.00288f
C2515 vdd.n227 gnd 0.006612f
C2516 vdd.n228 gnd 0.002797f
C2517 vdd.n229 gnd 0.002962f
C2518 vdd.n230 gnd 0.005206f
C2519 vdd.n231 gnd 0.002797f
C2520 vdd.n232 gnd 0.006612f
C2521 vdd.n233 gnd 0.002962f
C2522 vdd.n234 gnd 0.005206f
C2523 vdd.n235 gnd 0.002797f
C2524 vdd.n236 gnd 0.004959f
C2525 vdd.n237 gnd 0.004974f
C2526 vdd.t198 gnd 0.014206f
C2527 vdd.n238 gnd 0.031608f
C2528 vdd.n239 gnd 0.164495f
C2529 vdd.n240 gnd 0.002797f
C2530 vdd.n241 gnd 0.002962f
C2531 vdd.n242 gnd 0.006612f
C2532 vdd.n243 gnd 0.006612f
C2533 vdd.n244 gnd 0.002962f
C2534 vdd.n245 gnd 0.002797f
C2535 vdd.n246 gnd 0.005206f
C2536 vdd.n247 gnd 0.005206f
C2537 vdd.n248 gnd 0.002797f
C2538 vdd.n249 gnd 0.002962f
C2539 vdd.n250 gnd 0.006612f
C2540 vdd.n251 gnd 0.006612f
C2541 vdd.n252 gnd 0.002962f
C2542 vdd.n253 gnd 0.002797f
C2543 vdd.n254 gnd 0.005206f
C2544 vdd.n255 gnd 0.005206f
C2545 vdd.n256 gnd 0.002797f
C2546 vdd.n257 gnd 0.002962f
C2547 vdd.n258 gnd 0.006612f
C2548 vdd.n259 gnd 0.006612f
C2549 vdd.n260 gnd 0.015633f
C2550 vdd.n261 gnd 0.00288f
C2551 vdd.n262 gnd 0.002797f
C2552 vdd.n263 gnd 0.013456f
C2553 vdd.n264 gnd 0.009394f
C2554 vdd.t219 gnd 0.032912f
C2555 vdd.t135 gnd 0.032912f
C2556 vdd.n265 gnd 0.226192f
C2557 vdd.n266 gnd 0.177865f
C2558 vdd.t180 gnd 0.032912f
C2559 vdd.t184 gnd 0.032912f
C2560 vdd.n267 gnd 0.226192f
C2561 vdd.n268 gnd 0.143536f
C2562 vdd.t238 gnd 0.032912f
C2563 vdd.t175 gnd 0.032912f
C2564 vdd.n269 gnd 0.226192f
C2565 vdd.n270 gnd 0.143536f
C2566 vdd.t176 gnd 0.032912f
C2567 vdd.t236 gnd 0.032912f
C2568 vdd.n271 gnd 0.226192f
C2569 vdd.n272 gnd 0.143536f
C2570 vdd.t237 gnd 0.032912f
C2571 vdd.t151 gnd 0.032912f
C2572 vdd.n273 gnd 0.226192f
C2573 vdd.n274 gnd 0.143536f
C2574 vdd.t226 gnd 0.032912f
C2575 vdd.t233 gnd 0.032912f
C2576 vdd.n275 gnd 0.226192f
C2577 vdd.n276 gnd 0.143536f
C2578 vdd.t146 gnd 0.032912f
C2579 vdd.t199 gnd 0.032912f
C2580 vdd.n277 gnd 0.226192f
C2581 vdd.n278 gnd 0.143536f
C2582 vdd.n279 gnd 0.00561f
C2583 vdd.n280 gnd 0.005206f
C2584 vdd.n281 gnd 0.00288f
C2585 vdd.n282 gnd 0.006612f
C2586 vdd.n283 gnd 0.002797f
C2587 vdd.n284 gnd 0.002962f
C2588 vdd.n285 gnd 0.005206f
C2589 vdd.n286 gnd 0.002797f
C2590 vdd.n287 gnd 0.006612f
C2591 vdd.n288 gnd 0.002962f
C2592 vdd.n289 gnd 0.005206f
C2593 vdd.n290 gnd 0.002797f
C2594 vdd.n291 gnd 0.004959f
C2595 vdd.n292 gnd 0.004974f
C2596 vdd.t220 gnd 0.014206f
C2597 vdd.n293 gnd 0.031608f
C2598 vdd.n294 gnd 0.164495f
C2599 vdd.n295 gnd 0.002797f
C2600 vdd.n296 gnd 0.002962f
C2601 vdd.n297 gnd 0.006612f
C2602 vdd.n298 gnd 0.006612f
C2603 vdd.n299 gnd 0.002962f
C2604 vdd.n300 gnd 0.002797f
C2605 vdd.n301 gnd 0.005206f
C2606 vdd.n302 gnd 0.005206f
C2607 vdd.n303 gnd 0.002797f
C2608 vdd.n304 gnd 0.002962f
C2609 vdd.n305 gnd 0.006612f
C2610 vdd.n306 gnd 0.006612f
C2611 vdd.n307 gnd 0.002962f
C2612 vdd.n308 gnd 0.002797f
C2613 vdd.n309 gnd 0.005206f
C2614 vdd.n310 gnd 0.005206f
C2615 vdd.n311 gnd 0.002797f
C2616 vdd.n312 gnd 0.002962f
C2617 vdd.n313 gnd 0.006612f
C2618 vdd.n314 gnd 0.006612f
C2619 vdd.n315 gnd 0.015633f
C2620 vdd.n316 gnd 0.00288f
C2621 vdd.n317 gnd 0.002797f
C2622 vdd.n318 gnd 0.013456f
C2623 vdd.n319 gnd 0.0091f
C2624 vdd.n320 gnd 0.06353f
C2625 vdd.n321 gnd 0.256355f
C2626 vdd.n322 gnd 0.007857f
C2627 vdd.n323 gnd 0.010223f
C2628 vdd.n324 gnd 0.008228f
C2629 vdd.n325 gnd 0.008228f
C2630 vdd.n326 gnd 0.010223f
C2631 vdd.n327 gnd 0.010223f
C2632 vdd.n328 gnd 0.746958f
C2633 vdd.n329 gnd 0.010223f
C2634 vdd.n330 gnd 0.010223f
C2635 vdd.n331 gnd 0.010223f
C2636 vdd.n332 gnd 0.809639f
C2637 vdd.n333 gnd 0.010223f
C2638 vdd.n334 gnd 0.010223f
C2639 vdd.n335 gnd 0.010223f
C2640 vdd.n336 gnd 0.010223f
C2641 vdd.n337 gnd 0.008228f
C2642 vdd.n338 gnd 0.010223f
C2643 vdd.t129 gnd 0.522348f
C2644 vdd.n339 gnd 0.010223f
C2645 vdd.n340 gnd 0.010223f
C2646 vdd.n341 gnd 0.010223f
C2647 vdd.t205 gnd 0.522348f
C2648 vdd.n342 gnd 0.010223f
C2649 vdd.n343 gnd 0.010223f
C2650 vdd.n344 gnd 0.010223f
C2651 vdd.n345 gnd 0.010223f
C2652 vdd.n346 gnd 0.010223f
C2653 vdd.n347 gnd 0.008228f
C2654 vdd.n348 gnd 0.010223f
C2655 vdd.n349 gnd 0.590253f
C2656 vdd.n350 gnd 0.010223f
C2657 vdd.n351 gnd 0.010223f
C2658 vdd.n352 gnd 0.010223f
C2659 vdd.t181 gnd 0.522348f
C2660 vdd.n353 gnd 0.010223f
C2661 vdd.n354 gnd 0.010223f
C2662 vdd.n355 gnd 0.010223f
C2663 vdd.n356 gnd 0.010223f
C2664 vdd.n357 gnd 0.010223f
C2665 vdd.n358 gnd 0.008228f
C2666 vdd.n359 gnd 0.010223f
C2667 vdd.t171 gnd 0.522348f
C2668 vdd.n360 gnd 0.010223f
C2669 vdd.n361 gnd 0.010223f
C2670 vdd.n362 gnd 0.010223f
C2671 vdd.n363 gnd 0.882768f
C2672 vdd.n364 gnd 0.010223f
C2673 vdd.n365 gnd 0.010223f
C2674 vdd.n366 gnd 0.010223f
C2675 vdd.n367 gnd 0.010223f
C2676 vdd.n368 gnd 0.010223f
C2677 vdd.n369 gnd 0.006829f
C2678 vdd.n370 gnd 0.023279f
C2679 vdd.t46 gnd 0.522348f
C2680 vdd.n371 gnd 0.010223f
C2681 vdd.n372 gnd 0.023279f
C2682 vdd.n404 gnd 0.010223f
C2683 vdd.t48 gnd 0.125764f
C2684 vdd.t47 gnd 0.134407f
C2685 vdd.t45 gnd 0.164246f
C2686 vdd.n405 gnd 0.210541f
C2687 vdd.n406 gnd 0.177715f
C2688 vdd.n407 gnd 0.013494f
C2689 vdd.n408 gnd 0.010223f
C2690 vdd.n409 gnd 0.008228f
C2691 vdd.n410 gnd 0.010223f
C2692 vdd.n411 gnd 0.008228f
C2693 vdd.n412 gnd 0.010223f
C2694 vdd.n413 gnd 0.008228f
C2695 vdd.n414 gnd 0.010223f
C2696 vdd.n415 gnd 0.008228f
C2697 vdd.n416 gnd 0.010223f
C2698 vdd.n417 gnd 0.008228f
C2699 vdd.n418 gnd 0.010223f
C2700 vdd.t81 gnd 0.125764f
C2701 vdd.t80 gnd 0.134407f
C2702 vdd.t79 gnd 0.164246f
C2703 vdd.n419 gnd 0.210541f
C2704 vdd.n420 gnd 0.177715f
C2705 vdd.n421 gnd 0.008228f
C2706 vdd.n422 gnd 0.010223f
C2707 vdd.n423 gnd 0.008228f
C2708 vdd.n424 gnd 0.010223f
C2709 vdd.n425 gnd 0.008228f
C2710 vdd.n426 gnd 0.010223f
C2711 vdd.n427 gnd 0.008228f
C2712 vdd.n428 gnd 0.010223f
C2713 vdd.n429 gnd 0.008228f
C2714 vdd.n430 gnd 0.010223f
C2715 vdd.t87 gnd 0.125764f
C2716 vdd.t86 gnd 0.134407f
C2717 vdd.t85 gnd 0.164246f
C2718 vdd.n431 gnd 0.210541f
C2719 vdd.n432 gnd 0.177715f
C2720 vdd.n433 gnd 0.017608f
C2721 vdd.n434 gnd 0.010223f
C2722 vdd.n435 gnd 0.008228f
C2723 vdd.n436 gnd 0.010223f
C2724 vdd.n437 gnd 0.008228f
C2725 vdd.n438 gnd 0.010223f
C2726 vdd.n439 gnd 0.008228f
C2727 vdd.n440 gnd 0.010223f
C2728 vdd.n441 gnd 0.008228f
C2729 vdd.n442 gnd 0.010223f
C2730 vdd.n443 gnd 0.023279f
C2731 vdd.n444 gnd 0.023438f
C2732 vdd.n445 gnd 0.023438f
C2733 vdd.n446 gnd 0.006829f
C2734 vdd.n447 gnd 0.008228f
C2735 vdd.n448 gnd 0.010223f
C2736 vdd.n449 gnd 0.010223f
C2737 vdd.n450 gnd 0.008228f
C2738 vdd.n451 gnd 0.010223f
C2739 vdd.n452 gnd 0.010223f
C2740 vdd.n453 gnd 0.010223f
C2741 vdd.n454 gnd 0.010223f
C2742 vdd.n455 gnd 0.010223f
C2743 vdd.n456 gnd 0.008228f
C2744 vdd.n457 gnd 0.008228f
C2745 vdd.n458 gnd 0.010223f
C2746 vdd.n459 gnd 0.010223f
C2747 vdd.n460 gnd 0.008228f
C2748 vdd.n461 gnd 0.010223f
C2749 vdd.n462 gnd 0.010223f
C2750 vdd.n463 gnd 0.010223f
C2751 vdd.n464 gnd 0.010223f
C2752 vdd.n465 gnd 0.010223f
C2753 vdd.n466 gnd 0.008228f
C2754 vdd.n467 gnd 0.008228f
C2755 vdd.n468 gnd 0.010223f
C2756 vdd.n469 gnd 0.010223f
C2757 vdd.n470 gnd 0.008228f
C2758 vdd.n471 gnd 0.010223f
C2759 vdd.n472 gnd 0.010223f
C2760 vdd.n473 gnd 0.010223f
C2761 vdd.n474 gnd 0.010223f
C2762 vdd.n475 gnd 0.010223f
C2763 vdd.n476 gnd 0.008228f
C2764 vdd.n477 gnd 0.008228f
C2765 vdd.n478 gnd 0.010223f
C2766 vdd.n479 gnd 0.010223f
C2767 vdd.n480 gnd 0.008228f
C2768 vdd.n481 gnd 0.010223f
C2769 vdd.n482 gnd 0.010223f
C2770 vdd.n483 gnd 0.010223f
C2771 vdd.n484 gnd 0.010223f
C2772 vdd.n485 gnd 0.010223f
C2773 vdd.n486 gnd 0.008228f
C2774 vdd.n487 gnd 0.008228f
C2775 vdd.n488 gnd 0.010223f
C2776 vdd.n489 gnd 0.010223f
C2777 vdd.n490 gnd 0.00687f
C2778 vdd.n491 gnd 0.010223f
C2779 vdd.n492 gnd 0.010223f
C2780 vdd.n493 gnd 0.010223f
C2781 vdd.n494 gnd 0.010223f
C2782 vdd.n495 gnd 0.010223f
C2783 vdd.n496 gnd 0.00687f
C2784 vdd.n497 gnd 0.008228f
C2785 vdd.n498 gnd 0.010223f
C2786 vdd.n499 gnd 0.010223f
C2787 vdd.n500 gnd 0.008228f
C2788 vdd.n501 gnd 0.010223f
C2789 vdd.n502 gnd 0.010223f
C2790 vdd.n503 gnd 0.010223f
C2791 vdd.n504 gnd 0.010223f
C2792 vdd.n505 gnd 0.010223f
C2793 vdd.n506 gnd 0.008228f
C2794 vdd.n507 gnd 0.008228f
C2795 vdd.n508 gnd 0.010223f
C2796 vdd.n509 gnd 0.010223f
C2797 vdd.n510 gnd 0.008228f
C2798 vdd.n511 gnd 0.010223f
C2799 vdd.n512 gnd 0.010223f
C2800 vdd.n513 gnd 0.010223f
C2801 vdd.n514 gnd 0.010223f
C2802 vdd.n515 gnd 0.010223f
C2803 vdd.n516 gnd 0.008228f
C2804 vdd.n517 gnd 0.008228f
C2805 vdd.n518 gnd 0.010223f
C2806 vdd.n519 gnd 0.010223f
C2807 vdd.n520 gnd 0.008228f
C2808 vdd.n521 gnd 0.010223f
C2809 vdd.n522 gnd 0.010223f
C2810 vdd.n523 gnd 0.010223f
C2811 vdd.n524 gnd 0.010223f
C2812 vdd.n525 gnd 0.010223f
C2813 vdd.n526 gnd 0.008228f
C2814 vdd.n527 gnd 0.008228f
C2815 vdd.n528 gnd 0.010223f
C2816 vdd.n529 gnd 0.010223f
C2817 vdd.n530 gnd 0.008228f
C2818 vdd.n531 gnd 0.010223f
C2819 vdd.n532 gnd 0.010223f
C2820 vdd.n533 gnd 0.010223f
C2821 vdd.n534 gnd 0.010223f
C2822 vdd.n535 gnd 0.010223f
C2823 vdd.n536 gnd 0.008228f
C2824 vdd.n537 gnd 0.008228f
C2825 vdd.n538 gnd 0.010223f
C2826 vdd.n539 gnd 0.010223f
C2827 vdd.n540 gnd 0.008228f
C2828 vdd.n541 gnd 0.010223f
C2829 vdd.n542 gnd 0.010223f
C2830 vdd.n543 gnd 0.010223f
C2831 vdd.n544 gnd 0.010223f
C2832 vdd.n545 gnd 0.010223f
C2833 vdd.n546 gnd 0.005595f
C2834 vdd.n547 gnd 0.017608f
C2835 vdd.n548 gnd 0.010223f
C2836 vdd.n549 gnd 0.010223f
C2837 vdd.n550 gnd 0.008146f
C2838 vdd.n551 gnd 0.010223f
C2839 vdd.n552 gnd 0.010223f
C2840 vdd.n553 gnd 0.010223f
C2841 vdd.n554 gnd 0.010223f
C2842 vdd.n555 gnd 0.010223f
C2843 vdd.n556 gnd 0.008228f
C2844 vdd.n557 gnd 0.008228f
C2845 vdd.n558 gnd 0.010223f
C2846 vdd.n559 gnd 0.010223f
C2847 vdd.n560 gnd 0.008228f
C2848 vdd.n561 gnd 0.010223f
C2849 vdd.n562 gnd 0.010223f
C2850 vdd.n563 gnd 0.010223f
C2851 vdd.n564 gnd 0.010223f
C2852 vdd.n565 gnd 0.010223f
C2853 vdd.n566 gnd 0.008228f
C2854 vdd.n567 gnd 0.008228f
C2855 vdd.n568 gnd 0.010223f
C2856 vdd.n569 gnd 0.010223f
C2857 vdd.n570 gnd 0.008228f
C2858 vdd.n571 gnd 0.010223f
C2859 vdd.n572 gnd 0.010223f
C2860 vdd.n573 gnd 0.010223f
C2861 vdd.n574 gnd 0.010223f
C2862 vdd.n575 gnd 0.010223f
C2863 vdd.n576 gnd 0.008228f
C2864 vdd.n577 gnd 0.008228f
C2865 vdd.n578 gnd 0.010223f
C2866 vdd.n579 gnd 0.010223f
C2867 vdd.n580 gnd 0.008228f
C2868 vdd.n581 gnd 0.010223f
C2869 vdd.n582 gnd 0.010223f
C2870 vdd.n583 gnd 0.010223f
C2871 vdd.n584 gnd 0.010223f
C2872 vdd.n585 gnd 0.010223f
C2873 vdd.n586 gnd 0.008228f
C2874 vdd.n587 gnd 0.008228f
C2875 vdd.n588 gnd 0.010223f
C2876 vdd.n589 gnd 0.010223f
C2877 vdd.n590 gnd 0.008228f
C2878 vdd.n591 gnd 0.010223f
C2879 vdd.n592 gnd 0.010223f
C2880 vdd.n593 gnd 0.010223f
C2881 vdd.n594 gnd 0.010223f
C2882 vdd.n595 gnd 0.010223f
C2883 vdd.n596 gnd 0.008228f
C2884 vdd.n597 gnd 0.010223f
C2885 vdd.n598 gnd 0.008228f
C2886 vdd.n599 gnd 0.00432f
C2887 vdd.n600 gnd 0.010223f
C2888 vdd.n601 gnd 0.010223f
C2889 vdd.n602 gnd 0.008228f
C2890 vdd.n603 gnd 0.010223f
C2891 vdd.n604 gnd 0.008228f
C2892 vdd.n605 gnd 0.010223f
C2893 vdd.n606 gnd 0.008228f
C2894 vdd.n607 gnd 0.010223f
C2895 vdd.n608 gnd 0.008228f
C2896 vdd.n609 gnd 0.010223f
C2897 vdd.n610 gnd 0.008228f
C2898 vdd.n611 gnd 0.010223f
C2899 vdd.n612 gnd 0.010223f
C2900 vdd.n613 gnd 0.569359f
C2901 vdd.t133 gnd 0.522348f
C2902 vdd.n614 gnd 0.010223f
C2903 vdd.n615 gnd 0.008228f
C2904 vdd.n616 gnd 0.010223f
C2905 vdd.n617 gnd 0.008228f
C2906 vdd.n618 gnd 0.010223f
C2907 vdd.t121 gnd 0.522348f
C2908 vdd.n619 gnd 0.010223f
C2909 vdd.n620 gnd 0.008228f
C2910 vdd.n621 gnd 0.010223f
C2911 vdd.n622 gnd 0.008228f
C2912 vdd.n623 gnd 0.010223f
C2913 vdd.t164 gnd 0.522348f
C2914 vdd.n624 gnd 0.652935f
C2915 vdd.n625 gnd 0.010223f
C2916 vdd.n626 gnd 0.008228f
C2917 vdd.n627 gnd 0.010223f
C2918 vdd.n628 gnd 0.008228f
C2919 vdd.n629 gnd 0.010223f
C2920 vdd.t162 gnd 0.522348f
C2921 vdd.n630 gnd 0.010223f
C2922 vdd.n631 gnd 0.008228f
C2923 vdd.n632 gnd 0.010223f
C2924 vdd.n633 gnd 0.008228f
C2925 vdd.n634 gnd 0.010223f
C2926 vdd.n635 gnd 0.726064f
C2927 vdd.n636 gnd 0.867098f
C2928 vdd.t113 gnd 0.522348f
C2929 vdd.n637 gnd 0.010223f
C2930 vdd.n638 gnd 0.008228f
C2931 vdd.n639 gnd 0.010223f
C2932 vdd.n640 gnd 0.008228f
C2933 vdd.n641 gnd 0.010223f
C2934 vdd.n642 gnd 0.548465f
C2935 vdd.n643 gnd 0.010223f
C2936 vdd.n644 gnd 0.008228f
C2937 vdd.n645 gnd 0.010223f
C2938 vdd.n646 gnd 0.008228f
C2939 vdd.n647 gnd 0.010223f
C2940 vdd.n648 gnd 1.0447f
C2941 vdd.t152 gnd 0.522348f
C2942 vdd.n649 gnd 0.010223f
C2943 vdd.n650 gnd 0.008228f
C2944 vdd.n651 gnd 0.010223f
C2945 vdd.n652 gnd 0.008228f
C2946 vdd.n653 gnd 0.010223f
C2947 vdd.t21 gnd 0.522348f
C2948 vdd.n654 gnd 0.010223f
C2949 vdd.n655 gnd 0.008228f
C2950 vdd.n656 gnd 0.023438f
C2951 vdd.n657 gnd 0.023438f
C2952 vdd.n658 gnd 9.1202f
C2953 vdd.n659 gnd 0.579806f
C2954 vdd.n660 gnd 0.023438f
C2955 vdd.n661 gnd 0.008791f
C2956 vdd.n662 gnd 0.008228f
C2957 vdd.n667 gnd 0.006542f
C2958 vdd.n668 gnd 0.008228f
C2959 vdd.n669 gnd 0.010223f
C2960 vdd.n670 gnd 0.010223f
C2961 vdd.n671 gnd 0.010223f
C2962 vdd.n672 gnd 0.010223f
C2963 vdd.n673 gnd 0.010223f
C2964 vdd.n674 gnd 0.008228f
C2965 vdd.n675 gnd 0.010223f
C2966 vdd.n676 gnd 0.010223f
C2967 vdd.n677 gnd 0.010223f
C2968 vdd.n678 gnd 0.010223f
C2969 vdd.n679 gnd 0.010223f
C2970 vdd.n680 gnd 0.008228f
C2971 vdd.n681 gnd 0.010223f
C2972 vdd.n682 gnd 0.010223f
C2973 vdd.n683 gnd 0.010223f
C2974 vdd.n684 gnd 0.010223f
C2975 vdd.n685 gnd 0.010223f
C2976 vdd.t39 gnd 0.125764f
C2977 vdd.t40 gnd 0.134407f
C2978 vdd.t38 gnd 0.164246f
C2979 vdd.n686 gnd 0.210541f
C2980 vdd.n687 gnd 0.176892f
C2981 vdd.n688 gnd 0.016785f
C2982 vdd.n689 gnd 0.010223f
C2983 vdd.n690 gnd 0.010223f
C2984 vdd.n691 gnd 0.010223f
C2985 vdd.n692 gnd 0.010223f
C2986 vdd.n693 gnd 0.010223f
C2987 vdd.n694 gnd 0.008228f
C2988 vdd.n695 gnd 0.010223f
C2989 vdd.n696 gnd 0.010223f
C2990 vdd.n697 gnd 0.010223f
C2991 vdd.n698 gnd 0.010223f
C2992 vdd.n699 gnd 0.010223f
C2993 vdd.n700 gnd 0.008228f
C2994 vdd.n701 gnd 0.010223f
C2995 vdd.n702 gnd 0.010223f
C2996 vdd.n703 gnd 0.010223f
C2997 vdd.n704 gnd 0.010223f
C2998 vdd.n705 gnd 0.010223f
C2999 vdd.n706 gnd 0.008228f
C3000 vdd.n707 gnd 0.010223f
C3001 vdd.n708 gnd 0.010223f
C3002 vdd.n709 gnd 0.010223f
C3003 vdd.n710 gnd 0.010223f
C3004 vdd.n711 gnd 0.010223f
C3005 vdd.n712 gnd 0.008228f
C3006 vdd.n713 gnd 0.010223f
C3007 vdd.n714 gnd 0.010223f
C3008 vdd.n715 gnd 0.010223f
C3009 vdd.n716 gnd 0.010223f
C3010 vdd.n717 gnd 0.010223f
C3011 vdd.n718 gnd 0.008228f
C3012 vdd.n719 gnd 0.010223f
C3013 vdd.n720 gnd 0.010223f
C3014 vdd.n721 gnd 0.010223f
C3015 vdd.n722 gnd 0.008146f
C3016 vdd.t29 gnd 0.125764f
C3017 vdd.t30 gnd 0.134407f
C3018 vdd.t28 gnd 0.164246f
C3019 vdd.n723 gnd 0.210541f
C3020 vdd.n724 gnd 0.176892f
C3021 vdd.n725 gnd 0.010223f
C3022 vdd.n726 gnd 0.008228f
C3023 vdd.n728 gnd 0.010223f
C3024 vdd.n730 gnd 0.010223f
C3025 vdd.n731 gnd 0.010223f
C3026 vdd.n732 gnd 0.008228f
C3027 vdd.n733 gnd 0.010223f
C3028 vdd.n734 gnd 0.010223f
C3029 vdd.n735 gnd 0.010223f
C3030 vdd.n736 gnd 0.010223f
C3031 vdd.n737 gnd 0.010223f
C3032 vdd.n738 gnd 0.008228f
C3033 vdd.n739 gnd 0.010223f
C3034 vdd.n740 gnd 0.010223f
C3035 vdd.n741 gnd 0.010223f
C3036 vdd.n742 gnd 0.010223f
C3037 vdd.n743 gnd 0.010223f
C3038 vdd.n744 gnd 0.008228f
C3039 vdd.n745 gnd 0.010223f
C3040 vdd.n746 gnd 0.010223f
C3041 vdd.n747 gnd 0.010223f
C3042 vdd.n748 gnd 0.006542f
C3043 vdd.n753 gnd 0.006951f
C3044 vdd.n754 gnd 0.006951f
C3045 vdd.n755 gnd 0.006951f
C3046 vdd.n756 gnd 8.91126f
C3047 vdd.n757 gnd 0.006951f
C3048 vdd.n758 gnd 0.006951f
C3049 vdd.n759 gnd 0.006951f
C3050 vdd.n761 gnd 0.006951f
C3051 vdd.n762 gnd 0.006951f
C3052 vdd.n764 gnd 0.006951f
C3053 vdd.n765 gnd 0.00506f
C3054 vdd.n767 gnd 0.006951f
C3055 vdd.t15 gnd 0.280902f
C3056 vdd.t14 gnd 0.287539f
C3057 vdd.t12 gnd 0.183384f
C3058 vdd.n768 gnd 0.099109f
C3059 vdd.n769 gnd 0.056218f
C3060 vdd.n770 gnd 0.009935f
C3061 vdd.n771 gnd 0.01609f
C3062 vdd.n773 gnd 0.006951f
C3063 vdd.n774 gnd 0.710393f
C3064 vdd.n775 gnd 0.015227f
C3065 vdd.n776 gnd 0.015227f
C3066 vdd.n777 gnd 0.006951f
C3067 vdd.n778 gnd 0.016259f
C3068 vdd.n779 gnd 0.006951f
C3069 vdd.n780 gnd 0.006951f
C3070 vdd.n781 gnd 0.006951f
C3071 vdd.n782 gnd 0.006951f
C3072 vdd.n783 gnd 0.006951f
C3073 vdd.n785 gnd 0.006951f
C3074 vdd.n786 gnd 0.006951f
C3075 vdd.n788 gnd 0.006951f
C3076 vdd.n789 gnd 0.006951f
C3077 vdd.n791 gnd 0.006951f
C3078 vdd.n792 gnd 0.006951f
C3079 vdd.n794 gnd 0.006951f
C3080 vdd.n795 gnd 0.006951f
C3081 vdd.n797 gnd 0.006951f
C3082 vdd.n798 gnd 0.006951f
C3083 vdd.n800 gnd 0.006951f
C3084 vdd.n801 gnd 0.00506f
C3085 vdd.n803 gnd 0.006951f
C3086 vdd.t84 gnd 0.280902f
C3087 vdd.t83 gnd 0.287539f
C3088 vdd.t82 gnd 0.183384f
C3089 vdd.n804 gnd 0.099109f
C3090 vdd.n805 gnd 0.056218f
C3091 vdd.n806 gnd 0.009935f
C3092 vdd.n807 gnd 0.006951f
C3093 vdd.n808 gnd 0.006951f
C3094 vdd.t13 gnd 0.355197f
C3095 vdd.n809 gnd 0.006951f
C3096 vdd.n810 gnd 0.006951f
C3097 vdd.n811 gnd 0.006951f
C3098 vdd.n812 gnd 0.006951f
C3099 vdd.n813 gnd 0.006951f
C3100 vdd.n814 gnd 0.710393f
C3101 vdd.n815 gnd 0.006951f
C3102 vdd.n816 gnd 0.006951f
C3103 vdd.n817 gnd 0.6007f
C3104 vdd.n818 gnd 0.006951f
C3105 vdd.n819 gnd 0.006951f
C3106 vdd.n820 gnd 0.006951f
C3107 vdd.n821 gnd 0.006951f
C3108 vdd.n822 gnd 0.694723f
C3109 vdd.n823 gnd 0.006951f
C3110 vdd.n824 gnd 0.006951f
C3111 vdd.n825 gnd 0.006951f
C3112 vdd.n826 gnd 0.006951f
C3113 vdd.n827 gnd 0.006951f
C3114 vdd.n828 gnd 0.710393f
C3115 vdd.n829 gnd 0.006951f
C3116 vdd.n830 gnd 0.006951f
C3117 vdd.t104 gnd 0.355197f
C3118 vdd.n831 gnd 0.006951f
C3119 vdd.n832 gnd 0.006951f
C3120 vdd.n833 gnd 0.006951f
C3121 vdd.t89 gnd 0.355197f
C3122 vdd.n834 gnd 0.006951f
C3123 vdd.n835 gnd 0.006951f
C3124 vdd.n836 gnd 0.006951f
C3125 vdd.n837 gnd 0.006951f
C3126 vdd.n838 gnd 0.006951f
C3127 vdd.t35 gnd 0.297738f
C3128 vdd.n839 gnd 0.006951f
C3129 vdd.n840 gnd 0.006951f
C3130 vdd.n841 gnd 0.569359f
C3131 vdd.n842 gnd 0.006951f
C3132 vdd.t36 gnd 0.287539f
C3133 vdd.t34 gnd 0.183384f
C3134 vdd.t37 gnd 0.287539f
C3135 vdd.n843 gnd 0.161608f
C3136 vdd.n844 gnd 0.006951f
C3137 vdd.n845 gnd 0.006951f
C3138 vdd.n846 gnd 0.454443f
C3139 vdd.n847 gnd 0.006951f
C3140 vdd.n848 gnd 0.006951f
C3141 vdd.t92 gnd 0.10447f
C3142 vdd.n849 gnd 0.412655f
C3143 vdd.n850 gnd 0.006951f
C3144 vdd.n851 gnd 0.006951f
C3145 vdd.n852 gnd 0.006951f
C3146 vdd.n853 gnd 0.611147f
C3147 vdd.n854 gnd 0.006951f
C3148 vdd.n855 gnd 0.006951f
C3149 vdd.t111 gnd 0.355197f
C3150 vdd.n856 gnd 0.006951f
C3151 vdd.n857 gnd 0.006951f
C3152 vdd.n858 gnd 0.006951f
C3153 vdd.t266 gnd 0.355197f
C3154 vdd.n859 gnd 0.006951f
C3155 vdd.n860 gnd 0.006951f
C3156 vdd.t249 gnd 0.355197f
C3157 vdd.n861 gnd 0.006951f
C3158 vdd.n862 gnd 0.006951f
C3159 vdd.n863 gnd 0.006951f
C3160 vdd.t97 gnd 0.282068f
C3161 vdd.n864 gnd 0.006951f
C3162 vdd.n865 gnd 0.006951f
C3163 vdd.n866 gnd 0.58503f
C3164 vdd.n867 gnd 0.006951f
C3165 vdd.n868 gnd 0.006951f
C3166 vdd.n869 gnd 0.006951f
C3167 vdd.t96 gnd 0.355197f
C3168 vdd.n870 gnd 0.006951f
C3169 vdd.n871 gnd 0.006951f
C3170 vdd.t105 gnd 0.297738f
C3171 vdd.n872 gnd 0.428325f
C3172 vdd.n873 gnd 0.006951f
C3173 vdd.n874 gnd 0.006951f
C3174 vdd.n875 gnd 0.006951f
C3175 vdd.n876 gnd 0.370867f
C3176 vdd.n877 gnd 0.006951f
C3177 vdd.n878 gnd 0.006951f
C3178 vdd.t254 gnd 0.355197f
C3179 vdd.n879 gnd 0.006951f
C3180 vdd.n880 gnd 0.006951f
C3181 vdd.n881 gnd 0.006951f
C3182 vdd.n882 gnd 0.710393f
C3183 vdd.n883 gnd 0.006951f
C3184 vdd.n884 gnd 0.006951f
C3185 vdd.t107 gnd 0.24028f
C3186 vdd.t260 gnd 0.339526f
C3187 vdd.n885 gnd 0.006951f
C3188 vdd.n886 gnd 0.006951f
C3189 vdd.n887 gnd 0.006951f
C3190 vdd.n888 gnd 0.532795f
C3191 vdd.n889 gnd 0.006951f
C3192 vdd.n890 gnd 0.006951f
C3193 vdd.n891 gnd 0.006951f
C3194 vdd.n892 gnd 0.006951f
C3195 vdd.n893 gnd 0.006951f
C3196 vdd.t63 gnd 0.355197f
C3197 vdd.n894 gnd 0.006951f
C3198 vdd.n895 gnd 0.006951f
C3199 vdd.t98 gnd 0.355197f
C3200 vdd.n896 gnd 0.006951f
C3201 vdd.n897 gnd 0.015227f
C3202 vdd.n898 gnd 0.015227f
C3203 vdd.n899 gnd 0.846204f
C3204 vdd.n900 gnd 0.006951f
C3205 vdd.n901 gnd 0.006951f
C3206 vdd.t252 gnd 0.355197f
C3207 vdd.n902 gnd 0.015227f
C3208 vdd.n903 gnd 0.006951f
C3209 vdd.n904 gnd 0.006951f
C3210 vdd.t245 gnd 0.647711f
C3211 vdd.n922 gnd 0.016259f
C3212 vdd.n940 gnd 0.015227f
C3213 vdd.n941 gnd 0.006951f
C3214 vdd.n942 gnd 0.015227f
C3215 vdd.t78 gnd 0.280902f
C3216 vdd.t77 gnd 0.287539f
C3217 vdd.t76 gnd 0.183384f
C3218 vdd.n943 gnd 0.099109f
C3219 vdd.n944 gnd 0.056218f
C3220 vdd.n945 gnd 0.01609f
C3221 vdd.n946 gnd 0.006951f
C3222 vdd.n947 gnd 0.376091f
C3223 vdd.n948 gnd 0.015227f
C3224 vdd.n949 gnd 0.006951f
C3225 vdd.n950 gnd 0.016259f
C3226 vdd.n951 gnd 0.006951f
C3227 vdd.t61 gnd 0.280902f
C3228 vdd.t60 gnd 0.287539f
C3229 vdd.t58 gnd 0.183384f
C3230 vdd.n952 gnd 0.099109f
C3231 vdd.n953 gnd 0.056218f
C3232 vdd.n954 gnd 0.009935f
C3233 vdd.n955 gnd 0.006951f
C3234 vdd.n956 gnd 0.006951f
C3235 vdd.t59 gnd 0.355197f
C3236 vdd.n957 gnd 0.006951f
C3237 vdd.t243 gnd 0.355197f
C3238 vdd.n958 gnd 0.006951f
C3239 vdd.n959 gnd 0.006951f
C3240 vdd.n960 gnd 0.006951f
C3241 vdd.n961 gnd 0.006951f
C3242 vdd.n962 gnd 0.006951f
C3243 vdd.n963 gnd 0.710393f
C3244 vdd.n964 gnd 0.006951f
C3245 vdd.n965 gnd 0.006951f
C3246 vdd.t264 gnd 0.355197f
C3247 vdd.n966 gnd 0.006951f
C3248 vdd.n967 gnd 0.006951f
C3249 vdd.n968 gnd 0.006951f
C3250 vdd.n969 gnd 0.006951f
C3251 vdd.n970 gnd 0.470113f
C3252 vdd.n971 gnd 0.006951f
C3253 vdd.n972 gnd 0.006951f
C3254 vdd.n973 gnd 0.006951f
C3255 vdd.n974 gnd 0.006951f
C3256 vdd.n975 gnd 0.006951f
C3257 vdd.n976 gnd 0.626818f
C3258 vdd.n977 gnd 0.006951f
C3259 vdd.n978 gnd 0.006951f
C3260 vdd.t250 gnd 0.339526f
C3261 vdd.t112 gnd 0.24028f
C3262 vdd.n979 gnd 0.006951f
C3263 vdd.n980 gnd 0.006951f
C3264 vdd.n981 gnd 0.006951f
C3265 vdd.t110 gnd 0.355197f
C3266 vdd.n982 gnd 0.006951f
C3267 vdd.n983 gnd 0.006951f
C3268 vdd.t108 gnd 0.355197f
C3269 vdd.n984 gnd 0.006951f
C3270 vdd.n985 gnd 0.006951f
C3271 vdd.n986 gnd 0.006951f
C3272 vdd.t262 gnd 0.297738f
C3273 vdd.n987 gnd 0.006951f
C3274 vdd.n988 gnd 0.006951f
C3275 vdd.n989 gnd 0.569359f
C3276 vdd.n990 gnd 0.006951f
C3277 vdd.n991 gnd 0.006951f
C3278 vdd.n992 gnd 0.006951f
C3279 vdd.t256 gnd 0.355197f
C3280 vdd.n993 gnd 0.006951f
C3281 vdd.n994 gnd 0.006951f
C3282 vdd.t88 gnd 0.282068f
C3283 vdd.n995 gnd 0.412655f
C3284 vdd.n996 gnd 0.006951f
C3285 vdd.n997 gnd 0.006951f
C3286 vdd.n998 gnd 0.006951f
C3287 vdd.n999 gnd 0.611147f
C3288 vdd.n1000 gnd 0.006951f
C3289 vdd.n1001 gnd 0.006951f
C3290 vdd.t103 gnd 0.355197f
C3291 vdd.n1002 gnd 0.006951f
C3292 vdd.n1003 gnd 0.006951f
C3293 vdd.n1004 gnd 0.006951f
C3294 vdd.n1005 gnd 0.710393f
C3295 vdd.n1006 gnd 0.006951f
C3296 vdd.n1007 gnd 0.006951f
C3297 vdd.t100 gnd 0.355197f
C3298 vdd.n1008 gnd 0.006951f
C3299 vdd.n1009 gnd 0.006951f
C3300 vdd.n1010 gnd 0.006951f
C3301 vdd.t93 gnd 0.10447f
C3302 vdd.n1011 gnd 0.006951f
C3303 vdd.n1012 gnd 0.006951f
C3304 vdd.n1013 gnd 0.006951f
C3305 vdd.t68 gnd 0.287539f
C3306 vdd.t66 gnd 0.183384f
C3307 vdd.t69 gnd 0.287539f
C3308 vdd.n1014 gnd 0.161608f
C3309 vdd.n1015 gnd 0.006951f
C3310 vdd.n1016 gnd 0.006951f
C3311 vdd.t95 gnd 0.355197f
C3312 vdd.n1017 gnd 0.006951f
C3313 vdd.n1018 gnd 0.006951f
C3314 vdd.t67 gnd 0.297738f
C3315 vdd.n1019 gnd 0.605924f
C3316 vdd.n1020 gnd 0.006951f
C3317 vdd.n1021 gnd 0.006951f
C3318 vdd.n1022 gnd 0.006951f
C3319 vdd.n1023 gnd 0.370867f
C3320 vdd.n1024 gnd 0.006951f
C3321 vdd.n1025 gnd 0.006951f
C3322 vdd.n1026 gnd 0.496231f
C3323 vdd.n1027 gnd 0.006951f
C3324 vdd.n1028 gnd 0.006951f
C3325 vdd.n1029 gnd 0.006951f
C3326 vdd.n1030 gnd 0.710393f
C3327 vdd.n1031 gnd 0.006951f
C3328 vdd.n1032 gnd 0.006951f
C3329 vdd.t94 gnd 0.355197f
C3330 vdd.n1033 gnd 0.006951f
C3331 vdd.n1034 gnd 0.006951f
C3332 vdd.n1035 gnd 0.006951f
C3333 vdd.n1036 gnd 0.710393f
C3334 vdd.n1037 gnd 0.006951f
C3335 vdd.n1038 gnd 0.006951f
C3336 vdd.n1039 gnd 0.006951f
C3337 vdd.n1040 gnd 0.006951f
C3338 vdd.n1041 gnd 0.006951f
C3339 vdd.t17 gnd 0.355197f
C3340 vdd.n1042 gnd 0.006951f
C3341 vdd.n1043 gnd 0.006951f
C3342 vdd.n1044 gnd 0.006951f
C3343 vdd.n1045 gnd 0.015227f
C3344 vdd.n1046 gnd 0.015227f
C3345 vdd.n1047 gnd 1.00291f
C3346 vdd.n1048 gnd 0.006951f
C3347 vdd.n1049 gnd 0.006951f
C3348 vdd.n1050 gnd 0.46489f
C3349 vdd.n1051 gnd 0.015227f
C3350 vdd.n1052 gnd 0.006951f
C3351 vdd.n1053 gnd 0.006951f
C3352 vdd.n1054 gnd 9.1202f
C3353 vdd.n1087 gnd 0.016259f
C3354 vdd.n1088 gnd 0.006951f
C3355 vdd.n1089 gnd 0.006951f
C3356 vdd.n1090 gnd 0.006951f
C3357 vdd.n1091 gnd 0.006542f
C3358 vdd.n1094 gnd 0.023438f
C3359 vdd.n1095 gnd 0.006829f
C3360 vdd.n1096 gnd 0.008228f
C3361 vdd.n1098 gnd 0.010223f
C3362 vdd.n1099 gnd 0.010223f
C3363 vdd.n1100 gnd 0.008228f
C3364 vdd.n1102 gnd 0.010223f
C3365 vdd.n1103 gnd 0.010223f
C3366 vdd.n1104 gnd 0.010223f
C3367 vdd.n1105 gnd 0.010223f
C3368 vdd.n1106 gnd 0.010223f
C3369 vdd.n1107 gnd 0.008228f
C3370 vdd.n1109 gnd 0.010223f
C3371 vdd.n1110 gnd 0.010223f
C3372 vdd.n1111 gnd 0.010223f
C3373 vdd.n1112 gnd 0.010223f
C3374 vdd.n1113 gnd 0.010223f
C3375 vdd.n1114 gnd 0.008228f
C3376 vdd.n1116 gnd 0.010223f
C3377 vdd.n1117 gnd 0.010223f
C3378 vdd.n1118 gnd 0.010223f
C3379 vdd.n1119 gnd 0.010223f
C3380 vdd.n1120 gnd 0.00687f
C3381 vdd.t72 gnd 0.125764f
C3382 vdd.t71 gnd 0.134407f
C3383 vdd.t70 gnd 0.164246f
C3384 vdd.n1121 gnd 0.210541f
C3385 vdd.n1122 gnd 0.176892f
C3386 vdd.n1124 gnd 0.010223f
C3387 vdd.n1125 gnd 0.010223f
C3388 vdd.n1126 gnd 0.008228f
C3389 vdd.n1127 gnd 0.010223f
C3390 vdd.n1129 gnd 0.010223f
C3391 vdd.n1130 gnd 0.010223f
C3392 vdd.n1131 gnd 0.010223f
C3393 vdd.n1132 gnd 0.010223f
C3394 vdd.n1133 gnd 0.008228f
C3395 vdd.n1135 gnd 0.010223f
C3396 vdd.n1136 gnd 0.010223f
C3397 vdd.n1137 gnd 0.010223f
C3398 vdd.n1138 gnd 0.010223f
C3399 vdd.n1139 gnd 0.010223f
C3400 vdd.n1140 gnd 0.008228f
C3401 vdd.n1142 gnd 0.010223f
C3402 vdd.n1143 gnd 0.010223f
C3403 vdd.n1144 gnd 0.010223f
C3404 vdd.n1145 gnd 0.010223f
C3405 vdd.n1146 gnd 0.010223f
C3406 vdd.n1147 gnd 0.008228f
C3407 vdd.n1149 gnd 0.010223f
C3408 vdd.n1150 gnd 0.010223f
C3409 vdd.n1151 gnd 0.010223f
C3410 vdd.n1152 gnd 0.010223f
C3411 vdd.n1153 gnd 0.010223f
C3412 vdd.n1154 gnd 0.008228f
C3413 vdd.n1156 gnd 0.010223f
C3414 vdd.n1157 gnd 0.010223f
C3415 vdd.n1158 gnd 0.010223f
C3416 vdd.n1159 gnd 0.010223f
C3417 vdd.n1160 gnd 0.008146f
C3418 vdd.t57 gnd 0.125764f
C3419 vdd.t56 gnd 0.134407f
C3420 vdd.t55 gnd 0.164246f
C3421 vdd.n1161 gnd 0.210541f
C3422 vdd.n1162 gnd 0.176892f
C3423 vdd.n1164 gnd 0.010223f
C3424 vdd.n1165 gnd 0.010223f
C3425 vdd.n1166 gnd 0.008228f
C3426 vdd.n1167 gnd 0.010223f
C3427 vdd.n1169 gnd 0.010223f
C3428 vdd.n1170 gnd 0.010223f
C3429 vdd.n1171 gnd 0.010223f
C3430 vdd.n1172 gnd 0.010223f
C3431 vdd.n1173 gnd 0.008228f
C3432 vdd.n1175 gnd 0.010223f
C3433 vdd.n1176 gnd 0.010223f
C3434 vdd.n1177 gnd 0.010223f
C3435 vdd.n1178 gnd 0.010223f
C3436 vdd.n1179 gnd 0.010223f
C3437 vdd.n1180 gnd 0.008228f
C3438 vdd.n1182 gnd 0.010223f
C3439 vdd.n1183 gnd 0.010223f
C3440 vdd.n1184 gnd 0.010223f
C3441 vdd.n1185 gnd 0.010223f
C3442 vdd.n1186 gnd 0.010223f
C3443 vdd.n1187 gnd 0.008228f
C3444 vdd.n1189 gnd 0.010223f
C3445 vdd.n1190 gnd 0.010223f
C3446 vdd.n1191 gnd 0.006542f
C3447 vdd.n1192 gnd 0.008228f
C3448 vdd.n1193 gnd 0.006951f
C3449 vdd.n1194 gnd 0.006951f
C3450 vdd.n1195 gnd 0.006951f
C3451 vdd.n1196 gnd 0.006951f
C3452 vdd.n1197 gnd 0.006951f
C3453 vdd.n1198 gnd 0.006951f
C3454 vdd.n1199 gnd 0.006951f
C3455 vdd.n1200 gnd 0.006951f
C3456 vdd.n1201 gnd 0.006951f
C3457 vdd.n1202 gnd 0.006951f
C3458 vdd.n1203 gnd 0.006951f
C3459 vdd.n1204 gnd 0.006951f
C3460 vdd.n1205 gnd 0.006951f
C3461 vdd.n1206 gnd 0.006951f
C3462 vdd.n1207 gnd 0.006951f
C3463 vdd.n1208 gnd 0.006951f
C3464 vdd.n1209 gnd 0.006951f
C3465 vdd.n1210 gnd 0.006951f
C3466 vdd.n1211 gnd 0.006951f
C3467 vdd.n1212 gnd 0.006951f
C3468 vdd.n1213 gnd 0.006951f
C3469 vdd.n1214 gnd 0.006951f
C3470 vdd.n1215 gnd 0.006951f
C3471 vdd.n1216 gnd 0.006951f
C3472 vdd.n1217 gnd 0.006951f
C3473 vdd.n1218 gnd 0.006951f
C3474 vdd.n1219 gnd 0.006951f
C3475 vdd.n1220 gnd 0.006951f
C3476 vdd.n1221 gnd 0.006951f
C3477 vdd.n1222 gnd 0.006951f
C3478 vdd.n1223 gnd 0.006951f
C3479 vdd.t18 gnd 0.280902f
C3480 vdd.t19 gnd 0.287539f
C3481 vdd.t16 gnd 0.183384f
C3482 vdd.n1224 gnd 0.099109f
C3483 vdd.n1225 gnd 0.056218f
C3484 vdd.n1226 gnd 0.009935f
C3485 vdd.n1227 gnd 0.006951f
C3486 vdd.n1228 gnd 0.006951f
C3487 vdd.n1229 gnd 0.006951f
C3488 vdd.n1230 gnd 0.006951f
C3489 vdd.n1231 gnd 0.006951f
C3490 vdd.n1232 gnd 0.006951f
C3491 vdd.n1233 gnd 0.006951f
C3492 vdd.n1234 gnd 0.006951f
C3493 vdd.n1235 gnd 0.006951f
C3494 vdd.n1236 gnd 0.006951f
C3495 vdd.n1237 gnd 0.006951f
C3496 vdd.n1238 gnd 0.006951f
C3497 vdd.n1239 gnd 0.006951f
C3498 vdd.n1240 gnd 0.006951f
C3499 vdd.n1241 gnd 0.006951f
C3500 vdd.n1242 gnd 0.006951f
C3501 vdd.n1243 gnd 0.006951f
C3502 vdd.t32 gnd 0.280902f
C3503 vdd.t33 gnd 0.287539f
C3504 vdd.t31 gnd 0.183384f
C3505 vdd.n1244 gnd 0.099109f
C3506 vdd.n1245 gnd 0.056218f
C3507 vdd.n1246 gnd 0.006951f
C3508 vdd.n1247 gnd 0.006951f
C3509 vdd.n1248 gnd 0.006951f
C3510 vdd.n1249 gnd 0.006951f
C3511 vdd.n1250 gnd 0.006951f
C3512 vdd.n1251 gnd 0.006951f
C3513 vdd.n1252 gnd 0.006951f
C3514 vdd.n1253 gnd 0.006951f
C3515 vdd.n1254 gnd 0.006951f
C3516 vdd.n1255 gnd 0.006951f
C3517 vdd.n1256 gnd 0.006951f
C3518 vdd.n1257 gnd 0.006951f
C3519 vdd.n1258 gnd 0.006951f
C3520 vdd.n1259 gnd 0.006951f
C3521 vdd.n1260 gnd 0.006951f
C3522 vdd.n1261 gnd 0.006951f
C3523 vdd.n1262 gnd 0.006951f
C3524 vdd.n1263 gnd 0.006951f
C3525 vdd.n1264 gnd 0.006951f
C3526 vdd.n1265 gnd 0.006951f
C3527 vdd.n1266 gnd 0.006951f
C3528 vdd.n1267 gnd 0.006951f
C3529 vdd.n1268 gnd 0.006951f
C3530 vdd.n1269 gnd 0.006951f
C3531 vdd.n1270 gnd 0.006951f
C3532 vdd.n1271 gnd 0.006951f
C3533 vdd.n1272 gnd 0.00506f
C3534 vdd.n1273 gnd 0.009935f
C3535 vdd.n1274 gnd 0.005367f
C3536 vdd.n1275 gnd 0.006951f
C3537 vdd.n1276 gnd 0.006951f
C3538 vdd.n1277 gnd 0.006951f
C3539 vdd.n1278 gnd 0.016259f
C3540 vdd.n1279 gnd 0.016259f
C3541 vdd.n1280 gnd 0.015227f
C3542 vdd.n1281 gnd 0.015227f
C3543 vdd.n1282 gnd 0.006951f
C3544 vdd.n1283 gnd 0.006951f
C3545 vdd.n1284 gnd 0.006951f
C3546 vdd.n1285 gnd 0.006951f
C3547 vdd.n1286 gnd 0.006951f
C3548 vdd.n1287 gnd 0.006951f
C3549 vdd.n1288 gnd 0.006951f
C3550 vdd.n1289 gnd 0.006951f
C3551 vdd.n1290 gnd 0.006951f
C3552 vdd.n1291 gnd 0.006951f
C3553 vdd.n1292 gnd 0.006951f
C3554 vdd.n1293 gnd 0.006951f
C3555 vdd.n1294 gnd 0.006951f
C3556 vdd.n1295 gnd 0.006951f
C3557 vdd.n1296 gnd 0.006951f
C3558 vdd.n1297 gnd 0.006951f
C3559 vdd.n1298 gnd 0.006951f
C3560 vdd.n1299 gnd 0.006951f
C3561 vdd.n1300 gnd 0.006951f
C3562 vdd.n1301 gnd 0.006951f
C3563 vdd.n1302 gnd 0.006951f
C3564 vdd.n1303 gnd 0.006951f
C3565 vdd.n1304 gnd 0.006951f
C3566 vdd.n1305 gnd 0.006951f
C3567 vdd.n1306 gnd 0.006951f
C3568 vdd.n1307 gnd 0.006951f
C3569 vdd.n1308 gnd 0.006951f
C3570 vdd.n1309 gnd 0.423102f
C3571 vdd.n1310 gnd 0.006951f
C3572 vdd.n1311 gnd 0.006951f
C3573 vdd.n1312 gnd 0.006951f
C3574 vdd.n1313 gnd 0.006951f
C3575 vdd.n1314 gnd 0.006951f
C3576 vdd.n1315 gnd 0.006951f
C3577 vdd.n1316 gnd 0.006951f
C3578 vdd.n1317 gnd 0.006951f
C3579 vdd.n1318 gnd 0.006951f
C3580 vdd.n1319 gnd 0.006951f
C3581 vdd.n1320 gnd 0.006951f
C3582 vdd.n1321 gnd 0.006951f
C3583 vdd.n1322 gnd 0.006951f
C3584 vdd.n1323 gnd 0.006951f
C3585 vdd.n1324 gnd 0.006951f
C3586 vdd.n1325 gnd 0.006951f
C3587 vdd.n1326 gnd 0.006951f
C3588 vdd.n1327 gnd 0.006951f
C3589 vdd.n1328 gnd 0.006951f
C3590 vdd.n1329 gnd 0.006951f
C3591 vdd.n1330 gnd 0.22461f
C3592 vdd.n1331 gnd 0.006951f
C3593 vdd.n1332 gnd 0.006951f
C3594 vdd.n1333 gnd 0.006951f
C3595 vdd.n1334 gnd 0.006951f
C3596 vdd.n1335 gnd 0.006951f
C3597 vdd.n1336 gnd 0.006951f
C3598 vdd.n1337 gnd 0.006951f
C3599 vdd.n1338 gnd 0.006951f
C3600 vdd.n1339 gnd 0.006951f
C3601 vdd.n1340 gnd 0.006951f
C3602 vdd.n1341 gnd 0.006951f
C3603 vdd.n1342 gnd 0.006951f
C3604 vdd.n1343 gnd 0.006951f
C3605 vdd.n1344 gnd 0.006951f
C3606 vdd.n1345 gnd 0.006951f
C3607 vdd.n1346 gnd 0.006951f
C3608 vdd.n1347 gnd 0.006951f
C3609 vdd.n1348 gnd 0.006951f
C3610 vdd.n1349 gnd 0.006951f
C3611 vdd.n1350 gnd 0.006951f
C3612 vdd.n1351 gnd 0.006951f
C3613 vdd.n1352 gnd 0.006951f
C3614 vdd.n1353 gnd 0.006951f
C3615 vdd.n1354 gnd 0.006951f
C3616 vdd.n1355 gnd 0.006951f
C3617 vdd.n1356 gnd 0.006951f
C3618 vdd.n1357 gnd 0.006951f
C3619 vdd.n1358 gnd 0.015227f
C3620 vdd.n1359 gnd 0.015227f
C3621 vdd.n1360 gnd 0.016259f
C3622 vdd.n1361 gnd 0.006951f
C3623 vdd.n1362 gnd 0.006951f
C3624 vdd.n1363 gnd 0.005367f
C3625 vdd.n1364 gnd 0.006951f
C3626 vdd.n1365 gnd 0.006951f
C3627 vdd.n1366 gnd 0.00506f
C3628 vdd.n1367 gnd 0.006951f
C3629 vdd.n1368 gnd 0.006951f
C3630 vdd.n1369 gnd 0.006951f
C3631 vdd.n1370 gnd 0.006951f
C3632 vdd.n1371 gnd 0.006951f
C3633 vdd.n1372 gnd 0.006951f
C3634 vdd.n1373 gnd 0.006951f
C3635 vdd.n1374 gnd 0.006951f
C3636 vdd.n1375 gnd 0.006951f
C3637 vdd.n1376 gnd 0.006951f
C3638 vdd.n1377 gnd 0.006951f
C3639 vdd.n1378 gnd 0.006951f
C3640 vdd.n1379 gnd 0.006951f
C3641 vdd.n1380 gnd 0.006951f
C3642 vdd.n1381 gnd 0.006951f
C3643 vdd.n1382 gnd 0.006951f
C3644 vdd.n1383 gnd 0.006951f
C3645 vdd.n1384 gnd 0.006951f
C3646 vdd.n1385 gnd 0.006951f
C3647 vdd.n1386 gnd 0.006951f
C3648 vdd.n1387 gnd 0.006951f
C3649 vdd.n1388 gnd 0.006951f
C3650 vdd.n1389 gnd 0.006951f
C3651 vdd.n1390 gnd 0.006951f
C3652 vdd.n1391 gnd 0.006951f
C3653 vdd.n1392 gnd 0.006951f
C3654 vdd.n1393 gnd 0.027861f
C3655 vdd.n1395 gnd 0.023438f
C3656 vdd.n1396 gnd 0.008228f
C3657 vdd.n1398 gnd 0.010223f
C3658 vdd.n1399 gnd 0.008228f
C3659 vdd.n1400 gnd 0.010223f
C3660 vdd.n1402 gnd 0.010223f
C3661 vdd.n1403 gnd 0.010223f
C3662 vdd.n1405 gnd 0.010223f
C3663 vdd.n1406 gnd 0.006829f
C3664 vdd.n1407 gnd 0.579806f
C3665 vdd.n1408 gnd 0.010223f
C3666 vdd.n1409 gnd 0.023438f
C3667 vdd.n1410 gnd 0.008228f
C3668 vdd.n1411 gnd 0.010223f
C3669 vdd.n1412 gnd 0.008228f
C3670 vdd.n1413 gnd 0.010223f
C3671 vdd.n1414 gnd 1.0447f
C3672 vdd.n1415 gnd 0.010223f
C3673 vdd.n1416 gnd 0.008228f
C3674 vdd.n1417 gnd 0.008228f
C3675 vdd.n1418 gnd 0.010223f
C3676 vdd.n1419 gnd 0.008228f
C3677 vdd.n1420 gnd 0.010223f
C3678 vdd.t154 gnd 0.522348f
C3679 vdd.n1421 gnd 0.010223f
C3680 vdd.n1422 gnd 0.008228f
C3681 vdd.n1423 gnd 0.010223f
C3682 vdd.n1424 gnd 0.008228f
C3683 vdd.n1425 gnd 0.010223f
C3684 vdd.t117 gnd 0.522348f
C3685 vdd.n1426 gnd 0.010223f
C3686 vdd.n1427 gnd 0.008228f
C3687 vdd.n1428 gnd 0.010223f
C3688 vdd.n1429 gnd 0.008228f
C3689 vdd.n1430 gnd 0.010223f
C3690 vdd.t178 gnd 0.522348f
C3691 vdd.n1431 gnd 0.726064f
C3692 vdd.n1432 gnd 0.010223f
C3693 vdd.n1433 gnd 0.008228f
C3694 vdd.n1434 gnd 0.010223f
C3695 vdd.n1435 gnd 0.008228f
C3696 vdd.n1436 gnd 0.010223f
C3697 vdd.n1437 gnd 0.830533f
C3698 vdd.n1438 gnd 0.010223f
C3699 vdd.n1439 gnd 0.008228f
C3700 vdd.n1440 gnd 0.010223f
C3701 vdd.n1441 gnd 0.008228f
C3702 vdd.n1442 gnd 0.010223f
C3703 vdd.n1443 gnd 0.652935f
C3704 vdd.t196 gnd 0.522348f
C3705 vdd.n1444 gnd 0.010223f
C3706 vdd.n1445 gnd 0.008228f
C3707 vdd.n1446 gnd 0.010223f
C3708 vdd.n1447 gnd 0.008228f
C3709 vdd.n1448 gnd 0.010223f
C3710 vdd.t169 gnd 0.522348f
C3711 vdd.n1449 gnd 0.010223f
C3712 vdd.n1450 gnd 0.008228f
C3713 vdd.n1451 gnd 0.010223f
C3714 vdd.n1452 gnd 0.008228f
C3715 vdd.n1453 gnd 0.010223f
C3716 vdd.t131 gnd 0.522348f
C3717 vdd.n1454 gnd 0.569359f
C3718 vdd.n1455 gnd 0.010223f
C3719 vdd.n1456 gnd 0.008228f
C3720 vdd.n1457 gnd 0.010223f
C3721 vdd.n1458 gnd 0.008228f
C3722 vdd.n1459 gnd 0.010223f
C3723 vdd.t144 gnd 0.522348f
C3724 vdd.n1460 gnd 0.010223f
C3725 vdd.n1461 gnd 0.008228f
C3726 vdd.n1462 gnd 0.010223f
C3727 vdd.n1463 gnd 0.008228f
C3728 vdd.n1464 gnd 0.010223f
C3729 vdd.n1465 gnd 0.809639f
C3730 vdd.n1466 gnd 0.867098f
C3731 vdd.t190 gnd 0.522348f
C3732 vdd.n1467 gnd 0.010223f
C3733 vdd.n1468 gnd 0.008228f
C3734 vdd.n1469 gnd 0.010223f
C3735 vdd.n1470 gnd 0.008228f
C3736 vdd.n1471 gnd 0.010223f
C3737 vdd.n1472 gnd 0.632041f
C3738 vdd.n1473 gnd 0.010223f
C3739 vdd.n1474 gnd 0.008228f
C3740 vdd.n1475 gnd 0.010223f
C3741 vdd.n1476 gnd 0.008228f
C3742 vdd.n1477 gnd 0.010223f
C3743 vdd.t147 gnd 0.522348f
C3744 vdd.t123 gnd 0.522348f
C3745 vdd.n1478 gnd 0.010223f
C3746 vdd.n1479 gnd 0.008228f
C3747 vdd.n1480 gnd 0.010223f
C3748 vdd.n1481 gnd 0.008228f
C3749 vdd.n1482 gnd 0.010223f
C3750 vdd.t149 gnd 0.522348f
C3751 vdd.n1483 gnd 0.010223f
C3752 vdd.n1484 gnd 0.008228f
C3753 vdd.n1485 gnd 0.010223f
C3754 vdd.n1486 gnd 0.008228f
C3755 vdd.n1487 gnd 0.010223f
C3756 vdd.t115 gnd 0.522348f
C3757 vdd.n1488 gnd 0.767852f
C3758 vdd.n1489 gnd 0.010223f
C3759 vdd.n1490 gnd 0.008228f
C3760 vdd.n1491 gnd 0.010223f
C3761 vdd.n1492 gnd 0.008228f
C3762 vdd.n1493 gnd 0.010223f
C3763 vdd.n1494 gnd 1.0447f
C3764 vdd.n1495 gnd 0.010223f
C3765 vdd.n1496 gnd 0.008228f
C3766 vdd.n1497 gnd 0.010223f
C3767 vdd.n1498 gnd 0.008228f
C3768 vdd.n1499 gnd 0.010223f
C3769 vdd.n1500 gnd 0.882768f
C3770 vdd.n1501 gnd 0.010223f
C3771 vdd.n1502 gnd 0.008228f
C3772 vdd.n1503 gnd 0.023279f
C3773 vdd.n1504 gnd 0.006829f
C3774 vdd.n1505 gnd 0.023279f
C3775 vdd.n1506 gnd 1.379f
C3776 vdd.n1507 gnd 0.023279f
C3777 vdd.n1508 gnd 0.006829f
C3778 vdd.n1509 gnd 0.010223f
C3779 vdd.t50 gnd 0.125764f
C3780 vdd.t51 gnd 0.134407f
C3781 vdd.t49 gnd 0.164246f
C3782 vdd.n1510 gnd 0.210541f
C3783 vdd.n1511 gnd 0.177715f
C3784 vdd.n1512 gnd 0.013494f
C3785 vdd.n1513 gnd 0.010223f
C3786 vdd.n1544 gnd 0.010223f
C3787 vdd.n1545 gnd 0.010223f
C3788 vdd.n1546 gnd 0.023438f
C3789 vdd.n1547 gnd 0.008228f
C3790 vdd.n1548 gnd 0.010223f
C3791 vdd.n1549 gnd 0.010223f
C3792 vdd.n1550 gnd 0.010223f
C3793 vdd.n1551 gnd 0.010223f
C3794 vdd.n1552 gnd 0.008228f
C3795 vdd.n1553 gnd 0.010223f
C3796 vdd.n1554 gnd 0.010223f
C3797 vdd.n1555 gnd 0.010223f
C3798 vdd.n1556 gnd 0.010223f
C3799 vdd.n1557 gnd 0.010223f
C3800 vdd.n1558 gnd 0.008228f
C3801 vdd.n1559 gnd 0.010223f
C3802 vdd.n1560 gnd 0.010223f
C3803 vdd.n1561 gnd 0.010223f
C3804 vdd.n1562 gnd 0.010223f
C3805 vdd.n1563 gnd 0.010223f
C3806 vdd.n1564 gnd 0.008228f
C3807 vdd.n1565 gnd 0.010223f
C3808 vdd.n1566 gnd 0.010223f
C3809 vdd.n1567 gnd 0.010223f
C3810 vdd.n1568 gnd 0.010223f
C3811 vdd.n1569 gnd 0.010223f
C3812 vdd.n1570 gnd 0.00687f
C3813 vdd.n1571 gnd 0.010223f
C3814 vdd.n1572 gnd 0.010223f
C3815 vdd.n1573 gnd 0.010223f
C3816 vdd.n1574 gnd 0.008228f
C3817 vdd.n1575 gnd 0.010223f
C3818 vdd.n1576 gnd 0.010223f
C3819 vdd.n1577 gnd 0.010223f
C3820 vdd.n1578 gnd 0.010223f
C3821 vdd.n1579 gnd 0.010223f
C3822 vdd.n1580 gnd 0.008228f
C3823 vdd.n1581 gnd 0.010223f
C3824 vdd.n1582 gnd 0.010223f
C3825 vdd.n1583 gnd 0.010223f
C3826 vdd.n1584 gnd 0.010223f
C3827 vdd.n1585 gnd 0.010223f
C3828 vdd.n1586 gnd 0.008228f
C3829 vdd.n1587 gnd 0.010223f
C3830 vdd.n1588 gnd 0.010223f
C3831 vdd.n1589 gnd 0.010223f
C3832 vdd.n1590 gnd 0.010223f
C3833 vdd.n1591 gnd 0.010223f
C3834 vdd.n1592 gnd 0.008228f
C3835 vdd.n1593 gnd 0.010223f
C3836 vdd.n1594 gnd 0.010223f
C3837 vdd.n1595 gnd 0.010223f
C3838 vdd.n1596 gnd 0.010223f
C3839 vdd.n1597 gnd 0.010223f
C3840 vdd.n1598 gnd 0.008228f
C3841 vdd.n1599 gnd 0.010223f
C3842 vdd.n1600 gnd 0.010223f
C3843 vdd.n1601 gnd 0.010223f
C3844 vdd.n1602 gnd 0.010223f
C3845 vdd.n1603 gnd 0.008146f
C3846 vdd.n1604 gnd 0.010223f
C3847 vdd.n1605 gnd 0.010223f
C3848 vdd.n1606 gnd 0.010223f
C3849 vdd.n1607 gnd 0.010223f
C3850 vdd.n1608 gnd 0.010223f
C3851 vdd.n1609 gnd 0.008228f
C3852 vdd.n1610 gnd 0.010223f
C3853 vdd.n1611 gnd 0.010223f
C3854 vdd.n1612 gnd 0.010223f
C3855 vdd.n1613 gnd 0.010223f
C3856 vdd.n1614 gnd 0.010223f
C3857 vdd.n1615 gnd 0.008228f
C3858 vdd.n1616 gnd 0.010223f
C3859 vdd.n1617 gnd 0.010223f
C3860 vdd.n1618 gnd 0.010223f
C3861 vdd.n1619 gnd 0.010223f
C3862 vdd.n1620 gnd 0.010223f
C3863 vdd.n1621 gnd 0.008228f
C3864 vdd.n1622 gnd 0.010223f
C3865 vdd.n1623 gnd 0.010223f
C3866 vdd.n1624 gnd 0.010223f
C3867 vdd.n1625 gnd 0.010223f
C3868 vdd.n1626 gnd 0.010223f
C3869 vdd.n1627 gnd 0.008228f
C3870 vdd.n1628 gnd 0.010223f
C3871 vdd.n1629 gnd 0.010223f
C3872 vdd.n1630 gnd 0.010223f
C3873 vdd.n1631 gnd 0.010223f
C3874 vdd.n1632 gnd 0.010223f
C3875 vdd.n1633 gnd 0.00432f
C3876 vdd.n1634 gnd 0.010223f
C3877 vdd.n1635 gnd 0.008228f
C3878 vdd.n1636 gnd 0.008228f
C3879 vdd.n1637 gnd 0.008228f
C3880 vdd.n1638 gnd 0.010223f
C3881 vdd.n1639 gnd 0.010223f
C3882 vdd.n1640 gnd 0.010223f
C3883 vdd.n1641 gnd 0.008228f
C3884 vdd.n1642 gnd 0.008228f
C3885 vdd.n1643 gnd 0.008228f
C3886 vdd.n1644 gnd 0.010223f
C3887 vdd.n1645 gnd 0.010223f
C3888 vdd.n1646 gnd 0.010223f
C3889 vdd.n1647 gnd 0.008228f
C3890 vdd.n1648 gnd 0.008228f
C3891 vdd.n1649 gnd 0.008228f
C3892 vdd.n1650 gnd 0.010223f
C3893 vdd.n1651 gnd 0.010223f
C3894 vdd.n1652 gnd 0.010223f
C3895 vdd.n1653 gnd 0.008228f
C3896 vdd.n1654 gnd 0.008228f
C3897 vdd.n1655 gnd 0.008228f
C3898 vdd.n1656 gnd 0.010223f
C3899 vdd.n1657 gnd 0.010223f
C3900 vdd.n1658 gnd 0.010223f
C3901 vdd.n1659 gnd 0.008228f
C3902 vdd.n1660 gnd 0.008228f
C3903 vdd.n1661 gnd 0.008228f
C3904 vdd.n1662 gnd 0.010223f
C3905 vdd.n1663 gnd 0.010223f
C3906 vdd.n1664 gnd 0.010223f
C3907 vdd.n1665 gnd 0.010223f
C3908 vdd.t43 gnd 0.125764f
C3909 vdd.t44 gnd 0.134407f
C3910 vdd.t41 gnd 0.164246f
C3911 vdd.n1666 gnd 0.210541f
C3912 vdd.n1667 gnd 0.177715f
C3913 vdd.n1668 gnd 0.017608f
C3914 vdd.n1669 gnd 0.005595f
C3915 vdd.n1670 gnd 0.008228f
C3916 vdd.n1671 gnd 0.010223f
C3917 vdd.n1672 gnd 0.010223f
C3918 vdd.n1673 gnd 0.010223f
C3919 vdd.n1674 gnd 0.008228f
C3920 vdd.n1675 gnd 0.008228f
C3921 vdd.n1676 gnd 0.008228f
C3922 vdd.n1677 gnd 0.010223f
C3923 vdd.n1678 gnd 0.010223f
C3924 vdd.n1679 gnd 0.010223f
C3925 vdd.n1680 gnd 0.008228f
C3926 vdd.n1681 gnd 0.008228f
C3927 vdd.n1682 gnd 0.008228f
C3928 vdd.n1683 gnd 0.010223f
C3929 vdd.n1684 gnd 0.010223f
C3930 vdd.n1685 gnd 0.010223f
C3931 vdd.n1686 gnd 0.008228f
C3932 vdd.n1687 gnd 0.008228f
C3933 vdd.n1688 gnd 0.008228f
C3934 vdd.n1689 gnd 0.010223f
C3935 vdd.n1690 gnd 0.010223f
C3936 vdd.n1691 gnd 0.010223f
C3937 vdd.n1692 gnd 0.008228f
C3938 vdd.n1693 gnd 0.008228f
C3939 vdd.n1694 gnd 0.008228f
C3940 vdd.n1695 gnd 0.010223f
C3941 vdd.n1696 gnd 0.010223f
C3942 vdd.n1697 gnd 0.010223f
C3943 vdd.n1698 gnd 0.008228f
C3944 vdd.n1699 gnd 0.00687f
C3945 vdd.n1700 gnd 0.010223f
C3946 vdd.n1701 gnd 0.010223f
C3947 vdd.t53 gnd 0.125764f
C3948 vdd.t54 gnd 0.134407f
C3949 vdd.t52 gnd 0.164246f
C3950 vdd.n1702 gnd 0.210541f
C3951 vdd.n1703 gnd 0.177715f
C3952 vdd.n1704 gnd 0.017608f
C3953 vdd.n1705 gnd 0.010223f
C3954 vdd.n1706 gnd 0.010223f
C3955 vdd.n1707 gnd 0.010223f
C3956 vdd.n1708 gnd 0.008228f
C3957 vdd.n1709 gnd 0.008228f
C3958 vdd.n1710 gnd 0.008228f
C3959 vdd.n1711 gnd 0.010223f
C3960 vdd.n1712 gnd 0.010223f
C3961 vdd.n1713 gnd 0.010223f
C3962 vdd.n1714 gnd 0.008228f
C3963 vdd.n1715 gnd 0.008228f
C3964 vdd.n1716 gnd 0.008228f
C3965 vdd.n1717 gnd 0.010223f
C3966 vdd.n1718 gnd 0.010223f
C3967 vdd.n1719 gnd 0.010223f
C3968 vdd.n1720 gnd 0.008228f
C3969 vdd.n1721 gnd 0.008228f
C3970 vdd.n1722 gnd 0.008228f
C3971 vdd.n1723 gnd 0.010223f
C3972 vdd.n1724 gnd 0.010223f
C3973 vdd.n1725 gnd 0.010223f
C3974 vdd.n1726 gnd 0.008228f
C3975 vdd.n1727 gnd 0.008228f
C3976 vdd.n1728 gnd 0.008228f
C3977 vdd.n1729 gnd 0.010223f
C3978 vdd.n1730 gnd 0.010223f
C3979 vdd.n1731 gnd 0.010223f
C3980 vdd.n1732 gnd 0.008228f
C3981 vdd.n1733 gnd 0.006829f
C3982 vdd.n1734 gnd 0.023438f
C3983 vdd.n1736 gnd 2.30878f
C3984 vdd.n1737 gnd 0.023438f
C3985 vdd.n1738 gnd 0.003908f
C3986 vdd.n1739 gnd 0.023438f
C3987 vdd.n1740 gnd 0.023279f
C3988 vdd.n1741 gnd 0.010223f
C3989 vdd.n1742 gnd 0.008228f
C3990 vdd.n1743 gnd 0.010223f
C3991 vdd.t42 gnd 0.522348f
C3992 vdd.n1744 gnd 0.684276f
C3993 vdd.n1745 gnd 0.010223f
C3994 vdd.n1746 gnd 0.008228f
C3995 vdd.n1747 gnd 0.010223f
C3996 vdd.n1748 gnd 0.010223f
C3997 vdd.n1749 gnd 0.010223f
C3998 vdd.n1750 gnd 0.008228f
C3999 vdd.n1751 gnd 0.010223f
C4000 vdd.n1752 gnd 1.0447f
C4001 vdd.n1753 gnd 0.010223f
C4002 vdd.n1754 gnd 0.008228f
C4003 vdd.n1755 gnd 0.010223f
C4004 vdd.n1756 gnd 0.010223f
C4005 vdd.n1757 gnd 0.010223f
C4006 vdd.n1758 gnd 0.008228f
C4007 vdd.n1759 gnd 0.010223f
C4008 vdd.n1760 gnd 0.867098f
C4009 vdd.t119 gnd 0.522348f
C4010 vdd.n1761 gnd 0.6007f
C4011 vdd.n1762 gnd 0.010223f
C4012 vdd.n1763 gnd 0.008228f
C4013 vdd.n1764 gnd 0.010223f
C4014 vdd.n1765 gnd 0.010223f
C4015 vdd.n1766 gnd 0.010223f
C4016 vdd.n1767 gnd 0.008228f
C4017 vdd.n1768 gnd 0.010223f
C4018 vdd.n1769 gnd 0.621594f
C4019 vdd.n1770 gnd 0.010223f
C4020 vdd.n1771 gnd 0.008228f
C4021 vdd.n1772 gnd 0.010223f
C4022 vdd.n1773 gnd 0.010223f
C4023 vdd.n1774 gnd 0.010223f
C4024 vdd.n1775 gnd 0.008228f
C4025 vdd.n1776 gnd 0.010223f
C4026 vdd.n1777 gnd 0.590253f
C4027 vdd.n1778 gnd 0.799192f
C4028 vdd.n1779 gnd 0.010223f
C4029 vdd.n1780 gnd 0.008228f
C4030 vdd.n1781 gnd 0.010223f
C4031 vdd.n1782 gnd 0.010223f
C4032 vdd.n1783 gnd 0.010223f
C4033 vdd.n1784 gnd 0.008228f
C4034 vdd.n1785 gnd 0.010223f
C4035 vdd.n1786 gnd 0.867098f
C4036 vdd.n1787 gnd 0.010223f
C4037 vdd.n1788 gnd 0.008228f
C4038 vdd.n1789 gnd 0.010223f
C4039 vdd.n1790 gnd 0.010223f
C4040 vdd.n1791 gnd 0.010223f
C4041 vdd.n1792 gnd 0.008228f
C4042 vdd.n1793 gnd 0.010223f
C4043 vdd.t193 gnd 0.522348f
C4044 vdd.n1794 gnd 0.757405f
C4045 vdd.n1795 gnd 0.010223f
C4046 vdd.n1796 gnd 0.008228f
C4047 vdd.n1797 gnd 0.010223f
C4048 vdd.n1798 gnd 0.010223f
C4049 vdd.n1799 gnd 0.010223f
C4050 vdd.n1800 gnd 0.008228f
C4051 vdd.n1801 gnd 0.010223f
C4052 vdd.n1802 gnd 0.579806f
C4053 vdd.n1803 gnd 0.010223f
C4054 vdd.n1804 gnd 0.008228f
C4055 vdd.n1805 gnd 0.010223f
C4056 vdd.n1806 gnd 0.010223f
C4057 vdd.n1807 gnd 0.010223f
C4058 vdd.n1808 gnd 0.008228f
C4059 vdd.n1809 gnd 0.010223f
C4060 vdd.n1810 gnd 0.746958f
C4061 vdd.n1811 gnd 0.642488f
C4062 vdd.n1812 gnd 0.010223f
C4063 vdd.n1813 gnd 0.008228f
C4064 vdd.n1814 gnd 0.007857f
C4065 vdd.n1815 gnd 0.00561f
C4066 vdd.n1816 gnd 0.005206f
C4067 vdd.n1817 gnd 0.00288f
C4068 vdd.n1818 gnd 0.006612f
C4069 vdd.n1819 gnd 0.002797f
C4070 vdd.n1820 gnd 0.002962f
C4071 vdd.n1821 gnd 0.005206f
C4072 vdd.n1822 gnd 0.002797f
C4073 vdd.n1823 gnd 0.006612f
C4074 vdd.n1824 gnd 0.002962f
C4075 vdd.n1825 gnd 0.005206f
C4076 vdd.n1826 gnd 0.002797f
C4077 vdd.n1827 gnd 0.004959f
C4078 vdd.n1828 gnd 0.004974f
C4079 vdd.t155 gnd 0.014206f
C4080 vdd.n1829 gnd 0.031608f
C4081 vdd.n1830 gnd 0.164495f
C4082 vdd.n1831 gnd 0.002797f
C4083 vdd.n1832 gnd 0.002962f
C4084 vdd.n1833 gnd 0.006612f
C4085 vdd.n1834 gnd 0.006612f
C4086 vdd.n1835 gnd 0.002962f
C4087 vdd.n1836 gnd 0.002797f
C4088 vdd.n1837 gnd 0.005206f
C4089 vdd.n1838 gnd 0.005206f
C4090 vdd.n1839 gnd 0.002797f
C4091 vdd.n1840 gnd 0.002962f
C4092 vdd.n1841 gnd 0.006612f
C4093 vdd.n1842 gnd 0.006612f
C4094 vdd.n1843 gnd 0.002962f
C4095 vdd.n1844 gnd 0.002797f
C4096 vdd.n1845 gnd 0.005206f
C4097 vdd.n1846 gnd 0.005206f
C4098 vdd.n1847 gnd 0.002797f
C4099 vdd.n1848 gnd 0.002962f
C4100 vdd.n1849 gnd 0.006612f
C4101 vdd.n1850 gnd 0.006612f
C4102 vdd.n1851 gnd 0.015633f
C4103 vdd.n1852 gnd 0.00288f
C4104 vdd.n1853 gnd 0.002797f
C4105 vdd.n1854 gnd 0.013456f
C4106 vdd.n1855 gnd 0.009394f
C4107 vdd.t179 gnd 0.032912f
C4108 vdd.t225 gnd 0.032912f
C4109 vdd.n1856 gnd 0.226192f
C4110 vdd.n1857 gnd 0.177865f
C4111 vdd.t197 gnd 0.032912f
C4112 vdd.t235 gnd 0.032912f
C4113 vdd.n1858 gnd 0.226192f
C4114 vdd.n1859 gnd 0.143536f
C4115 vdd.t170 gnd 0.032912f
C4116 vdd.t126 gnd 0.032912f
C4117 vdd.n1860 gnd 0.226192f
C4118 vdd.n1861 gnd 0.143536f
C4119 vdd.t188 gnd 0.032912f
C4120 vdd.t132 gnd 0.032912f
C4121 vdd.n1862 gnd 0.226192f
C4122 vdd.n1863 gnd 0.143536f
C4123 vdd.t228 gnd 0.032912f
C4124 vdd.t239 gnd 0.032912f
C4125 vdd.n1864 gnd 0.226192f
C4126 vdd.n1865 gnd 0.143536f
C4127 vdd.t207 gnd 0.032912f
C4128 vdd.t138 gnd 0.032912f
C4129 vdd.n1866 gnd 0.226192f
C4130 vdd.n1867 gnd 0.143536f
C4131 vdd.t192 gnd 0.032912f
C4132 vdd.t150 gnd 0.032912f
C4133 vdd.n1868 gnd 0.226192f
C4134 vdd.n1869 gnd 0.143536f
C4135 vdd.n1870 gnd 0.00561f
C4136 vdd.n1871 gnd 0.005206f
C4137 vdd.n1872 gnd 0.00288f
C4138 vdd.n1873 gnd 0.006612f
C4139 vdd.n1874 gnd 0.002797f
C4140 vdd.n1875 gnd 0.002962f
C4141 vdd.n1876 gnd 0.005206f
C4142 vdd.n1877 gnd 0.002797f
C4143 vdd.n1878 gnd 0.006612f
C4144 vdd.n1879 gnd 0.002962f
C4145 vdd.n1880 gnd 0.005206f
C4146 vdd.n1881 gnd 0.002797f
C4147 vdd.n1882 gnd 0.004959f
C4148 vdd.n1883 gnd 0.004974f
C4149 vdd.t173 gnd 0.014206f
C4150 vdd.n1884 gnd 0.031608f
C4151 vdd.n1885 gnd 0.164495f
C4152 vdd.n1886 gnd 0.002797f
C4153 vdd.n1887 gnd 0.002962f
C4154 vdd.n1888 gnd 0.006612f
C4155 vdd.n1889 gnd 0.006612f
C4156 vdd.n1890 gnd 0.002962f
C4157 vdd.n1891 gnd 0.002797f
C4158 vdd.n1892 gnd 0.005206f
C4159 vdd.n1893 gnd 0.005206f
C4160 vdd.n1894 gnd 0.002797f
C4161 vdd.n1895 gnd 0.002962f
C4162 vdd.n1896 gnd 0.006612f
C4163 vdd.n1897 gnd 0.006612f
C4164 vdd.n1898 gnd 0.002962f
C4165 vdd.n1899 gnd 0.002797f
C4166 vdd.n1900 gnd 0.005206f
C4167 vdd.n1901 gnd 0.005206f
C4168 vdd.n1902 gnd 0.002797f
C4169 vdd.n1903 gnd 0.002962f
C4170 vdd.n1904 gnd 0.006612f
C4171 vdd.n1905 gnd 0.006612f
C4172 vdd.n1906 gnd 0.015633f
C4173 vdd.n1907 gnd 0.00288f
C4174 vdd.n1908 gnd 0.002797f
C4175 vdd.n1909 gnd 0.013456f
C4176 vdd.n1910 gnd 0.0091f
C4177 vdd.n1911 gnd 0.106792f
C4178 vdd.n1912 gnd 0.00561f
C4179 vdd.n1913 gnd 0.005206f
C4180 vdd.n1914 gnd 0.00288f
C4181 vdd.n1915 gnd 0.006612f
C4182 vdd.n1916 gnd 0.002797f
C4183 vdd.n1917 gnd 0.002962f
C4184 vdd.n1918 gnd 0.005206f
C4185 vdd.n1919 gnd 0.002797f
C4186 vdd.n1920 gnd 0.006612f
C4187 vdd.n1921 gnd 0.002962f
C4188 vdd.n1922 gnd 0.005206f
C4189 vdd.n1923 gnd 0.002797f
C4190 vdd.n1924 gnd 0.004959f
C4191 vdd.n1925 gnd 0.004974f
C4192 vdd.t221 gnd 0.014206f
C4193 vdd.n1926 gnd 0.031608f
C4194 vdd.n1927 gnd 0.164495f
C4195 vdd.n1928 gnd 0.002797f
C4196 vdd.n1929 gnd 0.002962f
C4197 vdd.n1930 gnd 0.006612f
C4198 vdd.n1931 gnd 0.006612f
C4199 vdd.n1932 gnd 0.002962f
C4200 vdd.n1933 gnd 0.002797f
C4201 vdd.n1934 gnd 0.005206f
C4202 vdd.n1935 gnd 0.005206f
C4203 vdd.n1936 gnd 0.002797f
C4204 vdd.n1937 gnd 0.002962f
C4205 vdd.n1938 gnd 0.006612f
C4206 vdd.n1939 gnd 0.006612f
C4207 vdd.n1940 gnd 0.002962f
C4208 vdd.n1941 gnd 0.002797f
C4209 vdd.n1942 gnd 0.005206f
C4210 vdd.n1943 gnd 0.005206f
C4211 vdd.n1944 gnd 0.002797f
C4212 vdd.n1945 gnd 0.002962f
C4213 vdd.n1946 gnd 0.006612f
C4214 vdd.n1947 gnd 0.006612f
C4215 vdd.n1948 gnd 0.015633f
C4216 vdd.n1949 gnd 0.00288f
C4217 vdd.n1950 gnd 0.002797f
C4218 vdd.n1951 gnd 0.013456f
C4219 vdd.n1952 gnd 0.009394f
C4220 vdd.t183 gnd 0.032912f
C4221 vdd.t118 gnd 0.032912f
C4222 vdd.n1953 gnd 0.226192f
C4223 vdd.n1954 gnd 0.177865f
C4224 vdd.t232 gnd 0.032912f
C4225 vdd.t209 gnd 0.032912f
C4226 vdd.n1955 gnd 0.226192f
C4227 vdd.n1956 gnd 0.143536f
C4228 vdd.t203 gnd 0.032912f
C4229 vdd.t156 gnd 0.032912f
C4230 vdd.n1957 gnd 0.226192f
C4231 vdd.n1958 gnd 0.143536f
C4232 vdd.t145 gnd 0.032912f
C4233 vdd.t204 gnd 0.032912f
C4234 vdd.n1959 gnd 0.226192f
C4235 vdd.n1960 gnd 0.143536f
C4236 vdd.t194 gnd 0.032912f
C4237 vdd.t191 gnd 0.032912f
C4238 vdd.n1961 gnd 0.226192f
C4239 vdd.n1962 gnd 0.143536f
C4240 vdd.t148 gnd 0.032912f
C4241 vdd.t124 gnd 0.032912f
C4242 vdd.n1963 gnd 0.226192f
C4243 vdd.n1964 gnd 0.143536f
C4244 vdd.t116 gnd 0.032912f
C4245 vdd.t189 gnd 0.032912f
C4246 vdd.n1965 gnd 0.226192f
C4247 vdd.n1966 gnd 0.143536f
C4248 vdd.n1967 gnd 0.00561f
C4249 vdd.n1968 gnd 0.005206f
C4250 vdd.n1969 gnd 0.00288f
C4251 vdd.n1970 gnd 0.006612f
C4252 vdd.n1971 gnd 0.002797f
C4253 vdd.n1972 gnd 0.002962f
C4254 vdd.n1973 gnd 0.005206f
C4255 vdd.n1974 gnd 0.002797f
C4256 vdd.n1975 gnd 0.006612f
C4257 vdd.n1976 gnd 0.002962f
C4258 vdd.n1977 gnd 0.005206f
C4259 vdd.n1978 gnd 0.002797f
C4260 vdd.n1979 gnd 0.004959f
C4261 vdd.n1980 gnd 0.004974f
C4262 vdd.t120 gnd 0.014206f
C4263 vdd.n1981 gnd 0.031608f
C4264 vdd.n1982 gnd 0.164495f
C4265 vdd.n1983 gnd 0.002797f
C4266 vdd.n1984 gnd 0.002962f
C4267 vdd.n1985 gnd 0.006612f
C4268 vdd.n1986 gnd 0.006612f
C4269 vdd.n1987 gnd 0.002962f
C4270 vdd.n1988 gnd 0.002797f
C4271 vdd.n1989 gnd 0.005206f
C4272 vdd.n1990 gnd 0.005206f
C4273 vdd.n1991 gnd 0.002797f
C4274 vdd.n1992 gnd 0.002962f
C4275 vdd.n1993 gnd 0.006612f
C4276 vdd.n1994 gnd 0.006612f
C4277 vdd.n1995 gnd 0.002962f
C4278 vdd.n1996 gnd 0.002797f
C4279 vdd.n1997 gnd 0.005206f
C4280 vdd.n1998 gnd 0.005206f
C4281 vdd.n1999 gnd 0.002797f
C4282 vdd.n2000 gnd 0.002962f
C4283 vdd.n2001 gnd 0.006612f
C4284 vdd.n2002 gnd 0.006612f
C4285 vdd.n2003 gnd 0.015633f
C4286 vdd.n2004 gnd 0.00288f
C4287 vdd.n2005 gnd 0.002797f
C4288 vdd.n2006 gnd 0.013456f
C4289 vdd.n2007 gnd 0.0091f
C4290 vdd.n2008 gnd 0.06353f
C4291 vdd.n2009 gnd 0.228916f
C4292 vdd.n2010 gnd 0.00561f
C4293 vdd.n2011 gnd 0.005206f
C4294 vdd.n2012 gnd 0.00288f
C4295 vdd.n2013 gnd 0.006612f
C4296 vdd.n2014 gnd 0.002797f
C4297 vdd.n2015 gnd 0.002962f
C4298 vdd.n2016 gnd 0.005206f
C4299 vdd.n2017 gnd 0.002797f
C4300 vdd.n2018 gnd 0.006612f
C4301 vdd.n2019 gnd 0.002962f
C4302 vdd.n2020 gnd 0.005206f
C4303 vdd.n2021 gnd 0.002797f
C4304 vdd.n2022 gnd 0.004959f
C4305 vdd.n2023 gnd 0.004974f
C4306 vdd.t231 gnd 0.014206f
C4307 vdd.n2024 gnd 0.031608f
C4308 vdd.n2025 gnd 0.164495f
C4309 vdd.n2026 gnd 0.002797f
C4310 vdd.n2027 gnd 0.002962f
C4311 vdd.n2028 gnd 0.006612f
C4312 vdd.n2029 gnd 0.006612f
C4313 vdd.n2030 gnd 0.002962f
C4314 vdd.n2031 gnd 0.002797f
C4315 vdd.n2032 gnd 0.005206f
C4316 vdd.n2033 gnd 0.005206f
C4317 vdd.n2034 gnd 0.002797f
C4318 vdd.n2035 gnd 0.002962f
C4319 vdd.n2036 gnd 0.006612f
C4320 vdd.n2037 gnd 0.006612f
C4321 vdd.n2038 gnd 0.002962f
C4322 vdd.n2039 gnd 0.002797f
C4323 vdd.n2040 gnd 0.005206f
C4324 vdd.n2041 gnd 0.005206f
C4325 vdd.n2042 gnd 0.002797f
C4326 vdd.n2043 gnd 0.002962f
C4327 vdd.n2044 gnd 0.006612f
C4328 vdd.n2045 gnd 0.006612f
C4329 vdd.n2046 gnd 0.015633f
C4330 vdd.n2047 gnd 0.00288f
C4331 vdd.n2048 gnd 0.002797f
C4332 vdd.n2049 gnd 0.013456f
C4333 vdd.n2050 gnd 0.009394f
C4334 vdd.t195 gnd 0.032912f
C4335 vdd.t140 gnd 0.032912f
C4336 vdd.n2051 gnd 0.226192f
C4337 vdd.n2052 gnd 0.177865f
C4338 vdd.t240 gnd 0.032912f
C4339 vdd.t216 gnd 0.032912f
C4340 vdd.n2053 gnd 0.226192f
C4341 vdd.n2054 gnd 0.143536f
C4342 vdd.t214 gnd 0.032912f
C4343 vdd.t174 gnd 0.032912f
C4344 vdd.n2055 gnd 0.226192f
C4345 vdd.n2056 gnd 0.143536f
C4346 vdd.t167 gnd 0.032912f
C4347 vdd.t215 gnd 0.032912f
C4348 vdd.n2057 gnd 0.226192f
C4349 vdd.n2058 gnd 0.143536f
C4350 vdd.t202 gnd 0.032912f
C4351 vdd.t201 gnd 0.032912f
C4352 vdd.n2059 gnd 0.226192f
C4353 vdd.n2060 gnd 0.143536f
C4354 vdd.t166 gnd 0.032912f
C4355 vdd.t142 gnd 0.032912f
C4356 vdd.n2061 gnd 0.226192f
C4357 vdd.n2062 gnd 0.143536f
C4358 vdd.t139 gnd 0.032912f
C4359 vdd.t200 gnd 0.032912f
C4360 vdd.n2063 gnd 0.226192f
C4361 vdd.n2064 gnd 0.143536f
C4362 vdd.n2065 gnd 0.00561f
C4363 vdd.n2066 gnd 0.005206f
C4364 vdd.n2067 gnd 0.00288f
C4365 vdd.n2068 gnd 0.006612f
C4366 vdd.n2069 gnd 0.002797f
C4367 vdd.n2070 gnd 0.002962f
C4368 vdd.n2071 gnd 0.005206f
C4369 vdd.n2072 gnd 0.002797f
C4370 vdd.n2073 gnd 0.006612f
C4371 vdd.n2074 gnd 0.002962f
C4372 vdd.n2075 gnd 0.005206f
C4373 vdd.n2076 gnd 0.002797f
C4374 vdd.n2077 gnd 0.004959f
C4375 vdd.n2078 gnd 0.004974f
C4376 vdd.t141 gnd 0.014206f
C4377 vdd.n2079 gnd 0.031608f
C4378 vdd.n2080 gnd 0.164495f
C4379 vdd.n2081 gnd 0.002797f
C4380 vdd.n2082 gnd 0.002962f
C4381 vdd.n2083 gnd 0.006612f
C4382 vdd.n2084 gnd 0.006612f
C4383 vdd.n2085 gnd 0.002962f
C4384 vdd.n2086 gnd 0.002797f
C4385 vdd.n2087 gnd 0.005206f
C4386 vdd.n2088 gnd 0.005206f
C4387 vdd.n2089 gnd 0.002797f
C4388 vdd.n2090 gnd 0.002962f
C4389 vdd.n2091 gnd 0.006612f
C4390 vdd.n2092 gnd 0.006612f
C4391 vdd.n2093 gnd 0.002962f
C4392 vdd.n2094 gnd 0.002797f
C4393 vdd.n2095 gnd 0.005206f
C4394 vdd.n2096 gnd 0.005206f
C4395 vdd.n2097 gnd 0.002797f
C4396 vdd.n2098 gnd 0.002962f
C4397 vdd.n2099 gnd 0.006612f
C4398 vdd.n2100 gnd 0.006612f
C4399 vdd.n2101 gnd 0.015633f
C4400 vdd.n2102 gnd 0.00288f
C4401 vdd.n2103 gnd 0.002797f
C4402 vdd.n2104 gnd 0.013456f
C4403 vdd.n2105 gnd 0.0091f
C4404 vdd.n2106 gnd 0.06353f
C4405 vdd.n2107 gnd 0.256355f
C4406 vdd.n2108 gnd 2.56885f
C4407 vdd.n2109 gnd 0.602965f
C4408 vdd.n2110 gnd 0.007857f
C4409 vdd.n2111 gnd 0.010223f
C4410 vdd.n2112 gnd 0.008228f
C4411 vdd.n2113 gnd 0.010223f
C4412 vdd.n2114 gnd 0.820086f
C4413 vdd.n2115 gnd 0.010223f
C4414 vdd.n2116 gnd 0.008228f
C4415 vdd.n2117 gnd 0.010223f
C4416 vdd.n2118 gnd 0.010223f
C4417 vdd.n2119 gnd 0.010223f
C4418 vdd.n2120 gnd 0.008228f
C4419 vdd.n2121 gnd 0.010223f
C4420 vdd.t125 gnd 0.522348f
C4421 vdd.n2122 gnd 0.867098f
C4422 vdd.n2123 gnd 0.010223f
C4423 vdd.n2124 gnd 0.008228f
C4424 vdd.n2125 gnd 0.010223f
C4425 vdd.n2126 gnd 0.010223f
C4426 vdd.n2127 gnd 0.010223f
C4427 vdd.n2128 gnd 0.008228f
C4428 vdd.n2129 gnd 0.010223f
C4429 vdd.n2130 gnd 0.736511f
C4430 vdd.n2131 gnd 0.010223f
C4431 vdd.n2132 gnd 0.008228f
C4432 vdd.n2133 gnd 0.010223f
C4433 vdd.n2134 gnd 0.010223f
C4434 vdd.n2135 gnd 0.010223f
C4435 vdd.n2136 gnd 0.008228f
C4436 vdd.n2137 gnd 0.010223f
C4437 vdd.n2138 gnd 0.867098f
C4438 vdd.t208 gnd 0.522348f
C4439 vdd.n2139 gnd 0.558912f
C4440 vdd.n2140 gnd 0.010223f
C4441 vdd.n2141 gnd 0.008228f
C4442 vdd.n2142 gnd 0.010223f
C4443 vdd.n2143 gnd 0.010223f
C4444 vdd.n2144 gnd 0.010223f
C4445 vdd.n2145 gnd 0.008228f
C4446 vdd.n2146 gnd 0.010223f
C4447 vdd.n2147 gnd 0.663382f
C4448 vdd.n2148 gnd 0.010223f
C4449 vdd.n2149 gnd 0.008228f
C4450 vdd.n2150 gnd 0.010223f
C4451 vdd.n2151 gnd 0.010223f
C4452 vdd.n2152 gnd 0.010223f
C4453 vdd.n2153 gnd 0.008228f
C4454 vdd.n2154 gnd 0.010223f
C4455 vdd.n2155 gnd 0.548465f
C4456 vdd.n2156 gnd 0.84098f
C4457 vdd.n2157 gnd 0.010223f
C4458 vdd.n2158 gnd 0.008228f
C4459 vdd.n2159 gnd 0.010223f
C4460 vdd.n2160 gnd 0.010223f
C4461 vdd.n2161 gnd 0.010223f
C4462 vdd.n2162 gnd 0.008228f
C4463 vdd.n2163 gnd 0.010223f
C4464 vdd.n2164 gnd 1.01858f
C4465 vdd.n2165 gnd 0.010223f
C4466 vdd.n2166 gnd 0.008228f
C4467 vdd.n2167 gnd 0.010223f
C4468 vdd.n2168 gnd 0.010223f
C4469 vdd.n2169 gnd 0.023279f
C4470 vdd.n2170 gnd 0.010223f
C4471 vdd.n2171 gnd 0.010223f
C4472 vdd.n2172 gnd 0.008228f
C4473 vdd.n2173 gnd 0.010223f
C4474 vdd.t25 gnd 0.522348f
C4475 vdd.n2174 gnd 0.987238f
C4476 vdd.n2175 gnd 0.010223f
C4477 vdd.n2176 gnd 0.008228f
C4478 vdd.n2177 gnd 0.010223f
C4479 vdd.n2178 gnd 0.010223f
C4480 vdd.n2179 gnd 0.023279f
C4481 vdd.n2180 gnd 0.006829f
C4482 vdd.n2181 gnd 0.023279f
C4483 vdd.n2182 gnd 1.379f
C4484 vdd.n2183 gnd 0.023279f
C4485 vdd.n2184 gnd 0.023438f
C4486 vdd.n2185 gnd 0.003908f
C4487 vdd.t27 gnd 0.125764f
C4488 vdd.t26 gnd 0.134407f
C4489 vdd.t24 gnd 0.164246f
C4490 vdd.n2186 gnd 0.210541f
C4491 vdd.n2187 gnd 0.176892f
C4492 vdd.n2188 gnd 0.012671f
C4493 vdd.n2189 gnd 0.00432f
C4494 vdd.n2190 gnd 0.008791f
C4495 vdd.n2191 gnd 0.773084f
C4496 vdd.n2193 gnd 0.008228f
C4497 vdd.n2194 gnd 0.008228f
C4498 vdd.n2195 gnd 0.010223f
C4499 vdd.n2197 gnd 0.010223f
C4500 vdd.n2198 gnd 0.010223f
C4501 vdd.n2199 gnd 0.008228f
C4502 vdd.n2200 gnd 0.008228f
C4503 vdd.n2201 gnd 0.008228f
C4504 vdd.n2202 gnd 0.010223f
C4505 vdd.n2204 gnd 0.010223f
C4506 vdd.n2205 gnd 0.010223f
C4507 vdd.n2206 gnd 0.008228f
C4508 vdd.n2207 gnd 0.008228f
C4509 vdd.n2208 gnd 0.008228f
C4510 vdd.n2209 gnd 0.010223f
C4511 vdd.n2211 gnd 0.010223f
C4512 vdd.n2212 gnd 0.010223f
C4513 vdd.n2213 gnd 0.008228f
C4514 vdd.n2214 gnd 0.008228f
C4515 vdd.n2215 gnd 0.008228f
C4516 vdd.n2216 gnd 0.010223f
C4517 vdd.n2218 gnd 0.010223f
C4518 vdd.n2219 gnd 0.010223f
C4519 vdd.n2220 gnd 0.008228f
C4520 vdd.n2221 gnd 0.010223f
C4521 vdd.n2222 gnd 0.010223f
C4522 vdd.n2223 gnd 0.010223f
C4523 vdd.n2224 gnd 0.016785f
C4524 vdd.n2225 gnd 0.005595f
C4525 vdd.n2226 gnd 0.008228f
C4526 vdd.n2227 gnd 0.010223f
C4527 vdd.n2229 gnd 0.010223f
C4528 vdd.n2230 gnd 0.010223f
C4529 vdd.n2231 gnd 0.008228f
C4530 vdd.n2232 gnd 0.008228f
C4531 vdd.n2233 gnd 0.008228f
C4532 vdd.n2234 gnd 0.010223f
C4533 vdd.n2236 gnd 0.010223f
C4534 vdd.n2237 gnd 0.010223f
C4535 vdd.n2238 gnd 0.008228f
C4536 vdd.n2239 gnd 0.008228f
C4537 vdd.n2240 gnd 0.008228f
C4538 vdd.n2241 gnd 0.010223f
C4539 vdd.n2243 gnd 0.010223f
C4540 vdd.n2244 gnd 0.010223f
C4541 vdd.n2245 gnd 0.008228f
C4542 vdd.n2246 gnd 0.008228f
C4543 vdd.n2247 gnd 0.008228f
C4544 vdd.n2248 gnd 0.010223f
C4545 vdd.n2250 gnd 0.010223f
C4546 vdd.n2251 gnd 0.010223f
C4547 vdd.n2252 gnd 0.008228f
C4548 vdd.n2253 gnd 0.008228f
C4549 vdd.n2254 gnd 0.008228f
C4550 vdd.n2255 gnd 0.010223f
C4551 vdd.n2257 gnd 0.010223f
C4552 vdd.n2258 gnd 0.010223f
C4553 vdd.n2259 gnd 0.008228f
C4554 vdd.n2260 gnd 0.010223f
C4555 vdd.n2261 gnd 0.010223f
C4556 vdd.n2262 gnd 0.010223f
C4557 vdd.n2263 gnd 0.016785f
C4558 vdd.n2264 gnd 0.00687f
C4559 vdd.n2265 gnd 0.008228f
C4560 vdd.n2266 gnd 0.010223f
C4561 vdd.n2268 gnd 0.010223f
C4562 vdd.n2269 gnd 0.010223f
C4563 vdd.n2270 gnd 0.008228f
C4564 vdd.n2271 gnd 0.008228f
C4565 vdd.n2272 gnd 0.008228f
C4566 vdd.n2273 gnd 0.010223f
C4567 vdd.n2275 gnd 0.010223f
C4568 vdd.n2276 gnd 0.010223f
C4569 vdd.n2277 gnd 0.008228f
C4570 vdd.n2278 gnd 0.008228f
C4571 vdd.n2279 gnd 0.008228f
C4572 vdd.n2280 gnd 0.010223f
C4573 vdd.n2282 gnd 0.010223f
C4574 vdd.n2283 gnd 0.010223f
C4575 vdd.n2284 gnd 0.008228f
C4576 vdd.n2285 gnd 0.008228f
C4577 vdd.n2286 gnd 0.008228f
C4578 vdd.n2287 gnd 0.010223f
C4579 vdd.n2289 gnd 0.010223f
C4580 vdd.n2290 gnd 0.008228f
C4581 vdd.n2291 gnd 0.008228f
C4582 vdd.n2292 gnd 0.010223f
C4583 vdd.n2294 gnd 0.010223f
C4584 vdd.n2295 gnd 0.010223f
C4585 vdd.n2296 gnd 0.008228f
C4586 vdd.n2297 gnd 0.008791f
C4587 vdd.n2298 gnd 0.773084f
C4588 vdd.n2299 gnd 0.027861f
C4589 vdd.n2300 gnd 0.006951f
C4590 vdd.n2301 gnd 0.006951f
C4591 vdd.n2302 gnd 0.006951f
C4592 vdd.n2303 gnd 0.006951f
C4593 vdd.n2304 gnd 0.006951f
C4594 vdd.n2305 gnd 0.006951f
C4595 vdd.n2306 gnd 0.006951f
C4596 vdd.n2307 gnd 0.006951f
C4597 vdd.n2308 gnd 0.006951f
C4598 vdd.n2309 gnd 0.006951f
C4599 vdd.n2310 gnd 0.006951f
C4600 vdd.n2311 gnd 0.006951f
C4601 vdd.n2312 gnd 0.006951f
C4602 vdd.n2313 gnd 0.006951f
C4603 vdd.n2314 gnd 0.006951f
C4604 vdd.n2315 gnd 0.006951f
C4605 vdd.n2316 gnd 0.006951f
C4606 vdd.n2317 gnd 0.006951f
C4607 vdd.n2318 gnd 0.006951f
C4608 vdd.n2319 gnd 0.006951f
C4609 vdd.n2320 gnd 0.006951f
C4610 vdd.n2321 gnd 0.006951f
C4611 vdd.n2322 gnd 0.006951f
C4612 vdd.n2323 gnd 0.006951f
C4613 vdd.n2324 gnd 0.006951f
C4614 vdd.n2325 gnd 0.006951f
C4615 vdd.n2326 gnd 0.006951f
C4616 vdd.n2327 gnd 0.006951f
C4617 vdd.n2328 gnd 0.006951f
C4618 vdd.n2329 gnd 0.006951f
C4619 vdd.n2330 gnd 0.006951f
C4620 vdd.n2331 gnd 0.016259f
C4621 vdd.n2332 gnd 0.016259f
C4622 vdd.n2334 gnd 8.91126f
C4623 vdd.n2336 gnd 0.016259f
C4624 vdd.n2337 gnd 0.016259f
C4625 vdd.n2338 gnd 0.015227f
C4626 vdd.n2339 gnd 0.006951f
C4627 vdd.n2340 gnd 0.006951f
C4628 vdd.n2341 gnd 0.710393f
C4629 vdd.n2342 gnd 0.006951f
C4630 vdd.n2343 gnd 0.006951f
C4631 vdd.n2344 gnd 0.006951f
C4632 vdd.n2345 gnd 0.006951f
C4633 vdd.n2346 gnd 0.006951f
C4634 vdd.n2347 gnd 0.6007f
C4635 vdd.n2348 gnd 0.006951f
C4636 vdd.n2349 gnd 0.006951f
C4637 vdd.n2350 gnd 0.006951f
C4638 vdd.n2351 gnd 0.006951f
C4639 vdd.n2352 gnd 0.006951f
C4640 vdd.n2353 gnd 0.710393f
C4641 vdd.n2354 gnd 0.006951f
C4642 vdd.n2355 gnd 0.006951f
C4643 vdd.n2356 gnd 0.006951f
C4644 vdd.n2357 gnd 0.006951f
C4645 vdd.n2358 gnd 0.006951f
C4646 vdd.n2359 gnd 0.694723f
C4647 vdd.n2360 gnd 0.006951f
C4648 vdd.n2361 gnd 0.006951f
C4649 vdd.n2362 gnd 0.006951f
C4650 vdd.n2363 gnd 0.006951f
C4651 vdd.n2364 gnd 0.006951f
C4652 vdd.n2365 gnd 0.710393f
C4653 vdd.n2366 gnd 0.006951f
C4654 vdd.n2367 gnd 0.006951f
C4655 vdd.n2368 gnd 0.006951f
C4656 vdd.n2369 gnd 0.006951f
C4657 vdd.n2370 gnd 0.006951f
C4658 vdd.n2371 gnd 0.569359f
C4659 vdd.n2372 gnd 0.006951f
C4660 vdd.n2373 gnd 0.006951f
C4661 vdd.n2374 gnd 0.005929f
C4662 vdd.n2375 gnd 0.020137f
C4663 vdd.n2376 gnd 0.004498f
C4664 vdd.n2377 gnd 0.006951f
C4665 vdd.n2378 gnd 0.412655f
C4666 vdd.n2379 gnd 0.006951f
C4667 vdd.n2380 gnd 0.006951f
C4668 vdd.n2381 gnd 0.006951f
C4669 vdd.n2382 gnd 0.006951f
C4670 vdd.n2383 gnd 0.006951f
C4671 vdd.n2384 gnd 0.454443f
C4672 vdd.n2385 gnd 0.006951f
C4673 vdd.n2386 gnd 0.006951f
C4674 vdd.n2387 gnd 0.006951f
C4675 vdd.n2388 gnd 0.006951f
C4676 vdd.n2389 gnd 0.006951f
C4677 vdd.n2390 gnd 0.611147f
C4678 vdd.n2391 gnd 0.006951f
C4679 vdd.n2392 gnd 0.006951f
C4680 vdd.n2393 gnd 0.006951f
C4681 vdd.n2394 gnd 0.006951f
C4682 vdd.n2395 gnd 0.006951f
C4683 vdd.n2396 gnd 0.58503f
C4684 vdd.n2397 gnd 0.006951f
C4685 vdd.n2398 gnd 0.006951f
C4686 vdd.n2399 gnd 0.006951f
C4687 vdd.n2400 gnd 0.006951f
C4688 vdd.n2401 gnd 0.006951f
C4689 vdd.n2402 gnd 0.428325f
C4690 vdd.n2403 gnd 0.006951f
C4691 vdd.n2404 gnd 0.006951f
C4692 vdd.n2405 gnd 0.006951f
C4693 vdd.n2406 gnd 0.006951f
C4694 vdd.n2407 gnd 0.006951f
C4695 vdd.n2408 gnd 0.22461f
C4696 vdd.n2409 gnd 0.006951f
C4697 vdd.n2410 gnd 0.006951f
C4698 vdd.n2411 gnd 0.006951f
C4699 vdd.n2412 gnd 0.006951f
C4700 vdd.n2413 gnd 0.006951f
C4701 vdd.n2414 gnd 0.370867f
C4702 vdd.n2415 gnd 0.006951f
C4703 vdd.n2416 gnd 0.006951f
C4704 vdd.n2417 gnd 0.006951f
C4705 vdd.n2418 gnd 0.006951f
C4706 vdd.n2419 gnd 0.006951f
C4707 vdd.n2420 gnd 0.710393f
C4708 vdd.n2421 gnd 0.006951f
C4709 vdd.n2422 gnd 0.006951f
C4710 vdd.n2423 gnd 0.006951f
C4711 vdd.n2424 gnd 0.006951f
C4712 vdd.n2425 gnd 0.006951f
C4713 vdd.n2426 gnd 0.006951f
C4714 vdd.n2427 gnd 0.006951f
C4715 vdd.n2428 gnd 0.532795f
C4716 vdd.n2429 gnd 0.006951f
C4717 vdd.n2430 gnd 0.006951f
C4718 vdd.n2431 gnd 0.006951f
C4719 vdd.n2432 gnd 0.006951f
C4720 vdd.n2433 gnd 0.006951f
C4721 vdd.n2434 gnd 0.006951f
C4722 vdd.n2435 gnd 0.443996f
C4723 vdd.n2436 gnd 0.006951f
C4724 vdd.n2437 gnd 0.006951f
C4725 vdd.n2438 gnd 0.006951f
C4726 vdd.n2439 gnd 0.01609f
C4727 vdd.n2440 gnd 0.015395f
C4728 vdd.n2441 gnd 0.006951f
C4729 vdd.n2442 gnd 0.006951f
C4730 vdd.n2443 gnd 0.005367f
C4731 vdd.n2444 gnd 0.006951f
C4732 vdd.n2445 gnd 0.006951f
C4733 vdd.n2446 gnd 0.00506f
C4734 vdd.n2447 gnd 0.006951f
C4735 vdd.n2448 gnd 0.006951f
C4736 vdd.n2449 gnd 0.006951f
C4737 vdd.n2450 gnd 0.006951f
C4738 vdd.n2451 gnd 0.006951f
C4739 vdd.n2452 gnd 0.006951f
C4740 vdd.n2453 gnd 0.006951f
C4741 vdd.n2454 gnd 0.006951f
C4742 vdd.n2455 gnd 0.006951f
C4743 vdd.n2456 gnd 0.006951f
C4744 vdd.n2457 gnd 0.006951f
C4745 vdd.n2458 gnd 0.006951f
C4746 vdd.n2459 gnd 0.006951f
C4747 vdd.n2460 gnd 0.006951f
C4748 vdd.n2461 gnd 0.006951f
C4749 vdd.n2462 gnd 0.006951f
C4750 vdd.n2463 gnd 0.006951f
C4751 vdd.n2464 gnd 0.006951f
C4752 vdd.n2465 gnd 0.006951f
C4753 vdd.n2466 gnd 0.006951f
C4754 vdd.n2467 gnd 0.006951f
C4755 vdd.n2468 gnd 0.006951f
C4756 vdd.n2469 gnd 0.006951f
C4757 vdd.n2470 gnd 0.006951f
C4758 vdd.n2471 gnd 0.006951f
C4759 vdd.n2472 gnd 0.006951f
C4760 vdd.n2473 gnd 0.006951f
C4761 vdd.n2474 gnd 0.006951f
C4762 vdd.n2475 gnd 0.006951f
C4763 vdd.n2476 gnd 0.006951f
C4764 vdd.n2477 gnd 0.006951f
C4765 vdd.n2478 gnd 0.006951f
C4766 vdd.n2479 gnd 0.006951f
C4767 vdd.n2480 gnd 0.006951f
C4768 vdd.n2481 gnd 0.006951f
C4769 vdd.n2482 gnd 0.006951f
C4770 vdd.n2483 gnd 0.006951f
C4771 vdd.n2484 gnd 0.006951f
C4772 vdd.n2485 gnd 0.006951f
C4773 vdd.n2486 gnd 0.006951f
C4774 vdd.n2487 gnd 0.006951f
C4775 vdd.n2488 gnd 0.006951f
C4776 vdd.n2489 gnd 0.006951f
C4777 vdd.n2490 gnd 0.006951f
C4778 vdd.n2491 gnd 0.006951f
C4779 vdd.n2492 gnd 0.006951f
C4780 vdd.n2493 gnd 0.006951f
C4781 vdd.n2494 gnd 0.006951f
C4782 vdd.n2495 gnd 0.006951f
C4783 vdd.n2496 gnd 0.006951f
C4784 vdd.n2497 gnd 0.006951f
C4785 vdd.n2498 gnd 0.006951f
C4786 vdd.n2499 gnd 0.006951f
C4787 vdd.n2500 gnd 0.006951f
C4788 vdd.n2501 gnd 0.006951f
C4789 vdd.n2502 gnd 0.006951f
C4790 vdd.n2503 gnd 0.006951f
C4791 vdd.n2504 gnd 0.006951f
C4792 vdd.n2505 gnd 0.006951f
C4793 vdd.n2506 gnd 0.006951f
C4794 vdd.n2507 gnd 0.016259f
C4795 vdd.n2508 gnd 0.015227f
C4796 vdd.n2509 gnd 0.015227f
C4797 vdd.n2510 gnd 0.846204f
C4798 vdd.n2511 gnd 0.015227f
C4799 vdd.n2512 gnd 0.016259f
C4800 vdd.n2513 gnd 0.015395f
C4801 vdd.n2514 gnd 0.006951f
C4802 vdd.n2515 gnd 0.006951f
C4803 vdd.n2516 gnd 0.006951f
C4804 vdd.n2517 gnd 0.005367f
C4805 vdd.n2518 gnd 0.009935f
C4806 vdd.n2519 gnd 0.00506f
C4807 vdd.n2520 gnd 0.006951f
C4808 vdd.n2521 gnd 0.006951f
C4809 vdd.n2522 gnd 0.006951f
C4810 vdd.n2523 gnd 0.006951f
C4811 vdd.n2524 gnd 0.006951f
C4812 vdd.n2525 gnd 0.006951f
C4813 vdd.n2526 gnd 0.006951f
C4814 vdd.n2527 gnd 0.006951f
C4815 vdd.n2528 gnd 0.006951f
C4816 vdd.n2529 gnd 0.006951f
C4817 vdd.n2530 gnd 0.006951f
C4818 vdd.n2531 gnd 0.006951f
C4819 vdd.n2532 gnd 0.006951f
C4820 vdd.n2533 gnd 0.006951f
C4821 vdd.n2534 gnd 0.006951f
C4822 vdd.n2535 gnd 0.006951f
C4823 vdd.n2536 gnd 0.006951f
C4824 vdd.n2537 gnd 0.006951f
C4825 vdd.n2538 gnd 0.006951f
C4826 vdd.n2539 gnd 0.006951f
C4827 vdd.n2540 gnd 0.006951f
C4828 vdd.n2541 gnd 0.006951f
C4829 vdd.n2542 gnd 0.006951f
C4830 vdd.n2543 gnd 0.006951f
C4831 vdd.n2544 gnd 0.006951f
C4832 vdd.n2545 gnd 0.006951f
C4833 vdd.n2546 gnd 0.006951f
C4834 vdd.n2547 gnd 0.006951f
C4835 vdd.n2548 gnd 0.006951f
C4836 vdd.n2549 gnd 0.006951f
C4837 vdd.n2550 gnd 0.006951f
C4838 vdd.n2551 gnd 0.006951f
C4839 vdd.n2552 gnd 0.006951f
C4840 vdd.n2553 gnd 0.006951f
C4841 vdd.n2554 gnd 0.006951f
C4842 vdd.n2555 gnd 0.006951f
C4843 vdd.n2556 gnd 0.006951f
C4844 vdd.n2557 gnd 0.006951f
C4845 vdd.n2558 gnd 0.006951f
C4846 vdd.n2559 gnd 0.006951f
C4847 vdd.n2560 gnd 0.006951f
C4848 vdd.n2561 gnd 0.006951f
C4849 vdd.n2562 gnd 0.006951f
C4850 vdd.n2563 gnd 0.006951f
C4851 vdd.n2564 gnd 0.006951f
C4852 vdd.n2565 gnd 0.006951f
C4853 vdd.n2566 gnd 0.006951f
C4854 vdd.n2567 gnd 0.006951f
C4855 vdd.n2568 gnd 0.006951f
C4856 vdd.n2569 gnd 0.006951f
C4857 vdd.n2570 gnd 0.006951f
C4858 vdd.n2571 gnd 0.006951f
C4859 vdd.n2572 gnd 0.006951f
C4860 vdd.n2573 gnd 0.006951f
C4861 vdd.n2574 gnd 0.006951f
C4862 vdd.n2575 gnd 0.006951f
C4863 vdd.n2576 gnd 0.006951f
C4864 vdd.n2577 gnd 0.006951f
C4865 vdd.n2578 gnd 0.006951f
C4866 vdd.n2579 gnd 0.006951f
C4867 vdd.n2580 gnd 0.016259f
C4868 vdd.n2581 gnd 0.016259f
C4869 vdd.n2582 gnd 0.867098f
C4870 vdd.t258 gnd 3.08185f
C4871 vdd.t101 gnd 3.08185f
C4872 vdd.n2615 gnd 0.016259f
C4873 vdd.t247 gnd 0.647711f
C4874 vdd.n2616 gnd 0.006951f
C4875 vdd.n2617 gnd 0.006951f
C4876 vdd.t64 gnd 0.280902f
C4877 vdd.t65 gnd 0.287539f
C4878 vdd.t62 gnd 0.183384f
C4879 vdd.n2618 gnd 0.099109f
C4880 vdd.n2619 gnd 0.056218f
C4881 vdd.n2620 gnd 0.006951f
C4882 vdd.t74 gnd 0.280902f
C4883 vdd.t75 gnd 0.287539f
C4884 vdd.t73 gnd 0.183384f
C4885 vdd.n2621 gnd 0.099109f
C4886 vdd.n2622 gnd 0.056218f
C4887 vdd.n2623 gnd 0.009935f
C4888 vdd.n2624 gnd 0.006951f
C4889 vdd.n2625 gnd 0.006951f
C4890 vdd.n2626 gnd 0.006951f
C4891 vdd.n2627 gnd 0.006951f
C4892 vdd.n2628 gnd 0.006951f
C4893 vdd.n2629 gnd 0.006951f
C4894 vdd.n2630 gnd 0.006951f
C4895 vdd.n2631 gnd 0.006951f
C4896 vdd.n2632 gnd 0.006951f
C4897 vdd.n2633 gnd 0.006951f
C4898 vdd.n2634 gnd 0.006951f
C4899 vdd.n2635 gnd 0.006951f
C4900 vdd.n2636 gnd 0.006951f
C4901 vdd.n2637 gnd 0.006951f
C4902 vdd.n2638 gnd 0.006951f
C4903 vdd.n2639 gnd 0.006951f
C4904 vdd.n2640 gnd 0.006951f
C4905 vdd.n2641 gnd 0.006951f
C4906 vdd.n2642 gnd 0.006951f
C4907 vdd.n2643 gnd 0.006951f
C4908 vdd.n2644 gnd 0.006951f
C4909 vdd.n2645 gnd 0.006951f
C4910 vdd.n2646 gnd 0.006951f
C4911 vdd.n2647 gnd 0.006951f
C4912 vdd.n2648 gnd 0.006951f
C4913 vdd.n2649 gnd 0.006951f
C4914 vdd.n2650 gnd 0.006951f
C4915 vdd.n2651 gnd 0.006951f
C4916 vdd.n2652 gnd 0.006951f
C4917 vdd.n2653 gnd 0.006951f
C4918 vdd.n2654 gnd 0.006951f
C4919 vdd.n2655 gnd 0.006951f
C4920 vdd.n2656 gnd 0.006951f
C4921 vdd.n2657 gnd 0.006951f
C4922 vdd.n2658 gnd 0.006951f
C4923 vdd.n2659 gnd 0.006951f
C4924 vdd.n2660 gnd 0.006951f
C4925 vdd.n2661 gnd 0.006951f
C4926 vdd.n2662 gnd 0.006951f
C4927 vdd.n2663 gnd 0.006951f
C4928 vdd.n2664 gnd 0.006951f
C4929 vdd.n2665 gnd 0.006951f
C4930 vdd.n2666 gnd 0.006951f
C4931 vdd.n2667 gnd 0.006951f
C4932 vdd.n2668 gnd 0.006951f
C4933 vdd.n2669 gnd 0.006951f
C4934 vdd.n2670 gnd 0.006951f
C4935 vdd.n2671 gnd 0.006951f
C4936 vdd.n2672 gnd 0.006951f
C4937 vdd.n2673 gnd 0.006951f
C4938 vdd.n2674 gnd 0.006951f
C4939 vdd.n2675 gnd 0.006951f
C4940 vdd.n2676 gnd 0.006951f
C4941 vdd.n2677 gnd 0.006951f
C4942 vdd.n2678 gnd 0.006951f
C4943 vdd.n2679 gnd 0.006951f
C4944 vdd.n2680 gnd 0.006951f
C4945 vdd.n2681 gnd 0.006951f
C4946 vdd.n2682 gnd 0.00506f
C4947 vdd.n2683 gnd 0.006951f
C4948 vdd.n2684 gnd 0.006951f
C4949 vdd.n2685 gnd 0.005367f
C4950 vdd.n2686 gnd 0.006951f
C4951 vdd.n2687 gnd 0.006951f
C4952 vdd.n2688 gnd 0.016259f
C4953 vdd.n2689 gnd 0.015227f
C4954 vdd.n2690 gnd 0.015227f
C4955 vdd.n2691 gnd 0.006951f
C4956 vdd.n2692 gnd 0.006951f
C4957 vdd.n2693 gnd 0.006951f
C4958 vdd.n2694 gnd 0.006951f
C4959 vdd.n2695 gnd 0.006951f
C4960 vdd.n2696 gnd 0.006951f
C4961 vdd.n2697 gnd 0.006951f
C4962 vdd.n2698 gnd 0.006951f
C4963 vdd.n2699 gnd 0.006951f
C4964 vdd.n2700 gnd 0.006951f
C4965 vdd.n2701 gnd 0.006951f
C4966 vdd.n2702 gnd 0.006951f
C4967 vdd.n2703 gnd 0.006951f
C4968 vdd.n2704 gnd 0.006951f
C4969 vdd.n2705 gnd 0.006951f
C4970 vdd.n2706 gnd 0.006951f
C4971 vdd.n2707 gnd 0.006951f
C4972 vdd.n2708 gnd 0.006951f
C4973 vdd.n2709 gnd 0.006951f
C4974 vdd.n2710 gnd 0.006951f
C4975 vdd.n2711 gnd 0.006951f
C4976 vdd.n2712 gnd 0.006951f
C4977 vdd.n2713 gnd 0.006951f
C4978 vdd.n2714 gnd 0.006951f
C4979 vdd.n2715 gnd 0.006951f
C4980 vdd.n2716 gnd 0.006951f
C4981 vdd.n2717 gnd 0.006951f
C4982 vdd.n2718 gnd 0.006951f
C4983 vdd.n2719 gnd 0.006951f
C4984 vdd.n2720 gnd 0.006951f
C4985 vdd.n2721 gnd 0.006951f
C4986 vdd.n2722 gnd 0.006951f
C4987 vdd.n2723 gnd 0.006951f
C4988 vdd.n2724 gnd 0.006951f
C4989 vdd.n2725 gnd 0.006951f
C4990 vdd.n2726 gnd 0.006951f
C4991 vdd.n2727 gnd 0.006951f
C4992 vdd.n2728 gnd 0.006951f
C4993 vdd.n2729 gnd 0.006951f
C4994 vdd.n2730 gnd 0.006951f
C4995 vdd.n2731 gnd 0.006951f
C4996 vdd.n2732 gnd 0.006951f
C4997 vdd.n2733 gnd 0.006951f
C4998 vdd.n2734 gnd 0.006951f
C4999 vdd.n2735 gnd 0.006951f
C5000 vdd.n2736 gnd 0.006951f
C5001 vdd.n2737 gnd 0.006951f
C5002 vdd.n2738 gnd 0.006951f
C5003 vdd.n2739 gnd 0.006951f
C5004 vdd.n2740 gnd 0.006951f
C5005 vdd.n2741 gnd 0.006951f
C5006 vdd.n2742 gnd 0.006951f
C5007 vdd.n2743 gnd 0.006951f
C5008 vdd.n2744 gnd 0.006951f
C5009 vdd.n2745 gnd 0.006951f
C5010 vdd.n2746 gnd 0.006951f
C5011 vdd.n2747 gnd 0.006951f
C5012 vdd.n2748 gnd 0.006951f
C5013 vdd.n2749 gnd 0.006951f
C5014 vdd.n2750 gnd 0.006951f
C5015 vdd.n2751 gnd 0.006951f
C5016 vdd.n2752 gnd 0.006951f
C5017 vdd.n2753 gnd 0.006951f
C5018 vdd.n2754 gnd 0.006951f
C5019 vdd.n2755 gnd 0.006951f
C5020 vdd.n2756 gnd 0.006951f
C5021 vdd.n2757 gnd 0.006951f
C5022 vdd.n2758 gnd 0.006951f
C5023 vdd.n2759 gnd 0.006951f
C5024 vdd.n2760 gnd 0.006951f
C5025 vdd.n2761 gnd 0.006951f
C5026 vdd.n2762 gnd 0.006951f
C5027 vdd.n2763 gnd 0.006951f
C5028 vdd.n2764 gnd 0.22461f
C5029 vdd.n2765 gnd 0.006951f
C5030 vdd.n2766 gnd 0.006951f
C5031 vdd.n2767 gnd 0.006951f
C5032 vdd.n2768 gnd 0.006951f
C5033 vdd.n2769 gnd 0.006951f
C5034 vdd.n2770 gnd 0.006951f
C5035 vdd.n2771 gnd 0.006951f
C5036 vdd.n2772 gnd 0.006951f
C5037 vdd.n2773 gnd 0.006951f
C5038 vdd.n2774 gnd 0.006951f
C5039 vdd.n2775 gnd 0.006951f
C5040 vdd.n2776 gnd 0.006951f
C5041 vdd.n2777 gnd 0.006951f
C5042 vdd.n2778 gnd 0.006951f
C5043 vdd.n2779 gnd 0.443996f
C5044 vdd.n2780 gnd 0.006951f
C5045 vdd.n2781 gnd 0.006951f
C5046 vdd.n2782 gnd 0.006951f
C5047 vdd.n2783 gnd 0.015227f
C5048 vdd.n2784 gnd 0.015227f
C5049 vdd.n2785 gnd 0.016259f
C5050 vdd.n2786 gnd 0.016259f
C5051 vdd.n2787 gnd 0.006951f
C5052 vdd.n2788 gnd 0.006951f
C5053 vdd.n2789 gnd 0.006951f
C5054 vdd.n2790 gnd 0.005367f
C5055 vdd.n2791 gnd 0.009935f
C5056 vdd.n2792 gnd 0.00506f
C5057 vdd.n2793 gnd 0.006951f
C5058 vdd.n2794 gnd 0.006951f
C5059 vdd.n2795 gnd 0.006951f
C5060 vdd.n2796 gnd 0.006951f
C5061 vdd.n2797 gnd 0.006951f
C5062 vdd.n2798 gnd 0.006951f
C5063 vdd.n2799 gnd 0.006951f
C5064 vdd.n2800 gnd 0.006951f
C5065 vdd.n2801 gnd 0.006951f
C5066 vdd.n2802 gnd 0.006951f
C5067 vdd.n2803 gnd 0.006951f
C5068 vdd.n2804 gnd 0.006951f
C5069 vdd.n2805 gnd 0.006951f
C5070 vdd.n2806 gnd 0.006951f
C5071 vdd.n2807 gnd 0.006951f
C5072 vdd.n2808 gnd 0.006951f
C5073 vdd.n2809 gnd 0.006951f
C5074 vdd.n2810 gnd 0.006951f
C5075 vdd.n2811 gnd 0.006951f
C5076 vdd.n2812 gnd 0.006951f
C5077 vdd.n2813 gnd 0.006951f
C5078 vdd.n2814 gnd 0.006951f
C5079 vdd.n2815 gnd 0.006951f
C5080 vdd.n2816 gnd 0.006951f
C5081 vdd.n2817 gnd 0.006951f
C5082 vdd.n2818 gnd 0.006951f
C5083 vdd.n2819 gnd 0.006951f
C5084 vdd.n2820 gnd 0.006951f
C5085 vdd.n2821 gnd 0.006951f
C5086 vdd.n2822 gnd 0.006951f
C5087 vdd.n2823 gnd 0.006951f
C5088 vdd.n2824 gnd 0.006951f
C5089 vdd.n2825 gnd 0.006951f
C5090 vdd.n2826 gnd 0.006951f
C5091 vdd.n2827 gnd 0.006951f
C5092 vdd.n2828 gnd 0.006951f
C5093 vdd.n2829 gnd 0.006951f
C5094 vdd.n2830 gnd 0.006951f
C5095 vdd.n2831 gnd 0.006951f
C5096 vdd.n2832 gnd 0.006951f
C5097 vdd.n2833 gnd 0.006951f
C5098 vdd.n2834 gnd 0.006951f
C5099 vdd.n2835 gnd 0.006951f
C5100 vdd.n2836 gnd 0.006951f
C5101 vdd.n2837 gnd 0.006951f
C5102 vdd.n2838 gnd 0.006951f
C5103 vdd.n2839 gnd 0.006951f
C5104 vdd.n2840 gnd 0.006951f
C5105 vdd.n2841 gnd 0.006951f
C5106 vdd.n2842 gnd 0.006951f
C5107 vdd.n2843 gnd 0.006951f
C5108 vdd.n2844 gnd 0.006951f
C5109 vdd.n2845 gnd 0.006951f
C5110 vdd.n2846 gnd 0.006951f
C5111 vdd.n2847 gnd 0.006951f
C5112 vdd.n2848 gnd 0.006951f
C5113 vdd.n2849 gnd 0.006951f
C5114 vdd.n2850 gnd 0.006951f
C5115 vdd.n2851 gnd 0.006951f
C5116 vdd.n2852 gnd 0.016259f
C5117 vdd.n2853 gnd 0.016259f
C5118 vdd.n2855 gnd 0.867098f
C5119 vdd.n2857 gnd 0.016259f
C5120 vdd.n2858 gnd 0.016259f
C5121 vdd.n2859 gnd 0.015227f
C5122 vdd.n2860 gnd 0.006951f
C5123 vdd.n2861 gnd 0.006951f
C5124 vdd.n2862 gnd 0.376091f
C5125 vdd.n2863 gnd 0.006951f
C5126 vdd.n2864 gnd 0.006951f
C5127 vdd.n2865 gnd 0.006951f
C5128 vdd.n2866 gnd 0.006951f
C5129 vdd.n2867 gnd 0.006951f
C5130 vdd.n2868 gnd 0.423102f
C5131 vdd.n2869 gnd 0.006951f
C5132 vdd.n2870 gnd 0.006951f
C5133 vdd.n2871 gnd 0.006951f
C5134 vdd.n2872 gnd 0.006951f
C5135 vdd.n2873 gnd 0.006951f
C5136 vdd.n2874 gnd 0.710393f
C5137 vdd.n2875 gnd 0.006951f
C5138 vdd.n2876 gnd 0.006951f
C5139 vdd.n2877 gnd 0.006951f
C5140 vdd.n2878 gnd 0.006951f
C5141 vdd.n2879 gnd 0.006951f
C5142 vdd.n2880 gnd 0.470113f
C5143 vdd.n2881 gnd 0.006951f
C5144 vdd.n2882 gnd 0.006951f
C5145 vdd.n2883 gnd 0.006951f
C5146 vdd.n2884 gnd 0.006951f
C5147 vdd.n2885 gnd 0.006951f
C5148 vdd.n2886 gnd 0.626818f
C5149 vdd.n2887 gnd 0.006951f
C5150 vdd.n2888 gnd 0.006951f
C5151 vdd.n2889 gnd 0.006951f
C5152 vdd.n2890 gnd 0.006951f
C5153 vdd.n2891 gnd 0.006951f
C5154 vdd.n2892 gnd 0.569359f
C5155 vdd.n2893 gnd 0.006951f
C5156 vdd.n2894 gnd 0.006951f
C5157 vdd.n2895 gnd 0.006951f
C5158 vdd.n2896 gnd 0.006951f
C5159 vdd.n2897 gnd 0.006951f
C5160 vdd.n2898 gnd 0.412655f
C5161 vdd.n2899 gnd 0.006951f
C5162 vdd.n2900 gnd 0.006951f
C5163 vdd.n2901 gnd 0.006951f
C5164 vdd.n2902 gnd 0.006951f
C5165 vdd.n2903 gnd 0.006951f
C5166 vdd.n2904 gnd 0.22461f
C5167 vdd.n2905 gnd 0.006951f
C5168 vdd.n2906 gnd 0.006951f
C5169 vdd.n2907 gnd 0.006951f
C5170 vdd.n2908 gnd 0.006951f
C5171 vdd.n2909 gnd 0.006951f
C5172 vdd.n2910 gnd 0.611147f
C5173 vdd.n2911 gnd 0.006951f
C5174 vdd.n2912 gnd 0.006951f
C5175 vdd.n2913 gnd 0.006951f
C5176 vdd.n2914 gnd 0.006951f
C5177 vdd.n2915 gnd 0.006951f
C5178 vdd.n2916 gnd 0.710393f
C5179 vdd.n2917 gnd 0.006951f
C5180 vdd.n2918 gnd 0.006951f
C5181 vdd.n2919 gnd 0.004498f
C5182 vdd.n2920 gnd 0.020137f
C5183 vdd.n2921 gnd 0.005929f
C5184 vdd.n2922 gnd 0.006951f
C5185 vdd.n2923 gnd 0.605924f
C5186 vdd.n2924 gnd 0.006951f
C5187 vdd.n2925 gnd 0.006951f
C5188 vdd.n2926 gnd 0.006951f
C5189 vdd.n2927 gnd 0.006951f
C5190 vdd.n2928 gnd 0.006951f
C5191 vdd.n2929 gnd 0.496231f
C5192 vdd.n2930 gnd 0.006951f
C5193 vdd.n2931 gnd 0.006951f
C5194 vdd.n2932 gnd 0.006951f
C5195 vdd.n2933 gnd 0.006951f
C5196 vdd.n2934 gnd 0.006951f
C5197 vdd.n2935 gnd 0.370867f
C5198 vdd.n2936 gnd 0.006951f
C5199 vdd.n2937 gnd 0.006951f
C5200 vdd.n2938 gnd 0.006951f
C5201 vdd.n2939 gnd 0.006951f
C5202 vdd.n2940 gnd 0.006951f
C5203 vdd.n2941 gnd 0.710393f
C5204 vdd.n2942 gnd 0.006951f
C5205 vdd.n2943 gnd 0.006951f
C5206 vdd.n2944 gnd 0.006951f
C5207 vdd.n2945 gnd 0.006951f
C5208 vdd.n2946 gnd 0.006951f
C5209 vdd.n2947 gnd 0.006951f
C5210 vdd.n2949 gnd 0.006951f
C5211 vdd.n2950 gnd 0.006951f
C5212 vdd.n2952 gnd 0.006951f
C5213 vdd.n2953 gnd 0.006951f
C5214 vdd.n2956 gnd 0.006951f
C5215 vdd.n2957 gnd 0.006951f
C5216 vdd.n2958 gnd 0.006951f
C5217 vdd.n2959 gnd 0.006951f
C5218 vdd.n2961 gnd 0.006951f
C5219 vdd.n2962 gnd 0.006951f
C5220 vdd.n2963 gnd 0.006951f
C5221 vdd.n2964 gnd 0.006951f
C5222 vdd.n2965 gnd 0.006951f
C5223 vdd.n2966 gnd 0.006951f
C5224 vdd.n2968 gnd 0.006951f
C5225 vdd.n2969 gnd 0.006951f
C5226 vdd.n2970 gnd 0.006951f
C5227 vdd.n2971 gnd 0.006951f
C5228 vdd.n2972 gnd 0.006951f
C5229 vdd.n2973 gnd 0.006951f
C5230 vdd.n2975 gnd 0.006951f
C5231 vdd.n2976 gnd 0.006951f
C5232 vdd.n2977 gnd 0.006951f
C5233 vdd.n2978 gnd 0.006951f
C5234 vdd.n2979 gnd 0.006951f
C5235 vdd.n2980 gnd 0.006951f
C5236 vdd.n2982 gnd 0.006951f
C5237 vdd.n2983 gnd 0.016259f
C5238 vdd.n2984 gnd 0.016259f
C5239 vdd.n2985 gnd 0.015227f
C5240 vdd.n2986 gnd 0.006951f
C5241 vdd.n2987 gnd 0.006951f
C5242 vdd.n2988 gnd 0.006951f
C5243 vdd.n2989 gnd 0.006951f
C5244 vdd.n2990 gnd 0.006951f
C5245 vdd.n2991 gnd 0.006951f
C5246 vdd.n2992 gnd 0.710393f
C5247 vdd.n2993 gnd 0.006951f
C5248 vdd.n2994 gnd 0.006951f
C5249 vdd.n2995 gnd 0.006951f
C5250 vdd.n2996 gnd 0.006951f
C5251 vdd.n2997 gnd 0.006951f
C5252 vdd.n2998 gnd 0.46489f
C5253 vdd.n2999 gnd 0.006951f
C5254 vdd.n3000 gnd 0.006951f
C5255 vdd.n3001 gnd 0.006951f
C5256 vdd.n3002 gnd 0.01609f
C5257 vdd.n3004 gnd 0.016259f
C5258 vdd.n3005 gnd 0.015395f
C5259 vdd.n3006 gnd 0.006951f
C5260 vdd.n3007 gnd 0.005367f
C5261 vdd.n3008 gnd 0.006951f
C5262 vdd.n3010 gnd 0.006951f
C5263 vdd.n3011 gnd 0.006951f
C5264 vdd.n3012 gnd 0.006951f
C5265 vdd.n3013 gnd 0.006951f
C5266 vdd.n3014 gnd 0.006951f
C5267 vdd.n3015 gnd 0.006951f
C5268 vdd.n3017 gnd 0.006951f
C5269 vdd.n3018 gnd 0.006951f
C5270 vdd.n3019 gnd 0.006951f
C5271 vdd.n3020 gnd 0.006951f
C5272 vdd.n3021 gnd 0.006951f
C5273 vdd.n3022 gnd 0.006951f
C5274 vdd.n3024 gnd 0.006951f
C5275 vdd.n3025 gnd 0.006951f
C5276 vdd.n3026 gnd 0.006951f
C5277 vdd.n3027 gnd 0.006951f
C5278 vdd.n3028 gnd 0.006951f
C5279 vdd.n3029 gnd 0.006951f
C5280 vdd.n3031 gnd 0.006951f
C5281 vdd.n3032 gnd 0.006951f
C5282 vdd.n3033 gnd 0.006951f
C5283 vdd.n3034 gnd 0.777072f
C5284 vdd.n3035 gnd 0.023873f
C5285 vdd.n3036 gnd 0.006951f
C5286 vdd.n3037 gnd 0.006951f
C5287 vdd.n3039 gnd 0.006951f
C5288 vdd.n3040 gnd 0.006951f
C5289 vdd.n3041 gnd 0.006951f
C5290 vdd.n3042 gnd 0.006951f
C5291 vdd.n3043 gnd 0.006951f
C5292 vdd.n3044 gnd 0.006951f
C5293 vdd.n3046 gnd 0.006951f
C5294 vdd.n3047 gnd 0.006951f
C5295 vdd.n3048 gnd 0.006951f
C5296 vdd.n3049 gnd 0.006951f
C5297 vdd.n3050 gnd 0.006951f
C5298 vdd.n3051 gnd 0.006951f
C5299 vdd.n3053 gnd 0.006951f
C5300 vdd.n3054 gnd 0.006951f
C5301 vdd.n3055 gnd 0.006951f
C5302 vdd.n3056 gnd 0.006951f
C5303 vdd.n3057 gnd 0.006951f
C5304 vdd.n3058 gnd 0.006951f
C5305 vdd.n3060 gnd 0.006951f
C5306 vdd.n3061 gnd 0.006951f
C5307 vdd.n3063 gnd 0.006951f
C5308 vdd.n3064 gnd 0.006951f
C5309 vdd.n3065 gnd 0.016259f
C5310 vdd.n3066 gnd 0.015227f
C5311 vdd.n3067 gnd 0.015227f
C5312 vdd.n3068 gnd 1.00291f
C5313 vdd.n3069 gnd 0.015227f
C5314 vdd.n3070 gnd 0.016259f
C5315 vdd.n3071 gnd 0.015395f
C5316 vdd.n3072 gnd 0.006951f
C5317 vdd.n3073 gnd 0.005367f
C5318 vdd.n3074 gnd 0.006951f
C5319 vdd.n3076 gnd 0.006951f
C5320 vdd.n3077 gnd 0.006951f
C5321 vdd.n3078 gnd 0.006951f
C5322 vdd.n3079 gnd 0.006951f
C5323 vdd.n3080 gnd 0.006951f
C5324 vdd.n3081 gnd 0.006951f
C5325 vdd.n3083 gnd 0.006951f
C5326 vdd.n3084 gnd 0.006951f
C5327 vdd.n3085 gnd 0.006951f
C5328 vdd.n3086 gnd 0.006951f
C5329 vdd.n3087 gnd 0.006951f
C5330 vdd.n3088 gnd 0.006951f
C5331 vdd.n3090 gnd 0.006951f
C5332 vdd.n3091 gnd 0.006951f
C5333 vdd.n3092 gnd 0.006951f
C5334 vdd.n3093 gnd 0.006951f
C5335 vdd.n3094 gnd 0.006951f
C5336 vdd.n3095 gnd 0.006951f
C5337 vdd.n3097 gnd 0.006951f
C5338 vdd.n3098 gnd 0.006951f
C5339 vdd.n3100 gnd 0.006951f
C5340 vdd.n3101 gnd 0.023873f
C5341 vdd.n3102 gnd 0.777072f
C5342 vdd.n3103 gnd 0.008791f
C5343 vdd.n3104 gnd 0.003908f
C5344 vdd.t22 gnd 0.125764f
C5345 vdd.t23 gnd 0.134407f
C5346 vdd.t20 gnd 0.164246f
C5347 vdd.n3105 gnd 0.210541f
C5348 vdd.n3106 gnd 0.176892f
C5349 vdd.n3107 gnd 0.012671f
C5350 vdd.n3108 gnd 0.010223f
C5351 vdd.n3109 gnd 0.00432f
C5352 vdd.n3110 gnd 0.008228f
C5353 vdd.n3111 gnd 0.010223f
C5354 vdd.n3112 gnd 0.010223f
C5355 vdd.n3113 gnd 0.008228f
C5356 vdd.n3114 gnd 0.008228f
C5357 vdd.n3115 gnd 0.010223f
C5358 vdd.n3117 gnd 0.010223f
C5359 vdd.n3118 gnd 0.008228f
C5360 vdd.n3119 gnd 0.008228f
C5361 vdd.n3120 gnd 0.008228f
C5362 vdd.n3121 gnd 0.010223f
C5363 vdd.n3123 gnd 0.010223f
C5364 vdd.n3125 gnd 0.010223f
C5365 vdd.n3126 gnd 0.008228f
C5366 vdd.n3127 gnd 0.008228f
C5367 vdd.n3128 gnd 0.008228f
C5368 vdd.n3129 gnd 0.010223f
C5369 vdd.n3131 gnd 0.010223f
C5370 vdd.n3133 gnd 0.010223f
C5371 vdd.n3134 gnd 0.008228f
C5372 vdd.n3135 gnd 0.008228f
C5373 vdd.n3136 gnd 0.008228f
C5374 vdd.n3137 gnd 0.010223f
C5375 vdd.n3139 gnd 0.010223f
C5376 vdd.n3140 gnd 0.010223f
C5377 vdd.n3141 gnd 0.008228f
C5378 vdd.n3142 gnd 0.008228f
C5379 vdd.n3143 gnd 0.010223f
C5380 vdd.n3144 gnd 0.010223f
C5381 vdd.n3146 gnd 0.010223f
C5382 vdd.n3147 gnd 0.008228f
C5383 vdd.n3148 gnd 0.010223f
C5384 vdd.n3149 gnd 0.010223f
C5385 vdd.n3150 gnd 0.010223f
C5386 vdd.n3151 gnd 0.016785f
C5387 vdd.n3152 gnd 0.005595f
C5388 vdd.n3153 gnd 0.010223f
C5389 vdd.n3155 gnd 0.010223f
C5390 vdd.n3157 gnd 0.010223f
C5391 vdd.n3158 gnd 0.008228f
C5392 vdd.n3159 gnd 0.008228f
C5393 vdd.n3160 gnd 0.008228f
C5394 vdd.n3161 gnd 0.010223f
C5395 vdd.n3163 gnd 0.010223f
C5396 vdd.n3165 gnd 0.010223f
C5397 vdd.n3166 gnd 0.008228f
C5398 vdd.n3167 gnd 0.008228f
C5399 vdd.n3168 gnd 0.008228f
C5400 vdd.n3169 gnd 0.010223f
C5401 vdd.n3171 gnd 0.010223f
C5402 vdd.n3173 gnd 0.010223f
C5403 vdd.n3174 gnd 0.008228f
C5404 vdd.n3175 gnd 0.008228f
C5405 vdd.n3176 gnd 0.008228f
C5406 vdd.n3177 gnd 0.010223f
C5407 vdd.n3179 gnd 0.010223f
C5408 vdd.n3181 gnd 0.010223f
C5409 vdd.n3182 gnd 0.008228f
C5410 vdd.n3183 gnd 0.008228f
C5411 vdd.n3184 gnd 0.008228f
C5412 vdd.n3185 gnd 0.010223f
C5413 vdd.n3187 gnd 0.010223f
C5414 vdd.n3189 gnd 0.010223f
C5415 vdd.n3190 gnd 0.008228f
C5416 vdd.n3191 gnd 0.008228f
C5417 vdd.n3192 gnd 0.00687f
C5418 vdd.n3193 gnd 0.010223f
C5419 vdd.n3195 gnd 0.010223f
C5420 vdd.n3197 gnd 0.010223f
C5421 vdd.n3198 gnd 0.00687f
C5422 vdd.n3199 gnd 0.008228f
C5423 vdd.n3200 gnd 0.008228f
C5424 vdd.n3201 gnd 0.010223f
C5425 vdd.n3203 gnd 0.010223f
C5426 vdd.n3205 gnd 0.010223f
C5427 vdd.n3206 gnd 0.008228f
C5428 vdd.n3207 gnd 0.008228f
C5429 vdd.n3208 gnd 0.008228f
C5430 vdd.n3209 gnd 0.010223f
C5431 vdd.n3211 gnd 0.010223f
C5432 vdd.n3213 gnd 0.010223f
C5433 vdd.n3214 gnd 0.008228f
C5434 vdd.n3215 gnd 0.008228f
C5435 vdd.n3216 gnd 0.008228f
C5436 vdd.n3217 gnd 0.010223f
C5437 vdd.n3219 gnd 0.010223f
C5438 vdd.n3220 gnd 0.010223f
C5439 vdd.n3221 gnd 0.008228f
C5440 vdd.n3222 gnd 0.008228f
C5441 vdd.n3223 gnd 0.010223f
C5442 vdd.n3224 gnd 0.010223f
C5443 vdd.n3225 gnd 0.008228f
C5444 vdd.n3226 gnd 0.008228f
C5445 vdd.n3227 gnd 0.010223f
C5446 vdd.n3228 gnd 0.010223f
C5447 vdd.n3230 gnd 0.010223f
C5448 vdd.n3231 gnd 0.008228f
C5449 vdd.n3232 gnd 0.006829f
C5450 vdd.n3233 gnd 0.023438f
C5451 vdd.n3234 gnd 0.023279f
C5452 vdd.n3235 gnd 0.006829f
C5453 vdd.n3236 gnd 0.023279f
C5454 vdd.n3237 gnd 1.379f
C5455 vdd.n3238 gnd 0.023279f
C5456 vdd.n3239 gnd 0.006829f
C5457 vdd.n3240 gnd 0.023279f
C5458 vdd.n3241 gnd 0.010223f
C5459 vdd.n3242 gnd 0.010223f
C5460 vdd.n3243 gnd 0.008228f
C5461 vdd.n3244 gnd 0.010223f
C5462 vdd.n3245 gnd 0.987238f
C5463 vdd.n3246 gnd 0.010223f
C5464 vdd.n3247 gnd 0.008228f
C5465 vdd.n3248 gnd 0.010223f
C5466 vdd.n3249 gnd 0.010223f
C5467 vdd.n3250 gnd 0.010223f
C5468 vdd.n3251 gnd 0.008228f
C5469 vdd.n3252 gnd 0.010223f
C5470 vdd.n3253 gnd 1.01858f
C5471 vdd.n3254 gnd 0.010223f
C5472 vdd.n3255 gnd 0.008228f
C5473 vdd.n3256 gnd 0.010223f
C5474 vdd.n3257 gnd 0.010223f
C5475 vdd.n3258 gnd 0.010223f
C5476 vdd.n3259 gnd 0.008228f
C5477 vdd.n3260 gnd 0.010223f
C5478 vdd.t211 gnd 0.522348f
C5479 vdd.n3261 gnd 0.84098f
C5480 vdd.n3262 gnd 0.010223f
C5481 vdd.n3263 gnd 0.008228f
C5482 vdd.n3264 gnd 0.010223f
C5483 vdd.n3265 gnd 0.010223f
C5484 vdd.n3266 gnd 0.010223f
C5485 vdd.n3267 gnd 0.008228f
C5486 vdd.n3268 gnd 0.010223f
C5487 vdd.n3269 gnd 0.663382f
C5488 vdd.n3270 gnd 0.010223f
C5489 vdd.n3271 gnd 0.008228f
C5490 vdd.n3272 gnd 0.010223f
C5491 vdd.n3273 gnd 0.010223f
C5492 vdd.n3274 gnd 0.010223f
C5493 vdd.n3275 gnd 0.008228f
C5494 vdd.n3276 gnd 0.010223f
C5495 vdd.n3277 gnd 0.830533f
C5496 vdd.n3278 gnd 0.558912f
C5497 vdd.n3279 gnd 0.010223f
C5498 vdd.n3280 gnd 0.008228f
C5499 vdd.n3281 gnd 0.010223f
C5500 vdd.n3282 gnd 0.010223f
C5501 vdd.n3283 gnd 0.010223f
C5502 vdd.n3284 gnd 0.008228f
C5503 vdd.n3285 gnd 0.010223f
C5504 vdd.n3286 gnd 0.736511f
C5505 vdd.n3287 gnd 0.010223f
C5506 vdd.n3288 gnd 0.008228f
C5507 vdd.n3289 gnd 0.010223f
C5508 vdd.n3290 gnd 0.010223f
C5509 vdd.n3291 gnd 0.010223f
C5510 vdd.n3292 gnd 0.010223f
C5511 vdd.n3293 gnd 0.010223f
C5512 vdd.n3294 gnd 0.008228f
C5513 vdd.n3295 gnd 0.008228f
C5514 vdd.n3296 gnd 0.010223f
C5515 vdd.t157 gnd 0.522348f
C5516 vdd.n3297 gnd 0.867098f
C5517 vdd.n3298 gnd 0.010223f
C5518 vdd.n3299 gnd 0.008228f
C5519 vdd.n3300 gnd 0.010223f
C5520 vdd.n3301 gnd 0.010223f
C5521 vdd.n3302 gnd 0.010223f
C5522 vdd.n3303 gnd 0.008228f
C5523 vdd.n3304 gnd 0.010223f
C5524 vdd.n3305 gnd 0.820086f
C5525 vdd.n3306 gnd 0.010223f
C5526 vdd.n3307 gnd 0.010223f
C5527 vdd.n3308 gnd 0.008228f
C5528 vdd.n3309 gnd 0.008228f
C5529 vdd.n3310 gnd 0.008228f
C5530 vdd.n3311 gnd 0.010223f
C5531 vdd.n3312 gnd 0.010223f
C5532 vdd.n3313 gnd 0.010223f
C5533 vdd.n3314 gnd 0.010223f
C5534 vdd.n3315 gnd 0.008228f
C5535 vdd.n3316 gnd 0.008228f
C5536 vdd.n3317 gnd 0.008228f
C5537 vdd.n3318 gnd 0.010223f
C5538 vdd.n3319 gnd 0.010223f
C5539 vdd.n3320 gnd 0.010223f
C5540 vdd.n3321 gnd 0.010223f
C5541 vdd.n3322 gnd 0.008228f
C5542 vdd.n3323 gnd 0.008228f
C5543 vdd.n3324 gnd 0.008228f
C5544 vdd.n3325 gnd 0.010223f
C5545 vdd.n3326 gnd 0.010223f
C5546 vdd.n3327 gnd 0.010223f
C5547 vdd.n3328 gnd 0.867098f
C5548 vdd.n3329 gnd 0.010223f
C5549 vdd.n3330 gnd 0.008228f
C5550 vdd.n3331 gnd 0.008228f
C5551 vdd.n3332 gnd 0.008228f
C5552 vdd.n3333 gnd 0.010223f
C5553 vdd.n3334 gnd 0.010223f
C5554 vdd.n3335 gnd 0.010223f
C5555 vdd.n3336 gnd 0.010223f
C5556 vdd.n3337 gnd 0.008228f
C5557 vdd.n3338 gnd 0.008228f
C5558 vdd.n3339 gnd 0.006829f
C5559 vdd.n3340 gnd 0.023279f
C5560 vdd.n3341 gnd 0.023438f
C5561 vdd.n3342 gnd 0.003908f
C5562 vdd.n3343 gnd 0.023438f
C5563 vdd.n3345 gnd 2.30878f
C5564 vdd.n3346 gnd 1.379f
C5565 vdd.n3347 gnd 0.684276f
C5566 vdd.n3348 gnd 0.010223f
C5567 vdd.n3349 gnd 0.008228f
C5568 vdd.n3350 gnd 0.008228f
C5569 vdd.n3351 gnd 0.008228f
C5570 vdd.n3352 gnd 0.010223f
C5571 vdd.n3353 gnd 1.0447f
C5572 vdd.n3354 gnd 1.0447f
C5573 vdd.n3355 gnd 0.6007f
C5574 vdd.n3356 gnd 0.010223f
C5575 vdd.n3357 gnd 0.008228f
C5576 vdd.n3358 gnd 0.008228f
C5577 vdd.n3359 gnd 0.008228f
C5578 vdd.n3360 gnd 0.010223f
C5579 vdd.n3361 gnd 0.621594f
C5580 vdd.n3362 gnd 0.767852f
C5581 vdd.t127 gnd 0.522348f
C5582 vdd.n3363 gnd 0.799192f
C5583 vdd.n3364 gnd 0.010223f
C5584 vdd.n3365 gnd 0.008228f
C5585 vdd.n3366 gnd 0.008228f
C5586 vdd.n3367 gnd 0.008228f
C5587 vdd.n3368 gnd 0.010223f
C5588 vdd.n3369 gnd 0.867098f
C5589 vdd.t136 gnd 0.522348f
C5590 vdd.n3370 gnd 0.632041f
C5591 vdd.n3371 gnd 0.757405f
C5592 vdd.n3372 gnd 0.010223f
C5593 vdd.n3373 gnd 0.008228f
C5594 vdd.n3374 gnd 0.008228f
C5595 vdd.n3375 gnd 0.008228f
C5596 vdd.n3376 gnd 0.010223f
C5597 vdd.n3377 gnd 0.579806f
C5598 vdd.t160 gnd 0.522348f
C5599 vdd.n3378 gnd 0.867098f
C5600 vdd.t186 gnd 0.522348f
C5601 vdd.n3379 gnd 0.642488f
C5602 vdd.n3380 gnd 0.010223f
C5603 vdd.n3381 gnd 0.008228f
C5604 vdd.n3382 gnd 0.007857f
C5605 vdd.n3383 gnd 0.602964f
C5606 vdd.n3384 gnd 2.55746f
C5607 a_n7636_8799.t26 gnd 0.112164f
C5608 a_n7636_8799.t21 gnd 0.112164f
C5609 a_n7636_8799.t20 gnd 0.112164f
C5610 a_n7636_8799.n0 gnd 0.993322f
C5611 a_n7636_8799.t33 gnd 0.144211f
C5612 a_n7636_8799.t7 gnd 0.144211f
C5613 a_n7636_8799.n1 gnd 1.13741f
C5614 a_n7636_8799.t4 gnd 0.144211f
C5615 a_n7636_8799.t8 gnd 0.144211f
C5616 a_n7636_8799.n2 gnd 1.13553f
C5617 a_n7636_8799.n3 gnd 1.02071f
C5618 a_n7636_8799.t35 gnd 0.144211f
C5619 a_n7636_8799.t3 gnd 0.144211f
C5620 a_n7636_8799.n4 gnd 1.13553f
C5621 a_n7636_8799.n5 gnd 0.503125f
C5622 a_n7636_8799.t0 gnd 0.144211f
C5623 a_n7636_8799.t31 gnd 0.144211f
C5624 a_n7636_8799.n6 gnd 1.13553f
C5625 a_n7636_8799.n7 gnd 3.19547f
C5626 a_n7636_8799.t5 gnd 0.144211f
C5627 a_n7636_8799.t9 gnd 0.144211f
C5628 a_n7636_8799.n8 gnd 1.13741f
C5629 a_n7636_8799.t10 gnd 0.144211f
C5630 a_n7636_8799.t32 gnd 0.144211f
C5631 a_n7636_8799.n9 gnd 1.13553f
C5632 a_n7636_8799.n10 gnd 1.02071f
C5633 a_n7636_8799.t34 gnd 0.144211f
C5634 a_n7636_8799.t1 gnd 0.144211f
C5635 a_n7636_8799.n11 gnd 1.13553f
C5636 a_n7636_8799.n12 gnd 0.503125f
C5637 a_n7636_8799.t2 gnd 0.144211f
C5638 a_n7636_8799.t6 gnd 0.144211f
C5639 a_n7636_8799.n13 gnd 1.13553f
C5640 a_n7636_8799.n14 gnd 2.04015f
C5641 a_n7636_8799.n15 gnd 6.34701f
C5642 a_n7636_8799.n16 gnd 0.051978f
C5643 a_n7636_8799.t78 gnd 0.597964f
C5644 a_n7636_8799.n17 gnd 0.267062f
C5645 a_n7636_8799.n18 gnd 0.051978f
C5646 a_n7636_8799.n19 gnd 0.011795f
C5647 a_n7636_8799.t36 gnd 0.597964f
C5648 a_n7636_8799.n20 gnd 0.051978f
C5649 a_n7636_8799.t61 gnd 0.597964f
C5650 a_n7636_8799.n21 gnd 0.266902f
C5651 a_n7636_8799.t62 gnd 0.597964f
C5652 a_n7636_8799.n22 gnd 0.051978f
C5653 a_n7636_8799.n23 gnd 0.011795f
C5654 a_n7636_8799.t72 gnd 0.597964f
C5655 a_n7636_8799.n24 gnd 0.051978f
C5656 a_n7636_8799.t98 gnd 0.597964f
C5657 a_n7636_8799.n25 gnd 0.262095f
C5658 a_n7636_8799.t114 gnd 0.597964f
C5659 a_n7636_8799.n26 gnd 0.051978f
C5660 a_n7636_8799.t117 gnd 0.597964f
C5661 a_n7636_8799.n27 gnd 0.266261f
C5662 a_n7636_8799.t115 gnd 0.609282f
C5663 a_n7636_8799.n28 gnd 0.250693f
C5664 a_n7636_8799.n29 gnd 0.16996f
C5665 a_n7636_8799.n30 gnd 0.011795f
C5666 a_n7636_8799.t73 gnd 0.597964f
C5667 a_n7636_8799.n31 gnd 0.267062f
C5668 a_n7636_8799.n32 gnd 0.011795f
C5669 a_n7636_8799.n33 gnd 0.051978f
C5670 a_n7636_8799.n34 gnd 0.051978f
C5671 a_n7636_8799.n35 gnd 0.051978f
C5672 a_n7636_8799.n36 gnd 0.266582f
C5673 a_n7636_8799.n37 gnd 0.011795f
C5674 a_n7636_8799.t71 gnd 0.597964f
C5675 a_n7636_8799.n38 gnd 0.267062f
C5676 a_n7636_8799.n39 gnd 0.051978f
C5677 a_n7636_8799.n40 gnd 0.051978f
C5678 a_n7636_8799.n41 gnd 0.051978f
C5679 a_n7636_8799.n42 gnd 0.261775f
C5680 a_n7636_8799.t96 gnd 0.597964f
C5681 a_n7636_8799.n43 gnd 0.266902f
C5682 a_n7636_8799.n44 gnd 0.011795f
C5683 a_n7636_8799.n45 gnd 0.051978f
C5684 a_n7636_8799.n46 gnd 0.051978f
C5685 a_n7636_8799.n47 gnd 0.051978f
C5686 a_n7636_8799.n48 gnd 0.261775f
C5687 a_n7636_8799.n49 gnd 0.011795f
C5688 a_n7636_8799.t93 gnd 0.597964f
C5689 a_n7636_8799.n50 gnd 0.267062f
C5690 a_n7636_8799.n51 gnd 0.051978f
C5691 a_n7636_8799.n52 gnd 0.051978f
C5692 a_n7636_8799.n53 gnd 0.051978f
C5693 a_n7636_8799.n54 gnd 0.266582f
C5694 a_n7636_8799.t60 gnd 0.597964f
C5695 a_n7636_8799.n55 gnd 0.262095f
C5696 a_n7636_8799.n56 gnd 0.011795f
C5697 a_n7636_8799.n57 gnd 0.051978f
C5698 a_n7636_8799.n58 gnd 0.051978f
C5699 a_n7636_8799.n59 gnd 0.051978f
C5700 a_n7636_8799.n60 gnd 0.011795f
C5701 a_n7636_8799.t116 gnd 0.597964f
C5702 a_n7636_8799.n61 gnd 0.266261f
C5703 a_n7636_8799.t45 gnd 0.597964f
C5704 a_n7636_8799.n62 gnd 0.261614f
C5705 a_n7636_8799.n63 gnd 0.299489f
C5706 a_n7636_8799.n64 gnd 0.051978f
C5707 a_n7636_8799.t87 gnd 0.597964f
C5708 a_n7636_8799.n65 gnd 0.267062f
C5709 a_n7636_8799.n66 gnd 0.051978f
C5710 a_n7636_8799.n67 gnd 0.011795f
C5711 a_n7636_8799.t44 gnd 0.597964f
C5712 a_n7636_8799.n68 gnd 0.051978f
C5713 a_n7636_8799.t69 gnd 0.597964f
C5714 a_n7636_8799.n69 gnd 0.266902f
C5715 a_n7636_8799.t70 gnd 0.597964f
C5716 a_n7636_8799.n70 gnd 0.051978f
C5717 a_n7636_8799.n71 gnd 0.011795f
C5718 a_n7636_8799.t80 gnd 0.597964f
C5719 a_n7636_8799.n72 gnd 0.051978f
C5720 a_n7636_8799.t111 gnd 0.597964f
C5721 a_n7636_8799.n73 gnd 0.262095f
C5722 a_n7636_8799.t126 gnd 0.597964f
C5723 a_n7636_8799.n74 gnd 0.051978f
C5724 a_n7636_8799.t130 gnd 0.597964f
C5725 a_n7636_8799.n75 gnd 0.266261f
C5726 a_n7636_8799.t128 gnd 0.609282f
C5727 a_n7636_8799.n76 gnd 0.250693f
C5728 a_n7636_8799.n77 gnd 0.16996f
C5729 a_n7636_8799.n78 gnd 0.011795f
C5730 a_n7636_8799.t81 gnd 0.597964f
C5731 a_n7636_8799.n79 gnd 0.267062f
C5732 a_n7636_8799.n80 gnd 0.011795f
C5733 a_n7636_8799.n81 gnd 0.051978f
C5734 a_n7636_8799.n82 gnd 0.051978f
C5735 a_n7636_8799.n83 gnd 0.051978f
C5736 a_n7636_8799.n84 gnd 0.266582f
C5737 a_n7636_8799.n85 gnd 0.011795f
C5738 a_n7636_8799.t79 gnd 0.597964f
C5739 a_n7636_8799.n86 gnd 0.267062f
C5740 a_n7636_8799.n87 gnd 0.051978f
C5741 a_n7636_8799.n88 gnd 0.051978f
C5742 a_n7636_8799.n89 gnd 0.051978f
C5743 a_n7636_8799.n90 gnd 0.261775f
C5744 a_n7636_8799.t109 gnd 0.597964f
C5745 a_n7636_8799.n91 gnd 0.266902f
C5746 a_n7636_8799.n92 gnd 0.011795f
C5747 a_n7636_8799.n93 gnd 0.051978f
C5748 a_n7636_8799.n94 gnd 0.051978f
C5749 a_n7636_8799.n95 gnd 0.051978f
C5750 a_n7636_8799.n96 gnd 0.261775f
C5751 a_n7636_8799.n97 gnd 0.011795f
C5752 a_n7636_8799.t105 gnd 0.597964f
C5753 a_n7636_8799.n98 gnd 0.267062f
C5754 a_n7636_8799.n99 gnd 0.051978f
C5755 a_n7636_8799.n100 gnd 0.051978f
C5756 a_n7636_8799.n101 gnd 0.051978f
C5757 a_n7636_8799.n102 gnd 0.266582f
C5758 a_n7636_8799.t66 gnd 0.597964f
C5759 a_n7636_8799.n103 gnd 0.262095f
C5760 a_n7636_8799.n104 gnd 0.011795f
C5761 a_n7636_8799.n105 gnd 0.051978f
C5762 a_n7636_8799.n106 gnd 0.051978f
C5763 a_n7636_8799.n107 gnd 0.051978f
C5764 a_n7636_8799.n108 gnd 0.011795f
C5765 a_n7636_8799.t129 gnd 0.597964f
C5766 a_n7636_8799.n109 gnd 0.266261f
C5767 a_n7636_8799.t55 gnd 0.597964f
C5768 a_n7636_8799.n110 gnd 0.261614f
C5769 a_n7636_8799.n111 gnd 0.134663f
C5770 a_n7636_8799.n112 gnd 0.9006f
C5771 a_n7636_8799.n113 gnd 0.051978f
C5772 a_n7636_8799.t89 gnd 0.597964f
C5773 a_n7636_8799.n114 gnd 0.267062f
C5774 a_n7636_8799.n115 gnd 0.051978f
C5775 a_n7636_8799.n116 gnd 0.011795f
C5776 a_n7636_8799.t77 gnd 0.597964f
C5777 a_n7636_8799.n117 gnd 0.051978f
C5778 a_n7636_8799.t121 gnd 0.597964f
C5779 a_n7636_8799.n118 gnd 0.266902f
C5780 a_n7636_8799.t97 gnd 0.597964f
C5781 a_n7636_8799.n119 gnd 0.051978f
C5782 a_n7636_8799.n120 gnd 0.011795f
C5783 a_n7636_8799.t37 gnd 0.597964f
C5784 a_n7636_8799.n121 gnd 0.051978f
C5785 a_n7636_8799.t67 gnd 0.597964f
C5786 a_n7636_8799.n122 gnd 0.262095f
C5787 a_n7636_8799.t118 gnd 0.597964f
C5788 a_n7636_8799.n123 gnd 0.051978f
C5789 a_n7636_8799.t76 gnd 0.597964f
C5790 a_n7636_8799.n124 gnd 0.266261f
C5791 a_n7636_8799.t94 gnd 0.609282f
C5792 a_n7636_8799.n125 gnd 0.250693f
C5793 a_n7636_8799.n126 gnd 0.16996f
C5794 a_n7636_8799.n127 gnd 0.011795f
C5795 a_n7636_8799.t110 gnd 0.597964f
C5796 a_n7636_8799.n128 gnd 0.267062f
C5797 a_n7636_8799.n129 gnd 0.011795f
C5798 a_n7636_8799.n130 gnd 0.051978f
C5799 a_n7636_8799.n131 gnd 0.051978f
C5800 a_n7636_8799.n132 gnd 0.051978f
C5801 a_n7636_8799.n133 gnd 0.266582f
C5802 a_n7636_8799.n134 gnd 0.011795f
C5803 a_n7636_8799.t49 gnd 0.597964f
C5804 a_n7636_8799.n135 gnd 0.267062f
C5805 a_n7636_8799.n136 gnd 0.051978f
C5806 a_n7636_8799.n137 gnd 0.051978f
C5807 a_n7636_8799.n138 gnd 0.051978f
C5808 a_n7636_8799.n139 gnd 0.261775f
C5809 a_n7636_8799.t82 gnd 0.597964f
C5810 a_n7636_8799.n140 gnd 0.266902f
C5811 a_n7636_8799.n141 gnd 0.011795f
C5812 a_n7636_8799.n142 gnd 0.051978f
C5813 a_n7636_8799.n143 gnd 0.051978f
C5814 a_n7636_8799.n144 gnd 0.051978f
C5815 a_n7636_8799.n145 gnd 0.261775f
C5816 a_n7636_8799.n146 gnd 0.011795f
C5817 a_n7636_8799.t125 gnd 0.597964f
C5818 a_n7636_8799.n147 gnd 0.267062f
C5819 a_n7636_8799.n148 gnd 0.051978f
C5820 a_n7636_8799.n149 gnd 0.051978f
C5821 a_n7636_8799.n150 gnd 0.051978f
C5822 a_n7636_8799.n151 gnd 0.266582f
C5823 a_n7636_8799.t41 gnd 0.597964f
C5824 a_n7636_8799.n152 gnd 0.262095f
C5825 a_n7636_8799.n153 gnd 0.011795f
C5826 a_n7636_8799.n154 gnd 0.051978f
C5827 a_n7636_8799.n155 gnd 0.051978f
C5828 a_n7636_8799.n156 gnd 0.051978f
C5829 a_n7636_8799.n157 gnd 0.011795f
C5830 a_n7636_8799.t53 gnd 0.597964f
C5831 a_n7636_8799.n158 gnd 0.266261f
C5832 a_n7636_8799.t106 gnd 0.597964f
C5833 a_n7636_8799.n159 gnd 0.261614f
C5834 a_n7636_8799.n160 gnd 0.134663f
C5835 a_n7636_8799.n161 gnd 1.5812f
C5836 a_n7636_8799.n162 gnd 0.051978f
C5837 a_n7636_8799.t75 gnd 0.597964f
C5838 a_n7636_8799.t57 gnd 0.597964f
C5839 a_n7636_8799.t120 gnd 0.597964f
C5840 a_n7636_8799.n163 gnd 0.267062f
C5841 a_n7636_8799.n164 gnd 0.051978f
C5842 a_n7636_8799.t88 gnd 0.597964f
C5843 a_n7636_8799.t86 gnd 0.597964f
C5844 a_n7636_8799.n165 gnd 0.051978f
C5845 a_n7636_8799.t38 gnd 0.597964f
C5846 a_n7636_8799.n166 gnd 0.267062f
C5847 a_n7636_8799.n167 gnd 0.051978f
C5848 a_n7636_8799.t92 gnd 0.597964f
C5849 a_n7636_8799.t91 gnd 0.597964f
C5850 a_n7636_8799.n168 gnd 0.051978f
C5851 a_n7636_8799.t40 gnd 0.597964f
C5852 a_n7636_8799.n169 gnd 0.266902f
C5853 a_n7636_8799.n170 gnd 0.051978f
C5854 a_n7636_8799.t39 gnd 0.597964f
C5855 a_n7636_8799.t108 gnd 0.597964f
C5856 a_n7636_8799.n171 gnd 0.051978f
C5857 a_n7636_8799.t52 gnd 0.597964f
C5858 a_n7636_8799.n172 gnd 0.266582f
C5859 a_n7636_8799.n173 gnd 0.051978f
C5860 a_n7636_8799.t43 gnd 0.597964f
C5861 a_n7636_8799.t112 gnd 0.597964f
C5862 a_n7636_8799.n174 gnd 0.051978f
C5863 a_n7636_8799.t74 gnd 0.597964f
C5864 a_n7636_8799.n175 gnd 0.266261f
C5865 a_n7636_8799.t56 gnd 0.609282f
C5866 a_n7636_8799.n176 gnd 0.250693f
C5867 a_n7636_8799.n177 gnd 0.16996f
C5868 a_n7636_8799.n178 gnd 0.011795f
C5869 a_n7636_8799.n179 gnd 0.267062f
C5870 a_n7636_8799.n180 gnd 0.011795f
C5871 a_n7636_8799.n181 gnd 0.262095f
C5872 a_n7636_8799.n182 gnd 0.051978f
C5873 a_n7636_8799.n183 gnd 0.051978f
C5874 a_n7636_8799.n184 gnd 0.051978f
C5875 a_n7636_8799.n185 gnd 0.011795f
C5876 a_n7636_8799.n186 gnd 0.267062f
C5877 a_n7636_8799.n187 gnd 0.011795f
C5878 a_n7636_8799.n188 gnd 0.261775f
C5879 a_n7636_8799.n189 gnd 0.051978f
C5880 a_n7636_8799.n190 gnd 0.051978f
C5881 a_n7636_8799.n191 gnd 0.051978f
C5882 a_n7636_8799.n192 gnd 0.011795f
C5883 a_n7636_8799.n193 gnd 0.266902f
C5884 a_n7636_8799.n194 gnd 0.261775f
C5885 a_n7636_8799.n195 gnd 0.011795f
C5886 a_n7636_8799.n196 gnd 0.051978f
C5887 a_n7636_8799.n197 gnd 0.051978f
C5888 a_n7636_8799.n198 gnd 0.051978f
C5889 a_n7636_8799.n199 gnd 0.011795f
C5890 a_n7636_8799.n200 gnd 0.266582f
C5891 a_n7636_8799.n201 gnd 0.262095f
C5892 a_n7636_8799.n202 gnd 0.011795f
C5893 a_n7636_8799.n203 gnd 0.051978f
C5894 a_n7636_8799.n204 gnd 0.051978f
C5895 a_n7636_8799.n205 gnd 0.051978f
C5896 a_n7636_8799.n206 gnd 0.011795f
C5897 a_n7636_8799.n207 gnd 0.266261f
C5898 a_n7636_8799.n208 gnd 0.261614f
C5899 a_n7636_8799.n209 gnd 0.299489f
C5900 a_n7636_8799.n210 gnd 0.051978f
C5901 a_n7636_8799.t84 gnd 0.597964f
C5902 a_n7636_8799.t64 gnd 0.597964f
C5903 a_n7636_8799.t131 gnd 0.597964f
C5904 a_n7636_8799.n211 gnd 0.267062f
C5905 a_n7636_8799.n212 gnd 0.051978f
C5906 a_n7636_8799.t101 gnd 0.597964f
C5907 a_n7636_8799.t100 gnd 0.597964f
C5908 a_n7636_8799.n213 gnd 0.051978f
C5909 a_n7636_8799.t46 gnd 0.597964f
C5910 a_n7636_8799.n214 gnd 0.267062f
C5911 a_n7636_8799.n215 gnd 0.051978f
C5912 a_n7636_8799.t104 gnd 0.597964f
C5913 a_n7636_8799.t103 gnd 0.597964f
C5914 a_n7636_8799.n216 gnd 0.051978f
C5915 a_n7636_8799.t48 gnd 0.597964f
C5916 a_n7636_8799.n217 gnd 0.266902f
C5917 a_n7636_8799.n218 gnd 0.051978f
C5918 a_n7636_8799.t47 gnd 0.597964f
C5919 a_n7636_8799.t123 gnd 0.597964f
C5920 a_n7636_8799.n219 gnd 0.051978f
C5921 a_n7636_8799.t63 gnd 0.597964f
C5922 a_n7636_8799.n220 gnd 0.266582f
C5923 a_n7636_8799.n221 gnd 0.051978f
C5924 a_n7636_8799.t51 gnd 0.597964f
C5925 a_n7636_8799.t124 gnd 0.597964f
C5926 a_n7636_8799.n222 gnd 0.051978f
C5927 a_n7636_8799.t85 gnd 0.597964f
C5928 a_n7636_8799.n223 gnd 0.266261f
C5929 a_n7636_8799.t65 gnd 0.609282f
C5930 a_n7636_8799.n224 gnd 0.250693f
C5931 a_n7636_8799.n225 gnd 0.16996f
C5932 a_n7636_8799.n226 gnd 0.011795f
C5933 a_n7636_8799.n227 gnd 0.267062f
C5934 a_n7636_8799.n228 gnd 0.011795f
C5935 a_n7636_8799.n229 gnd 0.262095f
C5936 a_n7636_8799.n230 gnd 0.051978f
C5937 a_n7636_8799.n231 gnd 0.051978f
C5938 a_n7636_8799.n232 gnd 0.051978f
C5939 a_n7636_8799.n233 gnd 0.011795f
C5940 a_n7636_8799.n234 gnd 0.267062f
C5941 a_n7636_8799.n235 gnd 0.011795f
C5942 a_n7636_8799.n236 gnd 0.261775f
C5943 a_n7636_8799.n237 gnd 0.051978f
C5944 a_n7636_8799.n238 gnd 0.051978f
C5945 a_n7636_8799.n239 gnd 0.051978f
C5946 a_n7636_8799.n240 gnd 0.011795f
C5947 a_n7636_8799.n241 gnd 0.266902f
C5948 a_n7636_8799.n242 gnd 0.261775f
C5949 a_n7636_8799.n243 gnd 0.011795f
C5950 a_n7636_8799.n244 gnd 0.051978f
C5951 a_n7636_8799.n245 gnd 0.051978f
C5952 a_n7636_8799.n246 gnd 0.051978f
C5953 a_n7636_8799.n247 gnd 0.011795f
C5954 a_n7636_8799.n248 gnd 0.266582f
C5955 a_n7636_8799.n249 gnd 0.262095f
C5956 a_n7636_8799.n250 gnd 0.011795f
C5957 a_n7636_8799.n251 gnd 0.051978f
C5958 a_n7636_8799.n252 gnd 0.051978f
C5959 a_n7636_8799.n253 gnd 0.051978f
C5960 a_n7636_8799.n254 gnd 0.011795f
C5961 a_n7636_8799.n255 gnd 0.266261f
C5962 a_n7636_8799.n256 gnd 0.261614f
C5963 a_n7636_8799.n257 gnd 0.134663f
C5964 a_n7636_8799.n258 gnd 0.9006f
C5965 a_n7636_8799.n259 gnd 0.051978f
C5966 a_n7636_8799.t107 gnd 0.597964f
C5967 a_n7636_8799.t54 gnd 0.597964f
C5968 a_n7636_8799.t90 gnd 0.597964f
C5969 a_n7636_8799.n260 gnd 0.267062f
C5970 a_n7636_8799.n261 gnd 0.051978f
C5971 a_n7636_8799.t42 gnd 0.597964f
C5972 a_n7636_8799.t59 gnd 0.597964f
C5973 a_n7636_8799.n262 gnd 0.051978f
C5974 a_n7636_8799.t127 gnd 0.597964f
C5975 a_n7636_8799.n263 gnd 0.267062f
C5976 a_n7636_8799.n264 gnd 0.051978f
C5977 a_n7636_8799.t99 gnd 0.597964f
C5978 a_n7636_8799.t122 gnd 0.597964f
C5979 a_n7636_8799.n265 gnd 0.051978f
C5980 a_n7636_8799.t83 gnd 0.597964f
C5981 a_n7636_8799.n266 gnd 0.266902f
C5982 a_n7636_8799.n267 gnd 0.051978f
C5983 a_n7636_8799.t102 gnd 0.597964f
C5984 a_n7636_8799.t50 gnd 0.597964f
C5985 a_n7636_8799.n268 gnd 0.051978f
C5986 a_n7636_8799.t119 gnd 0.597964f
C5987 a_n7636_8799.n269 gnd 0.266582f
C5988 a_n7636_8799.n270 gnd 0.051978f
C5989 a_n7636_8799.t68 gnd 0.597964f
C5990 a_n7636_8799.t113 gnd 0.597964f
C5991 a_n7636_8799.n271 gnd 0.051978f
C5992 a_n7636_8799.t58 gnd 0.597964f
C5993 a_n7636_8799.n272 gnd 0.266261f
C5994 a_n7636_8799.t95 gnd 0.609282f
C5995 a_n7636_8799.n273 gnd 0.250693f
C5996 a_n7636_8799.n274 gnd 0.16996f
C5997 a_n7636_8799.n275 gnd 0.011795f
C5998 a_n7636_8799.n276 gnd 0.267062f
C5999 a_n7636_8799.n277 gnd 0.011795f
C6000 a_n7636_8799.n278 gnd 0.262095f
C6001 a_n7636_8799.n279 gnd 0.051978f
C6002 a_n7636_8799.n280 gnd 0.051978f
C6003 a_n7636_8799.n281 gnd 0.051978f
C6004 a_n7636_8799.n282 gnd 0.011795f
C6005 a_n7636_8799.n283 gnd 0.267062f
C6006 a_n7636_8799.n284 gnd 0.011795f
C6007 a_n7636_8799.n285 gnd 0.261775f
C6008 a_n7636_8799.n286 gnd 0.051978f
C6009 a_n7636_8799.n287 gnd 0.051978f
C6010 a_n7636_8799.n288 gnd 0.051978f
C6011 a_n7636_8799.n289 gnd 0.011795f
C6012 a_n7636_8799.n290 gnd 0.266902f
C6013 a_n7636_8799.n291 gnd 0.261775f
C6014 a_n7636_8799.n292 gnd 0.011795f
C6015 a_n7636_8799.n293 gnd 0.051978f
C6016 a_n7636_8799.n294 gnd 0.051978f
C6017 a_n7636_8799.n295 gnd 0.051978f
C6018 a_n7636_8799.n296 gnd 0.011795f
C6019 a_n7636_8799.n297 gnd 0.266582f
C6020 a_n7636_8799.n298 gnd 0.262095f
C6021 a_n7636_8799.n299 gnd 0.011795f
C6022 a_n7636_8799.n300 gnd 0.051978f
C6023 a_n7636_8799.n301 gnd 0.051978f
C6024 a_n7636_8799.n302 gnd 0.051978f
C6025 a_n7636_8799.n303 gnd 0.011795f
C6026 a_n7636_8799.n304 gnd 0.266261f
C6027 a_n7636_8799.n305 gnd 0.261614f
C6028 a_n7636_8799.n306 gnd 0.134663f
C6029 a_n7636_8799.n307 gnd 1.21407f
C6030 a_n7636_8799.n308 gnd 13.9797f
C6031 a_n7636_8799.n309 gnd 4.37623f
C6032 a_n7636_8799.t17 gnd 0.112164f
C6033 a_n7636_8799.t18 gnd 0.112164f
C6034 a_n7636_8799.n310 gnd 0.993323f
C6035 a_n7636_8799.t13 gnd 0.112164f
C6036 a_n7636_8799.t14 gnd 0.112164f
C6037 a_n7636_8799.n311 gnd 0.991118f
C6038 a_n7636_8799.n312 gnd 0.789471f
C6039 a_n7636_8799.t12 gnd 0.112164f
C6040 a_n7636_8799.t27 gnd 0.112164f
C6041 a_n7636_8799.n313 gnd 0.991118f
C6042 a_n7636_8799.n314 gnd 0.742285f
C6043 a_n7636_8799.t28 gnd 0.112164f
C6044 a_n7636_8799.t23 gnd 0.112164f
C6045 a_n7636_8799.n315 gnd 0.991118f
C6046 a_n7636_8799.n316 gnd 0.387671f
C6047 a_n7636_8799.t25 gnd 0.112164f
C6048 a_n7636_8799.t11 gnd 0.112164f
C6049 a_n7636_8799.n317 gnd 0.991118f
C6050 a_n7636_8799.n318 gnd 2.71144f
C6051 a_n7636_8799.t24 gnd 0.112164f
C6052 a_n7636_8799.t22 gnd 0.112164f
C6053 a_n7636_8799.n319 gnd 0.993322f
C6054 a_n7636_8799.t15 gnd 0.112164f
C6055 a_n7636_8799.t19 gnd 0.112164f
C6056 a_n7636_8799.n320 gnd 0.991118f
C6057 a_n7636_8799.n321 gnd 0.789473f
C6058 a_n7636_8799.t29 gnd 0.112164f
C6059 a_n7636_8799.t16 gnd 0.112164f
C6060 a_n7636_8799.n322 gnd 0.991118f
C6061 a_n7636_8799.n323 gnd 2.46832f
C6062 a_n7636_8799.n324 gnd 0.789476f
C6063 a_n7636_8799.n325 gnd 0.991115f
C6064 a_n7636_8799.t30 gnd 0.112164f
C6065 a_n3827_n3924.n0 gnd 1.20073f
C6066 a_n3827_n3924.n1 gnd 1.70952f
C6067 a_n3827_n3924.n2 gnd 0.682766f
C6068 a_n3827_n3924.n3 gnd 1.54211f
C6069 a_n3827_n3924.n4 gnd 2.05091f
C6070 a_n3827_n3924.n5 gnd 1.58291f
C6071 a_n3827_n3924.n6 gnd 0.900145f
C6072 a_n3827_n3924.n7 gnd 1.67197f
C6073 a_n3827_n3924.n8 gnd 1.67197f
C6074 a_n3827_n3924.n9 gnd 2.84498f
C6075 a_n3827_n3924.n10 gnd 2.34829f
C6076 a_n3827_n3924.t24 gnd 0.091917f
C6077 a_n3827_n3924.t11 gnd 0.091917f
C6078 a_n3827_n3924.t15 gnd 0.091917f
C6079 a_n3827_n3924.n11 gnd 0.750697f
C6080 a_n3827_n3924.t49 gnd 1.19019f
C6081 a_n3827_n3924.t3 gnd 1.18694f
C6082 a_n3827_n3924.t13 gnd 0.955305f
C6083 a_n3827_n3924.t18 gnd 1.18864f
C6084 a_n3827_n3924.t16 gnd 1.18694f
C6085 a_n3827_n3924.t48 gnd 1.18694f
C6086 a_n3827_n3924.t17 gnd 1.18694f
C6087 a_n3827_n3924.t47 gnd 1.18694f
C6088 a_n3827_n3924.t9 gnd 1.18694f
C6089 a_n3827_n3924.t20 gnd 1.18694f
C6090 a_n3827_n3924.t10 gnd 1.18694f
C6091 a_n3827_n3924.n12 gnd 0.862207f
C6092 a_n3827_n3924.t43 gnd 0.955301f
C6093 a_n3827_n3924.t34 gnd 0.091917f
C6094 a_n3827_n3924.t40 gnd 0.091917f
C6095 a_n3827_n3924.n13 gnd 0.750696f
C6096 a_n3827_n3924.t37 gnd 0.091917f
C6097 a_n3827_n3924.t38 gnd 0.091917f
C6098 a_n3827_n3924.n14 gnd 0.750696f
C6099 a_n3827_n3924.t41 gnd 0.091917f
C6100 a_n3827_n3924.t33 gnd 0.091917f
C6101 a_n3827_n3924.n15 gnd 0.750696f
C6102 a_n3827_n3924.t30 gnd 0.091917f
C6103 a_n3827_n3924.t31 gnd 0.091917f
C6104 a_n3827_n3924.n16 gnd 0.750696f
C6105 a_n3827_n3924.t45 gnd 0.955301f
C6106 a_n3827_n3924.t8 gnd 0.955301f
C6107 a_n3827_n3924.t26 gnd 0.091917f
C6108 a_n3827_n3924.t12 gnd 0.091917f
C6109 a_n3827_n3924.n17 gnd 0.750696f
C6110 a_n3827_n3924.t2 gnd 0.091917f
C6111 a_n3827_n3924.t7 gnd 0.091917f
C6112 a_n3827_n3924.n18 gnd 0.750696f
C6113 a_n3827_n3924.t6 gnd 0.091917f
C6114 a_n3827_n3924.t5 gnd 0.091917f
C6115 a_n3827_n3924.n19 gnd 0.750696f
C6116 a_n3827_n3924.t21 gnd 0.091917f
C6117 a_n3827_n3924.t22 gnd 0.091917f
C6118 a_n3827_n3924.n20 gnd 0.750696f
C6119 a_n3827_n3924.t1 gnd 0.955301f
C6120 a_n3827_n3924.n21 gnd 0.862207f
C6121 a_n3827_n3924.t46 gnd 0.955301f
C6122 a_n3827_n3924.t39 gnd 0.091917f
C6123 a_n3827_n3924.t27 gnd 0.091917f
C6124 a_n3827_n3924.n22 gnd 0.750697f
C6125 a_n3827_n3924.t35 gnd 0.091917f
C6126 a_n3827_n3924.t36 gnd 0.091917f
C6127 a_n3827_n3924.n23 gnd 0.750697f
C6128 a_n3827_n3924.t42 gnd 0.091917f
C6129 a_n3827_n3924.t29 gnd 0.091917f
C6130 a_n3827_n3924.n24 gnd 0.750697f
C6131 a_n3827_n3924.t28 gnd 0.091917f
C6132 a_n3827_n3924.t44 gnd 0.091917f
C6133 a_n3827_n3924.n25 gnd 0.750697f
C6134 a_n3827_n3924.t32 gnd 0.955305f
C6135 a_n3827_n3924.t14 gnd 0.955305f
C6136 a_n3827_n3924.t19 gnd 0.091917f
C6137 a_n3827_n3924.t4 gnd 0.091917f
C6138 a_n3827_n3924.n26 gnd 0.750697f
C6139 a_n3827_n3924.t25 gnd 0.091917f
C6140 a_n3827_n3924.t23 gnd 0.091917f
C6141 a_n3827_n3924.n27 gnd 0.750697f
C6142 a_n3827_n3924.n28 gnd 0.750698f
C6143 a_n3827_n3924.t0 gnd 0.091917f
C6144 plus.n0 gnd 0.022377f
C6145 plus.t14 gnd 0.316499f
C6146 plus.n1 gnd 0.022377f
C6147 plus.t15 gnd 0.316499f
C6148 plus.t9 gnd 0.316499f
C6149 plus.n2 gnd 0.140599f
C6150 plus.n3 gnd 0.022377f
C6151 plus.t5 gnd 0.316499f
C6152 plus.t6 gnd 0.316499f
C6153 plus.n4 gnd 0.140599f
C6154 plus.n5 gnd 0.022377f
C6155 plus.t19 gnd 0.316499f
C6156 plus.t20 gnd 0.316499f
C6157 plus.n6 gnd 0.140599f
C6158 plus.n7 gnd 0.022377f
C6159 plus.t16 gnd 0.316499f
C6160 plus.t11 gnd 0.316499f
C6161 plus.n8 gnd 0.144342f
C6162 plus.t13 gnd 0.327587f
C6163 plus.n9 gnd 0.131117f
C6164 plus.n10 gnd 0.095513f
C6165 plus.n11 gnd 0.005078f
C6166 plus.n12 gnd 0.140599f
C6167 plus.n13 gnd 0.005078f
C6168 plus.n14 gnd 0.022377f
C6169 plus.n15 gnd 0.022377f
C6170 plus.n16 gnd 0.022377f
C6171 plus.n17 gnd 0.005078f
C6172 plus.n18 gnd 0.140599f
C6173 plus.n19 gnd 0.005078f
C6174 plus.n20 gnd 0.022377f
C6175 plus.n21 gnd 0.022377f
C6176 plus.n22 gnd 0.022377f
C6177 plus.n23 gnd 0.005078f
C6178 plus.n24 gnd 0.140599f
C6179 plus.n25 gnd 0.005078f
C6180 plus.n26 gnd 0.022377f
C6181 plus.n27 gnd 0.022377f
C6182 plus.n28 gnd 0.022377f
C6183 plus.n29 gnd 0.005078f
C6184 plus.n30 gnd 0.140599f
C6185 plus.n31 gnd 0.005078f
C6186 plus.n32 gnd 0.140392f
C6187 plus.n33 gnd 0.252782f
C6188 plus.n34 gnd 0.022377f
C6189 plus.n35 gnd 0.005078f
C6190 plus.t10 gnd 0.316499f
C6191 plus.n36 gnd 0.022377f
C6192 plus.n37 gnd 0.005078f
C6193 plus.t7 gnd 0.316499f
C6194 plus.n38 gnd 0.022377f
C6195 plus.n39 gnd 0.005078f
C6196 plus.t23 gnd 0.316499f
C6197 plus.n40 gnd 0.022377f
C6198 plus.n41 gnd 0.005078f
C6199 plus.t22 gnd 0.316499f
C6200 plus.t18 gnd 0.327587f
C6201 plus.t17 gnd 0.316499f
C6202 plus.n42 gnd 0.144342f
C6203 plus.n43 gnd 0.131117f
C6204 plus.n44 gnd 0.095513f
C6205 plus.n45 gnd 0.022377f
C6206 plus.n46 gnd 0.140599f
C6207 plus.n47 gnd 0.005078f
C6208 plus.t21 gnd 0.316499f
C6209 plus.n48 gnd 0.140599f
C6210 plus.n49 gnd 0.022377f
C6211 plus.n50 gnd 0.022377f
C6212 plus.n51 gnd 0.022377f
C6213 plus.n52 gnd 0.140599f
C6214 plus.n53 gnd 0.005078f
C6215 plus.t8 gnd 0.316499f
C6216 plus.n54 gnd 0.140599f
C6217 plus.n55 gnd 0.022377f
C6218 plus.n56 gnd 0.022377f
C6219 plus.n57 gnd 0.022377f
C6220 plus.n58 gnd 0.140599f
C6221 plus.n59 gnd 0.005078f
C6222 plus.t12 gnd 0.316499f
C6223 plus.n60 gnd 0.140599f
C6224 plus.n61 gnd 0.022377f
C6225 plus.n62 gnd 0.022377f
C6226 plus.n63 gnd 0.022377f
C6227 plus.n64 gnd 0.140599f
C6228 plus.n65 gnd 0.005078f
C6229 plus.t24 gnd 0.316499f
C6230 plus.n66 gnd 0.140392f
C6231 plus.n67 gnd 0.690234f
C6232 plus.n68 gnd 1.0438f
C6233 plus.t1 gnd 0.038629f
C6234 plus.t4 gnd 0.006898f
C6235 plus.t0 gnd 0.006898f
C6236 plus.n69 gnd 0.022372f
C6237 plus.n70 gnd 0.173674f
C6238 plus.t2 gnd 0.006898f
C6239 plus.t3 gnd 0.006898f
C6240 plus.n71 gnd 0.022372f
C6241 plus.n72 gnd 0.130363f
C6242 plus.n73 gnd 2.96826f
.ends

