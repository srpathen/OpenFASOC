* NGSPICE file created from opamp.ext - technology: sky130A

.subckt opamp output vdd plus minus commonsourceibias outputibias diffpairibias gnd CSoutput
Cload output gnd 0.0p
X0 CSoutput.t108 commonsourceibias.t48 gnd.t187 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X1 a_n5644_8799.t19 plus.t5 a_n2903_n3924.t17 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X2 vdd.t86 a_n5644_8799.t32 CSoutput.t115 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X3 a_n1986_8322.t19 a_n1996_n452.t44 vdd.t107 vdd.t106 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 a_n1808_13878.t11 a_n1996_n452.t26 a_n1996_n452.t27 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X5 CSoutput.t107 commonsourceibias.t49 gnd.t186 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X6 gnd.t185 commonsourceibias.t50 CSoutput.t106 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 CSoutput.t105 commonsourceibias.t51 gnd.t184 gnd.t108 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 gnd.t323 gnd.t321 plus.t4 gnd.t322 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X9 a_n2903_n3924.t16 plus.t6 a_n5644_8799.t18 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X10 a_n1996_n452.t21 a_n1996_n452.t20 a_n1808_13878.t10 vdd.t88 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X11 a_n1808_13878.t9 a_n1996_n452.t28 a_n1996_n452.t29 vdd.t108 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X12 vdd.t199 vdd.t197 vdd.t198 vdd.t172 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X13 a_n1808_13878.t19 a_n1996_n452.t45 vdd.t110 vdd.t109 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X14 output.t3 outputibias.t8 gnd.t46 gnd.t45 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X15 CSoutput.t24 a_n5644_8799.t33 vdd.t85 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X16 a_n2903_n3924.t25 minus.t5 a_n1996_n452.t2 gnd.t17 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X17 vdd.t196 vdd.t194 vdd.t195 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X18 gnd.t183 commonsourceibias.t52 CSoutput.t104 gnd.t90 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X19 CSoutput.t103 commonsourceibias.t53 gnd.t182 gnd.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 gnd.t181 commonsourceibias.t54 CSoutput.t102 gnd.t79 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X21 CSoutput.t101 commonsourceibias.t55 gnd.t180 gnd.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X22 a_n1996_n452.t9 minus.t6 a_n2903_n3924.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X23 gnd.t320 gnd.t317 gnd.t319 gnd.t318 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X24 CSoutput.t100 commonsourceibias.t56 gnd.t179 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X25 a_n1986_8322.t11 a_n1996_n452.t46 a_n5644_8799.t26 vdd.t87 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X26 CSoutput.t99 commonsourceibias.t57 gnd.t178 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X27 a_n1996_n452.t40 minus.t7 a_n2903_n3924.t39 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X28 gnd.t177 commonsourceibias.t58 CSoutput.t98 gnd.t120 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X29 CSoutput.t97 commonsourceibias.t59 gnd.t176 gnd.t100 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X30 CSoutput.t96 commonsourceibias.t60 gnd.t175 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X31 gnd.t316 gnd.t314 gnd.t315 gnd.t240 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X32 a_n2903_n3924.t28 minus.t8 a_n1996_n452.t5 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X33 CSoutput.t120 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X34 CSoutput.t2 a_n5644_8799.t34 vdd.t84 vdd.t42 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X35 vdd.t83 a_n5644_8799.t35 CSoutput.t21 vdd.t60 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X36 CSoutput.t95 commonsourceibias.t61 gnd.t174 gnd.t116 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 a_n5644_8799.t20 a_n1996_n452.t47 a_n1986_8322.t10 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X38 CSoutput.t13 a_n5644_8799.t36 vdd.t82 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X39 vdd.t81 a_n5644_8799.t37 CSoutput.t10 vdd.t76 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X40 gnd.t161 commonsourceibias.t62 CSoutput.t94 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X41 a_n2903_n3924.t41 diffpairibias.t16 gnd.t48 gnd.t47 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X42 CSoutput.t93 commonsourceibias.t63 gnd.t173 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X43 gnd.t172 commonsourceibias.t46 commonsourceibias.t47 gnd.t93 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X44 gnd.t313 gnd.t310 gnd.t312 gnd.t311 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X45 output.t19 CSoutput.t121 vdd.t99 gnd.t58 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X46 CSoutput.t92 commonsourceibias.t64 gnd.t171 gnd.t116 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X47 CSoutput.t119 a_n5644_8799.t38 vdd.t80 vdd.t38 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X48 vdd.t193 vdd.t191 vdd.t192 vdd.t125 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X49 a_n2903_n3924.t11 plus.t7 a_n5644_8799.t17 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X50 CSoutput.t91 commonsourceibias.t65 gnd.t170 gnd.t95 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X51 a_n5644_8799.t16 plus.t8 a_n2903_n3924.t7 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X52 outputibias.t7 outputibias.t6 gnd.t189 gnd.t188 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X53 gnd.t169 commonsourceibias.t66 CSoutput.t90 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X54 output.t18 CSoutput.t122 vdd.t92 gnd.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X55 CSoutput.t89 commonsourceibias.t67 gnd.t168 gnd.t95 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X56 gnd.t309 gnd.t307 gnd.t308 gnd.t240 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X57 CSoutput.t88 commonsourceibias.t68 gnd.t167 gnd.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X58 gnd.t166 commonsourceibias.t44 commonsourceibias.t45 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X59 gnd.t306 gnd.t304 gnd.t305 gnd.t215 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X60 a_n1808_13878.t8 a_n1996_n452.t24 a_n1996_n452.t25 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X61 vdd.t79 a_n5644_8799.t39 CSoutput.t111 vdd.t76 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X62 a_n1996_n452.t41 minus.t9 a_n2903_n3924.t40 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X63 diffpairibias.t15 diffpairibias.t14 gnd.t193 gnd.t192 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X64 a_n1996_n452.t23 a_n1996_n452.t22 a_n1808_13878.t7 vdd.t120 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X65 CSoutput.t1 a_n5644_8799.t40 vdd.t78 vdd.t54 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X66 CSoutput.t87 commonsourceibias.t69 gnd.t165 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X67 CSoutput.t86 commonsourceibias.t70 gnd.t164 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X68 vdd.t190 vdd.t188 vdd.t189 vdd.t157 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X69 gnd.t163 commonsourceibias.t71 CSoutput.t85 gnd.t103 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X70 gnd.t160 commonsourceibias.t72 CSoutput.t84 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X71 plus.t3 gnd.t301 gnd.t303 gnd.t302 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X72 CSoutput.t83 commonsourceibias.t73 gnd.t162 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X73 diffpairibias.t13 diffpairibias.t12 gnd.t195 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X74 gnd.t159 commonsourceibias.t26 commonsourceibias.t27 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X75 vdd.t187 vdd.t185 vdd.t186 vdd.t136 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X76 gnd.t300 gnd.t298 gnd.t299 gnd.t223 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X77 CSoutput.t82 commonsourceibias.t74 gnd.t158 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X78 gnd.t157 commonsourceibias.t75 CSoutput.t81 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X79 CSoutput.t80 commonsourceibias.t76 gnd.t156 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 vdd.t77 a_n5644_8799.t41 CSoutput.t12 vdd.t76 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 gnd.t155 commonsourceibias.t77 CSoutput.t79 gnd.t120 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X82 output.t17 CSoutput.t123 vdd.t90 gnd.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X83 vdd.t75 a_n5644_8799.t42 CSoutput.t110 vdd.t51 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X84 CSoutput.t27 a_n5644_8799.t43 vdd.t74 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X85 vdd.t73 a_n5644_8799.t44 CSoutput.t3 vdd.t27 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 a_n2903_n3924.t3 plus.t9 a_n5644_8799.t15 gnd.t55 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X87 gnd.t154 commonsourceibias.t78 CSoutput.t78 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 gnd.t297 gnd.t294 gnd.t296 gnd.t295 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X89 CSoutput.t22 a_n5644_8799.t45 vdd.t72 vdd.t38 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X90 CSoutput.t28 a_n5644_8799.t46 vdd.t71 vdd.t64 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X91 vdd.t89 CSoutput.t124 output.t16 gnd.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X92 a_n2903_n3924.t42 diffpairibias.t17 gnd.t52 gnd.t51 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X93 CSoutput.t33 a_n5644_8799.t47 vdd.t70 vdd.t64 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X94 gnd.t153 commonsourceibias.t79 CSoutput.t77 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X95 gnd.t293 gnd.t291 gnd.t292 gnd.t219 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X96 vdd.t69 a_n5644_8799.t48 CSoutput.t15 vdd.t62 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X97 gnd.t290 gnd.t288 gnd.t289 gnd.t219 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X98 a_n1996_n452.t37 a_n1996_n452.t36 a_n1808_13878.t6 vdd.t87 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X99 a_n1996_n452.t31 a_n1996_n452.t30 a_n1808_13878.t5 vdd.t9 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X100 vdd.t68 a_n5644_8799.t49 CSoutput.t19 vdd.t60 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X101 a_n5644_8799.t24 a_n1996_n452.t48 a_n1986_8322.t9 vdd.t20 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X102 gnd.t152 commonsourceibias.t80 CSoutput.t76 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X103 vdd.t67 a_n5644_8799.t50 CSoutput.t36 vdd.t62 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X104 a_n1996_n452.t4 minus.t10 a_n2903_n3924.t27 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X105 gnd.t151 commonsourceibias.t81 CSoutput.t75 gnd.t93 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X106 gnd.t150 commonsourceibias.t2 commonsourceibias.t3 gnd.t79 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X107 vdd.t91 CSoutput.t125 output.t15 gnd.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X108 vdd.t184 vdd.t182 vdd.t183 vdd.t136 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X109 a_n2903_n3924.t26 minus.t11 a_n1996_n452.t3 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X110 output.t14 CSoutput.t126 vdd.t100 gnd.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X111 CSoutput.t127 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X112 output.t2 outputibias.t9 gnd.t57 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X113 vdd.t66 a_n5644_8799.t51 CSoutput.t4 vdd.t51 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X114 vdd.t181 vdd.t179 vdd.t180 vdd.t165 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X115 vdd.t178 vdd.t175 vdd.t177 vdd.t176 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X116 gnd.t287 gnd.t285 gnd.t286 gnd.t233 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X117 CSoutput.t74 commonsourceibias.t82 gnd.t149 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X118 a_n2903_n3924.t46 diffpairibias.t18 gnd.t191 gnd.t190 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X119 outputibias.t5 outputibias.t4 gnd.t42 gnd.t41 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X120 vdd.t174 vdd.t171 vdd.t173 vdd.t172 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X121 gnd.t284 gnd.t282 gnd.t283 gnd.t215 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X122 CSoutput.t73 commonsourceibias.t83 gnd.t148 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X123 a_n2903_n3924.t38 minus.t12 a_n1996_n452.t39 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X124 output.t13 CSoutput.t128 vdd.t98 gnd.t24 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X125 vdd.t3 a_n1996_n452.t49 a_n1986_8322.t18 vdd.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X126 vdd.t170 vdd.t168 vdd.t169 vdd.t161 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X127 a_n1996_n452.t38 minus.t13 a_n2903_n3924.t37 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X128 CSoutput.t11 a_n5644_8799.t52 vdd.t65 vdd.t64 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X129 a_n1986_8322.t17 a_n1996_n452.t50 vdd.t123 vdd.t122 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X130 a_n2903_n3924.t12 plus.t10 a_n5644_8799.t14 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X131 a_n2903_n3924.t5 plus.t11 a_n5644_8799.t13 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X132 outputibias.t3 outputibias.t2 gnd.t66 gnd.t65 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X133 vdd.t63 a_n5644_8799.t53 CSoutput.t16 vdd.t62 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X134 gnd.t281 gnd.t279 gnd.t280 gnd.t219 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X135 vdd.t5 a_n1996_n452.t51 a_n1808_13878.t18 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X136 a_n5644_8799.t12 plus.t12 a_n2903_n3924.t1 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X137 a_n5644_8799.t11 plus.t13 a_n2903_n3924.t9 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X138 vdd.t167 vdd.t164 vdd.t166 vdd.t165 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X139 a_n1996_n452.t10 minus.t14 a_n2903_n3924.t33 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X140 diffpairibias.t11 diffpairibias.t10 gnd.t203 gnd.t202 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X141 vdd.t163 vdd.t160 vdd.t162 vdd.t161 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X142 vdd.t61 a_n5644_8799.t54 CSoutput.t0 vdd.t60 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X143 CSoutput.t72 commonsourceibias.t84 gnd.t147 gnd.t108 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X144 gnd.t278 gnd.t276 minus.t4 gnd.t277 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X145 gnd.t146 commonsourceibias.t85 CSoutput.t71 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X146 commonsourceibias.t1 commonsourceibias.t0 gnd.t145 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X147 a_n5644_8799.t27 a_n1996_n452.t52 a_n1986_8322.t8 vdd.t105 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X148 a_n1986_8322.t16 a_n1996_n452.t53 vdd.t114 vdd.t113 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X149 vdd.t159 vdd.t156 vdd.t158 vdd.t157 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X150 a_n2903_n3924.t35 minus.t15 a_n1996_n452.t12 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X151 vdd.t103 CSoutput.t129 output.t12 gnd.t25 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X152 a_n1996_n452.t35 a_n1996_n452.t34 a_n1808_13878.t4 vdd.t121 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X153 CSoutput.t130 a_n1986_8322.t23 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X154 a_n5644_8799.t25 a_n1996_n452.t54 a_n1986_8322.t7 vdd.t108 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X155 CSoutput.t70 commonsourceibias.t86 gnd.t144 gnd.t95 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X156 CSoutput.t131 a_n1986_8322.t22 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X157 a_n1808_13878.t3 a_n1996_n452.t14 a_n1996_n452.t15 vdd.t20 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X158 gnd.t142 commonsourceibias.t87 CSoutput.t69 gnd.t120 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X159 gnd.t143 commonsourceibias.t88 CSoutput.t68 gnd.t103 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X160 commonsourceibias.t37 commonsourceibias.t36 gnd.t141 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X161 gnd.t139 commonsourceibias.t89 CSoutput.t67 gnd.t90 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X162 vdd.t117 a_n1996_n452.t55 a_n1986_8322.t15 vdd.t116 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X163 gnd.t275 gnd.t273 minus.t3 gnd.t274 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X164 CSoutput.t66 commonsourceibias.t90 gnd.t138 gnd.t100 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 a_n2903_n3924.t14 plus.t14 a_n5644_8799.t10 gnd.t17 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X166 outputibias.t1 outputibias.t0 gnd.t199 gnd.t198 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X167 vdd.t155 vdd.t153 vdd.t154 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X168 gnd.t272 gnd.t269 gnd.t271 gnd.t270 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X169 a_n2903_n3924.t22 diffpairibias.t19 gnd.t11 gnd.t10 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X170 CSoutput.t25 a_n5644_8799.t55 vdd.t59 vdd.t54 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X171 a_n2903_n3924.t24 diffpairibias.t20 gnd.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X172 output.t1 outputibias.t10 gnd.t50 gnd.t49 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X173 commonsourceibias.t35 commonsourceibias.t34 gnd.t137 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X174 vdd.t58 a_n5644_8799.t56 CSoutput.t8 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X175 a_n5644_8799.t9 plus.t15 a_n2903_n3924.t0 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X176 gnd.t268 gnd.t266 gnd.t267 gnd.t240 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X177 gnd.t265 gnd.t262 gnd.t264 gnd.t263 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X178 CSoutput.t65 commonsourceibias.t91 gnd.t135 gnd.t108 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X179 CSoutput.t64 commonsourceibias.t92 gnd.t134 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X180 vdd.t57 a_n5644_8799.t57 CSoutput.t17 vdd.t40 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X181 output.t11 CSoutput.t132 vdd.t102 gnd.t59 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X182 gnd.t261 gnd.t259 gnd.t260 gnd.t208 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X183 commonsourceibias.t33 commonsourceibias.t32 gnd.t133 gnd.t116 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X184 diffpairibias.t9 diffpairibias.t8 gnd.t64 gnd.t63 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X185 CSoutput.t63 commonsourceibias.t93 gnd.t132 gnd.t100 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X186 CSoutput.t62 commonsourceibias.t94 gnd.t131 gnd.t72 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X187 output.t10 CSoutput.t133 vdd.t101 gnd.t60 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X188 gnd.t130 commonsourceibias.t30 commonsourceibias.t31 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X189 CSoutput.t20 a_n5644_8799.t58 vdd.t56 vdd.t44 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X190 commonsourceibias.t17 commonsourceibias.t16 gnd.t128 gnd.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X191 vdd.t152 vdd.t150 vdd.t151 vdd.t132 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X192 a_n1808_13878.t17 a_n1996_n452.t56 vdd.t22 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X193 vdd.t14 a_n1996_n452.t57 a_n1808_13878.t16 vdd.t13 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X194 gnd.t126 commonsourceibias.t95 CSoutput.t61 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X195 a_n2903_n3924.t30 minus.t16 a_n1996_n452.t7 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X196 commonsourceibias.t15 commonsourceibias.t14 gnd.t125 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X197 vdd.t149 vdd.t146 vdd.t148 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X198 gnd.t124 commonsourceibias.t12 commonsourceibias.t13 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X199 a_n1996_n452.t6 minus.t17 a_n2903_n3924.t29 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X200 gnd.t258 gnd.t256 gnd.t257 gnd.t208 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X201 diffpairibias.t7 diffpairibias.t6 gnd.t54 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X202 commonsourceibias.t11 commonsourceibias.t10 gnd.t123 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X203 CSoutput.t109 a_n5644_8799.t59 vdd.t55 vdd.t54 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X204 plus.t2 gnd.t253 gnd.t255 gnd.t254 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X205 a_n1996_n452.t11 minus.t18 a_n2903_n3924.t34 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X206 vdd.t53 a_n5644_8799.t60 CSoutput.t35 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X207 a_n5644_8799.t8 plus.t16 a_n2903_n3924.t8 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X208 a_n1986_8322.t6 a_n1996_n452.t58 a_n5644_8799.t29 vdd.t88 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X209 gnd.t252 gnd.t250 minus.t2 gnd.t251 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X210 gnd.t122 commonsourceibias.t96 CSoutput.t60 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X211 a_n2903_n3924.t20 minus.t19 a_n1996_n452.t0 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X212 vdd.t96 CSoutput.t134 output.t9 gnd.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X213 output.t0 outputibias.t11 gnd.t30 gnd.t29 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X214 vdd.t97 CSoutput.t135 output.t8 gnd.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X215 vdd.t52 a_n5644_8799.t61 CSoutput.t23 vdd.t51 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X216 CSoutput.t32 a_n5644_8799.t62 vdd.t50 vdd.t31 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X217 gnd.t121 commonsourceibias.t8 commonsourceibias.t9 gnd.t120 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X218 vdd.t49 a_n5644_8799.t63 CSoutput.t30 vdd.t40 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X219 vdd.t112 a_n1996_n452.t59 a_n1986_8322.t14 vdd.t111 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X220 a_n1808_13878.t15 a_n1996_n452.t60 vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X221 minus.t1 gnd.t247 gnd.t249 gnd.t248 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X222 gnd.t246 gnd.t243 gnd.t245 gnd.t244 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X223 a_n2903_n3924.t43 diffpairibias.t21 gnd.t62 gnd.t61 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X224 CSoutput.t116 a_n5644_8799.t64 vdd.t48 vdd.t44 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X225 gnd.t119 commonsourceibias.t6 commonsourceibias.t7 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X226 CSoutput.t114 a_n5644_8799.t65 vdd.t47 vdd.t42 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X227 CSoutput.t136 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X228 vdd.t145 vdd.t143 vdd.t144 vdd.t132 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X229 a_n5644_8799.t7 plus.t17 a_n2903_n3924.t2 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X230 a_n1986_8322.t5 a_n1996_n452.t61 a_n5644_8799.t30 vdd.t121 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X231 vdd.t16 a_n1996_n452.t62 a_n1986_8322.t13 vdd.t15 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X232 vdd.t46 a_n5644_8799.t66 CSoutput.t14 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X233 CSoutput.t7 a_n5644_8799.t67 vdd.t45 vdd.t44 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X234 a_n2903_n3924.t4 plus.t18 a_n5644_8799.t6 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X235 gnd.t118 commonsourceibias.t4 commonsourceibias.t5 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X236 CSoutput.t59 commonsourceibias.t97 gnd.t117 gnd.t116 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X237 vdd.t104 CSoutput.t137 output.t7 gnd.t26 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X238 diffpairibias.t5 diffpairibias.t4 gnd.t44 gnd.t43 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X239 output.t6 CSoutput.t138 vdd.t93 gnd.t27 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X240 vdd.t142 vdd.t139 vdd.t141 vdd.t140 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X241 vdd.t138 vdd.t135 vdd.t137 vdd.t136 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X242 gnd.t242 gnd.t239 gnd.t241 gnd.t240 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X243 a_n1808_13878.t2 a_n1996_n452.t16 a_n1996_n452.t17 vdd.t12 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X244 CSoutput.t58 commonsourceibias.t98 gnd.t115 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X245 a_n1986_8322.t4 a_n1996_n452.t63 a_n5644_8799.t31 vdd.t120 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X246 gnd.t113 commonsourceibias.t99 CSoutput.t57 gnd.t93 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X247 gnd.t238 gnd.t236 gnd.t237 gnd.t208 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X248 CSoutput.t31 a_n5644_8799.t68 vdd.t43 vdd.t42 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X249 a_n1986_8322.t12 a_n1996_n452.t64 vdd.t8 vdd.t7 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X250 gnd.t235 gnd.t232 gnd.t234 gnd.t233 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X251 minus.t0 gnd.t229 gnd.t231 gnd.t230 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X252 gnd.t112 commonsourceibias.t100 CSoutput.t56 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X253 gnd.t111 commonsourceibias.t101 CSoutput.t55 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X254 vdd.t18 a_n1996_n452.t65 a_n1808_13878.t14 vdd.t17 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X255 gnd.t228 gnd.t226 gnd.t227 gnd.t215 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X256 a_n2903_n3924.t36 minus.t20 a_n1996_n452.t13 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X257 commonsourceibias.t29 commonsourceibias.t28 gnd.t109 gnd.t108 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X258 gnd.t110 commonsourceibias.t102 CSoutput.t54 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X259 gnd.t225 gnd.t222 gnd.t224 gnd.t223 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X260 vdd.t94 CSoutput.t139 output.t5 gnd.t28 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X261 vdd.t134 vdd.t131 vdd.t133 vdd.t132 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X262 a_n1996_n452.t42 minus.t21 a_n2903_n3924.t44 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X263 a_n1986_8322.t3 a_n1996_n452.t66 a_n5644_8799.t28 vdd.t115 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X264 vdd.t130 vdd.t128 vdd.t129 vdd.t125 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X265 a_n5644_8799.t21 a_n1996_n452.t67 a_n1986_8322.t2 vdd.t12 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X266 a_n1808_13878.t13 a_n1996_n452.t68 vdd.t119 vdd.t118 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X267 vdd.t41 a_n5644_8799.t69 CSoutput.t18 vdd.t40 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X268 CSoutput.t117 a_n5644_8799.t70 vdd.t39 vdd.t38 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X269 gnd.t107 commonsourceibias.t103 CSoutput.t53 gnd.t103 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X270 a_n5644_8799.t5 plus.t19 a_n2903_n3924.t18 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X271 commonsourceibias.t19 commonsourceibias.t18 gnd.t96 gnd.t95 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X272 a_n2903_n3924.t45 minus.t22 a_n1996_n452.t43 gnd.t55 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X273 gnd.t106 commonsourceibias.t104 CSoutput.t52 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X274 gnd.t104 commonsourceibias.t24 commonsourceibias.t25 gnd.t103 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 a_n2903_n3924.t13 plus.t20 a_n5644_8799.t4 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X276 gnd.t102 commonsourceibias.t22 commonsourceibias.t23 gnd.t90 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X277 commonsourceibias.t21 commonsourceibias.t20 gnd.t101 gnd.t100 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 CSoutput.t112 a_n5644_8799.t71 vdd.t37 vdd.t31 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X279 a_n1808_13878.t1 a_n1996_n452.t32 a_n1996_n452.t33 vdd.t105 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X280 a_n2903_n3924.t47 diffpairibias.t22 gnd.t201 gnd.t200 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X281 gnd.t99 commonsourceibias.t105 CSoutput.t51 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X282 CSoutput.t50 commonsourceibias.t106 gnd.t97 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X283 gnd.t94 commonsourceibias.t107 CSoutput.t49 gnd.t93 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X284 gnd.t221 gnd.t218 gnd.t220 gnd.t219 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X285 gnd.t217 gnd.t214 gnd.t216 gnd.t215 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X286 a_n5644_8799.t3 plus.t21 a_n2903_n3924.t19 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X287 CSoutput.t6 a_n5644_8799.t72 vdd.t36 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X288 gnd.t213 gnd.t211 plus.t1 gnd.t212 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X289 CSoutput.t48 commonsourceibias.t108 gnd.t92 gnd.t72 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X290 gnd.t91 commonsourceibias.t109 CSoutput.t47 gnd.t90 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X291 commonsourceibias.t43 commonsourceibias.t42 gnd.t89 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X292 vdd.t35 a_n5644_8799.t73 CSoutput.t34 vdd.t27 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X293 gnd.t210 gnd.t207 gnd.t209 gnd.t208 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X294 diffpairibias.t3 diffpairibias.t2 gnd.t197 gnd.t196 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X295 a_n5644_8799.t22 a_n1996_n452.t69 a_n1986_8322.t1 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X296 a_n1996_n452.t19 a_n1996_n452.t18 a_n1808_13878.t0 vdd.t115 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X297 gnd.t206 gnd.t204 plus.t0 gnd.t205 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X298 gnd.t87 commonsourceibias.t110 CSoutput.t46 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X299 a_n2903_n3924.t15 plus.t22 a_n5644_8799.t2 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X300 vdd.t34 a_n5644_8799.t74 CSoutput.t29 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X301 vdd.t127 vdd.t124 vdd.t126 vdd.t125 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X302 CSoutput.t140 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X303 diffpairibias.t1 diffpairibias.t0 gnd.t40 gnd.t39 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X304 a_n2903_n3924.t6 plus.t23 a_n5644_8799.t1 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X305 gnd.t86 commonsourceibias.t111 CSoutput.t45 gnd.t79 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X306 commonsourceibias.t41 commonsourceibias.t40 gnd.t85 gnd.t72 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 CSoutput.t44 commonsourceibias.t112 gnd.t84 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X308 a_n5644_8799.t0 plus.t24 a_n2903_n3924.t10 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X309 a_n2903_n3924.t31 minus.t23 a_n1996_n452.t8 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X310 gnd.t82 commonsourceibias.t38 commonsourceibias.t39 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X311 vdd.t11 a_n1996_n452.t70 a_n1808_13878.t12 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X312 CSoutput.t118 a_n5644_8799.t75 vdd.t32 vdd.t31 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X313 a_n1996_n452.t1 minus.t24 a_n2903_n3924.t21 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X314 gnd.t80 commonsourceibias.t113 CSoutput.t43 gnd.t79 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X315 gnd.t78 commonsourceibias.t114 CSoutput.t42 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X316 vdd.t95 CSoutput.t141 output.t4 gnd.t67 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X317 gnd.t74 commonsourceibias.t115 CSoutput.t41 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X318 CSoutput.t5 a_n5644_8799.t76 vdd.t30 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X319 gnd.t76 commonsourceibias.t116 CSoutput.t40 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X320 vdd.t28 a_n5644_8799.t77 CSoutput.t113 vdd.t27 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X321 a_n1986_8322.t0 a_n1996_n452.t71 a_n5644_8799.t23 vdd.t9 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X322 CSoutput.t39 commonsourceibias.t117 gnd.t73 gnd.t72 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X323 gnd.t71 commonsourceibias.t118 CSoutput.t38 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X324 CSoutput.t37 commonsourceibias.t119 gnd.t69 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X325 vdd.t26 a_n5644_8799.t78 CSoutput.t26 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X326 CSoutput.t9 a_n5644_8799.t79 vdd.t24 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X327 a_n2903_n3924.t23 diffpairibias.t23 gnd.t14 gnd.t13 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
R0 commonsourceibias.n25 commonsourceibias.t10 230.006
R1 commonsourceibias.n91 commonsourceibias.t73 230.006
R2 commonsourceibias.n218 commonsourceibias.t98 230.006
R3 commonsourceibias.n154 commonsourceibias.t69 230.006
R4 commonsourceibias.n322 commonsourceibias.t2 230.006
R5 commonsourceibias.n281 commonsourceibias.t111 230.006
R6 commonsourceibias.n483 commonsourceibias.t113 230.006
R7 commonsourceibias.n419 commonsourceibias.t54 230.006
R8 commonsourceibias.n70 commonsourceibias.t22 207.983
R9 commonsourceibias.n136 commonsourceibias.t89 207.983
R10 commonsourceibias.n263 commonsourceibias.t109 207.983
R11 commonsourceibias.n199 commonsourceibias.t52 207.983
R12 commonsourceibias.n368 commonsourceibias.t14 207.983
R13 commonsourceibias.n402 commonsourceibias.t70 207.983
R14 commonsourceibias.n529 commonsourceibias.t63 207.983
R15 commonsourceibias.n465 commonsourceibias.t112 207.983
R16 commonsourceibias.n10 commonsourceibias.t0 168.701
R17 commonsourceibias.n63 commonsourceibias.t38 168.701
R18 commonsourceibias.n57 commonsourceibias.t20 168.701
R19 commonsourceibias.n16 commonsourceibias.t44 168.701
R20 commonsourceibias.n49 commonsourceibias.t18 168.701
R21 commonsourceibias.n43 commonsourceibias.t8 168.701
R22 commonsourceibias.n19 commonsourceibias.t40 168.701
R23 commonsourceibias.n21 commonsourceibias.t24 168.701
R24 commonsourceibias.n23 commonsourceibias.t34 168.701
R25 commonsourceibias.n26 commonsourceibias.t4 168.701
R26 commonsourceibias.n1 commonsourceibias.t49 168.701
R27 commonsourceibias.n129 commonsourceibias.t95 168.701
R28 commonsourceibias.n123 commonsourceibias.t90 168.701
R29 commonsourceibias.n7 commonsourceibias.t100 168.701
R30 commonsourceibias.n115 commonsourceibias.t86 168.701
R31 commonsourceibias.n109 commonsourceibias.t77 168.701
R32 commonsourceibias.n85 commonsourceibias.t94 168.701
R33 commonsourceibias.n87 commonsourceibias.t88 168.701
R34 commonsourceibias.n89 commonsourceibias.t60 168.701
R35 commonsourceibias.n92 commonsourceibias.t80 168.701
R36 commonsourceibias.n219 commonsourceibias.t102 168.701
R37 commonsourceibias.n216 commonsourceibias.t48 168.701
R38 commonsourceibias.n214 commonsourceibias.t103 168.701
R39 commonsourceibias.n212 commonsourceibias.t108 168.701
R40 commonsourceibias.n236 commonsourceibias.t87 168.701
R41 commonsourceibias.n242 commonsourceibias.t67 168.701
R42 commonsourceibias.n209 commonsourceibias.t115 168.701
R43 commonsourceibias.n250 commonsourceibias.t93 168.701
R44 commonsourceibias.n256 commonsourceibias.t96 168.701
R45 commonsourceibias.n203 commonsourceibias.t57 168.701
R46 commonsourceibias.n139 commonsourceibias.t119 168.701
R47 commonsourceibias.n192 commonsourceibias.t110 168.701
R48 commonsourceibias.n186 commonsourceibias.t59 168.701
R49 commonsourceibias.n145 commonsourceibias.t118 168.701
R50 commonsourceibias.n178 commonsourceibias.t65 168.701
R51 commonsourceibias.n172 commonsourceibias.t58 168.701
R52 commonsourceibias.n148 commonsourceibias.t117 168.701
R53 commonsourceibias.n150 commonsourceibias.t71 168.701
R54 commonsourceibias.n152 commonsourceibias.t83 168.701
R55 commonsourceibias.n155 commonsourceibias.t116 168.701
R56 commonsourceibias.n323 commonsourceibias.t32 168.701
R57 commonsourceibias.n320 commonsourceibias.t26 168.701
R58 commonsourceibias.n318 commonsourceibias.t16 168.701
R59 commonsourceibias.n316 commonsourceibias.t6 168.701
R60 commonsourceibias.n340 commonsourceibias.t36 168.701
R61 commonsourceibias.n346 commonsourceibias.t30 168.701
R62 commonsourceibias.n348 commonsourceibias.t42 168.701
R63 commonsourceibias.n355 commonsourceibias.t12 168.701
R64 commonsourceibias.n361 commonsourceibias.t28 168.701
R65 commonsourceibias.n308 commonsourceibias.t46 168.701
R66 commonsourceibias.n267 commonsourceibias.t99 168.701
R67 commonsourceibias.n395 commonsourceibias.t84 168.701
R68 commonsourceibias.n389 commonsourceibias.t72 168.701
R69 commonsourceibias.n382 commonsourceibias.t92 168.701
R70 commonsourceibias.n380 commonsourceibias.t66 168.701
R71 commonsourceibias.n282 commonsourceibias.t64 168.701
R72 commonsourceibias.n279 commonsourceibias.t104 168.701
R73 commonsourceibias.n277 commonsourceibias.t68 168.701
R74 commonsourceibias.n275 commonsourceibias.t79 168.701
R75 commonsourceibias.n299 commonsourceibias.t56 168.701
R76 commonsourceibias.n484 commonsourceibias.t97 168.701
R77 commonsourceibias.n481 commonsourceibias.t78 168.701
R78 commonsourceibias.n479 commonsourceibias.t53 168.701
R79 commonsourceibias.n477 commonsourceibias.t62 168.701
R80 commonsourceibias.n501 commonsourceibias.t82 168.701
R81 commonsourceibias.n507 commonsourceibias.t85 168.701
R82 commonsourceibias.n509 commonsourceibias.t74 168.701
R83 commonsourceibias.n516 commonsourceibias.t101 168.701
R84 commonsourceibias.n522 commonsourceibias.t91 168.701
R85 commonsourceibias.n469 commonsourceibias.t81 168.701
R86 commonsourceibias.n420 commonsourceibias.t61 168.701
R87 commonsourceibias.n417 commonsourceibias.t75 168.701
R88 commonsourceibias.n415 commonsourceibias.t55 168.701
R89 commonsourceibias.n413 commonsourceibias.t105 168.701
R90 commonsourceibias.n437 commonsourceibias.t76 168.701
R91 commonsourceibias.n443 commonsourceibias.t50 168.701
R92 commonsourceibias.n445 commonsourceibias.t106 168.701
R93 commonsourceibias.n452 commonsourceibias.t114 168.701
R94 commonsourceibias.n458 commonsourceibias.t51 168.701
R95 commonsourceibias.n405 commonsourceibias.t107 168.701
R96 commonsourceibias.n27 commonsourceibias.n24 161.3
R97 commonsourceibias.n29 commonsourceibias.n28 161.3
R98 commonsourceibias.n31 commonsourceibias.n30 161.3
R99 commonsourceibias.n32 commonsourceibias.n22 161.3
R100 commonsourceibias.n34 commonsourceibias.n33 161.3
R101 commonsourceibias.n36 commonsourceibias.n35 161.3
R102 commonsourceibias.n37 commonsourceibias.n20 161.3
R103 commonsourceibias.n39 commonsourceibias.n38 161.3
R104 commonsourceibias.n41 commonsourceibias.n40 161.3
R105 commonsourceibias.n42 commonsourceibias.n18 161.3
R106 commonsourceibias.n45 commonsourceibias.n44 161.3
R107 commonsourceibias.n46 commonsourceibias.n17 161.3
R108 commonsourceibias.n48 commonsourceibias.n47 161.3
R109 commonsourceibias.n50 commonsourceibias.n15 161.3
R110 commonsourceibias.n52 commonsourceibias.n51 161.3
R111 commonsourceibias.n53 commonsourceibias.n14 161.3
R112 commonsourceibias.n55 commonsourceibias.n54 161.3
R113 commonsourceibias.n56 commonsourceibias.n13 161.3
R114 commonsourceibias.n59 commonsourceibias.n58 161.3
R115 commonsourceibias.n60 commonsourceibias.n12 161.3
R116 commonsourceibias.n62 commonsourceibias.n61 161.3
R117 commonsourceibias.n64 commonsourceibias.n11 161.3
R118 commonsourceibias.n66 commonsourceibias.n65 161.3
R119 commonsourceibias.n68 commonsourceibias.n67 161.3
R120 commonsourceibias.n69 commonsourceibias.n9 161.3
R121 commonsourceibias.n93 commonsourceibias.n90 161.3
R122 commonsourceibias.n95 commonsourceibias.n94 161.3
R123 commonsourceibias.n97 commonsourceibias.n96 161.3
R124 commonsourceibias.n98 commonsourceibias.n88 161.3
R125 commonsourceibias.n100 commonsourceibias.n99 161.3
R126 commonsourceibias.n102 commonsourceibias.n101 161.3
R127 commonsourceibias.n103 commonsourceibias.n86 161.3
R128 commonsourceibias.n105 commonsourceibias.n104 161.3
R129 commonsourceibias.n107 commonsourceibias.n106 161.3
R130 commonsourceibias.n108 commonsourceibias.n84 161.3
R131 commonsourceibias.n111 commonsourceibias.n110 161.3
R132 commonsourceibias.n112 commonsourceibias.n8 161.3
R133 commonsourceibias.n114 commonsourceibias.n113 161.3
R134 commonsourceibias.n116 commonsourceibias.n6 161.3
R135 commonsourceibias.n118 commonsourceibias.n117 161.3
R136 commonsourceibias.n119 commonsourceibias.n5 161.3
R137 commonsourceibias.n121 commonsourceibias.n120 161.3
R138 commonsourceibias.n122 commonsourceibias.n4 161.3
R139 commonsourceibias.n125 commonsourceibias.n124 161.3
R140 commonsourceibias.n126 commonsourceibias.n3 161.3
R141 commonsourceibias.n128 commonsourceibias.n127 161.3
R142 commonsourceibias.n130 commonsourceibias.n2 161.3
R143 commonsourceibias.n132 commonsourceibias.n131 161.3
R144 commonsourceibias.n134 commonsourceibias.n133 161.3
R145 commonsourceibias.n135 commonsourceibias.n0 161.3
R146 commonsourceibias.n262 commonsourceibias.n202 161.3
R147 commonsourceibias.n261 commonsourceibias.n260 161.3
R148 commonsourceibias.n259 commonsourceibias.n258 161.3
R149 commonsourceibias.n257 commonsourceibias.n204 161.3
R150 commonsourceibias.n255 commonsourceibias.n254 161.3
R151 commonsourceibias.n253 commonsourceibias.n205 161.3
R152 commonsourceibias.n252 commonsourceibias.n251 161.3
R153 commonsourceibias.n249 commonsourceibias.n206 161.3
R154 commonsourceibias.n248 commonsourceibias.n247 161.3
R155 commonsourceibias.n246 commonsourceibias.n207 161.3
R156 commonsourceibias.n245 commonsourceibias.n244 161.3
R157 commonsourceibias.n243 commonsourceibias.n208 161.3
R158 commonsourceibias.n241 commonsourceibias.n240 161.3
R159 commonsourceibias.n239 commonsourceibias.n210 161.3
R160 commonsourceibias.n238 commonsourceibias.n237 161.3
R161 commonsourceibias.n235 commonsourceibias.n211 161.3
R162 commonsourceibias.n234 commonsourceibias.n233 161.3
R163 commonsourceibias.n232 commonsourceibias.n231 161.3
R164 commonsourceibias.n230 commonsourceibias.n213 161.3
R165 commonsourceibias.n229 commonsourceibias.n228 161.3
R166 commonsourceibias.n227 commonsourceibias.n226 161.3
R167 commonsourceibias.n225 commonsourceibias.n215 161.3
R168 commonsourceibias.n224 commonsourceibias.n223 161.3
R169 commonsourceibias.n222 commonsourceibias.n221 161.3
R170 commonsourceibias.n220 commonsourceibias.n217 161.3
R171 commonsourceibias.n156 commonsourceibias.n153 161.3
R172 commonsourceibias.n158 commonsourceibias.n157 161.3
R173 commonsourceibias.n160 commonsourceibias.n159 161.3
R174 commonsourceibias.n161 commonsourceibias.n151 161.3
R175 commonsourceibias.n163 commonsourceibias.n162 161.3
R176 commonsourceibias.n165 commonsourceibias.n164 161.3
R177 commonsourceibias.n166 commonsourceibias.n149 161.3
R178 commonsourceibias.n168 commonsourceibias.n167 161.3
R179 commonsourceibias.n170 commonsourceibias.n169 161.3
R180 commonsourceibias.n171 commonsourceibias.n147 161.3
R181 commonsourceibias.n174 commonsourceibias.n173 161.3
R182 commonsourceibias.n175 commonsourceibias.n146 161.3
R183 commonsourceibias.n177 commonsourceibias.n176 161.3
R184 commonsourceibias.n179 commonsourceibias.n144 161.3
R185 commonsourceibias.n181 commonsourceibias.n180 161.3
R186 commonsourceibias.n182 commonsourceibias.n143 161.3
R187 commonsourceibias.n184 commonsourceibias.n183 161.3
R188 commonsourceibias.n185 commonsourceibias.n142 161.3
R189 commonsourceibias.n188 commonsourceibias.n187 161.3
R190 commonsourceibias.n189 commonsourceibias.n141 161.3
R191 commonsourceibias.n191 commonsourceibias.n190 161.3
R192 commonsourceibias.n193 commonsourceibias.n140 161.3
R193 commonsourceibias.n195 commonsourceibias.n194 161.3
R194 commonsourceibias.n197 commonsourceibias.n196 161.3
R195 commonsourceibias.n198 commonsourceibias.n138 161.3
R196 commonsourceibias.n367 commonsourceibias.n307 161.3
R197 commonsourceibias.n366 commonsourceibias.n365 161.3
R198 commonsourceibias.n364 commonsourceibias.n363 161.3
R199 commonsourceibias.n362 commonsourceibias.n309 161.3
R200 commonsourceibias.n360 commonsourceibias.n359 161.3
R201 commonsourceibias.n358 commonsourceibias.n310 161.3
R202 commonsourceibias.n357 commonsourceibias.n356 161.3
R203 commonsourceibias.n354 commonsourceibias.n311 161.3
R204 commonsourceibias.n353 commonsourceibias.n352 161.3
R205 commonsourceibias.n351 commonsourceibias.n312 161.3
R206 commonsourceibias.n350 commonsourceibias.n349 161.3
R207 commonsourceibias.n347 commonsourceibias.n313 161.3
R208 commonsourceibias.n345 commonsourceibias.n344 161.3
R209 commonsourceibias.n343 commonsourceibias.n314 161.3
R210 commonsourceibias.n342 commonsourceibias.n341 161.3
R211 commonsourceibias.n339 commonsourceibias.n315 161.3
R212 commonsourceibias.n338 commonsourceibias.n337 161.3
R213 commonsourceibias.n336 commonsourceibias.n335 161.3
R214 commonsourceibias.n334 commonsourceibias.n317 161.3
R215 commonsourceibias.n333 commonsourceibias.n332 161.3
R216 commonsourceibias.n331 commonsourceibias.n330 161.3
R217 commonsourceibias.n329 commonsourceibias.n319 161.3
R218 commonsourceibias.n328 commonsourceibias.n327 161.3
R219 commonsourceibias.n326 commonsourceibias.n325 161.3
R220 commonsourceibias.n324 commonsourceibias.n321 161.3
R221 commonsourceibias.n301 commonsourceibias.n300 161.3
R222 commonsourceibias.n298 commonsourceibias.n274 161.3
R223 commonsourceibias.n297 commonsourceibias.n296 161.3
R224 commonsourceibias.n295 commonsourceibias.n294 161.3
R225 commonsourceibias.n293 commonsourceibias.n276 161.3
R226 commonsourceibias.n292 commonsourceibias.n291 161.3
R227 commonsourceibias.n290 commonsourceibias.n289 161.3
R228 commonsourceibias.n288 commonsourceibias.n278 161.3
R229 commonsourceibias.n287 commonsourceibias.n286 161.3
R230 commonsourceibias.n285 commonsourceibias.n284 161.3
R231 commonsourceibias.n283 commonsourceibias.n280 161.3
R232 commonsourceibias.n377 commonsourceibias.n273 161.3
R233 commonsourceibias.n401 commonsourceibias.n266 161.3
R234 commonsourceibias.n400 commonsourceibias.n399 161.3
R235 commonsourceibias.n398 commonsourceibias.n397 161.3
R236 commonsourceibias.n396 commonsourceibias.n268 161.3
R237 commonsourceibias.n394 commonsourceibias.n393 161.3
R238 commonsourceibias.n392 commonsourceibias.n269 161.3
R239 commonsourceibias.n391 commonsourceibias.n390 161.3
R240 commonsourceibias.n388 commonsourceibias.n270 161.3
R241 commonsourceibias.n387 commonsourceibias.n386 161.3
R242 commonsourceibias.n385 commonsourceibias.n271 161.3
R243 commonsourceibias.n384 commonsourceibias.n383 161.3
R244 commonsourceibias.n381 commonsourceibias.n272 161.3
R245 commonsourceibias.n379 commonsourceibias.n378 161.3
R246 commonsourceibias.n528 commonsourceibias.n468 161.3
R247 commonsourceibias.n527 commonsourceibias.n526 161.3
R248 commonsourceibias.n525 commonsourceibias.n524 161.3
R249 commonsourceibias.n523 commonsourceibias.n470 161.3
R250 commonsourceibias.n521 commonsourceibias.n520 161.3
R251 commonsourceibias.n519 commonsourceibias.n471 161.3
R252 commonsourceibias.n518 commonsourceibias.n517 161.3
R253 commonsourceibias.n515 commonsourceibias.n472 161.3
R254 commonsourceibias.n514 commonsourceibias.n513 161.3
R255 commonsourceibias.n512 commonsourceibias.n473 161.3
R256 commonsourceibias.n511 commonsourceibias.n510 161.3
R257 commonsourceibias.n508 commonsourceibias.n474 161.3
R258 commonsourceibias.n506 commonsourceibias.n505 161.3
R259 commonsourceibias.n504 commonsourceibias.n475 161.3
R260 commonsourceibias.n503 commonsourceibias.n502 161.3
R261 commonsourceibias.n500 commonsourceibias.n476 161.3
R262 commonsourceibias.n499 commonsourceibias.n498 161.3
R263 commonsourceibias.n497 commonsourceibias.n496 161.3
R264 commonsourceibias.n495 commonsourceibias.n478 161.3
R265 commonsourceibias.n494 commonsourceibias.n493 161.3
R266 commonsourceibias.n492 commonsourceibias.n491 161.3
R267 commonsourceibias.n490 commonsourceibias.n480 161.3
R268 commonsourceibias.n489 commonsourceibias.n488 161.3
R269 commonsourceibias.n487 commonsourceibias.n486 161.3
R270 commonsourceibias.n485 commonsourceibias.n482 161.3
R271 commonsourceibias.n464 commonsourceibias.n404 161.3
R272 commonsourceibias.n463 commonsourceibias.n462 161.3
R273 commonsourceibias.n461 commonsourceibias.n460 161.3
R274 commonsourceibias.n459 commonsourceibias.n406 161.3
R275 commonsourceibias.n457 commonsourceibias.n456 161.3
R276 commonsourceibias.n455 commonsourceibias.n407 161.3
R277 commonsourceibias.n454 commonsourceibias.n453 161.3
R278 commonsourceibias.n451 commonsourceibias.n408 161.3
R279 commonsourceibias.n450 commonsourceibias.n449 161.3
R280 commonsourceibias.n448 commonsourceibias.n409 161.3
R281 commonsourceibias.n447 commonsourceibias.n446 161.3
R282 commonsourceibias.n444 commonsourceibias.n410 161.3
R283 commonsourceibias.n442 commonsourceibias.n441 161.3
R284 commonsourceibias.n440 commonsourceibias.n411 161.3
R285 commonsourceibias.n439 commonsourceibias.n438 161.3
R286 commonsourceibias.n436 commonsourceibias.n412 161.3
R287 commonsourceibias.n435 commonsourceibias.n434 161.3
R288 commonsourceibias.n433 commonsourceibias.n432 161.3
R289 commonsourceibias.n431 commonsourceibias.n414 161.3
R290 commonsourceibias.n430 commonsourceibias.n429 161.3
R291 commonsourceibias.n428 commonsourceibias.n427 161.3
R292 commonsourceibias.n426 commonsourceibias.n416 161.3
R293 commonsourceibias.n425 commonsourceibias.n424 161.3
R294 commonsourceibias.n423 commonsourceibias.n422 161.3
R295 commonsourceibias.n421 commonsourceibias.n418 161.3
R296 commonsourceibias.n80 commonsourceibias.n78 81.5057
R297 commonsourceibias.n304 commonsourceibias.n302 81.5057
R298 commonsourceibias.n80 commonsourceibias.n79 80.9324
R299 commonsourceibias.n82 commonsourceibias.n81 80.9324
R300 commonsourceibias.n77 commonsourceibias.n76 80.9324
R301 commonsourceibias.n75 commonsourceibias.n74 80.9324
R302 commonsourceibias.n73 commonsourceibias.n72 80.9324
R303 commonsourceibias.n371 commonsourceibias.n370 80.9324
R304 commonsourceibias.n373 commonsourceibias.n372 80.9324
R305 commonsourceibias.n375 commonsourceibias.n374 80.9324
R306 commonsourceibias.n306 commonsourceibias.n305 80.9324
R307 commonsourceibias.n304 commonsourceibias.n303 80.9324
R308 commonsourceibias.n71 commonsourceibias.n70 80.6037
R309 commonsourceibias.n137 commonsourceibias.n136 80.6037
R310 commonsourceibias.n264 commonsourceibias.n263 80.6037
R311 commonsourceibias.n200 commonsourceibias.n199 80.6037
R312 commonsourceibias.n369 commonsourceibias.n368 80.6037
R313 commonsourceibias.n403 commonsourceibias.n402 80.6037
R314 commonsourceibias.n530 commonsourceibias.n529 80.6037
R315 commonsourceibias.n466 commonsourceibias.n465 80.6037
R316 commonsourceibias.n65 commonsourceibias.n64 56.5617
R317 commonsourceibias.n51 commonsourceibias.n50 56.5617
R318 commonsourceibias.n42 commonsourceibias.n41 56.5617
R319 commonsourceibias.n28 commonsourceibias.n27 56.5617
R320 commonsourceibias.n131 commonsourceibias.n130 56.5617
R321 commonsourceibias.n117 commonsourceibias.n116 56.5617
R322 commonsourceibias.n108 commonsourceibias.n107 56.5617
R323 commonsourceibias.n94 commonsourceibias.n93 56.5617
R324 commonsourceibias.n221 commonsourceibias.n220 56.5617
R325 commonsourceibias.n235 commonsourceibias.n234 56.5617
R326 commonsourceibias.n244 commonsourceibias.n243 56.5617
R327 commonsourceibias.n258 commonsourceibias.n257 56.5617
R328 commonsourceibias.n194 commonsourceibias.n193 56.5617
R329 commonsourceibias.n180 commonsourceibias.n179 56.5617
R330 commonsourceibias.n171 commonsourceibias.n170 56.5617
R331 commonsourceibias.n157 commonsourceibias.n156 56.5617
R332 commonsourceibias.n325 commonsourceibias.n324 56.5617
R333 commonsourceibias.n339 commonsourceibias.n338 56.5617
R334 commonsourceibias.n349 commonsourceibias.n347 56.5617
R335 commonsourceibias.n363 commonsourceibias.n362 56.5617
R336 commonsourceibias.n397 commonsourceibias.n396 56.5617
R337 commonsourceibias.n383 commonsourceibias.n381 56.5617
R338 commonsourceibias.n284 commonsourceibias.n283 56.5617
R339 commonsourceibias.n298 commonsourceibias.n297 56.5617
R340 commonsourceibias.n486 commonsourceibias.n485 56.5617
R341 commonsourceibias.n500 commonsourceibias.n499 56.5617
R342 commonsourceibias.n510 commonsourceibias.n508 56.5617
R343 commonsourceibias.n524 commonsourceibias.n523 56.5617
R344 commonsourceibias.n422 commonsourceibias.n421 56.5617
R345 commonsourceibias.n436 commonsourceibias.n435 56.5617
R346 commonsourceibias.n446 commonsourceibias.n444 56.5617
R347 commonsourceibias.n460 commonsourceibias.n459 56.5617
R348 commonsourceibias.n56 commonsourceibias.n55 56.0773
R349 commonsourceibias.n37 commonsourceibias.n36 56.0773
R350 commonsourceibias.n122 commonsourceibias.n121 56.0773
R351 commonsourceibias.n103 commonsourceibias.n102 56.0773
R352 commonsourceibias.n230 commonsourceibias.n229 56.0773
R353 commonsourceibias.n249 commonsourceibias.n248 56.0773
R354 commonsourceibias.n185 commonsourceibias.n184 56.0773
R355 commonsourceibias.n166 commonsourceibias.n165 56.0773
R356 commonsourceibias.n334 commonsourceibias.n333 56.0773
R357 commonsourceibias.n354 commonsourceibias.n353 56.0773
R358 commonsourceibias.n388 commonsourceibias.n387 56.0773
R359 commonsourceibias.n293 commonsourceibias.n292 56.0773
R360 commonsourceibias.n495 commonsourceibias.n494 56.0773
R361 commonsourceibias.n515 commonsourceibias.n514 56.0773
R362 commonsourceibias.n431 commonsourceibias.n430 56.0773
R363 commonsourceibias.n451 commonsourceibias.n450 56.0773
R364 commonsourceibias.n70 commonsourceibias.n69 46.0096
R365 commonsourceibias.n136 commonsourceibias.n135 46.0096
R366 commonsourceibias.n263 commonsourceibias.n262 46.0096
R367 commonsourceibias.n199 commonsourceibias.n198 46.0096
R368 commonsourceibias.n368 commonsourceibias.n367 46.0096
R369 commonsourceibias.n402 commonsourceibias.n401 46.0096
R370 commonsourceibias.n529 commonsourceibias.n528 46.0096
R371 commonsourceibias.n465 commonsourceibias.n464 46.0096
R372 commonsourceibias.n58 commonsourceibias.n12 41.5458
R373 commonsourceibias.n33 commonsourceibias.n32 41.5458
R374 commonsourceibias.n124 commonsourceibias.n3 41.5458
R375 commonsourceibias.n99 commonsourceibias.n98 41.5458
R376 commonsourceibias.n226 commonsourceibias.n225 41.5458
R377 commonsourceibias.n251 commonsourceibias.n205 41.5458
R378 commonsourceibias.n187 commonsourceibias.n141 41.5458
R379 commonsourceibias.n162 commonsourceibias.n161 41.5458
R380 commonsourceibias.n330 commonsourceibias.n329 41.5458
R381 commonsourceibias.n356 commonsourceibias.n310 41.5458
R382 commonsourceibias.n390 commonsourceibias.n269 41.5458
R383 commonsourceibias.n289 commonsourceibias.n288 41.5458
R384 commonsourceibias.n491 commonsourceibias.n490 41.5458
R385 commonsourceibias.n517 commonsourceibias.n471 41.5458
R386 commonsourceibias.n427 commonsourceibias.n426 41.5458
R387 commonsourceibias.n453 commonsourceibias.n407 41.5458
R388 commonsourceibias.n48 commonsourceibias.n17 40.577
R389 commonsourceibias.n44 commonsourceibias.n17 40.577
R390 commonsourceibias.n114 commonsourceibias.n8 40.577
R391 commonsourceibias.n110 commonsourceibias.n8 40.577
R392 commonsourceibias.n237 commonsourceibias.n210 40.577
R393 commonsourceibias.n241 commonsourceibias.n210 40.577
R394 commonsourceibias.n177 commonsourceibias.n146 40.577
R395 commonsourceibias.n173 commonsourceibias.n146 40.577
R396 commonsourceibias.n341 commonsourceibias.n314 40.577
R397 commonsourceibias.n345 commonsourceibias.n314 40.577
R398 commonsourceibias.n379 commonsourceibias.n273 40.577
R399 commonsourceibias.n300 commonsourceibias.n273 40.577
R400 commonsourceibias.n502 commonsourceibias.n475 40.577
R401 commonsourceibias.n506 commonsourceibias.n475 40.577
R402 commonsourceibias.n438 commonsourceibias.n411 40.577
R403 commonsourceibias.n442 commonsourceibias.n411 40.577
R404 commonsourceibias.n62 commonsourceibias.n12 39.6083
R405 commonsourceibias.n32 commonsourceibias.n31 39.6083
R406 commonsourceibias.n128 commonsourceibias.n3 39.6083
R407 commonsourceibias.n98 commonsourceibias.n97 39.6083
R408 commonsourceibias.n225 commonsourceibias.n224 39.6083
R409 commonsourceibias.n255 commonsourceibias.n205 39.6083
R410 commonsourceibias.n191 commonsourceibias.n141 39.6083
R411 commonsourceibias.n161 commonsourceibias.n160 39.6083
R412 commonsourceibias.n329 commonsourceibias.n328 39.6083
R413 commonsourceibias.n360 commonsourceibias.n310 39.6083
R414 commonsourceibias.n394 commonsourceibias.n269 39.6083
R415 commonsourceibias.n288 commonsourceibias.n287 39.6083
R416 commonsourceibias.n490 commonsourceibias.n489 39.6083
R417 commonsourceibias.n521 commonsourceibias.n471 39.6083
R418 commonsourceibias.n426 commonsourceibias.n425 39.6083
R419 commonsourceibias.n457 commonsourceibias.n407 39.6083
R420 commonsourceibias.n26 commonsourceibias.n25 33.0515
R421 commonsourceibias.n92 commonsourceibias.n91 33.0515
R422 commonsourceibias.n155 commonsourceibias.n154 33.0515
R423 commonsourceibias.n219 commonsourceibias.n218 33.0515
R424 commonsourceibias.n323 commonsourceibias.n322 33.0515
R425 commonsourceibias.n282 commonsourceibias.n281 33.0515
R426 commonsourceibias.n484 commonsourceibias.n483 33.0515
R427 commonsourceibias.n420 commonsourceibias.n419 33.0515
R428 commonsourceibias.n25 commonsourceibias.n24 28.5514
R429 commonsourceibias.n91 commonsourceibias.n90 28.5514
R430 commonsourceibias.n218 commonsourceibias.n217 28.5514
R431 commonsourceibias.n154 commonsourceibias.n153 28.5514
R432 commonsourceibias.n322 commonsourceibias.n321 28.5514
R433 commonsourceibias.n281 commonsourceibias.n280 28.5514
R434 commonsourceibias.n483 commonsourceibias.n482 28.5514
R435 commonsourceibias.n419 commonsourceibias.n418 28.5514
R436 commonsourceibias.n69 commonsourceibias.n68 26.0455
R437 commonsourceibias.n135 commonsourceibias.n134 26.0455
R438 commonsourceibias.n262 commonsourceibias.n261 26.0455
R439 commonsourceibias.n198 commonsourceibias.n197 26.0455
R440 commonsourceibias.n367 commonsourceibias.n366 26.0455
R441 commonsourceibias.n401 commonsourceibias.n400 26.0455
R442 commonsourceibias.n528 commonsourceibias.n527 26.0455
R443 commonsourceibias.n464 commonsourceibias.n463 26.0455
R444 commonsourceibias.n55 commonsourceibias.n14 25.0767
R445 commonsourceibias.n38 commonsourceibias.n37 25.0767
R446 commonsourceibias.n121 commonsourceibias.n5 25.0767
R447 commonsourceibias.n104 commonsourceibias.n103 25.0767
R448 commonsourceibias.n231 commonsourceibias.n230 25.0767
R449 commonsourceibias.n248 commonsourceibias.n207 25.0767
R450 commonsourceibias.n184 commonsourceibias.n143 25.0767
R451 commonsourceibias.n167 commonsourceibias.n166 25.0767
R452 commonsourceibias.n335 commonsourceibias.n334 25.0767
R453 commonsourceibias.n353 commonsourceibias.n312 25.0767
R454 commonsourceibias.n387 commonsourceibias.n271 25.0767
R455 commonsourceibias.n294 commonsourceibias.n293 25.0767
R456 commonsourceibias.n496 commonsourceibias.n495 25.0767
R457 commonsourceibias.n514 commonsourceibias.n473 25.0767
R458 commonsourceibias.n432 commonsourceibias.n431 25.0767
R459 commonsourceibias.n450 commonsourceibias.n409 25.0767
R460 commonsourceibias.n51 commonsourceibias.n16 24.3464
R461 commonsourceibias.n41 commonsourceibias.n19 24.3464
R462 commonsourceibias.n117 commonsourceibias.n7 24.3464
R463 commonsourceibias.n107 commonsourceibias.n85 24.3464
R464 commonsourceibias.n234 commonsourceibias.n212 24.3464
R465 commonsourceibias.n244 commonsourceibias.n209 24.3464
R466 commonsourceibias.n180 commonsourceibias.n145 24.3464
R467 commonsourceibias.n170 commonsourceibias.n148 24.3464
R468 commonsourceibias.n338 commonsourceibias.n316 24.3464
R469 commonsourceibias.n349 commonsourceibias.n348 24.3464
R470 commonsourceibias.n383 commonsourceibias.n382 24.3464
R471 commonsourceibias.n297 commonsourceibias.n275 24.3464
R472 commonsourceibias.n499 commonsourceibias.n477 24.3464
R473 commonsourceibias.n510 commonsourceibias.n509 24.3464
R474 commonsourceibias.n435 commonsourceibias.n413 24.3464
R475 commonsourceibias.n446 commonsourceibias.n445 24.3464
R476 commonsourceibias.n65 commonsourceibias.n10 23.8546
R477 commonsourceibias.n27 commonsourceibias.n26 23.8546
R478 commonsourceibias.n131 commonsourceibias.n1 23.8546
R479 commonsourceibias.n93 commonsourceibias.n92 23.8546
R480 commonsourceibias.n220 commonsourceibias.n219 23.8546
R481 commonsourceibias.n258 commonsourceibias.n203 23.8546
R482 commonsourceibias.n194 commonsourceibias.n139 23.8546
R483 commonsourceibias.n156 commonsourceibias.n155 23.8546
R484 commonsourceibias.n324 commonsourceibias.n323 23.8546
R485 commonsourceibias.n363 commonsourceibias.n308 23.8546
R486 commonsourceibias.n397 commonsourceibias.n267 23.8546
R487 commonsourceibias.n283 commonsourceibias.n282 23.8546
R488 commonsourceibias.n485 commonsourceibias.n484 23.8546
R489 commonsourceibias.n524 commonsourceibias.n469 23.8546
R490 commonsourceibias.n421 commonsourceibias.n420 23.8546
R491 commonsourceibias.n460 commonsourceibias.n405 23.8546
R492 commonsourceibias.n64 commonsourceibias.n63 16.9689
R493 commonsourceibias.n28 commonsourceibias.n23 16.9689
R494 commonsourceibias.n130 commonsourceibias.n129 16.9689
R495 commonsourceibias.n94 commonsourceibias.n89 16.9689
R496 commonsourceibias.n221 commonsourceibias.n216 16.9689
R497 commonsourceibias.n257 commonsourceibias.n256 16.9689
R498 commonsourceibias.n193 commonsourceibias.n192 16.9689
R499 commonsourceibias.n157 commonsourceibias.n152 16.9689
R500 commonsourceibias.n325 commonsourceibias.n320 16.9689
R501 commonsourceibias.n362 commonsourceibias.n361 16.9689
R502 commonsourceibias.n396 commonsourceibias.n395 16.9689
R503 commonsourceibias.n284 commonsourceibias.n279 16.9689
R504 commonsourceibias.n486 commonsourceibias.n481 16.9689
R505 commonsourceibias.n523 commonsourceibias.n522 16.9689
R506 commonsourceibias.n422 commonsourceibias.n417 16.9689
R507 commonsourceibias.n459 commonsourceibias.n458 16.9689
R508 commonsourceibias.n50 commonsourceibias.n49 16.477
R509 commonsourceibias.n43 commonsourceibias.n42 16.477
R510 commonsourceibias.n116 commonsourceibias.n115 16.477
R511 commonsourceibias.n109 commonsourceibias.n108 16.477
R512 commonsourceibias.n236 commonsourceibias.n235 16.477
R513 commonsourceibias.n243 commonsourceibias.n242 16.477
R514 commonsourceibias.n179 commonsourceibias.n178 16.477
R515 commonsourceibias.n172 commonsourceibias.n171 16.477
R516 commonsourceibias.n340 commonsourceibias.n339 16.477
R517 commonsourceibias.n347 commonsourceibias.n346 16.477
R518 commonsourceibias.n381 commonsourceibias.n380 16.477
R519 commonsourceibias.n299 commonsourceibias.n298 16.477
R520 commonsourceibias.n501 commonsourceibias.n500 16.477
R521 commonsourceibias.n508 commonsourceibias.n507 16.477
R522 commonsourceibias.n437 commonsourceibias.n436 16.477
R523 commonsourceibias.n444 commonsourceibias.n443 16.477
R524 commonsourceibias.n57 commonsourceibias.n56 15.9852
R525 commonsourceibias.n36 commonsourceibias.n21 15.9852
R526 commonsourceibias.n123 commonsourceibias.n122 15.9852
R527 commonsourceibias.n102 commonsourceibias.n87 15.9852
R528 commonsourceibias.n229 commonsourceibias.n214 15.9852
R529 commonsourceibias.n250 commonsourceibias.n249 15.9852
R530 commonsourceibias.n186 commonsourceibias.n185 15.9852
R531 commonsourceibias.n165 commonsourceibias.n150 15.9852
R532 commonsourceibias.n333 commonsourceibias.n318 15.9852
R533 commonsourceibias.n355 commonsourceibias.n354 15.9852
R534 commonsourceibias.n389 commonsourceibias.n388 15.9852
R535 commonsourceibias.n292 commonsourceibias.n277 15.9852
R536 commonsourceibias.n494 commonsourceibias.n479 15.9852
R537 commonsourceibias.n516 commonsourceibias.n515 15.9852
R538 commonsourceibias.n430 commonsourceibias.n415 15.9852
R539 commonsourceibias.n452 commonsourceibias.n451 15.9852
R540 commonsourceibias.n73 commonsourceibias.n71 13.2057
R541 commonsourceibias.n371 commonsourceibias.n369 13.2057
R542 commonsourceibias.n532 commonsourceibias.n265 10.122
R543 commonsourceibias.n112 commonsourceibias.n83 9.50363
R544 commonsourceibias.n377 commonsourceibias.n376 9.50363
R545 commonsourceibias.n201 commonsourceibias.n137 8.7339
R546 commonsourceibias.n467 commonsourceibias.n403 8.7339
R547 commonsourceibias.n58 commonsourceibias.n57 8.60764
R548 commonsourceibias.n33 commonsourceibias.n21 8.60764
R549 commonsourceibias.n124 commonsourceibias.n123 8.60764
R550 commonsourceibias.n99 commonsourceibias.n87 8.60764
R551 commonsourceibias.n226 commonsourceibias.n214 8.60764
R552 commonsourceibias.n251 commonsourceibias.n250 8.60764
R553 commonsourceibias.n187 commonsourceibias.n186 8.60764
R554 commonsourceibias.n162 commonsourceibias.n150 8.60764
R555 commonsourceibias.n330 commonsourceibias.n318 8.60764
R556 commonsourceibias.n356 commonsourceibias.n355 8.60764
R557 commonsourceibias.n390 commonsourceibias.n389 8.60764
R558 commonsourceibias.n289 commonsourceibias.n277 8.60764
R559 commonsourceibias.n491 commonsourceibias.n479 8.60764
R560 commonsourceibias.n517 commonsourceibias.n516 8.60764
R561 commonsourceibias.n427 commonsourceibias.n415 8.60764
R562 commonsourceibias.n453 commonsourceibias.n452 8.60764
R563 commonsourceibias.n532 commonsourceibias.n531 8.46921
R564 commonsourceibias.n49 commonsourceibias.n48 8.11581
R565 commonsourceibias.n44 commonsourceibias.n43 8.11581
R566 commonsourceibias.n115 commonsourceibias.n114 8.11581
R567 commonsourceibias.n110 commonsourceibias.n109 8.11581
R568 commonsourceibias.n237 commonsourceibias.n236 8.11581
R569 commonsourceibias.n242 commonsourceibias.n241 8.11581
R570 commonsourceibias.n178 commonsourceibias.n177 8.11581
R571 commonsourceibias.n173 commonsourceibias.n172 8.11581
R572 commonsourceibias.n341 commonsourceibias.n340 8.11581
R573 commonsourceibias.n346 commonsourceibias.n345 8.11581
R574 commonsourceibias.n380 commonsourceibias.n379 8.11581
R575 commonsourceibias.n300 commonsourceibias.n299 8.11581
R576 commonsourceibias.n502 commonsourceibias.n501 8.11581
R577 commonsourceibias.n507 commonsourceibias.n506 8.11581
R578 commonsourceibias.n438 commonsourceibias.n437 8.11581
R579 commonsourceibias.n443 commonsourceibias.n442 8.11581
R580 commonsourceibias.n63 commonsourceibias.n62 7.62397
R581 commonsourceibias.n31 commonsourceibias.n23 7.62397
R582 commonsourceibias.n129 commonsourceibias.n128 7.62397
R583 commonsourceibias.n97 commonsourceibias.n89 7.62397
R584 commonsourceibias.n224 commonsourceibias.n216 7.62397
R585 commonsourceibias.n256 commonsourceibias.n255 7.62397
R586 commonsourceibias.n192 commonsourceibias.n191 7.62397
R587 commonsourceibias.n160 commonsourceibias.n152 7.62397
R588 commonsourceibias.n328 commonsourceibias.n320 7.62397
R589 commonsourceibias.n361 commonsourceibias.n360 7.62397
R590 commonsourceibias.n395 commonsourceibias.n394 7.62397
R591 commonsourceibias.n287 commonsourceibias.n279 7.62397
R592 commonsourceibias.n489 commonsourceibias.n481 7.62397
R593 commonsourceibias.n522 commonsourceibias.n521 7.62397
R594 commonsourceibias.n425 commonsourceibias.n417 7.62397
R595 commonsourceibias.n458 commonsourceibias.n457 7.62397
R596 commonsourceibias.n265 commonsourceibias.n264 5.00473
R597 commonsourceibias.n201 commonsourceibias.n200 5.00473
R598 commonsourceibias.n531 commonsourceibias.n530 5.00473
R599 commonsourceibias.n467 commonsourceibias.n466 5.00473
R600 commonsourceibias commonsourceibias.n532 3.87639
R601 commonsourceibias.n265 commonsourceibias.n201 3.72967
R602 commonsourceibias.n531 commonsourceibias.n467 3.72967
R603 commonsourceibias.n78 commonsourceibias.t5 2.82907
R604 commonsourceibias.n78 commonsourceibias.t11 2.82907
R605 commonsourceibias.n79 commonsourceibias.t25 2.82907
R606 commonsourceibias.n79 commonsourceibias.t35 2.82907
R607 commonsourceibias.n81 commonsourceibias.t9 2.82907
R608 commonsourceibias.n81 commonsourceibias.t41 2.82907
R609 commonsourceibias.n76 commonsourceibias.t45 2.82907
R610 commonsourceibias.n76 commonsourceibias.t19 2.82907
R611 commonsourceibias.n74 commonsourceibias.t39 2.82907
R612 commonsourceibias.n74 commonsourceibias.t21 2.82907
R613 commonsourceibias.n72 commonsourceibias.t23 2.82907
R614 commonsourceibias.n72 commonsourceibias.t1 2.82907
R615 commonsourceibias.n370 commonsourceibias.t47 2.82907
R616 commonsourceibias.n370 commonsourceibias.t15 2.82907
R617 commonsourceibias.n372 commonsourceibias.t13 2.82907
R618 commonsourceibias.n372 commonsourceibias.t29 2.82907
R619 commonsourceibias.n374 commonsourceibias.t31 2.82907
R620 commonsourceibias.n374 commonsourceibias.t43 2.82907
R621 commonsourceibias.n305 commonsourceibias.t7 2.82907
R622 commonsourceibias.n305 commonsourceibias.t37 2.82907
R623 commonsourceibias.n303 commonsourceibias.t27 2.82907
R624 commonsourceibias.n303 commonsourceibias.t17 2.82907
R625 commonsourceibias.n302 commonsourceibias.t3 2.82907
R626 commonsourceibias.n302 commonsourceibias.t33 2.82907
R627 commonsourceibias.n68 commonsourceibias.n10 0.738255
R628 commonsourceibias.n134 commonsourceibias.n1 0.738255
R629 commonsourceibias.n261 commonsourceibias.n203 0.738255
R630 commonsourceibias.n197 commonsourceibias.n139 0.738255
R631 commonsourceibias.n366 commonsourceibias.n308 0.738255
R632 commonsourceibias.n400 commonsourceibias.n267 0.738255
R633 commonsourceibias.n527 commonsourceibias.n469 0.738255
R634 commonsourceibias.n463 commonsourceibias.n405 0.738255
R635 commonsourceibias.n75 commonsourceibias.n73 0.573776
R636 commonsourceibias.n77 commonsourceibias.n75 0.573776
R637 commonsourceibias.n82 commonsourceibias.n80 0.573776
R638 commonsourceibias.n306 commonsourceibias.n304 0.573776
R639 commonsourceibias.n375 commonsourceibias.n373 0.573776
R640 commonsourceibias.n373 commonsourceibias.n371 0.573776
R641 commonsourceibias.n83 commonsourceibias.n77 0.287138
R642 commonsourceibias.n83 commonsourceibias.n82 0.287138
R643 commonsourceibias.n376 commonsourceibias.n306 0.287138
R644 commonsourceibias.n376 commonsourceibias.n375 0.287138
R645 commonsourceibias.n71 commonsourceibias.n9 0.285035
R646 commonsourceibias.n137 commonsourceibias.n0 0.285035
R647 commonsourceibias.n264 commonsourceibias.n202 0.285035
R648 commonsourceibias.n200 commonsourceibias.n138 0.285035
R649 commonsourceibias.n369 commonsourceibias.n307 0.285035
R650 commonsourceibias.n403 commonsourceibias.n266 0.285035
R651 commonsourceibias.n530 commonsourceibias.n468 0.285035
R652 commonsourceibias.n466 commonsourceibias.n404 0.285035
R653 commonsourceibias.n16 commonsourceibias.n14 0.246418
R654 commonsourceibias.n38 commonsourceibias.n19 0.246418
R655 commonsourceibias.n7 commonsourceibias.n5 0.246418
R656 commonsourceibias.n104 commonsourceibias.n85 0.246418
R657 commonsourceibias.n231 commonsourceibias.n212 0.246418
R658 commonsourceibias.n209 commonsourceibias.n207 0.246418
R659 commonsourceibias.n145 commonsourceibias.n143 0.246418
R660 commonsourceibias.n167 commonsourceibias.n148 0.246418
R661 commonsourceibias.n335 commonsourceibias.n316 0.246418
R662 commonsourceibias.n348 commonsourceibias.n312 0.246418
R663 commonsourceibias.n382 commonsourceibias.n271 0.246418
R664 commonsourceibias.n294 commonsourceibias.n275 0.246418
R665 commonsourceibias.n496 commonsourceibias.n477 0.246418
R666 commonsourceibias.n509 commonsourceibias.n473 0.246418
R667 commonsourceibias.n432 commonsourceibias.n413 0.246418
R668 commonsourceibias.n445 commonsourceibias.n409 0.246418
R669 commonsourceibias.n67 commonsourceibias.n9 0.189894
R670 commonsourceibias.n67 commonsourceibias.n66 0.189894
R671 commonsourceibias.n66 commonsourceibias.n11 0.189894
R672 commonsourceibias.n61 commonsourceibias.n11 0.189894
R673 commonsourceibias.n61 commonsourceibias.n60 0.189894
R674 commonsourceibias.n60 commonsourceibias.n59 0.189894
R675 commonsourceibias.n59 commonsourceibias.n13 0.189894
R676 commonsourceibias.n54 commonsourceibias.n13 0.189894
R677 commonsourceibias.n54 commonsourceibias.n53 0.189894
R678 commonsourceibias.n53 commonsourceibias.n52 0.189894
R679 commonsourceibias.n52 commonsourceibias.n15 0.189894
R680 commonsourceibias.n47 commonsourceibias.n15 0.189894
R681 commonsourceibias.n47 commonsourceibias.n46 0.189894
R682 commonsourceibias.n46 commonsourceibias.n45 0.189894
R683 commonsourceibias.n45 commonsourceibias.n18 0.189894
R684 commonsourceibias.n40 commonsourceibias.n18 0.189894
R685 commonsourceibias.n40 commonsourceibias.n39 0.189894
R686 commonsourceibias.n39 commonsourceibias.n20 0.189894
R687 commonsourceibias.n35 commonsourceibias.n20 0.189894
R688 commonsourceibias.n35 commonsourceibias.n34 0.189894
R689 commonsourceibias.n34 commonsourceibias.n22 0.189894
R690 commonsourceibias.n30 commonsourceibias.n22 0.189894
R691 commonsourceibias.n30 commonsourceibias.n29 0.189894
R692 commonsourceibias.n29 commonsourceibias.n24 0.189894
R693 commonsourceibias.n111 commonsourceibias.n84 0.189894
R694 commonsourceibias.n106 commonsourceibias.n84 0.189894
R695 commonsourceibias.n106 commonsourceibias.n105 0.189894
R696 commonsourceibias.n105 commonsourceibias.n86 0.189894
R697 commonsourceibias.n101 commonsourceibias.n86 0.189894
R698 commonsourceibias.n101 commonsourceibias.n100 0.189894
R699 commonsourceibias.n100 commonsourceibias.n88 0.189894
R700 commonsourceibias.n96 commonsourceibias.n88 0.189894
R701 commonsourceibias.n96 commonsourceibias.n95 0.189894
R702 commonsourceibias.n95 commonsourceibias.n90 0.189894
R703 commonsourceibias.n133 commonsourceibias.n0 0.189894
R704 commonsourceibias.n133 commonsourceibias.n132 0.189894
R705 commonsourceibias.n132 commonsourceibias.n2 0.189894
R706 commonsourceibias.n127 commonsourceibias.n2 0.189894
R707 commonsourceibias.n127 commonsourceibias.n126 0.189894
R708 commonsourceibias.n126 commonsourceibias.n125 0.189894
R709 commonsourceibias.n125 commonsourceibias.n4 0.189894
R710 commonsourceibias.n120 commonsourceibias.n4 0.189894
R711 commonsourceibias.n120 commonsourceibias.n119 0.189894
R712 commonsourceibias.n119 commonsourceibias.n118 0.189894
R713 commonsourceibias.n118 commonsourceibias.n6 0.189894
R714 commonsourceibias.n113 commonsourceibias.n6 0.189894
R715 commonsourceibias.n260 commonsourceibias.n202 0.189894
R716 commonsourceibias.n260 commonsourceibias.n259 0.189894
R717 commonsourceibias.n259 commonsourceibias.n204 0.189894
R718 commonsourceibias.n254 commonsourceibias.n204 0.189894
R719 commonsourceibias.n254 commonsourceibias.n253 0.189894
R720 commonsourceibias.n253 commonsourceibias.n252 0.189894
R721 commonsourceibias.n252 commonsourceibias.n206 0.189894
R722 commonsourceibias.n247 commonsourceibias.n206 0.189894
R723 commonsourceibias.n247 commonsourceibias.n246 0.189894
R724 commonsourceibias.n246 commonsourceibias.n245 0.189894
R725 commonsourceibias.n245 commonsourceibias.n208 0.189894
R726 commonsourceibias.n240 commonsourceibias.n208 0.189894
R727 commonsourceibias.n240 commonsourceibias.n239 0.189894
R728 commonsourceibias.n239 commonsourceibias.n238 0.189894
R729 commonsourceibias.n238 commonsourceibias.n211 0.189894
R730 commonsourceibias.n233 commonsourceibias.n211 0.189894
R731 commonsourceibias.n233 commonsourceibias.n232 0.189894
R732 commonsourceibias.n232 commonsourceibias.n213 0.189894
R733 commonsourceibias.n228 commonsourceibias.n213 0.189894
R734 commonsourceibias.n228 commonsourceibias.n227 0.189894
R735 commonsourceibias.n227 commonsourceibias.n215 0.189894
R736 commonsourceibias.n223 commonsourceibias.n215 0.189894
R737 commonsourceibias.n223 commonsourceibias.n222 0.189894
R738 commonsourceibias.n222 commonsourceibias.n217 0.189894
R739 commonsourceibias.n196 commonsourceibias.n138 0.189894
R740 commonsourceibias.n196 commonsourceibias.n195 0.189894
R741 commonsourceibias.n195 commonsourceibias.n140 0.189894
R742 commonsourceibias.n190 commonsourceibias.n140 0.189894
R743 commonsourceibias.n190 commonsourceibias.n189 0.189894
R744 commonsourceibias.n189 commonsourceibias.n188 0.189894
R745 commonsourceibias.n188 commonsourceibias.n142 0.189894
R746 commonsourceibias.n183 commonsourceibias.n142 0.189894
R747 commonsourceibias.n183 commonsourceibias.n182 0.189894
R748 commonsourceibias.n182 commonsourceibias.n181 0.189894
R749 commonsourceibias.n181 commonsourceibias.n144 0.189894
R750 commonsourceibias.n176 commonsourceibias.n144 0.189894
R751 commonsourceibias.n176 commonsourceibias.n175 0.189894
R752 commonsourceibias.n175 commonsourceibias.n174 0.189894
R753 commonsourceibias.n174 commonsourceibias.n147 0.189894
R754 commonsourceibias.n169 commonsourceibias.n147 0.189894
R755 commonsourceibias.n169 commonsourceibias.n168 0.189894
R756 commonsourceibias.n168 commonsourceibias.n149 0.189894
R757 commonsourceibias.n164 commonsourceibias.n149 0.189894
R758 commonsourceibias.n164 commonsourceibias.n163 0.189894
R759 commonsourceibias.n163 commonsourceibias.n151 0.189894
R760 commonsourceibias.n159 commonsourceibias.n151 0.189894
R761 commonsourceibias.n159 commonsourceibias.n158 0.189894
R762 commonsourceibias.n158 commonsourceibias.n153 0.189894
R763 commonsourceibias.n326 commonsourceibias.n321 0.189894
R764 commonsourceibias.n327 commonsourceibias.n326 0.189894
R765 commonsourceibias.n327 commonsourceibias.n319 0.189894
R766 commonsourceibias.n331 commonsourceibias.n319 0.189894
R767 commonsourceibias.n332 commonsourceibias.n331 0.189894
R768 commonsourceibias.n332 commonsourceibias.n317 0.189894
R769 commonsourceibias.n336 commonsourceibias.n317 0.189894
R770 commonsourceibias.n337 commonsourceibias.n336 0.189894
R771 commonsourceibias.n337 commonsourceibias.n315 0.189894
R772 commonsourceibias.n342 commonsourceibias.n315 0.189894
R773 commonsourceibias.n343 commonsourceibias.n342 0.189894
R774 commonsourceibias.n344 commonsourceibias.n343 0.189894
R775 commonsourceibias.n344 commonsourceibias.n313 0.189894
R776 commonsourceibias.n350 commonsourceibias.n313 0.189894
R777 commonsourceibias.n351 commonsourceibias.n350 0.189894
R778 commonsourceibias.n352 commonsourceibias.n351 0.189894
R779 commonsourceibias.n352 commonsourceibias.n311 0.189894
R780 commonsourceibias.n357 commonsourceibias.n311 0.189894
R781 commonsourceibias.n358 commonsourceibias.n357 0.189894
R782 commonsourceibias.n359 commonsourceibias.n358 0.189894
R783 commonsourceibias.n359 commonsourceibias.n309 0.189894
R784 commonsourceibias.n364 commonsourceibias.n309 0.189894
R785 commonsourceibias.n365 commonsourceibias.n364 0.189894
R786 commonsourceibias.n365 commonsourceibias.n307 0.189894
R787 commonsourceibias.n285 commonsourceibias.n280 0.189894
R788 commonsourceibias.n286 commonsourceibias.n285 0.189894
R789 commonsourceibias.n286 commonsourceibias.n278 0.189894
R790 commonsourceibias.n290 commonsourceibias.n278 0.189894
R791 commonsourceibias.n291 commonsourceibias.n290 0.189894
R792 commonsourceibias.n291 commonsourceibias.n276 0.189894
R793 commonsourceibias.n295 commonsourceibias.n276 0.189894
R794 commonsourceibias.n296 commonsourceibias.n295 0.189894
R795 commonsourceibias.n296 commonsourceibias.n274 0.189894
R796 commonsourceibias.n301 commonsourceibias.n274 0.189894
R797 commonsourceibias.n378 commonsourceibias.n272 0.189894
R798 commonsourceibias.n384 commonsourceibias.n272 0.189894
R799 commonsourceibias.n385 commonsourceibias.n384 0.189894
R800 commonsourceibias.n386 commonsourceibias.n385 0.189894
R801 commonsourceibias.n386 commonsourceibias.n270 0.189894
R802 commonsourceibias.n391 commonsourceibias.n270 0.189894
R803 commonsourceibias.n392 commonsourceibias.n391 0.189894
R804 commonsourceibias.n393 commonsourceibias.n392 0.189894
R805 commonsourceibias.n393 commonsourceibias.n268 0.189894
R806 commonsourceibias.n398 commonsourceibias.n268 0.189894
R807 commonsourceibias.n399 commonsourceibias.n398 0.189894
R808 commonsourceibias.n399 commonsourceibias.n266 0.189894
R809 commonsourceibias.n487 commonsourceibias.n482 0.189894
R810 commonsourceibias.n488 commonsourceibias.n487 0.189894
R811 commonsourceibias.n488 commonsourceibias.n480 0.189894
R812 commonsourceibias.n492 commonsourceibias.n480 0.189894
R813 commonsourceibias.n493 commonsourceibias.n492 0.189894
R814 commonsourceibias.n493 commonsourceibias.n478 0.189894
R815 commonsourceibias.n497 commonsourceibias.n478 0.189894
R816 commonsourceibias.n498 commonsourceibias.n497 0.189894
R817 commonsourceibias.n498 commonsourceibias.n476 0.189894
R818 commonsourceibias.n503 commonsourceibias.n476 0.189894
R819 commonsourceibias.n504 commonsourceibias.n503 0.189894
R820 commonsourceibias.n505 commonsourceibias.n504 0.189894
R821 commonsourceibias.n505 commonsourceibias.n474 0.189894
R822 commonsourceibias.n511 commonsourceibias.n474 0.189894
R823 commonsourceibias.n512 commonsourceibias.n511 0.189894
R824 commonsourceibias.n513 commonsourceibias.n512 0.189894
R825 commonsourceibias.n513 commonsourceibias.n472 0.189894
R826 commonsourceibias.n518 commonsourceibias.n472 0.189894
R827 commonsourceibias.n519 commonsourceibias.n518 0.189894
R828 commonsourceibias.n520 commonsourceibias.n519 0.189894
R829 commonsourceibias.n520 commonsourceibias.n470 0.189894
R830 commonsourceibias.n525 commonsourceibias.n470 0.189894
R831 commonsourceibias.n526 commonsourceibias.n525 0.189894
R832 commonsourceibias.n526 commonsourceibias.n468 0.189894
R833 commonsourceibias.n423 commonsourceibias.n418 0.189894
R834 commonsourceibias.n424 commonsourceibias.n423 0.189894
R835 commonsourceibias.n424 commonsourceibias.n416 0.189894
R836 commonsourceibias.n428 commonsourceibias.n416 0.189894
R837 commonsourceibias.n429 commonsourceibias.n428 0.189894
R838 commonsourceibias.n429 commonsourceibias.n414 0.189894
R839 commonsourceibias.n433 commonsourceibias.n414 0.189894
R840 commonsourceibias.n434 commonsourceibias.n433 0.189894
R841 commonsourceibias.n434 commonsourceibias.n412 0.189894
R842 commonsourceibias.n439 commonsourceibias.n412 0.189894
R843 commonsourceibias.n440 commonsourceibias.n439 0.189894
R844 commonsourceibias.n441 commonsourceibias.n440 0.189894
R845 commonsourceibias.n441 commonsourceibias.n410 0.189894
R846 commonsourceibias.n447 commonsourceibias.n410 0.189894
R847 commonsourceibias.n448 commonsourceibias.n447 0.189894
R848 commonsourceibias.n449 commonsourceibias.n448 0.189894
R849 commonsourceibias.n449 commonsourceibias.n408 0.189894
R850 commonsourceibias.n454 commonsourceibias.n408 0.189894
R851 commonsourceibias.n455 commonsourceibias.n454 0.189894
R852 commonsourceibias.n456 commonsourceibias.n455 0.189894
R853 commonsourceibias.n456 commonsourceibias.n406 0.189894
R854 commonsourceibias.n461 commonsourceibias.n406 0.189894
R855 commonsourceibias.n462 commonsourceibias.n461 0.189894
R856 commonsourceibias.n462 commonsourceibias.n404 0.189894
R857 commonsourceibias.n112 commonsourceibias.n111 0.170955
R858 commonsourceibias.n113 commonsourceibias.n112 0.170955
R859 commonsourceibias.n377 commonsourceibias.n301 0.170955
R860 commonsourceibias.n378 commonsourceibias.n377 0.170955
R861 gnd.n6510 gnd.n687 1087.89
R862 gnd.n4071 gnd.n3735 939.716
R863 gnd.n6840 gnd.n166 838.452
R864 gnd.n198 gnd.n164 838.452
R865 gnd.n1558 gnd.n1446 838.452
R866 gnd.n5531 gnd.n1560 838.452
R867 gnd.n1145 gnd.n1133 838.452
R868 gnd.n4571 gnd.n4570 838.452
R869 gnd.n3911 gnd.n3772 838.452
R870 gnd.n3950 gnd.n2263 838.452
R871 gnd.n6842 gnd.n161 783.196
R872 gnd.n490 gnd.n163 783.196
R873 gnd.n5534 gnd.n5533 783.196
R874 gnd.n5651 gnd.n1492 783.196
R875 gnd.n5957 gnd.n1138 783.196
R876 gnd.n4520 gnd.n2126 783.196
R877 gnd.n4074 gnd.n4073 783.196
R878 gnd.n4069 gnd.n2259 783.196
R879 gnd.n4298 gnd.n4297 771.183
R880 gnd.n5720 gnd.n1382 771.183
R881 gnd.n4578 gnd.n2095 771.183
R882 gnd.n5722 gnd.n1377 771.183
R883 gnd.n3643 gnd.n2274 766.379
R884 gnd.n3646 gnd.n3645 766.379
R885 gnd.n2884 gnd.n2787 766.379
R886 gnd.n2880 gnd.n2785 766.379
R887 gnd.n3734 gnd.n2296 756.769
R888 gnd.n3637 gnd.n3636 756.769
R889 gnd.n2977 gnd.n2694 756.769
R890 gnd.n2975 gnd.n2697 756.769
R891 gnd.n6182 gnd.n879 655.866
R892 gnd.n6509 gnd.n688 655.866
R893 gnd.n6722 gnd.n6721 655.866
R894 gnd.n6014 gnd.n1049 655.866
R895 gnd.n6183 gnd.n6182 585
R896 gnd.n6182 gnd.n6181 585
R897 gnd.n883 gnd.n882 585
R898 gnd.n6180 gnd.n883 585
R899 gnd.n6178 gnd.n6177 585
R900 gnd.n6179 gnd.n6178 585
R901 gnd.n6176 gnd.n885 585
R902 gnd.n885 gnd.n884 585
R903 gnd.n6175 gnd.n6174 585
R904 gnd.n6174 gnd.n6173 585
R905 gnd.n890 gnd.n889 585
R906 gnd.n6172 gnd.n890 585
R907 gnd.n6170 gnd.n6169 585
R908 gnd.n6171 gnd.n6170 585
R909 gnd.n6168 gnd.n892 585
R910 gnd.n892 gnd.n891 585
R911 gnd.n6167 gnd.n6166 585
R912 gnd.n6166 gnd.n6165 585
R913 gnd.n898 gnd.n897 585
R914 gnd.n6164 gnd.n898 585
R915 gnd.n6162 gnd.n6161 585
R916 gnd.n6163 gnd.n6162 585
R917 gnd.n6160 gnd.n900 585
R918 gnd.n900 gnd.n899 585
R919 gnd.n6159 gnd.n6158 585
R920 gnd.n6158 gnd.n6157 585
R921 gnd.n906 gnd.n905 585
R922 gnd.n6156 gnd.n906 585
R923 gnd.n6154 gnd.n6153 585
R924 gnd.n6155 gnd.n6154 585
R925 gnd.n6152 gnd.n908 585
R926 gnd.n908 gnd.n907 585
R927 gnd.n6151 gnd.n6150 585
R928 gnd.n6150 gnd.n6149 585
R929 gnd.n914 gnd.n913 585
R930 gnd.n6148 gnd.n914 585
R931 gnd.n6146 gnd.n6145 585
R932 gnd.n6147 gnd.n6146 585
R933 gnd.n6144 gnd.n916 585
R934 gnd.n916 gnd.n915 585
R935 gnd.n6143 gnd.n6142 585
R936 gnd.n6142 gnd.n6141 585
R937 gnd.n922 gnd.n921 585
R938 gnd.n6140 gnd.n922 585
R939 gnd.n6138 gnd.n6137 585
R940 gnd.n6139 gnd.n6138 585
R941 gnd.n6136 gnd.n924 585
R942 gnd.n924 gnd.n923 585
R943 gnd.n6135 gnd.n6134 585
R944 gnd.n6134 gnd.n6133 585
R945 gnd.n930 gnd.n929 585
R946 gnd.n6132 gnd.n930 585
R947 gnd.n6130 gnd.n6129 585
R948 gnd.n6131 gnd.n6130 585
R949 gnd.n6128 gnd.n932 585
R950 gnd.n932 gnd.n931 585
R951 gnd.n6127 gnd.n6126 585
R952 gnd.n6126 gnd.n6125 585
R953 gnd.n938 gnd.n937 585
R954 gnd.n6124 gnd.n938 585
R955 gnd.n6122 gnd.n6121 585
R956 gnd.n6123 gnd.n6122 585
R957 gnd.n6120 gnd.n940 585
R958 gnd.n940 gnd.n939 585
R959 gnd.n6119 gnd.n6118 585
R960 gnd.n6118 gnd.n6117 585
R961 gnd.n946 gnd.n945 585
R962 gnd.n6116 gnd.n946 585
R963 gnd.n6114 gnd.n6113 585
R964 gnd.n6115 gnd.n6114 585
R965 gnd.n6112 gnd.n948 585
R966 gnd.n948 gnd.n947 585
R967 gnd.n6111 gnd.n6110 585
R968 gnd.n6110 gnd.n6109 585
R969 gnd.n954 gnd.n953 585
R970 gnd.n6108 gnd.n954 585
R971 gnd.n6106 gnd.n6105 585
R972 gnd.n6107 gnd.n6106 585
R973 gnd.n6104 gnd.n956 585
R974 gnd.n956 gnd.n955 585
R975 gnd.n6103 gnd.n6102 585
R976 gnd.n6102 gnd.n6101 585
R977 gnd.n962 gnd.n961 585
R978 gnd.n6100 gnd.n962 585
R979 gnd.n6098 gnd.n6097 585
R980 gnd.n6099 gnd.n6098 585
R981 gnd.n6096 gnd.n964 585
R982 gnd.n964 gnd.n963 585
R983 gnd.n6095 gnd.n6094 585
R984 gnd.n6094 gnd.n6093 585
R985 gnd.n970 gnd.n969 585
R986 gnd.n6092 gnd.n970 585
R987 gnd.n6090 gnd.n6089 585
R988 gnd.n6091 gnd.n6090 585
R989 gnd.n6088 gnd.n972 585
R990 gnd.n972 gnd.n971 585
R991 gnd.n6087 gnd.n6086 585
R992 gnd.n6086 gnd.n6085 585
R993 gnd.n978 gnd.n977 585
R994 gnd.n6084 gnd.n978 585
R995 gnd.n6082 gnd.n6081 585
R996 gnd.n6083 gnd.n6082 585
R997 gnd.n6080 gnd.n980 585
R998 gnd.n980 gnd.n979 585
R999 gnd.n6079 gnd.n6078 585
R1000 gnd.n6078 gnd.n6077 585
R1001 gnd.n986 gnd.n985 585
R1002 gnd.n6076 gnd.n986 585
R1003 gnd.n6074 gnd.n6073 585
R1004 gnd.n6075 gnd.n6074 585
R1005 gnd.n6072 gnd.n988 585
R1006 gnd.n988 gnd.n987 585
R1007 gnd.n6071 gnd.n6070 585
R1008 gnd.n6070 gnd.n6069 585
R1009 gnd.n994 gnd.n993 585
R1010 gnd.n6068 gnd.n994 585
R1011 gnd.n6066 gnd.n6065 585
R1012 gnd.n6067 gnd.n6066 585
R1013 gnd.n6064 gnd.n996 585
R1014 gnd.n996 gnd.n995 585
R1015 gnd.n6063 gnd.n6062 585
R1016 gnd.n6062 gnd.n6061 585
R1017 gnd.n1002 gnd.n1001 585
R1018 gnd.n6060 gnd.n1002 585
R1019 gnd.n6058 gnd.n6057 585
R1020 gnd.n6059 gnd.n6058 585
R1021 gnd.n6056 gnd.n1004 585
R1022 gnd.n1004 gnd.n1003 585
R1023 gnd.n6055 gnd.n6054 585
R1024 gnd.n6054 gnd.n6053 585
R1025 gnd.n1010 gnd.n1009 585
R1026 gnd.n6052 gnd.n1010 585
R1027 gnd.n6050 gnd.n6049 585
R1028 gnd.n6051 gnd.n6050 585
R1029 gnd.n6048 gnd.n1012 585
R1030 gnd.n1012 gnd.n1011 585
R1031 gnd.n6047 gnd.n6046 585
R1032 gnd.n6046 gnd.n6045 585
R1033 gnd.n1018 gnd.n1017 585
R1034 gnd.n6044 gnd.n1018 585
R1035 gnd.n6042 gnd.n6041 585
R1036 gnd.n6043 gnd.n6042 585
R1037 gnd.n6040 gnd.n1020 585
R1038 gnd.n1020 gnd.n1019 585
R1039 gnd.n6039 gnd.n6038 585
R1040 gnd.n6038 gnd.n6037 585
R1041 gnd.n1026 gnd.n1025 585
R1042 gnd.n6036 gnd.n1026 585
R1043 gnd.n6034 gnd.n6033 585
R1044 gnd.n6035 gnd.n6034 585
R1045 gnd.n6032 gnd.n1028 585
R1046 gnd.n1028 gnd.n1027 585
R1047 gnd.n6031 gnd.n6030 585
R1048 gnd.n6030 gnd.n6029 585
R1049 gnd.n1034 gnd.n1033 585
R1050 gnd.n6028 gnd.n1034 585
R1051 gnd.n6026 gnd.n6025 585
R1052 gnd.n6027 gnd.n6026 585
R1053 gnd.n6024 gnd.n1036 585
R1054 gnd.n1036 gnd.n1035 585
R1055 gnd.n6023 gnd.n6022 585
R1056 gnd.n6022 gnd.n6021 585
R1057 gnd.n1042 gnd.n1041 585
R1058 gnd.n6020 gnd.n1042 585
R1059 gnd.n6018 gnd.n6017 585
R1060 gnd.n6019 gnd.n6018 585
R1061 gnd.n6016 gnd.n1044 585
R1062 gnd.n1044 gnd.n1043 585
R1063 gnd.n880 gnd.n879 585
R1064 gnd.n879 gnd.n878 585
R1065 gnd.n6188 gnd.n6187 585
R1066 gnd.n6189 gnd.n6188 585
R1067 gnd.n877 gnd.n876 585
R1068 gnd.n6190 gnd.n877 585
R1069 gnd.n6193 gnd.n6192 585
R1070 gnd.n6192 gnd.n6191 585
R1071 gnd.n874 gnd.n873 585
R1072 gnd.n873 gnd.n872 585
R1073 gnd.n6198 gnd.n6197 585
R1074 gnd.n6199 gnd.n6198 585
R1075 gnd.n871 gnd.n870 585
R1076 gnd.n6200 gnd.n871 585
R1077 gnd.n6203 gnd.n6202 585
R1078 gnd.n6202 gnd.n6201 585
R1079 gnd.n868 gnd.n867 585
R1080 gnd.n867 gnd.n866 585
R1081 gnd.n6208 gnd.n6207 585
R1082 gnd.n6209 gnd.n6208 585
R1083 gnd.n865 gnd.n864 585
R1084 gnd.n6210 gnd.n865 585
R1085 gnd.n6213 gnd.n6212 585
R1086 gnd.n6212 gnd.n6211 585
R1087 gnd.n862 gnd.n861 585
R1088 gnd.n861 gnd.n860 585
R1089 gnd.n6218 gnd.n6217 585
R1090 gnd.n6219 gnd.n6218 585
R1091 gnd.n859 gnd.n858 585
R1092 gnd.n6220 gnd.n859 585
R1093 gnd.n6223 gnd.n6222 585
R1094 gnd.n6222 gnd.n6221 585
R1095 gnd.n856 gnd.n855 585
R1096 gnd.n855 gnd.n854 585
R1097 gnd.n6228 gnd.n6227 585
R1098 gnd.n6229 gnd.n6228 585
R1099 gnd.n853 gnd.n852 585
R1100 gnd.n6230 gnd.n853 585
R1101 gnd.n6233 gnd.n6232 585
R1102 gnd.n6232 gnd.n6231 585
R1103 gnd.n850 gnd.n849 585
R1104 gnd.n849 gnd.n848 585
R1105 gnd.n6238 gnd.n6237 585
R1106 gnd.n6239 gnd.n6238 585
R1107 gnd.n847 gnd.n846 585
R1108 gnd.n6240 gnd.n847 585
R1109 gnd.n6243 gnd.n6242 585
R1110 gnd.n6242 gnd.n6241 585
R1111 gnd.n844 gnd.n843 585
R1112 gnd.n843 gnd.n842 585
R1113 gnd.n6248 gnd.n6247 585
R1114 gnd.n6249 gnd.n6248 585
R1115 gnd.n841 gnd.n840 585
R1116 gnd.n6250 gnd.n841 585
R1117 gnd.n6253 gnd.n6252 585
R1118 gnd.n6252 gnd.n6251 585
R1119 gnd.n838 gnd.n837 585
R1120 gnd.n837 gnd.n836 585
R1121 gnd.n6258 gnd.n6257 585
R1122 gnd.n6259 gnd.n6258 585
R1123 gnd.n835 gnd.n834 585
R1124 gnd.n6260 gnd.n835 585
R1125 gnd.n6263 gnd.n6262 585
R1126 gnd.n6262 gnd.n6261 585
R1127 gnd.n832 gnd.n831 585
R1128 gnd.n831 gnd.n830 585
R1129 gnd.n6268 gnd.n6267 585
R1130 gnd.n6269 gnd.n6268 585
R1131 gnd.n829 gnd.n828 585
R1132 gnd.n6270 gnd.n829 585
R1133 gnd.n6273 gnd.n6272 585
R1134 gnd.n6272 gnd.n6271 585
R1135 gnd.n826 gnd.n825 585
R1136 gnd.n825 gnd.n824 585
R1137 gnd.n6278 gnd.n6277 585
R1138 gnd.n6279 gnd.n6278 585
R1139 gnd.n823 gnd.n822 585
R1140 gnd.n6280 gnd.n823 585
R1141 gnd.n6283 gnd.n6282 585
R1142 gnd.n6282 gnd.n6281 585
R1143 gnd.n820 gnd.n819 585
R1144 gnd.n819 gnd.n818 585
R1145 gnd.n6288 gnd.n6287 585
R1146 gnd.n6289 gnd.n6288 585
R1147 gnd.n817 gnd.n816 585
R1148 gnd.n6290 gnd.n817 585
R1149 gnd.n6293 gnd.n6292 585
R1150 gnd.n6292 gnd.n6291 585
R1151 gnd.n814 gnd.n813 585
R1152 gnd.n813 gnd.n812 585
R1153 gnd.n6298 gnd.n6297 585
R1154 gnd.n6299 gnd.n6298 585
R1155 gnd.n811 gnd.n810 585
R1156 gnd.n6300 gnd.n811 585
R1157 gnd.n6303 gnd.n6302 585
R1158 gnd.n6302 gnd.n6301 585
R1159 gnd.n808 gnd.n807 585
R1160 gnd.n807 gnd.n806 585
R1161 gnd.n6308 gnd.n6307 585
R1162 gnd.n6309 gnd.n6308 585
R1163 gnd.n805 gnd.n804 585
R1164 gnd.n6310 gnd.n805 585
R1165 gnd.n6313 gnd.n6312 585
R1166 gnd.n6312 gnd.n6311 585
R1167 gnd.n802 gnd.n801 585
R1168 gnd.n801 gnd.n800 585
R1169 gnd.n6318 gnd.n6317 585
R1170 gnd.n6319 gnd.n6318 585
R1171 gnd.n799 gnd.n798 585
R1172 gnd.n6320 gnd.n799 585
R1173 gnd.n6323 gnd.n6322 585
R1174 gnd.n6322 gnd.n6321 585
R1175 gnd.n796 gnd.n795 585
R1176 gnd.n795 gnd.n794 585
R1177 gnd.n6328 gnd.n6327 585
R1178 gnd.n6329 gnd.n6328 585
R1179 gnd.n793 gnd.n792 585
R1180 gnd.n6330 gnd.n793 585
R1181 gnd.n6333 gnd.n6332 585
R1182 gnd.n6332 gnd.n6331 585
R1183 gnd.n790 gnd.n789 585
R1184 gnd.n789 gnd.n788 585
R1185 gnd.n6338 gnd.n6337 585
R1186 gnd.n6339 gnd.n6338 585
R1187 gnd.n787 gnd.n786 585
R1188 gnd.n6340 gnd.n787 585
R1189 gnd.n6343 gnd.n6342 585
R1190 gnd.n6342 gnd.n6341 585
R1191 gnd.n784 gnd.n783 585
R1192 gnd.n783 gnd.n782 585
R1193 gnd.n6348 gnd.n6347 585
R1194 gnd.n6349 gnd.n6348 585
R1195 gnd.n781 gnd.n780 585
R1196 gnd.n6350 gnd.n781 585
R1197 gnd.n6353 gnd.n6352 585
R1198 gnd.n6352 gnd.n6351 585
R1199 gnd.n778 gnd.n777 585
R1200 gnd.n777 gnd.n776 585
R1201 gnd.n6358 gnd.n6357 585
R1202 gnd.n6359 gnd.n6358 585
R1203 gnd.n775 gnd.n774 585
R1204 gnd.n6360 gnd.n775 585
R1205 gnd.n6363 gnd.n6362 585
R1206 gnd.n6362 gnd.n6361 585
R1207 gnd.n772 gnd.n771 585
R1208 gnd.n771 gnd.n770 585
R1209 gnd.n6368 gnd.n6367 585
R1210 gnd.n6369 gnd.n6368 585
R1211 gnd.n769 gnd.n768 585
R1212 gnd.n6370 gnd.n769 585
R1213 gnd.n6373 gnd.n6372 585
R1214 gnd.n6372 gnd.n6371 585
R1215 gnd.n766 gnd.n765 585
R1216 gnd.n765 gnd.n764 585
R1217 gnd.n6378 gnd.n6377 585
R1218 gnd.n6379 gnd.n6378 585
R1219 gnd.n763 gnd.n762 585
R1220 gnd.n6380 gnd.n763 585
R1221 gnd.n6383 gnd.n6382 585
R1222 gnd.n6382 gnd.n6381 585
R1223 gnd.n760 gnd.n759 585
R1224 gnd.n759 gnd.n758 585
R1225 gnd.n6388 gnd.n6387 585
R1226 gnd.n6389 gnd.n6388 585
R1227 gnd.n757 gnd.n756 585
R1228 gnd.n6390 gnd.n757 585
R1229 gnd.n6393 gnd.n6392 585
R1230 gnd.n6392 gnd.n6391 585
R1231 gnd.n754 gnd.n753 585
R1232 gnd.n753 gnd.n752 585
R1233 gnd.n6398 gnd.n6397 585
R1234 gnd.n6399 gnd.n6398 585
R1235 gnd.n751 gnd.n750 585
R1236 gnd.n6400 gnd.n751 585
R1237 gnd.n6403 gnd.n6402 585
R1238 gnd.n6402 gnd.n6401 585
R1239 gnd.n748 gnd.n747 585
R1240 gnd.n747 gnd.n746 585
R1241 gnd.n6408 gnd.n6407 585
R1242 gnd.n6409 gnd.n6408 585
R1243 gnd.n745 gnd.n744 585
R1244 gnd.n6410 gnd.n745 585
R1245 gnd.n6413 gnd.n6412 585
R1246 gnd.n6412 gnd.n6411 585
R1247 gnd.n742 gnd.n741 585
R1248 gnd.n741 gnd.n740 585
R1249 gnd.n6418 gnd.n6417 585
R1250 gnd.n6419 gnd.n6418 585
R1251 gnd.n739 gnd.n738 585
R1252 gnd.n6420 gnd.n739 585
R1253 gnd.n6423 gnd.n6422 585
R1254 gnd.n6422 gnd.n6421 585
R1255 gnd.n736 gnd.n735 585
R1256 gnd.n735 gnd.n734 585
R1257 gnd.n6428 gnd.n6427 585
R1258 gnd.n6429 gnd.n6428 585
R1259 gnd.n733 gnd.n732 585
R1260 gnd.n6430 gnd.n733 585
R1261 gnd.n6433 gnd.n6432 585
R1262 gnd.n6432 gnd.n6431 585
R1263 gnd.n730 gnd.n729 585
R1264 gnd.n729 gnd.n728 585
R1265 gnd.n6438 gnd.n6437 585
R1266 gnd.n6439 gnd.n6438 585
R1267 gnd.n727 gnd.n726 585
R1268 gnd.n6440 gnd.n727 585
R1269 gnd.n6443 gnd.n6442 585
R1270 gnd.n6442 gnd.n6441 585
R1271 gnd.n724 gnd.n723 585
R1272 gnd.n723 gnd.n722 585
R1273 gnd.n6448 gnd.n6447 585
R1274 gnd.n6449 gnd.n6448 585
R1275 gnd.n721 gnd.n720 585
R1276 gnd.n6450 gnd.n721 585
R1277 gnd.n6453 gnd.n6452 585
R1278 gnd.n6452 gnd.n6451 585
R1279 gnd.n718 gnd.n717 585
R1280 gnd.n717 gnd.n716 585
R1281 gnd.n6458 gnd.n6457 585
R1282 gnd.n6459 gnd.n6458 585
R1283 gnd.n715 gnd.n714 585
R1284 gnd.n6460 gnd.n715 585
R1285 gnd.n6463 gnd.n6462 585
R1286 gnd.n6462 gnd.n6461 585
R1287 gnd.n712 gnd.n711 585
R1288 gnd.n711 gnd.n710 585
R1289 gnd.n6468 gnd.n6467 585
R1290 gnd.n6469 gnd.n6468 585
R1291 gnd.n709 gnd.n708 585
R1292 gnd.n6470 gnd.n709 585
R1293 gnd.n6473 gnd.n6472 585
R1294 gnd.n6472 gnd.n6471 585
R1295 gnd.n706 gnd.n705 585
R1296 gnd.n705 gnd.n704 585
R1297 gnd.n6478 gnd.n6477 585
R1298 gnd.n6479 gnd.n6478 585
R1299 gnd.n703 gnd.n702 585
R1300 gnd.n6480 gnd.n703 585
R1301 gnd.n6483 gnd.n6482 585
R1302 gnd.n6482 gnd.n6481 585
R1303 gnd.n700 gnd.n699 585
R1304 gnd.n699 gnd.n698 585
R1305 gnd.n6488 gnd.n6487 585
R1306 gnd.n6489 gnd.n6488 585
R1307 gnd.n697 gnd.n696 585
R1308 gnd.n6490 gnd.n697 585
R1309 gnd.n6493 gnd.n6492 585
R1310 gnd.n6492 gnd.n6491 585
R1311 gnd.n694 gnd.n693 585
R1312 gnd.n693 gnd.n692 585
R1313 gnd.n6499 gnd.n6498 585
R1314 gnd.n6500 gnd.n6499 585
R1315 gnd.n691 gnd.n690 585
R1316 gnd.n6501 gnd.n691 585
R1317 gnd.n6504 gnd.n6503 585
R1318 gnd.n6503 gnd.n6502 585
R1319 gnd.n6505 gnd.n688 585
R1320 gnd.n688 gnd.n687 585
R1321 gnd.n563 gnd.n562 585
R1322 gnd.n6712 gnd.n562 585
R1323 gnd.n6715 gnd.n6714 585
R1324 gnd.n6714 gnd.n6713 585
R1325 gnd.n566 gnd.n565 585
R1326 gnd.n6711 gnd.n566 585
R1327 gnd.n6709 gnd.n6708 585
R1328 gnd.n6710 gnd.n6709 585
R1329 gnd.n569 gnd.n568 585
R1330 gnd.n568 gnd.n567 585
R1331 gnd.n6704 gnd.n6703 585
R1332 gnd.n6703 gnd.n6702 585
R1333 gnd.n572 gnd.n571 585
R1334 gnd.n6701 gnd.n572 585
R1335 gnd.n6699 gnd.n6698 585
R1336 gnd.n6700 gnd.n6699 585
R1337 gnd.n575 gnd.n574 585
R1338 gnd.n574 gnd.n573 585
R1339 gnd.n6694 gnd.n6693 585
R1340 gnd.n6693 gnd.n6692 585
R1341 gnd.n578 gnd.n577 585
R1342 gnd.n6691 gnd.n578 585
R1343 gnd.n6689 gnd.n6688 585
R1344 gnd.n6690 gnd.n6689 585
R1345 gnd.n581 gnd.n580 585
R1346 gnd.n580 gnd.n579 585
R1347 gnd.n6684 gnd.n6683 585
R1348 gnd.n6683 gnd.n6682 585
R1349 gnd.n584 gnd.n583 585
R1350 gnd.n6681 gnd.n584 585
R1351 gnd.n6679 gnd.n6678 585
R1352 gnd.n6680 gnd.n6679 585
R1353 gnd.n587 gnd.n586 585
R1354 gnd.n586 gnd.n585 585
R1355 gnd.n6674 gnd.n6673 585
R1356 gnd.n6673 gnd.n6672 585
R1357 gnd.n590 gnd.n589 585
R1358 gnd.n6671 gnd.n590 585
R1359 gnd.n6669 gnd.n6668 585
R1360 gnd.n6670 gnd.n6669 585
R1361 gnd.n593 gnd.n592 585
R1362 gnd.n592 gnd.n591 585
R1363 gnd.n6664 gnd.n6663 585
R1364 gnd.n6663 gnd.n6662 585
R1365 gnd.n596 gnd.n595 585
R1366 gnd.n6661 gnd.n596 585
R1367 gnd.n6659 gnd.n6658 585
R1368 gnd.n6660 gnd.n6659 585
R1369 gnd.n599 gnd.n598 585
R1370 gnd.n598 gnd.n597 585
R1371 gnd.n6654 gnd.n6653 585
R1372 gnd.n6653 gnd.n6652 585
R1373 gnd.n602 gnd.n601 585
R1374 gnd.n6651 gnd.n602 585
R1375 gnd.n6649 gnd.n6648 585
R1376 gnd.n6650 gnd.n6649 585
R1377 gnd.n605 gnd.n604 585
R1378 gnd.n604 gnd.n603 585
R1379 gnd.n6644 gnd.n6643 585
R1380 gnd.n6643 gnd.n6642 585
R1381 gnd.n608 gnd.n607 585
R1382 gnd.n6641 gnd.n608 585
R1383 gnd.n6639 gnd.n6638 585
R1384 gnd.n6640 gnd.n6639 585
R1385 gnd.n611 gnd.n610 585
R1386 gnd.n610 gnd.n609 585
R1387 gnd.n6634 gnd.n6633 585
R1388 gnd.n6633 gnd.n6632 585
R1389 gnd.n614 gnd.n613 585
R1390 gnd.n6631 gnd.n614 585
R1391 gnd.n6629 gnd.n6628 585
R1392 gnd.n6630 gnd.n6629 585
R1393 gnd.n617 gnd.n616 585
R1394 gnd.n616 gnd.n615 585
R1395 gnd.n6624 gnd.n6623 585
R1396 gnd.n6623 gnd.n6622 585
R1397 gnd.n620 gnd.n619 585
R1398 gnd.n6621 gnd.n620 585
R1399 gnd.n6619 gnd.n6618 585
R1400 gnd.n6620 gnd.n6619 585
R1401 gnd.n623 gnd.n622 585
R1402 gnd.n622 gnd.n621 585
R1403 gnd.n6614 gnd.n6613 585
R1404 gnd.n6613 gnd.n6612 585
R1405 gnd.n626 gnd.n625 585
R1406 gnd.n6611 gnd.n626 585
R1407 gnd.n6609 gnd.n6608 585
R1408 gnd.n6610 gnd.n6609 585
R1409 gnd.n629 gnd.n628 585
R1410 gnd.n628 gnd.n627 585
R1411 gnd.n6604 gnd.n6603 585
R1412 gnd.n6603 gnd.n6602 585
R1413 gnd.n632 gnd.n631 585
R1414 gnd.n6601 gnd.n632 585
R1415 gnd.n6599 gnd.n6598 585
R1416 gnd.n6600 gnd.n6599 585
R1417 gnd.n635 gnd.n634 585
R1418 gnd.n634 gnd.n633 585
R1419 gnd.n6594 gnd.n6593 585
R1420 gnd.n6593 gnd.n6592 585
R1421 gnd.n638 gnd.n637 585
R1422 gnd.n6591 gnd.n638 585
R1423 gnd.n6589 gnd.n6588 585
R1424 gnd.n6590 gnd.n6589 585
R1425 gnd.n641 gnd.n640 585
R1426 gnd.n640 gnd.n639 585
R1427 gnd.n6584 gnd.n6583 585
R1428 gnd.n6583 gnd.n6582 585
R1429 gnd.n644 gnd.n643 585
R1430 gnd.n6581 gnd.n644 585
R1431 gnd.n6579 gnd.n6578 585
R1432 gnd.n6580 gnd.n6579 585
R1433 gnd.n647 gnd.n646 585
R1434 gnd.n646 gnd.n645 585
R1435 gnd.n6574 gnd.n6573 585
R1436 gnd.n6573 gnd.n6572 585
R1437 gnd.n650 gnd.n649 585
R1438 gnd.n6571 gnd.n650 585
R1439 gnd.n6569 gnd.n6568 585
R1440 gnd.n6570 gnd.n6569 585
R1441 gnd.n653 gnd.n652 585
R1442 gnd.n652 gnd.n651 585
R1443 gnd.n6564 gnd.n6563 585
R1444 gnd.n6563 gnd.n6562 585
R1445 gnd.n656 gnd.n655 585
R1446 gnd.n6561 gnd.n656 585
R1447 gnd.n6559 gnd.n6558 585
R1448 gnd.n6560 gnd.n6559 585
R1449 gnd.n659 gnd.n658 585
R1450 gnd.n658 gnd.n657 585
R1451 gnd.n6554 gnd.n6553 585
R1452 gnd.n6553 gnd.n6552 585
R1453 gnd.n662 gnd.n661 585
R1454 gnd.n6551 gnd.n662 585
R1455 gnd.n6549 gnd.n6548 585
R1456 gnd.n6550 gnd.n6549 585
R1457 gnd.n665 gnd.n664 585
R1458 gnd.n664 gnd.n663 585
R1459 gnd.n6544 gnd.n6543 585
R1460 gnd.n6543 gnd.n6542 585
R1461 gnd.n668 gnd.n667 585
R1462 gnd.n6541 gnd.n668 585
R1463 gnd.n6539 gnd.n6538 585
R1464 gnd.n6540 gnd.n6539 585
R1465 gnd.n671 gnd.n670 585
R1466 gnd.n670 gnd.n669 585
R1467 gnd.n6534 gnd.n6533 585
R1468 gnd.n6533 gnd.n6532 585
R1469 gnd.n674 gnd.n673 585
R1470 gnd.n6531 gnd.n674 585
R1471 gnd.n6529 gnd.n6528 585
R1472 gnd.n6530 gnd.n6529 585
R1473 gnd.n677 gnd.n676 585
R1474 gnd.n676 gnd.n675 585
R1475 gnd.n6524 gnd.n6523 585
R1476 gnd.n6523 gnd.n6522 585
R1477 gnd.n680 gnd.n679 585
R1478 gnd.n6521 gnd.n680 585
R1479 gnd.n6519 gnd.n6518 585
R1480 gnd.n6520 gnd.n6519 585
R1481 gnd.n683 gnd.n682 585
R1482 gnd.n682 gnd.n681 585
R1483 gnd.n6514 gnd.n6513 585
R1484 gnd.n6513 gnd.n6512 585
R1485 gnd.n686 gnd.n685 585
R1486 gnd.n6511 gnd.n686 585
R1487 gnd.n6509 gnd.n6508 585
R1488 gnd.n6510 gnd.n6509 585
R1489 gnd.n1133 gnd.n1132 585
R1490 gnd.n4569 gnd.n1133 585
R1491 gnd.n5966 gnd.n5965 585
R1492 gnd.n5965 gnd.n5964 585
R1493 gnd.n5967 gnd.n1128 585
R1494 gnd.n4529 gnd.n1128 585
R1495 gnd.n5969 gnd.n5968 585
R1496 gnd.n5970 gnd.n5969 585
R1497 gnd.n1112 gnd.n1111 585
R1498 gnd.n4267 gnd.n1112 585
R1499 gnd.n5978 gnd.n5977 585
R1500 gnd.n5977 gnd.n5976 585
R1501 gnd.n5979 gnd.n1107 585
R1502 gnd.n4542 gnd.n1107 585
R1503 gnd.n5981 gnd.n5980 585
R1504 gnd.n5982 gnd.n5981 585
R1505 gnd.n1093 gnd.n1092 585
R1506 gnd.n4260 gnd.n1093 585
R1507 gnd.n5990 gnd.n5989 585
R1508 gnd.n5989 gnd.n5988 585
R1509 gnd.n5991 gnd.n1088 585
R1510 gnd.n4252 gnd.n1088 585
R1511 gnd.n5993 gnd.n5992 585
R1512 gnd.n5994 gnd.n5993 585
R1513 gnd.n1072 gnd.n1071 585
R1514 gnd.n4217 gnd.n1072 585
R1515 gnd.n6002 gnd.n6001 585
R1516 gnd.n6001 gnd.n6000 585
R1517 gnd.n6003 gnd.n1066 585
R1518 gnd.n4225 gnd.n1066 585
R1519 gnd.n6005 gnd.n6004 585
R1520 gnd.n6006 gnd.n6005 585
R1521 gnd.n1067 gnd.n1065 585
R1522 gnd.n4206 gnd.n1065 585
R1523 gnd.n4182 gnd.n1054 585
R1524 gnd.n6012 gnd.n1054 585
R1525 gnd.n4184 gnd.n4183 585
R1526 gnd.n4183 gnd.n1050 585
R1527 gnd.n4185 gnd.n2165 585
R1528 gnd.n4197 gnd.n2165 585
R1529 gnd.n4186 gnd.n2174 585
R1530 gnd.n2174 gnd.n2172 585
R1531 gnd.n4188 gnd.n4187 585
R1532 gnd.n4189 gnd.n4188 585
R1533 gnd.n2175 gnd.n2173 585
R1534 gnd.n2173 gnd.n2169 585
R1535 gnd.n4158 gnd.n2184 585
R1536 gnd.n4170 gnd.n2184 585
R1537 gnd.n4159 gnd.n2192 585
R1538 gnd.n2192 gnd.n2182 585
R1539 gnd.n4161 gnd.n4160 585
R1540 gnd.n4162 gnd.n4161 585
R1541 gnd.n2193 gnd.n2191 585
R1542 gnd.n2191 gnd.n2188 585
R1543 gnd.n4137 gnd.n2199 585
R1544 gnd.n4150 gnd.n2199 585
R1545 gnd.n4138 gnd.n2210 585
R1546 gnd.n2210 gnd.n2208 585
R1547 gnd.n4140 gnd.n4139 585
R1548 gnd.n4141 gnd.n4140 585
R1549 gnd.n2211 gnd.n2209 585
R1550 gnd.n2209 gnd.n2205 585
R1551 gnd.n4117 gnd.n2218 585
R1552 gnd.n4129 gnd.n2218 585
R1553 gnd.n4118 gnd.n2228 585
R1554 gnd.n2228 gnd.n2216 585
R1555 gnd.n4120 gnd.n4119 585
R1556 gnd.n4121 gnd.n4120 585
R1557 gnd.n2229 gnd.n2227 585
R1558 gnd.n2227 gnd.n2224 585
R1559 gnd.n4097 gnd.n2235 585
R1560 gnd.n4109 gnd.n2235 585
R1561 gnd.n4098 gnd.n2246 585
R1562 gnd.n2246 gnd.n2244 585
R1563 gnd.n4100 gnd.n4099 585
R1564 gnd.n4101 gnd.n4100 585
R1565 gnd.n2247 gnd.n2245 585
R1566 gnd.n2245 gnd.n2241 585
R1567 gnd.n2268 gnd.n2254 585
R1568 gnd.n4089 gnd.n2254 585
R1569 gnd.n2266 gnd.n2264 585
R1570 gnd.n2264 gnd.n2252 585
R1571 gnd.n4080 gnd.n4079 585
R1572 gnd.n4081 gnd.n4080 585
R1573 gnd.n2265 gnd.n2263 585
R1574 gnd.n2263 gnd.n2260 585
R1575 gnd.n3951 gnd.n3950 585
R1576 gnd.n3949 gnd.n3948 585
R1577 gnd.n3947 gnd.n3946 585
R1578 gnd.n3945 gnd.n3944 585
R1579 gnd.n3943 gnd.n3942 585
R1580 gnd.n3941 gnd.n3940 585
R1581 gnd.n3939 gnd.n3938 585
R1582 gnd.n3937 gnd.n3936 585
R1583 gnd.n3935 gnd.n3934 585
R1584 gnd.n3933 gnd.n3932 585
R1585 gnd.n3931 gnd.n3930 585
R1586 gnd.n3929 gnd.n3928 585
R1587 gnd.n3927 gnd.n3926 585
R1588 gnd.n3925 gnd.n3924 585
R1589 gnd.n3923 gnd.n3922 585
R1590 gnd.n3921 gnd.n3920 585
R1591 gnd.n3919 gnd.n3918 585
R1592 gnd.n3856 gnd.n3853 585
R1593 gnd.n3914 gnd.n3772 585
R1594 gnd.n4071 gnd.n3772 585
R1595 gnd.n4572 gnd.n4571 585
R1596 gnd.n4366 gnd.n2124 585
R1597 gnd.n4378 gnd.n4367 585
R1598 gnd.n4379 gnd.n4365 585
R1599 gnd.n4364 gnd.n4356 585
R1600 gnd.n4386 gnd.n4355 585
R1601 gnd.n4387 gnd.n4354 585
R1602 gnd.n4348 gnd.n4347 585
R1603 gnd.n4394 gnd.n4346 585
R1604 gnd.n4395 gnd.n4345 585
R1605 gnd.n4344 gnd.n4336 585
R1606 gnd.n4402 gnd.n4335 585
R1607 gnd.n4403 gnd.n4334 585
R1608 gnd.n4328 gnd.n4327 585
R1609 gnd.n4410 gnd.n4326 585
R1610 gnd.n4411 gnd.n4325 585
R1611 gnd.n4324 gnd.n4316 585
R1612 gnd.n4418 gnd.n4315 585
R1613 gnd.n4419 gnd.n1145 585
R1614 gnd.n5956 gnd.n1145 585
R1615 gnd.n4570 gnd.n2125 585
R1616 gnd.n4570 gnd.n4569 585
R1617 gnd.n4531 gnd.n1136 585
R1618 gnd.n5964 gnd.n1136 585
R1619 gnd.n4534 gnd.n4530 585
R1620 gnd.n4530 gnd.n4529 585
R1621 gnd.n4535 gnd.n1126 585
R1622 gnd.n5970 gnd.n1126 585
R1623 gnd.n4536 gnd.n2142 585
R1624 gnd.n4267 gnd.n2142 585
R1625 gnd.n2139 gnd.n1115 585
R1626 gnd.n5976 gnd.n1115 585
R1627 gnd.n4541 gnd.n4540 585
R1628 gnd.n4542 gnd.n4541 585
R1629 gnd.n2138 gnd.n1106 585
R1630 gnd.n5982 gnd.n1106 585
R1631 gnd.n4259 gnd.n4258 585
R1632 gnd.n4260 gnd.n4259 585
R1633 gnd.n2145 gnd.n1095 585
R1634 gnd.n5988 gnd.n1095 585
R1635 gnd.n4254 gnd.n4253 585
R1636 gnd.n4253 gnd.n4252 585
R1637 gnd.n2147 gnd.n1086 585
R1638 gnd.n5994 gnd.n1086 585
R1639 gnd.n4219 gnd.n4218 585
R1640 gnd.n4218 gnd.n4217 585
R1641 gnd.n2156 gnd.n1075 585
R1642 gnd.n6000 gnd.n1075 585
R1643 gnd.n4224 gnd.n4223 585
R1644 gnd.n4225 gnd.n4224 585
R1645 gnd.n2155 gnd.n1064 585
R1646 gnd.n6006 gnd.n1064 585
R1647 gnd.n4205 gnd.n4204 585
R1648 gnd.n4206 gnd.n4205 585
R1649 gnd.n2160 gnd.n1052 585
R1650 gnd.n6012 gnd.n1052 585
R1651 gnd.n4200 gnd.n4199 585
R1652 gnd.n4199 gnd.n1050 585
R1653 gnd.n4198 gnd.n2162 585
R1654 gnd.n4198 gnd.n4197 585
R1655 gnd.n3877 gnd.n2163 585
R1656 gnd.n2172 gnd.n2163 585
R1657 gnd.n3880 gnd.n2171 585
R1658 gnd.n4189 gnd.n2171 585
R1659 gnd.n3882 gnd.n3881 585
R1660 gnd.n3881 gnd.n2169 585
R1661 gnd.n3883 gnd.n2183 585
R1662 gnd.n4170 gnd.n2183 585
R1663 gnd.n3885 gnd.n3884 585
R1664 gnd.n3884 gnd.n2182 585
R1665 gnd.n3886 gnd.n2190 585
R1666 gnd.n4162 gnd.n2190 585
R1667 gnd.n3888 gnd.n3887 585
R1668 gnd.n3887 gnd.n2188 585
R1669 gnd.n3889 gnd.n2198 585
R1670 gnd.n4150 gnd.n2198 585
R1671 gnd.n3891 gnd.n3890 585
R1672 gnd.n3890 gnd.n2208 585
R1673 gnd.n3892 gnd.n2207 585
R1674 gnd.n4141 gnd.n2207 585
R1675 gnd.n3894 gnd.n3893 585
R1676 gnd.n3893 gnd.n2205 585
R1677 gnd.n3895 gnd.n2217 585
R1678 gnd.n4129 gnd.n2217 585
R1679 gnd.n3897 gnd.n3896 585
R1680 gnd.n3896 gnd.n2216 585
R1681 gnd.n3898 gnd.n2226 585
R1682 gnd.n4121 gnd.n2226 585
R1683 gnd.n3900 gnd.n3899 585
R1684 gnd.n3899 gnd.n2224 585
R1685 gnd.n3901 gnd.n2234 585
R1686 gnd.n4109 gnd.n2234 585
R1687 gnd.n3903 gnd.n3902 585
R1688 gnd.n3902 gnd.n2244 585
R1689 gnd.n3904 gnd.n2243 585
R1690 gnd.n4101 gnd.n2243 585
R1691 gnd.n3906 gnd.n3905 585
R1692 gnd.n3905 gnd.n2241 585
R1693 gnd.n3907 gnd.n2253 585
R1694 gnd.n4089 gnd.n2253 585
R1695 gnd.n3909 gnd.n3908 585
R1696 gnd.n3908 gnd.n2252 585
R1697 gnd.n3910 gnd.n2262 585
R1698 gnd.n4081 gnd.n2262 585
R1699 gnd.n3912 gnd.n3911 585
R1700 gnd.n3911 gnd.n2260 585
R1701 gnd.n3643 gnd.n3642 585
R1702 gnd.n3644 gnd.n3643 585
R1703 gnd.n2349 gnd.n2348 585
R1704 gnd.n2355 gnd.n2348 585
R1705 gnd.n3618 gnd.n2367 585
R1706 gnd.n2367 gnd.n2354 585
R1707 gnd.n3620 gnd.n3619 585
R1708 gnd.n3621 gnd.n3620 585
R1709 gnd.n2368 gnd.n2366 585
R1710 gnd.n2366 gnd.n2362 585
R1711 gnd.n3352 gnd.n3351 585
R1712 gnd.n3351 gnd.n3350 585
R1713 gnd.n2373 gnd.n2372 585
R1714 gnd.n3320 gnd.n2373 585
R1715 gnd.n3340 gnd.n3339 585
R1716 gnd.n3339 gnd.n3338 585
R1717 gnd.n2380 gnd.n2379 585
R1718 gnd.n3326 gnd.n2380 585
R1719 gnd.n3296 gnd.n2400 585
R1720 gnd.n2400 gnd.n2399 585
R1721 gnd.n3298 gnd.n3297 585
R1722 gnd.n3299 gnd.n3298 585
R1723 gnd.n2401 gnd.n2398 585
R1724 gnd.n2409 gnd.n2398 585
R1725 gnd.n3274 gnd.n2421 585
R1726 gnd.n2421 gnd.n2408 585
R1727 gnd.n3276 gnd.n3275 585
R1728 gnd.n3277 gnd.n3276 585
R1729 gnd.n2422 gnd.n2420 585
R1730 gnd.n2420 gnd.n2416 585
R1731 gnd.n3262 gnd.n3261 585
R1732 gnd.n3261 gnd.n3260 585
R1733 gnd.n2427 gnd.n2426 585
R1734 gnd.n2437 gnd.n2427 585
R1735 gnd.n3251 gnd.n3250 585
R1736 gnd.n3250 gnd.n3249 585
R1737 gnd.n2434 gnd.n2433 585
R1738 gnd.n3237 gnd.n2434 585
R1739 gnd.n3211 gnd.n2455 585
R1740 gnd.n2455 gnd.n2444 585
R1741 gnd.n3213 gnd.n3212 585
R1742 gnd.n3214 gnd.n3213 585
R1743 gnd.n2456 gnd.n2454 585
R1744 gnd.n2464 gnd.n2454 585
R1745 gnd.n3189 gnd.n2476 585
R1746 gnd.n2476 gnd.n2463 585
R1747 gnd.n3191 gnd.n3190 585
R1748 gnd.n3192 gnd.n3191 585
R1749 gnd.n2477 gnd.n2475 585
R1750 gnd.n2475 gnd.n2471 585
R1751 gnd.n3177 gnd.n3176 585
R1752 gnd.n3176 gnd.n3175 585
R1753 gnd.n2482 gnd.n2481 585
R1754 gnd.n2491 gnd.n2482 585
R1755 gnd.n3166 gnd.n3165 585
R1756 gnd.n3165 gnd.n3164 585
R1757 gnd.n2489 gnd.n2488 585
R1758 gnd.n3152 gnd.n2489 585
R1759 gnd.n2590 gnd.n2589 585
R1760 gnd.n2590 gnd.n2498 585
R1761 gnd.n3109 gnd.n3108 585
R1762 gnd.n3108 gnd.n3107 585
R1763 gnd.n3110 gnd.n2584 585
R1764 gnd.n2595 gnd.n2584 585
R1765 gnd.n3112 gnd.n3111 585
R1766 gnd.n3113 gnd.n3112 585
R1767 gnd.n2585 gnd.n2583 585
R1768 gnd.n2608 gnd.n2583 585
R1769 gnd.n2568 gnd.n2567 585
R1770 gnd.n2571 gnd.n2568 585
R1771 gnd.n3123 gnd.n3122 585
R1772 gnd.n3122 gnd.n3121 585
R1773 gnd.n3124 gnd.n2562 585
R1774 gnd.n3083 gnd.n2562 585
R1775 gnd.n3126 gnd.n3125 585
R1776 gnd.n3127 gnd.n3126 585
R1777 gnd.n2563 gnd.n2561 585
R1778 gnd.n2622 gnd.n2561 585
R1779 gnd.n3075 gnd.n3074 585
R1780 gnd.n3074 gnd.n3073 585
R1781 gnd.n2619 gnd.n2618 585
R1782 gnd.n3057 gnd.n2619 585
R1783 gnd.n3044 gnd.n2638 585
R1784 gnd.n2638 gnd.n2637 585
R1785 gnd.n3046 gnd.n3045 585
R1786 gnd.n3047 gnd.n3046 585
R1787 gnd.n2639 gnd.n2636 585
R1788 gnd.n2645 gnd.n2636 585
R1789 gnd.n3025 gnd.n3024 585
R1790 gnd.n3026 gnd.n3025 585
R1791 gnd.n2656 gnd.n2655 585
R1792 gnd.n2655 gnd.n2651 585
R1793 gnd.n3015 gnd.n3014 585
R1794 gnd.n3016 gnd.n3015 585
R1795 gnd.n2666 gnd.n2665 585
R1796 gnd.n2671 gnd.n2665 585
R1797 gnd.n2993 gnd.n2684 585
R1798 gnd.n2684 gnd.n2670 585
R1799 gnd.n2995 gnd.n2994 585
R1800 gnd.n2996 gnd.n2995 585
R1801 gnd.n2685 gnd.n2683 585
R1802 gnd.n2683 gnd.n2679 585
R1803 gnd.n2984 gnd.n2983 585
R1804 gnd.n2985 gnd.n2984 585
R1805 gnd.n2692 gnd.n2691 585
R1806 gnd.n2696 gnd.n2691 585
R1807 gnd.n2961 gnd.n2713 585
R1808 gnd.n2713 gnd.n2695 585
R1809 gnd.n2963 gnd.n2962 585
R1810 gnd.n2964 gnd.n2963 585
R1811 gnd.n2714 gnd.n2712 585
R1812 gnd.n2712 gnd.n2703 585
R1813 gnd.n2956 gnd.n2955 585
R1814 gnd.n2955 gnd.n2954 585
R1815 gnd.n2761 gnd.n2760 585
R1816 gnd.n2762 gnd.n2761 585
R1817 gnd.n2915 gnd.n2914 585
R1818 gnd.n2916 gnd.n2915 585
R1819 gnd.n2771 gnd.n2770 585
R1820 gnd.n2770 gnd.n2769 585
R1821 gnd.n2910 gnd.n2909 585
R1822 gnd.n2909 gnd.n2908 585
R1823 gnd.n2774 gnd.n2773 585
R1824 gnd.n2775 gnd.n2774 585
R1825 gnd.n2899 gnd.n2898 585
R1826 gnd.n2900 gnd.n2899 585
R1827 gnd.n2782 gnd.n2781 585
R1828 gnd.n2891 gnd.n2781 585
R1829 gnd.n2894 gnd.n2893 585
R1830 gnd.n2893 gnd.n2892 585
R1831 gnd.n2785 gnd.n2784 585
R1832 gnd.n2786 gnd.n2785 585
R1833 gnd.n2880 gnd.n2879 585
R1834 gnd.n2878 gnd.n2804 585
R1835 gnd.n2877 gnd.n2803 585
R1836 gnd.n2882 gnd.n2803 585
R1837 gnd.n2876 gnd.n2875 585
R1838 gnd.n2874 gnd.n2873 585
R1839 gnd.n2872 gnd.n2871 585
R1840 gnd.n2870 gnd.n2869 585
R1841 gnd.n2868 gnd.n2867 585
R1842 gnd.n2866 gnd.n2865 585
R1843 gnd.n2864 gnd.n2863 585
R1844 gnd.n2862 gnd.n2861 585
R1845 gnd.n2860 gnd.n2859 585
R1846 gnd.n2858 gnd.n2857 585
R1847 gnd.n2856 gnd.n2855 585
R1848 gnd.n2854 gnd.n2853 585
R1849 gnd.n2852 gnd.n2851 585
R1850 gnd.n2850 gnd.n2849 585
R1851 gnd.n2848 gnd.n2847 585
R1852 gnd.n2846 gnd.n2845 585
R1853 gnd.n2844 gnd.n2843 585
R1854 gnd.n2842 gnd.n2841 585
R1855 gnd.n2840 gnd.n2839 585
R1856 gnd.n2838 gnd.n2837 585
R1857 gnd.n2836 gnd.n2835 585
R1858 gnd.n2834 gnd.n2833 585
R1859 gnd.n2791 gnd.n2790 585
R1860 gnd.n2885 gnd.n2884 585
R1861 gnd.n3647 gnd.n3646 585
R1862 gnd.n3649 gnd.n3648 585
R1863 gnd.n3651 gnd.n3650 585
R1864 gnd.n3653 gnd.n3652 585
R1865 gnd.n3655 gnd.n3654 585
R1866 gnd.n3657 gnd.n3656 585
R1867 gnd.n3659 gnd.n3658 585
R1868 gnd.n3661 gnd.n3660 585
R1869 gnd.n3663 gnd.n3662 585
R1870 gnd.n3665 gnd.n3664 585
R1871 gnd.n3667 gnd.n3666 585
R1872 gnd.n3669 gnd.n3668 585
R1873 gnd.n3671 gnd.n3670 585
R1874 gnd.n3673 gnd.n3672 585
R1875 gnd.n3675 gnd.n3674 585
R1876 gnd.n3677 gnd.n3676 585
R1877 gnd.n3679 gnd.n3678 585
R1878 gnd.n3681 gnd.n3680 585
R1879 gnd.n3683 gnd.n3682 585
R1880 gnd.n3685 gnd.n3684 585
R1881 gnd.n3687 gnd.n3686 585
R1882 gnd.n3689 gnd.n3688 585
R1883 gnd.n3691 gnd.n3690 585
R1884 gnd.n3693 gnd.n3692 585
R1885 gnd.n3695 gnd.n3694 585
R1886 gnd.n3696 gnd.n2316 585
R1887 gnd.n3697 gnd.n2274 585
R1888 gnd.n3735 gnd.n2274 585
R1889 gnd.n3645 gnd.n2346 585
R1890 gnd.n3645 gnd.n3644 585
R1891 gnd.n3313 gnd.n2345 585
R1892 gnd.n2355 gnd.n2345 585
R1893 gnd.n3315 gnd.n3314 585
R1894 gnd.n3314 gnd.n2354 585
R1895 gnd.n3316 gnd.n2364 585
R1896 gnd.n3621 gnd.n2364 585
R1897 gnd.n3318 gnd.n3317 585
R1898 gnd.n3317 gnd.n2362 585
R1899 gnd.n3319 gnd.n2375 585
R1900 gnd.n3350 gnd.n2375 585
R1901 gnd.n3322 gnd.n3321 585
R1902 gnd.n3321 gnd.n3320 585
R1903 gnd.n3323 gnd.n2382 585
R1904 gnd.n3338 gnd.n2382 585
R1905 gnd.n3325 gnd.n3324 585
R1906 gnd.n3326 gnd.n3325 585
R1907 gnd.n2392 gnd.n2391 585
R1908 gnd.n2399 gnd.n2391 585
R1909 gnd.n3301 gnd.n3300 585
R1910 gnd.n3300 gnd.n3299 585
R1911 gnd.n2395 gnd.n2394 585
R1912 gnd.n2409 gnd.n2395 585
R1913 gnd.n3227 gnd.n3226 585
R1914 gnd.n3226 gnd.n2408 585
R1915 gnd.n3228 gnd.n2418 585
R1916 gnd.n3277 gnd.n2418 585
R1917 gnd.n3230 gnd.n3229 585
R1918 gnd.n3229 gnd.n2416 585
R1919 gnd.n3231 gnd.n2429 585
R1920 gnd.n3260 gnd.n2429 585
R1921 gnd.n3233 gnd.n3232 585
R1922 gnd.n3232 gnd.n2437 585
R1923 gnd.n3234 gnd.n2436 585
R1924 gnd.n3249 gnd.n2436 585
R1925 gnd.n3236 gnd.n3235 585
R1926 gnd.n3237 gnd.n3236 585
R1927 gnd.n2448 gnd.n2447 585
R1928 gnd.n2447 gnd.n2444 585
R1929 gnd.n3216 gnd.n3215 585
R1930 gnd.n3215 gnd.n3214 585
R1931 gnd.n2451 gnd.n2450 585
R1932 gnd.n2464 gnd.n2451 585
R1933 gnd.n3140 gnd.n3139 585
R1934 gnd.n3139 gnd.n2463 585
R1935 gnd.n3141 gnd.n2473 585
R1936 gnd.n3192 gnd.n2473 585
R1937 gnd.n3143 gnd.n3142 585
R1938 gnd.n3142 gnd.n2471 585
R1939 gnd.n3144 gnd.n2484 585
R1940 gnd.n3175 gnd.n2484 585
R1941 gnd.n3146 gnd.n3145 585
R1942 gnd.n3145 gnd.n2491 585
R1943 gnd.n3147 gnd.n2490 585
R1944 gnd.n3164 gnd.n2490 585
R1945 gnd.n3149 gnd.n3148 585
R1946 gnd.n3152 gnd.n3149 585
R1947 gnd.n2501 gnd.n2500 585
R1948 gnd.n2500 gnd.n2498 585
R1949 gnd.n2592 gnd.n2591 585
R1950 gnd.n3107 gnd.n2591 585
R1951 gnd.n2594 gnd.n2593 585
R1952 gnd.n2595 gnd.n2594 585
R1953 gnd.n2605 gnd.n2581 585
R1954 gnd.n3113 gnd.n2581 585
R1955 gnd.n2607 gnd.n2606 585
R1956 gnd.n2608 gnd.n2607 585
R1957 gnd.n2604 gnd.n2603 585
R1958 gnd.n2604 gnd.n2571 585
R1959 gnd.n2602 gnd.n2569 585
R1960 gnd.n3121 gnd.n2569 585
R1961 gnd.n2558 gnd.n2556 585
R1962 gnd.n3083 gnd.n2558 585
R1963 gnd.n3129 gnd.n3128 585
R1964 gnd.n3128 gnd.n3127 585
R1965 gnd.n2557 gnd.n2555 585
R1966 gnd.n2622 gnd.n2557 585
R1967 gnd.n3054 gnd.n2621 585
R1968 gnd.n3073 gnd.n2621 585
R1969 gnd.n3056 gnd.n3055 585
R1970 gnd.n3057 gnd.n3056 585
R1971 gnd.n2631 gnd.n2630 585
R1972 gnd.n2637 gnd.n2630 585
R1973 gnd.n3049 gnd.n3048 585
R1974 gnd.n3048 gnd.n3047 585
R1975 gnd.n2634 gnd.n2633 585
R1976 gnd.n2645 gnd.n2634 585
R1977 gnd.n2934 gnd.n2653 585
R1978 gnd.n3026 gnd.n2653 585
R1979 gnd.n2936 gnd.n2935 585
R1980 gnd.n2935 gnd.n2651 585
R1981 gnd.n2937 gnd.n2664 585
R1982 gnd.n3016 gnd.n2664 585
R1983 gnd.n2939 gnd.n2938 585
R1984 gnd.n2939 gnd.n2671 585
R1985 gnd.n2941 gnd.n2940 585
R1986 gnd.n2940 gnd.n2670 585
R1987 gnd.n2942 gnd.n2681 585
R1988 gnd.n2996 gnd.n2681 585
R1989 gnd.n2944 gnd.n2943 585
R1990 gnd.n2943 gnd.n2679 585
R1991 gnd.n2945 gnd.n2690 585
R1992 gnd.n2985 gnd.n2690 585
R1993 gnd.n2947 gnd.n2946 585
R1994 gnd.n2947 gnd.n2696 585
R1995 gnd.n2949 gnd.n2948 585
R1996 gnd.n2948 gnd.n2695 585
R1997 gnd.n2950 gnd.n2711 585
R1998 gnd.n2964 gnd.n2711 585
R1999 gnd.n2951 gnd.n2764 585
R2000 gnd.n2764 gnd.n2703 585
R2001 gnd.n2953 gnd.n2952 585
R2002 gnd.n2954 gnd.n2953 585
R2003 gnd.n2765 gnd.n2763 585
R2004 gnd.n2763 gnd.n2762 585
R2005 gnd.n2918 gnd.n2917 585
R2006 gnd.n2917 gnd.n2916 585
R2007 gnd.n2768 gnd.n2767 585
R2008 gnd.n2769 gnd.n2768 585
R2009 gnd.n2907 gnd.n2906 585
R2010 gnd.n2908 gnd.n2907 585
R2011 gnd.n2777 gnd.n2776 585
R2012 gnd.n2776 gnd.n2775 585
R2013 gnd.n2902 gnd.n2901 585
R2014 gnd.n2901 gnd.n2900 585
R2015 gnd.n2780 gnd.n2779 585
R2016 gnd.n2891 gnd.n2780 585
R2017 gnd.n2890 gnd.n2889 585
R2018 gnd.n2892 gnd.n2890 585
R2019 gnd.n2788 gnd.n2787 585
R2020 gnd.n2787 gnd.n2786 585
R2021 gnd.n6840 gnd.n6839 585
R2022 gnd.n6841 gnd.n6840 585
R2023 gnd.n153 gnd.n152 585
R2024 gnd.n162 gnd.n153 585
R2025 gnd.n6849 gnd.n6848 585
R2026 gnd.n6848 gnd.n6847 585
R2027 gnd.n6850 gnd.n148 585
R2028 gnd.n148 gnd.n147 585
R2029 gnd.n6852 gnd.n6851 585
R2030 gnd.n6853 gnd.n6852 585
R2031 gnd.n133 gnd.n132 585
R2032 gnd.n144 gnd.n133 585
R2033 gnd.n6861 gnd.n6860 585
R2034 gnd.n6860 gnd.n6859 585
R2035 gnd.n6862 gnd.n128 585
R2036 gnd.n128 gnd.n127 585
R2037 gnd.n6864 gnd.n6863 585
R2038 gnd.n6865 gnd.n6864 585
R2039 gnd.n113 gnd.n112 585
R2040 gnd.n124 gnd.n113 585
R2041 gnd.n6873 gnd.n6872 585
R2042 gnd.n6872 gnd.n6871 585
R2043 gnd.n6874 gnd.n108 585
R2044 gnd.n114 gnd.n108 585
R2045 gnd.n6876 gnd.n6875 585
R2046 gnd.n6877 gnd.n6876 585
R2047 gnd.n96 gnd.n95 585
R2048 gnd.n99 gnd.n96 585
R2049 gnd.n6885 gnd.n6884 585
R2050 gnd.n6884 gnd.n6883 585
R2051 gnd.n6886 gnd.n90 585
R2052 gnd.n90 gnd.n88 585
R2053 gnd.n6888 gnd.n6887 585
R2054 gnd.n6889 gnd.n6888 585
R2055 gnd.n91 gnd.n89 585
R2056 gnd.n89 gnd.n85 585
R2057 gnd.n6804 gnd.n6803 585
R2058 gnd.n6803 gnd.n70 585
R2059 gnd.n6802 gnd.n71 585
R2060 gnd.n6897 gnd.n71 585
R2061 gnd.n6801 gnd.n6800 585
R2062 gnd.n6800 gnd.n6799 585
R2063 gnd.n498 gnd.n496 585
R2064 gnd.n499 gnd.n498 585
R2065 gnd.n6792 gnd.n6791 585
R2066 gnd.n6791 gnd.n6790 585
R2067 gnd.n504 gnd.n503 585
R2068 gnd.n6782 gnd.n504 585
R2069 gnd.n6765 gnd.n6764 585
R2070 gnd.n6764 gnd.n509 585
R2071 gnd.n6766 gnd.n519 585
R2072 gnd.n6774 gnd.n519 585
R2073 gnd.n6768 gnd.n6767 585
R2074 gnd.n6769 gnd.n6768 585
R2075 gnd.n525 gnd.n524 585
R2076 gnd.n6755 gnd.n524 585
R2077 gnd.n6731 gnd.n6730 585
R2078 gnd.n6730 gnd.n6729 585
R2079 gnd.n6732 gnd.n539 585
R2080 gnd.n6747 gnd.n539 585
R2081 gnd.n6733 gnd.n551 585
R2082 gnd.n1615 gnd.n551 585
R2083 gnd.n6735 gnd.n6734 585
R2084 gnd.n6736 gnd.n6735 585
R2085 gnd.n552 gnd.n550 585
R2086 gnd.n1622 gnd.n550 585
R2087 gnd.n5503 gnd.n1610 585
R2088 gnd.n5499 gnd.n1610 585
R2089 gnd.n5505 gnd.n5504 585
R2090 gnd.n5506 gnd.n5505 585
R2091 gnd.n1593 gnd.n1592 585
R2092 gnd.n5448 gnd.n1593 585
R2093 gnd.n5514 gnd.n5513 585
R2094 gnd.n5513 gnd.n5512 585
R2095 gnd.n5515 gnd.n1586 585
R2096 gnd.n5441 gnd.n1586 585
R2097 gnd.n5517 gnd.n5516 585
R2098 gnd.n5518 gnd.n5517 585
R2099 gnd.n1587 gnd.n1585 585
R2100 gnd.n5435 gnd.n1585 585
R2101 gnd.n1569 gnd.n1563 585
R2102 gnd.n5524 gnd.n1569 585
R2103 gnd.n5529 gnd.n1561 585
R2104 gnd.n5470 gnd.n1561 585
R2105 gnd.n5531 gnd.n5530 585
R2106 gnd.n5532 gnd.n5531 585
R2107 gnd.n1560 gnd.n1400 585
R2108 gnd.n5699 gnd.n1401 585
R2109 gnd.n5698 gnd.n1402 585
R2110 gnd.n1477 gnd.n1403 585
R2111 gnd.n5691 gnd.n1409 585
R2112 gnd.n5690 gnd.n1410 585
R2113 gnd.n1480 gnd.n1411 585
R2114 gnd.n5683 gnd.n1417 585
R2115 gnd.n5682 gnd.n1418 585
R2116 gnd.n1482 gnd.n1419 585
R2117 gnd.n5675 gnd.n1425 585
R2118 gnd.n5674 gnd.n1426 585
R2119 gnd.n1485 gnd.n1427 585
R2120 gnd.n5667 gnd.n1433 585
R2121 gnd.n5666 gnd.n1434 585
R2122 gnd.n1487 gnd.n1435 585
R2123 gnd.n5659 gnd.n1443 585
R2124 gnd.n5658 gnd.n5655 585
R2125 gnd.n1446 gnd.n1444 585
R2126 gnd.n5653 gnd.n1446 585
R2127 gnd.n199 gnd.n198 585
R2128 gnd.n250 gnd.n194 585
R2129 gnd.n252 gnd.n251 585
R2130 gnd.n254 gnd.n192 585
R2131 gnd.n256 gnd.n255 585
R2132 gnd.n257 gnd.n187 585
R2133 gnd.n259 gnd.n258 585
R2134 gnd.n261 gnd.n185 585
R2135 gnd.n263 gnd.n262 585
R2136 gnd.n264 gnd.n180 585
R2137 gnd.n266 gnd.n265 585
R2138 gnd.n268 gnd.n178 585
R2139 gnd.n270 gnd.n269 585
R2140 gnd.n271 gnd.n173 585
R2141 gnd.n273 gnd.n272 585
R2142 gnd.n275 gnd.n171 585
R2143 gnd.n277 gnd.n276 585
R2144 gnd.n278 gnd.n169 585
R2145 gnd.n279 gnd.n166 585
R2146 gnd.n166 gnd.n165 585
R2147 gnd.n246 gnd.n164 585
R2148 gnd.n6841 gnd.n164 585
R2149 gnd.n245 gnd.n244 585
R2150 gnd.n244 gnd.n162 585
R2151 gnd.n243 gnd.n155 585
R2152 gnd.n6847 gnd.n155 585
R2153 gnd.n204 gnd.n203 585
R2154 gnd.n203 gnd.n147 585
R2155 gnd.n239 gnd.n146 585
R2156 gnd.n6853 gnd.n146 585
R2157 gnd.n238 gnd.n237 585
R2158 gnd.n237 gnd.n144 585
R2159 gnd.n236 gnd.n135 585
R2160 gnd.n6859 gnd.n135 585
R2161 gnd.n207 gnd.n206 585
R2162 gnd.n206 gnd.n127 585
R2163 gnd.n232 gnd.n126 585
R2164 gnd.n6865 gnd.n126 585
R2165 gnd.n231 gnd.n230 585
R2166 gnd.n230 gnd.n124 585
R2167 gnd.n229 gnd.n116 585
R2168 gnd.n6871 gnd.n116 585
R2169 gnd.n210 gnd.n209 585
R2170 gnd.n209 gnd.n114 585
R2171 gnd.n225 gnd.n107 585
R2172 gnd.n6877 gnd.n107 585
R2173 gnd.n224 gnd.n223 585
R2174 gnd.n223 gnd.n99 585
R2175 gnd.n222 gnd.n98 585
R2176 gnd.n6883 gnd.n98 585
R2177 gnd.n213 gnd.n212 585
R2178 gnd.n212 gnd.n88 585
R2179 gnd.n218 gnd.n87 585
R2180 gnd.n6889 gnd.n87 585
R2181 gnd.n217 gnd.n216 585
R2182 gnd.n216 gnd.n85 585
R2183 gnd.n68 gnd.n67 585
R2184 gnd.n70 gnd.n68 585
R2185 gnd.n6899 gnd.n6898 585
R2186 gnd.n6898 gnd.n6897 585
R2187 gnd.n6900 gnd.n66 585
R2188 gnd.n6799 gnd.n66 585
R2189 gnd.n506 gnd.n64 585
R2190 gnd.n506 gnd.n499 585
R2191 gnd.n513 gnd.n507 585
R2192 gnd.n6790 gnd.n507 585
R2193 gnd.n6781 gnd.n6780 585
R2194 gnd.n6782 gnd.n6781 585
R2195 gnd.n512 gnd.n511 585
R2196 gnd.n511 gnd.n509 585
R2197 gnd.n6776 gnd.n6775 585
R2198 gnd.n6775 gnd.n6774 585
R2199 gnd.n516 gnd.n515 585
R2200 gnd.n6769 gnd.n516 585
R2201 gnd.n6754 gnd.n6753 585
R2202 gnd.n6755 gnd.n6754 585
R2203 gnd.n532 gnd.n531 585
R2204 gnd.n6729 gnd.n531 585
R2205 gnd.n6749 gnd.n6748 585
R2206 gnd.n6748 gnd.n6747 585
R2207 gnd.n535 gnd.n534 585
R2208 gnd.n1615 gnd.n535 585
R2209 gnd.n5452 gnd.n548 585
R2210 gnd.n6736 gnd.n548 585
R2211 gnd.n5451 gnd.n5450 585
R2212 gnd.n5450 gnd.n1622 585
R2213 gnd.n5456 gnd.n1621 585
R2214 gnd.n5499 gnd.n1621 585
R2215 gnd.n5457 gnd.n1608 585
R2216 gnd.n5506 gnd.n1608 585
R2217 gnd.n5458 gnd.n5449 585
R2218 gnd.n5449 gnd.n5448 585
R2219 gnd.n5438 gnd.n1596 585
R2220 gnd.n5512 gnd.n1596 585
R2221 gnd.n5462 gnd.n5437 585
R2222 gnd.n5441 gnd.n5437 585
R2223 gnd.n5463 gnd.n1583 585
R2224 gnd.n5518 gnd.n1583 585
R2225 gnd.n5464 gnd.n5436 585
R2226 gnd.n5436 gnd.n5435 585
R2227 gnd.n1635 gnd.n1567 585
R2228 gnd.n5524 gnd.n1567 585
R2229 gnd.n5469 gnd.n5468 585
R2230 gnd.n5470 gnd.n5469 585
R2231 gnd.n1634 gnd.n1558 585
R2232 gnd.n5532 gnd.n1558 585
R2233 gnd.n3630 gnd.n2296 585
R2234 gnd.n2296 gnd.n2273 585
R2235 gnd.n3631 gnd.n2357 585
R2236 gnd.n2357 gnd.n2347 585
R2237 gnd.n3633 gnd.n3632 585
R2238 gnd.n3634 gnd.n3633 585
R2239 gnd.n2358 gnd.n2356 585
R2240 gnd.n2365 gnd.n2356 585
R2241 gnd.n3624 gnd.n3623 585
R2242 gnd.n3623 gnd.n3622 585
R2243 gnd.n2361 gnd.n2360 585
R2244 gnd.n3349 gnd.n2361 585
R2245 gnd.n3334 gnd.n2384 585
R2246 gnd.n2384 gnd.n2374 585
R2247 gnd.n3336 gnd.n3335 585
R2248 gnd.n3337 gnd.n3336 585
R2249 gnd.n2385 gnd.n2383 585
R2250 gnd.n2383 gnd.n2381 585
R2251 gnd.n3329 gnd.n3328 585
R2252 gnd.n3328 gnd.n3327 585
R2253 gnd.n2388 gnd.n2387 585
R2254 gnd.n2397 gnd.n2388 585
R2255 gnd.n3285 gnd.n2411 585
R2256 gnd.n2411 gnd.n2396 585
R2257 gnd.n3287 gnd.n3286 585
R2258 gnd.n3288 gnd.n3287 585
R2259 gnd.n2412 gnd.n2410 585
R2260 gnd.n2419 gnd.n2410 585
R2261 gnd.n3280 gnd.n3279 585
R2262 gnd.n3279 gnd.n3278 585
R2263 gnd.n2415 gnd.n2414 585
R2264 gnd.n3259 gnd.n2415 585
R2265 gnd.n3245 gnd.n2439 585
R2266 gnd.n2439 gnd.n2428 585
R2267 gnd.n3247 gnd.n3246 585
R2268 gnd.n3248 gnd.n3247 585
R2269 gnd.n2440 gnd.n2438 585
R2270 gnd.n2438 gnd.n2435 585
R2271 gnd.n3240 gnd.n3239 585
R2272 gnd.n3239 gnd.n3238 585
R2273 gnd.n2443 gnd.n2442 585
R2274 gnd.n2453 gnd.n2443 585
R2275 gnd.n3200 gnd.n2466 585
R2276 gnd.n2466 gnd.n2452 585
R2277 gnd.n3202 gnd.n3201 585
R2278 gnd.n3203 gnd.n3202 585
R2279 gnd.n2467 gnd.n2465 585
R2280 gnd.n2474 gnd.n2465 585
R2281 gnd.n3195 gnd.n3194 585
R2282 gnd.n3194 gnd.n3193 585
R2283 gnd.n2470 gnd.n2469 585
R2284 gnd.n3174 gnd.n2470 585
R2285 gnd.n3160 gnd.n2493 585
R2286 gnd.n2493 gnd.n2483 585
R2287 gnd.n3162 gnd.n3161 585
R2288 gnd.n3163 gnd.n3162 585
R2289 gnd.n2494 gnd.n2492 585
R2290 gnd.n3151 gnd.n2492 585
R2291 gnd.n3155 gnd.n3154 585
R2292 gnd.n3154 gnd.n3153 585
R2293 gnd.n2497 gnd.n2496 585
R2294 gnd.n3106 gnd.n2497 585
R2295 gnd.n2599 gnd.n2598 585
R2296 gnd.n2600 gnd.n2599 585
R2297 gnd.n2579 gnd.n2578 585
R2298 gnd.n2582 gnd.n2579 585
R2299 gnd.n3116 gnd.n3115 585
R2300 gnd.n3115 gnd.n3114 585
R2301 gnd.n3117 gnd.n2573 585
R2302 gnd.n2609 gnd.n2573 585
R2303 gnd.n3119 gnd.n3118 585
R2304 gnd.n3120 gnd.n3119 585
R2305 gnd.n2574 gnd.n2572 585
R2306 gnd.n3084 gnd.n2572 585
R2307 gnd.n3068 gnd.n3067 585
R2308 gnd.n3067 gnd.n2560 585
R2309 gnd.n3069 gnd.n2624 585
R2310 gnd.n2624 gnd.n2559 585
R2311 gnd.n3071 gnd.n3070 585
R2312 gnd.n3072 gnd.n3071 585
R2313 gnd.n2625 gnd.n2623 585
R2314 gnd.n2623 gnd.n2620 585
R2315 gnd.n3060 gnd.n3059 585
R2316 gnd.n3059 gnd.n3058 585
R2317 gnd.n2628 gnd.n2627 585
R2318 gnd.n2635 gnd.n2628 585
R2319 gnd.n3034 gnd.n3033 585
R2320 gnd.n3035 gnd.n3034 585
R2321 gnd.n2647 gnd.n2646 585
R2322 gnd.n2654 gnd.n2646 585
R2323 gnd.n3029 gnd.n3028 585
R2324 gnd.n3028 gnd.n3027 585
R2325 gnd.n2650 gnd.n2649 585
R2326 gnd.n3017 gnd.n2650 585
R2327 gnd.n3004 gnd.n2674 585
R2328 gnd.n2674 gnd.n2673 585
R2329 gnd.n3006 gnd.n3005 585
R2330 gnd.n3007 gnd.n3006 585
R2331 gnd.n2675 gnd.n2672 585
R2332 gnd.n2682 gnd.n2672 585
R2333 gnd.n2999 gnd.n2998 585
R2334 gnd.n2998 gnd.n2997 585
R2335 gnd.n2678 gnd.n2677 585
R2336 gnd.n2986 gnd.n2678 585
R2337 gnd.n2973 gnd.n2699 585
R2338 gnd.n2699 gnd.n2698 585
R2339 gnd.n2975 gnd.n2974 585
R2340 gnd.n2976 gnd.n2975 585
R2341 gnd.n2969 gnd.n2697 585
R2342 gnd.n2968 gnd.n2967 585
R2343 gnd.n2702 gnd.n2701 585
R2344 gnd.n2965 gnd.n2702 585
R2345 gnd.n2724 gnd.n2723 585
R2346 gnd.n2727 gnd.n2726 585
R2347 gnd.n2725 gnd.n2720 585
R2348 gnd.n2732 gnd.n2731 585
R2349 gnd.n2734 gnd.n2733 585
R2350 gnd.n2737 gnd.n2736 585
R2351 gnd.n2735 gnd.n2718 585
R2352 gnd.n2742 gnd.n2741 585
R2353 gnd.n2744 gnd.n2743 585
R2354 gnd.n2747 gnd.n2746 585
R2355 gnd.n2745 gnd.n2716 585
R2356 gnd.n2752 gnd.n2751 585
R2357 gnd.n2756 gnd.n2753 585
R2358 gnd.n2757 gnd.n2694 585
R2359 gnd.n3636 gnd.n2311 585
R2360 gnd.n3703 gnd.n3702 585
R2361 gnd.n3705 gnd.n3704 585
R2362 gnd.n3707 gnd.n3706 585
R2363 gnd.n3709 gnd.n3708 585
R2364 gnd.n3711 gnd.n3710 585
R2365 gnd.n3713 gnd.n3712 585
R2366 gnd.n3715 gnd.n3714 585
R2367 gnd.n3717 gnd.n3716 585
R2368 gnd.n3719 gnd.n3718 585
R2369 gnd.n3721 gnd.n3720 585
R2370 gnd.n3723 gnd.n3722 585
R2371 gnd.n3725 gnd.n3724 585
R2372 gnd.n3728 gnd.n3727 585
R2373 gnd.n3726 gnd.n2299 585
R2374 gnd.n3732 gnd.n2297 585
R2375 gnd.n3734 gnd.n3733 585
R2376 gnd.n3735 gnd.n3734 585
R2377 gnd.n3637 gnd.n2352 585
R2378 gnd.n3637 gnd.n2273 585
R2379 gnd.n3639 gnd.n3638 585
R2380 gnd.n3638 gnd.n2347 585
R2381 gnd.n3635 gnd.n2351 585
R2382 gnd.n3635 gnd.n3634 585
R2383 gnd.n3614 gnd.n2353 585
R2384 gnd.n2365 gnd.n2353 585
R2385 gnd.n3613 gnd.n2363 585
R2386 gnd.n3622 gnd.n2363 585
R2387 gnd.n3347 gnd.n2370 585
R2388 gnd.n3349 gnd.n3347 585
R2389 gnd.n3346 gnd.n3345 585
R2390 gnd.n3346 gnd.n2374 585
R2391 gnd.n3344 gnd.n2376 585
R2392 gnd.n3337 gnd.n2376 585
R2393 gnd.n2389 gnd.n2377 585
R2394 gnd.n2389 gnd.n2381 585
R2395 gnd.n3293 gnd.n2390 585
R2396 gnd.n3327 gnd.n2390 585
R2397 gnd.n3292 gnd.n3291 585
R2398 gnd.n3291 gnd.n2397 585
R2399 gnd.n3290 gnd.n2405 585
R2400 gnd.n3290 gnd.n2396 585
R2401 gnd.n3289 gnd.n2407 585
R2402 gnd.n3289 gnd.n3288 585
R2403 gnd.n3268 gnd.n2406 585
R2404 gnd.n2419 gnd.n2406 585
R2405 gnd.n3267 gnd.n2417 585
R2406 gnd.n3278 gnd.n2417 585
R2407 gnd.n3258 gnd.n2424 585
R2408 gnd.n3259 gnd.n3258 585
R2409 gnd.n3257 gnd.n3256 585
R2410 gnd.n3257 gnd.n2428 585
R2411 gnd.n3255 gnd.n2430 585
R2412 gnd.n3248 gnd.n2430 585
R2413 gnd.n2445 gnd.n2431 585
R2414 gnd.n2445 gnd.n2435 585
R2415 gnd.n3208 gnd.n2446 585
R2416 gnd.n3238 gnd.n2446 585
R2417 gnd.n3207 gnd.n3206 585
R2418 gnd.n3206 gnd.n2453 585
R2419 gnd.n3205 gnd.n2460 585
R2420 gnd.n3205 gnd.n2452 585
R2421 gnd.n3204 gnd.n2462 585
R2422 gnd.n3204 gnd.n3203 585
R2423 gnd.n3183 gnd.n2461 585
R2424 gnd.n2474 gnd.n2461 585
R2425 gnd.n3182 gnd.n2472 585
R2426 gnd.n3193 gnd.n2472 585
R2427 gnd.n3173 gnd.n2479 585
R2428 gnd.n3174 gnd.n3173 585
R2429 gnd.n3172 gnd.n3171 585
R2430 gnd.n3172 gnd.n2483 585
R2431 gnd.n3170 gnd.n2485 585
R2432 gnd.n3163 gnd.n2485 585
R2433 gnd.n3150 gnd.n2486 585
R2434 gnd.n3151 gnd.n3150 585
R2435 gnd.n3103 gnd.n2499 585
R2436 gnd.n3153 gnd.n2499 585
R2437 gnd.n3105 gnd.n3104 585
R2438 gnd.n3106 gnd.n3105 585
R2439 gnd.n3098 gnd.n2601 585
R2440 gnd.n2601 gnd.n2600 585
R2441 gnd.n3096 gnd.n3095 585
R2442 gnd.n3095 gnd.n2582 585
R2443 gnd.n3093 gnd.n2580 585
R2444 gnd.n3114 gnd.n2580 585
R2445 gnd.n2611 gnd.n2610 585
R2446 gnd.n2610 gnd.n2609 585
R2447 gnd.n3087 gnd.n2570 585
R2448 gnd.n3120 gnd.n2570 585
R2449 gnd.n3086 gnd.n3085 585
R2450 gnd.n3085 gnd.n3084 585
R2451 gnd.n3082 gnd.n2613 585
R2452 gnd.n3082 gnd.n2560 585
R2453 gnd.n3081 gnd.n3080 585
R2454 gnd.n3081 gnd.n2559 585
R2455 gnd.n2616 gnd.n2615 585
R2456 gnd.n3072 gnd.n2615 585
R2457 gnd.n3040 gnd.n3039 585
R2458 gnd.n3039 gnd.n2620 585
R2459 gnd.n3041 gnd.n2629 585
R2460 gnd.n3058 gnd.n2629 585
R2461 gnd.n3038 gnd.n3037 585
R2462 gnd.n3037 gnd.n2635 585
R2463 gnd.n3036 gnd.n2643 585
R2464 gnd.n3036 gnd.n3035 585
R2465 gnd.n3021 gnd.n2644 585
R2466 gnd.n2654 gnd.n2644 585
R2467 gnd.n3020 gnd.n2652 585
R2468 gnd.n3027 gnd.n2652 585
R2469 gnd.n3019 gnd.n3018 585
R2470 gnd.n3018 gnd.n3017 585
R2471 gnd.n2663 gnd.n2660 585
R2472 gnd.n2673 gnd.n2663 585
R2473 gnd.n3009 gnd.n3008 585
R2474 gnd.n3008 gnd.n3007 585
R2475 gnd.n2669 gnd.n2668 585
R2476 gnd.n2682 gnd.n2669 585
R2477 gnd.n2989 gnd.n2680 585
R2478 gnd.n2997 gnd.n2680 585
R2479 gnd.n2988 gnd.n2987 585
R2480 gnd.n2987 gnd.n2986 585
R2481 gnd.n2689 gnd.n2687 585
R2482 gnd.n2698 gnd.n2689 585
R2483 gnd.n2978 gnd.n2977 585
R2484 gnd.n2977 gnd.n2976 585
R2485 gnd.n5347 gnd.n1714 585
R2486 gnd.n1714 gnd.n1700 585
R2487 gnd.n5349 gnd.n5348 585
R2488 gnd.n5350 gnd.n5349 585
R2489 gnd.n1715 gnd.n1713 585
R2490 gnd.n1713 gnd.n1708 585
R2491 gnd.n5218 gnd.n5217 585
R2492 gnd.n5219 gnd.n5218 585
R2493 gnd.n5216 gnd.n1788 585
R2494 gnd.n1793 gnd.n1788 585
R2495 gnd.n5215 gnd.n5214 585
R2496 gnd.n5214 gnd.n5213 585
R2497 gnd.n1790 gnd.n1789 585
R2498 gnd.n5190 gnd.n1790 585
R2499 gnd.n5202 gnd.n5201 585
R2500 gnd.n5203 gnd.n5202 585
R2501 gnd.n5200 gnd.n1803 585
R2502 gnd.n5196 gnd.n1803 585
R2503 gnd.n5199 gnd.n5198 585
R2504 gnd.n5198 gnd.n5197 585
R2505 gnd.n1805 gnd.n1804 585
R2506 gnd.n5184 gnd.n1805 585
R2507 gnd.n5170 gnd.n5169 585
R2508 gnd.n5169 gnd.n5168 585
R2509 gnd.n5171 gnd.n1822 585
R2510 gnd.n5167 gnd.n1822 585
R2511 gnd.n5173 gnd.n5172 585
R2512 gnd.n5174 gnd.n5173 585
R2513 gnd.n1823 gnd.n1821 585
R2514 gnd.n1821 gnd.n1816 585
R2515 gnd.n5159 gnd.n5158 585
R2516 gnd.n5160 gnd.n5159 585
R2517 gnd.n5157 gnd.n1827 585
R2518 gnd.n1832 gnd.n1827 585
R2519 gnd.n5156 gnd.n5155 585
R2520 gnd.n5155 gnd.n5154 585
R2521 gnd.n1829 gnd.n1828 585
R2522 gnd.n1841 gnd.n1829 585
R2523 gnd.n5143 gnd.n5142 585
R2524 gnd.n5144 gnd.n5143 585
R2525 gnd.n5141 gnd.n1842 585
R2526 gnd.n1842 gnd.n1838 585
R2527 gnd.n5140 gnd.n5139 585
R2528 gnd.n5139 gnd.n5138 585
R2529 gnd.n1844 gnd.n1843 585
R2530 gnd.n1845 gnd.n1844 585
R2531 gnd.n5079 gnd.n1868 585
R2532 gnd.n5079 gnd.n5078 585
R2533 gnd.n5081 gnd.n5080 585
R2534 gnd.n5080 gnd.n1853 585
R2535 gnd.n5082 gnd.n1866 585
R2536 gnd.n5062 gnd.n1866 585
R2537 gnd.n5084 gnd.n5083 585
R2538 gnd.n5085 gnd.n5084 585
R2539 gnd.n1867 gnd.n1865 585
R2540 gnd.n1865 gnd.n1861 585
R2541 gnd.n5056 gnd.n5055 585
R2542 gnd.n5057 gnd.n5056 585
R2543 gnd.n5054 gnd.n1874 585
R2544 gnd.n1880 gnd.n1874 585
R2545 gnd.n5053 gnd.n5052 585
R2546 gnd.n5052 gnd.n5051 585
R2547 gnd.n1876 gnd.n1875 585
R2548 gnd.n1877 gnd.n1876 585
R2549 gnd.n5040 gnd.n5039 585
R2550 gnd.n5041 gnd.n5040 585
R2551 gnd.n5038 gnd.n1890 585
R2552 gnd.n1890 gnd.n1887 585
R2553 gnd.n5037 gnd.n5036 585
R2554 gnd.n5036 gnd.n5035 585
R2555 gnd.n1892 gnd.n1891 585
R2556 gnd.n1899 gnd.n1892 585
R2557 gnd.n5022 gnd.n5021 585
R2558 gnd.n5023 gnd.n5022 585
R2559 gnd.n5020 gnd.n1902 585
R2560 gnd.n1902 gnd.n1898 585
R2561 gnd.n5019 gnd.n5018 585
R2562 gnd.n5018 gnd.n5017 585
R2563 gnd.n1904 gnd.n1903 585
R2564 gnd.n1916 gnd.n1904 585
R2565 gnd.n5004 gnd.n5003 585
R2566 gnd.n5005 gnd.n5004 585
R2567 gnd.n5002 gnd.n1917 585
R2568 gnd.n1917 gnd.n1913 585
R2569 gnd.n5001 gnd.n5000 585
R2570 gnd.n5000 gnd.n4999 585
R2571 gnd.n1919 gnd.n1918 585
R2572 gnd.n4939 gnd.n1919 585
R2573 gnd.n1942 gnd.n1941 585
R2574 gnd.n1942 gnd.n1928 585
R2575 gnd.n4947 gnd.n4946 585
R2576 gnd.n4946 gnd.n4945 585
R2577 gnd.n4948 gnd.n1939 585
R2578 gnd.n1939 gnd.n1937 585
R2579 gnd.n4950 gnd.n4949 585
R2580 gnd.n4951 gnd.n4950 585
R2581 gnd.n1940 gnd.n1938 585
R2582 gnd.n4927 gnd.n1938 585
R2583 gnd.n1970 gnd.n1969 585
R2584 gnd.n1969 gnd.n1948 585
R2585 gnd.n1972 gnd.n1971 585
R2586 gnd.n4897 gnd.n1972 585
R2587 gnd.n4900 gnd.n1968 585
R2588 gnd.n4900 gnd.n4899 585
R2589 gnd.n4902 gnd.n4901 585
R2590 gnd.n4901 gnd.n1955 585
R2591 gnd.n4903 gnd.n1966 585
R2592 gnd.n4890 gnd.n1966 585
R2593 gnd.n4905 gnd.n4904 585
R2594 gnd.n4906 gnd.n4905 585
R2595 gnd.n1967 gnd.n1965 585
R2596 gnd.n1965 gnd.n1962 585
R2597 gnd.n4881 gnd.n4880 585
R2598 gnd.n4882 gnd.n4881 585
R2599 gnd.n4879 gnd.n1977 585
R2600 gnd.n1982 gnd.n1977 585
R2601 gnd.n4878 gnd.n4877 585
R2602 gnd.n4877 gnd.n4876 585
R2603 gnd.n1979 gnd.n1978 585
R2604 gnd.n4853 gnd.n1979 585
R2605 gnd.n4865 gnd.n4864 585
R2606 gnd.n4866 gnd.n4865 585
R2607 gnd.n4863 gnd.n1991 585
R2608 gnd.n1991 gnd.n1988 585
R2609 gnd.n4862 gnd.n4861 585
R2610 gnd.n4861 gnd.n4860 585
R2611 gnd.n1993 gnd.n1992 585
R2612 gnd.n2006 gnd.n1993 585
R2613 gnd.n4823 gnd.n4822 585
R2614 gnd.n4822 gnd.n2005 585
R2615 gnd.n4824 gnd.n2016 585
R2616 gnd.n4766 gnd.n2016 585
R2617 gnd.n4826 gnd.n4825 585
R2618 gnd.n4827 gnd.n4826 585
R2619 gnd.n4821 gnd.n2015 585
R2620 gnd.n2015 gnd.n2012 585
R2621 gnd.n4820 gnd.n4819 585
R2622 gnd.n4819 gnd.n4818 585
R2623 gnd.n2018 gnd.n2017 585
R2624 gnd.n4760 gnd.n2018 585
R2625 gnd.n4789 gnd.n4788 585
R2626 gnd.n4789 gnd.n2027 585
R2627 gnd.n4791 gnd.n4790 585
R2628 gnd.n4790 gnd.n2026 585
R2629 gnd.n4792 gnd.n2041 585
R2630 gnd.n4777 gnd.n2041 585
R2631 gnd.n4794 gnd.n4793 585
R2632 gnd.n4795 gnd.n4794 585
R2633 gnd.n4787 gnd.n2040 585
R2634 gnd.n2040 gnd.n2036 585
R2635 gnd.n4786 gnd.n4785 585
R2636 gnd.n4785 gnd.n4784 585
R2637 gnd.n2043 gnd.n2042 585
R2638 gnd.n2050 gnd.n2043 585
R2639 gnd.n4753 gnd.n4752 585
R2640 gnd.n4754 gnd.n4753 585
R2641 gnd.n4751 gnd.n2052 585
R2642 gnd.n2052 gnd.n2049 585
R2643 gnd.n4750 gnd.n4749 585
R2644 gnd.n4749 gnd.n4748 585
R2645 gnd.n2054 gnd.n2053 585
R2646 gnd.n4672 gnd.n2054 585
R2647 gnd.n1275 gnd.n1274 585
R2648 gnd.n1279 gnd.n1275 585
R2649 gnd.n5834 gnd.n5833 585
R2650 gnd.n5833 gnd.n5832 585
R2651 gnd.n5835 gnd.n1253 585
R2652 gnd.n4739 gnd.n1253 585
R2653 gnd.n5900 gnd.n5899 585
R2654 gnd.n5898 gnd.n1252 585
R2655 gnd.n5897 gnd.n1251 585
R2656 gnd.n5902 gnd.n1251 585
R2657 gnd.n5896 gnd.n5895 585
R2658 gnd.n5894 gnd.n5893 585
R2659 gnd.n5892 gnd.n5891 585
R2660 gnd.n5890 gnd.n5889 585
R2661 gnd.n5888 gnd.n5887 585
R2662 gnd.n5886 gnd.n5885 585
R2663 gnd.n5884 gnd.n5883 585
R2664 gnd.n5882 gnd.n5881 585
R2665 gnd.n5880 gnd.n5879 585
R2666 gnd.n5878 gnd.n5877 585
R2667 gnd.n5876 gnd.n5875 585
R2668 gnd.n5874 gnd.n5873 585
R2669 gnd.n5872 gnd.n5871 585
R2670 gnd.n5870 gnd.n5869 585
R2671 gnd.n5868 gnd.n5867 585
R2672 gnd.n5866 gnd.n5865 585
R2673 gnd.n5864 gnd.n5863 585
R2674 gnd.n5862 gnd.n5861 585
R2675 gnd.n5860 gnd.n5859 585
R2676 gnd.n5858 gnd.n5857 585
R2677 gnd.n5856 gnd.n5855 585
R2678 gnd.n5854 gnd.n5853 585
R2679 gnd.n5852 gnd.n5851 585
R2680 gnd.n5850 gnd.n5849 585
R2681 gnd.n5848 gnd.n5847 585
R2682 gnd.n5846 gnd.n5845 585
R2683 gnd.n5844 gnd.n5843 585
R2684 gnd.n5842 gnd.n5841 585
R2685 gnd.n5840 gnd.n1215 585
R2686 gnd.n5905 gnd.n5904 585
R2687 gnd.n1217 gnd.n1214 585
R2688 gnd.n4677 gnd.n4676 585
R2689 gnd.n4679 gnd.n4678 585
R2690 gnd.n4682 gnd.n4681 585
R2691 gnd.n4684 gnd.n4683 585
R2692 gnd.n4686 gnd.n4685 585
R2693 gnd.n4688 gnd.n4687 585
R2694 gnd.n4690 gnd.n4689 585
R2695 gnd.n4692 gnd.n4691 585
R2696 gnd.n4694 gnd.n4693 585
R2697 gnd.n4696 gnd.n4695 585
R2698 gnd.n4698 gnd.n4697 585
R2699 gnd.n4700 gnd.n4699 585
R2700 gnd.n4702 gnd.n4701 585
R2701 gnd.n4704 gnd.n4703 585
R2702 gnd.n4706 gnd.n4705 585
R2703 gnd.n4708 gnd.n4707 585
R2704 gnd.n4710 gnd.n4709 585
R2705 gnd.n4712 gnd.n4711 585
R2706 gnd.n4714 gnd.n4713 585
R2707 gnd.n4716 gnd.n4715 585
R2708 gnd.n4718 gnd.n4717 585
R2709 gnd.n4720 gnd.n4719 585
R2710 gnd.n4722 gnd.n4721 585
R2711 gnd.n4724 gnd.n4723 585
R2712 gnd.n4726 gnd.n4725 585
R2713 gnd.n4728 gnd.n4727 585
R2714 gnd.n4730 gnd.n4729 585
R2715 gnd.n4732 gnd.n4731 585
R2716 gnd.n4734 gnd.n4733 585
R2717 gnd.n4736 gnd.n4735 585
R2718 gnd.n4738 gnd.n4737 585
R2719 gnd.n5228 gnd.n5227 585
R2720 gnd.n5229 gnd.n1784 585
R2721 gnd.n5231 gnd.n5230 585
R2722 gnd.n5233 gnd.n1782 585
R2723 gnd.n5235 gnd.n5234 585
R2724 gnd.n5236 gnd.n1781 585
R2725 gnd.n5238 gnd.n5237 585
R2726 gnd.n5240 gnd.n1779 585
R2727 gnd.n5242 gnd.n5241 585
R2728 gnd.n5243 gnd.n1778 585
R2729 gnd.n5245 gnd.n5244 585
R2730 gnd.n5247 gnd.n1776 585
R2731 gnd.n5249 gnd.n5248 585
R2732 gnd.n5250 gnd.n1775 585
R2733 gnd.n5252 gnd.n5251 585
R2734 gnd.n5254 gnd.n1773 585
R2735 gnd.n5256 gnd.n5255 585
R2736 gnd.n5257 gnd.n1772 585
R2737 gnd.n5259 gnd.n5258 585
R2738 gnd.n5261 gnd.n1770 585
R2739 gnd.n5263 gnd.n5262 585
R2740 gnd.n5264 gnd.n1769 585
R2741 gnd.n5266 gnd.n5265 585
R2742 gnd.n5268 gnd.n1767 585
R2743 gnd.n5270 gnd.n5269 585
R2744 gnd.n5271 gnd.n1766 585
R2745 gnd.n5273 gnd.n5272 585
R2746 gnd.n5275 gnd.n1764 585
R2747 gnd.n5277 gnd.n5276 585
R2748 gnd.n5279 gnd.n1761 585
R2749 gnd.n5281 gnd.n5280 585
R2750 gnd.n5283 gnd.n1760 585
R2751 gnd.n5284 gnd.n1702 585
R2752 gnd.n5287 gnd.n1521 585
R2753 gnd.n5289 gnd.n5288 585
R2754 gnd.n5291 gnd.n1758 585
R2755 gnd.n5293 gnd.n5292 585
R2756 gnd.n5295 gnd.n1755 585
R2757 gnd.n5297 gnd.n5296 585
R2758 gnd.n5299 gnd.n1753 585
R2759 gnd.n5301 gnd.n5300 585
R2760 gnd.n5302 gnd.n1752 585
R2761 gnd.n5304 gnd.n5303 585
R2762 gnd.n5306 gnd.n1750 585
R2763 gnd.n5308 gnd.n5307 585
R2764 gnd.n5309 gnd.n1749 585
R2765 gnd.n5311 gnd.n5310 585
R2766 gnd.n5313 gnd.n1747 585
R2767 gnd.n5315 gnd.n5314 585
R2768 gnd.n5316 gnd.n1746 585
R2769 gnd.n5318 gnd.n5317 585
R2770 gnd.n5320 gnd.n1744 585
R2771 gnd.n5322 gnd.n5321 585
R2772 gnd.n5323 gnd.n1743 585
R2773 gnd.n5325 gnd.n5324 585
R2774 gnd.n5327 gnd.n1741 585
R2775 gnd.n5329 gnd.n5328 585
R2776 gnd.n5330 gnd.n1740 585
R2777 gnd.n5332 gnd.n5331 585
R2778 gnd.n5334 gnd.n1738 585
R2779 gnd.n5336 gnd.n5335 585
R2780 gnd.n5337 gnd.n1737 585
R2781 gnd.n5339 gnd.n5338 585
R2782 gnd.n5341 gnd.n1736 585
R2783 gnd.n5342 gnd.n1735 585
R2784 gnd.n5345 gnd.n5344 585
R2785 gnd.n5226 gnd.n5224 585
R2786 gnd.n5226 gnd.n1700 585
R2787 gnd.n5223 gnd.n1710 585
R2788 gnd.n5350 gnd.n1710 585
R2789 gnd.n5222 gnd.n5221 585
R2790 gnd.n5221 gnd.n1708 585
R2791 gnd.n5220 gnd.n1785 585
R2792 gnd.n5220 gnd.n5219 585
R2793 gnd.n5188 gnd.n1786 585
R2794 gnd.n1793 gnd.n1786 585
R2795 gnd.n5189 gnd.n1791 585
R2796 gnd.n5213 gnd.n1791 585
R2797 gnd.n5192 gnd.n5191 585
R2798 gnd.n5191 gnd.n5190 585
R2799 gnd.n5193 gnd.n1800 585
R2800 gnd.n5203 gnd.n1800 585
R2801 gnd.n5195 gnd.n5194 585
R2802 gnd.n5196 gnd.n5195 585
R2803 gnd.n5187 gnd.n1807 585
R2804 gnd.n5197 gnd.n1807 585
R2805 gnd.n5186 gnd.n5185 585
R2806 gnd.n5185 gnd.n5184 585
R2807 gnd.n1809 gnd.n1808 585
R2808 gnd.n5168 gnd.n1809 585
R2809 gnd.n5166 gnd.n5165 585
R2810 gnd.n5167 gnd.n5166 585
R2811 gnd.n5164 gnd.n1818 585
R2812 gnd.n5174 gnd.n1818 585
R2813 gnd.n5163 gnd.n5162 585
R2814 gnd.n5162 gnd.n1816 585
R2815 gnd.n5161 gnd.n1824 585
R2816 gnd.n5161 gnd.n5160 585
R2817 gnd.n5066 gnd.n1825 585
R2818 gnd.n1832 gnd.n1825 585
R2819 gnd.n5067 gnd.n1830 585
R2820 gnd.n5154 gnd.n1830 585
R2821 gnd.n5069 gnd.n5068 585
R2822 gnd.n5068 gnd.n1841 585
R2823 gnd.n5070 gnd.n1840 585
R2824 gnd.n5144 gnd.n1840 585
R2825 gnd.n5072 gnd.n5071 585
R2826 gnd.n5071 gnd.n1838 585
R2827 gnd.n5073 gnd.n1846 585
R2828 gnd.n5138 gnd.n1846 585
R2829 gnd.n5074 gnd.n1870 585
R2830 gnd.n1870 gnd.n1845 585
R2831 gnd.n5076 gnd.n5075 585
R2832 gnd.n5078 gnd.n5076 585
R2833 gnd.n5065 gnd.n1869 585
R2834 gnd.n1869 gnd.n1853 585
R2835 gnd.n5064 gnd.n5063 585
R2836 gnd.n5063 gnd.n5062 585
R2837 gnd.n5061 gnd.n1863 585
R2838 gnd.n5085 gnd.n1863 585
R2839 gnd.n5060 gnd.n5059 585
R2840 gnd.n5059 gnd.n1861 585
R2841 gnd.n5058 gnd.n1871 585
R2842 gnd.n5058 gnd.n5057 585
R2843 gnd.n5027 gnd.n1872 585
R2844 gnd.n1880 gnd.n1872 585
R2845 gnd.n5028 gnd.n1878 585
R2846 gnd.n5051 gnd.n1878 585
R2847 gnd.n5030 gnd.n5029 585
R2848 gnd.n5029 gnd.n1877 585
R2849 gnd.n5031 gnd.n1889 585
R2850 gnd.n5041 gnd.n1889 585
R2851 gnd.n5032 gnd.n1895 585
R2852 gnd.n1895 gnd.n1887 585
R2853 gnd.n5034 gnd.n5033 585
R2854 gnd.n5035 gnd.n5034 585
R2855 gnd.n5026 gnd.n1894 585
R2856 gnd.n1899 gnd.n1894 585
R2857 gnd.n5025 gnd.n5024 585
R2858 gnd.n5024 gnd.n5023 585
R2859 gnd.n1897 gnd.n1896 585
R2860 gnd.n1898 gnd.n1897 585
R2861 gnd.n4932 gnd.n1905 585
R2862 gnd.n5017 gnd.n1905 585
R2863 gnd.n4934 gnd.n4933 585
R2864 gnd.n4933 gnd.n1916 585
R2865 gnd.n4935 gnd.n1915 585
R2866 gnd.n5005 gnd.n1915 585
R2867 gnd.n4937 gnd.n4936 585
R2868 gnd.n4936 gnd.n1913 585
R2869 gnd.n4938 gnd.n1921 585
R2870 gnd.n4999 gnd.n1921 585
R2871 gnd.n4941 gnd.n4940 585
R2872 gnd.n4940 gnd.n4939 585
R2873 gnd.n4942 gnd.n1945 585
R2874 gnd.n1945 gnd.n1928 585
R2875 gnd.n4944 gnd.n4943 585
R2876 gnd.n4945 gnd.n4944 585
R2877 gnd.n4931 gnd.n1944 585
R2878 gnd.n1944 gnd.n1937 585
R2879 gnd.n4930 gnd.n1936 585
R2880 gnd.n4951 gnd.n1936 585
R2881 gnd.n4929 gnd.n4928 585
R2882 gnd.n4928 gnd.n4927 585
R2883 gnd.n1947 gnd.n1946 585
R2884 gnd.n1948 gnd.n1947 585
R2885 gnd.n4896 gnd.n4895 585
R2886 gnd.n4897 gnd.n4896 585
R2887 gnd.n4894 gnd.n1973 585
R2888 gnd.n4899 gnd.n1973 585
R2889 gnd.n4893 gnd.n4892 585
R2890 gnd.n4892 gnd.n1955 585
R2891 gnd.n4891 gnd.n4887 585
R2892 gnd.n4891 gnd.n4890 585
R2893 gnd.n4886 gnd.n1964 585
R2894 gnd.n4906 gnd.n1964 585
R2895 gnd.n4885 gnd.n4884 585
R2896 gnd.n4884 gnd.n1962 585
R2897 gnd.n4883 gnd.n1974 585
R2898 gnd.n4883 gnd.n4882 585
R2899 gnd.n1998 gnd.n1975 585
R2900 gnd.n1982 gnd.n1975 585
R2901 gnd.n1999 gnd.n1980 585
R2902 gnd.n4876 gnd.n1980 585
R2903 gnd.n4855 gnd.n4854 585
R2904 gnd.n4854 gnd.n4853 585
R2905 gnd.n4856 gnd.n1990 585
R2906 gnd.n4866 gnd.n1990 585
R2907 gnd.n4857 gnd.n1996 585
R2908 gnd.n1996 gnd.n1988 585
R2909 gnd.n4859 gnd.n4858 585
R2910 gnd.n4860 gnd.n4859 585
R2911 gnd.n1997 gnd.n1995 585
R2912 gnd.n2006 gnd.n1995 585
R2913 gnd.n4763 gnd.n4762 585
R2914 gnd.n4763 gnd.n2005 585
R2915 gnd.n4768 gnd.n4767 585
R2916 gnd.n4767 gnd.n4766 585
R2917 gnd.n4769 gnd.n2014 585
R2918 gnd.n4827 gnd.n2014 585
R2919 gnd.n4771 gnd.n4770 585
R2920 gnd.n4770 gnd.n2012 585
R2921 gnd.n4772 gnd.n2019 585
R2922 gnd.n4818 gnd.n2019 585
R2923 gnd.n4773 gnd.n4761 585
R2924 gnd.n4761 gnd.n4760 585
R2925 gnd.n4775 gnd.n4774 585
R2926 gnd.n4775 gnd.n2027 585
R2927 gnd.n4776 gnd.n4758 585
R2928 gnd.n4776 gnd.n2026 585
R2929 gnd.n4779 gnd.n4778 585
R2930 gnd.n4778 gnd.n4777 585
R2931 gnd.n4780 gnd.n2038 585
R2932 gnd.n4795 gnd.n2038 585
R2933 gnd.n4781 gnd.n2046 585
R2934 gnd.n2046 gnd.n2036 585
R2935 gnd.n4783 gnd.n4782 585
R2936 gnd.n4784 gnd.n4783 585
R2937 gnd.n4757 gnd.n2045 585
R2938 gnd.n2050 gnd.n2045 585
R2939 gnd.n4756 gnd.n4755 585
R2940 gnd.n4755 gnd.n4754 585
R2941 gnd.n2048 gnd.n2047 585
R2942 gnd.n2049 gnd.n2048 585
R2943 gnd.n4747 gnd.n4746 585
R2944 gnd.n4748 gnd.n4747 585
R2945 gnd.n4745 gnd.n4673 585
R2946 gnd.n4673 gnd.n4672 585
R2947 gnd.n4744 gnd.n4743 585
R2948 gnd.n4743 gnd.n1279 585
R2949 gnd.n4742 gnd.n1277 585
R2950 gnd.n5832 gnd.n1277 585
R2951 gnd.n4741 gnd.n4740 585
R2952 gnd.n4740 gnd.n4739 585
R2953 gnd.n5961 gnd.n1138 585
R2954 gnd.n4569 gnd.n1138 585
R2955 gnd.n5963 gnd.n5962 585
R2956 gnd.n5964 gnd.n5963 585
R2957 gnd.n1123 gnd.n1122 585
R2958 gnd.n4529 gnd.n1123 585
R2959 gnd.n5972 gnd.n5971 585
R2960 gnd.n5971 gnd.n5970 585
R2961 gnd.n5973 gnd.n1117 585
R2962 gnd.n4267 gnd.n1117 585
R2963 gnd.n5975 gnd.n5974 585
R2964 gnd.n5976 gnd.n5975 585
R2965 gnd.n1103 gnd.n1102 585
R2966 gnd.n4542 gnd.n1103 585
R2967 gnd.n5984 gnd.n5983 585
R2968 gnd.n5983 gnd.n5982 585
R2969 gnd.n5985 gnd.n1097 585
R2970 gnd.n4260 gnd.n1097 585
R2971 gnd.n5987 gnd.n5986 585
R2972 gnd.n5988 gnd.n5987 585
R2973 gnd.n1083 gnd.n1082 585
R2974 gnd.n4252 gnd.n1083 585
R2975 gnd.n5996 gnd.n5995 585
R2976 gnd.n5995 gnd.n5994 585
R2977 gnd.n5997 gnd.n1077 585
R2978 gnd.n4217 gnd.n1077 585
R2979 gnd.n5999 gnd.n5998 585
R2980 gnd.n6000 gnd.n5999 585
R2981 gnd.n1061 gnd.n1060 585
R2982 gnd.n4225 gnd.n1061 585
R2983 gnd.n6008 gnd.n6007 585
R2984 gnd.n6007 gnd.n6006 585
R2985 gnd.n6009 gnd.n1056 585
R2986 gnd.n4206 gnd.n1056 585
R2987 gnd.n6011 gnd.n6010 585
R2988 gnd.n6012 gnd.n6011 585
R2989 gnd.n4194 gnd.n1055 585
R2990 gnd.n1055 gnd.n1050 585
R2991 gnd.n4196 gnd.n4195 585
R2992 gnd.n4197 gnd.n4196 585
R2993 gnd.n4192 gnd.n2166 585
R2994 gnd.n2172 gnd.n2166 585
R2995 gnd.n4191 gnd.n4190 585
R2996 gnd.n4190 gnd.n4189 585
R2997 gnd.n4167 gnd.n2168 585
R2998 gnd.n2169 gnd.n2168 585
R2999 gnd.n4169 gnd.n4168 585
R3000 gnd.n4170 gnd.n4169 585
R3001 gnd.n4165 gnd.n2185 585
R3002 gnd.n2185 gnd.n2182 585
R3003 gnd.n4164 gnd.n4163 585
R3004 gnd.n4163 gnd.n4162 585
R3005 gnd.n4147 gnd.n2187 585
R3006 gnd.n2188 gnd.n2187 585
R3007 gnd.n4149 gnd.n4148 585
R3008 gnd.n4150 gnd.n4149 585
R3009 gnd.n2201 gnd.n2200 585
R3010 gnd.n2208 gnd.n2200 585
R3011 gnd.n4143 gnd.n4142 585
R3012 gnd.n4142 gnd.n4141 585
R3013 gnd.n2204 gnd.n2203 585
R3014 gnd.n2205 gnd.n2204 585
R3015 gnd.n4128 gnd.n4127 585
R3016 gnd.n4129 gnd.n4128 585
R3017 gnd.n2220 gnd.n2219 585
R3018 gnd.n2219 gnd.n2216 585
R3019 gnd.n4123 gnd.n4122 585
R3020 gnd.n4122 gnd.n4121 585
R3021 gnd.n2223 gnd.n2222 585
R3022 gnd.n2224 gnd.n2223 585
R3023 gnd.n4108 gnd.n4107 585
R3024 gnd.n4109 gnd.n4108 585
R3025 gnd.n2237 gnd.n2236 585
R3026 gnd.n2244 gnd.n2236 585
R3027 gnd.n4103 gnd.n4102 585
R3028 gnd.n4102 gnd.n4101 585
R3029 gnd.n2240 gnd.n2239 585
R3030 gnd.n2241 gnd.n2240 585
R3031 gnd.n4088 gnd.n4087 585
R3032 gnd.n4089 gnd.n4088 585
R3033 gnd.n2256 gnd.n2255 585
R3034 gnd.n2255 gnd.n2252 585
R3035 gnd.n4083 gnd.n4082 585
R3036 gnd.n4082 gnd.n4081 585
R3037 gnd.n2259 gnd.n2258 585
R3038 gnd.n2260 gnd.n2259 585
R3039 gnd.n4069 gnd.n4068 585
R3040 gnd.n4067 gnd.n3774 585
R3041 gnd.n4066 gnd.n3773 585
R3042 gnd.n4071 gnd.n3773 585
R3043 gnd.n4065 gnd.n4064 585
R3044 gnd.n4063 gnd.n4062 585
R3045 gnd.n4061 gnd.n4060 585
R3046 gnd.n4059 gnd.n4058 585
R3047 gnd.n4057 gnd.n4056 585
R3048 gnd.n4055 gnd.n4054 585
R3049 gnd.n4053 gnd.n4052 585
R3050 gnd.n4051 gnd.n4050 585
R3051 gnd.n4049 gnd.n4048 585
R3052 gnd.n4047 gnd.n4046 585
R3053 gnd.n4045 gnd.n4044 585
R3054 gnd.n4043 gnd.n4042 585
R3055 gnd.n4041 gnd.n4040 585
R3056 gnd.n4039 gnd.n4038 585
R3057 gnd.n4037 gnd.n4036 585
R3058 gnd.n4034 gnd.n4033 585
R3059 gnd.n4032 gnd.n4031 585
R3060 gnd.n4030 gnd.n4029 585
R3061 gnd.n4028 gnd.n4027 585
R3062 gnd.n4026 gnd.n4025 585
R3063 gnd.n4024 gnd.n4023 585
R3064 gnd.n4022 gnd.n4021 585
R3065 gnd.n4020 gnd.n4019 585
R3066 gnd.n4018 gnd.n4017 585
R3067 gnd.n4016 gnd.n4015 585
R3068 gnd.n4014 gnd.n4013 585
R3069 gnd.n4012 gnd.n4011 585
R3070 gnd.n4010 gnd.n4009 585
R3071 gnd.n4008 gnd.n4007 585
R3072 gnd.n4006 gnd.n4005 585
R3073 gnd.n4004 gnd.n4003 585
R3074 gnd.n4002 gnd.n4001 585
R3075 gnd.n4000 gnd.n3999 585
R3076 gnd.n3998 gnd.n3997 585
R3077 gnd.n3996 gnd.n3995 585
R3078 gnd.n3994 gnd.n3993 585
R3079 gnd.n3992 gnd.n3991 585
R3080 gnd.n3990 gnd.n3989 585
R3081 gnd.n3988 gnd.n3987 585
R3082 gnd.n3986 gnd.n3985 585
R3083 gnd.n3984 gnd.n3983 585
R3084 gnd.n3982 gnd.n3981 585
R3085 gnd.n3980 gnd.n3979 585
R3086 gnd.n3978 gnd.n3977 585
R3087 gnd.n3976 gnd.n3975 585
R3088 gnd.n3974 gnd.n3973 585
R3089 gnd.n3972 gnd.n3971 585
R3090 gnd.n3970 gnd.n3969 585
R3091 gnd.n3968 gnd.n3967 585
R3092 gnd.n3966 gnd.n3965 585
R3093 gnd.n3964 gnd.n3963 585
R3094 gnd.n3962 gnd.n3961 585
R3095 gnd.n3960 gnd.n3959 585
R3096 gnd.n3958 gnd.n3957 585
R3097 gnd.n3956 gnd.n2272 585
R3098 gnd.n4073 gnd.n2271 585
R3099 gnd.n4521 gnd.n4520 585
R3100 gnd.n4519 gnd.n4430 585
R3101 gnd.n4518 gnd.n4517 585
R3102 gnd.n4511 gnd.n4431 585
R3103 gnd.n4513 gnd.n4512 585
R3104 gnd.n4510 gnd.n4509 585
R3105 gnd.n4508 gnd.n4507 585
R3106 gnd.n4501 gnd.n4433 585
R3107 gnd.n4503 gnd.n4502 585
R3108 gnd.n4500 gnd.n4499 585
R3109 gnd.n4498 gnd.n4497 585
R3110 gnd.n4491 gnd.n4435 585
R3111 gnd.n4493 gnd.n4492 585
R3112 gnd.n4490 gnd.n4489 585
R3113 gnd.n4488 gnd.n4487 585
R3114 gnd.n4481 gnd.n4437 585
R3115 gnd.n4483 gnd.n4482 585
R3116 gnd.n4480 gnd.n4479 585
R3117 gnd.n4478 gnd.n4477 585
R3118 gnd.n4471 gnd.n4439 585
R3119 gnd.n4473 gnd.n4472 585
R3120 gnd.n4470 gnd.n4443 585
R3121 gnd.n4469 gnd.n4468 585
R3122 gnd.n4462 gnd.n4444 585
R3123 gnd.n4464 gnd.n4463 585
R3124 gnd.n4461 gnd.n4460 585
R3125 gnd.n4459 gnd.n4458 585
R3126 gnd.n4452 gnd.n4446 585
R3127 gnd.n4454 gnd.n4453 585
R3128 gnd.n4451 gnd.n4450 585
R3129 gnd.n4449 gnd.n1211 585
R3130 gnd.n5908 gnd.n5907 585
R3131 gnd.n5910 gnd.n5909 585
R3132 gnd.n5912 gnd.n5911 585
R3133 gnd.n5914 gnd.n5913 585
R3134 gnd.n5916 gnd.n5915 585
R3135 gnd.n5918 gnd.n5917 585
R3136 gnd.n5920 gnd.n5919 585
R3137 gnd.n5922 gnd.n5921 585
R3138 gnd.n5925 gnd.n5924 585
R3139 gnd.n5927 gnd.n5926 585
R3140 gnd.n5929 gnd.n5928 585
R3141 gnd.n5931 gnd.n5930 585
R3142 gnd.n5933 gnd.n5932 585
R3143 gnd.n5935 gnd.n5934 585
R3144 gnd.n5937 gnd.n5936 585
R3145 gnd.n5939 gnd.n5938 585
R3146 gnd.n5941 gnd.n5940 585
R3147 gnd.n5943 gnd.n5942 585
R3148 gnd.n5945 gnd.n5944 585
R3149 gnd.n5947 gnd.n5946 585
R3150 gnd.n5949 gnd.n5948 585
R3151 gnd.n5951 gnd.n5950 585
R3152 gnd.n5952 gnd.n1184 585
R3153 gnd.n5954 gnd.n5953 585
R3154 gnd.n1143 gnd.n1142 585
R3155 gnd.n5958 gnd.n5957 585
R3156 gnd.n5957 gnd.n5956 585
R3157 gnd.n4525 gnd.n2126 585
R3158 gnd.n4569 gnd.n2126 585
R3159 gnd.n4526 gnd.n1135 585
R3160 gnd.n5964 gnd.n1135 585
R3161 gnd.n4528 gnd.n4527 585
R3162 gnd.n4529 gnd.n4528 585
R3163 gnd.n4270 gnd.n1125 585
R3164 gnd.n5970 gnd.n1125 585
R3165 gnd.n4269 gnd.n4268 585
R3166 gnd.n4268 gnd.n4267 585
R3167 gnd.n4265 gnd.n1114 585
R3168 gnd.n5976 gnd.n1114 585
R3169 gnd.n4264 gnd.n2137 585
R3170 gnd.n4542 gnd.n2137 585
R3171 gnd.n4263 gnd.n1105 585
R3172 gnd.n5982 gnd.n1105 585
R3173 gnd.n4262 gnd.n4261 585
R3174 gnd.n4261 gnd.n4260 585
R3175 gnd.n2143 gnd.n1094 585
R3176 gnd.n5988 gnd.n1094 585
R3177 gnd.n4213 gnd.n2148 585
R3178 gnd.n4252 gnd.n2148 585
R3179 gnd.n4214 gnd.n1085 585
R3180 gnd.n5994 gnd.n1085 585
R3181 gnd.n4216 gnd.n4215 585
R3182 gnd.n4217 gnd.n4216 585
R3183 gnd.n4211 gnd.n1074 585
R3184 gnd.n6000 gnd.n1074 585
R3185 gnd.n4210 gnd.n2154 585
R3186 gnd.n4225 gnd.n2154 585
R3187 gnd.n4209 gnd.n1063 585
R3188 gnd.n6006 gnd.n1063 585
R3189 gnd.n4208 gnd.n4207 585
R3190 gnd.n4207 gnd.n4206 585
R3191 gnd.n2158 gnd.n1051 585
R3192 gnd.n6012 gnd.n1051 585
R3193 gnd.n4179 gnd.n4178 585
R3194 gnd.n4178 gnd.n1050 585
R3195 gnd.n4177 gnd.n2164 585
R3196 gnd.n4197 gnd.n2164 585
R3197 gnd.n4176 gnd.n4175 585
R3198 gnd.n4175 gnd.n2172 585
R3199 gnd.n4174 gnd.n2170 585
R3200 gnd.n4189 gnd.n2170 585
R3201 gnd.n4173 gnd.n4172 585
R3202 gnd.n4172 gnd.n2169 585
R3203 gnd.n4171 gnd.n2179 585
R3204 gnd.n4171 gnd.n4170 585
R3205 gnd.n4155 gnd.n2181 585
R3206 gnd.n2182 gnd.n2181 585
R3207 gnd.n4154 gnd.n2189 585
R3208 gnd.n4162 gnd.n2189 585
R3209 gnd.n4153 gnd.n4152 585
R3210 gnd.n4152 gnd.n2188 585
R3211 gnd.n4151 gnd.n2195 585
R3212 gnd.n4151 gnd.n4150 585
R3213 gnd.n4134 gnd.n2197 585
R3214 gnd.n2208 gnd.n2197 585
R3215 gnd.n4133 gnd.n2206 585
R3216 gnd.n4141 gnd.n2206 585
R3217 gnd.n4132 gnd.n4131 585
R3218 gnd.n4131 gnd.n2205 585
R3219 gnd.n4130 gnd.n2213 585
R3220 gnd.n4130 gnd.n4129 585
R3221 gnd.n4114 gnd.n2215 585
R3222 gnd.n2216 gnd.n2215 585
R3223 gnd.n4113 gnd.n2225 585
R3224 gnd.n4121 gnd.n2225 585
R3225 gnd.n4112 gnd.n4111 585
R3226 gnd.n4111 gnd.n2224 585
R3227 gnd.n4110 gnd.n2231 585
R3228 gnd.n4110 gnd.n4109 585
R3229 gnd.n4094 gnd.n2233 585
R3230 gnd.n2244 gnd.n2233 585
R3231 gnd.n4093 gnd.n2242 585
R3232 gnd.n4101 gnd.n2242 585
R3233 gnd.n4092 gnd.n4091 585
R3234 gnd.n4091 gnd.n2241 585
R3235 gnd.n4090 gnd.n2249 585
R3236 gnd.n4090 gnd.n4089 585
R3237 gnd.n4076 gnd.n2251 585
R3238 gnd.n2252 gnd.n2251 585
R3239 gnd.n4077 gnd.n2261 585
R3240 gnd.n4081 gnd.n2261 585
R3241 gnd.n4075 gnd.n4074 585
R3242 gnd.n4074 gnd.n2260 585
R3243 gnd.n6843 gnd.n6842 585
R3244 gnd.n6842 gnd.n6841 585
R3245 gnd.n6844 gnd.n156 585
R3246 gnd.n162 gnd.n156 585
R3247 gnd.n6846 gnd.n6845 585
R3248 gnd.n6847 gnd.n6846 585
R3249 gnd.n143 gnd.n142 585
R3250 gnd.n147 gnd.n143 585
R3251 gnd.n6855 gnd.n6854 585
R3252 gnd.n6854 gnd.n6853 585
R3253 gnd.n6856 gnd.n137 585
R3254 gnd.n144 gnd.n137 585
R3255 gnd.n6858 gnd.n6857 585
R3256 gnd.n6859 gnd.n6858 585
R3257 gnd.n123 gnd.n122 585
R3258 gnd.n127 gnd.n123 585
R3259 gnd.n6867 gnd.n6866 585
R3260 gnd.n6866 gnd.n6865 585
R3261 gnd.n6868 gnd.n117 585
R3262 gnd.n124 gnd.n117 585
R3263 gnd.n6870 gnd.n6869 585
R3264 gnd.n6871 gnd.n6870 585
R3265 gnd.n105 gnd.n104 585
R3266 gnd.n114 gnd.n105 585
R3267 gnd.n6879 gnd.n6878 585
R3268 gnd.n6878 gnd.n6877 585
R3269 gnd.n6880 gnd.n100 585
R3270 gnd.n100 gnd.n99 585
R3271 gnd.n6882 gnd.n6881 585
R3272 gnd.n6883 gnd.n6882 585
R3273 gnd.n84 gnd.n82 585
R3274 gnd.n88 gnd.n84 585
R3275 gnd.n6891 gnd.n6890 585
R3276 gnd.n6890 gnd.n6889 585
R3277 gnd.n83 gnd.n75 585
R3278 gnd.n85 gnd.n83 585
R3279 gnd.n6894 gnd.n73 585
R3280 gnd.n73 gnd.n70 585
R3281 gnd.n6896 gnd.n6895 585
R3282 gnd.n6897 gnd.n6896 585
R3283 gnd.n6784 gnd.n72 585
R3284 gnd.n6799 gnd.n72 585
R3285 gnd.n6786 gnd.n6785 585
R3286 gnd.n6786 gnd.n499 585
R3287 gnd.n6789 gnd.n6788 585
R3288 gnd.n6790 gnd.n6789 585
R3289 gnd.n6787 gnd.n6783 585
R3290 gnd.n6783 gnd.n6782 585
R3291 gnd.n6771 gnd.n508 585
R3292 gnd.n509 gnd.n508 585
R3293 gnd.n6773 gnd.n6772 585
R3294 gnd.n6774 gnd.n6773 585
R3295 gnd.n6770 gnd.n521 585
R3296 gnd.n6770 gnd.n6769 585
R3297 gnd.n6743 gnd.n520 585
R3298 gnd.n6755 gnd.n520 585
R3299 gnd.n6744 gnd.n541 585
R3300 gnd.n6729 gnd.n541 585
R3301 gnd.n6746 gnd.n6745 585
R3302 gnd.n6747 gnd.n6746 585
R3303 gnd.n542 gnd.n540 585
R3304 gnd.n1615 gnd.n540 585
R3305 gnd.n6738 gnd.n6737 585
R3306 gnd.n6737 gnd.n6736 585
R3307 gnd.n545 gnd.n544 585
R3308 gnd.n1622 gnd.n545 585
R3309 gnd.n1605 gnd.n1604 585
R3310 gnd.n5499 gnd.n1605 585
R3311 gnd.n5508 gnd.n5507 585
R3312 gnd.n5507 gnd.n5506 585
R3313 gnd.n5509 gnd.n1598 585
R3314 gnd.n5448 gnd.n1598 585
R3315 gnd.n5511 gnd.n5510 585
R3316 gnd.n5512 gnd.n5511 585
R3317 gnd.n1580 gnd.n1579 585
R3318 gnd.n5441 gnd.n1580 585
R3319 gnd.n5520 gnd.n5519 585
R3320 gnd.n5519 gnd.n5518 585
R3321 gnd.n5521 gnd.n1571 585
R3322 gnd.n5435 gnd.n1571 585
R3323 gnd.n5523 gnd.n5522 585
R3324 gnd.n5524 gnd.n5523 585
R3325 gnd.n1572 gnd.n1570 585
R3326 gnd.n5470 gnd.n1570 585
R3327 gnd.n1573 gnd.n1492 585
R3328 gnd.n5532 gnd.n1492 585
R3329 gnd.n5651 gnd.n5650 585
R3330 gnd.n5649 gnd.n1491 585
R3331 gnd.n5648 gnd.n1490 585
R3332 gnd.n5653 gnd.n1490 585
R3333 gnd.n5647 gnd.n5646 585
R3334 gnd.n5645 gnd.n5644 585
R3335 gnd.n5643 gnd.n5642 585
R3336 gnd.n5641 gnd.n5640 585
R3337 gnd.n5639 gnd.n5638 585
R3338 gnd.n5637 gnd.n5636 585
R3339 gnd.n5635 gnd.n5634 585
R3340 gnd.n5633 gnd.n5632 585
R3341 gnd.n5631 gnd.n5630 585
R3342 gnd.n5629 gnd.n5628 585
R3343 gnd.n5627 gnd.n5626 585
R3344 gnd.n5625 gnd.n5624 585
R3345 gnd.n5623 gnd.n5622 585
R3346 gnd.n5621 gnd.n5620 585
R3347 gnd.n5619 gnd.n5618 585
R3348 gnd.n5616 gnd.n5615 585
R3349 gnd.n5614 gnd.n5613 585
R3350 gnd.n5612 gnd.n5611 585
R3351 gnd.n5610 gnd.n5609 585
R3352 gnd.n5608 gnd.n5607 585
R3353 gnd.n5606 gnd.n5605 585
R3354 gnd.n5604 gnd.n5603 585
R3355 gnd.n5602 gnd.n5601 585
R3356 gnd.n5599 gnd.n5598 585
R3357 gnd.n5597 gnd.n5596 585
R3358 gnd.n5595 gnd.n5594 585
R3359 gnd.n5593 gnd.n5592 585
R3360 gnd.n5591 gnd.n5590 585
R3361 gnd.n5589 gnd.n5588 585
R3362 gnd.n5587 gnd.n5586 585
R3363 gnd.n5585 gnd.n5584 585
R3364 gnd.n5583 gnd.n5582 585
R3365 gnd.n5581 gnd.n5580 585
R3366 gnd.n5579 gnd.n5578 585
R3367 gnd.n5577 gnd.n5576 585
R3368 gnd.n5575 gnd.n5574 585
R3369 gnd.n5573 gnd.n5572 585
R3370 gnd.n5571 gnd.n5570 585
R3371 gnd.n5569 gnd.n5568 585
R3372 gnd.n5567 gnd.n5566 585
R3373 gnd.n5565 gnd.n5564 585
R3374 gnd.n5563 gnd.n5562 585
R3375 gnd.n5561 gnd.n5560 585
R3376 gnd.n5559 gnd.n5558 585
R3377 gnd.n5557 gnd.n5556 585
R3378 gnd.n5555 gnd.n5554 585
R3379 gnd.n5553 gnd.n5552 585
R3380 gnd.n5551 gnd.n5550 585
R3381 gnd.n5549 gnd.n5548 585
R3382 gnd.n5547 gnd.n5546 585
R3383 gnd.n5545 gnd.n5544 585
R3384 gnd.n5543 gnd.n5542 585
R3385 gnd.n5541 gnd.n5540 585
R3386 gnd.n5535 gnd.n5534 585
R3387 gnd.n491 gnd.n490 585
R3388 gnd.n488 gnd.n284 585
R3389 gnd.n487 gnd.n486 585
R3390 gnd.n480 gnd.n286 585
R3391 gnd.n482 gnd.n481 585
R3392 gnd.n478 gnd.n288 585
R3393 gnd.n477 gnd.n476 585
R3394 gnd.n470 gnd.n290 585
R3395 gnd.n472 gnd.n471 585
R3396 gnd.n468 gnd.n292 585
R3397 gnd.n467 gnd.n466 585
R3398 gnd.n460 gnd.n294 585
R3399 gnd.n462 gnd.n461 585
R3400 gnd.n458 gnd.n296 585
R3401 gnd.n457 gnd.n456 585
R3402 gnd.n450 gnd.n298 585
R3403 gnd.n452 gnd.n451 585
R3404 gnd.n448 gnd.n300 585
R3405 gnd.n447 gnd.n446 585
R3406 gnd.n440 gnd.n302 585
R3407 gnd.n442 gnd.n441 585
R3408 gnd.n438 gnd.n306 585
R3409 gnd.n437 gnd.n436 585
R3410 gnd.n430 gnd.n308 585
R3411 gnd.n432 gnd.n431 585
R3412 gnd.n428 gnd.n310 585
R3413 gnd.n427 gnd.n426 585
R3414 gnd.n420 gnd.n312 585
R3415 gnd.n422 gnd.n421 585
R3416 gnd.n418 gnd.n314 585
R3417 gnd.n417 gnd.n416 585
R3418 gnd.n410 gnd.n316 585
R3419 gnd.n412 gnd.n411 585
R3420 gnd.n408 gnd.n318 585
R3421 gnd.n407 gnd.n406 585
R3422 gnd.n400 gnd.n320 585
R3423 gnd.n402 gnd.n401 585
R3424 gnd.n398 gnd.n322 585
R3425 gnd.n397 gnd.n396 585
R3426 gnd.n390 gnd.n324 585
R3427 gnd.n392 gnd.n391 585
R3428 gnd.n388 gnd.n387 585
R3429 gnd.n386 gnd.n329 585
R3430 gnd.n380 gnd.n330 585
R3431 gnd.n382 gnd.n381 585
R3432 gnd.n377 gnd.n332 585
R3433 gnd.n376 gnd.n375 585
R3434 gnd.n369 gnd.n334 585
R3435 gnd.n371 gnd.n370 585
R3436 gnd.n367 gnd.n336 585
R3437 gnd.n366 gnd.n365 585
R3438 gnd.n359 gnd.n338 585
R3439 gnd.n361 gnd.n360 585
R3440 gnd.n357 gnd.n340 585
R3441 gnd.n356 gnd.n355 585
R3442 gnd.n349 gnd.n342 585
R3443 gnd.n351 gnd.n350 585
R3444 gnd.n347 gnd.n346 585
R3445 gnd.n345 gnd.n161 585
R3446 gnd.n165 gnd.n161 585
R3447 gnd.n6837 gnd.n163 585
R3448 gnd.n6841 gnd.n163 585
R3449 gnd.n6836 gnd.n6835 585
R3450 gnd.n6835 gnd.n162 585
R3451 gnd.n6834 gnd.n154 585
R3452 gnd.n6847 gnd.n154 585
R3453 gnd.n6833 gnd.n6832 585
R3454 gnd.n6832 gnd.n147 585
R3455 gnd.n6831 gnd.n145 585
R3456 gnd.n6853 gnd.n145 585
R3457 gnd.n6830 gnd.n6829 585
R3458 gnd.n6829 gnd.n144 585
R3459 gnd.n6827 gnd.n134 585
R3460 gnd.n6859 gnd.n134 585
R3461 gnd.n6826 gnd.n6825 585
R3462 gnd.n6825 gnd.n127 585
R3463 gnd.n6824 gnd.n125 585
R3464 gnd.n6865 gnd.n125 585
R3465 gnd.n6823 gnd.n6822 585
R3466 gnd.n6822 gnd.n124 585
R3467 gnd.n6820 gnd.n115 585
R3468 gnd.n6871 gnd.n115 585
R3469 gnd.n6819 gnd.n6818 585
R3470 gnd.n6818 gnd.n114 585
R3471 gnd.n6817 gnd.n106 585
R3472 gnd.n6877 gnd.n106 585
R3473 gnd.n6816 gnd.n6815 585
R3474 gnd.n6815 gnd.n99 585
R3475 gnd.n6813 gnd.n97 585
R3476 gnd.n6883 gnd.n97 585
R3477 gnd.n6812 gnd.n6811 585
R3478 gnd.n6811 gnd.n88 585
R3479 gnd.n6810 gnd.n86 585
R3480 gnd.n6889 gnd.n86 585
R3481 gnd.n6809 gnd.n6808 585
R3482 gnd.n6808 gnd.n85 585
R3483 gnd.n6807 gnd.n494 585
R3484 gnd.n6807 gnd.n70 585
R3485 gnd.n6796 gnd.n69 585
R3486 gnd.n6897 gnd.n69 585
R3487 gnd.n6798 gnd.n6797 585
R3488 gnd.n6799 gnd.n6798 585
R3489 gnd.n6795 gnd.n500 585
R3490 gnd.n500 gnd.n499 585
R3491 gnd.n505 gnd.n501 585
R3492 gnd.n6790 gnd.n505 585
R3493 gnd.n6760 gnd.n510 585
R3494 gnd.n6782 gnd.n510 585
R3495 gnd.n6762 gnd.n6761 585
R3496 gnd.n6761 gnd.n509 585
R3497 gnd.n6759 gnd.n518 585
R3498 gnd.n6774 gnd.n518 585
R3499 gnd.n6758 gnd.n523 585
R3500 gnd.n6769 gnd.n523 585
R3501 gnd.n6757 gnd.n6756 585
R3502 gnd.n6756 gnd.n6755 585
R3503 gnd.n530 gnd.n528 585
R3504 gnd.n6729 gnd.n530 585
R3505 gnd.n1614 gnd.n537 585
R3506 gnd.n6747 gnd.n537 585
R3507 gnd.n1617 gnd.n1616 585
R3508 gnd.n1616 gnd.n1615 585
R3509 gnd.n1618 gnd.n547 585
R3510 gnd.n6736 gnd.n547 585
R3511 gnd.n1620 gnd.n1619 585
R3512 gnd.n1622 gnd.n1620 585
R3513 gnd.n5501 gnd.n5500 585
R3514 gnd.n5500 gnd.n5499 585
R3515 gnd.n1613 gnd.n1607 585
R3516 gnd.n5506 gnd.n1607 585
R3517 gnd.n5447 gnd.n5446 585
R3518 gnd.n5448 gnd.n5447 585
R3519 gnd.n5444 gnd.n1595 585
R3520 gnd.n5512 gnd.n1595 585
R3521 gnd.n5443 gnd.n5442 585
R3522 gnd.n5442 gnd.n5441 585
R3523 gnd.n5440 gnd.n1582 585
R3524 gnd.n5518 gnd.n1582 585
R3525 gnd.n1566 gnd.n1565 585
R3526 gnd.n5435 gnd.n1566 585
R3527 gnd.n5526 gnd.n5525 585
R3528 gnd.n5525 gnd.n5524 585
R3529 gnd.n5527 gnd.n1555 585
R3530 gnd.n5470 gnd.n1555 585
R3531 gnd.n5533 gnd.n1556 585
R3532 gnd.n5533 gnd.n5532 585
R3533 gnd.n6015 gnd.n6014 585
R3534 gnd.n6014 gnd.n6013 585
R3535 gnd.n6721 gnd.n6719 585
R3536 gnd.n6721 gnd.n6720 585
R3537 gnd.n6724 gnd.n6722 585
R3538 gnd.n6722 gnd.n517 585
R3539 gnd.n6725 gnd.n558 585
R3540 gnd.n558 gnd.n522 585
R3541 gnd.n6727 gnd.n6726 585
R3542 gnd.n6728 gnd.n6727 585
R3543 gnd.n559 gnd.n557 585
R3544 gnd.n557 gnd.n538 585
R3545 gnd.n5492 gnd.n5491 585
R3546 gnd.n5492 gnd.n536 585
R3547 gnd.n5494 gnd.n5493 585
R3548 gnd.n5493 gnd.n549 585
R3549 gnd.n5495 gnd.n1624 585
R3550 gnd.n1624 gnd.n546 585
R3551 gnd.n5497 gnd.n5496 585
R3552 gnd.n5498 gnd.n5497 585
R3553 gnd.n1625 gnd.n1623 585
R3554 gnd.n1623 gnd.n1609 585
R3555 gnd.n5483 gnd.n5482 585
R3556 gnd.n5482 gnd.n1606 585
R3557 gnd.n5481 gnd.n1627 585
R3558 gnd.n5481 gnd.n1597 585
R3559 gnd.n5480 gnd.n5479 585
R3560 gnd.n5480 gnd.n1594 585
R3561 gnd.n1629 gnd.n1628 585
R3562 gnd.n1628 gnd.n1584 585
R3563 gnd.n5475 gnd.n5474 585
R3564 gnd.n5474 gnd.n1581 585
R3565 gnd.n5473 gnd.n1631 585
R3566 gnd.n5473 gnd.n1568 585
R3567 gnd.n5472 gnd.n1633 585
R3568 gnd.n5472 gnd.n5471 585
R3569 gnd.n5417 gnd.n1632 585
R3570 gnd.n1632 gnd.n1559 585
R3571 gnd.n5419 gnd.n5418 585
R3572 gnd.n5419 gnd.n1557 585
R3573 gnd.n5420 gnd.n5412 585
R3574 gnd.n5420 gnd.n1489 585
R3575 gnd.n5422 gnd.n5421 585
R3576 gnd.n5421 gnd.n1447 585
R3577 gnd.n5423 gnd.n1664 585
R3578 gnd.n1664 gnd.n1662 585
R3579 gnd.n5425 gnd.n5424 585
R3580 gnd.n5426 gnd.n5425 585
R3581 gnd.n1665 gnd.n1663 585
R3582 gnd.n1663 gnd.n1380 585
R3583 gnd.n5406 gnd.n1379 585
R3584 gnd.n5721 gnd.n1379 585
R3585 gnd.n5405 gnd.n5404 585
R3586 gnd.n5404 gnd.n1378 585
R3587 gnd.n5403 gnd.n1667 585
R3588 gnd.n5403 gnd.n5402 585
R3589 gnd.n5391 gnd.n1668 585
R3590 gnd.n1669 gnd.n1668 585
R3591 gnd.n5393 gnd.n5392 585
R3592 gnd.n5394 gnd.n5393 585
R3593 gnd.n1678 gnd.n1677 585
R3594 gnd.n1677 gnd.n1676 585
R3595 gnd.n5385 gnd.n5384 585
R3596 gnd.n5384 gnd.n5383 585
R3597 gnd.n1681 gnd.n1680 585
R3598 gnd.n1689 gnd.n1681 585
R3599 gnd.n5374 gnd.n5373 585
R3600 gnd.n5375 gnd.n5374 585
R3601 gnd.n1691 gnd.n1690 585
R3602 gnd.n1690 gnd.n1688 585
R3603 gnd.n5369 gnd.n5368 585
R3604 gnd.n5368 gnd.n5367 585
R3605 gnd.n1694 gnd.n1693 585
R3606 gnd.n1701 gnd.n1694 585
R3607 gnd.n5358 gnd.n5357 585
R3608 gnd.n5359 gnd.n5358 585
R3609 gnd.n1704 gnd.n1703 585
R3610 gnd.n1712 gnd.n1703 585
R3611 gnd.n5353 gnd.n5352 585
R3612 gnd.n5352 gnd.n5351 585
R3613 gnd.n1707 gnd.n1706 585
R3614 gnd.n1787 gnd.n1707 585
R3615 gnd.n5211 gnd.n5210 585
R3616 gnd.n5212 gnd.n5211 585
R3617 gnd.n1795 gnd.n1794 585
R3618 gnd.n1802 gnd.n1794 585
R3619 gnd.n5206 gnd.n5205 585
R3620 gnd.n5205 gnd.n5204 585
R3621 gnd.n1798 gnd.n1797 585
R3622 gnd.n1806 gnd.n1798 585
R3623 gnd.n5182 gnd.n5181 585
R3624 gnd.n5183 gnd.n5182 585
R3625 gnd.n1812 gnd.n1811 585
R3626 gnd.n1820 gnd.n1811 585
R3627 gnd.n5177 gnd.n5176 585
R3628 gnd.n5176 gnd.n5175 585
R3629 gnd.n1815 gnd.n1814 585
R3630 gnd.n1826 gnd.n1815 585
R3631 gnd.n5152 gnd.n5151 585
R3632 gnd.n5153 gnd.n5152 585
R3633 gnd.n1834 gnd.n1833 585
R3634 gnd.n5103 gnd.n1833 585
R3635 gnd.n5147 gnd.n5146 585
R3636 gnd.n5146 gnd.n5145 585
R3637 gnd.n1837 gnd.n1836 585
R3638 gnd.n5137 gnd.n1837 585
R3639 gnd.n5093 gnd.n1856 585
R3640 gnd.n5077 gnd.n1856 585
R3641 gnd.n5095 gnd.n5094 585
R3642 gnd.n5096 gnd.n5095 585
R3643 gnd.n1857 gnd.n1855 585
R3644 gnd.n1864 gnd.n1855 585
R3645 gnd.n5088 gnd.n5087 585
R3646 gnd.n5087 gnd.n5086 585
R3647 gnd.n1860 gnd.n1859 585
R3648 gnd.n1873 gnd.n1860 585
R3649 gnd.n5049 gnd.n5048 585
R3650 gnd.n5050 gnd.n5049 585
R3651 gnd.n1883 gnd.n1882 585
R3652 gnd.n4975 gnd.n1882 585
R3653 gnd.n5044 gnd.n5043 585
R3654 gnd.n5043 gnd.n5042 585
R3655 gnd.n1886 gnd.n1885 585
R3656 gnd.n1893 gnd.n1886 585
R3657 gnd.n5013 gnd.n1908 585
R3658 gnd.n1908 gnd.n1901 585
R3659 gnd.n5015 gnd.n5014 585
R3660 gnd.n5016 gnd.n5015 585
R3661 gnd.n1909 gnd.n1907 585
R3662 gnd.n4969 gnd.n1907 585
R3663 gnd.n5008 gnd.n5007 585
R3664 gnd.n5007 gnd.n5006 585
R3665 gnd.n1912 gnd.n1911 585
R3666 gnd.n4998 gnd.n1912 585
R3667 gnd.n4960 gnd.n1930 585
R3668 gnd.n1930 gnd.n1920 585
R3669 gnd.n4962 gnd.n4961 585
R3670 gnd.n4963 gnd.n4962 585
R3671 gnd.n1931 gnd.n1929 585
R3672 gnd.n1943 gnd.n1929 585
R3673 gnd.n4955 gnd.n4954 585
R3674 gnd.n4954 gnd.n4953 585
R3675 gnd.n1934 gnd.n1933 585
R3676 gnd.n4926 gnd.n1934 585
R3677 gnd.n4914 gnd.n1957 585
R3678 gnd.n4898 gnd.n1957 585
R3679 gnd.n4916 gnd.n4915 585
R3680 gnd.n4917 gnd.n4916 585
R3681 gnd.n1958 gnd.n1956 585
R3682 gnd.n4889 gnd.n1956 585
R3683 gnd.n4909 gnd.n4908 585
R3684 gnd.n4908 gnd.n4907 585
R3685 gnd.n1961 gnd.n1960 585
R3686 gnd.n1976 gnd.n1961 585
R3687 gnd.n4874 gnd.n4873 585
R3688 gnd.n4875 gnd.n4874 585
R3689 gnd.n1984 gnd.n1983 585
R3690 gnd.n4852 gnd.n1983 585
R3691 gnd.n4869 gnd.n4868 585
R3692 gnd.n4868 gnd.n4867 585
R3693 gnd.n1987 gnd.n1986 585
R3694 gnd.n1994 gnd.n1987 585
R3695 gnd.n4835 gnd.n4834 585
R3696 gnd.n4836 gnd.n4835 585
R3697 gnd.n2008 gnd.n2007 585
R3698 gnd.n4765 gnd.n2007 585
R3699 gnd.n4830 gnd.n4829 585
R3700 gnd.n4829 gnd.n4828 585
R3701 gnd.n2011 gnd.n2010 585
R3702 gnd.n4817 gnd.n2011 585
R3703 gnd.n4803 gnd.n2030 585
R3704 gnd.n4759 gnd.n2030 585
R3705 gnd.n4805 gnd.n4804 585
R3706 gnd.n4806 gnd.n4805 585
R3707 gnd.n2031 gnd.n2029 585
R3708 gnd.n2039 gnd.n2029 585
R3709 gnd.n4798 gnd.n4797 585
R3710 gnd.n4797 gnd.n4796 585
R3711 gnd.n2035 gnd.n2034 585
R3712 gnd.n2044 gnd.n2035 585
R3713 gnd.n1288 gnd.n1287 585
R3714 gnd.n2051 gnd.n1288 585
R3715 gnd.n5827 gnd.n5826 585
R3716 gnd.n5826 gnd.n5825 585
R3717 gnd.n5828 gnd.n1282 585
R3718 gnd.n4671 gnd.n1282 585
R3719 gnd.n5830 gnd.n5829 585
R3720 gnd.n5831 gnd.n5830 585
R3721 gnd.n1283 gnd.n1281 585
R3722 gnd.n1281 gnd.n1276 585
R3723 gnd.n4640 gnd.n4639 585
R3724 gnd.n4640 gnd.n1250 585
R3725 gnd.n4642 gnd.n4641 585
R3726 gnd.n4641 gnd.n1218 585
R3727 gnd.n4643 gnd.n2068 585
R3728 gnd.n2068 gnd.n2065 585
R3729 gnd.n4645 gnd.n4644 585
R3730 gnd.n4646 gnd.n4645 585
R3731 gnd.n2069 gnd.n2067 585
R3732 gnd.n2067 gnd.n2064 585
R3733 gnd.n4631 gnd.n4630 585
R3734 gnd.n4630 gnd.n4629 585
R3735 gnd.n2072 gnd.n2071 585
R3736 gnd.n2083 gnd.n2072 585
R3737 gnd.n4603 gnd.n4602 585
R3738 gnd.n4604 gnd.n4603 585
R3739 gnd.n2085 gnd.n2084 585
R3740 gnd.n2084 gnd.n2081 585
R3741 gnd.n4598 gnd.n4597 585
R3742 gnd.n4597 gnd.n4596 585
R3743 gnd.n2088 gnd.n2087 585
R3744 gnd.n2089 gnd.n2088 585
R3745 gnd.n4587 gnd.n4586 585
R3746 gnd.n4588 gnd.n4587 585
R3747 gnd.n2099 gnd.n2098 585
R3748 gnd.n2098 gnd.n2096 585
R3749 gnd.n4582 gnd.n4581 585
R3750 gnd.n4581 gnd.n4580 585
R3751 gnd.n2102 gnd.n2101 585
R3752 gnd.n4579 gnd.n2102 585
R3753 gnd.n4562 gnd.n4561 585
R3754 gnd.n4562 gnd.n2103 585
R3755 gnd.n4564 gnd.n4563 585
R3756 gnd.n4563 gnd.n1155 585
R3757 gnd.n4565 gnd.n2128 585
R3758 gnd.n2128 gnd.n1144 585
R3759 gnd.n4567 gnd.n4566 585
R3760 gnd.n4568 gnd.n4567 585
R3761 gnd.n2129 gnd.n2127 585
R3762 gnd.n2127 gnd.n1137 585
R3763 gnd.n4554 gnd.n4553 585
R3764 gnd.n4553 gnd.n1134 585
R3765 gnd.n4552 gnd.n2131 585
R3766 gnd.n4552 gnd.n1127 585
R3767 gnd.n4551 gnd.n4550 585
R3768 gnd.n4551 gnd.n1124 585
R3769 gnd.n2133 gnd.n2132 585
R3770 gnd.n2132 gnd.n1116 585
R3771 gnd.n4546 gnd.n4545 585
R3772 gnd.n4545 gnd.n1113 585
R3773 gnd.n4544 gnd.n2135 585
R3774 gnd.n4544 gnd.n4543 585
R3775 gnd.n4247 gnd.n2136 585
R3776 gnd.n2136 gnd.n1104 585
R3777 gnd.n4248 gnd.n2150 585
R3778 gnd.n2150 gnd.n1096 585
R3779 gnd.n4250 gnd.n4249 585
R3780 gnd.n4251 gnd.n4250 585
R3781 gnd.n2151 gnd.n2149 585
R3782 gnd.n2149 gnd.n1087 585
R3783 gnd.n4241 gnd.n4240 585
R3784 gnd.n4240 gnd.n1084 585
R3785 gnd.n4239 gnd.n2153 585
R3786 gnd.n4239 gnd.n1076 585
R3787 gnd.n4238 gnd.n4237 585
R3788 gnd.n4238 gnd.n1073 585
R3789 gnd.n4228 gnd.n4227 585
R3790 gnd.n4227 gnd.n4226 585
R3791 gnd.n4233 gnd.n4232 585
R3792 gnd.n4232 gnd.n1062 585
R3793 gnd.n4231 gnd.n1049 585
R3794 gnd.n1053 gnd.n1049 585
R3795 gnd.n5720 gnd.n5719 585
R3796 gnd.n5721 gnd.n5720 585
R3797 gnd.n1383 gnd.n1381 585
R3798 gnd.n1381 gnd.n1378 585
R3799 gnd.n5401 gnd.n5400 585
R3800 gnd.n5402 gnd.n5401 585
R3801 gnd.n1671 gnd.n1670 585
R3802 gnd.n1670 gnd.n1669 585
R3803 gnd.n5396 gnd.n5395 585
R3804 gnd.n5395 gnd.n5394 585
R3805 gnd.n1674 gnd.n1673 585
R3806 gnd.n1676 gnd.n1674 585
R3807 gnd.n5382 gnd.n5381 585
R3808 gnd.n5383 gnd.n5382 585
R3809 gnd.n1683 gnd.n1682 585
R3810 gnd.n1689 gnd.n1682 585
R3811 gnd.n5377 gnd.n5376 585
R3812 gnd.n5376 gnd.n5375 585
R3813 gnd.n1686 gnd.n1685 585
R3814 gnd.n1688 gnd.n1686 585
R3815 gnd.n5366 gnd.n5365 585
R3816 gnd.n5367 gnd.n5366 585
R3817 gnd.n1696 gnd.n1695 585
R3818 gnd.n1701 gnd.n1695 585
R3819 gnd.n5361 gnd.n5360 585
R3820 gnd.n5360 gnd.n5359 585
R3821 gnd.n1699 gnd.n1698 585
R3822 gnd.n1712 gnd.n1699 585
R3823 gnd.n5114 gnd.n1709 585
R3824 gnd.n5351 gnd.n1709 585
R3825 gnd.n5117 gnd.n5113 585
R3826 gnd.n5113 gnd.n1787 585
R3827 gnd.n5118 gnd.n1792 585
R3828 gnd.n5212 gnd.n1792 585
R3829 gnd.n5119 gnd.n5112 585
R3830 gnd.n5112 gnd.n1802 585
R3831 gnd.n5110 gnd.n1799 585
R3832 gnd.n5204 gnd.n1799 585
R3833 gnd.n5123 gnd.n5109 585
R3834 gnd.n5109 gnd.n1806 585
R3835 gnd.n5124 gnd.n1810 585
R3836 gnd.n5183 gnd.n1810 585
R3837 gnd.n5125 gnd.n5108 585
R3838 gnd.n5108 gnd.n1820 585
R3839 gnd.n5106 gnd.n1817 585
R3840 gnd.n5175 gnd.n1817 585
R3841 gnd.n5129 gnd.n5105 585
R3842 gnd.n5105 gnd.n1826 585
R3843 gnd.n5130 gnd.n1831 585
R3844 gnd.n5153 gnd.n1831 585
R3845 gnd.n5131 gnd.n5104 585
R3846 gnd.n5104 gnd.n5103 585
R3847 gnd.n1849 gnd.n1839 585
R3848 gnd.n5145 gnd.n1839 585
R3849 gnd.n5136 gnd.n5135 585
R3850 gnd.n5137 gnd.n5136 585
R3851 gnd.n1848 gnd.n1847 585
R3852 gnd.n5077 gnd.n1847 585
R3853 gnd.n5098 gnd.n5097 585
R3854 gnd.n5097 gnd.n5096 585
R3855 gnd.n1852 gnd.n1851 585
R3856 gnd.n1864 gnd.n1852 585
R3857 gnd.n4979 gnd.n1862 585
R3858 gnd.n5086 gnd.n1862 585
R3859 gnd.n4978 gnd.n4977 585
R3860 gnd.n4977 gnd.n1873 585
R3861 gnd.n4983 gnd.n1879 585
R3862 gnd.n5050 gnd.n1879 585
R3863 gnd.n4984 gnd.n4976 585
R3864 gnd.n4976 gnd.n4975 585
R3865 gnd.n4985 gnd.n1888 585
R3866 gnd.n5042 gnd.n1888 585
R3867 gnd.n4973 gnd.n4972 585
R3868 gnd.n4972 gnd.n1893 585
R3869 gnd.n4989 gnd.n4971 585
R3870 gnd.n4971 gnd.n1901 585
R3871 gnd.n4990 gnd.n1906 585
R3872 gnd.n5016 gnd.n1906 585
R3873 gnd.n4991 gnd.n4970 585
R3874 gnd.n4970 gnd.n4969 585
R3875 gnd.n1924 gnd.n1914 585
R3876 gnd.n5006 gnd.n1914 585
R3877 gnd.n4996 gnd.n4995 585
R3878 gnd.n4998 gnd.n4996 585
R3879 gnd.n1923 gnd.n1922 585
R3880 gnd.n1922 gnd.n1920 585
R3881 gnd.n4965 gnd.n4964 585
R3882 gnd.n4964 gnd.n4963 585
R3883 gnd.n1927 gnd.n1926 585
R3884 gnd.n1943 gnd.n1927 585
R3885 gnd.n1951 gnd.n1935 585
R3886 gnd.n4953 gnd.n1935 585
R3887 gnd.n4925 gnd.n4924 585
R3888 gnd.n4926 gnd.n4925 585
R3889 gnd.n1950 gnd.n1949 585
R3890 gnd.n4898 gnd.n1949 585
R3891 gnd.n4919 gnd.n4918 585
R3892 gnd.n4918 gnd.n4917 585
R3893 gnd.n1954 gnd.n1953 585
R3894 gnd.n4889 gnd.n1954 585
R3895 gnd.n4844 gnd.n1963 585
R3896 gnd.n4907 gnd.n1963 585
R3897 gnd.n4845 gnd.n4843 585
R3898 gnd.n4843 gnd.n1976 585
R3899 gnd.n2001 gnd.n1981 585
R3900 gnd.n4875 gnd.n1981 585
R3901 gnd.n4850 gnd.n4849 585
R3902 gnd.n4852 gnd.n4850 585
R3903 gnd.n2000 gnd.n1989 585
R3904 gnd.n4867 gnd.n1989 585
R3905 gnd.n4839 gnd.n4838 585
R3906 gnd.n4838 gnd.n1994 585
R3907 gnd.n4837 gnd.n2003 585
R3908 gnd.n4837 gnd.n4836 585
R3909 gnd.n4811 gnd.n2004 585
R3910 gnd.n4765 gnd.n2004 585
R3911 gnd.n2022 gnd.n2013 585
R3912 gnd.n4828 gnd.n2013 585
R3913 gnd.n4816 gnd.n4815 585
R3914 gnd.n4817 gnd.n4816 585
R3915 gnd.n2021 gnd.n2020 585
R3916 gnd.n4759 gnd.n2020 585
R3917 gnd.n4808 gnd.n4807 585
R3918 gnd.n4807 gnd.n4806 585
R3919 gnd.n2025 gnd.n2024 585
R3920 gnd.n2039 gnd.n2025 585
R3921 gnd.n4663 gnd.n2037 585
R3922 gnd.n4796 gnd.n2037 585
R3923 gnd.n4664 gnd.n4661 585
R3924 gnd.n4661 gnd.n2044 585
R3925 gnd.n4665 gnd.n4660 585
R3926 gnd.n4660 gnd.n2051 585
R3927 gnd.n2056 gnd.n1289 585
R3928 gnd.n5825 gnd.n1289 585
R3929 gnd.n4670 gnd.n4669 585
R3930 gnd.n4671 gnd.n4670 585
R3931 gnd.n2055 gnd.n1278 585
R3932 gnd.n5831 gnd.n1278 585
R3933 gnd.n4656 gnd.n4655 585
R3934 gnd.n4655 gnd.n1276 585
R3935 gnd.n4654 gnd.n2058 585
R3936 gnd.n4654 gnd.n1250 585
R3937 gnd.n4653 gnd.n4652 585
R3938 gnd.n4653 gnd.n1218 585
R3939 gnd.n2060 gnd.n2059 585
R3940 gnd.n2065 gnd.n2059 585
R3941 gnd.n4648 gnd.n4647 585
R3942 gnd.n4647 gnd.n4646 585
R3943 gnd.n2063 gnd.n2062 585
R3944 gnd.n2064 gnd.n2063 585
R3945 gnd.n4285 gnd.n2073 585
R3946 gnd.n4629 gnd.n2073 585
R3947 gnd.n4286 gnd.n4284 585
R3948 gnd.n4284 gnd.n2083 585
R3949 gnd.n4282 gnd.n2082 585
R3950 gnd.n4604 gnd.n2082 585
R3951 gnd.n4290 gnd.n4281 585
R3952 gnd.n4281 gnd.n2081 585
R3953 gnd.n4291 gnd.n2090 585
R3954 gnd.n4596 gnd.n2090 585
R3955 gnd.n4292 gnd.n4280 585
R3956 gnd.n4280 gnd.n2089 585
R3957 gnd.n4278 gnd.n2097 585
R3958 gnd.n4588 gnd.n2097 585
R3959 gnd.n4297 gnd.n4296 585
R3960 gnd.n4297 gnd.n2096 585
R3961 gnd.n4299 gnd.n4298 585
R3962 gnd.n4301 gnd.n4300 585
R3963 gnd.n4303 gnd.n4302 585
R3964 gnd.n4274 gnd.n4273 585
R3965 gnd.n4307 gnd.n4275 585
R3966 gnd.n4309 gnd.n4308 585
R3967 gnd.n4424 gnd.n4310 585
R3968 gnd.n4423 gnd.n4311 585
R3969 gnd.n4422 gnd.n4312 585
R3970 gnd.n4318 gnd.n4313 585
R3971 gnd.n4415 gnd.n4319 585
R3972 gnd.n4414 gnd.n4320 585
R3973 gnd.n4322 gnd.n4321 585
R3974 gnd.n4407 gnd.n4330 585
R3975 gnd.n4406 gnd.n4331 585
R3976 gnd.n4338 gnd.n4332 585
R3977 gnd.n4399 gnd.n4339 585
R3978 gnd.n4398 gnd.n4340 585
R3979 gnd.n4342 gnd.n4341 585
R3980 gnd.n4391 gnd.n4350 585
R3981 gnd.n4390 gnd.n4351 585
R3982 gnd.n4358 gnd.n4352 585
R3983 gnd.n4383 gnd.n4359 585
R3984 gnd.n4382 gnd.n4360 585
R3985 gnd.n4362 gnd.n4361 585
R3986 gnd.n4375 gnd.n4372 585
R3987 gnd.n4374 gnd.n4373 585
R3988 gnd.n2119 gnd.n2118 585
R3989 gnd.n4578 gnd.n4577 585
R3990 gnd.n4579 gnd.n4578 585
R3991 gnd.n5723 gnd.n5722 585
R3992 gnd.n5722 gnd.n5721 585
R3993 gnd.n1376 gnd.n1374 585
R3994 gnd.n1378 gnd.n1376 585
R3995 gnd.n5727 gnd.n1373 585
R3996 gnd.n5402 gnd.n1373 585
R3997 gnd.n5728 gnd.n1372 585
R3998 gnd.n1669 gnd.n1372 585
R3999 gnd.n5729 gnd.n1371 585
R4000 gnd.n5394 gnd.n1371 585
R4001 gnd.n1675 gnd.n1369 585
R4002 gnd.n1676 gnd.n1675 585
R4003 gnd.n5733 gnd.n1368 585
R4004 gnd.n5383 gnd.n1368 585
R4005 gnd.n5734 gnd.n1367 585
R4006 gnd.n1689 gnd.n1367 585
R4007 gnd.n5735 gnd.n1366 585
R4008 gnd.n5375 gnd.n1366 585
R4009 gnd.n1687 gnd.n1364 585
R4010 gnd.n1688 gnd.n1687 585
R4011 gnd.n5739 gnd.n1363 585
R4012 gnd.n5367 gnd.n1363 585
R4013 gnd.n5740 gnd.n1362 585
R4014 gnd.n1701 gnd.n1362 585
R4015 gnd.n5741 gnd.n1361 585
R4016 gnd.n5359 gnd.n1361 585
R4017 gnd.n1711 gnd.n1359 585
R4018 gnd.n1712 gnd.n1711 585
R4019 gnd.n5745 gnd.n1358 585
R4020 gnd.n5351 gnd.n1358 585
R4021 gnd.n5746 gnd.n1357 585
R4022 gnd.n1787 gnd.n1357 585
R4023 gnd.n5747 gnd.n1356 585
R4024 gnd.n5212 gnd.n1356 585
R4025 gnd.n1801 gnd.n1354 585
R4026 gnd.n1802 gnd.n1801 585
R4027 gnd.n5751 gnd.n1353 585
R4028 gnd.n5204 gnd.n1353 585
R4029 gnd.n5752 gnd.n1352 585
R4030 gnd.n1806 gnd.n1352 585
R4031 gnd.n5753 gnd.n1351 585
R4032 gnd.n5183 gnd.n1351 585
R4033 gnd.n1819 gnd.n1349 585
R4034 gnd.n1820 gnd.n1819 585
R4035 gnd.n5757 gnd.n1348 585
R4036 gnd.n5175 gnd.n1348 585
R4037 gnd.n5758 gnd.n1347 585
R4038 gnd.n1826 gnd.n1347 585
R4039 gnd.n5759 gnd.n1346 585
R4040 gnd.n5153 gnd.n1346 585
R4041 gnd.n5102 gnd.n1344 585
R4042 gnd.n5103 gnd.n5102 585
R4043 gnd.n5763 gnd.n1343 585
R4044 gnd.n5145 gnd.n1343 585
R4045 gnd.n5764 gnd.n1342 585
R4046 gnd.n5137 gnd.n1342 585
R4047 gnd.n5765 gnd.n1341 585
R4048 gnd.n5077 gnd.n1341 585
R4049 gnd.n1854 gnd.n1339 585
R4050 gnd.n5096 gnd.n1854 585
R4051 gnd.n5769 gnd.n1338 585
R4052 gnd.n1864 gnd.n1338 585
R4053 gnd.n5770 gnd.n1337 585
R4054 gnd.n5086 gnd.n1337 585
R4055 gnd.n5771 gnd.n1336 585
R4056 gnd.n1873 gnd.n1336 585
R4057 gnd.n1881 gnd.n1334 585
R4058 gnd.n5050 gnd.n1881 585
R4059 gnd.n5775 gnd.n1333 585
R4060 gnd.n4975 gnd.n1333 585
R4061 gnd.n5776 gnd.n1332 585
R4062 gnd.n5042 gnd.n1332 585
R4063 gnd.n5777 gnd.n1331 585
R4064 gnd.n1893 gnd.n1331 585
R4065 gnd.n1900 gnd.n1329 585
R4066 gnd.n1901 gnd.n1900 585
R4067 gnd.n5781 gnd.n1328 585
R4068 gnd.n5016 gnd.n1328 585
R4069 gnd.n5782 gnd.n1327 585
R4070 gnd.n4969 gnd.n1327 585
R4071 gnd.n5783 gnd.n1326 585
R4072 gnd.n5006 gnd.n1326 585
R4073 gnd.n4997 gnd.n1324 585
R4074 gnd.n4998 gnd.n4997 585
R4075 gnd.n5787 gnd.n1323 585
R4076 gnd.n1920 gnd.n1323 585
R4077 gnd.n5788 gnd.n1322 585
R4078 gnd.n4963 gnd.n1322 585
R4079 gnd.n5789 gnd.n1321 585
R4080 gnd.n1943 gnd.n1321 585
R4081 gnd.n4952 gnd.n1319 585
R4082 gnd.n4953 gnd.n4952 585
R4083 gnd.n5793 gnd.n1318 585
R4084 gnd.n4926 gnd.n1318 585
R4085 gnd.n5794 gnd.n1317 585
R4086 gnd.n4898 gnd.n1317 585
R4087 gnd.n5795 gnd.n1316 585
R4088 gnd.n4917 gnd.n1316 585
R4089 gnd.n4888 gnd.n1314 585
R4090 gnd.n4889 gnd.n4888 585
R4091 gnd.n5799 gnd.n1313 585
R4092 gnd.n4907 gnd.n1313 585
R4093 gnd.n5800 gnd.n1312 585
R4094 gnd.n1976 gnd.n1312 585
R4095 gnd.n5801 gnd.n1311 585
R4096 gnd.n4875 gnd.n1311 585
R4097 gnd.n4851 gnd.n1309 585
R4098 gnd.n4852 gnd.n4851 585
R4099 gnd.n5805 gnd.n1308 585
R4100 gnd.n4867 gnd.n1308 585
R4101 gnd.n5806 gnd.n1307 585
R4102 gnd.n1994 gnd.n1307 585
R4103 gnd.n5807 gnd.n1306 585
R4104 gnd.n4836 gnd.n1306 585
R4105 gnd.n4764 gnd.n1304 585
R4106 gnd.n4765 gnd.n4764 585
R4107 gnd.n5811 gnd.n1303 585
R4108 gnd.n4828 gnd.n1303 585
R4109 gnd.n5812 gnd.n1302 585
R4110 gnd.n4817 gnd.n1302 585
R4111 gnd.n5813 gnd.n1301 585
R4112 gnd.n4759 gnd.n1301 585
R4113 gnd.n2028 gnd.n1299 585
R4114 gnd.n4806 gnd.n2028 585
R4115 gnd.n5817 gnd.n1298 585
R4116 gnd.n2039 gnd.n1298 585
R4117 gnd.n5818 gnd.n1297 585
R4118 gnd.n4796 gnd.n1297 585
R4119 gnd.n5819 gnd.n1296 585
R4120 gnd.n2044 gnd.n1296 585
R4121 gnd.n1293 gnd.n1291 585
R4122 gnd.n2051 gnd.n1291 585
R4123 gnd.n5824 gnd.n5823 585
R4124 gnd.n5825 gnd.n5824 585
R4125 gnd.n1292 gnd.n1290 585
R4126 gnd.n4671 gnd.n1290 585
R4127 gnd.n4616 gnd.n1280 585
R4128 gnd.n5831 gnd.n1280 585
R4129 gnd.n4617 gnd.n4615 585
R4130 gnd.n4615 gnd.n1276 585
R4131 gnd.n4614 gnd.n4612 585
R4132 gnd.n4614 gnd.n1250 585
R4133 gnd.n4621 gnd.n4611 585
R4134 gnd.n4611 gnd.n1218 585
R4135 gnd.n4622 gnd.n4610 585
R4136 gnd.n4610 gnd.n2065 585
R4137 gnd.n4623 gnd.n2066 585
R4138 gnd.n4646 gnd.n2066 585
R4139 gnd.n2077 gnd.n2075 585
R4140 gnd.n2075 gnd.n2064 585
R4141 gnd.n4628 gnd.n4627 585
R4142 gnd.n4629 gnd.n4628 585
R4143 gnd.n2076 gnd.n2074 585
R4144 gnd.n2083 gnd.n2074 585
R4145 gnd.n4606 gnd.n4605 585
R4146 gnd.n4605 gnd.n4604 585
R4147 gnd.n2080 gnd.n2079 585
R4148 gnd.n2081 gnd.n2080 585
R4149 gnd.n4595 gnd.n4594 585
R4150 gnd.n4596 gnd.n4595 585
R4151 gnd.n2092 gnd.n2091 585
R4152 gnd.n2091 gnd.n2089 585
R4153 gnd.n4590 gnd.n4589 585
R4154 gnd.n4589 gnd.n4588 585
R4155 gnd.n2095 gnd.n2094 585
R4156 gnd.n2096 gnd.n2095 585
R4157 gnd.n5662 gnd.n1438 585
R4158 gnd.n5663 gnd.n1437 585
R4159 gnd.n1657 gnd.n1431 585
R4160 gnd.n5670 gnd.n1430 585
R4161 gnd.n5671 gnd.n1429 585
R4162 gnd.n1654 gnd.n1423 585
R4163 gnd.n5678 gnd.n1422 585
R4164 gnd.n5679 gnd.n1421 585
R4165 gnd.n1652 gnd.n1415 585
R4166 gnd.n5686 gnd.n1414 585
R4167 gnd.n5687 gnd.n1413 585
R4168 gnd.n1649 gnd.n1407 585
R4169 gnd.n5694 gnd.n1406 585
R4170 gnd.n5695 gnd.n1405 585
R4171 gnd.n1647 gnd.n1398 585
R4172 gnd.n5702 gnd.n1397 585
R4173 gnd.n5703 gnd.n1396 585
R4174 gnd.n1644 gnd.n1393 585
R4175 gnd.n5708 gnd.n1392 585
R4176 gnd.n5709 gnd.n1391 585
R4177 gnd.n5710 gnd.n1390 585
R4178 gnd.n1641 gnd.n1388 585
R4179 gnd.n5714 gnd.n1387 585
R4180 gnd.n5715 gnd.n1386 585
R4181 gnd.n5716 gnd.n1382 585
R4182 gnd.n5429 gnd.n1377 585
R4183 gnd.n5426 gnd.n1377 585
R4184 gnd.n5430 gnd.n5428 585
R4185 gnd.n1639 gnd.n1638 585
R4186 gnd.n1660 gnd.n1659 585
R4187 gnd.n5344 gnd.n1714 473.281
R4188 gnd.n5227 gnd.n5226 473.281
R4189 gnd.n4740 gnd.n4738 473.281
R4190 gnd.n5900 gnd.n1253 473.281
R4191 gnd.n4674 gnd.t298 443.966
R4192 gnd.n1762 gnd.t232 443.966
R4193 gnd.n5837 gnd.t222 443.966
R4194 gnd.n1756 gnd.t285 443.966
R4195 gnd.n6181 gnd.n878 371.755
R4196 gnd.n4369 gnd.t269 371.625
R4197 gnd.n5656 gnd.t291 371.625
R4198 gnd.n2122 gnd.t314 371.625
R4199 gnd.n1511 gnd.t288 371.625
R4200 gnd.n1534 gnd.t279 371.625
R4201 gnd.n5536 gnd.t218 371.625
R4202 gnd.n282 gnd.t226 371.625
R4203 gnd.n304 gnd.t214 371.625
R4204 gnd.n326 gnd.t282 371.625
R4205 gnd.n200 gnd.t304 371.625
R4206 gnd.n3793 gnd.t256 371.625
R4207 gnd.n3815 gnd.t236 371.625
R4208 gnd.n3836 gnd.t259 371.625
R4209 gnd.n3854 gnd.t207 371.625
R4210 gnd.n1201 gnd.t307 371.625
R4211 gnd.n4428 gnd.t239 371.625
R4212 gnd.n4441 gnd.t266 371.625
R4213 gnd.n1439 gnd.t243 371.625
R4214 gnd.n2754 gnd.t262 323.425
R4215 gnd.n2312 gnd.t294 323.425
R4216 gnd.n3603 gnd.n3577 289.615
R4217 gnd.n3571 gnd.n3545 289.615
R4218 gnd.n3539 gnd.n3513 289.615
R4219 gnd.n3508 gnd.n3482 289.615
R4220 gnd.n3476 gnd.n3450 289.615
R4221 gnd.n3444 gnd.n3418 289.615
R4222 gnd.n3412 gnd.n3386 289.615
R4223 gnd.n3381 gnd.n3355 289.615
R4224 gnd.n2828 gnd.t317 279.217
R4225 gnd.n2338 gnd.t310 279.217
R4226 gnd.n1260 gnd.t213 260.649
R4227 gnd.n1727 gnd.t252 260.649
R4228 gnd.n5902 gnd.n5901 256.663
R4229 gnd.n5902 gnd.n1219 256.663
R4230 gnd.n5902 gnd.n1220 256.663
R4231 gnd.n5902 gnd.n1221 256.663
R4232 gnd.n5902 gnd.n1222 256.663
R4233 gnd.n5902 gnd.n1223 256.663
R4234 gnd.n5902 gnd.n1224 256.663
R4235 gnd.n5902 gnd.n1225 256.663
R4236 gnd.n5902 gnd.n1226 256.663
R4237 gnd.n5902 gnd.n1227 256.663
R4238 gnd.n5902 gnd.n1228 256.663
R4239 gnd.n5902 gnd.n1229 256.663
R4240 gnd.n5902 gnd.n1230 256.663
R4241 gnd.n5902 gnd.n1231 256.663
R4242 gnd.n5902 gnd.n1232 256.663
R4243 gnd.n5902 gnd.n1233 256.663
R4244 gnd.n5905 gnd.n1216 256.663
R4245 gnd.n5903 gnd.n5902 256.663
R4246 gnd.n5902 gnd.n1234 256.663
R4247 gnd.n5902 gnd.n1235 256.663
R4248 gnd.n5902 gnd.n1236 256.663
R4249 gnd.n5902 gnd.n1237 256.663
R4250 gnd.n5902 gnd.n1238 256.663
R4251 gnd.n5902 gnd.n1239 256.663
R4252 gnd.n5902 gnd.n1240 256.663
R4253 gnd.n5902 gnd.n1241 256.663
R4254 gnd.n5902 gnd.n1242 256.663
R4255 gnd.n5902 gnd.n1243 256.663
R4256 gnd.n5902 gnd.n1244 256.663
R4257 gnd.n5902 gnd.n1245 256.663
R4258 gnd.n5902 gnd.n1246 256.663
R4259 gnd.n5902 gnd.n1247 256.663
R4260 gnd.n5902 gnd.n1248 256.663
R4261 gnd.n5902 gnd.n1249 256.663
R4262 gnd.n5225 gnd.n1702 256.663
R4263 gnd.n5232 gnd.n1702 256.663
R4264 gnd.n1783 gnd.n1702 256.663
R4265 gnd.n5239 gnd.n1702 256.663
R4266 gnd.n1780 gnd.n1702 256.663
R4267 gnd.n5246 gnd.n1702 256.663
R4268 gnd.n1777 gnd.n1702 256.663
R4269 gnd.n5253 gnd.n1702 256.663
R4270 gnd.n1774 gnd.n1702 256.663
R4271 gnd.n5260 gnd.n1702 256.663
R4272 gnd.n1771 gnd.n1702 256.663
R4273 gnd.n5267 gnd.n1702 256.663
R4274 gnd.n1768 gnd.n1702 256.663
R4275 gnd.n5274 gnd.n1702 256.663
R4276 gnd.n1765 gnd.n1702 256.663
R4277 gnd.n5282 gnd.n1702 256.663
R4278 gnd.n5285 gnd.n1521 256.663
R4279 gnd.n5286 gnd.n1702 256.663
R4280 gnd.n5290 gnd.n1702 256.663
R4281 gnd.n1759 gnd.n1702 256.663
R4282 gnd.n5298 gnd.n1702 256.663
R4283 gnd.n1754 gnd.n1702 256.663
R4284 gnd.n5305 gnd.n1702 256.663
R4285 gnd.n1751 gnd.n1702 256.663
R4286 gnd.n5312 gnd.n1702 256.663
R4287 gnd.n1748 gnd.n1702 256.663
R4288 gnd.n5319 gnd.n1702 256.663
R4289 gnd.n1745 gnd.n1702 256.663
R4290 gnd.n5326 gnd.n1702 256.663
R4291 gnd.n1742 gnd.n1702 256.663
R4292 gnd.n5333 gnd.n1702 256.663
R4293 gnd.n1739 gnd.n1702 256.663
R4294 gnd.n5340 gnd.n1702 256.663
R4295 gnd.n5343 gnd.n1702 256.663
R4296 gnd.n4071 gnd.n3763 242.672
R4297 gnd.n4071 gnd.n3764 242.672
R4298 gnd.n4071 gnd.n3765 242.672
R4299 gnd.n4071 gnd.n3766 242.672
R4300 gnd.n4071 gnd.n3767 242.672
R4301 gnd.n4071 gnd.n3768 242.672
R4302 gnd.n4071 gnd.n3769 242.672
R4303 gnd.n4071 gnd.n3770 242.672
R4304 gnd.n4071 gnd.n3771 242.672
R4305 gnd.n5956 gnd.n1154 242.672
R4306 gnd.n5956 gnd.n1153 242.672
R4307 gnd.n5956 gnd.n1152 242.672
R4308 gnd.n5956 gnd.n1151 242.672
R4309 gnd.n5956 gnd.n1150 242.672
R4310 gnd.n5956 gnd.n1149 242.672
R4311 gnd.n5956 gnd.n1148 242.672
R4312 gnd.n5956 gnd.n1147 242.672
R4313 gnd.n5956 gnd.n1146 242.672
R4314 gnd.n2882 gnd.n2881 242.672
R4315 gnd.n2882 gnd.n2792 242.672
R4316 gnd.n2882 gnd.n2793 242.672
R4317 gnd.n2882 gnd.n2794 242.672
R4318 gnd.n2882 gnd.n2795 242.672
R4319 gnd.n2882 gnd.n2796 242.672
R4320 gnd.n2882 gnd.n2797 242.672
R4321 gnd.n2882 gnd.n2798 242.672
R4322 gnd.n2882 gnd.n2799 242.672
R4323 gnd.n2882 gnd.n2800 242.672
R4324 gnd.n2882 gnd.n2801 242.672
R4325 gnd.n2882 gnd.n2802 242.672
R4326 gnd.n2883 gnd.n2882 242.672
R4327 gnd.n3735 gnd.n2287 242.672
R4328 gnd.n3735 gnd.n2286 242.672
R4329 gnd.n3735 gnd.n2285 242.672
R4330 gnd.n3735 gnd.n2284 242.672
R4331 gnd.n3735 gnd.n2283 242.672
R4332 gnd.n3735 gnd.n2282 242.672
R4333 gnd.n3735 gnd.n2281 242.672
R4334 gnd.n3735 gnd.n2280 242.672
R4335 gnd.n3735 gnd.n2279 242.672
R4336 gnd.n3735 gnd.n2278 242.672
R4337 gnd.n3735 gnd.n2277 242.672
R4338 gnd.n3735 gnd.n2276 242.672
R4339 gnd.n3735 gnd.n2275 242.672
R4340 gnd.n5653 gnd.n1476 242.672
R4341 gnd.n5653 gnd.n1478 242.672
R4342 gnd.n5653 gnd.n1479 242.672
R4343 gnd.n5653 gnd.n1481 242.672
R4344 gnd.n5653 gnd.n1483 242.672
R4345 gnd.n5653 gnd.n1484 242.672
R4346 gnd.n5653 gnd.n1486 242.672
R4347 gnd.n5653 gnd.n1488 242.672
R4348 gnd.n5654 gnd.n5653 242.672
R4349 gnd.n197 gnd.n165 242.672
R4350 gnd.n253 gnd.n165 242.672
R4351 gnd.n193 gnd.n165 242.672
R4352 gnd.n260 gnd.n165 242.672
R4353 gnd.n186 gnd.n165 242.672
R4354 gnd.n267 gnd.n165 242.672
R4355 gnd.n179 gnd.n165 242.672
R4356 gnd.n274 gnd.n165 242.672
R4357 gnd.n172 gnd.n165 242.672
R4358 gnd.n2966 gnd.n2965 242.672
R4359 gnd.n2965 gnd.n2704 242.672
R4360 gnd.n2965 gnd.n2705 242.672
R4361 gnd.n2965 gnd.n2706 242.672
R4362 gnd.n2965 gnd.n2707 242.672
R4363 gnd.n2965 gnd.n2708 242.672
R4364 gnd.n2965 gnd.n2709 242.672
R4365 gnd.n2965 gnd.n2710 242.672
R4366 gnd.n3735 gnd.n2288 242.672
R4367 gnd.n3735 gnd.n2289 242.672
R4368 gnd.n3735 gnd.n2290 242.672
R4369 gnd.n3735 gnd.n2291 242.672
R4370 gnd.n3735 gnd.n2292 242.672
R4371 gnd.n3735 gnd.n2293 242.672
R4372 gnd.n3735 gnd.n2294 242.672
R4373 gnd.n3735 gnd.n2295 242.672
R4374 gnd.n4071 gnd.n4070 242.672
R4375 gnd.n4071 gnd.n3736 242.672
R4376 gnd.n4071 gnd.n3737 242.672
R4377 gnd.n4071 gnd.n3738 242.672
R4378 gnd.n4071 gnd.n3739 242.672
R4379 gnd.n4071 gnd.n3740 242.672
R4380 gnd.n4071 gnd.n3741 242.672
R4381 gnd.n4071 gnd.n3742 242.672
R4382 gnd.n4071 gnd.n3743 242.672
R4383 gnd.n4071 gnd.n3744 242.672
R4384 gnd.n4071 gnd.n3745 242.672
R4385 gnd.n4071 gnd.n3746 242.672
R4386 gnd.n4071 gnd.n3747 242.672
R4387 gnd.n4071 gnd.n3748 242.672
R4388 gnd.n4071 gnd.n3749 242.672
R4389 gnd.n4071 gnd.n3750 242.672
R4390 gnd.n4071 gnd.n3751 242.672
R4391 gnd.n4071 gnd.n3752 242.672
R4392 gnd.n4071 gnd.n3753 242.672
R4393 gnd.n4071 gnd.n3754 242.672
R4394 gnd.n4071 gnd.n3755 242.672
R4395 gnd.n4071 gnd.n3756 242.672
R4396 gnd.n4071 gnd.n3757 242.672
R4397 gnd.n4071 gnd.n3758 242.672
R4398 gnd.n4071 gnd.n3759 242.672
R4399 gnd.n4071 gnd.n3760 242.672
R4400 gnd.n4071 gnd.n3761 242.672
R4401 gnd.n4071 gnd.n3762 242.672
R4402 gnd.n4072 gnd.n4071 242.672
R4403 gnd.n5956 gnd.n1156 242.672
R4404 gnd.n5956 gnd.n1157 242.672
R4405 gnd.n5956 gnd.n1158 242.672
R4406 gnd.n5956 gnd.n1159 242.672
R4407 gnd.n5956 gnd.n1160 242.672
R4408 gnd.n5956 gnd.n1161 242.672
R4409 gnd.n5956 gnd.n1162 242.672
R4410 gnd.n5956 gnd.n1163 242.672
R4411 gnd.n5956 gnd.n1164 242.672
R4412 gnd.n5956 gnd.n1165 242.672
R4413 gnd.n5956 gnd.n1166 242.672
R4414 gnd.n5956 gnd.n1167 242.672
R4415 gnd.n5956 gnd.n1168 242.672
R4416 gnd.n5956 gnd.n1169 242.672
R4417 gnd.n5956 gnd.n1170 242.672
R4418 gnd.n5956 gnd.n1171 242.672
R4419 gnd.n5906 gnd.n1212 242.672
R4420 gnd.n5956 gnd.n1172 242.672
R4421 gnd.n5956 gnd.n1173 242.672
R4422 gnd.n5956 gnd.n1174 242.672
R4423 gnd.n5956 gnd.n1175 242.672
R4424 gnd.n5956 gnd.n1176 242.672
R4425 gnd.n5956 gnd.n1177 242.672
R4426 gnd.n5956 gnd.n1178 242.672
R4427 gnd.n5956 gnd.n1179 242.672
R4428 gnd.n5956 gnd.n1180 242.672
R4429 gnd.n5956 gnd.n1181 242.672
R4430 gnd.n5956 gnd.n1182 242.672
R4431 gnd.n5956 gnd.n1183 242.672
R4432 gnd.n5956 gnd.n5955 242.672
R4433 gnd.n5653 gnd.n5652 242.672
R4434 gnd.n5653 gnd.n1448 242.672
R4435 gnd.n5653 gnd.n1449 242.672
R4436 gnd.n5653 gnd.n1450 242.672
R4437 gnd.n5653 gnd.n1451 242.672
R4438 gnd.n5653 gnd.n1452 242.672
R4439 gnd.n5653 gnd.n1453 242.672
R4440 gnd.n5653 gnd.n1454 242.672
R4441 gnd.n5653 gnd.n1455 242.672
R4442 gnd.n5653 gnd.n1456 242.672
R4443 gnd.n5653 gnd.n1457 242.672
R4444 gnd.n5653 gnd.n1458 242.672
R4445 gnd.n5653 gnd.n1459 242.672
R4446 gnd.n5600 gnd.n1522 242.672
R4447 gnd.n5653 gnd.n1460 242.672
R4448 gnd.n5653 gnd.n1461 242.672
R4449 gnd.n5653 gnd.n1462 242.672
R4450 gnd.n5653 gnd.n1463 242.672
R4451 gnd.n5653 gnd.n1464 242.672
R4452 gnd.n5653 gnd.n1465 242.672
R4453 gnd.n5653 gnd.n1466 242.672
R4454 gnd.n5653 gnd.n1467 242.672
R4455 gnd.n5653 gnd.n1468 242.672
R4456 gnd.n5653 gnd.n1469 242.672
R4457 gnd.n5653 gnd.n1470 242.672
R4458 gnd.n5653 gnd.n1471 242.672
R4459 gnd.n5653 gnd.n1472 242.672
R4460 gnd.n5653 gnd.n1473 242.672
R4461 gnd.n5653 gnd.n1474 242.672
R4462 gnd.n5653 gnd.n1475 242.672
R4463 gnd.n489 gnd.n165 242.672
R4464 gnd.n285 gnd.n165 242.672
R4465 gnd.n479 gnd.n165 242.672
R4466 gnd.n289 gnd.n165 242.672
R4467 gnd.n469 gnd.n165 242.672
R4468 gnd.n293 gnd.n165 242.672
R4469 gnd.n459 gnd.n165 242.672
R4470 gnd.n297 gnd.n165 242.672
R4471 gnd.n449 gnd.n165 242.672
R4472 gnd.n301 gnd.n165 242.672
R4473 gnd.n439 gnd.n165 242.672
R4474 gnd.n307 gnd.n165 242.672
R4475 gnd.n429 gnd.n165 242.672
R4476 gnd.n311 gnd.n165 242.672
R4477 gnd.n419 gnd.n165 242.672
R4478 gnd.n315 gnd.n165 242.672
R4479 gnd.n409 gnd.n165 242.672
R4480 gnd.n319 gnd.n165 242.672
R4481 gnd.n399 gnd.n165 242.672
R4482 gnd.n323 gnd.n165 242.672
R4483 gnd.n389 gnd.n165 242.672
R4484 gnd.n379 gnd.n165 242.672
R4485 gnd.n378 gnd.n165 242.672
R4486 gnd.n333 gnd.n165 242.672
R4487 gnd.n368 gnd.n165 242.672
R4488 gnd.n337 gnd.n165 242.672
R4489 gnd.n358 gnd.n165 242.672
R4490 gnd.n341 gnd.n165 242.672
R4491 gnd.n348 gnd.n165 242.672
R4492 gnd.n4579 gnd.n2104 242.672
R4493 gnd.n4579 gnd.n2105 242.672
R4494 gnd.n4579 gnd.n2106 242.672
R4495 gnd.n4579 gnd.n2107 242.672
R4496 gnd.n4579 gnd.n2108 242.672
R4497 gnd.n4579 gnd.n2109 242.672
R4498 gnd.n4579 gnd.n2110 242.672
R4499 gnd.n4579 gnd.n2111 242.672
R4500 gnd.n4579 gnd.n2112 242.672
R4501 gnd.n4579 gnd.n2113 242.672
R4502 gnd.n4579 gnd.n2114 242.672
R4503 gnd.n4579 gnd.n2115 242.672
R4504 gnd.n4579 gnd.n2116 242.672
R4505 gnd.n4579 gnd.n2117 242.672
R4506 gnd.n5426 gnd.n1661 242.672
R4507 gnd.n5426 gnd.n1658 242.672
R4508 gnd.n5426 gnd.n1656 242.672
R4509 gnd.n5426 gnd.n1655 242.672
R4510 gnd.n5426 gnd.n1653 242.672
R4511 gnd.n5426 gnd.n1651 242.672
R4512 gnd.n5426 gnd.n1650 242.672
R4513 gnd.n5426 gnd.n1648 242.672
R4514 gnd.n5426 gnd.n1646 242.672
R4515 gnd.n5426 gnd.n1645 242.672
R4516 gnd.n5426 gnd.n1643 242.672
R4517 gnd.n5426 gnd.n1642 242.672
R4518 gnd.n5426 gnd.n1640 242.672
R4519 gnd.n5427 gnd.n5426 242.672
R4520 gnd.n347 gnd.n161 240.244
R4521 gnd.n350 gnd.n349 240.244
R4522 gnd.n357 gnd.n356 240.244
R4523 gnd.n360 gnd.n359 240.244
R4524 gnd.n367 gnd.n366 240.244
R4525 gnd.n370 gnd.n369 240.244
R4526 gnd.n377 gnd.n376 240.244
R4527 gnd.n381 gnd.n380 240.244
R4528 gnd.n388 gnd.n329 240.244
R4529 gnd.n391 gnd.n390 240.244
R4530 gnd.n398 gnd.n397 240.244
R4531 gnd.n401 gnd.n400 240.244
R4532 gnd.n408 gnd.n407 240.244
R4533 gnd.n411 gnd.n410 240.244
R4534 gnd.n418 gnd.n417 240.244
R4535 gnd.n421 gnd.n420 240.244
R4536 gnd.n428 gnd.n427 240.244
R4537 gnd.n431 gnd.n430 240.244
R4538 gnd.n438 gnd.n437 240.244
R4539 gnd.n441 gnd.n440 240.244
R4540 gnd.n448 gnd.n447 240.244
R4541 gnd.n451 gnd.n450 240.244
R4542 gnd.n458 gnd.n457 240.244
R4543 gnd.n461 gnd.n460 240.244
R4544 gnd.n468 gnd.n467 240.244
R4545 gnd.n471 gnd.n470 240.244
R4546 gnd.n478 gnd.n477 240.244
R4547 gnd.n481 gnd.n480 240.244
R4548 gnd.n488 gnd.n487 240.244
R4549 gnd.n5533 gnd.n1555 240.244
R4550 gnd.n5525 gnd.n1555 240.244
R4551 gnd.n5525 gnd.n1566 240.244
R4552 gnd.n1582 gnd.n1566 240.244
R4553 gnd.n5442 gnd.n1582 240.244
R4554 gnd.n5442 gnd.n1595 240.244
R4555 gnd.n5447 gnd.n1595 240.244
R4556 gnd.n5447 gnd.n1607 240.244
R4557 gnd.n5500 gnd.n1607 240.244
R4558 gnd.n5500 gnd.n1620 240.244
R4559 gnd.n1620 gnd.n547 240.244
R4560 gnd.n1616 gnd.n547 240.244
R4561 gnd.n1616 gnd.n537 240.244
R4562 gnd.n537 gnd.n530 240.244
R4563 gnd.n6756 gnd.n530 240.244
R4564 gnd.n6756 gnd.n523 240.244
R4565 gnd.n523 gnd.n518 240.244
R4566 gnd.n6761 gnd.n518 240.244
R4567 gnd.n6761 gnd.n510 240.244
R4568 gnd.n510 gnd.n505 240.244
R4569 gnd.n505 gnd.n500 240.244
R4570 gnd.n6798 gnd.n500 240.244
R4571 gnd.n6798 gnd.n69 240.244
R4572 gnd.n6807 gnd.n69 240.244
R4573 gnd.n6808 gnd.n6807 240.244
R4574 gnd.n6808 gnd.n86 240.244
R4575 gnd.n6811 gnd.n86 240.244
R4576 gnd.n6811 gnd.n97 240.244
R4577 gnd.n6815 gnd.n97 240.244
R4578 gnd.n6815 gnd.n106 240.244
R4579 gnd.n6818 gnd.n106 240.244
R4580 gnd.n6818 gnd.n115 240.244
R4581 gnd.n6822 gnd.n115 240.244
R4582 gnd.n6822 gnd.n125 240.244
R4583 gnd.n6825 gnd.n125 240.244
R4584 gnd.n6825 gnd.n134 240.244
R4585 gnd.n6829 gnd.n134 240.244
R4586 gnd.n6829 gnd.n145 240.244
R4587 gnd.n6832 gnd.n145 240.244
R4588 gnd.n6832 gnd.n154 240.244
R4589 gnd.n6835 gnd.n154 240.244
R4590 gnd.n6835 gnd.n163 240.244
R4591 gnd.n1491 gnd.n1490 240.244
R4592 gnd.n5646 gnd.n1490 240.244
R4593 gnd.n5644 gnd.n5643 240.244
R4594 gnd.n5640 gnd.n5639 240.244
R4595 gnd.n5636 gnd.n5635 240.244
R4596 gnd.n5632 gnd.n5631 240.244
R4597 gnd.n5628 gnd.n5627 240.244
R4598 gnd.n5624 gnd.n5623 240.244
R4599 gnd.n5620 gnd.n5619 240.244
R4600 gnd.n5615 gnd.n5614 240.244
R4601 gnd.n5611 gnd.n5610 240.244
R4602 gnd.n5607 gnd.n5606 240.244
R4603 gnd.n5603 gnd.n5602 240.244
R4604 gnd.n5598 gnd.n5597 240.244
R4605 gnd.n5594 gnd.n5593 240.244
R4606 gnd.n5590 gnd.n5589 240.244
R4607 gnd.n5586 gnd.n5585 240.244
R4608 gnd.n5582 gnd.n5581 240.244
R4609 gnd.n5578 gnd.n5577 240.244
R4610 gnd.n5574 gnd.n5573 240.244
R4611 gnd.n5570 gnd.n5569 240.244
R4612 gnd.n5566 gnd.n5565 240.244
R4613 gnd.n5562 gnd.n5561 240.244
R4614 gnd.n5558 gnd.n5557 240.244
R4615 gnd.n5554 gnd.n5553 240.244
R4616 gnd.n5550 gnd.n5549 240.244
R4617 gnd.n5546 gnd.n5545 240.244
R4618 gnd.n5542 gnd.n5541 240.244
R4619 gnd.n1570 gnd.n1492 240.244
R4620 gnd.n5523 gnd.n1570 240.244
R4621 gnd.n5523 gnd.n1571 240.244
R4622 gnd.n5519 gnd.n1571 240.244
R4623 gnd.n5519 gnd.n1580 240.244
R4624 gnd.n5511 gnd.n1580 240.244
R4625 gnd.n5511 gnd.n1598 240.244
R4626 gnd.n5507 gnd.n1598 240.244
R4627 gnd.n5507 gnd.n1605 240.244
R4628 gnd.n1605 gnd.n545 240.244
R4629 gnd.n6737 gnd.n545 240.244
R4630 gnd.n6737 gnd.n540 240.244
R4631 gnd.n6746 gnd.n540 240.244
R4632 gnd.n6746 gnd.n541 240.244
R4633 gnd.n541 gnd.n520 240.244
R4634 gnd.n6770 gnd.n520 240.244
R4635 gnd.n6773 gnd.n6770 240.244
R4636 gnd.n6773 gnd.n508 240.244
R4637 gnd.n6783 gnd.n508 240.244
R4638 gnd.n6789 gnd.n6783 240.244
R4639 gnd.n6789 gnd.n6786 240.244
R4640 gnd.n6786 gnd.n72 240.244
R4641 gnd.n6896 gnd.n72 240.244
R4642 gnd.n6896 gnd.n73 240.244
R4643 gnd.n83 gnd.n73 240.244
R4644 gnd.n6890 gnd.n83 240.244
R4645 gnd.n6890 gnd.n84 240.244
R4646 gnd.n6882 gnd.n84 240.244
R4647 gnd.n6882 gnd.n100 240.244
R4648 gnd.n6878 gnd.n100 240.244
R4649 gnd.n6878 gnd.n105 240.244
R4650 gnd.n6870 gnd.n105 240.244
R4651 gnd.n6870 gnd.n117 240.244
R4652 gnd.n6866 gnd.n117 240.244
R4653 gnd.n6866 gnd.n123 240.244
R4654 gnd.n6858 gnd.n123 240.244
R4655 gnd.n6858 gnd.n137 240.244
R4656 gnd.n6854 gnd.n137 240.244
R4657 gnd.n6854 gnd.n143 240.244
R4658 gnd.n6846 gnd.n143 240.244
R4659 gnd.n6846 gnd.n156 240.244
R4660 gnd.n6842 gnd.n156 240.244
R4661 gnd.n5957 gnd.n1143 240.244
R4662 gnd.n5954 gnd.n1184 240.244
R4663 gnd.n5950 gnd.n5949 240.244
R4664 gnd.n5946 gnd.n5945 240.244
R4665 gnd.n5942 gnd.n5941 240.244
R4666 gnd.n5938 gnd.n5937 240.244
R4667 gnd.n5934 gnd.n5933 240.244
R4668 gnd.n5930 gnd.n5929 240.244
R4669 gnd.n5926 gnd.n5925 240.244
R4670 gnd.n5921 gnd.n5920 240.244
R4671 gnd.n5917 gnd.n5916 240.244
R4672 gnd.n5913 gnd.n5912 240.244
R4673 gnd.n5909 gnd.n5908 240.244
R4674 gnd.n4450 gnd.n4449 240.244
R4675 gnd.n4453 gnd.n4452 240.244
R4676 gnd.n4460 gnd.n4459 240.244
R4677 gnd.n4463 gnd.n4462 240.244
R4678 gnd.n4468 gnd.n4443 240.244
R4679 gnd.n4472 gnd.n4471 240.244
R4680 gnd.n4479 gnd.n4478 240.244
R4681 gnd.n4482 gnd.n4481 240.244
R4682 gnd.n4489 gnd.n4488 240.244
R4683 gnd.n4492 gnd.n4491 240.244
R4684 gnd.n4499 gnd.n4498 240.244
R4685 gnd.n4502 gnd.n4501 240.244
R4686 gnd.n4509 gnd.n4508 240.244
R4687 gnd.n4512 gnd.n4511 240.244
R4688 gnd.n4517 gnd.n4430 240.244
R4689 gnd.n4074 gnd.n2261 240.244
R4690 gnd.n2261 gnd.n2251 240.244
R4691 gnd.n4090 gnd.n2251 240.244
R4692 gnd.n4091 gnd.n4090 240.244
R4693 gnd.n4091 gnd.n2242 240.244
R4694 gnd.n2242 gnd.n2233 240.244
R4695 gnd.n4110 gnd.n2233 240.244
R4696 gnd.n4111 gnd.n4110 240.244
R4697 gnd.n4111 gnd.n2225 240.244
R4698 gnd.n2225 gnd.n2215 240.244
R4699 gnd.n4130 gnd.n2215 240.244
R4700 gnd.n4131 gnd.n4130 240.244
R4701 gnd.n4131 gnd.n2206 240.244
R4702 gnd.n2206 gnd.n2197 240.244
R4703 gnd.n4151 gnd.n2197 240.244
R4704 gnd.n4152 gnd.n4151 240.244
R4705 gnd.n4152 gnd.n2189 240.244
R4706 gnd.n2189 gnd.n2181 240.244
R4707 gnd.n4171 gnd.n2181 240.244
R4708 gnd.n4172 gnd.n4171 240.244
R4709 gnd.n4172 gnd.n2170 240.244
R4710 gnd.n4175 gnd.n2170 240.244
R4711 gnd.n4175 gnd.n2164 240.244
R4712 gnd.n4178 gnd.n2164 240.244
R4713 gnd.n4178 gnd.n1051 240.244
R4714 gnd.n4207 gnd.n1051 240.244
R4715 gnd.n4207 gnd.n1063 240.244
R4716 gnd.n2154 gnd.n1063 240.244
R4717 gnd.n2154 gnd.n1074 240.244
R4718 gnd.n4216 gnd.n1074 240.244
R4719 gnd.n4216 gnd.n1085 240.244
R4720 gnd.n2148 gnd.n1085 240.244
R4721 gnd.n2148 gnd.n1094 240.244
R4722 gnd.n4261 gnd.n1094 240.244
R4723 gnd.n4261 gnd.n1105 240.244
R4724 gnd.n2137 gnd.n1105 240.244
R4725 gnd.n2137 gnd.n1114 240.244
R4726 gnd.n4268 gnd.n1114 240.244
R4727 gnd.n4268 gnd.n1125 240.244
R4728 gnd.n4528 gnd.n1125 240.244
R4729 gnd.n4528 gnd.n1135 240.244
R4730 gnd.n2126 gnd.n1135 240.244
R4731 gnd.n3774 gnd.n3773 240.244
R4732 gnd.n4064 gnd.n3773 240.244
R4733 gnd.n4062 gnd.n4061 240.244
R4734 gnd.n4058 gnd.n4057 240.244
R4735 gnd.n4054 gnd.n4053 240.244
R4736 gnd.n4050 gnd.n4049 240.244
R4737 gnd.n4046 gnd.n4045 240.244
R4738 gnd.n4042 gnd.n4041 240.244
R4739 gnd.n4038 gnd.n4037 240.244
R4740 gnd.n4033 gnd.n4032 240.244
R4741 gnd.n4029 gnd.n4028 240.244
R4742 gnd.n4025 gnd.n4024 240.244
R4743 gnd.n4021 gnd.n4020 240.244
R4744 gnd.n4017 gnd.n4016 240.244
R4745 gnd.n4013 gnd.n4012 240.244
R4746 gnd.n4009 gnd.n4008 240.244
R4747 gnd.n4005 gnd.n4004 240.244
R4748 gnd.n4001 gnd.n4000 240.244
R4749 gnd.n3997 gnd.n3996 240.244
R4750 gnd.n3993 gnd.n3992 240.244
R4751 gnd.n3989 gnd.n3988 240.244
R4752 gnd.n3985 gnd.n3984 240.244
R4753 gnd.n3981 gnd.n3980 240.244
R4754 gnd.n3977 gnd.n3976 240.244
R4755 gnd.n3973 gnd.n3972 240.244
R4756 gnd.n3969 gnd.n3968 240.244
R4757 gnd.n3965 gnd.n3964 240.244
R4758 gnd.n3961 gnd.n3960 240.244
R4759 gnd.n3957 gnd.n2272 240.244
R4760 gnd.n4082 gnd.n2259 240.244
R4761 gnd.n4082 gnd.n2255 240.244
R4762 gnd.n4088 gnd.n2255 240.244
R4763 gnd.n4088 gnd.n2240 240.244
R4764 gnd.n4102 gnd.n2240 240.244
R4765 gnd.n4102 gnd.n2236 240.244
R4766 gnd.n4108 gnd.n2236 240.244
R4767 gnd.n4108 gnd.n2223 240.244
R4768 gnd.n4122 gnd.n2223 240.244
R4769 gnd.n4122 gnd.n2219 240.244
R4770 gnd.n4128 gnd.n2219 240.244
R4771 gnd.n4128 gnd.n2204 240.244
R4772 gnd.n4142 gnd.n2204 240.244
R4773 gnd.n4142 gnd.n2200 240.244
R4774 gnd.n4149 gnd.n2200 240.244
R4775 gnd.n4149 gnd.n2187 240.244
R4776 gnd.n4163 gnd.n2187 240.244
R4777 gnd.n4163 gnd.n2185 240.244
R4778 gnd.n4169 gnd.n2185 240.244
R4779 gnd.n4169 gnd.n2168 240.244
R4780 gnd.n4190 gnd.n2168 240.244
R4781 gnd.n4190 gnd.n2166 240.244
R4782 gnd.n4196 gnd.n2166 240.244
R4783 gnd.n4196 gnd.n1055 240.244
R4784 gnd.n6011 gnd.n1055 240.244
R4785 gnd.n6011 gnd.n1056 240.244
R4786 gnd.n6007 gnd.n1056 240.244
R4787 gnd.n6007 gnd.n1061 240.244
R4788 gnd.n5999 gnd.n1061 240.244
R4789 gnd.n5999 gnd.n1077 240.244
R4790 gnd.n5995 gnd.n1077 240.244
R4791 gnd.n5995 gnd.n1083 240.244
R4792 gnd.n5987 gnd.n1083 240.244
R4793 gnd.n5987 gnd.n1097 240.244
R4794 gnd.n5983 gnd.n1097 240.244
R4795 gnd.n5983 gnd.n1103 240.244
R4796 gnd.n5975 gnd.n1103 240.244
R4797 gnd.n5975 gnd.n1117 240.244
R4798 gnd.n5971 gnd.n1117 240.244
R4799 gnd.n5971 gnd.n1123 240.244
R4800 gnd.n5963 gnd.n1123 240.244
R4801 gnd.n5963 gnd.n1138 240.244
R4802 gnd.n3734 gnd.n2297 240.244
R4803 gnd.n3727 gnd.n3726 240.244
R4804 gnd.n3724 gnd.n3723 240.244
R4805 gnd.n3720 gnd.n3719 240.244
R4806 gnd.n3716 gnd.n3715 240.244
R4807 gnd.n3712 gnd.n3711 240.244
R4808 gnd.n3708 gnd.n3707 240.244
R4809 gnd.n3704 gnd.n3703 240.244
R4810 gnd.n2977 gnd.n2689 240.244
R4811 gnd.n2987 gnd.n2689 240.244
R4812 gnd.n2987 gnd.n2680 240.244
R4813 gnd.n2680 gnd.n2669 240.244
R4814 gnd.n3008 gnd.n2669 240.244
R4815 gnd.n3008 gnd.n2663 240.244
R4816 gnd.n3018 gnd.n2663 240.244
R4817 gnd.n3018 gnd.n2652 240.244
R4818 gnd.n2652 gnd.n2644 240.244
R4819 gnd.n3036 gnd.n2644 240.244
R4820 gnd.n3037 gnd.n3036 240.244
R4821 gnd.n3037 gnd.n2629 240.244
R4822 gnd.n3039 gnd.n2629 240.244
R4823 gnd.n3039 gnd.n2615 240.244
R4824 gnd.n3081 gnd.n2615 240.244
R4825 gnd.n3082 gnd.n3081 240.244
R4826 gnd.n3085 gnd.n3082 240.244
R4827 gnd.n3085 gnd.n2570 240.244
R4828 gnd.n2610 gnd.n2570 240.244
R4829 gnd.n2610 gnd.n2580 240.244
R4830 gnd.n3095 gnd.n2580 240.244
R4831 gnd.n3095 gnd.n2601 240.244
R4832 gnd.n3105 gnd.n2601 240.244
R4833 gnd.n3105 gnd.n2499 240.244
R4834 gnd.n3150 gnd.n2499 240.244
R4835 gnd.n3150 gnd.n2485 240.244
R4836 gnd.n3172 gnd.n2485 240.244
R4837 gnd.n3173 gnd.n3172 240.244
R4838 gnd.n3173 gnd.n2472 240.244
R4839 gnd.n2472 gnd.n2461 240.244
R4840 gnd.n3204 gnd.n2461 240.244
R4841 gnd.n3205 gnd.n3204 240.244
R4842 gnd.n3206 gnd.n3205 240.244
R4843 gnd.n3206 gnd.n2446 240.244
R4844 gnd.n2446 gnd.n2445 240.244
R4845 gnd.n2445 gnd.n2430 240.244
R4846 gnd.n3257 gnd.n2430 240.244
R4847 gnd.n3258 gnd.n3257 240.244
R4848 gnd.n3258 gnd.n2417 240.244
R4849 gnd.n2417 gnd.n2406 240.244
R4850 gnd.n3289 gnd.n2406 240.244
R4851 gnd.n3290 gnd.n3289 240.244
R4852 gnd.n3291 gnd.n3290 240.244
R4853 gnd.n3291 gnd.n2390 240.244
R4854 gnd.n2390 gnd.n2389 240.244
R4855 gnd.n2389 gnd.n2376 240.244
R4856 gnd.n3346 gnd.n2376 240.244
R4857 gnd.n3347 gnd.n3346 240.244
R4858 gnd.n3347 gnd.n2363 240.244
R4859 gnd.n2363 gnd.n2353 240.244
R4860 gnd.n3635 gnd.n2353 240.244
R4861 gnd.n3638 gnd.n3635 240.244
R4862 gnd.n3638 gnd.n3637 240.244
R4863 gnd.n2967 gnd.n2702 240.244
R4864 gnd.n2723 gnd.n2702 240.244
R4865 gnd.n2726 gnd.n2725 240.244
R4866 gnd.n2733 gnd.n2732 240.244
R4867 gnd.n2736 gnd.n2735 240.244
R4868 gnd.n2743 gnd.n2742 240.244
R4869 gnd.n2746 gnd.n2745 240.244
R4870 gnd.n2753 gnd.n2752 240.244
R4871 gnd.n2975 gnd.n2699 240.244
R4872 gnd.n2699 gnd.n2678 240.244
R4873 gnd.n2998 gnd.n2678 240.244
R4874 gnd.n2998 gnd.n2672 240.244
R4875 gnd.n3006 gnd.n2672 240.244
R4876 gnd.n3006 gnd.n2674 240.244
R4877 gnd.n2674 gnd.n2650 240.244
R4878 gnd.n3028 gnd.n2650 240.244
R4879 gnd.n3028 gnd.n2646 240.244
R4880 gnd.n3034 gnd.n2646 240.244
R4881 gnd.n3034 gnd.n2628 240.244
R4882 gnd.n3059 gnd.n2628 240.244
R4883 gnd.n3059 gnd.n2623 240.244
R4884 gnd.n3071 gnd.n2623 240.244
R4885 gnd.n3071 gnd.n2624 240.244
R4886 gnd.n3067 gnd.n2624 240.244
R4887 gnd.n3067 gnd.n2572 240.244
R4888 gnd.n3119 gnd.n2572 240.244
R4889 gnd.n3119 gnd.n2573 240.244
R4890 gnd.n3115 gnd.n2573 240.244
R4891 gnd.n3115 gnd.n2579 240.244
R4892 gnd.n2599 gnd.n2579 240.244
R4893 gnd.n2599 gnd.n2497 240.244
R4894 gnd.n3154 gnd.n2497 240.244
R4895 gnd.n3154 gnd.n2492 240.244
R4896 gnd.n3162 gnd.n2492 240.244
R4897 gnd.n3162 gnd.n2493 240.244
R4898 gnd.n2493 gnd.n2470 240.244
R4899 gnd.n3194 gnd.n2470 240.244
R4900 gnd.n3194 gnd.n2465 240.244
R4901 gnd.n3202 gnd.n2465 240.244
R4902 gnd.n3202 gnd.n2466 240.244
R4903 gnd.n2466 gnd.n2443 240.244
R4904 gnd.n3239 gnd.n2443 240.244
R4905 gnd.n3239 gnd.n2438 240.244
R4906 gnd.n3247 gnd.n2438 240.244
R4907 gnd.n3247 gnd.n2439 240.244
R4908 gnd.n2439 gnd.n2415 240.244
R4909 gnd.n3279 gnd.n2415 240.244
R4910 gnd.n3279 gnd.n2410 240.244
R4911 gnd.n3287 gnd.n2410 240.244
R4912 gnd.n3287 gnd.n2411 240.244
R4913 gnd.n2411 gnd.n2388 240.244
R4914 gnd.n3328 gnd.n2388 240.244
R4915 gnd.n3328 gnd.n2383 240.244
R4916 gnd.n3336 gnd.n2383 240.244
R4917 gnd.n3336 gnd.n2384 240.244
R4918 gnd.n2384 gnd.n2361 240.244
R4919 gnd.n3623 gnd.n2361 240.244
R4920 gnd.n3623 gnd.n2356 240.244
R4921 gnd.n3633 gnd.n2356 240.244
R4922 gnd.n3633 gnd.n2357 240.244
R4923 gnd.n2357 gnd.n2296 240.244
R4924 gnd.n169 gnd.n166 240.244
R4925 gnd.n276 gnd.n275 240.244
R4926 gnd.n273 gnd.n173 240.244
R4927 gnd.n269 gnd.n268 240.244
R4928 gnd.n266 gnd.n180 240.244
R4929 gnd.n262 gnd.n261 240.244
R4930 gnd.n259 gnd.n187 240.244
R4931 gnd.n255 gnd.n254 240.244
R4932 gnd.n252 gnd.n194 240.244
R4933 gnd.n5469 gnd.n1558 240.244
R4934 gnd.n5469 gnd.n1567 240.244
R4935 gnd.n5436 gnd.n1567 240.244
R4936 gnd.n5436 gnd.n1583 240.244
R4937 gnd.n5437 gnd.n1583 240.244
R4938 gnd.n5437 gnd.n1596 240.244
R4939 gnd.n5449 gnd.n1596 240.244
R4940 gnd.n5449 gnd.n1608 240.244
R4941 gnd.n1621 gnd.n1608 240.244
R4942 gnd.n5450 gnd.n1621 240.244
R4943 gnd.n5450 gnd.n548 240.244
R4944 gnd.n548 gnd.n535 240.244
R4945 gnd.n6748 gnd.n535 240.244
R4946 gnd.n6748 gnd.n531 240.244
R4947 gnd.n6754 gnd.n531 240.244
R4948 gnd.n6754 gnd.n516 240.244
R4949 gnd.n6775 gnd.n516 240.244
R4950 gnd.n6775 gnd.n511 240.244
R4951 gnd.n6781 gnd.n511 240.244
R4952 gnd.n6781 gnd.n507 240.244
R4953 gnd.n507 gnd.n506 240.244
R4954 gnd.n506 gnd.n66 240.244
R4955 gnd.n6898 gnd.n66 240.244
R4956 gnd.n6898 gnd.n68 240.244
R4957 gnd.n216 gnd.n68 240.244
R4958 gnd.n216 gnd.n87 240.244
R4959 gnd.n212 gnd.n87 240.244
R4960 gnd.n212 gnd.n98 240.244
R4961 gnd.n223 gnd.n98 240.244
R4962 gnd.n223 gnd.n107 240.244
R4963 gnd.n209 gnd.n107 240.244
R4964 gnd.n209 gnd.n116 240.244
R4965 gnd.n230 gnd.n116 240.244
R4966 gnd.n230 gnd.n126 240.244
R4967 gnd.n206 gnd.n126 240.244
R4968 gnd.n206 gnd.n135 240.244
R4969 gnd.n237 gnd.n135 240.244
R4970 gnd.n237 gnd.n146 240.244
R4971 gnd.n203 gnd.n146 240.244
R4972 gnd.n203 gnd.n155 240.244
R4973 gnd.n244 gnd.n155 240.244
R4974 gnd.n244 gnd.n164 240.244
R4975 gnd.n1402 gnd.n1401 240.244
R4976 gnd.n1477 gnd.n1409 240.244
R4977 gnd.n1480 gnd.n1410 240.244
R4978 gnd.n1418 gnd.n1417 240.244
R4979 gnd.n1482 gnd.n1425 240.244
R4980 gnd.n1485 gnd.n1426 240.244
R4981 gnd.n1434 gnd.n1433 240.244
R4982 gnd.n1487 gnd.n1443 240.244
R4983 gnd.n5655 gnd.n1446 240.244
R4984 gnd.n5531 gnd.n1561 240.244
R4985 gnd.n1569 gnd.n1561 240.244
R4986 gnd.n1585 gnd.n1569 240.244
R4987 gnd.n5517 gnd.n1585 240.244
R4988 gnd.n5517 gnd.n1586 240.244
R4989 gnd.n5513 gnd.n1586 240.244
R4990 gnd.n5513 gnd.n1593 240.244
R4991 gnd.n5505 gnd.n1593 240.244
R4992 gnd.n5505 gnd.n1610 240.244
R4993 gnd.n1610 gnd.n550 240.244
R4994 gnd.n6735 gnd.n550 240.244
R4995 gnd.n6735 gnd.n551 240.244
R4996 gnd.n551 gnd.n539 240.244
R4997 gnd.n6730 gnd.n539 240.244
R4998 gnd.n6730 gnd.n524 240.244
R4999 gnd.n6768 gnd.n524 240.244
R5000 gnd.n6768 gnd.n519 240.244
R5001 gnd.n6764 gnd.n519 240.244
R5002 gnd.n6764 gnd.n504 240.244
R5003 gnd.n6791 gnd.n504 240.244
R5004 gnd.n6791 gnd.n498 240.244
R5005 gnd.n6800 gnd.n498 240.244
R5006 gnd.n6800 gnd.n71 240.244
R5007 gnd.n6803 gnd.n71 240.244
R5008 gnd.n6803 gnd.n89 240.244
R5009 gnd.n6888 gnd.n89 240.244
R5010 gnd.n6888 gnd.n90 240.244
R5011 gnd.n6884 gnd.n90 240.244
R5012 gnd.n6884 gnd.n96 240.244
R5013 gnd.n6876 gnd.n96 240.244
R5014 gnd.n6876 gnd.n108 240.244
R5015 gnd.n6872 gnd.n108 240.244
R5016 gnd.n6872 gnd.n113 240.244
R5017 gnd.n6864 gnd.n113 240.244
R5018 gnd.n6864 gnd.n128 240.244
R5019 gnd.n6860 gnd.n128 240.244
R5020 gnd.n6860 gnd.n133 240.244
R5021 gnd.n6852 gnd.n133 240.244
R5022 gnd.n6852 gnd.n148 240.244
R5023 gnd.n6848 gnd.n148 240.244
R5024 gnd.n6848 gnd.n153 240.244
R5025 gnd.n6840 gnd.n153 240.244
R5026 gnd.n2316 gnd.n2274 240.244
R5027 gnd.n3694 gnd.n3693 240.244
R5028 gnd.n3690 gnd.n3689 240.244
R5029 gnd.n3686 gnd.n3685 240.244
R5030 gnd.n3682 gnd.n3681 240.244
R5031 gnd.n3678 gnd.n3677 240.244
R5032 gnd.n3674 gnd.n3673 240.244
R5033 gnd.n3670 gnd.n3669 240.244
R5034 gnd.n3666 gnd.n3665 240.244
R5035 gnd.n3662 gnd.n3661 240.244
R5036 gnd.n3658 gnd.n3657 240.244
R5037 gnd.n3654 gnd.n3653 240.244
R5038 gnd.n3650 gnd.n3649 240.244
R5039 gnd.n2890 gnd.n2787 240.244
R5040 gnd.n2890 gnd.n2780 240.244
R5041 gnd.n2901 gnd.n2780 240.244
R5042 gnd.n2901 gnd.n2776 240.244
R5043 gnd.n2907 gnd.n2776 240.244
R5044 gnd.n2907 gnd.n2768 240.244
R5045 gnd.n2917 gnd.n2768 240.244
R5046 gnd.n2917 gnd.n2763 240.244
R5047 gnd.n2953 gnd.n2763 240.244
R5048 gnd.n2953 gnd.n2764 240.244
R5049 gnd.n2764 gnd.n2711 240.244
R5050 gnd.n2948 gnd.n2711 240.244
R5051 gnd.n2948 gnd.n2947 240.244
R5052 gnd.n2947 gnd.n2690 240.244
R5053 gnd.n2943 gnd.n2690 240.244
R5054 gnd.n2943 gnd.n2681 240.244
R5055 gnd.n2940 gnd.n2681 240.244
R5056 gnd.n2940 gnd.n2939 240.244
R5057 gnd.n2939 gnd.n2664 240.244
R5058 gnd.n2935 gnd.n2664 240.244
R5059 gnd.n2935 gnd.n2653 240.244
R5060 gnd.n2653 gnd.n2634 240.244
R5061 gnd.n3048 gnd.n2634 240.244
R5062 gnd.n3048 gnd.n2630 240.244
R5063 gnd.n3056 gnd.n2630 240.244
R5064 gnd.n3056 gnd.n2621 240.244
R5065 gnd.n2621 gnd.n2557 240.244
R5066 gnd.n3128 gnd.n2557 240.244
R5067 gnd.n3128 gnd.n2558 240.244
R5068 gnd.n2569 gnd.n2558 240.244
R5069 gnd.n2604 gnd.n2569 240.244
R5070 gnd.n2607 gnd.n2604 240.244
R5071 gnd.n2607 gnd.n2581 240.244
R5072 gnd.n2594 gnd.n2581 240.244
R5073 gnd.n2594 gnd.n2591 240.244
R5074 gnd.n2591 gnd.n2500 240.244
R5075 gnd.n3149 gnd.n2500 240.244
R5076 gnd.n3149 gnd.n2490 240.244
R5077 gnd.n3145 gnd.n2490 240.244
R5078 gnd.n3145 gnd.n2484 240.244
R5079 gnd.n3142 gnd.n2484 240.244
R5080 gnd.n3142 gnd.n2473 240.244
R5081 gnd.n3139 gnd.n2473 240.244
R5082 gnd.n3139 gnd.n2451 240.244
R5083 gnd.n3215 gnd.n2451 240.244
R5084 gnd.n3215 gnd.n2447 240.244
R5085 gnd.n3236 gnd.n2447 240.244
R5086 gnd.n3236 gnd.n2436 240.244
R5087 gnd.n3232 gnd.n2436 240.244
R5088 gnd.n3232 gnd.n2429 240.244
R5089 gnd.n3229 gnd.n2429 240.244
R5090 gnd.n3229 gnd.n2418 240.244
R5091 gnd.n3226 gnd.n2418 240.244
R5092 gnd.n3226 gnd.n2395 240.244
R5093 gnd.n3300 gnd.n2395 240.244
R5094 gnd.n3300 gnd.n2391 240.244
R5095 gnd.n3325 gnd.n2391 240.244
R5096 gnd.n3325 gnd.n2382 240.244
R5097 gnd.n3321 gnd.n2382 240.244
R5098 gnd.n3321 gnd.n2375 240.244
R5099 gnd.n3317 gnd.n2375 240.244
R5100 gnd.n3317 gnd.n2364 240.244
R5101 gnd.n3314 gnd.n2364 240.244
R5102 gnd.n3314 gnd.n2345 240.244
R5103 gnd.n3645 gnd.n2345 240.244
R5104 gnd.n2804 gnd.n2803 240.244
R5105 gnd.n2875 gnd.n2803 240.244
R5106 gnd.n2873 gnd.n2872 240.244
R5107 gnd.n2869 gnd.n2868 240.244
R5108 gnd.n2865 gnd.n2864 240.244
R5109 gnd.n2861 gnd.n2860 240.244
R5110 gnd.n2857 gnd.n2856 240.244
R5111 gnd.n2853 gnd.n2852 240.244
R5112 gnd.n2849 gnd.n2848 240.244
R5113 gnd.n2845 gnd.n2844 240.244
R5114 gnd.n2841 gnd.n2840 240.244
R5115 gnd.n2837 gnd.n2836 240.244
R5116 gnd.n2833 gnd.n2791 240.244
R5117 gnd.n2893 gnd.n2785 240.244
R5118 gnd.n2893 gnd.n2781 240.244
R5119 gnd.n2899 gnd.n2781 240.244
R5120 gnd.n2899 gnd.n2774 240.244
R5121 gnd.n2909 gnd.n2774 240.244
R5122 gnd.n2909 gnd.n2770 240.244
R5123 gnd.n2915 gnd.n2770 240.244
R5124 gnd.n2915 gnd.n2761 240.244
R5125 gnd.n2955 gnd.n2761 240.244
R5126 gnd.n2955 gnd.n2712 240.244
R5127 gnd.n2963 gnd.n2712 240.244
R5128 gnd.n2963 gnd.n2713 240.244
R5129 gnd.n2713 gnd.n2691 240.244
R5130 gnd.n2984 gnd.n2691 240.244
R5131 gnd.n2984 gnd.n2683 240.244
R5132 gnd.n2995 gnd.n2683 240.244
R5133 gnd.n2995 gnd.n2684 240.244
R5134 gnd.n2684 gnd.n2665 240.244
R5135 gnd.n3015 gnd.n2665 240.244
R5136 gnd.n3015 gnd.n2655 240.244
R5137 gnd.n3025 gnd.n2655 240.244
R5138 gnd.n3025 gnd.n2636 240.244
R5139 gnd.n3046 gnd.n2636 240.244
R5140 gnd.n3046 gnd.n2638 240.244
R5141 gnd.n2638 gnd.n2619 240.244
R5142 gnd.n3074 gnd.n2619 240.244
R5143 gnd.n3074 gnd.n2561 240.244
R5144 gnd.n3126 gnd.n2561 240.244
R5145 gnd.n3126 gnd.n2562 240.244
R5146 gnd.n3122 gnd.n2562 240.244
R5147 gnd.n3122 gnd.n2568 240.244
R5148 gnd.n2583 gnd.n2568 240.244
R5149 gnd.n3112 gnd.n2583 240.244
R5150 gnd.n3112 gnd.n2584 240.244
R5151 gnd.n3108 gnd.n2584 240.244
R5152 gnd.n3108 gnd.n2590 240.244
R5153 gnd.n2590 gnd.n2489 240.244
R5154 gnd.n3165 gnd.n2489 240.244
R5155 gnd.n3165 gnd.n2482 240.244
R5156 gnd.n3176 gnd.n2482 240.244
R5157 gnd.n3176 gnd.n2475 240.244
R5158 gnd.n3191 gnd.n2475 240.244
R5159 gnd.n3191 gnd.n2476 240.244
R5160 gnd.n2476 gnd.n2454 240.244
R5161 gnd.n3213 gnd.n2454 240.244
R5162 gnd.n3213 gnd.n2455 240.244
R5163 gnd.n2455 gnd.n2434 240.244
R5164 gnd.n3250 gnd.n2434 240.244
R5165 gnd.n3250 gnd.n2427 240.244
R5166 gnd.n3261 gnd.n2427 240.244
R5167 gnd.n3261 gnd.n2420 240.244
R5168 gnd.n3276 gnd.n2420 240.244
R5169 gnd.n3276 gnd.n2421 240.244
R5170 gnd.n2421 gnd.n2398 240.244
R5171 gnd.n3298 gnd.n2398 240.244
R5172 gnd.n3298 gnd.n2400 240.244
R5173 gnd.n2400 gnd.n2380 240.244
R5174 gnd.n3339 gnd.n2380 240.244
R5175 gnd.n3339 gnd.n2373 240.244
R5176 gnd.n3351 gnd.n2373 240.244
R5177 gnd.n3351 gnd.n2366 240.244
R5178 gnd.n3620 gnd.n2366 240.244
R5179 gnd.n3620 gnd.n2367 240.244
R5180 gnd.n2367 gnd.n2348 240.244
R5181 gnd.n3643 gnd.n2348 240.244
R5182 gnd.n4315 gnd.n1145 240.244
R5183 gnd.n4325 gnd.n4324 240.244
R5184 gnd.n4327 gnd.n4326 240.244
R5185 gnd.n4335 gnd.n4334 240.244
R5186 gnd.n4345 gnd.n4344 240.244
R5187 gnd.n4347 gnd.n4346 240.244
R5188 gnd.n4355 gnd.n4354 240.244
R5189 gnd.n4365 gnd.n4364 240.244
R5190 gnd.n4367 gnd.n4366 240.244
R5191 gnd.n3911 gnd.n2262 240.244
R5192 gnd.n3908 gnd.n2262 240.244
R5193 gnd.n3908 gnd.n2253 240.244
R5194 gnd.n3905 gnd.n2253 240.244
R5195 gnd.n3905 gnd.n2243 240.244
R5196 gnd.n3902 gnd.n2243 240.244
R5197 gnd.n3902 gnd.n2234 240.244
R5198 gnd.n3899 gnd.n2234 240.244
R5199 gnd.n3899 gnd.n2226 240.244
R5200 gnd.n3896 gnd.n2226 240.244
R5201 gnd.n3896 gnd.n2217 240.244
R5202 gnd.n3893 gnd.n2217 240.244
R5203 gnd.n3893 gnd.n2207 240.244
R5204 gnd.n3890 gnd.n2207 240.244
R5205 gnd.n3890 gnd.n2198 240.244
R5206 gnd.n3887 gnd.n2198 240.244
R5207 gnd.n3887 gnd.n2190 240.244
R5208 gnd.n3884 gnd.n2190 240.244
R5209 gnd.n3884 gnd.n2183 240.244
R5210 gnd.n3881 gnd.n2183 240.244
R5211 gnd.n3881 gnd.n2171 240.244
R5212 gnd.n2171 gnd.n2163 240.244
R5213 gnd.n4198 gnd.n2163 240.244
R5214 gnd.n4199 gnd.n4198 240.244
R5215 gnd.n4199 gnd.n1052 240.244
R5216 gnd.n4205 gnd.n1052 240.244
R5217 gnd.n4205 gnd.n1064 240.244
R5218 gnd.n4224 gnd.n1064 240.244
R5219 gnd.n4224 gnd.n1075 240.244
R5220 gnd.n4218 gnd.n1075 240.244
R5221 gnd.n4218 gnd.n1086 240.244
R5222 gnd.n4253 gnd.n1086 240.244
R5223 gnd.n4253 gnd.n1095 240.244
R5224 gnd.n4259 gnd.n1095 240.244
R5225 gnd.n4259 gnd.n1106 240.244
R5226 gnd.n4541 gnd.n1106 240.244
R5227 gnd.n4541 gnd.n1115 240.244
R5228 gnd.n2142 gnd.n1115 240.244
R5229 gnd.n2142 gnd.n1126 240.244
R5230 gnd.n4530 gnd.n1126 240.244
R5231 gnd.n4530 gnd.n1136 240.244
R5232 gnd.n4570 gnd.n1136 240.244
R5233 gnd.n3948 gnd.n3947 240.244
R5234 gnd.n3944 gnd.n3943 240.244
R5235 gnd.n3940 gnd.n3939 240.244
R5236 gnd.n3936 gnd.n3935 240.244
R5237 gnd.n3932 gnd.n3931 240.244
R5238 gnd.n3928 gnd.n3927 240.244
R5239 gnd.n3924 gnd.n3923 240.244
R5240 gnd.n3920 gnd.n3919 240.244
R5241 gnd.n3853 gnd.n3772 240.244
R5242 gnd.n4080 gnd.n2263 240.244
R5243 gnd.n4080 gnd.n2264 240.244
R5244 gnd.n2264 gnd.n2254 240.244
R5245 gnd.n2254 gnd.n2245 240.244
R5246 gnd.n4100 gnd.n2245 240.244
R5247 gnd.n4100 gnd.n2246 240.244
R5248 gnd.n2246 gnd.n2235 240.244
R5249 gnd.n2235 gnd.n2227 240.244
R5250 gnd.n4120 gnd.n2227 240.244
R5251 gnd.n4120 gnd.n2228 240.244
R5252 gnd.n2228 gnd.n2218 240.244
R5253 gnd.n2218 gnd.n2209 240.244
R5254 gnd.n4140 gnd.n2209 240.244
R5255 gnd.n4140 gnd.n2210 240.244
R5256 gnd.n2210 gnd.n2199 240.244
R5257 gnd.n2199 gnd.n2191 240.244
R5258 gnd.n4161 gnd.n2191 240.244
R5259 gnd.n4161 gnd.n2192 240.244
R5260 gnd.n2192 gnd.n2184 240.244
R5261 gnd.n2184 gnd.n2173 240.244
R5262 gnd.n4188 gnd.n2173 240.244
R5263 gnd.n4188 gnd.n2174 240.244
R5264 gnd.n2174 gnd.n2165 240.244
R5265 gnd.n4183 gnd.n2165 240.244
R5266 gnd.n4183 gnd.n1054 240.244
R5267 gnd.n1065 gnd.n1054 240.244
R5268 gnd.n6005 gnd.n1065 240.244
R5269 gnd.n6005 gnd.n1066 240.244
R5270 gnd.n6001 gnd.n1066 240.244
R5271 gnd.n6001 gnd.n1072 240.244
R5272 gnd.n5993 gnd.n1072 240.244
R5273 gnd.n5993 gnd.n1088 240.244
R5274 gnd.n5989 gnd.n1088 240.244
R5275 gnd.n5989 gnd.n1093 240.244
R5276 gnd.n5981 gnd.n1093 240.244
R5277 gnd.n5981 gnd.n1107 240.244
R5278 gnd.n5977 gnd.n1107 240.244
R5279 gnd.n5977 gnd.n1112 240.244
R5280 gnd.n5969 gnd.n1112 240.244
R5281 gnd.n5969 gnd.n1128 240.244
R5282 gnd.n5965 gnd.n1128 240.244
R5283 gnd.n5965 gnd.n1133 240.244
R5284 gnd.n6188 gnd.n879 240.244
R5285 gnd.n6188 gnd.n877 240.244
R5286 gnd.n6192 gnd.n877 240.244
R5287 gnd.n6192 gnd.n873 240.244
R5288 gnd.n6198 gnd.n873 240.244
R5289 gnd.n6198 gnd.n871 240.244
R5290 gnd.n6202 gnd.n871 240.244
R5291 gnd.n6202 gnd.n867 240.244
R5292 gnd.n6208 gnd.n867 240.244
R5293 gnd.n6208 gnd.n865 240.244
R5294 gnd.n6212 gnd.n865 240.244
R5295 gnd.n6212 gnd.n861 240.244
R5296 gnd.n6218 gnd.n861 240.244
R5297 gnd.n6218 gnd.n859 240.244
R5298 gnd.n6222 gnd.n859 240.244
R5299 gnd.n6222 gnd.n855 240.244
R5300 gnd.n6228 gnd.n855 240.244
R5301 gnd.n6228 gnd.n853 240.244
R5302 gnd.n6232 gnd.n853 240.244
R5303 gnd.n6232 gnd.n849 240.244
R5304 gnd.n6238 gnd.n849 240.244
R5305 gnd.n6238 gnd.n847 240.244
R5306 gnd.n6242 gnd.n847 240.244
R5307 gnd.n6242 gnd.n843 240.244
R5308 gnd.n6248 gnd.n843 240.244
R5309 gnd.n6248 gnd.n841 240.244
R5310 gnd.n6252 gnd.n841 240.244
R5311 gnd.n6252 gnd.n837 240.244
R5312 gnd.n6258 gnd.n837 240.244
R5313 gnd.n6258 gnd.n835 240.244
R5314 gnd.n6262 gnd.n835 240.244
R5315 gnd.n6262 gnd.n831 240.244
R5316 gnd.n6268 gnd.n831 240.244
R5317 gnd.n6268 gnd.n829 240.244
R5318 gnd.n6272 gnd.n829 240.244
R5319 gnd.n6272 gnd.n825 240.244
R5320 gnd.n6278 gnd.n825 240.244
R5321 gnd.n6278 gnd.n823 240.244
R5322 gnd.n6282 gnd.n823 240.244
R5323 gnd.n6282 gnd.n819 240.244
R5324 gnd.n6288 gnd.n819 240.244
R5325 gnd.n6288 gnd.n817 240.244
R5326 gnd.n6292 gnd.n817 240.244
R5327 gnd.n6292 gnd.n813 240.244
R5328 gnd.n6298 gnd.n813 240.244
R5329 gnd.n6298 gnd.n811 240.244
R5330 gnd.n6302 gnd.n811 240.244
R5331 gnd.n6302 gnd.n807 240.244
R5332 gnd.n6308 gnd.n807 240.244
R5333 gnd.n6308 gnd.n805 240.244
R5334 gnd.n6312 gnd.n805 240.244
R5335 gnd.n6312 gnd.n801 240.244
R5336 gnd.n6318 gnd.n801 240.244
R5337 gnd.n6318 gnd.n799 240.244
R5338 gnd.n6322 gnd.n799 240.244
R5339 gnd.n6322 gnd.n795 240.244
R5340 gnd.n6328 gnd.n795 240.244
R5341 gnd.n6328 gnd.n793 240.244
R5342 gnd.n6332 gnd.n793 240.244
R5343 gnd.n6332 gnd.n789 240.244
R5344 gnd.n6338 gnd.n789 240.244
R5345 gnd.n6338 gnd.n787 240.244
R5346 gnd.n6342 gnd.n787 240.244
R5347 gnd.n6342 gnd.n783 240.244
R5348 gnd.n6348 gnd.n783 240.244
R5349 gnd.n6348 gnd.n781 240.244
R5350 gnd.n6352 gnd.n781 240.244
R5351 gnd.n6352 gnd.n777 240.244
R5352 gnd.n6358 gnd.n777 240.244
R5353 gnd.n6358 gnd.n775 240.244
R5354 gnd.n6362 gnd.n775 240.244
R5355 gnd.n6362 gnd.n771 240.244
R5356 gnd.n6368 gnd.n771 240.244
R5357 gnd.n6368 gnd.n769 240.244
R5358 gnd.n6372 gnd.n769 240.244
R5359 gnd.n6372 gnd.n765 240.244
R5360 gnd.n6378 gnd.n765 240.244
R5361 gnd.n6378 gnd.n763 240.244
R5362 gnd.n6382 gnd.n763 240.244
R5363 gnd.n6382 gnd.n759 240.244
R5364 gnd.n6388 gnd.n759 240.244
R5365 gnd.n6388 gnd.n757 240.244
R5366 gnd.n6392 gnd.n757 240.244
R5367 gnd.n6392 gnd.n753 240.244
R5368 gnd.n6398 gnd.n753 240.244
R5369 gnd.n6398 gnd.n751 240.244
R5370 gnd.n6402 gnd.n751 240.244
R5371 gnd.n6402 gnd.n747 240.244
R5372 gnd.n6408 gnd.n747 240.244
R5373 gnd.n6408 gnd.n745 240.244
R5374 gnd.n6412 gnd.n745 240.244
R5375 gnd.n6412 gnd.n741 240.244
R5376 gnd.n6418 gnd.n741 240.244
R5377 gnd.n6418 gnd.n739 240.244
R5378 gnd.n6422 gnd.n739 240.244
R5379 gnd.n6422 gnd.n735 240.244
R5380 gnd.n6428 gnd.n735 240.244
R5381 gnd.n6428 gnd.n733 240.244
R5382 gnd.n6432 gnd.n733 240.244
R5383 gnd.n6432 gnd.n729 240.244
R5384 gnd.n6438 gnd.n729 240.244
R5385 gnd.n6438 gnd.n727 240.244
R5386 gnd.n6442 gnd.n727 240.244
R5387 gnd.n6442 gnd.n723 240.244
R5388 gnd.n6448 gnd.n723 240.244
R5389 gnd.n6448 gnd.n721 240.244
R5390 gnd.n6452 gnd.n721 240.244
R5391 gnd.n6452 gnd.n717 240.244
R5392 gnd.n6458 gnd.n717 240.244
R5393 gnd.n6458 gnd.n715 240.244
R5394 gnd.n6462 gnd.n715 240.244
R5395 gnd.n6462 gnd.n711 240.244
R5396 gnd.n6468 gnd.n711 240.244
R5397 gnd.n6468 gnd.n709 240.244
R5398 gnd.n6472 gnd.n709 240.244
R5399 gnd.n6472 gnd.n705 240.244
R5400 gnd.n6478 gnd.n705 240.244
R5401 gnd.n6478 gnd.n703 240.244
R5402 gnd.n6482 gnd.n703 240.244
R5403 gnd.n6482 gnd.n699 240.244
R5404 gnd.n6488 gnd.n699 240.244
R5405 gnd.n6488 gnd.n697 240.244
R5406 gnd.n6492 gnd.n697 240.244
R5407 gnd.n6492 gnd.n693 240.244
R5408 gnd.n6499 gnd.n693 240.244
R5409 gnd.n6499 gnd.n691 240.244
R5410 gnd.n6503 gnd.n691 240.244
R5411 gnd.n6503 gnd.n688 240.244
R5412 gnd.n6509 gnd.n686 240.244
R5413 gnd.n6513 gnd.n686 240.244
R5414 gnd.n6513 gnd.n682 240.244
R5415 gnd.n6519 gnd.n682 240.244
R5416 gnd.n6519 gnd.n680 240.244
R5417 gnd.n6523 gnd.n680 240.244
R5418 gnd.n6523 gnd.n676 240.244
R5419 gnd.n6529 gnd.n676 240.244
R5420 gnd.n6529 gnd.n674 240.244
R5421 gnd.n6533 gnd.n674 240.244
R5422 gnd.n6533 gnd.n670 240.244
R5423 gnd.n6539 gnd.n670 240.244
R5424 gnd.n6539 gnd.n668 240.244
R5425 gnd.n6543 gnd.n668 240.244
R5426 gnd.n6543 gnd.n664 240.244
R5427 gnd.n6549 gnd.n664 240.244
R5428 gnd.n6549 gnd.n662 240.244
R5429 gnd.n6553 gnd.n662 240.244
R5430 gnd.n6553 gnd.n658 240.244
R5431 gnd.n6559 gnd.n658 240.244
R5432 gnd.n6559 gnd.n656 240.244
R5433 gnd.n6563 gnd.n656 240.244
R5434 gnd.n6563 gnd.n652 240.244
R5435 gnd.n6569 gnd.n652 240.244
R5436 gnd.n6569 gnd.n650 240.244
R5437 gnd.n6573 gnd.n650 240.244
R5438 gnd.n6573 gnd.n646 240.244
R5439 gnd.n6579 gnd.n646 240.244
R5440 gnd.n6579 gnd.n644 240.244
R5441 gnd.n6583 gnd.n644 240.244
R5442 gnd.n6583 gnd.n640 240.244
R5443 gnd.n6589 gnd.n640 240.244
R5444 gnd.n6589 gnd.n638 240.244
R5445 gnd.n6593 gnd.n638 240.244
R5446 gnd.n6593 gnd.n634 240.244
R5447 gnd.n6599 gnd.n634 240.244
R5448 gnd.n6599 gnd.n632 240.244
R5449 gnd.n6603 gnd.n632 240.244
R5450 gnd.n6603 gnd.n628 240.244
R5451 gnd.n6609 gnd.n628 240.244
R5452 gnd.n6609 gnd.n626 240.244
R5453 gnd.n6613 gnd.n626 240.244
R5454 gnd.n6613 gnd.n622 240.244
R5455 gnd.n6619 gnd.n622 240.244
R5456 gnd.n6619 gnd.n620 240.244
R5457 gnd.n6623 gnd.n620 240.244
R5458 gnd.n6623 gnd.n616 240.244
R5459 gnd.n6629 gnd.n616 240.244
R5460 gnd.n6629 gnd.n614 240.244
R5461 gnd.n6633 gnd.n614 240.244
R5462 gnd.n6633 gnd.n610 240.244
R5463 gnd.n6639 gnd.n610 240.244
R5464 gnd.n6639 gnd.n608 240.244
R5465 gnd.n6643 gnd.n608 240.244
R5466 gnd.n6643 gnd.n604 240.244
R5467 gnd.n6649 gnd.n604 240.244
R5468 gnd.n6649 gnd.n602 240.244
R5469 gnd.n6653 gnd.n602 240.244
R5470 gnd.n6653 gnd.n598 240.244
R5471 gnd.n6659 gnd.n598 240.244
R5472 gnd.n6659 gnd.n596 240.244
R5473 gnd.n6663 gnd.n596 240.244
R5474 gnd.n6663 gnd.n592 240.244
R5475 gnd.n6669 gnd.n592 240.244
R5476 gnd.n6669 gnd.n590 240.244
R5477 gnd.n6673 gnd.n590 240.244
R5478 gnd.n6673 gnd.n586 240.244
R5479 gnd.n6679 gnd.n586 240.244
R5480 gnd.n6679 gnd.n584 240.244
R5481 gnd.n6683 gnd.n584 240.244
R5482 gnd.n6683 gnd.n580 240.244
R5483 gnd.n6689 gnd.n580 240.244
R5484 gnd.n6689 gnd.n578 240.244
R5485 gnd.n6693 gnd.n578 240.244
R5486 gnd.n6693 gnd.n574 240.244
R5487 gnd.n6699 gnd.n574 240.244
R5488 gnd.n6699 gnd.n572 240.244
R5489 gnd.n6703 gnd.n572 240.244
R5490 gnd.n6703 gnd.n568 240.244
R5491 gnd.n6709 gnd.n568 240.244
R5492 gnd.n6709 gnd.n566 240.244
R5493 gnd.n6714 gnd.n566 240.244
R5494 gnd.n6714 gnd.n562 240.244
R5495 gnd.n6721 gnd.n562 240.244
R5496 gnd.n4232 gnd.n1049 240.244
R5497 gnd.n4232 gnd.n4227 240.244
R5498 gnd.n4238 gnd.n4227 240.244
R5499 gnd.n4239 gnd.n4238 240.244
R5500 gnd.n4240 gnd.n4239 240.244
R5501 gnd.n4240 gnd.n2149 240.244
R5502 gnd.n4250 gnd.n2149 240.244
R5503 gnd.n4250 gnd.n2150 240.244
R5504 gnd.n2150 gnd.n2136 240.244
R5505 gnd.n4544 gnd.n2136 240.244
R5506 gnd.n4545 gnd.n4544 240.244
R5507 gnd.n4545 gnd.n2132 240.244
R5508 gnd.n4551 gnd.n2132 240.244
R5509 gnd.n4552 gnd.n4551 240.244
R5510 gnd.n4553 gnd.n4552 240.244
R5511 gnd.n4553 gnd.n2127 240.244
R5512 gnd.n4567 gnd.n2127 240.244
R5513 gnd.n4567 gnd.n2128 240.244
R5514 gnd.n4563 gnd.n2128 240.244
R5515 gnd.n4563 gnd.n4562 240.244
R5516 gnd.n4562 gnd.n2102 240.244
R5517 gnd.n4581 gnd.n2102 240.244
R5518 gnd.n4581 gnd.n2098 240.244
R5519 gnd.n4587 gnd.n2098 240.244
R5520 gnd.n4587 gnd.n2088 240.244
R5521 gnd.n4597 gnd.n2088 240.244
R5522 gnd.n4597 gnd.n2084 240.244
R5523 gnd.n4603 gnd.n2084 240.244
R5524 gnd.n4603 gnd.n2072 240.244
R5525 gnd.n4630 gnd.n2072 240.244
R5526 gnd.n4630 gnd.n2067 240.244
R5527 gnd.n4645 gnd.n2067 240.244
R5528 gnd.n4645 gnd.n2068 240.244
R5529 gnd.n4641 gnd.n2068 240.244
R5530 gnd.n4641 gnd.n4640 240.244
R5531 gnd.n4640 gnd.n1281 240.244
R5532 gnd.n5830 gnd.n1281 240.244
R5533 gnd.n5830 gnd.n1282 240.244
R5534 gnd.n5826 gnd.n1282 240.244
R5535 gnd.n5826 gnd.n1288 240.244
R5536 gnd.n2035 gnd.n1288 240.244
R5537 gnd.n4797 gnd.n2035 240.244
R5538 gnd.n4797 gnd.n2029 240.244
R5539 gnd.n4805 gnd.n2029 240.244
R5540 gnd.n4805 gnd.n2030 240.244
R5541 gnd.n2030 gnd.n2011 240.244
R5542 gnd.n4829 gnd.n2011 240.244
R5543 gnd.n4829 gnd.n2007 240.244
R5544 gnd.n4835 gnd.n2007 240.244
R5545 gnd.n4835 gnd.n1987 240.244
R5546 gnd.n4868 gnd.n1987 240.244
R5547 gnd.n4868 gnd.n1983 240.244
R5548 gnd.n4874 gnd.n1983 240.244
R5549 gnd.n4874 gnd.n1961 240.244
R5550 gnd.n4908 gnd.n1961 240.244
R5551 gnd.n4908 gnd.n1956 240.244
R5552 gnd.n4916 gnd.n1956 240.244
R5553 gnd.n4916 gnd.n1957 240.244
R5554 gnd.n1957 gnd.n1934 240.244
R5555 gnd.n4954 gnd.n1934 240.244
R5556 gnd.n4954 gnd.n1929 240.244
R5557 gnd.n4962 gnd.n1929 240.244
R5558 gnd.n4962 gnd.n1930 240.244
R5559 gnd.n1930 gnd.n1912 240.244
R5560 gnd.n5007 gnd.n1912 240.244
R5561 gnd.n5007 gnd.n1907 240.244
R5562 gnd.n5015 gnd.n1907 240.244
R5563 gnd.n5015 gnd.n1908 240.244
R5564 gnd.n1908 gnd.n1886 240.244
R5565 gnd.n5043 gnd.n1886 240.244
R5566 gnd.n5043 gnd.n1882 240.244
R5567 gnd.n5049 gnd.n1882 240.244
R5568 gnd.n5049 gnd.n1860 240.244
R5569 gnd.n5087 gnd.n1860 240.244
R5570 gnd.n5087 gnd.n1855 240.244
R5571 gnd.n5095 gnd.n1855 240.244
R5572 gnd.n5095 gnd.n1856 240.244
R5573 gnd.n1856 gnd.n1837 240.244
R5574 gnd.n5146 gnd.n1837 240.244
R5575 gnd.n5146 gnd.n1833 240.244
R5576 gnd.n5152 gnd.n1833 240.244
R5577 gnd.n5152 gnd.n1815 240.244
R5578 gnd.n5176 gnd.n1815 240.244
R5579 gnd.n5176 gnd.n1811 240.244
R5580 gnd.n5182 gnd.n1811 240.244
R5581 gnd.n5182 gnd.n1798 240.244
R5582 gnd.n5205 gnd.n1798 240.244
R5583 gnd.n5205 gnd.n1794 240.244
R5584 gnd.n5211 gnd.n1794 240.244
R5585 gnd.n5211 gnd.n1707 240.244
R5586 gnd.n5352 gnd.n1707 240.244
R5587 gnd.n5352 gnd.n1703 240.244
R5588 gnd.n5358 gnd.n1703 240.244
R5589 gnd.n5358 gnd.n1694 240.244
R5590 gnd.n5368 gnd.n1694 240.244
R5591 gnd.n5368 gnd.n1690 240.244
R5592 gnd.n5374 gnd.n1690 240.244
R5593 gnd.n5374 gnd.n1681 240.244
R5594 gnd.n5384 gnd.n1681 240.244
R5595 gnd.n5384 gnd.n1677 240.244
R5596 gnd.n5393 gnd.n1677 240.244
R5597 gnd.n5393 gnd.n1668 240.244
R5598 gnd.n5403 gnd.n1668 240.244
R5599 gnd.n5404 gnd.n5403 240.244
R5600 gnd.n5404 gnd.n1379 240.244
R5601 gnd.n1663 gnd.n1379 240.244
R5602 gnd.n5425 gnd.n1663 240.244
R5603 gnd.n5425 gnd.n1664 240.244
R5604 gnd.n5421 gnd.n1664 240.244
R5605 gnd.n5421 gnd.n5420 240.244
R5606 gnd.n5420 gnd.n5419 240.244
R5607 gnd.n5419 gnd.n1632 240.244
R5608 gnd.n5472 gnd.n1632 240.244
R5609 gnd.n5473 gnd.n5472 240.244
R5610 gnd.n5474 gnd.n5473 240.244
R5611 gnd.n5474 gnd.n1628 240.244
R5612 gnd.n5480 gnd.n1628 240.244
R5613 gnd.n5481 gnd.n5480 240.244
R5614 gnd.n5482 gnd.n5481 240.244
R5615 gnd.n5482 gnd.n1623 240.244
R5616 gnd.n5497 gnd.n1623 240.244
R5617 gnd.n5497 gnd.n1624 240.244
R5618 gnd.n5493 gnd.n1624 240.244
R5619 gnd.n5493 gnd.n5492 240.244
R5620 gnd.n5492 gnd.n557 240.244
R5621 gnd.n6727 gnd.n557 240.244
R5622 gnd.n6727 gnd.n558 240.244
R5623 gnd.n6722 gnd.n558 240.244
R5624 gnd.n6182 gnd.n883 240.244
R5625 gnd.n6178 gnd.n883 240.244
R5626 gnd.n6178 gnd.n885 240.244
R5627 gnd.n6174 gnd.n885 240.244
R5628 gnd.n6174 gnd.n890 240.244
R5629 gnd.n6170 gnd.n890 240.244
R5630 gnd.n6170 gnd.n892 240.244
R5631 gnd.n6166 gnd.n892 240.244
R5632 gnd.n6166 gnd.n898 240.244
R5633 gnd.n6162 gnd.n898 240.244
R5634 gnd.n6162 gnd.n900 240.244
R5635 gnd.n6158 gnd.n900 240.244
R5636 gnd.n6158 gnd.n906 240.244
R5637 gnd.n6154 gnd.n906 240.244
R5638 gnd.n6154 gnd.n908 240.244
R5639 gnd.n6150 gnd.n908 240.244
R5640 gnd.n6150 gnd.n914 240.244
R5641 gnd.n6146 gnd.n914 240.244
R5642 gnd.n6146 gnd.n916 240.244
R5643 gnd.n6142 gnd.n916 240.244
R5644 gnd.n6142 gnd.n922 240.244
R5645 gnd.n6138 gnd.n922 240.244
R5646 gnd.n6138 gnd.n924 240.244
R5647 gnd.n6134 gnd.n924 240.244
R5648 gnd.n6134 gnd.n930 240.244
R5649 gnd.n6130 gnd.n930 240.244
R5650 gnd.n6130 gnd.n932 240.244
R5651 gnd.n6126 gnd.n932 240.244
R5652 gnd.n6126 gnd.n938 240.244
R5653 gnd.n6122 gnd.n938 240.244
R5654 gnd.n6122 gnd.n940 240.244
R5655 gnd.n6118 gnd.n940 240.244
R5656 gnd.n6118 gnd.n946 240.244
R5657 gnd.n6114 gnd.n946 240.244
R5658 gnd.n6114 gnd.n948 240.244
R5659 gnd.n6110 gnd.n948 240.244
R5660 gnd.n6110 gnd.n954 240.244
R5661 gnd.n6106 gnd.n954 240.244
R5662 gnd.n6106 gnd.n956 240.244
R5663 gnd.n6102 gnd.n956 240.244
R5664 gnd.n6102 gnd.n962 240.244
R5665 gnd.n6098 gnd.n962 240.244
R5666 gnd.n6098 gnd.n964 240.244
R5667 gnd.n6094 gnd.n964 240.244
R5668 gnd.n6094 gnd.n970 240.244
R5669 gnd.n6090 gnd.n970 240.244
R5670 gnd.n6090 gnd.n972 240.244
R5671 gnd.n6086 gnd.n972 240.244
R5672 gnd.n6086 gnd.n978 240.244
R5673 gnd.n6082 gnd.n978 240.244
R5674 gnd.n6082 gnd.n980 240.244
R5675 gnd.n6078 gnd.n980 240.244
R5676 gnd.n6078 gnd.n986 240.244
R5677 gnd.n6074 gnd.n986 240.244
R5678 gnd.n6074 gnd.n988 240.244
R5679 gnd.n6070 gnd.n988 240.244
R5680 gnd.n6070 gnd.n994 240.244
R5681 gnd.n6066 gnd.n994 240.244
R5682 gnd.n6066 gnd.n996 240.244
R5683 gnd.n6062 gnd.n996 240.244
R5684 gnd.n6062 gnd.n1002 240.244
R5685 gnd.n6058 gnd.n1002 240.244
R5686 gnd.n6058 gnd.n1004 240.244
R5687 gnd.n6054 gnd.n1004 240.244
R5688 gnd.n6054 gnd.n1010 240.244
R5689 gnd.n6050 gnd.n1010 240.244
R5690 gnd.n6050 gnd.n1012 240.244
R5691 gnd.n6046 gnd.n1012 240.244
R5692 gnd.n6046 gnd.n1018 240.244
R5693 gnd.n6042 gnd.n1018 240.244
R5694 gnd.n6042 gnd.n1020 240.244
R5695 gnd.n6038 gnd.n1020 240.244
R5696 gnd.n6038 gnd.n1026 240.244
R5697 gnd.n6034 gnd.n1026 240.244
R5698 gnd.n6034 gnd.n1028 240.244
R5699 gnd.n6030 gnd.n1028 240.244
R5700 gnd.n6030 gnd.n1034 240.244
R5701 gnd.n6026 gnd.n1034 240.244
R5702 gnd.n6026 gnd.n1036 240.244
R5703 gnd.n6022 gnd.n1036 240.244
R5704 gnd.n6022 gnd.n1042 240.244
R5705 gnd.n6018 gnd.n1042 240.244
R5706 gnd.n6018 gnd.n1044 240.244
R5707 gnd.n6014 gnd.n1044 240.244
R5708 gnd.n4297 gnd.n2097 240.244
R5709 gnd.n4280 gnd.n2097 240.244
R5710 gnd.n4280 gnd.n2090 240.244
R5711 gnd.n4281 gnd.n2090 240.244
R5712 gnd.n4281 gnd.n2082 240.244
R5713 gnd.n4284 gnd.n2082 240.244
R5714 gnd.n4284 gnd.n2073 240.244
R5715 gnd.n2073 gnd.n2063 240.244
R5716 gnd.n4647 gnd.n2063 240.244
R5717 gnd.n4647 gnd.n2059 240.244
R5718 gnd.n4653 gnd.n2059 240.244
R5719 gnd.n4654 gnd.n4653 240.244
R5720 gnd.n4655 gnd.n4654 240.244
R5721 gnd.n4655 gnd.n1278 240.244
R5722 gnd.n4670 gnd.n1278 240.244
R5723 gnd.n4670 gnd.n1289 240.244
R5724 gnd.n4660 gnd.n1289 240.244
R5725 gnd.n4661 gnd.n4660 240.244
R5726 gnd.n4661 gnd.n2037 240.244
R5727 gnd.n2037 gnd.n2025 240.244
R5728 gnd.n4807 gnd.n2025 240.244
R5729 gnd.n4807 gnd.n2020 240.244
R5730 gnd.n4816 gnd.n2020 240.244
R5731 gnd.n4816 gnd.n2013 240.244
R5732 gnd.n2013 gnd.n2004 240.244
R5733 gnd.n4837 gnd.n2004 240.244
R5734 gnd.n4838 gnd.n4837 240.244
R5735 gnd.n4838 gnd.n1989 240.244
R5736 gnd.n4850 gnd.n1989 240.244
R5737 gnd.n4850 gnd.n1981 240.244
R5738 gnd.n4843 gnd.n1981 240.244
R5739 gnd.n4843 gnd.n1963 240.244
R5740 gnd.n1963 gnd.n1954 240.244
R5741 gnd.n4918 gnd.n1954 240.244
R5742 gnd.n4918 gnd.n1949 240.244
R5743 gnd.n4925 gnd.n1949 240.244
R5744 gnd.n4925 gnd.n1935 240.244
R5745 gnd.n1935 gnd.n1927 240.244
R5746 gnd.n4964 gnd.n1927 240.244
R5747 gnd.n4964 gnd.n1922 240.244
R5748 gnd.n4996 gnd.n1922 240.244
R5749 gnd.n4996 gnd.n1914 240.244
R5750 gnd.n4970 gnd.n1914 240.244
R5751 gnd.n4970 gnd.n1906 240.244
R5752 gnd.n4971 gnd.n1906 240.244
R5753 gnd.n4972 gnd.n4971 240.244
R5754 gnd.n4972 gnd.n1888 240.244
R5755 gnd.n4976 gnd.n1888 240.244
R5756 gnd.n4976 gnd.n1879 240.244
R5757 gnd.n4977 gnd.n1879 240.244
R5758 gnd.n4977 gnd.n1862 240.244
R5759 gnd.n1862 gnd.n1852 240.244
R5760 gnd.n5097 gnd.n1852 240.244
R5761 gnd.n5097 gnd.n1847 240.244
R5762 gnd.n5136 gnd.n1847 240.244
R5763 gnd.n5136 gnd.n1839 240.244
R5764 gnd.n5104 gnd.n1839 240.244
R5765 gnd.n5104 gnd.n1831 240.244
R5766 gnd.n5105 gnd.n1831 240.244
R5767 gnd.n5105 gnd.n1817 240.244
R5768 gnd.n5108 gnd.n1817 240.244
R5769 gnd.n5108 gnd.n1810 240.244
R5770 gnd.n5109 gnd.n1810 240.244
R5771 gnd.n5109 gnd.n1799 240.244
R5772 gnd.n5112 gnd.n1799 240.244
R5773 gnd.n5112 gnd.n1792 240.244
R5774 gnd.n5113 gnd.n1792 240.244
R5775 gnd.n5113 gnd.n1709 240.244
R5776 gnd.n1709 gnd.n1699 240.244
R5777 gnd.n5360 gnd.n1699 240.244
R5778 gnd.n5360 gnd.n1695 240.244
R5779 gnd.n5366 gnd.n1695 240.244
R5780 gnd.n5366 gnd.n1686 240.244
R5781 gnd.n5376 gnd.n1686 240.244
R5782 gnd.n5376 gnd.n1682 240.244
R5783 gnd.n5382 gnd.n1682 240.244
R5784 gnd.n5382 gnd.n1674 240.244
R5785 gnd.n5395 gnd.n1674 240.244
R5786 gnd.n5395 gnd.n1670 240.244
R5787 gnd.n5401 gnd.n1670 240.244
R5788 gnd.n5401 gnd.n1381 240.244
R5789 gnd.n5720 gnd.n1381 240.244
R5790 gnd.n4302 gnd.n4301 240.244
R5791 gnd.n4275 gnd.n4274 240.244
R5792 gnd.n4310 gnd.n4309 240.244
R5793 gnd.n4312 gnd.n4311 240.244
R5794 gnd.n4319 gnd.n4318 240.244
R5795 gnd.n4321 gnd.n4320 240.244
R5796 gnd.n4331 gnd.n4330 240.244
R5797 gnd.n4339 gnd.n4338 240.244
R5798 gnd.n4341 gnd.n4340 240.244
R5799 gnd.n4351 gnd.n4350 240.244
R5800 gnd.n4359 gnd.n4358 240.244
R5801 gnd.n4361 gnd.n4360 240.244
R5802 gnd.n4373 gnd.n4372 240.244
R5803 gnd.n4578 gnd.n2118 240.244
R5804 gnd.n4589 gnd.n2095 240.244
R5805 gnd.n4589 gnd.n2091 240.244
R5806 gnd.n4595 gnd.n2091 240.244
R5807 gnd.n4595 gnd.n2080 240.244
R5808 gnd.n4605 gnd.n2080 240.244
R5809 gnd.n4605 gnd.n2074 240.244
R5810 gnd.n4628 gnd.n2074 240.244
R5811 gnd.n4628 gnd.n2075 240.244
R5812 gnd.n2075 gnd.n2066 240.244
R5813 gnd.n4610 gnd.n2066 240.244
R5814 gnd.n4611 gnd.n4610 240.244
R5815 gnd.n4614 gnd.n4611 240.244
R5816 gnd.n4615 gnd.n4614 240.244
R5817 gnd.n4615 gnd.n1280 240.244
R5818 gnd.n1290 gnd.n1280 240.244
R5819 gnd.n5824 gnd.n1290 240.244
R5820 gnd.n5824 gnd.n1291 240.244
R5821 gnd.n1296 gnd.n1291 240.244
R5822 gnd.n1297 gnd.n1296 240.244
R5823 gnd.n1298 gnd.n1297 240.244
R5824 gnd.n2028 gnd.n1298 240.244
R5825 gnd.n2028 gnd.n1301 240.244
R5826 gnd.n1302 gnd.n1301 240.244
R5827 gnd.n1303 gnd.n1302 240.244
R5828 gnd.n4764 gnd.n1303 240.244
R5829 gnd.n4764 gnd.n1306 240.244
R5830 gnd.n1307 gnd.n1306 240.244
R5831 gnd.n1308 gnd.n1307 240.244
R5832 gnd.n4851 gnd.n1308 240.244
R5833 gnd.n4851 gnd.n1311 240.244
R5834 gnd.n1312 gnd.n1311 240.244
R5835 gnd.n1313 gnd.n1312 240.244
R5836 gnd.n4888 gnd.n1313 240.244
R5837 gnd.n4888 gnd.n1316 240.244
R5838 gnd.n1317 gnd.n1316 240.244
R5839 gnd.n1318 gnd.n1317 240.244
R5840 gnd.n4952 gnd.n1318 240.244
R5841 gnd.n4952 gnd.n1321 240.244
R5842 gnd.n1322 gnd.n1321 240.244
R5843 gnd.n1323 gnd.n1322 240.244
R5844 gnd.n4997 gnd.n1323 240.244
R5845 gnd.n4997 gnd.n1326 240.244
R5846 gnd.n1327 gnd.n1326 240.244
R5847 gnd.n1328 gnd.n1327 240.244
R5848 gnd.n1900 gnd.n1328 240.244
R5849 gnd.n1900 gnd.n1331 240.244
R5850 gnd.n1332 gnd.n1331 240.244
R5851 gnd.n1333 gnd.n1332 240.244
R5852 gnd.n1881 gnd.n1333 240.244
R5853 gnd.n1881 gnd.n1336 240.244
R5854 gnd.n1337 gnd.n1336 240.244
R5855 gnd.n1338 gnd.n1337 240.244
R5856 gnd.n1854 gnd.n1338 240.244
R5857 gnd.n1854 gnd.n1341 240.244
R5858 gnd.n1342 gnd.n1341 240.244
R5859 gnd.n1343 gnd.n1342 240.244
R5860 gnd.n5102 gnd.n1343 240.244
R5861 gnd.n5102 gnd.n1346 240.244
R5862 gnd.n1347 gnd.n1346 240.244
R5863 gnd.n1348 gnd.n1347 240.244
R5864 gnd.n1819 gnd.n1348 240.244
R5865 gnd.n1819 gnd.n1351 240.244
R5866 gnd.n1352 gnd.n1351 240.244
R5867 gnd.n1353 gnd.n1352 240.244
R5868 gnd.n1801 gnd.n1353 240.244
R5869 gnd.n1801 gnd.n1356 240.244
R5870 gnd.n1357 gnd.n1356 240.244
R5871 gnd.n1358 gnd.n1357 240.244
R5872 gnd.n1711 gnd.n1358 240.244
R5873 gnd.n1711 gnd.n1361 240.244
R5874 gnd.n1362 gnd.n1361 240.244
R5875 gnd.n1363 gnd.n1362 240.244
R5876 gnd.n1687 gnd.n1363 240.244
R5877 gnd.n1687 gnd.n1366 240.244
R5878 gnd.n1367 gnd.n1366 240.244
R5879 gnd.n1368 gnd.n1367 240.244
R5880 gnd.n1675 gnd.n1368 240.244
R5881 gnd.n1675 gnd.n1371 240.244
R5882 gnd.n1372 gnd.n1371 240.244
R5883 gnd.n1373 gnd.n1372 240.244
R5884 gnd.n1376 gnd.n1373 240.244
R5885 gnd.n5722 gnd.n1376 240.244
R5886 gnd.n1387 gnd.n1386 240.244
R5887 gnd.n1641 gnd.n1390 240.244
R5888 gnd.n1392 gnd.n1391 240.244
R5889 gnd.n1644 gnd.n1396 240.244
R5890 gnd.n1647 gnd.n1397 240.244
R5891 gnd.n1406 gnd.n1405 240.244
R5892 gnd.n1649 gnd.n1413 240.244
R5893 gnd.n1652 gnd.n1414 240.244
R5894 gnd.n1422 gnd.n1421 240.244
R5895 gnd.n1654 gnd.n1429 240.244
R5896 gnd.n1657 gnd.n1430 240.244
R5897 gnd.n1438 gnd.n1437 240.244
R5898 gnd.n1660 gnd.n1639 240.244
R5899 gnd.n5428 gnd.n1377 240.244
R5900 gnd.n1260 gnd.n1259 240.132
R5901 gnd.n1727 gnd.n1726 240.132
R5902 gnd.n6189 gnd.n878 225.874
R5903 gnd.n6190 gnd.n6189 225.874
R5904 gnd.n6191 gnd.n6190 225.874
R5905 gnd.n6191 gnd.n872 225.874
R5906 gnd.n6199 gnd.n872 225.874
R5907 gnd.n6200 gnd.n6199 225.874
R5908 gnd.n6201 gnd.n6200 225.874
R5909 gnd.n6201 gnd.n866 225.874
R5910 gnd.n6209 gnd.n866 225.874
R5911 gnd.n6210 gnd.n6209 225.874
R5912 gnd.n6211 gnd.n6210 225.874
R5913 gnd.n6211 gnd.n860 225.874
R5914 gnd.n6219 gnd.n860 225.874
R5915 gnd.n6220 gnd.n6219 225.874
R5916 gnd.n6221 gnd.n6220 225.874
R5917 gnd.n6221 gnd.n854 225.874
R5918 gnd.n6229 gnd.n854 225.874
R5919 gnd.n6230 gnd.n6229 225.874
R5920 gnd.n6231 gnd.n6230 225.874
R5921 gnd.n6231 gnd.n848 225.874
R5922 gnd.n6239 gnd.n848 225.874
R5923 gnd.n6240 gnd.n6239 225.874
R5924 gnd.n6241 gnd.n6240 225.874
R5925 gnd.n6241 gnd.n842 225.874
R5926 gnd.n6249 gnd.n842 225.874
R5927 gnd.n6250 gnd.n6249 225.874
R5928 gnd.n6251 gnd.n6250 225.874
R5929 gnd.n6251 gnd.n836 225.874
R5930 gnd.n6259 gnd.n836 225.874
R5931 gnd.n6260 gnd.n6259 225.874
R5932 gnd.n6261 gnd.n6260 225.874
R5933 gnd.n6261 gnd.n830 225.874
R5934 gnd.n6269 gnd.n830 225.874
R5935 gnd.n6270 gnd.n6269 225.874
R5936 gnd.n6271 gnd.n6270 225.874
R5937 gnd.n6271 gnd.n824 225.874
R5938 gnd.n6279 gnd.n824 225.874
R5939 gnd.n6280 gnd.n6279 225.874
R5940 gnd.n6281 gnd.n6280 225.874
R5941 gnd.n6281 gnd.n818 225.874
R5942 gnd.n6289 gnd.n818 225.874
R5943 gnd.n6290 gnd.n6289 225.874
R5944 gnd.n6291 gnd.n6290 225.874
R5945 gnd.n6291 gnd.n812 225.874
R5946 gnd.n6299 gnd.n812 225.874
R5947 gnd.n6300 gnd.n6299 225.874
R5948 gnd.n6301 gnd.n6300 225.874
R5949 gnd.n6301 gnd.n806 225.874
R5950 gnd.n6309 gnd.n806 225.874
R5951 gnd.n6310 gnd.n6309 225.874
R5952 gnd.n6311 gnd.n6310 225.874
R5953 gnd.n6311 gnd.n800 225.874
R5954 gnd.n6319 gnd.n800 225.874
R5955 gnd.n6320 gnd.n6319 225.874
R5956 gnd.n6321 gnd.n6320 225.874
R5957 gnd.n6321 gnd.n794 225.874
R5958 gnd.n6329 gnd.n794 225.874
R5959 gnd.n6330 gnd.n6329 225.874
R5960 gnd.n6331 gnd.n6330 225.874
R5961 gnd.n6331 gnd.n788 225.874
R5962 gnd.n6339 gnd.n788 225.874
R5963 gnd.n6340 gnd.n6339 225.874
R5964 gnd.n6341 gnd.n6340 225.874
R5965 gnd.n6341 gnd.n782 225.874
R5966 gnd.n6349 gnd.n782 225.874
R5967 gnd.n6350 gnd.n6349 225.874
R5968 gnd.n6351 gnd.n6350 225.874
R5969 gnd.n6351 gnd.n776 225.874
R5970 gnd.n6359 gnd.n776 225.874
R5971 gnd.n6360 gnd.n6359 225.874
R5972 gnd.n6361 gnd.n6360 225.874
R5973 gnd.n6361 gnd.n770 225.874
R5974 gnd.n6369 gnd.n770 225.874
R5975 gnd.n6370 gnd.n6369 225.874
R5976 gnd.n6371 gnd.n6370 225.874
R5977 gnd.n6371 gnd.n764 225.874
R5978 gnd.n6379 gnd.n764 225.874
R5979 gnd.n6380 gnd.n6379 225.874
R5980 gnd.n6381 gnd.n6380 225.874
R5981 gnd.n6381 gnd.n758 225.874
R5982 gnd.n6389 gnd.n758 225.874
R5983 gnd.n6390 gnd.n6389 225.874
R5984 gnd.n6391 gnd.n6390 225.874
R5985 gnd.n6391 gnd.n752 225.874
R5986 gnd.n6399 gnd.n752 225.874
R5987 gnd.n6400 gnd.n6399 225.874
R5988 gnd.n6401 gnd.n6400 225.874
R5989 gnd.n6401 gnd.n746 225.874
R5990 gnd.n6409 gnd.n746 225.874
R5991 gnd.n6410 gnd.n6409 225.874
R5992 gnd.n6411 gnd.n6410 225.874
R5993 gnd.n6411 gnd.n740 225.874
R5994 gnd.n6419 gnd.n740 225.874
R5995 gnd.n6420 gnd.n6419 225.874
R5996 gnd.n6421 gnd.n6420 225.874
R5997 gnd.n6421 gnd.n734 225.874
R5998 gnd.n6429 gnd.n734 225.874
R5999 gnd.n6430 gnd.n6429 225.874
R6000 gnd.n6431 gnd.n6430 225.874
R6001 gnd.n6431 gnd.n728 225.874
R6002 gnd.n6439 gnd.n728 225.874
R6003 gnd.n6440 gnd.n6439 225.874
R6004 gnd.n6441 gnd.n6440 225.874
R6005 gnd.n6441 gnd.n722 225.874
R6006 gnd.n6449 gnd.n722 225.874
R6007 gnd.n6450 gnd.n6449 225.874
R6008 gnd.n6451 gnd.n6450 225.874
R6009 gnd.n6451 gnd.n716 225.874
R6010 gnd.n6459 gnd.n716 225.874
R6011 gnd.n6460 gnd.n6459 225.874
R6012 gnd.n6461 gnd.n6460 225.874
R6013 gnd.n6461 gnd.n710 225.874
R6014 gnd.n6469 gnd.n710 225.874
R6015 gnd.n6470 gnd.n6469 225.874
R6016 gnd.n6471 gnd.n6470 225.874
R6017 gnd.n6471 gnd.n704 225.874
R6018 gnd.n6479 gnd.n704 225.874
R6019 gnd.n6480 gnd.n6479 225.874
R6020 gnd.n6481 gnd.n6480 225.874
R6021 gnd.n6481 gnd.n698 225.874
R6022 gnd.n6489 gnd.n698 225.874
R6023 gnd.n6490 gnd.n6489 225.874
R6024 gnd.n6491 gnd.n6490 225.874
R6025 gnd.n6491 gnd.n692 225.874
R6026 gnd.n6500 gnd.n692 225.874
R6027 gnd.n6501 gnd.n6500 225.874
R6028 gnd.n6502 gnd.n6501 225.874
R6029 gnd.n6502 gnd.n687 225.874
R6030 gnd.n2828 gnd.t320 224.174
R6031 gnd.n2338 gnd.t312 224.174
R6032 gnd.n1522 gnd.n1459 199.319
R6033 gnd.n1522 gnd.n1460 199.319
R6034 gnd.n1212 gnd.n1172 199.319
R6035 gnd.n1212 gnd.n1171 199.319
R6036 gnd.n1261 gnd.n1258 186.49
R6037 gnd.n1728 gnd.n1725 186.49
R6038 gnd.n3604 gnd.n3603 185
R6039 gnd.n3602 gnd.n3601 185
R6040 gnd.n3581 gnd.n3580 185
R6041 gnd.n3596 gnd.n3595 185
R6042 gnd.n3594 gnd.n3593 185
R6043 gnd.n3585 gnd.n3584 185
R6044 gnd.n3588 gnd.n3587 185
R6045 gnd.n3572 gnd.n3571 185
R6046 gnd.n3570 gnd.n3569 185
R6047 gnd.n3549 gnd.n3548 185
R6048 gnd.n3564 gnd.n3563 185
R6049 gnd.n3562 gnd.n3561 185
R6050 gnd.n3553 gnd.n3552 185
R6051 gnd.n3556 gnd.n3555 185
R6052 gnd.n3540 gnd.n3539 185
R6053 gnd.n3538 gnd.n3537 185
R6054 gnd.n3517 gnd.n3516 185
R6055 gnd.n3532 gnd.n3531 185
R6056 gnd.n3530 gnd.n3529 185
R6057 gnd.n3521 gnd.n3520 185
R6058 gnd.n3524 gnd.n3523 185
R6059 gnd.n3509 gnd.n3508 185
R6060 gnd.n3507 gnd.n3506 185
R6061 gnd.n3486 gnd.n3485 185
R6062 gnd.n3501 gnd.n3500 185
R6063 gnd.n3499 gnd.n3498 185
R6064 gnd.n3490 gnd.n3489 185
R6065 gnd.n3493 gnd.n3492 185
R6066 gnd.n3477 gnd.n3476 185
R6067 gnd.n3475 gnd.n3474 185
R6068 gnd.n3454 gnd.n3453 185
R6069 gnd.n3469 gnd.n3468 185
R6070 gnd.n3467 gnd.n3466 185
R6071 gnd.n3458 gnd.n3457 185
R6072 gnd.n3461 gnd.n3460 185
R6073 gnd.n3445 gnd.n3444 185
R6074 gnd.n3443 gnd.n3442 185
R6075 gnd.n3422 gnd.n3421 185
R6076 gnd.n3437 gnd.n3436 185
R6077 gnd.n3435 gnd.n3434 185
R6078 gnd.n3426 gnd.n3425 185
R6079 gnd.n3429 gnd.n3428 185
R6080 gnd.n3413 gnd.n3412 185
R6081 gnd.n3411 gnd.n3410 185
R6082 gnd.n3390 gnd.n3389 185
R6083 gnd.n3405 gnd.n3404 185
R6084 gnd.n3403 gnd.n3402 185
R6085 gnd.n3394 gnd.n3393 185
R6086 gnd.n3397 gnd.n3396 185
R6087 gnd.n3382 gnd.n3381 185
R6088 gnd.n3380 gnd.n3379 185
R6089 gnd.n3359 gnd.n3358 185
R6090 gnd.n3374 gnd.n3373 185
R6091 gnd.n3372 gnd.n3371 185
R6092 gnd.n3363 gnd.n3362 185
R6093 gnd.n3366 gnd.n3365 185
R6094 gnd.n2829 gnd.t319 178.987
R6095 gnd.n2339 gnd.t313 178.987
R6096 gnd.n1 gnd.t62 170.774
R6097 gnd.n7 gnd.t191 170.103
R6098 gnd.n6 gnd.t201 170.103
R6099 gnd.n5 gnd.t16 170.103
R6100 gnd.n4 gnd.t14 170.103
R6101 gnd.n3 gnd.t11 170.103
R6102 gnd.n2 gnd.t48 170.103
R6103 gnd.n1 gnd.t52 170.103
R6104 gnd.n5342 gnd.n5341 163.367
R6105 gnd.n5339 gnd.n1737 163.367
R6106 gnd.n5335 gnd.n5334 163.367
R6107 gnd.n5332 gnd.n1740 163.367
R6108 gnd.n5328 gnd.n5327 163.367
R6109 gnd.n5325 gnd.n1743 163.367
R6110 gnd.n5321 gnd.n5320 163.367
R6111 gnd.n5318 gnd.n1746 163.367
R6112 gnd.n5314 gnd.n5313 163.367
R6113 gnd.n5311 gnd.n1749 163.367
R6114 gnd.n5307 gnd.n5306 163.367
R6115 gnd.n5304 gnd.n1752 163.367
R6116 gnd.n5300 gnd.n5299 163.367
R6117 gnd.n5297 gnd.n1755 163.367
R6118 gnd.n5292 gnd.n5291 163.367
R6119 gnd.n5289 gnd.n5287 163.367
R6120 gnd.n5284 gnd.n5283 163.367
R6121 gnd.n5281 gnd.n1761 163.367
R6122 gnd.n5276 gnd.n5275 163.367
R6123 gnd.n5273 gnd.n1766 163.367
R6124 gnd.n5269 gnd.n5268 163.367
R6125 gnd.n5266 gnd.n1769 163.367
R6126 gnd.n5262 gnd.n5261 163.367
R6127 gnd.n5259 gnd.n1772 163.367
R6128 gnd.n5255 gnd.n5254 163.367
R6129 gnd.n5252 gnd.n1775 163.367
R6130 gnd.n5248 gnd.n5247 163.367
R6131 gnd.n5245 gnd.n1778 163.367
R6132 gnd.n5241 gnd.n5240 163.367
R6133 gnd.n5238 gnd.n1781 163.367
R6134 gnd.n5234 gnd.n5233 163.367
R6135 gnd.n5231 gnd.n1784 163.367
R6136 gnd.n4740 gnd.n1277 163.367
R6137 gnd.n4743 gnd.n1277 163.367
R6138 gnd.n4743 gnd.n4673 163.367
R6139 gnd.n4747 gnd.n4673 163.367
R6140 gnd.n4747 gnd.n2048 163.367
R6141 gnd.n4755 gnd.n2048 163.367
R6142 gnd.n4755 gnd.n2045 163.367
R6143 gnd.n4783 gnd.n2045 163.367
R6144 gnd.n4783 gnd.n2046 163.367
R6145 gnd.n2046 gnd.n2038 163.367
R6146 gnd.n4778 gnd.n2038 163.367
R6147 gnd.n4778 gnd.n4776 163.367
R6148 gnd.n4776 gnd.n4775 163.367
R6149 gnd.n4775 gnd.n4761 163.367
R6150 gnd.n4761 gnd.n2019 163.367
R6151 gnd.n4770 gnd.n2019 163.367
R6152 gnd.n4770 gnd.n2014 163.367
R6153 gnd.n4767 gnd.n2014 163.367
R6154 gnd.n4767 gnd.n4763 163.367
R6155 gnd.n4763 gnd.n1995 163.367
R6156 gnd.n4859 gnd.n1995 163.367
R6157 gnd.n4859 gnd.n1996 163.367
R6158 gnd.n1996 gnd.n1990 163.367
R6159 gnd.n4854 gnd.n1990 163.367
R6160 gnd.n4854 gnd.n1980 163.367
R6161 gnd.n1980 gnd.n1975 163.367
R6162 gnd.n4883 gnd.n1975 163.367
R6163 gnd.n4884 gnd.n4883 163.367
R6164 gnd.n4884 gnd.n1964 163.367
R6165 gnd.n4891 gnd.n1964 163.367
R6166 gnd.n4892 gnd.n4891 163.367
R6167 gnd.n4892 gnd.n1973 163.367
R6168 gnd.n4896 gnd.n1973 163.367
R6169 gnd.n4896 gnd.n1947 163.367
R6170 gnd.n4928 gnd.n1947 163.367
R6171 gnd.n4928 gnd.n1936 163.367
R6172 gnd.n1944 gnd.n1936 163.367
R6173 gnd.n4944 gnd.n1944 163.367
R6174 gnd.n4944 gnd.n1945 163.367
R6175 gnd.n4940 gnd.n1945 163.367
R6176 gnd.n4940 gnd.n1921 163.367
R6177 gnd.n4936 gnd.n1921 163.367
R6178 gnd.n4936 gnd.n1915 163.367
R6179 gnd.n4933 gnd.n1915 163.367
R6180 gnd.n4933 gnd.n1905 163.367
R6181 gnd.n1905 gnd.n1897 163.367
R6182 gnd.n5024 gnd.n1897 163.367
R6183 gnd.n5024 gnd.n1894 163.367
R6184 gnd.n5034 gnd.n1894 163.367
R6185 gnd.n5034 gnd.n1895 163.367
R6186 gnd.n1895 gnd.n1889 163.367
R6187 gnd.n5029 gnd.n1889 163.367
R6188 gnd.n5029 gnd.n1878 163.367
R6189 gnd.n1878 gnd.n1872 163.367
R6190 gnd.n5058 gnd.n1872 163.367
R6191 gnd.n5059 gnd.n5058 163.367
R6192 gnd.n5059 gnd.n1863 163.367
R6193 gnd.n5063 gnd.n1863 163.367
R6194 gnd.n5063 gnd.n1869 163.367
R6195 gnd.n5076 gnd.n1869 163.367
R6196 gnd.n5076 gnd.n1870 163.367
R6197 gnd.n1870 gnd.n1846 163.367
R6198 gnd.n5071 gnd.n1846 163.367
R6199 gnd.n5071 gnd.n1840 163.367
R6200 gnd.n5068 gnd.n1840 163.367
R6201 gnd.n5068 gnd.n1830 163.367
R6202 gnd.n1830 gnd.n1825 163.367
R6203 gnd.n5161 gnd.n1825 163.367
R6204 gnd.n5162 gnd.n5161 163.367
R6205 gnd.n5162 gnd.n1818 163.367
R6206 gnd.n5166 gnd.n1818 163.367
R6207 gnd.n5166 gnd.n1809 163.367
R6208 gnd.n5185 gnd.n1809 163.367
R6209 gnd.n5185 gnd.n1807 163.367
R6210 gnd.n5195 gnd.n1807 163.367
R6211 gnd.n5195 gnd.n1800 163.367
R6212 gnd.n5191 gnd.n1800 163.367
R6213 gnd.n5191 gnd.n1791 163.367
R6214 gnd.n1791 gnd.n1786 163.367
R6215 gnd.n5220 gnd.n1786 163.367
R6216 gnd.n5221 gnd.n5220 163.367
R6217 gnd.n5221 gnd.n1710 163.367
R6218 gnd.n5226 gnd.n1710 163.367
R6219 gnd.n1252 gnd.n1251 163.367
R6220 gnd.n5895 gnd.n1251 163.367
R6221 gnd.n5893 gnd.n5892 163.367
R6222 gnd.n5889 gnd.n5888 163.367
R6223 gnd.n5885 gnd.n5884 163.367
R6224 gnd.n5881 gnd.n5880 163.367
R6225 gnd.n5877 gnd.n5876 163.367
R6226 gnd.n5873 gnd.n5872 163.367
R6227 gnd.n5869 gnd.n5868 163.367
R6228 gnd.n5865 gnd.n5864 163.367
R6229 gnd.n5861 gnd.n5860 163.367
R6230 gnd.n5857 gnd.n5856 163.367
R6231 gnd.n5853 gnd.n5852 163.367
R6232 gnd.n5849 gnd.n5848 163.367
R6233 gnd.n5845 gnd.n5844 163.367
R6234 gnd.n5841 gnd.n5840 163.367
R6235 gnd.n5904 gnd.n1217 163.367
R6236 gnd.n4678 gnd.n4677 163.367
R6237 gnd.n4683 gnd.n4682 163.367
R6238 gnd.n4687 gnd.n4686 163.367
R6239 gnd.n4691 gnd.n4690 163.367
R6240 gnd.n4695 gnd.n4694 163.367
R6241 gnd.n4699 gnd.n4698 163.367
R6242 gnd.n4703 gnd.n4702 163.367
R6243 gnd.n4707 gnd.n4706 163.367
R6244 gnd.n4711 gnd.n4710 163.367
R6245 gnd.n4715 gnd.n4714 163.367
R6246 gnd.n4719 gnd.n4718 163.367
R6247 gnd.n4723 gnd.n4722 163.367
R6248 gnd.n4727 gnd.n4726 163.367
R6249 gnd.n4731 gnd.n4730 163.367
R6250 gnd.n4735 gnd.n4734 163.367
R6251 gnd.n5833 gnd.n1253 163.367
R6252 gnd.n5833 gnd.n1275 163.367
R6253 gnd.n2054 gnd.n1275 163.367
R6254 gnd.n4749 gnd.n2054 163.367
R6255 gnd.n4749 gnd.n2052 163.367
R6256 gnd.n4753 gnd.n2052 163.367
R6257 gnd.n4753 gnd.n2043 163.367
R6258 gnd.n4785 gnd.n2043 163.367
R6259 gnd.n4785 gnd.n2040 163.367
R6260 gnd.n4794 gnd.n2040 163.367
R6261 gnd.n4794 gnd.n2041 163.367
R6262 gnd.n4790 gnd.n2041 163.367
R6263 gnd.n4790 gnd.n4789 163.367
R6264 gnd.n4789 gnd.n2018 163.367
R6265 gnd.n4819 gnd.n2018 163.367
R6266 gnd.n4819 gnd.n2015 163.367
R6267 gnd.n4826 gnd.n2015 163.367
R6268 gnd.n4826 gnd.n2016 163.367
R6269 gnd.n4822 gnd.n2016 163.367
R6270 gnd.n4822 gnd.n1993 163.367
R6271 gnd.n4861 gnd.n1993 163.367
R6272 gnd.n4861 gnd.n1991 163.367
R6273 gnd.n4865 gnd.n1991 163.367
R6274 gnd.n4865 gnd.n1979 163.367
R6275 gnd.n4877 gnd.n1979 163.367
R6276 gnd.n4877 gnd.n1977 163.367
R6277 gnd.n4881 gnd.n1977 163.367
R6278 gnd.n4881 gnd.n1965 163.367
R6279 gnd.n4905 gnd.n1965 163.367
R6280 gnd.n4905 gnd.n1966 163.367
R6281 gnd.n4901 gnd.n1966 163.367
R6282 gnd.n4901 gnd.n4900 163.367
R6283 gnd.n4900 gnd.n1972 163.367
R6284 gnd.n1972 gnd.n1969 163.367
R6285 gnd.n1969 gnd.n1938 163.367
R6286 gnd.n4950 gnd.n1938 163.367
R6287 gnd.n4950 gnd.n1939 163.367
R6288 gnd.n4946 gnd.n1939 163.367
R6289 gnd.n4946 gnd.n1942 163.367
R6290 gnd.n1942 gnd.n1919 163.367
R6291 gnd.n5000 gnd.n1919 163.367
R6292 gnd.n5000 gnd.n1917 163.367
R6293 gnd.n5004 gnd.n1917 163.367
R6294 gnd.n5004 gnd.n1904 163.367
R6295 gnd.n5018 gnd.n1904 163.367
R6296 gnd.n5018 gnd.n1902 163.367
R6297 gnd.n5022 gnd.n1902 163.367
R6298 gnd.n5022 gnd.n1892 163.367
R6299 gnd.n5036 gnd.n1892 163.367
R6300 gnd.n5036 gnd.n1890 163.367
R6301 gnd.n5040 gnd.n1890 163.367
R6302 gnd.n5040 gnd.n1876 163.367
R6303 gnd.n5052 gnd.n1876 163.367
R6304 gnd.n5052 gnd.n1874 163.367
R6305 gnd.n5056 gnd.n1874 163.367
R6306 gnd.n5056 gnd.n1865 163.367
R6307 gnd.n5084 gnd.n1865 163.367
R6308 gnd.n5084 gnd.n1866 163.367
R6309 gnd.n5080 gnd.n1866 163.367
R6310 gnd.n5080 gnd.n5079 163.367
R6311 gnd.n5079 gnd.n1844 163.367
R6312 gnd.n5139 gnd.n1844 163.367
R6313 gnd.n5139 gnd.n1842 163.367
R6314 gnd.n5143 gnd.n1842 163.367
R6315 gnd.n5143 gnd.n1829 163.367
R6316 gnd.n5155 gnd.n1829 163.367
R6317 gnd.n5155 gnd.n1827 163.367
R6318 gnd.n5159 gnd.n1827 163.367
R6319 gnd.n5159 gnd.n1821 163.367
R6320 gnd.n5173 gnd.n1821 163.367
R6321 gnd.n5173 gnd.n1822 163.367
R6322 gnd.n5169 gnd.n1822 163.367
R6323 gnd.n5169 gnd.n1805 163.367
R6324 gnd.n5198 gnd.n1805 163.367
R6325 gnd.n5198 gnd.n1803 163.367
R6326 gnd.n5202 gnd.n1803 163.367
R6327 gnd.n5202 gnd.n1790 163.367
R6328 gnd.n5214 gnd.n1790 163.367
R6329 gnd.n5214 gnd.n1788 163.367
R6330 gnd.n5218 gnd.n1788 163.367
R6331 gnd.n5218 gnd.n1713 163.367
R6332 gnd.n5349 gnd.n1713 163.367
R6333 gnd.n5349 gnd.n1714 163.367
R6334 gnd.n1734 gnd.n1733 156.462
R6335 gnd.n3544 gnd.n3512 153.042
R6336 gnd.n3608 gnd.n3607 152.079
R6337 gnd.n3576 gnd.n3575 152.079
R6338 gnd.n3544 gnd.n3543 152.079
R6339 gnd.n1266 gnd.n1265 152
R6340 gnd.n1267 gnd.n1256 152
R6341 gnd.n1269 gnd.n1268 152
R6342 gnd.n1271 gnd.n1254 152
R6343 gnd.n1273 gnd.n1272 152
R6344 gnd.n1732 gnd.n1716 152
R6345 gnd.n1724 gnd.n1717 152
R6346 gnd.n1723 gnd.n1722 152
R6347 gnd.n1721 gnd.n1718 152
R6348 gnd.n1719 gnd.t250 150.546
R6349 gnd.t57 gnd.n3586 147.661
R6350 gnd.t50 gnd.n3554 147.661
R6351 gnd.t46 gnd.n3522 147.661
R6352 gnd.t30 gnd.n3491 147.661
R6353 gnd.t42 gnd.n3459 147.661
R6354 gnd.t189 gnd.n3427 147.661
R6355 gnd.t199 gnd.n3395 147.661
R6356 gnd.t66 gnd.n3364 147.661
R6357 gnd.n5286 gnd.n5285 143.351
R6358 gnd.n1233 gnd.n1216 143.351
R6359 gnd.n5903 gnd.n1216 143.351
R6360 gnd.n1263 gnd.t204 130.484
R6361 gnd.n1272 gnd.t211 126.766
R6362 gnd.n1270 gnd.t301 126.766
R6363 gnd.n1256 gnd.t321 126.766
R6364 gnd.n1264 gnd.t253 126.766
R6365 gnd.n1720 gnd.t229 126.766
R6366 gnd.n1722 gnd.t273 126.766
R6367 gnd.n1731 gnd.t247 126.766
R6368 gnd.n1733 gnd.t276 126.766
R6369 gnd.n6511 gnd.n6510 106.719
R6370 gnd.n6512 gnd.n6511 106.719
R6371 gnd.n6512 gnd.n681 106.719
R6372 gnd.n6520 gnd.n681 106.719
R6373 gnd.n6521 gnd.n6520 106.719
R6374 gnd.n6522 gnd.n6521 106.719
R6375 gnd.n6522 gnd.n675 106.719
R6376 gnd.n6530 gnd.n675 106.719
R6377 gnd.n6531 gnd.n6530 106.719
R6378 gnd.n6532 gnd.n6531 106.719
R6379 gnd.n6532 gnd.n669 106.719
R6380 gnd.n6540 gnd.n669 106.719
R6381 gnd.n6541 gnd.n6540 106.719
R6382 gnd.n6542 gnd.n6541 106.719
R6383 gnd.n6542 gnd.n663 106.719
R6384 gnd.n6550 gnd.n663 106.719
R6385 gnd.n6551 gnd.n6550 106.719
R6386 gnd.n6552 gnd.n6551 106.719
R6387 gnd.n6552 gnd.n657 106.719
R6388 gnd.n6560 gnd.n657 106.719
R6389 gnd.n6561 gnd.n6560 106.719
R6390 gnd.n6562 gnd.n6561 106.719
R6391 gnd.n6562 gnd.n651 106.719
R6392 gnd.n6570 gnd.n651 106.719
R6393 gnd.n6571 gnd.n6570 106.719
R6394 gnd.n6572 gnd.n6571 106.719
R6395 gnd.n6572 gnd.n645 106.719
R6396 gnd.n6580 gnd.n645 106.719
R6397 gnd.n6581 gnd.n6580 106.719
R6398 gnd.n6582 gnd.n6581 106.719
R6399 gnd.n6582 gnd.n639 106.719
R6400 gnd.n6590 gnd.n639 106.719
R6401 gnd.n6591 gnd.n6590 106.719
R6402 gnd.n6592 gnd.n6591 106.719
R6403 gnd.n6592 gnd.n633 106.719
R6404 gnd.n6600 gnd.n633 106.719
R6405 gnd.n6601 gnd.n6600 106.719
R6406 gnd.n6602 gnd.n6601 106.719
R6407 gnd.n6602 gnd.n627 106.719
R6408 gnd.n6610 gnd.n627 106.719
R6409 gnd.n6611 gnd.n6610 106.719
R6410 gnd.n6612 gnd.n6611 106.719
R6411 gnd.n6612 gnd.n621 106.719
R6412 gnd.n6620 gnd.n621 106.719
R6413 gnd.n6621 gnd.n6620 106.719
R6414 gnd.n6622 gnd.n6621 106.719
R6415 gnd.n6622 gnd.n615 106.719
R6416 gnd.n6630 gnd.n615 106.719
R6417 gnd.n6631 gnd.n6630 106.719
R6418 gnd.n6632 gnd.n6631 106.719
R6419 gnd.n6632 gnd.n609 106.719
R6420 gnd.n6640 gnd.n609 106.719
R6421 gnd.n6641 gnd.n6640 106.719
R6422 gnd.n6642 gnd.n6641 106.719
R6423 gnd.n6642 gnd.n603 106.719
R6424 gnd.n6650 gnd.n603 106.719
R6425 gnd.n6651 gnd.n6650 106.719
R6426 gnd.n6652 gnd.n6651 106.719
R6427 gnd.n6652 gnd.n597 106.719
R6428 gnd.n6660 gnd.n597 106.719
R6429 gnd.n6661 gnd.n6660 106.719
R6430 gnd.n6662 gnd.n6661 106.719
R6431 gnd.n6662 gnd.n591 106.719
R6432 gnd.n6670 gnd.n591 106.719
R6433 gnd.n6671 gnd.n6670 106.719
R6434 gnd.n6672 gnd.n6671 106.719
R6435 gnd.n6672 gnd.n585 106.719
R6436 gnd.n6680 gnd.n585 106.719
R6437 gnd.n6681 gnd.n6680 106.719
R6438 gnd.n6682 gnd.n6681 106.719
R6439 gnd.n6682 gnd.n579 106.719
R6440 gnd.n6690 gnd.n579 106.719
R6441 gnd.n6691 gnd.n6690 106.719
R6442 gnd.n6692 gnd.n6691 106.719
R6443 gnd.n6692 gnd.n573 106.719
R6444 gnd.n6700 gnd.n573 106.719
R6445 gnd.n6701 gnd.n6700 106.719
R6446 gnd.n6702 gnd.n6701 106.719
R6447 gnd.n6702 gnd.n567 106.719
R6448 gnd.n6710 gnd.n567 106.719
R6449 gnd.n6711 gnd.n6710 106.719
R6450 gnd.n6713 gnd.n6711 106.719
R6451 gnd.n6713 gnd.n6712 106.719
R6452 gnd.n5600 gnd.n1521 105.281
R6453 gnd.n5906 gnd.n5905 105.281
R6454 gnd.n3603 gnd.n3602 104.615
R6455 gnd.n3602 gnd.n3580 104.615
R6456 gnd.n3595 gnd.n3580 104.615
R6457 gnd.n3595 gnd.n3594 104.615
R6458 gnd.n3594 gnd.n3584 104.615
R6459 gnd.n3587 gnd.n3584 104.615
R6460 gnd.n3571 gnd.n3570 104.615
R6461 gnd.n3570 gnd.n3548 104.615
R6462 gnd.n3563 gnd.n3548 104.615
R6463 gnd.n3563 gnd.n3562 104.615
R6464 gnd.n3562 gnd.n3552 104.615
R6465 gnd.n3555 gnd.n3552 104.615
R6466 gnd.n3539 gnd.n3538 104.615
R6467 gnd.n3538 gnd.n3516 104.615
R6468 gnd.n3531 gnd.n3516 104.615
R6469 gnd.n3531 gnd.n3530 104.615
R6470 gnd.n3530 gnd.n3520 104.615
R6471 gnd.n3523 gnd.n3520 104.615
R6472 gnd.n3508 gnd.n3507 104.615
R6473 gnd.n3507 gnd.n3485 104.615
R6474 gnd.n3500 gnd.n3485 104.615
R6475 gnd.n3500 gnd.n3499 104.615
R6476 gnd.n3499 gnd.n3489 104.615
R6477 gnd.n3492 gnd.n3489 104.615
R6478 gnd.n3476 gnd.n3475 104.615
R6479 gnd.n3475 gnd.n3453 104.615
R6480 gnd.n3468 gnd.n3453 104.615
R6481 gnd.n3468 gnd.n3467 104.615
R6482 gnd.n3467 gnd.n3457 104.615
R6483 gnd.n3460 gnd.n3457 104.615
R6484 gnd.n3444 gnd.n3443 104.615
R6485 gnd.n3443 gnd.n3421 104.615
R6486 gnd.n3436 gnd.n3421 104.615
R6487 gnd.n3436 gnd.n3435 104.615
R6488 gnd.n3435 gnd.n3425 104.615
R6489 gnd.n3428 gnd.n3425 104.615
R6490 gnd.n3412 gnd.n3411 104.615
R6491 gnd.n3411 gnd.n3389 104.615
R6492 gnd.n3404 gnd.n3389 104.615
R6493 gnd.n3404 gnd.n3403 104.615
R6494 gnd.n3403 gnd.n3393 104.615
R6495 gnd.n3396 gnd.n3393 104.615
R6496 gnd.n3381 gnd.n3380 104.615
R6497 gnd.n3380 gnd.n3358 104.615
R6498 gnd.n3373 gnd.n3358 104.615
R6499 gnd.n3373 gnd.n3372 104.615
R6500 gnd.n3372 gnd.n3362 104.615
R6501 gnd.n3365 gnd.n3362 104.615
R6502 gnd.n2754 gnd.t265 100.632
R6503 gnd.n2312 gnd.t296 100.632
R6504 gnd.n350 gnd.n348 99.6594
R6505 gnd.n356 gnd.n341 99.6594
R6506 gnd.n360 gnd.n358 99.6594
R6507 gnd.n366 gnd.n337 99.6594
R6508 gnd.n370 gnd.n368 99.6594
R6509 gnd.n376 gnd.n333 99.6594
R6510 gnd.n381 gnd.n378 99.6594
R6511 gnd.n379 gnd.n329 99.6594
R6512 gnd.n391 gnd.n389 99.6594
R6513 gnd.n397 gnd.n323 99.6594
R6514 gnd.n401 gnd.n399 99.6594
R6515 gnd.n407 gnd.n319 99.6594
R6516 gnd.n411 gnd.n409 99.6594
R6517 gnd.n417 gnd.n315 99.6594
R6518 gnd.n421 gnd.n419 99.6594
R6519 gnd.n427 gnd.n311 99.6594
R6520 gnd.n431 gnd.n429 99.6594
R6521 gnd.n437 gnd.n307 99.6594
R6522 gnd.n441 gnd.n439 99.6594
R6523 gnd.n447 gnd.n301 99.6594
R6524 gnd.n451 gnd.n449 99.6594
R6525 gnd.n457 gnd.n297 99.6594
R6526 gnd.n461 gnd.n459 99.6594
R6527 gnd.n467 gnd.n293 99.6594
R6528 gnd.n471 gnd.n469 99.6594
R6529 gnd.n477 gnd.n289 99.6594
R6530 gnd.n481 gnd.n479 99.6594
R6531 gnd.n487 gnd.n285 99.6594
R6532 gnd.n490 gnd.n489 99.6594
R6533 gnd.n5652 gnd.n5651 99.6594
R6534 gnd.n5646 gnd.n1448 99.6594
R6535 gnd.n5643 gnd.n1449 99.6594
R6536 gnd.n5639 gnd.n1450 99.6594
R6537 gnd.n5635 gnd.n1451 99.6594
R6538 gnd.n5631 gnd.n1452 99.6594
R6539 gnd.n5627 gnd.n1453 99.6594
R6540 gnd.n5623 gnd.n1454 99.6594
R6541 gnd.n5619 gnd.n1455 99.6594
R6542 gnd.n5614 gnd.n1456 99.6594
R6543 gnd.n5610 gnd.n1457 99.6594
R6544 gnd.n5606 gnd.n1458 99.6594
R6545 gnd.n5602 gnd.n1459 99.6594
R6546 gnd.n5597 gnd.n1461 99.6594
R6547 gnd.n5593 gnd.n1462 99.6594
R6548 gnd.n5589 gnd.n1463 99.6594
R6549 gnd.n5585 gnd.n1464 99.6594
R6550 gnd.n5581 gnd.n1465 99.6594
R6551 gnd.n5577 gnd.n1466 99.6594
R6552 gnd.n5573 gnd.n1467 99.6594
R6553 gnd.n5569 gnd.n1468 99.6594
R6554 gnd.n5565 gnd.n1469 99.6594
R6555 gnd.n5561 gnd.n1470 99.6594
R6556 gnd.n5557 gnd.n1471 99.6594
R6557 gnd.n5553 gnd.n1472 99.6594
R6558 gnd.n5549 gnd.n1473 99.6594
R6559 gnd.n5545 gnd.n1474 99.6594
R6560 gnd.n5541 gnd.n1475 99.6594
R6561 gnd.n5955 gnd.n5954 99.6594
R6562 gnd.n5950 gnd.n1183 99.6594
R6563 gnd.n5946 gnd.n1182 99.6594
R6564 gnd.n5942 gnd.n1181 99.6594
R6565 gnd.n5938 gnd.n1180 99.6594
R6566 gnd.n5934 gnd.n1179 99.6594
R6567 gnd.n5930 gnd.n1178 99.6594
R6568 gnd.n5926 gnd.n1177 99.6594
R6569 gnd.n5921 gnd.n1176 99.6594
R6570 gnd.n5917 gnd.n1175 99.6594
R6571 gnd.n5913 gnd.n1174 99.6594
R6572 gnd.n5909 gnd.n1173 99.6594
R6573 gnd.n4449 gnd.n1171 99.6594
R6574 gnd.n4453 gnd.n1170 99.6594
R6575 gnd.n4459 gnd.n1169 99.6594
R6576 gnd.n4463 gnd.n1168 99.6594
R6577 gnd.n4468 gnd.n1167 99.6594
R6578 gnd.n4472 gnd.n1166 99.6594
R6579 gnd.n4478 gnd.n1165 99.6594
R6580 gnd.n4482 gnd.n1164 99.6594
R6581 gnd.n4488 gnd.n1163 99.6594
R6582 gnd.n4492 gnd.n1162 99.6594
R6583 gnd.n4498 gnd.n1161 99.6594
R6584 gnd.n4502 gnd.n1160 99.6594
R6585 gnd.n4508 gnd.n1159 99.6594
R6586 gnd.n4512 gnd.n1158 99.6594
R6587 gnd.n4517 gnd.n1157 99.6594
R6588 gnd.n4520 gnd.n1156 99.6594
R6589 gnd.n4070 gnd.n4069 99.6594
R6590 gnd.n4064 gnd.n3736 99.6594
R6591 gnd.n4061 gnd.n3737 99.6594
R6592 gnd.n4057 gnd.n3738 99.6594
R6593 gnd.n4053 gnd.n3739 99.6594
R6594 gnd.n4049 gnd.n3740 99.6594
R6595 gnd.n4045 gnd.n3741 99.6594
R6596 gnd.n4041 gnd.n3742 99.6594
R6597 gnd.n4037 gnd.n3743 99.6594
R6598 gnd.n4032 gnd.n3744 99.6594
R6599 gnd.n4028 gnd.n3745 99.6594
R6600 gnd.n4024 gnd.n3746 99.6594
R6601 gnd.n4020 gnd.n3747 99.6594
R6602 gnd.n4016 gnd.n3748 99.6594
R6603 gnd.n4012 gnd.n3749 99.6594
R6604 gnd.n4008 gnd.n3750 99.6594
R6605 gnd.n4004 gnd.n3751 99.6594
R6606 gnd.n4000 gnd.n3752 99.6594
R6607 gnd.n3996 gnd.n3753 99.6594
R6608 gnd.n3992 gnd.n3754 99.6594
R6609 gnd.n3988 gnd.n3755 99.6594
R6610 gnd.n3984 gnd.n3756 99.6594
R6611 gnd.n3980 gnd.n3757 99.6594
R6612 gnd.n3976 gnd.n3758 99.6594
R6613 gnd.n3972 gnd.n3759 99.6594
R6614 gnd.n3968 gnd.n3760 99.6594
R6615 gnd.n3964 gnd.n3761 99.6594
R6616 gnd.n3960 gnd.n3762 99.6594
R6617 gnd.n4072 gnd.n2272 99.6594
R6618 gnd.n3726 gnd.n2295 99.6594
R6619 gnd.n3724 gnd.n2294 99.6594
R6620 gnd.n3720 gnd.n2293 99.6594
R6621 gnd.n3716 gnd.n2292 99.6594
R6622 gnd.n3712 gnd.n2291 99.6594
R6623 gnd.n3708 gnd.n2290 99.6594
R6624 gnd.n3704 gnd.n2289 99.6594
R6625 gnd.n3636 gnd.n2288 99.6594
R6626 gnd.n2966 gnd.n2697 99.6594
R6627 gnd.n2723 gnd.n2704 99.6594
R6628 gnd.n2725 gnd.n2705 99.6594
R6629 gnd.n2733 gnd.n2706 99.6594
R6630 gnd.n2735 gnd.n2707 99.6594
R6631 gnd.n2743 gnd.n2708 99.6594
R6632 gnd.n2745 gnd.n2709 99.6594
R6633 gnd.n2753 gnd.n2710 99.6594
R6634 gnd.n276 gnd.n172 99.6594
R6635 gnd.n274 gnd.n273 99.6594
R6636 gnd.n269 gnd.n179 99.6594
R6637 gnd.n267 gnd.n266 99.6594
R6638 gnd.n262 gnd.n186 99.6594
R6639 gnd.n260 gnd.n259 99.6594
R6640 gnd.n255 gnd.n193 99.6594
R6641 gnd.n253 gnd.n252 99.6594
R6642 gnd.n198 gnd.n197 99.6594
R6643 gnd.n1560 gnd.n1476 99.6594
R6644 gnd.n1478 gnd.n1402 99.6594
R6645 gnd.n1479 gnd.n1409 99.6594
R6646 gnd.n1481 gnd.n1480 99.6594
R6647 gnd.n1483 gnd.n1418 99.6594
R6648 gnd.n1484 gnd.n1425 99.6594
R6649 gnd.n1486 gnd.n1485 99.6594
R6650 gnd.n1488 gnd.n1434 99.6594
R6651 gnd.n5654 gnd.n1443 99.6594
R6652 gnd.n3694 gnd.n2275 99.6594
R6653 gnd.n3690 gnd.n2276 99.6594
R6654 gnd.n3686 gnd.n2277 99.6594
R6655 gnd.n3682 gnd.n2278 99.6594
R6656 gnd.n3678 gnd.n2279 99.6594
R6657 gnd.n3674 gnd.n2280 99.6594
R6658 gnd.n3670 gnd.n2281 99.6594
R6659 gnd.n3666 gnd.n2282 99.6594
R6660 gnd.n3662 gnd.n2283 99.6594
R6661 gnd.n3658 gnd.n2284 99.6594
R6662 gnd.n3654 gnd.n2285 99.6594
R6663 gnd.n3650 gnd.n2286 99.6594
R6664 gnd.n3646 gnd.n2287 99.6594
R6665 gnd.n2881 gnd.n2880 99.6594
R6666 gnd.n2875 gnd.n2792 99.6594
R6667 gnd.n2872 gnd.n2793 99.6594
R6668 gnd.n2868 gnd.n2794 99.6594
R6669 gnd.n2864 gnd.n2795 99.6594
R6670 gnd.n2860 gnd.n2796 99.6594
R6671 gnd.n2856 gnd.n2797 99.6594
R6672 gnd.n2852 gnd.n2798 99.6594
R6673 gnd.n2848 gnd.n2799 99.6594
R6674 gnd.n2844 gnd.n2800 99.6594
R6675 gnd.n2840 gnd.n2801 99.6594
R6676 gnd.n2836 gnd.n2802 99.6594
R6677 gnd.n2883 gnd.n2791 99.6594
R6678 gnd.n4324 gnd.n1146 99.6594
R6679 gnd.n4326 gnd.n1147 99.6594
R6680 gnd.n4334 gnd.n1148 99.6594
R6681 gnd.n4344 gnd.n1149 99.6594
R6682 gnd.n4346 gnd.n1150 99.6594
R6683 gnd.n4354 gnd.n1151 99.6594
R6684 gnd.n4364 gnd.n1152 99.6594
R6685 gnd.n4367 gnd.n1153 99.6594
R6686 gnd.n4571 gnd.n1154 99.6594
R6687 gnd.n3950 gnd.n3763 99.6594
R6688 gnd.n3947 gnd.n3764 99.6594
R6689 gnd.n3943 gnd.n3765 99.6594
R6690 gnd.n3939 gnd.n3766 99.6594
R6691 gnd.n3935 gnd.n3767 99.6594
R6692 gnd.n3931 gnd.n3768 99.6594
R6693 gnd.n3927 gnd.n3769 99.6594
R6694 gnd.n3923 gnd.n3770 99.6594
R6695 gnd.n3919 gnd.n3771 99.6594
R6696 gnd.n3948 gnd.n3763 99.6594
R6697 gnd.n3944 gnd.n3764 99.6594
R6698 gnd.n3940 gnd.n3765 99.6594
R6699 gnd.n3936 gnd.n3766 99.6594
R6700 gnd.n3932 gnd.n3767 99.6594
R6701 gnd.n3928 gnd.n3768 99.6594
R6702 gnd.n3924 gnd.n3769 99.6594
R6703 gnd.n3920 gnd.n3770 99.6594
R6704 gnd.n3853 gnd.n3771 99.6594
R6705 gnd.n4366 gnd.n1154 99.6594
R6706 gnd.n4365 gnd.n1153 99.6594
R6707 gnd.n4355 gnd.n1152 99.6594
R6708 gnd.n4347 gnd.n1151 99.6594
R6709 gnd.n4345 gnd.n1150 99.6594
R6710 gnd.n4335 gnd.n1149 99.6594
R6711 gnd.n4327 gnd.n1148 99.6594
R6712 gnd.n4325 gnd.n1147 99.6594
R6713 gnd.n4315 gnd.n1146 99.6594
R6714 gnd.n2881 gnd.n2804 99.6594
R6715 gnd.n2873 gnd.n2792 99.6594
R6716 gnd.n2869 gnd.n2793 99.6594
R6717 gnd.n2865 gnd.n2794 99.6594
R6718 gnd.n2861 gnd.n2795 99.6594
R6719 gnd.n2857 gnd.n2796 99.6594
R6720 gnd.n2853 gnd.n2797 99.6594
R6721 gnd.n2849 gnd.n2798 99.6594
R6722 gnd.n2845 gnd.n2799 99.6594
R6723 gnd.n2841 gnd.n2800 99.6594
R6724 gnd.n2837 gnd.n2801 99.6594
R6725 gnd.n2833 gnd.n2802 99.6594
R6726 gnd.n2884 gnd.n2883 99.6594
R6727 gnd.n3649 gnd.n2287 99.6594
R6728 gnd.n3653 gnd.n2286 99.6594
R6729 gnd.n3657 gnd.n2285 99.6594
R6730 gnd.n3661 gnd.n2284 99.6594
R6731 gnd.n3665 gnd.n2283 99.6594
R6732 gnd.n3669 gnd.n2282 99.6594
R6733 gnd.n3673 gnd.n2281 99.6594
R6734 gnd.n3677 gnd.n2280 99.6594
R6735 gnd.n3681 gnd.n2279 99.6594
R6736 gnd.n3685 gnd.n2278 99.6594
R6737 gnd.n3689 gnd.n2277 99.6594
R6738 gnd.n3693 gnd.n2276 99.6594
R6739 gnd.n2316 gnd.n2275 99.6594
R6740 gnd.n1476 gnd.n1401 99.6594
R6741 gnd.n1478 gnd.n1477 99.6594
R6742 gnd.n1479 gnd.n1410 99.6594
R6743 gnd.n1481 gnd.n1417 99.6594
R6744 gnd.n1483 gnd.n1482 99.6594
R6745 gnd.n1484 gnd.n1426 99.6594
R6746 gnd.n1486 gnd.n1433 99.6594
R6747 gnd.n1488 gnd.n1487 99.6594
R6748 gnd.n5655 gnd.n5654 99.6594
R6749 gnd.n197 gnd.n194 99.6594
R6750 gnd.n254 gnd.n253 99.6594
R6751 gnd.n193 gnd.n187 99.6594
R6752 gnd.n261 gnd.n260 99.6594
R6753 gnd.n186 gnd.n180 99.6594
R6754 gnd.n268 gnd.n267 99.6594
R6755 gnd.n179 gnd.n173 99.6594
R6756 gnd.n275 gnd.n274 99.6594
R6757 gnd.n172 gnd.n169 99.6594
R6758 gnd.n2967 gnd.n2966 99.6594
R6759 gnd.n2726 gnd.n2704 99.6594
R6760 gnd.n2732 gnd.n2705 99.6594
R6761 gnd.n2736 gnd.n2706 99.6594
R6762 gnd.n2742 gnd.n2707 99.6594
R6763 gnd.n2746 gnd.n2708 99.6594
R6764 gnd.n2752 gnd.n2709 99.6594
R6765 gnd.n2710 gnd.n2694 99.6594
R6766 gnd.n3703 gnd.n2288 99.6594
R6767 gnd.n3707 gnd.n2289 99.6594
R6768 gnd.n3711 gnd.n2290 99.6594
R6769 gnd.n3715 gnd.n2291 99.6594
R6770 gnd.n3719 gnd.n2292 99.6594
R6771 gnd.n3723 gnd.n2293 99.6594
R6772 gnd.n3727 gnd.n2294 99.6594
R6773 gnd.n2297 gnd.n2295 99.6594
R6774 gnd.n4070 gnd.n3774 99.6594
R6775 gnd.n4062 gnd.n3736 99.6594
R6776 gnd.n4058 gnd.n3737 99.6594
R6777 gnd.n4054 gnd.n3738 99.6594
R6778 gnd.n4050 gnd.n3739 99.6594
R6779 gnd.n4046 gnd.n3740 99.6594
R6780 gnd.n4042 gnd.n3741 99.6594
R6781 gnd.n4038 gnd.n3742 99.6594
R6782 gnd.n4033 gnd.n3743 99.6594
R6783 gnd.n4029 gnd.n3744 99.6594
R6784 gnd.n4025 gnd.n3745 99.6594
R6785 gnd.n4021 gnd.n3746 99.6594
R6786 gnd.n4017 gnd.n3747 99.6594
R6787 gnd.n4013 gnd.n3748 99.6594
R6788 gnd.n4009 gnd.n3749 99.6594
R6789 gnd.n4005 gnd.n3750 99.6594
R6790 gnd.n4001 gnd.n3751 99.6594
R6791 gnd.n3997 gnd.n3752 99.6594
R6792 gnd.n3993 gnd.n3753 99.6594
R6793 gnd.n3989 gnd.n3754 99.6594
R6794 gnd.n3985 gnd.n3755 99.6594
R6795 gnd.n3981 gnd.n3756 99.6594
R6796 gnd.n3977 gnd.n3757 99.6594
R6797 gnd.n3973 gnd.n3758 99.6594
R6798 gnd.n3969 gnd.n3759 99.6594
R6799 gnd.n3965 gnd.n3760 99.6594
R6800 gnd.n3961 gnd.n3761 99.6594
R6801 gnd.n3957 gnd.n3762 99.6594
R6802 gnd.n4073 gnd.n4072 99.6594
R6803 gnd.n4430 gnd.n1156 99.6594
R6804 gnd.n4511 gnd.n1157 99.6594
R6805 gnd.n4509 gnd.n1158 99.6594
R6806 gnd.n4501 gnd.n1159 99.6594
R6807 gnd.n4499 gnd.n1160 99.6594
R6808 gnd.n4491 gnd.n1161 99.6594
R6809 gnd.n4489 gnd.n1162 99.6594
R6810 gnd.n4481 gnd.n1163 99.6594
R6811 gnd.n4479 gnd.n1164 99.6594
R6812 gnd.n4471 gnd.n1165 99.6594
R6813 gnd.n4443 gnd.n1166 99.6594
R6814 gnd.n4462 gnd.n1167 99.6594
R6815 gnd.n4460 gnd.n1168 99.6594
R6816 gnd.n4452 gnd.n1169 99.6594
R6817 gnd.n4450 gnd.n1170 99.6594
R6818 gnd.n5908 gnd.n1172 99.6594
R6819 gnd.n5912 gnd.n1173 99.6594
R6820 gnd.n5916 gnd.n1174 99.6594
R6821 gnd.n5920 gnd.n1175 99.6594
R6822 gnd.n5925 gnd.n1176 99.6594
R6823 gnd.n5929 gnd.n1177 99.6594
R6824 gnd.n5933 gnd.n1178 99.6594
R6825 gnd.n5937 gnd.n1179 99.6594
R6826 gnd.n5941 gnd.n1180 99.6594
R6827 gnd.n5945 gnd.n1181 99.6594
R6828 gnd.n5949 gnd.n1182 99.6594
R6829 gnd.n1184 gnd.n1183 99.6594
R6830 gnd.n5955 gnd.n1143 99.6594
R6831 gnd.n5652 gnd.n1491 99.6594
R6832 gnd.n5644 gnd.n1448 99.6594
R6833 gnd.n5640 gnd.n1449 99.6594
R6834 gnd.n5636 gnd.n1450 99.6594
R6835 gnd.n5632 gnd.n1451 99.6594
R6836 gnd.n5628 gnd.n1452 99.6594
R6837 gnd.n5624 gnd.n1453 99.6594
R6838 gnd.n5620 gnd.n1454 99.6594
R6839 gnd.n5615 gnd.n1455 99.6594
R6840 gnd.n5611 gnd.n1456 99.6594
R6841 gnd.n5607 gnd.n1457 99.6594
R6842 gnd.n5603 gnd.n1458 99.6594
R6843 gnd.n5598 gnd.n1460 99.6594
R6844 gnd.n5594 gnd.n1461 99.6594
R6845 gnd.n5590 gnd.n1462 99.6594
R6846 gnd.n5586 gnd.n1463 99.6594
R6847 gnd.n5582 gnd.n1464 99.6594
R6848 gnd.n5578 gnd.n1465 99.6594
R6849 gnd.n5574 gnd.n1466 99.6594
R6850 gnd.n5570 gnd.n1467 99.6594
R6851 gnd.n5566 gnd.n1468 99.6594
R6852 gnd.n5562 gnd.n1469 99.6594
R6853 gnd.n5558 gnd.n1470 99.6594
R6854 gnd.n5554 gnd.n1471 99.6594
R6855 gnd.n5550 gnd.n1472 99.6594
R6856 gnd.n5546 gnd.n1473 99.6594
R6857 gnd.n5542 gnd.n1474 99.6594
R6858 gnd.n5534 gnd.n1475 99.6594
R6859 gnd.n489 gnd.n488 99.6594
R6860 gnd.n480 gnd.n285 99.6594
R6861 gnd.n479 gnd.n478 99.6594
R6862 gnd.n470 gnd.n289 99.6594
R6863 gnd.n469 gnd.n468 99.6594
R6864 gnd.n460 gnd.n293 99.6594
R6865 gnd.n459 gnd.n458 99.6594
R6866 gnd.n450 gnd.n297 99.6594
R6867 gnd.n449 gnd.n448 99.6594
R6868 gnd.n440 gnd.n301 99.6594
R6869 gnd.n439 gnd.n438 99.6594
R6870 gnd.n430 gnd.n307 99.6594
R6871 gnd.n429 gnd.n428 99.6594
R6872 gnd.n420 gnd.n311 99.6594
R6873 gnd.n419 gnd.n418 99.6594
R6874 gnd.n410 gnd.n315 99.6594
R6875 gnd.n409 gnd.n408 99.6594
R6876 gnd.n400 gnd.n319 99.6594
R6877 gnd.n399 gnd.n398 99.6594
R6878 gnd.n390 gnd.n323 99.6594
R6879 gnd.n389 gnd.n388 99.6594
R6880 gnd.n380 gnd.n379 99.6594
R6881 gnd.n378 gnd.n377 99.6594
R6882 gnd.n369 gnd.n333 99.6594
R6883 gnd.n368 gnd.n367 99.6594
R6884 gnd.n359 gnd.n337 99.6594
R6885 gnd.n358 gnd.n357 99.6594
R6886 gnd.n349 gnd.n341 99.6594
R6887 gnd.n348 gnd.n347 99.6594
R6888 gnd.n4298 gnd.n2104 99.6594
R6889 gnd.n4302 gnd.n2105 99.6594
R6890 gnd.n4275 gnd.n2106 99.6594
R6891 gnd.n4310 gnd.n2107 99.6594
R6892 gnd.n4312 gnd.n2108 99.6594
R6893 gnd.n4319 gnd.n2109 99.6594
R6894 gnd.n4321 gnd.n2110 99.6594
R6895 gnd.n4331 gnd.n2111 99.6594
R6896 gnd.n4339 gnd.n2112 99.6594
R6897 gnd.n4341 gnd.n2113 99.6594
R6898 gnd.n4351 gnd.n2114 99.6594
R6899 gnd.n4359 gnd.n2115 99.6594
R6900 gnd.n4361 gnd.n2116 99.6594
R6901 gnd.n4373 gnd.n2117 99.6594
R6902 gnd.n4301 gnd.n2104 99.6594
R6903 gnd.n4274 gnd.n2105 99.6594
R6904 gnd.n4309 gnd.n2106 99.6594
R6905 gnd.n4311 gnd.n2107 99.6594
R6906 gnd.n4318 gnd.n2108 99.6594
R6907 gnd.n4320 gnd.n2109 99.6594
R6908 gnd.n4330 gnd.n2110 99.6594
R6909 gnd.n4338 gnd.n2111 99.6594
R6910 gnd.n4340 gnd.n2112 99.6594
R6911 gnd.n4350 gnd.n2113 99.6594
R6912 gnd.n4358 gnd.n2114 99.6594
R6913 gnd.n4360 gnd.n2115 99.6594
R6914 gnd.n4372 gnd.n2116 99.6594
R6915 gnd.n2118 gnd.n2117 99.6594
R6916 gnd.n1640 gnd.n1382 99.6594
R6917 gnd.n1642 gnd.n1387 99.6594
R6918 gnd.n1643 gnd.n1390 99.6594
R6919 gnd.n1645 gnd.n1392 99.6594
R6920 gnd.n1646 gnd.n1396 99.6594
R6921 gnd.n1648 gnd.n1647 99.6594
R6922 gnd.n1650 gnd.n1406 99.6594
R6923 gnd.n1651 gnd.n1413 99.6594
R6924 gnd.n1653 gnd.n1652 99.6594
R6925 gnd.n1655 gnd.n1422 99.6594
R6926 gnd.n1656 gnd.n1429 99.6594
R6927 gnd.n1658 gnd.n1657 99.6594
R6928 gnd.n1661 gnd.n1438 99.6594
R6929 gnd.n5427 gnd.n1639 99.6594
R6930 gnd.n1658 gnd.n1437 99.6594
R6931 gnd.n1656 gnd.n1430 99.6594
R6932 gnd.n1655 gnd.n1654 99.6594
R6933 gnd.n1653 gnd.n1421 99.6594
R6934 gnd.n1651 gnd.n1414 99.6594
R6935 gnd.n1650 gnd.n1649 99.6594
R6936 gnd.n1648 gnd.n1405 99.6594
R6937 gnd.n1646 gnd.n1397 99.6594
R6938 gnd.n1645 gnd.n1644 99.6594
R6939 gnd.n1643 gnd.n1391 99.6594
R6940 gnd.n1642 gnd.n1641 99.6594
R6941 gnd.n1640 gnd.n1386 99.6594
R6942 gnd.n5428 gnd.n5427 99.6594
R6943 gnd.n1661 gnd.n1660 99.6594
R6944 gnd.n4369 gnd.t272 98.63
R6945 gnd.n5656 gnd.t293 98.63
R6946 gnd.n2122 gnd.t315 98.63
R6947 gnd.n1511 gnd.t290 98.63
R6948 gnd.n1534 gnd.t281 98.63
R6949 gnd.n5536 gnd.t221 98.63
R6950 gnd.n282 gnd.t227 98.63
R6951 gnd.n304 gnd.t216 98.63
R6952 gnd.n326 gnd.t283 98.63
R6953 gnd.n200 gnd.t305 98.63
R6954 gnd.n3793 gnd.t258 98.63
R6955 gnd.n3815 gnd.t238 98.63
R6956 gnd.n3836 gnd.t261 98.63
R6957 gnd.n3854 gnd.t210 98.63
R6958 gnd.n1201 gnd.t308 98.63
R6959 gnd.n4428 gnd.t241 98.63
R6960 gnd.n4441 gnd.t267 98.63
R6961 gnd.n1439 gnd.t245 98.63
R6962 gnd.n4674 gnd.t300 92.8196
R6963 gnd.n1762 gnd.t234 92.8196
R6964 gnd.n5837 gnd.t225 92.8118
R6965 gnd.n1756 gnd.t286 92.8118
R6966 gnd.n1263 gnd.n1262 81.8399
R6967 gnd.n2755 gnd.t264 74.8376
R6968 gnd.n2313 gnd.t297 74.8376
R6969 gnd.n4675 gnd.t299 72.8438
R6970 gnd.n1763 gnd.t235 72.8438
R6971 gnd.n1264 gnd.n1257 72.8411
R6972 gnd.n1270 gnd.n1255 72.8411
R6973 gnd.n1731 gnd.n1730 72.8411
R6974 gnd.n4370 gnd.t271 72.836
R6975 gnd.n5838 gnd.t224 72.836
R6976 gnd.n1757 gnd.t287 72.836
R6977 gnd.n5657 gnd.t292 72.836
R6978 gnd.n2123 gnd.t316 72.836
R6979 gnd.n1512 gnd.t289 72.836
R6980 gnd.n1535 gnd.t280 72.836
R6981 gnd.n5537 gnd.t220 72.836
R6982 gnd.n283 gnd.t228 72.836
R6983 gnd.n305 gnd.t217 72.836
R6984 gnd.n327 gnd.t284 72.836
R6985 gnd.n201 gnd.t306 72.836
R6986 gnd.n3794 gnd.t257 72.836
R6987 gnd.n3816 gnd.t237 72.836
R6988 gnd.n3837 gnd.t260 72.836
R6989 gnd.n3855 gnd.t209 72.836
R6990 gnd.n1202 gnd.t309 72.836
R6991 gnd.n4429 gnd.t242 72.836
R6992 gnd.n4442 gnd.t268 72.836
R6993 gnd.n1440 gnd.t246 72.836
R6994 gnd.n5343 gnd.n5342 71.676
R6995 gnd.n5340 gnd.n5339 71.676
R6996 gnd.n5335 gnd.n1739 71.676
R6997 gnd.n5333 gnd.n5332 71.676
R6998 gnd.n5328 gnd.n1742 71.676
R6999 gnd.n5326 gnd.n5325 71.676
R7000 gnd.n5321 gnd.n1745 71.676
R7001 gnd.n5319 gnd.n5318 71.676
R7002 gnd.n5314 gnd.n1748 71.676
R7003 gnd.n5312 gnd.n5311 71.676
R7004 gnd.n5307 gnd.n1751 71.676
R7005 gnd.n5305 gnd.n5304 71.676
R7006 gnd.n5300 gnd.n1754 71.676
R7007 gnd.n5298 gnd.n5297 71.676
R7008 gnd.n5292 gnd.n1759 71.676
R7009 gnd.n5290 gnd.n5289 71.676
R7010 gnd.n5285 gnd.n5284 71.676
R7011 gnd.n5282 gnd.n5281 71.676
R7012 gnd.n5276 gnd.n1765 71.676
R7013 gnd.n5274 gnd.n5273 71.676
R7014 gnd.n5269 gnd.n1768 71.676
R7015 gnd.n5267 gnd.n5266 71.676
R7016 gnd.n5262 gnd.n1771 71.676
R7017 gnd.n5260 gnd.n5259 71.676
R7018 gnd.n5255 gnd.n1774 71.676
R7019 gnd.n5253 gnd.n5252 71.676
R7020 gnd.n5248 gnd.n1777 71.676
R7021 gnd.n5246 gnd.n5245 71.676
R7022 gnd.n5241 gnd.n1780 71.676
R7023 gnd.n5239 gnd.n5238 71.676
R7024 gnd.n5234 gnd.n1783 71.676
R7025 gnd.n5232 gnd.n5231 71.676
R7026 gnd.n5227 gnd.n5225 71.676
R7027 gnd.n5901 gnd.n5900 71.676
R7028 gnd.n5895 gnd.n1219 71.676
R7029 gnd.n5892 gnd.n1220 71.676
R7030 gnd.n5888 gnd.n1221 71.676
R7031 gnd.n5884 gnd.n1222 71.676
R7032 gnd.n5880 gnd.n1223 71.676
R7033 gnd.n5876 gnd.n1224 71.676
R7034 gnd.n5872 gnd.n1225 71.676
R7035 gnd.n5868 gnd.n1226 71.676
R7036 gnd.n5864 gnd.n1227 71.676
R7037 gnd.n5860 gnd.n1228 71.676
R7038 gnd.n5856 gnd.n1229 71.676
R7039 gnd.n5852 gnd.n1230 71.676
R7040 gnd.n5848 gnd.n1231 71.676
R7041 gnd.n5844 gnd.n1232 71.676
R7042 gnd.n5840 gnd.n1233 71.676
R7043 gnd.n1234 gnd.n1217 71.676
R7044 gnd.n4678 gnd.n1235 71.676
R7045 gnd.n4683 gnd.n1236 71.676
R7046 gnd.n4687 gnd.n1237 71.676
R7047 gnd.n4691 gnd.n1238 71.676
R7048 gnd.n4695 gnd.n1239 71.676
R7049 gnd.n4699 gnd.n1240 71.676
R7050 gnd.n4703 gnd.n1241 71.676
R7051 gnd.n4707 gnd.n1242 71.676
R7052 gnd.n4711 gnd.n1243 71.676
R7053 gnd.n4715 gnd.n1244 71.676
R7054 gnd.n4719 gnd.n1245 71.676
R7055 gnd.n4723 gnd.n1246 71.676
R7056 gnd.n4727 gnd.n1247 71.676
R7057 gnd.n4731 gnd.n1248 71.676
R7058 gnd.n4735 gnd.n1249 71.676
R7059 gnd.n5901 gnd.n1252 71.676
R7060 gnd.n5893 gnd.n1219 71.676
R7061 gnd.n5889 gnd.n1220 71.676
R7062 gnd.n5885 gnd.n1221 71.676
R7063 gnd.n5881 gnd.n1222 71.676
R7064 gnd.n5877 gnd.n1223 71.676
R7065 gnd.n5873 gnd.n1224 71.676
R7066 gnd.n5869 gnd.n1225 71.676
R7067 gnd.n5865 gnd.n1226 71.676
R7068 gnd.n5861 gnd.n1227 71.676
R7069 gnd.n5857 gnd.n1228 71.676
R7070 gnd.n5853 gnd.n1229 71.676
R7071 gnd.n5849 gnd.n1230 71.676
R7072 gnd.n5845 gnd.n1231 71.676
R7073 gnd.n5841 gnd.n1232 71.676
R7074 gnd.n5904 gnd.n5903 71.676
R7075 gnd.n4677 gnd.n1234 71.676
R7076 gnd.n4682 gnd.n1235 71.676
R7077 gnd.n4686 gnd.n1236 71.676
R7078 gnd.n4690 gnd.n1237 71.676
R7079 gnd.n4694 gnd.n1238 71.676
R7080 gnd.n4698 gnd.n1239 71.676
R7081 gnd.n4702 gnd.n1240 71.676
R7082 gnd.n4706 gnd.n1241 71.676
R7083 gnd.n4710 gnd.n1242 71.676
R7084 gnd.n4714 gnd.n1243 71.676
R7085 gnd.n4718 gnd.n1244 71.676
R7086 gnd.n4722 gnd.n1245 71.676
R7087 gnd.n4726 gnd.n1246 71.676
R7088 gnd.n4730 gnd.n1247 71.676
R7089 gnd.n4734 gnd.n1248 71.676
R7090 gnd.n4738 gnd.n1249 71.676
R7091 gnd.n5225 gnd.n1784 71.676
R7092 gnd.n5233 gnd.n5232 71.676
R7093 gnd.n1783 gnd.n1781 71.676
R7094 gnd.n5240 gnd.n5239 71.676
R7095 gnd.n1780 gnd.n1778 71.676
R7096 gnd.n5247 gnd.n5246 71.676
R7097 gnd.n1777 gnd.n1775 71.676
R7098 gnd.n5254 gnd.n5253 71.676
R7099 gnd.n1774 gnd.n1772 71.676
R7100 gnd.n5261 gnd.n5260 71.676
R7101 gnd.n1771 gnd.n1769 71.676
R7102 gnd.n5268 gnd.n5267 71.676
R7103 gnd.n1768 gnd.n1766 71.676
R7104 gnd.n5275 gnd.n5274 71.676
R7105 gnd.n1765 gnd.n1761 71.676
R7106 gnd.n5283 gnd.n5282 71.676
R7107 gnd.n5287 gnd.n5286 71.676
R7108 gnd.n5291 gnd.n5290 71.676
R7109 gnd.n1759 gnd.n1755 71.676
R7110 gnd.n5299 gnd.n5298 71.676
R7111 gnd.n1754 gnd.n1752 71.676
R7112 gnd.n5306 gnd.n5305 71.676
R7113 gnd.n1751 gnd.n1749 71.676
R7114 gnd.n5313 gnd.n5312 71.676
R7115 gnd.n1748 gnd.n1746 71.676
R7116 gnd.n5320 gnd.n5319 71.676
R7117 gnd.n1745 gnd.n1743 71.676
R7118 gnd.n5327 gnd.n5326 71.676
R7119 gnd.n1742 gnd.n1740 71.676
R7120 gnd.n5334 gnd.n5333 71.676
R7121 gnd.n1739 gnd.n1737 71.676
R7122 gnd.n5341 gnd.n5340 71.676
R7123 gnd.n5344 gnd.n5343 71.676
R7124 gnd.n8 gnd.t193 69.1507
R7125 gnd.n14 gnd.t40 68.4792
R7126 gnd.n13 gnd.t64 68.4792
R7127 gnd.n12 gnd.t203 68.4792
R7128 gnd.n11 gnd.t54 68.4792
R7129 gnd.n10 gnd.t197 68.4792
R7130 gnd.n9 gnd.t195 68.4792
R7131 gnd.n8 gnd.t44 68.4792
R7132 gnd.n2882 gnd.n2786 64.369
R7133 gnd.n6712 gnd.n136 64.0315
R7134 gnd.n4071 gnd.n2260 63.0944
R7135 gnd.n6841 gnd.n165 63.0944
R7136 gnd.n4680 gnd.n4675 59.5399
R7137 gnd.n5278 gnd.n1763 59.5399
R7138 gnd.n5839 gnd.n5838 59.5399
R7139 gnd.n5294 gnd.n1757 59.5399
R7140 gnd.n5836 gnd.n1273 59.1804
R7141 gnd.n3735 gnd.n2273 57.3586
R7142 gnd.n2541 gnd.t125 56.407
R7143 gnd.n2506 gnd.t173 56.407
R7144 gnd.n2517 gnd.t84 56.407
R7145 gnd.n2529 gnd.t164 56.407
R7146 gnd.n52 gnd.t102 56.407
R7147 gnd.n17 gnd.t91 56.407
R7148 gnd.n28 gnd.t183 56.407
R7149 gnd.n40 gnd.t139 56.407
R7150 gnd.n2550 gnd.t150 55.8337
R7151 gnd.n2515 gnd.t80 55.8337
R7152 gnd.n2526 gnd.t181 55.8337
R7153 gnd.n2538 gnd.t86 55.8337
R7154 gnd.n61 gnd.t123 55.8337
R7155 gnd.n26 gnd.t115 55.8337
R7156 gnd.n37 gnd.t165 55.8337
R7157 gnd.n49 gnd.t162 55.8337
R7158 gnd.n1261 gnd.n1260 54.358
R7159 gnd.n1728 gnd.n1727 54.358
R7160 gnd.n2541 gnd.n2540 53.0052
R7161 gnd.n2543 gnd.n2542 53.0052
R7162 gnd.n2545 gnd.n2544 53.0052
R7163 gnd.n2547 gnd.n2546 53.0052
R7164 gnd.n2549 gnd.n2548 53.0052
R7165 gnd.n2506 gnd.n2505 53.0052
R7166 gnd.n2508 gnd.n2507 53.0052
R7167 gnd.n2510 gnd.n2509 53.0052
R7168 gnd.n2512 gnd.n2511 53.0052
R7169 gnd.n2514 gnd.n2513 53.0052
R7170 gnd.n2517 gnd.n2516 53.0052
R7171 gnd.n2519 gnd.n2518 53.0052
R7172 gnd.n2521 gnd.n2520 53.0052
R7173 gnd.n2523 gnd.n2522 53.0052
R7174 gnd.n2525 gnd.n2524 53.0052
R7175 gnd.n2529 gnd.n2528 53.0052
R7176 gnd.n2531 gnd.n2530 53.0052
R7177 gnd.n2533 gnd.n2532 53.0052
R7178 gnd.n2535 gnd.n2534 53.0052
R7179 gnd.n2537 gnd.n2536 53.0052
R7180 gnd.n60 gnd.n59 53.0052
R7181 gnd.n58 gnd.n57 53.0052
R7182 gnd.n56 gnd.n55 53.0052
R7183 gnd.n54 gnd.n53 53.0052
R7184 gnd.n52 gnd.n51 53.0052
R7185 gnd.n25 gnd.n24 53.0052
R7186 gnd.n23 gnd.n22 53.0052
R7187 gnd.n21 gnd.n20 53.0052
R7188 gnd.n19 gnd.n18 53.0052
R7189 gnd.n17 gnd.n16 53.0052
R7190 gnd.n36 gnd.n35 53.0052
R7191 gnd.n34 gnd.n33 53.0052
R7192 gnd.n32 gnd.n31 53.0052
R7193 gnd.n30 gnd.n29 53.0052
R7194 gnd.n28 gnd.n27 53.0052
R7195 gnd.n48 gnd.n47 53.0052
R7196 gnd.n46 gnd.n45 53.0052
R7197 gnd.n44 gnd.n43 53.0052
R7198 gnd.n42 gnd.n41 53.0052
R7199 gnd.n40 gnd.n39 53.0052
R7200 gnd.n1719 gnd.n1718 52.4801
R7201 gnd.n3587 gnd.t57 52.3082
R7202 gnd.n3555 gnd.t50 52.3082
R7203 gnd.n3523 gnd.t46 52.3082
R7204 gnd.n3492 gnd.t30 52.3082
R7205 gnd.n3460 gnd.t42 52.3082
R7206 gnd.n3428 gnd.t189 52.3082
R7207 gnd.n3396 gnd.t199 52.3082
R7208 gnd.n3365 gnd.t66 52.3082
R7209 gnd.n3417 gnd.n3385 51.4173
R7210 gnd.n3481 gnd.n3480 50.455
R7211 gnd.n3449 gnd.n3448 50.455
R7212 gnd.n3417 gnd.n3416 50.455
R7213 gnd.n2829 gnd.n2828 45.1884
R7214 gnd.n2339 gnd.n2338 45.1884
R7215 gnd.n5346 gnd.n1734 44.3322
R7216 gnd.n1264 gnd.n1263 44.3189
R7217 gnd.n4371 gnd.n4370 42.2793
R7218 gnd.n5658 gnd.n5657 42.2793
R7219 gnd.n2830 gnd.n2829 42.2793
R7220 gnd.n2340 gnd.n2339 42.2793
R7221 gnd.n2756 gnd.n2755 42.2793
R7222 gnd.n3702 gnd.n2313 42.2793
R7223 gnd.n2124 gnd.n2123 42.2793
R7224 gnd.n5617 gnd.n1512 42.2793
R7225 gnd.n5580 gnd.n1535 42.2793
R7226 gnd.n5540 gnd.n5537 42.2793
R7227 gnd.n284 gnd.n283 42.2793
R7228 gnd.n306 gnd.n305 42.2793
R7229 gnd.n328 gnd.n327 42.2793
R7230 gnd.n250 gnd.n201 42.2793
R7231 gnd.n4035 gnd.n3794 42.2793
R7232 gnd.n3995 gnd.n3816 42.2793
R7233 gnd.n3956 gnd.n3837 42.2793
R7234 gnd.n3856 gnd.n3855 42.2793
R7235 gnd.n5923 gnd.n1202 42.2793
R7236 gnd.n4519 gnd.n4429 42.2793
R7237 gnd.n4470 gnd.n4442 42.2793
R7238 gnd.n1441 gnd.n1440 42.2793
R7239 gnd.n1262 gnd.n1261 41.6274
R7240 gnd.n1729 gnd.n1728 41.6274
R7241 gnd.n1271 gnd.n1270 40.8975
R7242 gnd.n1732 gnd.n1731 40.8975
R7243 gnd.n1270 gnd.n1269 35.055
R7244 gnd.n1265 gnd.n1264 35.055
R7245 gnd.n1721 gnd.n1720 35.055
R7246 gnd.n1731 gnd.n1717 35.055
R7247 gnd.n6181 gnd.n6180 34.6735
R7248 gnd.n6180 gnd.n6179 34.6735
R7249 gnd.n6179 gnd.n884 34.6735
R7250 gnd.n6173 gnd.n884 34.6735
R7251 gnd.n6173 gnd.n6172 34.6735
R7252 gnd.n6172 gnd.n6171 34.6735
R7253 gnd.n6171 gnd.n891 34.6735
R7254 gnd.n6165 gnd.n891 34.6735
R7255 gnd.n6165 gnd.n6164 34.6735
R7256 gnd.n6164 gnd.n6163 34.6735
R7257 gnd.n6163 gnd.n899 34.6735
R7258 gnd.n6157 gnd.n899 34.6735
R7259 gnd.n6157 gnd.n6156 34.6735
R7260 gnd.n6156 gnd.n6155 34.6735
R7261 gnd.n6155 gnd.n907 34.6735
R7262 gnd.n6149 gnd.n907 34.6735
R7263 gnd.n6149 gnd.n6148 34.6735
R7264 gnd.n6148 gnd.n6147 34.6735
R7265 gnd.n6147 gnd.n915 34.6735
R7266 gnd.n6141 gnd.n915 34.6735
R7267 gnd.n6141 gnd.n6140 34.6735
R7268 gnd.n6140 gnd.n6139 34.6735
R7269 gnd.n6139 gnd.n923 34.6735
R7270 gnd.n6133 gnd.n923 34.6735
R7271 gnd.n6133 gnd.n6132 34.6735
R7272 gnd.n6132 gnd.n6131 34.6735
R7273 gnd.n6131 gnd.n931 34.6735
R7274 gnd.n6125 gnd.n931 34.6735
R7275 gnd.n6125 gnd.n6124 34.6735
R7276 gnd.n6124 gnd.n6123 34.6735
R7277 gnd.n6123 gnd.n939 34.6735
R7278 gnd.n6117 gnd.n939 34.6735
R7279 gnd.n6117 gnd.n6116 34.6735
R7280 gnd.n6116 gnd.n6115 34.6735
R7281 gnd.n6115 gnd.n947 34.6735
R7282 gnd.n6109 gnd.n947 34.6735
R7283 gnd.n6109 gnd.n6108 34.6735
R7284 gnd.n6108 gnd.n6107 34.6735
R7285 gnd.n6107 gnd.n955 34.6735
R7286 gnd.n6101 gnd.n955 34.6735
R7287 gnd.n6101 gnd.n6100 34.6735
R7288 gnd.n6100 gnd.n6099 34.6735
R7289 gnd.n6099 gnd.n963 34.6735
R7290 gnd.n6093 gnd.n963 34.6735
R7291 gnd.n6093 gnd.n6092 34.6735
R7292 gnd.n6092 gnd.n6091 34.6735
R7293 gnd.n6091 gnd.n971 34.6735
R7294 gnd.n6085 gnd.n971 34.6735
R7295 gnd.n6085 gnd.n6084 34.6735
R7296 gnd.n6084 gnd.n6083 34.6735
R7297 gnd.n6083 gnd.n979 34.6735
R7298 gnd.n6077 gnd.n979 34.6735
R7299 gnd.n6077 gnd.n6076 34.6735
R7300 gnd.n6076 gnd.n6075 34.6735
R7301 gnd.n6075 gnd.n987 34.6735
R7302 gnd.n6069 gnd.n987 34.6735
R7303 gnd.n6069 gnd.n6068 34.6735
R7304 gnd.n6068 gnd.n6067 34.6735
R7305 gnd.n6067 gnd.n995 34.6735
R7306 gnd.n6061 gnd.n995 34.6735
R7307 gnd.n6061 gnd.n6060 34.6735
R7308 gnd.n6060 gnd.n6059 34.6735
R7309 gnd.n6059 gnd.n1003 34.6735
R7310 gnd.n6053 gnd.n1003 34.6735
R7311 gnd.n6053 gnd.n6052 34.6735
R7312 gnd.n6052 gnd.n6051 34.6735
R7313 gnd.n6051 gnd.n1011 34.6735
R7314 gnd.n6045 gnd.n1011 34.6735
R7315 gnd.n6045 gnd.n6044 34.6735
R7316 gnd.n6044 gnd.n6043 34.6735
R7317 gnd.n6043 gnd.n1019 34.6735
R7318 gnd.n6037 gnd.n1019 34.6735
R7319 gnd.n6037 gnd.n6036 34.6735
R7320 gnd.n6036 gnd.n6035 34.6735
R7321 gnd.n6035 gnd.n1027 34.6735
R7322 gnd.n6029 gnd.n1027 34.6735
R7323 gnd.n6029 gnd.n6028 34.6735
R7324 gnd.n6028 gnd.n6027 34.6735
R7325 gnd.n6027 gnd.n1035 34.6735
R7326 gnd.n6021 gnd.n1035 34.6735
R7327 gnd.n6021 gnd.n6020 34.6735
R7328 gnd.n6020 gnd.n6019 34.6735
R7329 gnd.n6019 gnd.n1043 34.6735
R7330 gnd.n2892 gnd.n2786 31.8661
R7331 gnd.n2892 gnd.n2891 31.8661
R7332 gnd.n2900 gnd.n2775 31.8661
R7333 gnd.n2908 gnd.n2775 31.8661
R7334 gnd.n2908 gnd.n2769 31.8661
R7335 gnd.n2916 gnd.n2769 31.8661
R7336 gnd.n2916 gnd.n2762 31.8661
R7337 gnd.n2954 gnd.n2762 31.8661
R7338 gnd.n2964 gnd.n2695 31.8661
R7339 gnd.n4081 gnd.n2260 31.8661
R7340 gnd.n4089 gnd.n2252 31.8661
R7341 gnd.n4089 gnd.n2241 31.8661
R7342 gnd.n4101 gnd.n2241 31.8661
R7343 gnd.n4101 gnd.n2244 31.8661
R7344 gnd.n4109 gnd.n2224 31.8661
R7345 gnd.n4121 gnd.n2224 31.8661
R7346 gnd.n4129 gnd.n2216 31.8661
R7347 gnd.n4141 gnd.n2205 31.8661
R7348 gnd.n4141 gnd.n2208 31.8661
R7349 gnd.n4150 gnd.n2188 31.8661
R7350 gnd.n4162 gnd.n2188 31.8661
R7351 gnd.n4170 gnd.n2182 31.8661
R7352 gnd.n4189 gnd.n2169 31.8661
R7353 gnd.n4189 gnd.n2172 31.8661
R7354 gnd.n4197 gnd.n1050 31.8661
R7355 gnd.n4568 gnd.n1144 31.8661
R7356 gnd.n2103 gnd.n1155 31.8661
R7357 gnd.n4579 gnd.n2103 31.8661
R7358 gnd.n4580 gnd.n4579 31.8661
R7359 gnd.n4580 gnd.n2096 31.8661
R7360 gnd.n4588 gnd.n2096 31.8661
R7361 gnd.n4596 gnd.n2089 31.8661
R7362 gnd.n4596 gnd.n2081 31.8661
R7363 gnd.n4604 gnd.n2081 31.8661
R7364 gnd.n4604 gnd.n2083 31.8661
R7365 gnd.n4629 gnd.n2064 31.8661
R7366 gnd.n4646 gnd.n2064 31.8661
R7367 gnd.n4646 gnd.n2065 31.8661
R7368 gnd.n5367 gnd.n1688 31.8661
R7369 gnd.n5375 gnd.n1688 31.8661
R7370 gnd.n5375 gnd.n1689 31.8661
R7371 gnd.n5383 gnd.n1676 31.8661
R7372 gnd.n5394 gnd.n1676 31.8661
R7373 gnd.n5394 gnd.n1669 31.8661
R7374 gnd.n5402 gnd.n1669 31.8661
R7375 gnd.n5721 gnd.n1378 31.8661
R7376 gnd.n5721 gnd.n1380 31.8661
R7377 gnd.n5426 gnd.n1380 31.8661
R7378 gnd.n5426 gnd.n1662 31.8661
R7379 gnd.n1662 gnd.n1447 31.8661
R7380 gnd.n1557 gnd.n1489 31.8661
R7381 gnd.n6782 gnd.n509 31.8661
R7382 gnd.n6790 gnd.n499 31.8661
R7383 gnd.n6799 gnd.n499 31.8661
R7384 gnd.n6897 gnd.n70 31.8661
R7385 gnd.n6889 gnd.n85 31.8661
R7386 gnd.n6889 gnd.n88 31.8661
R7387 gnd.n6883 gnd.n99 31.8661
R7388 gnd.n6877 gnd.n99 31.8661
R7389 gnd.n6871 gnd.n114 31.8661
R7390 gnd.n6865 gnd.n124 31.8661
R7391 gnd.n6865 gnd.n127 31.8661
R7392 gnd.n6853 gnd.n144 31.8661
R7393 gnd.n6853 gnd.n147 31.8661
R7394 gnd.n6847 gnd.n147 31.8661
R7395 gnd.n6841 gnd.n162 31.8661
R7396 gnd.t98 gnd.n2182 31.5474
R7397 gnd.t72 gnd.n70 31.5474
R7398 gnd.t116 gnd.n2216 30.9101
R7399 gnd.n2065 gnd.t192 30.9101
R7400 gnd.n5367 gnd.t190 30.9101
R7401 gnd.n6871 gnd.t75 30.9101
R7402 gnd.n5228 gnd.n5224 30.7517
R7403 gnd.n4741 gnd.n4737 30.7517
R7404 gnd.n6859 gnd.n136 28.6795
R7405 gnd.n5956 gnd.n1155 27.4049
R7406 gnd.n5653 gnd.n1447 27.4049
R7407 gnd.n6012 gnd.n1053 26.7676
R7408 gnd.n4206 gnd.n1062 26.7676
R7409 gnd.n4225 gnd.n1073 26.7676
R7410 gnd.n6000 gnd.n1076 26.7676
R7411 gnd.n5994 gnd.n1087 26.7676
R7412 gnd.n4252 gnd.n4251 26.7676
R7413 gnd.n5988 gnd.n1096 26.7676
R7414 gnd.n4260 gnd.n1104 26.7676
R7415 gnd.n4542 gnd.n1113 26.7676
R7416 gnd.n5976 gnd.n1116 26.7676
R7417 gnd.n4267 gnd.n1124 26.7676
R7418 gnd.n5970 gnd.n1127 26.7676
R7419 gnd.n5964 gnd.n1137 26.7676
R7420 gnd.n4569 gnd.n4568 26.7676
R7421 gnd.n5532 gnd.n1557 26.7676
R7422 gnd.n5470 gnd.n1559 26.7676
R7423 gnd.n5435 gnd.n1568 26.7676
R7424 gnd.n5518 gnd.n1581 26.7676
R7425 gnd.n5441 gnd.n1584 26.7676
R7426 gnd.n5512 gnd.n1594 26.7676
R7427 gnd.n5506 gnd.n1606 26.7676
R7428 gnd.n5499 gnd.n1609 26.7676
R7429 gnd.n5498 gnd.n1622 26.7676
R7430 gnd.n6736 gnd.n546 26.7676
R7431 gnd.n6747 gnd.n536 26.7676
R7432 gnd.n6729 gnd.n538 26.7676
R7433 gnd.n6769 gnd.n522 26.7676
R7434 gnd.n6774 gnd.n517 26.7676
R7435 gnd.n4370 gnd.n4369 25.7944
R7436 gnd.n5657 gnd.n5656 25.7944
R7437 gnd.n2755 gnd.n2754 25.7944
R7438 gnd.n2313 gnd.n2312 25.7944
R7439 gnd.n2123 gnd.n2122 25.7944
R7440 gnd.n1512 gnd.n1511 25.7944
R7441 gnd.n1535 gnd.n1534 25.7944
R7442 gnd.n5537 gnd.n5536 25.7944
R7443 gnd.n283 gnd.n282 25.7944
R7444 gnd.n305 gnd.n304 25.7944
R7445 gnd.n327 gnd.n326 25.7944
R7446 gnd.n201 gnd.n200 25.7944
R7447 gnd.n3794 gnd.n3793 25.7944
R7448 gnd.n3816 gnd.n3815 25.7944
R7449 gnd.n3837 gnd.n3836 25.7944
R7450 gnd.n3855 gnd.n3854 25.7944
R7451 gnd.n1202 gnd.n1201 25.7944
R7452 gnd.n4429 gnd.n4428 25.7944
R7453 gnd.n4442 gnd.n4441 25.7944
R7454 gnd.n1440 gnd.n1439 25.7944
R7455 gnd.n2976 gnd.n2696 24.8557
R7456 gnd.n2986 gnd.n2679 24.8557
R7457 gnd.n2682 gnd.n2670 24.8557
R7458 gnd.n3007 gnd.n2671 24.8557
R7459 gnd.n3017 gnd.n2651 24.8557
R7460 gnd.n3027 gnd.n3026 24.8557
R7461 gnd.n2637 gnd.n2635 24.8557
R7462 gnd.n3058 gnd.n3057 24.8557
R7463 gnd.n3073 gnd.n2620 24.8557
R7464 gnd.n3127 gnd.n2559 24.8557
R7465 gnd.n3083 gnd.n2560 24.8557
R7466 gnd.n3120 gnd.n2571 24.8557
R7467 gnd.n2609 gnd.n2608 24.8557
R7468 gnd.n3114 gnd.n3113 24.8557
R7469 gnd.n2595 gnd.n2582 24.8557
R7470 gnd.n3153 gnd.n3152 24.8557
R7471 gnd.n3163 gnd.n2491 24.8557
R7472 gnd.n3175 gnd.n2483 24.8557
R7473 gnd.n3174 gnd.n2471 24.8557
R7474 gnd.n3193 gnd.n3192 24.8557
R7475 gnd.n3203 gnd.n2464 24.8557
R7476 gnd.n3214 gnd.n2452 24.8557
R7477 gnd.n3238 gnd.n3237 24.8557
R7478 gnd.n3249 gnd.n2435 24.8557
R7479 gnd.n3248 gnd.n2437 24.8557
R7480 gnd.n3260 gnd.n2428 24.8557
R7481 gnd.n3278 gnd.n3277 24.8557
R7482 gnd.n2419 gnd.n2408 24.8557
R7483 gnd.n3299 gnd.n2396 24.8557
R7484 gnd.n3327 gnd.n3326 24.8557
R7485 gnd.n3338 gnd.n2381 24.8557
R7486 gnd.n3350 gnd.n2374 24.8557
R7487 gnd.n3622 gnd.n3621 24.8557
R7488 gnd.n3644 gnd.n2347 24.8557
R7489 gnd.n5359 gnd.n1700 24.8557
R7490 gnd.n2997 gnd.t65 23.2624
R7491 gnd.n2698 gnd.t263 22.6251
R7492 gnd.n4129 gnd.t105 21.9878
R7493 gnd.n114 gnd.t136 21.9878
R7494 gnd.n6013 gnd.t88 21.6691
R7495 gnd.n4754 gnd.n2049 21.6691
R7496 gnd.n4784 gnd.n2036 21.6691
R7497 gnd.n4766 gnd.n2005 21.6691
R7498 gnd.n4860 gnd.n1988 21.6691
R7499 gnd.n4882 gnd.n1962 21.6691
R7500 gnd.n4890 gnd.n1955 21.6691
R7501 gnd.n4897 gnd.n1948 21.6691
R7502 gnd.n4951 gnd.n1937 21.6691
R7503 gnd.n4939 gnd.n1928 21.6691
R7504 gnd.n5005 gnd.n1916 21.6691
R7505 gnd.n5023 gnd.n1898 21.6691
R7506 gnd.n5035 gnd.n1887 21.6691
R7507 gnd.n5051 gnd.n1877 21.6691
R7508 gnd.n5057 gnd.n1861 21.6691
R7509 gnd.n5138 gnd.n1845 21.6691
R7510 gnd.n5144 gnd.n1841 21.6691
R7511 gnd.n5197 gnd.n5196 21.6691
R7512 gnd.n6720 gnd.t70 21.6691
R7513 gnd.t29 gnd.n2703 21.3504
R7514 gnd.n4170 gnd.t140 21.3504
R7515 gnd.n4197 gnd.t129 21.3504
R7516 gnd.n6782 gnd.t95 21.3504
R7517 gnd.n6897 gnd.t120 21.3504
R7518 gnd.n4817 gnd.n2012 21.0318
R7519 gnd.n4999 gnd.n1920 21.0318
R7520 gnd.n5006 gnd.n1913 21.0318
R7521 gnd.n1832 gnd.n1826 21.0318
R7522 gnd.n3348 gnd.n1043 20.8043
R7523 gnd.t1 gnd.n2409 20.7131
R7524 gnd.n4150 gnd.t127 20.7131
R7525 gnd.n6006 gnd.t77 20.7131
R7526 gnd.n4629 gnd.t61 20.7131
R7527 gnd.n1689 gnd.t39 20.7131
R7528 gnd.n6755 gnd.t100 20.7131
R7529 gnd.t103 gnd.n88 20.7131
R7530 gnd.t8 gnd.n2444 20.0758
R7531 gnd.n4109 gnd.t79 20.0758
R7532 gnd.n5982 gnd.t83 20.0758
R7533 gnd.n5448 gnd.t90 20.0758
R7534 gnd.t114 gnd.n127 20.0758
R7535 gnd.n4675 gnd.n4674 19.9763
R7536 gnd.n1763 gnd.n1762 19.9763
R7537 gnd.n5838 gnd.n5837 19.9763
R7538 gnd.n1757 gnd.n1756 19.9763
R7539 gnd.n1259 gnd.t303 19.8005
R7540 gnd.n1259 gnd.t323 19.8005
R7541 gnd.n1258 gnd.t255 19.8005
R7542 gnd.n1258 gnd.t206 19.8005
R7543 gnd.n1726 gnd.t231 19.8005
R7544 gnd.n1726 gnd.t275 19.8005
R7545 gnd.n1725 gnd.t249 19.8005
R7546 gnd.n1725 gnd.t278 19.8005
R7547 gnd.n4806 gnd.n2027 19.7572
R7548 gnd.n4945 gnd.n1943 19.7572
R7549 gnd.n5017 gnd.n5016 19.7572
R7550 gnd.n5174 gnd.n1820 19.7572
R7551 gnd.t274 gnd.n1708 19.7572
R7552 gnd.n1255 gnd.n1254 19.5087
R7553 gnd.n1268 gnd.n1255 19.5087
R7554 gnd.n1266 gnd.n1257 19.5087
R7555 gnd.n1730 gnd.n1724 19.5087
R7556 gnd.n3164 gnd.t28 19.4385
R7557 gnd.n4590 gnd.n2094 19.3944
R7558 gnd.n4590 gnd.n2092 19.3944
R7559 gnd.n4594 gnd.n2092 19.3944
R7560 gnd.n4594 gnd.n2079 19.3944
R7561 gnd.n4606 gnd.n2079 19.3944
R7562 gnd.n4606 gnd.n2076 19.3944
R7563 gnd.n4627 gnd.n2076 19.3944
R7564 gnd.n4627 gnd.n2077 19.3944
R7565 gnd.n4623 gnd.n2077 19.3944
R7566 gnd.n4623 gnd.n4622 19.3944
R7567 gnd.n4622 gnd.n4621 19.3944
R7568 gnd.n4621 gnd.n4612 19.3944
R7569 gnd.n4617 gnd.n4612 19.3944
R7570 gnd.n4617 gnd.n4616 19.3944
R7571 gnd.n4616 gnd.n1292 19.3944
R7572 gnd.n5823 gnd.n1292 19.3944
R7573 gnd.n5823 gnd.n1293 19.3944
R7574 gnd.n5819 gnd.n1293 19.3944
R7575 gnd.n5819 gnd.n5818 19.3944
R7576 gnd.n5818 gnd.n5817 19.3944
R7577 gnd.n5817 gnd.n1299 19.3944
R7578 gnd.n5813 gnd.n1299 19.3944
R7579 gnd.n5813 gnd.n5812 19.3944
R7580 gnd.n5812 gnd.n5811 19.3944
R7581 gnd.n5811 gnd.n1304 19.3944
R7582 gnd.n5807 gnd.n1304 19.3944
R7583 gnd.n5807 gnd.n5806 19.3944
R7584 gnd.n5806 gnd.n5805 19.3944
R7585 gnd.n5805 gnd.n1309 19.3944
R7586 gnd.n5801 gnd.n1309 19.3944
R7587 gnd.n5801 gnd.n5800 19.3944
R7588 gnd.n5800 gnd.n5799 19.3944
R7589 gnd.n5799 gnd.n1314 19.3944
R7590 gnd.n5795 gnd.n1314 19.3944
R7591 gnd.n5795 gnd.n5794 19.3944
R7592 gnd.n5794 gnd.n5793 19.3944
R7593 gnd.n5793 gnd.n1319 19.3944
R7594 gnd.n5789 gnd.n1319 19.3944
R7595 gnd.n5789 gnd.n5788 19.3944
R7596 gnd.n5788 gnd.n5787 19.3944
R7597 gnd.n5787 gnd.n1324 19.3944
R7598 gnd.n5783 gnd.n1324 19.3944
R7599 gnd.n5783 gnd.n5782 19.3944
R7600 gnd.n5782 gnd.n5781 19.3944
R7601 gnd.n5781 gnd.n1329 19.3944
R7602 gnd.n5777 gnd.n1329 19.3944
R7603 gnd.n5777 gnd.n5776 19.3944
R7604 gnd.n5776 gnd.n5775 19.3944
R7605 gnd.n5775 gnd.n1334 19.3944
R7606 gnd.n5771 gnd.n1334 19.3944
R7607 gnd.n5771 gnd.n5770 19.3944
R7608 gnd.n5770 gnd.n5769 19.3944
R7609 gnd.n5769 gnd.n1339 19.3944
R7610 gnd.n5765 gnd.n1339 19.3944
R7611 gnd.n5765 gnd.n5764 19.3944
R7612 gnd.n5764 gnd.n5763 19.3944
R7613 gnd.n5763 gnd.n1344 19.3944
R7614 gnd.n5759 gnd.n1344 19.3944
R7615 gnd.n5759 gnd.n5758 19.3944
R7616 gnd.n5758 gnd.n5757 19.3944
R7617 gnd.n5757 gnd.n1349 19.3944
R7618 gnd.n5753 gnd.n1349 19.3944
R7619 gnd.n5753 gnd.n5752 19.3944
R7620 gnd.n5752 gnd.n5751 19.3944
R7621 gnd.n5751 gnd.n1354 19.3944
R7622 gnd.n5747 gnd.n1354 19.3944
R7623 gnd.n5747 gnd.n5746 19.3944
R7624 gnd.n5746 gnd.n5745 19.3944
R7625 gnd.n5745 gnd.n1359 19.3944
R7626 gnd.n5741 gnd.n1359 19.3944
R7627 gnd.n5741 gnd.n5740 19.3944
R7628 gnd.n5740 gnd.n5739 19.3944
R7629 gnd.n5739 gnd.n1364 19.3944
R7630 gnd.n5735 gnd.n1364 19.3944
R7631 gnd.n5735 gnd.n5734 19.3944
R7632 gnd.n5734 gnd.n5733 19.3944
R7633 gnd.n5733 gnd.n1369 19.3944
R7634 gnd.n5729 gnd.n1369 19.3944
R7635 gnd.n5729 gnd.n5728 19.3944
R7636 gnd.n5728 gnd.n5727 19.3944
R7637 gnd.n5727 gnd.n1374 19.3944
R7638 gnd.n5723 gnd.n1374 19.3944
R7639 gnd.n4375 gnd.n4374 19.3944
R7640 gnd.n4374 gnd.n2119 19.3944
R7641 gnd.n4577 gnd.n2119 19.3944
R7642 gnd.n4300 gnd.n4299 19.3944
R7643 gnd.n4303 gnd.n4300 19.3944
R7644 gnd.n4303 gnd.n4273 19.3944
R7645 gnd.n4307 gnd.n4273 19.3944
R7646 gnd.n4308 gnd.n4307 19.3944
R7647 gnd.n4424 gnd.n4308 19.3944
R7648 gnd.n4424 gnd.n4423 19.3944
R7649 gnd.n4423 gnd.n4422 19.3944
R7650 gnd.n4422 gnd.n4313 19.3944
R7651 gnd.n4415 gnd.n4313 19.3944
R7652 gnd.n4415 gnd.n4414 19.3944
R7653 gnd.n4414 gnd.n4322 19.3944
R7654 gnd.n4407 gnd.n4322 19.3944
R7655 gnd.n4407 gnd.n4406 19.3944
R7656 gnd.n4406 gnd.n4332 19.3944
R7657 gnd.n4399 gnd.n4332 19.3944
R7658 gnd.n4399 gnd.n4398 19.3944
R7659 gnd.n4398 gnd.n4342 19.3944
R7660 gnd.n4391 gnd.n4342 19.3944
R7661 gnd.n4391 gnd.n4390 19.3944
R7662 gnd.n4390 gnd.n4352 19.3944
R7663 gnd.n4383 gnd.n4352 19.3944
R7664 gnd.n4383 gnd.n4382 19.3944
R7665 gnd.n4382 gnd.n4362 19.3944
R7666 gnd.n5699 gnd.n1400 19.3944
R7667 gnd.n5699 gnd.n5698 19.3944
R7668 gnd.n5698 gnd.n1403 19.3944
R7669 gnd.n5691 gnd.n1403 19.3944
R7670 gnd.n5691 gnd.n5690 19.3944
R7671 gnd.n5690 gnd.n1411 19.3944
R7672 gnd.n5683 gnd.n1411 19.3944
R7673 gnd.n5683 gnd.n5682 19.3944
R7674 gnd.n5682 gnd.n1419 19.3944
R7675 gnd.n5675 gnd.n1419 19.3944
R7676 gnd.n5675 gnd.n5674 19.3944
R7677 gnd.n5674 gnd.n1427 19.3944
R7678 gnd.n5667 gnd.n1427 19.3944
R7679 gnd.n5667 gnd.n5666 19.3944
R7680 gnd.n5666 gnd.n1435 19.3944
R7681 gnd.n5659 gnd.n1435 19.3944
R7682 gnd.n2879 gnd.n2878 19.3944
R7683 gnd.n2878 gnd.n2877 19.3944
R7684 gnd.n2877 gnd.n2876 19.3944
R7685 gnd.n2876 gnd.n2874 19.3944
R7686 gnd.n2874 gnd.n2871 19.3944
R7687 gnd.n2871 gnd.n2870 19.3944
R7688 gnd.n2870 gnd.n2867 19.3944
R7689 gnd.n2867 gnd.n2866 19.3944
R7690 gnd.n2866 gnd.n2863 19.3944
R7691 gnd.n2863 gnd.n2862 19.3944
R7692 gnd.n2862 gnd.n2859 19.3944
R7693 gnd.n2859 gnd.n2858 19.3944
R7694 gnd.n2858 gnd.n2855 19.3944
R7695 gnd.n2855 gnd.n2854 19.3944
R7696 gnd.n2854 gnd.n2851 19.3944
R7697 gnd.n2851 gnd.n2850 19.3944
R7698 gnd.n2850 gnd.n2847 19.3944
R7699 gnd.n2847 gnd.n2846 19.3944
R7700 gnd.n2846 gnd.n2843 19.3944
R7701 gnd.n2843 gnd.n2842 19.3944
R7702 gnd.n2842 gnd.n2839 19.3944
R7703 gnd.n2839 gnd.n2838 19.3944
R7704 gnd.n2835 gnd.n2834 19.3944
R7705 gnd.n2834 gnd.n2790 19.3944
R7706 gnd.n2885 gnd.n2790 19.3944
R7707 gnd.n3652 gnd.n3651 19.3944
R7708 gnd.n3651 gnd.n3648 19.3944
R7709 gnd.n3648 gnd.n3647 19.3944
R7710 gnd.n3697 gnd.n3696 19.3944
R7711 gnd.n3696 gnd.n3695 19.3944
R7712 gnd.n3695 gnd.n3692 19.3944
R7713 gnd.n3692 gnd.n3691 19.3944
R7714 gnd.n3691 gnd.n3688 19.3944
R7715 gnd.n3688 gnd.n3687 19.3944
R7716 gnd.n3687 gnd.n3684 19.3944
R7717 gnd.n3684 gnd.n3683 19.3944
R7718 gnd.n3683 gnd.n3680 19.3944
R7719 gnd.n3680 gnd.n3679 19.3944
R7720 gnd.n3679 gnd.n3676 19.3944
R7721 gnd.n3676 gnd.n3675 19.3944
R7722 gnd.n3675 gnd.n3672 19.3944
R7723 gnd.n3672 gnd.n3671 19.3944
R7724 gnd.n3671 gnd.n3668 19.3944
R7725 gnd.n3668 gnd.n3667 19.3944
R7726 gnd.n3667 gnd.n3664 19.3944
R7727 gnd.n3664 gnd.n3663 19.3944
R7728 gnd.n3663 gnd.n3660 19.3944
R7729 gnd.n3660 gnd.n3659 19.3944
R7730 gnd.n3659 gnd.n3656 19.3944
R7731 gnd.n3656 gnd.n3655 19.3944
R7732 gnd.n2978 gnd.n2687 19.3944
R7733 gnd.n2988 gnd.n2687 19.3944
R7734 gnd.n2989 gnd.n2988 19.3944
R7735 gnd.n2989 gnd.n2668 19.3944
R7736 gnd.n3009 gnd.n2668 19.3944
R7737 gnd.n3009 gnd.n2660 19.3944
R7738 gnd.n3019 gnd.n2660 19.3944
R7739 gnd.n3020 gnd.n3019 19.3944
R7740 gnd.n3021 gnd.n3020 19.3944
R7741 gnd.n3021 gnd.n2643 19.3944
R7742 gnd.n3038 gnd.n2643 19.3944
R7743 gnd.n3041 gnd.n3038 19.3944
R7744 gnd.n3041 gnd.n3040 19.3944
R7745 gnd.n3040 gnd.n2616 19.3944
R7746 gnd.n3080 gnd.n2616 19.3944
R7747 gnd.n3080 gnd.n2613 19.3944
R7748 gnd.n3086 gnd.n2613 19.3944
R7749 gnd.n3087 gnd.n3086 19.3944
R7750 gnd.n3087 gnd.n2611 19.3944
R7751 gnd.n3093 gnd.n2611 19.3944
R7752 gnd.n3096 gnd.n3093 19.3944
R7753 gnd.n3098 gnd.n3096 19.3944
R7754 gnd.n3104 gnd.n3098 19.3944
R7755 gnd.n3104 gnd.n3103 19.3944
R7756 gnd.n3103 gnd.n2486 19.3944
R7757 gnd.n3170 gnd.n2486 19.3944
R7758 gnd.n3171 gnd.n3170 19.3944
R7759 gnd.n3171 gnd.n2479 19.3944
R7760 gnd.n3182 gnd.n2479 19.3944
R7761 gnd.n3183 gnd.n3182 19.3944
R7762 gnd.n3183 gnd.n2462 19.3944
R7763 gnd.n2462 gnd.n2460 19.3944
R7764 gnd.n3207 gnd.n2460 19.3944
R7765 gnd.n3208 gnd.n3207 19.3944
R7766 gnd.n3208 gnd.n2431 19.3944
R7767 gnd.n3255 gnd.n2431 19.3944
R7768 gnd.n3256 gnd.n3255 19.3944
R7769 gnd.n3256 gnd.n2424 19.3944
R7770 gnd.n3267 gnd.n2424 19.3944
R7771 gnd.n3268 gnd.n3267 19.3944
R7772 gnd.n3268 gnd.n2407 19.3944
R7773 gnd.n2407 gnd.n2405 19.3944
R7774 gnd.n3292 gnd.n2405 19.3944
R7775 gnd.n3293 gnd.n3292 19.3944
R7776 gnd.n3293 gnd.n2377 19.3944
R7777 gnd.n3344 gnd.n2377 19.3944
R7778 gnd.n3345 gnd.n3344 19.3944
R7779 gnd.n3345 gnd.n2370 19.3944
R7780 gnd.n3613 gnd.n2370 19.3944
R7781 gnd.n3614 gnd.n3613 19.3944
R7782 gnd.n3614 gnd.n2351 19.3944
R7783 gnd.n3639 gnd.n2351 19.3944
R7784 gnd.n3639 gnd.n2352 19.3944
R7785 gnd.n2969 gnd.n2968 19.3944
R7786 gnd.n2968 gnd.n2701 19.3944
R7787 gnd.n2724 gnd.n2701 19.3944
R7788 gnd.n2727 gnd.n2724 19.3944
R7789 gnd.n2727 gnd.n2720 19.3944
R7790 gnd.n2731 gnd.n2720 19.3944
R7791 gnd.n2734 gnd.n2731 19.3944
R7792 gnd.n2737 gnd.n2734 19.3944
R7793 gnd.n2737 gnd.n2718 19.3944
R7794 gnd.n2741 gnd.n2718 19.3944
R7795 gnd.n2744 gnd.n2741 19.3944
R7796 gnd.n2747 gnd.n2744 19.3944
R7797 gnd.n2747 gnd.n2716 19.3944
R7798 gnd.n2751 gnd.n2716 19.3944
R7799 gnd.n2974 gnd.n2973 19.3944
R7800 gnd.n2973 gnd.n2677 19.3944
R7801 gnd.n2999 gnd.n2677 19.3944
R7802 gnd.n2999 gnd.n2675 19.3944
R7803 gnd.n3005 gnd.n2675 19.3944
R7804 gnd.n3005 gnd.n3004 19.3944
R7805 gnd.n3004 gnd.n2649 19.3944
R7806 gnd.n3029 gnd.n2649 19.3944
R7807 gnd.n3029 gnd.n2647 19.3944
R7808 gnd.n3033 gnd.n2647 19.3944
R7809 gnd.n3033 gnd.n2627 19.3944
R7810 gnd.n3060 gnd.n2627 19.3944
R7811 gnd.n3060 gnd.n2625 19.3944
R7812 gnd.n3070 gnd.n2625 19.3944
R7813 gnd.n3070 gnd.n3069 19.3944
R7814 gnd.n3069 gnd.n3068 19.3944
R7815 gnd.n3068 gnd.n2574 19.3944
R7816 gnd.n3118 gnd.n2574 19.3944
R7817 gnd.n3118 gnd.n3117 19.3944
R7818 gnd.n3117 gnd.n3116 19.3944
R7819 gnd.n3116 gnd.n2578 19.3944
R7820 gnd.n2598 gnd.n2578 19.3944
R7821 gnd.n2598 gnd.n2496 19.3944
R7822 gnd.n3155 gnd.n2496 19.3944
R7823 gnd.n3155 gnd.n2494 19.3944
R7824 gnd.n3161 gnd.n2494 19.3944
R7825 gnd.n3161 gnd.n3160 19.3944
R7826 gnd.n3160 gnd.n2469 19.3944
R7827 gnd.n3195 gnd.n2469 19.3944
R7828 gnd.n3195 gnd.n2467 19.3944
R7829 gnd.n3201 gnd.n2467 19.3944
R7830 gnd.n3201 gnd.n3200 19.3944
R7831 gnd.n3200 gnd.n2442 19.3944
R7832 gnd.n3240 gnd.n2442 19.3944
R7833 gnd.n3240 gnd.n2440 19.3944
R7834 gnd.n3246 gnd.n2440 19.3944
R7835 gnd.n3246 gnd.n3245 19.3944
R7836 gnd.n3245 gnd.n2414 19.3944
R7837 gnd.n3280 gnd.n2414 19.3944
R7838 gnd.n3280 gnd.n2412 19.3944
R7839 gnd.n3286 gnd.n2412 19.3944
R7840 gnd.n3286 gnd.n3285 19.3944
R7841 gnd.n3285 gnd.n2387 19.3944
R7842 gnd.n3329 gnd.n2387 19.3944
R7843 gnd.n3329 gnd.n2385 19.3944
R7844 gnd.n3335 gnd.n2385 19.3944
R7845 gnd.n3335 gnd.n3334 19.3944
R7846 gnd.n3334 gnd.n2360 19.3944
R7847 gnd.n3624 gnd.n2360 19.3944
R7848 gnd.n3624 gnd.n2358 19.3944
R7849 gnd.n3632 gnd.n2358 19.3944
R7850 gnd.n3632 gnd.n3631 19.3944
R7851 gnd.n3631 gnd.n3630 19.3944
R7852 gnd.n3733 gnd.n3732 19.3944
R7853 gnd.n3732 gnd.n2299 19.3944
R7854 gnd.n3728 gnd.n2299 19.3944
R7855 gnd.n3728 gnd.n3725 19.3944
R7856 gnd.n3725 gnd.n3722 19.3944
R7857 gnd.n3722 gnd.n3721 19.3944
R7858 gnd.n3721 gnd.n3718 19.3944
R7859 gnd.n3718 gnd.n3717 19.3944
R7860 gnd.n3717 gnd.n3714 19.3944
R7861 gnd.n3714 gnd.n3713 19.3944
R7862 gnd.n3713 gnd.n3710 19.3944
R7863 gnd.n3710 gnd.n3709 19.3944
R7864 gnd.n3709 gnd.n3706 19.3944
R7865 gnd.n3706 gnd.n3705 19.3944
R7866 gnd.n2889 gnd.n2788 19.3944
R7867 gnd.n2889 gnd.n2779 19.3944
R7868 gnd.n2902 gnd.n2779 19.3944
R7869 gnd.n2902 gnd.n2777 19.3944
R7870 gnd.n2906 gnd.n2777 19.3944
R7871 gnd.n2906 gnd.n2767 19.3944
R7872 gnd.n2918 gnd.n2767 19.3944
R7873 gnd.n2918 gnd.n2765 19.3944
R7874 gnd.n2952 gnd.n2765 19.3944
R7875 gnd.n2952 gnd.n2951 19.3944
R7876 gnd.n2951 gnd.n2950 19.3944
R7877 gnd.n2950 gnd.n2949 19.3944
R7878 gnd.n2949 gnd.n2946 19.3944
R7879 gnd.n2946 gnd.n2945 19.3944
R7880 gnd.n2945 gnd.n2944 19.3944
R7881 gnd.n2944 gnd.n2942 19.3944
R7882 gnd.n2942 gnd.n2941 19.3944
R7883 gnd.n2941 gnd.n2938 19.3944
R7884 gnd.n2938 gnd.n2937 19.3944
R7885 gnd.n2937 gnd.n2936 19.3944
R7886 gnd.n2936 gnd.n2934 19.3944
R7887 gnd.n2934 gnd.n2633 19.3944
R7888 gnd.n3049 gnd.n2633 19.3944
R7889 gnd.n3049 gnd.n2631 19.3944
R7890 gnd.n3055 gnd.n2631 19.3944
R7891 gnd.n3055 gnd.n3054 19.3944
R7892 gnd.n3054 gnd.n2555 19.3944
R7893 gnd.n3129 gnd.n2555 19.3944
R7894 gnd.n3129 gnd.n2556 19.3944
R7895 gnd.n2603 gnd.n2602 19.3944
R7896 gnd.n2606 gnd.n2605 19.3944
R7897 gnd.n2593 gnd.n2592 19.3944
R7898 gnd.n3148 gnd.n2501 19.3944
R7899 gnd.n3148 gnd.n3147 19.3944
R7900 gnd.n3147 gnd.n3146 19.3944
R7901 gnd.n3146 gnd.n3144 19.3944
R7902 gnd.n3144 gnd.n3143 19.3944
R7903 gnd.n3143 gnd.n3141 19.3944
R7904 gnd.n3141 gnd.n3140 19.3944
R7905 gnd.n3140 gnd.n2450 19.3944
R7906 gnd.n3216 gnd.n2450 19.3944
R7907 gnd.n3216 gnd.n2448 19.3944
R7908 gnd.n3235 gnd.n2448 19.3944
R7909 gnd.n3235 gnd.n3234 19.3944
R7910 gnd.n3234 gnd.n3233 19.3944
R7911 gnd.n3233 gnd.n3231 19.3944
R7912 gnd.n3231 gnd.n3230 19.3944
R7913 gnd.n3230 gnd.n3228 19.3944
R7914 gnd.n3228 gnd.n3227 19.3944
R7915 gnd.n3227 gnd.n2394 19.3944
R7916 gnd.n3301 gnd.n2394 19.3944
R7917 gnd.n3301 gnd.n2392 19.3944
R7918 gnd.n3324 gnd.n2392 19.3944
R7919 gnd.n3324 gnd.n3323 19.3944
R7920 gnd.n3323 gnd.n3322 19.3944
R7921 gnd.n3322 gnd.n3319 19.3944
R7922 gnd.n3319 gnd.n3318 19.3944
R7923 gnd.n3318 gnd.n3316 19.3944
R7924 gnd.n3316 gnd.n3315 19.3944
R7925 gnd.n3315 gnd.n3313 19.3944
R7926 gnd.n3313 gnd.n2346 19.3944
R7927 gnd.n2894 gnd.n2784 19.3944
R7928 gnd.n2894 gnd.n2782 19.3944
R7929 gnd.n2898 gnd.n2782 19.3944
R7930 gnd.n2898 gnd.n2773 19.3944
R7931 gnd.n2910 gnd.n2773 19.3944
R7932 gnd.n2910 gnd.n2771 19.3944
R7933 gnd.n2914 gnd.n2771 19.3944
R7934 gnd.n2914 gnd.n2760 19.3944
R7935 gnd.n2956 gnd.n2760 19.3944
R7936 gnd.n2956 gnd.n2714 19.3944
R7937 gnd.n2962 gnd.n2714 19.3944
R7938 gnd.n2962 gnd.n2961 19.3944
R7939 gnd.n2961 gnd.n2692 19.3944
R7940 gnd.n2983 gnd.n2692 19.3944
R7941 gnd.n2983 gnd.n2685 19.3944
R7942 gnd.n2994 gnd.n2685 19.3944
R7943 gnd.n2994 gnd.n2993 19.3944
R7944 gnd.n2993 gnd.n2666 19.3944
R7945 gnd.n3014 gnd.n2666 19.3944
R7946 gnd.n3014 gnd.n2656 19.3944
R7947 gnd.n3024 gnd.n2656 19.3944
R7948 gnd.n3024 gnd.n2639 19.3944
R7949 gnd.n3045 gnd.n2639 19.3944
R7950 gnd.n3045 gnd.n3044 19.3944
R7951 gnd.n3044 gnd.n2618 19.3944
R7952 gnd.n3075 gnd.n2618 19.3944
R7953 gnd.n3075 gnd.n2563 19.3944
R7954 gnd.n3125 gnd.n2563 19.3944
R7955 gnd.n3125 gnd.n3124 19.3944
R7956 gnd.n3124 gnd.n3123 19.3944
R7957 gnd.n3123 gnd.n2567 19.3944
R7958 gnd.n2585 gnd.n2567 19.3944
R7959 gnd.n3111 gnd.n2585 19.3944
R7960 gnd.n3111 gnd.n3110 19.3944
R7961 gnd.n3110 gnd.n3109 19.3944
R7962 gnd.n3109 gnd.n2589 19.3944
R7963 gnd.n2589 gnd.n2488 19.3944
R7964 gnd.n3166 gnd.n2488 19.3944
R7965 gnd.n3166 gnd.n2481 19.3944
R7966 gnd.n3177 gnd.n2481 19.3944
R7967 gnd.n3177 gnd.n2477 19.3944
R7968 gnd.n3190 gnd.n2477 19.3944
R7969 gnd.n3190 gnd.n3189 19.3944
R7970 gnd.n3189 gnd.n2456 19.3944
R7971 gnd.n3212 gnd.n2456 19.3944
R7972 gnd.n3212 gnd.n3211 19.3944
R7973 gnd.n3211 gnd.n2433 19.3944
R7974 gnd.n3251 gnd.n2433 19.3944
R7975 gnd.n3251 gnd.n2426 19.3944
R7976 gnd.n3262 gnd.n2426 19.3944
R7977 gnd.n3262 gnd.n2422 19.3944
R7978 gnd.n3275 gnd.n2422 19.3944
R7979 gnd.n3275 gnd.n3274 19.3944
R7980 gnd.n3274 gnd.n2401 19.3944
R7981 gnd.n3297 gnd.n2401 19.3944
R7982 gnd.n3297 gnd.n3296 19.3944
R7983 gnd.n3296 gnd.n2379 19.3944
R7984 gnd.n3340 gnd.n2379 19.3944
R7985 gnd.n3340 gnd.n2372 19.3944
R7986 gnd.n3352 gnd.n2372 19.3944
R7987 gnd.n3352 gnd.n2368 19.3944
R7988 gnd.n3619 gnd.n2368 19.3944
R7989 gnd.n3619 gnd.n3618 19.3944
R7990 gnd.n3618 gnd.n2349 19.3944
R7991 gnd.n3642 gnd.n2349 19.3944
R7992 gnd.n4419 gnd.n4418 19.3944
R7993 gnd.n4418 gnd.n4316 19.3944
R7994 gnd.n4411 gnd.n4316 19.3944
R7995 gnd.n4411 gnd.n4410 19.3944
R7996 gnd.n4410 gnd.n4328 19.3944
R7997 gnd.n4403 gnd.n4328 19.3944
R7998 gnd.n4403 gnd.n4402 19.3944
R7999 gnd.n4402 gnd.n4336 19.3944
R8000 gnd.n4395 gnd.n4336 19.3944
R8001 gnd.n4395 gnd.n4394 19.3944
R8002 gnd.n4394 gnd.n4348 19.3944
R8003 gnd.n4387 gnd.n4348 19.3944
R8004 gnd.n4387 gnd.n4386 19.3944
R8005 gnd.n4386 gnd.n4356 19.3944
R8006 gnd.n4379 gnd.n4356 19.3944
R8007 gnd.n4379 gnd.n4378 19.3944
R8008 gnd.n4233 gnd.n4231 19.3944
R8009 gnd.n4233 gnd.n4228 19.3944
R8010 gnd.n4237 gnd.n4228 19.3944
R8011 gnd.n4237 gnd.n2153 19.3944
R8012 gnd.n4241 gnd.n2153 19.3944
R8013 gnd.n4241 gnd.n2151 19.3944
R8014 gnd.n4249 gnd.n2151 19.3944
R8015 gnd.n4249 gnd.n4248 19.3944
R8016 gnd.n4248 gnd.n4247 19.3944
R8017 gnd.n4247 gnd.n2135 19.3944
R8018 gnd.n4546 gnd.n2135 19.3944
R8019 gnd.n4546 gnd.n2133 19.3944
R8020 gnd.n4550 gnd.n2133 19.3944
R8021 gnd.n4550 gnd.n2131 19.3944
R8022 gnd.n4554 gnd.n2131 19.3944
R8023 gnd.n4554 gnd.n2129 19.3944
R8024 gnd.n4566 gnd.n2129 19.3944
R8025 gnd.n4566 gnd.n4565 19.3944
R8026 gnd.n4565 gnd.n4564 19.3944
R8027 gnd.n4564 gnd.n4561 19.3944
R8028 gnd.n4561 gnd.n2101 19.3944
R8029 gnd.n4582 gnd.n2101 19.3944
R8030 gnd.n4582 gnd.n2099 19.3944
R8031 gnd.n4586 gnd.n2099 19.3944
R8032 gnd.n4586 gnd.n2087 19.3944
R8033 gnd.n4598 gnd.n2087 19.3944
R8034 gnd.n4598 gnd.n2085 19.3944
R8035 gnd.n4602 gnd.n2085 19.3944
R8036 gnd.n4602 gnd.n2071 19.3944
R8037 gnd.n4631 gnd.n2071 19.3944
R8038 gnd.n4631 gnd.n2069 19.3944
R8039 gnd.n4644 gnd.n2069 19.3944
R8040 gnd.n4644 gnd.n4643 19.3944
R8041 gnd.n4643 gnd.n4642 19.3944
R8042 gnd.n4642 gnd.n4639 19.3944
R8043 gnd.n4639 gnd.n1283 19.3944
R8044 gnd.n5829 gnd.n1283 19.3944
R8045 gnd.n5829 gnd.n5828 19.3944
R8046 gnd.n5828 gnd.n5827 19.3944
R8047 gnd.n5827 gnd.n1287 19.3944
R8048 gnd.n2034 gnd.n1287 19.3944
R8049 gnd.n4798 gnd.n2034 19.3944
R8050 gnd.n4798 gnd.n2031 19.3944
R8051 gnd.n4804 gnd.n2031 19.3944
R8052 gnd.n4804 gnd.n4803 19.3944
R8053 gnd.n4803 gnd.n2010 19.3944
R8054 gnd.n4830 gnd.n2010 19.3944
R8055 gnd.n4830 gnd.n2008 19.3944
R8056 gnd.n4834 gnd.n2008 19.3944
R8057 gnd.n4834 gnd.n1986 19.3944
R8058 gnd.n4869 gnd.n1986 19.3944
R8059 gnd.n4869 gnd.n1984 19.3944
R8060 gnd.n4873 gnd.n1984 19.3944
R8061 gnd.n4873 gnd.n1960 19.3944
R8062 gnd.n4909 gnd.n1960 19.3944
R8063 gnd.n4909 gnd.n1958 19.3944
R8064 gnd.n4915 gnd.n1958 19.3944
R8065 gnd.n4915 gnd.n4914 19.3944
R8066 gnd.n4914 gnd.n1933 19.3944
R8067 gnd.n4955 gnd.n1933 19.3944
R8068 gnd.n4955 gnd.n1931 19.3944
R8069 gnd.n4961 gnd.n1931 19.3944
R8070 gnd.n4961 gnd.n4960 19.3944
R8071 gnd.n4960 gnd.n1911 19.3944
R8072 gnd.n5008 gnd.n1911 19.3944
R8073 gnd.n5008 gnd.n1909 19.3944
R8074 gnd.n5014 gnd.n1909 19.3944
R8075 gnd.n5014 gnd.n5013 19.3944
R8076 gnd.n5013 gnd.n1885 19.3944
R8077 gnd.n5044 gnd.n1885 19.3944
R8078 gnd.n5044 gnd.n1883 19.3944
R8079 gnd.n5048 gnd.n1883 19.3944
R8080 gnd.n5048 gnd.n1859 19.3944
R8081 gnd.n5088 gnd.n1859 19.3944
R8082 gnd.n5088 gnd.n1857 19.3944
R8083 gnd.n5094 gnd.n1857 19.3944
R8084 gnd.n5094 gnd.n5093 19.3944
R8085 gnd.n5093 gnd.n1836 19.3944
R8086 gnd.n5147 gnd.n1836 19.3944
R8087 gnd.n5147 gnd.n1834 19.3944
R8088 gnd.n5151 gnd.n1834 19.3944
R8089 gnd.n5151 gnd.n1814 19.3944
R8090 gnd.n5177 gnd.n1814 19.3944
R8091 gnd.n5177 gnd.n1812 19.3944
R8092 gnd.n5181 gnd.n1812 19.3944
R8093 gnd.n5181 gnd.n1797 19.3944
R8094 gnd.n5206 gnd.n1797 19.3944
R8095 gnd.n5206 gnd.n1795 19.3944
R8096 gnd.n5210 gnd.n1795 19.3944
R8097 gnd.n5210 gnd.n1706 19.3944
R8098 gnd.n5353 gnd.n1706 19.3944
R8099 gnd.n5353 gnd.n1704 19.3944
R8100 gnd.n5357 gnd.n1704 19.3944
R8101 gnd.n5357 gnd.n1693 19.3944
R8102 gnd.n5369 gnd.n1693 19.3944
R8103 gnd.n5369 gnd.n1691 19.3944
R8104 gnd.n5373 gnd.n1691 19.3944
R8105 gnd.n5373 gnd.n1680 19.3944
R8106 gnd.n5385 gnd.n1680 19.3944
R8107 gnd.n5385 gnd.n1678 19.3944
R8108 gnd.n5392 gnd.n1678 19.3944
R8109 gnd.n5392 gnd.n5391 19.3944
R8110 gnd.n5391 gnd.n1667 19.3944
R8111 gnd.n5405 gnd.n1667 19.3944
R8112 gnd.n5406 gnd.n5405 19.3944
R8113 gnd.n5406 gnd.n1665 19.3944
R8114 gnd.n5424 gnd.n1665 19.3944
R8115 gnd.n5424 gnd.n5423 19.3944
R8116 gnd.n5423 gnd.n5422 19.3944
R8117 gnd.n5422 gnd.n5412 19.3944
R8118 gnd.n5418 gnd.n5412 19.3944
R8119 gnd.n5418 gnd.n5417 19.3944
R8120 gnd.n5417 gnd.n1633 19.3944
R8121 gnd.n1633 gnd.n1631 19.3944
R8122 gnd.n5475 gnd.n1631 19.3944
R8123 gnd.n5475 gnd.n1629 19.3944
R8124 gnd.n5479 gnd.n1629 19.3944
R8125 gnd.n5479 gnd.n1627 19.3944
R8126 gnd.n5483 gnd.n1627 19.3944
R8127 gnd.n5483 gnd.n1625 19.3944
R8128 gnd.n5496 gnd.n1625 19.3944
R8129 gnd.n5496 gnd.n5495 19.3944
R8130 gnd.n5495 gnd.n5494 19.3944
R8131 gnd.n5494 gnd.n5491 19.3944
R8132 gnd.n5491 gnd.n559 19.3944
R8133 gnd.n6726 gnd.n559 19.3944
R8134 gnd.n6726 gnd.n6725 19.3944
R8135 gnd.n6725 gnd.n6724 19.3944
R8136 gnd.n6508 gnd.n685 19.3944
R8137 gnd.n6514 gnd.n685 19.3944
R8138 gnd.n6514 gnd.n683 19.3944
R8139 gnd.n6518 gnd.n683 19.3944
R8140 gnd.n6518 gnd.n679 19.3944
R8141 gnd.n6524 gnd.n679 19.3944
R8142 gnd.n6524 gnd.n677 19.3944
R8143 gnd.n6528 gnd.n677 19.3944
R8144 gnd.n6528 gnd.n673 19.3944
R8145 gnd.n6534 gnd.n673 19.3944
R8146 gnd.n6534 gnd.n671 19.3944
R8147 gnd.n6538 gnd.n671 19.3944
R8148 gnd.n6538 gnd.n667 19.3944
R8149 gnd.n6544 gnd.n667 19.3944
R8150 gnd.n6544 gnd.n665 19.3944
R8151 gnd.n6548 gnd.n665 19.3944
R8152 gnd.n6548 gnd.n661 19.3944
R8153 gnd.n6554 gnd.n661 19.3944
R8154 gnd.n6554 gnd.n659 19.3944
R8155 gnd.n6558 gnd.n659 19.3944
R8156 gnd.n6558 gnd.n655 19.3944
R8157 gnd.n6564 gnd.n655 19.3944
R8158 gnd.n6564 gnd.n653 19.3944
R8159 gnd.n6568 gnd.n653 19.3944
R8160 gnd.n6568 gnd.n649 19.3944
R8161 gnd.n6574 gnd.n649 19.3944
R8162 gnd.n6574 gnd.n647 19.3944
R8163 gnd.n6578 gnd.n647 19.3944
R8164 gnd.n6578 gnd.n643 19.3944
R8165 gnd.n6584 gnd.n643 19.3944
R8166 gnd.n6584 gnd.n641 19.3944
R8167 gnd.n6588 gnd.n641 19.3944
R8168 gnd.n6588 gnd.n637 19.3944
R8169 gnd.n6594 gnd.n637 19.3944
R8170 gnd.n6594 gnd.n635 19.3944
R8171 gnd.n6598 gnd.n635 19.3944
R8172 gnd.n6598 gnd.n631 19.3944
R8173 gnd.n6604 gnd.n631 19.3944
R8174 gnd.n6604 gnd.n629 19.3944
R8175 gnd.n6608 gnd.n629 19.3944
R8176 gnd.n6608 gnd.n625 19.3944
R8177 gnd.n6614 gnd.n625 19.3944
R8178 gnd.n6614 gnd.n623 19.3944
R8179 gnd.n6618 gnd.n623 19.3944
R8180 gnd.n6618 gnd.n619 19.3944
R8181 gnd.n6624 gnd.n619 19.3944
R8182 gnd.n6624 gnd.n617 19.3944
R8183 gnd.n6628 gnd.n617 19.3944
R8184 gnd.n6628 gnd.n613 19.3944
R8185 gnd.n6634 gnd.n613 19.3944
R8186 gnd.n6634 gnd.n611 19.3944
R8187 gnd.n6638 gnd.n611 19.3944
R8188 gnd.n6638 gnd.n607 19.3944
R8189 gnd.n6644 gnd.n607 19.3944
R8190 gnd.n6644 gnd.n605 19.3944
R8191 gnd.n6648 gnd.n605 19.3944
R8192 gnd.n6648 gnd.n601 19.3944
R8193 gnd.n6654 gnd.n601 19.3944
R8194 gnd.n6654 gnd.n599 19.3944
R8195 gnd.n6658 gnd.n599 19.3944
R8196 gnd.n6658 gnd.n595 19.3944
R8197 gnd.n6664 gnd.n595 19.3944
R8198 gnd.n6664 gnd.n593 19.3944
R8199 gnd.n6668 gnd.n593 19.3944
R8200 gnd.n6668 gnd.n589 19.3944
R8201 gnd.n6674 gnd.n589 19.3944
R8202 gnd.n6674 gnd.n587 19.3944
R8203 gnd.n6678 gnd.n587 19.3944
R8204 gnd.n6678 gnd.n583 19.3944
R8205 gnd.n6684 gnd.n583 19.3944
R8206 gnd.n6684 gnd.n581 19.3944
R8207 gnd.n6688 gnd.n581 19.3944
R8208 gnd.n6688 gnd.n577 19.3944
R8209 gnd.n6694 gnd.n577 19.3944
R8210 gnd.n6694 gnd.n575 19.3944
R8211 gnd.n6698 gnd.n575 19.3944
R8212 gnd.n6698 gnd.n571 19.3944
R8213 gnd.n6704 gnd.n571 19.3944
R8214 gnd.n6704 gnd.n569 19.3944
R8215 gnd.n6708 gnd.n569 19.3944
R8216 gnd.n6708 gnd.n565 19.3944
R8217 gnd.n6715 gnd.n565 19.3944
R8218 gnd.n6715 gnd.n563 19.3944
R8219 gnd.n6719 gnd.n563 19.3944
R8220 gnd.n6187 gnd.n880 19.3944
R8221 gnd.n6187 gnd.n876 19.3944
R8222 gnd.n6193 gnd.n876 19.3944
R8223 gnd.n6193 gnd.n874 19.3944
R8224 gnd.n6197 gnd.n874 19.3944
R8225 gnd.n6197 gnd.n870 19.3944
R8226 gnd.n6203 gnd.n870 19.3944
R8227 gnd.n6203 gnd.n868 19.3944
R8228 gnd.n6207 gnd.n868 19.3944
R8229 gnd.n6207 gnd.n864 19.3944
R8230 gnd.n6213 gnd.n864 19.3944
R8231 gnd.n6213 gnd.n862 19.3944
R8232 gnd.n6217 gnd.n862 19.3944
R8233 gnd.n6217 gnd.n858 19.3944
R8234 gnd.n6223 gnd.n858 19.3944
R8235 gnd.n6223 gnd.n856 19.3944
R8236 gnd.n6227 gnd.n856 19.3944
R8237 gnd.n6227 gnd.n852 19.3944
R8238 gnd.n6233 gnd.n852 19.3944
R8239 gnd.n6233 gnd.n850 19.3944
R8240 gnd.n6237 gnd.n850 19.3944
R8241 gnd.n6237 gnd.n846 19.3944
R8242 gnd.n6243 gnd.n846 19.3944
R8243 gnd.n6243 gnd.n844 19.3944
R8244 gnd.n6247 gnd.n844 19.3944
R8245 gnd.n6247 gnd.n840 19.3944
R8246 gnd.n6253 gnd.n840 19.3944
R8247 gnd.n6253 gnd.n838 19.3944
R8248 gnd.n6257 gnd.n838 19.3944
R8249 gnd.n6257 gnd.n834 19.3944
R8250 gnd.n6263 gnd.n834 19.3944
R8251 gnd.n6263 gnd.n832 19.3944
R8252 gnd.n6267 gnd.n832 19.3944
R8253 gnd.n6267 gnd.n828 19.3944
R8254 gnd.n6273 gnd.n828 19.3944
R8255 gnd.n6273 gnd.n826 19.3944
R8256 gnd.n6277 gnd.n826 19.3944
R8257 gnd.n6277 gnd.n822 19.3944
R8258 gnd.n6283 gnd.n822 19.3944
R8259 gnd.n6283 gnd.n820 19.3944
R8260 gnd.n6287 gnd.n820 19.3944
R8261 gnd.n6287 gnd.n816 19.3944
R8262 gnd.n6293 gnd.n816 19.3944
R8263 gnd.n6293 gnd.n814 19.3944
R8264 gnd.n6297 gnd.n814 19.3944
R8265 gnd.n6297 gnd.n810 19.3944
R8266 gnd.n6303 gnd.n810 19.3944
R8267 gnd.n6303 gnd.n808 19.3944
R8268 gnd.n6307 gnd.n808 19.3944
R8269 gnd.n6307 gnd.n804 19.3944
R8270 gnd.n6313 gnd.n804 19.3944
R8271 gnd.n6313 gnd.n802 19.3944
R8272 gnd.n6317 gnd.n802 19.3944
R8273 gnd.n6317 gnd.n798 19.3944
R8274 gnd.n6323 gnd.n798 19.3944
R8275 gnd.n6323 gnd.n796 19.3944
R8276 gnd.n6327 gnd.n796 19.3944
R8277 gnd.n6327 gnd.n792 19.3944
R8278 gnd.n6333 gnd.n792 19.3944
R8279 gnd.n6333 gnd.n790 19.3944
R8280 gnd.n6337 gnd.n790 19.3944
R8281 gnd.n6337 gnd.n786 19.3944
R8282 gnd.n6343 gnd.n786 19.3944
R8283 gnd.n6343 gnd.n784 19.3944
R8284 gnd.n6347 gnd.n784 19.3944
R8285 gnd.n6347 gnd.n780 19.3944
R8286 gnd.n6353 gnd.n780 19.3944
R8287 gnd.n6353 gnd.n778 19.3944
R8288 gnd.n6357 gnd.n778 19.3944
R8289 gnd.n6357 gnd.n774 19.3944
R8290 gnd.n6363 gnd.n774 19.3944
R8291 gnd.n6363 gnd.n772 19.3944
R8292 gnd.n6367 gnd.n772 19.3944
R8293 gnd.n6367 gnd.n768 19.3944
R8294 gnd.n6373 gnd.n768 19.3944
R8295 gnd.n6373 gnd.n766 19.3944
R8296 gnd.n6377 gnd.n766 19.3944
R8297 gnd.n6377 gnd.n762 19.3944
R8298 gnd.n6383 gnd.n762 19.3944
R8299 gnd.n6383 gnd.n760 19.3944
R8300 gnd.n6387 gnd.n760 19.3944
R8301 gnd.n6387 gnd.n756 19.3944
R8302 gnd.n6393 gnd.n756 19.3944
R8303 gnd.n6393 gnd.n754 19.3944
R8304 gnd.n6397 gnd.n754 19.3944
R8305 gnd.n6397 gnd.n750 19.3944
R8306 gnd.n6403 gnd.n750 19.3944
R8307 gnd.n6403 gnd.n748 19.3944
R8308 gnd.n6407 gnd.n748 19.3944
R8309 gnd.n6407 gnd.n744 19.3944
R8310 gnd.n6413 gnd.n744 19.3944
R8311 gnd.n6413 gnd.n742 19.3944
R8312 gnd.n6417 gnd.n742 19.3944
R8313 gnd.n6417 gnd.n738 19.3944
R8314 gnd.n6423 gnd.n738 19.3944
R8315 gnd.n6423 gnd.n736 19.3944
R8316 gnd.n6427 gnd.n736 19.3944
R8317 gnd.n6427 gnd.n732 19.3944
R8318 gnd.n6433 gnd.n732 19.3944
R8319 gnd.n6433 gnd.n730 19.3944
R8320 gnd.n6437 gnd.n730 19.3944
R8321 gnd.n6437 gnd.n726 19.3944
R8322 gnd.n6443 gnd.n726 19.3944
R8323 gnd.n6443 gnd.n724 19.3944
R8324 gnd.n6447 gnd.n724 19.3944
R8325 gnd.n6447 gnd.n720 19.3944
R8326 gnd.n6453 gnd.n720 19.3944
R8327 gnd.n6453 gnd.n718 19.3944
R8328 gnd.n6457 gnd.n718 19.3944
R8329 gnd.n6457 gnd.n714 19.3944
R8330 gnd.n6463 gnd.n714 19.3944
R8331 gnd.n6463 gnd.n712 19.3944
R8332 gnd.n6467 gnd.n712 19.3944
R8333 gnd.n6467 gnd.n708 19.3944
R8334 gnd.n6473 gnd.n708 19.3944
R8335 gnd.n6473 gnd.n706 19.3944
R8336 gnd.n6477 gnd.n706 19.3944
R8337 gnd.n6477 gnd.n702 19.3944
R8338 gnd.n6483 gnd.n702 19.3944
R8339 gnd.n6483 gnd.n700 19.3944
R8340 gnd.n6487 gnd.n700 19.3944
R8341 gnd.n6487 gnd.n696 19.3944
R8342 gnd.n6493 gnd.n696 19.3944
R8343 gnd.n6493 gnd.n694 19.3944
R8344 gnd.n6498 gnd.n694 19.3944
R8345 gnd.n6498 gnd.n690 19.3944
R8346 gnd.n6504 gnd.n690 19.3944
R8347 gnd.n6505 gnd.n6504 19.3944
R8348 gnd.n5650 gnd.n5649 19.3944
R8349 gnd.n5649 gnd.n5648 19.3944
R8350 gnd.n5648 gnd.n5647 19.3944
R8351 gnd.n5647 gnd.n5645 19.3944
R8352 gnd.n5645 gnd.n5642 19.3944
R8353 gnd.n5642 gnd.n5641 19.3944
R8354 gnd.n5641 gnd.n5638 19.3944
R8355 gnd.n5638 gnd.n5637 19.3944
R8356 gnd.n5637 gnd.n5634 19.3944
R8357 gnd.n5634 gnd.n5633 19.3944
R8358 gnd.n5633 gnd.n5630 19.3944
R8359 gnd.n5630 gnd.n5629 19.3944
R8360 gnd.n5629 gnd.n5626 19.3944
R8361 gnd.n5626 gnd.n5625 19.3944
R8362 gnd.n5625 gnd.n5622 19.3944
R8363 gnd.n5622 gnd.n5621 19.3944
R8364 gnd.n5621 gnd.n5618 19.3944
R8365 gnd.n5616 gnd.n5613 19.3944
R8366 gnd.n5613 gnd.n5612 19.3944
R8367 gnd.n5612 gnd.n5609 19.3944
R8368 gnd.n5609 gnd.n5608 19.3944
R8369 gnd.n5608 gnd.n5605 19.3944
R8370 gnd.n5605 gnd.n5604 19.3944
R8371 gnd.n5604 gnd.n5601 19.3944
R8372 gnd.n5599 gnd.n5596 19.3944
R8373 gnd.n5596 gnd.n5595 19.3944
R8374 gnd.n5595 gnd.n5592 19.3944
R8375 gnd.n5592 gnd.n5591 19.3944
R8376 gnd.n5591 gnd.n5588 19.3944
R8377 gnd.n5588 gnd.n5587 19.3944
R8378 gnd.n5587 gnd.n5584 19.3944
R8379 gnd.n5584 gnd.n5583 19.3944
R8380 gnd.n5579 gnd.n5576 19.3944
R8381 gnd.n5576 gnd.n5575 19.3944
R8382 gnd.n5575 gnd.n5572 19.3944
R8383 gnd.n5572 gnd.n5571 19.3944
R8384 gnd.n5571 gnd.n5568 19.3944
R8385 gnd.n5568 gnd.n5567 19.3944
R8386 gnd.n5567 gnd.n5564 19.3944
R8387 gnd.n5564 gnd.n5563 19.3944
R8388 gnd.n5563 gnd.n5560 19.3944
R8389 gnd.n5560 gnd.n5559 19.3944
R8390 gnd.n5559 gnd.n5556 19.3944
R8391 gnd.n5556 gnd.n5555 19.3944
R8392 gnd.n5555 gnd.n5552 19.3944
R8393 gnd.n5552 gnd.n5551 19.3944
R8394 gnd.n5551 gnd.n5548 19.3944
R8395 gnd.n5548 gnd.n5547 19.3944
R8396 gnd.n5547 gnd.n5544 19.3944
R8397 gnd.n5544 gnd.n5543 19.3944
R8398 gnd.n5527 gnd.n1556 19.3944
R8399 gnd.n5527 gnd.n5526 19.3944
R8400 gnd.n5526 gnd.n1565 19.3944
R8401 gnd.n5440 gnd.n1565 19.3944
R8402 gnd.n5443 gnd.n5440 19.3944
R8403 gnd.n5444 gnd.n5443 19.3944
R8404 gnd.n5446 gnd.n5444 19.3944
R8405 gnd.n5446 gnd.n1613 19.3944
R8406 gnd.n5501 gnd.n1613 19.3944
R8407 gnd.n5501 gnd.n1619 19.3944
R8408 gnd.n1619 gnd.n1618 19.3944
R8409 gnd.n1618 gnd.n1617 19.3944
R8410 gnd.n1617 gnd.n1614 19.3944
R8411 gnd.n1614 gnd.n528 19.3944
R8412 gnd.n6757 gnd.n528 19.3944
R8413 gnd.n6758 gnd.n6757 19.3944
R8414 gnd.n6759 gnd.n6758 19.3944
R8415 gnd.n6762 gnd.n6759 19.3944
R8416 gnd.n6762 gnd.n6760 19.3944
R8417 gnd.n6760 gnd.n501 19.3944
R8418 gnd.n6795 gnd.n501 19.3944
R8419 gnd.n6797 gnd.n6795 19.3944
R8420 gnd.n6797 gnd.n6796 19.3944
R8421 gnd.n6796 gnd.n494 19.3944
R8422 gnd.n6809 gnd.n494 19.3944
R8423 gnd.n6810 gnd.n6809 19.3944
R8424 gnd.n6812 gnd.n6810 19.3944
R8425 gnd.n6813 gnd.n6812 19.3944
R8426 gnd.n6816 gnd.n6813 19.3944
R8427 gnd.n6817 gnd.n6816 19.3944
R8428 gnd.n6819 gnd.n6817 19.3944
R8429 gnd.n6820 gnd.n6819 19.3944
R8430 gnd.n6823 gnd.n6820 19.3944
R8431 gnd.n6824 gnd.n6823 19.3944
R8432 gnd.n6826 gnd.n6824 19.3944
R8433 gnd.n6827 gnd.n6826 19.3944
R8434 gnd.n6830 gnd.n6827 19.3944
R8435 gnd.n6831 gnd.n6830 19.3944
R8436 gnd.n6833 gnd.n6831 19.3944
R8437 gnd.n6834 gnd.n6833 19.3944
R8438 gnd.n6836 gnd.n6834 19.3944
R8439 gnd.n6837 gnd.n6836 19.3944
R8440 gnd.n5530 gnd.n5529 19.3944
R8441 gnd.n5529 gnd.n1563 19.3944
R8442 gnd.n1587 gnd.n1563 19.3944
R8443 gnd.n5516 gnd.n1587 19.3944
R8444 gnd.n5516 gnd.n5515 19.3944
R8445 gnd.n5515 gnd.n5514 19.3944
R8446 gnd.n5514 gnd.n1592 19.3944
R8447 gnd.n5504 gnd.n1592 19.3944
R8448 gnd.n5504 gnd.n5503 19.3944
R8449 gnd.n5503 gnd.n552 19.3944
R8450 gnd.n6734 gnd.n552 19.3944
R8451 gnd.n6734 gnd.n6733 19.3944
R8452 gnd.n6733 gnd.n6732 19.3944
R8453 gnd.n6732 gnd.n6731 19.3944
R8454 gnd.n6731 gnd.n525 19.3944
R8455 gnd.n6767 gnd.n525 19.3944
R8456 gnd.n6767 gnd.n6766 19.3944
R8457 gnd.n6766 gnd.n6765 19.3944
R8458 gnd.n6765 gnd.n503 19.3944
R8459 gnd.n6792 gnd.n503 19.3944
R8460 gnd.n6792 gnd.n496 19.3944
R8461 gnd.n6801 gnd.n496 19.3944
R8462 gnd.n6802 gnd.n6801 19.3944
R8463 gnd.n6804 gnd.n6802 19.3944
R8464 gnd.n6804 gnd.n91 19.3944
R8465 gnd.n6887 gnd.n91 19.3944
R8466 gnd.n6887 gnd.n6886 19.3944
R8467 gnd.n6886 gnd.n6885 19.3944
R8468 gnd.n6885 gnd.n95 19.3944
R8469 gnd.n6875 gnd.n95 19.3944
R8470 gnd.n6875 gnd.n6874 19.3944
R8471 gnd.n6874 gnd.n6873 19.3944
R8472 gnd.n6873 gnd.n112 19.3944
R8473 gnd.n6863 gnd.n112 19.3944
R8474 gnd.n6863 gnd.n6862 19.3944
R8475 gnd.n6862 gnd.n6861 19.3944
R8476 gnd.n6861 gnd.n132 19.3944
R8477 gnd.n6851 gnd.n132 19.3944
R8478 gnd.n6851 gnd.n6850 19.3944
R8479 gnd.n6850 gnd.n6849 19.3944
R8480 gnd.n6849 gnd.n152 19.3944
R8481 gnd.n6839 gnd.n152 19.3944
R8482 gnd.n442 gnd.n302 19.3944
R8483 gnd.n446 gnd.n302 19.3944
R8484 gnd.n446 gnd.n300 19.3944
R8485 gnd.n452 gnd.n300 19.3944
R8486 gnd.n452 gnd.n298 19.3944
R8487 gnd.n456 gnd.n298 19.3944
R8488 gnd.n456 gnd.n296 19.3944
R8489 gnd.n462 gnd.n296 19.3944
R8490 gnd.n462 gnd.n294 19.3944
R8491 gnd.n466 gnd.n294 19.3944
R8492 gnd.n466 gnd.n292 19.3944
R8493 gnd.n472 gnd.n292 19.3944
R8494 gnd.n472 gnd.n290 19.3944
R8495 gnd.n476 gnd.n290 19.3944
R8496 gnd.n476 gnd.n288 19.3944
R8497 gnd.n482 gnd.n288 19.3944
R8498 gnd.n482 gnd.n286 19.3944
R8499 gnd.n486 gnd.n286 19.3944
R8500 gnd.n392 gnd.n324 19.3944
R8501 gnd.n396 gnd.n324 19.3944
R8502 gnd.n396 gnd.n322 19.3944
R8503 gnd.n402 gnd.n322 19.3944
R8504 gnd.n402 gnd.n320 19.3944
R8505 gnd.n406 gnd.n320 19.3944
R8506 gnd.n406 gnd.n318 19.3944
R8507 gnd.n412 gnd.n318 19.3944
R8508 gnd.n412 gnd.n316 19.3944
R8509 gnd.n416 gnd.n316 19.3944
R8510 gnd.n416 gnd.n314 19.3944
R8511 gnd.n422 gnd.n314 19.3944
R8512 gnd.n422 gnd.n312 19.3944
R8513 gnd.n426 gnd.n312 19.3944
R8514 gnd.n426 gnd.n310 19.3944
R8515 gnd.n432 gnd.n310 19.3944
R8516 gnd.n432 gnd.n308 19.3944
R8517 gnd.n436 gnd.n308 19.3944
R8518 gnd.n346 gnd.n345 19.3944
R8519 gnd.n351 gnd.n346 19.3944
R8520 gnd.n351 gnd.n342 19.3944
R8521 gnd.n355 gnd.n342 19.3944
R8522 gnd.n355 gnd.n340 19.3944
R8523 gnd.n361 gnd.n340 19.3944
R8524 gnd.n361 gnd.n338 19.3944
R8525 gnd.n365 gnd.n338 19.3944
R8526 gnd.n365 gnd.n336 19.3944
R8527 gnd.n371 gnd.n336 19.3944
R8528 gnd.n371 gnd.n334 19.3944
R8529 gnd.n375 gnd.n334 19.3944
R8530 gnd.n375 gnd.n332 19.3944
R8531 gnd.n382 gnd.n332 19.3944
R8532 gnd.n382 gnd.n330 19.3944
R8533 gnd.n386 gnd.n330 19.3944
R8534 gnd.n387 gnd.n386 19.3944
R8535 gnd.n279 gnd.n278 19.3944
R8536 gnd.n278 gnd.n277 19.3944
R8537 gnd.n277 gnd.n171 19.3944
R8538 gnd.n272 gnd.n171 19.3944
R8539 gnd.n272 gnd.n271 19.3944
R8540 gnd.n271 gnd.n270 19.3944
R8541 gnd.n270 gnd.n178 19.3944
R8542 gnd.n265 gnd.n178 19.3944
R8543 gnd.n265 gnd.n264 19.3944
R8544 gnd.n264 gnd.n263 19.3944
R8545 gnd.n263 gnd.n185 19.3944
R8546 gnd.n258 gnd.n185 19.3944
R8547 gnd.n258 gnd.n257 19.3944
R8548 gnd.n257 gnd.n256 19.3944
R8549 gnd.n256 gnd.n192 19.3944
R8550 gnd.n251 gnd.n192 19.3944
R8551 gnd.n5468 gnd.n1634 19.3944
R8552 gnd.n5468 gnd.n1635 19.3944
R8553 gnd.n5464 gnd.n1635 19.3944
R8554 gnd.n5464 gnd.n5463 19.3944
R8555 gnd.n5463 gnd.n5462 19.3944
R8556 gnd.n5462 gnd.n5438 19.3944
R8557 gnd.n5458 gnd.n5438 19.3944
R8558 gnd.n5458 gnd.n5457 19.3944
R8559 gnd.n5457 gnd.n5456 19.3944
R8560 gnd.n5456 gnd.n5451 19.3944
R8561 gnd.n5452 gnd.n5451 19.3944
R8562 gnd.n5452 gnd.n534 19.3944
R8563 gnd.n6749 gnd.n534 19.3944
R8564 gnd.n6749 gnd.n532 19.3944
R8565 gnd.n6753 gnd.n532 19.3944
R8566 gnd.n6753 gnd.n515 19.3944
R8567 gnd.n6776 gnd.n515 19.3944
R8568 gnd.n6776 gnd.n512 19.3944
R8569 gnd.n6780 gnd.n512 19.3944
R8570 gnd.n6780 gnd.n513 19.3944
R8571 gnd.n513 gnd.n64 19.3944
R8572 gnd.n6900 gnd.n64 19.3944
R8573 gnd.n6900 gnd.n6899 19.3944
R8574 gnd.n6899 gnd.n67 19.3944
R8575 gnd.n217 gnd.n67 19.3944
R8576 gnd.n218 gnd.n217 19.3944
R8577 gnd.n218 gnd.n213 19.3944
R8578 gnd.n222 gnd.n213 19.3944
R8579 gnd.n224 gnd.n222 19.3944
R8580 gnd.n225 gnd.n224 19.3944
R8581 gnd.n225 gnd.n210 19.3944
R8582 gnd.n229 gnd.n210 19.3944
R8583 gnd.n231 gnd.n229 19.3944
R8584 gnd.n232 gnd.n231 19.3944
R8585 gnd.n232 gnd.n207 19.3944
R8586 gnd.n236 gnd.n207 19.3944
R8587 gnd.n238 gnd.n236 19.3944
R8588 gnd.n239 gnd.n238 19.3944
R8589 gnd.n239 gnd.n204 19.3944
R8590 gnd.n243 gnd.n204 19.3944
R8591 gnd.n245 gnd.n243 19.3944
R8592 gnd.n246 gnd.n245 19.3944
R8593 gnd.n1573 gnd.n1572 19.3944
R8594 gnd.n5522 gnd.n1572 19.3944
R8595 gnd.n5522 gnd.n5521 19.3944
R8596 gnd.n5521 gnd.n5520 19.3944
R8597 gnd.n5520 gnd.n1579 19.3944
R8598 gnd.n5510 gnd.n1579 19.3944
R8599 gnd.n5510 gnd.n5509 19.3944
R8600 gnd.n5509 gnd.n5508 19.3944
R8601 gnd.n5508 gnd.n1604 19.3944
R8602 gnd.n1604 gnd.n544 19.3944
R8603 gnd.n6738 gnd.n544 19.3944
R8604 gnd.n6738 gnd.n542 19.3944
R8605 gnd.n6745 gnd.n542 19.3944
R8606 gnd.n6745 gnd.n6744 19.3944
R8607 gnd.n6744 gnd.n6743 19.3944
R8608 gnd.n6743 gnd.n521 19.3944
R8609 gnd.n6772 gnd.n6771 19.3944
R8610 gnd.n6788 gnd.n6787 19.3944
R8611 gnd.n6785 gnd.n6784 19.3944
R8612 gnd.n6895 gnd.n6894 19.3944
R8613 gnd.n6891 gnd.n75 19.3944
R8614 gnd.n6891 gnd.n82 19.3944
R8615 gnd.n6881 gnd.n82 19.3944
R8616 gnd.n6881 gnd.n6880 19.3944
R8617 gnd.n6880 gnd.n6879 19.3944
R8618 gnd.n6879 gnd.n104 19.3944
R8619 gnd.n6869 gnd.n104 19.3944
R8620 gnd.n6869 gnd.n6868 19.3944
R8621 gnd.n6868 gnd.n6867 19.3944
R8622 gnd.n6867 gnd.n122 19.3944
R8623 gnd.n6857 gnd.n122 19.3944
R8624 gnd.n6857 gnd.n6856 19.3944
R8625 gnd.n6856 gnd.n6855 19.3944
R8626 gnd.n6855 gnd.n142 19.3944
R8627 gnd.n6845 gnd.n142 19.3944
R8628 gnd.n6845 gnd.n6844 19.3944
R8629 gnd.n6844 gnd.n6843 19.3944
R8630 gnd.n4068 gnd.n4067 19.3944
R8631 gnd.n4067 gnd.n4066 19.3944
R8632 gnd.n4066 gnd.n4065 19.3944
R8633 gnd.n4065 gnd.n4063 19.3944
R8634 gnd.n4063 gnd.n4060 19.3944
R8635 gnd.n4060 gnd.n4059 19.3944
R8636 gnd.n4059 gnd.n4056 19.3944
R8637 gnd.n4056 gnd.n4055 19.3944
R8638 gnd.n4055 gnd.n4052 19.3944
R8639 gnd.n4052 gnd.n4051 19.3944
R8640 gnd.n4051 gnd.n4048 19.3944
R8641 gnd.n4048 gnd.n4047 19.3944
R8642 gnd.n4047 gnd.n4044 19.3944
R8643 gnd.n4044 gnd.n4043 19.3944
R8644 gnd.n4043 gnd.n4040 19.3944
R8645 gnd.n4040 gnd.n4039 19.3944
R8646 gnd.n4039 gnd.n4036 19.3944
R8647 gnd.n4034 gnd.n4031 19.3944
R8648 gnd.n4031 gnd.n4030 19.3944
R8649 gnd.n4030 gnd.n4027 19.3944
R8650 gnd.n4027 gnd.n4026 19.3944
R8651 gnd.n4026 gnd.n4023 19.3944
R8652 gnd.n4023 gnd.n4022 19.3944
R8653 gnd.n4022 gnd.n4019 19.3944
R8654 gnd.n4019 gnd.n4018 19.3944
R8655 gnd.n4018 gnd.n4015 19.3944
R8656 gnd.n4015 gnd.n4014 19.3944
R8657 gnd.n4014 gnd.n4011 19.3944
R8658 gnd.n4011 gnd.n4010 19.3944
R8659 gnd.n4010 gnd.n4007 19.3944
R8660 gnd.n4007 gnd.n4006 19.3944
R8661 gnd.n4006 gnd.n4003 19.3944
R8662 gnd.n4003 gnd.n4002 19.3944
R8663 gnd.n4002 gnd.n3999 19.3944
R8664 gnd.n3999 gnd.n3998 19.3944
R8665 gnd.n3994 gnd.n3991 19.3944
R8666 gnd.n3991 gnd.n3990 19.3944
R8667 gnd.n3990 gnd.n3987 19.3944
R8668 gnd.n3987 gnd.n3986 19.3944
R8669 gnd.n3986 gnd.n3983 19.3944
R8670 gnd.n3983 gnd.n3982 19.3944
R8671 gnd.n3982 gnd.n3979 19.3944
R8672 gnd.n3979 gnd.n3978 19.3944
R8673 gnd.n3978 gnd.n3975 19.3944
R8674 gnd.n3975 gnd.n3974 19.3944
R8675 gnd.n3974 gnd.n3971 19.3944
R8676 gnd.n3971 gnd.n3970 19.3944
R8677 gnd.n3970 gnd.n3967 19.3944
R8678 gnd.n3967 gnd.n3966 19.3944
R8679 gnd.n3966 gnd.n3963 19.3944
R8680 gnd.n3963 gnd.n3962 19.3944
R8681 gnd.n3962 gnd.n3959 19.3944
R8682 gnd.n3959 gnd.n3958 19.3944
R8683 gnd.n3951 gnd.n3949 19.3944
R8684 gnd.n3949 gnd.n3946 19.3944
R8685 gnd.n3946 gnd.n3945 19.3944
R8686 gnd.n3945 gnd.n3942 19.3944
R8687 gnd.n3942 gnd.n3941 19.3944
R8688 gnd.n3941 gnd.n3938 19.3944
R8689 gnd.n3938 gnd.n3937 19.3944
R8690 gnd.n3937 gnd.n3934 19.3944
R8691 gnd.n3934 gnd.n3933 19.3944
R8692 gnd.n3933 gnd.n3930 19.3944
R8693 gnd.n3930 gnd.n3929 19.3944
R8694 gnd.n3929 gnd.n3926 19.3944
R8695 gnd.n3926 gnd.n3925 19.3944
R8696 gnd.n3925 gnd.n3922 19.3944
R8697 gnd.n3922 gnd.n3921 19.3944
R8698 gnd.n3921 gnd.n3918 19.3944
R8699 gnd.n3912 gnd.n3910 19.3944
R8700 gnd.n3910 gnd.n3909 19.3944
R8701 gnd.n3909 gnd.n3907 19.3944
R8702 gnd.n3907 gnd.n3906 19.3944
R8703 gnd.n3906 gnd.n3904 19.3944
R8704 gnd.n3904 gnd.n3903 19.3944
R8705 gnd.n3903 gnd.n3901 19.3944
R8706 gnd.n3901 gnd.n3900 19.3944
R8707 gnd.n3900 gnd.n3898 19.3944
R8708 gnd.n3898 gnd.n3897 19.3944
R8709 gnd.n3897 gnd.n3895 19.3944
R8710 gnd.n3895 gnd.n3894 19.3944
R8711 gnd.n3894 gnd.n3892 19.3944
R8712 gnd.n3892 gnd.n3891 19.3944
R8713 gnd.n3891 gnd.n3889 19.3944
R8714 gnd.n3889 gnd.n3888 19.3944
R8715 gnd.n3888 gnd.n3886 19.3944
R8716 gnd.n3886 gnd.n3885 19.3944
R8717 gnd.n3885 gnd.n3883 19.3944
R8718 gnd.n3883 gnd.n3882 19.3944
R8719 gnd.n3882 gnd.n3880 19.3944
R8720 gnd.n3880 gnd.n3877 19.3944
R8721 gnd.n3877 gnd.n2162 19.3944
R8722 gnd.n4200 gnd.n2162 19.3944
R8723 gnd.n4200 gnd.n2160 19.3944
R8724 gnd.n4204 gnd.n2160 19.3944
R8725 gnd.n4204 gnd.n2155 19.3944
R8726 gnd.n4223 gnd.n2155 19.3944
R8727 gnd.n4223 gnd.n2156 19.3944
R8728 gnd.n4219 gnd.n2156 19.3944
R8729 gnd.n4219 gnd.n2147 19.3944
R8730 gnd.n4254 gnd.n2147 19.3944
R8731 gnd.n4254 gnd.n2145 19.3944
R8732 gnd.n4258 gnd.n2145 19.3944
R8733 gnd.n4258 gnd.n2138 19.3944
R8734 gnd.n4540 gnd.n2138 19.3944
R8735 gnd.n4540 gnd.n2139 19.3944
R8736 gnd.n4536 gnd.n2139 19.3944
R8737 gnd.n4536 gnd.n4535 19.3944
R8738 gnd.n4535 gnd.n4534 19.3944
R8739 gnd.n4534 gnd.n4531 19.3944
R8740 gnd.n4531 gnd.n2125 19.3944
R8741 gnd.n4077 gnd.n4075 19.3944
R8742 gnd.n4077 gnd.n4076 19.3944
R8743 gnd.n4076 gnd.n2249 19.3944
R8744 gnd.n4092 gnd.n2249 19.3944
R8745 gnd.n4093 gnd.n4092 19.3944
R8746 gnd.n4094 gnd.n4093 19.3944
R8747 gnd.n4094 gnd.n2231 19.3944
R8748 gnd.n4112 gnd.n2231 19.3944
R8749 gnd.n4113 gnd.n4112 19.3944
R8750 gnd.n4114 gnd.n4113 19.3944
R8751 gnd.n4114 gnd.n2213 19.3944
R8752 gnd.n4132 gnd.n2213 19.3944
R8753 gnd.n4133 gnd.n4132 19.3944
R8754 gnd.n4134 gnd.n4133 19.3944
R8755 gnd.n4134 gnd.n2195 19.3944
R8756 gnd.n4153 gnd.n2195 19.3944
R8757 gnd.n4154 gnd.n4153 19.3944
R8758 gnd.n4155 gnd.n4154 19.3944
R8759 gnd.n4155 gnd.n2179 19.3944
R8760 gnd.n4173 gnd.n2179 19.3944
R8761 gnd.n4174 gnd.n4173 19.3944
R8762 gnd.n4176 gnd.n4174 19.3944
R8763 gnd.n4177 gnd.n4176 19.3944
R8764 gnd.n4179 gnd.n4177 19.3944
R8765 gnd.n4179 gnd.n2158 19.3944
R8766 gnd.n4208 gnd.n2158 19.3944
R8767 gnd.n4209 gnd.n4208 19.3944
R8768 gnd.n4210 gnd.n4209 19.3944
R8769 gnd.n4211 gnd.n4210 19.3944
R8770 gnd.n4215 gnd.n4211 19.3944
R8771 gnd.n4215 gnd.n4214 19.3944
R8772 gnd.n4214 gnd.n4213 19.3944
R8773 gnd.n4213 gnd.n2143 19.3944
R8774 gnd.n4262 gnd.n2143 19.3944
R8775 gnd.n4263 gnd.n4262 19.3944
R8776 gnd.n4264 gnd.n4263 19.3944
R8777 gnd.n4265 gnd.n4264 19.3944
R8778 gnd.n4269 gnd.n4265 19.3944
R8779 gnd.n4270 gnd.n4269 19.3944
R8780 gnd.n4527 gnd.n4270 19.3944
R8781 gnd.n4527 gnd.n4526 19.3944
R8782 gnd.n4526 gnd.n4525 19.3944
R8783 gnd.n4079 gnd.n2265 19.3944
R8784 gnd.n4079 gnd.n2266 19.3944
R8785 gnd.n2268 gnd.n2266 19.3944
R8786 gnd.n2268 gnd.n2247 19.3944
R8787 gnd.n4099 gnd.n2247 19.3944
R8788 gnd.n4099 gnd.n4098 19.3944
R8789 gnd.n4098 gnd.n4097 19.3944
R8790 gnd.n4097 gnd.n2229 19.3944
R8791 gnd.n4119 gnd.n2229 19.3944
R8792 gnd.n4119 gnd.n4118 19.3944
R8793 gnd.n4118 gnd.n4117 19.3944
R8794 gnd.n4117 gnd.n2211 19.3944
R8795 gnd.n4139 gnd.n2211 19.3944
R8796 gnd.n4139 gnd.n4138 19.3944
R8797 gnd.n4138 gnd.n4137 19.3944
R8798 gnd.n4137 gnd.n2193 19.3944
R8799 gnd.n4160 gnd.n2193 19.3944
R8800 gnd.n4160 gnd.n4159 19.3944
R8801 gnd.n4159 gnd.n4158 19.3944
R8802 gnd.n4158 gnd.n2175 19.3944
R8803 gnd.n4187 gnd.n2175 19.3944
R8804 gnd.n4187 gnd.n4186 19.3944
R8805 gnd.n4186 gnd.n4185 19.3944
R8806 gnd.n4185 gnd.n4184 19.3944
R8807 gnd.n4184 gnd.n4182 19.3944
R8808 gnd.n4182 gnd.n1067 19.3944
R8809 gnd.n6004 gnd.n1067 19.3944
R8810 gnd.n6004 gnd.n6003 19.3944
R8811 gnd.n6003 gnd.n6002 19.3944
R8812 gnd.n6002 gnd.n1071 19.3944
R8813 gnd.n5992 gnd.n1071 19.3944
R8814 gnd.n5992 gnd.n5991 19.3944
R8815 gnd.n5991 gnd.n5990 19.3944
R8816 gnd.n5990 gnd.n1092 19.3944
R8817 gnd.n5980 gnd.n1092 19.3944
R8818 gnd.n5980 gnd.n5979 19.3944
R8819 gnd.n5979 gnd.n5978 19.3944
R8820 gnd.n5978 gnd.n1111 19.3944
R8821 gnd.n5968 gnd.n1111 19.3944
R8822 gnd.n5968 gnd.n5967 19.3944
R8823 gnd.n5967 gnd.n5966 19.3944
R8824 gnd.n5966 gnd.n1132 19.3944
R8825 gnd.n5958 gnd.n1142 19.3944
R8826 gnd.n5953 gnd.n1142 19.3944
R8827 gnd.n5953 gnd.n5952 19.3944
R8828 gnd.n5952 gnd.n5951 19.3944
R8829 gnd.n5951 gnd.n5948 19.3944
R8830 gnd.n5948 gnd.n5947 19.3944
R8831 gnd.n5947 gnd.n5944 19.3944
R8832 gnd.n5944 gnd.n5943 19.3944
R8833 gnd.n5943 gnd.n5940 19.3944
R8834 gnd.n5940 gnd.n5939 19.3944
R8835 gnd.n5939 gnd.n5936 19.3944
R8836 gnd.n5936 gnd.n5935 19.3944
R8837 gnd.n5935 gnd.n5932 19.3944
R8838 gnd.n5932 gnd.n5931 19.3944
R8839 gnd.n5931 gnd.n5928 19.3944
R8840 gnd.n5928 gnd.n5927 19.3944
R8841 gnd.n5927 gnd.n5924 19.3944
R8842 gnd.n4473 gnd.n4439 19.3944
R8843 gnd.n4477 gnd.n4439 19.3944
R8844 gnd.n4480 gnd.n4477 19.3944
R8845 gnd.n4483 gnd.n4480 19.3944
R8846 gnd.n4483 gnd.n4437 19.3944
R8847 gnd.n4487 gnd.n4437 19.3944
R8848 gnd.n4490 gnd.n4487 19.3944
R8849 gnd.n4493 gnd.n4490 19.3944
R8850 gnd.n4493 gnd.n4435 19.3944
R8851 gnd.n4497 gnd.n4435 19.3944
R8852 gnd.n4500 gnd.n4497 19.3944
R8853 gnd.n4503 gnd.n4500 19.3944
R8854 gnd.n4503 gnd.n4433 19.3944
R8855 gnd.n4507 gnd.n4433 19.3944
R8856 gnd.n4510 gnd.n4507 19.3944
R8857 gnd.n4513 gnd.n4510 19.3944
R8858 gnd.n4513 gnd.n4431 19.3944
R8859 gnd.n4518 gnd.n4431 19.3944
R8860 gnd.n4451 gnd.n1211 19.3944
R8861 gnd.n4454 gnd.n4451 19.3944
R8862 gnd.n4454 gnd.n4446 19.3944
R8863 gnd.n4458 gnd.n4446 19.3944
R8864 gnd.n4461 gnd.n4458 19.3944
R8865 gnd.n4464 gnd.n4461 19.3944
R8866 gnd.n4464 gnd.n4444 19.3944
R8867 gnd.n4469 gnd.n4444 19.3944
R8868 gnd.n5922 gnd.n5919 19.3944
R8869 gnd.n5919 gnd.n5918 19.3944
R8870 gnd.n5918 gnd.n5915 19.3944
R8871 gnd.n5915 gnd.n5914 19.3944
R8872 gnd.n5914 gnd.n5911 19.3944
R8873 gnd.n5911 gnd.n5910 19.3944
R8874 gnd.n5910 gnd.n5907 19.3944
R8875 gnd.n4083 gnd.n2258 19.3944
R8876 gnd.n4083 gnd.n2256 19.3944
R8877 gnd.n4087 gnd.n2256 19.3944
R8878 gnd.n4087 gnd.n2239 19.3944
R8879 gnd.n4103 gnd.n2239 19.3944
R8880 gnd.n4103 gnd.n2237 19.3944
R8881 gnd.n4107 gnd.n2237 19.3944
R8882 gnd.n4107 gnd.n2222 19.3944
R8883 gnd.n4123 gnd.n2222 19.3944
R8884 gnd.n4123 gnd.n2220 19.3944
R8885 gnd.n4127 gnd.n2220 19.3944
R8886 gnd.n4127 gnd.n2203 19.3944
R8887 gnd.n4143 gnd.n2203 19.3944
R8888 gnd.n4143 gnd.n2201 19.3944
R8889 gnd.n4148 gnd.n2201 19.3944
R8890 gnd.n4148 gnd.n4147 19.3944
R8891 gnd.n4165 gnd.n4164 19.3944
R8892 gnd.n4168 gnd.n4167 19.3944
R8893 gnd.n4192 gnd.n4191 19.3944
R8894 gnd.n4195 gnd.n4194 19.3944
R8895 gnd.n6010 gnd.n6009 19.3944
R8896 gnd.n6009 gnd.n6008 19.3944
R8897 gnd.n6008 gnd.n1060 19.3944
R8898 gnd.n5998 gnd.n1060 19.3944
R8899 gnd.n5998 gnd.n5997 19.3944
R8900 gnd.n5997 gnd.n5996 19.3944
R8901 gnd.n5996 gnd.n1082 19.3944
R8902 gnd.n5986 gnd.n1082 19.3944
R8903 gnd.n5986 gnd.n5985 19.3944
R8904 gnd.n5985 gnd.n5984 19.3944
R8905 gnd.n5984 gnd.n1102 19.3944
R8906 gnd.n5974 gnd.n1102 19.3944
R8907 gnd.n5974 gnd.n5973 19.3944
R8908 gnd.n5973 gnd.n5972 19.3944
R8909 gnd.n5972 gnd.n1122 19.3944
R8910 gnd.n5962 gnd.n1122 19.3944
R8911 gnd.n5962 gnd.n5961 19.3944
R8912 gnd.n6183 gnd.n882 19.3944
R8913 gnd.n6177 gnd.n882 19.3944
R8914 gnd.n6177 gnd.n6176 19.3944
R8915 gnd.n6176 gnd.n6175 19.3944
R8916 gnd.n6175 gnd.n889 19.3944
R8917 gnd.n6169 gnd.n889 19.3944
R8918 gnd.n6169 gnd.n6168 19.3944
R8919 gnd.n6168 gnd.n6167 19.3944
R8920 gnd.n6167 gnd.n897 19.3944
R8921 gnd.n6161 gnd.n897 19.3944
R8922 gnd.n6161 gnd.n6160 19.3944
R8923 gnd.n6160 gnd.n6159 19.3944
R8924 gnd.n6159 gnd.n905 19.3944
R8925 gnd.n6153 gnd.n905 19.3944
R8926 gnd.n6153 gnd.n6152 19.3944
R8927 gnd.n6152 gnd.n6151 19.3944
R8928 gnd.n6151 gnd.n913 19.3944
R8929 gnd.n6145 gnd.n913 19.3944
R8930 gnd.n6145 gnd.n6144 19.3944
R8931 gnd.n6144 gnd.n6143 19.3944
R8932 gnd.n6143 gnd.n921 19.3944
R8933 gnd.n6137 gnd.n921 19.3944
R8934 gnd.n6137 gnd.n6136 19.3944
R8935 gnd.n6136 gnd.n6135 19.3944
R8936 gnd.n6135 gnd.n929 19.3944
R8937 gnd.n6129 gnd.n929 19.3944
R8938 gnd.n6129 gnd.n6128 19.3944
R8939 gnd.n6128 gnd.n6127 19.3944
R8940 gnd.n6127 gnd.n937 19.3944
R8941 gnd.n6121 gnd.n937 19.3944
R8942 gnd.n6121 gnd.n6120 19.3944
R8943 gnd.n6120 gnd.n6119 19.3944
R8944 gnd.n6119 gnd.n945 19.3944
R8945 gnd.n6113 gnd.n945 19.3944
R8946 gnd.n6113 gnd.n6112 19.3944
R8947 gnd.n6112 gnd.n6111 19.3944
R8948 gnd.n6111 gnd.n953 19.3944
R8949 gnd.n6105 gnd.n953 19.3944
R8950 gnd.n6105 gnd.n6104 19.3944
R8951 gnd.n6104 gnd.n6103 19.3944
R8952 gnd.n6103 gnd.n961 19.3944
R8953 gnd.n6097 gnd.n961 19.3944
R8954 gnd.n6097 gnd.n6096 19.3944
R8955 gnd.n6096 gnd.n6095 19.3944
R8956 gnd.n6095 gnd.n969 19.3944
R8957 gnd.n6089 gnd.n969 19.3944
R8958 gnd.n6089 gnd.n6088 19.3944
R8959 gnd.n6088 gnd.n6087 19.3944
R8960 gnd.n6087 gnd.n977 19.3944
R8961 gnd.n6081 gnd.n977 19.3944
R8962 gnd.n6081 gnd.n6080 19.3944
R8963 gnd.n6080 gnd.n6079 19.3944
R8964 gnd.n6079 gnd.n985 19.3944
R8965 gnd.n6073 gnd.n985 19.3944
R8966 gnd.n6073 gnd.n6072 19.3944
R8967 gnd.n6072 gnd.n6071 19.3944
R8968 gnd.n6071 gnd.n993 19.3944
R8969 gnd.n6065 gnd.n993 19.3944
R8970 gnd.n6065 gnd.n6064 19.3944
R8971 gnd.n6064 gnd.n6063 19.3944
R8972 gnd.n6063 gnd.n1001 19.3944
R8973 gnd.n6057 gnd.n1001 19.3944
R8974 gnd.n6057 gnd.n6056 19.3944
R8975 gnd.n6056 gnd.n6055 19.3944
R8976 gnd.n6055 gnd.n1009 19.3944
R8977 gnd.n6049 gnd.n1009 19.3944
R8978 gnd.n6049 gnd.n6048 19.3944
R8979 gnd.n6048 gnd.n6047 19.3944
R8980 gnd.n6047 gnd.n1017 19.3944
R8981 gnd.n6041 gnd.n1017 19.3944
R8982 gnd.n6041 gnd.n6040 19.3944
R8983 gnd.n6040 gnd.n6039 19.3944
R8984 gnd.n6039 gnd.n1025 19.3944
R8985 gnd.n6033 gnd.n1025 19.3944
R8986 gnd.n6033 gnd.n6032 19.3944
R8987 gnd.n6032 gnd.n6031 19.3944
R8988 gnd.n6031 gnd.n1033 19.3944
R8989 gnd.n6025 gnd.n1033 19.3944
R8990 gnd.n6025 gnd.n6024 19.3944
R8991 gnd.n6024 gnd.n6023 19.3944
R8992 gnd.n6023 gnd.n1041 19.3944
R8993 gnd.n6017 gnd.n1041 19.3944
R8994 gnd.n6017 gnd.n6016 19.3944
R8995 gnd.n6016 gnd.n6015 19.3944
R8996 gnd.n4296 gnd.n4278 19.3944
R8997 gnd.n4292 gnd.n4278 19.3944
R8998 gnd.n4292 gnd.n4291 19.3944
R8999 gnd.n4291 gnd.n4290 19.3944
R9000 gnd.n4290 gnd.n4282 19.3944
R9001 gnd.n4286 gnd.n4282 19.3944
R9002 gnd.n4286 gnd.n4285 19.3944
R9003 gnd.n4285 gnd.n2062 19.3944
R9004 gnd.n4648 gnd.n2062 19.3944
R9005 gnd.n4648 gnd.n2060 19.3944
R9006 gnd.n4652 gnd.n2060 19.3944
R9007 gnd.n4652 gnd.n2058 19.3944
R9008 gnd.n4656 gnd.n2058 19.3944
R9009 gnd.n4656 gnd.n2055 19.3944
R9010 gnd.n4669 gnd.n2055 19.3944
R9011 gnd.n4669 gnd.n2056 19.3944
R9012 gnd.n4665 gnd.n2056 19.3944
R9013 gnd.n4665 gnd.n4664 19.3944
R9014 gnd.n4664 gnd.n4663 19.3944
R9015 gnd.n4663 gnd.n2024 19.3944
R9016 gnd.n4808 gnd.n2024 19.3944
R9017 gnd.n4808 gnd.n2021 19.3944
R9018 gnd.n4815 gnd.n2021 19.3944
R9019 gnd.n4815 gnd.n2022 19.3944
R9020 gnd.n4811 gnd.n2022 19.3944
R9021 gnd.n4811 gnd.n2003 19.3944
R9022 gnd.n4839 gnd.n2003 19.3944
R9023 gnd.n4839 gnd.n2000 19.3944
R9024 gnd.n4849 gnd.n2000 19.3944
R9025 gnd.n4849 gnd.n2001 19.3944
R9026 gnd.n4845 gnd.n2001 19.3944
R9027 gnd.n4845 gnd.n4844 19.3944
R9028 gnd.n4844 gnd.n1953 19.3944
R9029 gnd.n4919 gnd.n1953 19.3944
R9030 gnd.n4919 gnd.n1950 19.3944
R9031 gnd.n4924 gnd.n1950 19.3944
R9032 gnd.n4924 gnd.n1951 19.3944
R9033 gnd.n1951 gnd.n1926 19.3944
R9034 gnd.n4965 gnd.n1926 19.3944
R9035 gnd.n4965 gnd.n1923 19.3944
R9036 gnd.n4995 gnd.n1923 19.3944
R9037 gnd.n4995 gnd.n1924 19.3944
R9038 gnd.n4991 gnd.n1924 19.3944
R9039 gnd.n4991 gnd.n4990 19.3944
R9040 gnd.n4990 gnd.n4989 19.3944
R9041 gnd.n4989 gnd.n4973 19.3944
R9042 gnd.n4985 gnd.n4973 19.3944
R9043 gnd.n4985 gnd.n4984 19.3944
R9044 gnd.n4984 gnd.n4983 19.3944
R9045 gnd.n4983 gnd.n4978 19.3944
R9046 gnd.n4979 gnd.n4978 19.3944
R9047 gnd.n4979 gnd.n1851 19.3944
R9048 gnd.n5098 gnd.n1851 19.3944
R9049 gnd.n5098 gnd.n1848 19.3944
R9050 gnd.n5135 gnd.n1848 19.3944
R9051 gnd.n5135 gnd.n1849 19.3944
R9052 gnd.n5131 gnd.n1849 19.3944
R9053 gnd.n5131 gnd.n5130 19.3944
R9054 gnd.n5130 gnd.n5129 19.3944
R9055 gnd.n5129 gnd.n5106 19.3944
R9056 gnd.n5125 gnd.n5106 19.3944
R9057 gnd.n5125 gnd.n5124 19.3944
R9058 gnd.n5124 gnd.n5123 19.3944
R9059 gnd.n5123 gnd.n5110 19.3944
R9060 gnd.n5119 gnd.n5110 19.3944
R9061 gnd.n5119 gnd.n5118 19.3944
R9062 gnd.n5118 gnd.n5117 19.3944
R9063 gnd.n5117 gnd.n5114 19.3944
R9064 gnd.n5114 gnd.n1698 19.3944
R9065 gnd.n5361 gnd.n1698 19.3944
R9066 gnd.n5361 gnd.n1696 19.3944
R9067 gnd.n5365 gnd.n1696 19.3944
R9068 gnd.n5365 gnd.n1685 19.3944
R9069 gnd.n5377 gnd.n1685 19.3944
R9070 gnd.n5377 gnd.n1683 19.3944
R9071 gnd.n5381 gnd.n1683 19.3944
R9072 gnd.n5381 gnd.n1673 19.3944
R9073 gnd.n5396 gnd.n1673 19.3944
R9074 gnd.n5396 gnd.n1671 19.3944
R9075 gnd.n5400 gnd.n1671 19.3944
R9076 gnd.n5400 gnd.n1383 19.3944
R9077 gnd.n5719 gnd.n1383 19.3944
R9078 gnd.n5716 gnd.n5715 19.3944
R9079 gnd.n5715 gnd.n5714 19.3944
R9080 gnd.n5714 gnd.n1388 19.3944
R9081 gnd.n5710 gnd.n1388 19.3944
R9082 gnd.n5710 gnd.n5709 19.3944
R9083 gnd.n5709 gnd.n5708 19.3944
R9084 gnd.n5708 gnd.n1393 19.3944
R9085 gnd.n5703 gnd.n1393 19.3944
R9086 gnd.n5703 gnd.n5702 19.3944
R9087 gnd.n5702 gnd.n1398 19.3944
R9088 gnd.n5695 gnd.n1398 19.3944
R9089 gnd.n5695 gnd.n5694 19.3944
R9090 gnd.n5694 gnd.n1407 19.3944
R9091 gnd.n5687 gnd.n1407 19.3944
R9092 gnd.n5687 gnd.n5686 19.3944
R9093 gnd.n5686 gnd.n1415 19.3944
R9094 gnd.n5679 gnd.n1415 19.3944
R9095 gnd.n5679 gnd.n5678 19.3944
R9096 gnd.n5678 gnd.n1423 19.3944
R9097 gnd.n5671 gnd.n1423 19.3944
R9098 gnd.n5671 gnd.n5670 19.3944
R9099 gnd.n5670 gnd.n1431 19.3944
R9100 gnd.n5663 gnd.n1431 19.3944
R9101 gnd.n5663 gnd.n5662 19.3944
R9102 gnd.n1659 gnd.n1638 19.3944
R9103 gnd.n5430 gnd.n1638 19.3944
R9104 gnd.n5430 gnd.n5429 19.3944
R9105 gnd.t17 gnd.n2026 19.1199
R9106 gnd.t35 gnd.n5167 19.1199
R9107 gnd.n3121 gnd.t27 18.8012
R9108 gnd.n3106 gnd.t49 18.8012
R9109 gnd.n5902 gnd.n1218 18.8012
R9110 gnd.n5836 gnd.n5835 18.5761
R9111 gnd.n5347 gnd.n5346 18.5761
R9112 gnd.n2965 gnd.n2964 18.4825
R9113 gnd.t212 gnd.n1250 18.4825
R9114 gnd.n4672 gnd.t302 18.4825
R9115 gnd.n4818 gnd.t31 18.4825
R9116 gnd.n4927 gnd.n4926 18.4825
R9117 gnd.n1899 gnd.n1893 18.4825
R9118 gnd.n5160 gnd.t34 18.4825
R9119 gnd.n5184 gnd.n1806 18.4825
R9120 gnd.n5601 gnd.n5600 18.4247
R9121 gnd.n5907 gnd.n5906 18.4247
R9122 gnd.n5659 gnd.n5658 18.2308
R9123 gnd.n4378 gnd.n2124 18.2308
R9124 gnd.n251 gnd.n250 18.2308
R9125 gnd.n3918 gnd.n3856 18.2308
R9126 gnd.t4 gnd.n2645 18.1639
R9127 gnd.n2673 gnd.t60 17.5266
R9128 gnd.n3349 gnd.n3348 17.2079
R9129 gnd.n5832 gnd.n5831 17.2079
R9130 gnd.n2051 gnd.n2050 17.2079
R9131 gnd.n5203 gnd.n1802 17.2079
R9132 gnd.n5351 gnd.n5350 17.2079
R9133 gnd.n3072 gnd.t67 16.8893
R9134 gnd.n4081 gnd.t208 16.8893
R9135 gnd.t108 gnd.n1084 16.8893
R9136 gnd.t81 gnd.n549 16.8893
R9137 gnd.n162 gnd.t215 16.8893
R9138 gnd.n5583 gnd.n5580 16.6793
R9139 gnd.n436 gnd.n306 16.6793
R9140 gnd.n3998 gnd.n3995 16.6793
R9141 gnd.n4470 gnd.n4469 16.6793
R9142 gnd.n2900 gnd.t318 16.2519
R9143 gnd.n2600 gnd.t2 16.2519
R9144 gnd.n4588 gnd.t270 16.2519
R9145 gnd.t244 gnd.n1378 16.2519
R9146 gnd.n4748 gnd.n4671 15.9333
R9147 gnd.n4907 gnd.n4906 15.9333
R9148 gnd.n1880 gnd.n1873 15.9333
R9149 gnd.n1793 gnd.n1787 15.9333
R9150 gnd.n3588 gnd.n3586 15.6674
R9151 gnd.n3556 gnd.n3554 15.6674
R9152 gnd.n3524 gnd.n3522 15.6674
R9153 gnd.n3493 gnd.n3491 15.6674
R9154 gnd.n3461 gnd.n3459 15.6674
R9155 gnd.n3429 gnd.n3427 15.6674
R9156 gnd.n3397 gnd.n3395 15.6674
R9157 gnd.n3366 gnd.n3364 15.6674
R9158 gnd.n2891 gnd.t318 15.6146
R9159 gnd.t311 gnd.n2354 15.6146
R9160 gnd.t295 gnd.n2355 15.6146
R9161 gnd.t270 gnd.n2089 15.6146
R9162 gnd.n5402 gnd.t244 15.6146
R9163 gnd.n5540 gnd.n5535 15.3217
R9164 gnd.n491 gnd.n284 15.3217
R9165 gnd.n3956 gnd.n2271 15.3217
R9166 gnd.n4521 gnd.n4519 15.3217
R9167 gnd.t23 gnd.n1994 15.296
R9168 gnd.n5137 gnd.t21 15.296
R9169 gnd.n1720 gnd.n1719 15.0827
R9170 gnd.n1262 gnd.n1257 15.0481
R9171 gnd.n1730 gnd.n1729 15.0481
R9172 gnd.n3259 gnd.t59 14.9773
R9173 gnd.t208 gnd.n2252 14.9773
R9174 gnd.n4529 gnd.t240 14.9773
R9175 gnd.n4899 gnd.t10 14.9773
R9176 gnd.n5041 gnd.t53 14.9773
R9177 gnd.n5524 gnd.t219 14.9773
R9178 gnd.n6847 gnd.t215 14.9773
R9179 gnd.n5832 gnd.n1276 14.6587
R9180 gnd.n4875 gnd.n1982 14.6587
R9181 gnd.n5085 gnd.n1864 14.6587
R9182 gnd.n5204 gnd.n5203 14.6587
R9183 gnd.t41 gnd.n2397 14.34
R9184 gnd.n3337 gnd.t3 14.34
R9185 gnd.t254 gnd.n2044 14.0214
R9186 gnd.n5190 gnd.t230 14.0214
R9187 gnd.t277 gnd.n1701 14.0214
R9188 gnd.n3047 gnd.t45 13.7027
R9189 gnd.n2757 gnd.n2756 13.5763
R9190 gnd.n3702 gnd.n2311 13.5763
R9191 gnd.n2965 gnd.n2703 13.384
R9192 gnd.n4795 gnd.n2039 13.384
R9193 gnd.n4867 gnd.n4866 13.384
R9194 gnd.n4852 gnd.t5 13.384
R9195 gnd.n5096 gnd.t20 13.384
R9196 gnd.n5078 gnd.n5077 13.384
R9197 gnd.n5184 gnd.n5183 13.384
R9198 gnd.n1273 gnd.n1254 13.1884
R9199 gnd.n1268 gnd.n1267 13.1884
R9200 gnd.n1267 gnd.n1266 13.1884
R9201 gnd.n1723 gnd.n1718 13.1884
R9202 gnd.n1724 gnd.n1723 13.1884
R9203 gnd.n1269 gnd.n1256 13.146
R9204 gnd.n1265 gnd.n1256 13.146
R9205 gnd.n1722 gnd.n1721 13.146
R9206 gnd.n1722 gnd.n1717 13.146
R9207 gnd.n5902 gnd.n1250 13.0654
R9208 gnd.n5212 gnd.t63 13.0654
R9209 gnd.n5359 gnd.n1702 13.0654
R9210 gnd.n3589 gnd.n3585 12.8005
R9211 gnd.n3557 gnd.n3553 12.8005
R9212 gnd.n3525 gnd.n3521 12.8005
R9213 gnd.n3494 gnd.n3490 12.8005
R9214 gnd.n3462 gnd.n3458 12.8005
R9215 gnd.n3430 gnd.n3426 12.8005
R9216 gnd.n3398 gnd.n3394 12.8005
R9217 gnd.n3367 gnd.n3363 12.8005
R9218 gnd.n2756 gnd.n2751 12.4126
R9219 gnd.n3705 gnd.n3702 12.4126
R9220 gnd.n5899 gnd.n5836 12.1761
R9221 gnd.n5346 gnd.n5345 12.1761
R9222 gnd.n4759 gnd.n2027 12.1094
R9223 gnd.n4836 gnd.n2006 12.1094
R9224 gnd.n5145 gnd.n1838 12.1094
R9225 gnd.n5175 gnd.n5174 12.1094
R9226 gnd.n3593 gnd.n3592 12.0247
R9227 gnd.n3561 gnd.n3560 12.0247
R9228 gnd.n3529 gnd.n3528 12.0247
R9229 gnd.n3498 gnd.n3497 12.0247
R9230 gnd.n3466 gnd.n3465 12.0247
R9231 gnd.n3434 gnd.n3433 12.0247
R9232 gnd.n3402 gnd.n3401 12.0247
R9233 gnd.n3371 gnd.n3370 12.0247
R9234 gnd.n2244 gnd.t79 11.7908
R9235 gnd.t240 gnd.n1134 11.7908
R9236 gnd.t47 gnd.t55 11.7908
R9237 gnd.t202 gnd.t37 11.7908
R9238 gnd.n5471 gnd.t219 11.7908
R9239 gnd.n6859 gnd.t114 11.7908
R9240 gnd.t205 gnd.n4795 11.4721
R9241 gnd.t32 gnd.n1976 11.4721
R9242 gnd.n5086 gnd.t36 11.4721
R9243 gnd.n5350 gnd.t248 11.4721
R9244 gnd.n3596 gnd.n3583 11.249
R9245 gnd.n3564 gnd.n3551 11.249
R9246 gnd.n3532 gnd.n3519 11.249
R9247 gnd.n3501 gnd.n3488 11.249
R9248 gnd.n3469 gnd.n3456 11.249
R9249 gnd.n3437 gnd.n3424 11.249
R9250 gnd.n3405 gnd.n3392 11.249
R9251 gnd.n3374 gnd.n3361 11.249
R9252 gnd.n3035 gnd.t45 11.1535
R9253 gnd.n2208 gnd.t127 11.1535
R9254 gnd.n2083 gnd.t61 11.1535
R9255 gnd.n4853 gnd.t194 11.1535
R9256 gnd.t15 gnd.n1853 11.1535
R9257 gnd.n5383 gnd.t39 11.1535
R9258 gnd.n6883 gnd.t103 11.1535
R9259 gnd.n4828 gnd.n2012 10.8348
R9260 gnd.n4828 gnd.n4827 10.8348
R9261 gnd.n4999 gnd.n4998 10.8348
R9262 gnd.n4998 gnd.n1913 10.8348
R9263 gnd.n5154 gnd.n5153 10.8348
R9264 gnd.n5153 gnd.n1832 10.8348
R9265 gnd.n5543 gnd.n5540 10.6672
R9266 gnd.n486 gnd.n284 10.6672
R9267 gnd.n3958 gnd.n3956 10.6672
R9268 gnd.n4519 gnd.n4518 10.6672
R9269 gnd.n5280 gnd.n1760 10.6151
R9270 gnd.n5280 gnd.n5279 10.6151
R9271 gnd.n5277 gnd.n1764 10.6151
R9272 gnd.n5272 gnd.n1764 10.6151
R9273 gnd.n5272 gnd.n5271 10.6151
R9274 gnd.n5271 gnd.n5270 10.6151
R9275 gnd.n5270 gnd.n1767 10.6151
R9276 gnd.n5265 gnd.n1767 10.6151
R9277 gnd.n5265 gnd.n5264 10.6151
R9278 gnd.n5264 gnd.n5263 10.6151
R9279 gnd.n5263 gnd.n1770 10.6151
R9280 gnd.n5258 gnd.n1770 10.6151
R9281 gnd.n5258 gnd.n5257 10.6151
R9282 gnd.n5257 gnd.n5256 10.6151
R9283 gnd.n5256 gnd.n1773 10.6151
R9284 gnd.n5251 gnd.n1773 10.6151
R9285 gnd.n5251 gnd.n5250 10.6151
R9286 gnd.n5250 gnd.n5249 10.6151
R9287 gnd.n5249 gnd.n1776 10.6151
R9288 gnd.n5244 gnd.n1776 10.6151
R9289 gnd.n5244 gnd.n5243 10.6151
R9290 gnd.n5243 gnd.n5242 10.6151
R9291 gnd.n5242 gnd.n1779 10.6151
R9292 gnd.n5237 gnd.n1779 10.6151
R9293 gnd.n5237 gnd.n5236 10.6151
R9294 gnd.n5236 gnd.n5235 10.6151
R9295 gnd.n5235 gnd.n1782 10.6151
R9296 gnd.n5230 gnd.n1782 10.6151
R9297 gnd.n5230 gnd.n5229 10.6151
R9298 gnd.n5229 gnd.n5228 10.6151
R9299 gnd.n4742 gnd.n4741 10.6151
R9300 gnd.n4744 gnd.n4742 10.6151
R9301 gnd.n4745 gnd.n4744 10.6151
R9302 gnd.n4746 gnd.n4745 10.6151
R9303 gnd.n4746 gnd.n2047 10.6151
R9304 gnd.n4756 gnd.n2047 10.6151
R9305 gnd.n4757 gnd.n4756 10.6151
R9306 gnd.n4782 gnd.n4757 10.6151
R9307 gnd.n4782 gnd.n4781 10.6151
R9308 gnd.n4781 gnd.n4780 10.6151
R9309 gnd.n4780 gnd.n4779 10.6151
R9310 gnd.n4779 gnd.n4758 10.6151
R9311 gnd.n4774 gnd.n4758 10.6151
R9312 gnd.n4774 gnd.n4773 10.6151
R9313 gnd.n4773 gnd.n4772 10.6151
R9314 gnd.n4772 gnd.n4771 10.6151
R9315 gnd.n4771 gnd.n4769 10.6151
R9316 gnd.n4769 gnd.n4768 10.6151
R9317 gnd.n4768 gnd.n4762 10.6151
R9318 gnd.n4762 gnd.n1997 10.6151
R9319 gnd.n4858 gnd.n1997 10.6151
R9320 gnd.n4858 gnd.n4857 10.6151
R9321 gnd.n4857 gnd.n4856 10.6151
R9322 gnd.n4856 gnd.n4855 10.6151
R9323 gnd.n4855 gnd.n1999 10.6151
R9324 gnd.n1999 gnd.n1998 10.6151
R9325 gnd.n1998 gnd.n1974 10.6151
R9326 gnd.n4885 gnd.n1974 10.6151
R9327 gnd.n4886 gnd.n4885 10.6151
R9328 gnd.n4887 gnd.n4886 10.6151
R9329 gnd.n4893 gnd.n4887 10.6151
R9330 gnd.n4894 gnd.n4893 10.6151
R9331 gnd.n4895 gnd.n4894 10.6151
R9332 gnd.n4895 gnd.n1946 10.6151
R9333 gnd.n4929 gnd.n1946 10.6151
R9334 gnd.n4930 gnd.n4929 10.6151
R9335 gnd.n4931 gnd.n4930 10.6151
R9336 gnd.n4943 gnd.n4931 10.6151
R9337 gnd.n4943 gnd.n4942 10.6151
R9338 gnd.n4942 gnd.n4941 10.6151
R9339 gnd.n4941 gnd.n4938 10.6151
R9340 gnd.n4938 gnd.n4937 10.6151
R9341 gnd.n4937 gnd.n4935 10.6151
R9342 gnd.n4935 gnd.n4934 10.6151
R9343 gnd.n4934 gnd.n4932 10.6151
R9344 gnd.n4932 gnd.n1896 10.6151
R9345 gnd.n5025 gnd.n1896 10.6151
R9346 gnd.n5026 gnd.n5025 10.6151
R9347 gnd.n5033 gnd.n5026 10.6151
R9348 gnd.n5033 gnd.n5032 10.6151
R9349 gnd.n5032 gnd.n5031 10.6151
R9350 gnd.n5031 gnd.n5030 10.6151
R9351 gnd.n5030 gnd.n5028 10.6151
R9352 gnd.n5028 gnd.n5027 10.6151
R9353 gnd.n5027 gnd.n1871 10.6151
R9354 gnd.n5060 gnd.n1871 10.6151
R9355 gnd.n5061 gnd.n5060 10.6151
R9356 gnd.n5064 gnd.n5061 10.6151
R9357 gnd.n5065 gnd.n5064 10.6151
R9358 gnd.n5075 gnd.n5065 10.6151
R9359 gnd.n5075 gnd.n5074 10.6151
R9360 gnd.n5074 gnd.n5073 10.6151
R9361 gnd.n5073 gnd.n5072 10.6151
R9362 gnd.n5072 gnd.n5070 10.6151
R9363 gnd.n5070 gnd.n5069 10.6151
R9364 gnd.n5069 gnd.n5067 10.6151
R9365 gnd.n5067 gnd.n5066 10.6151
R9366 gnd.n5066 gnd.n1824 10.6151
R9367 gnd.n5163 gnd.n1824 10.6151
R9368 gnd.n5164 gnd.n5163 10.6151
R9369 gnd.n5165 gnd.n5164 10.6151
R9370 gnd.n5165 gnd.n1808 10.6151
R9371 gnd.n5186 gnd.n1808 10.6151
R9372 gnd.n5187 gnd.n5186 10.6151
R9373 gnd.n5194 gnd.n5187 10.6151
R9374 gnd.n5194 gnd.n5193 10.6151
R9375 gnd.n5193 gnd.n5192 10.6151
R9376 gnd.n5192 gnd.n5189 10.6151
R9377 gnd.n5189 gnd.n5188 10.6151
R9378 gnd.n5188 gnd.n1785 10.6151
R9379 gnd.n5222 gnd.n1785 10.6151
R9380 gnd.n5223 gnd.n5222 10.6151
R9381 gnd.n5224 gnd.n5223 10.6151
R9382 gnd.n4676 gnd.n1214 10.6151
R9383 gnd.n4679 gnd.n4676 10.6151
R9384 gnd.n4684 gnd.n4681 10.6151
R9385 gnd.n4685 gnd.n4684 10.6151
R9386 gnd.n4688 gnd.n4685 10.6151
R9387 gnd.n4689 gnd.n4688 10.6151
R9388 gnd.n4692 gnd.n4689 10.6151
R9389 gnd.n4693 gnd.n4692 10.6151
R9390 gnd.n4696 gnd.n4693 10.6151
R9391 gnd.n4697 gnd.n4696 10.6151
R9392 gnd.n4700 gnd.n4697 10.6151
R9393 gnd.n4701 gnd.n4700 10.6151
R9394 gnd.n4704 gnd.n4701 10.6151
R9395 gnd.n4705 gnd.n4704 10.6151
R9396 gnd.n4708 gnd.n4705 10.6151
R9397 gnd.n4709 gnd.n4708 10.6151
R9398 gnd.n4712 gnd.n4709 10.6151
R9399 gnd.n4713 gnd.n4712 10.6151
R9400 gnd.n4716 gnd.n4713 10.6151
R9401 gnd.n4717 gnd.n4716 10.6151
R9402 gnd.n4720 gnd.n4717 10.6151
R9403 gnd.n4721 gnd.n4720 10.6151
R9404 gnd.n4724 gnd.n4721 10.6151
R9405 gnd.n4725 gnd.n4724 10.6151
R9406 gnd.n4728 gnd.n4725 10.6151
R9407 gnd.n4729 gnd.n4728 10.6151
R9408 gnd.n4732 gnd.n4729 10.6151
R9409 gnd.n4733 gnd.n4732 10.6151
R9410 gnd.n4736 gnd.n4733 10.6151
R9411 gnd.n4737 gnd.n4736 10.6151
R9412 gnd.n5899 gnd.n5898 10.6151
R9413 gnd.n5898 gnd.n5897 10.6151
R9414 gnd.n5897 gnd.n5896 10.6151
R9415 gnd.n5896 gnd.n5894 10.6151
R9416 gnd.n5894 gnd.n5891 10.6151
R9417 gnd.n5891 gnd.n5890 10.6151
R9418 gnd.n5890 gnd.n5887 10.6151
R9419 gnd.n5887 gnd.n5886 10.6151
R9420 gnd.n5886 gnd.n5883 10.6151
R9421 gnd.n5883 gnd.n5882 10.6151
R9422 gnd.n5882 gnd.n5879 10.6151
R9423 gnd.n5879 gnd.n5878 10.6151
R9424 gnd.n5878 gnd.n5875 10.6151
R9425 gnd.n5875 gnd.n5874 10.6151
R9426 gnd.n5874 gnd.n5871 10.6151
R9427 gnd.n5871 gnd.n5870 10.6151
R9428 gnd.n5870 gnd.n5867 10.6151
R9429 gnd.n5867 gnd.n5866 10.6151
R9430 gnd.n5866 gnd.n5863 10.6151
R9431 gnd.n5863 gnd.n5862 10.6151
R9432 gnd.n5862 gnd.n5859 10.6151
R9433 gnd.n5859 gnd.n5858 10.6151
R9434 gnd.n5858 gnd.n5855 10.6151
R9435 gnd.n5855 gnd.n5854 10.6151
R9436 gnd.n5854 gnd.n5851 10.6151
R9437 gnd.n5851 gnd.n5850 10.6151
R9438 gnd.n5850 gnd.n5847 10.6151
R9439 gnd.n5847 gnd.n5846 10.6151
R9440 gnd.n5843 gnd.n5842 10.6151
R9441 gnd.n5842 gnd.n1215 10.6151
R9442 gnd.n5345 gnd.n1735 10.6151
R9443 gnd.n1736 gnd.n1735 10.6151
R9444 gnd.n5338 gnd.n1736 10.6151
R9445 gnd.n5338 gnd.n5337 10.6151
R9446 gnd.n5337 gnd.n5336 10.6151
R9447 gnd.n5336 gnd.n1738 10.6151
R9448 gnd.n5331 gnd.n1738 10.6151
R9449 gnd.n5331 gnd.n5330 10.6151
R9450 gnd.n5330 gnd.n5329 10.6151
R9451 gnd.n5329 gnd.n1741 10.6151
R9452 gnd.n5324 gnd.n1741 10.6151
R9453 gnd.n5324 gnd.n5323 10.6151
R9454 gnd.n5323 gnd.n5322 10.6151
R9455 gnd.n5322 gnd.n1744 10.6151
R9456 gnd.n5317 gnd.n1744 10.6151
R9457 gnd.n5317 gnd.n5316 10.6151
R9458 gnd.n5316 gnd.n5315 10.6151
R9459 gnd.n5315 gnd.n1747 10.6151
R9460 gnd.n5310 gnd.n1747 10.6151
R9461 gnd.n5310 gnd.n5309 10.6151
R9462 gnd.n5309 gnd.n5308 10.6151
R9463 gnd.n5308 gnd.n1750 10.6151
R9464 gnd.n5303 gnd.n1750 10.6151
R9465 gnd.n5303 gnd.n5302 10.6151
R9466 gnd.n5302 gnd.n5301 10.6151
R9467 gnd.n5301 gnd.n1753 10.6151
R9468 gnd.n5296 gnd.n1753 10.6151
R9469 gnd.n5296 gnd.n5295 10.6151
R9470 gnd.n5293 gnd.n1758 10.6151
R9471 gnd.n5288 gnd.n1758 10.6151
R9472 gnd.n5835 gnd.n5834 10.6151
R9473 gnd.n5834 gnd.n1274 10.6151
R9474 gnd.n2053 gnd.n1274 10.6151
R9475 gnd.n4750 gnd.n2053 10.6151
R9476 gnd.n4751 gnd.n4750 10.6151
R9477 gnd.n4752 gnd.n4751 10.6151
R9478 gnd.n4752 gnd.n2042 10.6151
R9479 gnd.n4786 gnd.n2042 10.6151
R9480 gnd.n4787 gnd.n4786 10.6151
R9481 gnd.n4793 gnd.n4787 10.6151
R9482 gnd.n4793 gnd.n4792 10.6151
R9483 gnd.n4792 gnd.n4791 10.6151
R9484 gnd.n4791 gnd.n4788 10.6151
R9485 gnd.n4788 gnd.n2017 10.6151
R9486 gnd.n4820 gnd.n2017 10.6151
R9487 gnd.n4821 gnd.n4820 10.6151
R9488 gnd.n4825 gnd.n4821 10.6151
R9489 gnd.n4825 gnd.n4824 10.6151
R9490 gnd.n4824 gnd.n4823 10.6151
R9491 gnd.n4823 gnd.n1992 10.6151
R9492 gnd.n4862 gnd.n1992 10.6151
R9493 gnd.n4863 gnd.n4862 10.6151
R9494 gnd.n4864 gnd.n4863 10.6151
R9495 gnd.n4864 gnd.n1978 10.6151
R9496 gnd.n4878 gnd.n1978 10.6151
R9497 gnd.n4879 gnd.n4878 10.6151
R9498 gnd.n4880 gnd.n4879 10.6151
R9499 gnd.n4880 gnd.n1967 10.6151
R9500 gnd.n4904 gnd.n1967 10.6151
R9501 gnd.n4904 gnd.n4903 10.6151
R9502 gnd.n4903 gnd.n4902 10.6151
R9503 gnd.n4902 gnd.n1968 10.6151
R9504 gnd.n1971 gnd.n1968 10.6151
R9505 gnd.n1971 gnd.n1970 10.6151
R9506 gnd.n1970 gnd.n1940 10.6151
R9507 gnd.n4949 gnd.n1940 10.6151
R9508 gnd.n4949 gnd.n4948 10.6151
R9509 gnd.n4948 gnd.n4947 10.6151
R9510 gnd.n4947 gnd.n1941 10.6151
R9511 gnd.n1941 gnd.n1918 10.6151
R9512 gnd.n5001 gnd.n1918 10.6151
R9513 gnd.n5002 gnd.n5001 10.6151
R9514 gnd.n5003 gnd.n5002 10.6151
R9515 gnd.n5003 gnd.n1903 10.6151
R9516 gnd.n5019 gnd.n1903 10.6151
R9517 gnd.n5020 gnd.n5019 10.6151
R9518 gnd.n5021 gnd.n5020 10.6151
R9519 gnd.n5021 gnd.n1891 10.6151
R9520 gnd.n5037 gnd.n1891 10.6151
R9521 gnd.n5038 gnd.n5037 10.6151
R9522 gnd.n5039 gnd.n5038 10.6151
R9523 gnd.n5039 gnd.n1875 10.6151
R9524 gnd.n5053 gnd.n1875 10.6151
R9525 gnd.n5054 gnd.n5053 10.6151
R9526 gnd.n5055 gnd.n5054 10.6151
R9527 gnd.n5055 gnd.n1867 10.6151
R9528 gnd.n5083 gnd.n1867 10.6151
R9529 gnd.n5083 gnd.n5082 10.6151
R9530 gnd.n5082 gnd.n5081 10.6151
R9531 gnd.n5081 gnd.n1868 10.6151
R9532 gnd.n1868 gnd.n1843 10.6151
R9533 gnd.n5140 gnd.n1843 10.6151
R9534 gnd.n5141 gnd.n5140 10.6151
R9535 gnd.n5142 gnd.n5141 10.6151
R9536 gnd.n5142 gnd.n1828 10.6151
R9537 gnd.n5156 gnd.n1828 10.6151
R9538 gnd.n5157 gnd.n5156 10.6151
R9539 gnd.n5158 gnd.n5157 10.6151
R9540 gnd.n5158 gnd.n1823 10.6151
R9541 gnd.n5172 gnd.n1823 10.6151
R9542 gnd.n5172 gnd.n5171 10.6151
R9543 gnd.n5171 gnd.n5170 10.6151
R9544 gnd.n5170 gnd.n1804 10.6151
R9545 gnd.n5199 gnd.n1804 10.6151
R9546 gnd.n5200 gnd.n5199 10.6151
R9547 gnd.n5201 gnd.n5200 10.6151
R9548 gnd.n5201 gnd.n1789 10.6151
R9549 gnd.n5215 gnd.n1789 10.6151
R9550 gnd.n5216 gnd.n5215 10.6151
R9551 gnd.n5217 gnd.n5216 10.6151
R9552 gnd.n5217 gnd.n1715 10.6151
R9553 gnd.n5348 gnd.n1715 10.6151
R9554 gnd.n5348 gnd.n5347 10.6151
R9555 gnd.n2954 gnd.t29 10.5161
R9556 gnd.n2399 gnd.t41 10.5161
R9557 gnd.n3320 gnd.t3 10.5161
R9558 gnd.t140 gnd.n2169 10.5161
R9559 gnd.n2172 gnd.t129 10.5161
R9560 gnd.n4876 gnd.t194 10.5161
R9561 gnd.n5062 gnd.t15 10.5161
R9562 gnd.n6790 gnd.t95 10.5161
R9563 gnd.n6799 gnd.t120 10.5161
R9564 gnd.n3597 gnd.n3581 10.4732
R9565 gnd.n3565 gnd.n3549 10.4732
R9566 gnd.n3533 gnd.n3517 10.4732
R9567 gnd.n3502 gnd.n3486 10.4732
R9568 gnd.n3470 gnd.n3454 10.4732
R9569 gnd.n3438 gnd.n3422 10.4732
R9570 gnd.n3406 gnd.n3390 10.4732
R9571 gnd.n3375 gnd.n3359 10.4732
R9572 gnd.t59 gnd.n2416 9.87883
R9573 gnd.t105 gnd.n2205 9.87883
R9574 gnd.n6013 gnd.n1050 9.87883
R9575 gnd.n4217 gnd.t108 9.87883
R9576 gnd.t51 gnd.t322 9.87883
R9577 gnd.n1615 gnd.t81 9.87883
R9578 gnd.n6720 gnd.n509 9.87883
R9579 gnd.n6877 gnd.t136 9.87883
R9580 gnd.n3601 gnd.n3600 9.69747
R9581 gnd.n3569 gnd.n3568 9.69747
R9582 gnd.n3537 gnd.n3536 9.69747
R9583 gnd.n3506 gnd.n3505 9.69747
R9584 gnd.n3474 gnd.n3473 9.69747
R9585 gnd.n3442 gnd.n3441 9.69747
R9586 gnd.n3410 gnd.n3409 9.69747
R9587 gnd.n3379 gnd.n3378 9.69747
R9588 gnd.n4760 gnd.n4759 9.56018
R9589 gnd.n4836 gnd.n2005 9.56018
R9590 gnd.n4889 gnd.t33 9.56018
R9591 gnd.n4963 gnd.n1928 9.56018
R9592 gnd.n4969 gnd.n1916 9.56018
R9593 gnd.n5050 gnd.t12 9.56018
R9594 gnd.n5145 gnd.n5144 9.56018
R9595 gnd.n5175 gnd.n1816 9.56018
R9596 gnd.n3607 gnd.n3606 9.45567
R9597 gnd.n3575 gnd.n3574 9.45567
R9598 gnd.n3543 gnd.n3542 9.45567
R9599 gnd.n3512 gnd.n3511 9.45567
R9600 gnd.n3480 gnd.n3479 9.45567
R9601 gnd.n3448 gnd.n3447 9.45567
R9602 gnd.n3416 gnd.n3415 9.45567
R9603 gnd.n3385 gnd.n3384 9.45567
R9604 gnd.n5580 gnd.n5579 9.30959
R9605 gnd.n442 gnd.n306 9.30959
R9606 gnd.n3995 gnd.n3994 9.30959
R9607 gnd.n4473 gnd.n4470 9.30959
R9608 gnd.n3606 gnd.n3605 9.3005
R9609 gnd.n3579 gnd.n3578 9.3005
R9610 gnd.n3600 gnd.n3599 9.3005
R9611 gnd.n3598 gnd.n3597 9.3005
R9612 gnd.n3583 gnd.n3582 9.3005
R9613 gnd.n3592 gnd.n3591 9.3005
R9614 gnd.n3590 gnd.n3589 9.3005
R9615 gnd.n3574 gnd.n3573 9.3005
R9616 gnd.n3547 gnd.n3546 9.3005
R9617 gnd.n3568 gnd.n3567 9.3005
R9618 gnd.n3566 gnd.n3565 9.3005
R9619 gnd.n3551 gnd.n3550 9.3005
R9620 gnd.n3560 gnd.n3559 9.3005
R9621 gnd.n3558 gnd.n3557 9.3005
R9622 gnd.n3542 gnd.n3541 9.3005
R9623 gnd.n3515 gnd.n3514 9.3005
R9624 gnd.n3536 gnd.n3535 9.3005
R9625 gnd.n3534 gnd.n3533 9.3005
R9626 gnd.n3519 gnd.n3518 9.3005
R9627 gnd.n3528 gnd.n3527 9.3005
R9628 gnd.n3526 gnd.n3525 9.3005
R9629 gnd.n3511 gnd.n3510 9.3005
R9630 gnd.n3484 gnd.n3483 9.3005
R9631 gnd.n3505 gnd.n3504 9.3005
R9632 gnd.n3503 gnd.n3502 9.3005
R9633 gnd.n3488 gnd.n3487 9.3005
R9634 gnd.n3497 gnd.n3496 9.3005
R9635 gnd.n3495 gnd.n3494 9.3005
R9636 gnd.n3479 gnd.n3478 9.3005
R9637 gnd.n3452 gnd.n3451 9.3005
R9638 gnd.n3473 gnd.n3472 9.3005
R9639 gnd.n3471 gnd.n3470 9.3005
R9640 gnd.n3456 gnd.n3455 9.3005
R9641 gnd.n3465 gnd.n3464 9.3005
R9642 gnd.n3463 gnd.n3462 9.3005
R9643 gnd.n3447 gnd.n3446 9.3005
R9644 gnd.n3420 gnd.n3419 9.3005
R9645 gnd.n3441 gnd.n3440 9.3005
R9646 gnd.n3439 gnd.n3438 9.3005
R9647 gnd.n3424 gnd.n3423 9.3005
R9648 gnd.n3433 gnd.n3432 9.3005
R9649 gnd.n3431 gnd.n3430 9.3005
R9650 gnd.n3415 gnd.n3414 9.3005
R9651 gnd.n3388 gnd.n3387 9.3005
R9652 gnd.n3409 gnd.n3408 9.3005
R9653 gnd.n3407 gnd.n3406 9.3005
R9654 gnd.n3392 gnd.n3391 9.3005
R9655 gnd.n3401 gnd.n3400 9.3005
R9656 gnd.n3399 gnd.n3398 9.3005
R9657 gnd.n3384 gnd.n3383 9.3005
R9658 gnd.n3357 gnd.n3356 9.3005
R9659 gnd.n3378 gnd.n3377 9.3005
R9660 gnd.n3376 gnd.n3375 9.3005
R9661 gnd.n3361 gnd.n3360 9.3005
R9662 gnd.n3370 gnd.n3369 9.3005
R9663 gnd.n3368 gnd.n3367 9.3005
R9664 gnd.n3732 gnd.n3731 9.3005
R9665 gnd.n3730 gnd.n2299 9.3005
R9666 gnd.n3729 gnd.n3728 9.3005
R9667 gnd.n3725 gnd.n2300 9.3005
R9668 gnd.n3722 gnd.n2301 9.3005
R9669 gnd.n3721 gnd.n2302 9.3005
R9670 gnd.n3718 gnd.n2303 9.3005
R9671 gnd.n3717 gnd.n2304 9.3005
R9672 gnd.n3714 gnd.n2305 9.3005
R9673 gnd.n3713 gnd.n2306 9.3005
R9674 gnd.n3710 gnd.n2307 9.3005
R9675 gnd.n3709 gnd.n2308 9.3005
R9676 gnd.n3706 gnd.n2309 9.3005
R9677 gnd.n3705 gnd.n2310 9.3005
R9678 gnd.n3702 gnd.n3701 9.3005
R9679 gnd.n3700 gnd.n2311 9.3005
R9680 gnd.n3733 gnd.n2298 9.3005
R9681 gnd.n2973 gnd.n2972 9.3005
R9682 gnd.n2677 gnd.n2676 9.3005
R9683 gnd.n3000 gnd.n2999 9.3005
R9684 gnd.n3001 gnd.n2675 9.3005
R9685 gnd.n3005 gnd.n3002 9.3005
R9686 gnd.n3004 gnd.n3003 9.3005
R9687 gnd.n2649 gnd.n2648 9.3005
R9688 gnd.n3030 gnd.n3029 9.3005
R9689 gnd.n3031 gnd.n2647 9.3005
R9690 gnd.n3033 gnd.n3032 9.3005
R9691 gnd.n2627 gnd.n2626 9.3005
R9692 gnd.n3061 gnd.n3060 9.3005
R9693 gnd.n3062 gnd.n2625 9.3005
R9694 gnd.n3070 gnd.n3063 9.3005
R9695 gnd.n3069 gnd.n3064 9.3005
R9696 gnd.n3068 gnd.n3066 9.3005
R9697 gnd.n3065 gnd.n2574 9.3005
R9698 gnd.n3118 gnd.n2575 9.3005
R9699 gnd.n3117 gnd.n2576 9.3005
R9700 gnd.n3116 gnd.n2577 9.3005
R9701 gnd.n2596 gnd.n2578 9.3005
R9702 gnd.n2598 gnd.n2597 9.3005
R9703 gnd.n2496 gnd.n2495 9.3005
R9704 gnd.n3156 gnd.n3155 9.3005
R9705 gnd.n3157 gnd.n2494 9.3005
R9706 gnd.n3161 gnd.n3158 9.3005
R9707 gnd.n3160 gnd.n3159 9.3005
R9708 gnd.n2469 gnd.n2468 9.3005
R9709 gnd.n3196 gnd.n3195 9.3005
R9710 gnd.n3197 gnd.n2467 9.3005
R9711 gnd.n3201 gnd.n3198 9.3005
R9712 gnd.n3200 gnd.n3199 9.3005
R9713 gnd.n2442 gnd.n2441 9.3005
R9714 gnd.n3241 gnd.n3240 9.3005
R9715 gnd.n3242 gnd.n2440 9.3005
R9716 gnd.n3246 gnd.n3243 9.3005
R9717 gnd.n3245 gnd.n3244 9.3005
R9718 gnd.n2414 gnd.n2413 9.3005
R9719 gnd.n3281 gnd.n3280 9.3005
R9720 gnd.n3282 gnd.n2412 9.3005
R9721 gnd.n3286 gnd.n3283 9.3005
R9722 gnd.n3285 gnd.n3284 9.3005
R9723 gnd.n2387 gnd.n2386 9.3005
R9724 gnd.n3330 gnd.n3329 9.3005
R9725 gnd.n3331 gnd.n2385 9.3005
R9726 gnd.n3335 gnd.n3332 9.3005
R9727 gnd.n3334 gnd.n3333 9.3005
R9728 gnd.n2360 gnd.n2359 9.3005
R9729 gnd.n3625 gnd.n3624 9.3005
R9730 gnd.n3626 gnd.n2358 9.3005
R9731 gnd.n3632 gnd.n3627 9.3005
R9732 gnd.n3631 gnd.n3628 9.3005
R9733 gnd.n3630 gnd.n3629 9.3005
R9734 gnd.n2974 gnd.n2971 9.3005
R9735 gnd.n2756 gnd.n2715 9.3005
R9736 gnd.n2751 gnd.n2750 9.3005
R9737 gnd.n2749 gnd.n2716 9.3005
R9738 gnd.n2748 gnd.n2747 9.3005
R9739 gnd.n2744 gnd.n2717 9.3005
R9740 gnd.n2741 gnd.n2740 9.3005
R9741 gnd.n2739 gnd.n2718 9.3005
R9742 gnd.n2738 gnd.n2737 9.3005
R9743 gnd.n2734 gnd.n2719 9.3005
R9744 gnd.n2731 gnd.n2730 9.3005
R9745 gnd.n2729 gnd.n2720 9.3005
R9746 gnd.n2728 gnd.n2727 9.3005
R9747 gnd.n2724 gnd.n2722 9.3005
R9748 gnd.n2721 gnd.n2701 9.3005
R9749 gnd.n2968 gnd.n2700 9.3005
R9750 gnd.n2970 gnd.n2969 9.3005
R9751 gnd.n2758 gnd.n2757 9.3005
R9752 gnd.n2981 gnd.n2687 9.3005
R9753 gnd.n2988 gnd.n2688 9.3005
R9754 gnd.n2990 gnd.n2989 9.3005
R9755 gnd.n2991 gnd.n2668 9.3005
R9756 gnd.n3010 gnd.n3009 9.3005
R9757 gnd.n3012 gnd.n2660 9.3005
R9758 gnd.n3019 gnd.n2662 9.3005
R9759 gnd.n3020 gnd.n2657 9.3005
R9760 gnd.n3022 gnd.n3021 9.3005
R9761 gnd.n2658 gnd.n2643 9.3005
R9762 gnd.n3038 gnd.n2641 9.3005
R9763 gnd.n3042 gnd.n3041 9.3005
R9764 gnd.n3040 gnd.n2617 9.3005
R9765 gnd.n3077 gnd.n2616 9.3005
R9766 gnd.n3080 gnd.n3079 9.3005
R9767 gnd.n2613 gnd.n2612 9.3005
R9768 gnd.n3086 gnd.n2614 9.3005
R9769 gnd.n3088 gnd.n3087 9.3005
R9770 gnd.n3090 gnd.n2611 9.3005
R9771 gnd.n3093 gnd.n3092 9.3005
R9772 gnd.n3096 gnd.n3094 9.3005
R9773 gnd.n3098 gnd.n3097 9.3005
R9774 gnd.n3104 gnd.n3099 9.3005
R9775 gnd.n3103 gnd.n3102 9.3005
R9776 gnd.n2487 gnd.n2486 9.3005
R9777 gnd.n3170 gnd.n3169 9.3005
R9778 gnd.n3171 gnd.n2480 9.3005
R9779 gnd.n3179 gnd.n2479 9.3005
R9780 gnd.n3182 gnd.n3181 9.3005
R9781 gnd.n3184 gnd.n3183 9.3005
R9782 gnd.n3187 gnd.n2462 9.3005
R9783 gnd.n3185 gnd.n2460 9.3005
R9784 gnd.n3207 gnd.n2458 9.3005
R9785 gnd.n3209 gnd.n3208 9.3005
R9786 gnd.n2432 gnd.n2431 9.3005
R9787 gnd.n3255 gnd.n3254 9.3005
R9788 gnd.n3256 gnd.n2425 9.3005
R9789 gnd.n3264 gnd.n2424 9.3005
R9790 gnd.n3267 gnd.n3266 9.3005
R9791 gnd.n3269 gnd.n3268 9.3005
R9792 gnd.n3272 gnd.n2407 9.3005
R9793 gnd.n3270 gnd.n2405 9.3005
R9794 gnd.n3292 gnd.n2403 9.3005
R9795 gnd.n3294 gnd.n3293 9.3005
R9796 gnd.n2378 gnd.n2377 9.3005
R9797 gnd.n3344 gnd.n3343 9.3005
R9798 gnd.n3345 gnd.n2371 9.3005
R9799 gnd.n3354 gnd.n2370 9.3005
R9800 gnd.n3613 gnd.n3612 9.3005
R9801 gnd.n3615 gnd.n3614 9.3005
R9802 gnd.n3616 gnd.n2351 9.3005
R9803 gnd.n3640 gnd.n3639 9.3005
R9804 gnd.n2352 gnd.n2314 9.3005
R9805 gnd.n2979 gnd.n2978 9.3005
R9806 gnd.n3696 gnd.n2315 9.3005
R9807 gnd.n3695 gnd.n2317 9.3005
R9808 gnd.n3692 gnd.n2318 9.3005
R9809 gnd.n3691 gnd.n2319 9.3005
R9810 gnd.n3688 gnd.n2320 9.3005
R9811 gnd.n3687 gnd.n2321 9.3005
R9812 gnd.n3684 gnd.n2322 9.3005
R9813 gnd.n3683 gnd.n2323 9.3005
R9814 gnd.n3680 gnd.n2324 9.3005
R9815 gnd.n3679 gnd.n2325 9.3005
R9816 gnd.n3676 gnd.n2326 9.3005
R9817 gnd.n3675 gnd.n2327 9.3005
R9818 gnd.n3672 gnd.n2328 9.3005
R9819 gnd.n3671 gnd.n2329 9.3005
R9820 gnd.n3668 gnd.n2330 9.3005
R9821 gnd.n3667 gnd.n2331 9.3005
R9822 gnd.n3664 gnd.n2332 9.3005
R9823 gnd.n3663 gnd.n2333 9.3005
R9824 gnd.n3660 gnd.n2334 9.3005
R9825 gnd.n3659 gnd.n2335 9.3005
R9826 gnd.n3656 gnd.n2336 9.3005
R9827 gnd.n3655 gnd.n2337 9.3005
R9828 gnd.n3652 gnd.n2341 9.3005
R9829 gnd.n3651 gnd.n2342 9.3005
R9830 gnd.n3648 gnd.n2343 9.3005
R9831 gnd.n3647 gnd.n2344 9.3005
R9832 gnd.n3698 gnd.n3697 9.3005
R9833 gnd.n3148 gnd.n3132 9.3005
R9834 gnd.n3147 gnd.n3133 9.3005
R9835 gnd.n3146 gnd.n3134 9.3005
R9836 gnd.n3144 gnd.n3135 9.3005
R9837 gnd.n3143 gnd.n3136 9.3005
R9838 gnd.n3141 gnd.n3137 9.3005
R9839 gnd.n3140 gnd.n3138 9.3005
R9840 gnd.n2450 gnd.n2449 9.3005
R9841 gnd.n3217 gnd.n3216 9.3005
R9842 gnd.n3218 gnd.n2448 9.3005
R9843 gnd.n3235 gnd.n3219 9.3005
R9844 gnd.n3234 gnd.n3220 9.3005
R9845 gnd.n3233 gnd.n3221 9.3005
R9846 gnd.n3231 gnd.n3222 9.3005
R9847 gnd.n3230 gnd.n3223 9.3005
R9848 gnd.n3228 gnd.n3224 9.3005
R9849 gnd.n3227 gnd.n3225 9.3005
R9850 gnd.n2394 gnd.n2393 9.3005
R9851 gnd.n3302 gnd.n3301 9.3005
R9852 gnd.n3303 gnd.n2392 9.3005
R9853 gnd.n3324 gnd.n3304 9.3005
R9854 gnd.n3323 gnd.n3305 9.3005
R9855 gnd.n3322 gnd.n3306 9.3005
R9856 gnd.n3319 gnd.n3307 9.3005
R9857 gnd.n3318 gnd.n3308 9.3005
R9858 gnd.n3316 gnd.n3309 9.3005
R9859 gnd.n3315 gnd.n3310 9.3005
R9860 gnd.n3313 gnd.n3312 9.3005
R9861 gnd.n3311 gnd.n2346 9.3005
R9862 gnd.n2889 gnd.n2888 9.3005
R9863 gnd.n2779 gnd.n2778 9.3005
R9864 gnd.n2903 gnd.n2902 9.3005
R9865 gnd.n2904 gnd.n2777 9.3005
R9866 gnd.n2906 gnd.n2905 9.3005
R9867 gnd.n2767 gnd.n2766 9.3005
R9868 gnd.n2919 gnd.n2918 9.3005
R9869 gnd.n2920 gnd.n2765 9.3005
R9870 gnd.n2952 gnd.n2921 9.3005
R9871 gnd.n2951 gnd.n2922 9.3005
R9872 gnd.n2950 gnd.n2923 9.3005
R9873 gnd.n2949 gnd.n2924 9.3005
R9874 gnd.n2946 gnd.n2925 9.3005
R9875 gnd.n2945 gnd.n2926 9.3005
R9876 gnd.n2944 gnd.n2927 9.3005
R9877 gnd.n2942 gnd.n2928 9.3005
R9878 gnd.n2941 gnd.n2929 9.3005
R9879 gnd.n2938 gnd.n2930 9.3005
R9880 gnd.n2937 gnd.n2931 9.3005
R9881 gnd.n2936 gnd.n2932 9.3005
R9882 gnd.n2934 gnd.n2933 9.3005
R9883 gnd.n2633 gnd.n2632 9.3005
R9884 gnd.n3050 gnd.n3049 9.3005
R9885 gnd.n3051 gnd.n2631 9.3005
R9886 gnd.n3055 gnd.n3052 9.3005
R9887 gnd.n3054 gnd.n3053 9.3005
R9888 gnd.n2555 gnd.n2554 9.3005
R9889 gnd.n3130 gnd.n3129 9.3005
R9890 gnd.n2887 gnd.n2788 9.3005
R9891 gnd.n2790 gnd.n2789 9.3005
R9892 gnd.n2834 gnd.n2832 9.3005
R9893 gnd.n2835 gnd.n2831 9.3005
R9894 gnd.n2838 gnd.n2827 9.3005
R9895 gnd.n2839 gnd.n2826 9.3005
R9896 gnd.n2842 gnd.n2825 9.3005
R9897 gnd.n2843 gnd.n2824 9.3005
R9898 gnd.n2846 gnd.n2823 9.3005
R9899 gnd.n2847 gnd.n2822 9.3005
R9900 gnd.n2850 gnd.n2821 9.3005
R9901 gnd.n2851 gnd.n2820 9.3005
R9902 gnd.n2854 gnd.n2819 9.3005
R9903 gnd.n2855 gnd.n2818 9.3005
R9904 gnd.n2858 gnd.n2817 9.3005
R9905 gnd.n2859 gnd.n2816 9.3005
R9906 gnd.n2862 gnd.n2815 9.3005
R9907 gnd.n2863 gnd.n2814 9.3005
R9908 gnd.n2866 gnd.n2813 9.3005
R9909 gnd.n2867 gnd.n2812 9.3005
R9910 gnd.n2870 gnd.n2811 9.3005
R9911 gnd.n2871 gnd.n2810 9.3005
R9912 gnd.n2874 gnd.n2809 9.3005
R9913 gnd.n2876 gnd.n2808 9.3005
R9914 gnd.n2877 gnd.n2807 9.3005
R9915 gnd.n2878 gnd.n2806 9.3005
R9916 gnd.n2879 gnd.n2805 9.3005
R9917 gnd.n2886 gnd.n2885 9.3005
R9918 gnd.n2895 gnd.n2894 9.3005
R9919 gnd.n2896 gnd.n2782 9.3005
R9920 gnd.n2898 gnd.n2897 9.3005
R9921 gnd.n2773 gnd.n2772 9.3005
R9922 gnd.n2911 gnd.n2910 9.3005
R9923 gnd.n2912 gnd.n2771 9.3005
R9924 gnd.n2914 gnd.n2913 9.3005
R9925 gnd.n2760 gnd.n2759 9.3005
R9926 gnd.n2957 gnd.n2956 9.3005
R9927 gnd.n2958 gnd.n2714 9.3005
R9928 gnd.n2962 gnd.n2960 9.3005
R9929 gnd.n2961 gnd.n2693 9.3005
R9930 gnd.n2980 gnd.n2692 9.3005
R9931 gnd.n2983 gnd.n2982 9.3005
R9932 gnd.n2686 gnd.n2685 9.3005
R9933 gnd.n2994 gnd.n2992 9.3005
R9934 gnd.n2993 gnd.n2667 9.3005
R9935 gnd.n3011 gnd.n2666 9.3005
R9936 gnd.n3014 gnd.n3013 9.3005
R9937 gnd.n2661 gnd.n2656 9.3005
R9938 gnd.n3024 gnd.n3023 9.3005
R9939 gnd.n2659 gnd.n2639 9.3005
R9940 gnd.n3045 gnd.n2640 9.3005
R9941 gnd.n3044 gnd.n3043 9.3005
R9942 gnd.n2642 gnd.n2618 9.3005
R9943 gnd.n3076 gnd.n3075 9.3005
R9944 gnd.n3078 gnd.n2563 9.3005
R9945 gnd.n3125 gnd.n2564 9.3005
R9946 gnd.n3124 gnd.n2565 9.3005
R9947 gnd.n3123 gnd.n2566 9.3005
R9948 gnd.n3089 gnd.n2567 9.3005
R9949 gnd.n3091 gnd.n2585 9.3005
R9950 gnd.n3111 gnd.n2586 9.3005
R9951 gnd.n3110 gnd.n2587 9.3005
R9952 gnd.n3109 gnd.n2588 9.3005
R9953 gnd.n3100 gnd.n2589 9.3005
R9954 gnd.n3101 gnd.n2488 9.3005
R9955 gnd.n3167 gnd.n3166 9.3005
R9956 gnd.n3168 gnd.n2481 9.3005
R9957 gnd.n3178 gnd.n3177 9.3005
R9958 gnd.n3180 gnd.n2477 9.3005
R9959 gnd.n3190 gnd.n2478 9.3005
R9960 gnd.n3189 gnd.n3188 9.3005
R9961 gnd.n3186 gnd.n2456 9.3005
R9962 gnd.n3212 gnd.n2457 9.3005
R9963 gnd.n3211 gnd.n3210 9.3005
R9964 gnd.n2459 gnd.n2433 9.3005
R9965 gnd.n3252 gnd.n3251 9.3005
R9966 gnd.n3253 gnd.n2426 9.3005
R9967 gnd.n3263 gnd.n3262 9.3005
R9968 gnd.n3265 gnd.n2422 9.3005
R9969 gnd.n3275 gnd.n2423 9.3005
R9970 gnd.n3274 gnd.n3273 9.3005
R9971 gnd.n3271 gnd.n2401 9.3005
R9972 gnd.n3297 gnd.n2402 9.3005
R9973 gnd.n3296 gnd.n3295 9.3005
R9974 gnd.n2404 gnd.n2379 9.3005
R9975 gnd.n3341 gnd.n3340 9.3005
R9976 gnd.n3342 gnd.n2372 9.3005
R9977 gnd.n3353 gnd.n3352 9.3005
R9978 gnd.n3611 gnd.n2368 9.3005
R9979 gnd.n3619 gnd.n2369 9.3005
R9980 gnd.n3618 gnd.n3617 9.3005
R9981 gnd.n2350 gnd.n2349 9.3005
R9982 gnd.n3642 gnd.n3641 9.3005
R9983 gnd.n2784 gnd.n2783 9.3005
R9984 gnd.n6185 gnd.n880 9.3005
R9985 gnd.n6187 gnd.n6186 9.3005
R9986 gnd.n876 gnd.n875 9.3005
R9987 gnd.n6194 gnd.n6193 9.3005
R9988 gnd.n6195 gnd.n874 9.3005
R9989 gnd.n6197 gnd.n6196 9.3005
R9990 gnd.n870 gnd.n869 9.3005
R9991 gnd.n6204 gnd.n6203 9.3005
R9992 gnd.n6205 gnd.n868 9.3005
R9993 gnd.n6207 gnd.n6206 9.3005
R9994 gnd.n864 gnd.n863 9.3005
R9995 gnd.n6214 gnd.n6213 9.3005
R9996 gnd.n6215 gnd.n862 9.3005
R9997 gnd.n6217 gnd.n6216 9.3005
R9998 gnd.n858 gnd.n857 9.3005
R9999 gnd.n6224 gnd.n6223 9.3005
R10000 gnd.n6225 gnd.n856 9.3005
R10001 gnd.n6227 gnd.n6226 9.3005
R10002 gnd.n852 gnd.n851 9.3005
R10003 gnd.n6234 gnd.n6233 9.3005
R10004 gnd.n6235 gnd.n850 9.3005
R10005 gnd.n6237 gnd.n6236 9.3005
R10006 gnd.n846 gnd.n845 9.3005
R10007 gnd.n6244 gnd.n6243 9.3005
R10008 gnd.n6245 gnd.n844 9.3005
R10009 gnd.n6247 gnd.n6246 9.3005
R10010 gnd.n840 gnd.n839 9.3005
R10011 gnd.n6254 gnd.n6253 9.3005
R10012 gnd.n6255 gnd.n838 9.3005
R10013 gnd.n6257 gnd.n6256 9.3005
R10014 gnd.n834 gnd.n833 9.3005
R10015 gnd.n6264 gnd.n6263 9.3005
R10016 gnd.n6265 gnd.n832 9.3005
R10017 gnd.n6267 gnd.n6266 9.3005
R10018 gnd.n828 gnd.n827 9.3005
R10019 gnd.n6274 gnd.n6273 9.3005
R10020 gnd.n6275 gnd.n826 9.3005
R10021 gnd.n6277 gnd.n6276 9.3005
R10022 gnd.n822 gnd.n821 9.3005
R10023 gnd.n6284 gnd.n6283 9.3005
R10024 gnd.n6285 gnd.n820 9.3005
R10025 gnd.n6287 gnd.n6286 9.3005
R10026 gnd.n816 gnd.n815 9.3005
R10027 gnd.n6294 gnd.n6293 9.3005
R10028 gnd.n6295 gnd.n814 9.3005
R10029 gnd.n6297 gnd.n6296 9.3005
R10030 gnd.n810 gnd.n809 9.3005
R10031 gnd.n6304 gnd.n6303 9.3005
R10032 gnd.n6305 gnd.n808 9.3005
R10033 gnd.n6307 gnd.n6306 9.3005
R10034 gnd.n804 gnd.n803 9.3005
R10035 gnd.n6314 gnd.n6313 9.3005
R10036 gnd.n6315 gnd.n802 9.3005
R10037 gnd.n6317 gnd.n6316 9.3005
R10038 gnd.n798 gnd.n797 9.3005
R10039 gnd.n6324 gnd.n6323 9.3005
R10040 gnd.n6325 gnd.n796 9.3005
R10041 gnd.n6327 gnd.n6326 9.3005
R10042 gnd.n792 gnd.n791 9.3005
R10043 gnd.n6334 gnd.n6333 9.3005
R10044 gnd.n6335 gnd.n790 9.3005
R10045 gnd.n6337 gnd.n6336 9.3005
R10046 gnd.n786 gnd.n785 9.3005
R10047 gnd.n6344 gnd.n6343 9.3005
R10048 gnd.n6345 gnd.n784 9.3005
R10049 gnd.n6347 gnd.n6346 9.3005
R10050 gnd.n780 gnd.n779 9.3005
R10051 gnd.n6354 gnd.n6353 9.3005
R10052 gnd.n6355 gnd.n778 9.3005
R10053 gnd.n6357 gnd.n6356 9.3005
R10054 gnd.n774 gnd.n773 9.3005
R10055 gnd.n6364 gnd.n6363 9.3005
R10056 gnd.n6365 gnd.n772 9.3005
R10057 gnd.n6367 gnd.n6366 9.3005
R10058 gnd.n768 gnd.n767 9.3005
R10059 gnd.n6374 gnd.n6373 9.3005
R10060 gnd.n6375 gnd.n766 9.3005
R10061 gnd.n6377 gnd.n6376 9.3005
R10062 gnd.n762 gnd.n761 9.3005
R10063 gnd.n6384 gnd.n6383 9.3005
R10064 gnd.n6385 gnd.n760 9.3005
R10065 gnd.n6387 gnd.n6386 9.3005
R10066 gnd.n756 gnd.n755 9.3005
R10067 gnd.n6394 gnd.n6393 9.3005
R10068 gnd.n6395 gnd.n754 9.3005
R10069 gnd.n6397 gnd.n6396 9.3005
R10070 gnd.n750 gnd.n749 9.3005
R10071 gnd.n6404 gnd.n6403 9.3005
R10072 gnd.n6405 gnd.n748 9.3005
R10073 gnd.n6407 gnd.n6406 9.3005
R10074 gnd.n744 gnd.n743 9.3005
R10075 gnd.n6414 gnd.n6413 9.3005
R10076 gnd.n6415 gnd.n742 9.3005
R10077 gnd.n6417 gnd.n6416 9.3005
R10078 gnd.n738 gnd.n737 9.3005
R10079 gnd.n6424 gnd.n6423 9.3005
R10080 gnd.n6425 gnd.n736 9.3005
R10081 gnd.n6427 gnd.n6426 9.3005
R10082 gnd.n732 gnd.n731 9.3005
R10083 gnd.n6434 gnd.n6433 9.3005
R10084 gnd.n6435 gnd.n730 9.3005
R10085 gnd.n6437 gnd.n6436 9.3005
R10086 gnd.n726 gnd.n725 9.3005
R10087 gnd.n6444 gnd.n6443 9.3005
R10088 gnd.n6445 gnd.n724 9.3005
R10089 gnd.n6447 gnd.n6446 9.3005
R10090 gnd.n720 gnd.n719 9.3005
R10091 gnd.n6454 gnd.n6453 9.3005
R10092 gnd.n6455 gnd.n718 9.3005
R10093 gnd.n6457 gnd.n6456 9.3005
R10094 gnd.n714 gnd.n713 9.3005
R10095 gnd.n6464 gnd.n6463 9.3005
R10096 gnd.n6465 gnd.n712 9.3005
R10097 gnd.n6467 gnd.n6466 9.3005
R10098 gnd.n708 gnd.n707 9.3005
R10099 gnd.n6474 gnd.n6473 9.3005
R10100 gnd.n6475 gnd.n706 9.3005
R10101 gnd.n6477 gnd.n6476 9.3005
R10102 gnd.n702 gnd.n701 9.3005
R10103 gnd.n6484 gnd.n6483 9.3005
R10104 gnd.n6485 gnd.n700 9.3005
R10105 gnd.n6487 gnd.n6486 9.3005
R10106 gnd.n696 gnd.n695 9.3005
R10107 gnd.n6494 gnd.n6493 9.3005
R10108 gnd.n6495 gnd.n694 9.3005
R10109 gnd.n6498 gnd.n6497 9.3005
R10110 gnd.n6496 gnd.n690 9.3005
R10111 gnd.n6504 gnd.n689 9.3005
R10112 gnd.n6506 gnd.n6505 9.3005
R10113 gnd.n685 gnd.n684 9.3005
R10114 gnd.n6515 gnd.n6514 9.3005
R10115 gnd.n6516 gnd.n683 9.3005
R10116 gnd.n6518 gnd.n6517 9.3005
R10117 gnd.n679 gnd.n678 9.3005
R10118 gnd.n6525 gnd.n6524 9.3005
R10119 gnd.n6526 gnd.n677 9.3005
R10120 gnd.n6528 gnd.n6527 9.3005
R10121 gnd.n673 gnd.n672 9.3005
R10122 gnd.n6535 gnd.n6534 9.3005
R10123 gnd.n6536 gnd.n671 9.3005
R10124 gnd.n6538 gnd.n6537 9.3005
R10125 gnd.n667 gnd.n666 9.3005
R10126 gnd.n6545 gnd.n6544 9.3005
R10127 gnd.n6546 gnd.n665 9.3005
R10128 gnd.n6548 gnd.n6547 9.3005
R10129 gnd.n661 gnd.n660 9.3005
R10130 gnd.n6555 gnd.n6554 9.3005
R10131 gnd.n6556 gnd.n659 9.3005
R10132 gnd.n6558 gnd.n6557 9.3005
R10133 gnd.n655 gnd.n654 9.3005
R10134 gnd.n6565 gnd.n6564 9.3005
R10135 gnd.n6566 gnd.n653 9.3005
R10136 gnd.n6568 gnd.n6567 9.3005
R10137 gnd.n649 gnd.n648 9.3005
R10138 gnd.n6575 gnd.n6574 9.3005
R10139 gnd.n6576 gnd.n647 9.3005
R10140 gnd.n6578 gnd.n6577 9.3005
R10141 gnd.n643 gnd.n642 9.3005
R10142 gnd.n6585 gnd.n6584 9.3005
R10143 gnd.n6586 gnd.n641 9.3005
R10144 gnd.n6588 gnd.n6587 9.3005
R10145 gnd.n637 gnd.n636 9.3005
R10146 gnd.n6595 gnd.n6594 9.3005
R10147 gnd.n6596 gnd.n635 9.3005
R10148 gnd.n6598 gnd.n6597 9.3005
R10149 gnd.n631 gnd.n630 9.3005
R10150 gnd.n6605 gnd.n6604 9.3005
R10151 gnd.n6606 gnd.n629 9.3005
R10152 gnd.n6608 gnd.n6607 9.3005
R10153 gnd.n625 gnd.n624 9.3005
R10154 gnd.n6615 gnd.n6614 9.3005
R10155 gnd.n6616 gnd.n623 9.3005
R10156 gnd.n6618 gnd.n6617 9.3005
R10157 gnd.n619 gnd.n618 9.3005
R10158 gnd.n6625 gnd.n6624 9.3005
R10159 gnd.n6626 gnd.n617 9.3005
R10160 gnd.n6628 gnd.n6627 9.3005
R10161 gnd.n613 gnd.n612 9.3005
R10162 gnd.n6635 gnd.n6634 9.3005
R10163 gnd.n6636 gnd.n611 9.3005
R10164 gnd.n6638 gnd.n6637 9.3005
R10165 gnd.n607 gnd.n606 9.3005
R10166 gnd.n6645 gnd.n6644 9.3005
R10167 gnd.n6646 gnd.n605 9.3005
R10168 gnd.n6648 gnd.n6647 9.3005
R10169 gnd.n601 gnd.n600 9.3005
R10170 gnd.n6655 gnd.n6654 9.3005
R10171 gnd.n6656 gnd.n599 9.3005
R10172 gnd.n6658 gnd.n6657 9.3005
R10173 gnd.n595 gnd.n594 9.3005
R10174 gnd.n6665 gnd.n6664 9.3005
R10175 gnd.n6666 gnd.n593 9.3005
R10176 gnd.n6668 gnd.n6667 9.3005
R10177 gnd.n589 gnd.n588 9.3005
R10178 gnd.n6675 gnd.n6674 9.3005
R10179 gnd.n6676 gnd.n587 9.3005
R10180 gnd.n6678 gnd.n6677 9.3005
R10181 gnd.n583 gnd.n582 9.3005
R10182 gnd.n6685 gnd.n6684 9.3005
R10183 gnd.n6686 gnd.n581 9.3005
R10184 gnd.n6688 gnd.n6687 9.3005
R10185 gnd.n577 gnd.n576 9.3005
R10186 gnd.n6695 gnd.n6694 9.3005
R10187 gnd.n6696 gnd.n575 9.3005
R10188 gnd.n6698 gnd.n6697 9.3005
R10189 gnd.n571 gnd.n570 9.3005
R10190 gnd.n6705 gnd.n6704 9.3005
R10191 gnd.n6706 gnd.n569 9.3005
R10192 gnd.n6708 gnd.n6707 9.3005
R10193 gnd.n565 gnd.n564 9.3005
R10194 gnd.n6716 gnd.n6715 9.3005
R10195 gnd.n6717 gnd.n563 9.3005
R10196 gnd.n6719 gnd.n6718 9.3005
R10197 gnd.n6508 gnd.n6507 9.3005
R10198 gnd.n6901 gnd.n6900 9.3005
R10199 gnd.n6899 gnd.n65 9.3005
R10200 gnd.n214 gnd.n67 9.3005
R10201 gnd.n217 gnd.n215 9.3005
R10202 gnd.n219 gnd.n218 9.3005
R10203 gnd.n220 gnd.n213 9.3005
R10204 gnd.n222 gnd.n221 9.3005
R10205 gnd.n224 gnd.n211 9.3005
R10206 gnd.n226 gnd.n225 9.3005
R10207 gnd.n227 gnd.n210 9.3005
R10208 gnd.n229 gnd.n228 9.3005
R10209 gnd.n231 gnd.n208 9.3005
R10210 gnd.n233 gnd.n232 9.3005
R10211 gnd.n234 gnd.n207 9.3005
R10212 gnd.n236 gnd.n235 9.3005
R10213 gnd.n238 gnd.n205 9.3005
R10214 gnd.n240 gnd.n239 9.3005
R10215 gnd.n241 gnd.n204 9.3005
R10216 gnd.n243 gnd.n242 9.3005
R10217 gnd.n245 gnd.n202 9.3005
R10218 gnd.n247 gnd.n246 9.3005
R10219 gnd.n278 gnd.n168 9.3005
R10220 gnd.n277 gnd.n170 9.3005
R10221 gnd.n174 gnd.n171 9.3005
R10222 gnd.n272 gnd.n175 9.3005
R10223 gnd.n271 gnd.n176 9.3005
R10224 gnd.n270 gnd.n177 9.3005
R10225 gnd.n181 gnd.n178 9.3005
R10226 gnd.n265 gnd.n182 9.3005
R10227 gnd.n264 gnd.n183 9.3005
R10228 gnd.n263 gnd.n184 9.3005
R10229 gnd.n188 gnd.n185 9.3005
R10230 gnd.n258 gnd.n189 9.3005
R10231 gnd.n257 gnd.n190 9.3005
R10232 gnd.n256 gnd.n191 9.3005
R10233 gnd.n195 gnd.n192 9.3005
R10234 gnd.n251 gnd.n196 9.3005
R10235 gnd.n250 gnd.n249 9.3005
R10236 gnd.n248 gnd.n199 9.3005
R10237 gnd.n280 gnd.n279 9.3005
R10238 gnd.n346 gnd.n343 9.3005
R10239 gnd.n352 gnd.n351 9.3005
R10240 gnd.n353 gnd.n342 9.3005
R10241 gnd.n355 gnd.n354 9.3005
R10242 gnd.n340 gnd.n339 9.3005
R10243 gnd.n362 gnd.n361 9.3005
R10244 gnd.n363 gnd.n338 9.3005
R10245 gnd.n365 gnd.n364 9.3005
R10246 gnd.n336 gnd.n335 9.3005
R10247 gnd.n372 gnd.n371 9.3005
R10248 gnd.n373 gnd.n334 9.3005
R10249 gnd.n375 gnd.n374 9.3005
R10250 gnd.n332 gnd.n331 9.3005
R10251 gnd.n383 gnd.n382 9.3005
R10252 gnd.n384 gnd.n330 9.3005
R10253 gnd.n386 gnd.n385 9.3005
R10254 gnd.n387 gnd.n325 9.3005
R10255 gnd.n393 gnd.n392 9.3005
R10256 gnd.n394 gnd.n324 9.3005
R10257 gnd.n396 gnd.n395 9.3005
R10258 gnd.n322 gnd.n321 9.3005
R10259 gnd.n403 gnd.n402 9.3005
R10260 gnd.n404 gnd.n320 9.3005
R10261 gnd.n406 gnd.n405 9.3005
R10262 gnd.n318 gnd.n317 9.3005
R10263 gnd.n413 gnd.n412 9.3005
R10264 gnd.n414 gnd.n316 9.3005
R10265 gnd.n416 gnd.n415 9.3005
R10266 gnd.n314 gnd.n313 9.3005
R10267 gnd.n423 gnd.n422 9.3005
R10268 gnd.n424 gnd.n312 9.3005
R10269 gnd.n426 gnd.n425 9.3005
R10270 gnd.n310 gnd.n309 9.3005
R10271 gnd.n433 gnd.n432 9.3005
R10272 gnd.n434 gnd.n308 9.3005
R10273 gnd.n436 gnd.n435 9.3005
R10274 gnd.n306 gnd.n303 9.3005
R10275 gnd.n443 gnd.n442 9.3005
R10276 gnd.n444 gnd.n302 9.3005
R10277 gnd.n446 gnd.n445 9.3005
R10278 gnd.n300 gnd.n299 9.3005
R10279 gnd.n453 gnd.n452 9.3005
R10280 gnd.n454 gnd.n298 9.3005
R10281 gnd.n456 gnd.n455 9.3005
R10282 gnd.n296 gnd.n295 9.3005
R10283 gnd.n463 gnd.n462 9.3005
R10284 gnd.n464 gnd.n294 9.3005
R10285 gnd.n466 gnd.n465 9.3005
R10286 gnd.n292 gnd.n291 9.3005
R10287 gnd.n473 gnd.n472 9.3005
R10288 gnd.n474 gnd.n290 9.3005
R10289 gnd.n476 gnd.n475 9.3005
R10290 gnd.n288 gnd.n287 9.3005
R10291 gnd.n483 gnd.n482 9.3005
R10292 gnd.n484 gnd.n286 9.3005
R10293 gnd.n486 gnd.n485 9.3005
R10294 gnd.n284 gnd.n281 9.3005
R10295 gnd.n492 gnd.n491 9.3005
R10296 gnd.n345 gnd.n344 9.3005
R10297 gnd.n5529 gnd.n5528 9.3005
R10298 gnd.n1564 gnd.n1563 9.3005
R10299 gnd.n1588 gnd.n1587 9.3005
R10300 gnd.n5516 gnd.n1589 9.3005
R10301 gnd.n5515 gnd.n1590 9.3005
R10302 gnd.n5514 gnd.n1591 9.3005
R10303 gnd.n5445 gnd.n1592 9.3005
R10304 gnd.n5504 gnd.n1611 9.3005
R10305 gnd.n5503 gnd.n5502 9.3005
R10306 gnd.n1612 gnd.n552 9.3005
R10307 gnd.n6734 gnd.n553 9.3005
R10308 gnd.n6733 gnd.n554 9.3005
R10309 gnd.n6732 gnd.n555 9.3005
R10310 gnd.n6731 gnd.n556 9.3005
R10311 gnd.n529 gnd.n525 9.3005
R10312 gnd.n6767 gnd.n526 9.3005
R10313 gnd.n6766 gnd.n527 9.3005
R10314 gnd.n6765 gnd.n6763 9.3005
R10315 gnd.n503 gnd.n502 9.3005
R10316 gnd.n6793 gnd.n6792 9.3005
R10317 gnd.n6794 gnd.n496 9.3005
R10318 gnd.n6801 gnd.n497 9.3005
R10319 gnd.n6802 gnd.n495 9.3005
R10320 gnd.n6805 gnd.n6804 9.3005
R10321 gnd.n6806 gnd.n91 9.3005
R10322 gnd.n6887 gnd.n92 9.3005
R10323 gnd.n6886 gnd.n93 9.3005
R10324 gnd.n6885 gnd.n94 9.3005
R10325 gnd.n6814 gnd.n95 9.3005
R10326 gnd.n6875 gnd.n109 9.3005
R10327 gnd.n6874 gnd.n110 9.3005
R10328 gnd.n6873 gnd.n111 9.3005
R10329 gnd.n6821 gnd.n112 9.3005
R10330 gnd.n6863 gnd.n129 9.3005
R10331 gnd.n6862 gnd.n130 9.3005
R10332 gnd.n6861 gnd.n131 9.3005
R10333 gnd.n6828 gnd.n132 9.3005
R10334 gnd.n6851 gnd.n149 9.3005
R10335 gnd.n6850 gnd.n150 9.3005
R10336 gnd.n6849 gnd.n151 9.3005
R10337 gnd.n167 gnd.n152 9.3005
R10338 gnd.n6839 gnd.n6838 9.3005
R10339 gnd.n5530 gnd.n1562 9.3005
R10340 gnd.n5528 gnd.n5527 9.3005
R10341 gnd.n5526 gnd.n1564 9.3005
R10342 gnd.n1588 gnd.n1565 9.3005
R10343 gnd.n5440 gnd.n1589 9.3005
R10344 gnd.n5443 gnd.n1590 9.3005
R10345 gnd.n5444 gnd.n1591 9.3005
R10346 gnd.n5446 gnd.n5445 9.3005
R10347 gnd.n1613 gnd.n1611 9.3005
R10348 gnd.n5502 gnd.n5501 9.3005
R10349 gnd.n1619 gnd.n1612 9.3005
R10350 gnd.n1618 gnd.n553 9.3005
R10351 gnd.n1617 gnd.n554 9.3005
R10352 gnd.n1614 gnd.n555 9.3005
R10353 gnd.n556 gnd.n528 9.3005
R10354 gnd.n6757 gnd.n529 9.3005
R10355 gnd.n6758 gnd.n526 9.3005
R10356 gnd.n6759 gnd.n527 9.3005
R10357 gnd.n6763 gnd.n6762 9.3005
R10358 gnd.n6760 gnd.n502 9.3005
R10359 gnd.n6793 gnd.n501 9.3005
R10360 gnd.n6795 gnd.n6794 9.3005
R10361 gnd.n6797 gnd.n497 9.3005
R10362 gnd.n6796 gnd.n495 9.3005
R10363 gnd.n6805 gnd.n494 9.3005
R10364 gnd.n6809 gnd.n6806 9.3005
R10365 gnd.n6810 gnd.n92 9.3005
R10366 gnd.n6812 gnd.n93 9.3005
R10367 gnd.n6813 gnd.n94 9.3005
R10368 gnd.n6816 gnd.n6814 9.3005
R10369 gnd.n6817 gnd.n109 9.3005
R10370 gnd.n6819 gnd.n110 9.3005
R10371 gnd.n6820 gnd.n111 9.3005
R10372 gnd.n6823 gnd.n6821 9.3005
R10373 gnd.n6824 gnd.n129 9.3005
R10374 gnd.n6826 gnd.n130 9.3005
R10375 gnd.n6827 gnd.n131 9.3005
R10376 gnd.n6830 gnd.n6828 9.3005
R10377 gnd.n6831 gnd.n149 9.3005
R10378 gnd.n6833 gnd.n150 9.3005
R10379 gnd.n6834 gnd.n151 9.3005
R10380 gnd.n6836 gnd.n167 9.3005
R10381 gnd.n6838 gnd.n6837 9.3005
R10382 gnd.n1562 gnd.n1556 9.3005
R10383 gnd.n5540 gnd.n5539 9.3005
R10384 gnd.n5543 gnd.n1554 9.3005
R10385 gnd.n5544 gnd.n1553 9.3005
R10386 gnd.n5547 gnd.n1552 9.3005
R10387 gnd.n5548 gnd.n1551 9.3005
R10388 gnd.n5551 gnd.n1550 9.3005
R10389 gnd.n5552 gnd.n1549 9.3005
R10390 gnd.n5555 gnd.n1548 9.3005
R10391 gnd.n5556 gnd.n1547 9.3005
R10392 gnd.n5559 gnd.n1546 9.3005
R10393 gnd.n5560 gnd.n1545 9.3005
R10394 gnd.n5563 gnd.n1544 9.3005
R10395 gnd.n5564 gnd.n1543 9.3005
R10396 gnd.n5567 gnd.n1542 9.3005
R10397 gnd.n5568 gnd.n1541 9.3005
R10398 gnd.n5571 gnd.n1540 9.3005
R10399 gnd.n5572 gnd.n1539 9.3005
R10400 gnd.n5575 gnd.n1538 9.3005
R10401 gnd.n5576 gnd.n1537 9.3005
R10402 gnd.n5579 gnd.n1536 9.3005
R10403 gnd.n5583 gnd.n1532 9.3005
R10404 gnd.n5584 gnd.n1531 9.3005
R10405 gnd.n5587 gnd.n1530 9.3005
R10406 gnd.n5588 gnd.n1529 9.3005
R10407 gnd.n5591 gnd.n1528 9.3005
R10408 gnd.n5592 gnd.n1527 9.3005
R10409 gnd.n5595 gnd.n1526 9.3005
R10410 gnd.n5596 gnd.n1525 9.3005
R10411 gnd.n5599 gnd.n1524 9.3005
R10412 gnd.n5601 gnd.n1520 9.3005
R10413 gnd.n5604 gnd.n1519 9.3005
R10414 gnd.n5605 gnd.n1518 9.3005
R10415 gnd.n5608 gnd.n1517 9.3005
R10416 gnd.n5609 gnd.n1516 9.3005
R10417 gnd.n5612 gnd.n1515 9.3005
R10418 gnd.n5613 gnd.n1514 9.3005
R10419 gnd.n5616 gnd.n1513 9.3005
R10420 gnd.n5618 gnd.n1510 9.3005
R10421 gnd.n5621 gnd.n1509 9.3005
R10422 gnd.n5622 gnd.n1508 9.3005
R10423 gnd.n5625 gnd.n1507 9.3005
R10424 gnd.n5626 gnd.n1506 9.3005
R10425 gnd.n5629 gnd.n1505 9.3005
R10426 gnd.n5630 gnd.n1504 9.3005
R10427 gnd.n5633 gnd.n1503 9.3005
R10428 gnd.n5634 gnd.n1502 9.3005
R10429 gnd.n5637 gnd.n1501 9.3005
R10430 gnd.n5638 gnd.n1500 9.3005
R10431 gnd.n5641 gnd.n1499 9.3005
R10432 gnd.n5642 gnd.n1498 9.3005
R10433 gnd.n5645 gnd.n1497 9.3005
R10434 gnd.n5647 gnd.n1496 9.3005
R10435 gnd.n5648 gnd.n1495 9.3005
R10436 gnd.n5649 gnd.n1494 9.3005
R10437 gnd.n5650 gnd.n1493 9.3005
R10438 gnd.n5580 gnd.n1533 9.3005
R10439 gnd.n5538 gnd.n5535 9.3005
R10440 gnd.n1575 gnd.n1572 9.3005
R10441 gnd.n5522 gnd.n1576 9.3005
R10442 gnd.n5521 gnd.n1577 9.3005
R10443 gnd.n5520 gnd.n1578 9.3005
R10444 gnd.n1599 gnd.n1579 9.3005
R10445 gnd.n5510 gnd.n1600 9.3005
R10446 gnd.n5509 gnd.n1601 9.3005
R10447 gnd.n5508 gnd.n1602 9.3005
R10448 gnd.n1604 gnd.n1603 9.3005
R10449 gnd.n544 gnd.n543 9.3005
R10450 gnd.n6739 gnd.n6738 9.3005
R10451 gnd.n6740 gnd.n542 9.3005
R10452 gnd.n6745 gnd.n6741 9.3005
R10453 gnd.n6744 gnd.n6742 9.3005
R10454 gnd.n6743 gnd.n77 9.3005
R10455 gnd.n82 gnd.n76 9.3005
R10456 gnd.n6881 gnd.n101 9.3005
R10457 gnd.n6880 gnd.n102 9.3005
R10458 gnd.n6879 gnd.n103 9.3005
R10459 gnd.n118 gnd.n104 9.3005
R10460 gnd.n6869 gnd.n119 9.3005
R10461 gnd.n6868 gnd.n120 9.3005
R10462 gnd.n6867 gnd.n121 9.3005
R10463 gnd.n138 gnd.n122 9.3005
R10464 gnd.n6857 gnd.n139 9.3005
R10465 gnd.n6856 gnd.n140 9.3005
R10466 gnd.n6855 gnd.n141 9.3005
R10467 gnd.n157 gnd.n142 9.3005
R10468 gnd.n6845 gnd.n158 9.3005
R10469 gnd.n6844 gnd.n159 9.3005
R10470 gnd.n6843 gnd.n160 9.3005
R10471 gnd.n1574 gnd.n1573 9.3005
R10472 gnd.n6892 gnd.n6891 9.3005
R10473 gnd.n6724 gnd.n6723 9.3005
R10474 gnd.n4234 gnd.n4233 9.3005
R10475 gnd.n4235 gnd.n4228 9.3005
R10476 gnd.n4237 gnd.n4236 9.3005
R10477 gnd.n2153 gnd.n2152 9.3005
R10478 gnd.n4242 gnd.n4241 9.3005
R10479 gnd.n4243 gnd.n2151 9.3005
R10480 gnd.n4249 gnd.n4244 9.3005
R10481 gnd.n4248 gnd.n4245 9.3005
R10482 gnd.n4247 gnd.n4246 9.3005
R10483 gnd.n2135 gnd.n2134 9.3005
R10484 gnd.n4547 gnd.n4546 9.3005
R10485 gnd.n4548 gnd.n2133 9.3005
R10486 gnd.n4550 gnd.n4549 9.3005
R10487 gnd.n2131 gnd.n2130 9.3005
R10488 gnd.n4555 gnd.n4554 9.3005
R10489 gnd.n4556 gnd.n2129 9.3005
R10490 gnd.n4566 gnd.n4557 9.3005
R10491 gnd.n4565 gnd.n4558 9.3005
R10492 gnd.n4564 gnd.n4559 9.3005
R10493 gnd.n4561 gnd.n4560 9.3005
R10494 gnd.n2101 gnd.n2100 9.3005
R10495 gnd.n4583 gnd.n4582 9.3005
R10496 gnd.n4584 gnd.n2099 9.3005
R10497 gnd.n4586 gnd.n4585 9.3005
R10498 gnd.n2087 gnd.n2086 9.3005
R10499 gnd.n4599 gnd.n4598 9.3005
R10500 gnd.n4600 gnd.n2085 9.3005
R10501 gnd.n4602 gnd.n4601 9.3005
R10502 gnd.n2071 gnd.n2070 9.3005
R10503 gnd.n4632 gnd.n4631 9.3005
R10504 gnd.n4633 gnd.n2069 9.3005
R10505 gnd.n4644 gnd.n4634 9.3005
R10506 gnd.n4643 gnd.n4635 9.3005
R10507 gnd.n4642 gnd.n4636 9.3005
R10508 gnd.n4639 gnd.n4638 9.3005
R10509 gnd.n4637 gnd.n1283 9.3005
R10510 gnd.n5829 gnd.n1284 9.3005
R10511 gnd.n5828 gnd.n1285 9.3005
R10512 gnd.n5827 gnd.n1286 9.3005
R10513 gnd.n2032 gnd.n1287 9.3005
R10514 gnd.n2034 gnd.n2033 9.3005
R10515 gnd.n4799 gnd.n4798 9.3005
R10516 gnd.n4800 gnd.n2031 9.3005
R10517 gnd.n4804 gnd.n4801 9.3005
R10518 gnd.n4803 gnd.n4802 9.3005
R10519 gnd.n2010 gnd.n2009 9.3005
R10520 gnd.n4831 gnd.n4830 9.3005
R10521 gnd.n4832 gnd.n2008 9.3005
R10522 gnd.n4834 gnd.n4833 9.3005
R10523 gnd.n1986 gnd.n1985 9.3005
R10524 gnd.n4870 gnd.n4869 9.3005
R10525 gnd.n4871 gnd.n1984 9.3005
R10526 gnd.n4873 gnd.n4872 9.3005
R10527 gnd.n1960 gnd.n1959 9.3005
R10528 gnd.n4910 gnd.n4909 9.3005
R10529 gnd.n4911 gnd.n1958 9.3005
R10530 gnd.n4915 gnd.n4912 9.3005
R10531 gnd.n4914 gnd.n4913 9.3005
R10532 gnd.n1933 gnd.n1932 9.3005
R10533 gnd.n4956 gnd.n4955 9.3005
R10534 gnd.n4957 gnd.n1931 9.3005
R10535 gnd.n4961 gnd.n4958 9.3005
R10536 gnd.n4960 gnd.n4959 9.3005
R10537 gnd.n1911 gnd.n1910 9.3005
R10538 gnd.n5009 gnd.n5008 9.3005
R10539 gnd.n5010 gnd.n1909 9.3005
R10540 gnd.n5014 gnd.n5011 9.3005
R10541 gnd.n5013 gnd.n5012 9.3005
R10542 gnd.n1885 gnd.n1884 9.3005
R10543 gnd.n5045 gnd.n5044 9.3005
R10544 gnd.n5046 gnd.n1883 9.3005
R10545 gnd.n5048 gnd.n5047 9.3005
R10546 gnd.n1859 gnd.n1858 9.3005
R10547 gnd.n5089 gnd.n5088 9.3005
R10548 gnd.n5090 gnd.n1857 9.3005
R10549 gnd.n5094 gnd.n5091 9.3005
R10550 gnd.n5093 gnd.n5092 9.3005
R10551 gnd.n1836 gnd.n1835 9.3005
R10552 gnd.n5148 gnd.n5147 9.3005
R10553 gnd.n5149 gnd.n1834 9.3005
R10554 gnd.n5151 gnd.n5150 9.3005
R10555 gnd.n1814 gnd.n1813 9.3005
R10556 gnd.n5178 gnd.n5177 9.3005
R10557 gnd.n5179 gnd.n1812 9.3005
R10558 gnd.n5181 gnd.n5180 9.3005
R10559 gnd.n1797 gnd.n1796 9.3005
R10560 gnd.n5207 gnd.n5206 9.3005
R10561 gnd.n5208 gnd.n1795 9.3005
R10562 gnd.n5210 gnd.n5209 9.3005
R10563 gnd.n1706 gnd.n1705 9.3005
R10564 gnd.n5354 gnd.n5353 9.3005
R10565 gnd.n5355 gnd.n1704 9.3005
R10566 gnd.n5357 gnd.n5356 9.3005
R10567 gnd.n1693 gnd.n1692 9.3005
R10568 gnd.n5370 gnd.n5369 9.3005
R10569 gnd.n5371 gnd.n1691 9.3005
R10570 gnd.n5373 gnd.n5372 9.3005
R10571 gnd.n1680 gnd.n1679 9.3005
R10572 gnd.n5386 gnd.n5385 9.3005
R10573 gnd.n5387 gnd.n1678 9.3005
R10574 gnd.n5392 gnd.n5388 9.3005
R10575 gnd.n5391 gnd.n5390 9.3005
R10576 gnd.n5389 gnd.n1667 9.3005
R10577 gnd.n5405 gnd.n1666 9.3005
R10578 gnd.n5407 gnd.n5406 9.3005
R10579 gnd.n5408 gnd.n1665 9.3005
R10580 gnd.n5424 gnd.n5409 9.3005
R10581 gnd.n5423 gnd.n5410 9.3005
R10582 gnd.n5422 gnd.n5411 9.3005
R10583 gnd.n5413 gnd.n5412 9.3005
R10584 gnd.n5418 gnd.n5414 9.3005
R10585 gnd.n5417 gnd.n5416 9.3005
R10586 gnd.n5415 gnd.n1633 9.3005
R10587 gnd.n1631 gnd.n1630 9.3005
R10588 gnd.n5476 gnd.n5475 9.3005
R10589 gnd.n5477 gnd.n1629 9.3005
R10590 gnd.n5479 gnd.n5478 9.3005
R10591 gnd.n1627 gnd.n1626 9.3005
R10592 gnd.n5484 gnd.n5483 9.3005
R10593 gnd.n5485 gnd.n1625 9.3005
R10594 gnd.n5496 gnd.n5486 9.3005
R10595 gnd.n5495 gnd.n5487 9.3005
R10596 gnd.n5494 gnd.n5488 9.3005
R10597 gnd.n5491 gnd.n5490 9.3005
R10598 gnd.n5489 gnd.n559 9.3005
R10599 gnd.n6726 gnd.n560 9.3005
R10600 gnd.n6725 gnd.n561 9.3005
R10601 gnd.n3880 gnd.n3879 9.3005
R10602 gnd.n3910 gnd.n3857 9.3005
R10603 gnd.n3909 gnd.n3858 9.3005
R10604 gnd.n3907 gnd.n3859 9.3005
R10605 gnd.n3906 gnd.n3860 9.3005
R10606 gnd.n3904 gnd.n3861 9.3005
R10607 gnd.n3903 gnd.n3862 9.3005
R10608 gnd.n3901 gnd.n3863 9.3005
R10609 gnd.n3900 gnd.n3864 9.3005
R10610 gnd.n3898 gnd.n3865 9.3005
R10611 gnd.n3897 gnd.n3866 9.3005
R10612 gnd.n3895 gnd.n3867 9.3005
R10613 gnd.n3894 gnd.n3868 9.3005
R10614 gnd.n3892 gnd.n3869 9.3005
R10615 gnd.n3891 gnd.n3870 9.3005
R10616 gnd.n3889 gnd.n3871 9.3005
R10617 gnd.n3888 gnd.n3872 9.3005
R10618 gnd.n3886 gnd.n3873 9.3005
R10619 gnd.n3885 gnd.n3874 9.3005
R10620 gnd.n3883 gnd.n3875 9.3005
R10621 gnd.n3882 gnd.n3876 9.3005
R10622 gnd.n3913 gnd.n3912 9.3005
R10623 gnd.n3918 gnd.n3917 9.3005
R10624 gnd.n3921 gnd.n3852 9.3005
R10625 gnd.n3922 gnd.n3851 9.3005
R10626 gnd.n3925 gnd.n3850 9.3005
R10627 gnd.n3926 gnd.n3849 9.3005
R10628 gnd.n3929 gnd.n3848 9.3005
R10629 gnd.n3930 gnd.n3847 9.3005
R10630 gnd.n3933 gnd.n3846 9.3005
R10631 gnd.n3934 gnd.n3845 9.3005
R10632 gnd.n3937 gnd.n3844 9.3005
R10633 gnd.n3938 gnd.n3843 9.3005
R10634 gnd.n3941 gnd.n3842 9.3005
R10635 gnd.n3942 gnd.n3841 9.3005
R10636 gnd.n3945 gnd.n3840 9.3005
R10637 gnd.n3946 gnd.n3839 9.3005
R10638 gnd.n3949 gnd.n3838 9.3005
R10639 gnd.n3952 gnd.n3951 9.3005
R10640 gnd.n3916 gnd.n3856 9.3005
R10641 gnd.n3915 gnd.n3914 9.3005
R10642 gnd.n5907 gnd.n1210 9.3005
R10643 gnd.n5910 gnd.n1209 9.3005
R10644 gnd.n5911 gnd.n1208 9.3005
R10645 gnd.n5914 gnd.n1207 9.3005
R10646 gnd.n5915 gnd.n1206 9.3005
R10647 gnd.n5918 gnd.n1205 9.3005
R10648 gnd.n5919 gnd.n1204 9.3005
R10649 gnd.n5922 gnd.n1203 9.3005
R10650 gnd.n5924 gnd.n1200 9.3005
R10651 gnd.n5927 gnd.n1199 9.3005
R10652 gnd.n5928 gnd.n1198 9.3005
R10653 gnd.n5931 gnd.n1197 9.3005
R10654 gnd.n5932 gnd.n1196 9.3005
R10655 gnd.n5935 gnd.n1195 9.3005
R10656 gnd.n5936 gnd.n1194 9.3005
R10657 gnd.n5939 gnd.n1193 9.3005
R10658 gnd.n5940 gnd.n1192 9.3005
R10659 gnd.n5943 gnd.n1191 9.3005
R10660 gnd.n5944 gnd.n1190 9.3005
R10661 gnd.n5947 gnd.n1189 9.3005
R10662 gnd.n5948 gnd.n1188 9.3005
R10663 gnd.n5951 gnd.n1187 9.3005
R10664 gnd.n5952 gnd.n1186 9.3005
R10665 gnd.n5953 gnd.n1185 9.3005
R10666 gnd.n1142 gnd.n1141 9.3005
R10667 gnd.n5959 gnd.n5958 9.3005
R10668 gnd.n4451 gnd.n4448 9.3005
R10669 gnd.n4455 gnd.n4454 9.3005
R10670 gnd.n4456 gnd.n4446 9.3005
R10671 gnd.n4458 gnd.n4457 9.3005
R10672 gnd.n4461 gnd.n4445 9.3005
R10673 gnd.n4465 gnd.n4464 9.3005
R10674 gnd.n4466 gnd.n4444 9.3005
R10675 gnd.n4469 gnd.n4467 9.3005
R10676 gnd.n4470 gnd.n4440 9.3005
R10677 gnd.n4474 gnd.n4473 9.3005
R10678 gnd.n4475 gnd.n4439 9.3005
R10679 gnd.n4477 gnd.n4476 9.3005
R10680 gnd.n4480 gnd.n4438 9.3005
R10681 gnd.n4484 gnd.n4483 9.3005
R10682 gnd.n4485 gnd.n4437 9.3005
R10683 gnd.n4487 gnd.n4486 9.3005
R10684 gnd.n4490 gnd.n4436 9.3005
R10685 gnd.n4494 gnd.n4493 9.3005
R10686 gnd.n4495 gnd.n4435 9.3005
R10687 gnd.n4497 gnd.n4496 9.3005
R10688 gnd.n4500 gnd.n4434 9.3005
R10689 gnd.n4504 gnd.n4503 9.3005
R10690 gnd.n4505 gnd.n4433 9.3005
R10691 gnd.n4507 gnd.n4506 9.3005
R10692 gnd.n4510 gnd.n4432 9.3005
R10693 gnd.n4514 gnd.n4513 9.3005
R10694 gnd.n4515 gnd.n4431 9.3005
R10695 gnd.n4518 gnd.n4516 9.3005
R10696 gnd.n4519 gnd.n4427 9.3005
R10697 gnd.n4522 gnd.n4521 9.3005
R10698 gnd.n4447 gnd.n1211 9.3005
R10699 gnd.n4079 gnd.n4078 9.3005
R10700 gnd.n2270 gnd.n2266 9.3005
R10701 gnd.n2269 gnd.n2268 9.3005
R10702 gnd.n2250 gnd.n2247 9.3005
R10703 gnd.n4099 gnd.n2248 9.3005
R10704 gnd.n4098 gnd.n4095 9.3005
R10705 gnd.n4097 gnd.n4096 9.3005
R10706 gnd.n2232 gnd.n2229 9.3005
R10707 gnd.n4119 gnd.n2230 9.3005
R10708 gnd.n4118 gnd.n4115 9.3005
R10709 gnd.n4117 gnd.n4116 9.3005
R10710 gnd.n2214 gnd.n2211 9.3005
R10711 gnd.n4139 gnd.n2212 9.3005
R10712 gnd.n4138 gnd.n4135 9.3005
R10713 gnd.n4137 gnd.n4136 9.3005
R10714 gnd.n2196 gnd.n2193 9.3005
R10715 gnd.n4160 gnd.n2194 9.3005
R10716 gnd.n4159 gnd.n4156 9.3005
R10717 gnd.n4158 gnd.n4157 9.3005
R10718 gnd.n2180 gnd.n2175 9.3005
R10719 gnd.n4187 gnd.n2176 9.3005
R10720 gnd.n4186 gnd.n2177 9.3005
R10721 gnd.n4185 gnd.n2178 9.3005
R10722 gnd.n4184 gnd.n4180 9.3005
R10723 gnd.n4182 gnd.n4181 9.3005
R10724 gnd.n2159 gnd.n1067 9.3005
R10725 gnd.n6004 gnd.n1068 9.3005
R10726 gnd.n6003 gnd.n1069 9.3005
R10727 gnd.n6002 gnd.n1070 9.3005
R10728 gnd.n4212 gnd.n1071 9.3005
R10729 gnd.n5992 gnd.n1089 9.3005
R10730 gnd.n5991 gnd.n1090 9.3005
R10731 gnd.n5990 gnd.n1091 9.3005
R10732 gnd.n2144 gnd.n1092 9.3005
R10733 gnd.n5980 gnd.n1108 9.3005
R10734 gnd.n5979 gnd.n1109 9.3005
R10735 gnd.n5978 gnd.n1110 9.3005
R10736 gnd.n4266 gnd.n1111 9.3005
R10737 gnd.n5968 gnd.n1129 9.3005
R10738 gnd.n5967 gnd.n1130 9.3005
R10739 gnd.n5966 gnd.n1131 9.3005
R10740 gnd.n4524 gnd.n1132 9.3005
R10741 gnd.n2267 gnd.n2265 9.3005
R10742 gnd.n4078 gnd.n4077 9.3005
R10743 gnd.n4076 gnd.n2270 9.3005
R10744 gnd.n2269 gnd.n2249 9.3005
R10745 gnd.n4092 gnd.n2250 9.3005
R10746 gnd.n4093 gnd.n2248 9.3005
R10747 gnd.n4095 gnd.n4094 9.3005
R10748 gnd.n4096 gnd.n2231 9.3005
R10749 gnd.n4112 gnd.n2232 9.3005
R10750 gnd.n4113 gnd.n2230 9.3005
R10751 gnd.n4115 gnd.n4114 9.3005
R10752 gnd.n4116 gnd.n2213 9.3005
R10753 gnd.n4132 gnd.n2214 9.3005
R10754 gnd.n4133 gnd.n2212 9.3005
R10755 gnd.n4135 gnd.n4134 9.3005
R10756 gnd.n4136 gnd.n2195 9.3005
R10757 gnd.n4153 gnd.n2196 9.3005
R10758 gnd.n4154 gnd.n2194 9.3005
R10759 gnd.n4156 gnd.n4155 9.3005
R10760 gnd.n4157 gnd.n2179 9.3005
R10761 gnd.n4173 gnd.n2180 9.3005
R10762 gnd.n4174 gnd.n2176 9.3005
R10763 gnd.n4176 gnd.n2177 9.3005
R10764 gnd.n4177 gnd.n2178 9.3005
R10765 gnd.n4180 gnd.n4179 9.3005
R10766 gnd.n4181 gnd.n2158 9.3005
R10767 gnd.n4208 gnd.n2159 9.3005
R10768 gnd.n4209 gnd.n1068 9.3005
R10769 gnd.n4210 gnd.n1069 9.3005
R10770 gnd.n4211 gnd.n1070 9.3005
R10771 gnd.n4215 gnd.n4212 9.3005
R10772 gnd.n4214 gnd.n1089 9.3005
R10773 gnd.n4213 gnd.n1090 9.3005
R10774 gnd.n2143 gnd.n1091 9.3005
R10775 gnd.n4262 gnd.n2144 9.3005
R10776 gnd.n4263 gnd.n1108 9.3005
R10777 gnd.n4264 gnd.n1109 9.3005
R10778 gnd.n4265 gnd.n1110 9.3005
R10779 gnd.n4269 gnd.n4266 9.3005
R10780 gnd.n4270 gnd.n1129 9.3005
R10781 gnd.n4527 gnd.n1130 9.3005
R10782 gnd.n4526 gnd.n1131 9.3005
R10783 gnd.n4525 gnd.n4524 9.3005
R10784 gnd.n4075 gnd.n2267 9.3005
R10785 gnd.n3956 gnd.n3955 9.3005
R10786 gnd.n3958 gnd.n3835 9.3005
R10787 gnd.n3959 gnd.n3834 9.3005
R10788 gnd.n3962 gnd.n3833 9.3005
R10789 gnd.n3963 gnd.n3832 9.3005
R10790 gnd.n3966 gnd.n3831 9.3005
R10791 gnd.n3967 gnd.n3830 9.3005
R10792 gnd.n3970 gnd.n3829 9.3005
R10793 gnd.n3971 gnd.n3828 9.3005
R10794 gnd.n3974 gnd.n3827 9.3005
R10795 gnd.n3975 gnd.n3826 9.3005
R10796 gnd.n3978 gnd.n3825 9.3005
R10797 gnd.n3979 gnd.n3824 9.3005
R10798 gnd.n3982 gnd.n3823 9.3005
R10799 gnd.n3983 gnd.n3822 9.3005
R10800 gnd.n3986 gnd.n3821 9.3005
R10801 gnd.n3987 gnd.n3820 9.3005
R10802 gnd.n3990 gnd.n3819 9.3005
R10803 gnd.n3991 gnd.n3818 9.3005
R10804 gnd.n3994 gnd.n3817 9.3005
R10805 gnd.n3998 gnd.n3813 9.3005
R10806 gnd.n3999 gnd.n3812 9.3005
R10807 gnd.n4002 gnd.n3811 9.3005
R10808 gnd.n4003 gnd.n3810 9.3005
R10809 gnd.n4006 gnd.n3809 9.3005
R10810 gnd.n4007 gnd.n3808 9.3005
R10811 gnd.n4010 gnd.n3807 9.3005
R10812 gnd.n4011 gnd.n3806 9.3005
R10813 gnd.n4014 gnd.n3805 9.3005
R10814 gnd.n4015 gnd.n3804 9.3005
R10815 gnd.n4018 gnd.n3803 9.3005
R10816 gnd.n4019 gnd.n3802 9.3005
R10817 gnd.n4022 gnd.n3801 9.3005
R10818 gnd.n4023 gnd.n3800 9.3005
R10819 gnd.n4026 gnd.n3799 9.3005
R10820 gnd.n4027 gnd.n3798 9.3005
R10821 gnd.n4030 gnd.n3797 9.3005
R10822 gnd.n4031 gnd.n3796 9.3005
R10823 gnd.n4034 gnd.n3795 9.3005
R10824 gnd.n4036 gnd.n3792 9.3005
R10825 gnd.n4039 gnd.n3791 9.3005
R10826 gnd.n4040 gnd.n3790 9.3005
R10827 gnd.n4043 gnd.n3789 9.3005
R10828 gnd.n4044 gnd.n3788 9.3005
R10829 gnd.n4047 gnd.n3787 9.3005
R10830 gnd.n4048 gnd.n3786 9.3005
R10831 gnd.n4051 gnd.n3785 9.3005
R10832 gnd.n4052 gnd.n3784 9.3005
R10833 gnd.n4055 gnd.n3783 9.3005
R10834 gnd.n4056 gnd.n3782 9.3005
R10835 gnd.n4059 gnd.n3781 9.3005
R10836 gnd.n4060 gnd.n3780 9.3005
R10837 gnd.n4063 gnd.n3779 9.3005
R10838 gnd.n4065 gnd.n3778 9.3005
R10839 gnd.n4066 gnd.n3777 9.3005
R10840 gnd.n4067 gnd.n3776 9.3005
R10841 gnd.n4068 gnd.n3775 9.3005
R10842 gnd.n3995 gnd.n3814 9.3005
R10843 gnd.n3954 gnd.n2271 9.3005
R10844 gnd.n4084 gnd.n4083 9.3005
R10845 gnd.n4085 gnd.n2256 9.3005
R10846 gnd.n4087 gnd.n4086 9.3005
R10847 gnd.n2239 gnd.n2238 9.3005
R10848 gnd.n4104 gnd.n4103 9.3005
R10849 gnd.n4105 gnd.n2237 9.3005
R10850 gnd.n4107 gnd.n4106 9.3005
R10851 gnd.n2222 gnd.n2221 9.3005
R10852 gnd.n4124 gnd.n4123 9.3005
R10853 gnd.n4125 gnd.n2220 9.3005
R10854 gnd.n4127 gnd.n4126 9.3005
R10855 gnd.n2203 gnd.n2202 9.3005
R10856 gnd.n4144 gnd.n4143 9.3005
R10857 gnd.n4145 gnd.n2201 9.3005
R10858 gnd.n4148 gnd.n4146 9.3005
R10859 gnd.n6008 gnd.n1059 9.3005
R10860 gnd.n1078 gnd.n1060 9.3005
R10861 gnd.n5998 gnd.n1079 9.3005
R10862 gnd.n5997 gnd.n1080 9.3005
R10863 gnd.n5996 gnd.n1081 9.3005
R10864 gnd.n1098 gnd.n1082 9.3005
R10865 gnd.n5986 gnd.n1099 9.3005
R10866 gnd.n5985 gnd.n1100 9.3005
R10867 gnd.n5984 gnd.n1101 9.3005
R10868 gnd.n1118 gnd.n1102 9.3005
R10869 gnd.n5974 gnd.n1119 9.3005
R10870 gnd.n5973 gnd.n1120 9.3005
R10871 gnd.n5972 gnd.n1121 9.3005
R10872 gnd.n1139 gnd.n1122 9.3005
R10873 gnd.n5962 gnd.n1140 9.3005
R10874 gnd.n5961 gnd.n5960 9.3005
R10875 gnd.n2258 gnd.n2257 9.3005
R10876 gnd.n6009 gnd.n1058 9.3005
R10877 gnd.n4231 gnd.n4230 9.3005
R10878 gnd.n6016 gnd.n1047 9.3005
R10879 gnd.n6017 gnd.n1046 9.3005
R10880 gnd.n1045 gnd.n1041 9.3005
R10881 gnd.n6023 gnd.n1040 9.3005
R10882 gnd.n6024 gnd.n1039 9.3005
R10883 gnd.n6025 gnd.n1038 9.3005
R10884 gnd.n1037 gnd.n1033 9.3005
R10885 gnd.n6031 gnd.n1032 9.3005
R10886 gnd.n6032 gnd.n1031 9.3005
R10887 gnd.n6033 gnd.n1030 9.3005
R10888 gnd.n1029 gnd.n1025 9.3005
R10889 gnd.n6039 gnd.n1024 9.3005
R10890 gnd.n6040 gnd.n1023 9.3005
R10891 gnd.n6041 gnd.n1022 9.3005
R10892 gnd.n1021 gnd.n1017 9.3005
R10893 gnd.n6047 gnd.n1016 9.3005
R10894 gnd.n6048 gnd.n1015 9.3005
R10895 gnd.n6049 gnd.n1014 9.3005
R10896 gnd.n1013 gnd.n1009 9.3005
R10897 gnd.n6055 gnd.n1008 9.3005
R10898 gnd.n6056 gnd.n1007 9.3005
R10899 gnd.n6057 gnd.n1006 9.3005
R10900 gnd.n1005 gnd.n1001 9.3005
R10901 gnd.n6063 gnd.n1000 9.3005
R10902 gnd.n6064 gnd.n999 9.3005
R10903 gnd.n6065 gnd.n998 9.3005
R10904 gnd.n997 gnd.n993 9.3005
R10905 gnd.n6071 gnd.n992 9.3005
R10906 gnd.n6072 gnd.n991 9.3005
R10907 gnd.n6073 gnd.n990 9.3005
R10908 gnd.n989 gnd.n985 9.3005
R10909 gnd.n6079 gnd.n984 9.3005
R10910 gnd.n6080 gnd.n983 9.3005
R10911 gnd.n6081 gnd.n982 9.3005
R10912 gnd.n981 gnd.n977 9.3005
R10913 gnd.n6087 gnd.n976 9.3005
R10914 gnd.n6088 gnd.n975 9.3005
R10915 gnd.n6089 gnd.n974 9.3005
R10916 gnd.n973 gnd.n969 9.3005
R10917 gnd.n6095 gnd.n968 9.3005
R10918 gnd.n6096 gnd.n967 9.3005
R10919 gnd.n6097 gnd.n966 9.3005
R10920 gnd.n965 gnd.n961 9.3005
R10921 gnd.n6103 gnd.n960 9.3005
R10922 gnd.n6104 gnd.n959 9.3005
R10923 gnd.n6105 gnd.n958 9.3005
R10924 gnd.n957 gnd.n953 9.3005
R10925 gnd.n6111 gnd.n952 9.3005
R10926 gnd.n6112 gnd.n951 9.3005
R10927 gnd.n6113 gnd.n950 9.3005
R10928 gnd.n949 gnd.n945 9.3005
R10929 gnd.n6119 gnd.n944 9.3005
R10930 gnd.n6120 gnd.n943 9.3005
R10931 gnd.n6121 gnd.n942 9.3005
R10932 gnd.n941 gnd.n937 9.3005
R10933 gnd.n6127 gnd.n936 9.3005
R10934 gnd.n6128 gnd.n935 9.3005
R10935 gnd.n6129 gnd.n934 9.3005
R10936 gnd.n933 gnd.n929 9.3005
R10937 gnd.n6135 gnd.n928 9.3005
R10938 gnd.n6136 gnd.n927 9.3005
R10939 gnd.n6137 gnd.n926 9.3005
R10940 gnd.n925 gnd.n921 9.3005
R10941 gnd.n6143 gnd.n920 9.3005
R10942 gnd.n6144 gnd.n919 9.3005
R10943 gnd.n6145 gnd.n918 9.3005
R10944 gnd.n917 gnd.n913 9.3005
R10945 gnd.n6151 gnd.n912 9.3005
R10946 gnd.n6152 gnd.n911 9.3005
R10947 gnd.n6153 gnd.n910 9.3005
R10948 gnd.n909 gnd.n905 9.3005
R10949 gnd.n6159 gnd.n904 9.3005
R10950 gnd.n6160 gnd.n903 9.3005
R10951 gnd.n6161 gnd.n902 9.3005
R10952 gnd.n901 gnd.n897 9.3005
R10953 gnd.n6167 gnd.n896 9.3005
R10954 gnd.n6168 gnd.n895 9.3005
R10955 gnd.n6169 gnd.n894 9.3005
R10956 gnd.n893 gnd.n889 9.3005
R10957 gnd.n6175 gnd.n888 9.3005
R10958 gnd.n6176 gnd.n887 9.3005
R10959 gnd.n6177 gnd.n886 9.3005
R10960 gnd.n882 gnd.n881 9.3005
R10961 gnd.n6184 gnd.n6183 9.3005
R10962 gnd.n6015 gnd.n1048 9.3005
R10963 gnd.n5429 gnd.n1375 9.3005
R10964 gnd.n4591 gnd.n4590 9.3005
R10965 gnd.n4592 gnd.n2092 9.3005
R10966 gnd.n4594 gnd.n4593 9.3005
R10967 gnd.n2079 gnd.n2078 9.3005
R10968 gnd.n4607 gnd.n4606 9.3005
R10969 gnd.n4608 gnd.n2076 9.3005
R10970 gnd.n4627 gnd.n4626 9.3005
R10971 gnd.n4625 gnd.n2077 9.3005
R10972 gnd.n4624 gnd.n4623 9.3005
R10973 gnd.n4622 gnd.n4609 9.3005
R10974 gnd.n4621 gnd.n4620 9.3005
R10975 gnd.n4619 gnd.n4612 9.3005
R10976 gnd.n4618 gnd.n4617 9.3005
R10977 gnd.n4616 gnd.n4613 9.3005
R10978 gnd.n1294 gnd.n1292 9.3005
R10979 gnd.n5823 gnd.n5822 9.3005
R10980 gnd.n5821 gnd.n1293 9.3005
R10981 gnd.n5820 gnd.n5819 9.3005
R10982 gnd.n5818 gnd.n1295 9.3005
R10983 gnd.n5817 gnd.n5816 9.3005
R10984 gnd.n5815 gnd.n1299 9.3005
R10985 gnd.n5814 gnd.n5813 9.3005
R10986 gnd.n5812 gnd.n1300 9.3005
R10987 gnd.n5811 gnd.n5810 9.3005
R10988 gnd.n5809 gnd.n1304 9.3005
R10989 gnd.n5808 gnd.n5807 9.3005
R10990 gnd.n5806 gnd.n1305 9.3005
R10991 gnd.n5805 gnd.n5804 9.3005
R10992 gnd.n5803 gnd.n1309 9.3005
R10993 gnd.n5802 gnd.n5801 9.3005
R10994 gnd.n5800 gnd.n1310 9.3005
R10995 gnd.n5799 gnd.n5798 9.3005
R10996 gnd.n5797 gnd.n1314 9.3005
R10997 gnd.n5796 gnd.n5795 9.3005
R10998 gnd.n5794 gnd.n1315 9.3005
R10999 gnd.n5793 gnd.n5792 9.3005
R11000 gnd.n5791 gnd.n1319 9.3005
R11001 gnd.n5790 gnd.n5789 9.3005
R11002 gnd.n5788 gnd.n1320 9.3005
R11003 gnd.n5787 gnd.n5786 9.3005
R11004 gnd.n5785 gnd.n1324 9.3005
R11005 gnd.n5784 gnd.n5783 9.3005
R11006 gnd.n5782 gnd.n1325 9.3005
R11007 gnd.n5781 gnd.n5780 9.3005
R11008 gnd.n5779 gnd.n1329 9.3005
R11009 gnd.n5778 gnd.n5777 9.3005
R11010 gnd.n5776 gnd.n1330 9.3005
R11011 gnd.n5775 gnd.n5774 9.3005
R11012 gnd.n5773 gnd.n1334 9.3005
R11013 gnd.n5772 gnd.n5771 9.3005
R11014 gnd.n5770 gnd.n1335 9.3005
R11015 gnd.n5769 gnd.n5768 9.3005
R11016 gnd.n5767 gnd.n1339 9.3005
R11017 gnd.n5766 gnd.n5765 9.3005
R11018 gnd.n5764 gnd.n1340 9.3005
R11019 gnd.n5763 gnd.n5762 9.3005
R11020 gnd.n5761 gnd.n1344 9.3005
R11021 gnd.n5760 gnd.n5759 9.3005
R11022 gnd.n5758 gnd.n1345 9.3005
R11023 gnd.n5757 gnd.n5756 9.3005
R11024 gnd.n5755 gnd.n1349 9.3005
R11025 gnd.n5754 gnd.n5753 9.3005
R11026 gnd.n5752 gnd.n1350 9.3005
R11027 gnd.n5751 gnd.n5750 9.3005
R11028 gnd.n5749 gnd.n1354 9.3005
R11029 gnd.n5748 gnd.n5747 9.3005
R11030 gnd.n5746 gnd.n1355 9.3005
R11031 gnd.n5745 gnd.n5744 9.3005
R11032 gnd.n5743 gnd.n1359 9.3005
R11033 gnd.n5742 gnd.n5741 9.3005
R11034 gnd.n5740 gnd.n1360 9.3005
R11035 gnd.n5739 gnd.n5738 9.3005
R11036 gnd.n5737 gnd.n1364 9.3005
R11037 gnd.n5736 gnd.n5735 9.3005
R11038 gnd.n5734 gnd.n1365 9.3005
R11039 gnd.n5733 gnd.n5732 9.3005
R11040 gnd.n5731 gnd.n1369 9.3005
R11041 gnd.n5730 gnd.n5729 9.3005
R11042 gnd.n5728 gnd.n1370 9.3005
R11043 gnd.n5727 gnd.n5726 9.3005
R11044 gnd.n5725 gnd.n1374 9.3005
R11045 gnd.n5724 gnd.n5723 9.3005
R11046 gnd.n2094 gnd.n2093 9.3005
R11047 gnd.n4577 gnd.n4576 9.3005
R11048 gnd.n3878 gnd.n3877 9.3005
R11049 gnd.n2162 gnd.n2161 9.3005
R11050 gnd.n4201 gnd.n4200 9.3005
R11051 gnd.n4202 gnd.n2160 9.3005
R11052 gnd.n4204 gnd.n4203 9.3005
R11053 gnd.n2157 gnd.n2155 9.3005
R11054 gnd.n4223 gnd.n4222 9.3005
R11055 gnd.n4221 gnd.n2156 9.3005
R11056 gnd.n4220 gnd.n4219 9.3005
R11057 gnd.n2147 gnd.n2146 9.3005
R11058 gnd.n4255 gnd.n4254 9.3005
R11059 gnd.n4256 gnd.n2145 9.3005
R11060 gnd.n4258 gnd.n4257 9.3005
R11061 gnd.n2140 gnd.n2138 9.3005
R11062 gnd.n4540 gnd.n4539 9.3005
R11063 gnd.n4538 gnd.n2139 9.3005
R11064 gnd.n4537 gnd.n4536 9.3005
R11065 gnd.n4535 gnd.n2141 9.3005
R11066 gnd.n4534 gnd.n4533 9.3005
R11067 gnd.n4532 gnd.n4531 9.3005
R11068 gnd.n2125 gnd.n2120 9.3005
R11069 gnd.n4418 gnd.n4417 9.3005
R11070 gnd.n4317 gnd.n4316 9.3005
R11071 gnd.n4412 gnd.n4411 9.3005
R11072 gnd.n4410 gnd.n4409 9.3005
R11073 gnd.n4329 gnd.n4328 9.3005
R11074 gnd.n4404 gnd.n4403 9.3005
R11075 gnd.n4402 gnd.n4401 9.3005
R11076 gnd.n4337 gnd.n4336 9.3005
R11077 gnd.n4396 gnd.n4395 9.3005
R11078 gnd.n4394 gnd.n4393 9.3005
R11079 gnd.n4349 gnd.n4348 9.3005
R11080 gnd.n4388 gnd.n4387 9.3005
R11081 gnd.n4386 gnd.n4385 9.3005
R11082 gnd.n4357 gnd.n4356 9.3005
R11083 gnd.n4380 gnd.n4379 9.3005
R11084 gnd.n4378 gnd.n4377 9.3005
R11085 gnd.n4368 gnd.n2124 9.3005
R11086 gnd.n4573 gnd.n4572 9.3005
R11087 gnd.n4420 gnd.n4419 9.3005
R11088 gnd.n4574 gnd.n2119 9.3005
R11089 gnd.n4374 gnd.n2121 9.3005
R11090 gnd.n4376 gnd.n4375 9.3005
R11091 gnd.n4363 gnd.n4362 9.3005
R11092 gnd.n4382 gnd.n4381 9.3005
R11093 gnd.n4384 gnd.n4383 9.3005
R11094 gnd.n4353 gnd.n4352 9.3005
R11095 gnd.n4390 gnd.n4389 9.3005
R11096 gnd.n4392 gnd.n4391 9.3005
R11097 gnd.n4343 gnd.n4342 9.3005
R11098 gnd.n4398 gnd.n4397 9.3005
R11099 gnd.n4400 gnd.n4399 9.3005
R11100 gnd.n4333 gnd.n4332 9.3005
R11101 gnd.n4406 gnd.n4405 9.3005
R11102 gnd.n4408 gnd.n4407 9.3005
R11103 gnd.n4323 gnd.n4322 9.3005
R11104 gnd.n4414 gnd.n4413 9.3005
R11105 gnd.n4416 gnd.n4415 9.3005
R11106 gnd.n4314 gnd.n4313 9.3005
R11107 gnd.n4422 gnd.n4421 9.3005
R11108 gnd.n4423 gnd.n4271 9.3005
R11109 gnd.n4425 gnd.n4424 9.3005
R11110 gnd.n4308 gnd.n4272 9.3005
R11111 gnd.n4307 gnd.n4306 9.3005
R11112 gnd.n4305 gnd.n4273 9.3005
R11113 gnd.n4304 gnd.n4303 9.3005
R11114 gnd.n4300 gnd.n4276 9.3005
R11115 gnd.n4299 gnd.n4277 9.3005
R11116 gnd.n4294 gnd.n4278 9.3005
R11117 gnd.n4293 gnd.n4292 9.3005
R11118 gnd.n4291 gnd.n4279 9.3005
R11119 gnd.n4290 gnd.n4289 9.3005
R11120 gnd.n4288 gnd.n4282 9.3005
R11121 gnd.n4287 gnd.n4286 9.3005
R11122 gnd.n4285 gnd.n4283 9.3005
R11123 gnd.n2062 gnd.n2061 9.3005
R11124 gnd.n4649 gnd.n4648 9.3005
R11125 gnd.n4650 gnd.n2060 9.3005
R11126 gnd.n4652 gnd.n4651 9.3005
R11127 gnd.n2058 gnd.n2057 9.3005
R11128 gnd.n4657 gnd.n4656 9.3005
R11129 gnd.n4658 gnd.n2055 9.3005
R11130 gnd.n4669 gnd.n4668 9.3005
R11131 gnd.n4667 gnd.n2056 9.3005
R11132 gnd.n4666 gnd.n4665 9.3005
R11133 gnd.n4664 gnd.n4659 9.3005
R11134 gnd.n4663 gnd.n4662 9.3005
R11135 gnd.n2024 gnd.n2023 9.3005
R11136 gnd.n4809 gnd.n4808 9.3005
R11137 gnd.n4810 gnd.n2021 9.3005
R11138 gnd.n4815 gnd.n4814 9.3005
R11139 gnd.n4813 gnd.n2022 9.3005
R11140 gnd.n4812 gnd.n4811 9.3005
R11141 gnd.n2003 gnd.n2002 9.3005
R11142 gnd.n4840 gnd.n4839 9.3005
R11143 gnd.n4841 gnd.n2000 9.3005
R11144 gnd.n4849 gnd.n4848 9.3005
R11145 gnd.n4847 gnd.n2001 9.3005
R11146 gnd.n4846 gnd.n4845 9.3005
R11147 gnd.n4844 gnd.n4842 9.3005
R11148 gnd.n1953 gnd.n1952 9.3005
R11149 gnd.n4920 gnd.n4919 9.3005
R11150 gnd.n4921 gnd.n1950 9.3005
R11151 gnd.n4924 gnd.n4923 9.3005
R11152 gnd.n4922 gnd.n1951 9.3005
R11153 gnd.n1926 gnd.n1925 9.3005
R11154 gnd.n4966 gnd.n4965 9.3005
R11155 gnd.n4967 gnd.n1923 9.3005
R11156 gnd.n4995 gnd.n4994 9.3005
R11157 gnd.n4993 gnd.n1924 9.3005
R11158 gnd.n4992 gnd.n4991 9.3005
R11159 gnd.n4990 gnd.n4968 9.3005
R11160 gnd.n4989 gnd.n4988 9.3005
R11161 gnd.n4987 gnd.n4973 9.3005
R11162 gnd.n4986 gnd.n4985 9.3005
R11163 gnd.n4984 gnd.n4974 9.3005
R11164 gnd.n4983 gnd.n4982 9.3005
R11165 gnd.n4981 gnd.n4978 9.3005
R11166 gnd.n4980 gnd.n4979 9.3005
R11167 gnd.n1851 gnd.n1850 9.3005
R11168 gnd.n5099 gnd.n5098 9.3005
R11169 gnd.n5100 gnd.n1848 9.3005
R11170 gnd.n5135 gnd.n5134 9.3005
R11171 gnd.n5133 gnd.n1849 9.3005
R11172 gnd.n5132 gnd.n5131 9.3005
R11173 gnd.n5130 gnd.n5101 9.3005
R11174 gnd.n5129 gnd.n5128 9.3005
R11175 gnd.n5127 gnd.n5106 9.3005
R11176 gnd.n5126 gnd.n5125 9.3005
R11177 gnd.n5124 gnd.n5107 9.3005
R11178 gnd.n5123 gnd.n5122 9.3005
R11179 gnd.n5121 gnd.n5110 9.3005
R11180 gnd.n5120 gnd.n5119 9.3005
R11181 gnd.n5118 gnd.n5111 9.3005
R11182 gnd.n5117 gnd.n5116 9.3005
R11183 gnd.n5115 gnd.n5114 9.3005
R11184 gnd.n1698 gnd.n1697 9.3005
R11185 gnd.n5362 gnd.n5361 9.3005
R11186 gnd.n5363 gnd.n1696 9.3005
R11187 gnd.n5365 gnd.n5364 9.3005
R11188 gnd.n1685 gnd.n1684 9.3005
R11189 gnd.n5378 gnd.n5377 9.3005
R11190 gnd.n5379 gnd.n1683 9.3005
R11191 gnd.n5381 gnd.n5380 9.3005
R11192 gnd.n1673 gnd.n1672 9.3005
R11193 gnd.n5397 gnd.n5396 9.3005
R11194 gnd.n5398 gnd.n1671 9.3005
R11195 gnd.n5400 gnd.n5399 9.3005
R11196 gnd.n1384 gnd.n1383 9.3005
R11197 gnd.n5719 gnd.n5718 9.3005
R11198 gnd.n4296 gnd.n4295 9.3005
R11199 gnd.n5715 gnd.n1385 9.3005
R11200 gnd.n5714 gnd.n5713 9.3005
R11201 gnd.n5712 gnd.n1388 9.3005
R11202 gnd.n5711 gnd.n5710 9.3005
R11203 gnd.n5709 gnd.n1389 9.3005
R11204 gnd.n5708 gnd.n5707 9.3005
R11205 gnd.n5717 gnd.n5716 9.3005
R11206 gnd.n5660 gnd.n5659 9.3005
R11207 gnd.n1436 gnd.n1435 9.3005
R11208 gnd.n5666 gnd.n5665 9.3005
R11209 gnd.n5668 gnd.n5667 9.3005
R11210 gnd.n1428 gnd.n1427 9.3005
R11211 gnd.n5674 gnd.n5673 9.3005
R11212 gnd.n5676 gnd.n5675 9.3005
R11213 gnd.n1420 gnd.n1419 9.3005
R11214 gnd.n5682 gnd.n5681 9.3005
R11215 gnd.n5684 gnd.n5683 9.3005
R11216 gnd.n1412 gnd.n1411 9.3005
R11217 gnd.n5690 gnd.n5689 9.3005
R11218 gnd.n5692 gnd.n5691 9.3005
R11219 gnd.n1404 gnd.n1403 9.3005
R11220 gnd.n5698 gnd.n5697 9.3005
R11221 gnd.n5700 gnd.n5699 9.3005
R11222 gnd.n1400 gnd.n1395 9.3005
R11223 gnd.n5658 gnd.n1445 9.3005
R11224 gnd.n1636 gnd.n1444 9.3005
R11225 gnd.n5705 gnd.n1393 9.3005
R11226 gnd.n5704 gnd.n5703 9.3005
R11227 gnd.n5702 gnd.n5701 9.3005
R11228 gnd.n1399 gnd.n1398 9.3005
R11229 gnd.n5696 gnd.n5695 9.3005
R11230 gnd.n5694 gnd.n5693 9.3005
R11231 gnd.n1408 gnd.n1407 9.3005
R11232 gnd.n5688 gnd.n5687 9.3005
R11233 gnd.n5686 gnd.n5685 9.3005
R11234 gnd.n1416 gnd.n1415 9.3005
R11235 gnd.n5680 gnd.n5679 9.3005
R11236 gnd.n5678 gnd.n5677 9.3005
R11237 gnd.n1424 gnd.n1423 9.3005
R11238 gnd.n5672 gnd.n5671 9.3005
R11239 gnd.n5670 gnd.n5669 9.3005
R11240 gnd.n1432 gnd.n1431 9.3005
R11241 gnd.n5664 gnd.n5663 9.3005
R11242 gnd.n5662 gnd.n5661 9.3005
R11243 gnd.n1659 gnd.n1442 9.3005
R11244 gnd.n1638 gnd.n1637 9.3005
R11245 gnd.n5431 gnd.n5430 9.3005
R11246 gnd.n5468 gnd.n5467 9.3005
R11247 gnd.n5466 gnd.n1635 9.3005
R11248 gnd.n5465 gnd.n5464 9.3005
R11249 gnd.n5463 gnd.n5434 9.3005
R11250 gnd.n5462 gnd.n5461 9.3005
R11251 gnd.n5460 gnd.n5438 9.3005
R11252 gnd.n5459 gnd.n5458 9.3005
R11253 gnd.n5457 gnd.n5439 9.3005
R11254 gnd.n5456 gnd.n5455 9.3005
R11255 gnd.n5454 gnd.n5451 9.3005
R11256 gnd.n5453 gnd.n5452 9.3005
R11257 gnd.n534 gnd.n533 9.3005
R11258 gnd.n6750 gnd.n6749 9.3005
R11259 gnd.n6751 gnd.n532 9.3005
R11260 gnd.n6753 gnd.n6752 9.3005
R11261 gnd.n515 gnd.n514 9.3005
R11262 gnd.n6777 gnd.n6776 9.3005
R11263 gnd.n6778 gnd.n512 9.3005
R11264 gnd.n6780 gnd.n6779 9.3005
R11265 gnd.n513 gnd.n63 9.3005
R11266 gnd.n5433 gnd.n1634 9.3005
R11267 gnd.n6902 gnd.n64 9.3005
R11268 gnd.t25 gnd.n2463 9.24152
R11269 gnd.n2365 gnd.t311 9.24152
R11270 gnd.n3634 gnd.t295 9.24152
R11271 gnd.t188 gnd.t25 8.92286
R11272 gnd.n3604 gnd.n3579 8.92171
R11273 gnd.n3572 gnd.n3547 8.92171
R11274 gnd.n3540 gnd.n3515 8.92171
R11275 gnd.n3509 gnd.n3484 8.92171
R11276 gnd.n3477 gnd.n3452 8.92171
R11277 gnd.n3445 gnd.n3420 8.92171
R11278 gnd.n3413 gnd.n3388 8.92171
R11279 gnd.n3382 gnd.n3357 8.92171
R11280 gnd.n1734 gnd.n1716 8.72777
R11281 gnd.n3107 gnd.t2 8.60421
R11282 gnd.n2527 gnd.n2515 8.43656
R11283 gnd.n38 gnd.n26 8.43656
R11284 gnd.n4867 gnd.n1988 8.28555
R11285 gnd.n4953 gnd.n4951 8.28555
R11286 gnd.n5023 gnd.n1901 8.28555
R11287 gnd.n5077 gnd.n1845 8.28555
R11288 gnd.n3605 gnd.n3577 8.14595
R11289 gnd.n3573 gnd.n3545 8.14595
R11290 gnd.n3541 gnd.n3513 8.14595
R11291 gnd.n3510 gnd.n3482 8.14595
R11292 gnd.n3478 gnd.n3450 8.14595
R11293 gnd.n3446 gnd.n3418 8.14595
R11294 gnd.n3414 gnd.n3386 8.14595
R11295 gnd.n3383 gnd.n3355 8.14595
R11296 gnd.n3879 gnd.n0 8.10675
R11297 gnd.n6903 gnd.n6902 8.10675
R11298 gnd.n3610 gnd.n3609 7.97301
R11299 gnd.t67 gnd.n2622 7.9669
R11300 gnd.n6903 gnd.n62 7.78567
R11301 gnd.n5658 gnd.n1444 7.75808
R11302 gnd.n4572 gnd.n2124 7.75808
R11303 gnd.n250 gnd.n199 7.75808
R11304 gnd.n3914 gnd.n3856 7.75808
R11305 gnd.n3348 gnd.n2362 7.64824
R11306 gnd.t0 gnd.n4898 7.64824
R11307 gnd.n4927 gnd.t22 7.64824
R11308 gnd.t38 gnd.n1899 7.64824
R11309 gnd.n5042 gnd.t18 7.64824
R11310 gnd.n5213 gnd.t230 7.64824
R11311 gnd.n2552 gnd.n2551 7.53171
R11312 gnd.n3016 gnd.t60 7.32958
R11313 gnd.n1272 gnd.n1271 7.30353
R11314 gnd.n1733 gnd.n1732 7.30353
R11315 gnd.n2976 gnd.n2695 7.01093
R11316 gnd.n2698 gnd.n2696 7.01093
R11317 gnd.n2986 gnd.n2985 7.01093
R11318 gnd.n2997 gnd.n2679 7.01093
R11319 gnd.n2996 gnd.n2682 7.01093
R11320 gnd.n3007 gnd.n2670 7.01093
R11321 gnd.n2673 gnd.n2671 7.01093
R11322 gnd.n3017 gnd.n3016 7.01093
R11323 gnd.n3027 gnd.n2651 7.01093
R11324 gnd.n3026 gnd.n2654 7.01093
R11325 gnd.n3035 gnd.n2645 7.01093
R11326 gnd.n3047 gnd.n2635 7.01093
R11327 gnd.n3057 gnd.n2620 7.01093
R11328 gnd.n3073 gnd.n3072 7.01093
R11329 gnd.n2622 gnd.n2559 7.01093
R11330 gnd.n3127 gnd.n2560 7.01093
R11331 gnd.n3121 gnd.n3120 7.01093
R11332 gnd.n2609 gnd.n2571 7.01093
R11333 gnd.n3113 gnd.n2582 7.01093
R11334 gnd.n2600 gnd.n2595 7.01093
R11335 gnd.n3107 gnd.n3106 7.01093
R11336 gnd.n3153 gnd.n2498 7.01093
R11337 gnd.n3152 gnd.n3151 7.01093
R11338 gnd.n3164 gnd.n3163 7.01093
R11339 gnd.n2491 gnd.n2483 7.01093
R11340 gnd.n3193 gnd.n2471 7.01093
R11341 gnd.n3192 gnd.n2474 7.01093
R11342 gnd.n3203 gnd.n2463 7.01093
R11343 gnd.n2464 gnd.n2452 7.01093
R11344 gnd.n3214 gnd.n2453 7.01093
R11345 gnd.n3238 gnd.n2444 7.01093
R11346 gnd.n3237 gnd.n2435 7.01093
R11347 gnd.n3260 gnd.n3259 7.01093
R11348 gnd.n3278 gnd.n2416 7.01093
R11349 gnd.n3277 gnd.n2419 7.01093
R11350 gnd.n3288 gnd.n2408 7.01093
R11351 gnd.n2409 gnd.n2396 7.01093
R11352 gnd.n3299 gnd.n2397 7.01093
R11353 gnd.n3326 gnd.n2381 7.01093
R11354 gnd.n3338 gnd.n3337 7.01093
R11355 gnd.n3320 gnd.n2374 7.01093
R11356 gnd.n3350 gnd.n3349 7.01093
R11357 gnd.n3622 gnd.n2362 7.01093
R11358 gnd.n3621 gnd.n2365 7.01093
R11359 gnd.n3634 gnd.n2354 7.01093
R11360 gnd.n2355 gnd.n2347 7.01093
R11361 gnd.n3644 gnd.n2273 7.01093
R11362 gnd.n4739 gnd.n1276 7.01093
R11363 gnd.n4784 gnd.n2044 7.01093
R11364 gnd.n4796 gnd.t205 7.01093
R11365 gnd.n4876 gnd.n4875 7.01093
R11366 gnd.n4899 gnd.t0 7.01093
R11367 gnd.n4898 gnd.n4897 7.01093
R11368 gnd.n5042 gnd.n1887 7.01093
R11369 gnd.t18 gnd.n5041 7.01093
R11370 gnd.n5062 gnd.n1864 7.01093
R11371 gnd.n1712 gnd.n1700 7.01093
R11372 gnd.n2654 gnd.t4 6.69227
R11373 gnd.n2474 gnd.t188 6.69227
R11374 gnd.n3327 gnd.t58 6.69227
R11375 gnd.n4543 gnd.t83 6.69227
R11376 gnd.t43 gnd.n2039 6.69227
R11377 gnd.n5183 gnd.t200 6.69227
R11378 gnd.t90 gnd.n1597 6.69227
R11379 gnd.n5279 gnd.n5278 6.5566
R11380 gnd.n4680 gnd.n4679 6.5566
R11381 gnd.n5843 gnd.n5839 6.5566
R11382 gnd.n5294 gnd.n5293 6.5566
R11383 gnd.n4739 gnd.t212 6.37362
R11384 gnd.n4906 gnd.t33 6.37362
R11385 gnd.t12 gnd.n1880 6.37362
R11386 gnd.n4375 gnd.n4371 6.20656
R11387 gnd.n1659 gnd.n1441 6.20656
R11388 gnd.t198 gnd.n3083 6.05496
R11389 gnd.n3084 gnd.t27 6.05496
R11390 gnd.t49 gnd.n2498 6.05496
R11391 gnd.t26 gnd.n3248 6.05496
R11392 gnd.n4226 gnd.t77 6.05496
R11393 gnd.t196 gnd.t6 6.05496
R11394 gnd.t19 gnd.t13 6.05496
R11395 gnd.n6728 gnd.t100 6.05496
R11396 gnd.n3607 gnd.n3577 5.81868
R11397 gnd.n3575 gnd.n3545 5.81868
R11398 gnd.n3543 gnd.n3513 5.81868
R11399 gnd.n3512 gnd.n3482 5.81868
R11400 gnd.n3480 gnd.n3450 5.81868
R11401 gnd.n3448 gnd.n3418 5.81868
R11402 gnd.n3416 gnd.n3386 5.81868
R11403 gnd.n3385 gnd.n3355 5.81868
R11404 gnd.n4672 gnd.n4671 5.73631
R11405 gnd.n1982 gnd.t32 5.73631
R11406 gnd.n4907 gnd.n1962 5.73631
R11407 gnd.n4890 gnd.n4889 5.73631
R11408 gnd.n4953 gnd.t22 5.73631
R11409 gnd.n1901 gnd.t38 5.73631
R11410 gnd.n5051 gnd.n5050 5.73631
R11411 gnd.n5057 gnd.n1873 5.73631
R11412 gnd.t36 gnd.n5085 5.73631
R11413 gnd.n5219 gnd.n1787 5.73631
R11414 gnd.n1760 gnd.n1521 5.62001
R11415 gnd.n5905 gnd.n1214 5.62001
R11416 gnd.n5905 gnd.n1215 5.62001
R11417 gnd.n5288 gnd.n1521 5.62001
R11418 gnd.n2835 gnd.n2830 5.4308
R11419 gnd.n3652 gnd.n2340 5.4308
R11420 gnd.n3151 gnd.t28 5.41765
R11421 gnd.t24 gnd.n3174 5.41765
R11422 gnd.t56 gnd.n2428 5.41765
R11423 gnd.n4765 gnd.t47 5.41765
R11424 gnd.n5103 gnd.t202 5.41765
R11425 gnd.n4206 gnd.n1053 5.09899
R11426 gnd.n6006 gnd.n1062 5.09899
R11427 gnd.n4226 gnd.n4225 5.09899
R11428 gnd.n6000 gnd.n1073 5.09899
R11429 gnd.n4217 gnd.n1076 5.09899
R11430 gnd.n5994 gnd.n1084 5.09899
R11431 gnd.n4252 gnd.n1087 5.09899
R11432 gnd.n4260 gnd.n1096 5.09899
R11433 gnd.n5982 gnd.n1104 5.09899
R11434 gnd.n4543 gnd.n4542 5.09899
R11435 gnd.n5976 gnd.n1113 5.09899
R11436 gnd.n4267 gnd.n1116 5.09899
R11437 gnd.n5970 gnd.n1124 5.09899
R11438 gnd.n4529 gnd.n1127 5.09899
R11439 gnd.n5964 gnd.n1134 5.09899
R11440 gnd.n4569 gnd.n1137 5.09899
R11441 gnd.n4866 gnd.t5 5.09899
R11442 gnd.n5078 gnd.t20 5.09899
R11443 gnd.n5532 gnd.n1559 5.09899
R11444 gnd.n5471 gnd.n5470 5.09899
R11445 gnd.n5524 gnd.n1568 5.09899
R11446 gnd.n5435 gnd.n1581 5.09899
R11447 gnd.n5518 gnd.n1584 5.09899
R11448 gnd.n5441 gnd.n1594 5.09899
R11449 gnd.n5512 gnd.n1597 5.09899
R11450 gnd.n5448 gnd.n1606 5.09899
R11451 gnd.n5506 gnd.n1609 5.09899
R11452 gnd.n1622 gnd.n546 5.09899
R11453 gnd.n6736 gnd.n549 5.09899
R11454 gnd.n1615 gnd.n536 5.09899
R11455 gnd.n6747 gnd.n538 5.09899
R11456 gnd.n6729 gnd.n6728 5.09899
R11457 gnd.n6755 gnd.n522 5.09899
R11458 gnd.n6769 gnd.n517 5.09899
R11459 gnd.n3605 gnd.n3604 5.04292
R11460 gnd.n3573 gnd.n3572 5.04292
R11461 gnd.n3541 gnd.n3540 5.04292
R11462 gnd.n3510 gnd.n3509 5.04292
R11463 gnd.n3478 gnd.n3477 5.04292
R11464 gnd.n3446 gnd.n3445 5.04292
R11465 gnd.n3414 gnd.n3413 5.04292
R11466 gnd.n3383 gnd.n3382 5.04292
R11467 gnd.n3114 gnd.t9 4.78034
R11468 gnd.n2453 gnd.t8 4.78034
R11469 gnd.n1702 gnd.t277 4.78034
R11470 gnd.n2556 gnd.n2553 4.74817
R11471 gnd.n2606 gnd.n2504 4.74817
R11472 gnd.n2593 gnd.n2503 4.74817
R11473 gnd.n2502 gnd.n2501 4.74817
R11474 gnd.n2602 gnd.n2553 4.74817
R11475 gnd.n2603 gnd.n2504 4.74817
R11476 gnd.n2605 gnd.n2503 4.74817
R11477 gnd.n2592 gnd.n2502 4.74817
R11478 gnd.n6772 gnd.n81 4.74817
R11479 gnd.n6787 gnd.n80 4.74817
R11480 gnd.n6785 gnd.n79 4.74817
R11481 gnd.n6895 gnd.n74 4.74817
R11482 gnd.n6893 gnd.n75 4.74817
R11483 gnd.n521 gnd.n81 4.74817
R11484 gnd.n6771 gnd.n80 4.74817
R11485 gnd.n6788 gnd.n79 4.74817
R11486 gnd.n6784 gnd.n74 4.74817
R11487 gnd.n6894 gnd.n6893 4.74817
R11488 gnd.n4164 gnd.n2186 4.74817
R11489 gnd.n4168 gnd.n4166 4.74817
R11490 gnd.n4191 gnd.n2167 4.74817
R11491 gnd.n4195 gnd.n4193 4.74817
R11492 gnd.n6010 gnd.n1057 4.74817
R11493 gnd.n4147 gnd.n2186 4.74817
R11494 gnd.n4166 gnd.n4165 4.74817
R11495 gnd.n4167 gnd.n2167 4.74817
R11496 gnd.n4193 gnd.n4192 4.74817
R11497 gnd.n4194 gnd.n1057 4.74817
R11498 gnd.n2551 gnd.n2550 4.74296
R11499 gnd.n62 gnd.n61 4.74296
R11500 gnd.n2527 gnd.n2526 4.7074
R11501 gnd.n2539 gnd.n2538 4.7074
R11502 gnd.n38 gnd.n37 4.7074
R11503 gnd.n50 gnd.n49 4.7074
R11504 gnd.n2551 gnd.n2539 4.65959
R11505 gnd.n62 gnd.n50 4.65959
R11506 gnd.n5600 gnd.n1523 4.6132
R11507 gnd.n5906 gnd.n1213 4.6132
R11508 gnd.n5956 gnd.n1144 4.46168
R11509 gnd.n5831 gnd.n1279 4.46168
R11510 gnd.n4754 gnd.n2051 4.46168
R11511 gnd.n2006 gnd.t23 4.46168
R11512 gnd.n4882 gnd.n1976 4.46168
R11513 gnd.n4917 gnd.n1955 4.46168
R11514 gnd.n4975 gnd.n1877 4.46168
R11515 gnd.n5086 gnd.n1861 4.46168
R11516 gnd.t21 gnd.n1838 4.46168
R11517 gnd.n5196 gnd.t251 4.46168
R11518 gnd.n5190 gnd.n1802 4.46168
R11519 gnd.n5351 gnd.n1708 4.46168
R11520 gnd.n5653 gnd.n1489 4.46168
R11521 gnd.n1729 gnd.n1716 4.46111
R11522 gnd.n3590 gnd.n3586 4.38594
R11523 gnd.n3558 gnd.n3554 4.38594
R11524 gnd.n3526 gnd.n3522 4.38594
R11525 gnd.n3495 gnd.n3491 4.38594
R11526 gnd.n3463 gnd.n3459 4.38594
R11527 gnd.n3431 gnd.n3427 4.38594
R11528 gnd.n3399 gnd.n3395 4.38594
R11529 gnd.n3368 gnd.n3364 4.38594
R11530 gnd.n3601 gnd.n3579 4.26717
R11531 gnd.n3569 gnd.n3547 4.26717
R11532 gnd.n3537 gnd.n3515 4.26717
R11533 gnd.n3506 gnd.n3484 4.26717
R11534 gnd.n3474 gnd.n3452 4.26717
R11535 gnd.n3442 gnd.n3420 4.26717
R11536 gnd.n3410 gnd.n3388 4.26717
R11537 gnd.n3379 gnd.n3357 4.26717
R11538 gnd.n3058 gnd.t7 4.14303
R11539 gnd.n3288 gnd.t1 4.14303
R11540 gnd.n4251 gnd.t93 4.14303
R11541 gnd.t68 gnd.n5498 4.14303
R11542 gnd.n3609 gnd.n3608 4.08274
R11543 gnd.n5278 gnd.n5277 4.05904
R11544 gnd.n4681 gnd.n4680 4.05904
R11545 gnd.n5846 gnd.n5839 4.05904
R11546 gnd.n5295 gnd.n5294 4.05904
R11547 gnd.n15 gnd.n7 3.99943
R11548 gnd.n4827 gnd.t55 3.82437
R11549 gnd.n4963 gnd.t6 3.82437
R11550 gnd.n4969 gnd.t19 3.82437
R11551 gnd.n5154 gnd.t37 3.82437
R11552 gnd.n3131 gnd.n2552 3.81325
R11553 gnd.n2539 gnd.n2527 3.72967
R11554 gnd.n50 gnd.n38 3.72967
R11555 gnd.n3609 gnd.n3481 3.70378
R11556 gnd.n15 gnd.n14 3.60163
R11557 gnd.n3600 gnd.n3581 3.49141
R11558 gnd.n3568 gnd.n3549 3.49141
R11559 gnd.n3536 gnd.n3517 3.49141
R11560 gnd.n3505 gnd.n3486 3.49141
R11561 gnd.n3473 gnd.n3454 3.49141
R11562 gnd.n3441 gnd.n3422 3.49141
R11563 gnd.n3409 gnd.n3390 3.49141
R11564 gnd.n3378 gnd.n3359 3.49141
R11565 gnd.n5618 gnd.n5617 3.29747
R11566 gnd.n5617 gnd.n5616 3.29747
R11567 gnd.n392 gnd.n328 3.29747
R11568 gnd.n387 gnd.n328 3.29747
R11569 gnd.n4036 gnd.n4035 3.29747
R11570 gnd.n4035 gnd.n4034 3.29747
R11571 gnd.n5924 gnd.n5923 3.29747
R11572 gnd.n5923 gnd.n5922 3.29747
R11573 gnd.t302 gnd.n1279 3.18706
R11574 gnd.n5825 gnd.t322 3.18706
R11575 gnd.n5825 gnd.t223 3.18706
R11576 gnd.n4796 gnd.n2036 3.18706
R11577 gnd.n4760 gnd.t31 3.18706
R11578 gnd.n4853 gnd.n4852 3.18706
R11579 gnd.n4926 gnd.n1948 3.18706
R11580 gnd.n5035 gnd.n1893 3.18706
R11581 gnd.n5096 gnd.n1853 3.18706
R11582 gnd.t34 gnd.n1816 3.18706
R11583 gnd.n5197 gnd.n1806 3.18706
R11584 gnd.t233 gnd.n5212 3.18706
R11585 gnd.t248 gnd.n1712 3.18706
R11586 gnd.n144 gnd.n136 3.18706
R11587 gnd.n2637 gnd.t7 2.8684
R11588 gnd.n4748 gnd.t51 2.8684
R11589 gnd.t63 gnd.n1793 2.8684
R11590 gnd.n2540 gnd.t109 2.82907
R11591 gnd.n2540 gnd.t172 2.82907
R11592 gnd.n2542 gnd.t89 2.82907
R11593 gnd.n2542 gnd.t124 2.82907
R11594 gnd.n2544 gnd.t141 2.82907
R11595 gnd.n2544 gnd.t130 2.82907
R11596 gnd.n2546 gnd.t128 2.82907
R11597 gnd.n2546 gnd.t119 2.82907
R11598 gnd.n2548 gnd.t133 2.82907
R11599 gnd.n2548 gnd.t159 2.82907
R11600 gnd.n2505 gnd.t135 2.82907
R11601 gnd.n2505 gnd.t151 2.82907
R11602 gnd.n2507 gnd.t158 2.82907
R11603 gnd.n2507 gnd.t111 2.82907
R11604 gnd.n2509 gnd.t149 2.82907
R11605 gnd.n2509 gnd.t146 2.82907
R11606 gnd.n2511 gnd.t182 2.82907
R11607 gnd.n2511 gnd.t161 2.82907
R11608 gnd.n2513 gnd.t117 2.82907
R11609 gnd.n2513 gnd.t154 2.82907
R11610 gnd.n2516 gnd.t184 2.82907
R11611 gnd.n2516 gnd.t94 2.82907
R11612 gnd.n2518 gnd.t97 2.82907
R11613 gnd.n2518 gnd.t78 2.82907
R11614 gnd.n2520 gnd.t156 2.82907
R11615 gnd.n2520 gnd.t185 2.82907
R11616 gnd.n2522 gnd.t180 2.82907
R11617 gnd.n2522 gnd.t99 2.82907
R11618 gnd.n2524 gnd.t174 2.82907
R11619 gnd.n2524 gnd.t157 2.82907
R11620 gnd.n2528 gnd.t147 2.82907
R11621 gnd.n2528 gnd.t113 2.82907
R11622 gnd.n2530 gnd.t134 2.82907
R11623 gnd.n2530 gnd.t160 2.82907
R11624 gnd.n2532 gnd.t179 2.82907
R11625 gnd.n2532 gnd.t169 2.82907
R11626 gnd.n2534 gnd.t167 2.82907
R11627 gnd.n2534 gnd.t153 2.82907
R11628 gnd.n2536 gnd.t171 2.82907
R11629 gnd.n2536 gnd.t106 2.82907
R11630 gnd.n59 gnd.t137 2.82907
R11631 gnd.n59 gnd.t118 2.82907
R11632 gnd.n57 gnd.t85 2.82907
R11633 gnd.n57 gnd.t104 2.82907
R11634 gnd.n55 gnd.t96 2.82907
R11635 gnd.n55 gnd.t121 2.82907
R11636 gnd.n53 gnd.t101 2.82907
R11637 gnd.n53 gnd.t166 2.82907
R11638 gnd.n51 gnd.t145 2.82907
R11639 gnd.n51 gnd.t82 2.82907
R11640 gnd.n24 gnd.t187 2.82907
R11641 gnd.n24 gnd.t110 2.82907
R11642 gnd.n22 gnd.t92 2.82907
R11643 gnd.n22 gnd.t107 2.82907
R11644 gnd.n20 gnd.t168 2.82907
R11645 gnd.n20 gnd.t142 2.82907
R11646 gnd.n18 gnd.t132 2.82907
R11647 gnd.n18 gnd.t74 2.82907
R11648 gnd.n16 gnd.t178 2.82907
R11649 gnd.n16 gnd.t122 2.82907
R11650 gnd.n35 gnd.t148 2.82907
R11651 gnd.n35 gnd.t76 2.82907
R11652 gnd.n33 gnd.t73 2.82907
R11653 gnd.n33 gnd.t163 2.82907
R11654 gnd.n31 gnd.t170 2.82907
R11655 gnd.n31 gnd.t177 2.82907
R11656 gnd.n29 gnd.t176 2.82907
R11657 gnd.n29 gnd.t71 2.82907
R11658 gnd.n27 gnd.t69 2.82907
R11659 gnd.n27 gnd.t87 2.82907
R11660 gnd.n47 gnd.t175 2.82907
R11661 gnd.n47 gnd.t152 2.82907
R11662 gnd.n45 gnd.t131 2.82907
R11663 gnd.n45 gnd.t143 2.82907
R11664 gnd.n43 gnd.t144 2.82907
R11665 gnd.n43 gnd.t155 2.82907
R11666 gnd.n41 gnd.t138 2.82907
R11667 gnd.n41 gnd.t112 2.82907
R11668 gnd.n39 gnd.t186 2.82907
R11669 gnd.n39 gnd.t126 2.82907
R11670 gnd.n3597 gnd.n3596 2.71565
R11671 gnd.n3565 gnd.n3564 2.71565
R11672 gnd.n3533 gnd.n3532 2.71565
R11673 gnd.n3502 gnd.n3501 2.71565
R11674 gnd.n3470 gnd.n3469 2.71565
R11675 gnd.n3438 gnd.n3437 2.71565
R11676 gnd.n3406 gnd.n3405 2.71565
R11677 gnd.n3375 gnd.n3374 2.71565
R11678 gnd.n2049 gnd.t223 2.54975
R11679 gnd.n4777 gnd.t17 2.54975
R11680 gnd.n5168 gnd.t35 2.54975
R11681 gnd.n5204 gnd.t251 2.54975
R11682 gnd.n5213 gnd.t233 2.54975
R11683 gnd.n3131 gnd.n2553 2.27742
R11684 gnd.n3131 gnd.n2504 2.27742
R11685 gnd.n3131 gnd.n2503 2.27742
R11686 gnd.n3131 gnd.n2502 2.27742
R11687 gnd.n6892 gnd.n81 2.27742
R11688 gnd.n6892 gnd.n80 2.27742
R11689 gnd.n6892 gnd.n79 2.27742
R11690 gnd.n6892 gnd.n74 2.27742
R11691 gnd.n6893 gnd.n6892 2.27742
R11692 gnd.n2186 gnd.n1058 2.27742
R11693 gnd.n4166 gnd.n1058 2.27742
R11694 gnd.n2167 gnd.n1058 2.27742
R11695 gnd.n4193 gnd.n1058 2.27742
R11696 gnd.n1058 gnd.n1057 2.27742
R11697 gnd.n2985 gnd.t263 2.23109
R11698 gnd.n2608 gnd.t9 2.23109
R11699 gnd.n4917 gnd.t10 2.23109
R11700 gnd.n4945 gnd.t196 2.23109
R11701 gnd.n5017 gnd.t13 2.23109
R11702 gnd.n4975 gnd.t53 2.23109
R11703 gnd.n3593 gnd.n3583 1.93989
R11704 gnd.n3561 gnd.n3551 1.93989
R11705 gnd.n3529 gnd.n3519 1.93989
R11706 gnd.n3498 gnd.n3488 1.93989
R11707 gnd.n3466 gnd.n3456 1.93989
R11708 gnd.n3434 gnd.n3424 1.93989
R11709 gnd.n3402 gnd.n3392 1.93989
R11710 gnd.n3371 gnd.n3361 1.93989
R11711 gnd.n4806 gnd.n2026 1.91244
R11712 gnd.n4860 gnd.n1994 1.91244
R11713 gnd.n1943 gnd.n1937 1.91244
R11714 gnd.n5016 gnd.n1898 1.91244
R11715 gnd.n5138 gnd.n5137 1.91244
R11716 gnd.n5167 gnd.n1820 1.91244
R11717 gnd.n5219 gnd.t274 1.91244
R11718 gnd.t65 gnd.n2996 1.59378
R11719 gnd.n3175 gnd.t24 1.59378
R11720 gnd.n2437 gnd.t56 1.59378
R11721 gnd.n4777 gnd.t43 1.59378
R11722 gnd.n5168 gnd.t200 1.59378
R11723 gnd.n2838 gnd.n2830 1.16414
R11724 gnd.n3655 gnd.n2340 1.16414
R11725 gnd.n3592 gnd.n3585 1.16414
R11726 gnd.n3560 gnd.n3553 1.16414
R11727 gnd.n3528 gnd.n3521 1.16414
R11728 gnd.n3497 gnd.n3490 1.16414
R11729 gnd.n3465 gnd.n3458 1.16414
R11730 gnd.n3433 gnd.n3426 1.16414
R11731 gnd.n3401 gnd.n3394 1.16414
R11732 gnd.n3370 gnd.n3363 1.16414
R11733 gnd.n5600 gnd.n5599 0.970197
R11734 gnd.n5906 gnd.n1211 0.970197
R11735 gnd.n3576 gnd.n3544 0.962709
R11736 gnd.n3608 gnd.n3576 0.962709
R11737 gnd.n3449 gnd.n3417 0.962709
R11738 gnd.n3481 gnd.n3449 0.962709
R11739 gnd.n3084 gnd.t198 0.956468
R11740 gnd.n3249 gnd.t26 0.956468
R11741 gnd.n4121 gnd.t116 0.956468
R11742 gnd.n5988 gnd.t93 0.956468
R11743 gnd.t192 gnd.n1218 0.956468
R11744 gnd.n1701 gnd.t190 0.956468
R11745 gnd.n5499 gnd.t68 0.956468
R11746 gnd.n124 gnd.t75 0.956468
R11747 gnd.n2 gnd.n1 0.672012
R11748 gnd.n3 gnd.n2 0.672012
R11749 gnd.n4 gnd.n3 0.672012
R11750 gnd.n5 gnd.n4 0.672012
R11751 gnd.n6 gnd.n5 0.672012
R11752 gnd.n7 gnd.n6 0.672012
R11753 gnd.n9 gnd.n8 0.672012
R11754 gnd.n10 gnd.n9 0.672012
R11755 gnd.n11 gnd.n10 0.672012
R11756 gnd.n12 gnd.n11 0.672012
R11757 gnd.n13 gnd.n12 0.672012
R11758 gnd.n14 gnd.n13 0.672012
R11759 gnd.n2050 gnd.t254 0.637812
R11760 gnd.n4818 gnd.n4817 0.637812
R11761 gnd.n4766 gnd.n4765 0.637812
R11762 gnd.n4939 gnd.n1920 0.637812
R11763 gnd.n5006 gnd.n5005 0.637812
R11764 gnd.n5103 gnd.n1841 0.637812
R11765 gnd.n5160 gnd.n1826 0.637812
R11766 gnd.n2550 gnd.n2549 0.573776
R11767 gnd.n2549 gnd.n2547 0.573776
R11768 gnd.n2547 gnd.n2545 0.573776
R11769 gnd.n2545 gnd.n2543 0.573776
R11770 gnd.n2543 gnd.n2541 0.573776
R11771 gnd.n2515 gnd.n2514 0.573776
R11772 gnd.n2514 gnd.n2512 0.573776
R11773 gnd.n2512 gnd.n2510 0.573776
R11774 gnd.n2510 gnd.n2508 0.573776
R11775 gnd.n2508 gnd.n2506 0.573776
R11776 gnd.n2526 gnd.n2525 0.573776
R11777 gnd.n2525 gnd.n2523 0.573776
R11778 gnd.n2523 gnd.n2521 0.573776
R11779 gnd.n2521 gnd.n2519 0.573776
R11780 gnd.n2519 gnd.n2517 0.573776
R11781 gnd.n2538 gnd.n2537 0.573776
R11782 gnd.n2537 gnd.n2535 0.573776
R11783 gnd.n2535 gnd.n2533 0.573776
R11784 gnd.n2533 gnd.n2531 0.573776
R11785 gnd.n2531 gnd.n2529 0.573776
R11786 gnd.n54 gnd.n52 0.573776
R11787 gnd.n56 gnd.n54 0.573776
R11788 gnd.n58 gnd.n56 0.573776
R11789 gnd.n60 gnd.n58 0.573776
R11790 gnd.n61 gnd.n60 0.573776
R11791 gnd.n19 gnd.n17 0.573776
R11792 gnd.n21 gnd.n19 0.573776
R11793 gnd.n23 gnd.n21 0.573776
R11794 gnd.n25 gnd.n23 0.573776
R11795 gnd.n26 gnd.n25 0.573776
R11796 gnd.n30 gnd.n28 0.573776
R11797 gnd.n32 gnd.n30 0.573776
R11798 gnd.n34 gnd.n32 0.573776
R11799 gnd.n36 gnd.n34 0.573776
R11800 gnd.n37 gnd.n36 0.573776
R11801 gnd.n42 gnd.n40 0.573776
R11802 gnd.n44 gnd.n42 0.573776
R11803 gnd.n46 gnd.n44 0.573776
R11804 gnd.n48 gnd.n46 0.573776
R11805 gnd.n49 gnd.n48 0.573776
R11806 gnd gnd.n0 0.551497
R11807 gnd.n248 gnd.n247 0.532512
R11808 gnd.n3915 gnd.n3913 0.532512
R11809 gnd.n344 gnd.n160 0.497451
R11810 gnd.n5960 gnd.n5959 0.497451
R11811 gnd.n1574 gnd.n1493 0.497451
R11812 gnd.n3775 gnd.n2257 0.497451
R11813 gnd.n5724 gnd.n1375 0.489829
R11814 gnd.n4576 gnd.n2093 0.489829
R11815 gnd.n4295 gnd.n4277 0.489829
R11816 gnd.n5718 gnd.n5717 0.489829
R11817 gnd.n3311 gnd.n2344 0.486781
R11818 gnd.n2887 gnd.n2886 0.48678
R11819 gnd.n3629 gnd.n2298 0.480683
R11820 gnd.n2971 gnd.n2970 0.480683
R11821 gnd.n6904 gnd.n6903 0.470187
R11822 gnd.n6892 gnd.n78 0.420375
R11823 gnd.n4229 gnd.n1058 0.420375
R11824 gnd.n6185 gnd.n6184 0.416659
R11825 gnd.n6507 gnd.n6506 0.416659
R11826 gnd.n4371 gnd.n4362 0.388379
R11827 gnd.n3589 gnd.n3588 0.388379
R11828 gnd.n3557 gnd.n3556 0.388379
R11829 gnd.n3525 gnd.n3524 0.388379
R11830 gnd.n3494 gnd.n3493 0.388379
R11831 gnd.n3462 gnd.n3461 0.388379
R11832 gnd.n3430 gnd.n3429 0.388379
R11833 gnd.n3398 gnd.n3397 0.388379
R11834 gnd.n3367 gnd.n3366 0.388379
R11835 gnd.n5662 gnd.n1441 0.388379
R11836 gnd.n6904 gnd.n15 0.374463
R11837 gnd.n2399 gnd.t58 0.319156
R11838 gnd.n4162 gnd.t98 0.319156
R11839 gnd.t88 gnd.n6012 0.319156
R11840 gnd.n6774 gnd.t70 0.319156
R11841 gnd.n85 gnd.t72 0.319156
R11842 gnd.n2805 gnd.n2783 0.311721
R11843 gnd.n4575 gnd.n2120 0.302329
R11844 gnd.n5433 gnd.n5432 0.302329
R11845 gnd gnd.n6904 0.295112
R11846 gnd.n493 gnd.n280 0.293183
R11847 gnd.n3953 gnd.n3952 0.293183
R11848 gnd.n6718 gnd.n78 0.280988
R11849 gnd.n4229 gnd.n1048 0.280988
R11850 gnd.n3700 gnd.n3699 0.268793
R11851 gnd.n493 gnd.n492 0.258122
R11852 gnd.n5538 gnd.n1394 0.258122
R11853 gnd.n4523 gnd.n4522 0.258122
R11854 gnd.n3954 gnd.n3953 0.258122
R11855 gnd.n3699 gnd.n3698 0.241354
R11856 gnd.n1523 gnd.n1520 0.229039
R11857 gnd.n1524 gnd.n1523 0.229039
R11858 gnd.n1213 gnd.n1210 0.229039
R11859 gnd.n4447 gnd.n1213 0.229039
R11860 gnd.n2959 gnd.n2758 0.206293
R11861 gnd.n3606 gnd.n3578 0.155672
R11862 gnd.n3599 gnd.n3578 0.155672
R11863 gnd.n3599 gnd.n3598 0.155672
R11864 gnd.n3598 gnd.n3582 0.155672
R11865 gnd.n3591 gnd.n3582 0.155672
R11866 gnd.n3591 gnd.n3590 0.155672
R11867 gnd.n3574 gnd.n3546 0.155672
R11868 gnd.n3567 gnd.n3546 0.155672
R11869 gnd.n3567 gnd.n3566 0.155672
R11870 gnd.n3566 gnd.n3550 0.155672
R11871 gnd.n3559 gnd.n3550 0.155672
R11872 gnd.n3559 gnd.n3558 0.155672
R11873 gnd.n3542 gnd.n3514 0.155672
R11874 gnd.n3535 gnd.n3514 0.155672
R11875 gnd.n3535 gnd.n3534 0.155672
R11876 gnd.n3534 gnd.n3518 0.155672
R11877 gnd.n3527 gnd.n3518 0.155672
R11878 gnd.n3527 gnd.n3526 0.155672
R11879 gnd.n3511 gnd.n3483 0.155672
R11880 gnd.n3504 gnd.n3483 0.155672
R11881 gnd.n3504 gnd.n3503 0.155672
R11882 gnd.n3503 gnd.n3487 0.155672
R11883 gnd.n3496 gnd.n3487 0.155672
R11884 gnd.n3496 gnd.n3495 0.155672
R11885 gnd.n3479 gnd.n3451 0.155672
R11886 gnd.n3472 gnd.n3451 0.155672
R11887 gnd.n3472 gnd.n3471 0.155672
R11888 gnd.n3471 gnd.n3455 0.155672
R11889 gnd.n3464 gnd.n3455 0.155672
R11890 gnd.n3464 gnd.n3463 0.155672
R11891 gnd.n3447 gnd.n3419 0.155672
R11892 gnd.n3440 gnd.n3419 0.155672
R11893 gnd.n3440 gnd.n3439 0.155672
R11894 gnd.n3439 gnd.n3423 0.155672
R11895 gnd.n3432 gnd.n3423 0.155672
R11896 gnd.n3432 gnd.n3431 0.155672
R11897 gnd.n3415 gnd.n3387 0.155672
R11898 gnd.n3408 gnd.n3387 0.155672
R11899 gnd.n3408 gnd.n3407 0.155672
R11900 gnd.n3407 gnd.n3391 0.155672
R11901 gnd.n3400 gnd.n3391 0.155672
R11902 gnd.n3400 gnd.n3399 0.155672
R11903 gnd.n3384 gnd.n3356 0.155672
R11904 gnd.n3377 gnd.n3356 0.155672
R11905 gnd.n3377 gnd.n3376 0.155672
R11906 gnd.n3376 gnd.n3360 0.155672
R11907 gnd.n3369 gnd.n3360 0.155672
R11908 gnd.n3369 gnd.n3368 0.155672
R11909 gnd.n3731 gnd.n2298 0.152939
R11910 gnd.n3731 gnd.n3730 0.152939
R11911 gnd.n3730 gnd.n3729 0.152939
R11912 gnd.n3729 gnd.n2300 0.152939
R11913 gnd.n2301 gnd.n2300 0.152939
R11914 gnd.n2302 gnd.n2301 0.152939
R11915 gnd.n2303 gnd.n2302 0.152939
R11916 gnd.n2304 gnd.n2303 0.152939
R11917 gnd.n2305 gnd.n2304 0.152939
R11918 gnd.n2306 gnd.n2305 0.152939
R11919 gnd.n2307 gnd.n2306 0.152939
R11920 gnd.n2308 gnd.n2307 0.152939
R11921 gnd.n2309 gnd.n2308 0.152939
R11922 gnd.n2310 gnd.n2309 0.152939
R11923 gnd.n3701 gnd.n2310 0.152939
R11924 gnd.n3701 gnd.n3700 0.152939
R11925 gnd.n2972 gnd.n2971 0.152939
R11926 gnd.n2972 gnd.n2676 0.152939
R11927 gnd.n3000 gnd.n2676 0.152939
R11928 gnd.n3001 gnd.n3000 0.152939
R11929 gnd.n3002 gnd.n3001 0.152939
R11930 gnd.n3003 gnd.n3002 0.152939
R11931 gnd.n3003 gnd.n2648 0.152939
R11932 gnd.n3030 gnd.n2648 0.152939
R11933 gnd.n3031 gnd.n3030 0.152939
R11934 gnd.n3032 gnd.n3031 0.152939
R11935 gnd.n3032 gnd.n2626 0.152939
R11936 gnd.n3061 gnd.n2626 0.152939
R11937 gnd.n3062 gnd.n3061 0.152939
R11938 gnd.n3063 gnd.n3062 0.152939
R11939 gnd.n3064 gnd.n3063 0.152939
R11940 gnd.n3066 gnd.n3064 0.152939
R11941 gnd.n3066 gnd.n3065 0.152939
R11942 gnd.n3065 gnd.n2575 0.152939
R11943 gnd.n2576 gnd.n2575 0.152939
R11944 gnd.n2577 gnd.n2576 0.152939
R11945 gnd.n2596 gnd.n2577 0.152939
R11946 gnd.n2597 gnd.n2596 0.152939
R11947 gnd.n2597 gnd.n2495 0.152939
R11948 gnd.n3156 gnd.n2495 0.152939
R11949 gnd.n3157 gnd.n3156 0.152939
R11950 gnd.n3158 gnd.n3157 0.152939
R11951 gnd.n3159 gnd.n3158 0.152939
R11952 gnd.n3159 gnd.n2468 0.152939
R11953 gnd.n3196 gnd.n2468 0.152939
R11954 gnd.n3197 gnd.n3196 0.152939
R11955 gnd.n3198 gnd.n3197 0.152939
R11956 gnd.n3199 gnd.n3198 0.152939
R11957 gnd.n3199 gnd.n2441 0.152939
R11958 gnd.n3241 gnd.n2441 0.152939
R11959 gnd.n3242 gnd.n3241 0.152939
R11960 gnd.n3243 gnd.n3242 0.152939
R11961 gnd.n3244 gnd.n3243 0.152939
R11962 gnd.n3244 gnd.n2413 0.152939
R11963 gnd.n3281 gnd.n2413 0.152939
R11964 gnd.n3282 gnd.n3281 0.152939
R11965 gnd.n3283 gnd.n3282 0.152939
R11966 gnd.n3284 gnd.n3283 0.152939
R11967 gnd.n3284 gnd.n2386 0.152939
R11968 gnd.n3330 gnd.n2386 0.152939
R11969 gnd.n3331 gnd.n3330 0.152939
R11970 gnd.n3332 gnd.n3331 0.152939
R11971 gnd.n3333 gnd.n3332 0.152939
R11972 gnd.n3333 gnd.n2359 0.152939
R11973 gnd.n3625 gnd.n2359 0.152939
R11974 gnd.n3626 gnd.n3625 0.152939
R11975 gnd.n3627 gnd.n3626 0.152939
R11976 gnd.n3628 gnd.n3627 0.152939
R11977 gnd.n3629 gnd.n3628 0.152939
R11978 gnd.n2970 gnd.n2700 0.152939
R11979 gnd.n2721 gnd.n2700 0.152939
R11980 gnd.n2722 gnd.n2721 0.152939
R11981 gnd.n2728 gnd.n2722 0.152939
R11982 gnd.n2729 gnd.n2728 0.152939
R11983 gnd.n2730 gnd.n2729 0.152939
R11984 gnd.n2730 gnd.n2719 0.152939
R11985 gnd.n2738 gnd.n2719 0.152939
R11986 gnd.n2739 gnd.n2738 0.152939
R11987 gnd.n2740 gnd.n2739 0.152939
R11988 gnd.n2740 gnd.n2717 0.152939
R11989 gnd.n2748 gnd.n2717 0.152939
R11990 gnd.n2749 gnd.n2748 0.152939
R11991 gnd.n2750 gnd.n2749 0.152939
R11992 gnd.n2750 gnd.n2715 0.152939
R11993 gnd.n2758 gnd.n2715 0.152939
R11994 gnd.n3698 gnd.n2315 0.152939
R11995 gnd.n2317 gnd.n2315 0.152939
R11996 gnd.n2318 gnd.n2317 0.152939
R11997 gnd.n2319 gnd.n2318 0.152939
R11998 gnd.n2320 gnd.n2319 0.152939
R11999 gnd.n2321 gnd.n2320 0.152939
R12000 gnd.n2322 gnd.n2321 0.152939
R12001 gnd.n2323 gnd.n2322 0.152939
R12002 gnd.n2324 gnd.n2323 0.152939
R12003 gnd.n2325 gnd.n2324 0.152939
R12004 gnd.n2326 gnd.n2325 0.152939
R12005 gnd.n2327 gnd.n2326 0.152939
R12006 gnd.n2328 gnd.n2327 0.152939
R12007 gnd.n2329 gnd.n2328 0.152939
R12008 gnd.n2330 gnd.n2329 0.152939
R12009 gnd.n2331 gnd.n2330 0.152939
R12010 gnd.n2332 gnd.n2331 0.152939
R12011 gnd.n2333 gnd.n2332 0.152939
R12012 gnd.n2334 gnd.n2333 0.152939
R12013 gnd.n2335 gnd.n2334 0.152939
R12014 gnd.n2336 gnd.n2335 0.152939
R12015 gnd.n2337 gnd.n2336 0.152939
R12016 gnd.n2341 gnd.n2337 0.152939
R12017 gnd.n2342 gnd.n2341 0.152939
R12018 gnd.n2343 gnd.n2342 0.152939
R12019 gnd.n2344 gnd.n2343 0.152939
R12020 gnd.n3133 gnd.n3132 0.152939
R12021 gnd.n3134 gnd.n3133 0.152939
R12022 gnd.n3135 gnd.n3134 0.152939
R12023 gnd.n3136 gnd.n3135 0.152939
R12024 gnd.n3137 gnd.n3136 0.152939
R12025 gnd.n3138 gnd.n3137 0.152939
R12026 gnd.n3138 gnd.n2449 0.152939
R12027 gnd.n3217 gnd.n2449 0.152939
R12028 gnd.n3218 gnd.n3217 0.152939
R12029 gnd.n3219 gnd.n3218 0.152939
R12030 gnd.n3220 gnd.n3219 0.152939
R12031 gnd.n3221 gnd.n3220 0.152939
R12032 gnd.n3222 gnd.n3221 0.152939
R12033 gnd.n3223 gnd.n3222 0.152939
R12034 gnd.n3224 gnd.n3223 0.152939
R12035 gnd.n3225 gnd.n3224 0.152939
R12036 gnd.n3225 gnd.n2393 0.152939
R12037 gnd.n3302 gnd.n2393 0.152939
R12038 gnd.n3303 gnd.n3302 0.152939
R12039 gnd.n3304 gnd.n3303 0.152939
R12040 gnd.n3305 gnd.n3304 0.152939
R12041 gnd.n3306 gnd.n3305 0.152939
R12042 gnd.n3307 gnd.n3306 0.152939
R12043 gnd.n3308 gnd.n3307 0.152939
R12044 gnd.n3309 gnd.n3308 0.152939
R12045 gnd.n3310 gnd.n3309 0.152939
R12046 gnd.n3312 gnd.n3310 0.152939
R12047 gnd.n3312 gnd.n3311 0.152939
R12048 gnd.n2888 gnd.n2887 0.152939
R12049 gnd.n2888 gnd.n2778 0.152939
R12050 gnd.n2903 gnd.n2778 0.152939
R12051 gnd.n2904 gnd.n2903 0.152939
R12052 gnd.n2905 gnd.n2904 0.152939
R12053 gnd.n2905 gnd.n2766 0.152939
R12054 gnd.n2919 gnd.n2766 0.152939
R12055 gnd.n2920 gnd.n2919 0.152939
R12056 gnd.n2921 gnd.n2920 0.152939
R12057 gnd.n2922 gnd.n2921 0.152939
R12058 gnd.n2923 gnd.n2922 0.152939
R12059 gnd.n2924 gnd.n2923 0.152939
R12060 gnd.n2925 gnd.n2924 0.152939
R12061 gnd.n2926 gnd.n2925 0.152939
R12062 gnd.n2927 gnd.n2926 0.152939
R12063 gnd.n2928 gnd.n2927 0.152939
R12064 gnd.n2929 gnd.n2928 0.152939
R12065 gnd.n2930 gnd.n2929 0.152939
R12066 gnd.n2931 gnd.n2930 0.152939
R12067 gnd.n2932 gnd.n2931 0.152939
R12068 gnd.n2933 gnd.n2932 0.152939
R12069 gnd.n2933 gnd.n2632 0.152939
R12070 gnd.n3050 gnd.n2632 0.152939
R12071 gnd.n3051 gnd.n3050 0.152939
R12072 gnd.n3052 gnd.n3051 0.152939
R12073 gnd.n3053 gnd.n3052 0.152939
R12074 gnd.n3053 gnd.n2554 0.152939
R12075 gnd.n3130 gnd.n2554 0.152939
R12076 gnd.n2806 gnd.n2805 0.152939
R12077 gnd.n2807 gnd.n2806 0.152939
R12078 gnd.n2808 gnd.n2807 0.152939
R12079 gnd.n2809 gnd.n2808 0.152939
R12080 gnd.n2810 gnd.n2809 0.152939
R12081 gnd.n2811 gnd.n2810 0.152939
R12082 gnd.n2812 gnd.n2811 0.152939
R12083 gnd.n2813 gnd.n2812 0.152939
R12084 gnd.n2814 gnd.n2813 0.152939
R12085 gnd.n2815 gnd.n2814 0.152939
R12086 gnd.n2816 gnd.n2815 0.152939
R12087 gnd.n2817 gnd.n2816 0.152939
R12088 gnd.n2818 gnd.n2817 0.152939
R12089 gnd.n2819 gnd.n2818 0.152939
R12090 gnd.n2820 gnd.n2819 0.152939
R12091 gnd.n2821 gnd.n2820 0.152939
R12092 gnd.n2822 gnd.n2821 0.152939
R12093 gnd.n2823 gnd.n2822 0.152939
R12094 gnd.n2824 gnd.n2823 0.152939
R12095 gnd.n2825 gnd.n2824 0.152939
R12096 gnd.n2826 gnd.n2825 0.152939
R12097 gnd.n2827 gnd.n2826 0.152939
R12098 gnd.n2831 gnd.n2827 0.152939
R12099 gnd.n2832 gnd.n2831 0.152939
R12100 gnd.n2832 gnd.n2789 0.152939
R12101 gnd.n2886 gnd.n2789 0.152939
R12102 gnd.n6186 gnd.n6185 0.152939
R12103 gnd.n6186 gnd.n875 0.152939
R12104 gnd.n6194 gnd.n875 0.152939
R12105 gnd.n6195 gnd.n6194 0.152939
R12106 gnd.n6196 gnd.n6195 0.152939
R12107 gnd.n6196 gnd.n869 0.152939
R12108 gnd.n6204 gnd.n869 0.152939
R12109 gnd.n6205 gnd.n6204 0.152939
R12110 gnd.n6206 gnd.n6205 0.152939
R12111 gnd.n6206 gnd.n863 0.152939
R12112 gnd.n6214 gnd.n863 0.152939
R12113 gnd.n6215 gnd.n6214 0.152939
R12114 gnd.n6216 gnd.n6215 0.152939
R12115 gnd.n6216 gnd.n857 0.152939
R12116 gnd.n6224 gnd.n857 0.152939
R12117 gnd.n6225 gnd.n6224 0.152939
R12118 gnd.n6226 gnd.n6225 0.152939
R12119 gnd.n6226 gnd.n851 0.152939
R12120 gnd.n6234 gnd.n851 0.152939
R12121 gnd.n6235 gnd.n6234 0.152939
R12122 gnd.n6236 gnd.n6235 0.152939
R12123 gnd.n6236 gnd.n845 0.152939
R12124 gnd.n6244 gnd.n845 0.152939
R12125 gnd.n6245 gnd.n6244 0.152939
R12126 gnd.n6246 gnd.n6245 0.152939
R12127 gnd.n6246 gnd.n839 0.152939
R12128 gnd.n6254 gnd.n839 0.152939
R12129 gnd.n6255 gnd.n6254 0.152939
R12130 gnd.n6256 gnd.n6255 0.152939
R12131 gnd.n6256 gnd.n833 0.152939
R12132 gnd.n6264 gnd.n833 0.152939
R12133 gnd.n6265 gnd.n6264 0.152939
R12134 gnd.n6266 gnd.n6265 0.152939
R12135 gnd.n6266 gnd.n827 0.152939
R12136 gnd.n6274 gnd.n827 0.152939
R12137 gnd.n6275 gnd.n6274 0.152939
R12138 gnd.n6276 gnd.n6275 0.152939
R12139 gnd.n6276 gnd.n821 0.152939
R12140 gnd.n6284 gnd.n821 0.152939
R12141 gnd.n6285 gnd.n6284 0.152939
R12142 gnd.n6286 gnd.n6285 0.152939
R12143 gnd.n6286 gnd.n815 0.152939
R12144 gnd.n6294 gnd.n815 0.152939
R12145 gnd.n6295 gnd.n6294 0.152939
R12146 gnd.n6296 gnd.n6295 0.152939
R12147 gnd.n6296 gnd.n809 0.152939
R12148 gnd.n6304 gnd.n809 0.152939
R12149 gnd.n6305 gnd.n6304 0.152939
R12150 gnd.n6306 gnd.n6305 0.152939
R12151 gnd.n6306 gnd.n803 0.152939
R12152 gnd.n6314 gnd.n803 0.152939
R12153 gnd.n6315 gnd.n6314 0.152939
R12154 gnd.n6316 gnd.n6315 0.152939
R12155 gnd.n6316 gnd.n797 0.152939
R12156 gnd.n6324 gnd.n797 0.152939
R12157 gnd.n6325 gnd.n6324 0.152939
R12158 gnd.n6326 gnd.n6325 0.152939
R12159 gnd.n6326 gnd.n791 0.152939
R12160 gnd.n6334 gnd.n791 0.152939
R12161 gnd.n6335 gnd.n6334 0.152939
R12162 gnd.n6336 gnd.n6335 0.152939
R12163 gnd.n6336 gnd.n785 0.152939
R12164 gnd.n6344 gnd.n785 0.152939
R12165 gnd.n6345 gnd.n6344 0.152939
R12166 gnd.n6346 gnd.n6345 0.152939
R12167 gnd.n6346 gnd.n779 0.152939
R12168 gnd.n6354 gnd.n779 0.152939
R12169 gnd.n6355 gnd.n6354 0.152939
R12170 gnd.n6356 gnd.n6355 0.152939
R12171 gnd.n6356 gnd.n773 0.152939
R12172 gnd.n6364 gnd.n773 0.152939
R12173 gnd.n6365 gnd.n6364 0.152939
R12174 gnd.n6366 gnd.n6365 0.152939
R12175 gnd.n6366 gnd.n767 0.152939
R12176 gnd.n6374 gnd.n767 0.152939
R12177 gnd.n6375 gnd.n6374 0.152939
R12178 gnd.n6376 gnd.n6375 0.152939
R12179 gnd.n6376 gnd.n761 0.152939
R12180 gnd.n6384 gnd.n761 0.152939
R12181 gnd.n6385 gnd.n6384 0.152939
R12182 gnd.n6386 gnd.n6385 0.152939
R12183 gnd.n6386 gnd.n755 0.152939
R12184 gnd.n6394 gnd.n755 0.152939
R12185 gnd.n6395 gnd.n6394 0.152939
R12186 gnd.n6396 gnd.n6395 0.152939
R12187 gnd.n6396 gnd.n749 0.152939
R12188 gnd.n6404 gnd.n749 0.152939
R12189 gnd.n6405 gnd.n6404 0.152939
R12190 gnd.n6406 gnd.n6405 0.152939
R12191 gnd.n6406 gnd.n743 0.152939
R12192 gnd.n6414 gnd.n743 0.152939
R12193 gnd.n6415 gnd.n6414 0.152939
R12194 gnd.n6416 gnd.n6415 0.152939
R12195 gnd.n6416 gnd.n737 0.152939
R12196 gnd.n6424 gnd.n737 0.152939
R12197 gnd.n6425 gnd.n6424 0.152939
R12198 gnd.n6426 gnd.n6425 0.152939
R12199 gnd.n6426 gnd.n731 0.152939
R12200 gnd.n6434 gnd.n731 0.152939
R12201 gnd.n6435 gnd.n6434 0.152939
R12202 gnd.n6436 gnd.n6435 0.152939
R12203 gnd.n6436 gnd.n725 0.152939
R12204 gnd.n6444 gnd.n725 0.152939
R12205 gnd.n6445 gnd.n6444 0.152939
R12206 gnd.n6446 gnd.n6445 0.152939
R12207 gnd.n6446 gnd.n719 0.152939
R12208 gnd.n6454 gnd.n719 0.152939
R12209 gnd.n6455 gnd.n6454 0.152939
R12210 gnd.n6456 gnd.n6455 0.152939
R12211 gnd.n6456 gnd.n713 0.152939
R12212 gnd.n6464 gnd.n713 0.152939
R12213 gnd.n6465 gnd.n6464 0.152939
R12214 gnd.n6466 gnd.n6465 0.152939
R12215 gnd.n6466 gnd.n707 0.152939
R12216 gnd.n6474 gnd.n707 0.152939
R12217 gnd.n6475 gnd.n6474 0.152939
R12218 gnd.n6476 gnd.n6475 0.152939
R12219 gnd.n6476 gnd.n701 0.152939
R12220 gnd.n6484 gnd.n701 0.152939
R12221 gnd.n6485 gnd.n6484 0.152939
R12222 gnd.n6486 gnd.n6485 0.152939
R12223 gnd.n6486 gnd.n695 0.152939
R12224 gnd.n6494 gnd.n695 0.152939
R12225 gnd.n6495 gnd.n6494 0.152939
R12226 gnd.n6497 gnd.n6495 0.152939
R12227 gnd.n6497 gnd.n6496 0.152939
R12228 gnd.n6496 gnd.n689 0.152939
R12229 gnd.n6506 gnd.n689 0.152939
R12230 gnd.n6507 gnd.n684 0.152939
R12231 gnd.n6515 gnd.n684 0.152939
R12232 gnd.n6516 gnd.n6515 0.152939
R12233 gnd.n6517 gnd.n6516 0.152939
R12234 gnd.n6517 gnd.n678 0.152939
R12235 gnd.n6525 gnd.n678 0.152939
R12236 gnd.n6526 gnd.n6525 0.152939
R12237 gnd.n6527 gnd.n6526 0.152939
R12238 gnd.n6527 gnd.n672 0.152939
R12239 gnd.n6535 gnd.n672 0.152939
R12240 gnd.n6536 gnd.n6535 0.152939
R12241 gnd.n6537 gnd.n6536 0.152939
R12242 gnd.n6537 gnd.n666 0.152939
R12243 gnd.n6545 gnd.n666 0.152939
R12244 gnd.n6546 gnd.n6545 0.152939
R12245 gnd.n6547 gnd.n6546 0.152939
R12246 gnd.n6547 gnd.n660 0.152939
R12247 gnd.n6555 gnd.n660 0.152939
R12248 gnd.n6556 gnd.n6555 0.152939
R12249 gnd.n6557 gnd.n6556 0.152939
R12250 gnd.n6557 gnd.n654 0.152939
R12251 gnd.n6565 gnd.n654 0.152939
R12252 gnd.n6566 gnd.n6565 0.152939
R12253 gnd.n6567 gnd.n6566 0.152939
R12254 gnd.n6567 gnd.n648 0.152939
R12255 gnd.n6575 gnd.n648 0.152939
R12256 gnd.n6576 gnd.n6575 0.152939
R12257 gnd.n6577 gnd.n6576 0.152939
R12258 gnd.n6577 gnd.n642 0.152939
R12259 gnd.n6585 gnd.n642 0.152939
R12260 gnd.n6586 gnd.n6585 0.152939
R12261 gnd.n6587 gnd.n6586 0.152939
R12262 gnd.n6587 gnd.n636 0.152939
R12263 gnd.n6595 gnd.n636 0.152939
R12264 gnd.n6596 gnd.n6595 0.152939
R12265 gnd.n6597 gnd.n6596 0.152939
R12266 gnd.n6597 gnd.n630 0.152939
R12267 gnd.n6605 gnd.n630 0.152939
R12268 gnd.n6606 gnd.n6605 0.152939
R12269 gnd.n6607 gnd.n6606 0.152939
R12270 gnd.n6607 gnd.n624 0.152939
R12271 gnd.n6615 gnd.n624 0.152939
R12272 gnd.n6616 gnd.n6615 0.152939
R12273 gnd.n6617 gnd.n6616 0.152939
R12274 gnd.n6617 gnd.n618 0.152939
R12275 gnd.n6625 gnd.n618 0.152939
R12276 gnd.n6626 gnd.n6625 0.152939
R12277 gnd.n6627 gnd.n6626 0.152939
R12278 gnd.n6627 gnd.n612 0.152939
R12279 gnd.n6635 gnd.n612 0.152939
R12280 gnd.n6636 gnd.n6635 0.152939
R12281 gnd.n6637 gnd.n6636 0.152939
R12282 gnd.n6637 gnd.n606 0.152939
R12283 gnd.n6645 gnd.n606 0.152939
R12284 gnd.n6646 gnd.n6645 0.152939
R12285 gnd.n6647 gnd.n6646 0.152939
R12286 gnd.n6647 gnd.n600 0.152939
R12287 gnd.n6655 gnd.n600 0.152939
R12288 gnd.n6656 gnd.n6655 0.152939
R12289 gnd.n6657 gnd.n6656 0.152939
R12290 gnd.n6657 gnd.n594 0.152939
R12291 gnd.n6665 gnd.n594 0.152939
R12292 gnd.n6666 gnd.n6665 0.152939
R12293 gnd.n6667 gnd.n6666 0.152939
R12294 gnd.n6667 gnd.n588 0.152939
R12295 gnd.n6675 gnd.n588 0.152939
R12296 gnd.n6676 gnd.n6675 0.152939
R12297 gnd.n6677 gnd.n6676 0.152939
R12298 gnd.n6677 gnd.n582 0.152939
R12299 gnd.n6685 gnd.n582 0.152939
R12300 gnd.n6686 gnd.n6685 0.152939
R12301 gnd.n6687 gnd.n6686 0.152939
R12302 gnd.n6687 gnd.n576 0.152939
R12303 gnd.n6695 gnd.n576 0.152939
R12304 gnd.n6696 gnd.n6695 0.152939
R12305 gnd.n6697 gnd.n6696 0.152939
R12306 gnd.n6697 gnd.n570 0.152939
R12307 gnd.n6705 gnd.n570 0.152939
R12308 gnd.n6706 gnd.n6705 0.152939
R12309 gnd.n6707 gnd.n6706 0.152939
R12310 gnd.n6707 gnd.n564 0.152939
R12311 gnd.n6716 gnd.n564 0.152939
R12312 gnd.n6717 gnd.n6716 0.152939
R12313 gnd.n6718 gnd.n6717 0.152939
R12314 gnd.n6892 gnd.n76 0.152939
R12315 gnd.n101 gnd.n76 0.152939
R12316 gnd.n102 gnd.n101 0.152939
R12317 gnd.n103 gnd.n102 0.152939
R12318 gnd.n118 gnd.n103 0.152939
R12319 gnd.n119 gnd.n118 0.152939
R12320 gnd.n120 gnd.n119 0.152939
R12321 gnd.n121 gnd.n120 0.152939
R12322 gnd.n138 gnd.n121 0.152939
R12323 gnd.n139 gnd.n138 0.152939
R12324 gnd.n140 gnd.n139 0.152939
R12325 gnd.n141 gnd.n140 0.152939
R12326 gnd.n157 gnd.n141 0.152939
R12327 gnd.n158 gnd.n157 0.152939
R12328 gnd.n159 gnd.n158 0.152939
R12329 gnd.n160 gnd.n159 0.152939
R12330 gnd.n6901 gnd.n65 0.152939
R12331 gnd.n214 gnd.n65 0.152939
R12332 gnd.n215 gnd.n214 0.152939
R12333 gnd.n219 gnd.n215 0.152939
R12334 gnd.n220 gnd.n219 0.152939
R12335 gnd.n221 gnd.n220 0.152939
R12336 gnd.n221 gnd.n211 0.152939
R12337 gnd.n226 gnd.n211 0.152939
R12338 gnd.n227 gnd.n226 0.152939
R12339 gnd.n228 gnd.n227 0.152939
R12340 gnd.n228 gnd.n208 0.152939
R12341 gnd.n233 gnd.n208 0.152939
R12342 gnd.n234 gnd.n233 0.152939
R12343 gnd.n235 gnd.n234 0.152939
R12344 gnd.n235 gnd.n205 0.152939
R12345 gnd.n240 gnd.n205 0.152939
R12346 gnd.n241 gnd.n240 0.152939
R12347 gnd.n242 gnd.n241 0.152939
R12348 gnd.n242 gnd.n202 0.152939
R12349 gnd.n247 gnd.n202 0.152939
R12350 gnd.n280 gnd.n168 0.152939
R12351 gnd.n170 gnd.n168 0.152939
R12352 gnd.n174 gnd.n170 0.152939
R12353 gnd.n175 gnd.n174 0.152939
R12354 gnd.n176 gnd.n175 0.152939
R12355 gnd.n177 gnd.n176 0.152939
R12356 gnd.n181 gnd.n177 0.152939
R12357 gnd.n182 gnd.n181 0.152939
R12358 gnd.n183 gnd.n182 0.152939
R12359 gnd.n184 gnd.n183 0.152939
R12360 gnd.n188 gnd.n184 0.152939
R12361 gnd.n189 gnd.n188 0.152939
R12362 gnd.n190 gnd.n189 0.152939
R12363 gnd.n191 gnd.n190 0.152939
R12364 gnd.n195 gnd.n191 0.152939
R12365 gnd.n196 gnd.n195 0.152939
R12366 gnd.n249 gnd.n196 0.152939
R12367 gnd.n249 gnd.n248 0.152939
R12368 gnd.n344 gnd.n343 0.152939
R12369 gnd.n352 gnd.n343 0.152939
R12370 gnd.n353 gnd.n352 0.152939
R12371 gnd.n354 gnd.n353 0.152939
R12372 gnd.n354 gnd.n339 0.152939
R12373 gnd.n362 gnd.n339 0.152939
R12374 gnd.n363 gnd.n362 0.152939
R12375 gnd.n364 gnd.n363 0.152939
R12376 gnd.n364 gnd.n335 0.152939
R12377 gnd.n372 gnd.n335 0.152939
R12378 gnd.n373 gnd.n372 0.152939
R12379 gnd.n374 gnd.n373 0.152939
R12380 gnd.n374 gnd.n331 0.152939
R12381 gnd.n383 gnd.n331 0.152939
R12382 gnd.n384 gnd.n383 0.152939
R12383 gnd.n385 gnd.n384 0.152939
R12384 gnd.n385 gnd.n325 0.152939
R12385 gnd.n393 gnd.n325 0.152939
R12386 gnd.n394 gnd.n393 0.152939
R12387 gnd.n395 gnd.n394 0.152939
R12388 gnd.n395 gnd.n321 0.152939
R12389 gnd.n403 gnd.n321 0.152939
R12390 gnd.n404 gnd.n403 0.152939
R12391 gnd.n405 gnd.n404 0.152939
R12392 gnd.n405 gnd.n317 0.152939
R12393 gnd.n413 gnd.n317 0.152939
R12394 gnd.n414 gnd.n413 0.152939
R12395 gnd.n415 gnd.n414 0.152939
R12396 gnd.n415 gnd.n313 0.152939
R12397 gnd.n423 gnd.n313 0.152939
R12398 gnd.n424 gnd.n423 0.152939
R12399 gnd.n425 gnd.n424 0.152939
R12400 gnd.n425 gnd.n309 0.152939
R12401 gnd.n433 gnd.n309 0.152939
R12402 gnd.n434 gnd.n433 0.152939
R12403 gnd.n435 gnd.n434 0.152939
R12404 gnd.n435 gnd.n303 0.152939
R12405 gnd.n443 gnd.n303 0.152939
R12406 gnd.n444 gnd.n443 0.152939
R12407 gnd.n445 gnd.n444 0.152939
R12408 gnd.n445 gnd.n299 0.152939
R12409 gnd.n453 gnd.n299 0.152939
R12410 gnd.n454 gnd.n453 0.152939
R12411 gnd.n455 gnd.n454 0.152939
R12412 gnd.n455 gnd.n295 0.152939
R12413 gnd.n463 gnd.n295 0.152939
R12414 gnd.n464 gnd.n463 0.152939
R12415 gnd.n465 gnd.n464 0.152939
R12416 gnd.n465 gnd.n291 0.152939
R12417 gnd.n473 gnd.n291 0.152939
R12418 gnd.n474 gnd.n473 0.152939
R12419 gnd.n475 gnd.n474 0.152939
R12420 gnd.n475 gnd.n287 0.152939
R12421 gnd.n483 gnd.n287 0.152939
R12422 gnd.n484 gnd.n483 0.152939
R12423 gnd.n485 gnd.n484 0.152939
R12424 gnd.n485 gnd.n281 0.152939
R12425 gnd.n492 gnd.n281 0.152939
R12426 gnd.n1494 gnd.n1493 0.152939
R12427 gnd.n1495 gnd.n1494 0.152939
R12428 gnd.n1496 gnd.n1495 0.152939
R12429 gnd.n1497 gnd.n1496 0.152939
R12430 gnd.n1498 gnd.n1497 0.152939
R12431 gnd.n1499 gnd.n1498 0.152939
R12432 gnd.n1500 gnd.n1499 0.152939
R12433 gnd.n1501 gnd.n1500 0.152939
R12434 gnd.n1502 gnd.n1501 0.152939
R12435 gnd.n1503 gnd.n1502 0.152939
R12436 gnd.n1504 gnd.n1503 0.152939
R12437 gnd.n1505 gnd.n1504 0.152939
R12438 gnd.n1506 gnd.n1505 0.152939
R12439 gnd.n1507 gnd.n1506 0.152939
R12440 gnd.n1508 gnd.n1507 0.152939
R12441 gnd.n1509 gnd.n1508 0.152939
R12442 gnd.n1510 gnd.n1509 0.152939
R12443 gnd.n1513 gnd.n1510 0.152939
R12444 gnd.n1514 gnd.n1513 0.152939
R12445 gnd.n1515 gnd.n1514 0.152939
R12446 gnd.n1516 gnd.n1515 0.152939
R12447 gnd.n1517 gnd.n1516 0.152939
R12448 gnd.n1518 gnd.n1517 0.152939
R12449 gnd.n1519 gnd.n1518 0.152939
R12450 gnd.n1520 gnd.n1519 0.152939
R12451 gnd.n1525 gnd.n1524 0.152939
R12452 gnd.n1526 gnd.n1525 0.152939
R12453 gnd.n1527 gnd.n1526 0.152939
R12454 gnd.n1528 gnd.n1527 0.152939
R12455 gnd.n1529 gnd.n1528 0.152939
R12456 gnd.n1530 gnd.n1529 0.152939
R12457 gnd.n1531 gnd.n1530 0.152939
R12458 gnd.n1532 gnd.n1531 0.152939
R12459 gnd.n1533 gnd.n1532 0.152939
R12460 gnd.n1536 gnd.n1533 0.152939
R12461 gnd.n1537 gnd.n1536 0.152939
R12462 gnd.n1538 gnd.n1537 0.152939
R12463 gnd.n1539 gnd.n1538 0.152939
R12464 gnd.n1540 gnd.n1539 0.152939
R12465 gnd.n1541 gnd.n1540 0.152939
R12466 gnd.n1542 gnd.n1541 0.152939
R12467 gnd.n1543 gnd.n1542 0.152939
R12468 gnd.n1544 gnd.n1543 0.152939
R12469 gnd.n1545 gnd.n1544 0.152939
R12470 gnd.n1546 gnd.n1545 0.152939
R12471 gnd.n1547 gnd.n1546 0.152939
R12472 gnd.n1548 gnd.n1547 0.152939
R12473 gnd.n1549 gnd.n1548 0.152939
R12474 gnd.n1550 gnd.n1549 0.152939
R12475 gnd.n1551 gnd.n1550 0.152939
R12476 gnd.n1552 gnd.n1551 0.152939
R12477 gnd.n1553 gnd.n1552 0.152939
R12478 gnd.n1554 gnd.n1553 0.152939
R12479 gnd.n5539 gnd.n1554 0.152939
R12480 gnd.n5539 gnd.n5538 0.152939
R12481 gnd.n1575 gnd.n1574 0.152939
R12482 gnd.n1576 gnd.n1575 0.152939
R12483 gnd.n1577 gnd.n1576 0.152939
R12484 gnd.n1578 gnd.n1577 0.152939
R12485 gnd.n1599 gnd.n1578 0.152939
R12486 gnd.n1600 gnd.n1599 0.152939
R12487 gnd.n1601 gnd.n1600 0.152939
R12488 gnd.n1602 gnd.n1601 0.152939
R12489 gnd.n1603 gnd.n1602 0.152939
R12490 gnd.n1603 gnd.n543 0.152939
R12491 gnd.n6739 gnd.n543 0.152939
R12492 gnd.n6740 gnd.n6739 0.152939
R12493 gnd.n6741 gnd.n6740 0.152939
R12494 gnd.n6742 gnd.n6741 0.152939
R12495 gnd.n6742 gnd.n77 0.152939
R12496 gnd.n6892 gnd.n77 0.152939
R12497 gnd.n6723 gnd.n561 0.152939
R12498 gnd.n4234 gnd.n4230 0.152939
R12499 gnd.n4235 gnd.n4234 0.152939
R12500 gnd.n4236 gnd.n4235 0.152939
R12501 gnd.n4236 gnd.n2152 0.152939
R12502 gnd.n4242 gnd.n2152 0.152939
R12503 gnd.n4243 gnd.n4242 0.152939
R12504 gnd.n4244 gnd.n4243 0.152939
R12505 gnd.n4245 gnd.n4244 0.152939
R12506 gnd.n4246 gnd.n4245 0.152939
R12507 gnd.n4246 gnd.n2134 0.152939
R12508 gnd.n4547 gnd.n2134 0.152939
R12509 gnd.n4548 gnd.n4547 0.152939
R12510 gnd.n4549 gnd.n4548 0.152939
R12511 gnd.n4549 gnd.n2130 0.152939
R12512 gnd.n4555 gnd.n2130 0.152939
R12513 gnd.n4556 gnd.n4555 0.152939
R12514 gnd.n4557 gnd.n4556 0.152939
R12515 gnd.n4558 gnd.n4557 0.152939
R12516 gnd.n4559 gnd.n4558 0.152939
R12517 gnd.n4560 gnd.n4559 0.152939
R12518 gnd.n4560 gnd.n2100 0.152939
R12519 gnd.n4583 gnd.n2100 0.152939
R12520 gnd.n4584 gnd.n4583 0.152939
R12521 gnd.n4585 gnd.n4584 0.152939
R12522 gnd.n4585 gnd.n2086 0.152939
R12523 gnd.n4599 gnd.n2086 0.152939
R12524 gnd.n4600 gnd.n4599 0.152939
R12525 gnd.n4601 gnd.n4600 0.152939
R12526 gnd.n4601 gnd.n2070 0.152939
R12527 gnd.n4632 gnd.n2070 0.152939
R12528 gnd.n4633 gnd.n4632 0.152939
R12529 gnd.n4634 gnd.n4633 0.152939
R12530 gnd.n4635 gnd.n4634 0.152939
R12531 gnd.n4636 gnd.n4635 0.152939
R12532 gnd.n4638 gnd.n4636 0.152939
R12533 gnd.n4638 gnd.n4637 0.152939
R12534 gnd.n4637 gnd.n1284 0.152939
R12535 gnd.n1285 gnd.n1284 0.152939
R12536 gnd.n1286 gnd.n1285 0.152939
R12537 gnd.n2032 gnd.n1286 0.152939
R12538 gnd.n2033 gnd.n2032 0.152939
R12539 gnd.n4799 gnd.n2033 0.152939
R12540 gnd.n4800 gnd.n4799 0.152939
R12541 gnd.n4801 gnd.n4800 0.152939
R12542 gnd.n4802 gnd.n4801 0.152939
R12543 gnd.n4802 gnd.n2009 0.152939
R12544 gnd.n4831 gnd.n2009 0.152939
R12545 gnd.n4832 gnd.n4831 0.152939
R12546 gnd.n4833 gnd.n4832 0.152939
R12547 gnd.n4833 gnd.n1985 0.152939
R12548 gnd.n4870 gnd.n1985 0.152939
R12549 gnd.n4871 gnd.n4870 0.152939
R12550 gnd.n4872 gnd.n4871 0.152939
R12551 gnd.n4872 gnd.n1959 0.152939
R12552 gnd.n4910 gnd.n1959 0.152939
R12553 gnd.n4911 gnd.n4910 0.152939
R12554 gnd.n4912 gnd.n4911 0.152939
R12555 gnd.n4913 gnd.n4912 0.152939
R12556 gnd.n4913 gnd.n1932 0.152939
R12557 gnd.n4956 gnd.n1932 0.152939
R12558 gnd.n4957 gnd.n4956 0.152939
R12559 gnd.n4958 gnd.n4957 0.152939
R12560 gnd.n4959 gnd.n4958 0.152939
R12561 gnd.n4959 gnd.n1910 0.152939
R12562 gnd.n5009 gnd.n1910 0.152939
R12563 gnd.n5010 gnd.n5009 0.152939
R12564 gnd.n5011 gnd.n5010 0.152939
R12565 gnd.n5012 gnd.n5011 0.152939
R12566 gnd.n5012 gnd.n1884 0.152939
R12567 gnd.n5045 gnd.n1884 0.152939
R12568 gnd.n5046 gnd.n5045 0.152939
R12569 gnd.n5047 gnd.n5046 0.152939
R12570 gnd.n5047 gnd.n1858 0.152939
R12571 gnd.n5089 gnd.n1858 0.152939
R12572 gnd.n5090 gnd.n5089 0.152939
R12573 gnd.n5091 gnd.n5090 0.152939
R12574 gnd.n5092 gnd.n5091 0.152939
R12575 gnd.n5092 gnd.n1835 0.152939
R12576 gnd.n5148 gnd.n1835 0.152939
R12577 gnd.n5149 gnd.n5148 0.152939
R12578 gnd.n5150 gnd.n5149 0.152939
R12579 gnd.n5150 gnd.n1813 0.152939
R12580 gnd.n5178 gnd.n1813 0.152939
R12581 gnd.n5179 gnd.n5178 0.152939
R12582 gnd.n5180 gnd.n5179 0.152939
R12583 gnd.n5180 gnd.n1796 0.152939
R12584 gnd.n5207 gnd.n1796 0.152939
R12585 gnd.n5208 gnd.n5207 0.152939
R12586 gnd.n5209 gnd.n5208 0.152939
R12587 gnd.n5209 gnd.n1705 0.152939
R12588 gnd.n5354 gnd.n1705 0.152939
R12589 gnd.n5355 gnd.n5354 0.152939
R12590 gnd.n5356 gnd.n5355 0.152939
R12591 gnd.n5356 gnd.n1692 0.152939
R12592 gnd.n5370 gnd.n1692 0.152939
R12593 gnd.n5371 gnd.n5370 0.152939
R12594 gnd.n5372 gnd.n5371 0.152939
R12595 gnd.n5372 gnd.n1679 0.152939
R12596 gnd.n5386 gnd.n1679 0.152939
R12597 gnd.n5387 gnd.n5386 0.152939
R12598 gnd.n5388 gnd.n5387 0.152939
R12599 gnd.n5390 gnd.n5388 0.152939
R12600 gnd.n5390 gnd.n5389 0.152939
R12601 gnd.n5389 gnd.n1666 0.152939
R12602 gnd.n5407 gnd.n1666 0.152939
R12603 gnd.n5408 gnd.n5407 0.152939
R12604 gnd.n5409 gnd.n5408 0.152939
R12605 gnd.n5410 gnd.n5409 0.152939
R12606 gnd.n5411 gnd.n5410 0.152939
R12607 gnd.n5413 gnd.n5411 0.152939
R12608 gnd.n5414 gnd.n5413 0.152939
R12609 gnd.n5416 gnd.n5414 0.152939
R12610 gnd.n5416 gnd.n5415 0.152939
R12611 gnd.n5415 gnd.n1630 0.152939
R12612 gnd.n5476 gnd.n1630 0.152939
R12613 gnd.n5477 gnd.n5476 0.152939
R12614 gnd.n5478 gnd.n5477 0.152939
R12615 gnd.n5478 gnd.n1626 0.152939
R12616 gnd.n5484 gnd.n1626 0.152939
R12617 gnd.n5485 gnd.n5484 0.152939
R12618 gnd.n5486 gnd.n5485 0.152939
R12619 gnd.n5487 gnd.n5486 0.152939
R12620 gnd.n5488 gnd.n5487 0.152939
R12621 gnd.n5490 gnd.n5488 0.152939
R12622 gnd.n5490 gnd.n5489 0.152939
R12623 gnd.n5489 gnd.n560 0.152939
R12624 gnd.n561 gnd.n560 0.152939
R12625 gnd.n3913 gnd.n3857 0.152939
R12626 gnd.n3858 gnd.n3857 0.152939
R12627 gnd.n3859 gnd.n3858 0.152939
R12628 gnd.n3860 gnd.n3859 0.152939
R12629 gnd.n3861 gnd.n3860 0.152939
R12630 gnd.n3862 gnd.n3861 0.152939
R12631 gnd.n3863 gnd.n3862 0.152939
R12632 gnd.n3864 gnd.n3863 0.152939
R12633 gnd.n3865 gnd.n3864 0.152939
R12634 gnd.n3866 gnd.n3865 0.152939
R12635 gnd.n3867 gnd.n3866 0.152939
R12636 gnd.n3868 gnd.n3867 0.152939
R12637 gnd.n3869 gnd.n3868 0.152939
R12638 gnd.n3870 gnd.n3869 0.152939
R12639 gnd.n3871 gnd.n3870 0.152939
R12640 gnd.n3872 gnd.n3871 0.152939
R12641 gnd.n3873 gnd.n3872 0.152939
R12642 gnd.n3874 gnd.n3873 0.152939
R12643 gnd.n3875 gnd.n3874 0.152939
R12644 gnd.n3876 gnd.n3875 0.152939
R12645 gnd.n3952 gnd.n3838 0.152939
R12646 gnd.n3839 gnd.n3838 0.152939
R12647 gnd.n3840 gnd.n3839 0.152939
R12648 gnd.n3841 gnd.n3840 0.152939
R12649 gnd.n3842 gnd.n3841 0.152939
R12650 gnd.n3843 gnd.n3842 0.152939
R12651 gnd.n3844 gnd.n3843 0.152939
R12652 gnd.n3845 gnd.n3844 0.152939
R12653 gnd.n3846 gnd.n3845 0.152939
R12654 gnd.n3847 gnd.n3846 0.152939
R12655 gnd.n3848 gnd.n3847 0.152939
R12656 gnd.n3849 gnd.n3848 0.152939
R12657 gnd.n3850 gnd.n3849 0.152939
R12658 gnd.n3851 gnd.n3850 0.152939
R12659 gnd.n3852 gnd.n3851 0.152939
R12660 gnd.n3917 gnd.n3852 0.152939
R12661 gnd.n3917 gnd.n3916 0.152939
R12662 gnd.n3916 gnd.n3915 0.152939
R12663 gnd.n1059 gnd.n1058 0.152939
R12664 gnd.n1078 gnd.n1059 0.152939
R12665 gnd.n1079 gnd.n1078 0.152939
R12666 gnd.n1080 gnd.n1079 0.152939
R12667 gnd.n1081 gnd.n1080 0.152939
R12668 gnd.n1098 gnd.n1081 0.152939
R12669 gnd.n1099 gnd.n1098 0.152939
R12670 gnd.n1100 gnd.n1099 0.152939
R12671 gnd.n1101 gnd.n1100 0.152939
R12672 gnd.n1118 gnd.n1101 0.152939
R12673 gnd.n1119 gnd.n1118 0.152939
R12674 gnd.n1120 gnd.n1119 0.152939
R12675 gnd.n1121 gnd.n1120 0.152939
R12676 gnd.n1139 gnd.n1121 0.152939
R12677 gnd.n1140 gnd.n1139 0.152939
R12678 gnd.n5960 gnd.n1140 0.152939
R12679 gnd.n5959 gnd.n1141 0.152939
R12680 gnd.n1185 gnd.n1141 0.152939
R12681 gnd.n1186 gnd.n1185 0.152939
R12682 gnd.n1187 gnd.n1186 0.152939
R12683 gnd.n1188 gnd.n1187 0.152939
R12684 gnd.n1189 gnd.n1188 0.152939
R12685 gnd.n1190 gnd.n1189 0.152939
R12686 gnd.n1191 gnd.n1190 0.152939
R12687 gnd.n1192 gnd.n1191 0.152939
R12688 gnd.n1193 gnd.n1192 0.152939
R12689 gnd.n1194 gnd.n1193 0.152939
R12690 gnd.n1195 gnd.n1194 0.152939
R12691 gnd.n1196 gnd.n1195 0.152939
R12692 gnd.n1197 gnd.n1196 0.152939
R12693 gnd.n1198 gnd.n1197 0.152939
R12694 gnd.n1199 gnd.n1198 0.152939
R12695 gnd.n1200 gnd.n1199 0.152939
R12696 gnd.n1203 gnd.n1200 0.152939
R12697 gnd.n1204 gnd.n1203 0.152939
R12698 gnd.n1205 gnd.n1204 0.152939
R12699 gnd.n1206 gnd.n1205 0.152939
R12700 gnd.n1207 gnd.n1206 0.152939
R12701 gnd.n1208 gnd.n1207 0.152939
R12702 gnd.n1209 gnd.n1208 0.152939
R12703 gnd.n1210 gnd.n1209 0.152939
R12704 gnd.n4448 gnd.n4447 0.152939
R12705 gnd.n4455 gnd.n4448 0.152939
R12706 gnd.n4456 gnd.n4455 0.152939
R12707 gnd.n4457 gnd.n4456 0.152939
R12708 gnd.n4457 gnd.n4445 0.152939
R12709 gnd.n4465 gnd.n4445 0.152939
R12710 gnd.n4466 gnd.n4465 0.152939
R12711 gnd.n4467 gnd.n4466 0.152939
R12712 gnd.n4467 gnd.n4440 0.152939
R12713 gnd.n4474 gnd.n4440 0.152939
R12714 gnd.n4475 gnd.n4474 0.152939
R12715 gnd.n4476 gnd.n4475 0.152939
R12716 gnd.n4476 gnd.n4438 0.152939
R12717 gnd.n4484 gnd.n4438 0.152939
R12718 gnd.n4485 gnd.n4484 0.152939
R12719 gnd.n4486 gnd.n4485 0.152939
R12720 gnd.n4486 gnd.n4436 0.152939
R12721 gnd.n4494 gnd.n4436 0.152939
R12722 gnd.n4495 gnd.n4494 0.152939
R12723 gnd.n4496 gnd.n4495 0.152939
R12724 gnd.n4496 gnd.n4434 0.152939
R12725 gnd.n4504 gnd.n4434 0.152939
R12726 gnd.n4505 gnd.n4504 0.152939
R12727 gnd.n4506 gnd.n4505 0.152939
R12728 gnd.n4506 gnd.n4432 0.152939
R12729 gnd.n4514 gnd.n4432 0.152939
R12730 gnd.n4515 gnd.n4514 0.152939
R12731 gnd.n4516 gnd.n4515 0.152939
R12732 gnd.n4516 gnd.n4427 0.152939
R12733 gnd.n4522 gnd.n4427 0.152939
R12734 gnd.n3776 gnd.n3775 0.152939
R12735 gnd.n3777 gnd.n3776 0.152939
R12736 gnd.n3778 gnd.n3777 0.152939
R12737 gnd.n3779 gnd.n3778 0.152939
R12738 gnd.n3780 gnd.n3779 0.152939
R12739 gnd.n3781 gnd.n3780 0.152939
R12740 gnd.n3782 gnd.n3781 0.152939
R12741 gnd.n3783 gnd.n3782 0.152939
R12742 gnd.n3784 gnd.n3783 0.152939
R12743 gnd.n3785 gnd.n3784 0.152939
R12744 gnd.n3786 gnd.n3785 0.152939
R12745 gnd.n3787 gnd.n3786 0.152939
R12746 gnd.n3788 gnd.n3787 0.152939
R12747 gnd.n3789 gnd.n3788 0.152939
R12748 gnd.n3790 gnd.n3789 0.152939
R12749 gnd.n3791 gnd.n3790 0.152939
R12750 gnd.n3792 gnd.n3791 0.152939
R12751 gnd.n3795 gnd.n3792 0.152939
R12752 gnd.n3796 gnd.n3795 0.152939
R12753 gnd.n3797 gnd.n3796 0.152939
R12754 gnd.n3798 gnd.n3797 0.152939
R12755 gnd.n3799 gnd.n3798 0.152939
R12756 gnd.n3800 gnd.n3799 0.152939
R12757 gnd.n3801 gnd.n3800 0.152939
R12758 gnd.n3802 gnd.n3801 0.152939
R12759 gnd.n3803 gnd.n3802 0.152939
R12760 gnd.n3804 gnd.n3803 0.152939
R12761 gnd.n3805 gnd.n3804 0.152939
R12762 gnd.n3806 gnd.n3805 0.152939
R12763 gnd.n3807 gnd.n3806 0.152939
R12764 gnd.n3808 gnd.n3807 0.152939
R12765 gnd.n3809 gnd.n3808 0.152939
R12766 gnd.n3810 gnd.n3809 0.152939
R12767 gnd.n3811 gnd.n3810 0.152939
R12768 gnd.n3812 gnd.n3811 0.152939
R12769 gnd.n3813 gnd.n3812 0.152939
R12770 gnd.n3814 gnd.n3813 0.152939
R12771 gnd.n3817 gnd.n3814 0.152939
R12772 gnd.n3818 gnd.n3817 0.152939
R12773 gnd.n3819 gnd.n3818 0.152939
R12774 gnd.n3820 gnd.n3819 0.152939
R12775 gnd.n3821 gnd.n3820 0.152939
R12776 gnd.n3822 gnd.n3821 0.152939
R12777 gnd.n3823 gnd.n3822 0.152939
R12778 gnd.n3824 gnd.n3823 0.152939
R12779 gnd.n3825 gnd.n3824 0.152939
R12780 gnd.n3826 gnd.n3825 0.152939
R12781 gnd.n3827 gnd.n3826 0.152939
R12782 gnd.n3828 gnd.n3827 0.152939
R12783 gnd.n3829 gnd.n3828 0.152939
R12784 gnd.n3830 gnd.n3829 0.152939
R12785 gnd.n3831 gnd.n3830 0.152939
R12786 gnd.n3832 gnd.n3831 0.152939
R12787 gnd.n3833 gnd.n3832 0.152939
R12788 gnd.n3834 gnd.n3833 0.152939
R12789 gnd.n3835 gnd.n3834 0.152939
R12790 gnd.n3955 gnd.n3835 0.152939
R12791 gnd.n3955 gnd.n3954 0.152939
R12792 gnd.n4084 gnd.n2257 0.152939
R12793 gnd.n4085 gnd.n4084 0.152939
R12794 gnd.n4086 gnd.n4085 0.152939
R12795 gnd.n4086 gnd.n2238 0.152939
R12796 gnd.n4104 gnd.n2238 0.152939
R12797 gnd.n4105 gnd.n4104 0.152939
R12798 gnd.n4106 gnd.n4105 0.152939
R12799 gnd.n4106 gnd.n2221 0.152939
R12800 gnd.n4124 gnd.n2221 0.152939
R12801 gnd.n4125 gnd.n4124 0.152939
R12802 gnd.n4126 gnd.n4125 0.152939
R12803 gnd.n4126 gnd.n2202 0.152939
R12804 gnd.n4144 gnd.n2202 0.152939
R12805 gnd.n4145 gnd.n4144 0.152939
R12806 gnd.n4146 gnd.n4145 0.152939
R12807 gnd.n4146 gnd.n1058 0.152939
R12808 gnd.n6184 gnd.n881 0.152939
R12809 gnd.n886 gnd.n881 0.152939
R12810 gnd.n887 gnd.n886 0.152939
R12811 gnd.n888 gnd.n887 0.152939
R12812 gnd.n893 gnd.n888 0.152939
R12813 gnd.n894 gnd.n893 0.152939
R12814 gnd.n895 gnd.n894 0.152939
R12815 gnd.n896 gnd.n895 0.152939
R12816 gnd.n901 gnd.n896 0.152939
R12817 gnd.n902 gnd.n901 0.152939
R12818 gnd.n903 gnd.n902 0.152939
R12819 gnd.n904 gnd.n903 0.152939
R12820 gnd.n909 gnd.n904 0.152939
R12821 gnd.n910 gnd.n909 0.152939
R12822 gnd.n911 gnd.n910 0.152939
R12823 gnd.n912 gnd.n911 0.152939
R12824 gnd.n917 gnd.n912 0.152939
R12825 gnd.n918 gnd.n917 0.152939
R12826 gnd.n919 gnd.n918 0.152939
R12827 gnd.n920 gnd.n919 0.152939
R12828 gnd.n925 gnd.n920 0.152939
R12829 gnd.n926 gnd.n925 0.152939
R12830 gnd.n927 gnd.n926 0.152939
R12831 gnd.n928 gnd.n927 0.152939
R12832 gnd.n933 gnd.n928 0.152939
R12833 gnd.n934 gnd.n933 0.152939
R12834 gnd.n935 gnd.n934 0.152939
R12835 gnd.n936 gnd.n935 0.152939
R12836 gnd.n941 gnd.n936 0.152939
R12837 gnd.n942 gnd.n941 0.152939
R12838 gnd.n943 gnd.n942 0.152939
R12839 gnd.n944 gnd.n943 0.152939
R12840 gnd.n949 gnd.n944 0.152939
R12841 gnd.n950 gnd.n949 0.152939
R12842 gnd.n951 gnd.n950 0.152939
R12843 gnd.n952 gnd.n951 0.152939
R12844 gnd.n957 gnd.n952 0.152939
R12845 gnd.n958 gnd.n957 0.152939
R12846 gnd.n959 gnd.n958 0.152939
R12847 gnd.n960 gnd.n959 0.152939
R12848 gnd.n965 gnd.n960 0.152939
R12849 gnd.n966 gnd.n965 0.152939
R12850 gnd.n967 gnd.n966 0.152939
R12851 gnd.n968 gnd.n967 0.152939
R12852 gnd.n973 gnd.n968 0.152939
R12853 gnd.n974 gnd.n973 0.152939
R12854 gnd.n975 gnd.n974 0.152939
R12855 gnd.n976 gnd.n975 0.152939
R12856 gnd.n981 gnd.n976 0.152939
R12857 gnd.n982 gnd.n981 0.152939
R12858 gnd.n983 gnd.n982 0.152939
R12859 gnd.n984 gnd.n983 0.152939
R12860 gnd.n989 gnd.n984 0.152939
R12861 gnd.n990 gnd.n989 0.152939
R12862 gnd.n991 gnd.n990 0.152939
R12863 gnd.n992 gnd.n991 0.152939
R12864 gnd.n997 gnd.n992 0.152939
R12865 gnd.n998 gnd.n997 0.152939
R12866 gnd.n999 gnd.n998 0.152939
R12867 gnd.n1000 gnd.n999 0.152939
R12868 gnd.n1005 gnd.n1000 0.152939
R12869 gnd.n1006 gnd.n1005 0.152939
R12870 gnd.n1007 gnd.n1006 0.152939
R12871 gnd.n1008 gnd.n1007 0.152939
R12872 gnd.n1013 gnd.n1008 0.152939
R12873 gnd.n1014 gnd.n1013 0.152939
R12874 gnd.n1015 gnd.n1014 0.152939
R12875 gnd.n1016 gnd.n1015 0.152939
R12876 gnd.n1021 gnd.n1016 0.152939
R12877 gnd.n1022 gnd.n1021 0.152939
R12878 gnd.n1023 gnd.n1022 0.152939
R12879 gnd.n1024 gnd.n1023 0.152939
R12880 gnd.n1029 gnd.n1024 0.152939
R12881 gnd.n1030 gnd.n1029 0.152939
R12882 gnd.n1031 gnd.n1030 0.152939
R12883 gnd.n1032 gnd.n1031 0.152939
R12884 gnd.n1037 gnd.n1032 0.152939
R12885 gnd.n1038 gnd.n1037 0.152939
R12886 gnd.n1039 gnd.n1038 0.152939
R12887 gnd.n1040 gnd.n1039 0.152939
R12888 gnd.n1045 gnd.n1040 0.152939
R12889 gnd.n1046 gnd.n1045 0.152939
R12890 gnd.n1047 gnd.n1046 0.152939
R12891 gnd.n1048 gnd.n1047 0.152939
R12892 gnd.n4591 gnd.n2093 0.152939
R12893 gnd.n4592 gnd.n4591 0.152939
R12894 gnd.n4593 gnd.n4592 0.152939
R12895 gnd.n4593 gnd.n2078 0.152939
R12896 gnd.n4607 gnd.n2078 0.152939
R12897 gnd.n4608 gnd.n4607 0.152939
R12898 gnd.n4626 gnd.n4608 0.152939
R12899 gnd.n4626 gnd.n4625 0.152939
R12900 gnd.n4625 gnd.n4624 0.152939
R12901 gnd.n4624 gnd.n4609 0.152939
R12902 gnd.n4620 gnd.n4609 0.152939
R12903 gnd.n4620 gnd.n4619 0.152939
R12904 gnd.n4619 gnd.n4618 0.152939
R12905 gnd.n4618 gnd.n4613 0.152939
R12906 gnd.n4613 gnd.n1294 0.152939
R12907 gnd.n5822 gnd.n1294 0.152939
R12908 gnd.n5822 gnd.n5821 0.152939
R12909 gnd.n5821 gnd.n5820 0.152939
R12910 gnd.n5820 gnd.n1295 0.152939
R12911 gnd.n5816 gnd.n1295 0.152939
R12912 gnd.n5816 gnd.n5815 0.152939
R12913 gnd.n5815 gnd.n5814 0.152939
R12914 gnd.n5814 gnd.n1300 0.152939
R12915 gnd.n5810 gnd.n1300 0.152939
R12916 gnd.n5810 gnd.n5809 0.152939
R12917 gnd.n5809 gnd.n5808 0.152939
R12918 gnd.n5808 gnd.n1305 0.152939
R12919 gnd.n5804 gnd.n1305 0.152939
R12920 gnd.n5804 gnd.n5803 0.152939
R12921 gnd.n5803 gnd.n5802 0.152939
R12922 gnd.n5802 gnd.n1310 0.152939
R12923 gnd.n5798 gnd.n1310 0.152939
R12924 gnd.n5798 gnd.n5797 0.152939
R12925 gnd.n5797 gnd.n5796 0.152939
R12926 gnd.n5796 gnd.n1315 0.152939
R12927 gnd.n5792 gnd.n1315 0.152939
R12928 gnd.n5792 gnd.n5791 0.152939
R12929 gnd.n5791 gnd.n5790 0.152939
R12930 gnd.n5790 gnd.n1320 0.152939
R12931 gnd.n5786 gnd.n1320 0.152939
R12932 gnd.n5786 gnd.n5785 0.152939
R12933 gnd.n5785 gnd.n5784 0.152939
R12934 gnd.n5784 gnd.n1325 0.152939
R12935 gnd.n5780 gnd.n1325 0.152939
R12936 gnd.n5780 gnd.n5779 0.152939
R12937 gnd.n5779 gnd.n5778 0.152939
R12938 gnd.n5778 gnd.n1330 0.152939
R12939 gnd.n5774 gnd.n1330 0.152939
R12940 gnd.n5774 gnd.n5773 0.152939
R12941 gnd.n5773 gnd.n5772 0.152939
R12942 gnd.n5772 gnd.n1335 0.152939
R12943 gnd.n5768 gnd.n1335 0.152939
R12944 gnd.n5768 gnd.n5767 0.152939
R12945 gnd.n5767 gnd.n5766 0.152939
R12946 gnd.n5766 gnd.n1340 0.152939
R12947 gnd.n5762 gnd.n1340 0.152939
R12948 gnd.n5762 gnd.n5761 0.152939
R12949 gnd.n5761 gnd.n5760 0.152939
R12950 gnd.n5760 gnd.n1345 0.152939
R12951 gnd.n5756 gnd.n1345 0.152939
R12952 gnd.n5756 gnd.n5755 0.152939
R12953 gnd.n5755 gnd.n5754 0.152939
R12954 gnd.n5754 gnd.n1350 0.152939
R12955 gnd.n5750 gnd.n1350 0.152939
R12956 gnd.n5750 gnd.n5749 0.152939
R12957 gnd.n5749 gnd.n5748 0.152939
R12958 gnd.n5748 gnd.n1355 0.152939
R12959 gnd.n5744 gnd.n1355 0.152939
R12960 gnd.n5744 gnd.n5743 0.152939
R12961 gnd.n5743 gnd.n5742 0.152939
R12962 gnd.n5742 gnd.n1360 0.152939
R12963 gnd.n5738 gnd.n1360 0.152939
R12964 gnd.n5738 gnd.n5737 0.152939
R12965 gnd.n5737 gnd.n5736 0.152939
R12966 gnd.n5736 gnd.n1365 0.152939
R12967 gnd.n5732 gnd.n1365 0.152939
R12968 gnd.n5732 gnd.n5731 0.152939
R12969 gnd.n5731 gnd.n5730 0.152939
R12970 gnd.n5730 gnd.n1370 0.152939
R12971 gnd.n5726 gnd.n1370 0.152939
R12972 gnd.n5726 gnd.n5725 0.152939
R12973 gnd.n5725 gnd.n5724 0.152939
R12974 gnd.n3878 gnd.n2161 0.152939
R12975 gnd.n4201 gnd.n2161 0.152939
R12976 gnd.n4202 gnd.n4201 0.152939
R12977 gnd.n4203 gnd.n4202 0.152939
R12978 gnd.n4203 gnd.n2157 0.152939
R12979 gnd.n4222 gnd.n2157 0.152939
R12980 gnd.n4222 gnd.n4221 0.152939
R12981 gnd.n4221 gnd.n4220 0.152939
R12982 gnd.n4220 gnd.n2146 0.152939
R12983 gnd.n4255 gnd.n2146 0.152939
R12984 gnd.n4256 gnd.n4255 0.152939
R12985 gnd.n4257 gnd.n4256 0.152939
R12986 gnd.n4257 gnd.n2140 0.152939
R12987 gnd.n4539 gnd.n2140 0.152939
R12988 gnd.n4539 gnd.n4538 0.152939
R12989 gnd.n4538 gnd.n4537 0.152939
R12990 gnd.n4537 gnd.n2141 0.152939
R12991 gnd.n4533 gnd.n2141 0.152939
R12992 gnd.n4533 gnd.n4532 0.152939
R12993 gnd.n4532 gnd.n2120 0.152939
R12994 gnd.n4277 gnd.n4276 0.152939
R12995 gnd.n4304 gnd.n4276 0.152939
R12996 gnd.n4305 gnd.n4304 0.152939
R12997 gnd.n4306 gnd.n4305 0.152939
R12998 gnd.n4306 gnd.n4272 0.152939
R12999 gnd.n4425 gnd.n4272 0.152939
R13000 gnd.n4295 gnd.n4294 0.152939
R13001 gnd.n4294 gnd.n4293 0.152939
R13002 gnd.n4293 gnd.n4279 0.152939
R13003 gnd.n4289 gnd.n4279 0.152939
R13004 gnd.n4289 gnd.n4288 0.152939
R13005 gnd.n4288 gnd.n4287 0.152939
R13006 gnd.n4287 gnd.n4283 0.152939
R13007 gnd.n4283 gnd.n2061 0.152939
R13008 gnd.n4649 gnd.n2061 0.152939
R13009 gnd.n4650 gnd.n4649 0.152939
R13010 gnd.n4651 gnd.n4650 0.152939
R13011 gnd.n4651 gnd.n2057 0.152939
R13012 gnd.n4657 gnd.n2057 0.152939
R13013 gnd.n4658 gnd.n4657 0.152939
R13014 gnd.n4668 gnd.n4658 0.152939
R13015 gnd.n4668 gnd.n4667 0.152939
R13016 gnd.n4667 gnd.n4666 0.152939
R13017 gnd.n4666 gnd.n4659 0.152939
R13018 gnd.n4662 gnd.n4659 0.152939
R13019 gnd.n4662 gnd.n2023 0.152939
R13020 gnd.n4809 gnd.n2023 0.152939
R13021 gnd.n4810 gnd.n4809 0.152939
R13022 gnd.n4814 gnd.n4810 0.152939
R13023 gnd.n4814 gnd.n4813 0.152939
R13024 gnd.n4813 gnd.n4812 0.152939
R13025 gnd.n4812 gnd.n2002 0.152939
R13026 gnd.n4840 gnd.n2002 0.152939
R13027 gnd.n4841 gnd.n4840 0.152939
R13028 gnd.n4848 gnd.n4841 0.152939
R13029 gnd.n4848 gnd.n4847 0.152939
R13030 gnd.n4847 gnd.n4846 0.152939
R13031 gnd.n4846 gnd.n4842 0.152939
R13032 gnd.n4842 gnd.n1952 0.152939
R13033 gnd.n4920 gnd.n1952 0.152939
R13034 gnd.n4921 gnd.n4920 0.152939
R13035 gnd.n4923 gnd.n4921 0.152939
R13036 gnd.n4923 gnd.n4922 0.152939
R13037 gnd.n4922 gnd.n1925 0.152939
R13038 gnd.n4966 gnd.n1925 0.152939
R13039 gnd.n4967 gnd.n4966 0.152939
R13040 gnd.n4994 gnd.n4967 0.152939
R13041 gnd.n4994 gnd.n4993 0.152939
R13042 gnd.n4993 gnd.n4992 0.152939
R13043 gnd.n4992 gnd.n4968 0.152939
R13044 gnd.n4988 gnd.n4968 0.152939
R13045 gnd.n4988 gnd.n4987 0.152939
R13046 gnd.n4987 gnd.n4986 0.152939
R13047 gnd.n4986 gnd.n4974 0.152939
R13048 gnd.n4982 gnd.n4974 0.152939
R13049 gnd.n4982 gnd.n4981 0.152939
R13050 gnd.n4981 gnd.n4980 0.152939
R13051 gnd.n4980 gnd.n1850 0.152939
R13052 gnd.n5099 gnd.n1850 0.152939
R13053 gnd.n5100 gnd.n5099 0.152939
R13054 gnd.n5134 gnd.n5100 0.152939
R13055 gnd.n5134 gnd.n5133 0.152939
R13056 gnd.n5133 gnd.n5132 0.152939
R13057 gnd.n5132 gnd.n5101 0.152939
R13058 gnd.n5128 gnd.n5101 0.152939
R13059 gnd.n5128 gnd.n5127 0.152939
R13060 gnd.n5127 gnd.n5126 0.152939
R13061 gnd.n5126 gnd.n5107 0.152939
R13062 gnd.n5122 gnd.n5107 0.152939
R13063 gnd.n5122 gnd.n5121 0.152939
R13064 gnd.n5121 gnd.n5120 0.152939
R13065 gnd.n5120 gnd.n5111 0.152939
R13066 gnd.n5116 gnd.n5111 0.152939
R13067 gnd.n5116 gnd.n5115 0.152939
R13068 gnd.n5115 gnd.n1697 0.152939
R13069 gnd.n5362 gnd.n1697 0.152939
R13070 gnd.n5363 gnd.n5362 0.152939
R13071 gnd.n5364 gnd.n5363 0.152939
R13072 gnd.n5364 gnd.n1684 0.152939
R13073 gnd.n5378 gnd.n1684 0.152939
R13074 gnd.n5379 gnd.n5378 0.152939
R13075 gnd.n5380 gnd.n5379 0.152939
R13076 gnd.n5380 gnd.n1672 0.152939
R13077 gnd.n5397 gnd.n1672 0.152939
R13078 gnd.n5398 gnd.n5397 0.152939
R13079 gnd.n5399 gnd.n5398 0.152939
R13080 gnd.n5399 gnd.n1384 0.152939
R13081 gnd.n5718 gnd.n1384 0.152939
R13082 gnd.n5717 gnd.n1385 0.152939
R13083 gnd.n5713 gnd.n1385 0.152939
R13084 gnd.n5713 gnd.n5712 0.152939
R13085 gnd.n5712 gnd.n5711 0.152939
R13086 gnd.n5711 gnd.n1389 0.152939
R13087 gnd.n5707 gnd.n1389 0.152939
R13088 gnd.n5467 gnd.n5433 0.152939
R13089 gnd.n5467 gnd.n5466 0.152939
R13090 gnd.n5466 gnd.n5465 0.152939
R13091 gnd.n5465 gnd.n5434 0.152939
R13092 gnd.n5461 gnd.n5434 0.152939
R13093 gnd.n5461 gnd.n5460 0.152939
R13094 gnd.n5460 gnd.n5459 0.152939
R13095 gnd.n5459 gnd.n5439 0.152939
R13096 gnd.n5455 gnd.n5439 0.152939
R13097 gnd.n5455 gnd.n5454 0.152939
R13098 gnd.n5454 gnd.n5453 0.152939
R13099 gnd.n5453 gnd.n533 0.152939
R13100 gnd.n6750 gnd.n533 0.152939
R13101 gnd.n6751 gnd.n6750 0.152939
R13102 gnd.n6752 gnd.n6751 0.152939
R13103 gnd.n6752 gnd.n514 0.152939
R13104 gnd.n6777 gnd.n514 0.152939
R13105 gnd.n6778 gnd.n6777 0.152939
R13106 gnd.n6779 gnd.n6778 0.152939
R13107 gnd.n6779 gnd.n63 0.152939
R13108 gnd.n6902 gnd.n6901 0.145814
R13109 gnd.n3879 gnd.n3876 0.145814
R13110 gnd.n3879 gnd.n3878 0.145814
R13111 gnd.n6902 gnd.n63 0.145814
R13112 gnd.n6723 gnd.n78 0.136171
R13113 gnd.n4230 gnd.n4229 0.136171
R13114 gnd.n4426 gnd.n4425 0.128549
R13115 gnd.n5707 gnd.n5706 0.128549
R13116 gnd.n2552 gnd.n0 0.127478
R13117 gnd.n3132 gnd.n3131 0.0767195
R13118 gnd.n3131 gnd.n3130 0.0767195
R13119 gnd.n4523 gnd.n4426 0.063
R13120 gnd.n5706 gnd.n1394 0.063
R13121 gnd.n1562 gnd.n1394 0.0538288
R13122 gnd.n6838 gnd.n493 0.0538288
R13123 gnd.n3953 gnd.n2267 0.0538288
R13124 gnd.n4524 gnd.n4523 0.0538288
R13125 gnd.n3699 gnd.n2314 0.0477147
R13126 gnd.n2895 gnd.n2783 0.0442063
R13127 gnd.n2896 gnd.n2895 0.0442063
R13128 gnd.n2897 gnd.n2896 0.0442063
R13129 gnd.n2897 gnd.n2772 0.0442063
R13130 gnd.n2911 gnd.n2772 0.0442063
R13131 gnd.n2912 gnd.n2911 0.0442063
R13132 gnd.n2913 gnd.n2912 0.0442063
R13133 gnd.n2913 gnd.n2759 0.0442063
R13134 gnd.n2957 gnd.n2759 0.0442063
R13135 gnd.n2958 gnd.n2957 0.0442063
R13136 gnd.n2960 gnd.n2693 0.0344674
R13137 gnd.n5528 gnd.n1562 0.0344674
R13138 gnd.n5528 gnd.n1564 0.0344674
R13139 gnd.n1588 gnd.n1564 0.0344674
R13140 gnd.n1589 gnd.n1588 0.0344674
R13141 gnd.n1590 gnd.n1589 0.0344674
R13142 gnd.n1591 gnd.n1590 0.0344674
R13143 gnd.n5445 gnd.n1591 0.0344674
R13144 gnd.n5445 gnd.n1611 0.0344674
R13145 gnd.n5502 gnd.n1611 0.0344674
R13146 gnd.n5502 gnd.n1612 0.0344674
R13147 gnd.n1612 gnd.n553 0.0344674
R13148 gnd.n554 gnd.n553 0.0344674
R13149 gnd.n555 gnd.n554 0.0344674
R13150 gnd.n556 gnd.n555 0.0344674
R13151 gnd.n556 gnd.n529 0.0344674
R13152 gnd.n529 gnd.n526 0.0344674
R13153 gnd.n527 gnd.n526 0.0344674
R13154 gnd.n6763 gnd.n527 0.0344674
R13155 gnd.n6763 gnd.n502 0.0344674
R13156 gnd.n6793 gnd.n502 0.0344674
R13157 gnd.n6794 gnd.n6793 0.0344674
R13158 gnd.n6794 gnd.n497 0.0344674
R13159 gnd.n497 gnd.n495 0.0344674
R13160 gnd.n6805 gnd.n495 0.0344674
R13161 gnd.n6806 gnd.n6805 0.0344674
R13162 gnd.n6806 gnd.n92 0.0344674
R13163 gnd.n93 gnd.n92 0.0344674
R13164 gnd.n94 gnd.n93 0.0344674
R13165 gnd.n6814 gnd.n94 0.0344674
R13166 gnd.n6814 gnd.n109 0.0344674
R13167 gnd.n110 gnd.n109 0.0344674
R13168 gnd.n111 gnd.n110 0.0344674
R13169 gnd.n6821 gnd.n111 0.0344674
R13170 gnd.n6821 gnd.n129 0.0344674
R13171 gnd.n130 gnd.n129 0.0344674
R13172 gnd.n131 gnd.n130 0.0344674
R13173 gnd.n6828 gnd.n131 0.0344674
R13174 gnd.n6828 gnd.n149 0.0344674
R13175 gnd.n150 gnd.n149 0.0344674
R13176 gnd.n151 gnd.n150 0.0344674
R13177 gnd.n167 gnd.n151 0.0344674
R13178 gnd.n6838 gnd.n167 0.0344674
R13179 gnd.n4078 gnd.n2267 0.0344674
R13180 gnd.n4078 gnd.n2270 0.0344674
R13181 gnd.n2270 gnd.n2269 0.0344674
R13182 gnd.n2269 gnd.n2250 0.0344674
R13183 gnd.n2250 gnd.n2248 0.0344674
R13184 gnd.n4095 gnd.n2248 0.0344674
R13185 gnd.n4096 gnd.n4095 0.0344674
R13186 gnd.n4096 gnd.n2232 0.0344674
R13187 gnd.n2232 gnd.n2230 0.0344674
R13188 gnd.n4115 gnd.n2230 0.0344674
R13189 gnd.n4116 gnd.n4115 0.0344674
R13190 gnd.n4116 gnd.n2214 0.0344674
R13191 gnd.n2214 gnd.n2212 0.0344674
R13192 gnd.n4135 gnd.n2212 0.0344674
R13193 gnd.n4136 gnd.n4135 0.0344674
R13194 gnd.n4136 gnd.n2196 0.0344674
R13195 gnd.n2196 gnd.n2194 0.0344674
R13196 gnd.n4156 gnd.n2194 0.0344674
R13197 gnd.n4157 gnd.n4156 0.0344674
R13198 gnd.n4157 gnd.n2180 0.0344674
R13199 gnd.n2180 gnd.n2176 0.0344674
R13200 gnd.n2177 gnd.n2176 0.0344674
R13201 gnd.n2178 gnd.n2177 0.0344674
R13202 gnd.n4180 gnd.n2178 0.0344674
R13203 gnd.n4181 gnd.n4180 0.0344674
R13204 gnd.n4181 gnd.n2159 0.0344674
R13205 gnd.n2159 gnd.n1068 0.0344674
R13206 gnd.n1069 gnd.n1068 0.0344674
R13207 gnd.n1070 gnd.n1069 0.0344674
R13208 gnd.n4212 gnd.n1070 0.0344674
R13209 gnd.n4212 gnd.n1089 0.0344674
R13210 gnd.n1090 gnd.n1089 0.0344674
R13211 gnd.n1091 gnd.n1090 0.0344674
R13212 gnd.n2144 gnd.n1091 0.0344674
R13213 gnd.n2144 gnd.n1108 0.0344674
R13214 gnd.n1109 gnd.n1108 0.0344674
R13215 gnd.n1110 gnd.n1109 0.0344674
R13216 gnd.n4266 gnd.n1110 0.0344674
R13217 gnd.n4266 gnd.n1129 0.0344674
R13218 gnd.n1130 gnd.n1129 0.0344674
R13219 gnd.n1131 gnd.n1130 0.0344674
R13220 gnd.n4524 gnd.n1131 0.0344674
R13221 gnd.n4421 gnd.n4271 0.0344674
R13222 gnd.n5705 gnd.n5704 0.0344674
R13223 gnd.n4575 gnd.n4574 0.029712
R13224 gnd.n5432 gnd.n5431 0.029712
R13225 gnd.n2980 gnd.n2979 0.0269946
R13226 gnd.n2982 gnd.n2981 0.0269946
R13227 gnd.n2688 gnd.n2686 0.0269946
R13228 gnd.n2992 gnd.n2990 0.0269946
R13229 gnd.n2991 gnd.n2667 0.0269946
R13230 gnd.n3011 gnd.n3010 0.0269946
R13231 gnd.n3013 gnd.n3012 0.0269946
R13232 gnd.n2662 gnd.n2661 0.0269946
R13233 gnd.n3023 gnd.n2657 0.0269946
R13234 gnd.n3022 gnd.n2659 0.0269946
R13235 gnd.n2658 gnd.n2640 0.0269946
R13236 gnd.n3043 gnd.n2641 0.0269946
R13237 gnd.n3042 gnd.n2642 0.0269946
R13238 gnd.n3076 gnd.n2617 0.0269946
R13239 gnd.n3078 gnd.n3077 0.0269946
R13240 gnd.n3079 gnd.n2564 0.0269946
R13241 gnd.n2612 gnd.n2565 0.0269946
R13242 gnd.n2614 gnd.n2566 0.0269946
R13243 gnd.n3089 gnd.n3088 0.0269946
R13244 gnd.n3091 gnd.n3090 0.0269946
R13245 gnd.n3092 gnd.n2586 0.0269946
R13246 gnd.n3094 gnd.n2587 0.0269946
R13247 gnd.n3097 gnd.n2588 0.0269946
R13248 gnd.n3100 gnd.n3099 0.0269946
R13249 gnd.n3102 gnd.n3101 0.0269946
R13250 gnd.n3167 gnd.n2487 0.0269946
R13251 gnd.n3169 gnd.n3168 0.0269946
R13252 gnd.n3178 gnd.n2480 0.0269946
R13253 gnd.n3180 gnd.n3179 0.0269946
R13254 gnd.n3181 gnd.n2478 0.0269946
R13255 gnd.n3188 gnd.n3184 0.0269946
R13256 gnd.n3187 gnd.n3186 0.0269946
R13257 gnd.n3185 gnd.n2457 0.0269946
R13258 gnd.n3210 gnd.n2458 0.0269946
R13259 gnd.n3209 gnd.n2459 0.0269946
R13260 gnd.n3252 gnd.n2432 0.0269946
R13261 gnd.n3254 gnd.n3253 0.0269946
R13262 gnd.n3263 gnd.n2425 0.0269946
R13263 gnd.n3265 gnd.n3264 0.0269946
R13264 gnd.n3266 gnd.n2423 0.0269946
R13265 gnd.n3273 gnd.n3269 0.0269946
R13266 gnd.n3272 gnd.n3271 0.0269946
R13267 gnd.n3270 gnd.n2402 0.0269946
R13268 gnd.n3295 gnd.n2403 0.0269946
R13269 gnd.n3294 gnd.n2404 0.0269946
R13270 gnd.n3341 gnd.n2378 0.0269946
R13271 gnd.n3343 gnd.n3342 0.0269946
R13272 gnd.n3353 gnd.n2371 0.0269946
R13273 gnd.n3612 gnd.n2369 0.0269946
R13274 gnd.n3617 gnd.n3615 0.0269946
R13275 gnd.n3616 gnd.n2350 0.0269946
R13276 gnd.n3641 gnd.n3640 0.0269946
R13277 gnd.n4420 gnd.n4314 0.0225788
R13278 gnd.n4417 gnd.n4416 0.0225788
R13279 gnd.n4413 gnd.n4317 0.0225788
R13280 gnd.n4412 gnd.n4323 0.0225788
R13281 gnd.n4409 gnd.n4408 0.0225788
R13282 gnd.n4405 gnd.n4329 0.0225788
R13283 gnd.n4404 gnd.n4333 0.0225788
R13284 gnd.n4401 gnd.n4400 0.0225788
R13285 gnd.n4397 gnd.n4337 0.0225788
R13286 gnd.n4396 gnd.n4343 0.0225788
R13287 gnd.n4393 gnd.n4392 0.0225788
R13288 gnd.n4389 gnd.n4349 0.0225788
R13289 gnd.n4388 gnd.n4353 0.0225788
R13290 gnd.n4385 gnd.n4384 0.0225788
R13291 gnd.n4381 gnd.n4357 0.0225788
R13292 gnd.n4380 gnd.n4363 0.0225788
R13293 gnd.n4377 gnd.n4376 0.0225788
R13294 gnd.n4368 gnd.n2121 0.0225788
R13295 gnd.n4574 gnd.n4573 0.0225788
R13296 gnd.n5701 gnd.n1395 0.0225788
R13297 gnd.n5700 gnd.n1399 0.0225788
R13298 gnd.n5697 gnd.n5696 0.0225788
R13299 gnd.n5693 gnd.n1404 0.0225788
R13300 gnd.n5692 gnd.n1408 0.0225788
R13301 gnd.n5689 gnd.n5688 0.0225788
R13302 gnd.n5685 gnd.n1412 0.0225788
R13303 gnd.n5684 gnd.n1416 0.0225788
R13304 gnd.n5681 gnd.n5680 0.0225788
R13305 gnd.n5677 gnd.n1420 0.0225788
R13306 gnd.n5676 gnd.n1424 0.0225788
R13307 gnd.n5673 gnd.n5672 0.0225788
R13308 gnd.n5669 gnd.n1428 0.0225788
R13309 gnd.n5668 gnd.n1432 0.0225788
R13310 gnd.n5665 gnd.n5664 0.0225788
R13311 gnd.n5661 gnd.n1436 0.0225788
R13312 gnd.n5660 gnd.n1442 0.0225788
R13313 gnd.n1637 gnd.n1445 0.0225788
R13314 gnd.n5431 gnd.n1636 0.0225788
R13315 gnd.n5432 gnd.n1375 0.0218415
R13316 gnd.n4576 gnd.n4575 0.0218415
R13317 gnd.n2960 gnd.n2959 0.0202011
R13318 gnd.n2959 gnd.n2958 0.0148637
R13319 gnd.n3610 gnd.n3354 0.0144266
R13320 gnd.n3611 gnd.n3610 0.0130679
R13321 gnd.n4421 gnd.n4420 0.0123886
R13322 gnd.n4417 gnd.n4314 0.0123886
R13323 gnd.n4416 gnd.n4317 0.0123886
R13324 gnd.n4413 gnd.n4412 0.0123886
R13325 gnd.n4409 gnd.n4323 0.0123886
R13326 gnd.n4408 gnd.n4329 0.0123886
R13327 gnd.n4405 gnd.n4404 0.0123886
R13328 gnd.n4401 gnd.n4333 0.0123886
R13329 gnd.n4400 gnd.n4337 0.0123886
R13330 gnd.n4397 gnd.n4396 0.0123886
R13331 gnd.n4393 gnd.n4343 0.0123886
R13332 gnd.n4392 gnd.n4349 0.0123886
R13333 gnd.n4389 gnd.n4388 0.0123886
R13334 gnd.n4385 gnd.n4353 0.0123886
R13335 gnd.n4384 gnd.n4357 0.0123886
R13336 gnd.n4381 gnd.n4380 0.0123886
R13337 gnd.n4377 gnd.n4363 0.0123886
R13338 gnd.n4376 gnd.n4368 0.0123886
R13339 gnd.n4573 gnd.n2121 0.0123886
R13340 gnd.n5704 gnd.n1395 0.0123886
R13341 gnd.n5701 gnd.n5700 0.0123886
R13342 gnd.n5697 gnd.n1399 0.0123886
R13343 gnd.n5696 gnd.n1404 0.0123886
R13344 gnd.n5693 gnd.n5692 0.0123886
R13345 gnd.n5689 gnd.n1408 0.0123886
R13346 gnd.n5688 gnd.n1412 0.0123886
R13347 gnd.n5685 gnd.n5684 0.0123886
R13348 gnd.n5681 gnd.n1416 0.0123886
R13349 gnd.n5680 gnd.n1420 0.0123886
R13350 gnd.n5677 gnd.n5676 0.0123886
R13351 gnd.n5673 gnd.n1424 0.0123886
R13352 gnd.n5672 gnd.n1428 0.0123886
R13353 gnd.n5669 gnd.n5668 0.0123886
R13354 gnd.n5665 gnd.n1432 0.0123886
R13355 gnd.n5664 gnd.n1436 0.0123886
R13356 gnd.n5661 gnd.n5660 0.0123886
R13357 gnd.n1445 gnd.n1442 0.0123886
R13358 gnd.n1637 gnd.n1636 0.0123886
R13359 gnd.n2979 gnd.n2693 0.00797283
R13360 gnd.n2981 gnd.n2980 0.00797283
R13361 gnd.n2982 gnd.n2688 0.00797283
R13362 gnd.n2990 gnd.n2686 0.00797283
R13363 gnd.n2992 gnd.n2991 0.00797283
R13364 gnd.n3010 gnd.n2667 0.00797283
R13365 gnd.n3012 gnd.n3011 0.00797283
R13366 gnd.n3013 gnd.n2662 0.00797283
R13367 gnd.n2661 gnd.n2657 0.00797283
R13368 gnd.n3023 gnd.n3022 0.00797283
R13369 gnd.n2659 gnd.n2658 0.00797283
R13370 gnd.n2641 gnd.n2640 0.00797283
R13371 gnd.n3043 gnd.n3042 0.00797283
R13372 gnd.n2642 gnd.n2617 0.00797283
R13373 gnd.n3077 gnd.n3076 0.00797283
R13374 gnd.n3079 gnd.n3078 0.00797283
R13375 gnd.n2612 gnd.n2564 0.00797283
R13376 gnd.n2614 gnd.n2565 0.00797283
R13377 gnd.n3088 gnd.n2566 0.00797283
R13378 gnd.n3090 gnd.n3089 0.00797283
R13379 gnd.n3092 gnd.n3091 0.00797283
R13380 gnd.n3094 gnd.n2586 0.00797283
R13381 gnd.n3097 gnd.n2587 0.00797283
R13382 gnd.n3099 gnd.n2588 0.00797283
R13383 gnd.n3102 gnd.n3100 0.00797283
R13384 gnd.n3101 gnd.n2487 0.00797283
R13385 gnd.n3169 gnd.n3167 0.00797283
R13386 gnd.n3168 gnd.n2480 0.00797283
R13387 gnd.n3179 gnd.n3178 0.00797283
R13388 gnd.n3181 gnd.n3180 0.00797283
R13389 gnd.n3184 gnd.n2478 0.00797283
R13390 gnd.n3188 gnd.n3187 0.00797283
R13391 gnd.n3186 gnd.n3185 0.00797283
R13392 gnd.n2458 gnd.n2457 0.00797283
R13393 gnd.n3210 gnd.n3209 0.00797283
R13394 gnd.n2459 gnd.n2432 0.00797283
R13395 gnd.n3254 gnd.n3252 0.00797283
R13396 gnd.n3253 gnd.n2425 0.00797283
R13397 gnd.n3264 gnd.n3263 0.00797283
R13398 gnd.n3266 gnd.n3265 0.00797283
R13399 gnd.n3269 gnd.n2423 0.00797283
R13400 gnd.n3273 gnd.n3272 0.00797283
R13401 gnd.n3271 gnd.n3270 0.00797283
R13402 gnd.n2403 gnd.n2402 0.00797283
R13403 gnd.n3295 gnd.n3294 0.00797283
R13404 gnd.n2404 gnd.n2378 0.00797283
R13405 gnd.n3343 gnd.n3341 0.00797283
R13406 gnd.n3342 gnd.n2371 0.00797283
R13407 gnd.n3354 gnd.n3353 0.00797283
R13408 gnd.n3612 gnd.n3611 0.00797283
R13409 gnd.n3615 gnd.n2369 0.00797283
R13410 gnd.n3617 gnd.n3616 0.00797283
R13411 gnd.n3640 gnd.n2350 0.00797283
R13412 gnd.n3641 gnd.n2314 0.00797283
R13413 gnd.n4426 gnd.n4271 0.00593478
R13414 gnd.n5706 gnd.n5705 0.00593478
R13415 CSoutput.n19 CSoutput.t133 184.661
R13416 CSoutput.n78 CSoutput.n77 165.8
R13417 CSoutput.n76 CSoutput.n0 165.8
R13418 CSoutput.n75 CSoutput.n74 165.8
R13419 CSoutput.n73 CSoutput.n72 165.8
R13420 CSoutput.n71 CSoutput.n2 165.8
R13421 CSoutput.n69 CSoutput.n68 165.8
R13422 CSoutput.n67 CSoutput.n3 165.8
R13423 CSoutput.n66 CSoutput.n65 165.8
R13424 CSoutput.n63 CSoutput.n4 165.8
R13425 CSoutput.n61 CSoutput.n60 165.8
R13426 CSoutput.n59 CSoutput.n5 165.8
R13427 CSoutput.n58 CSoutput.n57 165.8
R13428 CSoutput.n55 CSoutput.n6 165.8
R13429 CSoutput.n54 CSoutput.n53 165.8
R13430 CSoutput.n52 CSoutput.n51 165.8
R13431 CSoutput.n50 CSoutput.n8 165.8
R13432 CSoutput.n48 CSoutput.n47 165.8
R13433 CSoutput.n46 CSoutput.n9 165.8
R13434 CSoutput.n45 CSoutput.n44 165.8
R13435 CSoutput.n42 CSoutput.n10 165.8
R13436 CSoutput.n41 CSoutput.n40 165.8
R13437 CSoutput.n39 CSoutput.n38 165.8
R13438 CSoutput.n37 CSoutput.n12 165.8
R13439 CSoutput.n35 CSoutput.n34 165.8
R13440 CSoutput.n33 CSoutput.n13 165.8
R13441 CSoutput.n32 CSoutput.n31 165.8
R13442 CSoutput.n29 CSoutput.n14 165.8
R13443 CSoutput.n28 CSoutput.n27 165.8
R13444 CSoutput.n26 CSoutput.n25 165.8
R13445 CSoutput.n24 CSoutput.n16 165.8
R13446 CSoutput.n22 CSoutput.n21 165.8
R13447 CSoutput.n20 CSoutput.n17 165.8
R13448 CSoutput.n77 CSoutput.t134 162.194
R13449 CSoutput.n18 CSoutput.t135 120.501
R13450 CSoutput.n23 CSoutput.t122 120.501
R13451 CSoutput.n15 CSoutput.t141 120.501
R13452 CSoutput.n30 CSoutput.t138 120.501
R13453 CSoutput.n36 CSoutput.t124 120.501
R13454 CSoutput.n11 CSoutput.t126 120.501
R13455 CSoutput.n43 CSoutput.t139 120.501
R13456 CSoutput.n49 CSoutput.t128 120.501
R13457 CSoutput.n7 CSoutput.t129 120.501
R13458 CSoutput.n56 CSoutput.t123 120.501
R13459 CSoutput.n62 CSoutput.t137 120.501
R13460 CSoutput.n64 CSoutput.t132 120.501
R13461 CSoutput.n70 CSoutput.t125 120.501
R13462 CSoutput.n1 CSoutput.t121 120.501
R13463 CSoutput.n270 CSoutput.n268 103.469
R13464 CSoutput.n262 CSoutput.n260 103.469
R13465 CSoutput.n255 CSoutput.n253 103.469
R13466 CSoutput.n96 CSoutput.n94 103.469
R13467 CSoutput.n88 CSoutput.n86 103.469
R13468 CSoutput.n81 CSoutput.n79 103.469
R13469 CSoutput.n272 CSoutput.n271 103.111
R13470 CSoutput.n270 CSoutput.n269 103.111
R13471 CSoutput.n266 CSoutput.n265 103.111
R13472 CSoutput.n264 CSoutput.n263 103.111
R13473 CSoutput.n262 CSoutput.n261 103.111
R13474 CSoutput.n259 CSoutput.n258 103.111
R13475 CSoutput.n257 CSoutput.n256 103.111
R13476 CSoutput.n255 CSoutput.n254 103.111
R13477 CSoutput.n96 CSoutput.n95 103.111
R13478 CSoutput.n98 CSoutput.n97 103.111
R13479 CSoutput.n100 CSoutput.n99 103.111
R13480 CSoutput.n88 CSoutput.n87 103.111
R13481 CSoutput.n90 CSoutput.n89 103.111
R13482 CSoutput.n92 CSoutput.n91 103.111
R13483 CSoutput.n81 CSoutput.n80 103.111
R13484 CSoutput.n83 CSoutput.n82 103.111
R13485 CSoutput.n85 CSoutput.n84 103.111
R13486 CSoutput.n274 CSoutput.n273 103.111
R13487 CSoutput.n302 CSoutput.n300 81.5057
R13488 CSoutput.n290 CSoutput.n288 81.5057
R13489 CSoutput.n279 CSoutput.n277 81.5057
R13490 CSoutput.n338 CSoutput.n336 81.5057
R13491 CSoutput.n326 CSoutput.n324 81.5057
R13492 CSoutput.n315 CSoutput.n313 81.5057
R13493 CSoutput.n310 CSoutput.n309 80.9324
R13494 CSoutput.n308 CSoutput.n307 80.9324
R13495 CSoutput.n306 CSoutput.n305 80.9324
R13496 CSoutput.n304 CSoutput.n303 80.9324
R13497 CSoutput.n302 CSoutput.n301 80.9324
R13498 CSoutput.n298 CSoutput.n297 80.9324
R13499 CSoutput.n296 CSoutput.n295 80.9324
R13500 CSoutput.n294 CSoutput.n293 80.9324
R13501 CSoutput.n292 CSoutput.n291 80.9324
R13502 CSoutput.n290 CSoutput.n289 80.9324
R13503 CSoutput.n287 CSoutput.n286 80.9324
R13504 CSoutput.n285 CSoutput.n284 80.9324
R13505 CSoutput.n283 CSoutput.n282 80.9324
R13506 CSoutput.n281 CSoutput.n280 80.9324
R13507 CSoutput.n279 CSoutput.n278 80.9324
R13508 CSoutput.n338 CSoutput.n337 80.9324
R13509 CSoutput.n340 CSoutput.n339 80.9324
R13510 CSoutput.n342 CSoutput.n341 80.9324
R13511 CSoutput.n344 CSoutput.n343 80.9324
R13512 CSoutput.n346 CSoutput.n345 80.9324
R13513 CSoutput.n326 CSoutput.n325 80.9324
R13514 CSoutput.n328 CSoutput.n327 80.9324
R13515 CSoutput.n330 CSoutput.n329 80.9324
R13516 CSoutput.n332 CSoutput.n331 80.9324
R13517 CSoutput.n334 CSoutput.n333 80.9324
R13518 CSoutput.n315 CSoutput.n314 80.9324
R13519 CSoutput.n317 CSoutput.n316 80.9324
R13520 CSoutput.n319 CSoutput.n318 80.9324
R13521 CSoutput.n321 CSoutput.n320 80.9324
R13522 CSoutput.n323 CSoutput.n322 80.9324
R13523 CSoutput.n25 CSoutput.n24 48.1486
R13524 CSoutput.n69 CSoutput.n3 48.1486
R13525 CSoutput.n38 CSoutput.n37 48.1486
R13526 CSoutput.n42 CSoutput.n41 48.1486
R13527 CSoutput.n51 CSoutput.n50 48.1486
R13528 CSoutput.n55 CSoutput.n54 48.1486
R13529 CSoutput.n22 CSoutput.n17 46.462
R13530 CSoutput.n72 CSoutput.n71 46.462
R13531 CSoutput.n20 CSoutput.n19 44.9055
R13532 CSoutput.n29 CSoutput.n28 43.7635
R13533 CSoutput.n65 CSoutput.n63 43.7635
R13534 CSoutput.n35 CSoutput.n13 41.7396
R13535 CSoutput.n57 CSoutput.n5 41.7396
R13536 CSoutput.n44 CSoutput.n9 37.0171
R13537 CSoutput.n48 CSoutput.n9 37.0171
R13538 CSoutput.n76 CSoutput.n75 34.9932
R13539 CSoutput.n31 CSoutput.n13 32.2947
R13540 CSoutput.n61 CSoutput.n5 32.2947
R13541 CSoutput.n30 CSoutput.n29 29.6014
R13542 CSoutput.n63 CSoutput.n62 29.6014
R13543 CSoutput.n19 CSoutput.n18 28.4085
R13544 CSoutput.n18 CSoutput.n17 25.1176
R13545 CSoutput.n72 CSoutput.n1 25.1176
R13546 CSoutput.n43 CSoutput.n42 22.0922
R13547 CSoutput.n50 CSoutput.n49 22.0922
R13548 CSoutput.n77 CSoutput.n76 21.8586
R13549 CSoutput.n37 CSoutput.n36 18.9681
R13550 CSoutput.n56 CSoutput.n55 18.9681
R13551 CSoutput.n25 CSoutput.n15 17.6292
R13552 CSoutput.n64 CSoutput.n3 17.6292
R13553 CSoutput.n24 CSoutput.n23 15.844
R13554 CSoutput.n70 CSoutput.n69 15.844
R13555 CSoutput.n38 CSoutput.n11 14.5051
R13556 CSoutput.n54 CSoutput.n7 14.5051
R13557 CSoutput.n349 CSoutput.n78 11.4982
R13558 CSoutput.n41 CSoutput.n11 11.3811
R13559 CSoutput.n51 CSoutput.n7 11.3811
R13560 CSoutput.n23 CSoutput.n22 10.0422
R13561 CSoutput.n71 CSoutput.n70 10.0422
R13562 CSoutput.n267 CSoutput.n259 9.25285
R13563 CSoutput.n93 CSoutput.n85 9.25285
R13564 CSoutput.n299 CSoutput.n287 8.98182
R13565 CSoutput.n335 CSoutput.n323 8.98182
R13566 CSoutput.n312 CSoutput.n276 8.92829
R13567 CSoutput.n28 CSoutput.n15 8.25698
R13568 CSoutput.n65 CSoutput.n64 8.25698
R13569 CSoutput.n276 CSoutput.n275 7.12641
R13570 CSoutput.n102 CSoutput.n101 7.12641
R13571 CSoutput.n36 CSoutput.n35 6.91809
R13572 CSoutput.n57 CSoutput.n56 6.91809
R13573 CSoutput.n312 CSoutput.n311 6.02792
R13574 CSoutput.n348 CSoutput.n347 6.02792
R13575 CSoutput.n349 CSoutput.n102 5.33585
R13576 CSoutput.n311 CSoutput.n310 5.25266
R13577 CSoutput.n299 CSoutput.n298 5.25266
R13578 CSoutput.n347 CSoutput.n346 5.25266
R13579 CSoutput.n335 CSoutput.n334 5.25266
R13580 CSoutput.n275 CSoutput.n274 5.1449
R13581 CSoutput.n267 CSoutput.n266 5.1449
R13582 CSoutput.n101 CSoutput.n100 5.1449
R13583 CSoutput.n93 CSoutput.n92 5.1449
R13584 CSoutput.n193 CSoutput.n146 4.5005
R13585 CSoutput.n162 CSoutput.n146 4.5005
R13586 CSoutput.n157 CSoutput.n141 4.5005
R13587 CSoutput.n157 CSoutput.n143 4.5005
R13588 CSoutput.n157 CSoutput.n140 4.5005
R13589 CSoutput.n157 CSoutput.n144 4.5005
R13590 CSoutput.n157 CSoutput.n139 4.5005
R13591 CSoutput.n157 CSoutput.t127 4.5005
R13592 CSoutput.n157 CSoutput.n138 4.5005
R13593 CSoutput.n157 CSoutput.n145 4.5005
R13594 CSoutput.n157 CSoutput.n146 4.5005
R13595 CSoutput.n155 CSoutput.n141 4.5005
R13596 CSoutput.n155 CSoutput.n143 4.5005
R13597 CSoutput.n155 CSoutput.n140 4.5005
R13598 CSoutput.n155 CSoutput.n144 4.5005
R13599 CSoutput.n155 CSoutput.n139 4.5005
R13600 CSoutput.n155 CSoutput.t127 4.5005
R13601 CSoutput.n155 CSoutput.n138 4.5005
R13602 CSoutput.n155 CSoutput.n145 4.5005
R13603 CSoutput.n155 CSoutput.n146 4.5005
R13604 CSoutput.n154 CSoutput.n141 4.5005
R13605 CSoutput.n154 CSoutput.n143 4.5005
R13606 CSoutput.n154 CSoutput.n140 4.5005
R13607 CSoutput.n154 CSoutput.n144 4.5005
R13608 CSoutput.n154 CSoutput.n139 4.5005
R13609 CSoutput.n154 CSoutput.t127 4.5005
R13610 CSoutput.n154 CSoutput.n138 4.5005
R13611 CSoutput.n154 CSoutput.n145 4.5005
R13612 CSoutput.n154 CSoutput.n146 4.5005
R13613 CSoutput.n239 CSoutput.n141 4.5005
R13614 CSoutput.n239 CSoutput.n143 4.5005
R13615 CSoutput.n239 CSoutput.n140 4.5005
R13616 CSoutput.n239 CSoutput.n144 4.5005
R13617 CSoutput.n239 CSoutput.n139 4.5005
R13618 CSoutput.n239 CSoutput.t127 4.5005
R13619 CSoutput.n239 CSoutput.n138 4.5005
R13620 CSoutput.n239 CSoutput.n145 4.5005
R13621 CSoutput.n239 CSoutput.n146 4.5005
R13622 CSoutput.n237 CSoutput.n141 4.5005
R13623 CSoutput.n237 CSoutput.n143 4.5005
R13624 CSoutput.n237 CSoutput.n140 4.5005
R13625 CSoutput.n237 CSoutput.n144 4.5005
R13626 CSoutput.n237 CSoutput.n139 4.5005
R13627 CSoutput.n237 CSoutput.t127 4.5005
R13628 CSoutput.n237 CSoutput.n138 4.5005
R13629 CSoutput.n237 CSoutput.n145 4.5005
R13630 CSoutput.n235 CSoutput.n141 4.5005
R13631 CSoutput.n235 CSoutput.n143 4.5005
R13632 CSoutput.n235 CSoutput.n140 4.5005
R13633 CSoutput.n235 CSoutput.n144 4.5005
R13634 CSoutput.n235 CSoutput.n139 4.5005
R13635 CSoutput.n235 CSoutput.t127 4.5005
R13636 CSoutput.n235 CSoutput.n138 4.5005
R13637 CSoutput.n235 CSoutput.n145 4.5005
R13638 CSoutput.n165 CSoutput.n141 4.5005
R13639 CSoutput.n165 CSoutput.n143 4.5005
R13640 CSoutput.n165 CSoutput.n140 4.5005
R13641 CSoutput.n165 CSoutput.n144 4.5005
R13642 CSoutput.n165 CSoutput.n139 4.5005
R13643 CSoutput.n165 CSoutput.t127 4.5005
R13644 CSoutput.n165 CSoutput.n138 4.5005
R13645 CSoutput.n165 CSoutput.n145 4.5005
R13646 CSoutput.n165 CSoutput.n146 4.5005
R13647 CSoutput.n164 CSoutput.n141 4.5005
R13648 CSoutput.n164 CSoutput.n143 4.5005
R13649 CSoutput.n164 CSoutput.n140 4.5005
R13650 CSoutput.n164 CSoutput.n144 4.5005
R13651 CSoutput.n164 CSoutput.n139 4.5005
R13652 CSoutput.n164 CSoutput.t127 4.5005
R13653 CSoutput.n164 CSoutput.n138 4.5005
R13654 CSoutput.n164 CSoutput.n145 4.5005
R13655 CSoutput.n164 CSoutput.n146 4.5005
R13656 CSoutput.n168 CSoutput.n141 4.5005
R13657 CSoutput.n168 CSoutput.n143 4.5005
R13658 CSoutput.n168 CSoutput.n140 4.5005
R13659 CSoutput.n168 CSoutput.n144 4.5005
R13660 CSoutput.n168 CSoutput.n139 4.5005
R13661 CSoutput.n168 CSoutput.t127 4.5005
R13662 CSoutput.n168 CSoutput.n138 4.5005
R13663 CSoutput.n168 CSoutput.n145 4.5005
R13664 CSoutput.n168 CSoutput.n146 4.5005
R13665 CSoutput.n167 CSoutput.n141 4.5005
R13666 CSoutput.n167 CSoutput.n143 4.5005
R13667 CSoutput.n167 CSoutput.n140 4.5005
R13668 CSoutput.n167 CSoutput.n144 4.5005
R13669 CSoutput.n167 CSoutput.n139 4.5005
R13670 CSoutput.n167 CSoutput.t127 4.5005
R13671 CSoutput.n167 CSoutput.n138 4.5005
R13672 CSoutput.n167 CSoutput.n145 4.5005
R13673 CSoutput.n167 CSoutput.n146 4.5005
R13674 CSoutput.n150 CSoutput.n141 4.5005
R13675 CSoutput.n150 CSoutput.n143 4.5005
R13676 CSoutput.n150 CSoutput.n140 4.5005
R13677 CSoutput.n150 CSoutput.n144 4.5005
R13678 CSoutput.n150 CSoutput.n139 4.5005
R13679 CSoutput.n150 CSoutput.t127 4.5005
R13680 CSoutput.n150 CSoutput.n138 4.5005
R13681 CSoutput.n150 CSoutput.n145 4.5005
R13682 CSoutput.n150 CSoutput.n146 4.5005
R13683 CSoutput.n242 CSoutput.n141 4.5005
R13684 CSoutput.n242 CSoutput.n143 4.5005
R13685 CSoutput.n242 CSoutput.n140 4.5005
R13686 CSoutput.n242 CSoutput.n144 4.5005
R13687 CSoutput.n242 CSoutput.n139 4.5005
R13688 CSoutput.n242 CSoutput.t127 4.5005
R13689 CSoutput.n242 CSoutput.n138 4.5005
R13690 CSoutput.n242 CSoutput.n145 4.5005
R13691 CSoutput.n242 CSoutput.n146 4.5005
R13692 CSoutput.n229 CSoutput.n200 4.5005
R13693 CSoutput.n229 CSoutput.n206 4.5005
R13694 CSoutput.n187 CSoutput.n176 4.5005
R13695 CSoutput.n187 CSoutput.n178 4.5005
R13696 CSoutput.n187 CSoutput.n175 4.5005
R13697 CSoutput.n187 CSoutput.n179 4.5005
R13698 CSoutput.n187 CSoutput.n174 4.5005
R13699 CSoutput.n187 CSoutput.t120 4.5005
R13700 CSoutput.n187 CSoutput.n173 4.5005
R13701 CSoutput.n187 CSoutput.n180 4.5005
R13702 CSoutput.n229 CSoutput.n187 4.5005
R13703 CSoutput.n208 CSoutput.n176 4.5005
R13704 CSoutput.n208 CSoutput.n178 4.5005
R13705 CSoutput.n208 CSoutput.n175 4.5005
R13706 CSoutput.n208 CSoutput.n179 4.5005
R13707 CSoutput.n208 CSoutput.n174 4.5005
R13708 CSoutput.n208 CSoutput.t120 4.5005
R13709 CSoutput.n208 CSoutput.n173 4.5005
R13710 CSoutput.n208 CSoutput.n180 4.5005
R13711 CSoutput.n229 CSoutput.n208 4.5005
R13712 CSoutput.n186 CSoutput.n176 4.5005
R13713 CSoutput.n186 CSoutput.n178 4.5005
R13714 CSoutput.n186 CSoutput.n175 4.5005
R13715 CSoutput.n186 CSoutput.n179 4.5005
R13716 CSoutput.n186 CSoutput.n174 4.5005
R13717 CSoutput.n186 CSoutput.t120 4.5005
R13718 CSoutput.n186 CSoutput.n173 4.5005
R13719 CSoutput.n186 CSoutput.n180 4.5005
R13720 CSoutput.n229 CSoutput.n186 4.5005
R13721 CSoutput.n210 CSoutput.n176 4.5005
R13722 CSoutput.n210 CSoutput.n178 4.5005
R13723 CSoutput.n210 CSoutput.n175 4.5005
R13724 CSoutput.n210 CSoutput.n179 4.5005
R13725 CSoutput.n210 CSoutput.n174 4.5005
R13726 CSoutput.n210 CSoutput.t120 4.5005
R13727 CSoutput.n210 CSoutput.n173 4.5005
R13728 CSoutput.n210 CSoutput.n180 4.5005
R13729 CSoutput.n229 CSoutput.n210 4.5005
R13730 CSoutput.n176 CSoutput.n171 4.5005
R13731 CSoutput.n178 CSoutput.n171 4.5005
R13732 CSoutput.n175 CSoutput.n171 4.5005
R13733 CSoutput.n179 CSoutput.n171 4.5005
R13734 CSoutput.n174 CSoutput.n171 4.5005
R13735 CSoutput.t120 CSoutput.n171 4.5005
R13736 CSoutput.n173 CSoutput.n171 4.5005
R13737 CSoutput.n180 CSoutput.n171 4.5005
R13738 CSoutput.n232 CSoutput.n176 4.5005
R13739 CSoutput.n232 CSoutput.n178 4.5005
R13740 CSoutput.n232 CSoutput.n175 4.5005
R13741 CSoutput.n232 CSoutput.n179 4.5005
R13742 CSoutput.n232 CSoutput.n174 4.5005
R13743 CSoutput.n232 CSoutput.t120 4.5005
R13744 CSoutput.n232 CSoutput.n173 4.5005
R13745 CSoutput.n232 CSoutput.n180 4.5005
R13746 CSoutput.n230 CSoutput.n176 4.5005
R13747 CSoutput.n230 CSoutput.n178 4.5005
R13748 CSoutput.n230 CSoutput.n175 4.5005
R13749 CSoutput.n230 CSoutput.n179 4.5005
R13750 CSoutput.n230 CSoutput.n174 4.5005
R13751 CSoutput.n230 CSoutput.t120 4.5005
R13752 CSoutput.n230 CSoutput.n173 4.5005
R13753 CSoutput.n230 CSoutput.n180 4.5005
R13754 CSoutput.n230 CSoutput.n229 4.5005
R13755 CSoutput.n212 CSoutput.n176 4.5005
R13756 CSoutput.n212 CSoutput.n178 4.5005
R13757 CSoutput.n212 CSoutput.n175 4.5005
R13758 CSoutput.n212 CSoutput.n179 4.5005
R13759 CSoutput.n212 CSoutput.n174 4.5005
R13760 CSoutput.n212 CSoutput.t120 4.5005
R13761 CSoutput.n212 CSoutput.n173 4.5005
R13762 CSoutput.n212 CSoutput.n180 4.5005
R13763 CSoutput.n229 CSoutput.n212 4.5005
R13764 CSoutput.n184 CSoutput.n176 4.5005
R13765 CSoutput.n184 CSoutput.n178 4.5005
R13766 CSoutput.n184 CSoutput.n175 4.5005
R13767 CSoutput.n184 CSoutput.n179 4.5005
R13768 CSoutput.n184 CSoutput.n174 4.5005
R13769 CSoutput.n184 CSoutput.t120 4.5005
R13770 CSoutput.n184 CSoutput.n173 4.5005
R13771 CSoutput.n184 CSoutput.n180 4.5005
R13772 CSoutput.n229 CSoutput.n184 4.5005
R13773 CSoutput.n214 CSoutput.n176 4.5005
R13774 CSoutput.n214 CSoutput.n178 4.5005
R13775 CSoutput.n214 CSoutput.n175 4.5005
R13776 CSoutput.n214 CSoutput.n179 4.5005
R13777 CSoutput.n214 CSoutput.n174 4.5005
R13778 CSoutput.n214 CSoutput.t120 4.5005
R13779 CSoutput.n214 CSoutput.n173 4.5005
R13780 CSoutput.n214 CSoutput.n180 4.5005
R13781 CSoutput.n229 CSoutput.n214 4.5005
R13782 CSoutput.n183 CSoutput.n176 4.5005
R13783 CSoutput.n183 CSoutput.n178 4.5005
R13784 CSoutput.n183 CSoutput.n175 4.5005
R13785 CSoutput.n183 CSoutput.n179 4.5005
R13786 CSoutput.n183 CSoutput.n174 4.5005
R13787 CSoutput.n183 CSoutput.t120 4.5005
R13788 CSoutput.n183 CSoutput.n173 4.5005
R13789 CSoutput.n183 CSoutput.n180 4.5005
R13790 CSoutput.n229 CSoutput.n183 4.5005
R13791 CSoutput.n228 CSoutput.n176 4.5005
R13792 CSoutput.n228 CSoutput.n178 4.5005
R13793 CSoutput.n228 CSoutput.n175 4.5005
R13794 CSoutput.n228 CSoutput.n179 4.5005
R13795 CSoutput.n228 CSoutput.n174 4.5005
R13796 CSoutput.n228 CSoutput.t120 4.5005
R13797 CSoutput.n228 CSoutput.n173 4.5005
R13798 CSoutput.n228 CSoutput.n180 4.5005
R13799 CSoutput.n229 CSoutput.n228 4.5005
R13800 CSoutput.n227 CSoutput.n112 4.5005
R13801 CSoutput.n128 CSoutput.n112 4.5005
R13802 CSoutput.n123 CSoutput.n107 4.5005
R13803 CSoutput.n123 CSoutput.n109 4.5005
R13804 CSoutput.n123 CSoutput.n106 4.5005
R13805 CSoutput.n123 CSoutput.n110 4.5005
R13806 CSoutput.n123 CSoutput.n105 4.5005
R13807 CSoutput.n123 CSoutput.t140 4.5005
R13808 CSoutput.n123 CSoutput.n104 4.5005
R13809 CSoutput.n123 CSoutput.n111 4.5005
R13810 CSoutput.n123 CSoutput.n112 4.5005
R13811 CSoutput.n121 CSoutput.n107 4.5005
R13812 CSoutput.n121 CSoutput.n109 4.5005
R13813 CSoutput.n121 CSoutput.n106 4.5005
R13814 CSoutput.n121 CSoutput.n110 4.5005
R13815 CSoutput.n121 CSoutput.n105 4.5005
R13816 CSoutput.n121 CSoutput.t140 4.5005
R13817 CSoutput.n121 CSoutput.n104 4.5005
R13818 CSoutput.n121 CSoutput.n111 4.5005
R13819 CSoutput.n121 CSoutput.n112 4.5005
R13820 CSoutput.n120 CSoutput.n107 4.5005
R13821 CSoutput.n120 CSoutput.n109 4.5005
R13822 CSoutput.n120 CSoutput.n106 4.5005
R13823 CSoutput.n120 CSoutput.n110 4.5005
R13824 CSoutput.n120 CSoutput.n105 4.5005
R13825 CSoutput.n120 CSoutput.t140 4.5005
R13826 CSoutput.n120 CSoutput.n104 4.5005
R13827 CSoutput.n120 CSoutput.n111 4.5005
R13828 CSoutput.n120 CSoutput.n112 4.5005
R13829 CSoutput.n249 CSoutput.n107 4.5005
R13830 CSoutput.n249 CSoutput.n109 4.5005
R13831 CSoutput.n249 CSoutput.n106 4.5005
R13832 CSoutput.n249 CSoutput.n110 4.5005
R13833 CSoutput.n249 CSoutput.n105 4.5005
R13834 CSoutput.n249 CSoutput.t140 4.5005
R13835 CSoutput.n249 CSoutput.n104 4.5005
R13836 CSoutput.n249 CSoutput.n111 4.5005
R13837 CSoutput.n249 CSoutput.n112 4.5005
R13838 CSoutput.n247 CSoutput.n107 4.5005
R13839 CSoutput.n247 CSoutput.n109 4.5005
R13840 CSoutput.n247 CSoutput.n106 4.5005
R13841 CSoutput.n247 CSoutput.n110 4.5005
R13842 CSoutput.n247 CSoutput.n105 4.5005
R13843 CSoutput.n247 CSoutput.t140 4.5005
R13844 CSoutput.n247 CSoutput.n104 4.5005
R13845 CSoutput.n247 CSoutput.n111 4.5005
R13846 CSoutput.n245 CSoutput.n107 4.5005
R13847 CSoutput.n245 CSoutput.n109 4.5005
R13848 CSoutput.n245 CSoutput.n106 4.5005
R13849 CSoutput.n245 CSoutput.n110 4.5005
R13850 CSoutput.n245 CSoutput.n105 4.5005
R13851 CSoutput.n245 CSoutput.t140 4.5005
R13852 CSoutput.n245 CSoutput.n104 4.5005
R13853 CSoutput.n245 CSoutput.n111 4.5005
R13854 CSoutput.n131 CSoutput.n107 4.5005
R13855 CSoutput.n131 CSoutput.n109 4.5005
R13856 CSoutput.n131 CSoutput.n106 4.5005
R13857 CSoutput.n131 CSoutput.n110 4.5005
R13858 CSoutput.n131 CSoutput.n105 4.5005
R13859 CSoutput.n131 CSoutput.t140 4.5005
R13860 CSoutput.n131 CSoutput.n104 4.5005
R13861 CSoutput.n131 CSoutput.n111 4.5005
R13862 CSoutput.n131 CSoutput.n112 4.5005
R13863 CSoutput.n130 CSoutput.n107 4.5005
R13864 CSoutput.n130 CSoutput.n109 4.5005
R13865 CSoutput.n130 CSoutput.n106 4.5005
R13866 CSoutput.n130 CSoutput.n110 4.5005
R13867 CSoutput.n130 CSoutput.n105 4.5005
R13868 CSoutput.n130 CSoutput.t140 4.5005
R13869 CSoutput.n130 CSoutput.n104 4.5005
R13870 CSoutput.n130 CSoutput.n111 4.5005
R13871 CSoutput.n130 CSoutput.n112 4.5005
R13872 CSoutput.n134 CSoutput.n107 4.5005
R13873 CSoutput.n134 CSoutput.n109 4.5005
R13874 CSoutput.n134 CSoutput.n106 4.5005
R13875 CSoutput.n134 CSoutput.n110 4.5005
R13876 CSoutput.n134 CSoutput.n105 4.5005
R13877 CSoutput.n134 CSoutput.t140 4.5005
R13878 CSoutput.n134 CSoutput.n104 4.5005
R13879 CSoutput.n134 CSoutput.n111 4.5005
R13880 CSoutput.n134 CSoutput.n112 4.5005
R13881 CSoutput.n133 CSoutput.n107 4.5005
R13882 CSoutput.n133 CSoutput.n109 4.5005
R13883 CSoutput.n133 CSoutput.n106 4.5005
R13884 CSoutput.n133 CSoutput.n110 4.5005
R13885 CSoutput.n133 CSoutput.n105 4.5005
R13886 CSoutput.n133 CSoutput.t140 4.5005
R13887 CSoutput.n133 CSoutput.n104 4.5005
R13888 CSoutput.n133 CSoutput.n111 4.5005
R13889 CSoutput.n133 CSoutput.n112 4.5005
R13890 CSoutput.n116 CSoutput.n107 4.5005
R13891 CSoutput.n116 CSoutput.n109 4.5005
R13892 CSoutput.n116 CSoutput.n106 4.5005
R13893 CSoutput.n116 CSoutput.n110 4.5005
R13894 CSoutput.n116 CSoutput.n105 4.5005
R13895 CSoutput.n116 CSoutput.t140 4.5005
R13896 CSoutput.n116 CSoutput.n104 4.5005
R13897 CSoutput.n116 CSoutput.n111 4.5005
R13898 CSoutput.n116 CSoutput.n112 4.5005
R13899 CSoutput.n252 CSoutput.n107 4.5005
R13900 CSoutput.n252 CSoutput.n109 4.5005
R13901 CSoutput.n252 CSoutput.n106 4.5005
R13902 CSoutput.n252 CSoutput.n110 4.5005
R13903 CSoutput.n252 CSoutput.n105 4.5005
R13904 CSoutput.n252 CSoutput.t140 4.5005
R13905 CSoutput.n252 CSoutput.n104 4.5005
R13906 CSoutput.n252 CSoutput.n111 4.5005
R13907 CSoutput.n252 CSoutput.n112 4.5005
R13908 CSoutput.n275 CSoutput.n267 4.10845
R13909 CSoutput.n101 CSoutput.n93 4.10845
R13910 CSoutput.n273 CSoutput.t29 4.06363
R13911 CSoutput.n273 CSoutput.t114 4.06363
R13912 CSoutput.n271 CSoutput.t17 4.06363
R13913 CSoutput.n271 CSoutput.t33 4.06363
R13914 CSoutput.n269 CSoutput.t110 4.06363
R13915 CSoutput.n269 CSoutput.t6 4.06363
R13916 CSoutput.n268 CSoutput.t8 4.06363
R13917 CSoutput.n268 CSoutput.t25 4.06363
R13918 CSoutput.n265 CSoutput.t115 4.06363
R13919 CSoutput.n265 CSoutput.t31 4.06363
R13920 CSoutput.n263 CSoutput.t30 4.06363
R13921 CSoutput.n263 CSoutput.t11 4.06363
R13922 CSoutput.n261 CSoutput.t4 4.06363
R13923 CSoutput.n261 CSoutput.t5 4.06363
R13924 CSoutput.n260 CSoutput.t35 4.06363
R13925 CSoutput.n260 CSoutput.t109 4.06363
R13926 CSoutput.n258 CSoutput.t14 4.06363
R13927 CSoutput.n258 CSoutput.t2 4.06363
R13928 CSoutput.n256 CSoutput.t18 4.06363
R13929 CSoutput.n256 CSoutput.t28 4.06363
R13930 CSoutput.n254 CSoutput.t23 4.06363
R13931 CSoutput.n254 CSoutput.t24 4.06363
R13932 CSoutput.n253 CSoutput.t26 4.06363
R13933 CSoutput.n253 CSoutput.t1 4.06363
R13934 CSoutput.n94 CSoutput.t10 4.06363
R13935 CSoutput.n94 CSoutput.t13 4.06363
R13936 CSoutput.n95 CSoutput.t15 4.06363
R13937 CSoutput.n95 CSoutput.t112 4.06363
R13938 CSoutput.n97 CSoutput.t34 4.06363
R13939 CSoutput.n97 CSoutput.t119 4.06363
R13940 CSoutput.n99 CSoutput.t19 4.06363
R13941 CSoutput.n99 CSoutput.t20 4.06363
R13942 CSoutput.n86 CSoutput.t12 4.06363
R13943 CSoutput.n86 CSoutput.t27 4.06363
R13944 CSoutput.n87 CSoutput.t16 4.06363
R13945 CSoutput.n87 CSoutput.t118 4.06363
R13946 CSoutput.n89 CSoutput.t113 4.06363
R13947 CSoutput.n89 CSoutput.t22 4.06363
R13948 CSoutput.n91 CSoutput.t0 4.06363
R13949 CSoutput.n91 CSoutput.t116 4.06363
R13950 CSoutput.n79 CSoutput.t111 4.06363
R13951 CSoutput.n79 CSoutput.t9 4.06363
R13952 CSoutput.n80 CSoutput.t36 4.06363
R13953 CSoutput.n80 CSoutput.t32 4.06363
R13954 CSoutput.n82 CSoutput.t3 4.06363
R13955 CSoutput.n82 CSoutput.t117 4.06363
R13956 CSoutput.n84 CSoutput.t21 4.06363
R13957 CSoutput.n84 CSoutput.t7 4.06363
R13958 CSoutput.n44 CSoutput.n43 3.79402
R13959 CSoutput.n49 CSoutput.n48 3.79402
R13960 CSoutput.n311 CSoutput.n299 3.72967
R13961 CSoutput.n347 CSoutput.n335 3.72967
R13962 CSoutput.n349 CSoutput.n348 3.57343
R13963 CSoutput.n309 CSoutput.t54 2.82907
R13964 CSoutput.n309 CSoutput.t58 2.82907
R13965 CSoutput.n307 CSoutput.t53 2.82907
R13966 CSoutput.n307 CSoutput.t108 2.82907
R13967 CSoutput.n305 CSoutput.t69 2.82907
R13968 CSoutput.n305 CSoutput.t48 2.82907
R13969 CSoutput.n303 CSoutput.t41 2.82907
R13970 CSoutput.n303 CSoutput.t89 2.82907
R13971 CSoutput.n301 CSoutput.t60 2.82907
R13972 CSoutput.n301 CSoutput.t63 2.82907
R13973 CSoutput.n300 CSoutput.t47 2.82907
R13974 CSoutput.n300 CSoutput.t99 2.82907
R13975 CSoutput.n297 CSoutput.t40 2.82907
R13976 CSoutput.n297 CSoutput.t87 2.82907
R13977 CSoutput.n295 CSoutput.t85 2.82907
R13978 CSoutput.n295 CSoutput.t73 2.82907
R13979 CSoutput.n293 CSoutput.t98 2.82907
R13980 CSoutput.n293 CSoutput.t39 2.82907
R13981 CSoutput.n291 CSoutput.t38 2.82907
R13982 CSoutput.n291 CSoutput.t91 2.82907
R13983 CSoutput.n289 CSoutput.t46 2.82907
R13984 CSoutput.n289 CSoutput.t97 2.82907
R13985 CSoutput.n288 CSoutput.t104 2.82907
R13986 CSoutput.n288 CSoutput.t37 2.82907
R13987 CSoutput.n286 CSoutput.t76 2.82907
R13988 CSoutput.n286 CSoutput.t83 2.82907
R13989 CSoutput.n284 CSoutput.t68 2.82907
R13990 CSoutput.n284 CSoutput.t96 2.82907
R13991 CSoutput.n282 CSoutput.t79 2.82907
R13992 CSoutput.n282 CSoutput.t62 2.82907
R13993 CSoutput.n280 CSoutput.t56 2.82907
R13994 CSoutput.n280 CSoutput.t70 2.82907
R13995 CSoutput.n278 CSoutput.t61 2.82907
R13996 CSoutput.n278 CSoutput.t66 2.82907
R13997 CSoutput.n277 CSoutput.t67 2.82907
R13998 CSoutput.n277 CSoutput.t107 2.82907
R13999 CSoutput.n336 CSoutput.t75 2.82907
R14000 CSoutput.n336 CSoutput.t93 2.82907
R14001 CSoutput.n337 CSoutput.t55 2.82907
R14002 CSoutput.n337 CSoutput.t65 2.82907
R14003 CSoutput.n339 CSoutput.t71 2.82907
R14004 CSoutput.n339 CSoutput.t82 2.82907
R14005 CSoutput.n341 CSoutput.t94 2.82907
R14006 CSoutput.n341 CSoutput.t74 2.82907
R14007 CSoutput.n343 CSoutput.t78 2.82907
R14008 CSoutput.n343 CSoutput.t103 2.82907
R14009 CSoutput.n345 CSoutput.t43 2.82907
R14010 CSoutput.n345 CSoutput.t59 2.82907
R14011 CSoutput.n324 CSoutput.t49 2.82907
R14012 CSoutput.n324 CSoutput.t44 2.82907
R14013 CSoutput.n325 CSoutput.t42 2.82907
R14014 CSoutput.n325 CSoutput.t105 2.82907
R14015 CSoutput.n327 CSoutput.t106 2.82907
R14016 CSoutput.n327 CSoutput.t50 2.82907
R14017 CSoutput.n329 CSoutput.t51 2.82907
R14018 CSoutput.n329 CSoutput.t80 2.82907
R14019 CSoutput.n331 CSoutput.t81 2.82907
R14020 CSoutput.n331 CSoutput.t101 2.82907
R14021 CSoutput.n333 CSoutput.t102 2.82907
R14022 CSoutput.n333 CSoutput.t95 2.82907
R14023 CSoutput.n313 CSoutput.t57 2.82907
R14024 CSoutput.n313 CSoutput.t86 2.82907
R14025 CSoutput.n314 CSoutput.t84 2.82907
R14026 CSoutput.n314 CSoutput.t72 2.82907
R14027 CSoutput.n316 CSoutput.t90 2.82907
R14028 CSoutput.n316 CSoutput.t64 2.82907
R14029 CSoutput.n318 CSoutput.t77 2.82907
R14030 CSoutput.n318 CSoutput.t100 2.82907
R14031 CSoutput.n320 CSoutput.t52 2.82907
R14032 CSoutput.n320 CSoutput.t88 2.82907
R14033 CSoutput.n322 CSoutput.t45 2.82907
R14034 CSoutput.n322 CSoutput.t92 2.82907
R14035 CSoutput.n348 CSoutput.n312 2.75627
R14036 CSoutput.n75 CSoutput.n1 2.45513
R14037 CSoutput.n193 CSoutput.n191 2.251
R14038 CSoutput.n193 CSoutput.n190 2.251
R14039 CSoutput.n193 CSoutput.n189 2.251
R14040 CSoutput.n193 CSoutput.n188 2.251
R14041 CSoutput.n162 CSoutput.n161 2.251
R14042 CSoutput.n162 CSoutput.n160 2.251
R14043 CSoutput.n162 CSoutput.n159 2.251
R14044 CSoutput.n162 CSoutput.n158 2.251
R14045 CSoutput.n235 CSoutput.n234 2.251
R14046 CSoutput.n200 CSoutput.n198 2.251
R14047 CSoutput.n200 CSoutput.n197 2.251
R14048 CSoutput.n200 CSoutput.n196 2.251
R14049 CSoutput.n218 CSoutput.n200 2.251
R14050 CSoutput.n206 CSoutput.n205 2.251
R14051 CSoutput.n206 CSoutput.n204 2.251
R14052 CSoutput.n206 CSoutput.n203 2.251
R14053 CSoutput.n206 CSoutput.n202 2.251
R14054 CSoutput.n232 CSoutput.n172 2.251
R14055 CSoutput.n227 CSoutput.n225 2.251
R14056 CSoutput.n227 CSoutput.n224 2.251
R14057 CSoutput.n227 CSoutput.n223 2.251
R14058 CSoutput.n227 CSoutput.n222 2.251
R14059 CSoutput.n128 CSoutput.n127 2.251
R14060 CSoutput.n128 CSoutput.n126 2.251
R14061 CSoutput.n128 CSoutput.n125 2.251
R14062 CSoutput.n128 CSoutput.n124 2.251
R14063 CSoutput.n245 CSoutput.n244 2.251
R14064 CSoutput.n162 CSoutput.n142 2.2505
R14065 CSoutput.n157 CSoutput.n142 2.2505
R14066 CSoutput.n155 CSoutput.n142 2.2505
R14067 CSoutput.n154 CSoutput.n142 2.2505
R14068 CSoutput.n239 CSoutput.n142 2.2505
R14069 CSoutput.n237 CSoutput.n142 2.2505
R14070 CSoutput.n235 CSoutput.n142 2.2505
R14071 CSoutput.n165 CSoutput.n142 2.2505
R14072 CSoutput.n164 CSoutput.n142 2.2505
R14073 CSoutput.n168 CSoutput.n142 2.2505
R14074 CSoutput.n167 CSoutput.n142 2.2505
R14075 CSoutput.n150 CSoutput.n142 2.2505
R14076 CSoutput.n242 CSoutput.n142 2.2505
R14077 CSoutput.n242 CSoutput.n241 2.2505
R14078 CSoutput.n206 CSoutput.n177 2.2505
R14079 CSoutput.n187 CSoutput.n177 2.2505
R14080 CSoutput.n208 CSoutput.n177 2.2505
R14081 CSoutput.n186 CSoutput.n177 2.2505
R14082 CSoutput.n210 CSoutput.n177 2.2505
R14083 CSoutput.n177 CSoutput.n171 2.2505
R14084 CSoutput.n232 CSoutput.n177 2.2505
R14085 CSoutput.n230 CSoutput.n177 2.2505
R14086 CSoutput.n212 CSoutput.n177 2.2505
R14087 CSoutput.n184 CSoutput.n177 2.2505
R14088 CSoutput.n214 CSoutput.n177 2.2505
R14089 CSoutput.n183 CSoutput.n177 2.2505
R14090 CSoutput.n228 CSoutput.n177 2.2505
R14091 CSoutput.n228 CSoutput.n181 2.2505
R14092 CSoutput.n128 CSoutput.n108 2.2505
R14093 CSoutput.n123 CSoutput.n108 2.2505
R14094 CSoutput.n121 CSoutput.n108 2.2505
R14095 CSoutput.n120 CSoutput.n108 2.2505
R14096 CSoutput.n249 CSoutput.n108 2.2505
R14097 CSoutput.n247 CSoutput.n108 2.2505
R14098 CSoutput.n245 CSoutput.n108 2.2505
R14099 CSoutput.n131 CSoutput.n108 2.2505
R14100 CSoutput.n130 CSoutput.n108 2.2505
R14101 CSoutput.n134 CSoutput.n108 2.2505
R14102 CSoutput.n133 CSoutput.n108 2.2505
R14103 CSoutput.n116 CSoutput.n108 2.2505
R14104 CSoutput.n252 CSoutput.n108 2.2505
R14105 CSoutput.n252 CSoutput.n251 2.2505
R14106 CSoutput.n170 CSoutput.n163 2.25024
R14107 CSoutput.n170 CSoutput.n156 2.25024
R14108 CSoutput.n238 CSoutput.n170 2.25024
R14109 CSoutput.n170 CSoutput.n166 2.25024
R14110 CSoutput.n170 CSoutput.n169 2.25024
R14111 CSoutput.n170 CSoutput.n137 2.25024
R14112 CSoutput.n220 CSoutput.n217 2.25024
R14113 CSoutput.n220 CSoutput.n216 2.25024
R14114 CSoutput.n220 CSoutput.n215 2.25024
R14115 CSoutput.n220 CSoutput.n182 2.25024
R14116 CSoutput.n220 CSoutput.n219 2.25024
R14117 CSoutput.n221 CSoutput.n220 2.25024
R14118 CSoutput.n136 CSoutput.n129 2.25024
R14119 CSoutput.n136 CSoutput.n122 2.25024
R14120 CSoutput.n248 CSoutput.n136 2.25024
R14121 CSoutput.n136 CSoutput.n132 2.25024
R14122 CSoutput.n136 CSoutput.n135 2.25024
R14123 CSoutput.n136 CSoutput.n103 2.25024
R14124 CSoutput.n276 CSoutput.n102 1.95131
R14125 CSoutput.n237 CSoutput.n147 1.50111
R14126 CSoutput.n185 CSoutput.n171 1.50111
R14127 CSoutput.n247 CSoutput.n113 1.50111
R14128 CSoutput.n193 CSoutput.n192 1.501
R14129 CSoutput.n200 CSoutput.n199 1.501
R14130 CSoutput.n227 CSoutput.n226 1.501
R14131 CSoutput.n241 CSoutput.n152 1.12536
R14132 CSoutput.n241 CSoutput.n153 1.12536
R14133 CSoutput.n241 CSoutput.n240 1.12536
R14134 CSoutput.n201 CSoutput.n181 1.12536
R14135 CSoutput.n207 CSoutput.n181 1.12536
R14136 CSoutput.n209 CSoutput.n181 1.12536
R14137 CSoutput.n251 CSoutput.n118 1.12536
R14138 CSoutput.n251 CSoutput.n119 1.12536
R14139 CSoutput.n251 CSoutput.n250 1.12536
R14140 CSoutput.n241 CSoutput.n148 1.12536
R14141 CSoutput.n241 CSoutput.n149 1.12536
R14142 CSoutput.n241 CSoutput.n151 1.12536
R14143 CSoutput.n231 CSoutput.n181 1.12536
R14144 CSoutput.n211 CSoutput.n181 1.12536
R14145 CSoutput.n213 CSoutput.n181 1.12536
R14146 CSoutput.n251 CSoutput.n114 1.12536
R14147 CSoutput.n251 CSoutput.n115 1.12536
R14148 CSoutput.n251 CSoutput.n117 1.12536
R14149 CSoutput.n31 CSoutput.n30 0.669944
R14150 CSoutput.n62 CSoutput.n61 0.669944
R14151 CSoutput.n304 CSoutput.n302 0.573776
R14152 CSoutput.n306 CSoutput.n304 0.573776
R14153 CSoutput.n308 CSoutput.n306 0.573776
R14154 CSoutput.n310 CSoutput.n308 0.573776
R14155 CSoutput.n292 CSoutput.n290 0.573776
R14156 CSoutput.n294 CSoutput.n292 0.573776
R14157 CSoutput.n296 CSoutput.n294 0.573776
R14158 CSoutput.n298 CSoutput.n296 0.573776
R14159 CSoutput.n281 CSoutput.n279 0.573776
R14160 CSoutput.n283 CSoutput.n281 0.573776
R14161 CSoutput.n285 CSoutput.n283 0.573776
R14162 CSoutput.n287 CSoutput.n285 0.573776
R14163 CSoutput.n346 CSoutput.n344 0.573776
R14164 CSoutput.n344 CSoutput.n342 0.573776
R14165 CSoutput.n342 CSoutput.n340 0.573776
R14166 CSoutput.n340 CSoutput.n338 0.573776
R14167 CSoutput.n334 CSoutput.n332 0.573776
R14168 CSoutput.n332 CSoutput.n330 0.573776
R14169 CSoutput.n330 CSoutput.n328 0.573776
R14170 CSoutput.n328 CSoutput.n326 0.573776
R14171 CSoutput.n323 CSoutput.n321 0.573776
R14172 CSoutput.n321 CSoutput.n319 0.573776
R14173 CSoutput.n319 CSoutput.n317 0.573776
R14174 CSoutput.n317 CSoutput.n315 0.573776
R14175 CSoutput.n349 CSoutput.n252 0.53442
R14176 CSoutput.n272 CSoutput.n270 0.358259
R14177 CSoutput.n274 CSoutput.n272 0.358259
R14178 CSoutput.n264 CSoutput.n262 0.358259
R14179 CSoutput.n266 CSoutput.n264 0.358259
R14180 CSoutput.n257 CSoutput.n255 0.358259
R14181 CSoutput.n259 CSoutput.n257 0.358259
R14182 CSoutput.n100 CSoutput.n98 0.358259
R14183 CSoutput.n98 CSoutput.n96 0.358259
R14184 CSoutput.n92 CSoutput.n90 0.358259
R14185 CSoutput.n90 CSoutput.n88 0.358259
R14186 CSoutput.n85 CSoutput.n83 0.358259
R14187 CSoutput.n83 CSoutput.n81 0.358259
R14188 CSoutput.n21 CSoutput.n20 0.169105
R14189 CSoutput.n21 CSoutput.n16 0.169105
R14190 CSoutput.n26 CSoutput.n16 0.169105
R14191 CSoutput.n27 CSoutput.n26 0.169105
R14192 CSoutput.n27 CSoutput.n14 0.169105
R14193 CSoutput.n32 CSoutput.n14 0.169105
R14194 CSoutput.n33 CSoutput.n32 0.169105
R14195 CSoutput.n34 CSoutput.n33 0.169105
R14196 CSoutput.n34 CSoutput.n12 0.169105
R14197 CSoutput.n39 CSoutput.n12 0.169105
R14198 CSoutput.n40 CSoutput.n39 0.169105
R14199 CSoutput.n40 CSoutput.n10 0.169105
R14200 CSoutput.n45 CSoutput.n10 0.169105
R14201 CSoutput.n46 CSoutput.n45 0.169105
R14202 CSoutput.n47 CSoutput.n46 0.169105
R14203 CSoutput.n47 CSoutput.n8 0.169105
R14204 CSoutput.n52 CSoutput.n8 0.169105
R14205 CSoutput.n53 CSoutput.n52 0.169105
R14206 CSoutput.n53 CSoutput.n6 0.169105
R14207 CSoutput.n58 CSoutput.n6 0.169105
R14208 CSoutput.n59 CSoutput.n58 0.169105
R14209 CSoutput.n60 CSoutput.n59 0.169105
R14210 CSoutput.n60 CSoutput.n4 0.169105
R14211 CSoutput.n66 CSoutput.n4 0.169105
R14212 CSoutput.n67 CSoutput.n66 0.169105
R14213 CSoutput.n68 CSoutput.n67 0.169105
R14214 CSoutput.n68 CSoutput.n2 0.169105
R14215 CSoutput.n73 CSoutput.n2 0.169105
R14216 CSoutput.n74 CSoutput.n73 0.169105
R14217 CSoutput.n74 CSoutput.n0 0.169105
R14218 CSoutput.n78 CSoutput.n0 0.169105
R14219 CSoutput.n195 CSoutput.n194 0.0910737
R14220 CSoutput.n246 CSoutput.n243 0.0723685
R14221 CSoutput.n200 CSoutput.n195 0.0522944
R14222 CSoutput.n243 CSoutput.n242 0.0499135
R14223 CSoutput.n194 CSoutput.n193 0.0499135
R14224 CSoutput.n228 CSoutput.n227 0.0464294
R14225 CSoutput.n236 CSoutput.n233 0.0391444
R14226 CSoutput.n195 CSoutput.t131 0.023435
R14227 CSoutput.n243 CSoutput.t130 0.02262
R14228 CSoutput.n194 CSoutput.t136 0.02262
R14229 CSoutput CSoutput.n349 0.0052
R14230 CSoutput.n165 CSoutput.n148 0.00365111
R14231 CSoutput.n168 CSoutput.n149 0.00365111
R14232 CSoutput.n151 CSoutput.n150 0.00365111
R14233 CSoutput.n193 CSoutput.n152 0.00365111
R14234 CSoutput.n157 CSoutput.n153 0.00365111
R14235 CSoutput.n240 CSoutput.n154 0.00365111
R14236 CSoutput.n231 CSoutput.n230 0.00365111
R14237 CSoutput.n211 CSoutput.n184 0.00365111
R14238 CSoutput.n213 CSoutput.n183 0.00365111
R14239 CSoutput.n201 CSoutput.n200 0.00365111
R14240 CSoutput.n207 CSoutput.n187 0.00365111
R14241 CSoutput.n209 CSoutput.n186 0.00365111
R14242 CSoutput.n131 CSoutput.n114 0.00365111
R14243 CSoutput.n134 CSoutput.n115 0.00365111
R14244 CSoutput.n117 CSoutput.n116 0.00365111
R14245 CSoutput.n227 CSoutput.n118 0.00365111
R14246 CSoutput.n123 CSoutput.n119 0.00365111
R14247 CSoutput.n250 CSoutput.n120 0.00365111
R14248 CSoutput.n162 CSoutput.n152 0.00340054
R14249 CSoutput.n155 CSoutput.n153 0.00340054
R14250 CSoutput.n240 CSoutput.n239 0.00340054
R14251 CSoutput.n235 CSoutput.n148 0.00340054
R14252 CSoutput.n164 CSoutput.n149 0.00340054
R14253 CSoutput.n167 CSoutput.n151 0.00340054
R14254 CSoutput.n206 CSoutput.n201 0.00340054
R14255 CSoutput.n208 CSoutput.n207 0.00340054
R14256 CSoutput.n210 CSoutput.n209 0.00340054
R14257 CSoutput.n232 CSoutput.n231 0.00340054
R14258 CSoutput.n212 CSoutput.n211 0.00340054
R14259 CSoutput.n214 CSoutput.n213 0.00340054
R14260 CSoutput.n128 CSoutput.n118 0.00340054
R14261 CSoutput.n121 CSoutput.n119 0.00340054
R14262 CSoutput.n250 CSoutput.n249 0.00340054
R14263 CSoutput.n245 CSoutput.n114 0.00340054
R14264 CSoutput.n130 CSoutput.n115 0.00340054
R14265 CSoutput.n133 CSoutput.n117 0.00340054
R14266 CSoutput.n163 CSoutput.n157 0.00252698
R14267 CSoutput.n156 CSoutput.n154 0.00252698
R14268 CSoutput.n238 CSoutput.n237 0.00252698
R14269 CSoutput.n166 CSoutput.n164 0.00252698
R14270 CSoutput.n169 CSoutput.n167 0.00252698
R14271 CSoutput.n242 CSoutput.n137 0.00252698
R14272 CSoutput.n163 CSoutput.n162 0.00252698
R14273 CSoutput.n156 CSoutput.n155 0.00252698
R14274 CSoutput.n239 CSoutput.n238 0.00252698
R14275 CSoutput.n166 CSoutput.n165 0.00252698
R14276 CSoutput.n169 CSoutput.n168 0.00252698
R14277 CSoutput.n150 CSoutput.n137 0.00252698
R14278 CSoutput.n217 CSoutput.n187 0.00252698
R14279 CSoutput.n216 CSoutput.n186 0.00252698
R14280 CSoutput.n215 CSoutput.n171 0.00252698
R14281 CSoutput.n212 CSoutput.n182 0.00252698
R14282 CSoutput.n219 CSoutput.n214 0.00252698
R14283 CSoutput.n228 CSoutput.n221 0.00252698
R14284 CSoutput.n217 CSoutput.n206 0.00252698
R14285 CSoutput.n216 CSoutput.n208 0.00252698
R14286 CSoutput.n215 CSoutput.n210 0.00252698
R14287 CSoutput.n230 CSoutput.n182 0.00252698
R14288 CSoutput.n219 CSoutput.n184 0.00252698
R14289 CSoutput.n221 CSoutput.n183 0.00252698
R14290 CSoutput.n129 CSoutput.n123 0.00252698
R14291 CSoutput.n122 CSoutput.n120 0.00252698
R14292 CSoutput.n248 CSoutput.n247 0.00252698
R14293 CSoutput.n132 CSoutput.n130 0.00252698
R14294 CSoutput.n135 CSoutput.n133 0.00252698
R14295 CSoutput.n252 CSoutput.n103 0.00252698
R14296 CSoutput.n129 CSoutput.n128 0.00252698
R14297 CSoutput.n122 CSoutput.n121 0.00252698
R14298 CSoutput.n249 CSoutput.n248 0.00252698
R14299 CSoutput.n132 CSoutput.n131 0.00252698
R14300 CSoutput.n135 CSoutput.n134 0.00252698
R14301 CSoutput.n116 CSoutput.n103 0.00252698
R14302 CSoutput.n237 CSoutput.n236 0.0020275
R14303 CSoutput.n236 CSoutput.n235 0.0020275
R14304 CSoutput.n233 CSoutput.n171 0.0020275
R14305 CSoutput.n233 CSoutput.n232 0.0020275
R14306 CSoutput.n247 CSoutput.n246 0.0020275
R14307 CSoutput.n246 CSoutput.n245 0.0020275
R14308 CSoutput.n147 CSoutput.n146 0.00166668
R14309 CSoutput.n229 CSoutput.n185 0.00166668
R14310 CSoutput.n113 CSoutput.n112 0.00166668
R14311 CSoutput.n251 CSoutput.n113 0.00133328
R14312 CSoutput.n185 CSoutput.n181 0.00133328
R14313 CSoutput.n241 CSoutput.n147 0.00133328
R14314 CSoutput.n244 CSoutput.n136 0.001
R14315 CSoutput.n222 CSoutput.n136 0.001
R14316 CSoutput.n124 CSoutput.n104 0.001
R14317 CSoutput.n223 CSoutput.n104 0.001
R14318 CSoutput.n125 CSoutput.n105 0.001
R14319 CSoutput.n224 CSoutput.n105 0.001
R14320 CSoutput.n126 CSoutput.n106 0.001
R14321 CSoutput.n225 CSoutput.n106 0.001
R14322 CSoutput.n127 CSoutput.n107 0.001
R14323 CSoutput.n226 CSoutput.n107 0.001
R14324 CSoutput.n220 CSoutput.n172 0.001
R14325 CSoutput.n220 CSoutput.n218 0.001
R14326 CSoutput.n202 CSoutput.n173 0.001
R14327 CSoutput.n196 CSoutput.n173 0.001
R14328 CSoutput.n203 CSoutput.n174 0.001
R14329 CSoutput.n197 CSoutput.n174 0.001
R14330 CSoutput.n204 CSoutput.n175 0.001
R14331 CSoutput.n198 CSoutput.n175 0.001
R14332 CSoutput.n205 CSoutput.n176 0.001
R14333 CSoutput.n199 CSoutput.n176 0.001
R14334 CSoutput.n234 CSoutput.n170 0.001
R14335 CSoutput.n188 CSoutput.n170 0.001
R14336 CSoutput.n158 CSoutput.n138 0.001
R14337 CSoutput.n189 CSoutput.n138 0.001
R14338 CSoutput.n159 CSoutput.n139 0.001
R14339 CSoutput.n190 CSoutput.n139 0.001
R14340 CSoutput.n160 CSoutput.n140 0.001
R14341 CSoutput.n191 CSoutput.n140 0.001
R14342 CSoutput.n161 CSoutput.n141 0.001
R14343 CSoutput.n192 CSoutput.n141 0.001
R14344 CSoutput.n192 CSoutput.n142 0.001
R14345 CSoutput.n191 CSoutput.n143 0.001
R14346 CSoutput.n190 CSoutput.n144 0.001
R14347 CSoutput.n189 CSoutput.t127 0.001
R14348 CSoutput.n188 CSoutput.n145 0.001
R14349 CSoutput.n161 CSoutput.n143 0.001
R14350 CSoutput.n160 CSoutput.n144 0.001
R14351 CSoutput.n159 CSoutput.t127 0.001
R14352 CSoutput.n158 CSoutput.n145 0.001
R14353 CSoutput.n234 CSoutput.n146 0.001
R14354 CSoutput.n199 CSoutput.n177 0.001
R14355 CSoutput.n198 CSoutput.n178 0.001
R14356 CSoutput.n197 CSoutput.n179 0.001
R14357 CSoutput.n196 CSoutput.t120 0.001
R14358 CSoutput.n218 CSoutput.n180 0.001
R14359 CSoutput.n205 CSoutput.n178 0.001
R14360 CSoutput.n204 CSoutput.n179 0.001
R14361 CSoutput.n203 CSoutput.t120 0.001
R14362 CSoutput.n202 CSoutput.n180 0.001
R14363 CSoutput.n229 CSoutput.n172 0.001
R14364 CSoutput.n226 CSoutput.n108 0.001
R14365 CSoutput.n225 CSoutput.n109 0.001
R14366 CSoutput.n224 CSoutput.n110 0.001
R14367 CSoutput.n223 CSoutput.t140 0.001
R14368 CSoutput.n222 CSoutput.n111 0.001
R14369 CSoutput.n127 CSoutput.n109 0.001
R14370 CSoutput.n126 CSoutput.n110 0.001
R14371 CSoutput.n125 CSoutput.t140 0.001
R14372 CSoutput.n124 CSoutput.n111 0.001
R14373 CSoutput.n244 CSoutput.n112 0.001
R14374 plus.n43 plus.t18 322.512
R14375 plus.n9 plus.t13 322.512
R14376 plus.n42 plus.t17 297.12
R14377 plus.n46 plus.t22 297.12
R14378 plus.n48 plus.t21 297.12
R14379 plus.n52 plus.t23 297.12
R14380 plus.n54 plus.t8 297.12
R14381 plus.n58 plus.t7 297.12
R14382 plus.n60 plus.t12 297.12
R14383 plus.n64 plus.t10 297.12
R14384 plus.n66 plus.t24 297.12
R14385 plus.n32 plus.t14 297.12
R14386 plus.n30 plus.t15 297.12
R14387 plus.n2 plus.t9 297.12
R14388 plus.n24 plus.t5 297.12
R14389 plus.n4 plus.t6 297.12
R14390 plus.n18 plus.t19 297.12
R14391 plus.n6 plus.t20 297.12
R14392 plus.n12 plus.t16 297.12
R14393 plus.n8 plus.t11 297.12
R14394 plus.n70 plus.t0 243.97
R14395 plus.n70 plus.n69 223.454
R14396 plus.n72 plus.n71 223.454
R14397 plus.n67 plus.n66 161.3
R14398 plus.n65 plus.n34 161.3
R14399 plus.n64 plus.n63 161.3
R14400 plus.n62 plus.n35 161.3
R14401 plus.n61 plus.n60 161.3
R14402 plus.n59 plus.n36 161.3
R14403 plus.n58 plus.n57 161.3
R14404 plus.n56 plus.n37 161.3
R14405 plus.n55 plus.n54 161.3
R14406 plus.n53 plus.n38 161.3
R14407 plus.n52 plus.n51 161.3
R14408 plus.n50 plus.n39 161.3
R14409 plus.n49 plus.n48 161.3
R14410 plus.n47 plus.n40 161.3
R14411 plus.n46 plus.n45 161.3
R14412 plus.n44 plus.n41 161.3
R14413 plus.n11 plus.n10 161.3
R14414 plus.n12 plus.n7 161.3
R14415 plus.n14 plus.n13 161.3
R14416 plus.n15 plus.n6 161.3
R14417 plus.n17 plus.n16 161.3
R14418 plus.n18 plus.n5 161.3
R14419 plus.n20 plus.n19 161.3
R14420 plus.n21 plus.n4 161.3
R14421 plus.n23 plus.n22 161.3
R14422 plus.n24 plus.n3 161.3
R14423 plus.n26 plus.n25 161.3
R14424 plus.n27 plus.n2 161.3
R14425 plus.n29 plus.n28 161.3
R14426 plus.n30 plus.n1 161.3
R14427 plus.n31 plus.n0 161.3
R14428 plus.n33 plus.n32 161.3
R14429 plus.n44 plus.n43 45.0031
R14430 plus.n10 plus.n9 45.0031
R14431 plus.n66 plus.n65 41.6278
R14432 plus.n32 plus.n31 41.6278
R14433 plus.n42 plus.n41 37.246
R14434 plus.n64 plus.n35 37.246
R14435 plus.n30 plus.n29 37.246
R14436 plus.n11 plus.n8 37.246
R14437 plus.n47 plus.n46 32.8641
R14438 plus.n60 plus.n59 32.8641
R14439 plus.n25 plus.n2 32.8641
R14440 plus.n13 plus.n12 32.8641
R14441 plus.n68 plus.n67 31.6047
R14442 plus.n48 plus.n39 28.4823
R14443 plus.n58 plus.n37 28.4823
R14444 plus.n24 plus.n23 28.4823
R14445 plus.n17 plus.n6 28.4823
R14446 plus.n53 plus.n52 24.1005
R14447 plus.n54 plus.n53 24.1005
R14448 plus.n19 plus.n4 24.1005
R14449 plus.n19 plus.n18 24.1005
R14450 plus.n69 plus.t4 19.8005
R14451 plus.n69 plus.t2 19.8005
R14452 plus.n71 plus.t1 19.8005
R14453 plus.n71 plus.t3 19.8005
R14454 plus.n52 plus.n39 19.7187
R14455 plus.n54 plus.n37 19.7187
R14456 plus.n23 plus.n4 19.7187
R14457 plus.n18 plus.n17 19.7187
R14458 plus.n43 plus.n42 15.6319
R14459 plus.n9 plus.n8 15.6319
R14460 plus.n48 plus.n47 15.3369
R14461 plus.n59 plus.n58 15.3369
R14462 plus.n25 plus.n24 15.3369
R14463 plus.n13 plus.n6 15.3369
R14464 plus plus.n73 14.1121
R14465 plus.n68 plus.n33 11.866
R14466 plus.n46 plus.n41 10.955
R14467 plus.n60 plus.n35 10.955
R14468 plus.n29 plus.n2 10.955
R14469 plus.n12 plus.n11 10.955
R14470 plus.n65 plus.n64 6.57323
R14471 plus.n31 plus.n30 6.57323
R14472 plus.n73 plus.n72 5.40567
R14473 plus.n73 plus.n68 1.188
R14474 plus.n72 plus.n70 0.716017
R14475 plus.n45 plus.n44 0.189894
R14476 plus.n45 plus.n40 0.189894
R14477 plus.n49 plus.n40 0.189894
R14478 plus.n50 plus.n49 0.189894
R14479 plus.n51 plus.n50 0.189894
R14480 plus.n51 plus.n38 0.189894
R14481 plus.n55 plus.n38 0.189894
R14482 plus.n56 plus.n55 0.189894
R14483 plus.n57 plus.n56 0.189894
R14484 plus.n57 plus.n36 0.189894
R14485 plus.n61 plus.n36 0.189894
R14486 plus.n62 plus.n61 0.189894
R14487 plus.n63 plus.n62 0.189894
R14488 plus.n63 plus.n34 0.189894
R14489 plus.n67 plus.n34 0.189894
R14490 plus.n33 plus.n0 0.189894
R14491 plus.n1 plus.n0 0.189894
R14492 plus.n28 plus.n1 0.189894
R14493 plus.n28 plus.n27 0.189894
R14494 plus.n27 plus.n26 0.189894
R14495 plus.n26 plus.n3 0.189894
R14496 plus.n22 plus.n3 0.189894
R14497 plus.n22 plus.n21 0.189894
R14498 plus.n21 plus.n20 0.189894
R14499 plus.n20 plus.n5 0.189894
R14500 plus.n16 plus.n5 0.189894
R14501 plus.n16 plus.n15 0.189894
R14502 plus.n15 plus.n14 0.189894
R14503 plus.n14 plus.n7 0.189894
R14504 plus.n10 plus.n7 0.189894
R14505 a_n2903_n3924.n8 a_n2903_n3924.t43 214.944
R14506 a_n2903_n3924.n11 a_n2903_n3924.t46 214.413
R14507 a_n2903_n3924.n11 a_n2903_n3924.t47 214.321
R14508 a_n2903_n3924.n10 a_n2903_n3924.t24 214.321
R14509 a_n2903_n3924.n10 a_n2903_n3924.t23 214.321
R14510 a_n2903_n3924.n9 a_n2903_n3924.t22 214.321
R14511 a_n2903_n3924.n9 a_n2903_n3924.t41 214.321
R14512 a_n2903_n3924.n8 a_n2903_n3924.t42 214.321
R14513 a_n2903_n3924.n5 a_n2903_n3924.t4 55.8337
R14514 a_n2903_n3924.n5 a_n2903_n3924.t21 55.8337
R14515 a_n2903_n3924.n7 a_n2903_n3924.t25 55.8337
R14516 a_n2903_n3924.n4 a_n2903_n3924.t10 55.8335
R14517 a_n2903_n3924.n0 a_n2903_n3924.t37 55.8335
R14518 a_n2903_n3924.n1 a_n2903_n3924.t28 55.8335
R14519 a_n2903_n3924.n1 a_n2903_n3924.t9 55.8335
R14520 a_n2903_n3924.n3 a_n2903_n3924.t14 55.8335
R14521 a_n2903_n3924.n29 a_n2903_n3924.n3 53.0054
R14522 a_n2903_n3924.n4 a_n2903_n3924.n12 53.0052
R14523 a_n2903_n3924.n5 a_n2903_n3924.n13 53.0052
R14524 a_n2903_n3924.n5 a_n2903_n3924.n14 53.0052
R14525 a_n2903_n3924.n5 a_n2903_n3924.n15 53.0052
R14526 a_n2903_n3924.n6 a_n2903_n3924.n16 53.0052
R14527 a_n2903_n3924.n6 a_n2903_n3924.n17 53.0052
R14528 a_n2903_n3924.n7 a_n2903_n3924.n18 53.0052
R14529 a_n2903_n3924.n7 a_n2903_n3924.n19 53.0052
R14530 a_n2903_n3924.n0 a_n2903_n3924.n22 53.0051
R14531 a_n2903_n3924.n1 a_n2903_n3924.n23 53.0051
R14532 a_n2903_n3924.n1 a_n2903_n3924.n24 53.0051
R14533 a_n2903_n3924.n1 a_n2903_n3924.n25 53.0051
R14534 a_n2903_n3924.n2 a_n2903_n3924.n26 53.0051
R14535 a_n2903_n3924.n2 a_n2903_n3924.n27 53.0051
R14536 a_n2903_n3924.n3 a_n2903_n3924.n28 53.0051
R14537 a_n2903_n3924.n20 a_n2903_n3924.n7 12.1986
R14538 a_n2903_n3924.n21 a_n2903_n3924.n4 12.1986
R14539 a_n2903_n3924.n20 a_n2903_n3924.n3 5.11903
R14540 a_n2903_n3924.n0 a_n2903_n3924.n21 5.11903
R14541 a_n2903_n3924.n22 a_n2903_n3924.t44 2.82907
R14542 a_n2903_n3924.n22 a_n2903_n3924.t36 2.82907
R14543 a_n2903_n3924.n23 a_n2903_n3924.t29 2.82907
R14544 a_n2903_n3924.n23 a_n2903_n3924.t30 2.82907
R14545 a_n2903_n3924.n24 a_n2903_n3924.t27 2.82907
R14546 a_n2903_n3924.n24 a_n2903_n3924.t38 2.82907
R14547 a_n2903_n3924.n25 a_n2903_n3924.t39 2.82907
R14548 a_n2903_n3924.n25 a_n2903_n3924.t26 2.82907
R14549 a_n2903_n3924.n26 a_n2903_n3924.t8 2.82907
R14550 a_n2903_n3924.n26 a_n2903_n3924.t5 2.82907
R14551 a_n2903_n3924.n27 a_n2903_n3924.t18 2.82907
R14552 a_n2903_n3924.n27 a_n2903_n3924.t13 2.82907
R14553 a_n2903_n3924.n28 a_n2903_n3924.t17 2.82907
R14554 a_n2903_n3924.n28 a_n2903_n3924.t16 2.82907
R14555 a_n2903_n3924.n12 a_n2903_n3924.t1 2.82907
R14556 a_n2903_n3924.n12 a_n2903_n3924.t12 2.82907
R14557 a_n2903_n3924.n13 a_n2903_n3924.t7 2.82907
R14558 a_n2903_n3924.n13 a_n2903_n3924.t11 2.82907
R14559 a_n2903_n3924.n14 a_n2903_n3924.t19 2.82907
R14560 a_n2903_n3924.n14 a_n2903_n3924.t6 2.82907
R14561 a_n2903_n3924.n15 a_n2903_n3924.t2 2.82907
R14562 a_n2903_n3924.n15 a_n2903_n3924.t15 2.82907
R14563 a_n2903_n3924.n16 a_n2903_n3924.t40 2.82907
R14564 a_n2903_n3924.n16 a_n2903_n3924.t31 2.82907
R14565 a_n2903_n3924.n17 a_n2903_n3924.t33 2.82907
R14566 a_n2903_n3924.n17 a_n2903_n3924.t35 2.82907
R14567 a_n2903_n3924.n18 a_n2903_n3924.t34 2.82907
R14568 a_n2903_n3924.n18 a_n2903_n3924.t20 2.82907
R14569 a_n2903_n3924.n19 a_n2903_n3924.t32 2.82907
R14570 a_n2903_n3924.n19 a_n2903_n3924.t45 2.82907
R14571 a_n2903_n3924.t0 a_n2903_n3924.n29 2.82907
R14572 a_n2903_n3924.n29 a_n2903_n3924.t3 2.82907
R14573 a_n2903_n3924.n8 a_n2903_n3924.n20 1.95694
R14574 a_n2903_n3924.n21 a_n2903_n3924.n11 1.95694
R14575 a_n2903_n3924.n7 a_n2903_n3924.n6 1.77636
R14576 a_n2903_n3924.n5 a_n2903_n3924.n4 1.77636
R14577 a_n2903_n3924.n3 a_n2903_n3924.n2 1.77636
R14578 a_n2903_n3924.n1 a_n2903_n3924.n0 1.77636
R14579 a_n2903_n3924.n9 a_n2903_n3924.n8 1.39367
R14580 a_n2903_n3924.n10 a_n2903_n3924.n9 1.34352
R14581 a_n2903_n3924.n11 a_n2903_n3924.n10 1.25123
R14582 a_n2903_n3924.n2 a_n2903_n3924.n1 1.12334
R14583 a_n2903_n3924.n6 a_n2903_n3924.n5 1.12334
R14584 a_n5644_8799.n85 a_n5644_8799.t65 485.149
R14585 a_n5644_8799.n107 a_n5644_8799.t68 485.149
R14586 a_n5644_8799.n130 a_n5644_8799.t34 485.149
R14587 a_n5644_8799.n17 a_n5644_8799.t49 485.149
R14588 a_n5644_8799.n39 a_n5644_8799.t54 485.149
R14589 a_n5644_8799.n62 a_n5644_8799.t35 485.149
R14590 a_n5644_8799.n100 a_n5644_8799.t56 464.166
R14591 a_n5644_8799.n99 a_n5644_8799.t55 464.166
R14592 a_n5644_8799.n81 a_n5644_8799.t42 464.166
R14593 a_n5644_8799.n93 a_n5644_8799.t72 464.166
R14594 a_n5644_8799.n92 a_n5644_8799.t57 464.166
R14595 a_n5644_8799.n84 a_n5644_8799.t47 464.166
R14596 a_n5644_8799.n86 a_n5644_8799.t74 464.166
R14597 a_n5644_8799.n122 a_n5644_8799.t60 464.166
R14598 a_n5644_8799.n121 a_n5644_8799.t59 464.166
R14599 a_n5644_8799.n103 a_n5644_8799.t51 464.166
R14600 a_n5644_8799.n115 a_n5644_8799.t76 464.166
R14601 a_n5644_8799.n114 a_n5644_8799.t63 464.166
R14602 a_n5644_8799.n106 a_n5644_8799.t52 464.166
R14603 a_n5644_8799.n108 a_n5644_8799.t32 464.166
R14604 a_n5644_8799.n145 a_n5644_8799.t78 464.166
R14605 a_n5644_8799.n144 a_n5644_8799.t40 464.166
R14606 a_n5644_8799.n126 a_n5644_8799.t61 464.166
R14607 a_n5644_8799.n138 a_n5644_8799.t33 464.166
R14608 a_n5644_8799.n137 a_n5644_8799.t69 464.166
R14609 a_n5644_8799.n129 a_n5644_8799.t46 464.166
R14610 a_n5644_8799.n131 a_n5644_8799.t66 464.166
R14611 a_n5644_8799.n18 a_n5644_8799.t58 464.166
R14612 a_n5644_8799.n20 a_n5644_8799.t73 464.166
R14613 a_n5644_8799.n24 a_n5644_8799.t38 464.166
R14614 a_n5644_8799.n25 a_n5644_8799.t48 464.166
R14615 a_n5644_8799.n13 a_n5644_8799.t71 464.166
R14616 a_n5644_8799.n31 a_n5644_8799.t37 464.166
R14617 a_n5644_8799.n32 a_n5644_8799.t36 464.166
R14618 a_n5644_8799.n40 a_n5644_8799.t64 464.166
R14619 a_n5644_8799.n42 a_n5644_8799.t77 464.166
R14620 a_n5644_8799.n46 a_n5644_8799.t45 464.166
R14621 a_n5644_8799.n47 a_n5644_8799.t53 464.166
R14622 a_n5644_8799.n35 a_n5644_8799.t75 464.166
R14623 a_n5644_8799.n53 a_n5644_8799.t41 464.166
R14624 a_n5644_8799.n54 a_n5644_8799.t43 464.166
R14625 a_n5644_8799.n63 a_n5644_8799.t67 464.166
R14626 a_n5644_8799.n65 a_n5644_8799.t44 464.166
R14627 a_n5644_8799.n69 a_n5644_8799.t70 464.166
R14628 a_n5644_8799.n70 a_n5644_8799.t50 464.166
R14629 a_n5644_8799.n58 a_n5644_8799.t62 464.166
R14630 a_n5644_8799.n76 a_n5644_8799.t39 464.166
R14631 a_n5644_8799.n77 a_n5644_8799.t79 464.166
R14632 a_n5644_8799.n88 a_n5644_8799.n87 161.3
R14633 a_n5644_8799.n89 a_n5644_8799.n84 161.3
R14634 a_n5644_8799.n91 a_n5644_8799.n90 161.3
R14635 a_n5644_8799.n92 a_n5644_8799.n83 161.3
R14636 a_n5644_8799.n93 a_n5644_8799.n82 161.3
R14637 a_n5644_8799.n95 a_n5644_8799.n94 161.3
R14638 a_n5644_8799.n96 a_n5644_8799.n81 161.3
R14639 a_n5644_8799.n98 a_n5644_8799.n97 161.3
R14640 a_n5644_8799.n99 a_n5644_8799.n80 161.3
R14641 a_n5644_8799.n101 a_n5644_8799.n100 161.3
R14642 a_n5644_8799.n110 a_n5644_8799.n109 161.3
R14643 a_n5644_8799.n111 a_n5644_8799.n106 161.3
R14644 a_n5644_8799.n113 a_n5644_8799.n112 161.3
R14645 a_n5644_8799.n114 a_n5644_8799.n105 161.3
R14646 a_n5644_8799.n115 a_n5644_8799.n104 161.3
R14647 a_n5644_8799.n117 a_n5644_8799.n116 161.3
R14648 a_n5644_8799.n118 a_n5644_8799.n103 161.3
R14649 a_n5644_8799.n120 a_n5644_8799.n119 161.3
R14650 a_n5644_8799.n121 a_n5644_8799.n102 161.3
R14651 a_n5644_8799.n123 a_n5644_8799.n122 161.3
R14652 a_n5644_8799.n133 a_n5644_8799.n132 161.3
R14653 a_n5644_8799.n134 a_n5644_8799.n129 161.3
R14654 a_n5644_8799.n136 a_n5644_8799.n135 161.3
R14655 a_n5644_8799.n137 a_n5644_8799.n128 161.3
R14656 a_n5644_8799.n138 a_n5644_8799.n127 161.3
R14657 a_n5644_8799.n140 a_n5644_8799.n139 161.3
R14658 a_n5644_8799.n141 a_n5644_8799.n126 161.3
R14659 a_n5644_8799.n143 a_n5644_8799.n142 161.3
R14660 a_n5644_8799.n144 a_n5644_8799.n125 161.3
R14661 a_n5644_8799.n146 a_n5644_8799.n145 161.3
R14662 a_n5644_8799.n33 a_n5644_8799.n32 161.3
R14663 a_n5644_8799.n31 a_n5644_8799.n12 161.3
R14664 a_n5644_8799.n30 a_n5644_8799.n29 161.3
R14665 a_n5644_8799.n28 a_n5644_8799.n13 161.3
R14666 a_n5644_8799.n27 a_n5644_8799.n26 161.3
R14667 a_n5644_8799.n25 a_n5644_8799.n14 161.3
R14668 a_n5644_8799.n24 a_n5644_8799.n23 161.3
R14669 a_n5644_8799.n22 a_n5644_8799.n15 161.3
R14670 a_n5644_8799.n21 a_n5644_8799.n20 161.3
R14671 a_n5644_8799.n19 a_n5644_8799.n16 161.3
R14672 a_n5644_8799.n55 a_n5644_8799.n54 161.3
R14673 a_n5644_8799.n53 a_n5644_8799.n34 161.3
R14674 a_n5644_8799.n52 a_n5644_8799.n51 161.3
R14675 a_n5644_8799.n50 a_n5644_8799.n35 161.3
R14676 a_n5644_8799.n49 a_n5644_8799.n48 161.3
R14677 a_n5644_8799.n47 a_n5644_8799.n36 161.3
R14678 a_n5644_8799.n46 a_n5644_8799.n45 161.3
R14679 a_n5644_8799.n44 a_n5644_8799.n37 161.3
R14680 a_n5644_8799.n43 a_n5644_8799.n42 161.3
R14681 a_n5644_8799.n41 a_n5644_8799.n38 161.3
R14682 a_n5644_8799.n78 a_n5644_8799.n77 161.3
R14683 a_n5644_8799.n76 a_n5644_8799.n57 161.3
R14684 a_n5644_8799.n75 a_n5644_8799.n74 161.3
R14685 a_n5644_8799.n73 a_n5644_8799.n58 161.3
R14686 a_n5644_8799.n72 a_n5644_8799.n71 161.3
R14687 a_n5644_8799.n70 a_n5644_8799.n59 161.3
R14688 a_n5644_8799.n69 a_n5644_8799.n68 161.3
R14689 a_n5644_8799.n67 a_n5644_8799.n60 161.3
R14690 a_n5644_8799.n66 a_n5644_8799.n65 161.3
R14691 a_n5644_8799.n64 a_n5644_8799.n61 161.3
R14692 a_n5644_8799.n8 a_n5644_8799.n6 98.9633
R14693 a_n5644_8799.n3 a_n5644_8799.n1 98.9631
R14694 a_n5644_8799.n10 a_n5644_8799.n9 98.6055
R14695 a_n5644_8799.n8 a_n5644_8799.n7 98.6055
R14696 a_n5644_8799.n3 a_n5644_8799.n2 98.6055
R14697 a_n5644_8799.n5 a_n5644_8799.n4 98.6055
R14698 a_n5644_8799.n152 a_n5644_8799.n150 81.3764
R14699 a_n5644_8799.n161 a_n5644_8799.n159 81.3764
R14700 a_n5644_8799.n164 a_n5644_8799.n0 81.3764
R14701 a_n5644_8799.n165 a_n5644_8799.n164 80.9326
R14702 a_n5644_8799.n158 a_n5644_8799.n157 80.9324
R14703 a_n5644_8799.n156 a_n5644_8799.n155 80.9324
R14704 a_n5644_8799.n154 a_n5644_8799.n153 80.9324
R14705 a_n5644_8799.n152 a_n5644_8799.n151 80.9324
R14706 a_n5644_8799.n161 a_n5644_8799.n160 80.9324
R14707 a_n5644_8799.n163 a_n5644_8799.n162 80.9324
R14708 a_n5644_8799.n88 a_n5644_8799.n85 70.4033
R14709 a_n5644_8799.n110 a_n5644_8799.n107 70.4033
R14710 a_n5644_8799.n133 a_n5644_8799.n130 70.4033
R14711 a_n5644_8799.n17 a_n5644_8799.n16 70.4033
R14712 a_n5644_8799.n39 a_n5644_8799.n38 70.4033
R14713 a_n5644_8799.n62 a_n5644_8799.n61 70.4033
R14714 a_n5644_8799.n100 a_n5644_8799.n99 48.2005
R14715 a_n5644_8799.n93 a_n5644_8799.n92 48.2005
R14716 a_n5644_8799.n122 a_n5644_8799.n121 48.2005
R14717 a_n5644_8799.n115 a_n5644_8799.n114 48.2005
R14718 a_n5644_8799.n145 a_n5644_8799.n144 48.2005
R14719 a_n5644_8799.n138 a_n5644_8799.n137 48.2005
R14720 a_n5644_8799.n25 a_n5644_8799.n24 48.2005
R14721 a_n5644_8799.n32 a_n5644_8799.n31 48.2005
R14722 a_n5644_8799.n47 a_n5644_8799.n46 48.2005
R14723 a_n5644_8799.n54 a_n5644_8799.n53 48.2005
R14724 a_n5644_8799.n70 a_n5644_8799.n69 48.2005
R14725 a_n5644_8799.n77 a_n5644_8799.n76 48.2005
R14726 a_n5644_8799.n98 a_n5644_8799.n81 37.246
R14727 a_n5644_8799.n87 a_n5644_8799.n84 37.246
R14728 a_n5644_8799.n120 a_n5644_8799.n103 37.246
R14729 a_n5644_8799.n109 a_n5644_8799.n106 37.246
R14730 a_n5644_8799.n143 a_n5644_8799.n126 37.246
R14731 a_n5644_8799.n132 a_n5644_8799.n129 37.246
R14732 a_n5644_8799.n20 a_n5644_8799.n19 37.246
R14733 a_n5644_8799.n30 a_n5644_8799.n13 37.246
R14734 a_n5644_8799.n42 a_n5644_8799.n41 37.246
R14735 a_n5644_8799.n52 a_n5644_8799.n35 37.246
R14736 a_n5644_8799.n65 a_n5644_8799.n64 37.246
R14737 a_n5644_8799.n75 a_n5644_8799.n58 37.246
R14738 a_n5644_8799.n94 a_n5644_8799.n81 35.7853
R14739 a_n5644_8799.n91 a_n5644_8799.n84 35.7853
R14740 a_n5644_8799.n116 a_n5644_8799.n103 35.7853
R14741 a_n5644_8799.n113 a_n5644_8799.n106 35.7853
R14742 a_n5644_8799.n139 a_n5644_8799.n126 35.7853
R14743 a_n5644_8799.n136 a_n5644_8799.n129 35.7853
R14744 a_n5644_8799.n20 a_n5644_8799.n15 35.7853
R14745 a_n5644_8799.n26 a_n5644_8799.n13 35.7853
R14746 a_n5644_8799.n42 a_n5644_8799.n37 35.7853
R14747 a_n5644_8799.n48 a_n5644_8799.n35 35.7853
R14748 a_n5644_8799.n65 a_n5644_8799.n60 35.7853
R14749 a_n5644_8799.n71 a_n5644_8799.n58 35.7853
R14750 a_n5644_8799.n163 a_n5644_8799.n158 32.7526
R14751 a_n5644_8799.n11 a_n5644_8799.n5 30.7135
R14752 a_n5644_8799.n86 a_n5644_8799.n85 20.9576
R14753 a_n5644_8799.n108 a_n5644_8799.n107 20.9576
R14754 a_n5644_8799.n131 a_n5644_8799.n130 20.9576
R14755 a_n5644_8799.n18 a_n5644_8799.n17 20.9576
R14756 a_n5644_8799.n40 a_n5644_8799.n39 20.9576
R14757 a_n5644_8799.n63 a_n5644_8799.n62 20.9576
R14758 a_n5644_8799.n11 a_n5644_8799.n10 17.7361
R14759 a_n5644_8799.n94 a_n5644_8799.n93 12.4157
R14760 a_n5644_8799.n92 a_n5644_8799.n91 12.4157
R14761 a_n5644_8799.n116 a_n5644_8799.n115 12.4157
R14762 a_n5644_8799.n114 a_n5644_8799.n113 12.4157
R14763 a_n5644_8799.n139 a_n5644_8799.n138 12.4157
R14764 a_n5644_8799.n137 a_n5644_8799.n136 12.4157
R14765 a_n5644_8799.n24 a_n5644_8799.n15 12.4157
R14766 a_n5644_8799.n26 a_n5644_8799.n25 12.4157
R14767 a_n5644_8799.n46 a_n5644_8799.n37 12.4157
R14768 a_n5644_8799.n48 a_n5644_8799.n47 12.4157
R14769 a_n5644_8799.n69 a_n5644_8799.n60 12.4157
R14770 a_n5644_8799.n71 a_n5644_8799.n70 12.4157
R14771 a_n5644_8799.n154 a_n5644_8799.n149 12.3339
R14772 a_n5644_8799.n149 a_n5644_8799.n11 11.4887
R14773 a_n5644_8799.n99 a_n5644_8799.n98 10.955
R14774 a_n5644_8799.n87 a_n5644_8799.n86 10.955
R14775 a_n5644_8799.n121 a_n5644_8799.n120 10.955
R14776 a_n5644_8799.n109 a_n5644_8799.n108 10.955
R14777 a_n5644_8799.n144 a_n5644_8799.n143 10.955
R14778 a_n5644_8799.n132 a_n5644_8799.n131 10.955
R14779 a_n5644_8799.n19 a_n5644_8799.n18 10.955
R14780 a_n5644_8799.n31 a_n5644_8799.n30 10.955
R14781 a_n5644_8799.n41 a_n5644_8799.n40 10.955
R14782 a_n5644_8799.n53 a_n5644_8799.n52 10.955
R14783 a_n5644_8799.n64 a_n5644_8799.n63 10.955
R14784 a_n5644_8799.n76 a_n5644_8799.n75 10.955
R14785 a_n5644_8799.n124 a_n5644_8799.n101 9.05164
R14786 a_n5644_8799.n56 a_n5644_8799.n33 9.05164
R14787 a_n5644_8799.n148 a_n5644_8799.n79 6.86985
R14788 a_n5644_8799.n148 a_n5644_8799.n147 6.51296
R14789 a_n5644_8799.n124 a_n5644_8799.n123 4.94368
R14790 a_n5644_8799.n147 a_n5644_8799.n146 4.94368
R14791 a_n5644_8799.n56 a_n5644_8799.n55 4.94368
R14792 a_n5644_8799.n79 a_n5644_8799.n78 4.94368
R14793 a_n5644_8799.n147 a_n5644_8799.n124 4.10845
R14794 a_n5644_8799.n79 a_n5644_8799.n56 4.10845
R14795 a_n5644_8799.n9 a_n5644_8799.t31 3.61217
R14796 a_n5644_8799.n9 a_n5644_8799.t22 3.61217
R14797 a_n5644_8799.n7 a_n5644_8799.t29 3.61217
R14798 a_n5644_8799.n7 a_n5644_8799.t24 3.61217
R14799 a_n5644_8799.n6 a_n5644_8799.t23 3.61217
R14800 a_n5644_8799.n6 a_n5644_8799.t25 3.61217
R14801 a_n5644_8799.n1 a_n5644_8799.t30 3.61217
R14802 a_n5644_8799.n1 a_n5644_8799.t20 3.61217
R14803 a_n5644_8799.n2 a_n5644_8799.t26 3.61217
R14804 a_n5644_8799.n2 a_n5644_8799.t27 3.61217
R14805 a_n5644_8799.n4 a_n5644_8799.t28 3.61217
R14806 a_n5644_8799.n4 a_n5644_8799.t21 3.61217
R14807 a_n5644_8799.n149 a_n5644_8799.n148 3.4105
R14808 a_n5644_8799.n159 a_n5644_8799.t13 2.82907
R14809 a_n5644_8799.n159 a_n5644_8799.t11 2.82907
R14810 a_n5644_8799.n160 a_n5644_8799.t4 2.82907
R14811 a_n5644_8799.n160 a_n5644_8799.t8 2.82907
R14812 a_n5644_8799.n162 a_n5644_8799.t18 2.82907
R14813 a_n5644_8799.n162 a_n5644_8799.t5 2.82907
R14814 a_n5644_8799.n157 a_n5644_8799.t14 2.82907
R14815 a_n5644_8799.n157 a_n5644_8799.t0 2.82907
R14816 a_n5644_8799.n155 a_n5644_8799.t17 2.82907
R14817 a_n5644_8799.n155 a_n5644_8799.t12 2.82907
R14818 a_n5644_8799.n153 a_n5644_8799.t1 2.82907
R14819 a_n5644_8799.n153 a_n5644_8799.t16 2.82907
R14820 a_n5644_8799.n151 a_n5644_8799.t2 2.82907
R14821 a_n5644_8799.n151 a_n5644_8799.t3 2.82907
R14822 a_n5644_8799.n150 a_n5644_8799.t6 2.82907
R14823 a_n5644_8799.n150 a_n5644_8799.t7 2.82907
R14824 a_n5644_8799.n0 a_n5644_8799.t10 2.82907
R14825 a_n5644_8799.n0 a_n5644_8799.t9 2.82907
R14826 a_n5644_8799.n165 a_n5644_8799.t15 2.82907
R14827 a_n5644_8799.t19 a_n5644_8799.n165 2.82907
R14828 a_n5644_8799.n154 a_n5644_8799.n152 0.444466
R14829 a_n5644_8799.n156 a_n5644_8799.n154 0.444466
R14830 a_n5644_8799.n158 a_n5644_8799.n156 0.444466
R14831 a_n5644_8799.n164 a_n5644_8799.n163 0.444466
R14832 a_n5644_8799.n163 a_n5644_8799.n161 0.444466
R14833 a_n5644_8799.n10 a_n5644_8799.n8 0.358259
R14834 a_n5644_8799.n5 a_n5644_8799.n3 0.358259
R14835 a_n5644_8799.n101 a_n5644_8799.n80 0.189894
R14836 a_n5644_8799.n97 a_n5644_8799.n80 0.189894
R14837 a_n5644_8799.n97 a_n5644_8799.n96 0.189894
R14838 a_n5644_8799.n96 a_n5644_8799.n95 0.189894
R14839 a_n5644_8799.n95 a_n5644_8799.n82 0.189894
R14840 a_n5644_8799.n83 a_n5644_8799.n82 0.189894
R14841 a_n5644_8799.n90 a_n5644_8799.n83 0.189894
R14842 a_n5644_8799.n90 a_n5644_8799.n89 0.189894
R14843 a_n5644_8799.n89 a_n5644_8799.n88 0.189894
R14844 a_n5644_8799.n123 a_n5644_8799.n102 0.189894
R14845 a_n5644_8799.n119 a_n5644_8799.n102 0.189894
R14846 a_n5644_8799.n119 a_n5644_8799.n118 0.189894
R14847 a_n5644_8799.n118 a_n5644_8799.n117 0.189894
R14848 a_n5644_8799.n117 a_n5644_8799.n104 0.189894
R14849 a_n5644_8799.n105 a_n5644_8799.n104 0.189894
R14850 a_n5644_8799.n112 a_n5644_8799.n105 0.189894
R14851 a_n5644_8799.n112 a_n5644_8799.n111 0.189894
R14852 a_n5644_8799.n111 a_n5644_8799.n110 0.189894
R14853 a_n5644_8799.n146 a_n5644_8799.n125 0.189894
R14854 a_n5644_8799.n142 a_n5644_8799.n125 0.189894
R14855 a_n5644_8799.n142 a_n5644_8799.n141 0.189894
R14856 a_n5644_8799.n141 a_n5644_8799.n140 0.189894
R14857 a_n5644_8799.n140 a_n5644_8799.n127 0.189894
R14858 a_n5644_8799.n128 a_n5644_8799.n127 0.189894
R14859 a_n5644_8799.n135 a_n5644_8799.n128 0.189894
R14860 a_n5644_8799.n135 a_n5644_8799.n134 0.189894
R14861 a_n5644_8799.n134 a_n5644_8799.n133 0.189894
R14862 a_n5644_8799.n21 a_n5644_8799.n16 0.189894
R14863 a_n5644_8799.n22 a_n5644_8799.n21 0.189894
R14864 a_n5644_8799.n23 a_n5644_8799.n22 0.189894
R14865 a_n5644_8799.n23 a_n5644_8799.n14 0.189894
R14866 a_n5644_8799.n27 a_n5644_8799.n14 0.189894
R14867 a_n5644_8799.n28 a_n5644_8799.n27 0.189894
R14868 a_n5644_8799.n29 a_n5644_8799.n28 0.189894
R14869 a_n5644_8799.n29 a_n5644_8799.n12 0.189894
R14870 a_n5644_8799.n33 a_n5644_8799.n12 0.189894
R14871 a_n5644_8799.n43 a_n5644_8799.n38 0.189894
R14872 a_n5644_8799.n44 a_n5644_8799.n43 0.189894
R14873 a_n5644_8799.n45 a_n5644_8799.n44 0.189894
R14874 a_n5644_8799.n45 a_n5644_8799.n36 0.189894
R14875 a_n5644_8799.n49 a_n5644_8799.n36 0.189894
R14876 a_n5644_8799.n50 a_n5644_8799.n49 0.189894
R14877 a_n5644_8799.n51 a_n5644_8799.n50 0.189894
R14878 a_n5644_8799.n51 a_n5644_8799.n34 0.189894
R14879 a_n5644_8799.n55 a_n5644_8799.n34 0.189894
R14880 a_n5644_8799.n66 a_n5644_8799.n61 0.189894
R14881 a_n5644_8799.n67 a_n5644_8799.n66 0.189894
R14882 a_n5644_8799.n68 a_n5644_8799.n67 0.189894
R14883 a_n5644_8799.n68 a_n5644_8799.n59 0.189894
R14884 a_n5644_8799.n72 a_n5644_8799.n59 0.189894
R14885 a_n5644_8799.n73 a_n5644_8799.n72 0.189894
R14886 a_n5644_8799.n74 a_n5644_8799.n73 0.189894
R14887 a_n5644_8799.n74 a_n5644_8799.n57 0.189894
R14888 a_n5644_8799.n78 a_n5644_8799.n57 0.189894
R14889 vdd.n291 vdd.n255 756.745
R14890 vdd.n244 vdd.n208 756.745
R14891 vdd.n201 vdd.n165 756.745
R14892 vdd.n154 vdd.n118 756.745
R14893 vdd.n112 vdd.n76 756.745
R14894 vdd.n65 vdd.n29 756.745
R14895 vdd.n1106 vdd.n1070 756.745
R14896 vdd.n1153 vdd.n1117 756.745
R14897 vdd.n1016 vdd.n980 756.745
R14898 vdd.n1063 vdd.n1027 756.745
R14899 vdd.n927 vdd.n891 756.745
R14900 vdd.n974 vdd.n938 756.745
R14901 vdd.n1791 vdd.t171 640.208
R14902 vdd.n755 vdd.t156 640.208
R14903 vdd.n1765 vdd.t197 640.208
R14904 vdd.n747 vdd.t188 640.208
R14905 vdd.n2536 vdd.t139 640.208
R14906 vdd.n2256 vdd.t179 640.208
R14907 vdd.n622 vdd.t160 640.208
R14908 vdd.n2253 vdd.t164 640.208
R14909 vdd.n589 vdd.t168 640.208
R14910 vdd.n817 vdd.t175 640.208
R14911 vdd.n1320 vdd.t135 592.009
R14912 vdd.n1358 vdd.t182 592.009
R14913 vdd.n1254 vdd.t185 592.009
R14914 vdd.n1947 vdd.t131 592.009
R14915 vdd.n1584 vdd.t143 592.009
R14916 vdd.n1544 vdd.t150 592.009
R14917 vdd.n2908 vdd.t194 592.009
R14918 vdd.n405 vdd.t146 592.009
R14919 vdd.n365 vdd.t153 592.009
R14920 vdd.n557 vdd.t124 592.009
R14921 vdd.n2804 vdd.t128 592.009
R14922 vdd.n2711 vdd.t191 592.009
R14923 vdd.n292 vdd.n291 585
R14924 vdd.n290 vdd.n257 585
R14925 vdd.n289 vdd.n288 585
R14926 vdd.n260 vdd.n258 585
R14927 vdd.n283 vdd.n282 585
R14928 vdd.n281 vdd.n280 585
R14929 vdd.n264 vdd.n263 585
R14930 vdd.n275 vdd.n274 585
R14931 vdd.n273 vdd.n272 585
R14932 vdd.n268 vdd.n267 585
R14933 vdd.n245 vdd.n244 585
R14934 vdd.n243 vdd.n210 585
R14935 vdd.n242 vdd.n241 585
R14936 vdd.n213 vdd.n211 585
R14937 vdd.n236 vdd.n235 585
R14938 vdd.n234 vdd.n233 585
R14939 vdd.n217 vdd.n216 585
R14940 vdd.n228 vdd.n227 585
R14941 vdd.n226 vdd.n225 585
R14942 vdd.n221 vdd.n220 585
R14943 vdd.n202 vdd.n201 585
R14944 vdd.n200 vdd.n167 585
R14945 vdd.n199 vdd.n198 585
R14946 vdd.n170 vdd.n168 585
R14947 vdd.n193 vdd.n192 585
R14948 vdd.n191 vdd.n190 585
R14949 vdd.n174 vdd.n173 585
R14950 vdd.n185 vdd.n184 585
R14951 vdd.n183 vdd.n182 585
R14952 vdd.n178 vdd.n177 585
R14953 vdd.n155 vdd.n154 585
R14954 vdd.n153 vdd.n120 585
R14955 vdd.n152 vdd.n151 585
R14956 vdd.n123 vdd.n121 585
R14957 vdd.n146 vdd.n145 585
R14958 vdd.n144 vdd.n143 585
R14959 vdd.n127 vdd.n126 585
R14960 vdd.n138 vdd.n137 585
R14961 vdd.n136 vdd.n135 585
R14962 vdd.n131 vdd.n130 585
R14963 vdd.n113 vdd.n112 585
R14964 vdd.n111 vdd.n78 585
R14965 vdd.n110 vdd.n109 585
R14966 vdd.n81 vdd.n79 585
R14967 vdd.n104 vdd.n103 585
R14968 vdd.n102 vdd.n101 585
R14969 vdd.n85 vdd.n84 585
R14970 vdd.n96 vdd.n95 585
R14971 vdd.n94 vdd.n93 585
R14972 vdd.n89 vdd.n88 585
R14973 vdd.n66 vdd.n65 585
R14974 vdd.n64 vdd.n31 585
R14975 vdd.n63 vdd.n62 585
R14976 vdd.n34 vdd.n32 585
R14977 vdd.n57 vdd.n56 585
R14978 vdd.n55 vdd.n54 585
R14979 vdd.n38 vdd.n37 585
R14980 vdd.n49 vdd.n48 585
R14981 vdd.n47 vdd.n46 585
R14982 vdd.n42 vdd.n41 585
R14983 vdd.n1107 vdd.n1106 585
R14984 vdd.n1105 vdd.n1072 585
R14985 vdd.n1104 vdd.n1103 585
R14986 vdd.n1075 vdd.n1073 585
R14987 vdd.n1098 vdd.n1097 585
R14988 vdd.n1096 vdd.n1095 585
R14989 vdd.n1079 vdd.n1078 585
R14990 vdd.n1090 vdd.n1089 585
R14991 vdd.n1088 vdd.n1087 585
R14992 vdd.n1083 vdd.n1082 585
R14993 vdd.n1154 vdd.n1153 585
R14994 vdd.n1152 vdd.n1119 585
R14995 vdd.n1151 vdd.n1150 585
R14996 vdd.n1122 vdd.n1120 585
R14997 vdd.n1145 vdd.n1144 585
R14998 vdd.n1143 vdd.n1142 585
R14999 vdd.n1126 vdd.n1125 585
R15000 vdd.n1137 vdd.n1136 585
R15001 vdd.n1135 vdd.n1134 585
R15002 vdd.n1130 vdd.n1129 585
R15003 vdd.n1017 vdd.n1016 585
R15004 vdd.n1015 vdd.n982 585
R15005 vdd.n1014 vdd.n1013 585
R15006 vdd.n985 vdd.n983 585
R15007 vdd.n1008 vdd.n1007 585
R15008 vdd.n1006 vdd.n1005 585
R15009 vdd.n989 vdd.n988 585
R15010 vdd.n1000 vdd.n999 585
R15011 vdd.n998 vdd.n997 585
R15012 vdd.n993 vdd.n992 585
R15013 vdd.n1064 vdd.n1063 585
R15014 vdd.n1062 vdd.n1029 585
R15015 vdd.n1061 vdd.n1060 585
R15016 vdd.n1032 vdd.n1030 585
R15017 vdd.n1055 vdd.n1054 585
R15018 vdd.n1053 vdd.n1052 585
R15019 vdd.n1036 vdd.n1035 585
R15020 vdd.n1047 vdd.n1046 585
R15021 vdd.n1045 vdd.n1044 585
R15022 vdd.n1040 vdd.n1039 585
R15023 vdd.n928 vdd.n927 585
R15024 vdd.n926 vdd.n893 585
R15025 vdd.n925 vdd.n924 585
R15026 vdd.n896 vdd.n894 585
R15027 vdd.n919 vdd.n918 585
R15028 vdd.n917 vdd.n916 585
R15029 vdd.n900 vdd.n899 585
R15030 vdd.n911 vdd.n910 585
R15031 vdd.n909 vdd.n908 585
R15032 vdd.n904 vdd.n903 585
R15033 vdd.n975 vdd.n974 585
R15034 vdd.n973 vdd.n940 585
R15035 vdd.n972 vdd.n971 585
R15036 vdd.n943 vdd.n941 585
R15037 vdd.n966 vdd.n965 585
R15038 vdd.n964 vdd.n963 585
R15039 vdd.n947 vdd.n946 585
R15040 vdd.n958 vdd.n957 585
R15041 vdd.n956 vdd.n955 585
R15042 vdd.n951 vdd.n950 585
R15043 vdd.n3024 vdd.n330 515.122
R15044 vdd.n2906 vdd.n328 515.122
R15045 vdd.n515 vdd.n478 515.122
R15046 vdd.n2842 vdd.n479 515.122
R15047 vdd.n1942 vdd.n865 515.122
R15048 vdd.n1945 vdd.n1944 515.122
R15049 vdd.n1227 vdd.n1191 515.122
R15050 vdd.n1423 vdd.n1192 515.122
R15051 vdd.n269 vdd.t47 329.043
R15052 vdd.n222 vdd.t58 329.043
R15053 vdd.n179 vdd.t43 329.043
R15054 vdd.n132 vdd.t53 329.043
R15055 vdd.n90 vdd.t84 329.043
R15056 vdd.n43 vdd.t26 329.043
R15057 vdd.n1084 vdd.t82 329.043
R15058 vdd.n1131 vdd.t68 329.043
R15059 vdd.n994 vdd.t74 329.043
R15060 vdd.n1041 vdd.t61 329.043
R15061 vdd.n905 vdd.t24 329.043
R15062 vdd.n952 vdd.t83 329.043
R15063 vdd.n1320 vdd.t138 319.788
R15064 vdd.n1358 vdd.t184 319.788
R15065 vdd.n1254 vdd.t187 319.788
R15066 vdd.n1947 vdd.t133 319.788
R15067 vdd.n1584 vdd.t144 319.788
R15068 vdd.n1544 vdd.t151 319.788
R15069 vdd.n2908 vdd.t195 319.788
R15070 vdd.n405 vdd.t148 319.788
R15071 vdd.n365 vdd.t154 319.788
R15072 vdd.n557 vdd.t127 319.788
R15073 vdd.n2804 vdd.t130 319.788
R15074 vdd.n2711 vdd.t193 319.788
R15075 vdd.n1321 vdd.t137 303.69
R15076 vdd.n1359 vdd.t183 303.69
R15077 vdd.n1255 vdd.t186 303.69
R15078 vdd.n1948 vdd.t134 303.69
R15079 vdd.n1585 vdd.t145 303.69
R15080 vdd.n1545 vdd.t152 303.69
R15081 vdd.n2909 vdd.t196 303.69
R15082 vdd.n406 vdd.t149 303.69
R15083 vdd.n366 vdd.t155 303.69
R15084 vdd.n558 vdd.t126 303.69
R15085 vdd.n2805 vdd.t129 303.69
R15086 vdd.n2712 vdd.t192 303.69
R15087 vdd.n2479 vdd.n703 297.074
R15088 vdd.n2672 vdd.n599 297.074
R15089 vdd.n2609 vdd.n596 297.074
R15090 vdd.n2402 vdd.n704 297.074
R15091 vdd.n2217 vdd.n744 297.074
R15092 vdd.n2148 vdd.n2147 297.074
R15093 vdd.n1894 vdd.n840 297.074
R15094 vdd.n1990 vdd.n838 297.074
R15095 vdd.n2588 vdd.n597 297.074
R15096 vdd.n2675 vdd.n2674 297.074
R15097 vdd.n2251 vdd.n705 297.074
R15098 vdd.n2477 vdd.n706 297.074
R15099 vdd.n2145 vdd.n753 297.074
R15100 vdd.n751 vdd.n726 297.074
R15101 vdd.n1831 vdd.n841 297.074
R15102 vdd.n1988 vdd.n842 297.074
R15103 vdd.n2590 vdd.n597 185
R15104 vdd.n2673 vdd.n597 185
R15105 vdd.n2592 vdd.n2591 185
R15106 vdd.n2591 vdd.n595 185
R15107 vdd.n2593 vdd.n629 185
R15108 vdd.n2603 vdd.n629 185
R15109 vdd.n2594 vdd.n638 185
R15110 vdd.n638 vdd.n636 185
R15111 vdd.n2596 vdd.n2595 185
R15112 vdd.n2597 vdd.n2596 185
R15113 vdd.n2549 vdd.n637 185
R15114 vdd.n637 vdd.n633 185
R15115 vdd.n2548 vdd.n2547 185
R15116 vdd.n2547 vdd.n2546 185
R15117 vdd.n640 vdd.n639 185
R15118 vdd.n641 vdd.n640 185
R15119 vdd.n2539 vdd.n2538 185
R15120 vdd.n2540 vdd.n2539 185
R15121 vdd.n2535 vdd.n650 185
R15122 vdd.n650 vdd.n647 185
R15123 vdd.n2534 vdd.n2533 185
R15124 vdd.n2533 vdd.n2532 185
R15125 vdd.n652 vdd.n651 185
R15126 vdd.n660 vdd.n652 185
R15127 vdd.n2525 vdd.n2524 185
R15128 vdd.n2526 vdd.n2525 185
R15129 vdd.n2523 vdd.n661 185
R15130 vdd.n2374 vdd.n661 185
R15131 vdd.n2522 vdd.n2521 185
R15132 vdd.n2521 vdd.n2520 185
R15133 vdd.n663 vdd.n662 185
R15134 vdd.n664 vdd.n663 185
R15135 vdd.n2513 vdd.n2512 185
R15136 vdd.n2514 vdd.n2513 185
R15137 vdd.n2511 vdd.n673 185
R15138 vdd.n673 vdd.n670 185
R15139 vdd.n2510 vdd.n2509 185
R15140 vdd.n2509 vdd.n2508 185
R15141 vdd.n675 vdd.n674 185
R15142 vdd.n683 vdd.n675 185
R15143 vdd.n2501 vdd.n2500 185
R15144 vdd.n2502 vdd.n2501 185
R15145 vdd.n2499 vdd.n684 185
R15146 vdd.n690 vdd.n684 185
R15147 vdd.n2498 vdd.n2497 185
R15148 vdd.n2497 vdd.n2496 185
R15149 vdd.n686 vdd.n685 185
R15150 vdd.n687 vdd.n686 185
R15151 vdd.n2489 vdd.n2488 185
R15152 vdd.n2490 vdd.n2489 185
R15153 vdd.n2487 vdd.n696 185
R15154 vdd.n2395 vdd.n696 185
R15155 vdd.n2486 vdd.n2485 185
R15156 vdd.n2485 vdd.n2484 185
R15157 vdd.n698 vdd.n697 185
R15158 vdd.t21 vdd.n698 185
R15159 vdd.n2477 vdd.n2476 185
R15160 vdd.n2478 vdd.n2477 185
R15161 vdd.n2475 vdd.n706 185
R15162 vdd.n2474 vdd.n2473 185
R15163 vdd.n708 vdd.n707 185
R15164 vdd.n2260 vdd.n2259 185
R15165 vdd.n2262 vdd.n2261 185
R15166 vdd.n2264 vdd.n2263 185
R15167 vdd.n2266 vdd.n2265 185
R15168 vdd.n2268 vdd.n2267 185
R15169 vdd.n2270 vdd.n2269 185
R15170 vdd.n2272 vdd.n2271 185
R15171 vdd.n2274 vdd.n2273 185
R15172 vdd.n2276 vdd.n2275 185
R15173 vdd.n2278 vdd.n2277 185
R15174 vdd.n2280 vdd.n2279 185
R15175 vdd.n2282 vdd.n2281 185
R15176 vdd.n2284 vdd.n2283 185
R15177 vdd.n2286 vdd.n2285 185
R15178 vdd.n2288 vdd.n2287 185
R15179 vdd.n2290 vdd.n2289 185
R15180 vdd.n2292 vdd.n2291 185
R15181 vdd.n2294 vdd.n2293 185
R15182 vdd.n2296 vdd.n2295 185
R15183 vdd.n2298 vdd.n2297 185
R15184 vdd.n2300 vdd.n2299 185
R15185 vdd.n2302 vdd.n2301 185
R15186 vdd.n2304 vdd.n2303 185
R15187 vdd.n2306 vdd.n2305 185
R15188 vdd.n2308 vdd.n2307 185
R15189 vdd.n2310 vdd.n2309 185
R15190 vdd.n2312 vdd.n2311 185
R15191 vdd.n2314 vdd.n2313 185
R15192 vdd.n2316 vdd.n2315 185
R15193 vdd.n2318 vdd.n2317 185
R15194 vdd.n2320 vdd.n2319 185
R15195 vdd.n2321 vdd.n2251 185
R15196 vdd.n2471 vdd.n2251 185
R15197 vdd.n2676 vdd.n2675 185
R15198 vdd.n2677 vdd.n588 185
R15199 vdd.n2679 vdd.n2678 185
R15200 vdd.n2681 vdd.n586 185
R15201 vdd.n2683 vdd.n2682 185
R15202 vdd.n2684 vdd.n585 185
R15203 vdd.n2686 vdd.n2685 185
R15204 vdd.n2688 vdd.n583 185
R15205 vdd.n2690 vdd.n2689 185
R15206 vdd.n2691 vdd.n582 185
R15207 vdd.n2693 vdd.n2692 185
R15208 vdd.n2695 vdd.n580 185
R15209 vdd.n2697 vdd.n2696 185
R15210 vdd.n2698 vdd.n579 185
R15211 vdd.n2700 vdd.n2699 185
R15212 vdd.n2702 vdd.n578 185
R15213 vdd.n2703 vdd.n576 185
R15214 vdd.n2706 vdd.n2705 185
R15215 vdd.n577 vdd.n575 185
R15216 vdd.n2562 vdd.n2561 185
R15217 vdd.n2564 vdd.n2563 185
R15218 vdd.n2566 vdd.n2558 185
R15219 vdd.n2568 vdd.n2567 185
R15220 vdd.n2569 vdd.n2557 185
R15221 vdd.n2571 vdd.n2570 185
R15222 vdd.n2573 vdd.n2555 185
R15223 vdd.n2575 vdd.n2574 185
R15224 vdd.n2576 vdd.n2554 185
R15225 vdd.n2578 vdd.n2577 185
R15226 vdd.n2580 vdd.n2552 185
R15227 vdd.n2582 vdd.n2581 185
R15228 vdd.n2583 vdd.n2551 185
R15229 vdd.n2585 vdd.n2584 185
R15230 vdd.n2587 vdd.n2550 185
R15231 vdd.n2589 vdd.n2588 185
R15232 vdd.n2588 vdd.n484 185
R15233 vdd.n2674 vdd.n592 185
R15234 vdd.n2674 vdd.n2673 185
R15235 vdd.n2326 vdd.n594 185
R15236 vdd.n595 vdd.n594 185
R15237 vdd.n2327 vdd.n628 185
R15238 vdd.n2603 vdd.n628 185
R15239 vdd.n2329 vdd.n2328 185
R15240 vdd.n2328 vdd.n636 185
R15241 vdd.n2330 vdd.n635 185
R15242 vdd.n2597 vdd.n635 185
R15243 vdd.n2332 vdd.n2331 185
R15244 vdd.n2331 vdd.n633 185
R15245 vdd.n2333 vdd.n643 185
R15246 vdd.n2546 vdd.n643 185
R15247 vdd.n2335 vdd.n2334 185
R15248 vdd.n2334 vdd.n641 185
R15249 vdd.n2336 vdd.n649 185
R15250 vdd.n2540 vdd.n649 185
R15251 vdd.n2338 vdd.n2337 185
R15252 vdd.n2337 vdd.n647 185
R15253 vdd.n2339 vdd.n654 185
R15254 vdd.n2532 vdd.n654 185
R15255 vdd.n2341 vdd.n2340 185
R15256 vdd.n2340 vdd.n660 185
R15257 vdd.n2342 vdd.n659 185
R15258 vdd.n2526 vdd.n659 185
R15259 vdd.n2376 vdd.n2375 185
R15260 vdd.n2375 vdd.n2374 185
R15261 vdd.n2377 vdd.n666 185
R15262 vdd.n2520 vdd.n666 185
R15263 vdd.n2379 vdd.n2378 185
R15264 vdd.n2378 vdd.n664 185
R15265 vdd.n2380 vdd.n672 185
R15266 vdd.n2514 vdd.n672 185
R15267 vdd.n2382 vdd.n2381 185
R15268 vdd.n2381 vdd.n670 185
R15269 vdd.n2383 vdd.n677 185
R15270 vdd.n2508 vdd.n677 185
R15271 vdd.n2385 vdd.n2384 185
R15272 vdd.n2384 vdd.n683 185
R15273 vdd.n2386 vdd.n682 185
R15274 vdd.n2502 vdd.n682 185
R15275 vdd.n2388 vdd.n2387 185
R15276 vdd.n2387 vdd.n690 185
R15277 vdd.n2389 vdd.n689 185
R15278 vdd.n2496 vdd.n689 185
R15279 vdd.n2391 vdd.n2390 185
R15280 vdd.n2390 vdd.n687 185
R15281 vdd.n2392 vdd.n695 185
R15282 vdd.n2490 vdd.n695 185
R15283 vdd.n2394 vdd.n2393 185
R15284 vdd.n2395 vdd.n2394 185
R15285 vdd.n2325 vdd.n700 185
R15286 vdd.n2484 vdd.n700 185
R15287 vdd.n2324 vdd.n2323 185
R15288 vdd.n2323 vdd.t21 185
R15289 vdd.n2322 vdd.n705 185
R15290 vdd.n2478 vdd.n705 185
R15291 vdd.n1942 vdd.n1941 185
R15292 vdd.n1943 vdd.n1942 185
R15293 vdd.n866 vdd.n864 185
R15294 vdd.n1508 vdd.n864 185
R15295 vdd.n1511 vdd.n1510 185
R15296 vdd.n1510 vdd.n1509 185
R15297 vdd.n869 vdd.n868 185
R15298 vdd.n870 vdd.n869 185
R15299 vdd.n1497 vdd.n1496 185
R15300 vdd.n1498 vdd.n1497 185
R15301 vdd.n878 vdd.n877 185
R15302 vdd.n1489 vdd.n877 185
R15303 vdd.n1492 vdd.n1491 185
R15304 vdd.n1491 vdd.n1490 185
R15305 vdd.n881 vdd.n880 185
R15306 vdd.n888 vdd.n881 185
R15307 vdd.n1480 vdd.n1479 185
R15308 vdd.n1481 vdd.n1480 185
R15309 vdd.n890 vdd.n889 185
R15310 vdd.n889 vdd.n887 185
R15311 vdd.n1475 vdd.n1474 185
R15312 vdd.n1474 vdd.n1473 185
R15313 vdd.n1163 vdd.n1162 185
R15314 vdd.n1164 vdd.n1163 185
R15315 vdd.n1464 vdd.n1463 185
R15316 vdd.n1465 vdd.n1464 185
R15317 vdd.n1171 vdd.n1170 185
R15318 vdd.n1455 vdd.n1170 185
R15319 vdd.n1458 vdd.n1457 185
R15320 vdd.n1457 vdd.n1456 185
R15321 vdd.n1174 vdd.n1173 185
R15322 vdd.n1180 vdd.n1174 185
R15323 vdd.n1446 vdd.n1445 185
R15324 vdd.n1447 vdd.n1446 185
R15325 vdd.n1182 vdd.n1181 185
R15326 vdd.n1438 vdd.n1181 185
R15327 vdd.n1441 vdd.n1440 185
R15328 vdd.n1440 vdd.n1439 185
R15329 vdd.n1185 vdd.n1184 185
R15330 vdd.n1186 vdd.n1185 185
R15331 vdd.n1429 vdd.n1428 185
R15332 vdd.n1430 vdd.n1429 185
R15333 vdd.n1193 vdd.n1192 185
R15334 vdd.n1228 vdd.n1192 185
R15335 vdd.n1424 vdd.n1423 185
R15336 vdd.n1196 vdd.n1195 185
R15337 vdd.n1420 vdd.n1419 185
R15338 vdd.n1421 vdd.n1420 185
R15339 vdd.n1230 vdd.n1229 185
R15340 vdd.n1415 vdd.n1232 185
R15341 vdd.n1414 vdd.n1233 185
R15342 vdd.n1413 vdd.n1234 185
R15343 vdd.n1236 vdd.n1235 185
R15344 vdd.n1409 vdd.n1238 185
R15345 vdd.n1408 vdd.n1239 185
R15346 vdd.n1407 vdd.n1240 185
R15347 vdd.n1242 vdd.n1241 185
R15348 vdd.n1403 vdd.n1244 185
R15349 vdd.n1402 vdd.n1245 185
R15350 vdd.n1401 vdd.n1246 185
R15351 vdd.n1248 vdd.n1247 185
R15352 vdd.n1397 vdd.n1250 185
R15353 vdd.n1396 vdd.n1251 185
R15354 vdd.n1395 vdd.n1252 185
R15355 vdd.n1256 vdd.n1253 185
R15356 vdd.n1391 vdd.n1258 185
R15357 vdd.n1390 vdd.n1259 185
R15358 vdd.n1389 vdd.n1260 185
R15359 vdd.n1262 vdd.n1261 185
R15360 vdd.n1385 vdd.n1264 185
R15361 vdd.n1384 vdd.n1265 185
R15362 vdd.n1383 vdd.n1266 185
R15363 vdd.n1268 vdd.n1267 185
R15364 vdd.n1379 vdd.n1270 185
R15365 vdd.n1378 vdd.n1271 185
R15366 vdd.n1377 vdd.n1272 185
R15367 vdd.n1274 vdd.n1273 185
R15368 vdd.n1373 vdd.n1276 185
R15369 vdd.n1372 vdd.n1277 185
R15370 vdd.n1371 vdd.n1278 185
R15371 vdd.n1280 vdd.n1279 185
R15372 vdd.n1367 vdd.n1282 185
R15373 vdd.n1366 vdd.n1283 185
R15374 vdd.n1365 vdd.n1284 185
R15375 vdd.n1286 vdd.n1285 185
R15376 vdd.n1361 vdd.n1288 185
R15377 vdd.n1360 vdd.n1357 185
R15378 vdd.n1356 vdd.n1289 185
R15379 vdd.n1291 vdd.n1290 185
R15380 vdd.n1352 vdd.n1293 185
R15381 vdd.n1351 vdd.n1294 185
R15382 vdd.n1350 vdd.n1295 185
R15383 vdd.n1297 vdd.n1296 185
R15384 vdd.n1346 vdd.n1299 185
R15385 vdd.n1345 vdd.n1300 185
R15386 vdd.n1344 vdd.n1301 185
R15387 vdd.n1303 vdd.n1302 185
R15388 vdd.n1340 vdd.n1305 185
R15389 vdd.n1339 vdd.n1306 185
R15390 vdd.n1338 vdd.n1307 185
R15391 vdd.n1309 vdd.n1308 185
R15392 vdd.n1334 vdd.n1311 185
R15393 vdd.n1333 vdd.n1312 185
R15394 vdd.n1332 vdd.n1313 185
R15395 vdd.n1315 vdd.n1314 185
R15396 vdd.n1328 vdd.n1317 185
R15397 vdd.n1327 vdd.n1318 185
R15398 vdd.n1326 vdd.n1319 185
R15399 vdd.n1323 vdd.n1227 185
R15400 vdd.n1421 vdd.n1227 185
R15401 vdd.n1946 vdd.n1945 185
R15402 vdd.n1950 vdd.n859 185
R15403 vdd.n1613 vdd.n858 185
R15404 vdd.n1616 vdd.n1615 185
R15405 vdd.n1618 vdd.n1617 185
R15406 vdd.n1621 vdd.n1620 185
R15407 vdd.n1623 vdd.n1622 185
R15408 vdd.n1625 vdd.n1611 185
R15409 vdd.n1627 vdd.n1626 185
R15410 vdd.n1628 vdd.n1605 185
R15411 vdd.n1630 vdd.n1629 185
R15412 vdd.n1632 vdd.n1603 185
R15413 vdd.n1634 vdd.n1633 185
R15414 vdd.n1635 vdd.n1598 185
R15415 vdd.n1637 vdd.n1636 185
R15416 vdd.n1639 vdd.n1596 185
R15417 vdd.n1641 vdd.n1640 185
R15418 vdd.n1642 vdd.n1592 185
R15419 vdd.n1644 vdd.n1643 185
R15420 vdd.n1646 vdd.n1589 185
R15421 vdd.n1648 vdd.n1647 185
R15422 vdd.n1590 vdd.n1583 185
R15423 vdd.n1652 vdd.n1587 185
R15424 vdd.n1653 vdd.n1579 185
R15425 vdd.n1655 vdd.n1654 185
R15426 vdd.n1657 vdd.n1577 185
R15427 vdd.n1659 vdd.n1658 185
R15428 vdd.n1660 vdd.n1572 185
R15429 vdd.n1662 vdd.n1661 185
R15430 vdd.n1664 vdd.n1570 185
R15431 vdd.n1666 vdd.n1665 185
R15432 vdd.n1667 vdd.n1565 185
R15433 vdd.n1669 vdd.n1668 185
R15434 vdd.n1671 vdd.n1563 185
R15435 vdd.n1673 vdd.n1672 185
R15436 vdd.n1674 vdd.n1558 185
R15437 vdd.n1676 vdd.n1675 185
R15438 vdd.n1678 vdd.n1556 185
R15439 vdd.n1680 vdd.n1679 185
R15440 vdd.n1681 vdd.n1552 185
R15441 vdd.n1683 vdd.n1682 185
R15442 vdd.n1685 vdd.n1549 185
R15443 vdd.n1687 vdd.n1686 185
R15444 vdd.n1550 vdd.n1543 185
R15445 vdd.n1691 vdd.n1547 185
R15446 vdd.n1692 vdd.n1539 185
R15447 vdd.n1694 vdd.n1693 185
R15448 vdd.n1696 vdd.n1537 185
R15449 vdd.n1698 vdd.n1697 185
R15450 vdd.n1699 vdd.n1532 185
R15451 vdd.n1701 vdd.n1700 185
R15452 vdd.n1703 vdd.n1530 185
R15453 vdd.n1705 vdd.n1704 185
R15454 vdd.n1706 vdd.n1525 185
R15455 vdd.n1708 vdd.n1707 185
R15456 vdd.n1710 vdd.n1524 185
R15457 vdd.n1711 vdd.n1521 185
R15458 vdd.n1714 vdd.n1713 185
R15459 vdd.n1523 vdd.n1519 185
R15460 vdd.n1931 vdd.n1517 185
R15461 vdd.n1933 vdd.n1932 185
R15462 vdd.n1935 vdd.n1515 185
R15463 vdd.n1937 vdd.n1936 185
R15464 vdd.n1938 vdd.n865 185
R15465 vdd.n1944 vdd.n862 185
R15466 vdd.n1944 vdd.n1943 185
R15467 vdd.n873 vdd.n861 185
R15468 vdd.n1508 vdd.n861 185
R15469 vdd.n1507 vdd.n1506 185
R15470 vdd.n1509 vdd.n1507 185
R15471 vdd.n872 vdd.n871 185
R15472 vdd.n871 vdd.n870 185
R15473 vdd.n1500 vdd.n1499 185
R15474 vdd.n1499 vdd.n1498 185
R15475 vdd.n876 vdd.n875 185
R15476 vdd.n1489 vdd.n876 185
R15477 vdd.n1488 vdd.n1487 185
R15478 vdd.n1490 vdd.n1488 185
R15479 vdd.n883 vdd.n882 185
R15480 vdd.n888 vdd.n882 185
R15481 vdd.n1483 vdd.n1482 185
R15482 vdd.n1482 vdd.n1481 185
R15483 vdd.n886 vdd.n885 185
R15484 vdd.n887 vdd.n886 185
R15485 vdd.n1472 vdd.n1471 185
R15486 vdd.n1473 vdd.n1472 185
R15487 vdd.n1166 vdd.n1165 185
R15488 vdd.n1165 vdd.n1164 185
R15489 vdd.n1467 vdd.n1466 185
R15490 vdd.n1466 vdd.n1465 185
R15491 vdd.n1169 vdd.n1168 185
R15492 vdd.n1455 vdd.n1169 185
R15493 vdd.n1454 vdd.n1453 185
R15494 vdd.n1456 vdd.n1454 185
R15495 vdd.n1176 vdd.n1175 185
R15496 vdd.n1180 vdd.n1175 185
R15497 vdd.n1449 vdd.n1448 185
R15498 vdd.n1448 vdd.n1447 185
R15499 vdd.n1179 vdd.n1178 185
R15500 vdd.n1438 vdd.n1179 185
R15501 vdd.n1437 vdd.n1436 185
R15502 vdd.n1439 vdd.n1437 185
R15503 vdd.n1188 vdd.n1187 185
R15504 vdd.n1187 vdd.n1186 185
R15505 vdd.n1432 vdd.n1431 185
R15506 vdd.n1431 vdd.n1430 185
R15507 vdd.n1191 vdd.n1190 185
R15508 vdd.n1228 vdd.n1191 185
R15509 vdd.n746 vdd.n744 185
R15510 vdd.n2146 vdd.n744 185
R15511 vdd.n2068 vdd.n763 185
R15512 vdd.n763 vdd.t2 185
R15513 vdd.n2070 vdd.n2069 185
R15514 vdd.n2071 vdd.n2070 185
R15515 vdd.n2067 vdd.n762 185
R15516 vdd.n1770 vdd.n762 185
R15517 vdd.n2066 vdd.n2065 185
R15518 vdd.n2065 vdd.n2064 185
R15519 vdd.n765 vdd.n764 185
R15520 vdd.n766 vdd.n765 185
R15521 vdd.n2055 vdd.n2054 185
R15522 vdd.n2056 vdd.n2055 185
R15523 vdd.n2053 vdd.n776 185
R15524 vdd.n776 vdd.n773 185
R15525 vdd.n2052 vdd.n2051 185
R15526 vdd.n2051 vdd.n2050 185
R15527 vdd.n778 vdd.n777 185
R15528 vdd.n779 vdd.n778 185
R15529 vdd.n2043 vdd.n2042 185
R15530 vdd.n2044 vdd.n2043 185
R15531 vdd.n2041 vdd.n787 185
R15532 vdd.n792 vdd.n787 185
R15533 vdd.n2040 vdd.n2039 185
R15534 vdd.n2039 vdd.n2038 185
R15535 vdd.n789 vdd.n788 185
R15536 vdd.n798 vdd.n789 185
R15537 vdd.n2031 vdd.n2030 185
R15538 vdd.n2032 vdd.n2031 185
R15539 vdd.n2029 vdd.n799 185
R15540 vdd.n1871 vdd.n799 185
R15541 vdd.n2028 vdd.n2027 185
R15542 vdd.n2027 vdd.n2026 185
R15543 vdd.n801 vdd.n800 185
R15544 vdd.n802 vdd.n801 185
R15545 vdd.n2019 vdd.n2018 185
R15546 vdd.n2020 vdd.n2019 185
R15547 vdd.n2017 vdd.n811 185
R15548 vdd.n811 vdd.n808 185
R15549 vdd.n2016 vdd.n2015 185
R15550 vdd.n2015 vdd.n2014 185
R15551 vdd.n813 vdd.n812 185
R15552 vdd.n823 vdd.n813 185
R15553 vdd.n2006 vdd.n2005 185
R15554 vdd.n2007 vdd.n2006 185
R15555 vdd.n2004 vdd.n824 185
R15556 vdd.n824 vdd.n820 185
R15557 vdd.n2003 vdd.n2002 185
R15558 vdd.n2002 vdd.n2001 185
R15559 vdd.n826 vdd.n825 185
R15560 vdd.n827 vdd.n826 185
R15561 vdd.n1994 vdd.n1993 185
R15562 vdd.n1995 vdd.n1994 185
R15563 vdd.n1992 vdd.n836 185
R15564 vdd.n836 vdd.n833 185
R15565 vdd.n1991 vdd.n1990 185
R15566 vdd.n1990 vdd.n1989 185
R15567 vdd.n838 vdd.n837 185
R15568 vdd.n1726 vdd.n1725 185
R15569 vdd.n1727 vdd.n1723 185
R15570 vdd.n1723 vdd.n839 185
R15571 vdd.n1729 vdd.n1728 185
R15572 vdd.n1731 vdd.n1722 185
R15573 vdd.n1734 vdd.n1733 185
R15574 vdd.n1735 vdd.n1721 185
R15575 vdd.n1737 vdd.n1736 185
R15576 vdd.n1739 vdd.n1720 185
R15577 vdd.n1742 vdd.n1741 185
R15578 vdd.n1743 vdd.n1719 185
R15579 vdd.n1745 vdd.n1744 185
R15580 vdd.n1747 vdd.n1718 185
R15581 vdd.n1750 vdd.n1749 185
R15582 vdd.n1751 vdd.n1717 185
R15583 vdd.n1753 vdd.n1752 185
R15584 vdd.n1755 vdd.n1716 185
R15585 vdd.n1928 vdd.n1756 185
R15586 vdd.n1927 vdd.n1926 185
R15587 vdd.n1924 vdd.n1757 185
R15588 vdd.n1922 vdd.n1921 185
R15589 vdd.n1920 vdd.n1758 185
R15590 vdd.n1919 vdd.n1918 185
R15591 vdd.n1916 vdd.n1759 185
R15592 vdd.n1914 vdd.n1913 185
R15593 vdd.n1912 vdd.n1760 185
R15594 vdd.n1911 vdd.n1910 185
R15595 vdd.n1908 vdd.n1761 185
R15596 vdd.n1906 vdd.n1905 185
R15597 vdd.n1904 vdd.n1762 185
R15598 vdd.n1903 vdd.n1902 185
R15599 vdd.n1900 vdd.n1763 185
R15600 vdd.n1898 vdd.n1897 185
R15601 vdd.n1896 vdd.n1764 185
R15602 vdd.n1895 vdd.n1894 185
R15603 vdd.n2149 vdd.n2148 185
R15604 vdd.n2151 vdd.n2150 185
R15605 vdd.n2153 vdd.n2152 185
R15606 vdd.n2156 vdd.n2155 185
R15607 vdd.n2158 vdd.n2157 185
R15608 vdd.n2160 vdd.n2159 185
R15609 vdd.n2162 vdd.n2161 185
R15610 vdd.n2164 vdd.n2163 185
R15611 vdd.n2166 vdd.n2165 185
R15612 vdd.n2168 vdd.n2167 185
R15613 vdd.n2170 vdd.n2169 185
R15614 vdd.n2172 vdd.n2171 185
R15615 vdd.n2174 vdd.n2173 185
R15616 vdd.n2176 vdd.n2175 185
R15617 vdd.n2178 vdd.n2177 185
R15618 vdd.n2180 vdd.n2179 185
R15619 vdd.n2182 vdd.n2181 185
R15620 vdd.n2184 vdd.n2183 185
R15621 vdd.n2186 vdd.n2185 185
R15622 vdd.n2188 vdd.n2187 185
R15623 vdd.n2190 vdd.n2189 185
R15624 vdd.n2192 vdd.n2191 185
R15625 vdd.n2194 vdd.n2193 185
R15626 vdd.n2196 vdd.n2195 185
R15627 vdd.n2198 vdd.n2197 185
R15628 vdd.n2200 vdd.n2199 185
R15629 vdd.n2202 vdd.n2201 185
R15630 vdd.n2204 vdd.n2203 185
R15631 vdd.n2206 vdd.n2205 185
R15632 vdd.n2208 vdd.n2207 185
R15633 vdd.n2210 vdd.n2209 185
R15634 vdd.n2212 vdd.n2211 185
R15635 vdd.n2214 vdd.n2213 185
R15636 vdd.n2215 vdd.n745 185
R15637 vdd.n2217 vdd.n2216 185
R15638 vdd.n2218 vdd.n2217 185
R15639 vdd.n2147 vdd.n749 185
R15640 vdd.n2147 vdd.n2146 185
R15641 vdd.n1768 vdd.n750 185
R15642 vdd.t2 vdd.n750 185
R15643 vdd.n1769 vdd.n760 185
R15644 vdd.n2071 vdd.n760 185
R15645 vdd.n1772 vdd.n1771 185
R15646 vdd.n1771 vdd.n1770 185
R15647 vdd.n1773 vdd.n767 185
R15648 vdd.n2064 vdd.n767 185
R15649 vdd.n1775 vdd.n1774 185
R15650 vdd.n1774 vdd.n766 185
R15651 vdd.n1776 vdd.n774 185
R15652 vdd.n2056 vdd.n774 185
R15653 vdd.n1778 vdd.n1777 185
R15654 vdd.n1777 vdd.n773 185
R15655 vdd.n1779 vdd.n780 185
R15656 vdd.n2050 vdd.n780 185
R15657 vdd.n1781 vdd.n1780 185
R15658 vdd.n1780 vdd.n779 185
R15659 vdd.n1782 vdd.n785 185
R15660 vdd.n2044 vdd.n785 185
R15661 vdd.n1784 vdd.n1783 185
R15662 vdd.n1783 vdd.n792 185
R15663 vdd.n1785 vdd.n790 185
R15664 vdd.n2038 vdd.n790 185
R15665 vdd.n1787 vdd.n1786 185
R15666 vdd.n1786 vdd.n798 185
R15667 vdd.n1788 vdd.n796 185
R15668 vdd.n2032 vdd.n796 185
R15669 vdd.n1873 vdd.n1872 185
R15670 vdd.n1872 vdd.n1871 185
R15671 vdd.n1874 vdd.n803 185
R15672 vdd.n2026 vdd.n803 185
R15673 vdd.n1876 vdd.n1875 185
R15674 vdd.n1875 vdd.n802 185
R15675 vdd.n1877 vdd.n809 185
R15676 vdd.n2020 vdd.n809 185
R15677 vdd.n1879 vdd.n1878 185
R15678 vdd.n1878 vdd.n808 185
R15679 vdd.n1880 vdd.n814 185
R15680 vdd.n2014 vdd.n814 185
R15681 vdd.n1882 vdd.n1881 185
R15682 vdd.n1881 vdd.n823 185
R15683 vdd.n1883 vdd.n821 185
R15684 vdd.n2007 vdd.n821 185
R15685 vdd.n1885 vdd.n1884 185
R15686 vdd.n1884 vdd.n820 185
R15687 vdd.n1886 vdd.n828 185
R15688 vdd.n2001 vdd.n828 185
R15689 vdd.n1888 vdd.n1887 185
R15690 vdd.n1887 vdd.n827 185
R15691 vdd.n1889 vdd.n834 185
R15692 vdd.n1995 vdd.n834 185
R15693 vdd.n1891 vdd.n1890 185
R15694 vdd.n1890 vdd.n833 185
R15695 vdd.n1892 vdd.n840 185
R15696 vdd.n1989 vdd.n840 185
R15697 vdd.n3024 vdd.n3023 185
R15698 vdd.n3025 vdd.n3024 185
R15699 vdd.n325 vdd.n324 185
R15700 vdd.n3026 vdd.n325 185
R15701 vdd.n3029 vdd.n3028 185
R15702 vdd.n3028 vdd.n3027 185
R15703 vdd.n3030 vdd.n319 185
R15704 vdd.n319 vdd.n318 185
R15705 vdd.n3032 vdd.n3031 185
R15706 vdd.n3033 vdd.n3032 185
R15707 vdd.n314 vdd.n313 185
R15708 vdd.n3034 vdd.n314 185
R15709 vdd.n3037 vdd.n3036 185
R15710 vdd.n3036 vdd.n3035 185
R15711 vdd.n3038 vdd.n309 185
R15712 vdd.n309 vdd.n308 185
R15713 vdd.n3040 vdd.n3039 185
R15714 vdd.n3041 vdd.n3040 185
R15715 vdd.n303 vdd.n301 185
R15716 vdd.n3042 vdd.n303 185
R15717 vdd.n3045 vdd.n3044 185
R15718 vdd.n3044 vdd.n3043 185
R15719 vdd.n302 vdd.n300 185
R15720 vdd.n304 vdd.n302 185
R15721 vdd.n2881 vdd.n2880 185
R15722 vdd.n2882 vdd.n2881 185
R15723 vdd.n458 vdd.n457 185
R15724 vdd.n457 vdd.n456 185
R15725 vdd.n2876 vdd.n2875 185
R15726 vdd.n2875 vdd.n2874 185
R15727 vdd.n461 vdd.n460 185
R15728 vdd.n467 vdd.n461 185
R15729 vdd.n2865 vdd.n2864 185
R15730 vdd.n2866 vdd.n2865 185
R15731 vdd.n469 vdd.n468 185
R15732 vdd.n2857 vdd.n468 185
R15733 vdd.n2860 vdd.n2859 185
R15734 vdd.n2859 vdd.n2858 185
R15735 vdd.n472 vdd.n471 185
R15736 vdd.n473 vdd.n472 185
R15737 vdd.n2848 vdd.n2847 185
R15738 vdd.n2849 vdd.n2848 185
R15739 vdd.n480 vdd.n479 185
R15740 vdd.n516 vdd.n479 185
R15741 vdd.n2843 vdd.n2842 185
R15742 vdd.n483 vdd.n482 185
R15743 vdd.n2839 vdd.n2838 185
R15744 vdd.n2840 vdd.n2839 185
R15745 vdd.n518 vdd.n517 185
R15746 vdd.n522 vdd.n521 185
R15747 vdd.n2834 vdd.n523 185
R15748 vdd.n2833 vdd.n2832 185
R15749 vdd.n2831 vdd.n2830 185
R15750 vdd.n2829 vdd.n2828 185
R15751 vdd.n2827 vdd.n2826 185
R15752 vdd.n2825 vdd.n2824 185
R15753 vdd.n2823 vdd.n2822 185
R15754 vdd.n2821 vdd.n2820 185
R15755 vdd.n2819 vdd.n2818 185
R15756 vdd.n2817 vdd.n2816 185
R15757 vdd.n2815 vdd.n2814 185
R15758 vdd.n2813 vdd.n2812 185
R15759 vdd.n2811 vdd.n2810 185
R15760 vdd.n2809 vdd.n2808 185
R15761 vdd.n2807 vdd.n2806 185
R15762 vdd.n2798 vdd.n536 185
R15763 vdd.n2800 vdd.n2799 185
R15764 vdd.n2797 vdd.n2796 185
R15765 vdd.n2795 vdd.n2794 185
R15766 vdd.n2793 vdd.n2792 185
R15767 vdd.n2791 vdd.n2790 185
R15768 vdd.n2789 vdd.n2788 185
R15769 vdd.n2787 vdd.n2786 185
R15770 vdd.n2785 vdd.n2784 185
R15771 vdd.n2783 vdd.n2782 185
R15772 vdd.n2781 vdd.n2780 185
R15773 vdd.n2779 vdd.n2778 185
R15774 vdd.n2777 vdd.n2776 185
R15775 vdd.n2775 vdd.n2774 185
R15776 vdd.n2773 vdd.n2772 185
R15777 vdd.n2771 vdd.n2770 185
R15778 vdd.n2769 vdd.n2768 185
R15779 vdd.n2767 vdd.n2766 185
R15780 vdd.n2765 vdd.n2764 185
R15781 vdd.n2763 vdd.n2762 185
R15782 vdd.n2761 vdd.n2760 185
R15783 vdd.n2759 vdd.n2758 185
R15784 vdd.n2752 vdd.n556 185
R15785 vdd.n2754 vdd.n2753 185
R15786 vdd.n2751 vdd.n2750 185
R15787 vdd.n2749 vdd.n2748 185
R15788 vdd.n2747 vdd.n2746 185
R15789 vdd.n2745 vdd.n2744 185
R15790 vdd.n2743 vdd.n2742 185
R15791 vdd.n2741 vdd.n2740 185
R15792 vdd.n2739 vdd.n2738 185
R15793 vdd.n2737 vdd.n2736 185
R15794 vdd.n2735 vdd.n2734 185
R15795 vdd.n2733 vdd.n2732 185
R15796 vdd.n2731 vdd.n2730 185
R15797 vdd.n2729 vdd.n2728 185
R15798 vdd.n2727 vdd.n2726 185
R15799 vdd.n2725 vdd.n2724 185
R15800 vdd.n2723 vdd.n2722 185
R15801 vdd.n2721 vdd.n2720 185
R15802 vdd.n2719 vdd.n2718 185
R15803 vdd.n2717 vdd.n2716 185
R15804 vdd.n2715 vdd.n2714 185
R15805 vdd.n2710 vdd.n515 185
R15806 vdd.n2840 vdd.n515 185
R15807 vdd.n2907 vdd.n2906 185
R15808 vdd.n2911 vdd.n440 185
R15809 vdd.n2913 vdd.n2912 185
R15810 vdd.n2915 vdd.n438 185
R15811 vdd.n2917 vdd.n2916 185
R15812 vdd.n2918 vdd.n433 185
R15813 vdd.n2920 vdd.n2919 185
R15814 vdd.n2922 vdd.n431 185
R15815 vdd.n2924 vdd.n2923 185
R15816 vdd.n2925 vdd.n426 185
R15817 vdd.n2927 vdd.n2926 185
R15818 vdd.n2929 vdd.n424 185
R15819 vdd.n2931 vdd.n2930 185
R15820 vdd.n2932 vdd.n419 185
R15821 vdd.n2934 vdd.n2933 185
R15822 vdd.n2936 vdd.n417 185
R15823 vdd.n2938 vdd.n2937 185
R15824 vdd.n2939 vdd.n413 185
R15825 vdd.n2941 vdd.n2940 185
R15826 vdd.n2943 vdd.n410 185
R15827 vdd.n2945 vdd.n2944 185
R15828 vdd.n411 vdd.n404 185
R15829 vdd.n2949 vdd.n408 185
R15830 vdd.n2950 vdd.n400 185
R15831 vdd.n2952 vdd.n2951 185
R15832 vdd.n2954 vdd.n398 185
R15833 vdd.n2956 vdd.n2955 185
R15834 vdd.n2957 vdd.n393 185
R15835 vdd.n2959 vdd.n2958 185
R15836 vdd.n2961 vdd.n391 185
R15837 vdd.n2963 vdd.n2962 185
R15838 vdd.n2964 vdd.n386 185
R15839 vdd.n2966 vdd.n2965 185
R15840 vdd.n2968 vdd.n384 185
R15841 vdd.n2970 vdd.n2969 185
R15842 vdd.n2971 vdd.n379 185
R15843 vdd.n2973 vdd.n2972 185
R15844 vdd.n2975 vdd.n377 185
R15845 vdd.n2977 vdd.n2976 185
R15846 vdd.n2978 vdd.n373 185
R15847 vdd.n2980 vdd.n2979 185
R15848 vdd.n2982 vdd.n370 185
R15849 vdd.n2984 vdd.n2983 185
R15850 vdd.n371 vdd.n364 185
R15851 vdd.n2988 vdd.n368 185
R15852 vdd.n2989 vdd.n360 185
R15853 vdd.n2991 vdd.n2990 185
R15854 vdd.n2993 vdd.n358 185
R15855 vdd.n2995 vdd.n2994 185
R15856 vdd.n2996 vdd.n353 185
R15857 vdd.n2998 vdd.n2997 185
R15858 vdd.n3000 vdd.n351 185
R15859 vdd.n3002 vdd.n3001 185
R15860 vdd.n3003 vdd.n346 185
R15861 vdd.n3005 vdd.n3004 185
R15862 vdd.n3007 vdd.n344 185
R15863 vdd.n3009 vdd.n3008 185
R15864 vdd.n3010 vdd.n338 185
R15865 vdd.n3012 vdd.n3011 185
R15866 vdd.n3014 vdd.n337 185
R15867 vdd.n3015 vdd.n336 185
R15868 vdd.n3018 vdd.n3017 185
R15869 vdd.n3019 vdd.n334 185
R15870 vdd.n3020 vdd.n330 185
R15871 vdd.n2902 vdd.n328 185
R15872 vdd.n3025 vdd.n328 185
R15873 vdd.n2901 vdd.n327 185
R15874 vdd.n3026 vdd.n327 185
R15875 vdd.n2900 vdd.n326 185
R15876 vdd.n3027 vdd.n326 185
R15877 vdd.n446 vdd.n445 185
R15878 vdd.n445 vdd.n318 185
R15879 vdd.n2896 vdd.n317 185
R15880 vdd.n3033 vdd.n317 185
R15881 vdd.n2895 vdd.n316 185
R15882 vdd.n3034 vdd.n316 185
R15883 vdd.n2894 vdd.n315 185
R15884 vdd.n3035 vdd.n315 185
R15885 vdd.n449 vdd.n448 185
R15886 vdd.n448 vdd.n308 185
R15887 vdd.n2890 vdd.n307 185
R15888 vdd.n3041 vdd.n307 185
R15889 vdd.n2889 vdd.n306 185
R15890 vdd.n3042 vdd.n306 185
R15891 vdd.n2888 vdd.n305 185
R15892 vdd.n3043 vdd.n305 185
R15893 vdd.n455 vdd.n451 185
R15894 vdd.n455 vdd.n304 185
R15895 vdd.n2884 vdd.n2883 185
R15896 vdd.n2883 vdd.n2882 185
R15897 vdd.n454 vdd.n453 185
R15898 vdd.n456 vdd.n454 185
R15899 vdd.n2873 vdd.n2872 185
R15900 vdd.n2874 vdd.n2873 185
R15901 vdd.n463 vdd.n462 185
R15902 vdd.n467 vdd.n462 185
R15903 vdd.n2868 vdd.n2867 185
R15904 vdd.n2867 vdd.n2866 185
R15905 vdd.n466 vdd.n465 185
R15906 vdd.n2857 vdd.n466 185
R15907 vdd.n2856 vdd.n2855 185
R15908 vdd.n2858 vdd.n2856 185
R15909 vdd.n475 vdd.n474 185
R15910 vdd.n474 vdd.n473 185
R15911 vdd.n2851 vdd.n2850 185
R15912 vdd.n2850 vdd.n2849 185
R15913 vdd.n478 vdd.n477 185
R15914 vdd.n516 vdd.n478 185
R15915 vdd.n703 vdd.n702 185
R15916 vdd.n2469 vdd.n2468 185
R15917 vdd.n2467 vdd.n2252 185
R15918 vdd.n2471 vdd.n2252 185
R15919 vdd.n2466 vdd.n2465 185
R15920 vdd.n2464 vdd.n2463 185
R15921 vdd.n2462 vdd.n2461 185
R15922 vdd.n2460 vdd.n2459 185
R15923 vdd.n2458 vdd.n2457 185
R15924 vdd.n2456 vdd.n2455 185
R15925 vdd.n2454 vdd.n2453 185
R15926 vdd.n2452 vdd.n2451 185
R15927 vdd.n2450 vdd.n2449 185
R15928 vdd.n2448 vdd.n2447 185
R15929 vdd.n2446 vdd.n2445 185
R15930 vdd.n2444 vdd.n2443 185
R15931 vdd.n2442 vdd.n2441 185
R15932 vdd.n2440 vdd.n2439 185
R15933 vdd.n2438 vdd.n2437 185
R15934 vdd.n2436 vdd.n2435 185
R15935 vdd.n2434 vdd.n2433 185
R15936 vdd.n2432 vdd.n2431 185
R15937 vdd.n2430 vdd.n2429 185
R15938 vdd.n2428 vdd.n2427 185
R15939 vdd.n2426 vdd.n2425 185
R15940 vdd.n2424 vdd.n2423 185
R15941 vdd.n2422 vdd.n2421 185
R15942 vdd.n2420 vdd.n2419 185
R15943 vdd.n2418 vdd.n2417 185
R15944 vdd.n2416 vdd.n2415 185
R15945 vdd.n2414 vdd.n2413 185
R15946 vdd.n2412 vdd.n2411 185
R15947 vdd.n2410 vdd.n2409 185
R15948 vdd.n2407 vdd.n2406 185
R15949 vdd.n2405 vdd.n2404 185
R15950 vdd.n2403 vdd.n2402 185
R15951 vdd.n2609 vdd.n2608 185
R15952 vdd.n2611 vdd.n624 185
R15953 vdd.n2613 vdd.n2612 185
R15954 vdd.n2615 vdd.n621 185
R15955 vdd.n2617 vdd.n2616 185
R15956 vdd.n2619 vdd.n619 185
R15957 vdd.n2621 vdd.n2620 185
R15958 vdd.n2622 vdd.n618 185
R15959 vdd.n2624 vdd.n2623 185
R15960 vdd.n2626 vdd.n616 185
R15961 vdd.n2628 vdd.n2627 185
R15962 vdd.n2629 vdd.n615 185
R15963 vdd.n2631 vdd.n2630 185
R15964 vdd.n2633 vdd.n613 185
R15965 vdd.n2635 vdd.n2634 185
R15966 vdd.n2636 vdd.n612 185
R15967 vdd.n2638 vdd.n2637 185
R15968 vdd.n2640 vdd.n520 185
R15969 vdd.n2642 vdd.n2641 185
R15970 vdd.n2644 vdd.n610 185
R15971 vdd.n2646 vdd.n2645 185
R15972 vdd.n2647 vdd.n609 185
R15973 vdd.n2649 vdd.n2648 185
R15974 vdd.n2651 vdd.n607 185
R15975 vdd.n2653 vdd.n2652 185
R15976 vdd.n2654 vdd.n606 185
R15977 vdd.n2656 vdd.n2655 185
R15978 vdd.n2658 vdd.n604 185
R15979 vdd.n2660 vdd.n2659 185
R15980 vdd.n2661 vdd.n603 185
R15981 vdd.n2663 vdd.n2662 185
R15982 vdd.n2665 vdd.n602 185
R15983 vdd.n2666 vdd.n601 185
R15984 vdd.n2669 vdd.n2668 185
R15985 vdd.n2670 vdd.n599 185
R15986 vdd.n599 vdd.n484 185
R15987 vdd.n2607 vdd.n596 185
R15988 vdd.n2673 vdd.n596 185
R15989 vdd.n2606 vdd.n2605 185
R15990 vdd.n2605 vdd.n595 185
R15991 vdd.n2604 vdd.n626 185
R15992 vdd.n2604 vdd.n2603 185
R15993 vdd.n2358 vdd.n627 185
R15994 vdd.n636 vdd.n627 185
R15995 vdd.n2359 vdd.n634 185
R15996 vdd.n2597 vdd.n634 185
R15997 vdd.n2361 vdd.n2360 185
R15998 vdd.n2360 vdd.n633 185
R15999 vdd.n2362 vdd.n642 185
R16000 vdd.n2546 vdd.n642 185
R16001 vdd.n2364 vdd.n2363 185
R16002 vdd.n2363 vdd.n641 185
R16003 vdd.n2365 vdd.n648 185
R16004 vdd.n2540 vdd.n648 185
R16005 vdd.n2367 vdd.n2366 185
R16006 vdd.n2366 vdd.n647 185
R16007 vdd.n2368 vdd.n653 185
R16008 vdd.n2532 vdd.n653 185
R16009 vdd.n2370 vdd.n2369 185
R16010 vdd.n2369 vdd.n660 185
R16011 vdd.n2371 vdd.n658 185
R16012 vdd.n2526 vdd.n658 185
R16013 vdd.n2373 vdd.n2372 185
R16014 vdd.n2374 vdd.n2373 185
R16015 vdd.n2357 vdd.n665 185
R16016 vdd.n2520 vdd.n665 185
R16017 vdd.n2356 vdd.n2355 185
R16018 vdd.n2355 vdd.n664 185
R16019 vdd.n2354 vdd.n671 185
R16020 vdd.n2514 vdd.n671 185
R16021 vdd.n2353 vdd.n2352 185
R16022 vdd.n2352 vdd.n670 185
R16023 vdd.n2351 vdd.n676 185
R16024 vdd.n2508 vdd.n676 185
R16025 vdd.n2350 vdd.n2349 185
R16026 vdd.n2349 vdd.n683 185
R16027 vdd.n2348 vdd.n681 185
R16028 vdd.n2502 vdd.n681 185
R16029 vdd.n2347 vdd.n2346 185
R16030 vdd.n2346 vdd.n690 185
R16031 vdd.n2345 vdd.n688 185
R16032 vdd.n2496 vdd.n688 185
R16033 vdd.n2344 vdd.n2343 185
R16034 vdd.n2343 vdd.n687 185
R16035 vdd.n2255 vdd.n694 185
R16036 vdd.n2490 vdd.n694 185
R16037 vdd.n2397 vdd.n2396 185
R16038 vdd.n2396 vdd.n2395 185
R16039 vdd.n2398 vdd.n699 185
R16040 vdd.n2484 vdd.n699 185
R16041 vdd.n2400 vdd.n2399 185
R16042 vdd.n2399 vdd.t21 185
R16043 vdd.n2401 vdd.n704 185
R16044 vdd.n2478 vdd.n704 185
R16045 vdd.n2480 vdd.n2479 185
R16046 vdd.n2479 vdd.n2478 185
R16047 vdd.n2481 vdd.n701 185
R16048 vdd.n701 vdd.t21 185
R16049 vdd.n2483 vdd.n2482 185
R16050 vdd.n2484 vdd.n2483 185
R16051 vdd.n693 vdd.n692 185
R16052 vdd.n2395 vdd.n693 185
R16053 vdd.n2492 vdd.n2491 185
R16054 vdd.n2491 vdd.n2490 185
R16055 vdd.n2493 vdd.n691 185
R16056 vdd.n691 vdd.n687 185
R16057 vdd.n2495 vdd.n2494 185
R16058 vdd.n2496 vdd.n2495 185
R16059 vdd.n680 vdd.n679 185
R16060 vdd.n690 vdd.n680 185
R16061 vdd.n2504 vdd.n2503 185
R16062 vdd.n2503 vdd.n2502 185
R16063 vdd.n2505 vdd.n678 185
R16064 vdd.n683 vdd.n678 185
R16065 vdd.n2507 vdd.n2506 185
R16066 vdd.n2508 vdd.n2507 185
R16067 vdd.n669 vdd.n668 185
R16068 vdd.n670 vdd.n669 185
R16069 vdd.n2516 vdd.n2515 185
R16070 vdd.n2515 vdd.n2514 185
R16071 vdd.n2517 vdd.n667 185
R16072 vdd.n667 vdd.n664 185
R16073 vdd.n2519 vdd.n2518 185
R16074 vdd.n2520 vdd.n2519 185
R16075 vdd.n657 vdd.n656 185
R16076 vdd.n2374 vdd.n657 185
R16077 vdd.n2528 vdd.n2527 185
R16078 vdd.n2527 vdd.n2526 185
R16079 vdd.n2529 vdd.n655 185
R16080 vdd.n660 vdd.n655 185
R16081 vdd.n2531 vdd.n2530 185
R16082 vdd.n2532 vdd.n2531 185
R16083 vdd.n646 vdd.n645 185
R16084 vdd.n647 vdd.n646 185
R16085 vdd.n2542 vdd.n2541 185
R16086 vdd.n2541 vdd.n2540 185
R16087 vdd.n2543 vdd.n644 185
R16088 vdd.n644 vdd.n641 185
R16089 vdd.n2545 vdd.n2544 185
R16090 vdd.n2546 vdd.n2545 185
R16091 vdd.n632 vdd.n631 185
R16092 vdd.n633 vdd.n632 185
R16093 vdd.n2599 vdd.n2598 185
R16094 vdd.n2598 vdd.n2597 185
R16095 vdd.n2600 vdd.n630 185
R16096 vdd.n636 vdd.n630 185
R16097 vdd.n2602 vdd.n2601 185
R16098 vdd.n2603 vdd.n2602 185
R16099 vdd.n600 vdd.n598 185
R16100 vdd.n598 vdd.n595 185
R16101 vdd.n2672 vdd.n2671 185
R16102 vdd.n2673 vdd.n2672 185
R16103 vdd.n2145 vdd.n2144 185
R16104 vdd.n2146 vdd.n2145 185
R16105 vdd.n754 vdd.n752 185
R16106 vdd.n752 vdd.t2 185
R16107 vdd.n2060 vdd.n761 185
R16108 vdd.n2071 vdd.n761 185
R16109 vdd.n2061 vdd.n770 185
R16110 vdd.n1770 vdd.n770 185
R16111 vdd.n2063 vdd.n2062 185
R16112 vdd.n2064 vdd.n2063 185
R16113 vdd.n2059 vdd.n769 185
R16114 vdd.n769 vdd.n766 185
R16115 vdd.n2058 vdd.n2057 185
R16116 vdd.n2057 vdd.n2056 185
R16117 vdd.n772 vdd.n771 185
R16118 vdd.n773 vdd.n772 185
R16119 vdd.n2049 vdd.n2048 185
R16120 vdd.n2050 vdd.n2049 185
R16121 vdd.n2047 vdd.n782 185
R16122 vdd.n782 vdd.n779 185
R16123 vdd.n2046 vdd.n2045 185
R16124 vdd.n2045 vdd.n2044 185
R16125 vdd.n784 vdd.n783 185
R16126 vdd.n792 vdd.n784 185
R16127 vdd.n2037 vdd.n2036 185
R16128 vdd.n2038 vdd.n2037 185
R16129 vdd.n2035 vdd.n793 185
R16130 vdd.n798 vdd.n793 185
R16131 vdd.n2034 vdd.n2033 185
R16132 vdd.n2033 vdd.n2032 185
R16133 vdd.n795 vdd.n794 185
R16134 vdd.n1871 vdd.n795 185
R16135 vdd.n2025 vdd.n2024 185
R16136 vdd.n2026 vdd.n2025 185
R16137 vdd.n2023 vdd.n805 185
R16138 vdd.n805 vdd.n802 185
R16139 vdd.n2022 vdd.n2021 185
R16140 vdd.n2021 vdd.n2020 185
R16141 vdd.n807 vdd.n806 185
R16142 vdd.n808 vdd.n807 185
R16143 vdd.n2013 vdd.n2012 185
R16144 vdd.n2014 vdd.n2013 185
R16145 vdd.n2010 vdd.n816 185
R16146 vdd.n823 vdd.n816 185
R16147 vdd.n2009 vdd.n2008 185
R16148 vdd.n2008 vdd.n2007 185
R16149 vdd.n819 vdd.n818 185
R16150 vdd.n820 vdd.n819 185
R16151 vdd.n2000 vdd.n1999 185
R16152 vdd.n2001 vdd.n2000 185
R16153 vdd.n1998 vdd.n830 185
R16154 vdd.n830 vdd.n827 185
R16155 vdd.n1997 vdd.n1996 185
R16156 vdd.n1996 vdd.n1995 185
R16157 vdd.n832 vdd.n831 185
R16158 vdd.n833 vdd.n832 185
R16159 vdd.n1988 vdd.n1987 185
R16160 vdd.n1989 vdd.n1988 185
R16161 vdd.n2076 vdd.n726 185
R16162 vdd.n2218 vdd.n726 185
R16163 vdd.n2078 vdd.n2077 185
R16164 vdd.n2080 vdd.n2079 185
R16165 vdd.n2082 vdd.n2081 185
R16166 vdd.n2084 vdd.n2083 185
R16167 vdd.n2086 vdd.n2085 185
R16168 vdd.n2088 vdd.n2087 185
R16169 vdd.n2090 vdd.n2089 185
R16170 vdd.n2092 vdd.n2091 185
R16171 vdd.n2094 vdd.n2093 185
R16172 vdd.n2096 vdd.n2095 185
R16173 vdd.n2098 vdd.n2097 185
R16174 vdd.n2100 vdd.n2099 185
R16175 vdd.n2102 vdd.n2101 185
R16176 vdd.n2104 vdd.n2103 185
R16177 vdd.n2106 vdd.n2105 185
R16178 vdd.n2108 vdd.n2107 185
R16179 vdd.n2110 vdd.n2109 185
R16180 vdd.n2112 vdd.n2111 185
R16181 vdd.n2114 vdd.n2113 185
R16182 vdd.n2116 vdd.n2115 185
R16183 vdd.n2118 vdd.n2117 185
R16184 vdd.n2120 vdd.n2119 185
R16185 vdd.n2122 vdd.n2121 185
R16186 vdd.n2124 vdd.n2123 185
R16187 vdd.n2126 vdd.n2125 185
R16188 vdd.n2128 vdd.n2127 185
R16189 vdd.n2130 vdd.n2129 185
R16190 vdd.n2132 vdd.n2131 185
R16191 vdd.n2134 vdd.n2133 185
R16192 vdd.n2136 vdd.n2135 185
R16193 vdd.n2138 vdd.n2137 185
R16194 vdd.n2140 vdd.n2139 185
R16195 vdd.n2142 vdd.n2141 185
R16196 vdd.n2143 vdd.n753 185
R16197 vdd.n2075 vdd.n751 185
R16198 vdd.n2146 vdd.n751 185
R16199 vdd.n2074 vdd.n2073 185
R16200 vdd.n2073 vdd.t2 185
R16201 vdd.n2072 vdd.n758 185
R16202 vdd.n2072 vdd.n2071 185
R16203 vdd.n1852 vdd.n759 185
R16204 vdd.n1770 vdd.n759 185
R16205 vdd.n1853 vdd.n768 185
R16206 vdd.n2064 vdd.n768 185
R16207 vdd.n1855 vdd.n1854 185
R16208 vdd.n1854 vdd.n766 185
R16209 vdd.n1856 vdd.n775 185
R16210 vdd.n2056 vdd.n775 185
R16211 vdd.n1858 vdd.n1857 185
R16212 vdd.n1857 vdd.n773 185
R16213 vdd.n1859 vdd.n781 185
R16214 vdd.n2050 vdd.n781 185
R16215 vdd.n1861 vdd.n1860 185
R16216 vdd.n1860 vdd.n779 185
R16217 vdd.n1862 vdd.n786 185
R16218 vdd.n2044 vdd.n786 185
R16219 vdd.n1864 vdd.n1863 185
R16220 vdd.n1863 vdd.n792 185
R16221 vdd.n1865 vdd.n791 185
R16222 vdd.n2038 vdd.n791 185
R16223 vdd.n1867 vdd.n1866 185
R16224 vdd.n1866 vdd.n798 185
R16225 vdd.n1868 vdd.n797 185
R16226 vdd.n2032 vdd.n797 185
R16227 vdd.n1870 vdd.n1869 185
R16228 vdd.n1871 vdd.n1870 185
R16229 vdd.n1851 vdd.n804 185
R16230 vdd.n2026 vdd.n804 185
R16231 vdd.n1850 vdd.n1849 185
R16232 vdd.n1849 vdd.n802 185
R16233 vdd.n1848 vdd.n810 185
R16234 vdd.n2020 vdd.n810 185
R16235 vdd.n1847 vdd.n1846 185
R16236 vdd.n1846 vdd.n808 185
R16237 vdd.n1845 vdd.n815 185
R16238 vdd.n2014 vdd.n815 185
R16239 vdd.n1844 vdd.n1843 185
R16240 vdd.n1843 vdd.n823 185
R16241 vdd.n1842 vdd.n822 185
R16242 vdd.n2007 vdd.n822 185
R16243 vdd.n1841 vdd.n1840 185
R16244 vdd.n1840 vdd.n820 185
R16245 vdd.n1839 vdd.n829 185
R16246 vdd.n2001 vdd.n829 185
R16247 vdd.n1838 vdd.n1837 185
R16248 vdd.n1837 vdd.n827 185
R16249 vdd.n1836 vdd.n835 185
R16250 vdd.n1995 vdd.n835 185
R16251 vdd.n1835 vdd.n1834 185
R16252 vdd.n1834 vdd.n833 185
R16253 vdd.n1833 vdd.n841 185
R16254 vdd.n1989 vdd.n841 185
R16255 vdd.n1986 vdd.n842 185
R16256 vdd.n1985 vdd.n1984 185
R16257 vdd.n1982 vdd.n843 185
R16258 vdd.n1980 vdd.n1979 185
R16259 vdd.n1978 vdd.n844 185
R16260 vdd.n1977 vdd.n1976 185
R16261 vdd.n1974 vdd.n845 185
R16262 vdd.n1972 vdd.n1971 185
R16263 vdd.n1970 vdd.n846 185
R16264 vdd.n1969 vdd.n1968 185
R16265 vdd.n1966 vdd.n847 185
R16266 vdd.n1964 vdd.n1963 185
R16267 vdd.n1962 vdd.n848 185
R16268 vdd.n1961 vdd.n1960 185
R16269 vdd.n1958 vdd.n849 185
R16270 vdd.n1956 vdd.n1955 185
R16271 vdd.n1954 vdd.n850 185
R16272 vdd.n1953 vdd.n852 185
R16273 vdd.n1798 vdd.n853 185
R16274 vdd.n1801 vdd.n1800 185
R16275 vdd.n1803 vdd.n1802 185
R16276 vdd.n1805 vdd.n1797 185
R16277 vdd.n1808 vdd.n1807 185
R16278 vdd.n1809 vdd.n1796 185
R16279 vdd.n1811 vdd.n1810 185
R16280 vdd.n1813 vdd.n1795 185
R16281 vdd.n1816 vdd.n1815 185
R16282 vdd.n1817 vdd.n1794 185
R16283 vdd.n1819 vdd.n1818 185
R16284 vdd.n1821 vdd.n1793 185
R16285 vdd.n1824 vdd.n1823 185
R16286 vdd.n1825 vdd.n1790 185
R16287 vdd.n1828 vdd.n1827 185
R16288 vdd.n1830 vdd.n1789 185
R16289 vdd.n1832 vdd.n1831 185
R16290 vdd.n1831 vdd.n839 185
R16291 vdd.n291 vdd.n290 171.744
R16292 vdd.n290 vdd.n289 171.744
R16293 vdd.n289 vdd.n258 171.744
R16294 vdd.n282 vdd.n258 171.744
R16295 vdd.n282 vdd.n281 171.744
R16296 vdd.n281 vdd.n263 171.744
R16297 vdd.n274 vdd.n263 171.744
R16298 vdd.n274 vdd.n273 171.744
R16299 vdd.n273 vdd.n267 171.744
R16300 vdd.n244 vdd.n243 171.744
R16301 vdd.n243 vdd.n242 171.744
R16302 vdd.n242 vdd.n211 171.744
R16303 vdd.n235 vdd.n211 171.744
R16304 vdd.n235 vdd.n234 171.744
R16305 vdd.n234 vdd.n216 171.744
R16306 vdd.n227 vdd.n216 171.744
R16307 vdd.n227 vdd.n226 171.744
R16308 vdd.n226 vdd.n220 171.744
R16309 vdd.n201 vdd.n200 171.744
R16310 vdd.n200 vdd.n199 171.744
R16311 vdd.n199 vdd.n168 171.744
R16312 vdd.n192 vdd.n168 171.744
R16313 vdd.n192 vdd.n191 171.744
R16314 vdd.n191 vdd.n173 171.744
R16315 vdd.n184 vdd.n173 171.744
R16316 vdd.n184 vdd.n183 171.744
R16317 vdd.n183 vdd.n177 171.744
R16318 vdd.n154 vdd.n153 171.744
R16319 vdd.n153 vdd.n152 171.744
R16320 vdd.n152 vdd.n121 171.744
R16321 vdd.n145 vdd.n121 171.744
R16322 vdd.n145 vdd.n144 171.744
R16323 vdd.n144 vdd.n126 171.744
R16324 vdd.n137 vdd.n126 171.744
R16325 vdd.n137 vdd.n136 171.744
R16326 vdd.n136 vdd.n130 171.744
R16327 vdd.n112 vdd.n111 171.744
R16328 vdd.n111 vdd.n110 171.744
R16329 vdd.n110 vdd.n79 171.744
R16330 vdd.n103 vdd.n79 171.744
R16331 vdd.n103 vdd.n102 171.744
R16332 vdd.n102 vdd.n84 171.744
R16333 vdd.n95 vdd.n84 171.744
R16334 vdd.n95 vdd.n94 171.744
R16335 vdd.n94 vdd.n88 171.744
R16336 vdd.n65 vdd.n64 171.744
R16337 vdd.n64 vdd.n63 171.744
R16338 vdd.n63 vdd.n32 171.744
R16339 vdd.n56 vdd.n32 171.744
R16340 vdd.n56 vdd.n55 171.744
R16341 vdd.n55 vdd.n37 171.744
R16342 vdd.n48 vdd.n37 171.744
R16343 vdd.n48 vdd.n47 171.744
R16344 vdd.n47 vdd.n41 171.744
R16345 vdd.n1106 vdd.n1105 171.744
R16346 vdd.n1105 vdd.n1104 171.744
R16347 vdd.n1104 vdd.n1073 171.744
R16348 vdd.n1097 vdd.n1073 171.744
R16349 vdd.n1097 vdd.n1096 171.744
R16350 vdd.n1096 vdd.n1078 171.744
R16351 vdd.n1089 vdd.n1078 171.744
R16352 vdd.n1089 vdd.n1088 171.744
R16353 vdd.n1088 vdd.n1082 171.744
R16354 vdd.n1153 vdd.n1152 171.744
R16355 vdd.n1152 vdd.n1151 171.744
R16356 vdd.n1151 vdd.n1120 171.744
R16357 vdd.n1144 vdd.n1120 171.744
R16358 vdd.n1144 vdd.n1143 171.744
R16359 vdd.n1143 vdd.n1125 171.744
R16360 vdd.n1136 vdd.n1125 171.744
R16361 vdd.n1136 vdd.n1135 171.744
R16362 vdd.n1135 vdd.n1129 171.744
R16363 vdd.n1016 vdd.n1015 171.744
R16364 vdd.n1015 vdd.n1014 171.744
R16365 vdd.n1014 vdd.n983 171.744
R16366 vdd.n1007 vdd.n983 171.744
R16367 vdd.n1007 vdd.n1006 171.744
R16368 vdd.n1006 vdd.n988 171.744
R16369 vdd.n999 vdd.n988 171.744
R16370 vdd.n999 vdd.n998 171.744
R16371 vdd.n998 vdd.n992 171.744
R16372 vdd.n1063 vdd.n1062 171.744
R16373 vdd.n1062 vdd.n1061 171.744
R16374 vdd.n1061 vdd.n1030 171.744
R16375 vdd.n1054 vdd.n1030 171.744
R16376 vdd.n1054 vdd.n1053 171.744
R16377 vdd.n1053 vdd.n1035 171.744
R16378 vdd.n1046 vdd.n1035 171.744
R16379 vdd.n1046 vdd.n1045 171.744
R16380 vdd.n1045 vdd.n1039 171.744
R16381 vdd.n927 vdd.n926 171.744
R16382 vdd.n926 vdd.n925 171.744
R16383 vdd.n925 vdd.n894 171.744
R16384 vdd.n918 vdd.n894 171.744
R16385 vdd.n918 vdd.n917 171.744
R16386 vdd.n917 vdd.n899 171.744
R16387 vdd.n910 vdd.n899 171.744
R16388 vdd.n910 vdd.n909 171.744
R16389 vdd.n909 vdd.n903 171.744
R16390 vdd.n974 vdd.n973 171.744
R16391 vdd.n973 vdd.n972 171.744
R16392 vdd.n972 vdd.n941 171.744
R16393 vdd.n965 vdd.n941 171.744
R16394 vdd.n965 vdd.n964 171.744
R16395 vdd.n964 vdd.n946 171.744
R16396 vdd.n957 vdd.n946 171.744
R16397 vdd.n957 vdd.n956 171.744
R16398 vdd.n956 vdd.n950 171.744
R16399 vdd.n3017 vdd.n334 146.341
R16400 vdd.n3015 vdd.n3014 146.341
R16401 vdd.n3012 vdd.n338 146.341
R16402 vdd.n3008 vdd.n3007 146.341
R16403 vdd.n3005 vdd.n346 146.341
R16404 vdd.n3001 vdd.n3000 146.341
R16405 vdd.n2998 vdd.n353 146.341
R16406 vdd.n2994 vdd.n2993 146.341
R16407 vdd.n2991 vdd.n360 146.341
R16408 vdd.n371 vdd.n368 146.341
R16409 vdd.n2983 vdd.n2982 146.341
R16410 vdd.n2980 vdd.n373 146.341
R16411 vdd.n2976 vdd.n2975 146.341
R16412 vdd.n2973 vdd.n379 146.341
R16413 vdd.n2969 vdd.n2968 146.341
R16414 vdd.n2966 vdd.n386 146.341
R16415 vdd.n2962 vdd.n2961 146.341
R16416 vdd.n2959 vdd.n393 146.341
R16417 vdd.n2955 vdd.n2954 146.341
R16418 vdd.n2952 vdd.n400 146.341
R16419 vdd.n411 vdd.n408 146.341
R16420 vdd.n2944 vdd.n2943 146.341
R16421 vdd.n2941 vdd.n413 146.341
R16422 vdd.n2937 vdd.n2936 146.341
R16423 vdd.n2934 vdd.n419 146.341
R16424 vdd.n2930 vdd.n2929 146.341
R16425 vdd.n2927 vdd.n426 146.341
R16426 vdd.n2923 vdd.n2922 146.341
R16427 vdd.n2920 vdd.n433 146.341
R16428 vdd.n2916 vdd.n2915 146.341
R16429 vdd.n2913 vdd.n440 146.341
R16430 vdd.n2850 vdd.n478 146.341
R16431 vdd.n2850 vdd.n474 146.341
R16432 vdd.n2856 vdd.n474 146.341
R16433 vdd.n2856 vdd.n466 146.341
R16434 vdd.n2867 vdd.n466 146.341
R16435 vdd.n2867 vdd.n462 146.341
R16436 vdd.n2873 vdd.n462 146.341
R16437 vdd.n2873 vdd.n454 146.341
R16438 vdd.n2883 vdd.n454 146.341
R16439 vdd.n2883 vdd.n455 146.341
R16440 vdd.n455 vdd.n305 146.341
R16441 vdd.n306 vdd.n305 146.341
R16442 vdd.n307 vdd.n306 146.341
R16443 vdd.n448 vdd.n307 146.341
R16444 vdd.n448 vdd.n315 146.341
R16445 vdd.n316 vdd.n315 146.341
R16446 vdd.n317 vdd.n316 146.341
R16447 vdd.n445 vdd.n317 146.341
R16448 vdd.n445 vdd.n326 146.341
R16449 vdd.n327 vdd.n326 146.341
R16450 vdd.n328 vdd.n327 146.341
R16451 vdd.n2839 vdd.n483 146.341
R16452 vdd.n2839 vdd.n517 146.341
R16453 vdd.n523 vdd.n522 146.341
R16454 vdd.n2832 vdd.n2831 146.341
R16455 vdd.n2828 vdd.n2827 146.341
R16456 vdd.n2824 vdd.n2823 146.341
R16457 vdd.n2820 vdd.n2819 146.341
R16458 vdd.n2816 vdd.n2815 146.341
R16459 vdd.n2812 vdd.n2811 146.341
R16460 vdd.n2808 vdd.n2807 146.341
R16461 vdd.n2799 vdd.n2798 146.341
R16462 vdd.n2796 vdd.n2795 146.341
R16463 vdd.n2792 vdd.n2791 146.341
R16464 vdd.n2788 vdd.n2787 146.341
R16465 vdd.n2784 vdd.n2783 146.341
R16466 vdd.n2780 vdd.n2779 146.341
R16467 vdd.n2776 vdd.n2775 146.341
R16468 vdd.n2772 vdd.n2771 146.341
R16469 vdd.n2768 vdd.n2767 146.341
R16470 vdd.n2764 vdd.n2763 146.341
R16471 vdd.n2760 vdd.n2759 146.341
R16472 vdd.n2753 vdd.n2752 146.341
R16473 vdd.n2750 vdd.n2749 146.341
R16474 vdd.n2746 vdd.n2745 146.341
R16475 vdd.n2742 vdd.n2741 146.341
R16476 vdd.n2738 vdd.n2737 146.341
R16477 vdd.n2734 vdd.n2733 146.341
R16478 vdd.n2730 vdd.n2729 146.341
R16479 vdd.n2726 vdd.n2725 146.341
R16480 vdd.n2722 vdd.n2721 146.341
R16481 vdd.n2718 vdd.n2717 146.341
R16482 vdd.n2714 vdd.n515 146.341
R16483 vdd.n2848 vdd.n479 146.341
R16484 vdd.n2848 vdd.n472 146.341
R16485 vdd.n2859 vdd.n472 146.341
R16486 vdd.n2859 vdd.n468 146.341
R16487 vdd.n2865 vdd.n468 146.341
R16488 vdd.n2865 vdd.n461 146.341
R16489 vdd.n2875 vdd.n461 146.341
R16490 vdd.n2875 vdd.n457 146.341
R16491 vdd.n2881 vdd.n457 146.341
R16492 vdd.n2881 vdd.n302 146.341
R16493 vdd.n3044 vdd.n302 146.341
R16494 vdd.n3044 vdd.n303 146.341
R16495 vdd.n3040 vdd.n303 146.341
R16496 vdd.n3040 vdd.n309 146.341
R16497 vdd.n3036 vdd.n309 146.341
R16498 vdd.n3036 vdd.n314 146.341
R16499 vdd.n3032 vdd.n314 146.341
R16500 vdd.n3032 vdd.n319 146.341
R16501 vdd.n3028 vdd.n319 146.341
R16502 vdd.n3028 vdd.n325 146.341
R16503 vdd.n3024 vdd.n325 146.341
R16504 vdd.n1936 vdd.n1935 146.341
R16505 vdd.n1933 vdd.n1517 146.341
R16506 vdd.n1713 vdd.n1523 146.341
R16507 vdd.n1711 vdd.n1710 146.341
R16508 vdd.n1708 vdd.n1525 146.341
R16509 vdd.n1704 vdd.n1703 146.341
R16510 vdd.n1701 vdd.n1532 146.341
R16511 vdd.n1697 vdd.n1696 146.341
R16512 vdd.n1694 vdd.n1539 146.341
R16513 vdd.n1550 vdd.n1547 146.341
R16514 vdd.n1686 vdd.n1685 146.341
R16515 vdd.n1683 vdd.n1552 146.341
R16516 vdd.n1679 vdd.n1678 146.341
R16517 vdd.n1676 vdd.n1558 146.341
R16518 vdd.n1672 vdd.n1671 146.341
R16519 vdd.n1669 vdd.n1565 146.341
R16520 vdd.n1665 vdd.n1664 146.341
R16521 vdd.n1662 vdd.n1572 146.341
R16522 vdd.n1658 vdd.n1657 146.341
R16523 vdd.n1655 vdd.n1579 146.341
R16524 vdd.n1590 vdd.n1587 146.341
R16525 vdd.n1647 vdd.n1646 146.341
R16526 vdd.n1644 vdd.n1592 146.341
R16527 vdd.n1640 vdd.n1639 146.341
R16528 vdd.n1637 vdd.n1598 146.341
R16529 vdd.n1633 vdd.n1632 146.341
R16530 vdd.n1630 vdd.n1605 146.341
R16531 vdd.n1626 vdd.n1625 146.341
R16532 vdd.n1623 vdd.n1620 146.341
R16533 vdd.n1618 vdd.n1615 146.341
R16534 vdd.n1613 vdd.n859 146.341
R16535 vdd.n1431 vdd.n1191 146.341
R16536 vdd.n1431 vdd.n1187 146.341
R16537 vdd.n1437 vdd.n1187 146.341
R16538 vdd.n1437 vdd.n1179 146.341
R16539 vdd.n1448 vdd.n1179 146.341
R16540 vdd.n1448 vdd.n1175 146.341
R16541 vdd.n1454 vdd.n1175 146.341
R16542 vdd.n1454 vdd.n1169 146.341
R16543 vdd.n1466 vdd.n1169 146.341
R16544 vdd.n1466 vdd.n1165 146.341
R16545 vdd.n1472 vdd.n1165 146.341
R16546 vdd.n1472 vdd.n886 146.341
R16547 vdd.n1482 vdd.n886 146.341
R16548 vdd.n1482 vdd.n882 146.341
R16549 vdd.n1488 vdd.n882 146.341
R16550 vdd.n1488 vdd.n876 146.341
R16551 vdd.n1499 vdd.n876 146.341
R16552 vdd.n1499 vdd.n871 146.341
R16553 vdd.n1507 vdd.n871 146.341
R16554 vdd.n1507 vdd.n861 146.341
R16555 vdd.n1944 vdd.n861 146.341
R16556 vdd.n1420 vdd.n1196 146.341
R16557 vdd.n1420 vdd.n1229 146.341
R16558 vdd.n1233 vdd.n1232 146.341
R16559 vdd.n1235 vdd.n1234 146.341
R16560 vdd.n1239 vdd.n1238 146.341
R16561 vdd.n1241 vdd.n1240 146.341
R16562 vdd.n1245 vdd.n1244 146.341
R16563 vdd.n1247 vdd.n1246 146.341
R16564 vdd.n1251 vdd.n1250 146.341
R16565 vdd.n1253 vdd.n1252 146.341
R16566 vdd.n1259 vdd.n1258 146.341
R16567 vdd.n1261 vdd.n1260 146.341
R16568 vdd.n1265 vdd.n1264 146.341
R16569 vdd.n1267 vdd.n1266 146.341
R16570 vdd.n1271 vdd.n1270 146.341
R16571 vdd.n1273 vdd.n1272 146.341
R16572 vdd.n1277 vdd.n1276 146.341
R16573 vdd.n1279 vdd.n1278 146.341
R16574 vdd.n1283 vdd.n1282 146.341
R16575 vdd.n1285 vdd.n1284 146.341
R16576 vdd.n1357 vdd.n1288 146.341
R16577 vdd.n1290 vdd.n1289 146.341
R16578 vdd.n1294 vdd.n1293 146.341
R16579 vdd.n1296 vdd.n1295 146.341
R16580 vdd.n1300 vdd.n1299 146.341
R16581 vdd.n1302 vdd.n1301 146.341
R16582 vdd.n1306 vdd.n1305 146.341
R16583 vdd.n1308 vdd.n1307 146.341
R16584 vdd.n1312 vdd.n1311 146.341
R16585 vdd.n1314 vdd.n1313 146.341
R16586 vdd.n1318 vdd.n1317 146.341
R16587 vdd.n1319 vdd.n1227 146.341
R16588 vdd.n1429 vdd.n1192 146.341
R16589 vdd.n1429 vdd.n1185 146.341
R16590 vdd.n1440 vdd.n1185 146.341
R16591 vdd.n1440 vdd.n1181 146.341
R16592 vdd.n1446 vdd.n1181 146.341
R16593 vdd.n1446 vdd.n1174 146.341
R16594 vdd.n1457 vdd.n1174 146.341
R16595 vdd.n1457 vdd.n1170 146.341
R16596 vdd.n1464 vdd.n1170 146.341
R16597 vdd.n1464 vdd.n1163 146.341
R16598 vdd.n1474 vdd.n1163 146.341
R16599 vdd.n1474 vdd.n889 146.341
R16600 vdd.n1480 vdd.n889 146.341
R16601 vdd.n1480 vdd.n881 146.341
R16602 vdd.n1491 vdd.n881 146.341
R16603 vdd.n1491 vdd.n877 146.341
R16604 vdd.n1497 vdd.n877 146.341
R16605 vdd.n1497 vdd.n869 146.341
R16606 vdd.n1510 vdd.n869 146.341
R16607 vdd.n1510 vdd.n864 146.341
R16608 vdd.n1942 vdd.n864 146.341
R16609 vdd.n863 vdd.n839 141.707
R16610 vdd.n2840 vdd.n484 141.707
R16611 vdd.n1791 vdd.t174 127.284
R16612 vdd.n755 vdd.t158 127.284
R16613 vdd.n1765 vdd.t199 127.284
R16614 vdd.n747 vdd.t189 127.284
R16615 vdd.n2536 vdd.t141 127.284
R16616 vdd.n2536 vdd.t142 127.284
R16617 vdd.n2256 vdd.t181 127.284
R16618 vdd.n622 vdd.t162 127.284
R16619 vdd.n2253 vdd.t167 127.284
R16620 vdd.n589 vdd.t169 127.284
R16621 vdd.n817 vdd.t177 127.284
R16622 vdd.n817 vdd.t178 127.284
R16623 vdd.n22 vdd.n20 117.314
R16624 vdd.n17 vdd.n15 117.314
R16625 vdd.n27 vdd.n26 116.927
R16626 vdd.n24 vdd.n23 116.927
R16627 vdd.n22 vdd.n21 116.927
R16628 vdd.n17 vdd.n16 116.927
R16629 vdd.n19 vdd.n18 116.927
R16630 vdd.n27 vdd.n25 116.927
R16631 vdd.n1792 vdd.t173 111.188
R16632 vdd.n756 vdd.t159 111.188
R16633 vdd.n1766 vdd.t198 111.188
R16634 vdd.n748 vdd.t190 111.188
R16635 vdd.n2257 vdd.t180 111.188
R16636 vdd.n623 vdd.t163 111.188
R16637 vdd.n2254 vdd.t166 111.188
R16638 vdd.n590 vdd.t170 111.188
R16639 vdd.n2479 vdd.n701 99.5127
R16640 vdd.n2483 vdd.n701 99.5127
R16641 vdd.n2483 vdd.n693 99.5127
R16642 vdd.n2491 vdd.n693 99.5127
R16643 vdd.n2491 vdd.n691 99.5127
R16644 vdd.n2495 vdd.n691 99.5127
R16645 vdd.n2495 vdd.n680 99.5127
R16646 vdd.n2503 vdd.n680 99.5127
R16647 vdd.n2503 vdd.n678 99.5127
R16648 vdd.n2507 vdd.n678 99.5127
R16649 vdd.n2507 vdd.n669 99.5127
R16650 vdd.n2515 vdd.n669 99.5127
R16651 vdd.n2515 vdd.n667 99.5127
R16652 vdd.n2519 vdd.n667 99.5127
R16653 vdd.n2519 vdd.n657 99.5127
R16654 vdd.n2527 vdd.n657 99.5127
R16655 vdd.n2527 vdd.n655 99.5127
R16656 vdd.n2531 vdd.n655 99.5127
R16657 vdd.n2531 vdd.n646 99.5127
R16658 vdd.n2541 vdd.n646 99.5127
R16659 vdd.n2541 vdd.n644 99.5127
R16660 vdd.n2545 vdd.n644 99.5127
R16661 vdd.n2545 vdd.n632 99.5127
R16662 vdd.n2598 vdd.n632 99.5127
R16663 vdd.n2598 vdd.n630 99.5127
R16664 vdd.n2602 vdd.n630 99.5127
R16665 vdd.n2602 vdd.n598 99.5127
R16666 vdd.n2672 vdd.n598 99.5127
R16667 vdd.n2668 vdd.n599 99.5127
R16668 vdd.n2666 vdd.n2665 99.5127
R16669 vdd.n2663 vdd.n603 99.5127
R16670 vdd.n2659 vdd.n2658 99.5127
R16671 vdd.n2656 vdd.n606 99.5127
R16672 vdd.n2652 vdd.n2651 99.5127
R16673 vdd.n2649 vdd.n609 99.5127
R16674 vdd.n2645 vdd.n2644 99.5127
R16675 vdd.n2642 vdd.n2640 99.5127
R16676 vdd.n2638 vdd.n612 99.5127
R16677 vdd.n2634 vdd.n2633 99.5127
R16678 vdd.n2631 vdd.n615 99.5127
R16679 vdd.n2627 vdd.n2626 99.5127
R16680 vdd.n2624 vdd.n618 99.5127
R16681 vdd.n2620 vdd.n2619 99.5127
R16682 vdd.n2617 vdd.n621 99.5127
R16683 vdd.n2612 vdd.n2611 99.5127
R16684 vdd.n2399 vdd.n704 99.5127
R16685 vdd.n2399 vdd.n699 99.5127
R16686 vdd.n2396 vdd.n699 99.5127
R16687 vdd.n2396 vdd.n694 99.5127
R16688 vdd.n2343 vdd.n694 99.5127
R16689 vdd.n2343 vdd.n688 99.5127
R16690 vdd.n2346 vdd.n688 99.5127
R16691 vdd.n2346 vdd.n681 99.5127
R16692 vdd.n2349 vdd.n681 99.5127
R16693 vdd.n2349 vdd.n676 99.5127
R16694 vdd.n2352 vdd.n676 99.5127
R16695 vdd.n2352 vdd.n671 99.5127
R16696 vdd.n2355 vdd.n671 99.5127
R16697 vdd.n2355 vdd.n665 99.5127
R16698 vdd.n2373 vdd.n665 99.5127
R16699 vdd.n2373 vdd.n658 99.5127
R16700 vdd.n2369 vdd.n658 99.5127
R16701 vdd.n2369 vdd.n653 99.5127
R16702 vdd.n2366 vdd.n653 99.5127
R16703 vdd.n2366 vdd.n648 99.5127
R16704 vdd.n2363 vdd.n648 99.5127
R16705 vdd.n2363 vdd.n642 99.5127
R16706 vdd.n2360 vdd.n642 99.5127
R16707 vdd.n2360 vdd.n634 99.5127
R16708 vdd.n634 vdd.n627 99.5127
R16709 vdd.n2604 vdd.n627 99.5127
R16710 vdd.n2605 vdd.n2604 99.5127
R16711 vdd.n2605 vdd.n596 99.5127
R16712 vdd.n2469 vdd.n2252 99.5127
R16713 vdd.n2465 vdd.n2252 99.5127
R16714 vdd.n2463 vdd.n2462 99.5127
R16715 vdd.n2459 vdd.n2458 99.5127
R16716 vdd.n2455 vdd.n2454 99.5127
R16717 vdd.n2451 vdd.n2450 99.5127
R16718 vdd.n2447 vdd.n2446 99.5127
R16719 vdd.n2443 vdd.n2442 99.5127
R16720 vdd.n2439 vdd.n2438 99.5127
R16721 vdd.n2435 vdd.n2434 99.5127
R16722 vdd.n2431 vdd.n2430 99.5127
R16723 vdd.n2427 vdd.n2426 99.5127
R16724 vdd.n2423 vdd.n2422 99.5127
R16725 vdd.n2419 vdd.n2418 99.5127
R16726 vdd.n2415 vdd.n2414 99.5127
R16727 vdd.n2411 vdd.n2410 99.5127
R16728 vdd.n2406 vdd.n2405 99.5127
R16729 vdd.n2217 vdd.n745 99.5127
R16730 vdd.n2213 vdd.n2212 99.5127
R16731 vdd.n2209 vdd.n2208 99.5127
R16732 vdd.n2205 vdd.n2204 99.5127
R16733 vdd.n2201 vdd.n2200 99.5127
R16734 vdd.n2197 vdd.n2196 99.5127
R16735 vdd.n2193 vdd.n2192 99.5127
R16736 vdd.n2189 vdd.n2188 99.5127
R16737 vdd.n2185 vdd.n2184 99.5127
R16738 vdd.n2181 vdd.n2180 99.5127
R16739 vdd.n2177 vdd.n2176 99.5127
R16740 vdd.n2173 vdd.n2172 99.5127
R16741 vdd.n2169 vdd.n2168 99.5127
R16742 vdd.n2165 vdd.n2164 99.5127
R16743 vdd.n2161 vdd.n2160 99.5127
R16744 vdd.n2157 vdd.n2156 99.5127
R16745 vdd.n2152 vdd.n2151 99.5127
R16746 vdd.n1890 vdd.n840 99.5127
R16747 vdd.n1890 vdd.n834 99.5127
R16748 vdd.n1887 vdd.n834 99.5127
R16749 vdd.n1887 vdd.n828 99.5127
R16750 vdd.n1884 vdd.n828 99.5127
R16751 vdd.n1884 vdd.n821 99.5127
R16752 vdd.n1881 vdd.n821 99.5127
R16753 vdd.n1881 vdd.n814 99.5127
R16754 vdd.n1878 vdd.n814 99.5127
R16755 vdd.n1878 vdd.n809 99.5127
R16756 vdd.n1875 vdd.n809 99.5127
R16757 vdd.n1875 vdd.n803 99.5127
R16758 vdd.n1872 vdd.n803 99.5127
R16759 vdd.n1872 vdd.n796 99.5127
R16760 vdd.n1786 vdd.n796 99.5127
R16761 vdd.n1786 vdd.n790 99.5127
R16762 vdd.n1783 vdd.n790 99.5127
R16763 vdd.n1783 vdd.n785 99.5127
R16764 vdd.n1780 vdd.n785 99.5127
R16765 vdd.n1780 vdd.n780 99.5127
R16766 vdd.n1777 vdd.n780 99.5127
R16767 vdd.n1777 vdd.n774 99.5127
R16768 vdd.n1774 vdd.n774 99.5127
R16769 vdd.n1774 vdd.n767 99.5127
R16770 vdd.n1771 vdd.n767 99.5127
R16771 vdd.n1771 vdd.n760 99.5127
R16772 vdd.n760 vdd.n750 99.5127
R16773 vdd.n2147 vdd.n750 99.5127
R16774 vdd.n1725 vdd.n1723 99.5127
R16775 vdd.n1729 vdd.n1723 99.5127
R16776 vdd.n1733 vdd.n1731 99.5127
R16777 vdd.n1737 vdd.n1721 99.5127
R16778 vdd.n1741 vdd.n1739 99.5127
R16779 vdd.n1745 vdd.n1719 99.5127
R16780 vdd.n1749 vdd.n1747 99.5127
R16781 vdd.n1753 vdd.n1717 99.5127
R16782 vdd.n1756 vdd.n1755 99.5127
R16783 vdd.n1926 vdd.n1924 99.5127
R16784 vdd.n1922 vdd.n1758 99.5127
R16785 vdd.n1918 vdd.n1916 99.5127
R16786 vdd.n1914 vdd.n1760 99.5127
R16787 vdd.n1910 vdd.n1908 99.5127
R16788 vdd.n1906 vdd.n1762 99.5127
R16789 vdd.n1902 vdd.n1900 99.5127
R16790 vdd.n1898 vdd.n1764 99.5127
R16791 vdd.n1990 vdd.n836 99.5127
R16792 vdd.n1994 vdd.n836 99.5127
R16793 vdd.n1994 vdd.n826 99.5127
R16794 vdd.n2002 vdd.n826 99.5127
R16795 vdd.n2002 vdd.n824 99.5127
R16796 vdd.n2006 vdd.n824 99.5127
R16797 vdd.n2006 vdd.n813 99.5127
R16798 vdd.n2015 vdd.n813 99.5127
R16799 vdd.n2015 vdd.n811 99.5127
R16800 vdd.n2019 vdd.n811 99.5127
R16801 vdd.n2019 vdd.n801 99.5127
R16802 vdd.n2027 vdd.n801 99.5127
R16803 vdd.n2027 vdd.n799 99.5127
R16804 vdd.n2031 vdd.n799 99.5127
R16805 vdd.n2031 vdd.n789 99.5127
R16806 vdd.n2039 vdd.n789 99.5127
R16807 vdd.n2039 vdd.n787 99.5127
R16808 vdd.n2043 vdd.n787 99.5127
R16809 vdd.n2043 vdd.n778 99.5127
R16810 vdd.n2051 vdd.n778 99.5127
R16811 vdd.n2051 vdd.n776 99.5127
R16812 vdd.n2055 vdd.n776 99.5127
R16813 vdd.n2055 vdd.n765 99.5127
R16814 vdd.n2065 vdd.n765 99.5127
R16815 vdd.n2065 vdd.n762 99.5127
R16816 vdd.n2070 vdd.n762 99.5127
R16817 vdd.n2070 vdd.n763 99.5127
R16818 vdd.n763 vdd.n744 99.5127
R16819 vdd.n2588 vdd.n2587 99.5127
R16820 vdd.n2585 vdd.n2551 99.5127
R16821 vdd.n2581 vdd.n2580 99.5127
R16822 vdd.n2578 vdd.n2554 99.5127
R16823 vdd.n2574 vdd.n2573 99.5127
R16824 vdd.n2571 vdd.n2557 99.5127
R16825 vdd.n2567 vdd.n2566 99.5127
R16826 vdd.n2564 vdd.n2561 99.5127
R16827 vdd.n2705 vdd.n577 99.5127
R16828 vdd.n2703 vdd.n2702 99.5127
R16829 vdd.n2700 vdd.n579 99.5127
R16830 vdd.n2696 vdd.n2695 99.5127
R16831 vdd.n2693 vdd.n582 99.5127
R16832 vdd.n2689 vdd.n2688 99.5127
R16833 vdd.n2686 vdd.n585 99.5127
R16834 vdd.n2682 vdd.n2681 99.5127
R16835 vdd.n2679 vdd.n588 99.5127
R16836 vdd.n2323 vdd.n705 99.5127
R16837 vdd.n2323 vdd.n700 99.5127
R16838 vdd.n2394 vdd.n700 99.5127
R16839 vdd.n2394 vdd.n695 99.5127
R16840 vdd.n2390 vdd.n695 99.5127
R16841 vdd.n2390 vdd.n689 99.5127
R16842 vdd.n2387 vdd.n689 99.5127
R16843 vdd.n2387 vdd.n682 99.5127
R16844 vdd.n2384 vdd.n682 99.5127
R16845 vdd.n2384 vdd.n677 99.5127
R16846 vdd.n2381 vdd.n677 99.5127
R16847 vdd.n2381 vdd.n672 99.5127
R16848 vdd.n2378 vdd.n672 99.5127
R16849 vdd.n2378 vdd.n666 99.5127
R16850 vdd.n2375 vdd.n666 99.5127
R16851 vdd.n2375 vdd.n659 99.5127
R16852 vdd.n2340 vdd.n659 99.5127
R16853 vdd.n2340 vdd.n654 99.5127
R16854 vdd.n2337 vdd.n654 99.5127
R16855 vdd.n2337 vdd.n649 99.5127
R16856 vdd.n2334 vdd.n649 99.5127
R16857 vdd.n2334 vdd.n643 99.5127
R16858 vdd.n2331 vdd.n643 99.5127
R16859 vdd.n2331 vdd.n635 99.5127
R16860 vdd.n2328 vdd.n635 99.5127
R16861 vdd.n2328 vdd.n628 99.5127
R16862 vdd.n628 vdd.n594 99.5127
R16863 vdd.n2674 vdd.n594 99.5127
R16864 vdd.n2473 vdd.n708 99.5127
R16865 vdd.n2261 vdd.n2260 99.5127
R16866 vdd.n2265 vdd.n2264 99.5127
R16867 vdd.n2269 vdd.n2268 99.5127
R16868 vdd.n2273 vdd.n2272 99.5127
R16869 vdd.n2277 vdd.n2276 99.5127
R16870 vdd.n2281 vdd.n2280 99.5127
R16871 vdd.n2285 vdd.n2284 99.5127
R16872 vdd.n2289 vdd.n2288 99.5127
R16873 vdd.n2293 vdd.n2292 99.5127
R16874 vdd.n2297 vdd.n2296 99.5127
R16875 vdd.n2301 vdd.n2300 99.5127
R16876 vdd.n2305 vdd.n2304 99.5127
R16877 vdd.n2309 vdd.n2308 99.5127
R16878 vdd.n2313 vdd.n2312 99.5127
R16879 vdd.n2317 vdd.n2316 99.5127
R16880 vdd.n2319 vdd.n2251 99.5127
R16881 vdd.n2477 vdd.n698 99.5127
R16882 vdd.n2485 vdd.n698 99.5127
R16883 vdd.n2485 vdd.n696 99.5127
R16884 vdd.n2489 vdd.n696 99.5127
R16885 vdd.n2489 vdd.n686 99.5127
R16886 vdd.n2497 vdd.n686 99.5127
R16887 vdd.n2497 vdd.n684 99.5127
R16888 vdd.n2501 vdd.n684 99.5127
R16889 vdd.n2501 vdd.n675 99.5127
R16890 vdd.n2509 vdd.n675 99.5127
R16891 vdd.n2509 vdd.n673 99.5127
R16892 vdd.n2513 vdd.n673 99.5127
R16893 vdd.n2513 vdd.n663 99.5127
R16894 vdd.n2521 vdd.n663 99.5127
R16895 vdd.n2521 vdd.n661 99.5127
R16896 vdd.n2525 vdd.n661 99.5127
R16897 vdd.n2525 vdd.n652 99.5127
R16898 vdd.n2533 vdd.n652 99.5127
R16899 vdd.n2533 vdd.n650 99.5127
R16900 vdd.n2539 vdd.n650 99.5127
R16901 vdd.n2539 vdd.n640 99.5127
R16902 vdd.n2547 vdd.n640 99.5127
R16903 vdd.n2547 vdd.n637 99.5127
R16904 vdd.n2596 vdd.n637 99.5127
R16905 vdd.n2596 vdd.n638 99.5127
R16906 vdd.n638 vdd.n629 99.5127
R16907 vdd.n2591 vdd.n629 99.5127
R16908 vdd.n2591 vdd.n597 99.5127
R16909 vdd.n2141 vdd.n2140 99.5127
R16910 vdd.n2137 vdd.n2136 99.5127
R16911 vdd.n2133 vdd.n2132 99.5127
R16912 vdd.n2129 vdd.n2128 99.5127
R16913 vdd.n2125 vdd.n2124 99.5127
R16914 vdd.n2121 vdd.n2120 99.5127
R16915 vdd.n2117 vdd.n2116 99.5127
R16916 vdd.n2113 vdd.n2112 99.5127
R16917 vdd.n2109 vdd.n2108 99.5127
R16918 vdd.n2105 vdd.n2104 99.5127
R16919 vdd.n2101 vdd.n2100 99.5127
R16920 vdd.n2097 vdd.n2096 99.5127
R16921 vdd.n2093 vdd.n2092 99.5127
R16922 vdd.n2089 vdd.n2088 99.5127
R16923 vdd.n2085 vdd.n2084 99.5127
R16924 vdd.n2081 vdd.n2080 99.5127
R16925 vdd.n2077 vdd.n726 99.5127
R16926 vdd.n1834 vdd.n841 99.5127
R16927 vdd.n1834 vdd.n835 99.5127
R16928 vdd.n1837 vdd.n835 99.5127
R16929 vdd.n1837 vdd.n829 99.5127
R16930 vdd.n1840 vdd.n829 99.5127
R16931 vdd.n1840 vdd.n822 99.5127
R16932 vdd.n1843 vdd.n822 99.5127
R16933 vdd.n1843 vdd.n815 99.5127
R16934 vdd.n1846 vdd.n815 99.5127
R16935 vdd.n1846 vdd.n810 99.5127
R16936 vdd.n1849 vdd.n810 99.5127
R16937 vdd.n1849 vdd.n804 99.5127
R16938 vdd.n1870 vdd.n804 99.5127
R16939 vdd.n1870 vdd.n797 99.5127
R16940 vdd.n1866 vdd.n797 99.5127
R16941 vdd.n1866 vdd.n791 99.5127
R16942 vdd.n1863 vdd.n791 99.5127
R16943 vdd.n1863 vdd.n786 99.5127
R16944 vdd.n1860 vdd.n786 99.5127
R16945 vdd.n1860 vdd.n781 99.5127
R16946 vdd.n1857 vdd.n781 99.5127
R16947 vdd.n1857 vdd.n775 99.5127
R16948 vdd.n1854 vdd.n775 99.5127
R16949 vdd.n1854 vdd.n768 99.5127
R16950 vdd.n768 vdd.n759 99.5127
R16951 vdd.n2072 vdd.n759 99.5127
R16952 vdd.n2073 vdd.n2072 99.5127
R16953 vdd.n2073 vdd.n751 99.5127
R16954 vdd.n1984 vdd.n1982 99.5127
R16955 vdd.n1980 vdd.n844 99.5127
R16956 vdd.n1976 vdd.n1974 99.5127
R16957 vdd.n1972 vdd.n846 99.5127
R16958 vdd.n1968 vdd.n1966 99.5127
R16959 vdd.n1964 vdd.n848 99.5127
R16960 vdd.n1960 vdd.n1958 99.5127
R16961 vdd.n1956 vdd.n850 99.5127
R16962 vdd.n1798 vdd.n852 99.5127
R16963 vdd.n1803 vdd.n1800 99.5127
R16964 vdd.n1807 vdd.n1805 99.5127
R16965 vdd.n1811 vdd.n1796 99.5127
R16966 vdd.n1815 vdd.n1813 99.5127
R16967 vdd.n1819 vdd.n1794 99.5127
R16968 vdd.n1823 vdd.n1821 99.5127
R16969 vdd.n1828 vdd.n1790 99.5127
R16970 vdd.n1831 vdd.n1830 99.5127
R16971 vdd.n1988 vdd.n832 99.5127
R16972 vdd.n1996 vdd.n832 99.5127
R16973 vdd.n1996 vdd.n830 99.5127
R16974 vdd.n2000 vdd.n830 99.5127
R16975 vdd.n2000 vdd.n819 99.5127
R16976 vdd.n2008 vdd.n819 99.5127
R16977 vdd.n2008 vdd.n816 99.5127
R16978 vdd.n2013 vdd.n816 99.5127
R16979 vdd.n2013 vdd.n807 99.5127
R16980 vdd.n2021 vdd.n807 99.5127
R16981 vdd.n2021 vdd.n805 99.5127
R16982 vdd.n2025 vdd.n805 99.5127
R16983 vdd.n2025 vdd.n795 99.5127
R16984 vdd.n2033 vdd.n795 99.5127
R16985 vdd.n2033 vdd.n793 99.5127
R16986 vdd.n2037 vdd.n793 99.5127
R16987 vdd.n2037 vdd.n784 99.5127
R16988 vdd.n2045 vdd.n784 99.5127
R16989 vdd.n2045 vdd.n782 99.5127
R16990 vdd.n2049 vdd.n782 99.5127
R16991 vdd.n2049 vdd.n772 99.5127
R16992 vdd.n2057 vdd.n772 99.5127
R16993 vdd.n2057 vdd.n769 99.5127
R16994 vdd.n2063 vdd.n769 99.5127
R16995 vdd.n2063 vdd.n770 99.5127
R16996 vdd.n770 vdd.n761 99.5127
R16997 vdd.n761 vdd.n752 99.5127
R16998 vdd.n2145 vdd.n752 99.5127
R16999 vdd.n9 vdd.n7 98.9633
R17000 vdd.n2 vdd.n0 98.9633
R17001 vdd.n9 vdd.n8 98.6055
R17002 vdd.n11 vdd.n10 98.6055
R17003 vdd.n13 vdd.n12 98.6055
R17004 vdd.n6 vdd.n5 98.6055
R17005 vdd.n4 vdd.n3 98.6055
R17006 vdd.n2 vdd.n1 98.6055
R17007 vdd.t47 vdd.n267 85.8723
R17008 vdd.t58 vdd.n220 85.8723
R17009 vdd.t43 vdd.n177 85.8723
R17010 vdd.t53 vdd.n130 85.8723
R17011 vdd.t84 vdd.n88 85.8723
R17012 vdd.t26 vdd.n41 85.8723
R17013 vdd.t82 vdd.n1082 85.8723
R17014 vdd.t68 vdd.n1129 85.8723
R17015 vdd.t74 vdd.n992 85.8723
R17016 vdd.t61 vdd.n1039 85.8723
R17017 vdd.t24 vdd.n903 85.8723
R17018 vdd.t83 vdd.n950 85.8723
R17019 vdd.n2537 vdd.n2536 78.546
R17020 vdd.n2011 vdd.n817 78.546
R17021 vdd.n254 vdd.n253 75.1835
R17022 vdd.n252 vdd.n251 75.1835
R17023 vdd.n250 vdd.n249 75.1835
R17024 vdd.n164 vdd.n163 75.1835
R17025 vdd.n162 vdd.n161 75.1835
R17026 vdd.n160 vdd.n159 75.1835
R17027 vdd.n75 vdd.n74 75.1835
R17028 vdd.n73 vdd.n72 75.1835
R17029 vdd.n71 vdd.n70 75.1835
R17030 vdd.n1112 vdd.n1111 75.1835
R17031 vdd.n1114 vdd.n1113 75.1835
R17032 vdd.n1116 vdd.n1115 75.1835
R17033 vdd.n1022 vdd.n1021 75.1835
R17034 vdd.n1024 vdd.n1023 75.1835
R17035 vdd.n1026 vdd.n1025 75.1835
R17036 vdd.n933 vdd.n932 75.1835
R17037 vdd.n935 vdd.n934 75.1835
R17038 vdd.n937 vdd.n936 75.1835
R17039 vdd.n2472 vdd.n2471 72.8958
R17040 vdd.n2471 vdd.n2235 72.8958
R17041 vdd.n2471 vdd.n2236 72.8958
R17042 vdd.n2471 vdd.n2237 72.8958
R17043 vdd.n2471 vdd.n2238 72.8958
R17044 vdd.n2471 vdd.n2239 72.8958
R17045 vdd.n2471 vdd.n2240 72.8958
R17046 vdd.n2471 vdd.n2241 72.8958
R17047 vdd.n2471 vdd.n2242 72.8958
R17048 vdd.n2471 vdd.n2243 72.8958
R17049 vdd.n2471 vdd.n2244 72.8958
R17050 vdd.n2471 vdd.n2245 72.8958
R17051 vdd.n2471 vdd.n2246 72.8958
R17052 vdd.n2471 vdd.n2247 72.8958
R17053 vdd.n2471 vdd.n2248 72.8958
R17054 vdd.n2471 vdd.n2249 72.8958
R17055 vdd.n2471 vdd.n2250 72.8958
R17056 vdd.n593 vdd.n484 72.8958
R17057 vdd.n2680 vdd.n484 72.8958
R17058 vdd.n587 vdd.n484 72.8958
R17059 vdd.n2687 vdd.n484 72.8958
R17060 vdd.n584 vdd.n484 72.8958
R17061 vdd.n2694 vdd.n484 72.8958
R17062 vdd.n581 vdd.n484 72.8958
R17063 vdd.n2701 vdd.n484 72.8958
R17064 vdd.n2704 vdd.n484 72.8958
R17065 vdd.n2560 vdd.n484 72.8958
R17066 vdd.n2565 vdd.n484 72.8958
R17067 vdd.n2559 vdd.n484 72.8958
R17068 vdd.n2572 vdd.n484 72.8958
R17069 vdd.n2556 vdd.n484 72.8958
R17070 vdd.n2579 vdd.n484 72.8958
R17071 vdd.n2553 vdd.n484 72.8958
R17072 vdd.n2586 vdd.n484 72.8958
R17073 vdd.n1724 vdd.n839 72.8958
R17074 vdd.n1730 vdd.n839 72.8958
R17075 vdd.n1732 vdd.n839 72.8958
R17076 vdd.n1738 vdd.n839 72.8958
R17077 vdd.n1740 vdd.n839 72.8958
R17078 vdd.n1746 vdd.n839 72.8958
R17079 vdd.n1748 vdd.n839 72.8958
R17080 vdd.n1754 vdd.n839 72.8958
R17081 vdd.n1925 vdd.n839 72.8958
R17082 vdd.n1923 vdd.n839 72.8958
R17083 vdd.n1917 vdd.n839 72.8958
R17084 vdd.n1915 vdd.n839 72.8958
R17085 vdd.n1909 vdd.n839 72.8958
R17086 vdd.n1907 vdd.n839 72.8958
R17087 vdd.n1901 vdd.n839 72.8958
R17088 vdd.n1899 vdd.n839 72.8958
R17089 vdd.n1893 vdd.n839 72.8958
R17090 vdd.n2218 vdd.n727 72.8958
R17091 vdd.n2218 vdd.n728 72.8958
R17092 vdd.n2218 vdd.n729 72.8958
R17093 vdd.n2218 vdd.n730 72.8958
R17094 vdd.n2218 vdd.n731 72.8958
R17095 vdd.n2218 vdd.n732 72.8958
R17096 vdd.n2218 vdd.n733 72.8958
R17097 vdd.n2218 vdd.n734 72.8958
R17098 vdd.n2218 vdd.n735 72.8958
R17099 vdd.n2218 vdd.n736 72.8958
R17100 vdd.n2218 vdd.n737 72.8958
R17101 vdd.n2218 vdd.n738 72.8958
R17102 vdd.n2218 vdd.n739 72.8958
R17103 vdd.n2218 vdd.n740 72.8958
R17104 vdd.n2218 vdd.n741 72.8958
R17105 vdd.n2218 vdd.n742 72.8958
R17106 vdd.n2218 vdd.n743 72.8958
R17107 vdd.n2471 vdd.n2470 72.8958
R17108 vdd.n2471 vdd.n2219 72.8958
R17109 vdd.n2471 vdd.n2220 72.8958
R17110 vdd.n2471 vdd.n2221 72.8958
R17111 vdd.n2471 vdd.n2222 72.8958
R17112 vdd.n2471 vdd.n2223 72.8958
R17113 vdd.n2471 vdd.n2224 72.8958
R17114 vdd.n2471 vdd.n2225 72.8958
R17115 vdd.n2471 vdd.n2226 72.8958
R17116 vdd.n2471 vdd.n2227 72.8958
R17117 vdd.n2471 vdd.n2228 72.8958
R17118 vdd.n2471 vdd.n2229 72.8958
R17119 vdd.n2471 vdd.n2230 72.8958
R17120 vdd.n2471 vdd.n2231 72.8958
R17121 vdd.n2471 vdd.n2232 72.8958
R17122 vdd.n2471 vdd.n2233 72.8958
R17123 vdd.n2471 vdd.n2234 72.8958
R17124 vdd.n2610 vdd.n484 72.8958
R17125 vdd.n625 vdd.n484 72.8958
R17126 vdd.n2618 vdd.n484 72.8958
R17127 vdd.n620 vdd.n484 72.8958
R17128 vdd.n2625 vdd.n484 72.8958
R17129 vdd.n617 vdd.n484 72.8958
R17130 vdd.n2632 vdd.n484 72.8958
R17131 vdd.n614 vdd.n484 72.8958
R17132 vdd.n2639 vdd.n484 72.8958
R17133 vdd.n2643 vdd.n484 72.8958
R17134 vdd.n611 vdd.n484 72.8958
R17135 vdd.n2650 vdd.n484 72.8958
R17136 vdd.n608 vdd.n484 72.8958
R17137 vdd.n2657 vdd.n484 72.8958
R17138 vdd.n605 vdd.n484 72.8958
R17139 vdd.n2664 vdd.n484 72.8958
R17140 vdd.n2667 vdd.n484 72.8958
R17141 vdd.n2218 vdd.n725 72.8958
R17142 vdd.n2218 vdd.n724 72.8958
R17143 vdd.n2218 vdd.n723 72.8958
R17144 vdd.n2218 vdd.n722 72.8958
R17145 vdd.n2218 vdd.n721 72.8958
R17146 vdd.n2218 vdd.n720 72.8958
R17147 vdd.n2218 vdd.n719 72.8958
R17148 vdd.n2218 vdd.n718 72.8958
R17149 vdd.n2218 vdd.n717 72.8958
R17150 vdd.n2218 vdd.n716 72.8958
R17151 vdd.n2218 vdd.n715 72.8958
R17152 vdd.n2218 vdd.n714 72.8958
R17153 vdd.n2218 vdd.n713 72.8958
R17154 vdd.n2218 vdd.n712 72.8958
R17155 vdd.n2218 vdd.n711 72.8958
R17156 vdd.n2218 vdd.n710 72.8958
R17157 vdd.n2218 vdd.n709 72.8958
R17158 vdd.n1983 vdd.n839 72.8958
R17159 vdd.n1981 vdd.n839 72.8958
R17160 vdd.n1975 vdd.n839 72.8958
R17161 vdd.n1973 vdd.n839 72.8958
R17162 vdd.n1967 vdd.n839 72.8958
R17163 vdd.n1965 vdd.n839 72.8958
R17164 vdd.n1959 vdd.n839 72.8958
R17165 vdd.n1957 vdd.n839 72.8958
R17166 vdd.n851 vdd.n839 72.8958
R17167 vdd.n1799 vdd.n839 72.8958
R17168 vdd.n1804 vdd.n839 72.8958
R17169 vdd.n1806 vdd.n839 72.8958
R17170 vdd.n1812 vdd.n839 72.8958
R17171 vdd.n1814 vdd.n839 72.8958
R17172 vdd.n1820 vdd.n839 72.8958
R17173 vdd.n1822 vdd.n839 72.8958
R17174 vdd.n1829 vdd.n839 72.8958
R17175 vdd.n1422 vdd.n1421 66.2847
R17176 vdd.n1421 vdd.n1197 66.2847
R17177 vdd.n1421 vdd.n1198 66.2847
R17178 vdd.n1421 vdd.n1199 66.2847
R17179 vdd.n1421 vdd.n1200 66.2847
R17180 vdd.n1421 vdd.n1201 66.2847
R17181 vdd.n1421 vdd.n1202 66.2847
R17182 vdd.n1421 vdd.n1203 66.2847
R17183 vdd.n1421 vdd.n1204 66.2847
R17184 vdd.n1421 vdd.n1205 66.2847
R17185 vdd.n1421 vdd.n1206 66.2847
R17186 vdd.n1421 vdd.n1207 66.2847
R17187 vdd.n1421 vdd.n1208 66.2847
R17188 vdd.n1421 vdd.n1209 66.2847
R17189 vdd.n1421 vdd.n1210 66.2847
R17190 vdd.n1421 vdd.n1211 66.2847
R17191 vdd.n1421 vdd.n1212 66.2847
R17192 vdd.n1421 vdd.n1213 66.2847
R17193 vdd.n1421 vdd.n1214 66.2847
R17194 vdd.n1421 vdd.n1215 66.2847
R17195 vdd.n1421 vdd.n1216 66.2847
R17196 vdd.n1421 vdd.n1217 66.2847
R17197 vdd.n1421 vdd.n1218 66.2847
R17198 vdd.n1421 vdd.n1219 66.2847
R17199 vdd.n1421 vdd.n1220 66.2847
R17200 vdd.n1421 vdd.n1221 66.2847
R17201 vdd.n1421 vdd.n1222 66.2847
R17202 vdd.n1421 vdd.n1223 66.2847
R17203 vdd.n1421 vdd.n1224 66.2847
R17204 vdd.n1421 vdd.n1225 66.2847
R17205 vdd.n1421 vdd.n1226 66.2847
R17206 vdd.n863 vdd.n860 66.2847
R17207 vdd.n1614 vdd.n863 66.2847
R17208 vdd.n1619 vdd.n863 66.2847
R17209 vdd.n1624 vdd.n863 66.2847
R17210 vdd.n1612 vdd.n863 66.2847
R17211 vdd.n1631 vdd.n863 66.2847
R17212 vdd.n1604 vdd.n863 66.2847
R17213 vdd.n1638 vdd.n863 66.2847
R17214 vdd.n1597 vdd.n863 66.2847
R17215 vdd.n1645 vdd.n863 66.2847
R17216 vdd.n1591 vdd.n863 66.2847
R17217 vdd.n1586 vdd.n863 66.2847
R17218 vdd.n1656 vdd.n863 66.2847
R17219 vdd.n1578 vdd.n863 66.2847
R17220 vdd.n1663 vdd.n863 66.2847
R17221 vdd.n1571 vdd.n863 66.2847
R17222 vdd.n1670 vdd.n863 66.2847
R17223 vdd.n1564 vdd.n863 66.2847
R17224 vdd.n1677 vdd.n863 66.2847
R17225 vdd.n1557 vdd.n863 66.2847
R17226 vdd.n1684 vdd.n863 66.2847
R17227 vdd.n1551 vdd.n863 66.2847
R17228 vdd.n1546 vdd.n863 66.2847
R17229 vdd.n1695 vdd.n863 66.2847
R17230 vdd.n1538 vdd.n863 66.2847
R17231 vdd.n1702 vdd.n863 66.2847
R17232 vdd.n1531 vdd.n863 66.2847
R17233 vdd.n1709 vdd.n863 66.2847
R17234 vdd.n1712 vdd.n863 66.2847
R17235 vdd.n1522 vdd.n863 66.2847
R17236 vdd.n1934 vdd.n863 66.2847
R17237 vdd.n1516 vdd.n863 66.2847
R17238 vdd.n2841 vdd.n2840 66.2847
R17239 vdd.n2840 vdd.n485 66.2847
R17240 vdd.n2840 vdd.n486 66.2847
R17241 vdd.n2840 vdd.n487 66.2847
R17242 vdd.n2840 vdd.n488 66.2847
R17243 vdd.n2840 vdd.n489 66.2847
R17244 vdd.n2840 vdd.n490 66.2847
R17245 vdd.n2840 vdd.n491 66.2847
R17246 vdd.n2840 vdd.n492 66.2847
R17247 vdd.n2840 vdd.n493 66.2847
R17248 vdd.n2840 vdd.n494 66.2847
R17249 vdd.n2840 vdd.n495 66.2847
R17250 vdd.n2840 vdd.n496 66.2847
R17251 vdd.n2840 vdd.n497 66.2847
R17252 vdd.n2840 vdd.n498 66.2847
R17253 vdd.n2840 vdd.n499 66.2847
R17254 vdd.n2840 vdd.n500 66.2847
R17255 vdd.n2840 vdd.n501 66.2847
R17256 vdd.n2840 vdd.n502 66.2847
R17257 vdd.n2840 vdd.n503 66.2847
R17258 vdd.n2840 vdd.n504 66.2847
R17259 vdd.n2840 vdd.n505 66.2847
R17260 vdd.n2840 vdd.n506 66.2847
R17261 vdd.n2840 vdd.n507 66.2847
R17262 vdd.n2840 vdd.n508 66.2847
R17263 vdd.n2840 vdd.n509 66.2847
R17264 vdd.n2840 vdd.n510 66.2847
R17265 vdd.n2840 vdd.n511 66.2847
R17266 vdd.n2840 vdd.n512 66.2847
R17267 vdd.n2840 vdd.n513 66.2847
R17268 vdd.n2840 vdd.n514 66.2847
R17269 vdd.n2905 vdd.n329 66.2847
R17270 vdd.n2914 vdd.n329 66.2847
R17271 vdd.n439 vdd.n329 66.2847
R17272 vdd.n2921 vdd.n329 66.2847
R17273 vdd.n432 vdd.n329 66.2847
R17274 vdd.n2928 vdd.n329 66.2847
R17275 vdd.n425 vdd.n329 66.2847
R17276 vdd.n2935 vdd.n329 66.2847
R17277 vdd.n418 vdd.n329 66.2847
R17278 vdd.n2942 vdd.n329 66.2847
R17279 vdd.n412 vdd.n329 66.2847
R17280 vdd.n407 vdd.n329 66.2847
R17281 vdd.n2953 vdd.n329 66.2847
R17282 vdd.n399 vdd.n329 66.2847
R17283 vdd.n2960 vdd.n329 66.2847
R17284 vdd.n392 vdd.n329 66.2847
R17285 vdd.n2967 vdd.n329 66.2847
R17286 vdd.n385 vdd.n329 66.2847
R17287 vdd.n2974 vdd.n329 66.2847
R17288 vdd.n378 vdd.n329 66.2847
R17289 vdd.n2981 vdd.n329 66.2847
R17290 vdd.n372 vdd.n329 66.2847
R17291 vdd.n367 vdd.n329 66.2847
R17292 vdd.n2992 vdd.n329 66.2847
R17293 vdd.n359 vdd.n329 66.2847
R17294 vdd.n2999 vdd.n329 66.2847
R17295 vdd.n352 vdd.n329 66.2847
R17296 vdd.n3006 vdd.n329 66.2847
R17297 vdd.n345 vdd.n329 66.2847
R17298 vdd.n3013 vdd.n329 66.2847
R17299 vdd.n3016 vdd.n329 66.2847
R17300 vdd.n333 vdd.n329 66.2847
R17301 vdd.n334 vdd.n333 52.4337
R17302 vdd.n3016 vdd.n3015 52.4337
R17303 vdd.n3013 vdd.n3012 52.4337
R17304 vdd.n3008 vdd.n345 52.4337
R17305 vdd.n3006 vdd.n3005 52.4337
R17306 vdd.n3001 vdd.n352 52.4337
R17307 vdd.n2999 vdd.n2998 52.4337
R17308 vdd.n2994 vdd.n359 52.4337
R17309 vdd.n2992 vdd.n2991 52.4337
R17310 vdd.n368 vdd.n367 52.4337
R17311 vdd.n2983 vdd.n372 52.4337
R17312 vdd.n2981 vdd.n2980 52.4337
R17313 vdd.n2976 vdd.n378 52.4337
R17314 vdd.n2974 vdd.n2973 52.4337
R17315 vdd.n2969 vdd.n385 52.4337
R17316 vdd.n2967 vdd.n2966 52.4337
R17317 vdd.n2962 vdd.n392 52.4337
R17318 vdd.n2960 vdd.n2959 52.4337
R17319 vdd.n2955 vdd.n399 52.4337
R17320 vdd.n2953 vdd.n2952 52.4337
R17321 vdd.n408 vdd.n407 52.4337
R17322 vdd.n2944 vdd.n412 52.4337
R17323 vdd.n2942 vdd.n2941 52.4337
R17324 vdd.n2937 vdd.n418 52.4337
R17325 vdd.n2935 vdd.n2934 52.4337
R17326 vdd.n2930 vdd.n425 52.4337
R17327 vdd.n2928 vdd.n2927 52.4337
R17328 vdd.n2923 vdd.n432 52.4337
R17329 vdd.n2921 vdd.n2920 52.4337
R17330 vdd.n2916 vdd.n439 52.4337
R17331 vdd.n2914 vdd.n2913 52.4337
R17332 vdd.n2906 vdd.n2905 52.4337
R17333 vdd.n2842 vdd.n2841 52.4337
R17334 vdd.n517 vdd.n485 52.4337
R17335 vdd.n523 vdd.n486 52.4337
R17336 vdd.n2831 vdd.n487 52.4337
R17337 vdd.n2827 vdd.n488 52.4337
R17338 vdd.n2823 vdd.n489 52.4337
R17339 vdd.n2819 vdd.n490 52.4337
R17340 vdd.n2815 vdd.n491 52.4337
R17341 vdd.n2811 vdd.n492 52.4337
R17342 vdd.n2807 vdd.n493 52.4337
R17343 vdd.n2799 vdd.n494 52.4337
R17344 vdd.n2795 vdd.n495 52.4337
R17345 vdd.n2791 vdd.n496 52.4337
R17346 vdd.n2787 vdd.n497 52.4337
R17347 vdd.n2783 vdd.n498 52.4337
R17348 vdd.n2779 vdd.n499 52.4337
R17349 vdd.n2775 vdd.n500 52.4337
R17350 vdd.n2771 vdd.n501 52.4337
R17351 vdd.n2767 vdd.n502 52.4337
R17352 vdd.n2763 vdd.n503 52.4337
R17353 vdd.n2759 vdd.n504 52.4337
R17354 vdd.n2753 vdd.n505 52.4337
R17355 vdd.n2749 vdd.n506 52.4337
R17356 vdd.n2745 vdd.n507 52.4337
R17357 vdd.n2741 vdd.n508 52.4337
R17358 vdd.n2737 vdd.n509 52.4337
R17359 vdd.n2733 vdd.n510 52.4337
R17360 vdd.n2729 vdd.n511 52.4337
R17361 vdd.n2725 vdd.n512 52.4337
R17362 vdd.n2721 vdd.n513 52.4337
R17363 vdd.n2717 vdd.n514 52.4337
R17364 vdd.n1936 vdd.n1516 52.4337
R17365 vdd.n1934 vdd.n1933 52.4337
R17366 vdd.n1523 vdd.n1522 52.4337
R17367 vdd.n1712 vdd.n1711 52.4337
R17368 vdd.n1709 vdd.n1708 52.4337
R17369 vdd.n1704 vdd.n1531 52.4337
R17370 vdd.n1702 vdd.n1701 52.4337
R17371 vdd.n1697 vdd.n1538 52.4337
R17372 vdd.n1695 vdd.n1694 52.4337
R17373 vdd.n1547 vdd.n1546 52.4337
R17374 vdd.n1686 vdd.n1551 52.4337
R17375 vdd.n1684 vdd.n1683 52.4337
R17376 vdd.n1679 vdd.n1557 52.4337
R17377 vdd.n1677 vdd.n1676 52.4337
R17378 vdd.n1672 vdd.n1564 52.4337
R17379 vdd.n1670 vdd.n1669 52.4337
R17380 vdd.n1665 vdd.n1571 52.4337
R17381 vdd.n1663 vdd.n1662 52.4337
R17382 vdd.n1658 vdd.n1578 52.4337
R17383 vdd.n1656 vdd.n1655 52.4337
R17384 vdd.n1587 vdd.n1586 52.4337
R17385 vdd.n1647 vdd.n1591 52.4337
R17386 vdd.n1645 vdd.n1644 52.4337
R17387 vdd.n1640 vdd.n1597 52.4337
R17388 vdd.n1638 vdd.n1637 52.4337
R17389 vdd.n1633 vdd.n1604 52.4337
R17390 vdd.n1631 vdd.n1630 52.4337
R17391 vdd.n1626 vdd.n1612 52.4337
R17392 vdd.n1624 vdd.n1623 52.4337
R17393 vdd.n1619 vdd.n1618 52.4337
R17394 vdd.n1614 vdd.n1613 52.4337
R17395 vdd.n1945 vdd.n860 52.4337
R17396 vdd.n1423 vdd.n1422 52.4337
R17397 vdd.n1229 vdd.n1197 52.4337
R17398 vdd.n1233 vdd.n1198 52.4337
R17399 vdd.n1235 vdd.n1199 52.4337
R17400 vdd.n1239 vdd.n1200 52.4337
R17401 vdd.n1241 vdd.n1201 52.4337
R17402 vdd.n1245 vdd.n1202 52.4337
R17403 vdd.n1247 vdd.n1203 52.4337
R17404 vdd.n1251 vdd.n1204 52.4337
R17405 vdd.n1253 vdd.n1205 52.4337
R17406 vdd.n1259 vdd.n1206 52.4337
R17407 vdd.n1261 vdd.n1207 52.4337
R17408 vdd.n1265 vdd.n1208 52.4337
R17409 vdd.n1267 vdd.n1209 52.4337
R17410 vdd.n1271 vdd.n1210 52.4337
R17411 vdd.n1273 vdd.n1211 52.4337
R17412 vdd.n1277 vdd.n1212 52.4337
R17413 vdd.n1279 vdd.n1213 52.4337
R17414 vdd.n1283 vdd.n1214 52.4337
R17415 vdd.n1285 vdd.n1215 52.4337
R17416 vdd.n1357 vdd.n1216 52.4337
R17417 vdd.n1290 vdd.n1217 52.4337
R17418 vdd.n1294 vdd.n1218 52.4337
R17419 vdd.n1296 vdd.n1219 52.4337
R17420 vdd.n1300 vdd.n1220 52.4337
R17421 vdd.n1302 vdd.n1221 52.4337
R17422 vdd.n1306 vdd.n1222 52.4337
R17423 vdd.n1308 vdd.n1223 52.4337
R17424 vdd.n1312 vdd.n1224 52.4337
R17425 vdd.n1314 vdd.n1225 52.4337
R17426 vdd.n1318 vdd.n1226 52.4337
R17427 vdd.n1422 vdd.n1196 52.4337
R17428 vdd.n1232 vdd.n1197 52.4337
R17429 vdd.n1234 vdd.n1198 52.4337
R17430 vdd.n1238 vdd.n1199 52.4337
R17431 vdd.n1240 vdd.n1200 52.4337
R17432 vdd.n1244 vdd.n1201 52.4337
R17433 vdd.n1246 vdd.n1202 52.4337
R17434 vdd.n1250 vdd.n1203 52.4337
R17435 vdd.n1252 vdd.n1204 52.4337
R17436 vdd.n1258 vdd.n1205 52.4337
R17437 vdd.n1260 vdd.n1206 52.4337
R17438 vdd.n1264 vdd.n1207 52.4337
R17439 vdd.n1266 vdd.n1208 52.4337
R17440 vdd.n1270 vdd.n1209 52.4337
R17441 vdd.n1272 vdd.n1210 52.4337
R17442 vdd.n1276 vdd.n1211 52.4337
R17443 vdd.n1278 vdd.n1212 52.4337
R17444 vdd.n1282 vdd.n1213 52.4337
R17445 vdd.n1284 vdd.n1214 52.4337
R17446 vdd.n1288 vdd.n1215 52.4337
R17447 vdd.n1289 vdd.n1216 52.4337
R17448 vdd.n1293 vdd.n1217 52.4337
R17449 vdd.n1295 vdd.n1218 52.4337
R17450 vdd.n1299 vdd.n1219 52.4337
R17451 vdd.n1301 vdd.n1220 52.4337
R17452 vdd.n1305 vdd.n1221 52.4337
R17453 vdd.n1307 vdd.n1222 52.4337
R17454 vdd.n1311 vdd.n1223 52.4337
R17455 vdd.n1313 vdd.n1224 52.4337
R17456 vdd.n1317 vdd.n1225 52.4337
R17457 vdd.n1319 vdd.n1226 52.4337
R17458 vdd.n860 vdd.n859 52.4337
R17459 vdd.n1615 vdd.n1614 52.4337
R17460 vdd.n1620 vdd.n1619 52.4337
R17461 vdd.n1625 vdd.n1624 52.4337
R17462 vdd.n1612 vdd.n1605 52.4337
R17463 vdd.n1632 vdd.n1631 52.4337
R17464 vdd.n1604 vdd.n1598 52.4337
R17465 vdd.n1639 vdd.n1638 52.4337
R17466 vdd.n1597 vdd.n1592 52.4337
R17467 vdd.n1646 vdd.n1645 52.4337
R17468 vdd.n1591 vdd.n1590 52.4337
R17469 vdd.n1586 vdd.n1579 52.4337
R17470 vdd.n1657 vdd.n1656 52.4337
R17471 vdd.n1578 vdd.n1572 52.4337
R17472 vdd.n1664 vdd.n1663 52.4337
R17473 vdd.n1571 vdd.n1565 52.4337
R17474 vdd.n1671 vdd.n1670 52.4337
R17475 vdd.n1564 vdd.n1558 52.4337
R17476 vdd.n1678 vdd.n1677 52.4337
R17477 vdd.n1557 vdd.n1552 52.4337
R17478 vdd.n1685 vdd.n1684 52.4337
R17479 vdd.n1551 vdd.n1550 52.4337
R17480 vdd.n1546 vdd.n1539 52.4337
R17481 vdd.n1696 vdd.n1695 52.4337
R17482 vdd.n1538 vdd.n1532 52.4337
R17483 vdd.n1703 vdd.n1702 52.4337
R17484 vdd.n1531 vdd.n1525 52.4337
R17485 vdd.n1710 vdd.n1709 52.4337
R17486 vdd.n1713 vdd.n1712 52.4337
R17487 vdd.n1522 vdd.n1517 52.4337
R17488 vdd.n1935 vdd.n1934 52.4337
R17489 vdd.n1516 vdd.n865 52.4337
R17490 vdd.n2841 vdd.n483 52.4337
R17491 vdd.n522 vdd.n485 52.4337
R17492 vdd.n2832 vdd.n486 52.4337
R17493 vdd.n2828 vdd.n487 52.4337
R17494 vdd.n2824 vdd.n488 52.4337
R17495 vdd.n2820 vdd.n489 52.4337
R17496 vdd.n2816 vdd.n490 52.4337
R17497 vdd.n2812 vdd.n491 52.4337
R17498 vdd.n2808 vdd.n492 52.4337
R17499 vdd.n2798 vdd.n493 52.4337
R17500 vdd.n2796 vdd.n494 52.4337
R17501 vdd.n2792 vdd.n495 52.4337
R17502 vdd.n2788 vdd.n496 52.4337
R17503 vdd.n2784 vdd.n497 52.4337
R17504 vdd.n2780 vdd.n498 52.4337
R17505 vdd.n2776 vdd.n499 52.4337
R17506 vdd.n2772 vdd.n500 52.4337
R17507 vdd.n2768 vdd.n501 52.4337
R17508 vdd.n2764 vdd.n502 52.4337
R17509 vdd.n2760 vdd.n503 52.4337
R17510 vdd.n2752 vdd.n504 52.4337
R17511 vdd.n2750 vdd.n505 52.4337
R17512 vdd.n2746 vdd.n506 52.4337
R17513 vdd.n2742 vdd.n507 52.4337
R17514 vdd.n2738 vdd.n508 52.4337
R17515 vdd.n2734 vdd.n509 52.4337
R17516 vdd.n2730 vdd.n510 52.4337
R17517 vdd.n2726 vdd.n511 52.4337
R17518 vdd.n2722 vdd.n512 52.4337
R17519 vdd.n2718 vdd.n513 52.4337
R17520 vdd.n2714 vdd.n514 52.4337
R17521 vdd.n2905 vdd.n440 52.4337
R17522 vdd.n2915 vdd.n2914 52.4337
R17523 vdd.n439 vdd.n433 52.4337
R17524 vdd.n2922 vdd.n2921 52.4337
R17525 vdd.n432 vdd.n426 52.4337
R17526 vdd.n2929 vdd.n2928 52.4337
R17527 vdd.n425 vdd.n419 52.4337
R17528 vdd.n2936 vdd.n2935 52.4337
R17529 vdd.n418 vdd.n413 52.4337
R17530 vdd.n2943 vdd.n2942 52.4337
R17531 vdd.n412 vdd.n411 52.4337
R17532 vdd.n407 vdd.n400 52.4337
R17533 vdd.n2954 vdd.n2953 52.4337
R17534 vdd.n399 vdd.n393 52.4337
R17535 vdd.n2961 vdd.n2960 52.4337
R17536 vdd.n392 vdd.n386 52.4337
R17537 vdd.n2968 vdd.n2967 52.4337
R17538 vdd.n385 vdd.n379 52.4337
R17539 vdd.n2975 vdd.n2974 52.4337
R17540 vdd.n378 vdd.n373 52.4337
R17541 vdd.n2982 vdd.n2981 52.4337
R17542 vdd.n372 vdd.n371 52.4337
R17543 vdd.n367 vdd.n360 52.4337
R17544 vdd.n2993 vdd.n2992 52.4337
R17545 vdd.n359 vdd.n353 52.4337
R17546 vdd.n3000 vdd.n2999 52.4337
R17547 vdd.n352 vdd.n346 52.4337
R17548 vdd.n3007 vdd.n3006 52.4337
R17549 vdd.n345 vdd.n338 52.4337
R17550 vdd.n3014 vdd.n3013 52.4337
R17551 vdd.n3017 vdd.n3016 52.4337
R17552 vdd.n333 vdd.n330 52.4337
R17553 vdd.t118 vdd.t111 51.4683
R17554 vdd.n250 vdd.n248 42.0461
R17555 vdd.n160 vdd.n158 42.0461
R17556 vdd.n71 vdd.n69 42.0461
R17557 vdd.n1112 vdd.n1110 42.0461
R17558 vdd.n1022 vdd.n1020 42.0461
R17559 vdd.n933 vdd.n931 42.0461
R17560 vdd.n296 vdd.n295 41.6884
R17561 vdd.n206 vdd.n205 41.6884
R17562 vdd.n117 vdd.n116 41.6884
R17563 vdd.n1158 vdd.n1157 41.6884
R17564 vdd.n1068 vdd.n1067 41.6884
R17565 vdd.n979 vdd.n978 41.6884
R17566 vdd.n1322 vdd.n1321 41.1157
R17567 vdd.n1360 vdd.n1359 41.1157
R17568 vdd.n1256 vdd.n1255 41.1157
R17569 vdd.n2910 vdd.n2909 41.1157
R17570 vdd.n2949 vdd.n406 41.1157
R17571 vdd.n2988 vdd.n366 41.1157
R17572 vdd.n2667 vdd.n2666 39.2114
R17573 vdd.n2664 vdd.n2663 39.2114
R17574 vdd.n2659 vdd.n605 39.2114
R17575 vdd.n2657 vdd.n2656 39.2114
R17576 vdd.n2652 vdd.n608 39.2114
R17577 vdd.n2650 vdd.n2649 39.2114
R17578 vdd.n2645 vdd.n611 39.2114
R17579 vdd.n2643 vdd.n2642 39.2114
R17580 vdd.n2639 vdd.n2638 39.2114
R17581 vdd.n2634 vdd.n614 39.2114
R17582 vdd.n2632 vdd.n2631 39.2114
R17583 vdd.n2627 vdd.n617 39.2114
R17584 vdd.n2625 vdd.n2624 39.2114
R17585 vdd.n2620 vdd.n620 39.2114
R17586 vdd.n2618 vdd.n2617 39.2114
R17587 vdd.n2612 vdd.n625 39.2114
R17588 vdd.n2610 vdd.n2609 39.2114
R17589 vdd.n2470 vdd.n703 39.2114
R17590 vdd.n2465 vdd.n2219 39.2114
R17591 vdd.n2462 vdd.n2220 39.2114
R17592 vdd.n2458 vdd.n2221 39.2114
R17593 vdd.n2454 vdd.n2222 39.2114
R17594 vdd.n2450 vdd.n2223 39.2114
R17595 vdd.n2446 vdd.n2224 39.2114
R17596 vdd.n2442 vdd.n2225 39.2114
R17597 vdd.n2438 vdd.n2226 39.2114
R17598 vdd.n2434 vdd.n2227 39.2114
R17599 vdd.n2430 vdd.n2228 39.2114
R17600 vdd.n2426 vdd.n2229 39.2114
R17601 vdd.n2422 vdd.n2230 39.2114
R17602 vdd.n2418 vdd.n2231 39.2114
R17603 vdd.n2414 vdd.n2232 39.2114
R17604 vdd.n2410 vdd.n2233 39.2114
R17605 vdd.n2405 vdd.n2234 39.2114
R17606 vdd.n2213 vdd.n743 39.2114
R17607 vdd.n2209 vdd.n742 39.2114
R17608 vdd.n2205 vdd.n741 39.2114
R17609 vdd.n2201 vdd.n740 39.2114
R17610 vdd.n2197 vdd.n739 39.2114
R17611 vdd.n2193 vdd.n738 39.2114
R17612 vdd.n2189 vdd.n737 39.2114
R17613 vdd.n2185 vdd.n736 39.2114
R17614 vdd.n2181 vdd.n735 39.2114
R17615 vdd.n2177 vdd.n734 39.2114
R17616 vdd.n2173 vdd.n733 39.2114
R17617 vdd.n2169 vdd.n732 39.2114
R17618 vdd.n2165 vdd.n731 39.2114
R17619 vdd.n2161 vdd.n730 39.2114
R17620 vdd.n2157 vdd.n729 39.2114
R17621 vdd.n2152 vdd.n728 39.2114
R17622 vdd.n2148 vdd.n727 39.2114
R17623 vdd.n1724 vdd.n838 39.2114
R17624 vdd.n1730 vdd.n1729 39.2114
R17625 vdd.n1733 vdd.n1732 39.2114
R17626 vdd.n1738 vdd.n1737 39.2114
R17627 vdd.n1741 vdd.n1740 39.2114
R17628 vdd.n1746 vdd.n1745 39.2114
R17629 vdd.n1749 vdd.n1748 39.2114
R17630 vdd.n1754 vdd.n1753 39.2114
R17631 vdd.n1925 vdd.n1756 39.2114
R17632 vdd.n1924 vdd.n1923 39.2114
R17633 vdd.n1917 vdd.n1758 39.2114
R17634 vdd.n1916 vdd.n1915 39.2114
R17635 vdd.n1909 vdd.n1760 39.2114
R17636 vdd.n1908 vdd.n1907 39.2114
R17637 vdd.n1901 vdd.n1762 39.2114
R17638 vdd.n1900 vdd.n1899 39.2114
R17639 vdd.n1893 vdd.n1764 39.2114
R17640 vdd.n2586 vdd.n2585 39.2114
R17641 vdd.n2581 vdd.n2553 39.2114
R17642 vdd.n2579 vdd.n2578 39.2114
R17643 vdd.n2574 vdd.n2556 39.2114
R17644 vdd.n2572 vdd.n2571 39.2114
R17645 vdd.n2567 vdd.n2559 39.2114
R17646 vdd.n2565 vdd.n2564 39.2114
R17647 vdd.n2560 vdd.n577 39.2114
R17648 vdd.n2704 vdd.n2703 39.2114
R17649 vdd.n2701 vdd.n2700 39.2114
R17650 vdd.n2696 vdd.n581 39.2114
R17651 vdd.n2694 vdd.n2693 39.2114
R17652 vdd.n2689 vdd.n584 39.2114
R17653 vdd.n2687 vdd.n2686 39.2114
R17654 vdd.n2682 vdd.n587 39.2114
R17655 vdd.n2680 vdd.n2679 39.2114
R17656 vdd.n2675 vdd.n593 39.2114
R17657 vdd.n2472 vdd.n706 39.2114
R17658 vdd.n2235 vdd.n708 39.2114
R17659 vdd.n2261 vdd.n2236 39.2114
R17660 vdd.n2265 vdd.n2237 39.2114
R17661 vdd.n2269 vdd.n2238 39.2114
R17662 vdd.n2273 vdd.n2239 39.2114
R17663 vdd.n2277 vdd.n2240 39.2114
R17664 vdd.n2281 vdd.n2241 39.2114
R17665 vdd.n2285 vdd.n2242 39.2114
R17666 vdd.n2289 vdd.n2243 39.2114
R17667 vdd.n2293 vdd.n2244 39.2114
R17668 vdd.n2297 vdd.n2245 39.2114
R17669 vdd.n2301 vdd.n2246 39.2114
R17670 vdd.n2305 vdd.n2247 39.2114
R17671 vdd.n2309 vdd.n2248 39.2114
R17672 vdd.n2313 vdd.n2249 39.2114
R17673 vdd.n2317 vdd.n2250 39.2114
R17674 vdd.n2473 vdd.n2472 39.2114
R17675 vdd.n2260 vdd.n2235 39.2114
R17676 vdd.n2264 vdd.n2236 39.2114
R17677 vdd.n2268 vdd.n2237 39.2114
R17678 vdd.n2272 vdd.n2238 39.2114
R17679 vdd.n2276 vdd.n2239 39.2114
R17680 vdd.n2280 vdd.n2240 39.2114
R17681 vdd.n2284 vdd.n2241 39.2114
R17682 vdd.n2288 vdd.n2242 39.2114
R17683 vdd.n2292 vdd.n2243 39.2114
R17684 vdd.n2296 vdd.n2244 39.2114
R17685 vdd.n2300 vdd.n2245 39.2114
R17686 vdd.n2304 vdd.n2246 39.2114
R17687 vdd.n2308 vdd.n2247 39.2114
R17688 vdd.n2312 vdd.n2248 39.2114
R17689 vdd.n2316 vdd.n2249 39.2114
R17690 vdd.n2319 vdd.n2250 39.2114
R17691 vdd.n593 vdd.n588 39.2114
R17692 vdd.n2681 vdd.n2680 39.2114
R17693 vdd.n587 vdd.n585 39.2114
R17694 vdd.n2688 vdd.n2687 39.2114
R17695 vdd.n584 vdd.n582 39.2114
R17696 vdd.n2695 vdd.n2694 39.2114
R17697 vdd.n581 vdd.n579 39.2114
R17698 vdd.n2702 vdd.n2701 39.2114
R17699 vdd.n2705 vdd.n2704 39.2114
R17700 vdd.n2561 vdd.n2560 39.2114
R17701 vdd.n2566 vdd.n2565 39.2114
R17702 vdd.n2559 vdd.n2557 39.2114
R17703 vdd.n2573 vdd.n2572 39.2114
R17704 vdd.n2556 vdd.n2554 39.2114
R17705 vdd.n2580 vdd.n2579 39.2114
R17706 vdd.n2553 vdd.n2551 39.2114
R17707 vdd.n2587 vdd.n2586 39.2114
R17708 vdd.n1725 vdd.n1724 39.2114
R17709 vdd.n1731 vdd.n1730 39.2114
R17710 vdd.n1732 vdd.n1721 39.2114
R17711 vdd.n1739 vdd.n1738 39.2114
R17712 vdd.n1740 vdd.n1719 39.2114
R17713 vdd.n1747 vdd.n1746 39.2114
R17714 vdd.n1748 vdd.n1717 39.2114
R17715 vdd.n1755 vdd.n1754 39.2114
R17716 vdd.n1926 vdd.n1925 39.2114
R17717 vdd.n1923 vdd.n1922 39.2114
R17718 vdd.n1918 vdd.n1917 39.2114
R17719 vdd.n1915 vdd.n1914 39.2114
R17720 vdd.n1910 vdd.n1909 39.2114
R17721 vdd.n1907 vdd.n1906 39.2114
R17722 vdd.n1902 vdd.n1901 39.2114
R17723 vdd.n1899 vdd.n1898 39.2114
R17724 vdd.n1894 vdd.n1893 39.2114
R17725 vdd.n2151 vdd.n727 39.2114
R17726 vdd.n2156 vdd.n728 39.2114
R17727 vdd.n2160 vdd.n729 39.2114
R17728 vdd.n2164 vdd.n730 39.2114
R17729 vdd.n2168 vdd.n731 39.2114
R17730 vdd.n2172 vdd.n732 39.2114
R17731 vdd.n2176 vdd.n733 39.2114
R17732 vdd.n2180 vdd.n734 39.2114
R17733 vdd.n2184 vdd.n735 39.2114
R17734 vdd.n2188 vdd.n736 39.2114
R17735 vdd.n2192 vdd.n737 39.2114
R17736 vdd.n2196 vdd.n738 39.2114
R17737 vdd.n2200 vdd.n739 39.2114
R17738 vdd.n2204 vdd.n740 39.2114
R17739 vdd.n2208 vdd.n741 39.2114
R17740 vdd.n2212 vdd.n742 39.2114
R17741 vdd.n745 vdd.n743 39.2114
R17742 vdd.n2470 vdd.n2469 39.2114
R17743 vdd.n2463 vdd.n2219 39.2114
R17744 vdd.n2459 vdd.n2220 39.2114
R17745 vdd.n2455 vdd.n2221 39.2114
R17746 vdd.n2451 vdd.n2222 39.2114
R17747 vdd.n2447 vdd.n2223 39.2114
R17748 vdd.n2443 vdd.n2224 39.2114
R17749 vdd.n2439 vdd.n2225 39.2114
R17750 vdd.n2435 vdd.n2226 39.2114
R17751 vdd.n2431 vdd.n2227 39.2114
R17752 vdd.n2427 vdd.n2228 39.2114
R17753 vdd.n2423 vdd.n2229 39.2114
R17754 vdd.n2419 vdd.n2230 39.2114
R17755 vdd.n2415 vdd.n2231 39.2114
R17756 vdd.n2411 vdd.n2232 39.2114
R17757 vdd.n2406 vdd.n2233 39.2114
R17758 vdd.n2402 vdd.n2234 39.2114
R17759 vdd.n2611 vdd.n2610 39.2114
R17760 vdd.n625 vdd.n621 39.2114
R17761 vdd.n2619 vdd.n2618 39.2114
R17762 vdd.n620 vdd.n618 39.2114
R17763 vdd.n2626 vdd.n2625 39.2114
R17764 vdd.n617 vdd.n615 39.2114
R17765 vdd.n2633 vdd.n2632 39.2114
R17766 vdd.n614 vdd.n612 39.2114
R17767 vdd.n2640 vdd.n2639 39.2114
R17768 vdd.n2644 vdd.n2643 39.2114
R17769 vdd.n611 vdd.n609 39.2114
R17770 vdd.n2651 vdd.n2650 39.2114
R17771 vdd.n608 vdd.n606 39.2114
R17772 vdd.n2658 vdd.n2657 39.2114
R17773 vdd.n605 vdd.n603 39.2114
R17774 vdd.n2665 vdd.n2664 39.2114
R17775 vdd.n2668 vdd.n2667 39.2114
R17776 vdd.n753 vdd.n709 39.2114
R17777 vdd.n2140 vdd.n710 39.2114
R17778 vdd.n2136 vdd.n711 39.2114
R17779 vdd.n2132 vdd.n712 39.2114
R17780 vdd.n2128 vdd.n713 39.2114
R17781 vdd.n2124 vdd.n714 39.2114
R17782 vdd.n2120 vdd.n715 39.2114
R17783 vdd.n2116 vdd.n716 39.2114
R17784 vdd.n2112 vdd.n717 39.2114
R17785 vdd.n2108 vdd.n718 39.2114
R17786 vdd.n2104 vdd.n719 39.2114
R17787 vdd.n2100 vdd.n720 39.2114
R17788 vdd.n2096 vdd.n721 39.2114
R17789 vdd.n2092 vdd.n722 39.2114
R17790 vdd.n2088 vdd.n723 39.2114
R17791 vdd.n2084 vdd.n724 39.2114
R17792 vdd.n2080 vdd.n725 39.2114
R17793 vdd.n1983 vdd.n842 39.2114
R17794 vdd.n1982 vdd.n1981 39.2114
R17795 vdd.n1975 vdd.n844 39.2114
R17796 vdd.n1974 vdd.n1973 39.2114
R17797 vdd.n1967 vdd.n846 39.2114
R17798 vdd.n1966 vdd.n1965 39.2114
R17799 vdd.n1959 vdd.n848 39.2114
R17800 vdd.n1958 vdd.n1957 39.2114
R17801 vdd.n851 vdd.n850 39.2114
R17802 vdd.n1799 vdd.n1798 39.2114
R17803 vdd.n1804 vdd.n1803 39.2114
R17804 vdd.n1807 vdd.n1806 39.2114
R17805 vdd.n1812 vdd.n1811 39.2114
R17806 vdd.n1815 vdd.n1814 39.2114
R17807 vdd.n1820 vdd.n1819 39.2114
R17808 vdd.n1823 vdd.n1822 39.2114
R17809 vdd.n1829 vdd.n1828 39.2114
R17810 vdd.n2077 vdd.n725 39.2114
R17811 vdd.n2081 vdd.n724 39.2114
R17812 vdd.n2085 vdd.n723 39.2114
R17813 vdd.n2089 vdd.n722 39.2114
R17814 vdd.n2093 vdd.n721 39.2114
R17815 vdd.n2097 vdd.n720 39.2114
R17816 vdd.n2101 vdd.n719 39.2114
R17817 vdd.n2105 vdd.n718 39.2114
R17818 vdd.n2109 vdd.n717 39.2114
R17819 vdd.n2113 vdd.n716 39.2114
R17820 vdd.n2117 vdd.n715 39.2114
R17821 vdd.n2121 vdd.n714 39.2114
R17822 vdd.n2125 vdd.n713 39.2114
R17823 vdd.n2129 vdd.n712 39.2114
R17824 vdd.n2133 vdd.n711 39.2114
R17825 vdd.n2137 vdd.n710 39.2114
R17826 vdd.n2141 vdd.n709 39.2114
R17827 vdd.n1984 vdd.n1983 39.2114
R17828 vdd.n1981 vdd.n1980 39.2114
R17829 vdd.n1976 vdd.n1975 39.2114
R17830 vdd.n1973 vdd.n1972 39.2114
R17831 vdd.n1968 vdd.n1967 39.2114
R17832 vdd.n1965 vdd.n1964 39.2114
R17833 vdd.n1960 vdd.n1959 39.2114
R17834 vdd.n1957 vdd.n1956 39.2114
R17835 vdd.n852 vdd.n851 39.2114
R17836 vdd.n1800 vdd.n1799 39.2114
R17837 vdd.n1805 vdd.n1804 39.2114
R17838 vdd.n1806 vdd.n1796 39.2114
R17839 vdd.n1813 vdd.n1812 39.2114
R17840 vdd.n1814 vdd.n1794 39.2114
R17841 vdd.n1821 vdd.n1820 39.2114
R17842 vdd.n1822 vdd.n1790 39.2114
R17843 vdd.n1830 vdd.n1829 39.2114
R17844 vdd.n1949 vdd.n1948 37.2369
R17845 vdd.n1652 vdd.n1585 37.2369
R17846 vdd.n1691 vdd.n1545 37.2369
R17847 vdd.n2758 vdd.n558 37.2369
R17848 vdd.n2806 vdd.n2805 37.2369
R17849 vdd.n2713 vdd.n2712 37.2369
R17850 vdd.n1991 vdd.n837 31.6883
R17851 vdd.n2216 vdd.n746 31.6883
R17852 vdd.n2149 vdd.n749 31.6883
R17853 vdd.n1895 vdd.n1892 31.6883
R17854 vdd.n2403 vdd.n2401 31.6883
R17855 vdd.n2608 vdd.n2607 31.6883
R17856 vdd.n2480 vdd.n702 31.6883
R17857 vdd.n2671 vdd.n2670 31.6883
R17858 vdd.n2590 vdd.n2589 31.6883
R17859 vdd.n2676 vdd.n592 31.6883
R17860 vdd.n2322 vdd.n2321 31.6883
R17861 vdd.n2476 vdd.n2475 31.6883
R17862 vdd.n1987 vdd.n1986 31.6883
R17863 vdd.n2144 vdd.n2143 31.6883
R17864 vdd.n2076 vdd.n2075 31.6883
R17865 vdd.n1833 vdd.n1832 31.6883
R17866 vdd.n1826 vdd.n1792 30.449
R17867 vdd.n757 vdd.n756 30.449
R17868 vdd.n1767 vdd.n1766 30.449
R17869 vdd.n2154 vdd.n748 30.449
R17870 vdd.n2258 vdd.n2257 30.449
R17871 vdd.n2614 vdd.n623 30.449
R17872 vdd.n2408 vdd.n2254 30.449
R17873 vdd.n591 vdd.n590 30.449
R17874 vdd.n1421 vdd.n1228 22.6735
R17875 vdd.n1943 vdd.n863 22.6735
R17876 vdd.n2840 vdd.n516 22.6735
R17877 vdd.n3025 vdd.n329 22.6735
R17878 vdd.n1432 vdd.n1190 19.3944
R17879 vdd.n1432 vdd.n1188 19.3944
R17880 vdd.n1436 vdd.n1188 19.3944
R17881 vdd.n1436 vdd.n1178 19.3944
R17882 vdd.n1449 vdd.n1178 19.3944
R17883 vdd.n1449 vdd.n1176 19.3944
R17884 vdd.n1453 vdd.n1176 19.3944
R17885 vdd.n1453 vdd.n1168 19.3944
R17886 vdd.n1467 vdd.n1168 19.3944
R17887 vdd.n1467 vdd.n1166 19.3944
R17888 vdd.n1471 vdd.n1166 19.3944
R17889 vdd.n1471 vdd.n885 19.3944
R17890 vdd.n1483 vdd.n885 19.3944
R17891 vdd.n1483 vdd.n883 19.3944
R17892 vdd.n1487 vdd.n883 19.3944
R17893 vdd.n1487 vdd.n875 19.3944
R17894 vdd.n1500 vdd.n875 19.3944
R17895 vdd.n1500 vdd.n872 19.3944
R17896 vdd.n1506 vdd.n872 19.3944
R17897 vdd.n1506 vdd.n873 19.3944
R17898 vdd.n873 vdd.n862 19.3944
R17899 vdd.n1356 vdd.n1291 19.3944
R17900 vdd.n1352 vdd.n1291 19.3944
R17901 vdd.n1352 vdd.n1351 19.3944
R17902 vdd.n1351 vdd.n1350 19.3944
R17903 vdd.n1350 vdd.n1297 19.3944
R17904 vdd.n1346 vdd.n1297 19.3944
R17905 vdd.n1346 vdd.n1345 19.3944
R17906 vdd.n1345 vdd.n1344 19.3944
R17907 vdd.n1344 vdd.n1303 19.3944
R17908 vdd.n1340 vdd.n1303 19.3944
R17909 vdd.n1340 vdd.n1339 19.3944
R17910 vdd.n1339 vdd.n1338 19.3944
R17911 vdd.n1338 vdd.n1309 19.3944
R17912 vdd.n1334 vdd.n1309 19.3944
R17913 vdd.n1334 vdd.n1333 19.3944
R17914 vdd.n1333 vdd.n1332 19.3944
R17915 vdd.n1332 vdd.n1315 19.3944
R17916 vdd.n1328 vdd.n1315 19.3944
R17917 vdd.n1328 vdd.n1327 19.3944
R17918 vdd.n1327 vdd.n1326 19.3944
R17919 vdd.n1391 vdd.n1390 19.3944
R17920 vdd.n1390 vdd.n1389 19.3944
R17921 vdd.n1389 vdd.n1262 19.3944
R17922 vdd.n1385 vdd.n1262 19.3944
R17923 vdd.n1385 vdd.n1384 19.3944
R17924 vdd.n1384 vdd.n1383 19.3944
R17925 vdd.n1383 vdd.n1268 19.3944
R17926 vdd.n1379 vdd.n1268 19.3944
R17927 vdd.n1379 vdd.n1378 19.3944
R17928 vdd.n1378 vdd.n1377 19.3944
R17929 vdd.n1377 vdd.n1274 19.3944
R17930 vdd.n1373 vdd.n1274 19.3944
R17931 vdd.n1373 vdd.n1372 19.3944
R17932 vdd.n1372 vdd.n1371 19.3944
R17933 vdd.n1371 vdd.n1280 19.3944
R17934 vdd.n1367 vdd.n1280 19.3944
R17935 vdd.n1367 vdd.n1366 19.3944
R17936 vdd.n1366 vdd.n1365 19.3944
R17937 vdd.n1365 vdd.n1286 19.3944
R17938 vdd.n1361 vdd.n1286 19.3944
R17939 vdd.n1424 vdd.n1195 19.3944
R17940 vdd.n1419 vdd.n1195 19.3944
R17941 vdd.n1419 vdd.n1230 19.3944
R17942 vdd.n1415 vdd.n1230 19.3944
R17943 vdd.n1415 vdd.n1414 19.3944
R17944 vdd.n1414 vdd.n1413 19.3944
R17945 vdd.n1413 vdd.n1236 19.3944
R17946 vdd.n1409 vdd.n1236 19.3944
R17947 vdd.n1409 vdd.n1408 19.3944
R17948 vdd.n1408 vdd.n1407 19.3944
R17949 vdd.n1407 vdd.n1242 19.3944
R17950 vdd.n1403 vdd.n1242 19.3944
R17951 vdd.n1403 vdd.n1402 19.3944
R17952 vdd.n1402 vdd.n1401 19.3944
R17953 vdd.n1401 vdd.n1248 19.3944
R17954 vdd.n1397 vdd.n1248 19.3944
R17955 vdd.n1397 vdd.n1396 19.3944
R17956 vdd.n1396 vdd.n1395 19.3944
R17957 vdd.n1648 vdd.n1583 19.3944
R17958 vdd.n1648 vdd.n1589 19.3944
R17959 vdd.n1643 vdd.n1589 19.3944
R17960 vdd.n1643 vdd.n1642 19.3944
R17961 vdd.n1642 vdd.n1641 19.3944
R17962 vdd.n1641 vdd.n1596 19.3944
R17963 vdd.n1636 vdd.n1596 19.3944
R17964 vdd.n1636 vdd.n1635 19.3944
R17965 vdd.n1635 vdd.n1634 19.3944
R17966 vdd.n1634 vdd.n1603 19.3944
R17967 vdd.n1629 vdd.n1603 19.3944
R17968 vdd.n1629 vdd.n1628 19.3944
R17969 vdd.n1628 vdd.n1627 19.3944
R17970 vdd.n1627 vdd.n1611 19.3944
R17971 vdd.n1622 vdd.n1611 19.3944
R17972 vdd.n1622 vdd.n1621 19.3944
R17973 vdd.n1617 vdd.n1616 19.3944
R17974 vdd.n1950 vdd.n858 19.3944
R17975 vdd.n1687 vdd.n1543 19.3944
R17976 vdd.n1687 vdd.n1549 19.3944
R17977 vdd.n1682 vdd.n1549 19.3944
R17978 vdd.n1682 vdd.n1681 19.3944
R17979 vdd.n1681 vdd.n1680 19.3944
R17980 vdd.n1680 vdd.n1556 19.3944
R17981 vdd.n1675 vdd.n1556 19.3944
R17982 vdd.n1675 vdd.n1674 19.3944
R17983 vdd.n1674 vdd.n1673 19.3944
R17984 vdd.n1673 vdd.n1563 19.3944
R17985 vdd.n1668 vdd.n1563 19.3944
R17986 vdd.n1668 vdd.n1667 19.3944
R17987 vdd.n1667 vdd.n1666 19.3944
R17988 vdd.n1666 vdd.n1570 19.3944
R17989 vdd.n1661 vdd.n1570 19.3944
R17990 vdd.n1661 vdd.n1660 19.3944
R17991 vdd.n1660 vdd.n1659 19.3944
R17992 vdd.n1659 vdd.n1577 19.3944
R17993 vdd.n1654 vdd.n1577 19.3944
R17994 vdd.n1654 vdd.n1653 19.3944
R17995 vdd.n1938 vdd.n1937 19.3944
R17996 vdd.n1937 vdd.n1515 19.3944
R17997 vdd.n1932 vdd.n1931 19.3944
R17998 vdd.n1714 vdd.n1519 19.3944
R17999 vdd.n1714 vdd.n1521 19.3944
R18000 vdd.n1524 vdd.n1521 19.3944
R18001 vdd.n1707 vdd.n1524 19.3944
R18002 vdd.n1707 vdd.n1706 19.3944
R18003 vdd.n1706 vdd.n1705 19.3944
R18004 vdd.n1705 vdd.n1530 19.3944
R18005 vdd.n1700 vdd.n1530 19.3944
R18006 vdd.n1700 vdd.n1699 19.3944
R18007 vdd.n1699 vdd.n1698 19.3944
R18008 vdd.n1698 vdd.n1537 19.3944
R18009 vdd.n1693 vdd.n1537 19.3944
R18010 vdd.n1693 vdd.n1692 19.3944
R18011 vdd.n1428 vdd.n1193 19.3944
R18012 vdd.n1428 vdd.n1184 19.3944
R18013 vdd.n1441 vdd.n1184 19.3944
R18014 vdd.n1441 vdd.n1182 19.3944
R18015 vdd.n1445 vdd.n1182 19.3944
R18016 vdd.n1445 vdd.n1173 19.3944
R18017 vdd.n1458 vdd.n1173 19.3944
R18018 vdd.n1458 vdd.n1171 19.3944
R18019 vdd.n1463 vdd.n1171 19.3944
R18020 vdd.n1463 vdd.n1162 19.3944
R18021 vdd.n1475 vdd.n1162 19.3944
R18022 vdd.n1475 vdd.n890 19.3944
R18023 vdd.n1479 vdd.n890 19.3944
R18024 vdd.n1479 vdd.n880 19.3944
R18025 vdd.n1492 vdd.n880 19.3944
R18026 vdd.n1492 vdd.n878 19.3944
R18027 vdd.n1496 vdd.n878 19.3944
R18028 vdd.n1496 vdd.n868 19.3944
R18029 vdd.n1511 vdd.n868 19.3944
R18030 vdd.n1511 vdd.n866 19.3944
R18031 vdd.n1941 vdd.n866 19.3944
R18032 vdd.n2851 vdd.n477 19.3944
R18033 vdd.n2851 vdd.n475 19.3944
R18034 vdd.n2855 vdd.n475 19.3944
R18035 vdd.n2855 vdd.n465 19.3944
R18036 vdd.n2868 vdd.n465 19.3944
R18037 vdd.n2868 vdd.n463 19.3944
R18038 vdd.n2872 vdd.n463 19.3944
R18039 vdd.n2872 vdd.n453 19.3944
R18040 vdd.n2884 vdd.n453 19.3944
R18041 vdd.n2884 vdd.n451 19.3944
R18042 vdd.n2888 vdd.n451 19.3944
R18043 vdd.n2889 vdd.n2888 19.3944
R18044 vdd.n2890 vdd.n2889 19.3944
R18045 vdd.n2890 vdd.n449 19.3944
R18046 vdd.n2894 vdd.n449 19.3944
R18047 vdd.n2895 vdd.n2894 19.3944
R18048 vdd.n2896 vdd.n2895 19.3944
R18049 vdd.n2896 vdd.n446 19.3944
R18050 vdd.n2900 vdd.n446 19.3944
R18051 vdd.n2901 vdd.n2900 19.3944
R18052 vdd.n2902 vdd.n2901 19.3944
R18053 vdd.n2945 vdd.n404 19.3944
R18054 vdd.n2945 vdd.n410 19.3944
R18055 vdd.n2940 vdd.n410 19.3944
R18056 vdd.n2940 vdd.n2939 19.3944
R18057 vdd.n2939 vdd.n2938 19.3944
R18058 vdd.n2938 vdd.n417 19.3944
R18059 vdd.n2933 vdd.n417 19.3944
R18060 vdd.n2933 vdd.n2932 19.3944
R18061 vdd.n2932 vdd.n2931 19.3944
R18062 vdd.n2931 vdd.n424 19.3944
R18063 vdd.n2926 vdd.n424 19.3944
R18064 vdd.n2926 vdd.n2925 19.3944
R18065 vdd.n2925 vdd.n2924 19.3944
R18066 vdd.n2924 vdd.n431 19.3944
R18067 vdd.n2919 vdd.n431 19.3944
R18068 vdd.n2919 vdd.n2918 19.3944
R18069 vdd.n2918 vdd.n2917 19.3944
R18070 vdd.n2917 vdd.n438 19.3944
R18071 vdd.n2912 vdd.n438 19.3944
R18072 vdd.n2912 vdd.n2911 19.3944
R18073 vdd.n2984 vdd.n364 19.3944
R18074 vdd.n2984 vdd.n370 19.3944
R18075 vdd.n2979 vdd.n370 19.3944
R18076 vdd.n2979 vdd.n2978 19.3944
R18077 vdd.n2978 vdd.n2977 19.3944
R18078 vdd.n2977 vdd.n377 19.3944
R18079 vdd.n2972 vdd.n377 19.3944
R18080 vdd.n2972 vdd.n2971 19.3944
R18081 vdd.n2971 vdd.n2970 19.3944
R18082 vdd.n2970 vdd.n384 19.3944
R18083 vdd.n2965 vdd.n384 19.3944
R18084 vdd.n2965 vdd.n2964 19.3944
R18085 vdd.n2964 vdd.n2963 19.3944
R18086 vdd.n2963 vdd.n391 19.3944
R18087 vdd.n2958 vdd.n391 19.3944
R18088 vdd.n2958 vdd.n2957 19.3944
R18089 vdd.n2957 vdd.n2956 19.3944
R18090 vdd.n2956 vdd.n398 19.3944
R18091 vdd.n2951 vdd.n398 19.3944
R18092 vdd.n2951 vdd.n2950 19.3944
R18093 vdd.n3020 vdd.n3019 19.3944
R18094 vdd.n3019 vdd.n3018 19.3944
R18095 vdd.n3018 vdd.n336 19.3944
R18096 vdd.n337 vdd.n336 19.3944
R18097 vdd.n3011 vdd.n337 19.3944
R18098 vdd.n3011 vdd.n3010 19.3944
R18099 vdd.n3010 vdd.n3009 19.3944
R18100 vdd.n3009 vdd.n344 19.3944
R18101 vdd.n3004 vdd.n344 19.3944
R18102 vdd.n3004 vdd.n3003 19.3944
R18103 vdd.n3003 vdd.n3002 19.3944
R18104 vdd.n3002 vdd.n351 19.3944
R18105 vdd.n2997 vdd.n351 19.3944
R18106 vdd.n2997 vdd.n2996 19.3944
R18107 vdd.n2996 vdd.n2995 19.3944
R18108 vdd.n2995 vdd.n358 19.3944
R18109 vdd.n2990 vdd.n358 19.3944
R18110 vdd.n2990 vdd.n2989 19.3944
R18111 vdd.n2847 vdd.n480 19.3944
R18112 vdd.n2847 vdd.n471 19.3944
R18113 vdd.n2860 vdd.n471 19.3944
R18114 vdd.n2860 vdd.n469 19.3944
R18115 vdd.n2864 vdd.n469 19.3944
R18116 vdd.n2864 vdd.n460 19.3944
R18117 vdd.n2876 vdd.n460 19.3944
R18118 vdd.n2876 vdd.n458 19.3944
R18119 vdd.n2880 vdd.n458 19.3944
R18120 vdd.n2880 vdd.n300 19.3944
R18121 vdd.n3045 vdd.n300 19.3944
R18122 vdd.n3045 vdd.n301 19.3944
R18123 vdd.n3039 vdd.n301 19.3944
R18124 vdd.n3039 vdd.n3038 19.3944
R18125 vdd.n3038 vdd.n3037 19.3944
R18126 vdd.n3037 vdd.n313 19.3944
R18127 vdd.n3031 vdd.n313 19.3944
R18128 vdd.n3031 vdd.n3030 19.3944
R18129 vdd.n3030 vdd.n3029 19.3944
R18130 vdd.n3029 vdd.n324 19.3944
R18131 vdd.n3023 vdd.n324 19.3944
R18132 vdd.n2800 vdd.n536 19.3944
R18133 vdd.n2800 vdd.n2797 19.3944
R18134 vdd.n2797 vdd.n2794 19.3944
R18135 vdd.n2794 vdd.n2793 19.3944
R18136 vdd.n2793 vdd.n2790 19.3944
R18137 vdd.n2790 vdd.n2789 19.3944
R18138 vdd.n2789 vdd.n2786 19.3944
R18139 vdd.n2786 vdd.n2785 19.3944
R18140 vdd.n2785 vdd.n2782 19.3944
R18141 vdd.n2782 vdd.n2781 19.3944
R18142 vdd.n2781 vdd.n2778 19.3944
R18143 vdd.n2778 vdd.n2777 19.3944
R18144 vdd.n2777 vdd.n2774 19.3944
R18145 vdd.n2774 vdd.n2773 19.3944
R18146 vdd.n2773 vdd.n2770 19.3944
R18147 vdd.n2770 vdd.n2769 19.3944
R18148 vdd.n2769 vdd.n2766 19.3944
R18149 vdd.n2766 vdd.n2765 19.3944
R18150 vdd.n2765 vdd.n2762 19.3944
R18151 vdd.n2762 vdd.n2761 19.3944
R18152 vdd.n2843 vdd.n482 19.3944
R18153 vdd.n2838 vdd.n482 19.3944
R18154 vdd.n521 vdd.n518 19.3944
R18155 vdd.n2834 vdd.n2833 19.3944
R18156 vdd.n2833 vdd.n2830 19.3944
R18157 vdd.n2830 vdd.n2829 19.3944
R18158 vdd.n2829 vdd.n2826 19.3944
R18159 vdd.n2826 vdd.n2825 19.3944
R18160 vdd.n2825 vdd.n2822 19.3944
R18161 vdd.n2822 vdd.n2821 19.3944
R18162 vdd.n2821 vdd.n2818 19.3944
R18163 vdd.n2818 vdd.n2817 19.3944
R18164 vdd.n2817 vdd.n2814 19.3944
R18165 vdd.n2814 vdd.n2813 19.3944
R18166 vdd.n2813 vdd.n2810 19.3944
R18167 vdd.n2810 vdd.n2809 19.3944
R18168 vdd.n2754 vdd.n556 19.3944
R18169 vdd.n2754 vdd.n2751 19.3944
R18170 vdd.n2751 vdd.n2748 19.3944
R18171 vdd.n2748 vdd.n2747 19.3944
R18172 vdd.n2747 vdd.n2744 19.3944
R18173 vdd.n2744 vdd.n2743 19.3944
R18174 vdd.n2743 vdd.n2740 19.3944
R18175 vdd.n2740 vdd.n2739 19.3944
R18176 vdd.n2739 vdd.n2736 19.3944
R18177 vdd.n2736 vdd.n2735 19.3944
R18178 vdd.n2735 vdd.n2732 19.3944
R18179 vdd.n2732 vdd.n2731 19.3944
R18180 vdd.n2731 vdd.n2728 19.3944
R18181 vdd.n2728 vdd.n2727 19.3944
R18182 vdd.n2727 vdd.n2724 19.3944
R18183 vdd.n2724 vdd.n2723 19.3944
R18184 vdd.n2720 vdd.n2719 19.3944
R18185 vdd.n2716 vdd.n2715 19.3944
R18186 vdd.n1360 vdd.n1356 19.0066
R18187 vdd.n1652 vdd.n1583 19.0066
R18188 vdd.n2949 vdd.n404 19.0066
R18189 vdd.n2758 vdd.n556 19.0066
R18190 vdd.n1792 vdd.n1791 16.0975
R18191 vdd.n756 vdd.n755 16.0975
R18192 vdd.n1321 vdd.n1320 16.0975
R18193 vdd.n1359 vdd.n1358 16.0975
R18194 vdd.n1255 vdd.n1254 16.0975
R18195 vdd.n1948 vdd.n1947 16.0975
R18196 vdd.n1585 vdd.n1584 16.0975
R18197 vdd.n1545 vdd.n1544 16.0975
R18198 vdd.n1766 vdd.n1765 16.0975
R18199 vdd.n748 vdd.n747 16.0975
R18200 vdd.n2257 vdd.n2256 16.0975
R18201 vdd.n2909 vdd.n2908 16.0975
R18202 vdd.n406 vdd.n405 16.0975
R18203 vdd.n366 vdd.n365 16.0975
R18204 vdd.n558 vdd.n557 16.0975
R18205 vdd.n2805 vdd.n2804 16.0975
R18206 vdd.n623 vdd.n622 16.0975
R18207 vdd.n2254 vdd.n2253 16.0975
R18208 vdd.n2712 vdd.n2711 16.0975
R18209 vdd.n590 vdd.n589 16.0975
R18210 vdd.t111 vdd.n2218 15.4182
R18211 vdd.n2471 vdd.t118 15.4182
R18212 vdd.n1989 vdd.n839 14.5112
R18213 vdd.n2673 vdd.n484 14.5112
R18214 vdd.n28 vdd.n27 14.4007
R18215 vdd.n292 vdd.n257 13.1884
R18216 vdd.n245 vdd.n210 13.1884
R18217 vdd.n202 vdd.n167 13.1884
R18218 vdd.n155 vdd.n120 13.1884
R18219 vdd.n113 vdd.n78 13.1884
R18220 vdd.n66 vdd.n31 13.1884
R18221 vdd.n1107 vdd.n1072 13.1884
R18222 vdd.n1154 vdd.n1119 13.1884
R18223 vdd.n1017 vdd.n982 13.1884
R18224 vdd.n1064 vdd.n1029 13.1884
R18225 vdd.n928 vdd.n893 13.1884
R18226 vdd.n975 vdd.n940 13.1884
R18227 vdd.n1391 vdd.n1256 12.9944
R18228 vdd.n1395 vdd.n1256 12.9944
R18229 vdd.n1691 vdd.n1543 12.9944
R18230 vdd.n1692 vdd.n1691 12.9944
R18231 vdd.n2988 vdd.n364 12.9944
R18232 vdd.n2989 vdd.n2988 12.9944
R18233 vdd.n2806 vdd.n536 12.9944
R18234 vdd.n2809 vdd.n2806 12.9944
R18235 vdd.n293 vdd.n255 12.8005
R18236 vdd.n288 vdd.n259 12.8005
R18237 vdd.n246 vdd.n208 12.8005
R18238 vdd.n241 vdd.n212 12.8005
R18239 vdd.n203 vdd.n165 12.8005
R18240 vdd.n198 vdd.n169 12.8005
R18241 vdd.n156 vdd.n118 12.8005
R18242 vdd.n151 vdd.n122 12.8005
R18243 vdd.n114 vdd.n76 12.8005
R18244 vdd.n109 vdd.n80 12.8005
R18245 vdd.n67 vdd.n29 12.8005
R18246 vdd.n62 vdd.n33 12.8005
R18247 vdd.n1108 vdd.n1070 12.8005
R18248 vdd.n1103 vdd.n1074 12.8005
R18249 vdd.n1155 vdd.n1117 12.8005
R18250 vdd.n1150 vdd.n1121 12.8005
R18251 vdd.n1018 vdd.n980 12.8005
R18252 vdd.n1013 vdd.n984 12.8005
R18253 vdd.n1065 vdd.n1027 12.8005
R18254 vdd.n1060 vdd.n1031 12.8005
R18255 vdd.n929 vdd.n891 12.8005
R18256 vdd.n924 vdd.n895 12.8005
R18257 vdd.n976 vdd.n938 12.8005
R18258 vdd.n971 vdd.n942 12.8005
R18259 vdd.n287 vdd.n260 12.0247
R18260 vdd.n240 vdd.n213 12.0247
R18261 vdd.n197 vdd.n170 12.0247
R18262 vdd.n150 vdd.n123 12.0247
R18263 vdd.n108 vdd.n81 12.0247
R18264 vdd.n61 vdd.n34 12.0247
R18265 vdd.n1102 vdd.n1075 12.0247
R18266 vdd.n1149 vdd.n1122 12.0247
R18267 vdd.n1012 vdd.n985 12.0247
R18268 vdd.n1059 vdd.n1032 12.0247
R18269 vdd.n923 vdd.n896 12.0247
R18270 vdd.n970 vdd.n943 12.0247
R18271 vdd.n1430 vdd.n1186 11.337
R18272 vdd.n1439 vdd.n1186 11.337
R18273 vdd.n1439 vdd.n1438 11.337
R18274 vdd.n1447 vdd.n1180 11.337
R18275 vdd.n1456 vdd.n1455 11.337
R18276 vdd.n1473 vdd.n1164 11.337
R18277 vdd.n1481 vdd.n887 11.337
R18278 vdd.n1490 vdd.n1489 11.337
R18279 vdd.n1498 vdd.n870 11.337
R18280 vdd.n1509 vdd.n870 11.337
R18281 vdd.n1509 vdd.n1508 11.337
R18282 vdd.n2849 vdd.n473 11.337
R18283 vdd.n2858 vdd.n473 11.337
R18284 vdd.n2858 vdd.n2857 11.337
R18285 vdd.n2866 vdd.n467 11.337
R18286 vdd.n2882 vdd.n456 11.337
R18287 vdd.n3043 vdd.n304 11.337
R18288 vdd.n3041 vdd.n308 11.337
R18289 vdd.n3035 vdd.n3034 11.337
R18290 vdd.n3033 vdd.n318 11.337
R18291 vdd.n3027 vdd.n318 11.337
R18292 vdd.n3027 vdd.n3026 11.337
R18293 vdd.n284 vdd.n283 11.249
R18294 vdd.n237 vdd.n236 11.249
R18295 vdd.n194 vdd.n193 11.249
R18296 vdd.n147 vdd.n146 11.249
R18297 vdd.n105 vdd.n104 11.249
R18298 vdd.n58 vdd.n57 11.249
R18299 vdd.n1099 vdd.n1098 11.249
R18300 vdd.n1146 vdd.n1145 11.249
R18301 vdd.n1009 vdd.n1008 11.249
R18302 vdd.n1056 vdd.n1055 11.249
R18303 vdd.n920 vdd.n919 11.249
R18304 vdd.n967 vdd.n966 11.249
R18305 vdd.n2146 vdd.t122 11.1103
R18306 vdd.n2478 vdd.t13 11.1103
R18307 vdd.n1228 vdd.t136 10.7702
R18308 vdd.t147 vdd.n3025 10.7702
R18309 vdd.n269 vdd.n268 10.7238
R18310 vdd.n222 vdd.n221 10.7238
R18311 vdd.n179 vdd.n178 10.7238
R18312 vdd.n132 vdd.n131 10.7238
R18313 vdd.n90 vdd.n89 10.7238
R18314 vdd.n43 vdd.n42 10.7238
R18315 vdd.n1084 vdd.n1083 10.7238
R18316 vdd.n1131 vdd.n1130 10.7238
R18317 vdd.n994 vdd.n993 10.7238
R18318 vdd.n1041 vdd.n1040 10.7238
R18319 vdd.n905 vdd.n904 10.7238
R18320 vdd.n952 vdd.n951 10.7238
R18321 vdd.n1992 vdd.n1991 10.6151
R18322 vdd.n1993 vdd.n1992 10.6151
R18323 vdd.n1993 vdd.n825 10.6151
R18324 vdd.n2003 vdd.n825 10.6151
R18325 vdd.n2004 vdd.n2003 10.6151
R18326 vdd.n2005 vdd.n2004 10.6151
R18327 vdd.n2005 vdd.n812 10.6151
R18328 vdd.n2016 vdd.n812 10.6151
R18329 vdd.n2017 vdd.n2016 10.6151
R18330 vdd.n2018 vdd.n2017 10.6151
R18331 vdd.n2018 vdd.n800 10.6151
R18332 vdd.n2028 vdd.n800 10.6151
R18333 vdd.n2029 vdd.n2028 10.6151
R18334 vdd.n2030 vdd.n2029 10.6151
R18335 vdd.n2030 vdd.n788 10.6151
R18336 vdd.n2040 vdd.n788 10.6151
R18337 vdd.n2041 vdd.n2040 10.6151
R18338 vdd.n2042 vdd.n2041 10.6151
R18339 vdd.n2042 vdd.n777 10.6151
R18340 vdd.n2052 vdd.n777 10.6151
R18341 vdd.n2053 vdd.n2052 10.6151
R18342 vdd.n2054 vdd.n2053 10.6151
R18343 vdd.n2054 vdd.n764 10.6151
R18344 vdd.n2066 vdd.n764 10.6151
R18345 vdd.n2067 vdd.n2066 10.6151
R18346 vdd.n2069 vdd.n2067 10.6151
R18347 vdd.n2069 vdd.n2068 10.6151
R18348 vdd.n2068 vdd.n746 10.6151
R18349 vdd.n2216 vdd.n2215 10.6151
R18350 vdd.n2215 vdd.n2214 10.6151
R18351 vdd.n2214 vdd.n2211 10.6151
R18352 vdd.n2211 vdd.n2210 10.6151
R18353 vdd.n2210 vdd.n2207 10.6151
R18354 vdd.n2207 vdd.n2206 10.6151
R18355 vdd.n2206 vdd.n2203 10.6151
R18356 vdd.n2203 vdd.n2202 10.6151
R18357 vdd.n2202 vdd.n2199 10.6151
R18358 vdd.n2199 vdd.n2198 10.6151
R18359 vdd.n2198 vdd.n2195 10.6151
R18360 vdd.n2195 vdd.n2194 10.6151
R18361 vdd.n2194 vdd.n2191 10.6151
R18362 vdd.n2191 vdd.n2190 10.6151
R18363 vdd.n2190 vdd.n2187 10.6151
R18364 vdd.n2187 vdd.n2186 10.6151
R18365 vdd.n2186 vdd.n2183 10.6151
R18366 vdd.n2183 vdd.n2182 10.6151
R18367 vdd.n2182 vdd.n2179 10.6151
R18368 vdd.n2179 vdd.n2178 10.6151
R18369 vdd.n2178 vdd.n2175 10.6151
R18370 vdd.n2175 vdd.n2174 10.6151
R18371 vdd.n2174 vdd.n2171 10.6151
R18372 vdd.n2171 vdd.n2170 10.6151
R18373 vdd.n2170 vdd.n2167 10.6151
R18374 vdd.n2167 vdd.n2166 10.6151
R18375 vdd.n2166 vdd.n2163 10.6151
R18376 vdd.n2163 vdd.n2162 10.6151
R18377 vdd.n2162 vdd.n2159 10.6151
R18378 vdd.n2159 vdd.n2158 10.6151
R18379 vdd.n2158 vdd.n2155 10.6151
R18380 vdd.n2153 vdd.n2150 10.6151
R18381 vdd.n2150 vdd.n2149 10.6151
R18382 vdd.n1892 vdd.n1891 10.6151
R18383 vdd.n1891 vdd.n1889 10.6151
R18384 vdd.n1889 vdd.n1888 10.6151
R18385 vdd.n1888 vdd.n1886 10.6151
R18386 vdd.n1886 vdd.n1885 10.6151
R18387 vdd.n1885 vdd.n1883 10.6151
R18388 vdd.n1883 vdd.n1882 10.6151
R18389 vdd.n1882 vdd.n1880 10.6151
R18390 vdd.n1880 vdd.n1879 10.6151
R18391 vdd.n1879 vdd.n1877 10.6151
R18392 vdd.n1877 vdd.n1876 10.6151
R18393 vdd.n1876 vdd.n1874 10.6151
R18394 vdd.n1874 vdd.n1873 10.6151
R18395 vdd.n1873 vdd.n1788 10.6151
R18396 vdd.n1788 vdd.n1787 10.6151
R18397 vdd.n1787 vdd.n1785 10.6151
R18398 vdd.n1785 vdd.n1784 10.6151
R18399 vdd.n1784 vdd.n1782 10.6151
R18400 vdd.n1782 vdd.n1781 10.6151
R18401 vdd.n1781 vdd.n1779 10.6151
R18402 vdd.n1779 vdd.n1778 10.6151
R18403 vdd.n1778 vdd.n1776 10.6151
R18404 vdd.n1776 vdd.n1775 10.6151
R18405 vdd.n1775 vdd.n1773 10.6151
R18406 vdd.n1773 vdd.n1772 10.6151
R18407 vdd.n1772 vdd.n1769 10.6151
R18408 vdd.n1769 vdd.n1768 10.6151
R18409 vdd.n1768 vdd.n749 10.6151
R18410 vdd.n1726 vdd.n837 10.6151
R18411 vdd.n1727 vdd.n1726 10.6151
R18412 vdd.n1728 vdd.n1727 10.6151
R18413 vdd.n1728 vdd.n1722 10.6151
R18414 vdd.n1734 vdd.n1722 10.6151
R18415 vdd.n1735 vdd.n1734 10.6151
R18416 vdd.n1736 vdd.n1735 10.6151
R18417 vdd.n1736 vdd.n1720 10.6151
R18418 vdd.n1742 vdd.n1720 10.6151
R18419 vdd.n1743 vdd.n1742 10.6151
R18420 vdd.n1744 vdd.n1743 10.6151
R18421 vdd.n1744 vdd.n1718 10.6151
R18422 vdd.n1750 vdd.n1718 10.6151
R18423 vdd.n1751 vdd.n1750 10.6151
R18424 vdd.n1752 vdd.n1751 10.6151
R18425 vdd.n1752 vdd.n1716 10.6151
R18426 vdd.n1928 vdd.n1716 10.6151
R18427 vdd.n1928 vdd.n1927 10.6151
R18428 vdd.n1927 vdd.n1757 10.6151
R18429 vdd.n1921 vdd.n1757 10.6151
R18430 vdd.n1921 vdd.n1920 10.6151
R18431 vdd.n1920 vdd.n1919 10.6151
R18432 vdd.n1919 vdd.n1759 10.6151
R18433 vdd.n1913 vdd.n1759 10.6151
R18434 vdd.n1913 vdd.n1912 10.6151
R18435 vdd.n1912 vdd.n1911 10.6151
R18436 vdd.n1911 vdd.n1761 10.6151
R18437 vdd.n1905 vdd.n1761 10.6151
R18438 vdd.n1905 vdd.n1904 10.6151
R18439 vdd.n1904 vdd.n1903 10.6151
R18440 vdd.n1903 vdd.n1763 10.6151
R18441 vdd.n1897 vdd.n1896 10.6151
R18442 vdd.n1896 vdd.n1895 10.6151
R18443 vdd.n2401 vdd.n2400 10.6151
R18444 vdd.n2400 vdd.n2398 10.6151
R18445 vdd.n2398 vdd.n2397 10.6151
R18446 vdd.n2397 vdd.n2255 10.6151
R18447 vdd.n2344 vdd.n2255 10.6151
R18448 vdd.n2345 vdd.n2344 10.6151
R18449 vdd.n2347 vdd.n2345 10.6151
R18450 vdd.n2348 vdd.n2347 10.6151
R18451 vdd.n2350 vdd.n2348 10.6151
R18452 vdd.n2351 vdd.n2350 10.6151
R18453 vdd.n2353 vdd.n2351 10.6151
R18454 vdd.n2354 vdd.n2353 10.6151
R18455 vdd.n2356 vdd.n2354 10.6151
R18456 vdd.n2357 vdd.n2356 10.6151
R18457 vdd.n2372 vdd.n2357 10.6151
R18458 vdd.n2372 vdd.n2371 10.6151
R18459 vdd.n2371 vdd.n2370 10.6151
R18460 vdd.n2370 vdd.n2368 10.6151
R18461 vdd.n2368 vdd.n2367 10.6151
R18462 vdd.n2367 vdd.n2365 10.6151
R18463 vdd.n2365 vdd.n2364 10.6151
R18464 vdd.n2364 vdd.n2362 10.6151
R18465 vdd.n2362 vdd.n2361 10.6151
R18466 vdd.n2361 vdd.n2359 10.6151
R18467 vdd.n2359 vdd.n2358 10.6151
R18468 vdd.n2358 vdd.n626 10.6151
R18469 vdd.n2606 vdd.n626 10.6151
R18470 vdd.n2607 vdd.n2606 10.6151
R18471 vdd.n2468 vdd.n702 10.6151
R18472 vdd.n2468 vdd.n2467 10.6151
R18473 vdd.n2467 vdd.n2466 10.6151
R18474 vdd.n2466 vdd.n2464 10.6151
R18475 vdd.n2464 vdd.n2461 10.6151
R18476 vdd.n2461 vdd.n2460 10.6151
R18477 vdd.n2460 vdd.n2457 10.6151
R18478 vdd.n2457 vdd.n2456 10.6151
R18479 vdd.n2456 vdd.n2453 10.6151
R18480 vdd.n2453 vdd.n2452 10.6151
R18481 vdd.n2452 vdd.n2449 10.6151
R18482 vdd.n2449 vdd.n2448 10.6151
R18483 vdd.n2448 vdd.n2445 10.6151
R18484 vdd.n2445 vdd.n2444 10.6151
R18485 vdd.n2444 vdd.n2441 10.6151
R18486 vdd.n2441 vdd.n2440 10.6151
R18487 vdd.n2440 vdd.n2437 10.6151
R18488 vdd.n2437 vdd.n2436 10.6151
R18489 vdd.n2436 vdd.n2433 10.6151
R18490 vdd.n2433 vdd.n2432 10.6151
R18491 vdd.n2432 vdd.n2429 10.6151
R18492 vdd.n2429 vdd.n2428 10.6151
R18493 vdd.n2428 vdd.n2425 10.6151
R18494 vdd.n2425 vdd.n2424 10.6151
R18495 vdd.n2424 vdd.n2421 10.6151
R18496 vdd.n2421 vdd.n2420 10.6151
R18497 vdd.n2420 vdd.n2417 10.6151
R18498 vdd.n2417 vdd.n2416 10.6151
R18499 vdd.n2416 vdd.n2413 10.6151
R18500 vdd.n2413 vdd.n2412 10.6151
R18501 vdd.n2412 vdd.n2409 10.6151
R18502 vdd.n2407 vdd.n2404 10.6151
R18503 vdd.n2404 vdd.n2403 10.6151
R18504 vdd.n2481 vdd.n2480 10.6151
R18505 vdd.n2482 vdd.n2481 10.6151
R18506 vdd.n2482 vdd.n692 10.6151
R18507 vdd.n2492 vdd.n692 10.6151
R18508 vdd.n2493 vdd.n2492 10.6151
R18509 vdd.n2494 vdd.n2493 10.6151
R18510 vdd.n2494 vdd.n679 10.6151
R18511 vdd.n2504 vdd.n679 10.6151
R18512 vdd.n2505 vdd.n2504 10.6151
R18513 vdd.n2506 vdd.n2505 10.6151
R18514 vdd.n2506 vdd.n668 10.6151
R18515 vdd.n2516 vdd.n668 10.6151
R18516 vdd.n2517 vdd.n2516 10.6151
R18517 vdd.n2518 vdd.n2517 10.6151
R18518 vdd.n2518 vdd.n656 10.6151
R18519 vdd.n2528 vdd.n656 10.6151
R18520 vdd.n2529 vdd.n2528 10.6151
R18521 vdd.n2530 vdd.n2529 10.6151
R18522 vdd.n2530 vdd.n645 10.6151
R18523 vdd.n2542 vdd.n645 10.6151
R18524 vdd.n2543 vdd.n2542 10.6151
R18525 vdd.n2544 vdd.n2543 10.6151
R18526 vdd.n2544 vdd.n631 10.6151
R18527 vdd.n2599 vdd.n631 10.6151
R18528 vdd.n2600 vdd.n2599 10.6151
R18529 vdd.n2601 vdd.n2600 10.6151
R18530 vdd.n2601 vdd.n600 10.6151
R18531 vdd.n2671 vdd.n600 10.6151
R18532 vdd.n2670 vdd.n2669 10.6151
R18533 vdd.n2669 vdd.n601 10.6151
R18534 vdd.n602 vdd.n601 10.6151
R18535 vdd.n2662 vdd.n602 10.6151
R18536 vdd.n2662 vdd.n2661 10.6151
R18537 vdd.n2661 vdd.n2660 10.6151
R18538 vdd.n2660 vdd.n604 10.6151
R18539 vdd.n2655 vdd.n604 10.6151
R18540 vdd.n2655 vdd.n2654 10.6151
R18541 vdd.n2654 vdd.n2653 10.6151
R18542 vdd.n2653 vdd.n607 10.6151
R18543 vdd.n2648 vdd.n607 10.6151
R18544 vdd.n2648 vdd.n2647 10.6151
R18545 vdd.n2647 vdd.n2646 10.6151
R18546 vdd.n2646 vdd.n610 10.6151
R18547 vdd.n2641 vdd.n610 10.6151
R18548 vdd.n2641 vdd.n520 10.6151
R18549 vdd.n2637 vdd.n520 10.6151
R18550 vdd.n2637 vdd.n2636 10.6151
R18551 vdd.n2636 vdd.n2635 10.6151
R18552 vdd.n2635 vdd.n613 10.6151
R18553 vdd.n2630 vdd.n613 10.6151
R18554 vdd.n2630 vdd.n2629 10.6151
R18555 vdd.n2629 vdd.n2628 10.6151
R18556 vdd.n2628 vdd.n616 10.6151
R18557 vdd.n2623 vdd.n616 10.6151
R18558 vdd.n2623 vdd.n2622 10.6151
R18559 vdd.n2622 vdd.n2621 10.6151
R18560 vdd.n2621 vdd.n619 10.6151
R18561 vdd.n2616 vdd.n619 10.6151
R18562 vdd.n2616 vdd.n2615 10.6151
R18563 vdd.n2613 vdd.n624 10.6151
R18564 vdd.n2608 vdd.n624 10.6151
R18565 vdd.n2589 vdd.n2550 10.6151
R18566 vdd.n2584 vdd.n2550 10.6151
R18567 vdd.n2584 vdd.n2583 10.6151
R18568 vdd.n2583 vdd.n2582 10.6151
R18569 vdd.n2582 vdd.n2552 10.6151
R18570 vdd.n2577 vdd.n2552 10.6151
R18571 vdd.n2577 vdd.n2576 10.6151
R18572 vdd.n2576 vdd.n2575 10.6151
R18573 vdd.n2575 vdd.n2555 10.6151
R18574 vdd.n2570 vdd.n2555 10.6151
R18575 vdd.n2570 vdd.n2569 10.6151
R18576 vdd.n2569 vdd.n2568 10.6151
R18577 vdd.n2568 vdd.n2558 10.6151
R18578 vdd.n2563 vdd.n2558 10.6151
R18579 vdd.n2563 vdd.n2562 10.6151
R18580 vdd.n2562 vdd.n575 10.6151
R18581 vdd.n2706 vdd.n575 10.6151
R18582 vdd.n2706 vdd.n576 10.6151
R18583 vdd.n578 vdd.n576 10.6151
R18584 vdd.n2699 vdd.n578 10.6151
R18585 vdd.n2699 vdd.n2698 10.6151
R18586 vdd.n2698 vdd.n2697 10.6151
R18587 vdd.n2697 vdd.n580 10.6151
R18588 vdd.n2692 vdd.n580 10.6151
R18589 vdd.n2692 vdd.n2691 10.6151
R18590 vdd.n2691 vdd.n2690 10.6151
R18591 vdd.n2690 vdd.n583 10.6151
R18592 vdd.n2685 vdd.n583 10.6151
R18593 vdd.n2685 vdd.n2684 10.6151
R18594 vdd.n2684 vdd.n2683 10.6151
R18595 vdd.n2683 vdd.n586 10.6151
R18596 vdd.n2678 vdd.n2677 10.6151
R18597 vdd.n2677 vdd.n2676 10.6151
R18598 vdd.n2324 vdd.n2322 10.6151
R18599 vdd.n2325 vdd.n2324 10.6151
R18600 vdd.n2393 vdd.n2325 10.6151
R18601 vdd.n2393 vdd.n2392 10.6151
R18602 vdd.n2392 vdd.n2391 10.6151
R18603 vdd.n2391 vdd.n2389 10.6151
R18604 vdd.n2389 vdd.n2388 10.6151
R18605 vdd.n2388 vdd.n2386 10.6151
R18606 vdd.n2386 vdd.n2385 10.6151
R18607 vdd.n2385 vdd.n2383 10.6151
R18608 vdd.n2383 vdd.n2382 10.6151
R18609 vdd.n2382 vdd.n2380 10.6151
R18610 vdd.n2380 vdd.n2379 10.6151
R18611 vdd.n2379 vdd.n2377 10.6151
R18612 vdd.n2377 vdd.n2376 10.6151
R18613 vdd.n2376 vdd.n2342 10.6151
R18614 vdd.n2342 vdd.n2341 10.6151
R18615 vdd.n2341 vdd.n2339 10.6151
R18616 vdd.n2339 vdd.n2338 10.6151
R18617 vdd.n2338 vdd.n2336 10.6151
R18618 vdd.n2336 vdd.n2335 10.6151
R18619 vdd.n2335 vdd.n2333 10.6151
R18620 vdd.n2333 vdd.n2332 10.6151
R18621 vdd.n2332 vdd.n2330 10.6151
R18622 vdd.n2330 vdd.n2329 10.6151
R18623 vdd.n2329 vdd.n2327 10.6151
R18624 vdd.n2327 vdd.n2326 10.6151
R18625 vdd.n2326 vdd.n592 10.6151
R18626 vdd.n2475 vdd.n2474 10.6151
R18627 vdd.n2474 vdd.n707 10.6151
R18628 vdd.n2259 vdd.n707 10.6151
R18629 vdd.n2262 vdd.n2259 10.6151
R18630 vdd.n2263 vdd.n2262 10.6151
R18631 vdd.n2266 vdd.n2263 10.6151
R18632 vdd.n2267 vdd.n2266 10.6151
R18633 vdd.n2270 vdd.n2267 10.6151
R18634 vdd.n2271 vdd.n2270 10.6151
R18635 vdd.n2274 vdd.n2271 10.6151
R18636 vdd.n2275 vdd.n2274 10.6151
R18637 vdd.n2278 vdd.n2275 10.6151
R18638 vdd.n2279 vdd.n2278 10.6151
R18639 vdd.n2282 vdd.n2279 10.6151
R18640 vdd.n2283 vdd.n2282 10.6151
R18641 vdd.n2286 vdd.n2283 10.6151
R18642 vdd.n2287 vdd.n2286 10.6151
R18643 vdd.n2290 vdd.n2287 10.6151
R18644 vdd.n2291 vdd.n2290 10.6151
R18645 vdd.n2294 vdd.n2291 10.6151
R18646 vdd.n2295 vdd.n2294 10.6151
R18647 vdd.n2298 vdd.n2295 10.6151
R18648 vdd.n2299 vdd.n2298 10.6151
R18649 vdd.n2302 vdd.n2299 10.6151
R18650 vdd.n2303 vdd.n2302 10.6151
R18651 vdd.n2306 vdd.n2303 10.6151
R18652 vdd.n2307 vdd.n2306 10.6151
R18653 vdd.n2310 vdd.n2307 10.6151
R18654 vdd.n2311 vdd.n2310 10.6151
R18655 vdd.n2314 vdd.n2311 10.6151
R18656 vdd.n2315 vdd.n2314 10.6151
R18657 vdd.n2320 vdd.n2318 10.6151
R18658 vdd.n2321 vdd.n2320 10.6151
R18659 vdd.n2476 vdd.n697 10.6151
R18660 vdd.n2486 vdd.n697 10.6151
R18661 vdd.n2487 vdd.n2486 10.6151
R18662 vdd.n2488 vdd.n2487 10.6151
R18663 vdd.n2488 vdd.n685 10.6151
R18664 vdd.n2498 vdd.n685 10.6151
R18665 vdd.n2499 vdd.n2498 10.6151
R18666 vdd.n2500 vdd.n2499 10.6151
R18667 vdd.n2500 vdd.n674 10.6151
R18668 vdd.n2510 vdd.n674 10.6151
R18669 vdd.n2511 vdd.n2510 10.6151
R18670 vdd.n2512 vdd.n2511 10.6151
R18671 vdd.n2512 vdd.n662 10.6151
R18672 vdd.n2522 vdd.n662 10.6151
R18673 vdd.n2523 vdd.n2522 10.6151
R18674 vdd.n2524 vdd.n2523 10.6151
R18675 vdd.n2524 vdd.n651 10.6151
R18676 vdd.n2534 vdd.n651 10.6151
R18677 vdd.n2535 vdd.n2534 10.6151
R18678 vdd.n2538 vdd.n2535 10.6151
R18679 vdd.n2548 vdd.n639 10.6151
R18680 vdd.n2549 vdd.n2548 10.6151
R18681 vdd.n2595 vdd.n2549 10.6151
R18682 vdd.n2595 vdd.n2594 10.6151
R18683 vdd.n2594 vdd.n2593 10.6151
R18684 vdd.n2593 vdd.n2592 10.6151
R18685 vdd.n2592 vdd.n2590 10.6151
R18686 vdd.n1987 vdd.n831 10.6151
R18687 vdd.n1997 vdd.n831 10.6151
R18688 vdd.n1998 vdd.n1997 10.6151
R18689 vdd.n1999 vdd.n1998 10.6151
R18690 vdd.n1999 vdd.n818 10.6151
R18691 vdd.n2009 vdd.n818 10.6151
R18692 vdd.n2010 vdd.n2009 10.6151
R18693 vdd.n2012 vdd.n806 10.6151
R18694 vdd.n2022 vdd.n806 10.6151
R18695 vdd.n2023 vdd.n2022 10.6151
R18696 vdd.n2024 vdd.n2023 10.6151
R18697 vdd.n2024 vdd.n794 10.6151
R18698 vdd.n2034 vdd.n794 10.6151
R18699 vdd.n2035 vdd.n2034 10.6151
R18700 vdd.n2036 vdd.n2035 10.6151
R18701 vdd.n2036 vdd.n783 10.6151
R18702 vdd.n2046 vdd.n783 10.6151
R18703 vdd.n2047 vdd.n2046 10.6151
R18704 vdd.n2048 vdd.n2047 10.6151
R18705 vdd.n2048 vdd.n771 10.6151
R18706 vdd.n2058 vdd.n771 10.6151
R18707 vdd.n2059 vdd.n2058 10.6151
R18708 vdd.n2062 vdd.n2059 10.6151
R18709 vdd.n2062 vdd.n2061 10.6151
R18710 vdd.n2061 vdd.n2060 10.6151
R18711 vdd.n2060 vdd.n754 10.6151
R18712 vdd.n2144 vdd.n754 10.6151
R18713 vdd.n2143 vdd.n2142 10.6151
R18714 vdd.n2142 vdd.n2139 10.6151
R18715 vdd.n2139 vdd.n2138 10.6151
R18716 vdd.n2138 vdd.n2135 10.6151
R18717 vdd.n2135 vdd.n2134 10.6151
R18718 vdd.n2134 vdd.n2131 10.6151
R18719 vdd.n2131 vdd.n2130 10.6151
R18720 vdd.n2130 vdd.n2127 10.6151
R18721 vdd.n2127 vdd.n2126 10.6151
R18722 vdd.n2126 vdd.n2123 10.6151
R18723 vdd.n2123 vdd.n2122 10.6151
R18724 vdd.n2122 vdd.n2119 10.6151
R18725 vdd.n2119 vdd.n2118 10.6151
R18726 vdd.n2118 vdd.n2115 10.6151
R18727 vdd.n2115 vdd.n2114 10.6151
R18728 vdd.n2114 vdd.n2111 10.6151
R18729 vdd.n2111 vdd.n2110 10.6151
R18730 vdd.n2110 vdd.n2107 10.6151
R18731 vdd.n2107 vdd.n2106 10.6151
R18732 vdd.n2106 vdd.n2103 10.6151
R18733 vdd.n2103 vdd.n2102 10.6151
R18734 vdd.n2102 vdd.n2099 10.6151
R18735 vdd.n2099 vdd.n2098 10.6151
R18736 vdd.n2098 vdd.n2095 10.6151
R18737 vdd.n2095 vdd.n2094 10.6151
R18738 vdd.n2094 vdd.n2091 10.6151
R18739 vdd.n2091 vdd.n2090 10.6151
R18740 vdd.n2090 vdd.n2087 10.6151
R18741 vdd.n2087 vdd.n2086 10.6151
R18742 vdd.n2086 vdd.n2083 10.6151
R18743 vdd.n2083 vdd.n2082 10.6151
R18744 vdd.n2079 vdd.n2078 10.6151
R18745 vdd.n2078 vdd.n2076 10.6151
R18746 vdd.n1835 vdd.n1833 10.6151
R18747 vdd.n1836 vdd.n1835 10.6151
R18748 vdd.n1838 vdd.n1836 10.6151
R18749 vdd.n1839 vdd.n1838 10.6151
R18750 vdd.n1841 vdd.n1839 10.6151
R18751 vdd.n1842 vdd.n1841 10.6151
R18752 vdd.n1844 vdd.n1842 10.6151
R18753 vdd.n1845 vdd.n1844 10.6151
R18754 vdd.n1847 vdd.n1845 10.6151
R18755 vdd.n1848 vdd.n1847 10.6151
R18756 vdd.n1850 vdd.n1848 10.6151
R18757 vdd.n1851 vdd.n1850 10.6151
R18758 vdd.n1869 vdd.n1851 10.6151
R18759 vdd.n1869 vdd.n1868 10.6151
R18760 vdd.n1868 vdd.n1867 10.6151
R18761 vdd.n1867 vdd.n1865 10.6151
R18762 vdd.n1865 vdd.n1864 10.6151
R18763 vdd.n1864 vdd.n1862 10.6151
R18764 vdd.n1862 vdd.n1861 10.6151
R18765 vdd.n1861 vdd.n1859 10.6151
R18766 vdd.n1859 vdd.n1858 10.6151
R18767 vdd.n1858 vdd.n1856 10.6151
R18768 vdd.n1856 vdd.n1855 10.6151
R18769 vdd.n1855 vdd.n1853 10.6151
R18770 vdd.n1853 vdd.n1852 10.6151
R18771 vdd.n1852 vdd.n758 10.6151
R18772 vdd.n2074 vdd.n758 10.6151
R18773 vdd.n2075 vdd.n2074 10.6151
R18774 vdd.n1986 vdd.n1985 10.6151
R18775 vdd.n1985 vdd.n843 10.6151
R18776 vdd.n1979 vdd.n843 10.6151
R18777 vdd.n1979 vdd.n1978 10.6151
R18778 vdd.n1978 vdd.n1977 10.6151
R18779 vdd.n1977 vdd.n845 10.6151
R18780 vdd.n1971 vdd.n845 10.6151
R18781 vdd.n1971 vdd.n1970 10.6151
R18782 vdd.n1970 vdd.n1969 10.6151
R18783 vdd.n1969 vdd.n847 10.6151
R18784 vdd.n1963 vdd.n847 10.6151
R18785 vdd.n1963 vdd.n1962 10.6151
R18786 vdd.n1962 vdd.n1961 10.6151
R18787 vdd.n1961 vdd.n849 10.6151
R18788 vdd.n1955 vdd.n849 10.6151
R18789 vdd.n1955 vdd.n1954 10.6151
R18790 vdd.n1954 vdd.n1953 10.6151
R18791 vdd.n1953 vdd.n853 10.6151
R18792 vdd.n1801 vdd.n853 10.6151
R18793 vdd.n1802 vdd.n1801 10.6151
R18794 vdd.n1802 vdd.n1797 10.6151
R18795 vdd.n1808 vdd.n1797 10.6151
R18796 vdd.n1809 vdd.n1808 10.6151
R18797 vdd.n1810 vdd.n1809 10.6151
R18798 vdd.n1810 vdd.n1795 10.6151
R18799 vdd.n1816 vdd.n1795 10.6151
R18800 vdd.n1817 vdd.n1816 10.6151
R18801 vdd.n1818 vdd.n1817 10.6151
R18802 vdd.n1818 vdd.n1793 10.6151
R18803 vdd.n1824 vdd.n1793 10.6151
R18804 vdd.n1825 vdd.n1824 10.6151
R18805 vdd.n1827 vdd.n1789 10.6151
R18806 vdd.n1832 vdd.n1789 10.6151
R18807 vdd.n280 vdd.n262 10.4732
R18808 vdd.n233 vdd.n215 10.4732
R18809 vdd.n190 vdd.n172 10.4732
R18810 vdd.n143 vdd.n125 10.4732
R18811 vdd.n101 vdd.n83 10.4732
R18812 vdd.n54 vdd.n36 10.4732
R18813 vdd.n1095 vdd.n1077 10.4732
R18814 vdd.n1142 vdd.n1124 10.4732
R18815 vdd.n1005 vdd.n987 10.4732
R18816 vdd.n1052 vdd.n1034 10.4732
R18817 vdd.n916 vdd.n898 10.4732
R18818 vdd.n963 vdd.n945 10.4732
R18819 vdd.t31 vdd.n888 10.3167
R18820 vdd.n2874 vdd.t51 10.3167
R18821 vdd.n1465 vdd.t27 10.09
R18822 vdd.n3042 vdd.t64 10.09
R18823 vdd.n279 vdd.n264 9.69747
R18824 vdd.n232 vdd.n217 9.69747
R18825 vdd.n189 vdd.n174 9.69747
R18826 vdd.n142 vdd.n127 9.69747
R18827 vdd.n100 vdd.n85 9.69747
R18828 vdd.n53 vdd.n38 9.69747
R18829 vdd.n1094 vdd.n1079 9.69747
R18830 vdd.n1141 vdd.n1126 9.69747
R18831 vdd.n1004 vdd.n989 9.69747
R18832 vdd.n1051 vdd.n1036 9.69747
R18833 vdd.n915 vdd.n900 9.69747
R18834 vdd.n962 vdd.n947 9.69747
R18835 vdd.n1929 vdd.n1928 9.67831
R18836 vdd.n2836 vdd.n520 9.67831
R18837 vdd.n2707 vdd.n2706 9.67831
R18838 vdd.n1953 vdd.n1952 9.67831
R18839 vdd.n295 vdd.n294 9.45567
R18840 vdd.n248 vdd.n247 9.45567
R18841 vdd.n205 vdd.n204 9.45567
R18842 vdd.n158 vdd.n157 9.45567
R18843 vdd.n116 vdd.n115 9.45567
R18844 vdd.n69 vdd.n68 9.45567
R18845 vdd.n1110 vdd.n1109 9.45567
R18846 vdd.n1157 vdd.n1156 9.45567
R18847 vdd.n1020 vdd.n1019 9.45567
R18848 vdd.n1067 vdd.n1066 9.45567
R18849 vdd.n931 vdd.n930 9.45567
R18850 vdd.n978 vdd.n977 9.45567
R18851 vdd.n1689 vdd.n1543 9.3005
R18852 vdd.n1688 vdd.n1687 9.3005
R18853 vdd.n1549 vdd.n1548 9.3005
R18854 vdd.n1682 vdd.n1553 9.3005
R18855 vdd.n1681 vdd.n1554 9.3005
R18856 vdd.n1680 vdd.n1555 9.3005
R18857 vdd.n1559 vdd.n1556 9.3005
R18858 vdd.n1675 vdd.n1560 9.3005
R18859 vdd.n1674 vdd.n1561 9.3005
R18860 vdd.n1673 vdd.n1562 9.3005
R18861 vdd.n1566 vdd.n1563 9.3005
R18862 vdd.n1668 vdd.n1567 9.3005
R18863 vdd.n1667 vdd.n1568 9.3005
R18864 vdd.n1666 vdd.n1569 9.3005
R18865 vdd.n1573 vdd.n1570 9.3005
R18866 vdd.n1661 vdd.n1574 9.3005
R18867 vdd.n1660 vdd.n1575 9.3005
R18868 vdd.n1659 vdd.n1576 9.3005
R18869 vdd.n1580 vdd.n1577 9.3005
R18870 vdd.n1654 vdd.n1581 9.3005
R18871 vdd.n1653 vdd.n1582 9.3005
R18872 vdd.n1652 vdd.n1651 9.3005
R18873 vdd.n1650 vdd.n1583 9.3005
R18874 vdd.n1649 vdd.n1648 9.3005
R18875 vdd.n1589 vdd.n1588 9.3005
R18876 vdd.n1643 vdd.n1593 9.3005
R18877 vdd.n1642 vdd.n1594 9.3005
R18878 vdd.n1641 vdd.n1595 9.3005
R18879 vdd.n1599 vdd.n1596 9.3005
R18880 vdd.n1636 vdd.n1600 9.3005
R18881 vdd.n1635 vdd.n1601 9.3005
R18882 vdd.n1634 vdd.n1602 9.3005
R18883 vdd.n1606 vdd.n1603 9.3005
R18884 vdd.n1629 vdd.n1607 9.3005
R18885 vdd.n1628 vdd.n1608 9.3005
R18886 vdd.n1627 vdd.n1609 9.3005
R18887 vdd.n1611 vdd.n1610 9.3005
R18888 vdd.n1622 vdd.n854 9.3005
R18889 vdd.n1691 vdd.n1690 9.3005
R18890 vdd.n1715 vdd.n1714 9.3005
R18891 vdd.n1521 vdd.n1520 9.3005
R18892 vdd.n1526 vdd.n1524 9.3005
R18893 vdd.n1707 vdd.n1527 9.3005
R18894 vdd.n1706 vdd.n1528 9.3005
R18895 vdd.n1705 vdd.n1529 9.3005
R18896 vdd.n1533 vdd.n1530 9.3005
R18897 vdd.n1700 vdd.n1534 9.3005
R18898 vdd.n1699 vdd.n1535 9.3005
R18899 vdd.n1698 vdd.n1536 9.3005
R18900 vdd.n1540 vdd.n1537 9.3005
R18901 vdd.n1693 vdd.n1541 9.3005
R18902 vdd.n1692 vdd.n1542 9.3005
R18903 vdd.n1937 vdd.n1514 9.3005
R18904 vdd.n1939 vdd.n1938 9.3005
R18905 vdd.n1476 vdd.n1475 9.3005
R18906 vdd.n1477 vdd.n890 9.3005
R18907 vdd.n1479 vdd.n1478 9.3005
R18908 vdd.n880 vdd.n879 9.3005
R18909 vdd.n1493 vdd.n1492 9.3005
R18910 vdd.n1494 vdd.n878 9.3005
R18911 vdd.n1496 vdd.n1495 9.3005
R18912 vdd.n868 vdd.n867 9.3005
R18913 vdd.n1512 vdd.n1511 9.3005
R18914 vdd.n1513 vdd.n866 9.3005
R18915 vdd.n1941 vdd.n1940 9.3005
R18916 vdd.n271 vdd.n270 9.3005
R18917 vdd.n266 vdd.n265 9.3005
R18918 vdd.n277 vdd.n276 9.3005
R18919 vdd.n279 vdd.n278 9.3005
R18920 vdd.n262 vdd.n261 9.3005
R18921 vdd.n285 vdd.n284 9.3005
R18922 vdd.n287 vdd.n286 9.3005
R18923 vdd.n259 vdd.n256 9.3005
R18924 vdd.n294 vdd.n293 9.3005
R18925 vdd.n224 vdd.n223 9.3005
R18926 vdd.n219 vdd.n218 9.3005
R18927 vdd.n230 vdd.n229 9.3005
R18928 vdd.n232 vdd.n231 9.3005
R18929 vdd.n215 vdd.n214 9.3005
R18930 vdd.n238 vdd.n237 9.3005
R18931 vdd.n240 vdd.n239 9.3005
R18932 vdd.n212 vdd.n209 9.3005
R18933 vdd.n247 vdd.n246 9.3005
R18934 vdd.n181 vdd.n180 9.3005
R18935 vdd.n176 vdd.n175 9.3005
R18936 vdd.n187 vdd.n186 9.3005
R18937 vdd.n189 vdd.n188 9.3005
R18938 vdd.n172 vdd.n171 9.3005
R18939 vdd.n195 vdd.n194 9.3005
R18940 vdd.n197 vdd.n196 9.3005
R18941 vdd.n169 vdd.n166 9.3005
R18942 vdd.n204 vdd.n203 9.3005
R18943 vdd.n134 vdd.n133 9.3005
R18944 vdd.n129 vdd.n128 9.3005
R18945 vdd.n140 vdd.n139 9.3005
R18946 vdd.n142 vdd.n141 9.3005
R18947 vdd.n125 vdd.n124 9.3005
R18948 vdd.n148 vdd.n147 9.3005
R18949 vdd.n150 vdd.n149 9.3005
R18950 vdd.n122 vdd.n119 9.3005
R18951 vdd.n157 vdd.n156 9.3005
R18952 vdd.n92 vdd.n91 9.3005
R18953 vdd.n87 vdd.n86 9.3005
R18954 vdd.n98 vdd.n97 9.3005
R18955 vdd.n100 vdd.n99 9.3005
R18956 vdd.n83 vdd.n82 9.3005
R18957 vdd.n106 vdd.n105 9.3005
R18958 vdd.n108 vdd.n107 9.3005
R18959 vdd.n80 vdd.n77 9.3005
R18960 vdd.n115 vdd.n114 9.3005
R18961 vdd.n45 vdd.n44 9.3005
R18962 vdd.n40 vdd.n39 9.3005
R18963 vdd.n51 vdd.n50 9.3005
R18964 vdd.n53 vdd.n52 9.3005
R18965 vdd.n36 vdd.n35 9.3005
R18966 vdd.n59 vdd.n58 9.3005
R18967 vdd.n61 vdd.n60 9.3005
R18968 vdd.n33 vdd.n30 9.3005
R18969 vdd.n68 vdd.n67 9.3005
R18970 vdd.n2758 vdd.n2757 9.3005
R18971 vdd.n2761 vdd.n555 9.3005
R18972 vdd.n2762 vdd.n554 9.3005
R18973 vdd.n2765 vdd.n553 9.3005
R18974 vdd.n2766 vdd.n552 9.3005
R18975 vdd.n2769 vdd.n551 9.3005
R18976 vdd.n2770 vdd.n550 9.3005
R18977 vdd.n2773 vdd.n549 9.3005
R18978 vdd.n2774 vdd.n548 9.3005
R18979 vdd.n2777 vdd.n547 9.3005
R18980 vdd.n2778 vdd.n546 9.3005
R18981 vdd.n2781 vdd.n545 9.3005
R18982 vdd.n2782 vdd.n544 9.3005
R18983 vdd.n2785 vdd.n543 9.3005
R18984 vdd.n2786 vdd.n542 9.3005
R18985 vdd.n2789 vdd.n541 9.3005
R18986 vdd.n2790 vdd.n540 9.3005
R18987 vdd.n2793 vdd.n539 9.3005
R18988 vdd.n2794 vdd.n538 9.3005
R18989 vdd.n2797 vdd.n537 9.3005
R18990 vdd.n2801 vdd.n2800 9.3005
R18991 vdd.n2802 vdd.n536 9.3005
R18992 vdd.n2806 vdd.n2803 9.3005
R18993 vdd.n2809 vdd.n535 9.3005
R18994 vdd.n2810 vdd.n534 9.3005
R18995 vdd.n2813 vdd.n533 9.3005
R18996 vdd.n2814 vdd.n532 9.3005
R18997 vdd.n2817 vdd.n531 9.3005
R18998 vdd.n2818 vdd.n530 9.3005
R18999 vdd.n2821 vdd.n529 9.3005
R19000 vdd.n2822 vdd.n528 9.3005
R19001 vdd.n2825 vdd.n527 9.3005
R19002 vdd.n2826 vdd.n526 9.3005
R19003 vdd.n2829 vdd.n525 9.3005
R19004 vdd.n2830 vdd.n524 9.3005
R19005 vdd.n2833 vdd.n519 9.3005
R19006 vdd.n482 vdd.n481 9.3005
R19007 vdd.n2844 vdd.n2843 9.3005
R19008 vdd.n2847 vdd.n2846 9.3005
R19009 vdd.n471 vdd.n470 9.3005
R19010 vdd.n2861 vdd.n2860 9.3005
R19011 vdd.n2862 vdd.n469 9.3005
R19012 vdd.n2864 vdd.n2863 9.3005
R19013 vdd.n460 vdd.n459 9.3005
R19014 vdd.n2877 vdd.n2876 9.3005
R19015 vdd.n2878 vdd.n458 9.3005
R19016 vdd.n2880 vdd.n2879 9.3005
R19017 vdd.n300 vdd.n298 9.3005
R19018 vdd.n2845 vdd.n480 9.3005
R19019 vdd.n3046 vdd.n3045 9.3005
R19020 vdd.n301 vdd.n299 9.3005
R19021 vdd.n3039 vdd.n310 9.3005
R19022 vdd.n3038 vdd.n311 9.3005
R19023 vdd.n3037 vdd.n312 9.3005
R19024 vdd.n320 vdd.n313 9.3005
R19025 vdd.n3031 vdd.n321 9.3005
R19026 vdd.n3030 vdd.n322 9.3005
R19027 vdd.n3029 vdd.n323 9.3005
R19028 vdd.n331 vdd.n324 9.3005
R19029 vdd.n3023 vdd.n3022 9.3005
R19030 vdd.n3019 vdd.n332 9.3005
R19031 vdd.n3018 vdd.n335 9.3005
R19032 vdd.n339 vdd.n336 9.3005
R19033 vdd.n340 vdd.n337 9.3005
R19034 vdd.n3011 vdd.n341 9.3005
R19035 vdd.n3010 vdd.n342 9.3005
R19036 vdd.n3009 vdd.n343 9.3005
R19037 vdd.n347 vdd.n344 9.3005
R19038 vdd.n3004 vdd.n348 9.3005
R19039 vdd.n3003 vdd.n349 9.3005
R19040 vdd.n3002 vdd.n350 9.3005
R19041 vdd.n354 vdd.n351 9.3005
R19042 vdd.n2997 vdd.n355 9.3005
R19043 vdd.n2996 vdd.n356 9.3005
R19044 vdd.n2995 vdd.n357 9.3005
R19045 vdd.n361 vdd.n358 9.3005
R19046 vdd.n2990 vdd.n362 9.3005
R19047 vdd.n2989 vdd.n363 9.3005
R19048 vdd.n2988 vdd.n2987 9.3005
R19049 vdd.n2986 vdd.n364 9.3005
R19050 vdd.n2985 vdd.n2984 9.3005
R19051 vdd.n370 vdd.n369 9.3005
R19052 vdd.n2979 vdd.n374 9.3005
R19053 vdd.n2978 vdd.n375 9.3005
R19054 vdd.n2977 vdd.n376 9.3005
R19055 vdd.n380 vdd.n377 9.3005
R19056 vdd.n2972 vdd.n381 9.3005
R19057 vdd.n2971 vdd.n382 9.3005
R19058 vdd.n2970 vdd.n383 9.3005
R19059 vdd.n387 vdd.n384 9.3005
R19060 vdd.n2965 vdd.n388 9.3005
R19061 vdd.n2964 vdd.n389 9.3005
R19062 vdd.n2963 vdd.n390 9.3005
R19063 vdd.n394 vdd.n391 9.3005
R19064 vdd.n2958 vdd.n395 9.3005
R19065 vdd.n2957 vdd.n396 9.3005
R19066 vdd.n2956 vdd.n397 9.3005
R19067 vdd.n401 vdd.n398 9.3005
R19068 vdd.n2951 vdd.n402 9.3005
R19069 vdd.n2950 vdd.n403 9.3005
R19070 vdd.n2949 vdd.n2948 9.3005
R19071 vdd.n2947 vdd.n404 9.3005
R19072 vdd.n2946 vdd.n2945 9.3005
R19073 vdd.n410 vdd.n409 9.3005
R19074 vdd.n2940 vdd.n414 9.3005
R19075 vdd.n2939 vdd.n415 9.3005
R19076 vdd.n2938 vdd.n416 9.3005
R19077 vdd.n420 vdd.n417 9.3005
R19078 vdd.n2933 vdd.n421 9.3005
R19079 vdd.n2932 vdd.n422 9.3005
R19080 vdd.n2931 vdd.n423 9.3005
R19081 vdd.n427 vdd.n424 9.3005
R19082 vdd.n2926 vdd.n428 9.3005
R19083 vdd.n2925 vdd.n429 9.3005
R19084 vdd.n2924 vdd.n430 9.3005
R19085 vdd.n434 vdd.n431 9.3005
R19086 vdd.n2919 vdd.n435 9.3005
R19087 vdd.n2918 vdd.n436 9.3005
R19088 vdd.n2917 vdd.n437 9.3005
R19089 vdd.n441 vdd.n438 9.3005
R19090 vdd.n2912 vdd.n442 9.3005
R19091 vdd.n2911 vdd.n443 9.3005
R19092 vdd.n2907 vdd.n2904 9.3005
R19093 vdd.n3021 vdd.n3020 9.3005
R19094 vdd.n2852 vdd.n2851 9.3005
R19095 vdd.n2853 vdd.n475 9.3005
R19096 vdd.n2855 vdd.n2854 9.3005
R19097 vdd.n465 vdd.n464 9.3005
R19098 vdd.n2869 vdd.n2868 9.3005
R19099 vdd.n2870 vdd.n463 9.3005
R19100 vdd.n2872 vdd.n2871 9.3005
R19101 vdd.n453 vdd.n452 9.3005
R19102 vdd.n2885 vdd.n2884 9.3005
R19103 vdd.n2886 vdd.n451 9.3005
R19104 vdd.n2888 vdd.n2887 9.3005
R19105 vdd.n2889 vdd.n450 9.3005
R19106 vdd.n2891 vdd.n2890 9.3005
R19107 vdd.n2892 vdd.n449 9.3005
R19108 vdd.n2894 vdd.n2893 9.3005
R19109 vdd.n2895 vdd.n447 9.3005
R19110 vdd.n2897 vdd.n2896 9.3005
R19111 vdd.n2898 vdd.n446 9.3005
R19112 vdd.n2900 vdd.n2899 9.3005
R19113 vdd.n2901 vdd.n444 9.3005
R19114 vdd.n2903 vdd.n2902 9.3005
R19115 vdd.n477 vdd.n476 9.3005
R19116 vdd.n2710 vdd.n2709 9.3005
R19117 vdd.n2715 vdd.n2708 9.3005
R19118 vdd.n2724 vdd.n572 9.3005
R19119 vdd.n2727 vdd.n571 9.3005
R19120 vdd.n2728 vdd.n570 9.3005
R19121 vdd.n2731 vdd.n569 9.3005
R19122 vdd.n2732 vdd.n568 9.3005
R19123 vdd.n2735 vdd.n567 9.3005
R19124 vdd.n2736 vdd.n566 9.3005
R19125 vdd.n2739 vdd.n565 9.3005
R19126 vdd.n2740 vdd.n564 9.3005
R19127 vdd.n2743 vdd.n563 9.3005
R19128 vdd.n2744 vdd.n562 9.3005
R19129 vdd.n2747 vdd.n561 9.3005
R19130 vdd.n2748 vdd.n560 9.3005
R19131 vdd.n2751 vdd.n559 9.3005
R19132 vdd.n2755 vdd.n2754 9.3005
R19133 vdd.n2756 vdd.n556 9.3005
R19134 vdd.n1951 vdd.n1950 9.3005
R19135 vdd.n1946 vdd.n857 9.3005
R19136 vdd.n1433 vdd.n1432 9.3005
R19137 vdd.n1434 vdd.n1188 9.3005
R19138 vdd.n1436 vdd.n1435 9.3005
R19139 vdd.n1178 vdd.n1177 9.3005
R19140 vdd.n1450 vdd.n1449 9.3005
R19141 vdd.n1451 vdd.n1176 9.3005
R19142 vdd.n1453 vdd.n1452 9.3005
R19143 vdd.n1168 vdd.n1167 9.3005
R19144 vdd.n1468 vdd.n1467 9.3005
R19145 vdd.n1469 vdd.n1166 9.3005
R19146 vdd.n1471 vdd.n1470 9.3005
R19147 vdd.n885 vdd.n884 9.3005
R19148 vdd.n1484 vdd.n1483 9.3005
R19149 vdd.n1485 vdd.n883 9.3005
R19150 vdd.n1487 vdd.n1486 9.3005
R19151 vdd.n875 vdd.n874 9.3005
R19152 vdd.n1501 vdd.n1500 9.3005
R19153 vdd.n1502 vdd.n872 9.3005
R19154 vdd.n1506 vdd.n1505 9.3005
R19155 vdd.n1504 vdd.n873 9.3005
R19156 vdd.n1503 vdd.n862 9.3005
R19157 vdd.n1190 vdd.n1189 9.3005
R19158 vdd.n1326 vdd.n1325 9.3005
R19159 vdd.n1327 vdd.n1316 9.3005
R19160 vdd.n1329 vdd.n1328 9.3005
R19161 vdd.n1330 vdd.n1315 9.3005
R19162 vdd.n1332 vdd.n1331 9.3005
R19163 vdd.n1333 vdd.n1310 9.3005
R19164 vdd.n1335 vdd.n1334 9.3005
R19165 vdd.n1336 vdd.n1309 9.3005
R19166 vdd.n1338 vdd.n1337 9.3005
R19167 vdd.n1339 vdd.n1304 9.3005
R19168 vdd.n1341 vdd.n1340 9.3005
R19169 vdd.n1342 vdd.n1303 9.3005
R19170 vdd.n1344 vdd.n1343 9.3005
R19171 vdd.n1345 vdd.n1298 9.3005
R19172 vdd.n1347 vdd.n1346 9.3005
R19173 vdd.n1348 vdd.n1297 9.3005
R19174 vdd.n1350 vdd.n1349 9.3005
R19175 vdd.n1351 vdd.n1292 9.3005
R19176 vdd.n1353 vdd.n1352 9.3005
R19177 vdd.n1354 vdd.n1291 9.3005
R19178 vdd.n1356 vdd.n1355 9.3005
R19179 vdd.n1360 vdd.n1287 9.3005
R19180 vdd.n1362 vdd.n1361 9.3005
R19181 vdd.n1363 vdd.n1286 9.3005
R19182 vdd.n1365 vdd.n1364 9.3005
R19183 vdd.n1366 vdd.n1281 9.3005
R19184 vdd.n1368 vdd.n1367 9.3005
R19185 vdd.n1369 vdd.n1280 9.3005
R19186 vdd.n1371 vdd.n1370 9.3005
R19187 vdd.n1372 vdd.n1275 9.3005
R19188 vdd.n1374 vdd.n1373 9.3005
R19189 vdd.n1375 vdd.n1274 9.3005
R19190 vdd.n1377 vdd.n1376 9.3005
R19191 vdd.n1378 vdd.n1269 9.3005
R19192 vdd.n1380 vdd.n1379 9.3005
R19193 vdd.n1381 vdd.n1268 9.3005
R19194 vdd.n1383 vdd.n1382 9.3005
R19195 vdd.n1384 vdd.n1263 9.3005
R19196 vdd.n1386 vdd.n1385 9.3005
R19197 vdd.n1387 vdd.n1262 9.3005
R19198 vdd.n1389 vdd.n1388 9.3005
R19199 vdd.n1390 vdd.n1257 9.3005
R19200 vdd.n1392 vdd.n1391 9.3005
R19201 vdd.n1393 vdd.n1256 9.3005
R19202 vdd.n1395 vdd.n1394 9.3005
R19203 vdd.n1396 vdd.n1249 9.3005
R19204 vdd.n1398 vdd.n1397 9.3005
R19205 vdd.n1399 vdd.n1248 9.3005
R19206 vdd.n1401 vdd.n1400 9.3005
R19207 vdd.n1402 vdd.n1243 9.3005
R19208 vdd.n1404 vdd.n1403 9.3005
R19209 vdd.n1405 vdd.n1242 9.3005
R19210 vdd.n1407 vdd.n1406 9.3005
R19211 vdd.n1408 vdd.n1237 9.3005
R19212 vdd.n1410 vdd.n1409 9.3005
R19213 vdd.n1411 vdd.n1236 9.3005
R19214 vdd.n1413 vdd.n1412 9.3005
R19215 vdd.n1414 vdd.n1231 9.3005
R19216 vdd.n1416 vdd.n1415 9.3005
R19217 vdd.n1417 vdd.n1230 9.3005
R19218 vdd.n1419 vdd.n1418 9.3005
R19219 vdd.n1195 vdd.n1194 9.3005
R19220 vdd.n1425 vdd.n1424 9.3005
R19221 vdd.n1324 vdd.n1323 9.3005
R19222 vdd.n1428 vdd.n1427 9.3005
R19223 vdd.n1184 vdd.n1183 9.3005
R19224 vdd.n1442 vdd.n1441 9.3005
R19225 vdd.n1443 vdd.n1182 9.3005
R19226 vdd.n1445 vdd.n1444 9.3005
R19227 vdd.n1173 vdd.n1172 9.3005
R19228 vdd.n1459 vdd.n1458 9.3005
R19229 vdd.n1460 vdd.n1171 9.3005
R19230 vdd.n1463 vdd.n1462 9.3005
R19231 vdd.n1461 vdd.n1162 9.3005
R19232 vdd.n1426 vdd.n1193 9.3005
R19233 vdd.n1086 vdd.n1085 9.3005
R19234 vdd.n1081 vdd.n1080 9.3005
R19235 vdd.n1092 vdd.n1091 9.3005
R19236 vdd.n1094 vdd.n1093 9.3005
R19237 vdd.n1077 vdd.n1076 9.3005
R19238 vdd.n1100 vdd.n1099 9.3005
R19239 vdd.n1102 vdd.n1101 9.3005
R19240 vdd.n1074 vdd.n1071 9.3005
R19241 vdd.n1109 vdd.n1108 9.3005
R19242 vdd.n1133 vdd.n1132 9.3005
R19243 vdd.n1128 vdd.n1127 9.3005
R19244 vdd.n1139 vdd.n1138 9.3005
R19245 vdd.n1141 vdd.n1140 9.3005
R19246 vdd.n1124 vdd.n1123 9.3005
R19247 vdd.n1147 vdd.n1146 9.3005
R19248 vdd.n1149 vdd.n1148 9.3005
R19249 vdd.n1121 vdd.n1118 9.3005
R19250 vdd.n1156 vdd.n1155 9.3005
R19251 vdd.n996 vdd.n995 9.3005
R19252 vdd.n991 vdd.n990 9.3005
R19253 vdd.n1002 vdd.n1001 9.3005
R19254 vdd.n1004 vdd.n1003 9.3005
R19255 vdd.n987 vdd.n986 9.3005
R19256 vdd.n1010 vdd.n1009 9.3005
R19257 vdd.n1012 vdd.n1011 9.3005
R19258 vdd.n984 vdd.n981 9.3005
R19259 vdd.n1019 vdd.n1018 9.3005
R19260 vdd.n1043 vdd.n1042 9.3005
R19261 vdd.n1038 vdd.n1037 9.3005
R19262 vdd.n1049 vdd.n1048 9.3005
R19263 vdd.n1051 vdd.n1050 9.3005
R19264 vdd.n1034 vdd.n1033 9.3005
R19265 vdd.n1057 vdd.n1056 9.3005
R19266 vdd.n1059 vdd.n1058 9.3005
R19267 vdd.n1031 vdd.n1028 9.3005
R19268 vdd.n1066 vdd.n1065 9.3005
R19269 vdd.n907 vdd.n906 9.3005
R19270 vdd.n902 vdd.n901 9.3005
R19271 vdd.n913 vdd.n912 9.3005
R19272 vdd.n915 vdd.n914 9.3005
R19273 vdd.n898 vdd.n897 9.3005
R19274 vdd.n921 vdd.n920 9.3005
R19275 vdd.n923 vdd.n922 9.3005
R19276 vdd.n895 vdd.n892 9.3005
R19277 vdd.n930 vdd.n929 9.3005
R19278 vdd.n954 vdd.n953 9.3005
R19279 vdd.n949 vdd.n948 9.3005
R19280 vdd.n960 vdd.n959 9.3005
R19281 vdd.n962 vdd.n961 9.3005
R19282 vdd.n945 vdd.n944 9.3005
R19283 vdd.n968 vdd.n967 9.3005
R19284 vdd.n970 vdd.n969 9.3005
R19285 vdd.n942 vdd.n939 9.3005
R19286 vdd.n977 vdd.n976 9.3005
R19287 vdd.n1438 vdd.t60 8.95635
R19288 vdd.t42 vdd.n3033 8.95635
R19289 vdd.n276 vdd.n275 8.92171
R19290 vdd.n229 vdd.n228 8.92171
R19291 vdd.n186 vdd.n185 8.92171
R19292 vdd.n139 vdd.n138 8.92171
R19293 vdd.n97 vdd.n96 8.92171
R19294 vdd.n50 vdd.n49 8.92171
R19295 vdd.n1091 vdd.n1090 8.92171
R19296 vdd.n1138 vdd.n1137 8.92171
R19297 vdd.n1001 vdd.n1000 8.92171
R19298 vdd.n1048 vdd.n1047 8.92171
R19299 vdd.n912 vdd.n911 8.92171
R19300 vdd.n959 vdd.n958 8.92171
R19301 vdd.n207 vdd.n117 8.81535
R19302 vdd.n1069 vdd.n979 8.81535
R19303 vdd.n1465 vdd.t38 8.72962
R19304 vdd.t40 vdd.n3042 8.72962
R19305 vdd.n888 vdd.t76 8.50289
R19306 vdd.n1943 vdd.t132 8.50289
R19307 vdd.n516 vdd.t125 8.50289
R19308 vdd.n2874 vdd.t54 8.50289
R19309 vdd.n28 vdd.n14 8.42249
R19310 vdd.n3048 vdd.n3047 8.16225
R19311 vdd.n1161 vdd.n1160 8.16225
R19312 vdd.n272 vdd.n266 8.14595
R19313 vdd.n225 vdd.n219 8.14595
R19314 vdd.n182 vdd.n176 8.14595
R19315 vdd.n135 vdd.n129 8.14595
R19316 vdd.n93 vdd.n87 8.14595
R19317 vdd.n46 vdd.n40 8.14595
R19318 vdd.n1087 vdd.n1081 8.14595
R19319 vdd.n1134 vdd.n1128 8.14595
R19320 vdd.n997 vdd.n991 8.14595
R19321 vdd.n1044 vdd.n1038 8.14595
R19322 vdd.n908 vdd.n902 8.14595
R19323 vdd.n955 vdd.n949 8.14595
R19324 vdd.n2537 vdd.n639 8.11757
R19325 vdd.n2011 vdd.n2010 8.11757
R19326 vdd.n1989 vdd.n833 7.70933
R19327 vdd.n1995 vdd.n833 7.70933
R19328 vdd.n2001 vdd.n827 7.70933
R19329 vdd.n2001 vdd.n820 7.70933
R19330 vdd.n2007 vdd.n820 7.70933
R19331 vdd.n2007 vdd.n823 7.70933
R19332 vdd.n2014 vdd.n808 7.70933
R19333 vdd.n2020 vdd.n808 7.70933
R19334 vdd.n2026 vdd.n802 7.70933
R19335 vdd.n2032 vdd.n798 7.70933
R19336 vdd.n2038 vdd.n792 7.70933
R19337 vdd.n2050 vdd.n779 7.70933
R19338 vdd.n2056 vdd.n773 7.70933
R19339 vdd.n2056 vdd.n766 7.70933
R19340 vdd.n2064 vdd.n766 7.70933
R19341 vdd.n2071 vdd.t2 7.70933
R19342 vdd.n2146 vdd.t2 7.70933
R19343 vdd.n2478 vdd.t21 7.70933
R19344 vdd.n2484 vdd.t21 7.70933
R19345 vdd.n2490 vdd.n687 7.70933
R19346 vdd.n2496 vdd.n687 7.70933
R19347 vdd.n2496 vdd.n690 7.70933
R19348 vdd.n2502 vdd.n683 7.70933
R19349 vdd.n2514 vdd.n670 7.70933
R19350 vdd.n2520 vdd.n664 7.70933
R19351 vdd.n2526 vdd.n660 7.70933
R19352 vdd.n2532 vdd.n647 7.70933
R19353 vdd.n2540 vdd.n647 7.70933
R19354 vdd.n2546 vdd.n641 7.70933
R19355 vdd.n2546 vdd.n633 7.70933
R19356 vdd.n2597 vdd.n633 7.70933
R19357 vdd.n2597 vdd.n636 7.70933
R19358 vdd.n2603 vdd.n595 7.70933
R19359 vdd.n2673 vdd.n595 7.70933
R19360 vdd.n271 vdd.n268 7.3702
R19361 vdd.n224 vdd.n221 7.3702
R19362 vdd.n181 vdd.n178 7.3702
R19363 vdd.n134 vdd.n131 7.3702
R19364 vdd.n92 vdd.n89 7.3702
R19365 vdd.n45 vdd.n42 7.3702
R19366 vdd.n1086 vdd.n1083 7.3702
R19367 vdd.n1133 vdd.n1130 7.3702
R19368 vdd.n996 vdd.n993 7.3702
R19369 vdd.n1043 vdd.n1040 7.3702
R19370 vdd.n907 vdd.n904 7.3702
R19371 vdd.n954 vdd.n951 7.3702
R19372 vdd.n1361 vdd.n1360 6.98232
R19373 vdd.n1653 vdd.n1652 6.98232
R19374 vdd.n2950 vdd.n2949 6.98232
R19375 vdd.n2761 vdd.n2758 6.98232
R19376 vdd.n1498 vdd.t23 6.68904
R19377 vdd.n2857 vdd.t25 6.68904
R19378 vdd.t62 vdd.n887 6.46231
R19379 vdd.n2882 vdd.t29 6.46231
R19380 vdd.n1456 vdd.t44 6.23558
R19381 vdd.t33 vdd.n308 6.23558
R19382 vdd.n3048 vdd.n297 6.22547
R19383 vdd.n1160 vdd.n1159 6.22547
R19384 vdd.n2026 vdd.t87 6.00885
R19385 vdd.n2526 vdd.t20 6.00885
R19386 vdd.n823 vdd.t176 5.89549
R19387 vdd.t140 vdd.n641 5.89549
R19388 vdd.n272 vdd.n271 5.81868
R19389 vdd.n225 vdd.n224 5.81868
R19390 vdd.n182 vdd.n181 5.81868
R19391 vdd.n135 vdd.n134 5.81868
R19392 vdd.n93 vdd.n92 5.81868
R19393 vdd.n46 vdd.n45 5.81868
R19394 vdd.n1087 vdd.n1086 5.81868
R19395 vdd.n1134 vdd.n1133 5.81868
R19396 vdd.n997 vdd.n996 5.81868
R19397 vdd.n1044 vdd.n1043 5.81868
R19398 vdd.n908 vdd.n907 5.81868
R19399 vdd.n955 vdd.n954 5.81868
R19400 vdd.t172 vdd.n827 5.78212
R19401 vdd.n1770 vdd.t157 5.78212
R19402 vdd.n2395 vdd.t165 5.78212
R19403 vdd.n636 vdd.t161 5.78212
R19404 vdd.n2154 vdd.n2153 5.77611
R19405 vdd.n1897 vdd.n1767 5.77611
R19406 vdd.n2408 vdd.n2407 5.77611
R19407 vdd.n2614 vdd.n2613 5.77611
R19408 vdd.n2678 vdd.n591 5.77611
R19409 vdd.n2318 vdd.n2258 5.77611
R19410 vdd.n2079 vdd.n757 5.77611
R19411 vdd.n1827 vdd.n1826 5.77611
R19412 vdd.n1323 vdd.n1322 5.62474
R19413 vdd.n1949 vdd.n1946 5.62474
R19414 vdd.n2910 vdd.n2907 5.62474
R19415 vdd.n2713 vdd.n2710 5.62474
R19416 vdd.t106 vdd.n779 5.44203
R19417 vdd.n683 vdd.t4 5.44203
R19418 vdd.n1180 vdd.t44 5.10193
R19419 vdd.t12 vdd.n802 5.10193
R19420 vdd.n792 vdd.t121 5.10193
R19421 vdd.t108 vdd.n670 5.10193
R19422 vdd.n660 vdd.t120 5.10193
R19423 vdd.n3035 vdd.t33 5.10193
R19424 vdd.n275 vdd.n266 5.04292
R19425 vdd.n228 vdd.n219 5.04292
R19426 vdd.n185 vdd.n176 5.04292
R19427 vdd.n138 vdd.n129 5.04292
R19428 vdd.n96 vdd.n87 5.04292
R19429 vdd.n49 vdd.n40 5.04292
R19430 vdd.n1090 vdd.n1081 5.04292
R19431 vdd.n1137 vdd.n1128 5.04292
R19432 vdd.n1000 vdd.n991 5.04292
R19433 vdd.n1047 vdd.n1038 5.04292
R19434 vdd.n911 vdd.n902 5.04292
R19435 vdd.n958 vdd.n949 5.04292
R19436 vdd.n1473 vdd.t62 4.8752
R19437 vdd.t105 vdd.t15 4.8752
R19438 vdd.t6 vdd.t116 4.8752
R19439 vdd.t0 vdd.t9 4.8752
R19440 vdd.t109 vdd.t88 4.8752
R19441 vdd.t29 vdd.n304 4.8752
R19442 vdd.n2155 vdd.n2154 4.83952
R19443 vdd.n1767 vdd.n1763 4.83952
R19444 vdd.n2409 vdd.n2408 4.83952
R19445 vdd.n2615 vdd.n2614 4.83952
R19446 vdd.n591 vdd.n586 4.83952
R19447 vdd.n2315 vdd.n2258 4.83952
R19448 vdd.n2082 vdd.n757 4.83952
R19449 vdd.n1826 vdd.n1825 4.83952
R19450 vdd.n1621 vdd.n855 4.74817
R19451 vdd.n1616 vdd.n856 4.74817
R19452 vdd.n1518 vdd.n1515 4.74817
R19453 vdd.n1930 vdd.n1519 4.74817
R19454 vdd.n1932 vdd.n1518 4.74817
R19455 vdd.n1931 vdd.n1930 4.74817
R19456 vdd.n2838 vdd.n2837 4.74817
R19457 vdd.n2835 vdd.n2834 4.74817
R19458 vdd.n2835 vdd.n521 4.74817
R19459 vdd.n2837 vdd.n518 4.74817
R19460 vdd.n2720 vdd.n573 4.74817
R19461 vdd.n2716 vdd.n574 4.74817
R19462 vdd.n2719 vdd.n574 4.74817
R19463 vdd.n2723 vdd.n573 4.74817
R19464 vdd.n1617 vdd.n855 4.74817
R19465 vdd.n858 vdd.n856 4.74817
R19466 vdd.n297 vdd.n296 4.7074
R19467 vdd.n207 vdd.n206 4.7074
R19468 vdd.n1159 vdd.n1158 4.7074
R19469 vdd.n1069 vdd.n1068 4.7074
R19470 vdd.n1489 vdd.t23 4.64847
R19471 vdd.n2866 vdd.t25 4.64847
R19472 vdd.n2032 vdd.t113 4.53511
R19473 vdd.n2520 vdd.t17 4.53511
R19474 vdd.n2064 vdd.t7 4.30838
R19475 vdd.n2490 vdd.t10 4.30838
R19476 vdd.n276 vdd.n264 4.26717
R19477 vdd.n229 vdd.n217 4.26717
R19478 vdd.n186 vdd.n174 4.26717
R19479 vdd.n139 vdd.n127 4.26717
R19480 vdd.n97 vdd.n85 4.26717
R19481 vdd.n50 vdd.n38 4.26717
R19482 vdd.n1091 vdd.n1079 4.26717
R19483 vdd.n1138 vdd.n1126 4.26717
R19484 vdd.n1001 vdd.n989 4.26717
R19485 vdd.n1048 vdd.n1036 4.26717
R19486 vdd.n912 vdd.n900 4.26717
R19487 vdd.n959 vdd.n947 4.26717
R19488 vdd.n297 vdd.n207 4.10845
R19489 vdd.n1159 vdd.n1069 4.10845
R19490 vdd.n253 vdd.t70 4.06363
R19491 vdd.n253 vdd.t34 4.06363
R19492 vdd.n251 vdd.t36 4.06363
R19493 vdd.n251 vdd.t57 4.06363
R19494 vdd.n249 vdd.t59 4.06363
R19495 vdd.n249 vdd.t75 4.06363
R19496 vdd.n163 vdd.t65 4.06363
R19497 vdd.n163 vdd.t86 4.06363
R19498 vdd.n161 vdd.t30 4.06363
R19499 vdd.n161 vdd.t49 4.06363
R19500 vdd.n159 vdd.t55 4.06363
R19501 vdd.n159 vdd.t66 4.06363
R19502 vdd.n74 vdd.t71 4.06363
R19503 vdd.n74 vdd.t46 4.06363
R19504 vdd.n72 vdd.t85 4.06363
R19505 vdd.n72 vdd.t41 4.06363
R19506 vdd.n70 vdd.t78 4.06363
R19507 vdd.n70 vdd.t52 4.06363
R19508 vdd.n1111 vdd.t37 4.06363
R19509 vdd.n1111 vdd.t81 4.06363
R19510 vdd.n1113 vdd.t80 4.06363
R19511 vdd.n1113 vdd.t69 4.06363
R19512 vdd.n1115 vdd.t56 4.06363
R19513 vdd.n1115 vdd.t35 4.06363
R19514 vdd.n1021 vdd.t32 4.06363
R19515 vdd.n1021 vdd.t77 4.06363
R19516 vdd.n1023 vdd.t72 4.06363
R19517 vdd.n1023 vdd.t63 4.06363
R19518 vdd.n1025 vdd.t48 4.06363
R19519 vdd.n1025 vdd.t28 4.06363
R19520 vdd.n932 vdd.t50 4.06363
R19521 vdd.n932 vdd.t79 4.06363
R19522 vdd.n934 vdd.t39 4.06363
R19523 vdd.n934 vdd.t67 4.06363
R19524 vdd.n936 vdd.t45 4.06363
R19525 vdd.n936 vdd.t73 4.06363
R19526 vdd.n26 vdd.t98 3.9605
R19527 vdd.n26 vdd.t103 3.9605
R19528 vdd.n23 vdd.t93 3.9605
R19529 vdd.n23 vdd.t89 3.9605
R19530 vdd.n21 vdd.t92 3.9605
R19531 vdd.n21 vdd.t95 3.9605
R19532 vdd.n20 vdd.t101 3.9605
R19533 vdd.n20 vdd.t97 3.9605
R19534 vdd.n15 vdd.t99 3.9605
R19535 vdd.n15 vdd.t96 3.9605
R19536 vdd.n16 vdd.t102 3.9605
R19537 vdd.n16 vdd.t91 3.9605
R19538 vdd.n18 vdd.t90 3.9605
R19539 vdd.n18 vdd.t104 3.9605
R19540 vdd.n25 vdd.t100 3.9605
R19541 vdd.n25 vdd.t94 3.9605
R19542 vdd.n7 vdd.t110 3.61217
R19543 vdd.n7 vdd.t18 3.61217
R19544 vdd.n8 vdd.t1 3.61217
R19545 vdd.n8 vdd.t5 3.61217
R19546 vdd.n10 vdd.t22 3.61217
R19547 vdd.n10 vdd.t11 3.61217
R19548 vdd.n12 vdd.t119 3.61217
R19549 vdd.n12 vdd.t14 3.61217
R19550 vdd.n5 vdd.t123 3.61217
R19551 vdd.n5 vdd.t112 3.61217
R19552 vdd.n3 vdd.t8 3.61217
R19553 vdd.n3 vdd.t3 3.61217
R19554 vdd.n1 vdd.t107 3.61217
R19555 vdd.n1 vdd.t117 3.61217
R19556 vdd.n0 vdd.t114 3.61217
R19557 vdd.n0 vdd.t16 3.61217
R19558 vdd.n280 vdd.n279 3.49141
R19559 vdd.n233 vdd.n232 3.49141
R19560 vdd.n190 vdd.n189 3.49141
R19561 vdd.n143 vdd.n142 3.49141
R19562 vdd.n101 vdd.n100 3.49141
R19563 vdd.n54 vdd.n53 3.49141
R19564 vdd.n1095 vdd.n1094 3.49141
R19565 vdd.n1142 vdd.n1141 3.49141
R19566 vdd.n1005 vdd.n1004 3.49141
R19567 vdd.n1052 vdd.n1051 3.49141
R19568 vdd.n916 vdd.n915 3.49141
R19569 vdd.n963 vdd.n962 3.49141
R19570 vdd.n1770 vdd.t7 3.40145
R19571 vdd.n2218 vdd.t122 3.40145
R19572 vdd.n2471 vdd.t13 3.40145
R19573 vdd.n2395 vdd.t10 3.40145
R19574 vdd.n1871 vdd.t113 3.17472
R19575 vdd.n2374 vdd.t17 3.17472
R19576 vdd.n1490 vdd.t76 2.83463
R19577 vdd.n1508 vdd.t132 2.83463
R19578 vdd.n2849 vdd.t125 2.83463
R19579 vdd.n467 vdd.t54 2.83463
R19580 vdd.n283 vdd.n262 2.71565
R19581 vdd.n236 vdd.n215 2.71565
R19582 vdd.n193 vdd.n172 2.71565
R19583 vdd.n146 vdd.n125 2.71565
R19584 vdd.n104 vdd.n83 2.71565
R19585 vdd.n57 vdd.n36 2.71565
R19586 vdd.n1098 vdd.n1077 2.71565
R19587 vdd.n1145 vdd.n1124 2.71565
R19588 vdd.n1008 vdd.n987 2.71565
R19589 vdd.n1055 vdd.n1034 2.71565
R19590 vdd.n919 vdd.n898 2.71565
R19591 vdd.n966 vdd.n945 2.71565
R19592 vdd.t38 vdd.n1164 2.6079
R19593 vdd.n2020 vdd.t12 2.6079
R19594 vdd.n2044 vdd.t121 2.6079
R19595 vdd.n2508 vdd.t108 2.6079
R19596 vdd.n2532 vdd.t120 2.6079
R19597 vdd.n3043 vdd.t40 2.6079
R19598 vdd.n2538 vdd.n2537 2.49806
R19599 vdd.n2012 vdd.n2011 2.49806
R19600 vdd.n270 vdd.n269 2.4129
R19601 vdd.n223 vdd.n222 2.4129
R19602 vdd.n180 vdd.n179 2.4129
R19603 vdd.n133 vdd.n132 2.4129
R19604 vdd.n91 vdd.n90 2.4129
R19605 vdd.n44 vdd.n43 2.4129
R19606 vdd.n1085 vdd.n1084 2.4129
R19607 vdd.n1132 vdd.n1131 2.4129
R19608 vdd.n995 vdd.n994 2.4129
R19609 vdd.n1042 vdd.n1041 2.4129
R19610 vdd.n906 vdd.n905 2.4129
R19611 vdd.n953 vdd.n952 2.4129
R19612 vdd.n1447 vdd.t60 2.38117
R19613 vdd.n3034 vdd.t42 2.38117
R19614 vdd.n1929 vdd.n1518 2.27742
R19615 vdd.n1930 vdd.n1929 2.27742
R19616 vdd.n2836 vdd.n2835 2.27742
R19617 vdd.n2837 vdd.n2836 2.27742
R19618 vdd.n2707 vdd.n574 2.27742
R19619 vdd.n2707 vdd.n573 2.27742
R19620 vdd.n1952 vdd.n855 2.27742
R19621 vdd.n1952 vdd.n856 2.27742
R19622 vdd.n2044 vdd.t106 2.2678
R19623 vdd.n2508 vdd.t4 2.2678
R19624 vdd.t116 vdd.n773 2.04107
R19625 vdd.n690 vdd.t0 2.04107
R19626 vdd.n284 vdd.n260 1.93989
R19627 vdd.n237 vdd.n213 1.93989
R19628 vdd.n194 vdd.n170 1.93989
R19629 vdd.n147 vdd.n123 1.93989
R19630 vdd.n105 vdd.n81 1.93989
R19631 vdd.n58 vdd.n34 1.93989
R19632 vdd.n1099 vdd.n1075 1.93989
R19633 vdd.n1146 vdd.n1122 1.93989
R19634 vdd.n1009 vdd.n985 1.93989
R19635 vdd.n1056 vdd.n1032 1.93989
R19636 vdd.n920 vdd.n896 1.93989
R19637 vdd.n967 vdd.n943 1.93989
R19638 vdd.n1995 vdd.t172 1.92771
R19639 vdd.n2071 vdd.t157 1.92771
R19640 vdd.n2484 vdd.t165 1.92771
R19641 vdd.n2603 vdd.t161 1.92771
R19642 vdd.n1871 vdd.t87 1.70098
R19643 vdd.n798 vdd.t105 1.70098
R19644 vdd.t88 vdd.n664 1.70098
R19645 vdd.n2374 vdd.t20 1.70098
R19646 vdd.n1455 vdd.t27 1.24752
R19647 vdd.t64 vdd.n3041 1.24752
R19648 vdd.n295 vdd.n255 1.16414
R19649 vdd.n288 vdd.n287 1.16414
R19650 vdd.n248 vdd.n208 1.16414
R19651 vdd.n241 vdd.n240 1.16414
R19652 vdd.n205 vdd.n165 1.16414
R19653 vdd.n198 vdd.n197 1.16414
R19654 vdd.n158 vdd.n118 1.16414
R19655 vdd.n151 vdd.n150 1.16414
R19656 vdd.n116 vdd.n76 1.16414
R19657 vdd.n109 vdd.n108 1.16414
R19658 vdd.n69 vdd.n29 1.16414
R19659 vdd.n62 vdd.n61 1.16414
R19660 vdd.n1110 vdd.n1070 1.16414
R19661 vdd.n1103 vdd.n1102 1.16414
R19662 vdd.n1157 vdd.n1117 1.16414
R19663 vdd.n1150 vdd.n1149 1.16414
R19664 vdd.n1020 vdd.n980 1.16414
R19665 vdd.n1013 vdd.n1012 1.16414
R19666 vdd.n1067 vdd.n1027 1.16414
R19667 vdd.n1060 vdd.n1059 1.16414
R19668 vdd.n931 vdd.n891 1.16414
R19669 vdd.n924 vdd.n923 1.16414
R19670 vdd.n978 vdd.n938 1.16414
R19671 vdd.n971 vdd.n970 1.16414
R19672 vdd.n2038 vdd.t15 1.13415
R19673 vdd.n2514 vdd.t109 1.13415
R19674 vdd.n1481 vdd.t31 1.02079
R19675 vdd.t176 vdd.t115 1.02079
R19676 vdd.t19 vdd.t140 1.02079
R19677 vdd.t51 vdd.n456 1.02079
R19678 vdd.n1326 vdd.n1322 0.970197
R19679 vdd.n1950 vdd.n1949 0.970197
R19680 vdd.n2911 vdd.n2910 0.970197
R19681 vdd.n2715 vdd.n2713 0.970197
R19682 vdd.n2014 vdd.t115 0.794056
R19683 vdd.n2050 vdd.t6 0.794056
R19684 vdd.n2502 vdd.t9 0.794056
R19685 vdd.n2540 vdd.t19 0.794056
R19686 vdd.n1160 vdd.n28 0.74827
R19687 vdd vdd.n3048 0.740437
R19688 vdd.n1430 vdd.t136 0.567326
R19689 vdd.n3026 vdd.t147 0.567326
R19690 vdd.n1940 vdd.n1939 0.537085
R19691 vdd.n2845 vdd.n2844 0.537085
R19692 vdd.n3022 vdd.n3021 0.537085
R19693 vdd.n2904 vdd.n2903 0.537085
R19694 vdd.n2709 vdd.n476 0.537085
R19695 vdd.n1503 vdd.n857 0.537085
R19696 vdd.n1324 vdd.n1189 0.537085
R19697 vdd.n1426 vdd.n1425 0.537085
R19698 vdd.n4 vdd.n2 0.459552
R19699 vdd.n11 vdd.n9 0.459552
R19700 vdd.n293 vdd.n292 0.388379
R19701 vdd.n259 vdd.n257 0.388379
R19702 vdd.n246 vdd.n245 0.388379
R19703 vdd.n212 vdd.n210 0.388379
R19704 vdd.n203 vdd.n202 0.388379
R19705 vdd.n169 vdd.n167 0.388379
R19706 vdd.n156 vdd.n155 0.388379
R19707 vdd.n122 vdd.n120 0.388379
R19708 vdd.n114 vdd.n113 0.388379
R19709 vdd.n80 vdd.n78 0.388379
R19710 vdd.n67 vdd.n66 0.388379
R19711 vdd.n33 vdd.n31 0.388379
R19712 vdd.n1108 vdd.n1107 0.388379
R19713 vdd.n1074 vdd.n1072 0.388379
R19714 vdd.n1155 vdd.n1154 0.388379
R19715 vdd.n1121 vdd.n1119 0.388379
R19716 vdd.n1018 vdd.n1017 0.388379
R19717 vdd.n984 vdd.n982 0.388379
R19718 vdd.n1065 vdd.n1064 0.388379
R19719 vdd.n1031 vdd.n1029 0.388379
R19720 vdd.n929 vdd.n928 0.388379
R19721 vdd.n895 vdd.n893 0.388379
R19722 vdd.n976 vdd.n975 0.388379
R19723 vdd.n942 vdd.n940 0.388379
R19724 vdd.n19 vdd.n17 0.387128
R19725 vdd.n24 vdd.n22 0.387128
R19726 vdd.n6 vdd.n4 0.358259
R19727 vdd.n13 vdd.n11 0.358259
R19728 vdd.n252 vdd.n250 0.358259
R19729 vdd.n254 vdd.n252 0.358259
R19730 vdd.n296 vdd.n254 0.358259
R19731 vdd.n162 vdd.n160 0.358259
R19732 vdd.n164 vdd.n162 0.358259
R19733 vdd.n206 vdd.n164 0.358259
R19734 vdd.n73 vdd.n71 0.358259
R19735 vdd.n75 vdd.n73 0.358259
R19736 vdd.n117 vdd.n75 0.358259
R19737 vdd.n1158 vdd.n1116 0.358259
R19738 vdd.n1116 vdd.n1114 0.358259
R19739 vdd.n1114 vdd.n1112 0.358259
R19740 vdd.n1068 vdd.n1026 0.358259
R19741 vdd.n1026 vdd.n1024 0.358259
R19742 vdd.n1024 vdd.n1022 0.358259
R19743 vdd.n979 vdd.n937 0.358259
R19744 vdd.n937 vdd.n935 0.358259
R19745 vdd.n935 vdd.n933 0.358259
R19746 vdd.n14 vdd.n6 0.334552
R19747 vdd.n14 vdd.n13 0.334552
R19748 vdd.n27 vdd.n19 0.21707
R19749 vdd.n27 vdd.n24 0.21707
R19750 vdd.n294 vdd.n256 0.155672
R19751 vdd.n286 vdd.n256 0.155672
R19752 vdd.n286 vdd.n285 0.155672
R19753 vdd.n285 vdd.n261 0.155672
R19754 vdd.n278 vdd.n261 0.155672
R19755 vdd.n278 vdd.n277 0.155672
R19756 vdd.n277 vdd.n265 0.155672
R19757 vdd.n270 vdd.n265 0.155672
R19758 vdd.n247 vdd.n209 0.155672
R19759 vdd.n239 vdd.n209 0.155672
R19760 vdd.n239 vdd.n238 0.155672
R19761 vdd.n238 vdd.n214 0.155672
R19762 vdd.n231 vdd.n214 0.155672
R19763 vdd.n231 vdd.n230 0.155672
R19764 vdd.n230 vdd.n218 0.155672
R19765 vdd.n223 vdd.n218 0.155672
R19766 vdd.n204 vdd.n166 0.155672
R19767 vdd.n196 vdd.n166 0.155672
R19768 vdd.n196 vdd.n195 0.155672
R19769 vdd.n195 vdd.n171 0.155672
R19770 vdd.n188 vdd.n171 0.155672
R19771 vdd.n188 vdd.n187 0.155672
R19772 vdd.n187 vdd.n175 0.155672
R19773 vdd.n180 vdd.n175 0.155672
R19774 vdd.n157 vdd.n119 0.155672
R19775 vdd.n149 vdd.n119 0.155672
R19776 vdd.n149 vdd.n148 0.155672
R19777 vdd.n148 vdd.n124 0.155672
R19778 vdd.n141 vdd.n124 0.155672
R19779 vdd.n141 vdd.n140 0.155672
R19780 vdd.n140 vdd.n128 0.155672
R19781 vdd.n133 vdd.n128 0.155672
R19782 vdd.n115 vdd.n77 0.155672
R19783 vdd.n107 vdd.n77 0.155672
R19784 vdd.n107 vdd.n106 0.155672
R19785 vdd.n106 vdd.n82 0.155672
R19786 vdd.n99 vdd.n82 0.155672
R19787 vdd.n99 vdd.n98 0.155672
R19788 vdd.n98 vdd.n86 0.155672
R19789 vdd.n91 vdd.n86 0.155672
R19790 vdd.n68 vdd.n30 0.155672
R19791 vdd.n60 vdd.n30 0.155672
R19792 vdd.n60 vdd.n59 0.155672
R19793 vdd.n59 vdd.n35 0.155672
R19794 vdd.n52 vdd.n35 0.155672
R19795 vdd.n52 vdd.n51 0.155672
R19796 vdd.n51 vdd.n39 0.155672
R19797 vdd.n44 vdd.n39 0.155672
R19798 vdd.n1109 vdd.n1071 0.155672
R19799 vdd.n1101 vdd.n1071 0.155672
R19800 vdd.n1101 vdd.n1100 0.155672
R19801 vdd.n1100 vdd.n1076 0.155672
R19802 vdd.n1093 vdd.n1076 0.155672
R19803 vdd.n1093 vdd.n1092 0.155672
R19804 vdd.n1092 vdd.n1080 0.155672
R19805 vdd.n1085 vdd.n1080 0.155672
R19806 vdd.n1156 vdd.n1118 0.155672
R19807 vdd.n1148 vdd.n1118 0.155672
R19808 vdd.n1148 vdd.n1147 0.155672
R19809 vdd.n1147 vdd.n1123 0.155672
R19810 vdd.n1140 vdd.n1123 0.155672
R19811 vdd.n1140 vdd.n1139 0.155672
R19812 vdd.n1139 vdd.n1127 0.155672
R19813 vdd.n1132 vdd.n1127 0.155672
R19814 vdd.n1019 vdd.n981 0.155672
R19815 vdd.n1011 vdd.n981 0.155672
R19816 vdd.n1011 vdd.n1010 0.155672
R19817 vdd.n1010 vdd.n986 0.155672
R19818 vdd.n1003 vdd.n986 0.155672
R19819 vdd.n1003 vdd.n1002 0.155672
R19820 vdd.n1002 vdd.n990 0.155672
R19821 vdd.n995 vdd.n990 0.155672
R19822 vdd.n1066 vdd.n1028 0.155672
R19823 vdd.n1058 vdd.n1028 0.155672
R19824 vdd.n1058 vdd.n1057 0.155672
R19825 vdd.n1057 vdd.n1033 0.155672
R19826 vdd.n1050 vdd.n1033 0.155672
R19827 vdd.n1050 vdd.n1049 0.155672
R19828 vdd.n1049 vdd.n1037 0.155672
R19829 vdd.n1042 vdd.n1037 0.155672
R19830 vdd.n930 vdd.n892 0.155672
R19831 vdd.n922 vdd.n892 0.155672
R19832 vdd.n922 vdd.n921 0.155672
R19833 vdd.n921 vdd.n897 0.155672
R19834 vdd.n914 vdd.n897 0.155672
R19835 vdd.n914 vdd.n913 0.155672
R19836 vdd.n913 vdd.n901 0.155672
R19837 vdd.n906 vdd.n901 0.155672
R19838 vdd.n977 vdd.n939 0.155672
R19839 vdd.n969 vdd.n939 0.155672
R19840 vdd.n969 vdd.n968 0.155672
R19841 vdd.n968 vdd.n944 0.155672
R19842 vdd.n961 vdd.n944 0.155672
R19843 vdd.n961 vdd.n960 0.155672
R19844 vdd.n960 vdd.n948 0.155672
R19845 vdd.n953 vdd.n948 0.155672
R19846 vdd.n1715 vdd.n1520 0.152939
R19847 vdd.n1526 vdd.n1520 0.152939
R19848 vdd.n1527 vdd.n1526 0.152939
R19849 vdd.n1528 vdd.n1527 0.152939
R19850 vdd.n1529 vdd.n1528 0.152939
R19851 vdd.n1533 vdd.n1529 0.152939
R19852 vdd.n1534 vdd.n1533 0.152939
R19853 vdd.n1535 vdd.n1534 0.152939
R19854 vdd.n1536 vdd.n1535 0.152939
R19855 vdd.n1540 vdd.n1536 0.152939
R19856 vdd.n1541 vdd.n1540 0.152939
R19857 vdd.n1542 vdd.n1541 0.152939
R19858 vdd.n1690 vdd.n1542 0.152939
R19859 vdd.n1690 vdd.n1689 0.152939
R19860 vdd.n1689 vdd.n1688 0.152939
R19861 vdd.n1688 vdd.n1548 0.152939
R19862 vdd.n1553 vdd.n1548 0.152939
R19863 vdd.n1554 vdd.n1553 0.152939
R19864 vdd.n1555 vdd.n1554 0.152939
R19865 vdd.n1559 vdd.n1555 0.152939
R19866 vdd.n1560 vdd.n1559 0.152939
R19867 vdd.n1561 vdd.n1560 0.152939
R19868 vdd.n1562 vdd.n1561 0.152939
R19869 vdd.n1566 vdd.n1562 0.152939
R19870 vdd.n1567 vdd.n1566 0.152939
R19871 vdd.n1568 vdd.n1567 0.152939
R19872 vdd.n1569 vdd.n1568 0.152939
R19873 vdd.n1573 vdd.n1569 0.152939
R19874 vdd.n1574 vdd.n1573 0.152939
R19875 vdd.n1575 vdd.n1574 0.152939
R19876 vdd.n1576 vdd.n1575 0.152939
R19877 vdd.n1580 vdd.n1576 0.152939
R19878 vdd.n1581 vdd.n1580 0.152939
R19879 vdd.n1582 vdd.n1581 0.152939
R19880 vdd.n1651 vdd.n1582 0.152939
R19881 vdd.n1651 vdd.n1650 0.152939
R19882 vdd.n1650 vdd.n1649 0.152939
R19883 vdd.n1649 vdd.n1588 0.152939
R19884 vdd.n1593 vdd.n1588 0.152939
R19885 vdd.n1594 vdd.n1593 0.152939
R19886 vdd.n1595 vdd.n1594 0.152939
R19887 vdd.n1599 vdd.n1595 0.152939
R19888 vdd.n1600 vdd.n1599 0.152939
R19889 vdd.n1601 vdd.n1600 0.152939
R19890 vdd.n1602 vdd.n1601 0.152939
R19891 vdd.n1606 vdd.n1602 0.152939
R19892 vdd.n1607 vdd.n1606 0.152939
R19893 vdd.n1608 vdd.n1607 0.152939
R19894 vdd.n1609 vdd.n1608 0.152939
R19895 vdd.n1610 vdd.n1609 0.152939
R19896 vdd.n1610 vdd.n854 0.152939
R19897 vdd.n1939 vdd.n1514 0.152939
R19898 vdd.n1477 vdd.n1476 0.152939
R19899 vdd.n1478 vdd.n1477 0.152939
R19900 vdd.n1478 vdd.n879 0.152939
R19901 vdd.n1493 vdd.n879 0.152939
R19902 vdd.n1494 vdd.n1493 0.152939
R19903 vdd.n1495 vdd.n1494 0.152939
R19904 vdd.n1495 vdd.n867 0.152939
R19905 vdd.n1512 vdd.n867 0.152939
R19906 vdd.n1513 vdd.n1512 0.152939
R19907 vdd.n1940 vdd.n1513 0.152939
R19908 vdd.n524 vdd.n519 0.152939
R19909 vdd.n525 vdd.n524 0.152939
R19910 vdd.n526 vdd.n525 0.152939
R19911 vdd.n527 vdd.n526 0.152939
R19912 vdd.n528 vdd.n527 0.152939
R19913 vdd.n529 vdd.n528 0.152939
R19914 vdd.n530 vdd.n529 0.152939
R19915 vdd.n531 vdd.n530 0.152939
R19916 vdd.n532 vdd.n531 0.152939
R19917 vdd.n533 vdd.n532 0.152939
R19918 vdd.n534 vdd.n533 0.152939
R19919 vdd.n535 vdd.n534 0.152939
R19920 vdd.n2803 vdd.n535 0.152939
R19921 vdd.n2803 vdd.n2802 0.152939
R19922 vdd.n2802 vdd.n2801 0.152939
R19923 vdd.n2801 vdd.n537 0.152939
R19924 vdd.n538 vdd.n537 0.152939
R19925 vdd.n539 vdd.n538 0.152939
R19926 vdd.n540 vdd.n539 0.152939
R19927 vdd.n541 vdd.n540 0.152939
R19928 vdd.n542 vdd.n541 0.152939
R19929 vdd.n543 vdd.n542 0.152939
R19930 vdd.n544 vdd.n543 0.152939
R19931 vdd.n545 vdd.n544 0.152939
R19932 vdd.n546 vdd.n545 0.152939
R19933 vdd.n547 vdd.n546 0.152939
R19934 vdd.n548 vdd.n547 0.152939
R19935 vdd.n549 vdd.n548 0.152939
R19936 vdd.n550 vdd.n549 0.152939
R19937 vdd.n551 vdd.n550 0.152939
R19938 vdd.n552 vdd.n551 0.152939
R19939 vdd.n553 vdd.n552 0.152939
R19940 vdd.n554 vdd.n553 0.152939
R19941 vdd.n555 vdd.n554 0.152939
R19942 vdd.n2757 vdd.n555 0.152939
R19943 vdd.n2757 vdd.n2756 0.152939
R19944 vdd.n2756 vdd.n2755 0.152939
R19945 vdd.n2755 vdd.n559 0.152939
R19946 vdd.n560 vdd.n559 0.152939
R19947 vdd.n561 vdd.n560 0.152939
R19948 vdd.n562 vdd.n561 0.152939
R19949 vdd.n563 vdd.n562 0.152939
R19950 vdd.n564 vdd.n563 0.152939
R19951 vdd.n565 vdd.n564 0.152939
R19952 vdd.n566 vdd.n565 0.152939
R19953 vdd.n567 vdd.n566 0.152939
R19954 vdd.n568 vdd.n567 0.152939
R19955 vdd.n569 vdd.n568 0.152939
R19956 vdd.n570 vdd.n569 0.152939
R19957 vdd.n571 vdd.n570 0.152939
R19958 vdd.n572 vdd.n571 0.152939
R19959 vdd.n2844 vdd.n481 0.152939
R19960 vdd.n2846 vdd.n2845 0.152939
R19961 vdd.n2846 vdd.n470 0.152939
R19962 vdd.n2861 vdd.n470 0.152939
R19963 vdd.n2862 vdd.n2861 0.152939
R19964 vdd.n2863 vdd.n2862 0.152939
R19965 vdd.n2863 vdd.n459 0.152939
R19966 vdd.n2877 vdd.n459 0.152939
R19967 vdd.n2878 vdd.n2877 0.152939
R19968 vdd.n2879 vdd.n2878 0.152939
R19969 vdd.n2879 vdd.n298 0.152939
R19970 vdd.n3046 vdd.n299 0.152939
R19971 vdd.n310 vdd.n299 0.152939
R19972 vdd.n311 vdd.n310 0.152939
R19973 vdd.n312 vdd.n311 0.152939
R19974 vdd.n320 vdd.n312 0.152939
R19975 vdd.n321 vdd.n320 0.152939
R19976 vdd.n322 vdd.n321 0.152939
R19977 vdd.n323 vdd.n322 0.152939
R19978 vdd.n331 vdd.n323 0.152939
R19979 vdd.n3022 vdd.n331 0.152939
R19980 vdd.n3021 vdd.n332 0.152939
R19981 vdd.n335 vdd.n332 0.152939
R19982 vdd.n339 vdd.n335 0.152939
R19983 vdd.n340 vdd.n339 0.152939
R19984 vdd.n341 vdd.n340 0.152939
R19985 vdd.n342 vdd.n341 0.152939
R19986 vdd.n343 vdd.n342 0.152939
R19987 vdd.n347 vdd.n343 0.152939
R19988 vdd.n348 vdd.n347 0.152939
R19989 vdd.n349 vdd.n348 0.152939
R19990 vdd.n350 vdd.n349 0.152939
R19991 vdd.n354 vdd.n350 0.152939
R19992 vdd.n355 vdd.n354 0.152939
R19993 vdd.n356 vdd.n355 0.152939
R19994 vdd.n357 vdd.n356 0.152939
R19995 vdd.n361 vdd.n357 0.152939
R19996 vdd.n362 vdd.n361 0.152939
R19997 vdd.n363 vdd.n362 0.152939
R19998 vdd.n2987 vdd.n363 0.152939
R19999 vdd.n2987 vdd.n2986 0.152939
R20000 vdd.n2986 vdd.n2985 0.152939
R20001 vdd.n2985 vdd.n369 0.152939
R20002 vdd.n374 vdd.n369 0.152939
R20003 vdd.n375 vdd.n374 0.152939
R20004 vdd.n376 vdd.n375 0.152939
R20005 vdd.n380 vdd.n376 0.152939
R20006 vdd.n381 vdd.n380 0.152939
R20007 vdd.n382 vdd.n381 0.152939
R20008 vdd.n383 vdd.n382 0.152939
R20009 vdd.n387 vdd.n383 0.152939
R20010 vdd.n388 vdd.n387 0.152939
R20011 vdd.n389 vdd.n388 0.152939
R20012 vdd.n390 vdd.n389 0.152939
R20013 vdd.n394 vdd.n390 0.152939
R20014 vdd.n395 vdd.n394 0.152939
R20015 vdd.n396 vdd.n395 0.152939
R20016 vdd.n397 vdd.n396 0.152939
R20017 vdd.n401 vdd.n397 0.152939
R20018 vdd.n402 vdd.n401 0.152939
R20019 vdd.n403 vdd.n402 0.152939
R20020 vdd.n2948 vdd.n403 0.152939
R20021 vdd.n2948 vdd.n2947 0.152939
R20022 vdd.n2947 vdd.n2946 0.152939
R20023 vdd.n2946 vdd.n409 0.152939
R20024 vdd.n414 vdd.n409 0.152939
R20025 vdd.n415 vdd.n414 0.152939
R20026 vdd.n416 vdd.n415 0.152939
R20027 vdd.n420 vdd.n416 0.152939
R20028 vdd.n421 vdd.n420 0.152939
R20029 vdd.n422 vdd.n421 0.152939
R20030 vdd.n423 vdd.n422 0.152939
R20031 vdd.n427 vdd.n423 0.152939
R20032 vdd.n428 vdd.n427 0.152939
R20033 vdd.n429 vdd.n428 0.152939
R20034 vdd.n430 vdd.n429 0.152939
R20035 vdd.n434 vdd.n430 0.152939
R20036 vdd.n435 vdd.n434 0.152939
R20037 vdd.n436 vdd.n435 0.152939
R20038 vdd.n437 vdd.n436 0.152939
R20039 vdd.n441 vdd.n437 0.152939
R20040 vdd.n442 vdd.n441 0.152939
R20041 vdd.n443 vdd.n442 0.152939
R20042 vdd.n2904 vdd.n443 0.152939
R20043 vdd.n2852 vdd.n476 0.152939
R20044 vdd.n2853 vdd.n2852 0.152939
R20045 vdd.n2854 vdd.n2853 0.152939
R20046 vdd.n2854 vdd.n464 0.152939
R20047 vdd.n2869 vdd.n464 0.152939
R20048 vdd.n2870 vdd.n2869 0.152939
R20049 vdd.n2871 vdd.n2870 0.152939
R20050 vdd.n2871 vdd.n452 0.152939
R20051 vdd.n2885 vdd.n452 0.152939
R20052 vdd.n2886 vdd.n2885 0.152939
R20053 vdd.n2887 vdd.n2886 0.152939
R20054 vdd.n2887 vdd.n450 0.152939
R20055 vdd.n2891 vdd.n450 0.152939
R20056 vdd.n2892 vdd.n2891 0.152939
R20057 vdd.n2893 vdd.n2892 0.152939
R20058 vdd.n2893 vdd.n447 0.152939
R20059 vdd.n2897 vdd.n447 0.152939
R20060 vdd.n2898 vdd.n2897 0.152939
R20061 vdd.n2899 vdd.n2898 0.152939
R20062 vdd.n2899 vdd.n444 0.152939
R20063 vdd.n2903 vdd.n444 0.152939
R20064 vdd.n2709 vdd.n2708 0.152939
R20065 vdd.n1951 vdd.n857 0.152939
R20066 vdd.n1433 vdd.n1189 0.152939
R20067 vdd.n1434 vdd.n1433 0.152939
R20068 vdd.n1435 vdd.n1434 0.152939
R20069 vdd.n1435 vdd.n1177 0.152939
R20070 vdd.n1450 vdd.n1177 0.152939
R20071 vdd.n1451 vdd.n1450 0.152939
R20072 vdd.n1452 vdd.n1451 0.152939
R20073 vdd.n1452 vdd.n1167 0.152939
R20074 vdd.n1468 vdd.n1167 0.152939
R20075 vdd.n1469 vdd.n1468 0.152939
R20076 vdd.n1470 vdd.n1469 0.152939
R20077 vdd.n1470 vdd.n884 0.152939
R20078 vdd.n1484 vdd.n884 0.152939
R20079 vdd.n1485 vdd.n1484 0.152939
R20080 vdd.n1486 vdd.n1485 0.152939
R20081 vdd.n1486 vdd.n874 0.152939
R20082 vdd.n1501 vdd.n874 0.152939
R20083 vdd.n1502 vdd.n1501 0.152939
R20084 vdd.n1505 vdd.n1502 0.152939
R20085 vdd.n1505 vdd.n1504 0.152939
R20086 vdd.n1504 vdd.n1503 0.152939
R20087 vdd.n1425 vdd.n1194 0.152939
R20088 vdd.n1418 vdd.n1194 0.152939
R20089 vdd.n1418 vdd.n1417 0.152939
R20090 vdd.n1417 vdd.n1416 0.152939
R20091 vdd.n1416 vdd.n1231 0.152939
R20092 vdd.n1412 vdd.n1231 0.152939
R20093 vdd.n1412 vdd.n1411 0.152939
R20094 vdd.n1411 vdd.n1410 0.152939
R20095 vdd.n1410 vdd.n1237 0.152939
R20096 vdd.n1406 vdd.n1237 0.152939
R20097 vdd.n1406 vdd.n1405 0.152939
R20098 vdd.n1405 vdd.n1404 0.152939
R20099 vdd.n1404 vdd.n1243 0.152939
R20100 vdd.n1400 vdd.n1243 0.152939
R20101 vdd.n1400 vdd.n1399 0.152939
R20102 vdd.n1399 vdd.n1398 0.152939
R20103 vdd.n1398 vdd.n1249 0.152939
R20104 vdd.n1394 vdd.n1249 0.152939
R20105 vdd.n1394 vdd.n1393 0.152939
R20106 vdd.n1393 vdd.n1392 0.152939
R20107 vdd.n1392 vdd.n1257 0.152939
R20108 vdd.n1388 vdd.n1257 0.152939
R20109 vdd.n1388 vdd.n1387 0.152939
R20110 vdd.n1387 vdd.n1386 0.152939
R20111 vdd.n1386 vdd.n1263 0.152939
R20112 vdd.n1382 vdd.n1263 0.152939
R20113 vdd.n1382 vdd.n1381 0.152939
R20114 vdd.n1381 vdd.n1380 0.152939
R20115 vdd.n1380 vdd.n1269 0.152939
R20116 vdd.n1376 vdd.n1269 0.152939
R20117 vdd.n1376 vdd.n1375 0.152939
R20118 vdd.n1375 vdd.n1374 0.152939
R20119 vdd.n1374 vdd.n1275 0.152939
R20120 vdd.n1370 vdd.n1275 0.152939
R20121 vdd.n1370 vdd.n1369 0.152939
R20122 vdd.n1369 vdd.n1368 0.152939
R20123 vdd.n1368 vdd.n1281 0.152939
R20124 vdd.n1364 vdd.n1281 0.152939
R20125 vdd.n1364 vdd.n1363 0.152939
R20126 vdd.n1363 vdd.n1362 0.152939
R20127 vdd.n1362 vdd.n1287 0.152939
R20128 vdd.n1355 vdd.n1287 0.152939
R20129 vdd.n1355 vdd.n1354 0.152939
R20130 vdd.n1354 vdd.n1353 0.152939
R20131 vdd.n1353 vdd.n1292 0.152939
R20132 vdd.n1349 vdd.n1292 0.152939
R20133 vdd.n1349 vdd.n1348 0.152939
R20134 vdd.n1348 vdd.n1347 0.152939
R20135 vdd.n1347 vdd.n1298 0.152939
R20136 vdd.n1343 vdd.n1298 0.152939
R20137 vdd.n1343 vdd.n1342 0.152939
R20138 vdd.n1342 vdd.n1341 0.152939
R20139 vdd.n1341 vdd.n1304 0.152939
R20140 vdd.n1337 vdd.n1304 0.152939
R20141 vdd.n1337 vdd.n1336 0.152939
R20142 vdd.n1336 vdd.n1335 0.152939
R20143 vdd.n1335 vdd.n1310 0.152939
R20144 vdd.n1331 vdd.n1310 0.152939
R20145 vdd.n1331 vdd.n1330 0.152939
R20146 vdd.n1330 vdd.n1329 0.152939
R20147 vdd.n1329 vdd.n1316 0.152939
R20148 vdd.n1325 vdd.n1316 0.152939
R20149 vdd.n1325 vdd.n1324 0.152939
R20150 vdd.n1427 vdd.n1426 0.152939
R20151 vdd.n1427 vdd.n1183 0.152939
R20152 vdd.n1442 vdd.n1183 0.152939
R20153 vdd.n1443 vdd.n1442 0.152939
R20154 vdd.n1444 vdd.n1443 0.152939
R20155 vdd.n1444 vdd.n1172 0.152939
R20156 vdd.n1459 vdd.n1172 0.152939
R20157 vdd.n1460 vdd.n1459 0.152939
R20158 vdd.n1462 vdd.n1460 0.152939
R20159 vdd.n1462 vdd.n1461 0.152939
R20160 vdd.n1929 vdd.n1514 0.110256
R20161 vdd.n2836 vdd.n481 0.110256
R20162 vdd.n2708 vdd.n2707 0.110256
R20163 vdd.n1952 vdd.n1951 0.110256
R20164 vdd.n1476 vdd.n1161 0.0695946
R20165 vdd.n3047 vdd.n298 0.0695946
R20166 vdd.n3047 vdd.n3046 0.0695946
R20167 vdd.n1461 vdd.n1161 0.0695946
R20168 vdd.n1929 vdd.n1715 0.0431829
R20169 vdd.n1952 vdd.n854 0.0431829
R20170 vdd.n2836 vdd.n519 0.0431829
R20171 vdd.n2707 vdd.n572 0.0431829
R20172 vdd vdd.n28 0.00833333
R20173 a_n1996_n452.n82 a_n1996_n452.t60 512.366
R20174 a_n1996_n452.n81 a_n1996_n452.t51 512.366
R20175 a_n1996_n452.n80 a_n1996_n452.t45 512.366
R20176 a_n1996_n452.n84 a_n1996_n452.t68 512.366
R20177 a_n1996_n452.n83 a_n1996_n452.t57 512.366
R20178 a_n1996_n452.n79 a_n1996_n452.t56 512.366
R20179 a_n1996_n452.n86 a_n1996_n452.t64 512.366
R20180 a_n1996_n452.n85 a_n1996_n452.t49 512.366
R20181 a_n1996_n452.n78 a_n1996_n452.t50 512.366
R20182 a_n1996_n452.n88 a_n1996_n452.t53 512.366
R20183 a_n1996_n452.n87 a_n1996_n452.t62 512.366
R20184 a_n1996_n452.n77 a_n1996_n452.t44 512.366
R20185 a_n1996_n452.n25 a_n1996_n452.t71 539.01
R20186 a_n1996_n452.n69 a_n1996_n452.t54 512.366
R20187 a_n1996_n452.n68 a_n1996_n452.t58 512.366
R20188 a_n1996_n452.n66 a_n1996_n452.t48 512.366
R20189 a_n1996_n452.n67 a_n1996_n452.t63 512.366
R20190 a_n1996_n452.n21 a_n1996_n452.t18 539.01
R20191 a_n1996_n452.n72 a_n1996_n452.t16 512.366
R20192 a_n1996_n452.n71 a_n1996_n452.t36 512.366
R20193 a_n1996_n452.n55 a_n1996_n452.t32 512.366
R20194 a_n1996_n452.n70 a_n1996_n452.t34 512.366
R20195 a_n1996_n452.n15 a_n1996_n452.t30 539.01
R20196 a_n1996_n452.n93 a_n1996_n452.t28 512.366
R20197 a_n1996_n452.n94 a_n1996_n452.t20 512.366
R20198 a_n1996_n452.n53 a_n1996_n452.t14 512.366
R20199 a_n1996_n452.n95 a_n1996_n452.t22 512.366
R20200 a_n1996_n452.n19 a_n1996_n452.t66 539.01
R20201 a_n1996_n452.n90 a_n1996_n452.t67 512.366
R20202 a_n1996_n452.n91 a_n1996_n452.t46 512.366
R20203 a_n1996_n452.n54 a_n1996_n452.t52 512.366
R20204 a_n1996_n452.n92 a_n1996_n452.t61 512.366
R20205 a_n1996_n452.n4 a_n1996_n452.n50 70.1674
R20206 a_n1996_n452.n6 a_n1996_n452.n48 70.1674
R20207 a_n1996_n452.n8 a_n1996_n452.n46 70.1674
R20208 a_n1996_n452.n10 a_n1996_n452.n44 70.1674
R20209 a_n1996_n452.n33 a_n1996_n452.n23 70.3058
R20210 a_n1996_n452.n51 a_n1996_n452.n29 70.3058
R20211 a_n1996_n452.n24 a_n1996_n452.n31 70.1674
R20212 a_n1996_n452.n31 a_n1996_n452.n66 20.9683
R20213 a_n1996_n452.n30 a_n1996_n452.n24 75.0448
R20214 a_n1996_n452.n68 a_n1996_n452.n30 11.2134
R20215 a_n1996_n452.n22 a_n1996_n452.n25 44.8194
R20216 a_n1996_n452.n29 a_n1996_n452.n36 70.1674
R20217 a_n1996_n452.n36 a_n1996_n452.n55 20.9683
R20218 a_n1996_n452.n35 a_n1996_n452.n34 75.0448
R20219 a_n1996_n452.n71 a_n1996_n452.n35 11.2134
R20220 a_n1996_n452.n20 a_n1996_n452.n21 44.8194
R20221 a_n1996_n452.n12 a_n1996_n452.n42 70.3058
R20222 a_n1996_n452.n16 a_n1996_n452.n39 70.3058
R20223 a_n1996_n452.n38 a_n1996_n452.n17 70.1674
R20224 a_n1996_n452.n38 a_n1996_n452.n54 20.9683
R20225 a_n1996_n452.n17 a_n1996_n452.n37 75.0448
R20226 a_n1996_n452.n91 a_n1996_n452.n37 11.2134
R20227 a_n1996_n452.n18 a_n1996_n452.n19 44.8194
R20228 a_n1996_n452.n41 a_n1996_n452.n13 70.1674
R20229 a_n1996_n452.n41 a_n1996_n452.n53 20.9683
R20230 a_n1996_n452.n13 a_n1996_n452.n40 75.0448
R20231 a_n1996_n452.n94 a_n1996_n452.n40 11.2134
R20232 a_n1996_n452.n14 a_n1996_n452.n15 44.8194
R20233 a_n1996_n452.n44 a_n1996_n452.n77 20.9683
R20234 a_n1996_n452.n43 a_n1996_n452.n11 75.0448
R20235 a_n1996_n452.n87 a_n1996_n452.n43 11.2134
R20236 a_n1996_n452.n11 a_n1996_n452.n88 161.3
R20237 a_n1996_n452.n46 a_n1996_n452.n78 20.9683
R20238 a_n1996_n452.n45 a_n1996_n452.n9 75.0448
R20239 a_n1996_n452.n85 a_n1996_n452.n45 11.2134
R20240 a_n1996_n452.n9 a_n1996_n452.n86 161.3
R20241 a_n1996_n452.n48 a_n1996_n452.n79 20.9683
R20242 a_n1996_n452.n47 a_n1996_n452.n7 75.0448
R20243 a_n1996_n452.n83 a_n1996_n452.n47 11.2134
R20244 a_n1996_n452.n7 a_n1996_n452.n84 161.3
R20245 a_n1996_n452.n50 a_n1996_n452.n80 20.9683
R20246 a_n1996_n452.n49 a_n1996_n452.n5 75.0448
R20247 a_n1996_n452.n81 a_n1996_n452.n49 11.2134
R20248 a_n1996_n452.n5 a_n1996_n452.n82 161.3
R20249 a_n1996_n452.n3 a_n1996_n452.n64 81.3764
R20250 a_n1996_n452.n1 a_n1996_n452.n59 81.3764
R20251 a_n1996_n452.n0 a_n1996_n452.n56 81.3764
R20252 a_n1996_n452.n3 a_n1996_n452.n65 80.9324
R20253 a_n1996_n452.n3 a_n1996_n452.n63 80.9324
R20254 a_n1996_n452.n2 a_n1996_n452.n62 80.9324
R20255 a_n1996_n452.n2 a_n1996_n452.n61 80.9324
R20256 a_n1996_n452.n1 a_n1996_n452.n60 80.9324
R20257 a_n1996_n452.n1 a_n1996_n452.n58 80.9324
R20258 a_n1996_n452.n0 a_n1996_n452.n57 80.9324
R20259 a_n1996_n452.n27 a_n1996_n452.t31 74.6477
R20260 a_n1996_n452.n26 a_n1996_n452.t27 74.6477
R20261 a_n1996_n452.n75 a_n1996_n452.t19 74.2899
R20262 a_n1996_n452.n28 a_n1996_n452.t25 74.2897
R20263 a_n1996_n452.n27 a_n1996_n452.n52 70.6783
R20264 a_n1996_n452.n26 a_n1996_n452.n73 70.6783
R20265 a_n1996_n452.n26 a_n1996_n452.n74 70.6783
R20266 a_n1996_n452.n97 a_n1996_n452.n28 70.6782
R20267 a_n1996_n452.n82 a_n1996_n452.n81 48.2005
R20268 a_n1996_n452.t65 a_n1996_n452.n50 533.335
R20269 a_n1996_n452.n84 a_n1996_n452.n83 48.2005
R20270 a_n1996_n452.t70 a_n1996_n452.n48 533.335
R20271 a_n1996_n452.n86 a_n1996_n452.n85 48.2005
R20272 a_n1996_n452.t59 a_n1996_n452.n46 533.335
R20273 a_n1996_n452.n88 a_n1996_n452.n87 48.2005
R20274 a_n1996_n452.t55 a_n1996_n452.n44 533.335
R20275 a_n1996_n452.n69 a_n1996_n452.n68 48.2005
R20276 a_n1996_n452.n67 a_n1996_n452.n31 20.9683
R20277 a_n1996_n452.n72 a_n1996_n452.n71 48.2005
R20278 a_n1996_n452.n70 a_n1996_n452.n36 20.9683
R20279 a_n1996_n452.n94 a_n1996_n452.n93 48.2005
R20280 a_n1996_n452.n95 a_n1996_n452.n41 20.9683
R20281 a_n1996_n452.n91 a_n1996_n452.n90 48.2005
R20282 a_n1996_n452.n92 a_n1996_n452.n38 20.9683
R20283 a_n1996_n452.n33 a_n1996_n452.t69 533.058
R20284 a_n1996_n452.n51 a_n1996_n452.t26 533.058
R20285 a_n1996_n452.t24 a_n1996_n452.n42 533.058
R20286 a_n1996_n452.t47 a_n1996_n452.n39 533.058
R20287 a_n1996_n452.n2 a_n1996_n452.n1 32.0139
R20288 a_n1996_n452.n49 a_n1996_n452.n80 35.3134
R20289 a_n1996_n452.n47 a_n1996_n452.n79 35.3134
R20290 a_n1996_n452.n45 a_n1996_n452.n78 35.3134
R20291 a_n1996_n452.n43 a_n1996_n452.n77 35.3134
R20292 a_n1996_n452.n30 a_n1996_n452.n66 35.3134
R20293 a_n1996_n452.n35 a_n1996_n452.n55 35.3134
R20294 a_n1996_n452.n53 a_n1996_n452.n40 35.3134
R20295 a_n1996_n452.n54 a_n1996_n452.n37 35.3134
R20296 a_n1996_n452.n29 a_n1996_n452.n3 23.891
R20297 a_n1996_n452.n18 a_n1996_n452.n89 12.046
R20298 a_n1996_n452.n23 a_n1996_n452.n32 11.8414
R20299 a_n1996_n452.n76 a_n1996_n452.n20 10.5365
R20300 a_n1996_n452.n28 a_n1996_n452.n96 9.50122
R20301 a_n1996_n452.n89 a_n1996_n452.n11 7.47588
R20302 a_n1996_n452.n4 a_n1996_n452.n32 7.47588
R20303 a_n1996_n452.n96 a_n1996_n452.n12 6.70126
R20304 a_n1996_n452.n76 a_n1996_n452.n75 5.65783
R20305 a_n1996_n452.n96 a_n1996_n452.n32 5.3452
R20306 a_n1996_n452.n29 a_n1996_n452.n22 3.95126
R20307 a_n1996_n452.n14 a_n1996_n452.n16 3.95126
R20308 a_n1996_n452.n52 a_n1996_n452.t29 3.61217
R20309 a_n1996_n452.n52 a_n1996_n452.t21 3.61217
R20310 a_n1996_n452.n73 a_n1996_n452.t33 3.61217
R20311 a_n1996_n452.n73 a_n1996_n452.t35 3.61217
R20312 a_n1996_n452.n74 a_n1996_n452.t17 3.61217
R20313 a_n1996_n452.n74 a_n1996_n452.t37 3.61217
R20314 a_n1996_n452.t15 a_n1996_n452.n97 3.61217
R20315 a_n1996_n452.n97 a_n1996_n452.t23 3.61217
R20316 a_n1996_n452.n64 a_n1996_n452.t8 2.82907
R20317 a_n1996_n452.n64 a_n1996_n452.t1 2.82907
R20318 a_n1996_n452.n65 a_n1996_n452.t12 2.82907
R20319 a_n1996_n452.n65 a_n1996_n452.t41 2.82907
R20320 a_n1996_n452.n63 a_n1996_n452.t0 2.82907
R20321 a_n1996_n452.n63 a_n1996_n452.t10 2.82907
R20322 a_n1996_n452.n62 a_n1996_n452.t43 2.82907
R20323 a_n1996_n452.n62 a_n1996_n452.t11 2.82907
R20324 a_n1996_n452.n61 a_n1996_n452.t2 2.82907
R20325 a_n1996_n452.n61 a_n1996_n452.t9 2.82907
R20326 a_n1996_n452.n59 a_n1996_n452.t13 2.82907
R20327 a_n1996_n452.n59 a_n1996_n452.t38 2.82907
R20328 a_n1996_n452.n60 a_n1996_n452.t7 2.82907
R20329 a_n1996_n452.n60 a_n1996_n452.t42 2.82907
R20330 a_n1996_n452.n58 a_n1996_n452.t39 2.82907
R20331 a_n1996_n452.n58 a_n1996_n452.t6 2.82907
R20332 a_n1996_n452.n57 a_n1996_n452.t3 2.82907
R20333 a_n1996_n452.n57 a_n1996_n452.t4 2.82907
R20334 a_n1996_n452.n56 a_n1996_n452.t5 2.82907
R20335 a_n1996_n452.n56 a_n1996_n452.t40 2.82907
R20336 a_n1996_n452.n89 a_n1996_n452.n76 1.30542
R20337 a_n1996_n452.n8 a_n1996_n452.n7 1.04595
R20338 a_n1996_n452.n25 a_n1996_n452.n69 13.657
R20339 a_n1996_n452.n67 a_n1996_n452.n33 21.4216
R20340 a_n1996_n452.n21 a_n1996_n452.n72 13.657
R20341 a_n1996_n452.n70 a_n1996_n452.n51 21.4216
R20342 a_n1996_n452.n93 a_n1996_n452.n15 13.657
R20343 a_n1996_n452.n42 a_n1996_n452.n95 21.4216
R20344 a_n1996_n452.n90 a_n1996_n452.n19 13.657
R20345 a_n1996_n452.n39 a_n1996_n452.n92 21.4216
R20346 a_n1996_n452.n3 a_n1996_n452.n2 1.3324
R20347 a_n1996_n452.n1 a_n1996_n452.n0 0.888431
R20348 a_n1996_n452.n24 a_n1996_n452.n22 0.758076
R20349 a_n1996_n452.n24 a_n1996_n452.n23 0.758076
R20350 a_n1996_n452.n34 a_n1996_n452.n20 0.758076
R20351 a_n1996_n452.n18 a_n1996_n452.n17 0.758076
R20352 a_n1996_n452.n17 a_n1996_n452.n16 0.758076
R20353 a_n1996_n452.n14 a_n1996_n452.n13 0.758076
R20354 a_n1996_n452.n13 a_n1996_n452.n12 0.758076
R20355 a_n1996_n452.n11 a_n1996_n452.n10 0.758076
R20356 a_n1996_n452.n9 a_n1996_n452.n8 0.758076
R20357 a_n1996_n452.n7 a_n1996_n452.n6 0.758076
R20358 a_n1996_n452.n5 a_n1996_n452.n4 0.758076
R20359 a_n1996_n452.n34 a_n1996_n452.n29 0.720197
R20360 a_n1996_n452.n28 a_n1996_n452.n27 0.716017
R20361 a_n1996_n452.n75 a_n1996_n452.n26 0.716017
R20362 a_n1996_n452.n10 a_n1996_n452.n9 0.67853
R20363 a_n1996_n452.n6 a_n1996_n452.n5 0.67853
R20364 a_n1986_8322.n6 a_n1986_8322.t14 74.6477
R20365 a_n1986_8322.n1 a_n1986_8322.t1 74.6477
R20366 a_n1986_8322.n16 a_n1986_8322.t10 74.6474
R20367 a_n1986_8322.n14 a_n1986_8322.t3 74.2899
R20368 a_n1986_8322.n7 a_n1986_8322.t12 74.2899
R20369 a_n1986_8322.n8 a_n1986_8322.t15 74.2899
R20370 a_n1986_8322.n11 a_n1986_8322.t16 74.2899
R20371 a_n1986_8322.n4 a_n1986_8322.t0 74.2899
R20372 a_n1986_8322.n16 a_n1986_8322.n15 70.6783
R20373 a_n1986_8322.n6 a_n1986_8322.n5 70.6783
R20374 a_n1986_8322.n10 a_n1986_8322.n9 70.6783
R20375 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R20376 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R20377 a_n1986_8322.n18 a_n1986_8322.n17 70.6782
R20378 a_n1986_8322.n12 a_n1986_8322.n4 22.7556
R20379 a_n1986_8322.n13 a_n1986_8322.t22 9.7972
R20380 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R20381 a_n1986_8322.n14 a_n1986_8322.n13 5.83671
R20382 a_n1986_8322.n13 a_n1986_8322.n12 5.3452
R20383 a_n1986_8322.n15 a_n1986_8322.t8 3.61217
R20384 a_n1986_8322.n15 a_n1986_8322.t5 3.61217
R20385 a_n1986_8322.n5 a_n1986_8322.t18 3.61217
R20386 a_n1986_8322.n5 a_n1986_8322.t17 3.61217
R20387 a_n1986_8322.n9 a_n1986_8322.t13 3.61217
R20388 a_n1986_8322.n9 a_n1986_8322.t19 3.61217
R20389 a_n1986_8322.n0 a_n1986_8322.t9 3.61217
R20390 a_n1986_8322.n0 a_n1986_8322.t4 3.61217
R20391 a_n1986_8322.n2 a_n1986_8322.t7 3.61217
R20392 a_n1986_8322.n2 a_n1986_8322.t6 3.61217
R20393 a_n1986_8322.n18 a_n1986_8322.t2 3.61217
R20394 a_n1986_8322.t11 a_n1986_8322.n18 3.61217
R20395 a_n1986_8322.n11 a_n1986_8322.n10 0.358259
R20396 a_n1986_8322.n10 a_n1986_8322.n8 0.358259
R20397 a_n1986_8322.n7 a_n1986_8322.n6 0.358259
R20398 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R20399 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R20400 a_n1986_8322.n17 a_n1986_8322.n14 0.358259
R20401 a_n1986_8322.n17 a_n1986_8322.n16 0.358259
R20402 a_n1986_8322.n8 a_n1986_8322.n7 0.101793
R20403 a_n1986_8322.t23 a_n1986_8322.t20 0.0788333
R20404 a_n1986_8322.t21 a_n1986_8322.t23 0.0631667
R20405 a_n1986_8322.t22 a_n1986_8322.t21 0.0471944
R20406 a_n1986_8322.t22 a_n1986_8322.t20 0.0453889
R20407 a_n1808_13878.n5 a_n1808_13878.n3 98.9633
R20408 a_n1808_13878.n2 a_n1808_13878.n0 98.7517
R20409 a_n1808_13878.n2 a_n1808_13878.n1 98.6055
R20410 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R20411 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R20412 a_n1808_13878.n7 a_n1808_13878.n6 98.6054
R20413 a_n1808_13878.n9 a_n1808_13878.t13 74.6477
R20414 a_n1808_13878.n14 a_n1808_13878.t14 74.2899
R20415 a_n1808_13878.n11 a_n1808_13878.t15 74.2899
R20416 a_n1808_13878.n10 a_n1808_13878.t12 74.2899
R20417 a_n1808_13878.n13 a_n1808_13878.n12 70.6783
R20418 a_n1808_13878.n9 a_n1808_13878.n8 70.6783
R20419 a_n1808_13878.n16 a_n1808_13878.n15 13.5694
R20420 a_n1808_13878.n15 a_n1808_13878.n7 11.5762
R20421 a_n1808_13878.n15 a_n1808_13878.n14 6.2408
R20422 a_n1808_13878.n1 a_n1808_13878.t6 3.61217
R20423 a_n1808_13878.n1 a_n1808_13878.t1 3.61217
R20424 a_n1808_13878.n0 a_n1808_13878.t0 3.61217
R20425 a_n1808_13878.n0 a_n1808_13878.t2 3.61217
R20426 a_n1808_13878.n6 a_n1808_13878.t7 3.61217
R20427 a_n1808_13878.n6 a_n1808_13878.t8 3.61217
R20428 a_n1808_13878.n4 a_n1808_13878.t10 3.61217
R20429 a_n1808_13878.n4 a_n1808_13878.t3 3.61217
R20430 a_n1808_13878.n3 a_n1808_13878.t5 3.61217
R20431 a_n1808_13878.n3 a_n1808_13878.t9 3.61217
R20432 a_n1808_13878.n12 a_n1808_13878.t18 3.61217
R20433 a_n1808_13878.n12 a_n1808_13878.t19 3.61217
R20434 a_n1808_13878.n8 a_n1808_13878.t16 3.61217
R20435 a_n1808_13878.n8 a_n1808_13878.t17 3.61217
R20436 a_n1808_13878.n17 a_n1808_13878.t4 3.61217
R20437 a_n1808_13878.t11 a_n1808_13878.n17 3.61217
R20438 a_n1808_13878.n7 a_n1808_13878.n5 0.358259
R20439 a_n1808_13878.n10 a_n1808_13878.n9 0.358259
R20440 a_n1808_13878.n13 a_n1808_13878.n11 0.358259
R20441 a_n1808_13878.n14 a_n1808_13878.n13 0.358259
R20442 a_n1808_13878.n16 a_n1808_13878.n2 0.146627
R20443 a_n1808_13878.n11 a_n1808_13878.n10 0.101793
R20444 outputibias.n27 outputibias.n1 289.615
R20445 outputibias.n58 outputibias.n32 289.615
R20446 outputibias.n90 outputibias.n64 289.615
R20447 outputibias.n122 outputibias.n96 289.615
R20448 outputibias.n28 outputibias.n27 185
R20449 outputibias.n26 outputibias.n25 185
R20450 outputibias.n5 outputibias.n4 185
R20451 outputibias.n20 outputibias.n19 185
R20452 outputibias.n18 outputibias.n17 185
R20453 outputibias.n9 outputibias.n8 185
R20454 outputibias.n12 outputibias.n11 185
R20455 outputibias.n59 outputibias.n58 185
R20456 outputibias.n57 outputibias.n56 185
R20457 outputibias.n36 outputibias.n35 185
R20458 outputibias.n51 outputibias.n50 185
R20459 outputibias.n49 outputibias.n48 185
R20460 outputibias.n40 outputibias.n39 185
R20461 outputibias.n43 outputibias.n42 185
R20462 outputibias.n91 outputibias.n90 185
R20463 outputibias.n89 outputibias.n88 185
R20464 outputibias.n68 outputibias.n67 185
R20465 outputibias.n83 outputibias.n82 185
R20466 outputibias.n81 outputibias.n80 185
R20467 outputibias.n72 outputibias.n71 185
R20468 outputibias.n75 outputibias.n74 185
R20469 outputibias.n123 outputibias.n122 185
R20470 outputibias.n121 outputibias.n120 185
R20471 outputibias.n100 outputibias.n99 185
R20472 outputibias.n115 outputibias.n114 185
R20473 outputibias.n113 outputibias.n112 185
R20474 outputibias.n104 outputibias.n103 185
R20475 outputibias.n107 outputibias.n106 185
R20476 outputibias.n0 outputibias.t9 178.945
R20477 outputibias.n133 outputibias.t8 177.018
R20478 outputibias.n132 outputibias.t11 177.018
R20479 outputibias.n0 outputibias.t10 177.018
R20480 outputibias.t5 outputibias.n10 147.661
R20481 outputibias.t7 outputibias.n41 147.661
R20482 outputibias.t1 outputibias.n73 147.661
R20483 outputibias.t3 outputibias.n105 147.661
R20484 outputibias.n128 outputibias.t4 132.363
R20485 outputibias.n128 outputibias.t6 130.436
R20486 outputibias.n129 outputibias.t0 130.436
R20487 outputibias.n130 outputibias.t2 130.436
R20488 outputibias.n27 outputibias.n26 104.615
R20489 outputibias.n26 outputibias.n4 104.615
R20490 outputibias.n19 outputibias.n4 104.615
R20491 outputibias.n19 outputibias.n18 104.615
R20492 outputibias.n18 outputibias.n8 104.615
R20493 outputibias.n11 outputibias.n8 104.615
R20494 outputibias.n58 outputibias.n57 104.615
R20495 outputibias.n57 outputibias.n35 104.615
R20496 outputibias.n50 outputibias.n35 104.615
R20497 outputibias.n50 outputibias.n49 104.615
R20498 outputibias.n49 outputibias.n39 104.615
R20499 outputibias.n42 outputibias.n39 104.615
R20500 outputibias.n90 outputibias.n89 104.615
R20501 outputibias.n89 outputibias.n67 104.615
R20502 outputibias.n82 outputibias.n67 104.615
R20503 outputibias.n82 outputibias.n81 104.615
R20504 outputibias.n81 outputibias.n71 104.615
R20505 outputibias.n74 outputibias.n71 104.615
R20506 outputibias.n122 outputibias.n121 104.615
R20507 outputibias.n121 outputibias.n99 104.615
R20508 outputibias.n114 outputibias.n99 104.615
R20509 outputibias.n114 outputibias.n113 104.615
R20510 outputibias.n113 outputibias.n103 104.615
R20511 outputibias.n106 outputibias.n103 104.615
R20512 outputibias.n63 outputibias.n31 95.6354
R20513 outputibias.n63 outputibias.n62 94.6732
R20514 outputibias.n95 outputibias.n94 94.6732
R20515 outputibias.n127 outputibias.n126 94.6732
R20516 outputibias.n11 outputibias.t5 52.3082
R20517 outputibias.n42 outputibias.t7 52.3082
R20518 outputibias.n74 outputibias.t1 52.3082
R20519 outputibias.n106 outputibias.t3 52.3082
R20520 outputibias.n12 outputibias.n10 15.6674
R20521 outputibias.n43 outputibias.n41 15.6674
R20522 outputibias.n75 outputibias.n73 15.6674
R20523 outputibias.n107 outputibias.n105 15.6674
R20524 outputibias.n13 outputibias.n9 12.8005
R20525 outputibias.n44 outputibias.n40 12.8005
R20526 outputibias.n76 outputibias.n72 12.8005
R20527 outputibias.n108 outputibias.n104 12.8005
R20528 outputibias.n17 outputibias.n16 12.0247
R20529 outputibias.n48 outputibias.n47 12.0247
R20530 outputibias.n80 outputibias.n79 12.0247
R20531 outputibias.n112 outputibias.n111 12.0247
R20532 outputibias.n20 outputibias.n7 11.249
R20533 outputibias.n51 outputibias.n38 11.249
R20534 outputibias.n83 outputibias.n70 11.249
R20535 outputibias.n115 outputibias.n102 11.249
R20536 outputibias.n21 outputibias.n5 10.4732
R20537 outputibias.n52 outputibias.n36 10.4732
R20538 outputibias.n84 outputibias.n68 10.4732
R20539 outputibias.n116 outputibias.n100 10.4732
R20540 outputibias.n25 outputibias.n24 9.69747
R20541 outputibias.n56 outputibias.n55 9.69747
R20542 outputibias.n88 outputibias.n87 9.69747
R20543 outputibias.n120 outputibias.n119 9.69747
R20544 outputibias.n31 outputibias.n30 9.45567
R20545 outputibias.n62 outputibias.n61 9.45567
R20546 outputibias.n94 outputibias.n93 9.45567
R20547 outputibias.n126 outputibias.n125 9.45567
R20548 outputibias.n30 outputibias.n29 9.3005
R20549 outputibias.n3 outputibias.n2 9.3005
R20550 outputibias.n24 outputibias.n23 9.3005
R20551 outputibias.n22 outputibias.n21 9.3005
R20552 outputibias.n7 outputibias.n6 9.3005
R20553 outputibias.n16 outputibias.n15 9.3005
R20554 outputibias.n14 outputibias.n13 9.3005
R20555 outputibias.n61 outputibias.n60 9.3005
R20556 outputibias.n34 outputibias.n33 9.3005
R20557 outputibias.n55 outputibias.n54 9.3005
R20558 outputibias.n53 outputibias.n52 9.3005
R20559 outputibias.n38 outputibias.n37 9.3005
R20560 outputibias.n47 outputibias.n46 9.3005
R20561 outputibias.n45 outputibias.n44 9.3005
R20562 outputibias.n93 outputibias.n92 9.3005
R20563 outputibias.n66 outputibias.n65 9.3005
R20564 outputibias.n87 outputibias.n86 9.3005
R20565 outputibias.n85 outputibias.n84 9.3005
R20566 outputibias.n70 outputibias.n69 9.3005
R20567 outputibias.n79 outputibias.n78 9.3005
R20568 outputibias.n77 outputibias.n76 9.3005
R20569 outputibias.n125 outputibias.n124 9.3005
R20570 outputibias.n98 outputibias.n97 9.3005
R20571 outputibias.n119 outputibias.n118 9.3005
R20572 outputibias.n117 outputibias.n116 9.3005
R20573 outputibias.n102 outputibias.n101 9.3005
R20574 outputibias.n111 outputibias.n110 9.3005
R20575 outputibias.n109 outputibias.n108 9.3005
R20576 outputibias.n28 outputibias.n3 8.92171
R20577 outputibias.n59 outputibias.n34 8.92171
R20578 outputibias.n91 outputibias.n66 8.92171
R20579 outputibias.n123 outputibias.n98 8.92171
R20580 outputibias.n29 outputibias.n1 8.14595
R20581 outputibias.n60 outputibias.n32 8.14595
R20582 outputibias.n92 outputibias.n64 8.14595
R20583 outputibias.n124 outputibias.n96 8.14595
R20584 outputibias.n31 outputibias.n1 5.81868
R20585 outputibias.n62 outputibias.n32 5.81868
R20586 outputibias.n94 outputibias.n64 5.81868
R20587 outputibias.n126 outputibias.n96 5.81868
R20588 outputibias.n131 outputibias.n130 5.20947
R20589 outputibias.n29 outputibias.n28 5.04292
R20590 outputibias.n60 outputibias.n59 5.04292
R20591 outputibias.n92 outputibias.n91 5.04292
R20592 outputibias.n124 outputibias.n123 5.04292
R20593 outputibias.n131 outputibias.n127 4.42209
R20594 outputibias.n14 outputibias.n10 4.38594
R20595 outputibias.n45 outputibias.n41 4.38594
R20596 outputibias.n77 outputibias.n73 4.38594
R20597 outputibias.n109 outputibias.n105 4.38594
R20598 outputibias.n132 outputibias.n131 4.28454
R20599 outputibias.n25 outputibias.n3 4.26717
R20600 outputibias.n56 outputibias.n34 4.26717
R20601 outputibias.n88 outputibias.n66 4.26717
R20602 outputibias.n120 outputibias.n98 4.26717
R20603 outputibias.n24 outputibias.n5 3.49141
R20604 outputibias.n55 outputibias.n36 3.49141
R20605 outputibias.n87 outputibias.n68 3.49141
R20606 outputibias.n119 outputibias.n100 3.49141
R20607 outputibias.n21 outputibias.n20 2.71565
R20608 outputibias.n52 outputibias.n51 2.71565
R20609 outputibias.n84 outputibias.n83 2.71565
R20610 outputibias.n116 outputibias.n115 2.71565
R20611 outputibias.n17 outputibias.n7 1.93989
R20612 outputibias.n48 outputibias.n38 1.93989
R20613 outputibias.n80 outputibias.n70 1.93989
R20614 outputibias.n112 outputibias.n102 1.93989
R20615 outputibias.n130 outputibias.n129 1.9266
R20616 outputibias.n129 outputibias.n128 1.9266
R20617 outputibias.n133 outputibias.n132 1.92658
R20618 outputibias.n134 outputibias.n133 1.29913
R20619 outputibias.n16 outputibias.n9 1.16414
R20620 outputibias.n47 outputibias.n40 1.16414
R20621 outputibias.n79 outputibias.n72 1.16414
R20622 outputibias.n111 outputibias.n104 1.16414
R20623 outputibias.n127 outputibias.n95 0.962709
R20624 outputibias.n95 outputibias.n63 0.962709
R20625 outputibias.n13 outputibias.n12 0.388379
R20626 outputibias.n44 outputibias.n43 0.388379
R20627 outputibias.n76 outputibias.n75 0.388379
R20628 outputibias.n108 outputibias.n107 0.388379
R20629 outputibias.n134 outputibias.n0 0.337251
R20630 outputibias outputibias.n134 0.302375
R20631 outputibias.n30 outputibias.n2 0.155672
R20632 outputibias.n23 outputibias.n2 0.155672
R20633 outputibias.n23 outputibias.n22 0.155672
R20634 outputibias.n22 outputibias.n6 0.155672
R20635 outputibias.n15 outputibias.n6 0.155672
R20636 outputibias.n15 outputibias.n14 0.155672
R20637 outputibias.n61 outputibias.n33 0.155672
R20638 outputibias.n54 outputibias.n33 0.155672
R20639 outputibias.n54 outputibias.n53 0.155672
R20640 outputibias.n53 outputibias.n37 0.155672
R20641 outputibias.n46 outputibias.n37 0.155672
R20642 outputibias.n46 outputibias.n45 0.155672
R20643 outputibias.n93 outputibias.n65 0.155672
R20644 outputibias.n86 outputibias.n65 0.155672
R20645 outputibias.n86 outputibias.n85 0.155672
R20646 outputibias.n85 outputibias.n69 0.155672
R20647 outputibias.n78 outputibias.n69 0.155672
R20648 outputibias.n78 outputibias.n77 0.155672
R20649 outputibias.n125 outputibias.n97 0.155672
R20650 outputibias.n118 outputibias.n97 0.155672
R20651 outputibias.n118 outputibias.n117 0.155672
R20652 outputibias.n117 outputibias.n101 0.155672
R20653 outputibias.n110 outputibias.n101 0.155672
R20654 outputibias.n110 outputibias.n109 0.155672
R20655 output.n41 output.n15 289.615
R20656 output.n72 output.n46 289.615
R20657 output.n104 output.n78 289.615
R20658 output.n136 output.n110 289.615
R20659 output.n77 output.n45 197.26
R20660 output.n77 output.n76 196.298
R20661 output.n109 output.n108 196.298
R20662 output.n141 output.n140 196.298
R20663 output.n42 output.n41 185
R20664 output.n40 output.n39 185
R20665 output.n19 output.n18 185
R20666 output.n34 output.n33 185
R20667 output.n32 output.n31 185
R20668 output.n23 output.n22 185
R20669 output.n26 output.n25 185
R20670 output.n73 output.n72 185
R20671 output.n71 output.n70 185
R20672 output.n50 output.n49 185
R20673 output.n65 output.n64 185
R20674 output.n63 output.n62 185
R20675 output.n54 output.n53 185
R20676 output.n57 output.n56 185
R20677 output.n105 output.n104 185
R20678 output.n103 output.n102 185
R20679 output.n82 output.n81 185
R20680 output.n97 output.n96 185
R20681 output.n95 output.n94 185
R20682 output.n86 output.n85 185
R20683 output.n89 output.n88 185
R20684 output.n137 output.n136 185
R20685 output.n135 output.n134 185
R20686 output.n114 output.n113 185
R20687 output.n129 output.n128 185
R20688 output.n127 output.n126 185
R20689 output.n118 output.n117 185
R20690 output.n121 output.n120 185
R20691 output.t2 output.n24 147.661
R20692 output.t1 output.n55 147.661
R20693 output.t3 output.n87 147.661
R20694 output.t0 output.n119 147.661
R20695 output.n41 output.n40 104.615
R20696 output.n40 output.n18 104.615
R20697 output.n33 output.n18 104.615
R20698 output.n33 output.n32 104.615
R20699 output.n32 output.n22 104.615
R20700 output.n25 output.n22 104.615
R20701 output.n72 output.n71 104.615
R20702 output.n71 output.n49 104.615
R20703 output.n64 output.n49 104.615
R20704 output.n64 output.n63 104.615
R20705 output.n63 output.n53 104.615
R20706 output.n56 output.n53 104.615
R20707 output.n104 output.n103 104.615
R20708 output.n103 output.n81 104.615
R20709 output.n96 output.n81 104.615
R20710 output.n96 output.n95 104.615
R20711 output.n95 output.n85 104.615
R20712 output.n88 output.n85 104.615
R20713 output.n136 output.n135 104.615
R20714 output.n135 output.n113 104.615
R20715 output.n128 output.n113 104.615
R20716 output.n128 output.n127 104.615
R20717 output.n127 output.n117 104.615
R20718 output.n120 output.n117 104.615
R20719 output.n1 output.t9 77.056
R20720 output.n14 output.t10 76.6694
R20721 output.n1 output.n0 72.7095
R20722 output.n3 output.n2 72.7095
R20723 output.n5 output.n4 72.7095
R20724 output.n7 output.n6 72.7095
R20725 output.n9 output.n8 72.7095
R20726 output.n11 output.n10 72.7095
R20727 output.n13 output.n12 72.7095
R20728 output.n25 output.t2 52.3082
R20729 output.n56 output.t1 52.3082
R20730 output.n88 output.t3 52.3082
R20731 output.n120 output.t0 52.3082
R20732 output.n26 output.n24 15.6674
R20733 output.n57 output.n55 15.6674
R20734 output.n89 output.n87 15.6674
R20735 output.n121 output.n119 15.6674
R20736 output.n27 output.n23 12.8005
R20737 output.n58 output.n54 12.8005
R20738 output.n90 output.n86 12.8005
R20739 output.n122 output.n118 12.8005
R20740 output.n31 output.n30 12.0247
R20741 output.n62 output.n61 12.0247
R20742 output.n94 output.n93 12.0247
R20743 output.n126 output.n125 12.0247
R20744 output.n34 output.n21 11.249
R20745 output.n65 output.n52 11.249
R20746 output.n97 output.n84 11.249
R20747 output.n129 output.n116 11.249
R20748 output.n35 output.n19 10.4732
R20749 output.n66 output.n50 10.4732
R20750 output.n98 output.n82 10.4732
R20751 output.n130 output.n114 10.4732
R20752 output.n39 output.n38 9.69747
R20753 output.n70 output.n69 9.69747
R20754 output.n102 output.n101 9.69747
R20755 output.n134 output.n133 9.69747
R20756 output.n45 output.n44 9.45567
R20757 output.n76 output.n75 9.45567
R20758 output.n108 output.n107 9.45567
R20759 output.n140 output.n139 9.45567
R20760 output.n44 output.n43 9.3005
R20761 output.n17 output.n16 9.3005
R20762 output.n38 output.n37 9.3005
R20763 output.n36 output.n35 9.3005
R20764 output.n21 output.n20 9.3005
R20765 output.n30 output.n29 9.3005
R20766 output.n28 output.n27 9.3005
R20767 output.n75 output.n74 9.3005
R20768 output.n48 output.n47 9.3005
R20769 output.n69 output.n68 9.3005
R20770 output.n67 output.n66 9.3005
R20771 output.n52 output.n51 9.3005
R20772 output.n61 output.n60 9.3005
R20773 output.n59 output.n58 9.3005
R20774 output.n107 output.n106 9.3005
R20775 output.n80 output.n79 9.3005
R20776 output.n101 output.n100 9.3005
R20777 output.n99 output.n98 9.3005
R20778 output.n84 output.n83 9.3005
R20779 output.n93 output.n92 9.3005
R20780 output.n91 output.n90 9.3005
R20781 output.n139 output.n138 9.3005
R20782 output.n112 output.n111 9.3005
R20783 output.n133 output.n132 9.3005
R20784 output.n131 output.n130 9.3005
R20785 output.n116 output.n115 9.3005
R20786 output.n125 output.n124 9.3005
R20787 output.n123 output.n122 9.3005
R20788 output.n42 output.n17 8.92171
R20789 output.n73 output.n48 8.92171
R20790 output.n105 output.n80 8.92171
R20791 output.n137 output.n112 8.92171
R20792 output output.n141 8.15037
R20793 output.n43 output.n15 8.14595
R20794 output.n74 output.n46 8.14595
R20795 output.n106 output.n78 8.14595
R20796 output.n138 output.n110 8.14595
R20797 output.n45 output.n15 5.81868
R20798 output.n76 output.n46 5.81868
R20799 output.n108 output.n78 5.81868
R20800 output.n140 output.n110 5.81868
R20801 output.n43 output.n42 5.04292
R20802 output.n74 output.n73 5.04292
R20803 output.n106 output.n105 5.04292
R20804 output.n138 output.n137 5.04292
R20805 output.n28 output.n24 4.38594
R20806 output.n59 output.n55 4.38594
R20807 output.n91 output.n87 4.38594
R20808 output.n123 output.n119 4.38594
R20809 output.n39 output.n17 4.26717
R20810 output.n70 output.n48 4.26717
R20811 output.n102 output.n80 4.26717
R20812 output.n134 output.n112 4.26717
R20813 output.n0 output.t15 3.9605
R20814 output.n0 output.t19 3.9605
R20815 output.n2 output.t7 3.9605
R20816 output.n2 output.t11 3.9605
R20817 output.n4 output.t12 3.9605
R20818 output.n4 output.t17 3.9605
R20819 output.n6 output.t5 3.9605
R20820 output.n6 output.t13 3.9605
R20821 output.n8 output.t16 3.9605
R20822 output.n8 output.t14 3.9605
R20823 output.n10 output.t4 3.9605
R20824 output.n10 output.t6 3.9605
R20825 output.n12 output.t8 3.9605
R20826 output.n12 output.t18 3.9605
R20827 output.n38 output.n19 3.49141
R20828 output.n69 output.n50 3.49141
R20829 output.n101 output.n82 3.49141
R20830 output.n133 output.n114 3.49141
R20831 output.n35 output.n34 2.71565
R20832 output.n66 output.n65 2.71565
R20833 output.n98 output.n97 2.71565
R20834 output.n130 output.n129 2.71565
R20835 output.n31 output.n21 1.93989
R20836 output.n62 output.n52 1.93989
R20837 output.n94 output.n84 1.93989
R20838 output.n126 output.n116 1.93989
R20839 output.n30 output.n23 1.16414
R20840 output.n61 output.n54 1.16414
R20841 output.n93 output.n86 1.16414
R20842 output.n125 output.n118 1.16414
R20843 output.n141 output.n109 0.962709
R20844 output.n109 output.n77 0.962709
R20845 output.n27 output.n26 0.388379
R20846 output.n58 output.n57 0.388379
R20847 output.n90 output.n89 0.388379
R20848 output.n122 output.n121 0.388379
R20849 output.n14 output.n13 0.387128
R20850 output.n13 output.n11 0.387128
R20851 output.n11 output.n9 0.387128
R20852 output.n9 output.n7 0.387128
R20853 output.n7 output.n5 0.387128
R20854 output.n5 output.n3 0.387128
R20855 output.n3 output.n1 0.387128
R20856 output.n44 output.n16 0.155672
R20857 output.n37 output.n16 0.155672
R20858 output.n37 output.n36 0.155672
R20859 output.n36 output.n20 0.155672
R20860 output.n29 output.n20 0.155672
R20861 output.n29 output.n28 0.155672
R20862 output.n75 output.n47 0.155672
R20863 output.n68 output.n47 0.155672
R20864 output.n68 output.n67 0.155672
R20865 output.n67 output.n51 0.155672
R20866 output.n60 output.n51 0.155672
R20867 output.n60 output.n59 0.155672
R20868 output.n107 output.n79 0.155672
R20869 output.n100 output.n79 0.155672
R20870 output.n100 output.n99 0.155672
R20871 output.n99 output.n83 0.155672
R20872 output.n92 output.n83 0.155672
R20873 output.n92 output.n91 0.155672
R20874 output.n139 output.n111 0.155672
R20875 output.n132 output.n111 0.155672
R20876 output.n132 output.n131 0.155672
R20877 output.n131 output.n115 0.155672
R20878 output.n124 output.n115 0.155672
R20879 output.n124 output.n123 0.155672
R20880 output output.n14 0.126227
R20881 minus.n43 minus.t24 322.512
R20882 minus.n9 minus.t8 322.512
R20883 minus.n66 minus.t5 297.12
R20884 minus.n64 minus.t6 297.12
R20885 minus.n36 minus.t22 297.12
R20886 minus.n58 minus.t18 297.12
R20887 minus.n38 minus.t19 297.12
R20888 minus.n52 minus.t14 297.12
R20889 minus.n40 minus.t15 297.12
R20890 minus.n46 minus.t9 297.12
R20891 minus.n42 minus.t23 297.12
R20892 minus.n8 minus.t7 297.12
R20893 minus.n12 minus.t11 297.12
R20894 minus.n14 minus.t10 297.12
R20895 minus.n18 minus.t12 297.12
R20896 minus.n20 minus.t17 297.12
R20897 minus.n24 minus.t16 297.12
R20898 minus.n26 minus.t21 297.12
R20899 minus.n30 minus.t20 297.12
R20900 minus.n32 minus.t13 297.12
R20901 minus.n72 minus.t4 243.255
R20902 minus.n71 minus.n69 224.169
R20903 minus.n71 minus.n70 223.454
R20904 minus.n45 minus.n44 161.3
R20905 minus.n46 minus.n41 161.3
R20906 minus.n48 minus.n47 161.3
R20907 minus.n49 minus.n40 161.3
R20908 minus.n51 minus.n50 161.3
R20909 minus.n52 minus.n39 161.3
R20910 minus.n54 minus.n53 161.3
R20911 minus.n55 minus.n38 161.3
R20912 minus.n57 minus.n56 161.3
R20913 minus.n58 minus.n37 161.3
R20914 minus.n60 minus.n59 161.3
R20915 minus.n61 minus.n36 161.3
R20916 minus.n63 minus.n62 161.3
R20917 minus.n64 minus.n35 161.3
R20918 minus.n65 minus.n34 161.3
R20919 minus.n67 minus.n66 161.3
R20920 minus.n33 minus.n32 161.3
R20921 minus.n31 minus.n0 161.3
R20922 minus.n30 minus.n29 161.3
R20923 minus.n28 minus.n1 161.3
R20924 minus.n27 minus.n26 161.3
R20925 minus.n25 minus.n2 161.3
R20926 minus.n24 minus.n23 161.3
R20927 minus.n22 minus.n3 161.3
R20928 minus.n21 minus.n20 161.3
R20929 minus.n19 minus.n4 161.3
R20930 minus.n18 minus.n17 161.3
R20931 minus.n16 minus.n5 161.3
R20932 minus.n15 minus.n14 161.3
R20933 minus.n13 minus.n6 161.3
R20934 minus.n12 minus.n11 161.3
R20935 minus.n10 minus.n7 161.3
R20936 minus.n44 minus.n43 45.0031
R20937 minus.n10 minus.n9 45.0031
R20938 minus.n66 minus.n65 41.6278
R20939 minus.n32 minus.n31 41.6278
R20940 minus.n64 minus.n63 37.246
R20941 minus.n45 minus.n42 37.246
R20942 minus.n8 minus.n7 37.246
R20943 minus.n30 minus.n1 37.246
R20944 minus.n59 minus.n36 32.8641
R20945 minus.n47 minus.n46 32.8641
R20946 minus.n13 minus.n12 32.8641
R20947 minus.n26 minus.n25 32.8641
R20948 minus.n68 minus.n67 31.8206
R20949 minus.n58 minus.n57 28.4823
R20950 minus.n51 minus.n40 28.4823
R20951 minus.n14 minus.n5 28.4823
R20952 minus.n24 minus.n3 28.4823
R20953 minus.n53 minus.n38 24.1005
R20954 minus.n53 minus.n52 24.1005
R20955 minus.n19 minus.n18 24.1005
R20956 minus.n20 minus.n19 24.1005
R20957 minus.n70 minus.t3 19.8005
R20958 minus.n70 minus.t1 19.8005
R20959 minus.n69 minus.t2 19.8005
R20960 minus.n69 minus.t0 19.8005
R20961 minus.n57 minus.n38 19.7187
R20962 minus.n52 minus.n51 19.7187
R20963 minus.n18 minus.n5 19.7187
R20964 minus.n20 minus.n3 19.7187
R20965 minus.n43 minus.n42 15.6319
R20966 minus.n9 minus.n8 15.6319
R20967 minus.n59 minus.n58 15.3369
R20968 minus.n47 minus.n40 15.3369
R20969 minus.n14 minus.n13 15.3369
R20970 minus.n25 minus.n24 15.3369
R20971 minus.n68 minus.n33 12.0819
R20972 minus minus.n73 11.2074
R20973 minus.n63 minus.n36 10.955
R20974 minus.n46 minus.n45 10.955
R20975 minus.n12 minus.n7 10.955
R20976 minus.n26 minus.n1 10.955
R20977 minus.n65 minus.n64 6.57323
R20978 minus.n31 minus.n30 6.57323
R20979 minus.n73 minus.n72 4.80222
R20980 minus.n73 minus.n68 0.972091
R20981 minus.n72 minus.n71 0.716017
R20982 minus.n67 minus.n34 0.189894
R20983 minus.n35 minus.n34 0.189894
R20984 minus.n62 minus.n35 0.189894
R20985 minus.n62 minus.n61 0.189894
R20986 minus.n61 minus.n60 0.189894
R20987 minus.n60 minus.n37 0.189894
R20988 minus.n56 minus.n37 0.189894
R20989 minus.n56 minus.n55 0.189894
R20990 minus.n55 minus.n54 0.189894
R20991 minus.n54 minus.n39 0.189894
R20992 minus.n50 minus.n39 0.189894
R20993 minus.n50 minus.n49 0.189894
R20994 minus.n49 minus.n48 0.189894
R20995 minus.n48 minus.n41 0.189894
R20996 minus.n44 minus.n41 0.189894
R20997 minus.n11 minus.n10 0.189894
R20998 minus.n11 minus.n6 0.189894
R20999 minus.n15 minus.n6 0.189894
R21000 minus.n16 minus.n15 0.189894
R21001 minus.n17 minus.n16 0.189894
R21002 minus.n17 minus.n4 0.189894
R21003 minus.n21 minus.n4 0.189894
R21004 minus.n22 minus.n21 0.189894
R21005 minus.n23 minus.n22 0.189894
R21006 minus.n23 minus.n2 0.189894
R21007 minus.n27 minus.n2 0.189894
R21008 minus.n28 minus.n27 0.189894
R21009 minus.n29 minus.n28 0.189894
R21010 minus.n29 minus.n0 0.189894
R21011 minus.n33 minus.n0 0.189894
R21012 diffpairibias.n0 diffpairibias.t18 436.822
R21013 diffpairibias.n21 diffpairibias.t19 435.479
R21014 diffpairibias.n20 diffpairibias.t16 435.479
R21015 diffpairibias.n19 diffpairibias.t17 435.479
R21016 diffpairibias.n18 diffpairibias.t21 435.479
R21017 diffpairibias.n0 diffpairibias.t22 435.479
R21018 diffpairibias.n1 diffpairibias.t20 435.479
R21019 diffpairibias.n2 diffpairibias.t23 435.479
R21020 diffpairibias.n10 diffpairibias.t0 377.536
R21021 diffpairibias.n10 diffpairibias.t8 376.193
R21022 diffpairibias.n11 diffpairibias.t10 376.193
R21023 diffpairibias.n12 diffpairibias.t6 376.193
R21024 diffpairibias.n13 diffpairibias.t2 376.193
R21025 diffpairibias.n14 diffpairibias.t12 376.193
R21026 diffpairibias.n15 diffpairibias.t4 376.193
R21027 diffpairibias.n16 diffpairibias.t14 376.193
R21028 diffpairibias.n3 diffpairibias.t1 113.368
R21029 diffpairibias.n3 diffpairibias.t9 112.698
R21030 diffpairibias.n4 diffpairibias.t11 112.698
R21031 diffpairibias.n5 diffpairibias.t7 112.698
R21032 diffpairibias.n6 diffpairibias.t3 112.698
R21033 diffpairibias.n7 diffpairibias.t13 112.698
R21034 diffpairibias.n8 diffpairibias.t5 112.698
R21035 diffpairibias.n9 diffpairibias.t15 112.698
R21036 diffpairibias.n17 diffpairibias.n16 4.77242
R21037 diffpairibias.n17 diffpairibias.n9 4.30807
R21038 diffpairibias.n18 diffpairibias.n17 4.13945
R21039 diffpairibias.n16 diffpairibias.n15 1.34352
R21040 diffpairibias.n15 diffpairibias.n14 1.34352
R21041 diffpairibias.n14 diffpairibias.n13 1.34352
R21042 diffpairibias.n13 diffpairibias.n12 1.34352
R21043 diffpairibias.n12 diffpairibias.n11 1.34352
R21044 diffpairibias.n11 diffpairibias.n10 1.34352
R21045 diffpairibias.n2 diffpairibias.n1 1.34352
R21046 diffpairibias.n1 diffpairibias.n0 1.34352
R21047 diffpairibias.n19 diffpairibias.n18 1.34352
R21048 diffpairibias.n20 diffpairibias.n19 1.34352
R21049 diffpairibias.n21 diffpairibias.n20 1.34352
R21050 diffpairibias.n22 diffpairibias.n21 0.862419
R21051 diffpairibias diffpairibias.n22 0.684875
R21052 diffpairibias.n9 diffpairibias.n8 0.672012
R21053 diffpairibias.n8 diffpairibias.n7 0.672012
R21054 diffpairibias.n7 diffpairibias.n6 0.672012
R21055 diffpairibias.n6 diffpairibias.n5 0.672012
R21056 diffpairibias.n5 diffpairibias.n4 0.672012
R21057 diffpairibias.n4 diffpairibias.n3 0.672012
R21058 diffpairibias.n22 diffpairibias.n2 0.190907
C0 commonsourceibias outputibias 0.003832f
C1 plus diffpairibias 3.42e-19
C2 vdd commonsourceibias 0.004218f
C3 CSoutput plus 0.839035f
C4 commonsourceibias diffpairibias 0.06482f
C5 CSoutput commonsourceibias 41.846302f
C6 minus plus 8.845019f
C7 minus commonsourceibias 0.323913f
C8 plus commonsourceibias 0.278362f
C9 output outputibias 2.34152f
C10 vdd output 7.23429f
C11 CSoutput output 6.13881f
C12 CSoutput outputibias 0.032386f
C13 vdd CSoutput 67.6707f
C14 minus diffpairibias 3.4e-19
C15 commonsourceibias output 0.006808f
C16 CSoutput minus 2.48853f
C17 vdd plus 0.066355f
C18 diffpairibias gnd 48.980137f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.144416p
C22 plus gnd 32.641903f
C23 minus gnd 26.354519f
C24 CSoutput gnd 0.107008p
C25 vdd gnd 0.344772p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 minus.n0 gnd 0.032421f
C74 minus.n1 gnd 0.007357f
C75 minus.n2 gnd 0.032421f
C76 minus.n3 gnd 0.007357f
C77 minus.n4 gnd 0.032421f
C78 minus.n5 gnd 0.007357f
C79 minus.n6 gnd 0.032421f
C80 minus.n7 gnd 0.007357f
C81 minus.t8 gnd 0.474624f
C82 minus.t7 gnd 0.458559f
C83 minus.n8 gnd 0.209129f
C84 minus.n9 gnd 0.189969f
C85 minus.n10 gnd 0.138384f
C86 minus.n11 gnd 0.032421f
C87 minus.t11 gnd 0.458559f
C88 minus.n12 gnd 0.203706f
C89 minus.n13 gnd 0.007357f
C90 minus.t10 gnd 0.458559f
C91 minus.n14 gnd 0.203706f
C92 minus.n15 gnd 0.032421f
C93 minus.n16 gnd 0.032421f
C94 minus.n17 gnd 0.032421f
C95 minus.t12 gnd 0.458559f
C96 minus.n18 gnd 0.203706f
C97 minus.n19 gnd 0.007357f
C98 minus.t17 gnd 0.458559f
C99 minus.n20 gnd 0.203706f
C100 minus.n21 gnd 0.032421f
C101 minus.n22 gnd 0.032421f
C102 minus.n23 gnd 0.032421f
C103 minus.t16 gnd 0.458559f
C104 minus.n24 gnd 0.203706f
C105 minus.n25 gnd 0.007357f
C106 minus.t21 gnd 0.458559f
C107 minus.n26 gnd 0.203706f
C108 minus.n27 gnd 0.032421f
C109 minus.n28 gnd 0.032421f
C110 minus.n29 gnd 0.032421f
C111 minus.t20 gnd 0.458559f
C112 minus.n30 gnd 0.203706f
C113 minus.n31 gnd 0.007357f
C114 minus.t13 gnd 0.458559f
C115 minus.n32 gnd 0.203407f
C116 minus.n33 gnd 0.374594f
C117 minus.n34 gnd 0.032421f
C118 minus.t5 gnd 0.458559f
C119 minus.t6 gnd 0.458559f
C120 minus.n35 gnd 0.032421f
C121 minus.t22 gnd 0.458559f
C122 minus.n36 gnd 0.203706f
C123 minus.n37 gnd 0.032421f
C124 minus.t18 gnd 0.458559f
C125 minus.t19 gnd 0.458559f
C126 minus.n38 gnd 0.203706f
C127 minus.n39 gnd 0.032421f
C128 minus.t14 gnd 0.458559f
C129 minus.t15 gnd 0.458559f
C130 minus.n40 gnd 0.203706f
C131 minus.n41 gnd 0.032421f
C132 minus.t9 gnd 0.458559f
C133 minus.t23 gnd 0.458559f
C134 minus.n42 gnd 0.209129f
C135 minus.t24 gnd 0.474624f
C136 minus.n43 gnd 0.189969f
C137 minus.n44 gnd 0.138384f
C138 minus.n45 gnd 0.007357f
C139 minus.n46 gnd 0.203706f
C140 minus.n47 gnd 0.007357f
C141 minus.n48 gnd 0.032421f
C142 minus.n49 gnd 0.032421f
C143 minus.n50 gnd 0.032421f
C144 minus.n51 gnd 0.007357f
C145 minus.n52 gnd 0.203706f
C146 minus.n53 gnd 0.007357f
C147 minus.n54 gnd 0.032421f
C148 minus.n55 gnd 0.032421f
C149 minus.n56 gnd 0.032421f
C150 minus.n57 gnd 0.007357f
C151 minus.n58 gnd 0.203706f
C152 minus.n59 gnd 0.007357f
C153 minus.n60 gnd 0.032421f
C154 minus.n61 gnd 0.032421f
C155 minus.n62 gnd 0.032421f
C156 minus.n63 gnd 0.007357f
C157 minus.n64 gnd 0.203706f
C158 minus.n65 gnd 0.007357f
C159 minus.n66 gnd 0.203407f
C160 minus.n67 gnd 1.01305f
C161 minus.n68 gnd 1.52513f
C162 minus.t2 gnd 0.009994f
C163 minus.t0 gnd 0.009994f
C164 minus.n69 gnd 0.032864f
C165 minus.t3 gnd 0.009994f
C166 minus.t1 gnd 0.009994f
C167 minus.n70 gnd 0.032413f
C168 minus.n71 gnd 0.276633f
C169 minus.t4 gnd 0.055627f
C170 minus.n72 gnd 0.150956f
C171 minus.n73 gnd 1.81817f
C172 output.t9 gnd 0.464308f
C173 output.t15 gnd 0.044422f
C174 output.t19 gnd 0.044422f
C175 output.n0 gnd 0.364624f
C176 output.n1 gnd 0.614102f
C177 output.t7 gnd 0.044422f
C178 output.t11 gnd 0.044422f
C179 output.n2 gnd 0.364624f
C180 output.n3 gnd 0.350265f
C181 output.t12 gnd 0.044422f
C182 output.t17 gnd 0.044422f
C183 output.n4 gnd 0.364624f
C184 output.n5 gnd 0.350265f
C185 output.t5 gnd 0.044422f
C186 output.t13 gnd 0.044422f
C187 output.n6 gnd 0.364624f
C188 output.n7 gnd 0.350265f
C189 output.t16 gnd 0.044422f
C190 output.t14 gnd 0.044422f
C191 output.n8 gnd 0.364624f
C192 output.n9 gnd 0.350265f
C193 output.t4 gnd 0.044422f
C194 output.t6 gnd 0.044422f
C195 output.n10 gnd 0.364624f
C196 output.n11 gnd 0.350265f
C197 output.t8 gnd 0.044422f
C198 output.t18 gnd 0.044422f
C199 output.n12 gnd 0.364624f
C200 output.n13 gnd 0.350265f
C201 output.t10 gnd 0.462979f
C202 output.n14 gnd 0.28994f
C203 output.n15 gnd 0.015803f
C204 output.n16 gnd 0.011243f
C205 output.n17 gnd 0.006041f
C206 output.n18 gnd 0.01428f
C207 output.n19 gnd 0.006397f
C208 output.n20 gnd 0.011243f
C209 output.n21 gnd 0.006041f
C210 output.n22 gnd 0.01428f
C211 output.n23 gnd 0.006397f
C212 output.n24 gnd 0.048111f
C213 output.t2 gnd 0.023274f
C214 output.n25 gnd 0.01071f
C215 output.n26 gnd 0.008435f
C216 output.n27 gnd 0.006041f
C217 output.n28 gnd 0.267512f
C218 output.n29 gnd 0.011243f
C219 output.n30 gnd 0.006041f
C220 output.n31 gnd 0.006397f
C221 output.n32 gnd 0.01428f
C222 output.n33 gnd 0.01428f
C223 output.n34 gnd 0.006397f
C224 output.n35 gnd 0.006041f
C225 output.n36 gnd 0.011243f
C226 output.n37 gnd 0.011243f
C227 output.n38 gnd 0.006041f
C228 output.n39 gnd 0.006397f
C229 output.n40 gnd 0.01428f
C230 output.n41 gnd 0.030913f
C231 output.n42 gnd 0.006397f
C232 output.n43 gnd 0.006041f
C233 output.n44 gnd 0.025987f
C234 output.n45 gnd 0.097665f
C235 output.n46 gnd 0.015803f
C236 output.n47 gnd 0.011243f
C237 output.n48 gnd 0.006041f
C238 output.n49 gnd 0.01428f
C239 output.n50 gnd 0.006397f
C240 output.n51 gnd 0.011243f
C241 output.n52 gnd 0.006041f
C242 output.n53 gnd 0.01428f
C243 output.n54 gnd 0.006397f
C244 output.n55 gnd 0.048111f
C245 output.t1 gnd 0.023274f
C246 output.n56 gnd 0.01071f
C247 output.n57 gnd 0.008435f
C248 output.n58 gnd 0.006041f
C249 output.n59 gnd 0.267512f
C250 output.n60 gnd 0.011243f
C251 output.n61 gnd 0.006041f
C252 output.n62 gnd 0.006397f
C253 output.n63 gnd 0.01428f
C254 output.n64 gnd 0.01428f
C255 output.n65 gnd 0.006397f
C256 output.n66 gnd 0.006041f
C257 output.n67 gnd 0.011243f
C258 output.n68 gnd 0.011243f
C259 output.n69 gnd 0.006041f
C260 output.n70 gnd 0.006397f
C261 output.n71 gnd 0.01428f
C262 output.n72 gnd 0.030913f
C263 output.n73 gnd 0.006397f
C264 output.n74 gnd 0.006041f
C265 output.n75 gnd 0.025987f
C266 output.n76 gnd 0.09306f
C267 output.n77 gnd 1.65264f
C268 output.n78 gnd 0.015803f
C269 output.n79 gnd 0.011243f
C270 output.n80 gnd 0.006041f
C271 output.n81 gnd 0.01428f
C272 output.n82 gnd 0.006397f
C273 output.n83 gnd 0.011243f
C274 output.n84 gnd 0.006041f
C275 output.n85 gnd 0.01428f
C276 output.n86 gnd 0.006397f
C277 output.n87 gnd 0.048111f
C278 output.t3 gnd 0.023274f
C279 output.n88 gnd 0.01071f
C280 output.n89 gnd 0.008435f
C281 output.n90 gnd 0.006041f
C282 output.n91 gnd 0.267512f
C283 output.n92 gnd 0.011243f
C284 output.n93 gnd 0.006041f
C285 output.n94 gnd 0.006397f
C286 output.n95 gnd 0.01428f
C287 output.n96 gnd 0.01428f
C288 output.n97 gnd 0.006397f
C289 output.n98 gnd 0.006041f
C290 output.n99 gnd 0.011243f
C291 output.n100 gnd 0.011243f
C292 output.n101 gnd 0.006041f
C293 output.n102 gnd 0.006397f
C294 output.n103 gnd 0.01428f
C295 output.n104 gnd 0.030913f
C296 output.n105 gnd 0.006397f
C297 output.n106 gnd 0.006041f
C298 output.n107 gnd 0.025987f
C299 output.n108 gnd 0.09306f
C300 output.n109 gnd 0.713089f
C301 output.n110 gnd 0.015803f
C302 output.n111 gnd 0.011243f
C303 output.n112 gnd 0.006041f
C304 output.n113 gnd 0.01428f
C305 output.n114 gnd 0.006397f
C306 output.n115 gnd 0.011243f
C307 output.n116 gnd 0.006041f
C308 output.n117 gnd 0.01428f
C309 output.n118 gnd 0.006397f
C310 output.n119 gnd 0.048111f
C311 output.t0 gnd 0.023274f
C312 output.n120 gnd 0.01071f
C313 output.n121 gnd 0.008435f
C314 output.n122 gnd 0.006041f
C315 output.n123 gnd 0.267512f
C316 output.n124 gnd 0.011243f
C317 output.n125 gnd 0.006041f
C318 output.n126 gnd 0.006397f
C319 output.n127 gnd 0.01428f
C320 output.n128 gnd 0.01428f
C321 output.n129 gnd 0.006397f
C322 output.n130 gnd 0.006041f
C323 output.n131 gnd 0.011243f
C324 output.n132 gnd 0.011243f
C325 output.n133 gnd 0.006041f
C326 output.n134 gnd 0.006397f
C327 output.n135 gnd 0.01428f
C328 output.n136 gnd 0.030913f
C329 output.n137 gnd 0.006397f
C330 output.n138 gnd 0.006041f
C331 output.n139 gnd 0.025987f
C332 output.n140 gnd 0.09306f
C333 output.n141 gnd 1.67353f
C334 outputibias.t10 gnd 0.11477f
C335 outputibias.t9 gnd 0.115567f
C336 outputibias.n0 gnd 0.130108f
C337 outputibias.n1 gnd 0.001372f
C338 outputibias.n2 gnd 9.76e-19
C339 outputibias.n3 gnd 5.24e-19
C340 outputibias.n4 gnd 0.001239f
C341 outputibias.n5 gnd 5.55e-19
C342 outputibias.n6 gnd 9.76e-19
C343 outputibias.n7 gnd 5.24e-19
C344 outputibias.n8 gnd 0.001239f
C345 outputibias.n9 gnd 5.55e-19
C346 outputibias.n10 gnd 0.004176f
C347 outputibias.t5 gnd 0.00202f
C348 outputibias.n11 gnd 9.3e-19
C349 outputibias.n12 gnd 7.32e-19
C350 outputibias.n13 gnd 5.24e-19
C351 outputibias.n14 gnd 0.02322f
C352 outputibias.n15 gnd 9.76e-19
C353 outputibias.n16 gnd 5.24e-19
C354 outputibias.n17 gnd 5.55e-19
C355 outputibias.n18 gnd 0.001239f
C356 outputibias.n19 gnd 0.001239f
C357 outputibias.n20 gnd 5.55e-19
C358 outputibias.n21 gnd 5.24e-19
C359 outputibias.n22 gnd 9.76e-19
C360 outputibias.n23 gnd 9.76e-19
C361 outputibias.n24 gnd 5.24e-19
C362 outputibias.n25 gnd 5.55e-19
C363 outputibias.n26 gnd 0.001239f
C364 outputibias.n27 gnd 0.002683f
C365 outputibias.n28 gnd 5.55e-19
C366 outputibias.n29 gnd 5.24e-19
C367 outputibias.n30 gnd 0.002256f
C368 outputibias.n31 gnd 0.005781f
C369 outputibias.n32 gnd 0.001372f
C370 outputibias.n33 gnd 9.76e-19
C371 outputibias.n34 gnd 5.24e-19
C372 outputibias.n35 gnd 0.001239f
C373 outputibias.n36 gnd 5.55e-19
C374 outputibias.n37 gnd 9.76e-19
C375 outputibias.n38 gnd 5.24e-19
C376 outputibias.n39 gnd 0.001239f
C377 outputibias.n40 gnd 5.55e-19
C378 outputibias.n41 gnd 0.004176f
C379 outputibias.t7 gnd 0.00202f
C380 outputibias.n42 gnd 9.3e-19
C381 outputibias.n43 gnd 7.32e-19
C382 outputibias.n44 gnd 5.24e-19
C383 outputibias.n45 gnd 0.02322f
C384 outputibias.n46 gnd 9.76e-19
C385 outputibias.n47 gnd 5.24e-19
C386 outputibias.n48 gnd 5.55e-19
C387 outputibias.n49 gnd 0.001239f
C388 outputibias.n50 gnd 0.001239f
C389 outputibias.n51 gnd 5.55e-19
C390 outputibias.n52 gnd 5.24e-19
C391 outputibias.n53 gnd 9.76e-19
C392 outputibias.n54 gnd 9.76e-19
C393 outputibias.n55 gnd 5.24e-19
C394 outputibias.n56 gnd 5.55e-19
C395 outputibias.n57 gnd 0.001239f
C396 outputibias.n58 gnd 0.002683f
C397 outputibias.n59 gnd 5.55e-19
C398 outputibias.n60 gnd 5.24e-19
C399 outputibias.n61 gnd 0.002256f
C400 outputibias.n62 gnd 0.005197f
C401 outputibias.n63 gnd 0.121892f
C402 outputibias.n64 gnd 0.001372f
C403 outputibias.n65 gnd 9.76e-19
C404 outputibias.n66 gnd 5.24e-19
C405 outputibias.n67 gnd 0.001239f
C406 outputibias.n68 gnd 5.55e-19
C407 outputibias.n69 gnd 9.76e-19
C408 outputibias.n70 gnd 5.24e-19
C409 outputibias.n71 gnd 0.001239f
C410 outputibias.n72 gnd 5.55e-19
C411 outputibias.n73 gnd 0.004176f
C412 outputibias.t1 gnd 0.00202f
C413 outputibias.n74 gnd 9.3e-19
C414 outputibias.n75 gnd 7.32e-19
C415 outputibias.n76 gnd 5.24e-19
C416 outputibias.n77 gnd 0.02322f
C417 outputibias.n78 gnd 9.76e-19
C418 outputibias.n79 gnd 5.24e-19
C419 outputibias.n80 gnd 5.55e-19
C420 outputibias.n81 gnd 0.001239f
C421 outputibias.n82 gnd 0.001239f
C422 outputibias.n83 gnd 5.55e-19
C423 outputibias.n84 gnd 5.24e-19
C424 outputibias.n85 gnd 9.76e-19
C425 outputibias.n86 gnd 9.76e-19
C426 outputibias.n87 gnd 5.24e-19
C427 outputibias.n88 gnd 5.55e-19
C428 outputibias.n89 gnd 0.001239f
C429 outputibias.n90 gnd 0.002683f
C430 outputibias.n91 gnd 5.55e-19
C431 outputibias.n92 gnd 5.24e-19
C432 outputibias.n93 gnd 0.002256f
C433 outputibias.n94 gnd 0.005197f
C434 outputibias.n95 gnd 0.064513f
C435 outputibias.n96 gnd 0.001372f
C436 outputibias.n97 gnd 9.76e-19
C437 outputibias.n98 gnd 5.24e-19
C438 outputibias.n99 gnd 0.001239f
C439 outputibias.n100 gnd 5.55e-19
C440 outputibias.n101 gnd 9.76e-19
C441 outputibias.n102 gnd 5.24e-19
C442 outputibias.n103 gnd 0.001239f
C443 outputibias.n104 gnd 5.55e-19
C444 outputibias.n105 gnd 0.004176f
C445 outputibias.t3 gnd 0.00202f
C446 outputibias.n106 gnd 9.3e-19
C447 outputibias.n107 gnd 7.32e-19
C448 outputibias.n108 gnd 5.24e-19
C449 outputibias.n109 gnd 0.02322f
C450 outputibias.n110 gnd 9.76e-19
C451 outputibias.n111 gnd 5.24e-19
C452 outputibias.n112 gnd 5.55e-19
C453 outputibias.n113 gnd 0.001239f
C454 outputibias.n114 gnd 0.001239f
C455 outputibias.n115 gnd 5.55e-19
C456 outputibias.n116 gnd 5.24e-19
C457 outputibias.n117 gnd 9.76e-19
C458 outputibias.n118 gnd 9.76e-19
C459 outputibias.n119 gnd 5.24e-19
C460 outputibias.n120 gnd 5.55e-19
C461 outputibias.n121 gnd 0.001239f
C462 outputibias.n122 gnd 0.002683f
C463 outputibias.n123 gnd 5.55e-19
C464 outputibias.n124 gnd 5.24e-19
C465 outputibias.n125 gnd 0.002256f
C466 outputibias.n126 gnd 0.005197f
C467 outputibias.n127 gnd 0.084814f
C468 outputibias.t2 gnd 0.108319f
C469 outputibias.t0 gnd 0.108319f
C470 outputibias.t6 gnd 0.108319f
C471 outputibias.t4 gnd 0.109238f
C472 outputibias.n128 gnd 0.134674f
C473 outputibias.n129 gnd 0.07244f
C474 outputibias.n130 gnd 0.079818f
C475 outputibias.n131 gnd 0.164901f
C476 outputibias.t11 gnd 0.11477f
C477 outputibias.n132 gnd 0.067481f
C478 outputibias.t8 gnd 0.11477f
C479 outputibias.n133 gnd 0.065115f
C480 outputibias.n134 gnd 0.029159f
C481 a_n1808_13878.t4 gnd 0.185683f
C482 a_n1808_13878.t0 gnd 0.185683f
C483 a_n1808_13878.t2 gnd 0.185683f
C484 a_n1808_13878.n0 gnd 1.46364f
C485 a_n1808_13878.t6 gnd 0.185683f
C486 a_n1808_13878.t1 gnd 0.185683f
C487 a_n1808_13878.n1 gnd 1.46209f
C488 a_n1808_13878.n2 gnd 2.04299f
C489 a_n1808_13878.t5 gnd 0.185683f
C490 a_n1808_13878.t9 gnd 0.185683f
C491 a_n1808_13878.n3 gnd 1.46451f
C492 a_n1808_13878.t10 gnd 0.185683f
C493 a_n1808_13878.t3 gnd 0.185683f
C494 a_n1808_13878.n4 gnd 1.46209f
C495 a_n1808_13878.n5 gnd 1.31424f
C496 a_n1808_13878.t7 gnd 0.185683f
C497 a_n1808_13878.t8 gnd 0.185683f
C498 a_n1808_13878.n6 gnd 1.46209f
C499 a_n1808_13878.n7 gnd 1.80499f
C500 a_n1808_13878.t13 gnd 1.73864f
C501 a_n1808_13878.t16 gnd 0.185683f
C502 a_n1808_13878.t17 gnd 0.185683f
C503 a_n1808_13878.n8 gnd 1.30795f
C504 a_n1808_13878.n9 gnd 1.46144f
C505 a_n1808_13878.t12 gnd 1.73518f
C506 a_n1808_13878.n10 gnd 0.735417f
C507 a_n1808_13878.t15 gnd 1.73518f
C508 a_n1808_13878.n11 gnd 0.735417f
C509 a_n1808_13878.t18 gnd 0.185683f
C510 a_n1808_13878.t19 gnd 0.185683f
C511 a_n1808_13878.n12 gnd 1.30795f
C512 a_n1808_13878.n13 gnd 0.742539f
C513 a_n1808_13878.t14 gnd 1.73518f
C514 a_n1808_13878.n14 gnd 1.73174f
C515 a_n1808_13878.n15 gnd 2.52099f
C516 a_n1808_13878.n16 gnd 3.70273f
C517 a_n1808_13878.n17 gnd 1.46209f
C518 a_n1808_13878.t11 gnd 0.185683f
C519 a_n1986_8322.t20 gnd 38.672398f
C520 a_n1986_8322.t22 gnd 27.512402f
C521 a_n1986_8322.t23 gnd 19.268198f
C522 a_n1986_8322.t21 gnd 38.672398f
C523 a_n1986_8322.t2 gnd 0.093533f
C524 a_n1986_8322.t1 gnd 0.875792f
C525 a_n1986_8322.t9 gnd 0.093533f
C526 a_n1986_8322.t4 gnd 0.093533f
C527 a_n1986_8322.n0 gnd 0.658844f
C528 a_n1986_8322.n1 gnd 0.736161f
C529 a_n1986_8322.t7 gnd 0.093533f
C530 a_n1986_8322.t6 gnd 0.093533f
C531 a_n1986_8322.n2 gnd 0.658844f
C532 a_n1986_8322.n3 gnd 0.374034f
C533 a_n1986_8322.t0 gnd 0.874048f
C534 a_n1986_8322.n4 gnd 1.39896f
C535 a_n1986_8322.t14 gnd 0.875792f
C536 a_n1986_8322.t18 gnd 0.093533f
C537 a_n1986_8322.t17 gnd 0.093533f
C538 a_n1986_8322.n5 gnd 0.658844f
C539 a_n1986_8322.n6 gnd 0.736161f
C540 a_n1986_8322.t12 gnd 0.874048f
C541 a_n1986_8322.n7 gnd 0.370446f
C542 a_n1986_8322.t15 gnd 0.874048f
C543 a_n1986_8322.n8 gnd 0.370446f
C544 a_n1986_8322.t13 gnd 0.093533f
C545 a_n1986_8322.t19 gnd 0.093533f
C546 a_n1986_8322.n9 gnd 0.658844f
C547 a_n1986_8322.n10 gnd 0.374034f
C548 a_n1986_8322.t16 gnd 0.874048f
C549 a_n1986_8322.n11 gnd 0.872317f
C550 a_n1986_8322.n12 gnd 1.59071f
C551 a_n1986_8322.n13 gnd 3.20172f
C552 a_n1986_8322.t3 gnd 0.874048f
C553 a_n1986_8322.n14 gnd 0.76652f
C554 a_n1986_8322.t10 gnd 0.875789f
C555 a_n1986_8322.t8 gnd 0.093533f
C556 a_n1986_8322.t5 gnd 0.093533f
C557 a_n1986_8322.n15 gnd 0.658844f
C558 a_n1986_8322.n16 gnd 0.736163f
C559 a_n1986_8322.n17 gnd 0.374032f
C560 a_n1986_8322.n18 gnd 0.658845f
C561 a_n1986_8322.t11 gnd 0.093533f
C562 a_n1996_n452.n0 gnd 0.822727f
C563 a_n1996_n452.n1 gnd 3.34433f
C564 a_n1996_n452.n2 gnd 3.17111f
C565 a_n1996_n452.n3 gnd 3.91594f
C566 a_n1996_n452.n4 gnd 0.527811f
C567 a_n1996_n452.n5 gnd 0.205584f
C568 a_n1996_n452.n6 gnd 0.151417f
C569 a_n1996_n452.n7 gnd 0.237979f
C570 a_n1996_n452.n8 gnd 0.183812f
C571 a_n1996_n452.n9 gnd 0.205584f
C572 a_n1996_n452.n10 gnd 0.151417f
C573 a_n1996_n452.n11 gnd 0.581979f
C574 a_n1996_n452.n12 gnd 0.433746f
C575 a_n1996_n452.n13 gnd 0.21667f
C576 a_n1996_n452.n14 gnd 0.494132f
C577 a_n1996_n452.n15 gnd 0.283464f
C578 a_n1996_n452.n16 gnd 0.439964f
C579 a_n1996_n452.n17 gnd 0.21667f
C580 a_n1996_n452.n18 gnd 0.734001f
C581 a_n1996_n452.n19 gnd 0.283464f
C582 a_n1996_n452.n20 gnd 0.641354f
C583 a_n1996_n452.n21 gnd 0.283464f
C584 a_n1996_n452.n22 gnd 0.494132f
C585 a_n1996_n452.n23 gnd 0.666675f
C586 a_n1996_n452.n24 gnd 0.21667f
C587 a_n1996_n452.n25 gnd 0.283464f
C588 a_n1996_n452.n26 gnd 1.78382f
C589 a_n1996_n452.n27 gnd 1.18284f
C590 a_n1996_n452.n28 gnd 1.92214f
C591 a_n1996_n452.n29 gnd 3.22512f
C592 a_n1996_n452.n30 gnd 0.008389f
C593 a_n1996_n452.n32 gnd 1.34296f
C594 a_n1996_n452.n33 gnd 0.286629f
C595 a_n1996_n452.n34 gnd 0.108335f
C596 a_n1996_n452.n35 gnd 0.008389f
C597 a_n1996_n452.n37 gnd 0.008389f
C598 a_n1996_n452.n39 gnd 0.286629f
C599 a_n1996_n452.n40 gnd 0.008389f
C600 a_n1996_n452.n42 gnd 0.286629f
C601 a_n1996_n452.n43 gnd 0.008389f
C602 a_n1996_n452.n44 gnd 0.286221f
C603 a_n1996_n452.n45 gnd 0.008389f
C604 a_n1996_n452.n46 gnd 0.286221f
C605 a_n1996_n452.n47 gnd 0.008389f
C606 a_n1996_n452.n48 gnd 0.286221f
C607 a_n1996_n452.n49 gnd 0.008389f
C608 a_n1996_n452.n50 gnd 0.286221f
C609 a_n1996_n452.n51 gnd 0.286629f
C610 a_n1996_n452.t23 gnd 0.150285f
C611 a_n1996_n452.t31 gnd 1.40719f
C612 a_n1996_n452.t29 gnd 0.150285f
C613 a_n1996_n452.t21 gnd 0.150285f
C614 a_n1996_n452.n52 gnd 1.05861f
C615 a_n1996_n452.t14 gnd 0.699053f
C616 a_n1996_n452.n53 gnd 0.307348f
C617 a_n1996_n452.t22 gnd 0.699053f
C618 a_n1996_n452.t28 gnd 0.699053f
C619 a_n1996_n452.t52 gnd 0.699053f
C620 a_n1996_n452.n54 gnd 0.307348f
C621 a_n1996_n452.t61 gnd 0.699053f
C622 a_n1996_n452.t67 gnd 0.699053f
C623 a_n1996_n452.t18 gnd 0.713776f
C624 a_n1996_n452.t16 gnd 0.699053f
C625 a_n1996_n452.t36 gnd 0.699053f
C626 a_n1996_n452.t32 gnd 0.699053f
C627 a_n1996_n452.n55 gnd 0.307348f
C628 a_n1996_n452.t34 gnd 0.699053f
C629 a_n1996_n452.t26 gnd 0.710611f
C630 a_n1996_n452.t5 gnd 0.116888f
C631 a_n1996_n452.t40 gnd 0.116888f
C632 a_n1996_n452.n56 gnd 1.03516f
C633 a_n1996_n452.t3 gnd 0.116888f
C634 a_n1996_n452.t4 gnd 0.116888f
C635 a_n1996_n452.n57 gnd 1.03287f
C636 a_n1996_n452.t39 gnd 0.116888f
C637 a_n1996_n452.t6 gnd 0.116888f
C638 a_n1996_n452.n58 gnd 1.03287f
C639 a_n1996_n452.t13 gnd 0.116888f
C640 a_n1996_n452.t38 gnd 0.116888f
C641 a_n1996_n452.n59 gnd 1.03516f
C642 a_n1996_n452.t7 gnd 0.116888f
C643 a_n1996_n452.t42 gnd 0.116888f
C644 a_n1996_n452.n60 gnd 1.03287f
C645 a_n1996_n452.t2 gnd 0.116888f
C646 a_n1996_n452.t9 gnd 0.116888f
C647 a_n1996_n452.n61 gnd 1.03287f
C648 a_n1996_n452.t43 gnd 0.116888f
C649 a_n1996_n452.t11 gnd 0.116888f
C650 a_n1996_n452.n62 gnd 1.03287f
C651 a_n1996_n452.t0 gnd 0.116888f
C652 a_n1996_n452.t10 gnd 0.116888f
C653 a_n1996_n452.n63 gnd 1.03287f
C654 a_n1996_n452.t8 gnd 0.116888f
C655 a_n1996_n452.t1 gnd 0.116888f
C656 a_n1996_n452.n64 gnd 1.03516f
C657 a_n1996_n452.t12 gnd 0.116888f
C658 a_n1996_n452.t41 gnd 0.116888f
C659 a_n1996_n452.n65 gnd 1.03287f
C660 a_n1996_n452.t71 gnd 0.713776f
C661 a_n1996_n452.t54 gnd 0.699053f
C662 a_n1996_n452.t58 gnd 0.699053f
C663 a_n1996_n452.t48 gnd 0.699053f
C664 a_n1996_n452.n66 gnd 0.307348f
C665 a_n1996_n452.t63 gnd 0.699053f
C666 a_n1996_n452.t69 gnd 0.710611f
C667 a_n1996_n452.n67 gnd 0.309974f
C668 a_n1996_n452.n68 gnd 0.303445f
C669 a_n1996_n452.n69 gnd 0.309974f
C670 a_n1996_n452.n70 gnd 0.309974f
C671 a_n1996_n452.n71 gnd 0.303445f
C672 a_n1996_n452.n72 gnd 0.309974f
C673 a_n1996_n452.t27 gnd 1.40719f
C674 a_n1996_n452.t33 gnd 0.150285f
C675 a_n1996_n452.t35 gnd 0.150285f
C676 a_n1996_n452.n73 gnd 1.05861f
C677 a_n1996_n452.t17 gnd 0.150285f
C678 a_n1996_n452.t37 gnd 0.150285f
C679 a_n1996_n452.n74 gnd 1.05861f
C680 a_n1996_n452.t19 gnd 1.40439f
C681 a_n1996_n452.n75 gnd 1.14844f
C682 a_n1996_n452.n76 gnd 0.789587f
C683 a_n1996_n452.t53 gnd 0.699053f
C684 a_n1996_n452.t62 gnd 0.699053f
C685 a_n1996_n452.t44 gnd 0.699053f
C686 a_n1996_n452.n77 gnd 0.307348f
C687 a_n1996_n452.t64 gnd 0.699053f
C688 a_n1996_n452.t49 gnd 0.699053f
C689 a_n1996_n452.t50 gnd 0.699053f
C690 a_n1996_n452.n78 gnd 0.307348f
C691 a_n1996_n452.t68 gnd 0.699053f
C692 a_n1996_n452.t57 gnd 0.699053f
C693 a_n1996_n452.t56 gnd 0.699053f
C694 a_n1996_n452.n79 gnd 0.307348f
C695 a_n1996_n452.t60 gnd 0.699053f
C696 a_n1996_n452.t51 gnd 0.699053f
C697 a_n1996_n452.t45 gnd 0.699053f
C698 a_n1996_n452.n80 gnd 0.307348f
C699 a_n1996_n452.t65 gnd 0.710766f
C700 a_n1996_n452.n81 gnd 0.303445f
C701 a_n1996_n452.n82 gnd 0.297934f
C702 a_n1996_n452.t70 gnd 0.710766f
C703 a_n1996_n452.n83 gnd 0.303445f
C704 a_n1996_n452.n84 gnd 0.297934f
C705 a_n1996_n452.t59 gnd 0.710766f
C706 a_n1996_n452.n85 gnd 0.303445f
C707 a_n1996_n452.n86 gnd 0.297934f
C708 a_n1996_n452.t55 gnd 0.710766f
C709 a_n1996_n452.n87 gnd 0.303445f
C710 a_n1996_n452.n88 gnd 0.297934f
C711 a_n1996_n452.n89 gnd 1.00969f
C712 a_n1996_n452.t66 gnd 0.713776f
C713 a_n1996_n452.n90 gnd 0.309974f
C714 a_n1996_n452.t46 gnd 0.699053f
C715 a_n1996_n452.n91 gnd 0.303445f
C716 a_n1996_n452.n92 gnd 0.309974f
C717 a_n1996_n452.t47 gnd 0.710611f
C718 a_n1996_n452.t30 gnd 0.713776f
C719 a_n1996_n452.n93 gnd 0.309974f
C720 a_n1996_n452.t20 gnd 0.699053f
C721 a_n1996_n452.n94 gnd 0.303445f
C722 a_n1996_n452.n95 gnd 0.309974f
C723 a_n1996_n452.t24 gnd 0.710611f
C724 a_n1996_n452.n96 gnd 1.13585f
C725 a_n1996_n452.t25 gnd 1.40439f
C726 a_n1996_n452.n97 gnd 1.05861f
C727 a_n1996_n452.t15 gnd 0.150285f
C728 vdd.t114 gnd 0.032933f
C729 vdd.t16 gnd 0.032933f
C730 vdd.n0 gnd 0.259746f
C731 vdd.t107 gnd 0.032933f
C732 vdd.t117 gnd 0.032933f
C733 vdd.n1 gnd 0.259317f
C734 vdd.n2 gnd 0.23914f
C735 vdd.t8 gnd 0.032933f
C736 vdd.t3 gnd 0.032933f
C737 vdd.n3 gnd 0.259317f
C738 vdd.n4 gnd 0.120942f
C739 vdd.t123 gnd 0.032933f
C740 vdd.t112 gnd 0.032933f
C741 vdd.n5 gnd 0.259317f
C742 vdd.n6 gnd 0.113482f
C743 vdd.t110 gnd 0.032933f
C744 vdd.t18 gnd 0.032933f
C745 vdd.n7 gnd 0.259746f
C746 vdd.t1 gnd 0.032933f
C747 vdd.t5 gnd 0.032933f
C748 vdd.n8 gnd 0.259317f
C749 vdd.n9 gnd 0.23914f
C750 vdd.t22 gnd 0.032933f
C751 vdd.t11 gnd 0.032933f
C752 vdd.n10 gnd 0.259317f
C753 vdd.n11 gnd 0.120942f
C754 vdd.t119 gnd 0.032933f
C755 vdd.t14 gnd 0.032933f
C756 vdd.n12 gnd 0.259317f
C757 vdd.n13 gnd 0.113482f
C758 vdd.n14 gnd 0.080229f
C759 vdd.t99 gnd 0.018296f
C760 vdd.t96 gnd 0.018296f
C761 vdd.n15 gnd 0.168407f
C762 vdd.t102 gnd 0.018296f
C763 vdd.t91 gnd 0.018296f
C764 vdd.n16 gnd 0.167914f
C765 vdd.n17 gnd 0.292223f
C766 vdd.t90 gnd 0.018296f
C767 vdd.t104 gnd 0.018296f
C768 vdd.n18 gnd 0.167914f
C769 vdd.n19 gnd 0.120896f
C770 vdd.t101 gnd 0.018296f
C771 vdd.t97 gnd 0.018296f
C772 vdd.n20 gnd 0.168407f
C773 vdd.t92 gnd 0.018296f
C774 vdd.t95 gnd 0.018296f
C775 vdd.n21 gnd 0.167914f
C776 vdd.n22 gnd 0.292223f
C777 vdd.t93 gnd 0.018296f
C778 vdd.t89 gnd 0.018296f
C779 vdd.n23 gnd 0.167914f
C780 vdd.n24 gnd 0.120896f
C781 vdd.t100 gnd 0.018296f
C782 vdd.t94 gnd 0.018296f
C783 vdd.n25 gnd 0.167914f
C784 vdd.t98 gnd 0.018296f
C785 vdd.t103 gnd 0.018296f
C786 vdd.n26 gnd 0.167914f
C787 vdd.n27 gnd 18.208302f
C788 vdd.n28 gnd 6.72294f
C789 vdd.n29 gnd 0.00499f
C790 vdd.n30 gnd 0.004631f
C791 vdd.n31 gnd 0.002561f
C792 vdd.n32 gnd 0.005881f
C793 vdd.n33 gnd 0.002488f
C794 vdd.n34 gnd 0.002635f
C795 vdd.n35 gnd 0.004631f
C796 vdd.n36 gnd 0.002488f
C797 vdd.n37 gnd 0.005881f
C798 vdd.n38 gnd 0.002635f
C799 vdd.n39 gnd 0.004631f
C800 vdd.n40 gnd 0.002488f
C801 vdd.n41 gnd 0.004411f
C802 vdd.n42 gnd 0.004424f
C803 vdd.t26 gnd 0.012636f
C804 vdd.n43 gnd 0.028114f
C805 vdd.n44 gnd 0.146311f
C806 vdd.n45 gnd 0.002488f
C807 vdd.n46 gnd 0.002635f
C808 vdd.n47 gnd 0.005881f
C809 vdd.n48 gnd 0.005881f
C810 vdd.n49 gnd 0.002635f
C811 vdd.n50 gnd 0.002488f
C812 vdd.n51 gnd 0.004631f
C813 vdd.n52 gnd 0.004631f
C814 vdd.n53 gnd 0.002488f
C815 vdd.n54 gnd 0.002635f
C816 vdd.n55 gnd 0.005881f
C817 vdd.n56 gnd 0.005881f
C818 vdd.n57 gnd 0.002635f
C819 vdd.n58 gnd 0.002488f
C820 vdd.n59 gnd 0.004631f
C821 vdd.n60 gnd 0.004631f
C822 vdd.n61 gnd 0.002488f
C823 vdd.n62 gnd 0.002635f
C824 vdd.n63 gnd 0.005881f
C825 vdd.n64 gnd 0.005881f
C826 vdd.n65 gnd 0.013905f
C827 vdd.n66 gnd 0.002561f
C828 vdd.n67 gnd 0.002488f
C829 vdd.n68 gnd 0.011968f
C830 vdd.n69 gnd 0.008356f
C831 vdd.t78 gnd 0.029274f
C832 vdd.t52 gnd 0.029274f
C833 vdd.n70 gnd 0.201188f
C834 vdd.n71 gnd 0.158204f
C835 vdd.t85 gnd 0.029274f
C836 vdd.t41 gnd 0.029274f
C837 vdd.n72 gnd 0.201188f
C838 vdd.n73 gnd 0.127669f
C839 vdd.t71 gnd 0.029274f
C840 vdd.t46 gnd 0.029274f
C841 vdd.n74 gnd 0.201188f
C842 vdd.n75 gnd 0.127669f
C843 vdd.n76 gnd 0.00499f
C844 vdd.n77 gnd 0.004631f
C845 vdd.n78 gnd 0.002561f
C846 vdd.n79 gnd 0.005881f
C847 vdd.n80 gnd 0.002488f
C848 vdd.n81 gnd 0.002635f
C849 vdd.n82 gnd 0.004631f
C850 vdd.n83 gnd 0.002488f
C851 vdd.n84 gnd 0.005881f
C852 vdd.n85 gnd 0.002635f
C853 vdd.n86 gnd 0.004631f
C854 vdd.n87 gnd 0.002488f
C855 vdd.n88 gnd 0.004411f
C856 vdd.n89 gnd 0.004424f
C857 vdd.t84 gnd 0.012636f
C858 vdd.n90 gnd 0.028114f
C859 vdd.n91 gnd 0.146311f
C860 vdd.n92 gnd 0.002488f
C861 vdd.n93 gnd 0.002635f
C862 vdd.n94 gnd 0.005881f
C863 vdd.n95 gnd 0.005881f
C864 vdd.n96 gnd 0.002635f
C865 vdd.n97 gnd 0.002488f
C866 vdd.n98 gnd 0.004631f
C867 vdd.n99 gnd 0.004631f
C868 vdd.n100 gnd 0.002488f
C869 vdd.n101 gnd 0.002635f
C870 vdd.n102 gnd 0.005881f
C871 vdd.n103 gnd 0.005881f
C872 vdd.n104 gnd 0.002635f
C873 vdd.n105 gnd 0.002488f
C874 vdd.n106 gnd 0.004631f
C875 vdd.n107 gnd 0.004631f
C876 vdd.n108 gnd 0.002488f
C877 vdd.n109 gnd 0.002635f
C878 vdd.n110 gnd 0.005881f
C879 vdd.n111 gnd 0.005881f
C880 vdd.n112 gnd 0.013905f
C881 vdd.n113 gnd 0.002561f
C882 vdd.n114 gnd 0.002488f
C883 vdd.n115 gnd 0.011968f
C884 vdd.n116 gnd 0.008094f
C885 vdd.n117 gnd 0.094987f
C886 vdd.n118 gnd 0.00499f
C887 vdd.n119 gnd 0.004631f
C888 vdd.n120 gnd 0.002561f
C889 vdd.n121 gnd 0.005881f
C890 vdd.n122 gnd 0.002488f
C891 vdd.n123 gnd 0.002635f
C892 vdd.n124 gnd 0.004631f
C893 vdd.n125 gnd 0.002488f
C894 vdd.n126 gnd 0.005881f
C895 vdd.n127 gnd 0.002635f
C896 vdd.n128 gnd 0.004631f
C897 vdd.n129 gnd 0.002488f
C898 vdd.n130 gnd 0.004411f
C899 vdd.n131 gnd 0.004424f
C900 vdd.t53 gnd 0.012636f
C901 vdd.n132 gnd 0.028114f
C902 vdd.n133 gnd 0.146311f
C903 vdd.n134 gnd 0.002488f
C904 vdd.n135 gnd 0.002635f
C905 vdd.n136 gnd 0.005881f
C906 vdd.n137 gnd 0.005881f
C907 vdd.n138 gnd 0.002635f
C908 vdd.n139 gnd 0.002488f
C909 vdd.n140 gnd 0.004631f
C910 vdd.n141 gnd 0.004631f
C911 vdd.n142 gnd 0.002488f
C912 vdd.n143 gnd 0.002635f
C913 vdd.n144 gnd 0.005881f
C914 vdd.n145 gnd 0.005881f
C915 vdd.n146 gnd 0.002635f
C916 vdd.n147 gnd 0.002488f
C917 vdd.n148 gnd 0.004631f
C918 vdd.n149 gnd 0.004631f
C919 vdd.n150 gnd 0.002488f
C920 vdd.n151 gnd 0.002635f
C921 vdd.n152 gnd 0.005881f
C922 vdd.n153 gnd 0.005881f
C923 vdd.n154 gnd 0.013905f
C924 vdd.n155 gnd 0.002561f
C925 vdd.n156 gnd 0.002488f
C926 vdd.n157 gnd 0.011968f
C927 vdd.n158 gnd 0.008356f
C928 vdd.t55 gnd 0.029274f
C929 vdd.t66 gnd 0.029274f
C930 vdd.n159 gnd 0.201188f
C931 vdd.n160 gnd 0.158204f
C932 vdd.t30 gnd 0.029274f
C933 vdd.t49 gnd 0.029274f
C934 vdd.n161 gnd 0.201188f
C935 vdd.n162 gnd 0.127669f
C936 vdd.t65 gnd 0.029274f
C937 vdd.t86 gnd 0.029274f
C938 vdd.n163 gnd 0.201188f
C939 vdd.n164 gnd 0.127669f
C940 vdd.n165 gnd 0.00499f
C941 vdd.n166 gnd 0.004631f
C942 vdd.n167 gnd 0.002561f
C943 vdd.n168 gnd 0.005881f
C944 vdd.n169 gnd 0.002488f
C945 vdd.n170 gnd 0.002635f
C946 vdd.n171 gnd 0.004631f
C947 vdd.n172 gnd 0.002488f
C948 vdd.n173 gnd 0.005881f
C949 vdd.n174 gnd 0.002635f
C950 vdd.n175 gnd 0.004631f
C951 vdd.n176 gnd 0.002488f
C952 vdd.n177 gnd 0.004411f
C953 vdd.n178 gnd 0.004424f
C954 vdd.t43 gnd 0.012636f
C955 vdd.n179 gnd 0.028114f
C956 vdd.n180 gnd 0.146311f
C957 vdd.n181 gnd 0.002488f
C958 vdd.n182 gnd 0.002635f
C959 vdd.n183 gnd 0.005881f
C960 vdd.n184 gnd 0.005881f
C961 vdd.n185 gnd 0.002635f
C962 vdd.n186 gnd 0.002488f
C963 vdd.n187 gnd 0.004631f
C964 vdd.n188 gnd 0.004631f
C965 vdd.n189 gnd 0.002488f
C966 vdd.n190 gnd 0.002635f
C967 vdd.n191 gnd 0.005881f
C968 vdd.n192 gnd 0.005881f
C969 vdd.n193 gnd 0.002635f
C970 vdd.n194 gnd 0.002488f
C971 vdd.n195 gnd 0.004631f
C972 vdd.n196 gnd 0.004631f
C973 vdd.n197 gnd 0.002488f
C974 vdd.n198 gnd 0.002635f
C975 vdd.n199 gnd 0.005881f
C976 vdd.n200 gnd 0.005881f
C977 vdd.n201 gnd 0.013905f
C978 vdd.n202 gnd 0.002561f
C979 vdd.n203 gnd 0.002488f
C980 vdd.n204 gnd 0.011968f
C981 vdd.n205 gnd 0.008094f
C982 vdd.n206 gnd 0.056507f
C983 vdd.n207 gnd 0.203611f
C984 vdd.n208 gnd 0.00499f
C985 vdd.n209 gnd 0.004631f
C986 vdd.n210 gnd 0.002561f
C987 vdd.n211 gnd 0.005881f
C988 vdd.n212 gnd 0.002488f
C989 vdd.n213 gnd 0.002635f
C990 vdd.n214 gnd 0.004631f
C991 vdd.n215 gnd 0.002488f
C992 vdd.n216 gnd 0.005881f
C993 vdd.n217 gnd 0.002635f
C994 vdd.n218 gnd 0.004631f
C995 vdd.n219 gnd 0.002488f
C996 vdd.n220 gnd 0.004411f
C997 vdd.n221 gnd 0.004424f
C998 vdd.t58 gnd 0.012636f
C999 vdd.n222 gnd 0.028114f
C1000 vdd.n223 gnd 0.146311f
C1001 vdd.n224 gnd 0.002488f
C1002 vdd.n225 gnd 0.002635f
C1003 vdd.n226 gnd 0.005881f
C1004 vdd.n227 gnd 0.005881f
C1005 vdd.n228 gnd 0.002635f
C1006 vdd.n229 gnd 0.002488f
C1007 vdd.n230 gnd 0.004631f
C1008 vdd.n231 gnd 0.004631f
C1009 vdd.n232 gnd 0.002488f
C1010 vdd.n233 gnd 0.002635f
C1011 vdd.n234 gnd 0.005881f
C1012 vdd.n235 gnd 0.005881f
C1013 vdd.n236 gnd 0.002635f
C1014 vdd.n237 gnd 0.002488f
C1015 vdd.n238 gnd 0.004631f
C1016 vdd.n239 gnd 0.004631f
C1017 vdd.n240 gnd 0.002488f
C1018 vdd.n241 gnd 0.002635f
C1019 vdd.n242 gnd 0.005881f
C1020 vdd.n243 gnd 0.005881f
C1021 vdd.n244 gnd 0.013905f
C1022 vdd.n245 gnd 0.002561f
C1023 vdd.n246 gnd 0.002488f
C1024 vdd.n247 gnd 0.011968f
C1025 vdd.n248 gnd 0.008356f
C1026 vdd.t59 gnd 0.029274f
C1027 vdd.t75 gnd 0.029274f
C1028 vdd.n249 gnd 0.201188f
C1029 vdd.n250 gnd 0.158204f
C1030 vdd.t36 gnd 0.029274f
C1031 vdd.t57 gnd 0.029274f
C1032 vdd.n251 gnd 0.201188f
C1033 vdd.n252 gnd 0.127669f
C1034 vdd.t70 gnd 0.029274f
C1035 vdd.t34 gnd 0.029274f
C1036 vdd.n253 gnd 0.201188f
C1037 vdd.n254 gnd 0.127669f
C1038 vdd.n255 gnd 0.00499f
C1039 vdd.n256 gnd 0.004631f
C1040 vdd.n257 gnd 0.002561f
C1041 vdd.n258 gnd 0.005881f
C1042 vdd.n259 gnd 0.002488f
C1043 vdd.n260 gnd 0.002635f
C1044 vdd.n261 gnd 0.004631f
C1045 vdd.n262 gnd 0.002488f
C1046 vdd.n263 gnd 0.005881f
C1047 vdd.n264 gnd 0.002635f
C1048 vdd.n265 gnd 0.004631f
C1049 vdd.n266 gnd 0.002488f
C1050 vdd.n267 gnd 0.004411f
C1051 vdd.n268 gnd 0.004424f
C1052 vdd.t47 gnd 0.012636f
C1053 vdd.n269 gnd 0.028114f
C1054 vdd.n270 gnd 0.146311f
C1055 vdd.n271 gnd 0.002488f
C1056 vdd.n272 gnd 0.002635f
C1057 vdd.n273 gnd 0.005881f
C1058 vdd.n274 gnd 0.005881f
C1059 vdd.n275 gnd 0.002635f
C1060 vdd.n276 gnd 0.002488f
C1061 vdd.n277 gnd 0.004631f
C1062 vdd.n278 gnd 0.004631f
C1063 vdd.n279 gnd 0.002488f
C1064 vdd.n280 gnd 0.002635f
C1065 vdd.n281 gnd 0.005881f
C1066 vdd.n282 gnd 0.005881f
C1067 vdd.n283 gnd 0.002635f
C1068 vdd.n284 gnd 0.002488f
C1069 vdd.n285 gnd 0.004631f
C1070 vdd.n286 gnd 0.004631f
C1071 vdd.n287 gnd 0.002488f
C1072 vdd.n288 gnd 0.002635f
C1073 vdd.n289 gnd 0.005881f
C1074 vdd.n290 gnd 0.005881f
C1075 vdd.n291 gnd 0.013905f
C1076 vdd.n292 gnd 0.002561f
C1077 vdd.n293 gnd 0.002488f
C1078 vdd.n294 gnd 0.011968f
C1079 vdd.n295 gnd 0.008094f
C1080 vdd.n296 gnd 0.056507f
C1081 vdd.n297 gnd 0.220385f
C1082 vdd.n298 gnd 0.006988f
C1083 vdd.n299 gnd 0.009093f
C1084 vdd.n300 gnd 0.007318f
C1085 vdd.n301 gnd 0.007318f
C1086 vdd.n302 gnd 0.009093f
C1087 vdd.n303 gnd 0.009093f
C1088 vdd.n304 gnd 0.664388f
C1089 vdd.n305 gnd 0.009093f
C1090 vdd.n306 gnd 0.009093f
C1091 vdd.n307 gnd 0.009093f
C1092 vdd.n308 gnd 0.720141f
C1093 vdd.n309 gnd 0.009093f
C1094 vdd.n310 gnd 0.009093f
C1095 vdd.n311 gnd 0.009093f
C1096 vdd.n312 gnd 0.009093f
C1097 vdd.n313 gnd 0.007318f
C1098 vdd.n314 gnd 0.009093f
C1099 vdd.t33 gnd 0.464607f
C1100 vdd.n315 gnd 0.009093f
C1101 vdd.n316 gnd 0.009093f
C1102 vdd.n317 gnd 0.009093f
C1103 vdd.n318 gnd 0.929214f
C1104 vdd.n319 gnd 0.009093f
C1105 vdd.n320 gnd 0.009093f
C1106 vdd.n321 gnd 0.009093f
C1107 vdd.n322 gnd 0.009093f
C1108 vdd.n323 gnd 0.009093f
C1109 vdd.n324 gnd 0.007318f
C1110 vdd.n325 gnd 0.009093f
C1111 vdd.n326 gnd 0.009093f
C1112 vdd.n327 gnd 0.009093f
C1113 vdd.n328 gnd 0.022159f
C1114 vdd.n329 gnd 2.22082f
C1115 vdd.n330 gnd 0.022667f
C1116 vdd.n331 gnd 0.009093f
C1117 vdd.n332 gnd 0.009093f
C1118 vdd.n334 gnd 0.009093f
C1119 vdd.n335 gnd 0.009093f
C1120 vdd.n336 gnd 0.007318f
C1121 vdd.n337 gnd 0.007318f
C1122 vdd.n338 gnd 0.009093f
C1123 vdd.n339 gnd 0.009093f
C1124 vdd.n340 gnd 0.009093f
C1125 vdd.n341 gnd 0.009093f
C1126 vdd.n342 gnd 0.009093f
C1127 vdd.n343 gnd 0.009093f
C1128 vdd.n344 gnd 0.007318f
C1129 vdd.n346 gnd 0.009093f
C1130 vdd.n347 gnd 0.009093f
C1131 vdd.n348 gnd 0.009093f
C1132 vdd.n349 gnd 0.009093f
C1133 vdd.n350 gnd 0.009093f
C1134 vdd.n351 gnd 0.007318f
C1135 vdd.n353 gnd 0.009093f
C1136 vdd.n354 gnd 0.009093f
C1137 vdd.n355 gnd 0.009093f
C1138 vdd.n356 gnd 0.009093f
C1139 vdd.n357 gnd 0.009093f
C1140 vdd.n358 gnd 0.007318f
C1141 vdd.n360 gnd 0.009093f
C1142 vdd.n361 gnd 0.009093f
C1143 vdd.n362 gnd 0.009093f
C1144 vdd.n363 gnd 0.009093f
C1145 vdd.n364 gnd 0.006111f
C1146 vdd.t155 gnd 0.111862f
C1147 vdd.t154 gnd 0.11955f
C1148 vdd.t153 gnd 0.14609f
C1149 vdd.n365 gnd 0.187267f
C1150 vdd.n366 gnd 0.15807f
C1151 vdd.n368 gnd 0.009093f
C1152 vdd.n369 gnd 0.009093f
C1153 vdd.n370 gnd 0.007318f
C1154 vdd.n371 gnd 0.009093f
C1155 vdd.n373 gnd 0.009093f
C1156 vdd.n374 gnd 0.009093f
C1157 vdd.n375 gnd 0.009093f
C1158 vdd.n376 gnd 0.009093f
C1159 vdd.n377 gnd 0.007318f
C1160 vdd.n379 gnd 0.009093f
C1161 vdd.n380 gnd 0.009093f
C1162 vdd.n381 gnd 0.009093f
C1163 vdd.n382 gnd 0.009093f
C1164 vdd.n383 gnd 0.009093f
C1165 vdd.n384 gnd 0.007318f
C1166 vdd.n386 gnd 0.009093f
C1167 vdd.n387 gnd 0.009093f
C1168 vdd.n388 gnd 0.009093f
C1169 vdd.n389 gnd 0.009093f
C1170 vdd.n390 gnd 0.009093f
C1171 vdd.n391 gnd 0.007318f
C1172 vdd.n393 gnd 0.009093f
C1173 vdd.n394 gnd 0.009093f
C1174 vdd.n395 gnd 0.009093f
C1175 vdd.n396 gnd 0.009093f
C1176 vdd.n397 gnd 0.009093f
C1177 vdd.n398 gnd 0.007318f
C1178 vdd.n400 gnd 0.009093f
C1179 vdd.n401 gnd 0.009093f
C1180 vdd.n402 gnd 0.009093f
C1181 vdd.n403 gnd 0.009093f
C1182 vdd.n404 gnd 0.007245f
C1183 vdd.t149 gnd 0.111862f
C1184 vdd.t148 gnd 0.11955f
C1185 vdd.t146 gnd 0.14609f
C1186 vdd.n405 gnd 0.187267f
C1187 vdd.n406 gnd 0.15807f
C1188 vdd.n408 gnd 0.009093f
C1189 vdd.n409 gnd 0.009093f
C1190 vdd.n410 gnd 0.007318f
C1191 vdd.n411 gnd 0.009093f
C1192 vdd.n413 gnd 0.009093f
C1193 vdd.n414 gnd 0.009093f
C1194 vdd.n415 gnd 0.009093f
C1195 vdd.n416 gnd 0.009093f
C1196 vdd.n417 gnd 0.007318f
C1197 vdd.n419 gnd 0.009093f
C1198 vdd.n420 gnd 0.009093f
C1199 vdd.n421 gnd 0.009093f
C1200 vdd.n422 gnd 0.009093f
C1201 vdd.n423 gnd 0.009093f
C1202 vdd.n424 gnd 0.007318f
C1203 vdd.n426 gnd 0.009093f
C1204 vdd.n427 gnd 0.009093f
C1205 vdd.n428 gnd 0.009093f
C1206 vdd.n429 gnd 0.009093f
C1207 vdd.n430 gnd 0.009093f
C1208 vdd.n431 gnd 0.007318f
C1209 vdd.n433 gnd 0.009093f
C1210 vdd.n434 gnd 0.009093f
C1211 vdd.n435 gnd 0.009093f
C1212 vdd.n436 gnd 0.009093f
C1213 vdd.n437 gnd 0.009093f
C1214 vdd.n438 gnd 0.007318f
C1215 vdd.n440 gnd 0.009093f
C1216 vdd.n441 gnd 0.009093f
C1217 vdd.n442 gnd 0.009093f
C1218 vdd.n443 gnd 0.009093f
C1219 vdd.n444 gnd 0.009093f
C1220 vdd.n445 gnd 0.009093f
C1221 vdd.n446 gnd 0.007318f
C1222 vdd.n447 gnd 0.009093f
C1223 vdd.n448 gnd 0.009093f
C1224 vdd.n449 gnd 0.007318f
C1225 vdd.n450 gnd 0.009093f
C1226 vdd.n451 gnd 0.007318f
C1227 vdd.n452 gnd 0.009093f
C1228 vdd.n453 gnd 0.007318f
C1229 vdd.n454 gnd 0.009093f
C1230 vdd.n455 gnd 0.009093f
C1231 vdd.n456 gnd 0.506422f
C1232 vdd.t29 gnd 0.464607f
C1233 vdd.n457 gnd 0.009093f
C1234 vdd.n458 gnd 0.007318f
C1235 vdd.n459 gnd 0.009093f
C1236 vdd.n460 gnd 0.007318f
C1237 vdd.n461 gnd 0.009093f
C1238 vdd.t54 gnd 0.464607f
C1239 vdd.n462 gnd 0.009093f
C1240 vdd.n463 gnd 0.007318f
C1241 vdd.n464 gnd 0.009093f
C1242 vdd.n465 gnd 0.007318f
C1243 vdd.n466 gnd 0.009093f
C1244 vdd.t25 gnd 0.464607f
C1245 vdd.n467 gnd 0.580759f
C1246 vdd.n468 gnd 0.009093f
C1247 vdd.n469 gnd 0.007318f
C1248 vdd.n470 gnd 0.009093f
C1249 vdd.n471 gnd 0.007318f
C1250 vdd.n472 gnd 0.009093f
C1251 vdd.n473 gnd 0.929214f
C1252 vdd.n474 gnd 0.009093f
C1253 vdd.n475 gnd 0.007318f
C1254 vdd.n476 gnd 0.022159f
C1255 vdd.n477 gnd 0.006074f
C1256 vdd.n478 gnd 0.022159f
C1257 vdd.t125 gnd 0.464607f
C1258 vdd.n479 gnd 0.022159f
C1259 vdd.n480 gnd 0.006074f
C1260 vdd.n481 gnd 0.00782f
C1261 vdd.n482 gnd 0.007318f
C1262 vdd.n483 gnd 0.009093f
C1263 vdd.n484 gnd 6.40228f
C1264 vdd.n515 gnd 0.022667f
C1265 vdd.n516 gnd 1.27767f
C1266 vdd.n517 gnd 0.009093f
C1267 vdd.n518 gnd 0.007318f
C1268 vdd.n519 gnd 0.005819f
C1269 vdd.n520 gnd 0.014858f
C1270 vdd.n521 gnd 0.007318f
C1271 vdd.n522 gnd 0.009093f
C1272 vdd.n523 gnd 0.009093f
C1273 vdd.n524 gnd 0.009093f
C1274 vdd.n525 gnd 0.009093f
C1275 vdd.n526 gnd 0.009093f
C1276 vdd.n527 gnd 0.009093f
C1277 vdd.n528 gnd 0.009093f
C1278 vdd.n529 gnd 0.009093f
C1279 vdd.n530 gnd 0.009093f
C1280 vdd.n531 gnd 0.009093f
C1281 vdd.n532 gnd 0.009093f
C1282 vdd.n533 gnd 0.009093f
C1283 vdd.n534 gnd 0.009093f
C1284 vdd.n535 gnd 0.009093f
C1285 vdd.n536 gnd 0.006111f
C1286 vdd.n537 gnd 0.009093f
C1287 vdd.n538 gnd 0.009093f
C1288 vdd.n539 gnd 0.009093f
C1289 vdd.n540 gnd 0.009093f
C1290 vdd.n541 gnd 0.009093f
C1291 vdd.n542 gnd 0.009093f
C1292 vdd.n543 gnd 0.009093f
C1293 vdd.n544 gnd 0.009093f
C1294 vdd.n545 gnd 0.009093f
C1295 vdd.n546 gnd 0.009093f
C1296 vdd.n547 gnd 0.009093f
C1297 vdd.n548 gnd 0.009093f
C1298 vdd.n549 gnd 0.009093f
C1299 vdd.n550 gnd 0.009093f
C1300 vdd.n551 gnd 0.009093f
C1301 vdd.n552 gnd 0.009093f
C1302 vdd.n553 gnd 0.009093f
C1303 vdd.n554 gnd 0.009093f
C1304 vdd.n555 gnd 0.009093f
C1305 vdd.n556 gnd 0.007245f
C1306 vdd.t126 gnd 0.111862f
C1307 vdd.t127 gnd 0.11955f
C1308 vdd.t124 gnd 0.14609f
C1309 vdd.n557 gnd 0.187267f
C1310 vdd.n558 gnd 0.157338f
C1311 vdd.n559 gnd 0.009093f
C1312 vdd.n560 gnd 0.009093f
C1313 vdd.n561 gnd 0.009093f
C1314 vdd.n562 gnd 0.009093f
C1315 vdd.n563 gnd 0.009093f
C1316 vdd.n564 gnd 0.009093f
C1317 vdd.n565 gnd 0.009093f
C1318 vdd.n566 gnd 0.009093f
C1319 vdd.n567 gnd 0.009093f
C1320 vdd.n568 gnd 0.009093f
C1321 vdd.n569 gnd 0.009093f
C1322 vdd.n570 gnd 0.009093f
C1323 vdd.n571 gnd 0.009093f
C1324 vdd.n572 gnd 0.005819f
C1325 vdd.n575 gnd 0.006183f
C1326 vdd.n576 gnd 0.006183f
C1327 vdd.n577 gnd 0.006183f
C1328 vdd.n578 gnd 0.006183f
C1329 vdd.n579 gnd 0.006183f
C1330 vdd.n580 gnd 0.006183f
C1331 vdd.n582 gnd 0.006183f
C1332 vdd.n583 gnd 0.006183f
C1333 vdd.n585 gnd 0.006183f
C1334 vdd.n586 gnd 0.004501f
C1335 vdd.n588 gnd 0.006183f
C1336 vdd.t170 gnd 0.249851f
C1337 vdd.t169 gnd 0.255754f
C1338 vdd.t168 gnd 0.163112f
C1339 vdd.n589 gnd 0.088153f
C1340 vdd.n590 gnd 0.050003f
C1341 vdd.n591 gnd 0.008836f
C1342 vdd.n592 gnd 0.014451f
C1343 vdd.n594 gnd 0.006183f
C1344 vdd.n595 gnd 0.631866f
C1345 vdd.n596 gnd 0.013698f
C1346 vdd.n597 gnd 0.013698f
C1347 vdd.n598 gnd 0.006183f
C1348 vdd.n599 gnd 0.014671f
C1349 vdd.n600 gnd 0.006183f
C1350 vdd.n601 gnd 0.006183f
C1351 vdd.n602 gnd 0.006183f
C1352 vdd.n603 gnd 0.006183f
C1353 vdd.n604 gnd 0.006183f
C1354 vdd.n606 gnd 0.006183f
C1355 vdd.n607 gnd 0.006183f
C1356 vdd.n609 gnd 0.006183f
C1357 vdd.n610 gnd 0.006183f
C1358 vdd.n612 gnd 0.006183f
C1359 vdd.n613 gnd 0.006183f
C1360 vdd.n615 gnd 0.006183f
C1361 vdd.n616 gnd 0.006183f
C1362 vdd.n618 gnd 0.006183f
C1363 vdd.n619 gnd 0.006183f
C1364 vdd.n621 gnd 0.006183f
C1365 vdd.t163 gnd 0.249851f
C1366 vdd.t162 gnd 0.255754f
C1367 vdd.t160 gnd 0.163112f
C1368 vdd.n622 gnd 0.088153f
C1369 vdd.n623 gnd 0.050003f
C1370 vdd.n624 gnd 0.006183f
C1371 vdd.n626 gnd 0.006183f
C1372 vdd.n627 gnd 0.006183f
C1373 vdd.t161 gnd 0.315933f
C1374 vdd.n628 gnd 0.006183f
C1375 vdd.n629 gnd 0.006183f
C1376 vdd.n630 gnd 0.006183f
C1377 vdd.n631 gnd 0.006183f
C1378 vdd.n632 gnd 0.006183f
C1379 vdd.n633 gnd 0.631866f
C1380 vdd.n634 gnd 0.006183f
C1381 vdd.n635 gnd 0.006183f
C1382 vdd.n636 gnd 0.552882f
C1383 vdd.n637 gnd 0.006183f
C1384 vdd.n638 gnd 0.006183f
C1385 vdd.n639 gnd 0.005456f
C1386 vdd.n640 gnd 0.006183f
C1387 vdd.n641 gnd 0.557528f
C1388 vdd.n642 gnd 0.006183f
C1389 vdd.n643 gnd 0.006183f
C1390 vdd.n644 gnd 0.006183f
C1391 vdd.n645 gnd 0.006183f
C1392 vdd.n646 gnd 0.006183f
C1393 vdd.n647 gnd 0.631866f
C1394 vdd.n648 gnd 0.006183f
C1395 vdd.n649 gnd 0.006183f
C1396 vdd.t140 gnd 0.28341f
C1397 vdd.t19 gnd 0.074337f
C1398 vdd.n650 gnd 0.006183f
C1399 vdd.n651 gnd 0.006183f
C1400 vdd.n652 gnd 0.006183f
C1401 vdd.t120 gnd 0.315933f
C1402 vdd.n653 gnd 0.006183f
C1403 vdd.n654 gnd 0.006183f
C1404 vdd.n655 gnd 0.006183f
C1405 vdd.n656 gnd 0.006183f
C1406 vdd.n657 gnd 0.006183f
C1407 vdd.t20 gnd 0.315933f
C1408 vdd.n658 gnd 0.006183f
C1409 vdd.n659 gnd 0.006183f
C1410 vdd.n660 gnd 0.525006f
C1411 vdd.n661 gnd 0.006183f
C1412 vdd.n662 gnd 0.006183f
C1413 vdd.n663 gnd 0.006183f
C1414 vdd.n664 gnd 0.385624f
C1415 vdd.n665 gnd 0.006183f
C1416 vdd.n666 gnd 0.006183f
C1417 vdd.t17 gnd 0.315933f
C1418 vdd.n667 gnd 0.006183f
C1419 vdd.n668 gnd 0.006183f
C1420 vdd.n669 gnd 0.006183f
C1421 vdd.n670 gnd 0.525006f
C1422 vdd.n671 gnd 0.006183f
C1423 vdd.n672 gnd 0.006183f
C1424 vdd.t88 gnd 0.269472f
C1425 vdd.t109 gnd 0.246242f
C1426 vdd.n673 gnd 0.006183f
C1427 vdd.n674 gnd 0.006183f
C1428 vdd.n675 gnd 0.006183f
C1429 vdd.t4 gnd 0.315933f
C1430 vdd.n676 gnd 0.006183f
C1431 vdd.n677 gnd 0.006183f
C1432 vdd.t108 gnd 0.315933f
C1433 vdd.n678 gnd 0.006183f
C1434 vdd.n679 gnd 0.006183f
C1435 vdd.n680 gnd 0.006183f
C1436 vdd.t9 gnd 0.232304f
C1437 vdd.n681 gnd 0.006183f
C1438 vdd.n682 gnd 0.006183f
C1439 vdd.n683 gnd 0.538944f
C1440 vdd.n684 gnd 0.006183f
C1441 vdd.n685 gnd 0.006183f
C1442 vdd.n686 gnd 0.006183f
C1443 vdd.n687 gnd 0.631866f
C1444 vdd.n688 gnd 0.006183f
C1445 vdd.n689 gnd 0.006183f
C1446 vdd.t0 gnd 0.28341f
C1447 vdd.n690 gnd 0.399562f
C1448 vdd.n691 gnd 0.006183f
C1449 vdd.n692 gnd 0.006183f
C1450 vdd.n693 gnd 0.006183f
C1451 vdd.t10 gnd 0.315933f
C1452 vdd.n694 gnd 0.006183f
C1453 vdd.n695 gnd 0.006183f
C1454 vdd.n696 gnd 0.006183f
C1455 vdd.n697 gnd 0.006183f
C1456 vdd.n698 gnd 0.006183f
C1457 vdd.t21 gnd 0.631866f
C1458 vdd.n699 gnd 0.006183f
C1459 vdd.n700 gnd 0.006183f
C1460 vdd.t165 gnd 0.315933f
C1461 vdd.n701 gnd 0.006183f
C1462 vdd.n702 gnd 0.014671f
C1463 vdd.n703 gnd 0.014671f
C1464 vdd.t13 gnd 0.594697f
C1465 vdd.n704 gnd 0.013698f
C1466 vdd.n705 gnd 0.013698f
C1467 vdd.n706 gnd 0.014671f
C1468 vdd.n707 gnd 0.006183f
C1469 vdd.n708 gnd 0.006183f
C1470 vdd.t122 gnd 0.594697f
C1471 vdd.n726 gnd 0.014671f
C1472 vdd.n744 gnd 0.013698f
C1473 vdd.n745 gnd 0.006183f
C1474 vdd.n746 gnd 0.013698f
C1475 vdd.t190 gnd 0.249851f
C1476 vdd.t189 gnd 0.255754f
C1477 vdd.t188 gnd 0.163112f
C1478 vdd.n747 gnd 0.088153f
C1479 vdd.n748 gnd 0.050003f
C1480 vdd.n749 gnd 0.014451f
C1481 vdd.n750 gnd 0.006183f
C1482 vdd.t2 gnd 0.631866f
C1483 vdd.n751 gnd 0.013698f
C1484 vdd.n752 gnd 0.006183f
C1485 vdd.n753 gnd 0.014671f
C1486 vdd.n754 gnd 0.006183f
C1487 vdd.t159 gnd 0.249851f
C1488 vdd.t158 gnd 0.255754f
C1489 vdd.t156 gnd 0.163112f
C1490 vdd.n755 gnd 0.088153f
C1491 vdd.n756 gnd 0.050003f
C1492 vdd.n757 gnd 0.008836f
C1493 vdd.n758 gnd 0.006183f
C1494 vdd.n759 gnd 0.006183f
C1495 vdd.t157 gnd 0.315933f
C1496 vdd.n760 gnd 0.006183f
C1497 vdd.n761 gnd 0.006183f
C1498 vdd.n762 gnd 0.006183f
C1499 vdd.n763 gnd 0.006183f
C1500 vdd.n764 gnd 0.006183f
C1501 vdd.n765 gnd 0.006183f
C1502 vdd.n766 gnd 0.631866f
C1503 vdd.n767 gnd 0.006183f
C1504 vdd.n768 gnd 0.006183f
C1505 vdd.t7 gnd 0.315933f
C1506 vdd.n769 gnd 0.006183f
C1507 vdd.n770 gnd 0.006183f
C1508 vdd.n771 gnd 0.006183f
C1509 vdd.n772 gnd 0.006183f
C1510 vdd.n773 gnd 0.399562f
C1511 vdd.n774 gnd 0.006183f
C1512 vdd.n775 gnd 0.006183f
C1513 vdd.n776 gnd 0.006183f
C1514 vdd.n777 gnd 0.006183f
C1515 vdd.n778 gnd 0.006183f
C1516 vdd.n779 gnd 0.538944f
C1517 vdd.n780 gnd 0.006183f
C1518 vdd.n781 gnd 0.006183f
C1519 vdd.t116 gnd 0.28341f
C1520 vdd.t6 gnd 0.232304f
C1521 vdd.n782 gnd 0.006183f
C1522 vdd.n783 gnd 0.006183f
C1523 vdd.n784 gnd 0.006183f
C1524 vdd.t121 gnd 0.315933f
C1525 vdd.n785 gnd 0.006183f
C1526 vdd.n786 gnd 0.006183f
C1527 vdd.t106 gnd 0.315933f
C1528 vdd.n787 gnd 0.006183f
C1529 vdd.n788 gnd 0.006183f
C1530 vdd.n789 gnd 0.006183f
C1531 vdd.t15 gnd 0.246242f
C1532 vdd.n790 gnd 0.006183f
C1533 vdd.n791 gnd 0.006183f
C1534 vdd.n792 gnd 0.525006f
C1535 vdd.n793 gnd 0.006183f
C1536 vdd.n794 gnd 0.006183f
C1537 vdd.n795 gnd 0.006183f
C1538 vdd.t113 gnd 0.315933f
C1539 vdd.n796 gnd 0.006183f
C1540 vdd.n797 gnd 0.006183f
C1541 vdd.t105 gnd 0.269472f
C1542 vdd.n798 gnd 0.385624f
C1543 vdd.n799 gnd 0.006183f
C1544 vdd.n800 gnd 0.006183f
C1545 vdd.n801 gnd 0.006183f
C1546 vdd.n802 gnd 0.525006f
C1547 vdd.n803 gnd 0.006183f
C1548 vdd.n804 gnd 0.006183f
C1549 vdd.t87 gnd 0.315933f
C1550 vdd.n805 gnd 0.006183f
C1551 vdd.n806 gnd 0.006183f
C1552 vdd.n807 gnd 0.006183f
C1553 vdd.n808 gnd 0.631866f
C1554 vdd.n809 gnd 0.006183f
C1555 vdd.n810 gnd 0.006183f
C1556 vdd.t12 gnd 0.315933f
C1557 vdd.n811 gnd 0.006183f
C1558 vdd.n812 gnd 0.006183f
C1559 vdd.n813 gnd 0.006183f
C1560 vdd.t115 gnd 0.074337f
C1561 vdd.n814 gnd 0.006183f
C1562 vdd.n815 gnd 0.006183f
C1563 vdd.n816 gnd 0.006183f
C1564 vdd.t177 gnd 0.255754f
C1565 vdd.t175 gnd 0.163112f
C1566 vdd.t178 gnd 0.255754f
C1567 vdd.n817 gnd 0.143744f
C1568 vdd.n818 gnd 0.006183f
C1569 vdd.n819 gnd 0.006183f
C1570 vdd.n820 gnd 0.631866f
C1571 vdd.n821 gnd 0.006183f
C1572 vdd.n822 gnd 0.006183f
C1573 vdd.t176 gnd 0.28341f
C1574 vdd.n823 gnd 0.557528f
C1575 vdd.n824 gnd 0.006183f
C1576 vdd.n825 gnd 0.006183f
C1577 vdd.n826 gnd 0.006183f
C1578 vdd.n827 gnd 0.552882f
C1579 vdd.n828 gnd 0.006183f
C1580 vdd.n829 gnd 0.006183f
C1581 vdd.n830 gnd 0.006183f
C1582 vdd.n831 gnd 0.006183f
C1583 vdd.n832 gnd 0.006183f
C1584 vdd.n833 gnd 0.631866f
C1585 vdd.n834 gnd 0.006183f
C1586 vdd.n835 gnd 0.006183f
C1587 vdd.t172 gnd 0.315933f
C1588 vdd.n836 gnd 0.006183f
C1589 vdd.n837 gnd 0.014671f
C1590 vdd.n838 gnd 0.014671f
C1591 vdd.n839 gnd 6.40228f
C1592 vdd.n840 gnd 0.013698f
C1593 vdd.n841 gnd 0.013698f
C1594 vdd.n842 gnd 0.014671f
C1595 vdd.n843 gnd 0.006183f
C1596 vdd.n844 gnd 0.006183f
C1597 vdd.n845 gnd 0.006183f
C1598 vdd.n846 gnd 0.006183f
C1599 vdd.n847 gnd 0.006183f
C1600 vdd.n848 gnd 0.006183f
C1601 vdd.n849 gnd 0.006183f
C1602 vdd.n850 gnd 0.006183f
C1603 vdd.n852 gnd 0.006183f
C1604 vdd.n853 gnd 0.006183f
C1605 vdd.n854 gnd 0.005819f
C1606 vdd.n857 gnd 0.022667f
C1607 vdd.n858 gnd 0.007318f
C1608 vdd.n859 gnd 0.009093f
C1609 vdd.n861 gnd 0.009093f
C1610 vdd.n862 gnd 0.006074f
C1611 vdd.t132 gnd 0.464607f
C1612 vdd.n863 gnd 6.7368f
C1613 vdd.n864 gnd 0.009093f
C1614 vdd.n865 gnd 0.022667f
C1615 vdd.n866 gnd 0.007318f
C1616 vdd.n867 gnd 0.009093f
C1617 vdd.n868 gnd 0.007318f
C1618 vdd.n869 gnd 0.009093f
C1619 vdd.n870 gnd 0.929214f
C1620 vdd.n871 gnd 0.009093f
C1621 vdd.n872 gnd 0.007318f
C1622 vdd.n873 gnd 0.007318f
C1623 vdd.n874 gnd 0.009093f
C1624 vdd.n875 gnd 0.007318f
C1625 vdd.n876 gnd 0.009093f
C1626 vdd.t23 gnd 0.464607f
C1627 vdd.n877 gnd 0.009093f
C1628 vdd.n878 gnd 0.007318f
C1629 vdd.n879 gnd 0.009093f
C1630 vdd.n880 gnd 0.007318f
C1631 vdd.n881 gnd 0.009093f
C1632 vdd.t76 gnd 0.464607f
C1633 vdd.n882 gnd 0.009093f
C1634 vdd.n883 gnd 0.007318f
C1635 vdd.n884 gnd 0.009093f
C1636 vdd.n885 gnd 0.007318f
C1637 vdd.n886 gnd 0.009093f
C1638 vdd.n887 gnd 0.729433f
C1639 vdd.n888 gnd 0.771248f
C1640 vdd.t31 gnd 0.464607f
C1641 vdd.n889 gnd 0.009093f
C1642 vdd.n890 gnd 0.007318f
C1643 vdd.n891 gnd 0.00499f
C1644 vdd.n892 gnd 0.004631f
C1645 vdd.n893 gnd 0.002561f
C1646 vdd.n894 gnd 0.005881f
C1647 vdd.n895 gnd 0.002488f
C1648 vdd.n896 gnd 0.002635f
C1649 vdd.n897 gnd 0.004631f
C1650 vdd.n898 gnd 0.002488f
C1651 vdd.n899 gnd 0.005881f
C1652 vdd.n900 gnd 0.002635f
C1653 vdd.n901 gnd 0.004631f
C1654 vdd.n902 gnd 0.002488f
C1655 vdd.n903 gnd 0.004411f
C1656 vdd.n904 gnd 0.004424f
C1657 vdd.t24 gnd 0.012636f
C1658 vdd.n905 gnd 0.028114f
C1659 vdd.n906 gnd 0.146311f
C1660 vdd.n907 gnd 0.002488f
C1661 vdd.n908 gnd 0.002635f
C1662 vdd.n909 gnd 0.005881f
C1663 vdd.n910 gnd 0.005881f
C1664 vdd.n911 gnd 0.002635f
C1665 vdd.n912 gnd 0.002488f
C1666 vdd.n913 gnd 0.004631f
C1667 vdd.n914 gnd 0.004631f
C1668 vdd.n915 gnd 0.002488f
C1669 vdd.n916 gnd 0.002635f
C1670 vdd.n917 gnd 0.005881f
C1671 vdd.n918 gnd 0.005881f
C1672 vdd.n919 gnd 0.002635f
C1673 vdd.n920 gnd 0.002488f
C1674 vdd.n921 gnd 0.004631f
C1675 vdd.n922 gnd 0.004631f
C1676 vdd.n923 gnd 0.002488f
C1677 vdd.n924 gnd 0.002635f
C1678 vdd.n925 gnd 0.005881f
C1679 vdd.n926 gnd 0.005881f
C1680 vdd.n927 gnd 0.013905f
C1681 vdd.n928 gnd 0.002561f
C1682 vdd.n929 gnd 0.002488f
C1683 vdd.n930 gnd 0.011968f
C1684 vdd.n931 gnd 0.008356f
C1685 vdd.t50 gnd 0.029274f
C1686 vdd.t79 gnd 0.029274f
C1687 vdd.n932 gnd 0.201188f
C1688 vdd.n933 gnd 0.158204f
C1689 vdd.t39 gnd 0.029274f
C1690 vdd.t67 gnd 0.029274f
C1691 vdd.n934 gnd 0.201188f
C1692 vdd.n935 gnd 0.127669f
C1693 vdd.t45 gnd 0.029274f
C1694 vdd.t73 gnd 0.029274f
C1695 vdd.n936 gnd 0.201188f
C1696 vdd.n937 gnd 0.127669f
C1697 vdd.n938 gnd 0.00499f
C1698 vdd.n939 gnd 0.004631f
C1699 vdd.n940 gnd 0.002561f
C1700 vdd.n941 gnd 0.005881f
C1701 vdd.n942 gnd 0.002488f
C1702 vdd.n943 gnd 0.002635f
C1703 vdd.n944 gnd 0.004631f
C1704 vdd.n945 gnd 0.002488f
C1705 vdd.n946 gnd 0.005881f
C1706 vdd.n947 gnd 0.002635f
C1707 vdd.n948 gnd 0.004631f
C1708 vdd.n949 gnd 0.002488f
C1709 vdd.n950 gnd 0.004411f
C1710 vdd.n951 gnd 0.004424f
C1711 vdd.t83 gnd 0.012636f
C1712 vdd.n952 gnd 0.028114f
C1713 vdd.n953 gnd 0.146311f
C1714 vdd.n954 gnd 0.002488f
C1715 vdd.n955 gnd 0.002635f
C1716 vdd.n956 gnd 0.005881f
C1717 vdd.n957 gnd 0.005881f
C1718 vdd.n958 gnd 0.002635f
C1719 vdd.n959 gnd 0.002488f
C1720 vdd.n960 gnd 0.004631f
C1721 vdd.n961 gnd 0.004631f
C1722 vdd.n962 gnd 0.002488f
C1723 vdd.n963 gnd 0.002635f
C1724 vdd.n964 gnd 0.005881f
C1725 vdd.n965 gnd 0.005881f
C1726 vdd.n966 gnd 0.002635f
C1727 vdd.n967 gnd 0.002488f
C1728 vdd.n968 gnd 0.004631f
C1729 vdd.n969 gnd 0.004631f
C1730 vdd.n970 gnd 0.002488f
C1731 vdd.n971 gnd 0.002635f
C1732 vdd.n972 gnd 0.005881f
C1733 vdd.n973 gnd 0.005881f
C1734 vdd.n974 gnd 0.013905f
C1735 vdd.n975 gnd 0.002561f
C1736 vdd.n976 gnd 0.002488f
C1737 vdd.n977 gnd 0.011968f
C1738 vdd.n978 gnd 0.008094f
C1739 vdd.n979 gnd 0.094987f
C1740 vdd.n980 gnd 0.00499f
C1741 vdd.n981 gnd 0.004631f
C1742 vdd.n982 gnd 0.002561f
C1743 vdd.n983 gnd 0.005881f
C1744 vdd.n984 gnd 0.002488f
C1745 vdd.n985 gnd 0.002635f
C1746 vdd.n986 gnd 0.004631f
C1747 vdd.n987 gnd 0.002488f
C1748 vdd.n988 gnd 0.005881f
C1749 vdd.n989 gnd 0.002635f
C1750 vdd.n990 gnd 0.004631f
C1751 vdd.n991 gnd 0.002488f
C1752 vdd.n992 gnd 0.004411f
C1753 vdd.n993 gnd 0.004424f
C1754 vdd.t74 gnd 0.012636f
C1755 vdd.n994 gnd 0.028114f
C1756 vdd.n995 gnd 0.146311f
C1757 vdd.n996 gnd 0.002488f
C1758 vdd.n997 gnd 0.002635f
C1759 vdd.n998 gnd 0.005881f
C1760 vdd.n999 gnd 0.005881f
C1761 vdd.n1000 gnd 0.002635f
C1762 vdd.n1001 gnd 0.002488f
C1763 vdd.n1002 gnd 0.004631f
C1764 vdd.n1003 gnd 0.004631f
C1765 vdd.n1004 gnd 0.002488f
C1766 vdd.n1005 gnd 0.002635f
C1767 vdd.n1006 gnd 0.005881f
C1768 vdd.n1007 gnd 0.005881f
C1769 vdd.n1008 gnd 0.002635f
C1770 vdd.n1009 gnd 0.002488f
C1771 vdd.n1010 gnd 0.004631f
C1772 vdd.n1011 gnd 0.004631f
C1773 vdd.n1012 gnd 0.002488f
C1774 vdd.n1013 gnd 0.002635f
C1775 vdd.n1014 gnd 0.005881f
C1776 vdd.n1015 gnd 0.005881f
C1777 vdd.n1016 gnd 0.013905f
C1778 vdd.n1017 gnd 0.002561f
C1779 vdd.n1018 gnd 0.002488f
C1780 vdd.n1019 gnd 0.011968f
C1781 vdd.n1020 gnd 0.008356f
C1782 vdd.t32 gnd 0.029274f
C1783 vdd.t77 gnd 0.029274f
C1784 vdd.n1021 gnd 0.201188f
C1785 vdd.n1022 gnd 0.158204f
C1786 vdd.t72 gnd 0.029274f
C1787 vdd.t63 gnd 0.029274f
C1788 vdd.n1023 gnd 0.201188f
C1789 vdd.n1024 gnd 0.127669f
C1790 vdd.t48 gnd 0.029274f
C1791 vdd.t28 gnd 0.029274f
C1792 vdd.n1025 gnd 0.201188f
C1793 vdd.n1026 gnd 0.127669f
C1794 vdd.n1027 gnd 0.00499f
C1795 vdd.n1028 gnd 0.004631f
C1796 vdd.n1029 gnd 0.002561f
C1797 vdd.n1030 gnd 0.005881f
C1798 vdd.n1031 gnd 0.002488f
C1799 vdd.n1032 gnd 0.002635f
C1800 vdd.n1033 gnd 0.004631f
C1801 vdd.n1034 gnd 0.002488f
C1802 vdd.n1035 gnd 0.005881f
C1803 vdd.n1036 gnd 0.002635f
C1804 vdd.n1037 gnd 0.004631f
C1805 vdd.n1038 gnd 0.002488f
C1806 vdd.n1039 gnd 0.004411f
C1807 vdd.n1040 gnd 0.004424f
C1808 vdd.t61 gnd 0.012636f
C1809 vdd.n1041 gnd 0.028114f
C1810 vdd.n1042 gnd 0.146311f
C1811 vdd.n1043 gnd 0.002488f
C1812 vdd.n1044 gnd 0.002635f
C1813 vdd.n1045 gnd 0.005881f
C1814 vdd.n1046 gnd 0.005881f
C1815 vdd.n1047 gnd 0.002635f
C1816 vdd.n1048 gnd 0.002488f
C1817 vdd.n1049 gnd 0.004631f
C1818 vdd.n1050 gnd 0.004631f
C1819 vdd.n1051 gnd 0.002488f
C1820 vdd.n1052 gnd 0.002635f
C1821 vdd.n1053 gnd 0.005881f
C1822 vdd.n1054 gnd 0.005881f
C1823 vdd.n1055 gnd 0.002635f
C1824 vdd.n1056 gnd 0.002488f
C1825 vdd.n1057 gnd 0.004631f
C1826 vdd.n1058 gnd 0.004631f
C1827 vdd.n1059 gnd 0.002488f
C1828 vdd.n1060 gnd 0.002635f
C1829 vdd.n1061 gnd 0.005881f
C1830 vdd.n1062 gnd 0.005881f
C1831 vdd.n1063 gnd 0.013905f
C1832 vdd.n1064 gnd 0.002561f
C1833 vdd.n1065 gnd 0.002488f
C1834 vdd.n1066 gnd 0.011968f
C1835 vdd.n1067 gnd 0.008094f
C1836 vdd.n1068 gnd 0.056507f
C1837 vdd.n1069 gnd 0.203611f
C1838 vdd.n1070 gnd 0.00499f
C1839 vdd.n1071 gnd 0.004631f
C1840 vdd.n1072 gnd 0.002561f
C1841 vdd.n1073 gnd 0.005881f
C1842 vdd.n1074 gnd 0.002488f
C1843 vdd.n1075 gnd 0.002635f
C1844 vdd.n1076 gnd 0.004631f
C1845 vdd.n1077 gnd 0.002488f
C1846 vdd.n1078 gnd 0.005881f
C1847 vdd.n1079 gnd 0.002635f
C1848 vdd.n1080 gnd 0.004631f
C1849 vdd.n1081 gnd 0.002488f
C1850 vdd.n1082 gnd 0.004411f
C1851 vdd.n1083 gnd 0.004424f
C1852 vdd.t82 gnd 0.012636f
C1853 vdd.n1084 gnd 0.028114f
C1854 vdd.n1085 gnd 0.146311f
C1855 vdd.n1086 gnd 0.002488f
C1856 vdd.n1087 gnd 0.002635f
C1857 vdd.n1088 gnd 0.005881f
C1858 vdd.n1089 gnd 0.005881f
C1859 vdd.n1090 gnd 0.002635f
C1860 vdd.n1091 gnd 0.002488f
C1861 vdd.n1092 gnd 0.004631f
C1862 vdd.n1093 gnd 0.004631f
C1863 vdd.n1094 gnd 0.002488f
C1864 vdd.n1095 gnd 0.002635f
C1865 vdd.n1096 gnd 0.005881f
C1866 vdd.n1097 gnd 0.005881f
C1867 vdd.n1098 gnd 0.002635f
C1868 vdd.n1099 gnd 0.002488f
C1869 vdd.n1100 gnd 0.004631f
C1870 vdd.n1101 gnd 0.004631f
C1871 vdd.n1102 gnd 0.002488f
C1872 vdd.n1103 gnd 0.002635f
C1873 vdd.n1104 gnd 0.005881f
C1874 vdd.n1105 gnd 0.005881f
C1875 vdd.n1106 gnd 0.013905f
C1876 vdd.n1107 gnd 0.002561f
C1877 vdd.n1108 gnd 0.002488f
C1878 vdd.n1109 gnd 0.011968f
C1879 vdd.n1110 gnd 0.008356f
C1880 vdd.t37 gnd 0.029274f
C1881 vdd.t81 gnd 0.029274f
C1882 vdd.n1111 gnd 0.201188f
C1883 vdd.n1112 gnd 0.158204f
C1884 vdd.t80 gnd 0.029274f
C1885 vdd.t69 gnd 0.029274f
C1886 vdd.n1113 gnd 0.201188f
C1887 vdd.n1114 gnd 0.127669f
C1888 vdd.t56 gnd 0.029274f
C1889 vdd.t35 gnd 0.029274f
C1890 vdd.n1115 gnd 0.201188f
C1891 vdd.n1116 gnd 0.127669f
C1892 vdd.n1117 gnd 0.00499f
C1893 vdd.n1118 gnd 0.004631f
C1894 vdd.n1119 gnd 0.002561f
C1895 vdd.n1120 gnd 0.005881f
C1896 vdd.n1121 gnd 0.002488f
C1897 vdd.n1122 gnd 0.002635f
C1898 vdd.n1123 gnd 0.004631f
C1899 vdd.n1124 gnd 0.002488f
C1900 vdd.n1125 gnd 0.005881f
C1901 vdd.n1126 gnd 0.002635f
C1902 vdd.n1127 gnd 0.004631f
C1903 vdd.n1128 gnd 0.002488f
C1904 vdd.n1129 gnd 0.004411f
C1905 vdd.n1130 gnd 0.004424f
C1906 vdd.t68 gnd 0.012636f
C1907 vdd.n1131 gnd 0.028114f
C1908 vdd.n1132 gnd 0.146311f
C1909 vdd.n1133 gnd 0.002488f
C1910 vdd.n1134 gnd 0.002635f
C1911 vdd.n1135 gnd 0.005881f
C1912 vdd.n1136 gnd 0.005881f
C1913 vdd.n1137 gnd 0.002635f
C1914 vdd.n1138 gnd 0.002488f
C1915 vdd.n1139 gnd 0.004631f
C1916 vdd.n1140 gnd 0.004631f
C1917 vdd.n1141 gnd 0.002488f
C1918 vdd.n1142 gnd 0.002635f
C1919 vdd.n1143 gnd 0.005881f
C1920 vdd.n1144 gnd 0.005881f
C1921 vdd.n1145 gnd 0.002635f
C1922 vdd.n1146 gnd 0.002488f
C1923 vdd.n1147 gnd 0.004631f
C1924 vdd.n1148 gnd 0.004631f
C1925 vdd.n1149 gnd 0.002488f
C1926 vdd.n1150 gnd 0.002635f
C1927 vdd.n1151 gnd 0.005881f
C1928 vdd.n1152 gnd 0.005881f
C1929 vdd.n1153 gnd 0.013905f
C1930 vdd.n1154 gnd 0.002561f
C1931 vdd.n1155 gnd 0.002488f
C1932 vdd.n1156 gnd 0.011968f
C1933 vdd.n1157 gnd 0.008094f
C1934 vdd.n1158 gnd 0.056507f
C1935 vdd.n1159 gnd 0.220385f
C1936 vdd.n1160 gnd 1.85217f
C1937 vdd.n1161 gnd 0.536312f
C1938 vdd.n1162 gnd 0.007318f
C1939 vdd.n1163 gnd 0.009093f
C1940 vdd.n1164 gnd 0.571467f
C1941 vdd.n1165 gnd 0.009093f
C1942 vdd.n1166 gnd 0.007318f
C1943 vdd.n1167 gnd 0.009093f
C1944 vdd.n1168 gnd 0.007318f
C1945 vdd.n1169 gnd 0.009093f
C1946 vdd.t27 gnd 0.464607f
C1947 vdd.t38 gnd 0.464607f
C1948 vdd.n1170 gnd 0.009093f
C1949 vdd.n1171 gnd 0.007318f
C1950 vdd.n1172 gnd 0.009093f
C1951 vdd.n1173 gnd 0.007318f
C1952 vdd.n1174 gnd 0.009093f
C1953 vdd.t44 gnd 0.464607f
C1954 vdd.n1175 gnd 0.009093f
C1955 vdd.n1176 gnd 0.007318f
C1956 vdd.n1177 gnd 0.009093f
C1957 vdd.n1178 gnd 0.007318f
C1958 vdd.n1179 gnd 0.009093f
C1959 vdd.t60 gnd 0.464607f
C1960 vdd.n1180 gnd 0.67368f
C1961 vdd.n1181 gnd 0.009093f
C1962 vdd.n1182 gnd 0.007318f
C1963 vdd.n1183 gnd 0.009093f
C1964 vdd.n1184 gnd 0.007318f
C1965 vdd.n1185 gnd 0.009093f
C1966 vdd.n1186 gnd 0.929214f
C1967 vdd.n1187 gnd 0.009093f
C1968 vdd.n1188 gnd 0.007318f
C1969 vdd.n1189 gnd 0.022159f
C1970 vdd.n1190 gnd 0.006074f
C1971 vdd.n1191 gnd 0.022159f
C1972 vdd.t136 gnd 0.464607f
C1973 vdd.n1192 gnd 0.022159f
C1974 vdd.n1193 gnd 0.006074f
C1975 vdd.n1194 gnd 0.009093f
C1976 vdd.n1195 gnd 0.007318f
C1977 vdd.n1196 gnd 0.009093f
C1978 vdd.n1227 gnd 0.022667f
C1979 vdd.n1228 gnd 1.37059f
C1980 vdd.n1229 gnd 0.009093f
C1981 vdd.n1230 gnd 0.007318f
C1982 vdd.n1231 gnd 0.009093f
C1983 vdd.n1232 gnd 0.009093f
C1984 vdd.n1233 gnd 0.009093f
C1985 vdd.n1234 gnd 0.009093f
C1986 vdd.n1235 gnd 0.009093f
C1987 vdd.n1236 gnd 0.007318f
C1988 vdd.n1237 gnd 0.009093f
C1989 vdd.n1238 gnd 0.009093f
C1990 vdd.n1239 gnd 0.009093f
C1991 vdd.n1240 gnd 0.009093f
C1992 vdd.n1241 gnd 0.009093f
C1993 vdd.n1242 gnd 0.007318f
C1994 vdd.n1243 gnd 0.009093f
C1995 vdd.n1244 gnd 0.009093f
C1996 vdd.n1245 gnd 0.009093f
C1997 vdd.n1246 gnd 0.009093f
C1998 vdd.n1247 gnd 0.009093f
C1999 vdd.n1248 gnd 0.007318f
C2000 vdd.n1249 gnd 0.009093f
C2001 vdd.n1250 gnd 0.009093f
C2002 vdd.n1251 gnd 0.009093f
C2003 vdd.n1252 gnd 0.009093f
C2004 vdd.n1253 gnd 0.009093f
C2005 vdd.t186 gnd 0.111862f
C2006 vdd.t187 gnd 0.11955f
C2007 vdd.t185 gnd 0.14609f
C2008 vdd.n1254 gnd 0.187267f
C2009 vdd.n1255 gnd 0.15807f
C2010 vdd.n1256 gnd 0.015661f
C2011 vdd.n1257 gnd 0.009093f
C2012 vdd.n1258 gnd 0.009093f
C2013 vdd.n1259 gnd 0.009093f
C2014 vdd.n1260 gnd 0.009093f
C2015 vdd.n1261 gnd 0.009093f
C2016 vdd.n1262 gnd 0.007318f
C2017 vdd.n1263 gnd 0.009093f
C2018 vdd.n1264 gnd 0.009093f
C2019 vdd.n1265 gnd 0.009093f
C2020 vdd.n1266 gnd 0.009093f
C2021 vdd.n1267 gnd 0.009093f
C2022 vdd.n1268 gnd 0.007318f
C2023 vdd.n1269 gnd 0.009093f
C2024 vdd.n1270 gnd 0.009093f
C2025 vdd.n1271 gnd 0.009093f
C2026 vdd.n1272 gnd 0.009093f
C2027 vdd.n1273 gnd 0.009093f
C2028 vdd.n1274 gnd 0.007318f
C2029 vdd.n1275 gnd 0.009093f
C2030 vdd.n1276 gnd 0.009093f
C2031 vdd.n1277 gnd 0.009093f
C2032 vdd.n1278 gnd 0.009093f
C2033 vdd.n1279 gnd 0.009093f
C2034 vdd.n1280 gnd 0.007318f
C2035 vdd.n1281 gnd 0.009093f
C2036 vdd.n1282 gnd 0.009093f
C2037 vdd.n1283 gnd 0.009093f
C2038 vdd.n1284 gnd 0.009093f
C2039 vdd.n1285 gnd 0.009093f
C2040 vdd.n1286 gnd 0.007318f
C2041 vdd.n1287 gnd 0.009093f
C2042 vdd.n1288 gnd 0.009093f
C2043 vdd.n1289 gnd 0.009093f
C2044 vdd.n1290 gnd 0.009093f
C2045 vdd.n1291 gnd 0.007318f
C2046 vdd.n1292 gnd 0.009093f
C2047 vdd.n1293 gnd 0.009093f
C2048 vdd.n1294 gnd 0.009093f
C2049 vdd.n1295 gnd 0.009093f
C2050 vdd.n1296 gnd 0.009093f
C2051 vdd.n1297 gnd 0.007318f
C2052 vdd.n1298 gnd 0.009093f
C2053 vdd.n1299 gnd 0.009093f
C2054 vdd.n1300 gnd 0.009093f
C2055 vdd.n1301 gnd 0.009093f
C2056 vdd.n1302 gnd 0.009093f
C2057 vdd.n1303 gnd 0.007318f
C2058 vdd.n1304 gnd 0.009093f
C2059 vdd.n1305 gnd 0.009093f
C2060 vdd.n1306 gnd 0.009093f
C2061 vdd.n1307 gnd 0.009093f
C2062 vdd.n1308 gnd 0.009093f
C2063 vdd.n1309 gnd 0.007318f
C2064 vdd.n1310 gnd 0.009093f
C2065 vdd.n1311 gnd 0.009093f
C2066 vdd.n1312 gnd 0.009093f
C2067 vdd.n1313 gnd 0.009093f
C2068 vdd.n1314 gnd 0.009093f
C2069 vdd.n1315 gnd 0.007318f
C2070 vdd.n1316 gnd 0.009093f
C2071 vdd.n1317 gnd 0.009093f
C2072 vdd.n1318 gnd 0.009093f
C2073 vdd.n1319 gnd 0.009093f
C2074 vdd.t137 gnd 0.111862f
C2075 vdd.t138 gnd 0.11955f
C2076 vdd.t135 gnd 0.14609f
C2077 vdd.n1320 gnd 0.187267f
C2078 vdd.n1321 gnd 0.15807f
C2079 vdd.n1322 gnd 0.012002f
C2080 vdd.n1323 gnd 0.003476f
C2081 vdd.n1324 gnd 0.022667f
C2082 vdd.n1325 gnd 0.009093f
C2083 vdd.n1326 gnd 0.003842f
C2084 vdd.n1327 gnd 0.007318f
C2085 vdd.n1328 gnd 0.007318f
C2086 vdd.n1329 gnd 0.009093f
C2087 vdd.n1330 gnd 0.009093f
C2088 vdd.n1331 gnd 0.009093f
C2089 vdd.n1332 gnd 0.007318f
C2090 vdd.n1333 gnd 0.007318f
C2091 vdd.n1334 gnd 0.007318f
C2092 vdd.n1335 gnd 0.009093f
C2093 vdd.n1336 gnd 0.009093f
C2094 vdd.n1337 gnd 0.009093f
C2095 vdd.n1338 gnd 0.007318f
C2096 vdd.n1339 gnd 0.007318f
C2097 vdd.n1340 gnd 0.007318f
C2098 vdd.n1341 gnd 0.009093f
C2099 vdd.n1342 gnd 0.009093f
C2100 vdd.n1343 gnd 0.009093f
C2101 vdd.n1344 gnd 0.007318f
C2102 vdd.n1345 gnd 0.007318f
C2103 vdd.n1346 gnd 0.007318f
C2104 vdd.n1347 gnd 0.009093f
C2105 vdd.n1348 gnd 0.009093f
C2106 vdd.n1349 gnd 0.009093f
C2107 vdd.n1350 gnd 0.007318f
C2108 vdd.n1351 gnd 0.007318f
C2109 vdd.n1352 gnd 0.007318f
C2110 vdd.n1353 gnd 0.009093f
C2111 vdd.n1354 gnd 0.009093f
C2112 vdd.n1355 gnd 0.009093f
C2113 vdd.n1356 gnd 0.007245f
C2114 vdd.n1357 gnd 0.009093f
C2115 vdd.t183 gnd 0.111862f
C2116 vdd.t184 gnd 0.11955f
C2117 vdd.t182 gnd 0.14609f
C2118 vdd.n1358 gnd 0.187267f
C2119 vdd.n1359 gnd 0.15807f
C2120 vdd.n1360 gnd 0.015661f
C2121 vdd.n1361 gnd 0.004977f
C2122 vdd.n1362 gnd 0.009093f
C2123 vdd.n1363 gnd 0.009093f
C2124 vdd.n1364 gnd 0.009093f
C2125 vdd.n1365 gnd 0.007318f
C2126 vdd.n1366 gnd 0.007318f
C2127 vdd.n1367 gnd 0.007318f
C2128 vdd.n1368 gnd 0.009093f
C2129 vdd.n1369 gnd 0.009093f
C2130 vdd.n1370 gnd 0.009093f
C2131 vdd.n1371 gnd 0.007318f
C2132 vdd.n1372 gnd 0.007318f
C2133 vdd.n1373 gnd 0.007318f
C2134 vdd.n1374 gnd 0.009093f
C2135 vdd.n1375 gnd 0.009093f
C2136 vdd.n1376 gnd 0.009093f
C2137 vdd.n1377 gnd 0.007318f
C2138 vdd.n1378 gnd 0.007318f
C2139 vdd.n1379 gnd 0.007318f
C2140 vdd.n1380 gnd 0.009093f
C2141 vdd.n1381 gnd 0.009093f
C2142 vdd.n1382 gnd 0.009093f
C2143 vdd.n1383 gnd 0.007318f
C2144 vdd.n1384 gnd 0.007318f
C2145 vdd.n1385 gnd 0.007318f
C2146 vdd.n1386 gnd 0.009093f
C2147 vdd.n1387 gnd 0.009093f
C2148 vdd.n1388 gnd 0.009093f
C2149 vdd.n1389 gnd 0.007318f
C2150 vdd.n1390 gnd 0.007318f
C2151 vdd.n1391 gnd 0.006111f
C2152 vdd.n1392 gnd 0.009093f
C2153 vdd.n1393 gnd 0.009093f
C2154 vdd.n1394 gnd 0.009093f
C2155 vdd.n1395 gnd 0.006111f
C2156 vdd.n1396 gnd 0.007318f
C2157 vdd.n1397 gnd 0.007318f
C2158 vdd.n1398 gnd 0.009093f
C2159 vdd.n1399 gnd 0.009093f
C2160 vdd.n1400 gnd 0.009093f
C2161 vdd.n1401 gnd 0.007318f
C2162 vdd.n1402 gnd 0.007318f
C2163 vdd.n1403 gnd 0.007318f
C2164 vdd.n1404 gnd 0.009093f
C2165 vdd.n1405 gnd 0.009093f
C2166 vdd.n1406 gnd 0.009093f
C2167 vdd.n1407 gnd 0.007318f
C2168 vdd.n1408 gnd 0.007318f
C2169 vdd.n1409 gnd 0.007318f
C2170 vdd.n1410 gnd 0.009093f
C2171 vdd.n1411 gnd 0.009093f
C2172 vdd.n1412 gnd 0.009093f
C2173 vdd.n1413 gnd 0.007318f
C2174 vdd.n1414 gnd 0.007318f
C2175 vdd.n1415 gnd 0.007318f
C2176 vdd.n1416 gnd 0.009093f
C2177 vdd.n1417 gnd 0.009093f
C2178 vdd.n1418 gnd 0.009093f
C2179 vdd.n1419 gnd 0.007318f
C2180 vdd.n1420 gnd 0.009093f
C2181 vdd.n1421 gnd 2.22082f
C2182 vdd.n1423 gnd 0.022667f
C2183 vdd.n1424 gnd 0.006074f
C2184 vdd.n1425 gnd 0.022667f
C2185 vdd.n1426 gnd 0.022159f
C2186 vdd.n1427 gnd 0.009093f
C2187 vdd.n1428 gnd 0.007318f
C2188 vdd.n1429 gnd 0.009093f
C2189 vdd.n1430 gnd 0.487837f
C2190 vdd.n1431 gnd 0.009093f
C2191 vdd.n1432 gnd 0.007318f
C2192 vdd.n1433 gnd 0.009093f
C2193 vdd.n1434 gnd 0.009093f
C2194 vdd.n1435 gnd 0.009093f
C2195 vdd.n1436 gnd 0.007318f
C2196 vdd.n1437 gnd 0.009093f
C2197 vdd.n1438 gnd 0.831647f
C2198 vdd.n1439 gnd 0.929214f
C2199 vdd.n1440 gnd 0.009093f
C2200 vdd.n1441 gnd 0.007318f
C2201 vdd.n1442 gnd 0.009093f
C2202 vdd.n1443 gnd 0.009093f
C2203 vdd.n1444 gnd 0.009093f
C2204 vdd.n1445 gnd 0.007318f
C2205 vdd.n1446 gnd 0.009093f
C2206 vdd.n1447 gnd 0.562174f
C2207 vdd.n1448 gnd 0.009093f
C2208 vdd.n1449 gnd 0.007318f
C2209 vdd.n1450 gnd 0.009093f
C2210 vdd.n1451 gnd 0.009093f
C2211 vdd.n1452 gnd 0.009093f
C2212 vdd.n1453 gnd 0.007318f
C2213 vdd.n1454 gnd 0.009093f
C2214 vdd.n1455 gnd 0.515714f
C2215 vdd.n1456 gnd 0.720141f
C2216 vdd.n1457 gnd 0.009093f
C2217 vdd.n1458 gnd 0.007318f
C2218 vdd.n1459 gnd 0.009093f
C2219 vdd.n1460 gnd 0.009093f
C2220 vdd.n1461 gnd 0.006988f
C2221 vdd.n1462 gnd 0.009093f
C2222 vdd.n1463 gnd 0.007318f
C2223 vdd.n1464 gnd 0.009093f
C2224 vdd.n1465 gnd 0.771248f
C2225 vdd.n1466 gnd 0.009093f
C2226 vdd.n1467 gnd 0.007318f
C2227 vdd.n1468 gnd 0.009093f
C2228 vdd.n1469 gnd 0.009093f
C2229 vdd.n1470 gnd 0.009093f
C2230 vdd.n1471 gnd 0.007318f
C2231 vdd.n1472 gnd 0.009093f
C2232 vdd.t62 gnd 0.464607f
C2233 vdd.n1473 gnd 0.664388f
C2234 vdd.n1474 gnd 0.009093f
C2235 vdd.n1475 gnd 0.007318f
C2236 vdd.n1476 gnd 0.006988f
C2237 vdd.n1477 gnd 0.009093f
C2238 vdd.n1478 gnd 0.009093f
C2239 vdd.n1479 gnd 0.007318f
C2240 vdd.n1480 gnd 0.009093f
C2241 vdd.n1481 gnd 0.506422f
C2242 vdd.n1482 gnd 0.009093f
C2243 vdd.n1483 gnd 0.007318f
C2244 vdd.n1484 gnd 0.009093f
C2245 vdd.n1485 gnd 0.009093f
C2246 vdd.n1486 gnd 0.009093f
C2247 vdd.n1487 gnd 0.007318f
C2248 vdd.n1488 gnd 0.009093f
C2249 vdd.n1489 gnd 0.655096f
C2250 vdd.n1490 gnd 0.580759f
C2251 vdd.n1491 gnd 0.009093f
C2252 vdd.n1492 gnd 0.007318f
C2253 vdd.n1493 gnd 0.009093f
C2254 vdd.n1494 gnd 0.009093f
C2255 vdd.n1495 gnd 0.009093f
C2256 vdd.n1496 gnd 0.007318f
C2257 vdd.n1497 gnd 0.009093f
C2258 vdd.n1498 gnd 0.738725f
C2259 vdd.n1499 gnd 0.009093f
C2260 vdd.n1500 gnd 0.007318f
C2261 vdd.n1501 gnd 0.009093f
C2262 vdd.n1502 gnd 0.009093f
C2263 vdd.n1503 gnd 0.022159f
C2264 vdd.n1504 gnd 0.009093f
C2265 vdd.n1505 gnd 0.009093f
C2266 vdd.n1506 gnd 0.007318f
C2267 vdd.n1507 gnd 0.009093f
C2268 vdd.n1508 gnd 0.580759f
C2269 vdd.n1509 gnd 0.929214f
C2270 vdd.n1510 gnd 0.009093f
C2271 vdd.n1511 gnd 0.007318f
C2272 vdd.n1512 gnd 0.009093f
C2273 vdd.n1513 gnd 0.009093f
C2274 vdd.n1514 gnd 0.00782f
C2275 vdd.n1515 gnd 0.007318f
C2276 vdd.n1517 gnd 0.009093f
C2277 vdd.n1519 gnd 0.007318f
C2278 vdd.n1520 gnd 0.009093f
C2279 vdd.n1521 gnd 0.007318f
C2280 vdd.n1523 gnd 0.009093f
C2281 vdd.n1524 gnd 0.007318f
C2282 vdd.n1525 gnd 0.009093f
C2283 vdd.n1526 gnd 0.009093f
C2284 vdd.n1527 gnd 0.009093f
C2285 vdd.n1528 gnd 0.009093f
C2286 vdd.n1529 gnd 0.009093f
C2287 vdd.n1530 gnd 0.007318f
C2288 vdd.n1532 gnd 0.009093f
C2289 vdd.n1533 gnd 0.009093f
C2290 vdd.n1534 gnd 0.009093f
C2291 vdd.n1535 gnd 0.009093f
C2292 vdd.n1536 gnd 0.009093f
C2293 vdd.n1537 gnd 0.007318f
C2294 vdd.n1539 gnd 0.009093f
C2295 vdd.n1540 gnd 0.009093f
C2296 vdd.n1541 gnd 0.009093f
C2297 vdd.n1542 gnd 0.009093f
C2298 vdd.n1543 gnd 0.006111f
C2299 vdd.t152 gnd 0.111862f
C2300 vdd.t151 gnd 0.11955f
C2301 vdd.t150 gnd 0.14609f
C2302 vdd.n1544 gnd 0.187267f
C2303 vdd.n1545 gnd 0.157338f
C2304 vdd.n1547 gnd 0.009093f
C2305 vdd.n1548 gnd 0.009093f
C2306 vdd.n1549 gnd 0.007318f
C2307 vdd.n1550 gnd 0.009093f
C2308 vdd.n1552 gnd 0.009093f
C2309 vdd.n1553 gnd 0.009093f
C2310 vdd.n1554 gnd 0.009093f
C2311 vdd.n1555 gnd 0.009093f
C2312 vdd.n1556 gnd 0.007318f
C2313 vdd.n1558 gnd 0.009093f
C2314 vdd.n1559 gnd 0.009093f
C2315 vdd.n1560 gnd 0.009093f
C2316 vdd.n1561 gnd 0.009093f
C2317 vdd.n1562 gnd 0.009093f
C2318 vdd.n1563 gnd 0.007318f
C2319 vdd.n1565 gnd 0.009093f
C2320 vdd.n1566 gnd 0.009093f
C2321 vdd.n1567 gnd 0.009093f
C2322 vdd.n1568 gnd 0.009093f
C2323 vdd.n1569 gnd 0.009093f
C2324 vdd.n1570 gnd 0.007318f
C2325 vdd.n1572 gnd 0.009093f
C2326 vdd.n1573 gnd 0.009093f
C2327 vdd.n1574 gnd 0.009093f
C2328 vdd.n1575 gnd 0.009093f
C2329 vdd.n1576 gnd 0.009093f
C2330 vdd.n1577 gnd 0.007318f
C2331 vdd.n1579 gnd 0.009093f
C2332 vdd.n1580 gnd 0.009093f
C2333 vdd.n1581 gnd 0.009093f
C2334 vdd.n1582 gnd 0.009093f
C2335 vdd.n1583 gnd 0.007245f
C2336 vdd.t145 gnd 0.111862f
C2337 vdd.t144 gnd 0.11955f
C2338 vdd.t143 gnd 0.14609f
C2339 vdd.n1584 gnd 0.187267f
C2340 vdd.n1585 gnd 0.157338f
C2341 vdd.n1587 gnd 0.009093f
C2342 vdd.n1588 gnd 0.009093f
C2343 vdd.n1589 gnd 0.007318f
C2344 vdd.n1590 gnd 0.009093f
C2345 vdd.n1592 gnd 0.009093f
C2346 vdd.n1593 gnd 0.009093f
C2347 vdd.n1594 gnd 0.009093f
C2348 vdd.n1595 gnd 0.009093f
C2349 vdd.n1596 gnd 0.007318f
C2350 vdd.n1598 gnd 0.009093f
C2351 vdd.n1599 gnd 0.009093f
C2352 vdd.n1600 gnd 0.009093f
C2353 vdd.n1601 gnd 0.009093f
C2354 vdd.n1602 gnd 0.009093f
C2355 vdd.n1603 gnd 0.007318f
C2356 vdd.n1605 gnd 0.009093f
C2357 vdd.n1606 gnd 0.009093f
C2358 vdd.n1607 gnd 0.009093f
C2359 vdd.n1608 gnd 0.009093f
C2360 vdd.n1609 gnd 0.009093f
C2361 vdd.n1610 gnd 0.009093f
C2362 vdd.n1611 gnd 0.007318f
C2363 vdd.n1613 gnd 0.009093f
C2364 vdd.n1615 gnd 0.009093f
C2365 vdd.n1616 gnd 0.007318f
C2366 vdd.n1617 gnd 0.007318f
C2367 vdd.n1618 gnd 0.009093f
C2368 vdd.n1620 gnd 0.009093f
C2369 vdd.n1621 gnd 0.007318f
C2370 vdd.n1622 gnd 0.007318f
C2371 vdd.n1623 gnd 0.009093f
C2372 vdd.n1625 gnd 0.009093f
C2373 vdd.n1626 gnd 0.009093f
C2374 vdd.n1627 gnd 0.007318f
C2375 vdd.n1628 gnd 0.007318f
C2376 vdd.n1629 gnd 0.007318f
C2377 vdd.n1630 gnd 0.009093f
C2378 vdd.n1632 gnd 0.009093f
C2379 vdd.n1633 gnd 0.009093f
C2380 vdd.n1634 gnd 0.007318f
C2381 vdd.n1635 gnd 0.007318f
C2382 vdd.n1636 gnd 0.007318f
C2383 vdd.n1637 gnd 0.009093f
C2384 vdd.n1639 gnd 0.009093f
C2385 vdd.n1640 gnd 0.009093f
C2386 vdd.n1641 gnd 0.007318f
C2387 vdd.n1642 gnd 0.007318f
C2388 vdd.n1643 gnd 0.007318f
C2389 vdd.n1644 gnd 0.009093f
C2390 vdd.n1646 gnd 0.009093f
C2391 vdd.n1647 gnd 0.009093f
C2392 vdd.n1648 gnd 0.007318f
C2393 vdd.n1649 gnd 0.009093f
C2394 vdd.n1650 gnd 0.009093f
C2395 vdd.n1651 gnd 0.009093f
C2396 vdd.n1652 gnd 0.01493f
C2397 vdd.n1653 gnd 0.004977f
C2398 vdd.n1654 gnd 0.007318f
C2399 vdd.n1655 gnd 0.009093f
C2400 vdd.n1657 gnd 0.009093f
C2401 vdd.n1658 gnd 0.009093f
C2402 vdd.n1659 gnd 0.007318f
C2403 vdd.n1660 gnd 0.007318f
C2404 vdd.n1661 gnd 0.007318f
C2405 vdd.n1662 gnd 0.009093f
C2406 vdd.n1664 gnd 0.009093f
C2407 vdd.n1665 gnd 0.009093f
C2408 vdd.n1666 gnd 0.007318f
C2409 vdd.n1667 gnd 0.007318f
C2410 vdd.n1668 gnd 0.007318f
C2411 vdd.n1669 gnd 0.009093f
C2412 vdd.n1671 gnd 0.009093f
C2413 vdd.n1672 gnd 0.009093f
C2414 vdd.n1673 gnd 0.007318f
C2415 vdd.n1674 gnd 0.007318f
C2416 vdd.n1675 gnd 0.007318f
C2417 vdd.n1676 gnd 0.009093f
C2418 vdd.n1678 gnd 0.009093f
C2419 vdd.n1679 gnd 0.009093f
C2420 vdd.n1680 gnd 0.007318f
C2421 vdd.n1681 gnd 0.007318f
C2422 vdd.n1682 gnd 0.007318f
C2423 vdd.n1683 gnd 0.009093f
C2424 vdd.n1685 gnd 0.009093f
C2425 vdd.n1686 gnd 0.009093f
C2426 vdd.n1687 gnd 0.007318f
C2427 vdd.n1688 gnd 0.009093f
C2428 vdd.n1689 gnd 0.009093f
C2429 vdd.n1690 gnd 0.009093f
C2430 vdd.n1691 gnd 0.01493f
C2431 vdd.n1692 gnd 0.006111f
C2432 vdd.n1693 gnd 0.007318f
C2433 vdd.n1694 gnd 0.009093f
C2434 vdd.n1696 gnd 0.009093f
C2435 vdd.n1697 gnd 0.009093f
C2436 vdd.n1698 gnd 0.007318f
C2437 vdd.n1699 gnd 0.007318f
C2438 vdd.n1700 gnd 0.007318f
C2439 vdd.n1701 gnd 0.009093f
C2440 vdd.n1703 gnd 0.009093f
C2441 vdd.n1704 gnd 0.009093f
C2442 vdd.n1705 gnd 0.007318f
C2443 vdd.n1706 gnd 0.007318f
C2444 vdd.n1707 gnd 0.007318f
C2445 vdd.n1708 gnd 0.009093f
C2446 vdd.n1710 gnd 0.009093f
C2447 vdd.n1711 gnd 0.009093f
C2448 vdd.n1713 gnd 0.009093f
C2449 vdd.n1714 gnd 0.007318f
C2450 vdd.n1715 gnd 0.005819f
C2451 vdd.n1716 gnd 0.006183f
C2452 vdd.n1717 gnd 0.006183f
C2453 vdd.n1718 gnd 0.006183f
C2454 vdd.n1719 gnd 0.006183f
C2455 vdd.n1720 gnd 0.006183f
C2456 vdd.n1721 gnd 0.006183f
C2457 vdd.n1722 gnd 0.006183f
C2458 vdd.n1723 gnd 0.006183f
C2459 vdd.n1725 gnd 0.006183f
C2460 vdd.n1726 gnd 0.006183f
C2461 vdd.n1727 gnd 0.006183f
C2462 vdd.n1728 gnd 0.006183f
C2463 vdd.n1729 gnd 0.006183f
C2464 vdd.n1731 gnd 0.006183f
C2465 vdd.n1733 gnd 0.006183f
C2466 vdd.n1734 gnd 0.006183f
C2467 vdd.n1735 gnd 0.006183f
C2468 vdd.n1736 gnd 0.006183f
C2469 vdd.n1737 gnd 0.006183f
C2470 vdd.n1739 gnd 0.006183f
C2471 vdd.n1741 gnd 0.006183f
C2472 vdd.n1742 gnd 0.006183f
C2473 vdd.n1743 gnd 0.006183f
C2474 vdd.n1744 gnd 0.006183f
C2475 vdd.n1745 gnd 0.006183f
C2476 vdd.n1747 gnd 0.006183f
C2477 vdd.n1749 gnd 0.006183f
C2478 vdd.n1750 gnd 0.006183f
C2479 vdd.n1751 gnd 0.006183f
C2480 vdd.n1752 gnd 0.006183f
C2481 vdd.n1753 gnd 0.006183f
C2482 vdd.n1755 gnd 0.006183f
C2483 vdd.n1756 gnd 0.006183f
C2484 vdd.n1757 gnd 0.006183f
C2485 vdd.n1758 gnd 0.006183f
C2486 vdd.n1759 gnd 0.006183f
C2487 vdd.n1760 gnd 0.006183f
C2488 vdd.n1761 gnd 0.006183f
C2489 vdd.n1762 gnd 0.006183f
C2490 vdd.n1763 gnd 0.004501f
C2491 vdd.n1764 gnd 0.006183f
C2492 vdd.t198 gnd 0.249851f
C2493 vdd.t199 gnd 0.255754f
C2494 vdd.t197 gnd 0.163112f
C2495 vdd.n1765 gnd 0.088153f
C2496 vdd.n1766 gnd 0.050003f
C2497 vdd.n1767 gnd 0.008836f
C2498 vdd.n1768 gnd 0.006183f
C2499 vdd.n1769 gnd 0.006183f
C2500 vdd.n1770 gnd 0.376332f
C2501 vdd.n1771 gnd 0.006183f
C2502 vdd.n1772 gnd 0.006183f
C2503 vdd.n1773 gnd 0.006183f
C2504 vdd.n1774 gnd 0.006183f
C2505 vdd.n1775 gnd 0.006183f
C2506 vdd.n1776 gnd 0.006183f
C2507 vdd.n1777 gnd 0.006183f
C2508 vdd.n1778 gnd 0.006183f
C2509 vdd.n1779 gnd 0.006183f
C2510 vdd.n1780 gnd 0.006183f
C2511 vdd.n1781 gnd 0.006183f
C2512 vdd.n1782 gnd 0.006183f
C2513 vdd.n1783 gnd 0.006183f
C2514 vdd.n1784 gnd 0.006183f
C2515 vdd.n1785 gnd 0.006183f
C2516 vdd.n1786 gnd 0.006183f
C2517 vdd.n1787 gnd 0.006183f
C2518 vdd.n1788 gnd 0.006183f
C2519 vdd.n1789 gnd 0.006183f
C2520 vdd.n1790 gnd 0.006183f
C2521 vdd.t173 gnd 0.249851f
C2522 vdd.t174 gnd 0.255754f
C2523 vdd.t171 gnd 0.163112f
C2524 vdd.n1791 gnd 0.088153f
C2525 vdd.n1792 gnd 0.050003f
C2526 vdd.n1793 gnd 0.006183f
C2527 vdd.n1794 gnd 0.006183f
C2528 vdd.n1795 gnd 0.006183f
C2529 vdd.n1796 gnd 0.006183f
C2530 vdd.n1797 gnd 0.006183f
C2531 vdd.n1798 gnd 0.006183f
C2532 vdd.n1800 gnd 0.006183f
C2533 vdd.n1801 gnd 0.006183f
C2534 vdd.n1802 gnd 0.006183f
C2535 vdd.n1803 gnd 0.006183f
C2536 vdd.n1805 gnd 0.006183f
C2537 vdd.n1807 gnd 0.006183f
C2538 vdd.n1808 gnd 0.006183f
C2539 vdd.n1809 gnd 0.006183f
C2540 vdd.n1810 gnd 0.006183f
C2541 vdd.n1811 gnd 0.006183f
C2542 vdd.n1813 gnd 0.006183f
C2543 vdd.n1815 gnd 0.006183f
C2544 vdd.n1816 gnd 0.006183f
C2545 vdd.n1817 gnd 0.006183f
C2546 vdd.n1818 gnd 0.006183f
C2547 vdd.n1819 gnd 0.006183f
C2548 vdd.n1821 gnd 0.006183f
C2549 vdd.n1823 gnd 0.006183f
C2550 vdd.n1824 gnd 0.006183f
C2551 vdd.n1825 gnd 0.004501f
C2552 vdd.n1826 gnd 0.008836f
C2553 vdd.n1827 gnd 0.004774f
C2554 vdd.n1828 gnd 0.006183f
C2555 vdd.n1830 gnd 0.006183f
C2556 vdd.n1831 gnd 0.014671f
C2557 vdd.n1832 gnd 0.014671f
C2558 vdd.n1833 gnd 0.013698f
C2559 vdd.n1834 gnd 0.006183f
C2560 vdd.n1835 gnd 0.006183f
C2561 vdd.n1836 gnd 0.006183f
C2562 vdd.n1837 gnd 0.006183f
C2563 vdd.n1838 gnd 0.006183f
C2564 vdd.n1839 gnd 0.006183f
C2565 vdd.n1840 gnd 0.006183f
C2566 vdd.n1841 gnd 0.006183f
C2567 vdd.n1842 gnd 0.006183f
C2568 vdd.n1843 gnd 0.006183f
C2569 vdd.n1844 gnd 0.006183f
C2570 vdd.n1845 gnd 0.006183f
C2571 vdd.n1846 gnd 0.006183f
C2572 vdd.n1847 gnd 0.006183f
C2573 vdd.n1848 gnd 0.006183f
C2574 vdd.n1849 gnd 0.006183f
C2575 vdd.n1850 gnd 0.006183f
C2576 vdd.n1851 gnd 0.006183f
C2577 vdd.n1852 gnd 0.006183f
C2578 vdd.n1853 gnd 0.006183f
C2579 vdd.n1854 gnd 0.006183f
C2580 vdd.n1855 gnd 0.006183f
C2581 vdd.n1856 gnd 0.006183f
C2582 vdd.n1857 gnd 0.006183f
C2583 vdd.n1858 gnd 0.006183f
C2584 vdd.n1859 gnd 0.006183f
C2585 vdd.n1860 gnd 0.006183f
C2586 vdd.n1861 gnd 0.006183f
C2587 vdd.n1862 gnd 0.006183f
C2588 vdd.n1863 gnd 0.006183f
C2589 vdd.n1864 gnd 0.006183f
C2590 vdd.n1865 gnd 0.006183f
C2591 vdd.n1866 gnd 0.006183f
C2592 vdd.n1867 gnd 0.006183f
C2593 vdd.n1868 gnd 0.006183f
C2594 vdd.n1869 gnd 0.006183f
C2595 vdd.n1870 gnd 0.006183f
C2596 vdd.n1871 gnd 0.199781f
C2597 vdd.n1872 gnd 0.006183f
C2598 vdd.n1873 gnd 0.006183f
C2599 vdd.n1874 gnd 0.006183f
C2600 vdd.n1875 gnd 0.006183f
C2601 vdd.n1876 gnd 0.006183f
C2602 vdd.n1877 gnd 0.006183f
C2603 vdd.n1878 gnd 0.006183f
C2604 vdd.n1879 gnd 0.006183f
C2605 vdd.n1880 gnd 0.006183f
C2606 vdd.n1881 gnd 0.006183f
C2607 vdd.n1882 gnd 0.006183f
C2608 vdd.n1883 gnd 0.006183f
C2609 vdd.n1884 gnd 0.006183f
C2610 vdd.n1885 gnd 0.006183f
C2611 vdd.n1886 gnd 0.006183f
C2612 vdd.n1887 gnd 0.006183f
C2613 vdd.n1888 gnd 0.006183f
C2614 vdd.n1889 gnd 0.006183f
C2615 vdd.n1890 gnd 0.006183f
C2616 vdd.n1891 gnd 0.006183f
C2617 vdd.n1892 gnd 0.013698f
C2618 vdd.n1894 gnd 0.014671f
C2619 vdd.n1895 gnd 0.014671f
C2620 vdd.n1896 gnd 0.006183f
C2621 vdd.n1897 gnd 0.004774f
C2622 vdd.n1898 gnd 0.006183f
C2623 vdd.n1900 gnd 0.006183f
C2624 vdd.n1902 gnd 0.006183f
C2625 vdd.n1903 gnd 0.006183f
C2626 vdd.n1904 gnd 0.006183f
C2627 vdd.n1905 gnd 0.006183f
C2628 vdd.n1906 gnd 0.006183f
C2629 vdd.n1908 gnd 0.006183f
C2630 vdd.n1910 gnd 0.006183f
C2631 vdd.n1911 gnd 0.006183f
C2632 vdd.n1912 gnd 0.006183f
C2633 vdd.n1913 gnd 0.006183f
C2634 vdd.n1914 gnd 0.006183f
C2635 vdd.n1916 gnd 0.006183f
C2636 vdd.n1918 gnd 0.006183f
C2637 vdd.n1919 gnd 0.006183f
C2638 vdd.n1920 gnd 0.006183f
C2639 vdd.n1921 gnd 0.006183f
C2640 vdd.n1922 gnd 0.006183f
C2641 vdd.n1924 gnd 0.006183f
C2642 vdd.n1926 gnd 0.006183f
C2643 vdd.n1927 gnd 0.006183f
C2644 vdd.n1928 gnd 0.018442f
C2645 vdd.n1929 gnd 0.546711f
C2646 vdd.n1931 gnd 0.007318f
C2647 vdd.n1932 gnd 0.007318f
C2648 vdd.n1933 gnd 0.009093f
C2649 vdd.n1935 gnd 0.009093f
C2650 vdd.n1936 gnd 0.009093f
C2651 vdd.n1937 gnd 0.007318f
C2652 vdd.n1938 gnd 0.006074f
C2653 vdd.n1939 gnd 0.022667f
C2654 vdd.n1940 gnd 0.022159f
C2655 vdd.n1941 gnd 0.006074f
C2656 vdd.n1942 gnd 0.022159f
C2657 vdd.n1943 gnd 1.27767f
C2658 vdd.n1944 gnd 0.022159f
C2659 vdd.n1945 gnd 0.022667f
C2660 vdd.n1946 gnd 0.003476f
C2661 vdd.t134 gnd 0.111862f
C2662 vdd.t133 gnd 0.11955f
C2663 vdd.t131 gnd 0.14609f
C2664 vdd.n1947 gnd 0.187267f
C2665 vdd.n1948 gnd 0.157338f
C2666 vdd.n1949 gnd 0.01127f
C2667 vdd.n1950 gnd 0.003842f
C2668 vdd.n1951 gnd 0.00782f
C2669 vdd.n1952 gnd 0.546711f
C2670 vdd.n1953 gnd 0.018442f
C2671 vdd.n1954 gnd 0.006183f
C2672 vdd.n1955 gnd 0.006183f
C2673 vdd.n1956 gnd 0.006183f
C2674 vdd.n1958 gnd 0.006183f
C2675 vdd.n1960 gnd 0.006183f
C2676 vdd.n1961 gnd 0.006183f
C2677 vdd.n1962 gnd 0.006183f
C2678 vdd.n1963 gnd 0.006183f
C2679 vdd.n1964 gnd 0.006183f
C2680 vdd.n1966 gnd 0.006183f
C2681 vdd.n1968 gnd 0.006183f
C2682 vdd.n1969 gnd 0.006183f
C2683 vdd.n1970 gnd 0.006183f
C2684 vdd.n1971 gnd 0.006183f
C2685 vdd.n1972 gnd 0.006183f
C2686 vdd.n1974 gnd 0.006183f
C2687 vdd.n1976 gnd 0.006183f
C2688 vdd.n1977 gnd 0.006183f
C2689 vdd.n1978 gnd 0.006183f
C2690 vdd.n1979 gnd 0.006183f
C2691 vdd.n1980 gnd 0.006183f
C2692 vdd.n1982 gnd 0.006183f
C2693 vdd.n1984 gnd 0.006183f
C2694 vdd.n1985 gnd 0.006183f
C2695 vdd.n1986 gnd 0.014671f
C2696 vdd.n1987 gnd 0.013698f
C2697 vdd.n1988 gnd 0.013698f
C2698 vdd.n1989 gnd 0.91063f
C2699 vdd.n1990 gnd 0.013698f
C2700 vdd.n1991 gnd 0.013698f
C2701 vdd.n1992 gnd 0.006183f
C2702 vdd.n1993 gnd 0.006183f
C2703 vdd.n1994 gnd 0.006183f
C2704 vdd.n1995 gnd 0.394916f
C2705 vdd.n1996 gnd 0.006183f
C2706 vdd.n1997 gnd 0.006183f
C2707 vdd.n1998 gnd 0.006183f
C2708 vdd.n1999 gnd 0.006183f
C2709 vdd.n2000 gnd 0.006183f
C2710 vdd.n2001 gnd 0.631866f
C2711 vdd.n2002 gnd 0.006183f
C2712 vdd.n2003 gnd 0.006183f
C2713 vdd.n2004 gnd 0.006183f
C2714 vdd.n2005 gnd 0.006183f
C2715 vdd.n2006 gnd 0.006183f
C2716 vdd.n2007 gnd 0.631866f
C2717 vdd.n2008 gnd 0.006183f
C2718 vdd.n2009 gnd 0.006183f
C2719 vdd.n2010 gnd 0.005456f
C2720 vdd.n2011 gnd 0.017911f
C2721 vdd.n2012 gnd 0.003819f
C2722 vdd.n2013 gnd 0.006183f
C2723 vdd.n2014 gnd 0.348455f
C2724 vdd.n2015 gnd 0.006183f
C2725 vdd.n2016 gnd 0.006183f
C2726 vdd.n2017 gnd 0.006183f
C2727 vdd.n2018 gnd 0.006183f
C2728 vdd.n2019 gnd 0.006183f
C2729 vdd.n2020 gnd 0.422792f
C2730 vdd.n2021 gnd 0.006183f
C2731 vdd.n2022 gnd 0.006183f
C2732 vdd.n2023 gnd 0.006183f
C2733 vdd.n2024 gnd 0.006183f
C2734 vdd.n2025 gnd 0.006183f
C2735 vdd.n2026 gnd 0.562174f
C2736 vdd.n2027 gnd 0.006183f
C2737 vdd.n2028 gnd 0.006183f
C2738 vdd.n2029 gnd 0.006183f
C2739 vdd.n2030 gnd 0.006183f
C2740 vdd.n2031 gnd 0.006183f
C2741 vdd.n2032 gnd 0.501776f
C2742 vdd.n2033 gnd 0.006183f
C2743 vdd.n2034 gnd 0.006183f
C2744 vdd.n2035 gnd 0.006183f
C2745 vdd.n2036 gnd 0.006183f
C2746 vdd.n2037 gnd 0.006183f
C2747 vdd.n2038 gnd 0.362393f
C2748 vdd.n2039 gnd 0.006183f
C2749 vdd.n2040 gnd 0.006183f
C2750 vdd.n2041 gnd 0.006183f
C2751 vdd.n2042 gnd 0.006183f
C2752 vdd.n2043 gnd 0.006183f
C2753 vdd.n2044 gnd 0.199781f
C2754 vdd.n2045 gnd 0.006183f
C2755 vdd.n2046 gnd 0.006183f
C2756 vdd.n2047 gnd 0.006183f
C2757 vdd.n2048 gnd 0.006183f
C2758 vdd.n2049 gnd 0.006183f
C2759 vdd.n2050 gnd 0.348455f
C2760 vdd.n2051 gnd 0.006183f
C2761 vdd.n2052 gnd 0.006183f
C2762 vdd.n2053 gnd 0.006183f
C2763 vdd.n2054 gnd 0.006183f
C2764 vdd.n2055 gnd 0.006183f
C2765 vdd.n2056 gnd 0.631866f
C2766 vdd.n2057 gnd 0.006183f
C2767 vdd.n2058 gnd 0.006183f
C2768 vdd.n2059 gnd 0.006183f
C2769 vdd.n2060 gnd 0.006183f
C2770 vdd.n2061 gnd 0.006183f
C2771 vdd.n2062 gnd 0.006183f
C2772 vdd.n2063 gnd 0.006183f
C2773 vdd.n2064 gnd 0.492483f
C2774 vdd.n2065 gnd 0.006183f
C2775 vdd.n2066 gnd 0.006183f
C2776 vdd.n2067 gnd 0.006183f
C2777 vdd.n2068 gnd 0.006183f
C2778 vdd.n2069 gnd 0.006183f
C2779 vdd.n2070 gnd 0.006183f
C2780 vdd.n2071 gnd 0.394916f
C2781 vdd.n2072 gnd 0.006183f
C2782 vdd.n2073 gnd 0.006183f
C2783 vdd.n2074 gnd 0.006183f
C2784 vdd.n2075 gnd 0.014451f
C2785 vdd.n2076 gnd 0.013918f
C2786 vdd.n2077 gnd 0.006183f
C2787 vdd.n2078 gnd 0.006183f
C2788 vdd.n2079 gnd 0.004774f
C2789 vdd.n2080 gnd 0.006183f
C2790 vdd.n2081 gnd 0.006183f
C2791 vdd.n2082 gnd 0.004501f
C2792 vdd.n2083 gnd 0.006183f
C2793 vdd.n2084 gnd 0.006183f
C2794 vdd.n2085 gnd 0.006183f
C2795 vdd.n2086 gnd 0.006183f
C2796 vdd.n2087 gnd 0.006183f
C2797 vdd.n2088 gnd 0.006183f
C2798 vdd.n2089 gnd 0.006183f
C2799 vdd.n2090 gnd 0.006183f
C2800 vdd.n2091 gnd 0.006183f
C2801 vdd.n2092 gnd 0.006183f
C2802 vdd.n2093 gnd 0.006183f
C2803 vdd.n2094 gnd 0.006183f
C2804 vdd.n2095 gnd 0.006183f
C2805 vdd.n2096 gnd 0.006183f
C2806 vdd.n2097 gnd 0.006183f
C2807 vdd.n2098 gnd 0.006183f
C2808 vdd.n2099 gnd 0.006183f
C2809 vdd.n2100 gnd 0.006183f
C2810 vdd.n2101 gnd 0.006183f
C2811 vdd.n2102 gnd 0.006183f
C2812 vdd.n2103 gnd 0.006183f
C2813 vdd.n2104 gnd 0.006183f
C2814 vdd.n2105 gnd 0.006183f
C2815 vdd.n2106 gnd 0.006183f
C2816 vdd.n2107 gnd 0.006183f
C2817 vdd.n2108 gnd 0.006183f
C2818 vdd.n2109 gnd 0.006183f
C2819 vdd.n2110 gnd 0.006183f
C2820 vdd.n2111 gnd 0.006183f
C2821 vdd.n2112 gnd 0.006183f
C2822 vdd.n2113 gnd 0.006183f
C2823 vdd.n2114 gnd 0.006183f
C2824 vdd.n2115 gnd 0.006183f
C2825 vdd.n2116 gnd 0.006183f
C2826 vdd.n2117 gnd 0.006183f
C2827 vdd.n2118 gnd 0.006183f
C2828 vdd.n2119 gnd 0.006183f
C2829 vdd.n2120 gnd 0.006183f
C2830 vdd.n2121 gnd 0.006183f
C2831 vdd.n2122 gnd 0.006183f
C2832 vdd.n2123 gnd 0.006183f
C2833 vdd.n2124 gnd 0.006183f
C2834 vdd.n2125 gnd 0.006183f
C2835 vdd.n2126 gnd 0.006183f
C2836 vdd.n2127 gnd 0.006183f
C2837 vdd.n2128 gnd 0.006183f
C2838 vdd.n2129 gnd 0.006183f
C2839 vdd.n2130 gnd 0.006183f
C2840 vdd.n2131 gnd 0.006183f
C2841 vdd.n2132 gnd 0.006183f
C2842 vdd.n2133 gnd 0.006183f
C2843 vdd.n2134 gnd 0.006183f
C2844 vdd.n2135 gnd 0.006183f
C2845 vdd.n2136 gnd 0.006183f
C2846 vdd.n2137 gnd 0.006183f
C2847 vdd.n2138 gnd 0.006183f
C2848 vdd.n2139 gnd 0.006183f
C2849 vdd.n2140 gnd 0.006183f
C2850 vdd.n2141 gnd 0.006183f
C2851 vdd.n2142 gnd 0.006183f
C2852 vdd.n2143 gnd 0.014671f
C2853 vdd.n2144 gnd 0.013698f
C2854 vdd.n2145 gnd 0.013698f
C2855 vdd.n2146 gnd 0.771248f
C2856 vdd.n2147 gnd 0.013698f
C2857 vdd.n2148 gnd 0.014671f
C2858 vdd.n2149 gnd 0.013918f
C2859 vdd.n2150 gnd 0.006183f
C2860 vdd.n2151 gnd 0.006183f
C2861 vdd.n2152 gnd 0.006183f
C2862 vdd.n2153 gnd 0.004774f
C2863 vdd.n2154 gnd 0.008836f
C2864 vdd.n2155 gnd 0.004501f
C2865 vdd.n2156 gnd 0.006183f
C2866 vdd.n2157 gnd 0.006183f
C2867 vdd.n2158 gnd 0.006183f
C2868 vdd.n2159 gnd 0.006183f
C2869 vdd.n2160 gnd 0.006183f
C2870 vdd.n2161 gnd 0.006183f
C2871 vdd.n2162 gnd 0.006183f
C2872 vdd.n2163 gnd 0.006183f
C2873 vdd.n2164 gnd 0.006183f
C2874 vdd.n2165 gnd 0.006183f
C2875 vdd.n2166 gnd 0.006183f
C2876 vdd.n2167 gnd 0.006183f
C2877 vdd.n2168 gnd 0.006183f
C2878 vdd.n2169 gnd 0.006183f
C2879 vdd.n2170 gnd 0.006183f
C2880 vdd.n2171 gnd 0.006183f
C2881 vdd.n2172 gnd 0.006183f
C2882 vdd.n2173 gnd 0.006183f
C2883 vdd.n2174 gnd 0.006183f
C2884 vdd.n2175 gnd 0.006183f
C2885 vdd.n2176 gnd 0.006183f
C2886 vdd.n2177 gnd 0.006183f
C2887 vdd.n2178 gnd 0.006183f
C2888 vdd.n2179 gnd 0.006183f
C2889 vdd.n2180 gnd 0.006183f
C2890 vdd.n2181 gnd 0.006183f
C2891 vdd.n2182 gnd 0.006183f
C2892 vdd.n2183 gnd 0.006183f
C2893 vdd.n2184 gnd 0.006183f
C2894 vdd.n2185 gnd 0.006183f
C2895 vdd.n2186 gnd 0.006183f
C2896 vdd.n2187 gnd 0.006183f
C2897 vdd.n2188 gnd 0.006183f
C2898 vdd.n2189 gnd 0.006183f
C2899 vdd.n2190 gnd 0.006183f
C2900 vdd.n2191 gnd 0.006183f
C2901 vdd.n2192 gnd 0.006183f
C2902 vdd.n2193 gnd 0.006183f
C2903 vdd.n2194 gnd 0.006183f
C2904 vdd.n2195 gnd 0.006183f
C2905 vdd.n2196 gnd 0.006183f
C2906 vdd.n2197 gnd 0.006183f
C2907 vdd.n2198 gnd 0.006183f
C2908 vdd.n2199 gnd 0.006183f
C2909 vdd.n2200 gnd 0.006183f
C2910 vdd.n2201 gnd 0.006183f
C2911 vdd.n2202 gnd 0.006183f
C2912 vdd.n2203 gnd 0.006183f
C2913 vdd.n2204 gnd 0.006183f
C2914 vdd.n2205 gnd 0.006183f
C2915 vdd.n2206 gnd 0.006183f
C2916 vdd.n2207 gnd 0.006183f
C2917 vdd.n2208 gnd 0.006183f
C2918 vdd.n2209 gnd 0.006183f
C2919 vdd.n2210 gnd 0.006183f
C2920 vdd.n2211 gnd 0.006183f
C2921 vdd.n2212 gnd 0.006183f
C2922 vdd.n2213 gnd 0.006183f
C2923 vdd.n2214 gnd 0.006183f
C2924 vdd.n2215 gnd 0.006183f
C2925 vdd.n2216 gnd 0.014671f
C2926 vdd.n2217 gnd 0.014671f
C2927 vdd.n2218 gnd 0.771248f
C2928 vdd.t111 gnd 2.74118f
C2929 vdd.t118 gnd 2.74118f
C2930 vdd.n2251 gnd 0.014671f
C2931 vdd.n2252 gnd 0.006183f
C2932 vdd.t166 gnd 0.249851f
C2933 vdd.t167 gnd 0.255754f
C2934 vdd.t164 gnd 0.163112f
C2935 vdd.n2253 gnd 0.088153f
C2936 vdd.n2254 gnd 0.050003f
C2937 vdd.n2255 gnd 0.006183f
C2938 vdd.t180 gnd 0.249851f
C2939 vdd.t181 gnd 0.255754f
C2940 vdd.t179 gnd 0.163112f
C2941 vdd.n2256 gnd 0.088153f
C2942 vdd.n2257 gnd 0.050003f
C2943 vdd.n2258 gnd 0.008836f
C2944 vdd.n2259 gnd 0.006183f
C2945 vdd.n2260 gnd 0.006183f
C2946 vdd.n2261 gnd 0.006183f
C2947 vdd.n2262 gnd 0.006183f
C2948 vdd.n2263 gnd 0.006183f
C2949 vdd.n2264 gnd 0.006183f
C2950 vdd.n2265 gnd 0.006183f
C2951 vdd.n2266 gnd 0.006183f
C2952 vdd.n2267 gnd 0.006183f
C2953 vdd.n2268 gnd 0.006183f
C2954 vdd.n2269 gnd 0.006183f
C2955 vdd.n2270 gnd 0.006183f
C2956 vdd.n2271 gnd 0.006183f
C2957 vdd.n2272 gnd 0.006183f
C2958 vdd.n2273 gnd 0.006183f
C2959 vdd.n2274 gnd 0.006183f
C2960 vdd.n2275 gnd 0.006183f
C2961 vdd.n2276 gnd 0.006183f
C2962 vdd.n2277 gnd 0.006183f
C2963 vdd.n2278 gnd 0.006183f
C2964 vdd.n2279 gnd 0.006183f
C2965 vdd.n2280 gnd 0.006183f
C2966 vdd.n2281 gnd 0.006183f
C2967 vdd.n2282 gnd 0.006183f
C2968 vdd.n2283 gnd 0.006183f
C2969 vdd.n2284 gnd 0.006183f
C2970 vdd.n2285 gnd 0.006183f
C2971 vdd.n2286 gnd 0.006183f
C2972 vdd.n2287 gnd 0.006183f
C2973 vdd.n2288 gnd 0.006183f
C2974 vdd.n2289 gnd 0.006183f
C2975 vdd.n2290 gnd 0.006183f
C2976 vdd.n2291 gnd 0.006183f
C2977 vdd.n2292 gnd 0.006183f
C2978 vdd.n2293 gnd 0.006183f
C2979 vdd.n2294 gnd 0.006183f
C2980 vdd.n2295 gnd 0.006183f
C2981 vdd.n2296 gnd 0.006183f
C2982 vdd.n2297 gnd 0.006183f
C2983 vdd.n2298 gnd 0.006183f
C2984 vdd.n2299 gnd 0.006183f
C2985 vdd.n2300 gnd 0.006183f
C2986 vdd.n2301 gnd 0.006183f
C2987 vdd.n2302 gnd 0.006183f
C2988 vdd.n2303 gnd 0.006183f
C2989 vdd.n2304 gnd 0.006183f
C2990 vdd.n2305 gnd 0.006183f
C2991 vdd.n2306 gnd 0.006183f
C2992 vdd.n2307 gnd 0.006183f
C2993 vdd.n2308 gnd 0.006183f
C2994 vdd.n2309 gnd 0.006183f
C2995 vdd.n2310 gnd 0.006183f
C2996 vdd.n2311 gnd 0.006183f
C2997 vdd.n2312 gnd 0.006183f
C2998 vdd.n2313 gnd 0.006183f
C2999 vdd.n2314 gnd 0.006183f
C3000 vdd.n2315 gnd 0.004501f
C3001 vdd.n2316 gnd 0.006183f
C3002 vdd.n2317 gnd 0.006183f
C3003 vdd.n2318 gnd 0.004774f
C3004 vdd.n2319 gnd 0.006183f
C3005 vdd.n2320 gnd 0.006183f
C3006 vdd.n2321 gnd 0.014671f
C3007 vdd.n2322 gnd 0.013698f
C3008 vdd.n2323 gnd 0.006183f
C3009 vdd.n2324 gnd 0.006183f
C3010 vdd.n2325 gnd 0.006183f
C3011 vdd.n2326 gnd 0.006183f
C3012 vdd.n2327 gnd 0.006183f
C3013 vdd.n2328 gnd 0.006183f
C3014 vdd.n2329 gnd 0.006183f
C3015 vdd.n2330 gnd 0.006183f
C3016 vdd.n2331 gnd 0.006183f
C3017 vdd.n2332 gnd 0.006183f
C3018 vdd.n2333 gnd 0.006183f
C3019 vdd.n2334 gnd 0.006183f
C3020 vdd.n2335 gnd 0.006183f
C3021 vdd.n2336 gnd 0.006183f
C3022 vdd.n2337 gnd 0.006183f
C3023 vdd.n2338 gnd 0.006183f
C3024 vdd.n2339 gnd 0.006183f
C3025 vdd.n2340 gnd 0.006183f
C3026 vdd.n2341 gnd 0.006183f
C3027 vdd.n2342 gnd 0.006183f
C3028 vdd.n2343 gnd 0.006183f
C3029 vdd.n2344 gnd 0.006183f
C3030 vdd.n2345 gnd 0.006183f
C3031 vdd.n2346 gnd 0.006183f
C3032 vdd.n2347 gnd 0.006183f
C3033 vdd.n2348 gnd 0.006183f
C3034 vdd.n2349 gnd 0.006183f
C3035 vdd.n2350 gnd 0.006183f
C3036 vdd.n2351 gnd 0.006183f
C3037 vdd.n2352 gnd 0.006183f
C3038 vdd.n2353 gnd 0.006183f
C3039 vdd.n2354 gnd 0.006183f
C3040 vdd.n2355 gnd 0.006183f
C3041 vdd.n2356 gnd 0.006183f
C3042 vdd.n2357 gnd 0.006183f
C3043 vdd.n2358 gnd 0.006183f
C3044 vdd.n2359 gnd 0.006183f
C3045 vdd.n2360 gnd 0.006183f
C3046 vdd.n2361 gnd 0.006183f
C3047 vdd.n2362 gnd 0.006183f
C3048 vdd.n2363 gnd 0.006183f
C3049 vdd.n2364 gnd 0.006183f
C3050 vdd.n2365 gnd 0.006183f
C3051 vdd.n2366 gnd 0.006183f
C3052 vdd.n2367 gnd 0.006183f
C3053 vdd.n2368 gnd 0.006183f
C3054 vdd.n2369 gnd 0.006183f
C3055 vdd.n2370 gnd 0.006183f
C3056 vdd.n2371 gnd 0.006183f
C3057 vdd.n2372 gnd 0.006183f
C3058 vdd.n2373 gnd 0.006183f
C3059 vdd.n2374 gnd 0.199781f
C3060 vdd.n2375 gnd 0.006183f
C3061 vdd.n2376 gnd 0.006183f
C3062 vdd.n2377 gnd 0.006183f
C3063 vdd.n2378 gnd 0.006183f
C3064 vdd.n2379 gnd 0.006183f
C3065 vdd.n2380 gnd 0.006183f
C3066 vdd.n2381 gnd 0.006183f
C3067 vdd.n2382 gnd 0.006183f
C3068 vdd.n2383 gnd 0.006183f
C3069 vdd.n2384 gnd 0.006183f
C3070 vdd.n2385 gnd 0.006183f
C3071 vdd.n2386 gnd 0.006183f
C3072 vdd.n2387 gnd 0.006183f
C3073 vdd.n2388 gnd 0.006183f
C3074 vdd.n2389 gnd 0.006183f
C3075 vdd.n2390 gnd 0.006183f
C3076 vdd.n2391 gnd 0.006183f
C3077 vdd.n2392 gnd 0.006183f
C3078 vdd.n2393 gnd 0.006183f
C3079 vdd.n2394 gnd 0.006183f
C3080 vdd.n2395 gnd 0.376332f
C3081 vdd.n2396 gnd 0.006183f
C3082 vdd.n2397 gnd 0.006183f
C3083 vdd.n2398 gnd 0.006183f
C3084 vdd.n2399 gnd 0.006183f
C3085 vdd.n2400 gnd 0.006183f
C3086 vdd.n2401 gnd 0.013698f
C3087 vdd.n2402 gnd 0.014671f
C3088 vdd.n2403 gnd 0.014671f
C3089 vdd.n2404 gnd 0.006183f
C3090 vdd.n2405 gnd 0.006183f
C3091 vdd.n2406 gnd 0.006183f
C3092 vdd.n2407 gnd 0.004774f
C3093 vdd.n2408 gnd 0.008836f
C3094 vdd.n2409 gnd 0.004501f
C3095 vdd.n2410 gnd 0.006183f
C3096 vdd.n2411 gnd 0.006183f
C3097 vdd.n2412 gnd 0.006183f
C3098 vdd.n2413 gnd 0.006183f
C3099 vdd.n2414 gnd 0.006183f
C3100 vdd.n2415 gnd 0.006183f
C3101 vdd.n2416 gnd 0.006183f
C3102 vdd.n2417 gnd 0.006183f
C3103 vdd.n2418 gnd 0.006183f
C3104 vdd.n2419 gnd 0.006183f
C3105 vdd.n2420 gnd 0.006183f
C3106 vdd.n2421 gnd 0.006183f
C3107 vdd.n2422 gnd 0.006183f
C3108 vdd.n2423 gnd 0.006183f
C3109 vdd.n2424 gnd 0.006183f
C3110 vdd.n2425 gnd 0.006183f
C3111 vdd.n2426 gnd 0.006183f
C3112 vdd.n2427 gnd 0.006183f
C3113 vdd.n2428 gnd 0.006183f
C3114 vdd.n2429 gnd 0.006183f
C3115 vdd.n2430 gnd 0.006183f
C3116 vdd.n2431 gnd 0.006183f
C3117 vdd.n2432 gnd 0.006183f
C3118 vdd.n2433 gnd 0.006183f
C3119 vdd.n2434 gnd 0.006183f
C3120 vdd.n2435 gnd 0.006183f
C3121 vdd.n2436 gnd 0.006183f
C3122 vdd.n2437 gnd 0.006183f
C3123 vdd.n2438 gnd 0.006183f
C3124 vdd.n2439 gnd 0.006183f
C3125 vdd.n2440 gnd 0.006183f
C3126 vdd.n2441 gnd 0.006183f
C3127 vdd.n2442 gnd 0.006183f
C3128 vdd.n2443 gnd 0.006183f
C3129 vdd.n2444 gnd 0.006183f
C3130 vdd.n2445 gnd 0.006183f
C3131 vdd.n2446 gnd 0.006183f
C3132 vdd.n2447 gnd 0.006183f
C3133 vdd.n2448 gnd 0.006183f
C3134 vdd.n2449 gnd 0.006183f
C3135 vdd.n2450 gnd 0.006183f
C3136 vdd.n2451 gnd 0.006183f
C3137 vdd.n2452 gnd 0.006183f
C3138 vdd.n2453 gnd 0.006183f
C3139 vdd.n2454 gnd 0.006183f
C3140 vdd.n2455 gnd 0.006183f
C3141 vdd.n2456 gnd 0.006183f
C3142 vdd.n2457 gnd 0.006183f
C3143 vdd.n2458 gnd 0.006183f
C3144 vdd.n2459 gnd 0.006183f
C3145 vdd.n2460 gnd 0.006183f
C3146 vdd.n2461 gnd 0.006183f
C3147 vdd.n2462 gnd 0.006183f
C3148 vdd.n2463 gnd 0.006183f
C3149 vdd.n2464 gnd 0.006183f
C3150 vdd.n2465 gnd 0.006183f
C3151 vdd.n2466 gnd 0.006183f
C3152 vdd.n2467 gnd 0.006183f
C3153 vdd.n2468 gnd 0.006183f
C3154 vdd.n2469 gnd 0.006183f
C3155 vdd.n2471 gnd 0.771248f
C3156 vdd.n2473 gnd 0.006183f
C3157 vdd.n2474 gnd 0.006183f
C3158 vdd.n2475 gnd 0.014671f
C3159 vdd.n2476 gnd 0.013698f
C3160 vdd.n2477 gnd 0.013698f
C3161 vdd.n2478 gnd 0.771248f
C3162 vdd.n2479 gnd 0.013698f
C3163 vdd.n2480 gnd 0.013698f
C3164 vdd.n2481 gnd 0.006183f
C3165 vdd.n2482 gnd 0.006183f
C3166 vdd.n2483 gnd 0.006183f
C3167 vdd.n2484 gnd 0.394916f
C3168 vdd.n2485 gnd 0.006183f
C3169 vdd.n2486 gnd 0.006183f
C3170 vdd.n2487 gnd 0.006183f
C3171 vdd.n2488 gnd 0.006183f
C3172 vdd.n2489 gnd 0.006183f
C3173 vdd.n2490 gnd 0.492483f
C3174 vdd.n2491 gnd 0.006183f
C3175 vdd.n2492 gnd 0.006183f
C3176 vdd.n2493 gnd 0.006183f
C3177 vdd.n2494 gnd 0.006183f
C3178 vdd.n2495 gnd 0.006183f
C3179 vdd.n2496 gnd 0.631866f
C3180 vdd.n2497 gnd 0.006183f
C3181 vdd.n2498 gnd 0.006183f
C3182 vdd.n2499 gnd 0.006183f
C3183 vdd.n2500 gnd 0.006183f
C3184 vdd.n2501 gnd 0.006183f
C3185 vdd.n2502 gnd 0.348455f
C3186 vdd.n2503 gnd 0.006183f
C3187 vdd.n2504 gnd 0.006183f
C3188 vdd.n2505 gnd 0.006183f
C3189 vdd.n2506 gnd 0.006183f
C3190 vdd.n2507 gnd 0.006183f
C3191 vdd.n2508 gnd 0.199781f
C3192 vdd.n2509 gnd 0.006183f
C3193 vdd.n2510 gnd 0.006183f
C3194 vdd.n2511 gnd 0.006183f
C3195 vdd.n2512 gnd 0.006183f
C3196 vdd.n2513 gnd 0.006183f
C3197 vdd.n2514 gnd 0.362393f
C3198 vdd.n2515 gnd 0.006183f
C3199 vdd.n2516 gnd 0.006183f
C3200 vdd.n2517 gnd 0.006183f
C3201 vdd.n2518 gnd 0.006183f
C3202 vdd.n2519 gnd 0.006183f
C3203 vdd.n2520 gnd 0.501776f
C3204 vdd.n2521 gnd 0.006183f
C3205 vdd.n2522 gnd 0.006183f
C3206 vdd.n2523 gnd 0.006183f
C3207 vdd.n2524 gnd 0.006183f
C3208 vdd.n2525 gnd 0.006183f
C3209 vdd.n2526 gnd 0.562174f
C3210 vdd.n2527 gnd 0.006183f
C3211 vdd.n2528 gnd 0.006183f
C3212 vdd.n2529 gnd 0.006183f
C3213 vdd.n2530 gnd 0.006183f
C3214 vdd.n2531 gnd 0.006183f
C3215 vdd.n2532 gnd 0.422792f
C3216 vdd.n2533 gnd 0.006183f
C3217 vdd.n2534 gnd 0.006183f
C3218 vdd.n2535 gnd 0.006183f
C3219 vdd.t141 gnd 0.255754f
C3220 vdd.t139 gnd 0.163112f
C3221 vdd.t142 gnd 0.255754f
C3222 vdd.n2536 gnd 0.143744f
C3223 vdd.n2537 gnd 0.017911f
C3224 vdd.n2538 gnd 0.003819f
C3225 vdd.n2539 gnd 0.006183f
C3226 vdd.n2540 gnd 0.348455f
C3227 vdd.n2541 gnd 0.006183f
C3228 vdd.n2542 gnd 0.006183f
C3229 vdd.n2543 gnd 0.006183f
C3230 vdd.n2544 gnd 0.006183f
C3231 vdd.n2545 gnd 0.006183f
C3232 vdd.n2546 gnd 0.631866f
C3233 vdd.n2547 gnd 0.006183f
C3234 vdd.n2548 gnd 0.006183f
C3235 vdd.n2549 gnd 0.006183f
C3236 vdd.n2550 gnd 0.006183f
C3237 vdd.n2551 gnd 0.006183f
C3238 vdd.n2552 gnd 0.006183f
C3239 vdd.n2554 gnd 0.006183f
C3240 vdd.n2555 gnd 0.006183f
C3241 vdd.n2557 gnd 0.006183f
C3242 vdd.n2558 gnd 0.006183f
C3243 vdd.n2561 gnd 0.006183f
C3244 vdd.n2562 gnd 0.006183f
C3245 vdd.n2563 gnd 0.006183f
C3246 vdd.n2564 gnd 0.006183f
C3247 vdd.n2566 gnd 0.006183f
C3248 vdd.n2567 gnd 0.006183f
C3249 vdd.n2568 gnd 0.006183f
C3250 vdd.n2569 gnd 0.006183f
C3251 vdd.n2570 gnd 0.006183f
C3252 vdd.n2571 gnd 0.006183f
C3253 vdd.n2573 gnd 0.006183f
C3254 vdd.n2574 gnd 0.006183f
C3255 vdd.n2575 gnd 0.006183f
C3256 vdd.n2576 gnd 0.006183f
C3257 vdd.n2577 gnd 0.006183f
C3258 vdd.n2578 gnd 0.006183f
C3259 vdd.n2580 gnd 0.006183f
C3260 vdd.n2581 gnd 0.006183f
C3261 vdd.n2582 gnd 0.006183f
C3262 vdd.n2583 gnd 0.006183f
C3263 vdd.n2584 gnd 0.006183f
C3264 vdd.n2585 gnd 0.006183f
C3265 vdd.n2587 gnd 0.006183f
C3266 vdd.n2588 gnd 0.014671f
C3267 vdd.n2589 gnd 0.014671f
C3268 vdd.n2590 gnd 0.013698f
C3269 vdd.n2591 gnd 0.006183f
C3270 vdd.n2592 gnd 0.006183f
C3271 vdd.n2593 gnd 0.006183f
C3272 vdd.n2594 gnd 0.006183f
C3273 vdd.n2595 gnd 0.006183f
C3274 vdd.n2596 gnd 0.006183f
C3275 vdd.n2597 gnd 0.631866f
C3276 vdd.n2598 gnd 0.006183f
C3277 vdd.n2599 gnd 0.006183f
C3278 vdd.n2600 gnd 0.006183f
C3279 vdd.n2601 gnd 0.006183f
C3280 vdd.n2602 gnd 0.006183f
C3281 vdd.n2603 gnd 0.394916f
C3282 vdd.n2604 gnd 0.006183f
C3283 vdd.n2605 gnd 0.006183f
C3284 vdd.n2606 gnd 0.006183f
C3285 vdd.n2607 gnd 0.014451f
C3286 vdd.n2608 gnd 0.013918f
C3287 vdd.n2609 gnd 0.014671f
C3288 vdd.n2611 gnd 0.006183f
C3289 vdd.n2612 gnd 0.006183f
C3290 vdd.n2613 gnd 0.004774f
C3291 vdd.n2614 gnd 0.008836f
C3292 vdd.n2615 gnd 0.004501f
C3293 vdd.n2616 gnd 0.006183f
C3294 vdd.n2617 gnd 0.006183f
C3295 vdd.n2619 gnd 0.006183f
C3296 vdd.n2620 gnd 0.006183f
C3297 vdd.n2621 gnd 0.006183f
C3298 vdd.n2622 gnd 0.006183f
C3299 vdd.n2623 gnd 0.006183f
C3300 vdd.n2624 gnd 0.006183f
C3301 vdd.n2626 gnd 0.006183f
C3302 vdd.n2627 gnd 0.006183f
C3303 vdd.n2628 gnd 0.006183f
C3304 vdd.n2629 gnd 0.006183f
C3305 vdd.n2630 gnd 0.006183f
C3306 vdd.n2631 gnd 0.006183f
C3307 vdd.n2633 gnd 0.006183f
C3308 vdd.n2634 gnd 0.006183f
C3309 vdd.n2635 gnd 0.006183f
C3310 vdd.n2636 gnd 0.006183f
C3311 vdd.n2637 gnd 0.006183f
C3312 vdd.n2638 gnd 0.006183f
C3313 vdd.n2640 gnd 0.006183f
C3314 vdd.n2641 gnd 0.006183f
C3315 vdd.n2642 gnd 0.006183f
C3316 vdd.n2644 gnd 0.006183f
C3317 vdd.n2645 gnd 0.006183f
C3318 vdd.n2646 gnd 0.006183f
C3319 vdd.n2647 gnd 0.006183f
C3320 vdd.n2648 gnd 0.006183f
C3321 vdd.n2649 gnd 0.006183f
C3322 vdd.n2651 gnd 0.006183f
C3323 vdd.n2652 gnd 0.006183f
C3324 vdd.n2653 gnd 0.006183f
C3325 vdd.n2654 gnd 0.006183f
C3326 vdd.n2655 gnd 0.006183f
C3327 vdd.n2656 gnd 0.006183f
C3328 vdd.n2658 gnd 0.006183f
C3329 vdd.n2659 gnd 0.006183f
C3330 vdd.n2660 gnd 0.006183f
C3331 vdd.n2661 gnd 0.006183f
C3332 vdd.n2662 gnd 0.006183f
C3333 vdd.n2663 gnd 0.006183f
C3334 vdd.n2665 gnd 0.006183f
C3335 vdd.n2666 gnd 0.006183f
C3336 vdd.n2668 gnd 0.006183f
C3337 vdd.n2669 gnd 0.006183f
C3338 vdd.n2670 gnd 0.014671f
C3339 vdd.n2671 gnd 0.013698f
C3340 vdd.n2672 gnd 0.013698f
C3341 vdd.n2673 gnd 0.91063f
C3342 vdd.n2674 gnd 0.013698f
C3343 vdd.n2675 gnd 0.014671f
C3344 vdd.n2676 gnd 0.013918f
C3345 vdd.n2677 gnd 0.006183f
C3346 vdd.n2678 gnd 0.004774f
C3347 vdd.n2679 gnd 0.006183f
C3348 vdd.n2681 gnd 0.006183f
C3349 vdd.n2682 gnd 0.006183f
C3350 vdd.n2683 gnd 0.006183f
C3351 vdd.n2684 gnd 0.006183f
C3352 vdd.n2685 gnd 0.006183f
C3353 vdd.n2686 gnd 0.006183f
C3354 vdd.n2688 gnd 0.006183f
C3355 vdd.n2689 gnd 0.006183f
C3356 vdd.n2690 gnd 0.006183f
C3357 vdd.n2691 gnd 0.006183f
C3358 vdd.n2692 gnd 0.006183f
C3359 vdd.n2693 gnd 0.006183f
C3360 vdd.n2695 gnd 0.006183f
C3361 vdd.n2696 gnd 0.006183f
C3362 vdd.n2697 gnd 0.006183f
C3363 vdd.n2698 gnd 0.006183f
C3364 vdd.n2699 gnd 0.006183f
C3365 vdd.n2700 gnd 0.006183f
C3366 vdd.n2702 gnd 0.006183f
C3367 vdd.n2703 gnd 0.006183f
C3368 vdd.n2705 gnd 0.006183f
C3369 vdd.n2706 gnd 0.014858f
C3370 vdd.n2707 gnd 0.550295f
C3371 vdd.n2708 gnd 0.00782f
C3372 vdd.n2709 gnd 0.022667f
C3373 vdd.n2710 gnd 0.003476f
C3374 vdd.t192 gnd 0.111862f
C3375 vdd.t193 gnd 0.11955f
C3376 vdd.t191 gnd 0.14609f
C3377 vdd.n2711 gnd 0.187267f
C3378 vdd.n2712 gnd 0.157338f
C3379 vdd.n2713 gnd 0.01127f
C3380 vdd.n2714 gnd 0.009093f
C3381 vdd.n2715 gnd 0.003842f
C3382 vdd.n2716 gnd 0.007318f
C3383 vdd.n2717 gnd 0.009093f
C3384 vdd.n2718 gnd 0.009093f
C3385 vdd.n2719 gnd 0.007318f
C3386 vdd.n2720 gnd 0.007318f
C3387 vdd.n2721 gnd 0.009093f
C3388 vdd.n2722 gnd 0.009093f
C3389 vdd.n2723 gnd 0.007318f
C3390 vdd.n2724 gnd 0.007318f
C3391 vdd.n2725 gnd 0.009093f
C3392 vdd.n2726 gnd 0.009093f
C3393 vdd.n2727 gnd 0.007318f
C3394 vdd.n2728 gnd 0.007318f
C3395 vdd.n2729 gnd 0.009093f
C3396 vdd.n2730 gnd 0.009093f
C3397 vdd.n2731 gnd 0.007318f
C3398 vdd.n2732 gnd 0.007318f
C3399 vdd.n2733 gnd 0.009093f
C3400 vdd.n2734 gnd 0.009093f
C3401 vdd.n2735 gnd 0.007318f
C3402 vdd.n2736 gnd 0.007318f
C3403 vdd.n2737 gnd 0.009093f
C3404 vdd.n2738 gnd 0.009093f
C3405 vdd.n2739 gnd 0.007318f
C3406 vdd.n2740 gnd 0.007318f
C3407 vdd.n2741 gnd 0.009093f
C3408 vdd.n2742 gnd 0.009093f
C3409 vdd.n2743 gnd 0.007318f
C3410 vdd.n2744 gnd 0.007318f
C3411 vdd.n2745 gnd 0.009093f
C3412 vdd.n2746 gnd 0.009093f
C3413 vdd.n2747 gnd 0.007318f
C3414 vdd.n2748 gnd 0.007318f
C3415 vdd.n2749 gnd 0.009093f
C3416 vdd.n2750 gnd 0.009093f
C3417 vdd.n2751 gnd 0.007318f
C3418 vdd.n2752 gnd 0.009093f
C3419 vdd.n2753 gnd 0.009093f
C3420 vdd.n2754 gnd 0.007318f
C3421 vdd.n2755 gnd 0.009093f
C3422 vdd.n2756 gnd 0.009093f
C3423 vdd.n2757 gnd 0.009093f
C3424 vdd.n2758 gnd 0.01493f
C3425 vdd.n2759 gnd 0.009093f
C3426 vdd.n2760 gnd 0.009093f
C3427 vdd.n2761 gnd 0.004977f
C3428 vdd.n2762 gnd 0.007318f
C3429 vdd.n2763 gnd 0.009093f
C3430 vdd.n2764 gnd 0.009093f
C3431 vdd.n2765 gnd 0.007318f
C3432 vdd.n2766 gnd 0.007318f
C3433 vdd.n2767 gnd 0.009093f
C3434 vdd.n2768 gnd 0.009093f
C3435 vdd.n2769 gnd 0.007318f
C3436 vdd.n2770 gnd 0.007318f
C3437 vdd.n2771 gnd 0.009093f
C3438 vdd.n2772 gnd 0.009093f
C3439 vdd.n2773 gnd 0.007318f
C3440 vdd.n2774 gnd 0.007318f
C3441 vdd.n2775 gnd 0.009093f
C3442 vdd.n2776 gnd 0.009093f
C3443 vdd.n2777 gnd 0.007318f
C3444 vdd.n2778 gnd 0.007318f
C3445 vdd.n2779 gnd 0.009093f
C3446 vdd.n2780 gnd 0.009093f
C3447 vdd.n2781 gnd 0.007318f
C3448 vdd.n2782 gnd 0.007318f
C3449 vdd.n2783 gnd 0.009093f
C3450 vdd.n2784 gnd 0.009093f
C3451 vdd.n2785 gnd 0.007318f
C3452 vdd.n2786 gnd 0.007318f
C3453 vdd.n2787 gnd 0.009093f
C3454 vdd.n2788 gnd 0.009093f
C3455 vdd.n2789 gnd 0.007318f
C3456 vdd.n2790 gnd 0.007318f
C3457 vdd.n2791 gnd 0.009093f
C3458 vdd.n2792 gnd 0.009093f
C3459 vdd.n2793 gnd 0.007318f
C3460 vdd.n2794 gnd 0.007318f
C3461 vdd.n2795 gnd 0.009093f
C3462 vdd.n2796 gnd 0.009093f
C3463 vdd.n2797 gnd 0.007318f
C3464 vdd.n2798 gnd 0.009093f
C3465 vdd.n2799 gnd 0.009093f
C3466 vdd.n2800 gnd 0.007318f
C3467 vdd.n2801 gnd 0.009093f
C3468 vdd.n2802 gnd 0.009093f
C3469 vdd.n2803 gnd 0.009093f
C3470 vdd.t129 gnd 0.111862f
C3471 vdd.t130 gnd 0.11955f
C3472 vdd.t128 gnd 0.14609f
C3473 vdd.n2804 gnd 0.187267f
C3474 vdd.n2805 gnd 0.157338f
C3475 vdd.n2806 gnd 0.01493f
C3476 vdd.n2807 gnd 0.009093f
C3477 vdd.n2808 gnd 0.009093f
C3478 vdd.n2809 gnd 0.006111f
C3479 vdd.n2810 gnd 0.007318f
C3480 vdd.n2811 gnd 0.009093f
C3481 vdd.n2812 gnd 0.009093f
C3482 vdd.n2813 gnd 0.007318f
C3483 vdd.n2814 gnd 0.007318f
C3484 vdd.n2815 gnd 0.009093f
C3485 vdd.n2816 gnd 0.009093f
C3486 vdd.n2817 gnd 0.007318f
C3487 vdd.n2818 gnd 0.007318f
C3488 vdd.n2819 gnd 0.009093f
C3489 vdd.n2820 gnd 0.009093f
C3490 vdd.n2821 gnd 0.007318f
C3491 vdd.n2822 gnd 0.007318f
C3492 vdd.n2823 gnd 0.009093f
C3493 vdd.n2824 gnd 0.009093f
C3494 vdd.n2825 gnd 0.007318f
C3495 vdd.n2826 gnd 0.007318f
C3496 vdd.n2827 gnd 0.009093f
C3497 vdd.n2828 gnd 0.009093f
C3498 vdd.n2829 gnd 0.007318f
C3499 vdd.n2830 gnd 0.007318f
C3500 vdd.n2831 gnd 0.009093f
C3501 vdd.n2832 gnd 0.009093f
C3502 vdd.n2833 gnd 0.007318f
C3503 vdd.n2834 gnd 0.007318f
C3504 vdd.n2836 gnd 0.550295f
C3505 vdd.n2838 gnd 0.007318f
C3506 vdd.n2839 gnd 0.009093f
C3507 vdd.n2840 gnd 6.7368f
C3508 vdd.n2842 gnd 0.022667f
C3509 vdd.n2843 gnd 0.006074f
C3510 vdd.n2844 gnd 0.022667f
C3511 vdd.n2845 gnd 0.022159f
C3512 vdd.n2846 gnd 0.009093f
C3513 vdd.n2847 gnd 0.007318f
C3514 vdd.n2848 gnd 0.009093f
C3515 vdd.n2849 gnd 0.580759f
C3516 vdd.n2850 gnd 0.009093f
C3517 vdd.n2851 gnd 0.007318f
C3518 vdd.n2852 gnd 0.009093f
C3519 vdd.n2853 gnd 0.009093f
C3520 vdd.n2854 gnd 0.009093f
C3521 vdd.n2855 gnd 0.007318f
C3522 vdd.n2856 gnd 0.009093f
C3523 vdd.n2857 gnd 0.738725f
C3524 vdd.n2858 gnd 0.929214f
C3525 vdd.n2859 gnd 0.009093f
C3526 vdd.n2860 gnd 0.007318f
C3527 vdd.n2861 gnd 0.009093f
C3528 vdd.n2862 gnd 0.009093f
C3529 vdd.n2863 gnd 0.009093f
C3530 vdd.n2864 gnd 0.007318f
C3531 vdd.n2865 gnd 0.009093f
C3532 vdd.n2866 gnd 0.655096f
C3533 vdd.n2867 gnd 0.009093f
C3534 vdd.n2868 gnd 0.007318f
C3535 vdd.n2869 gnd 0.009093f
C3536 vdd.n2870 gnd 0.009093f
C3537 vdd.n2871 gnd 0.009093f
C3538 vdd.n2872 gnd 0.007318f
C3539 vdd.n2873 gnd 0.009093f
C3540 vdd.t51 gnd 0.464607f
C3541 vdd.n2874 gnd 0.771248f
C3542 vdd.n2875 gnd 0.009093f
C3543 vdd.n2876 gnd 0.007318f
C3544 vdd.n2877 gnd 0.009093f
C3545 vdd.n2878 gnd 0.009093f
C3546 vdd.n2879 gnd 0.009093f
C3547 vdd.n2880 gnd 0.007318f
C3548 vdd.n2881 gnd 0.009093f
C3549 vdd.n2882 gnd 0.729433f
C3550 vdd.n2883 gnd 0.009093f
C3551 vdd.n2884 gnd 0.007318f
C3552 vdd.n2885 gnd 0.009093f
C3553 vdd.n2886 gnd 0.009093f
C3554 vdd.n2887 gnd 0.009093f
C3555 vdd.n2888 gnd 0.007318f
C3556 vdd.n2889 gnd 0.007318f
C3557 vdd.n2890 gnd 0.007318f
C3558 vdd.n2891 gnd 0.009093f
C3559 vdd.n2892 gnd 0.009093f
C3560 vdd.n2893 gnd 0.009093f
C3561 vdd.n2894 gnd 0.007318f
C3562 vdd.n2895 gnd 0.007318f
C3563 vdd.n2896 gnd 0.007318f
C3564 vdd.n2897 gnd 0.009093f
C3565 vdd.n2898 gnd 0.009093f
C3566 vdd.n2899 gnd 0.009093f
C3567 vdd.n2900 gnd 0.007318f
C3568 vdd.n2901 gnd 0.007318f
C3569 vdd.n2902 gnd 0.006074f
C3570 vdd.n2903 gnd 0.022159f
C3571 vdd.n2904 gnd 0.022667f
C3572 vdd.n2906 gnd 0.022667f
C3573 vdd.n2907 gnd 0.003476f
C3574 vdd.t196 gnd 0.111862f
C3575 vdd.t195 gnd 0.11955f
C3576 vdd.t194 gnd 0.14609f
C3577 vdd.n2908 gnd 0.187267f
C3578 vdd.n2909 gnd 0.15807f
C3579 vdd.n2910 gnd 0.012002f
C3580 vdd.n2911 gnd 0.003842f
C3581 vdd.n2912 gnd 0.007318f
C3582 vdd.n2913 gnd 0.009093f
C3583 vdd.n2915 gnd 0.009093f
C3584 vdd.n2916 gnd 0.009093f
C3585 vdd.n2917 gnd 0.007318f
C3586 vdd.n2918 gnd 0.007318f
C3587 vdd.n2919 gnd 0.007318f
C3588 vdd.n2920 gnd 0.009093f
C3589 vdd.n2922 gnd 0.009093f
C3590 vdd.n2923 gnd 0.009093f
C3591 vdd.n2924 gnd 0.007318f
C3592 vdd.n2925 gnd 0.007318f
C3593 vdd.n2926 gnd 0.007318f
C3594 vdd.n2927 gnd 0.009093f
C3595 vdd.n2929 gnd 0.009093f
C3596 vdd.n2930 gnd 0.009093f
C3597 vdd.n2931 gnd 0.007318f
C3598 vdd.n2932 gnd 0.007318f
C3599 vdd.n2933 gnd 0.007318f
C3600 vdd.n2934 gnd 0.009093f
C3601 vdd.n2936 gnd 0.009093f
C3602 vdd.n2937 gnd 0.009093f
C3603 vdd.n2938 gnd 0.007318f
C3604 vdd.n2939 gnd 0.007318f
C3605 vdd.n2940 gnd 0.007318f
C3606 vdd.n2941 gnd 0.009093f
C3607 vdd.n2943 gnd 0.009093f
C3608 vdd.n2944 gnd 0.009093f
C3609 vdd.n2945 gnd 0.007318f
C3610 vdd.n2946 gnd 0.009093f
C3611 vdd.n2947 gnd 0.009093f
C3612 vdd.n2948 gnd 0.009093f
C3613 vdd.n2949 gnd 0.015661f
C3614 vdd.n2950 gnd 0.004977f
C3615 vdd.n2951 gnd 0.007318f
C3616 vdd.n2952 gnd 0.009093f
C3617 vdd.n2954 gnd 0.009093f
C3618 vdd.n2955 gnd 0.009093f
C3619 vdd.n2956 gnd 0.007318f
C3620 vdd.n2957 gnd 0.007318f
C3621 vdd.n2958 gnd 0.007318f
C3622 vdd.n2959 gnd 0.009093f
C3623 vdd.n2961 gnd 0.009093f
C3624 vdd.n2962 gnd 0.009093f
C3625 vdd.n2963 gnd 0.007318f
C3626 vdd.n2964 gnd 0.007318f
C3627 vdd.n2965 gnd 0.007318f
C3628 vdd.n2966 gnd 0.009093f
C3629 vdd.n2968 gnd 0.009093f
C3630 vdd.n2969 gnd 0.009093f
C3631 vdd.n2970 gnd 0.007318f
C3632 vdd.n2971 gnd 0.007318f
C3633 vdd.n2972 gnd 0.007318f
C3634 vdd.n2973 gnd 0.009093f
C3635 vdd.n2975 gnd 0.009093f
C3636 vdd.n2976 gnd 0.009093f
C3637 vdd.n2977 gnd 0.007318f
C3638 vdd.n2978 gnd 0.007318f
C3639 vdd.n2979 gnd 0.007318f
C3640 vdd.n2980 gnd 0.009093f
C3641 vdd.n2982 gnd 0.009093f
C3642 vdd.n2983 gnd 0.009093f
C3643 vdd.n2984 gnd 0.007318f
C3644 vdd.n2985 gnd 0.009093f
C3645 vdd.n2986 gnd 0.009093f
C3646 vdd.n2987 gnd 0.009093f
C3647 vdd.n2988 gnd 0.015661f
C3648 vdd.n2989 gnd 0.006111f
C3649 vdd.n2990 gnd 0.007318f
C3650 vdd.n2991 gnd 0.009093f
C3651 vdd.n2993 gnd 0.009093f
C3652 vdd.n2994 gnd 0.009093f
C3653 vdd.n2995 gnd 0.007318f
C3654 vdd.n2996 gnd 0.007318f
C3655 vdd.n2997 gnd 0.007318f
C3656 vdd.n2998 gnd 0.009093f
C3657 vdd.n3000 gnd 0.009093f
C3658 vdd.n3001 gnd 0.009093f
C3659 vdd.n3002 gnd 0.007318f
C3660 vdd.n3003 gnd 0.007318f
C3661 vdd.n3004 gnd 0.007318f
C3662 vdd.n3005 gnd 0.009093f
C3663 vdd.n3007 gnd 0.009093f
C3664 vdd.n3008 gnd 0.009093f
C3665 vdd.n3009 gnd 0.007318f
C3666 vdd.n3010 gnd 0.007318f
C3667 vdd.n3011 gnd 0.007318f
C3668 vdd.n3012 gnd 0.009093f
C3669 vdd.n3014 gnd 0.009093f
C3670 vdd.n3015 gnd 0.009093f
C3671 vdd.n3017 gnd 0.009093f
C3672 vdd.n3018 gnd 0.007318f
C3673 vdd.n3019 gnd 0.007318f
C3674 vdd.n3020 gnd 0.006074f
C3675 vdd.n3021 gnd 0.022667f
C3676 vdd.n3022 gnd 0.022159f
C3677 vdd.n3023 gnd 0.006074f
C3678 vdd.n3024 gnd 0.022159f
C3679 vdd.n3025 gnd 1.37059f
C3680 vdd.t147 gnd 0.464607f
C3681 vdd.n3026 gnd 0.487837f
C3682 vdd.n3027 gnd 0.929214f
C3683 vdd.n3028 gnd 0.009093f
C3684 vdd.n3029 gnd 0.007318f
C3685 vdd.n3030 gnd 0.007318f
C3686 vdd.n3031 gnd 0.007318f
C3687 vdd.n3032 gnd 0.009093f
C3688 vdd.n3033 gnd 0.831647f
C3689 vdd.t42 gnd 0.464607f
C3690 vdd.n3034 gnd 0.562174f
C3691 vdd.n3035 gnd 0.67368f
C3692 vdd.n3036 gnd 0.009093f
C3693 vdd.n3037 gnd 0.007318f
C3694 vdd.n3038 gnd 0.007318f
C3695 vdd.n3039 gnd 0.007318f
C3696 vdd.n3040 gnd 0.009093f
C3697 vdd.n3041 gnd 0.515714f
C3698 vdd.t64 gnd 0.464607f
C3699 vdd.n3042 gnd 0.771248f
C3700 vdd.t40 gnd 0.464607f
C3701 vdd.n3043 gnd 0.571467f
C3702 vdd.n3044 gnd 0.009093f
C3703 vdd.n3045 gnd 0.007318f
C3704 vdd.n3046 gnd 0.006988f
C3705 vdd.n3047 gnd 0.536312f
C3706 vdd.n3048 gnd 1.84155f
C3707 a_n5644_8799.t15 gnd 0.111879f
C3708 a_n5644_8799.t10 gnd 0.111879f
C3709 a_n5644_8799.t9 gnd 0.111879f
C3710 a_n5644_8799.n0 gnd 0.990799f
C3711 a_n5644_8799.t30 gnd 0.143844f
C3712 a_n5644_8799.t20 gnd 0.143844f
C3713 a_n5644_8799.n1 gnd 1.13452f
C3714 a_n5644_8799.t26 gnd 0.143844f
C3715 a_n5644_8799.t27 gnd 0.143844f
C3716 a_n5644_8799.n2 gnd 1.13265f
C3717 a_n5644_8799.n3 gnd 1.01812f
C3718 a_n5644_8799.t28 gnd 0.143844f
C3719 a_n5644_8799.t21 gnd 0.143844f
C3720 a_n5644_8799.n4 gnd 1.13265f
C3721 a_n5644_8799.n5 gnd 2.94695f
C3722 a_n5644_8799.t23 gnd 0.143844f
C3723 a_n5644_8799.t25 gnd 0.143844f
C3724 a_n5644_8799.n6 gnd 1.13452f
C3725 a_n5644_8799.t29 gnd 0.143844f
C3726 a_n5644_8799.t24 gnd 0.143844f
C3727 a_n5644_8799.n7 gnd 1.13265f
C3728 a_n5644_8799.n8 gnd 1.01811f
C3729 a_n5644_8799.t31 gnd 0.143844f
C3730 a_n5644_8799.t22 gnd 0.143844f
C3731 a_n5644_8799.n9 gnd 1.13265f
C3732 a_n5644_8799.n10 gnd 1.80867f
C3733 a_n5644_8799.n11 gnd 5.67846f
C3734 a_n5644_8799.n12 gnd 0.051846f
C3735 a_n5644_8799.t71 gnd 0.596445f
C3736 a_n5644_8799.n13 gnd 0.266384f
C3737 a_n5644_8799.n14 gnd 0.051846f
C3738 a_n5644_8799.n15 gnd 0.011765f
C3739 a_n5644_8799.t38 gnd 0.596445f
C3740 a_n5644_8799.n16 gnd 0.16507f
C3741 a_n5644_8799.t58 gnd 0.596445f
C3742 a_n5644_8799.t49 gnd 0.607734f
C3743 a_n5644_8799.n17 gnd 0.250039f
C3744 a_n5644_8799.n18 gnd 0.263347f
C3745 a_n5644_8799.n19 gnd 0.011765f
C3746 a_n5644_8799.t73 gnd 0.596445f
C3747 a_n5644_8799.n20 gnd 0.266384f
C3748 a_n5644_8799.n21 gnd 0.051846f
C3749 a_n5644_8799.n22 gnd 0.051846f
C3750 a_n5644_8799.n23 gnd 0.051846f
C3751 a_n5644_8799.n24 gnd 0.263667f
C3752 a_n5644_8799.t48 gnd 0.596445f
C3753 a_n5644_8799.n25 gnd 0.263667f
C3754 a_n5644_8799.n26 gnd 0.011765f
C3755 a_n5644_8799.n27 gnd 0.051846f
C3756 a_n5644_8799.n28 gnd 0.051846f
C3757 a_n5644_8799.n29 gnd 0.051846f
C3758 a_n5644_8799.n30 gnd 0.011765f
C3759 a_n5644_8799.t37 gnd 0.596445f
C3760 a_n5644_8799.n31 gnd 0.263347f
C3761 a_n5644_8799.t36 gnd 0.596445f
C3762 a_n5644_8799.n32 gnd 0.26095f
C3763 a_n5644_8799.n33 gnd 0.295016f
C3764 a_n5644_8799.n34 gnd 0.051846f
C3765 a_n5644_8799.t75 gnd 0.596445f
C3766 a_n5644_8799.n35 gnd 0.266384f
C3767 a_n5644_8799.n36 gnd 0.051846f
C3768 a_n5644_8799.n37 gnd 0.011765f
C3769 a_n5644_8799.t45 gnd 0.596445f
C3770 a_n5644_8799.n38 gnd 0.16507f
C3771 a_n5644_8799.t64 gnd 0.596445f
C3772 a_n5644_8799.t54 gnd 0.607734f
C3773 a_n5644_8799.n39 gnd 0.250039f
C3774 a_n5644_8799.n40 gnd 0.263347f
C3775 a_n5644_8799.n41 gnd 0.011765f
C3776 a_n5644_8799.t77 gnd 0.596445f
C3777 a_n5644_8799.n42 gnd 0.266384f
C3778 a_n5644_8799.n43 gnd 0.051846f
C3779 a_n5644_8799.n44 gnd 0.051846f
C3780 a_n5644_8799.n45 gnd 0.051846f
C3781 a_n5644_8799.n46 gnd 0.263667f
C3782 a_n5644_8799.t53 gnd 0.596445f
C3783 a_n5644_8799.n47 gnd 0.263667f
C3784 a_n5644_8799.n48 gnd 0.011765f
C3785 a_n5644_8799.n49 gnd 0.051846f
C3786 a_n5644_8799.n50 gnd 0.051846f
C3787 a_n5644_8799.n51 gnd 0.051846f
C3788 a_n5644_8799.n52 gnd 0.011765f
C3789 a_n5644_8799.t41 gnd 0.596445f
C3790 a_n5644_8799.n53 gnd 0.263347f
C3791 a_n5644_8799.t43 gnd 0.596445f
C3792 a_n5644_8799.n54 gnd 0.26095f
C3793 a_n5644_8799.n55 gnd 0.130362f
C3794 a_n5644_8799.n56 gnd 0.897033f
C3795 a_n5644_8799.n57 gnd 0.051846f
C3796 a_n5644_8799.t62 gnd 0.596445f
C3797 a_n5644_8799.n58 gnd 0.266384f
C3798 a_n5644_8799.n59 gnd 0.051846f
C3799 a_n5644_8799.n60 gnd 0.011765f
C3800 a_n5644_8799.t70 gnd 0.596445f
C3801 a_n5644_8799.n61 gnd 0.16507f
C3802 a_n5644_8799.t67 gnd 0.596445f
C3803 a_n5644_8799.t35 gnd 0.607734f
C3804 a_n5644_8799.n62 gnd 0.250039f
C3805 a_n5644_8799.n63 gnd 0.263347f
C3806 a_n5644_8799.n64 gnd 0.011765f
C3807 a_n5644_8799.t44 gnd 0.596445f
C3808 a_n5644_8799.n65 gnd 0.266384f
C3809 a_n5644_8799.n66 gnd 0.051846f
C3810 a_n5644_8799.n67 gnd 0.051846f
C3811 a_n5644_8799.n68 gnd 0.051846f
C3812 a_n5644_8799.n69 gnd 0.263667f
C3813 a_n5644_8799.t50 gnd 0.596445f
C3814 a_n5644_8799.n70 gnd 0.263667f
C3815 a_n5644_8799.n71 gnd 0.011765f
C3816 a_n5644_8799.n72 gnd 0.051846f
C3817 a_n5644_8799.n73 gnd 0.051846f
C3818 a_n5644_8799.n74 gnd 0.051846f
C3819 a_n5644_8799.n75 gnd 0.011765f
C3820 a_n5644_8799.t39 gnd 0.596445f
C3821 a_n5644_8799.n76 gnd 0.263347f
C3822 a_n5644_8799.t79 gnd 0.596445f
C3823 a_n5644_8799.n77 gnd 0.26095f
C3824 a_n5644_8799.n78 gnd 0.130362f
C3825 a_n5644_8799.n79 gnd 1.4561f
C3826 a_n5644_8799.n80 gnd 0.051846f
C3827 a_n5644_8799.t56 gnd 0.596445f
C3828 a_n5644_8799.t55 gnd 0.596445f
C3829 a_n5644_8799.t42 gnd 0.596445f
C3830 a_n5644_8799.n81 gnd 0.266384f
C3831 a_n5644_8799.n82 gnd 0.051846f
C3832 a_n5644_8799.t72 gnd 0.596445f
C3833 a_n5644_8799.t57 gnd 0.596445f
C3834 a_n5644_8799.n83 gnd 0.051846f
C3835 a_n5644_8799.t47 gnd 0.596445f
C3836 a_n5644_8799.n84 gnd 0.266384f
C3837 a_n5644_8799.t65 gnd 0.607734f
C3838 a_n5644_8799.n85 gnd 0.250039f
C3839 a_n5644_8799.t74 gnd 0.596445f
C3840 a_n5644_8799.n86 gnd 0.263347f
C3841 a_n5644_8799.n87 gnd 0.011765f
C3842 a_n5644_8799.n88 gnd 0.16507f
C3843 a_n5644_8799.n89 gnd 0.051846f
C3844 a_n5644_8799.n90 gnd 0.051846f
C3845 a_n5644_8799.n91 gnd 0.011765f
C3846 a_n5644_8799.n92 gnd 0.263667f
C3847 a_n5644_8799.n93 gnd 0.263667f
C3848 a_n5644_8799.n94 gnd 0.011765f
C3849 a_n5644_8799.n95 gnd 0.051846f
C3850 a_n5644_8799.n96 gnd 0.051846f
C3851 a_n5644_8799.n97 gnd 0.051846f
C3852 a_n5644_8799.n98 gnd 0.011765f
C3853 a_n5644_8799.n99 gnd 0.263347f
C3854 a_n5644_8799.n100 gnd 0.26095f
C3855 a_n5644_8799.n101 gnd 0.295016f
C3856 a_n5644_8799.n102 gnd 0.051846f
C3857 a_n5644_8799.t60 gnd 0.596445f
C3858 a_n5644_8799.t59 gnd 0.596445f
C3859 a_n5644_8799.t51 gnd 0.596445f
C3860 a_n5644_8799.n103 gnd 0.266384f
C3861 a_n5644_8799.n104 gnd 0.051846f
C3862 a_n5644_8799.t76 gnd 0.596445f
C3863 a_n5644_8799.t63 gnd 0.596445f
C3864 a_n5644_8799.n105 gnd 0.051846f
C3865 a_n5644_8799.t52 gnd 0.596445f
C3866 a_n5644_8799.n106 gnd 0.266384f
C3867 a_n5644_8799.t68 gnd 0.607734f
C3868 a_n5644_8799.n107 gnd 0.250039f
C3869 a_n5644_8799.t32 gnd 0.596445f
C3870 a_n5644_8799.n108 gnd 0.263347f
C3871 a_n5644_8799.n109 gnd 0.011765f
C3872 a_n5644_8799.n110 gnd 0.16507f
C3873 a_n5644_8799.n111 gnd 0.051846f
C3874 a_n5644_8799.n112 gnd 0.051846f
C3875 a_n5644_8799.n113 gnd 0.011765f
C3876 a_n5644_8799.n114 gnd 0.263667f
C3877 a_n5644_8799.n115 gnd 0.263667f
C3878 a_n5644_8799.n116 gnd 0.011765f
C3879 a_n5644_8799.n117 gnd 0.051846f
C3880 a_n5644_8799.n118 gnd 0.051846f
C3881 a_n5644_8799.n119 gnd 0.051846f
C3882 a_n5644_8799.n120 gnd 0.011765f
C3883 a_n5644_8799.n121 gnd 0.263347f
C3884 a_n5644_8799.n122 gnd 0.26095f
C3885 a_n5644_8799.n123 gnd 0.130362f
C3886 a_n5644_8799.n124 gnd 0.897033f
C3887 a_n5644_8799.n125 gnd 0.051846f
C3888 a_n5644_8799.t78 gnd 0.596445f
C3889 a_n5644_8799.t40 gnd 0.596445f
C3890 a_n5644_8799.t61 gnd 0.596445f
C3891 a_n5644_8799.n126 gnd 0.266384f
C3892 a_n5644_8799.n127 gnd 0.051846f
C3893 a_n5644_8799.t33 gnd 0.596445f
C3894 a_n5644_8799.t69 gnd 0.596445f
C3895 a_n5644_8799.n128 gnd 0.051846f
C3896 a_n5644_8799.t46 gnd 0.596445f
C3897 a_n5644_8799.n129 gnd 0.266384f
C3898 a_n5644_8799.t34 gnd 0.607734f
C3899 a_n5644_8799.n130 gnd 0.250039f
C3900 a_n5644_8799.t66 gnd 0.596445f
C3901 a_n5644_8799.n131 gnd 0.263347f
C3902 a_n5644_8799.n132 gnd 0.011765f
C3903 a_n5644_8799.n133 gnd 0.16507f
C3904 a_n5644_8799.n134 gnd 0.051846f
C3905 a_n5644_8799.n135 gnd 0.051846f
C3906 a_n5644_8799.n136 gnd 0.011765f
C3907 a_n5644_8799.n137 gnd 0.263667f
C3908 a_n5644_8799.n138 gnd 0.263667f
C3909 a_n5644_8799.n139 gnd 0.011765f
C3910 a_n5644_8799.n140 gnd 0.051846f
C3911 a_n5644_8799.n141 gnd 0.051846f
C3912 a_n5644_8799.n142 gnd 0.051846f
C3913 a_n5644_8799.n143 gnd 0.011765f
C3914 a_n5644_8799.n144 gnd 0.263347f
C3915 a_n5644_8799.n145 gnd 0.26095f
C3916 a_n5644_8799.n146 gnd 0.130362f
C3917 a_n5644_8799.n147 gnd 1.13032f
C3918 a_n5644_8799.n148 gnd 12.2154f
C3919 a_n5644_8799.n149 gnd 4.36511f
C3920 a_n5644_8799.t6 gnd 0.111879f
C3921 a_n5644_8799.t7 gnd 0.111879f
C3922 a_n5644_8799.n150 gnd 0.990799f
C3923 a_n5644_8799.t2 gnd 0.111879f
C3924 a_n5644_8799.t3 gnd 0.111879f
C3925 a_n5644_8799.n151 gnd 0.988601f
C3926 a_n5644_8799.n152 gnd 0.787466f
C3927 a_n5644_8799.t1 gnd 0.111879f
C3928 a_n5644_8799.t16 gnd 0.111879f
C3929 a_n5644_8799.n153 gnd 0.988601f
C3930 a_n5644_8799.n154 gnd 0.740399f
C3931 a_n5644_8799.t17 gnd 0.111879f
C3932 a_n5644_8799.t12 gnd 0.111879f
C3933 a_n5644_8799.n155 gnd 0.988601f
C3934 a_n5644_8799.n156 gnd 0.386686f
C3935 a_n5644_8799.t14 gnd 0.111879f
C3936 a_n5644_8799.t0 gnd 0.111879f
C3937 a_n5644_8799.n157 gnd 0.988601f
C3938 a_n5644_8799.n158 gnd 2.70455f
C3939 a_n5644_8799.t13 gnd 0.111879f
C3940 a_n5644_8799.t11 gnd 0.111879f
C3941 a_n5644_8799.n159 gnd 0.990799f
C3942 a_n5644_8799.t4 gnd 0.111879f
C3943 a_n5644_8799.t8 gnd 0.111879f
C3944 a_n5644_8799.n160 gnd 0.9886f
C3945 a_n5644_8799.n161 gnd 0.787468f
C3946 a_n5644_8799.t18 gnd 0.111879f
C3947 a_n5644_8799.t5 gnd 0.111879f
C3948 a_n5644_8799.n162 gnd 0.9886f
C3949 a_n5644_8799.n163 gnd 2.46205f
C3950 a_n5644_8799.n164 gnd 0.78747f
C3951 a_n5644_8799.n165 gnd 0.988597f
C3952 a_n5644_8799.t19 gnd 0.111879f
C3953 a_n2903_n3924.n0 gnd 0.954594f
C3954 a_n2903_n3924.n1 gnd 1.81294f
C3955 a_n2903_n3924.n2 gnd 0.724068f
C3956 a_n2903_n3924.n3 gnd 1.31663f
C3957 a_n2903_n3924.n4 gnd 1.27336f
C3958 a_n2903_n3924.n5 gnd 1.81293f
C3959 a_n2903_n3924.n6 gnd 0.724066f
C3960 a_n2903_n3924.n7 gnd 1.63539f
C3961 a_n2903_n3924.n8 gnd 1.60399f
C3962 a_n2903_n3924.n9 gnd 1.7731f
C3963 a_n2903_n3924.n10 gnd 1.7731f
C3964 a_n2903_n3924.n11 gnd 2.13362f
C3965 a_n2903_n3924.t14 gnd 1.01309f
C3966 a_n2903_n3924.t10 gnd 1.01309f
C3967 a_n2903_n3924.t1 gnd 0.097476f
C3968 a_n2903_n3924.t12 gnd 0.097476f
C3969 a_n2903_n3924.n12 gnd 0.796106f
C3970 a_n2903_n3924.t7 gnd 0.097476f
C3971 a_n2903_n3924.t11 gnd 0.097476f
C3972 a_n2903_n3924.n13 gnd 0.796106f
C3973 a_n2903_n3924.t19 gnd 0.097476f
C3974 a_n2903_n3924.t6 gnd 0.097476f
C3975 a_n2903_n3924.n14 gnd 0.796106f
C3976 a_n2903_n3924.t2 gnd 0.097476f
C3977 a_n2903_n3924.t15 gnd 0.097476f
C3978 a_n2903_n3924.n15 gnd 0.796106f
C3979 a_n2903_n3924.t4 gnd 1.01309f
C3980 a_n2903_n3924.t21 gnd 1.01309f
C3981 a_n2903_n3924.t40 gnd 0.097476f
C3982 a_n2903_n3924.t31 gnd 0.097476f
C3983 a_n2903_n3924.n16 gnd 0.796106f
C3984 a_n2903_n3924.t33 gnd 0.097476f
C3985 a_n2903_n3924.t35 gnd 0.097476f
C3986 a_n2903_n3924.n17 gnd 0.796106f
C3987 a_n2903_n3924.t34 gnd 0.097476f
C3988 a_n2903_n3924.t20 gnd 0.097476f
C3989 a_n2903_n3924.n18 gnd 0.796106f
C3990 a_n2903_n3924.t32 gnd 0.097476f
C3991 a_n2903_n3924.t45 gnd 0.097476f
C3992 a_n2903_n3924.n19 gnd 0.796106f
C3993 a_n2903_n3924.t25 gnd 1.01309f
C3994 a_n2903_n3924.n20 gnd 0.914361f
C3995 a_n2903_n3924.t43 gnd 1.26033f
C3996 a_n2903_n3924.t42 gnd 1.25874f
C3997 a_n2903_n3924.t41 gnd 1.25874f
C3998 a_n2903_n3924.t22 gnd 1.25874f
C3999 a_n2903_n3924.t23 gnd 1.25874f
C4000 a_n2903_n3924.t24 gnd 1.25874f
C4001 a_n2903_n3924.t47 gnd 1.25874f
C4002 a_n2903_n3924.t46 gnd 1.25909f
C4003 a_n2903_n3924.n21 gnd 0.914361f
C4004 a_n2903_n3924.t37 gnd 1.01309f
C4005 a_n2903_n3924.t44 gnd 0.097476f
C4006 a_n2903_n3924.t36 gnd 0.097476f
C4007 a_n2903_n3924.n22 gnd 0.796105f
C4008 a_n2903_n3924.t29 gnd 0.097476f
C4009 a_n2903_n3924.t30 gnd 0.097476f
C4010 a_n2903_n3924.n23 gnd 0.796105f
C4011 a_n2903_n3924.t27 gnd 0.097476f
C4012 a_n2903_n3924.t38 gnd 0.097476f
C4013 a_n2903_n3924.n24 gnd 0.796105f
C4014 a_n2903_n3924.t39 gnd 0.097476f
C4015 a_n2903_n3924.t26 gnd 0.097476f
C4016 a_n2903_n3924.n25 gnd 0.796105f
C4017 a_n2903_n3924.t28 gnd 1.01309f
C4018 a_n2903_n3924.t9 gnd 1.01309f
C4019 a_n2903_n3924.t8 gnd 0.097476f
C4020 a_n2903_n3924.t5 gnd 0.097476f
C4021 a_n2903_n3924.n26 gnd 0.796105f
C4022 a_n2903_n3924.t18 gnd 0.097476f
C4023 a_n2903_n3924.t13 gnd 0.097476f
C4024 a_n2903_n3924.n27 gnd 0.796105f
C4025 a_n2903_n3924.t17 gnd 0.097476f
C4026 a_n2903_n3924.t16 gnd 0.097476f
C4027 a_n2903_n3924.n28 gnd 0.796105f
C4028 a_n2903_n3924.t3 gnd 0.097476f
C4029 a_n2903_n3924.n29 gnd 0.796102f
C4030 a_n2903_n3924.t0 gnd 0.097476f
C4031 plus.n0 gnd 0.023626f
C4032 plus.t14 gnd 0.334167f
C4033 plus.n1 gnd 0.023626f
C4034 plus.t15 gnd 0.334167f
C4035 plus.t9 gnd 0.334167f
C4036 plus.n2 gnd 0.148448f
C4037 plus.n3 gnd 0.023626f
C4038 plus.t5 gnd 0.334167f
C4039 plus.t6 gnd 0.334167f
C4040 plus.n4 gnd 0.148448f
C4041 plus.n5 gnd 0.023626f
C4042 plus.t19 gnd 0.334167f
C4043 plus.t20 gnd 0.334167f
C4044 plus.n6 gnd 0.148448f
C4045 plus.n7 gnd 0.023626f
C4046 plus.t16 gnd 0.334167f
C4047 plus.t11 gnd 0.334167f
C4048 plus.n8 gnd 0.152399f
C4049 plus.t13 gnd 0.345875f
C4050 plus.n9 gnd 0.138437f
C4051 plus.n10 gnd 0.100845f
C4052 plus.n11 gnd 0.005361f
C4053 plus.n12 gnd 0.148448f
C4054 plus.n13 gnd 0.005361f
C4055 plus.n14 gnd 0.023626f
C4056 plus.n15 gnd 0.023626f
C4057 plus.n16 gnd 0.023626f
C4058 plus.n17 gnd 0.005361f
C4059 plus.n18 gnd 0.148448f
C4060 plus.n19 gnd 0.005361f
C4061 plus.n20 gnd 0.023626f
C4062 plus.n21 gnd 0.023626f
C4063 plus.n22 gnd 0.023626f
C4064 plus.n23 gnd 0.005361f
C4065 plus.n24 gnd 0.148448f
C4066 plus.n25 gnd 0.005361f
C4067 plus.n26 gnd 0.023626f
C4068 plus.n27 gnd 0.023626f
C4069 plus.n28 gnd 0.023626f
C4070 plus.n29 gnd 0.005361f
C4071 plus.n30 gnd 0.148448f
C4072 plus.n31 gnd 0.005361f
C4073 plus.n32 gnd 0.148229f
C4074 plus.n33 gnd 0.266893f
C4075 plus.n34 gnd 0.023626f
C4076 plus.n35 gnd 0.005361f
C4077 plus.t10 gnd 0.334167f
C4078 plus.n36 gnd 0.023626f
C4079 plus.n37 gnd 0.005361f
C4080 plus.t7 gnd 0.334167f
C4081 plus.n38 gnd 0.023626f
C4082 plus.n39 gnd 0.005361f
C4083 plus.t23 gnd 0.334167f
C4084 plus.n40 gnd 0.023626f
C4085 plus.n41 gnd 0.005361f
C4086 plus.t22 gnd 0.334167f
C4087 plus.t18 gnd 0.345875f
C4088 plus.t17 gnd 0.334167f
C4089 plus.n42 gnd 0.152399f
C4090 plus.n43 gnd 0.138437f
C4091 plus.n44 gnd 0.100845f
C4092 plus.n45 gnd 0.023626f
C4093 plus.n46 gnd 0.148448f
C4094 plus.n47 gnd 0.005361f
C4095 plus.t21 gnd 0.334167f
C4096 plus.n48 gnd 0.148448f
C4097 plus.n49 gnd 0.023626f
C4098 plus.n50 gnd 0.023626f
C4099 plus.n51 gnd 0.023626f
C4100 plus.n52 gnd 0.148448f
C4101 plus.n53 gnd 0.005361f
C4102 plus.t8 gnd 0.334167f
C4103 plus.n54 gnd 0.148448f
C4104 plus.n55 gnd 0.023626f
C4105 plus.n56 gnd 0.023626f
C4106 plus.n57 gnd 0.023626f
C4107 plus.n58 gnd 0.148448f
C4108 plus.n59 gnd 0.005361f
C4109 plus.t12 gnd 0.334167f
C4110 plus.n60 gnd 0.148448f
C4111 plus.n61 gnd 0.023626f
C4112 plus.n62 gnd 0.023626f
C4113 plus.n63 gnd 0.023626f
C4114 plus.n64 gnd 0.148448f
C4115 plus.n65 gnd 0.005361f
C4116 plus.t24 gnd 0.334167f
C4117 plus.n66 gnd 0.148229f
C4118 plus.n67 gnd 0.728767f
C4119 plus.n68 gnd 1.10207f
C4120 plus.t0 gnd 0.040785f
C4121 plus.t4 gnd 0.007283f
C4122 plus.t2 gnd 0.007283f
C4123 plus.n69 gnd 0.023621f
C4124 plus.n70 gnd 0.183369f
C4125 plus.t1 gnd 0.007283f
C4126 plus.t3 gnd 0.007283f
C4127 plus.n71 gnd 0.023621f
C4128 plus.n72 gnd 0.137641f
C4129 plus.n73 gnd 2.4365f
C4130 CSoutput.n0 gnd 0.037257f
C4131 CSoutput.t121 gnd 0.246449f
C4132 CSoutput.n1 gnd 0.111284f
C4133 CSoutput.n2 gnd 0.037257f
C4134 CSoutput.t125 gnd 0.246449f
C4135 CSoutput.n3 gnd 0.029529f
C4136 CSoutput.n4 gnd 0.037257f
C4137 CSoutput.t137 gnd 0.246449f
C4138 CSoutput.n5 gnd 0.025463f
C4139 CSoutput.n6 gnd 0.037257f
C4140 CSoutput.t123 gnd 0.246449f
C4141 CSoutput.t129 gnd 0.246449f
C4142 CSoutput.n7 gnd 0.110071f
C4143 CSoutput.n8 gnd 0.037257f
C4144 CSoutput.t128 gnd 0.246449f
C4145 CSoutput.n9 gnd 0.024278f
C4146 CSoutput.n10 gnd 0.037257f
C4147 CSoutput.t139 gnd 0.246449f
C4148 CSoutput.t126 gnd 0.246449f
C4149 CSoutput.n11 gnd 0.110071f
C4150 CSoutput.n12 gnd 0.037257f
C4151 CSoutput.t124 gnd 0.246449f
C4152 CSoutput.n13 gnd 0.025463f
C4153 CSoutput.n14 gnd 0.037257f
C4154 CSoutput.t138 gnd 0.246449f
C4155 CSoutput.t141 gnd 0.246449f
C4156 CSoutput.n15 gnd 0.110071f
C4157 CSoutput.n16 gnd 0.037257f
C4158 CSoutput.t122 gnd 0.246449f
C4159 CSoutput.n17 gnd 0.027196f
C4160 CSoutput.t133 gnd 0.294513f
C4161 CSoutput.t135 gnd 0.246449f
C4162 CSoutput.n18 gnd 0.140518f
C4163 CSoutput.n19 gnd 0.136351f
C4164 CSoutput.n20 gnd 0.158184f
C4165 CSoutput.n21 gnd 0.037257f
C4166 CSoutput.n22 gnd 0.031095f
C4167 CSoutput.n23 gnd 0.110071f
C4168 CSoutput.n24 gnd 0.029975f
C4169 CSoutput.n25 gnd 0.029529f
C4170 CSoutput.n26 gnd 0.037257f
C4171 CSoutput.n27 gnd 0.037257f
C4172 CSoutput.n28 gnd 0.030856f
C4173 CSoutput.n29 gnd 0.026198f
C4174 CSoutput.n30 gnd 0.112521f
C4175 CSoutput.n31 gnd 0.026559f
C4176 CSoutput.n32 gnd 0.037257f
C4177 CSoutput.n33 gnd 0.037257f
C4178 CSoutput.n34 gnd 0.037257f
C4179 CSoutput.n35 gnd 0.030528f
C4180 CSoutput.n36 gnd 0.110071f
C4181 CSoutput.n37 gnd 0.029195f
C4182 CSoutput.n38 gnd 0.030309f
C4183 CSoutput.n39 gnd 0.037257f
C4184 CSoutput.n40 gnd 0.037257f
C4185 CSoutput.n41 gnd 0.031089f
C4186 CSoutput.n42 gnd 0.028416f
C4187 CSoutput.n43 gnd 0.110071f
C4188 CSoutput.n44 gnd 0.029136f
C4189 CSoutput.n45 gnd 0.037257f
C4190 CSoutput.n46 gnd 0.037257f
C4191 CSoutput.n47 gnd 0.037257f
C4192 CSoutput.n48 gnd 0.029136f
C4193 CSoutput.n49 gnd 0.110071f
C4194 CSoutput.n50 gnd 0.028416f
C4195 CSoutput.n51 gnd 0.031089f
C4196 CSoutput.n52 gnd 0.037257f
C4197 CSoutput.n53 gnd 0.037257f
C4198 CSoutput.n54 gnd 0.030309f
C4199 CSoutput.n55 gnd 0.029195f
C4200 CSoutput.n56 gnd 0.110071f
C4201 CSoutput.n57 gnd 0.030528f
C4202 CSoutput.n58 gnd 0.037257f
C4203 CSoutput.n59 gnd 0.037257f
C4204 CSoutput.n60 gnd 0.037257f
C4205 CSoutput.n61 gnd 0.026559f
C4206 CSoutput.n62 gnd 0.112521f
C4207 CSoutput.n63 gnd 0.026198f
C4208 CSoutput.t132 gnd 0.246449f
C4209 CSoutput.n64 gnd 0.110071f
C4210 CSoutput.n65 gnd 0.030856f
C4211 CSoutput.n66 gnd 0.037257f
C4212 CSoutput.n67 gnd 0.037257f
C4213 CSoutput.n68 gnd 0.037257f
C4214 CSoutput.n69 gnd 0.029975f
C4215 CSoutput.n70 gnd 0.110071f
C4216 CSoutput.n71 gnd 0.031095f
C4217 CSoutput.n72 gnd 0.027196f
C4218 CSoutput.n73 gnd 0.037257f
C4219 CSoutput.n74 gnd 0.037257f
C4220 CSoutput.n75 gnd 0.028205f
C4221 CSoutput.n76 gnd 0.016751f
C4222 CSoutput.t134 gnd 0.276903f
C4223 CSoutput.n77 gnd 0.137554f
C4224 CSoutput.n78 gnd 0.562728f
C4225 CSoutput.t111 gnd 0.046473f
C4226 CSoutput.t9 gnd 0.046473f
C4227 CSoutput.n79 gnd 0.359811f
C4228 CSoutput.t36 gnd 0.046473f
C4229 CSoutput.t32 gnd 0.046473f
C4230 CSoutput.n80 gnd 0.35917f
C4231 CSoutput.n81 gnd 0.364557f
C4232 CSoutput.t3 gnd 0.046473f
C4233 CSoutput.t117 gnd 0.046473f
C4234 CSoutput.n82 gnd 0.35917f
C4235 CSoutput.n83 gnd 0.179638f
C4236 CSoutput.t21 gnd 0.046473f
C4237 CSoutput.t7 gnd 0.046473f
C4238 CSoutput.n84 gnd 0.35917f
C4239 CSoutput.n85 gnd 0.329415f
C4240 CSoutput.t12 gnd 0.046473f
C4241 CSoutput.t27 gnd 0.046473f
C4242 CSoutput.n86 gnd 0.359811f
C4243 CSoutput.t16 gnd 0.046473f
C4244 CSoutput.t118 gnd 0.046473f
C4245 CSoutput.n87 gnd 0.35917f
C4246 CSoutput.n88 gnd 0.364557f
C4247 CSoutput.t113 gnd 0.046473f
C4248 CSoutput.t22 gnd 0.046473f
C4249 CSoutput.n89 gnd 0.35917f
C4250 CSoutput.n90 gnd 0.179638f
C4251 CSoutput.t0 gnd 0.046473f
C4252 CSoutput.t116 gnd 0.046473f
C4253 CSoutput.n91 gnd 0.35917f
C4254 CSoutput.n92 gnd 0.267886f
C4255 CSoutput.n93 gnd 0.337802f
C4256 CSoutput.t10 gnd 0.046473f
C4257 CSoutput.t13 gnd 0.046473f
C4258 CSoutput.n94 gnd 0.359811f
C4259 CSoutput.t15 gnd 0.046473f
C4260 CSoutput.t112 gnd 0.046473f
C4261 CSoutput.n95 gnd 0.35917f
C4262 CSoutput.n96 gnd 0.364557f
C4263 CSoutput.t34 gnd 0.046473f
C4264 CSoutput.t119 gnd 0.046473f
C4265 CSoutput.n97 gnd 0.35917f
C4266 CSoutput.n98 gnd 0.179638f
C4267 CSoutput.t19 gnd 0.046473f
C4268 CSoutput.t20 gnd 0.046473f
C4269 CSoutput.n99 gnd 0.35917f
C4270 CSoutput.n100 gnd 0.267886f
C4271 CSoutput.n101 gnd 0.377576f
C4272 CSoutput.n102 gnd 6.34822f
C4273 CSoutput.n104 gnd 0.659075f
C4274 CSoutput.n105 gnd 0.494306f
C4275 CSoutput.n106 gnd 0.659075f
C4276 CSoutput.n107 gnd 0.659075f
C4277 CSoutput.n108 gnd 1.77443f
C4278 CSoutput.n109 gnd 0.659075f
C4279 CSoutput.n110 gnd 0.659075f
C4280 CSoutput.t140 gnd 0.823844f
C4281 CSoutput.n111 gnd 0.659075f
C4282 CSoutput.n112 gnd 0.659075f
C4283 CSoutput.n116 gnd 0.659075f
C4284 CSoutput.n120 gnd 0.659075f
C4285 CSoutput.n121 gnd 0.659075f
C4286 CSoutput.n123 gnd 0.659075f
C4287 CSoutput.n128 gnd 0.659075f
C4288 CSoutput.n130 gnd 0.659075f
C4289 CSoutput.n131 gnd 0.659075f
C4290 CSoutput.n133 gnd 0.659075f
C4291 CSoutput.n134 gnd 0.659075f
C4292 CSoutput.n136 gnd 0.659075f
C4293 CSoutput.t130 gnd 11.0131f
C4294 CSoutput.n138 gnd 0.659075f
C4295 CSoutput.n139 gnd 0.494306f
C4296 CSoutput.n140 gnd 0.659075f
C4297 CSoutput.n141 gnd 0.659075f
C4298 CSoutput.n142 gnd 1.77443f
C4299 CSoutput.n143 gnd 0.659075f
C4300 CSoutput.n144 gnd 0.659075f
C4301 CSoutput.t127 gnd 0.823844f
C4302 CSoutput.n145 gnd 0.659075f
C4303 CSoutput.n146 gnd 0.659075f
C4304 CSoutput.n150 gnd 0.659075f
C4305 CSoutput.n154 gnd 0.659075f
C4306 CSoutput.n155 gnd 0.659075f
C4307 CSoutput.n157 gnd 0.659075f
C4308 CSoutput.n162 gnd 0.659075f
C4309 CSoutput.n164 gnd 0.659075f
C4310 CSoutput.n165 gnd 0.659075f
C4311 CSoutput.n167 gnd 0.659075f
C4312 CSoutput.n168 gnd 0.659075f
C4313 CSoutput.n170 gnd 0.659075f
C4314 CSoutput.n171 gnd 0.494306f
C4315 CSoutput.n173 gnd 0.659075f
C4316 CSoutput.n174 gnd 0.494306f
C4317 CSoutput.n175 gnd 0.659075f
C4318 CSoutput.n176 gnd 0.659075f
C4319 CSoutput.n177 gnd 1.77443f
C4320 CSoutput.n178 gnd 0.659075f
C4321 CSoutput.n179 gnd 0.659075f
C4322 CSoutput.t120 gnd 0.823844f
C4323 CSoutput.n180 gnd 0.659075f
C4324 CSoutput.n181 gnd 1.77443f
C4325 CSoutput.n183 gnd 0.659075f
C4326 CSoutput.n184 gnd 0.659075f
C4327 CSoutput.n186 gnd 0.659075f
C4328 CSoutput.n187 gnd 0.659075f
C4329 CSoutput.t131 gnd 10.8336f
C4330 CSoutput.t136 gnd 11.0131f
C4331 CSoutput.n193 gnd 2.06762f
C4332 CSoutput.n194 gnd 8.42271f
C4333 CSoutput.n195 gnd 8.775161f
C4334 CSoutput.n200 gnd 2.23978f
C4335 CSoutput.n206 gnd 0.659075f
C4336 CSoutput.n208 gnd 0.659075f
C4337 CSoutput.n210 gnd 0.659075f
C4338 CSoutput.n212 gnd 0.659075f
C4339 CSoutput.n214 gnd 0.659075f
C4340 CSoutput.n220 gnd 0.659075f
C4341 CSoutput.n227 gnd 1.20915f
C4342 CSoutput.n228 gnd 1.20915f
C4343 CSoutput.n229 gnd 0.659075f
C4344 CSoutput.n230 gnd 0.659075f
C4345 CSoutput.n232 gnd 0.494306f
C4346 CSoutput.n233 gnd 0.423329f
C4347 CSoutput.n235 gnd 0.494306f
C4348 CSoutput.n236 gnd 0.423329f
C4349 CSoutput.n237 gnd 0.494306f
C4350 CSoutput.n239 gnd 0.659075f
C4351 CSoutput.n241 gnd 1.77443f
C4352 CSoutput.n242 gnd 2.06762f
C4353 CSoutput.n243 gnd 7.74673f
C4354 CSoutput.n245 gnd 0.494306f
C4355 CSoutput.n246 gnd 1.27188f
C4356 CSoutput.n247 gnd 0.494306f
C4357 CSoutput.n249 gnd 0.659075f
C4358 CSoutput.n251 gnd 1.77443f
C4359 CSoutput.n252 gnd 3.865f
C4360 CSoutput.t26 gnd 0.046473f
C4361 CSoutput.t1 gnd 0.046473f
C4362 CSoutput.n253 gnd 0.359811f
C4363 CSoutput.t23 gnd 0.046473f
C4364 CSoutput.t24 gnd 0.046473f
C4365 CSoutput.n254 gnd 0.35917f
C4366 CSoutput.n255 gnd 0.364557f
C4367 CSoutput.t18 gnd 0.046473f
C4368 CSoutput.t28 gnd 0.046473f
C4369 CSoutput.n256 gnd 0.35917f
C4370 CSoutput.n257 gnd 0.179638f
C4371 CSoutput.t14 gnd 0.046473f
C4372 CSoutput.t2 gnd 0.046473f
C4373 CSoutput.n258 gnd 0.35917f
C4374 CSoutput.n259 gnd 0.329415f
C4375 CSoutput.t35 gnd 0.046473f
C4376 CSoutput.t109 gnd 0.046473f
C4377 CSoutput.n260 gnd 0.359811f
C4378 CSoutput.t4 gnd 0.046473f
C4379 CSoutput.t5 gnd 0.046473f
C4380 CSoutput.n261 gnd 0.35917f
C4381 CSoutput.n262 gnd 0.364557f
C4382 CSoutput.t30 gnd 0.046473f
C4383 CSoutput.t11 gnd 0.046473f
C4384 CSoutput.n263 gnd 0.35917f
C4385 CSoutput.n264 gnd 0.179638f
C4386 CSoutput.t115 gnd 0.046473f
C4387 CSoutput.t31 gnd 0.046473f
C4388 CSoutput.n265 gnd 0.35917f
C4389 CSoutput.n266 gnd 0.267886f
C4390 CSoutput.n267 gnd 0.337802f
C4391 CSoutput.t8 gnd 0.046473f
C4392 CSoutput.t25 gnd 0.046473f
C4393 CSoutput.n268 gnd 0.359811f
C4394 CSoutput.t110 gnd 0.046473f
C4395 CSoutput.t6 gnd 0.046473f
C4396 CSoutput.n269 gnd 0.35917f
C4397 CSoutput.n270 gnd 0.364557f
C4398 CSoutput.t17 gnd 0.046473f
C4399 CSoutput.t33 gnd 0.046473f
C4400 CSoutput.n271 gnd 0.35917f
C4401 CSoutput.n272 gnd 0.179638f
C4402 CSoutput.t29 gnd 0.046473f
C4403 CSoutput.t114 gnd 0.046473f
C4404 CSoutput.n273 gnd 0.359168f
C4405 CSoutput.n274 gnd 0.267887f
C4406 CSoutput.n275 gnd 0.377576f
C4407 CSoutput.n276 gnd 9.32377f
C4408 CSoutput.t67 gnd 0.040664f
C4409 CSoutput.t107 gnd 0.040664f
C4410 CSoutput.n277 gnd 0.360525f
C4411 CSoutput.t61 gnd 0.040664f
C4412 CSoutput.t66 gnd 0.040664f
C4413 CSoutput.n278 gnd 0.359322f
C4414 CSoutput.n279 gnd 0.334821f
C4415 CSoutput.t56 gnd 0.040664f
C4416 CSoutput.t70 gnd 0.040664f
C4417 CSoutput.n280 gnd 0.359322f
C4418 CSoutput.n281 gnd 0.165051f
C4419 CSoutput.t79 gnd 0.040664f
C4420 CSoutput.t62 gnd 0.040664f
C4421 CSoutput.n282 gnd 0.359322f
C4422 CSoutput.n283 gnd 0.165051f
C4423 CSoutput.t68 gnd 0.040664f
C4424 CSoutput.t96 gnd 0.040664f
C4425 CSoutput.n284 gnd 0.359322f
C4426 CSoutput.n285 gnd 0.165051f
C4427 CSoutput.t76 gnd 0.040664f
C4428 CSoutput.t83 gnd 0.040664f
C4429 CSoutput.n286 gnd 0.359322f
C4430 CSoutput.n287 gnd 0.304428f
C4431 CSoutput.t104 gnd 0.040664f
C4432 CSoutput.t37 gnd 0.040664f
C4433 CSoutput.n288 gnd 0.360525f
C4434 CSoutput.t46 gnd 0.040664f
C4435 CSoutput.t97 gnd 0.040664f
C4436 CSoutput.n289 gnd 0.359322f
C4437 CSoutput.n290 gnd 0.334821f
C4438 CSoutput.t38 gnd 0.040664f
C4439 CSoutput.t91 gnd 0.040664f
C4440 CSoutput.n291 gnd 0.359322f
C4441 CSoutput.n292 gnd 0.165051f
C4442 CSoutput.t98 gnd 0.040664f
C4443 CSoutput.t39 gnd 0.040664f
C4444 CSoutput.n293 gnd 0.359322f
C4445 CSoutput.n294 gnd 0.165051f
C4446 CSoutput.t85 gnd 0.040664f
C4447 CSoutput.t73 gnd 0.040664f
C4448 CSoutput.n295 gnd 0.359322f
C4449 CSoutput.n296 gnd 0.165051f
C4450 CSoutput.t40 gnd 0.040664f
C4451 CSoutput.t87 gnd 0.040664f
C4452 CSoutput.n297 gnd 0.359322f
C4453 CSoutput.n298 gnd 0.250583f
C4454 CSoutput.n299 gnd 0.316063f
C4455 CSoutput.t47 gnd 0.040664f
C4456 CSoutput.t99 gnd 0.040664f
C4457 CSoutput.n300 gnd 0.360525f
C4458 CSoutput.t60 gnd 0.040664f
C4459 CSoutput.t63 gnd 0.040664f
C4460 CSoutput.n301 gnd 0.359322f
C4461 CSoutput.n302 gnd 0.334821f
C4462 CSoutput.t41 gnd 0.040664f
C4463 CSoutput.t89 gnd 0.040664f
C4464 CSoutput.n303 gnd 0.359322f
C4465 CSoutput.n304 gnd 0.165051f
C4466 CSoutput.t69 gnd 0.040664f
C4467 CSoutput.t48 gnd 0.040664f
C4468 CSoutput.n305 gnd 0.359322f
C4469 CSoutput.n306 gnd 0.165051f
C4470 CSoutput.t53 gnd 0.040664f
C4471 CSoutput.t108 gnd 0.040664f
C4472 CSoutput.n307 gnd 0.359322f
C4473 CSoutput.n308 gnd 0.165051f
C4474 CSoutput.t54 gnd 0.040664f
C4475 CSoutput.t58 gnd 0.040664f
C4476 CSoutput.n309 gnd 0.359322f
C4477 CSoutput.n310 gnd 0.250583f
C4478 CSoutput.n311 gnd 0.339402f
C4479 CSoutput.n312 gnd 9.778309f
C4480 CSoutput.t57 gnd 0.040664f
C4481 CSoutput.t86 gnd 0.040664f
C4482 CSoutput.n313 gnd 0.360525f
C4483 CSoutput.t84 gnd 0.040664f
C4484 CSoutput.t72 gnd 0.040664f
C4485 CSoutput.n314 gnd 0.359322f
C4486 CSoutput.n315 gnd 0.334821f
C4487 CSoutput.t90 gnd 0.040664f
C4488 CSoutput.t64 gnd 0.040664f
C4489 CSoutput.n316 gnd 0.359322f
C4490 CSoutput.n317 gnd 0.165051f
C4491 CSoutput.t77 gnd 0.040664f
C4492 CSoutput.t100 gnd 0.040664f
C4493 CSoutput.n318 gnd 0.359322f
C4494 CSoutput.n319 gnd 0.165051f
C4495 CSoutput.t52 gnd 0.040664f
C4496 CSoutput.t88 gnd 0.040664f
C4497 CSoutput.n320 gnd 0.359322f
C4498 CSoutput.n321 gnd 0.165051f
C4499 CSoutput.t45 gnd 0.040664f
C4500 CSoutput.t92 gnd 0.040664f
C4501 CSoutput.n322 gnd 0.359322f
C4502 CSoutput.n323 gnd 0.304428f
C4503 CSoutput.t49 gnd 0.040664f
C4504 CSoutput.t44 gnd 0.040664f
C4505 CSoutput.n324 gnd 0.360525f
C4506 CSoutput.t42 gnd 0.040664f
C4507 CSoutput.t105 gnd 0.040664f
C4508 CSoutput.n325 gnd 0.359322f
C4509 CSoutput.n326 gnd 0.334821f
C4510 CSoutput.t106 gnd 0.040664f
C4511 CSoutput.t50 gnd 0.040664f
C4512 CSoutput.n327 gnd 0.359322f
C4513 CSoutput.n328 gnd 0.165051f
C4514 CSoutput.t51 gnd 0.040664f
C4515 CSoutput.t80 gnd 0.040664f
C4516 CSoutput.n329 gnd 0.359322f
C4517 CSoutput.n330 gnd 0.165051f
C4518 CSoutput.t81 gnd 0.040664f
C4519 CSoutput.t101 gnd 0.040664f
C4520 CSoutput.n331 gnd 0.359322f
C4521 CSoutput.n332 gnd 0.165051f
C4522 CSoutput.t102 gnd 0.040664f
C4523 CSoutput.t95 gnd 0.040664f
C4524 CSoutput.n333 gnd 0.359322f
C4525 CSoutput.n334 gnd 0.250583f
C4526 CSoutput.n335 gnd 0.316063f
C4527 CSoutput.t75 gnd 0.040664f
C4528 CSoutput.t93 gnd 0.040664f
C4529 CSoutput.n336 gnd 0.360525f
C4530 CSoutput.t55 gnd 0.040664f
C4531 CSoutput.t65 gnd 0.040664f
C4532 CSoutput.n337 gnd 0.359322f
C4533 CSoutput.n338 gnd 0.334821f
C4534 CSoutput.t71 gnd 0.040664f
C4535 CSoutput.t82 gnd 0.040664f
C4536 CSoutput.n339 gnd 0.359322f
C4537 CSoutput.n340 gnd 0.165051f
C4538 CSoutput.t94 gnd 0.040664f
C4539 CSoutput.t74 gnd 0.040664f
C4540 CSoutput.n341 gnd 0.359322f
C4541 CSoutput.n342 gnd 0.165051f
C4542 CSoutput.t78 gnd 0.040664f
C4543 CSoutput.t103 gnd 0.040664f
C4544 CSoutput.n343 gnd 0.359322f
C4545 CSoutput.n344 gnd 0.165051f
C4546 CSoutput.t43 gnd 0.040664f
C4547 CSoutput.t59 gnd 0.040664f
C4548 CSoutput.n345 gnd 0.359322f
C4549 CSoutput.n346 gnd 0.250583f
C4550 CSoutput.n347 gnd 0.339402f
C4551 CSoutput.n348 gnd 5.3586f
C4552 CSoutput.n349 gnd 11.3806f
C4553 commonsourceibias.n0 gnd 0.012292f
C4554 commonsourceibias.t89 gnd 0.186134f
C4555 commonsourceibias.t49 gnd 0.172107f
C4556 commonsourceibias.n1 gnd 0.068671f
C4557 commonsourceibias.n2 gnd 0.009212f
C4558 commonsourceibias.t95 gnd 0.172107f
C4559 commonsourceibias.n3 gnd 0.007452f
C4560 commonsourceibias.n4 gnd 0.009212f
C4561 commonsourceibias.t90 gnd 0.172107f
C4562 commonsourceibias.n5 gnd 0.008893f
C4563 commonsourceibias.n6 gnd 0.009212f
C4564 commonsourceibias.t100 gnd 0.172107f
C4565 commonsourceibias.n7 gnd 0.068671f
C4566 commonsourceibias.t86 gnd 0.172107f
C4567 commonsourceibias.n8 gnd 0.00744f
C4568 commonsourceibias.n9 gnd 0.012292f
C4569 commonsourceibias.t22 gnd 0.186134f
C4570 commonsourceibias.t0 gnd 0.172107f
C4571 commonsourceibias.n10 gnd 0.068671f
C4572 commonsourceibias.n11 gnd 0.009212f
C4573 commonsourceibias.t38 gnd 0.172107f
C4574 commonsourceibias.n12 gnd 0.007452f
C4575 commonsourceibias.n13 gnd 0.009212f
C4576 commonsourceibias.t20 gnd 0.172107f
C4577 commonsourceibias.n14 gnd 0.008893f
C4578 commonsourceibias.n15 gnd 0.009212f
C4579 commonsourceibias.t44 gnd 0.172107f
C4580 commonsourceibias.n16 gnd 0.068671f
C4581 commonsourceibias.t18 gnd 0.172107f
C4582 commonsourceibias.n17 gnd 0.00744f
C4583 commonsourceibias.n18 gnd 0.009212f
C4584 commonsourceibias.t8 gnd 0.172107f
C4585 commonsourceibias.t40 gnd 0.172107f
C4586 commonsourceibias.n19 gnd 0.068671f
C4587 commonsourceibias.n20 gnd 0.009212f
C4588 commonsourceibias.t24 gnd 0.172107f
C4589 commonsourceibias.n21 gnd 0.068671f
C4590 commonsourceibias.n22 gnd 0.009212f
C4591 commonsourceibias.t34 gnd 0.172107f
C4592 commonsourceibias.n23 gnd 0.068671f
C4593 commonsourceibias.n24 gnd 0.046375f
C4594 commonsourceibias.t4 gnd 0.172107f
C4595 commonsourceibias.t10 gnd 0.194203f
C4596 commonsourceibias.n25 gnd 0.079692f
C4597 commonsourceibias.n26 gnd 0.082502f
C4598 commonsourceibias.n27 gnd 0.011354f
C4599 commonsourceibias.n28 gnd 0.012561f
C4600 commonsourceibias.n29 gnd 0.009212f
C4601 commonsourceibias.n30 gnd 0.009212f
C4602 commonsourceibias.n31 gnd 0.012479f
C4603 commonsourceibias.n32 gnd 0.007452f
C4604 commonsourceibias.n33 gnd 0.012633f
C4605 commonsourceibias.n34 gnd 0.009212f
C4606 commonsourceibias.n35 gnd 0.009212f
C4607 commonsourceibias.n36 gnd 0.01271f
C4608 commonsourceibias.n37 gnd 0.01096f
C4609 commonsourceibias.n38 gnd 0.008893f
C4610 commonsourceibias.n39 gnd 0.009212f
C4611 commonsourceibias.n40 gnd 0.009212f
C4612 commonsourceibias.n41 gnd 0.011268f
C4613 commonsourceibias.n42 gnd 0.012647f
C4614 commonsourceibias.n43 gnd 0.068671f
C4615 commonsourceibias.n44 gnd 0.012562f
C4616 commonsourceibias.n45 gnd 0.009212f
C4617 commonsourceibias.n46 gnd 0.009212f
C4618 commonsourceibias.n47 gnd 0.009212f
C4619 commonsourceibias.n48 gnd 0.012562f
C4620 commonsourceibias.n49 gnd 0.068671f
C4621 commonsourceibias.n50 gnd 0.012647f
C4622 commonsourceibias.n51 gnd 0.011268f
C4623 commonsourceibias.n52 gnd 0.009212f
C4624 commonsourceibias.n53 gnd 0.009212f
C4625 commonsourceibias.n54 gnd 0.009212f
C4626 commonsourceibias.n55 gnd 0.01096f
C4627 commonsourceibias.n56 gnd 0.01271f
C4628 commonsourceibias.n57 gnd 0.068671f
C4629 commonsourceibias.n58 gnd 0.012633f
C4630 commonsourceibias.n59 gnd 0.009212f
C4631 commonsourceibias.n60 gnd 0.009212f
C4632 commonsourceibias.n61 gnd 0.009212f
C4633 commonsourceibias.n62 gnd 0.012479f
C4634 commonsourceibias.n63 gnd 0.068671f
C4635 commonsourceibias.n64 gnd 0.012561f
C4636 commonsourceibias.n65 gnd 0.011354f
C4637 commonsourceibias.n66 gnd 0.009212f
C4638 commonsourceibias.n67 gnd 0.009212f
C4639 commonsourceibias.n68 gnd 0.009345f
C4640 commonsourceibias.n69 gnd 0.009661f
C4641 commonsourceibias.n70 gnd 0.082165f
C4642 commonsourceibias.n71 gnd 0.09115f
C4643 commonsourceibias.t23 gnd 0.019878f
C4644 commonsourceibias.t1 gnd 0.019878f
C4645 commonsourceibias.n72 gnd 0.175652f
C4646 commonsourceibias.n73 gnd 0.151777f
C4647 commonsourceibias.t39 gnd 0.019878f
C4648 commonsourceibias.t21 gnd 0.019878f
C4649 commonsourceibias.n74 gnd 0.175652f
C4650 commonsourceibias.n75 gnd 0.080684f
C4651 commonsourceibias.t45 gnd 0.019878f
C4652 commonsourceibias.t19 gnd 0.019878f
C4653 commonsourceibias.n76 gnd 0.175652f
C4654 commonsourceibias.n77 gnd 0.067408f
C4655 commonsourceibias.t5 gnd 0.019878f
C4656 commonsourceibias.t11 gnd 0.019878f
C4657 commonsourceibias.n78 gnd 0.17624f
C4658 commonsourceibias.t25 gnd 0.019878f
C4659 commonsourceibias.t35 gnd 0.019878f
C4660 commonsourceibias.n79 gnd 0.175652f
C4661 commonsourceibias.n80 gnd 0.163675f
C4662 commonsourceibias.t9 gnd 0.019878f
C4663 commonsourceibias.t41 gnd 0.019878f
C4664 commonsourceibias.n81 gnd 0.175652f
C4665 commonsourceibias.n82 gnd 0.067408f
C4666 commonsourceibias.n83 gnd 0.081623f
C4667 commonsourceibias.n84 gnd 0.009212f
C4668 commonsourceibias.t77 gnd 0.172107f
C4669 commonsourceibias.t94 gnd 0.172107f
C4670 commonsourceibias.n85 gnd 0.068671f
C4671 commonsourceibias.n86 gnd 0.009212f
C4672 commonsourceibias.t88 gnd 0.172107f
C4673 commonsourceibias.n87 gnd 0.068671f
C4674 commonsourceibias.n88 gnd 0.009212f
C4675 commonsourceibias.t60 gnd 0.172107f
C4676 commonsourceibias.n89 gnd 0.068671f
C4677 commonsourceibias.n90 gnd 0.046375f
C4678 commonsourceibias.t80 gnd 0.172107f
C4679 commonsourceibias.t73 gnd 0.194203f
C4680 commonsourceibias.n91 gnd 0.079692f
C4681 commonsourceibias.n92 gnd 0.082502f
C4682 commonsourceibias.n93 gnd 0.011354f
C4683 commonsourceibias.n94 gnd 0.012561f
C4684 commonsourceibias.n95 gnd 0.009212f
C4685 commonsourceibias.n96 gnd 0.009212f
C4686 commonsourceibias.n97 gnd 0.012479f
C4687 commonsourceibias.n98 gnd 0.007452f
C4688 commonsourceibias.n99 gnd 0.012633f
C4689 commonsourceibias.n100 gnd 0.009212f
C4690 commonsourceibias.n101 gnd 0.009212f
C4691 commonsourceibias.n102 gnd 0.01271f
C4692 commonsourceibias.n103 gnd 0.01096f
C4693 commonsourceibias.n104 gnd 0.008893f
C4694 commonsourceibias.n105 gnd 0.009212f
C4695 commonsourceibias.n106 gnd 0.009212f
C4696 commonsourceibias.n107 gnd 0.011268f
C4697 commonsourceibias.n108 gnd 0.012647f
C4698 commonsourceibias.n109 gnd 0.068671f
C4699 commonsourceibias.n110 gnd 0.012562f
C4700 commonsourceibias.n111 gnd 0.009168f
C4701 commonsourceibias.n112 gnd 0.066591f
C4702 commonsourceibias.n113 gnd 0.009168f
C4703 commonsourceibias.n114 gnd 0.012562f
C4704 commonsourceibias.n115 gnd 0.068671f
C4705 commonsourceibias.n116 gnd 0.012647f
C4706 commonsourceibias.n117 gnd 0.011268f
C4707 commonsourceibias.n118 gnd 0.009212f
C4708 commonsourceibias.n119 gnd 0.009212f
C4709 commonsourceibias.n120 gnd 0.009212f
C4710 commonsourceibias.n121 gnd 0.01096f
C4711 commonsourceibias.n122 gnd 0.01271f
C4712 commonsourceibias.n123 gnd 0.068671f
C4713 commonsourceibias.n124 gnd 0.012633f
C4714 commonsourceibias.n125 gnd 0.009212f
C4715 commonsourceibias.n126 gnd 0.009212f
C4716 commonsourceibias.n127 gnd 0.009212f
C4717 commonsourceibias.n128 gnd 0.012479f
C4718 commonsourceibias.n129 gnd 0.068671f
C4719 commonsourceibias.n130 gnd 0.012561f
C4720 commonsourceibias.n131 gnd 0.011354f
C4721 commonsourceibias.n132 gnd 0.009212f
C4722 commonsourceibias.n133 gnd 0.009212f
C4723 commonsourceibias.n134 gnd 0.009345f
C4724 commonsourceibias.n135 gnd 0.009661f
C4725 commonsourceibias.n136 gnd 0.082165f
C4726 commonsourceibias.n137 gnd 0.053193f
C4727 commonsourceibias.n138 gnd 0.012292f
C4728 commonsourceibias.t52 gnd 0.186134f
C4729 commonsourceibias.t119 gnd 0.172107f
C4730 commonsourceibias.n139 gnd 0.068671f
C4731 commonsourceibias.n140 gnd 0.009212f
C4732 commonsourceibias.t110 gnd 0.172107f
C4733 commonsourceibias.n141 gnd 0.007452f
C4734 commonsourceibias.n142 gnd 0.009212f
C4735 commonsourceibias.t59 gnd 0.172107f
C4736 commonsourceibias.n143 gnd 0.008893f
C4737 commonsourceibias.n144 gnd 0.009212f
C4738 commonsourceibias.t118 gnd 0.172107f
C4739 commonsourceibias.n145 gnd 0.068671f
C4740 commonsourceibias.t65 gnd 0.172107f
C4741 commonsourceibias.n146 gnd 0.00744f
C4742 commonsourceibias.n147 gnd 0.009212f
C4743 commonsourceibias.t58 gnd 0.172107f
C4744 commonsourceibias.t117 gnd 0.172107f
C4745 commonsourceibias.n148 gnd 0.068671f
C4746 commonsourceibias.n149 gnd 0.009212f
C4747 commonsourceibias.t71 gnd 0.172107f
C4748 commonsourceibias.n150 gnd 0.068671f
C4749 commonsourceibias.n151 gnd 0.009212f
C4750 commonsourceibias.t83 gnd 0.172107f
C4751 commonsourceibias.n152 gnd 0.068671f
C4752 commonsourceibias.n153 gnd 0.046375f
C4753 commonsourceibias.t116 gnd 0.172107f
C4754 commonsourceibias.t69 gnd 0.194203f
C4755 commonsourceibias.n154 gnd 0.079692f
C4756 commonsourceibias.n155 gnd 0.082502f
C4757 commonsourceibias.n156 gnd 0.011354f
C4758 commonsourceibias.n157 gnd 0.012561f
C4759 commonsourceibias.n158 gnd 0.009212f
C4760 commonsourceibias.n159 gnd 0.009212f
C4761 commonsourceibias.n160 gnd 0.012479f
C4762 commonsourceibias.n161 gnd 0.007452f
C4763 commonsourceibias.n162 gnd 0.012633f
C4764 commonsourceibias.n163 gnd 0.009212f
C4765 commonsourceibias.n164 gnd 0.009212f
C4766 commonsourceibias.n165 gnd 0.01271f
C4767 commonsourceibias.n166 gnd 0.01096f
C4768 commonsourceibias.n167 gnd 0.008893f
C4769 commonsourceibias.n168 gnd 0.009212f
C4770 commonsourceibias.n169 gnd 0.009212f
C4771 commonsourceibias.n170 gnd 0.011268f
C4772 commonsourceibias.n171 gnd 0.012647f
C4773 commonsourceibias.n172 gnd 0.068671f
C4774 commonsourceibias.n173 gnd 0.012562f
C4775 commonsourceibias.n174 gnd 0.009212f
C4776 commonsourceibias.n175 gnd 0.009212f
C4777 commonsourceibias.n176 gnd 0.009212f
C4778 commonsourceibias.n177 gnd 0.012562f
C4779 commonsourceibias.n178 gnd 0.068671f
C4780 commonsourceibias.n179 gnd 0.012647f
C4781 commonsourceibias.n180 gnd 0.011268f
C4782 commonsourceibias.n181 gnd 0.009212f
C4783 commonsourceibias.n182 gnd 0.009212f
C4784 commonsourceibias.n183 gnd 0.009212f
C4785 commonsourceibias.n184 gnd 0.01096f
C4786 commonsourceibias.n185 gnd 0.01271f
C4787 commonsourceibias.n186 gnd 0.068671f
C4788 commonsourceibias.n187 gnd 0.012633f
C4789 commonsourceibias.n188 gnd 0.009212f
C4790 commonsourceibias.n189 gnd 0.009212f
C4791 commonsourceibias.n190 gnd 0.009212f
C4792 commonsourceibias.n191 gnd 0.012479f
C4793 commonsourceibias.n192 gnd 0.068671f
C4794 commonsourceibias.n193 gnd 0.012561f
C4795 commonsourceibias.n194 gnd 0.011354f
C4796 commonsourceibias.n195 gnd 0.009212f
C4797 commonsourceibias.n196 gnd 0.009212f
C4798 commonsourceibias.n197 gnd 0.009345f
C4799 commonsourceibias.n198 gnd 0.009661f
C4800 commonsourceibias.n199 gnd 0.082165f
C4801 commonsourceibias.n200 gnd 0.027962f
C4802 commonsourceibias.n201 gnd 0.146988f
C4803 commonsourceibias.n202 gnd 0.012292f
C4804 commonsourceibias.t57 gnd 0.172107f
C4805 commonsourceibias.n203 gnd 0.068671f
C4806 commonsourceibias.n204 gnd 0.009212f
C4807 commonsourceibias.t96 gnd 0.172107f
C4808 commonsourceibias.n205 gnd 0.007452f
C4809 commonsourceibias.n206 gnd 0.009212f
C4810 commonsourceibias.t93 gnd 0.172107f
C4811 commonsourceibias.n207 gnd 0.008893f
C4812 commonsourceibias.n208 gnd 0.009212f
C4813 commonsourceibias.t115 gnd 0.172107f
C4814 commonsourceibias.n209 gnd 0.068671f
C4815 commonsourceibias.t67 gnd 0.172107f
C4816 commonsourceibias.n210 gnd 0.00744f
C4817 commonsourceibias.n211 gnd 0.009212f
C4818 commonsourceibias.t87 gnd 0.172107f
C4819 commonsourceibias.t108 gnd 0.172107f
C4820 commonsourceibias.n212 gnd 0.068671f
C4821 commonsourceibias.n213 gnd 0.009212f
C4822 commonsourceibias.t103 gnd 0.172107f
C4823 commonsourceibias.n214 gnd 0.068671f
C4824 commonsourceibias.n215 gnd 0.009212f
C4825 commonsourceibias.t48 gnd 0.172107f
C4826 commonsourceibias.n216 gnd 0.068671f
C4827 commonsourceibias.n217 gnd 0.046375f
C4828 commonsourceibias.t102 gnd 0.172107f
C4829 commonsourceibias.t98 gnd 0.194203f
C4830 commonsourceibias.n218 gnd 0.079692f
C4831 commonsourceibias.n219 gnd 0.082502f
C4832 commonsourceibias.n220 gnd 0.011354f
C4833 commonsourceibias.n221 gnd 0.012561f
C4834 commonsourceibias.n222 gnd 0.009212f
C4835 commonsourceibias.n223 gnd 0.009212f
C4836 commonsourceibias.n224 gnd 0.012479f
C4837 commonsourceibias.n225 gnd 0.007452f
C4838 commonsourceibias.n226 gnd 0.012633f
C4839 commonsourceibias.n227 gnd 0.009212f
C4840 commonsourceibias.n228 gnd 0.009212f
C4841 commonsourceibias.n229 gnd 0.01271f
C4842 commonsourceibias.n230 gnd 0.01096f
C4843 commonsourceibias.n231 gnd 0.008893f
C4844 commonsourceibias.n232 gnd 0.009212f
C4845 commonsourceibias.n233 gnd 0.009212f
C4846 commonsourceibias.n234 gnd 0.011268f
C4847 commonsourceibias.n235 gnd 0.012647f
C4848 commonsourceibias.n236 gnd 0.068671f
C4849 commonsourceibias.n237 gnd 0.012562f
C4850 commonsourceibias.n238 gnd 0.009212f
C4851 commonsourceibias.n239 gnd 0.009212f
C4852 commonsourceibias.n240 gnd 0.009212f
C4853 commonsourceibias.n241 gnd 0.012562f
C4854 commonsourceibias.n242 gnd 0.068671f
C4855 commonsourceibias.n243 gnd 0.012647f
C4856 commonsourceibias.n244 gnd 0.011268f
C4857 commonsourceibias.n245 gnd 0.009212f
C4858 commonsourceibias.n246 gnd 0.009212f
C4859 commonsourceibias.n247 gnd 0.009212f
C4860 commonsourceibias.n248 gnd 0.01096f
C4861 commonsourceibias.n249 gnd 0.01271f
C4862 commonsourceibias.n250 gnd 0.068671f
C4863 commonsourceibias.n251 gnd 0.012633f
C4864 commonsourceibias.n252 gnd 0.009212f
C4865 commonsourceibias.n253 gnd 0.009212f
C4866 commonsourceibias.n254 gnd 0.009212f
C4867 commonsourceibias.n255 gnd 0.012479f
C4868 commonsourceibias.n256 gnd 0.068671f
C4869 commonsourceibias.n257 gnd 0.012561f
C4870 commonsourceibias.n258 gnd 0.011354f
C4871 commonsourceibias.n259 gnd 0.009212f
C4872 commonsourceibias.n260 gnd 0.009212f
C4873 commonsourceibias.n261 gnd 0.009345f
C4874 commonsourceibias.n262 gnd 0.009661f
C4875 commonsourceibias.t109 gnd 0.186134f
C4876 commonsourceibias.n263 gnd 0.082165f
C4877 commonsourceibias.n264 gnd 0.027962f
C4878 commonsourceibias.n265 gnd 0.437625f
C4879 commonsourceibias.n266 gnd 0.012292f
C4880 commonsourceibias.t70 gnd 0.186134f
C4881 commonsourceibias.t99 gnd 0.172107f
C4882 commonsourceibias.n267 gnd 0.068671f
C4883 commonsourceibias.n268 gnd 0.009212f
C4884 commonsourceibias.t84 gnd 0.172107f
C4885 commonsourceibias.n269 gnd 0.007452f
C4886 commonsourceibias.n270 gnd 0.009212f
C4887 commonsourceibias.t72 gnd 0.172107f
C4888 commonsourceibias.n271 gnd 0.008893f
C4889 commonsourceibias.n272 gnd 0.009212f
C4890 commonsourceibias.t66 gnd 0.172107f
C4891 commonsourceibias.n273 gnd 0.00744f
C4892 commonsourceibias.n274 gnd 0.009212f
C4893 commonsourceibias.t56 gnd 0.172107f
C4894 commonsourceibias.t79 gnd 0.172107f
C4895 commonsourceibias.n275 gnd 0.068671f
C4896 commonsourceibias.n276 gnd 0.009212f
C4897 commonsourceibias.t68 gnd 0.172107f
C4898 commonsourceibias.n277 gnd 0.068671f
C4899 commonsourceibias.n278 gnd 0.009212f
C4900 commonsourceibias.t104 gnd 0.172107f
C4901 commonsourceibias.n279 gnd 0.068671f
C4902 commonsourceibias.n280 gnd 0.046375f
C4903 commonsourceibias.t64 gnd 0.172107f
C4904 commonsourceibias.t111 gnd 0.194203f
C4905 commonsourceibias.n281 gnd 0.079692f
C4906 commonsourceibias.n282 gnd 0.082502f
C4907 commonsourceibias.n283 gnd 0.011354f
C4908 commonsourceibias.n284 gnd 0.012561f
C4909 commonsourceibias.n285 gnd 0.009212f
C4910 commonsourceibias.n286 gnd 0.009212f
C4911 commonsourceibias.n287 gnd 0.012479f
C4912 commonsourceibias.n288 gnd 0.007452f
C4913 commonsourceibias.n289 gnd 0.012633f
C4914 commonsourceibias.n290 gnd 0.009212f
C4915 commonsourceibias.n291 gnd 0.009212f
C4916 commonsourceibias.n292 gnd 0.01271f
C4917 commonsourceibias.n293 gnd 0.01096f
C4918 commonsourceibias.n294 gnd 0.008893f
C4919 commonsourceibias.n295 gnd 0.009212f
C4920 commonsourceibias.n296 gnd 0.009212f
C4921 commonsourceibias.n297 gnd 0.011268f
C4922 commonsourceibias.n298 gnd 0.012647f
C4923 commonsourceibias.n299 gnd 0.068671f
C4924 commonsourceibias.n300 gnd 0.012562f
C4925 commonsourceibias.n301 gnd 0.009168f
C4926 commonsourceibias.t3 gnd 0.019878f
C4927 commonsourceibias.t33 gnd 0.019878f
C4928 commonsourceibias.n302 gnd 0.17624f
C4929 commonsourceibias.t27 gnd 0.019878f
C4930 commonsourceibias.t17 gnd 0.019878f
C4931 commonsourceibias.n303 gnd 0.175652f
C4932 commonsourceibias.n304 gnd 0.163675f
C4933 commonsourceibias.t7 gnd 0.019878f
C4934 commonsourceibias.t37 gnd 0.019878f
C4935 commonsourceibias.n305 gnd 0.175652f
C4936 commonsourceibias.n306 gnd 0.067408f
C4937 commonsourceibias.n307 gnd 0.012292f
C4938 commonsourceibias.t46 gnd 0.172107f
C4939 commonsourceibias.n308 gnd 0.068671f
C4940 commonsourceibias.n309 gnd 0.009212f
C4941 commonsourceibias.t28 gnd 0.172107f
C4942 commonsourceibias.n310 gnd 0.007452f
C4943 commonsourceibias.n311 gnd 0.009212f
C4944 commonsourceibias.t12 gnd 0.172107f
C4945 commonsourceibias.n312 gnd 0.008893f
C4946 commonsourceibias.n313 gnd 0.009212f
C4947 commonsourceibias.t30 gnd 0.172107f
C4948 commonsourceibias.n314 gnd 0.00744f
C4949 commonsourceibias.n315 gnd 0.009212f
C4950 commonsourceibias.t36 gnd 0.172107f
C4951 commonsourceibias.t6 gnd 0.172107f
C4952 commonsourceibias.n316 gnd 0.068671f
C4953 commonsourceibias.n317 gnd 0.009212f
C4954 commonsourceibias.t16 gnd 0.172107f
C4955 commonsourceibias.n318 gnd 0.068671f
C4956 commonsourceibias.n319 gnd 0.009212f
C4957 commonsourceibias.t26 gnd 0.172107f
C4958 commonsourceibias.n320 gnd 0.068671f
C4959 commonsourceibias.n321 gnd 0.046375f
C4960 commonsourceibias.t32 gnd 0.172107f
C4961 commonsourceibias.t2 gnd 0.194203f
C4962 commonsourceibias.n322 gnd 0.079692f
C4963 commonsourceibias.n323 gnd 0.082502f
C4964 commonsourceibias.n324 gnd 0.011354f
C4965 commonsourceibias.n325 gnd 0.012561f
C4966 commonsourceibias.n326 gnd 0.009212f
C4967 commonsourceibias.n327 gnd 0.009212f
C4968 commonsourceibias.n328 gnd 0.012479f
C4969 commonsourceibias.n329 gnd 0.007452f
C4970 commonsourceibias.n330 gnd 0.012633f
C4971 commonsourceibias.n331 gnd 0.009212f
C4972 commonsourceibias.n332 gnd 0.009212f
C4973 commonsourceibias.n333 gnd 0.01271f
C4974 commonsourceibias.n334 gnd 0.01096f
C4975 commonsourceibias.n335 gnd 0.008893f
C4976 commonsourceibias.n336 gnd 0.009212f
C4977 commonsourceibias.n337 gnd 0.009212f
C4978 commonsourceibias.n338 gnd 0.011268f
C4979 commonsourceibias.n339 gnd 0.012647f
C4980 commonsourceibias.n340 gnd 0.068671f
C4981 commonsourceibias.n341 gnd 0.012562f
C4982 commonsourceibias.n342 gnd 0.009212f
C4983 commonsourceibias.n343 gnd 0.009212f
C4984 commonsourceibias.n344 gnd 0.009212f
C4985 commonsourceibias.n345 gnd 0.012562f
C4986 commonsourceibias.n346 gnd 0.068671f
C4987 commonsourceibias.n347 gnd 0.012647f
C4988 commonsourceibias.t42 gnd 0.172107f
C4989 commonsourceibias.n348 gnd 0.068671f
C4990 commonsourceibias.n349 gnd 0.011268f
C4991 commonsourceibias.n350 gnd 0.009212f
C4992 commonsourceibias.n351 gnd 0.009212f
C4993 commonsourceibias.n352 gnd 0.009212f
C4994 commonsourceibias.n353 gnd 0.01096f
C4995 commonsourceibias.n354 gnd 0.01271f
C4996 commonsourceibias.n355 gnd 0.068671f
C4997 commonsourceibias.n356 gnd 0.012633f
C4998 commonsourceibias.n357 gnd 0.009212f
C4999 commonsourceibias.n358 gnd 0.009212f
C5000 commonsourceibias.n359 gnd 0.009212f
C5001 commonsourceibias.n360 gnd 0.012479f
C5002 commonsourceibias.n361 gnd 0.068671f
C5003 commonsourceibias.n362 gnd 0.012561f
C5004 commonsourceibias.n363 gnd 0.011354f
C5005 commonsourceibias.n364 gnd 0.009212f
C5006 commonsourceibias.n365 gnd 0.009212f
C5007 commonsourceibias.n366 gnd 0.009345f
C5008 commonsourceibias.n367 gnd 0.009661f
C5009 commonsourceibias.t14 gnd 0.186134f
C5010 commonsourceibias.n368 gnd 0.082165f
C5011 commonsourceibias.n369 gnd 0.09115f
C5012 commonsourceibias.t47 gnd 0.019878f
C5013 commonsourceibias.t15 gnd 0.019878f
C5014 commonsourceibias.n370 gnd 0.175652f
C5015 commonsourceibias.n371 gnd 0.151777f
C5016 commonsourceibias.t13 gnd 0.019878f
C5017 commonsourceibias.t29 gnd 0.019878f
C5018 commonsourceibias.n372 gnd 0.175652f
C5019 commonsourceibias.n373 gnd 0.080684f
C5020 commonsourceibias.t31 gnd 0.019878f
C5021 commonsourceibias.t43 gnd 0.019878f
C5022 commonsourceibias.n374 gnd 0.175652f
C5023 commonsourceibias.n375 gnd 0.067408f
C5024 commonsourceibias.n376 gnd 0.081623f
C5025 commonsourceibias.n377 gnd 0.066591f
C5026 commonsourceibias.n378 gnd 0.009168f
C5027 commonsourceibias.n379 gnd 0.012562f
C5028 commonsourceibias.n380 gnd 0.068671f
C5029 commonsourceibias.n381 gnd 0.012647f
C5030 commonsourceibias.t92 gnd 0.172107f
C5031 commonsourceibias.n382 gnd 0.068671f
C5032 commonsourceibias.n383 gnd 0.011268f
C5033 commonsourceibias.n384 gnd 0.009212f
C5034 commonsourceibias.n385 gnd 0.009212f
C5035 commonsourceibias.n386 gnd 0.009212f
C5036 commonsourceibias.n387 gnd 0.01096f
C5037 commonsourceibias.n388 gnd 0.01271f
C5038 commonsourceibias.n389 gnd 0.068671f
C5039 commonsourceibias.n390 gnd 0.012633f
C5040 commonsourceibias.n391 gnd 0.009212f
C5041 commonsourceibias.n392 gnd 0.009212f
C5042 commonsourceibias.n393 gnd 0.009212f
C5043 commonsourceibias.n394 gnd 0.012479f
C5044 commonsourceibias.n395 gnd 0.068671f
C5045 commonsourceibias.n396 gnd 0.012561f
C5046 commonsourceibias.n397 gnd 0.011354f
C5047 commonsourceibias.n398 gnd 0.009212f
C5048 commonsourceibias.n399 gnd 0.009212f
C5049 commonsourceibias.n400 gnd 0.009345f
C5050 commonsourceibias.n401 gnd 0.009661f
C5051 commonsourceibias.n402 gnd 0.082165f
C5052 commonsourceibias.n403 gnd 0.053193f
C5053 commonsourceibias.n404 gnd 0.012292f
C5054 commonsourceibias.t107 gnd 0.172107f
C5055 commonsourceibias.n405 gnd 0.068671f
C5056 commonsourceibias.n406 gnd 0.009212f
C5057 commonsourceibias.t51 gnd 0.172107f
C5058 commonsourceibias.n407 gnd 0.007452f
C5059 commonsourceibias.n408 gnd 0.009212f
C5060 commonsourceibias.t114 gnd 0.172107f
C5061 commonsourceibias.n409 gnd 0.008893f
C5062 commonsourceibias.n410 gnd 0.009212f
C5063 commonsourceibias.t50 gnd 0.172107f
C5064 commonsourceibias.n411 gnd 0.00744f
C5065 commonsourceibias.n412 gnd 0.009212f
C5066 commonsourceibias.t76 gnd 0.172107f
C5067 commonsourceibias.t105 gnd 0.172107f
C5068 commonsourceibias.n413 gnd 0.068671f
C5069 commonsourceibias.n414 gnd 0.009212f
C5070 commonsourceibias.t55 gnd 0.172107f
C5071 commonsourceibias.n415 gnd 0.068671f
C5072 commonsourceibias.n416 gnd 0.009212f
C5073 commonsourceibias.t75 gnd 0.172107f
C5074 commonsourceibias.n417 gnd 0.068671f
C5075 commonsourceibias.n418 gnd 0.046375f
C5076 commonsourceibias.t61 gnd 0.172107f
C5077 commonsourceibias.t54 gnd 0.194203f
C5078 commonsourceibias.n419 gnd 0.079692f
C5079 commonsourceibias.n420 gnd 0.082502f
C5080 commonsourceibias.n421 gnd 0.011354f
C5081 commonsourceibias.n422 gnd 0.012561f
C5082 commonsourceibias.n423 gnd 0.009212f
C5083 commonsourceibias.n424 gnd 0.009212f
C5084 commonsourceibias.n425 gnd 0.012479f
C5085 commonsourceibias.n426 gnd 0.007452f
C5086 commonsourceibias.n427 gnd 0.012633f
C5087 commonsourceibias.n428 gnd 0.009212f
C5088 commonsourceibias.n429 gnd 0.009212f
C5089 commonsourceibias.n430 gnd 0.01271f
C5090 commonsourceibias.n431 gnd 0.01096f
C5091 commonsourceibias.n432 gnd 0.008893f
C5092 commonsourceibias.n433 gnd 0.009212f
C5093 commonsourceibias.n434 gnd 0.009212f
C5094 commonsourceibias.n435 gnd 0.011268f
C5095 commonsourceibias.n436 gnd 0.012647f
C5096 commonsourceibias.n437 gnd 0.068671f
C5097 commonsourceibias.n438 gnd 0.012562f
C5098 commonsourceibias.n439 gnd 0.009212f
C5099 commonsourceibias.n440 gnd 0.009212f
C5100 commonsourceibias.n441 gnd 0.009212f
C5101 commonsourceibias.n442 gnd 0.012562f
C5102 commonsourceibias.n443 gnd 0.068671f
C5103 commonsourceibias.n444 gnd 0.012647f
C5104 commonsourceibias.t106 gnd 0.172107f
C5105 commonsourceibias.n445 gnd 0.068671f
C5106 commonsourceibias.n446 gnd 0.011268f
C5107 commonsourceibias.n447 gnd 0.009212f
C5108 commonsourceibias.n448 gnd 0.009212f
C5109 commonsourceibias.n449 gnd 0.009212f
C5110 commonsourceibias.n450 gnd 0.01096f
C5111 commonsourceibias.n451 gnd 0.01271f
C5112 commonsourceibias.n452 gnd 0.068671f
C5113 commonsourceibias.n453 gnd 0.012633f
C5114 commonsourceibias.n454 gnd 0.009212f
C5115 commonsourceibias.n455 gnd 0.009212f
C5116 commonsourceibias.n456 gnd 0.009212f
C5117 commonsourceibias.n457 gnd 0.012479f
C5118 commonsourceibias.n458 gnd 0.068671f
C5119 commonsourceibias.n459 gnd 0.012561f
C5120 commonsourceibias.n460 gnd 0.011354f
C5121 commonsourceibias.n461 gnd 0.009212f
C5122 commonsourceibias.n462 gnd 0.009212f
C5123 commonsourceibias.n463 gnd 0.009345f
C5124 commonsourceibias.n464 gnd 0.009661f
C5125 commonsourceibias.t112 gnd 0.186134f
C5126 commonsourceibias.n465 gnd 0.082165f
C5127 commonsourceibias.n466 gnd 0.027962f
C5128 commonsourceibias.n467 gnd 0.146988f
C5129 commonsourceibias.n468 gnd 0.012292f
C5130 commonsourceibias.t81 gnd 0.172107f
C5131 commonsourceibias.n469 gnd 0.068671f
C5132 commonsourceibias.n470 gnd 0.009212f
C5133 commonsourceibias.t91 gnd 0.172107f
C5134 commonsourceibias.n471 gnd 0.007452f
C5135 commonsourceibias.n472 gnd 0.009212f
C5136 commonsourceibias.t101 gnd 0.172107f
C5137 commonsourceibias.n473 gnd 0.008893f
C5138 commonsourceibias.n474 gnd 0.009212f
C5139 commonsourceibias.t85 gnd 0.172107f
C5140 commonsourceibias.n475 gnd 0.00744f
C5141 commonsourceibias.n476 gnd 0.009212f
C5142 commonsourceibias.t82 gnd 0.172107f
C5143 commonsourceibias.t62 gnd 0.172107f
C5144 commonsourceibias.n477 gnd 0.068671f
C5145 commonsourceibias.n478 gnd 0.009212f
C5146 commonsourceibias.t53 gnd 0.172107f
C5147 commonsourceibias.n479 gnd 0.068671f
C5148 commonsourceibias.n480 gnd 0.009212f
C5149 commonsourceibias.t78 gnd 0.172107f
C5150 commonsourceibias.n481 gnd 0.068671f
C5151 commonsourceibias.n482 gnd 0.046375f
C5152 commonsourceibias.t97 gnd 0.172107f
C5153 commonsourceibias.t113 gnd 0.194203f
C5154 commonsourceibias.n483 gnd 0.079692f
C5155 commonsourceibias.n484 gnd 0.082502f
C5156 commonsourceibias.n485 gnd 0.011354f
C5157 commonsourceibias.n486 gnd 0.012561f
C5158 commonsourceibias.n487 gnd 0.009212f
C5159 commonsourceibias.n488 gnd 0.009212f
C5160 commonsourceibias.n489 gnd 0.012479f
C5161 commonsourceibias.n490 gnd 0.007452f
C5162 commonsourceibias.n491 gnd 0.012633f
C5163 commonsourceibias.n492 gnd 0.009212f
C5164 commonsourceibias.n493 gnd 0.009212f
C5165 commonsourceibias.n494 gnd 0.01271f
C5166 commonsourceibias.n495 gnd 0.01096f
C5167 commonsourceibias.n496 gnd 0.008893f
C5168 commonsourceibias.n497 gnd 0.009212f
C5169 commonsourceibias.n498 gnd 0.009212f
C5170 commonsourceibias.n499 gnd 0.011268f
C5171 commonsourceibias.n500 gnd 0.012647f
C5172 commonsourceibias.n501 gnd 0.068671f
C5173 commonsourceibias.n502 gnd 0.012562f
C5174 commonsourceibias.n503 gnd 0.009212f
C5175 commonsourceibias.n504 gnd 0.009212f
C5176 commonsourceibias.n505 gnd 0.009212f
C5177 commonsourceibias.n506 gnd 0.012562f
C5178 commonsourceibias.n507 gnd 0.068671f
C5179 commonsourceibias.n508 gnd 0.012647f
C5180 commonsourceibias.t74 gnd 0.172107f
C5181 commonsourceibias.n509 gnd 0.068671f
C5182 commonsourceibias.n510 gnd 0.011268f
C5183 commonsourceibias.n511 gnd 0.009212f
C5184 commonsourceibias.n512 gnd 0.009212f
C5185 commonsourceibias.n513 gnd 0.009212f
C5186 commonsourceibias.n514 gnd 0.01096f
C5187 commonsourceibias.n515 gnd 0.01271f
C5188 commonsourceibias.n516 gnd 0.068671f
C5189 commonsourceibias.n517 gnd 0.012633f
C5190 commonsourceibias.n518 gnd 0.009212f
C5191 commonsourceibias.n519 gnd 0.009212f
C5192 commonsourceibias.n520 gnd 0.009212f
C5193 commonsourceibias.n521 gnd 0.012479f
C5194 commonsourceibias.n522 gnd 0.068671f
C5195 commonsourceibias.n523 gnd 0.012561f
C5196 commonsourceibias.n524 gnd 0.011354f
C5197 commonsourceibias.n525 gnd 0.009212f
C5198 commonsourceibias.n526 gnd 0.009212f
C5199 commonsourceibias.n527 gnd 0.009345f
C5200 commonsourceibias.n528 gnd 0.009661f
C5201 commonsourceibias.t63 gnd 0.186134f
C5202 commonsourceibias.n529 gnd 0.082165f
C5203 commonsourceibias.n530 gnd 0.027962f
C5204 commonsourceibias.n531 gnd 0.194173f
C5205 commonsourceibias.n532 gnd 4.69557f
.ends

