* NGSPICE file created from opamp.ext - technology: sky130A

.subckt opamp output vdd plus minus commonsourceibias outputibias diffpairibias gnd CSoutput
Cload output gnd 0.0p
X0 CSoutput.t135 commonsourceibias.t64 gnd.t355 gnd.t286 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X1 CSoutput.t144 a_n1986_8322.t8 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X2 vdd.t64 a_n5644_8799.t32 CSoutput.t139 vdd.t11 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X3 a_n1986_8322.t9 a_n2356_n452.t44 vdd.t178 vdd.t177 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 a_n1808_13878.t11 a_n2356_n452.t18 a_n2356_n452.t19 vdd.t197 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X5 CSoutput.t134 commonsourceibias.t65 gnd.t354 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X6 a_n5644_8799.t15 plus.t5 a_n2903_n3924.t26 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X7 CSoutput.t133 commonsourceibias.t66 gnd.t353 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 gnd.t350 commonsourceibias.t67 CSoutput.t132 gnd.t277 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X9 a_n2903_n3924.t25 plus.t6 a_n5644_8799.t21 gnd.t193 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X10 a_n2356_n452.t21 a_n2356_n452.t20 a_n1808_13878.t10 vdd.t156 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X11 a_n1808_13878.t9 a_n2356_n452.t14 a_n2356_n452.t15 vdd.t153 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X12 vdd.t140 vdd.t138 vdd.t139 vdd.t113 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X13 a_n1808_13878.t19 a_n2356_n452.t45 vdd.t199 vdd.t198 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X14 CSoutput.t30 a_n5644_8799.t33 vdd.t63 vdd.t7 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X15 vdd.t137 vdd.t135 vdd.t136 vdd.t88 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X16 gnd.t352 commonsourceibias.t68 CSoutput.t131 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X17 CSoutput.t130 commonsourceibias.t69 gnd.t351 gnd.t275 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X18 CSoutput.t129 commonsourceibias.t70 gnd.t349 gnd.t275 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 CSoutput.t128 commonsourceibias.t71 gnd.t348 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 gnd.t347 commonsourceibias.t72 CSoutput.t127 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X21 gnd.t346 commonsourceibias.t73 CSoutput.t126 gnd.t256 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X22 vdd.t160 CSoutput.t145 output.t18 gnd.t181 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X23 commonsourceibias.t9 commonsourceibias.t8 gnd.t345 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X24 CSoutput.t125 commonsourceibias.t74 gnd.t344 gnd.t290 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X25 a_n1986_8322.t20 a_n2356_n452.t46 a_n5644_8799.t30 vdd.t145 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X26 CSoutput.t124 commonsourceibias.t75 gnd.t343 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X27 a_n2356_n452.t32 minus.t5 a_n2903_n3924.t34 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X28 a_n5644_8799.t3 plus.t7 a_n2903_n3924.t24 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X29 a_n2356_n452.t35 minus.t6 a_n2903_n3924.t37 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X30 gnd.t172 gnd.t169 gnd.t171 gnd.t170 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X31 CSoutput.t146 a_n1986_8322.t8 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X32 CSoutput.t123 commonsourceibias.t76 gnd.t340 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X33 gnd.t342 commonsourceibias.t77 CSoutput.t122 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X34 CSoutput.t121 commonsourceibias.t78 gnd.t341 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 CSoutput.t120 commonsourceibias.t79 gnd.t339 gnd.t286 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X36 gnd.t168 gnd.t166 gnd.t167 gnd.t91 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X37 gnd.t165 gnd.t163 gnd.t164 gnd.t74 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X38 CSoutput.t22 a_n5644_8799.t34 vdd.t62 vdd.t20 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X39 vdd.t61 a_n5644_8799.t35 CSoutput.t20 vdd.t38 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X40 a_n2903_n3924.t23 plus.t8 a_n5644_8799.t27 gnd.t357 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X41 CSoutput.t119 commonsourceibias.t80 gnd.t338 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X42 a_n5644_8799.t25 a_n2356_n452.t47 a_n1986_8322.t18 vdd.t197 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X43 CSoutput.t11 a_n5644_8799.t36 vdd.t60 vdd.t1 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X44 vdd.t59 a_n5644_8799.t37 CSoutput.t9 vdd.t54 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X45 a_n2903_n3924.t28 minus.t7 a_n2356_n452.t29 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X46 gnd.t337 commonsourceibias.t81 CSoutput.t118 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X47 a_n2903_n3924.t30 diffpairibias.t16 gnd.t49 gnd.t48 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X48 CSoutput.t117 commonsourceibias.t82 gnd.t336 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X49 gnd.t335 commonsourceibias.t10 commonsourceibias.t11 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X50 output.t19 outputibias.t8 gnd.t180 gnd.t179 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X51 CSoutput.t116 commonsourceibias.t83 gnd.t334 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 CSoutput.t19 a_n5644_8799.t38 vdd.t58 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X53 vdd.t134 vdd.t132 vdd.t133 vdd.t66 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X54 gnd.t333 commonsourceibias.t84 CSoutput.t115 gnd.t282 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X55 CSoutput.t114 commonsourceibias.t85 gnd.t332 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X56 CSoutput.t113 commonsourceibias.t86 gnd.t331 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X57 gnd.t330 commonsourceibias.t87 CSoutput.t112 gnd.t282 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X58 output.t17 CSoutput.t147 vdd.t161 gnd.t194 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X59 gnd.t327 commonsourceibias.t88 CSoutput.t111 gnd.t277 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X60 plus.t4 gnd.t160 gnd.t162 gnd.t161 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X61 CSoutput.t110 commonsourceibias.t89 gnd.t329 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X62 a_n2903_n3924.t22 plus.t9 a_n5644_8799.t18 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X63 gnd.t159 gnd.t157 gnd.t158 gnd.t91 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X64 CSoutput.t109 commonsourceibias.t90 gnd.t328 gnd.t275 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X65 gnd.t326 commonsourceibias.t14 commonsourceibias.t15 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X66 a_n1808_13878.t8 a_n2356_n452.t24 a_n2356_n452.t25 vdd.t179 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X67 vdd.t57 a_n5644_8799.t39 CSoutput.t7 vdd.t54 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X68 gnd.t156 gnd.t154 gnd.t155 gnd.t111 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X69 a_n2903_n3924.t21 plus.t10 a_n5644_8799.t24 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X70 diffpairibias.t15 diffpairibias.t14 gnd.t12 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X71 a_n2356_n452.t11 a_n2356_n452.t10 a_n1808_13878.t7 vdd.t182 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X72 CSoutput.t31 a_n5644_8799.t40 vdd.t56 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X73 gnd.t325 commonsourceibias.t91 CSoutput.t108 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X74 CSoutput.t107 commonsourceibias.t92 gnd.t324 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X75 CSoutput.t106 commonsourceibias.t93 gnd.t323 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X76 vdd.t131 vdd.t129 vdd.t130 vdd.t98 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X77 gnd.t322 commonsourceibias.t94 CSoutput.t105 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X78 gnd.t320 commonsourceibias.t95 CSoutput.t104 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X79 CSoutput.t103 commonsourceibias.t96 gnd.t321 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 diffpairibias.t13 diffpairibias.t12 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X81 gnd.t319 commonsourceibias.t12 commonsourceibias.t13 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X82 vdd.t128 vdd.t126 vdd.t127 vdd.t77 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X83 CSoutput.t102 commonsourceibias.t97 gnd.t318 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X84 CSoutput.t101 commonsourceibias.t98 gnd.t317 gnd.t290 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 gnd.t153 gnd.t151 gnd.t152 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X86 gnd.t316 commonsourceibias.t99 CSoutput.t100 gnd.t256 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X87 CSoutput.t99 commonsourceibias.t100 gnd.t315 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 gnd.t314 commonsourceibias.t101 CSoutput.t98 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 vdd.t55 a_n5644_8799.t41 CSoutput.t142 vdd.t54 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X90 gnd.t313 commonsourceibias.t102 CSoutput.t97 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 output.t16 CSoutput.t148 vdd.t170 gnd.t195 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X92 vdd.t53 a_n5644_8799.t42 CSoutput.t12 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X93 CSoutput.t27 a_n5644_8799.t43 vdd.t52 vdd.t1 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X94 a_n2903_n3924.t32 minus.t8 a_n2356_n452.t31 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X95 CSoutput.t149 a_n1986_8322.t8 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X96 a_n2903_n3924.t20 plus.t11 a_n5644_8799.t22 gnd.t13 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X97 gnd.t312 commonsourceibias.t18 commonsourceibias.t19 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X98 vdd.t51 a_n5644_8799.t44 CSoutput.t29 vdd.t5 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X99 gnd.t150 gnd.t148 minus.t4 gnd.t149 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X100 a_n5644_8799.t29 plus.t12 a_n2903_n3924.t19 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X101 gnd.t147 gnd.t145 gnd.t146 gnd.t70 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X102 gnd.t311 commonsourceibias.t103 CSoutput.t96 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X103 CSoutput.t34 a_n5644_8799.t45 vdd.t50 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X104 CSoutput.t26 a_n5644_8799.t46 vdd.t49 vdd.t42 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X105 vdd.t174 CSoutput.t150 output.t15 gnd.t182 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X106 output.t14 CSoutput.t151 vdd.t173 gnd.t183 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X107 a_n2903_n3924.t46 diffpairibias.t17 gnd.t359 gnd.t358 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X108 CSoutput.t140 a_n5644_8799.t47 vdd.t48 vdd.t42 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X109 a_n2903_n3924.t18 plus.t13 a_n5644_8799.t11 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X110 gnd.t310 commonsourceibias.t104 CSoutput.t95 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X111 gnd.t144 gnd.t142 gnd.t143 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X112 vdd.t47 a_n5644_8799.t48 CSoutput.t143 vdd.t40 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X113 gnd.t141 gnd.t139 gnd.t140 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X114 CSoutput.t94 commonsourceibias.t105 gnd.t308 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X115 a_n2356_n452.t7 a_n2356_n452.t6 a_n1808_13878.t6 vdd.t145 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X116 a_n2356_n452.t23 a_n2356_n452.t22 a_n1808_13878.t5 vdd.t186 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X117 vdd.t46 a_n5644_8799.t49 CSoutput.t3 vdd.t38 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X118 a_n5644_8799.t26 a_n2356_n452.t48 a_n1986_8322.t19 vdd.t185 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X119 gnd.t307 commonsourceibias.t106 CSoutput.t93 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X120 vdd.t45 a_n5644_8799.t50 CSoutput.t136 vdd.t40 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X121 gnd.t309 commonsourceibias.t107 CSoutput.t92 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X122 gnd.t306 commonsourceibias.t16 commonsourceibias.t17 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X123 output.t2 outputibias.t9 gnd.t42 gnd.t41 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X124 vdd.t125 vdd.t123 vdd.t124 vdd.t77 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X125 output.t13 CSoutput.t152 vdd.t172 gnd.t184 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X126 CSoutput.t153 a_n1986_8322.t8 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X127 vdd.t44 a_n5644_8799.t51 CSoutput.t6 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X128 vdd.t122 vdd.t120 vdd.t121 vdd.t106 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X129 vdd.t119 vdd.t116 vdd.t118 vdd.t117 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X130 CSoutput.t91 commonsourceibias.t108 gnd.t305 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X131 gnd.t304 commonsourceibias.t109 CSoutput.t90 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X132 CSoutput.t89 commonsourceibias.t110 gnd.t303 gnd.t290 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X133 gnd.t302 commonsourceibias.t111 CSoutput.t88 gnd.t282 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X134 gnd.t138 gnd.t135 gnd.t137 gnd.t136 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X135 a_n2903_n3924.t4 diffpairibias.t18 gnd.t10 gnd.t9 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X136 gnd.t300 commonsourceibias.t112 CSoutput.t87 gnd.t256 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X137 gnd.t301 commonsourceibias.t22 commonsourceibias.t23 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X138 vdd.t115 vdd.t112 vdd.t114 vdd.t113 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X139 CSoutput.t86 commonsourceibias.t113 gnd.t299 gnd.t286 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X140 output.t12 CSoutput.t154 vdd.t168 gnd.t185 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X141 CSoutput.t155 a_n1986_8322.t8 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X142 vdd.t190 a_n2356_n452.t49 a_n1986_8322.t15 vdd.t189 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X143 vdd.t111 vdd.t109 vdd.t110 vdd.t102 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X144 CSoutput.t14 a_n5644_8799.t52 vdd.t43 vdd.t42 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X145 a_n1986_8322.t16 a_n2356_n452.t50 vdd.t192 vdd.t191 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X146 vdd.t41 a_n5644_8799.t53 CSoutput.t28 vdd.t40 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X147 plus.t3 gnd.t132 gnd.t134 gnd.t133 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X148 gnd.t131 gnd.t129 gnd.t130 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X149 vdd.t158 a_n2356_n452.t51 a_n1808_13878.t18 vdd.t157 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X150 gnd.t128 gnd.t126 minus.t3 gnd.t127 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X151 a_n2356_n452.t34 minus.t9 a_n2903_n3924.t36 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X152 a_n5644_8799.t4 plus.t14 a_n2903_n3924.t17 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X153 vdd.t108 vdd.t105 vdd.t107 vdd.t106 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X154 a_n5644_8799.t14 plus.t15 a_n2903_n3924.t16 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X155 diffpairibias.t11 diffpairibias.t10 gnd.t25 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X156 vdd.t104 vdd.t101 vdd.t103 vdd.t102 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X157 vdd.t39 a_n5644_8799.t54 CSoutput.t1 vdd.t38 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X158 CSoutput.t85 commonsourceibias.t114 gnd.t297 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X159 gnd.t296 commonsourceibias.t115 CSoutput.t84 gnd.t277 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X160 commonsourceibias.t21 commonsourceibias.t20 gnd.t298 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X161 a_n5644_8799.t6 a_n2356_n452.t52 a_n1986_8322.t7 vdd.t159 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X162 a_n1986_8322.t4 a_n2356_n452.t53 vdd.t152 vdd.t151 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X163 vdd.t100 vdd.t97 vdd.t99 vdd.t98 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X164 CSoutput.t83 commonsourceibias.t116 gnd.t295 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 vdd.t169 CSoutput.t156 output.t11 gnd.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X166 a_n2356_n452.t17 a_n2356_n452.t16 a_n1808_13878.t4 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X167 a_n5644_8799.t2 a_n2356_n452.t54 a_n1986_8322.t5 vdd.t153 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X168 gnd.t125 gnd.t123 minus.t2 gnd.t124 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X169 gnd.t122 gnd.t120 gnd.t121 gnd.t74 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X170 CSoutput.t82 commonsourceibias.t117 gnd.t294 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X171 a_n1808_13878.t3 a_n2356_n452.t2 a_n2356_n452.t3 vdd.t185 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X172 gnd.t293 commonsourceibias.t118 CSoutput.t81 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X173 gnd.t292 commonsourceibias.t119 CSoutput.t80 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X174 a_n2903_n3924.t15 plus.t16 a_n5644_8799.t7 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X175 a_n2356_n452.t33 minus.t10 a_n2903_n3924.t35 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X176 outputibias.t7 outputibias.t6 gnd.t38 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X177 vdd.t175 CSoutput.t157 output.t10 gnd.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X178 commonsourceibias.t31 commonsourceibias.t30 gnd.t291 gnd.t290 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X179 gnd.t289 commonsourceibias.t120 CSoutput.t79 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X180 outputibias.t5 outputibias.t4 gnd.t44 gnd.t43 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X181 vdd.t194 a_n2356_n452.t55 a_n1986_8322.t17 vdd.t193 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X182 CSoutput.t78 commonsourceibias.t121 gnd.t288 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X183 vdd.t96 vdd.t94 vdd.t95 vdd.t88 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X184 gnd.t86 gnd.t83 gnd.t85 gnd.t84 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X185 a_n2903_n3924.t1 diffpairibias.t19 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X186 CSoutput.t141 a_n5644_8799.t55 vdd.t37 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X187 a_n5644_8799.t31 plus.t17 a_n2903_n3924.t14 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X188 a_n2903_n3924.t33 diffpairibias.t20 gnd.t175 gnd.t174 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X189 commonsourceibias.t29 commonsourceibias.t28 gnd.t287 gnd.t286 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X190 vdd.t36 a_n5644_8799.t56 CSoutput.t24 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X191 gnd.t119 gnd.t117 gnd.t118 gnd.t91 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X192 gnd.t116 gnd.t114 gnd.t115 gnd.t74 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X193 a_n5644_8799.t9 plus.t18 a_n2903_n3924.t13 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X194 CSoutput.t77 commonsourceibias.t122 gnd.t285 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X195 CSoutput.t76 commonsourceibias.t123 gnd.t281 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 vdd.t35 a_n5644_8799.t57 CSoutput.t37 vdd.t18 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X197 commonsourceibias.t27 commonsourceibias.t26 gnd.t284 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X198 gnd.t283 commonsourceibias.t24 commonsourceibias.t25 gnd.t282 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X199 diffpairibias.t9 diffpairibias.t8 gnd.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X200 CSoutput.t75 commonsourceibias.t124 gnd.t280 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X201 CSoutput.t74 commonsourceibias.t125 gnd.t279 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X202 a_n2356_n452.t28 minus.t11 a_n2903_n3924.t27 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X203 output.t9 CSoutput.t158 vdd.t163 gnd.t21 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X204 a_n2903_n3924.t12 plus.t19 a_n5644_8799.t28 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X205 gnd.t278 commonsourceibias.t42 commonsourceibias.t43 gnd.t277 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X206 CSoutput.t137 a_n5644_8799.t58 vdd.t34 vdd.t22 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X207 commonsourceibias.t41 commonsourceibias.t40 gnd.t276 gnd.t275 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X208 outputibias.t3 outputibias.t2 gnd.t40 gnd.t39 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X209 vdd.t93 vdd.t91 vdd.t92 vdd.t73 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X210 a_n1808_13878.t17 a_n2356_n452.t56 vdd.t196 vdd.t195 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X211 vdd.t155 a_n2356_n452.t57 a_n1808_13878.t16 vdd.t154 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X212 gnd.t273 commonsourceibias.t126 CSoutput.t73 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X213 commonsourceibias.t39 commonsourceibias.t38 gnd.t274 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X214 vdd.t90 vdd.t87 vdd.t89 vdd.t88 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X215 a_n2903_n3924.t45 minus.t12 a_n2356_n452.t43 gnd.t356 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X216 gnd.t272 commonsourceibias.t36 commonsourceibias.t37 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X217 diffpairibias.t7 diffpairibias.t6 gnd.t177 gnd.t176 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X218 CSoutput.t72 commonsourceibias.t127 gnd.t271 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X219 commonsourceibias.t35 commonsourceibias.t34 gnd.t270 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X220 CSoutput.t36 a_n5644_8799.t59 vdd.t33 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X221 vdd.t31 a_n5644_8799.t60 CSoutput.t32 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X222 gnd.t113 gnd.t110 gnd.t112 gnd.t111 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X223 a_n2903_n3924.t38 minus.t13 a_n2356_n452.t36 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X224 a_n1986_8322.t6 a_n2356_n452.t58 a_n5644_8799.t5 vdd.t156 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X225 minus.t1 gnd.t107 gnd.t109 gnd.t108 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X226 gnd.t106 gnd.t104 plus.t2 gnd.t105 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X227 gnd.t269 commonsourceibias.t128 CSoutput.t71 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X228 a_n2903_n3924.t42 minus.t14 a_n2356_n452.t40 gnd.t193 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X229 vdd.t165 CSoutput.t159 output.t8 gnd.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X230 vdd.t30 a_n5644_8799.t61 CSoutput.t23 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X231 CSoutput.t38 a_n5644_8799.t62 vdd.t28 vdd.t9 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X232 CSoutput.t70 commonsourceibias.t129 gnd.t268 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X233 gnd.t267 commonsourceibias.t32 commonsourceibias.t33 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X234 vdd.t27 a_n5644_8799.t63 CSoutput.t25 vdd.t18 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X235 vdd.t142 a_n2356_n452.t59 a_n1986_8322.t0 vdd.t141 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X236 gnd.t265 commonsourceibias.t130 CSoutput.t69 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X237 a_n1808_13878.t15 a_n2356_n452.t60 vdd.t144 vdd.t143 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X238 output.t7 CSoutput.t160 vdd.t167 gnd.t7 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X239 gnd.t103 gnd.t100 gnd.t102 gnd.t101 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X240 a_n2903_n3924.t47 diffpairibias.t21 gnd.t363 gnd.t362 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X241 CSoutput.t35 a_n5644_8799.t64 vdd.t26 vdd.t22 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X242 a_n5644_8799.t19 plus.t20 a_n2903_n3924.t11 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X243 a_n2356_n452.t0 minus.t15 a_n2903_n3924.t2 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X244 gnd.t264 commonsourceibias.t50 commonsourceibias.t51 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X245 CSoutput.t0 a_n5644_8799.t65 vdd.t25 vdd.t20 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X246 a_n2903_n3924.t5 minus.t16 a_n2356_n452.t26 gnd.t13 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X247 vdd.t86 vdd.t84 vdd.t85 vdd.t73 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X248 a_n1986_8322.t2 a_n2356_n452.t61 a_n5644_8799.t1 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X249 vdd.t150 a_n2356_n452.t62 a_n1986_8322.t3 vdd.t149 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X250 vdd.t24 a_n5644_8799.t66 CSoutput.t39 vdd.t11 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X251 CSoutput.t15 a_n5644_8799.t67 vdd.t23 vdd.t22 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X252 gnd.t99 gnd.t97 gnd.t98 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X253 output.t1 outputibias.t10 gnd.t36 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X254 a_n2903_n3924.t43 minus.t17 a_n2356_n452.t41 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X255 CSoutput.t68 commonsourceibias.t131 gnd.t263 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X256 gnd.t262 commonsourceibias.t48 commonsourceibias.t49 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X257 gnd.t96 gnd.t94 gnd.t95 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X258 a_n2903_n3924.t44 minus.t18 a_n2356_n452.t42 gnd.t357 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X259 CSoutput.t67 commonsourceibias.t132 gnd.t261 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X260 output.t0 outputibias.t11 gnd.t30 gnd.t29 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X261 vdd.t171 CSoutput.t161 output.t6 gnd.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X262 output.t5 CSoutput.t162 vdd.t164 gnd.t187 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X263 diffpairibias.t5 diffpairibias.t4 gnd.t51 gnd.t50 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X264 vdd.t83 vdd.t80 vdd.t82 vdd.t81 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X265 vdd.t79 vdd.t76 vdd.t78 vdd.t77 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X266 gnd.t93 gnd.t90 gnd.t92 gnd.t91 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X267 a_n1808_13878.t2 a_n2356_n452.t12 a_n2356_n452.t13 vdd.t146 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X268 CSoutput.t66 commonsourceibias.t133 gnd.t259 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X269 gnd.t257 commonsourceibias.t46 commonsourceibias.t47 gnd.t256 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X270 a_n1986_8322.t11 a_n2356_n452.t63 a_n5644_8799.t13 vdd.t182 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X271 gnd.t89 gnd.t87 plus.t1 gnd.t88 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X272 a_n2903_n3924.t41 minus.t19 a_n2356_n452.t39 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X273 gnd.t255 commonsourceibias.t134 CSoutput.t65 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X274 CSoutput.t17 a_n5644_8799.t68 vdd.t21 vdd.t20 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X275 a_n1986_8322.t12 a_n2356_n452.t64 vdd.t184 vdd.t183 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X276 gnd.t254 commonsourceibias.t135 CSoutput.t64 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X277 gnd.t253 commonsourceibias.t136 CSoutput.t63 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 vdd.t188 a_n2356_n452.t65 a_n1808_13878.t14 vdd.t187 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X279 commonsourceibias.t45 commonsourceibias.t44 gnd.t252 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X280 gnd.t250 commonsourceibias.t137 CSoutput.t62 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X281 vdd.t166 CSoutput.t163 output.t4 gnd.t188 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X282 vdd.t75 vdd.t72 vdd.t74 vdd.t73 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X283 commonsourceibias.t61 commonsourceibias.t60 gnd.t249 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X284 a_n1986_8322.t14 a_n2356_n452.t66 a_n5644_8799.t17 vdd.t176 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X285 minus.t0 gnd.t80 gnd.t82 gnd.t81 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X286 gnd.t79 gnd.t77 plus.t0 gnd.t78 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X287 gnd.t76 gnd.t73 gnd.t75 gnd.t74 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X288 a_n2903_n3924.t10 plus.t21 a_n5644_8799.t8 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X289 vdd.t71 vdd.t69 vdd.t70 vdd.t66 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X290 a_n5644_8799.t0 a_n2356_n452.t67 a_n1986_8322.t1 vdd.t146 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X291 a_n1808_13878.t13 a_n2356_n452.t68 vdd.t148 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X292 vdd.t19 a_n5644_8799.t69 CSoutput.t5 vdd.t18 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X293 CSoutput.t8 a_n5644_8799.t70 vdd.t17 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X294 gnd.t247 commonsourceibias.t138 CSoutput.t61 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X295 a_n2356_n452.t30 minus.t20 a_n2903_n3924.t31 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X296 commonsourceibias.t59 commonsourceibias.t58 gnd.t246 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X297 CSoutput.t60 commonsourceibias.t139 gnd.t244 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X298 a_n2356_n452.t1 minus.t21 a_n2903_n3924.t3 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X299 gnd.t72 gnd.t69 gnd.t71 gnd.t70 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X300 gnd.t243 commonsourceibias.t140 CSoutput.t59 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X301 gnd.t241 commonsourceibias.t56 commonsourceibias.t57 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X302 gnd.t68 gnd.t65 gnd.t67 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X303 gnd.t239 commonsourceibias.t54 commonsourceibias.t55 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X304 commonsourceibias.t53 commonsourceibias.t52 gnd.t238 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X305 gnd.t236 commonsourceibias.t141 CSoutput.t58 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X306 CSoutput.t21 a_n5644_8799.t71 vdd.t15 vdd.t9 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X307 a_n1808_13878.t1 a_n2356_n452.t4 a_n2356_n452.t5 vdd.t159 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X308 a_n2903_n3924.t39 minus.t22 a_n2356_n452.t37 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X309 gnd.t235 commonsourceibias.t142 CSoutput.t57 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X310 CSoutput.t56 commonsourceibias.t143 gnd.t233 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X311 gnd.t232 commonsourceibias.t144 CSoutput.t55 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X312 a_n2903_n3924.t0 diffpairibias.t22 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X313 gnd.t64 gnd.t61 gnd.t63 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X314 CSoutput.t54 commonsourceibias.t145 gnd.t199 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X315 CSoutput.t2 a_n5644_8799.t72 vdd.t14 vdd.t7 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X316 CSoutput.t53 commonsourceibias.t146 gnd.t230 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X317 gnd.t229 commonsourceibias.t147 CSoutput.t52 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X318 commonsourceibias.t1 commonsourceibias.t0 gnd.t227 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X319 vdd.t13 a_n5644_8799.t73 CSoutput.t138 vdd.t5 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X320 CSoutput.t164 a_n1986_8322.t8 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X321 diffpairibias.t3 diffpairibias.t2 gnd.t361 gnd.t360 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X322 a_n5644_8799.t12 a_n2356_n452.t69 a_n1986_8322.t10 vdd.t179 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X323 a_n2356_n452.t9 a_n2356_n452.t8 a_n1808_13878.t0 vdd.t176 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X324 gnd.t225 commonsourceibias.t148 CSoutput.t51 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X325 a_n2356_n452.t27 minus.t23 a_n2903_n3924.t6 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X326 vdd.t12 a_n5644_8799.t74 CSoutput.t33 vdd.t11 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X327 gnd.t60 gnd.t57 gnd.t59 gnd.t58 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X328 vdd.t68 vdd.t65 vdd.t67 vdd.t66 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X329 gnd.t224 commonsourceibias.t149 CSoutput.t50 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 diffpairibias.t1 diffpairibias.t0 gnd.t27 gnd.t26 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X331 CSoutput.t49 commonsourceibias.t150 gnd.t222 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X332 gnd.t220 commonsourceibias.t151 CSoutput.t48 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X333 commonsourceibias.t7 commonsourceibias.t6 gnd.t219 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X334 gnd.t218 commonsourceibias.t4 commonsourceibias.t5 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X335 gnd.t216 commonsourceibias.t152 CSoutput.t47 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X336 a_n5644_8799.t23 plus.t22 a_n2903_n3924.t9 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X337 vdd.t181 a_n2356_n452.t70 a_n1808_13878.t12 vdd.t180 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X338 CSoutput.t18 a_n5644_8799.t75 vdd.t10 vdd.t9 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X339 a_n5644_8799.t10 plus.t23 a_n2903_n3924.t8 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X340 a_n2356_n452.t38 minus.t24 a_n2903_n3924.t40 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X341 gnd.t214 commonsourceibias.t153 CSoutput.t46 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X342 gnd.t212 commonsourceibias.t154 CSoutput.t45 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X343 commonsourceibias.t3 commonsourceibias.t2 gnd.t210 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X344 gnd.t56 gnd.t53 gnd.t55 gnd.t54 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X345 vdd.t162 CSoutput.t165 output.t3 gnd.t45 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X346 gnd.t208 commonsourceibias.t155 CSoutput.t44 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X347 CSoutput.t4 a_n5644_8799.t76 vdd.t8 vdd.t7 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X348 gnd.t207 commonsourceibias.t156 CSoutput.t43 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X349 vdd.t6 a_n5644_8799.t77 CSoutput.t13 vdd.t5 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X350 a_n1986_8322.t13 a_n2356_n452.t71 a_n5644_8799.t16 vdd.t186 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X351 CSoutput.t42 commonsourceibias.t157 gnd.t205 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X352 gnd.t203 commonsourceibias.t158 CSoutput.t41 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X353 CSoutput.t40 commonsourceibias.t159 gnd.t201 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X354 a_n2903_n3924.t7 plus.t24 a_n5644_8799.t20 gnd.t356 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X355 outputibias.t1 outputibias.t0 gnd.t191 gnd.t190 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X356 commonsourceibias.t63 commonsourceibias.t62 gnd.t197 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X357 vdd.t4 a_n5644_8799.t78 CSoutput.t10 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X358 CSoutput.t16 a_n5644_8799.t79 vdd.t2 vdd.t1 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X359 a_n2903_n3924.t29 diffpairibias.t23 gnd.t23 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
R0 commonsourceibias.n35 commonsourceibias.t62 223.028
R1 commonsourceibias.n128 commonsourceibias.t129 223.028
R2 commonsourceibias.n307 commonsourceibias.t139 223.028
R3 commonsourceibias.n217 commonsourceibias.t108 223.028
R4 commonsourceibias.n454 commonsourceibias.t46 223.028
R5 commonsourceibias.n395 commonsourceibias.t112 223.028
R6 commonsourceibias.n679 commonsourceibias.t73 223.028
R7 commonsourceibias.n589 commonsourceibias.t99 223.028
R8 commonsourceibias.n99 commonsourceibias.t54 207.983
R9 commonsourceibias.n192 commonsourceibias.t120 207.983
R10 commonsourceibias.n371 commonsourceibias.t147 207.983
R11 commonsourceibias.n281 commonsourceibias.t68 207.983
R12 commonsourceibias.n520 commonsourceibias.t38 207.983
R13 commonsourceibias.n566 commonsourceibias.t93 207.983
R14 commonsourceibias.n745 commonsourceibias.t82 207.983
R15 commonsourceibias.n655 commonsourceibias.t150 207.983
R16 commonsourceibias.n97 commonsourceibias.t20 168.701
R17 commonsourceibias.n91 commonsourceibias.t4 168.701
R18 commonsourceibias.n17 commonsourceibias.t52 168.701
R19 commonsourceibias.n83 commonsourceibias.t14 168.701
R20 commonsourceibias.n77 commonsourceibias.t58 168.701
R21 commonsourceibias.n22 commonsourceibias.t32 168.701
R22 commonsourceibias.n69 commonsourceibias.t6 168.701
R23 commonsourceibias.n63 commonsourceibias.t56 168.701
R24 commonsourceibias.n25 commonsourceibias.t28 168.701
R25 commonsourceibias.n27 commonsourceibias.t48 168.701
R26 commonsourceibias.n29 commonsourceibias.t34 168.701
R27 commonsourceibias.n46 commonsourceibias.t18 168.701
R28 commonsourceibias.n40 commonsourceibias.t60 168.701
R29 commonsourceibias.n34 commonsourceibias.t22 168.701
R30 commonsourceibias.n190 commonsourceibias.t65 168.701
R31 commonsourceibias.n184 commonsourceibias.t126 168.701
R32 commonsourceibias.n5 commonsourceibias.t121 168.701
R33 commonsourceibias.n176 commonsourceibias.t135 168.701
R34 commonsourceibias.n170 commonsourceibias.t117 168.701
R35 commonsourceibias.n10 commonsourceibias.t102 168.701
R36 commonsourceibias.n162 commonsourceibias.t125 168.701
R37 commonsourceibias.n156 commonsourceibias.t119 168.701
R38 commonsourceibias.n118 commonsourceibias.t79 168.701
R39 commonsourceibias.n120 commonsourceibias.t106 168.701
R40 commonsourceibias.n122 commonsourceibias.t96 168.701
R41 commonsourceibias.n139 commonsourceibias.t141 168.701
R42 commonsourceibias.n133 commonsourceibias.t116 168.701
R43 commonsourceibias.n127 commonsourceibias.t152 168.701
R44 commonsourceibias.n306 commonsourceibias.t130 168.701
R45 commonsourceibias.n312 commonsourceibias.t76 168.701
R46 commonsourceibias.n318 commonsourceibias.t149 168.701
R47 commonsourceibias.n301 commonsourceibias.t133 168.701
R48 commonsourceibias.n299 commonsourceibias.t137 168.701
R49 commonsourceibias.n297 commonsourceibias.t64 168.701
R50 commonsourceibias.n335 commonsourceibias.t138 168.701
R51 commonsourceibias.n341 commonsourceibias.t146 168.701
R52 commonsourceibias.n294 commonsourceibias.t118 168.701
R53 commonsourceibias.n349 commonsourceibias.t89 168.701
R54 commonsourceibias.n355 commonsourceibias.t155 168.701
R55 commonsourceibias.n289 commonsourceibias.t124 168.701
R56 commonsourceibias.n363 commonsourceibias.t128 168.701
R57 commonsourceibias.n369 commonsourceibias.t75 168.701
R58 commonsourceibias.n279 commonsourceibias.t159 168.701
R59 commonsourceibias.n273 commonsourceibias.t148 168.701
R60 commonsourceibias.n199 commonsourceibias.t78 168.701
R61 commonsourceibias.n265 commonsourceibias.t158 168.701
R62 commonsourceibias.n259 commonsourceibias.t85 168.701
R63 commonsourceibias.n204 commonsourceibias.t77 168.701
R64 commonsourceibias.n251 commonsourceibias.t157 168.701
R65 commonsourceibias.n245 commonsourceibias.t94 168.701
R66 commonsourceibias.n207 commonsourceibias.t113 168.701
R67 commonsourceibias.n209 commonsourceibias.t156 168.701
R68 commonsourceibias.n211 commonsourceibias.t92 168.701
R69 commonsourceibias.n228 commonsourceibias.t109 168.701
R70 commonsourceibias.n222 commonsourceibias.t105 168.701
R71 commonsourceibias.n216 commonsourceibias.t91 168.701
R72 commonsourceibias.n453 commonsourceibias.t8 168.701
R73 commonsourceibias.n459 commonsourceibias.t24 168.701
R74 commonsourceibias.n465 commonsourceibias.t2 168.701
R75 commonsourceibias.n448 commonsourceibias.t16 168.701
R76 commonsourceibias.n446 commonsourceibias.t26 168.701
R77 commonsourceibias.n444 commonsourceibias.t12 168.701
R78 commonsourceibias.n482 commonsourceibias.t40 168.701
R79 commonsourceibias.n488 commonsourceibias.t50 168.701
R80 commonsourceibias.n490 commonsourceibias.t30 168.701
R81 commonsourceibias.n497 commonsourceibias.t42 168.701
R82 commonsourceibias.n503 commonsourceibias.t0 168.701
R83 commonsourceibias.n505 commonsourceibias.t36 168.701
R84 commonsourceibias.n512 commonsourceibias.t44 168.701
R85 commonsourceibias.n518 commonsourceibias.t10 168.701
R86 commonsourceibias.n564 commonsourceibias.t134 168.701
R87 commonsourceibias.n558 commonsourceibias.t114 168.701
R88 commonsourceibias.n551 commonsourceibias.t95 168.701
R89 commonsourceibias.n549 commonsourceibias.t123 168.701
R90 commonsourceibias.n543 commonsourceibias.t88 168.701
R91 commonsourceibias.n536 commonsourceibias.t74 168.701
R92 commonsourceibias.n534 commonsourceibias.t104 168.701
R93 commonsourceibias.n394 commonsourceibias.t131 168.701
R94 commonsourceibias.n400 commonsourceibias.t84 168.701
R95 commonsourceibias.n406 commonsourceibias.t127 168.701
R96 commonsourceibias.n389 commonsourceibias.t151 168.701
R97 commonsourceibias.n387 commonsourceibias.t83 168.701
R98 commonsourceibias.n385 commonsourceibias.t140 168.701
R99 commonsourceibias.n423 commonsourceibias.t90 168.701
R100 commonsourceibias.n678 commonsourceibias.t145 168.701
R101 commonsourceibias.n684 commonsourceibias.t111 168.701
R102 commonsourceibias.n690 commonsourceibias.t86 168.701
R103 commonsourceibias.n673 commonsourceibias.t153 168.701
R104 commonsourceibias.n671 commonsourceibias.t132 168.701
R105 commonsourceibias.n669 commonsourceibias.t103 168.701
R106 commonsourceibias.n707 commonsourceibias.t69 168.701
R107 commonsourceibias.n713 commonsourceibias.t81 168.701
R108 commonsourceibias.n715 commonsourceibias.t110 168.701
R109 commonsourceibias.n722 commonsourceibias.t115 168.701
R110 commonsourceibias.n728 commonsourceibias.t97 168.701
R111 commonsourceibias.n730 commonsourceibias.t136 168.701
R112 commonsourceibias.n737 commonsourceibias.t122 168.701
R113 commonsourceibias.n743 commonsourceibias.t107 168.701
R114 commonsourceibias.n588 commonsourceibias.t71 168.701
R115 commonsourceibias.n594 commonsourceibias.t87 168.701
R116 commonsourceibias.n600 commonsourceibias.t100 168.701
R117 commonsourceibias.n583 commonsourceibias.t72 168.701
R118 commonsourceibias.n581 commonsourceibias.t80 168.701
R119 commonsourceibias.n579 commonsourceibias.t101 168.701
R120 commonsourceibias.n617 commonsourceibias.t70 168.701
R121 commonsourceibias.n623 commonsourceibias.t144 168.701
R122 commonsourceibias.n625 commonsourceibias.t98 168.701
R123 commonsourceibias.n632 commonsourceibias.t67 168.701
R124 commonsourceibias.n638 commonsourceibias.t143 168.701
R125 commonsourceibias.n640 commonsourceibias.t154 168.701
R126 commonsourceibias.n647 commonsourceibias.t66 168.701
R127 commonsourceibias.n653 commonsourceibias.t142 168.701
R128 commonsourceibias.n36 commonsourceibias.n33 161.3
R129 commonsourceibias.n38 commonsourceibias.n37 161.3
R130 commonsourceibias.n39 commonsourceibias.n32 161.3
R131 commonsourceibias.n42 commonsourceibias.n41 161.3
R132 commonsourceibias.n43 commonsourceibias.n31 161.3
R133 commonsourceibias.n45 commonsourceibias.n44 161.3
R134 commonsourceibias.n47 commonsourceibias.n30 161.3
R135 commonsourceibias.n49 commonsourceibias.n48 161.3
R136 commonsourceibias.n51 commonsourceibias.n50 161.3
R137 commonsourceibias.n52 commonsourceibias.n28 161.3
R138 commonsourceibias.n54 commonsourceibias.n53 161.3
R139 commonsourceibias.n56 commonsourceibias.n55 161.3
R140 commonsourceibias.n57 commonsourceibias.n26 161.3
R141 commonsourceibias.n59 commonsourceibias.n58 161.3
R142 commonsourceibias.n61 commonsourceibias.n60 161.3
R143 commonsourceibias.n62 commonsourceibias.n24 161.3
R144 commonsourceibias.n65 commonsourceibias.n64 161.3
R145 commonsourceibias.n66 commonsourceibias.n23 161.3
R146 commonsourceibias.n68 commonsourceibias.n67 161.3
R147 commonsourceibias.n70 commonsourceibias.n21 161.3
R148 commonsourceibias.n72 commonsourceibias.n71 161.3
R149 commonsourceibias.n73 commonsourceibias.n20 161.3
R150 commonsourceibias.n75 commonsourceibias.n74 161.3
R151 commonsourceibias.n76 commonsourceibias.n19 161.3
R152 commonsourceibias.n79 commonsourceibias.n78 161.3
R153 commonsourceibias.n80 commonsourceibias.n18 161.3
R154 commonsourceibias.n82 commonsourceibias.n81 161.3
R155 commonsourceibias.n84 commonsourceibias.n16 161.3
R156 commonsourceibias.n86 commonsourceibias.n85 161.3
R157 commonsourceibias.n87 commonsourceibias.n15 161.3
R158 commonsourceibias.n89 commonsourceibias.n88 161.3
R159 commonsourceibias.n90 commonsourceibias.n14 161.3
R160 commonsourceibias.n93 commonsourceibias.n92 161.3
R161 commonsourceibias.n94 commonsourceibias.n13 161.3
R162 commonsourceibias.n96 commonsourceibias.n95 161.3
R163 commonsourceibias.n98 commonsourceibias.n12 161.3
R164 commonsourceibias.n129 commonsourceibias.n126 161.3
R165 commonsourceibias.n131 commonsourceibias.n130 161.3
R166 commonsourceibias.n132 commonsourceibias.n125 161.3
R167 commonsourceibias.n135 commonsourceibias.n134 161.3
R168 commonsourceibias.n136 commonsourceibias.n124 161.3
R169 commonsourceibias.n138 commonsourceibias.n137 161.3
R170 commonsourceibias.n140 commonsourceibias.n123 161.3
R171 commonsourceibias.n142 commonsourceibias.n141 161.3
R172 commonsourceibias.n144 commonsourceibias.n143 161.3
R173 commonsourceibias.n145 commonsourceibias.n121 161.3
R174 commonsourceibias.n147 commonsourceibias.n146 161.3
R175 commonsourceibias.n149 commonsourceibias.n148 161.3
R176 commonsourceibias.n150 commonsourceibias.n119 161.3
R177 commonsourceibias.n152 commonsourceibias.n151 161.3
R178 commonsourceibias.n154 commonsourceibias.n153 161.3
R179 commonsourceibias.n155 commonsourceibias.n117 161.3
R180 commonsourceibias.n158 commonsourceibias.n157 161.3
R181 commonsourceibias.n159 commonsourceibias.n11 161.3
R182 commonsourceibias.n161 commonsourceibias.n160 161.3
R183 commonsourceibias.n163 commonsourceibias.n9 161.3
R184 commonsourceibias.n165 commonsourceibias.n164 161.3
R185 commonsourceibias.n166 commonsourceibias.n8 161.3
R186 commonsourceibias.n168 commonsourceibias.n167 161.3
R187 commonsourceibias.n169 commonsourceibias.n7 161.3
R188 commonsourceibias.n172 commonsourceibias.n171 161.3
R189 commonsourceibias.n173 commonsourceibias.n6 161.3
R190 commonsourceibias.n175 commonsourceibias.n174 161.3
R191 commonsourceibias.n177 commonsourceibias.n4 161.3
R192 commonsourceibias.n179 commonsourceibias.n178 161.3
R193 commonsourceibias.n180 commonsourceibias.n3 161.3
R194 commonsourceibias.n182 commonsourceibias.n181 161.3
R195 commonsourceibias.n183 commonsourceibias.n2 161.3
R196 commonsourceibias.n186 commonsourceibias.n185 161.3
R197 commonsourceibias.n187 commonsourceibias.n1 161.3
R198 commonsourceibias.n189 commonsourceibias.n188 161.3
R199 commonsourceibias.n191 commonsourceibias.n0 161.3
R200 commonsourceibias.n370 commonsourceibias.n284 161.3
R201 commonsourceibias.n368 commonsourceibias.n367 161.3
R202 commonsourceibias.n366 commonsourceibias.n285 161.3
R203 commonsourceibias.n365 commonsourceibias.n364 161.3
R204 commonsourceibias.n362 commonsourceibias.n286 161.3
R205 commonsourceibias.n361 commonsourceibias.n360 161.3
R206 commonsourceibias.n359 commonsourceibias.n287 161.3
R207 commonsourceibias.n358 commonsourceibias.n357 161.3
R208 commonsourceibias.n356 commonsourceibias.n288 161.3
R209 commonsourceibias.n354 commonsourceibias.n353 161.3
R210 commonsourceibias.n352 commonsourceibias.n290 161.3
R211 commonsourceibias.n351 commonsourceibias.n350 161.3
R212 commonsourceibias.n348 commonsourceibias.n291 161.3
R213 commonsourceibias.n347 commonsourceibias.n346 161.3
R214 commonsourceibias.n345 commonsourceibias.n292 161.3
R215 commonsourceibias.n344 commonsourceibias.n343 161.3
R216 commonsourceibias.n342 commonsourceibias.n293 161.3
R217 commonsourceibias.n340 commonsourceibias.n339 161.3
R218 commonsourceibias.n338 commonsourceibias.n295 161.3
R219 commonsourceibias.n337 commonsourceibias.n336 161.3
R220 commonsourceibias.n334 commonsourceibias.n296 161.3
R221 commonsourceibias.n333 commonsourceibias.n332 161.3
R222 commonsourceibias.n331 commonsourceibias.n330 161.3
R223 commonsourceibias.n329 commonsourceibias.n298 161.3
R224 commonsourceibias.n328 commonsourceibias.n327 161.3
R225 commonsourceibias.n326 commonsourceibias.n325 161.3
R226 commonsourceibias.n324 commonsourceibias.n300 161.3
R227 commonsourceibias.n323 commonsourceibias.n322 161.3
R228 commonsourceibias.n321 commonsourceibias.n320 161.3
R229 commonsourceibias.n319 commonsourceibias.n302 161.3
R230 commonsourceibias.n317 commonsourceibias.n316 161.3
R231 commonsourceibias.n315 commonsourceibias.n303 161.3
R232 commonsourceibias.n314 commonsourceibias.n313 161.3
R233 commonsourceibias.n311 commonsourceibias.n304 161.3
R234 commonsourceibias.n310 commonsourceibias.n309 161.3
R235 commonsourceibias.n308 commonsourceibias.n305 161.3
R236 commonsourceibias.n218 commonsourceibias.n215 161.3
R237 commonsourceibias.n220 commonsourceibias.n219 161.3
R238 commonsourceibias.n221 commonsourceibias.n214 161.3
R239 commonsourceibias.n224 commonsourceibias.n223 161.3
R240 commonsourceibias.n225 commonsourceibias.n213 161.3
R241 commonsourceibias.n227 commonsourceibias.n226 161.3
R242 commonsourceibias.n229 commonsourceibias.n212 161.3
R243 commonsourceibias.n231 commonsourceibias.n230 161.3
R244 commonsourceibias.n233 commonsourceibias.n232 161.3
R245 commonsourceibias.n234 commonsourceibias.n210 161.3
R246 commonsourceibias.n236 commonsourceibias.n235 161.3
R247 commonsourceibias.n238 commonsourceibias.n237 161.3
R248 commonsourceibias.n239 commonsourceibias.n208 161.3
R249 commonsourceibias.n241 commonsourceibias.n240 161.3
R250 commonsourceibias.n243 commonsourceibias.n242 161.3
R251 commonsourceibias.n244 commonsourceibias.n206 161.3
R252 commonsourceibias.n247 commonsourceibias.n246 161.3
R253 commonsourceibias.n248 commonsourceibias.n205 161.3
R254 commonsourceibias.n250 commonsourceibias.n249 161.3
R255 commonsourceibias.n252 commonsourceibias.n203 161.3
R256 commonsourceibias.n254 commonsourceibias.n253 161.3
R257 commonsourceibias.n255 commonsourceibias.n202 161.3
R258 commonsourceibias.n257 commonsourceibias.n256 161.3
R259 commonsourceibias.n258 commonsourceibias.n201 161.3
R260 commonsourceibias.n261 commonsourceibias.n260 161.3
R261 commonsourceibias.n262 commonsourceibias.n200 161.3
R262 commonsourceibias.n264 commonsourceibias.n263 161.3
R263 commonsourceibias.n266 commonsourceibias.n198 161.3
R264 commonsourceibias.n268 commonsourceibias.n267 161.3
R265 commonsourceibias.n269 commonsourceibias.n197 161.3
R266 commonsourceibias.n271 commonsourceibias.n270 161.3
R267 commonsourceibias.n272 commonsourceibias.n196 161.3
R268 commonsourceibias.n275 commonsourceibias.n274 161.3
R269 commonsourceibias.n276 commonsourceibias.n195 161.3
R270 commonsourceibias.n278 commonsourceibias.n277 161.3
R271 commonsourceibias.n280 commonsourceibias.n194 161.3
R272 commonsourceibias.n519 commonsourceibias.n433 161.3
R273 commonsourceibias.n517 commonsourceibias.n516 161.3
R274 commonsourceibias.n515 commonsourceibias.n434 161.3
R275 commonsourceibias.n514 commonsourceibias.n513 161.3
R276 commonsourceibias.n511 commonsourceibias.n435 161.3
R277 commonsourceibias.n510 commonsourceibias.n509 161.3
R278 commonsourceibias.n508 commonsourceibias.n436 161.3
R279 commonsourceibias.n507 commonsourceibias.n506 161.3
R280 commonsourceibias.n504 commonsourceibias.n437 161.3
R281 commonsourceibias.n502 commonsourceibias.n501 161.3
R282 commonsourceibias.n500 commonsourceibias.n438 161.3
R283 commonsourceibias.n499 commonsourceibias.n498 161.3
R284 commonsourceibias.n496 commonsourceibias.n439 161.3
R285 commonsourceibias.n495 commonsourceibias.n494 161.3
R286 commonsourceibias.n493 commonsourceibias.n440 161.3
R287 commonsourceibias.n492 commonsourceibias.n491 161.3
R288 commonsourceibias.n489 commonsourceibias.n441 161.3
R289 commonsourceibias.n487 commonsourceibias.n486 161.3
R290 commonsourceibias.n485 commonsourceibias.n442 161.3
R291 commonsourceibias.n484 commonsourceibias.n483 161.3
R292 commonsourceibias.n481 commonsourceibias.n443 161.3
R293 commonsourceibias.n480 commonsourceibias.n479 161.3
R294 commonsourceibias.n478 commonsourceibias.n477 161.3
R295 commonsourceibias.n476 commonsourceibias.n445 161.3
R296 commonsourceibias.n475 commonsourceibias.n474 161.3
R297 commonsourceibias.n473 commonsourceibias.n472 161.3
R298 commonsourceibias.n471 commonsourceibias.n447 161.3
R299 commonsourceibias.n470 commonsourceibias.n469 161.3
R300 commonsourceibias.n468 commonsourceibias.n467 161.3
R301 commonsourceibias.n466 commonsourceibias.n449 161.3
R302 commonsourceibias.n464 commonsourceibias.n463 161.3
R303 commonsourceibias.n462 commonsourceibias.n450 161.3
R304 commonsourceibias.n461 commonsourceibias.n460 161.3
R305 commonsourceibias.n458 commonsourceibias.n451 161.3
R306 commonsourceibias.n457 commonsourceibias.n456 161.3
R307 commonsourceibias.n455 commonsourceibias.n452 161.3
R308 commonsourceibias.n425 commonsourceibias.n424 161.3
R309 commonsourceibias.n422 commonsourceibias.n384 161.3
R310 commonsourceibias.n421 commonsourceibias.n420 161.3
R311 commonsourceibias.n419 commonsourceibias.n418 161.3
R312 commonsourceibias.n417 commonsourceibias.n386 161.3
R313 commonsourceibias.n416 commonsourceibias.n415 161.3
R314 commonsourceibias.n414 commonsourceibias.n413 161.3
R315 commonsourceibias.n412 commonsourceibias.n388 161.3
R316 commonsourceibias.n411 commonsourceibias.n410 161.3
R317 commonsourceibias.n409 commonsourceibias.n408 161.3
R318 commonsourceibias.n407 commonsourceibias.n390 161.3
R319 commonsourceibias.n405 commonsourceibias.n404 161.3
R320 commonsourceibias.n403 commonsourceibias.n391 161.3
R321 commonsourceibias.n402 commonsourceibias.n401 161.3
R322 commonsourceibias.n399 commonsourceibias.n392 161.3
R323 commonsourceibias.n398 commonsourceibias.n397 161.3
R324 commonsourceibias.n396 commonsourceibias.n393 161.3
R325 commonsourceibias.n531 commonsourceibias.n383 161.3
R326 commonsourceibias.n565 commonsourceibias.n374 161.3
R327 commonsourceibias.n563 commonsourceibias.n562 161.3
R328 commonsourceibias.n561 commonsourceibias.n375 161.3
R329 commonsourceibias.n560 commonsourceibias.n559 161.3
R330 commonsourceibias.n557 commonsourceibias.n376 161.3
R331 commonsourceibias.n556 commonsourceibias.n555 161.3
R332 commonsourceibias.n554 commonsourceibias.n377 161.3
R333 commonsourceibias.n553 commonsourceibias.n552 161.3
R334 commonsourceibias.n550 commonsourceibias.n378 161.3
R335 commonsourceibias.n548 commonsourceibias.n547 161.3
R336 commonsourceibias.n546 commonsourceibias.n379 161.3
R337 commonsourceibias.n545 commonsourceibias.n544 161.3
R338 commonsourceibias.n542 commonsourceibias.n380 161.3
R339 commonsourceibias.n541 commonsourceibias.n540 161.3
R340 commonsourceibias.n539 commonsourceibias.n381 161.3
R341 commonsourceibias.n538 commonsourceibias.n537 161.3
R342 commonsourceibias.n535 commonsourceibias.n382 161.3
R343 commonsourceibias.n533 commonsourceibias.n532 161.3
R344 commonsourceibias.n744 commonsourceibias.n658 161.3
R345 commonsourceibias.n742 commonsourceibias.n741 161.3
R346 commonsourceibias.n740 commonsourceibias.n659 161.3
R347 commonsourceibias.n739 commonsourceibias.n738 161.3
R348 commonsourceibias.n736 commonsourceibias.n660 161.3
R349 commonsourceibias.n735 commonsourceibias.n734 161.3
R350 commonsourceibias.n733 commonsourceibias.n661 161.3
R351 commonsourceibias.n732 commonsourceibias.n731 161.3
R352 commonsourceibias.n729 commonsourceibias.n662 161.3
R353 commonsourceibias.n727 commonsourceibias.n726 161.3
R354 commonsourceibias.n725 commonsourceibias.n663 161.3
R355 commonsourceibias.n724 commonsourceibias.n723 161.3
R356 commonsourceibias.n721 commonsourceibias.n664 161.3
R357 commonsourceibias.n720 commonsourceibias.n719 161.3
R358 commonsourceibias.n718 commonsourceibias.n665 161.3
R359 commonsourceibias.n717 commonsourceibias.n716 161.3
R360 commonsourceibias.n714 commonsourceibias.n666 161.3
R361 commonsourceibias.n712 commonsourceibias.n711 161.3
R362 commonsourceibias.n710 commonsourceibias.n667 161.3
R363 commonsourceibias.n709 commonsourceibias.n708 161.3
R364 commonsourceibias.n706 commonsourceibias.n668 161.3
R365 commonsourceibias.n705 commonsourceibias.n704 161.3
R366 commonsourceibias.n703 commonsourceibias.n702 161.3
R367 commonsourceibias.n701 commonsourceibias.n670 161.3
R368 commonsourceibias.n700 commonsourceibias.n699 161.3
R369 commonsourceibias.n698 commonsourceibias.n697 161.3
R370 commonsourceibias.n696 commonsourceibias.n672 161.3
R371 commonsourceibias.n695 commonsourceibias.n694 161.3
R372 commonsourceibias.n693 commonsourceibias.n692 161.3
R373 commonsourceibias.n691 commonsourceibias.n674 161.3
R374 commonsourceibias.n689 commonsourceibias.n688 161.3
R375 commonsourceibias.n687 commonsourceibias.n675 161.3
R376 commonsourceibias.n686 commonsourceibias.n685 161.3
R377 commonsourceibias.n683 commonsourceibias.n676 161.3
R378 commonsourceibias.n682 commonsourceibias.n681 161.3
R379 commonsourceibias.n680 commonsourceibias.n677 161.3
R380 commonsourceibias.n654 commonsourceibias.n568 161.3
R381 commonsourceibias.n652 commonsourceibias.n651 161.3
R382 commonsourceibias.n650 commonsourceibias.n569 161.3
R383 commonsourceibias.n649 commonsourceibias.n648 161.3
R384 commonsourceibias.n646 commonsourceibias.n570 161.3
R385 commonsourceibias.n645 commonsourceibias.n644 161.3
R386 commonsourceibias.n643 commonsourceibias.n571 161.3
R387 commonsourceibias.n642 commonsourceibias.n641 161.3
R388 commonsourceibias.n639 commonsourceibias.n572 161.3
R389 commonsourceibias.n637 commonsourceibias.n636 161.3
R390 commonsourceibias.n635 commonsourceibias.n573 161.3
R391 commonsourceibias.n634 commonsourceibias.n633 161.3
R392 commonsourceibias.n631 commonsourceibias.n574 161.3
R393 commonsourceibias.n630 commonsourceibias.n629 161.3
R394 commonsourceibias.n628 commonsourceibias.n575 161.3
R395 commonsourceibias.n627 commonsourceibias.n626 161.3
R396 commonsourceibias.n624 commonsourceibias.n576 161.3
R397 commonsourceibias.n622 commonsourceibias.n621 161.3
R398 commonsourceibias.n620 commonsourceibias.n577 161.3
R399 commonsourceibias.n619 commonsourceibias.n618 161.3
R400 commonsourceibias.n616 commonsourceibias.n578 161.3
R401 commonsourceibias.n615 commonsourceibias.n614 161.3
R402 commonsourceibias.n613 commonsourceibias.n612 161.3
R403 commonsourceibias.n611 commonsourceibias.n580 161.3
R404 commonsourceibias.n610 commonsourceibias.n609 161.3
R405 commonsourceibias.n608 commonsourceibias.n607 161.3
R406 commonsourceibias.n606 commonsourceibias.n582 161.3
R407 commonsourceibias.n605 commonsourceibias.n604 161.3
R408 commonsourceibias.n603 commonsourceibias.n602 161.3
R409 commonsourceibias.n601 commonsourceibias.n584 161.3
R410 commonsourceibias.n599 commonsourceibias.n598 161.3
R411 commonsourceibias.n597 commonsourceibias.n585 161.3
R412 commonsourceibias.n596 commonsourceibias.n595 161.3
R413 commonsourceibias.n593 commonsourceibias.n586 161.3
R414 commonsourceibias.n592 commonsourceibias.n591 161.3
R415 commonsourceibias.n590 commonsourceibias.n587 161.3
R416 commonsourceibias.n111 commonsourceibias.n109 81.5057
R417 commonsourceibias.n428 commonsourceibias.n426 81.5057
R418 commonsourceibias.n111 commonsourceibias.n110 80.9324
R419 commonsourceibias.n113 commonsourceibias.n112 80.9324
R420 commonsourceibias.n115 commonsourceibias.n114 80.9324
R421 commonsourceibias.n108 commonsourceibias.n107 80.9324
R422 commonsourceibias.n106 commonsourceibias.n105 80.9324
R423 commonsourceibias.n104 commonsourceibias.n103 80.9324
R424 commonsourceibias.n102 commonsourceibias.n101 80.9324
R425 commonsourceibias.n523 commonsourceibias.n522 80.9324
R426 commonsourceibias.n525 commonsourceibias.n524 80.9324
R427 commonsourceibias.n527 commonsourceibias.n526 80.9324
R428 commonsourceibias.n529 commonsourceibias.n528 80.9324
R429 commonsourceibias.n432 commonsourceibias.n431 80.9324
R430 commonsourceibias.n430 commonsourceibias.n429 80.9324
R431 commonsourceibias.n428 commonsourceibias.n427 80.9324
R432 commonsourceibias.n100 commonsourceibias.n99 80.6037
R433 commonsourceibias.n193 commonsourceibias.n192 80.6037
R434 commonsourceibias.n372 commonsourceibias.n371 80.6037
R435 commonsourceibias.n282 commonsourceibias.n281 80.6037
R436 commonsourceibias.n521 commonsourceibias.n520 80.6037
R437 commonsourceibias.n567 commonsourceibias.n566 80.6037
R438 commonsourceibias.n746 commonsourceibias.n745 80.6037
R439 commonsourceibias.n656 commonsourceibias.n655 80.6037
R440 commonsourceibias.n85 commonsourceibias.n84 56.5617
R441 commonsourceibias.n71 commonsourceibias.n70 56.5617
R442 commonsourceibias.n62 commonsourceibias.n61 56.5617
R443 commonsourceibias.n48 commonsourceibias.n47 56.5617
R444 commonsourceibias.n178 commonsourceibias.n177 56.5617
R445 commonsourceibias.n164 commonsourceibias.n163 56.5617
R446 commonsourceibias.n155 commonsourceibias.n154 56.5617
R447 commonsourceibias.n141 commonsourceibias.n140 56.5617
R448 commonsourceibias.n320 commonsourceibias.n319 56.5617
R449 commonsourceibias.n334 commonsourceibias.n333 56.5617
R450 commonsourceibias.n343 commonsourceibias.n342 56.5617
R451 commonsourceibias.n357 commonsourceibias.n356 56.5617
R452 commonsourceibias.n267 commonsourceibias.n266 56.5617
R453 commonsourceibias.n253 commonsourceibias.n252 56.5617
R454 commonsourceibias.n244 commonsourceibias.n243 56.5617
R455 commonsourceibias.n230 commonsourceibias.n229 56.5617
R456 commonsourceibias.n467 commonsourceibias.n466 56.5617
R457 commonsourceibias.n481 commonsourceibias.n480 56.5617
R458 commonsourceibias.n491 commonsourceibias.n489 56.5617
R459 commonsourceibias.n506 commonsourceibias.n504 56.5617
R460 commonsourceibias.n552 commonsourceibias.n550 56.5617
R461 commonsourceibias.n537 commonsourceibias.n535 56.5617
R462 commonsourceibias.n408 commonsourceibias.n407 56.5617
R463 commonsourceibias.n422 commonsourceibias.n421 56.5617
R464 commonsourceibias.n692 commonsourceibias.n691 56.5617
R465 commonsourceibias.n706 commonsourceibias.n705 56.5617
R466 commonsourceibias.n716 commonsourceibias.n714 56.5617
R467 commonsourceibias.n731 commonsourceibias.n729 56.5617
R468 commonsourceibias.n602 commonsourceibias.n601 56.5617
R469 commonsourceibias.n616 commonsourceibias.n615 56.5617
R470 commonsourceibias.n626 commonsourceibias.n624 56.5617
R471 commonsourceibias.n641 commonsourceibias.n639 56.5617
R472 commonsourceibias.n76 commonsourceibias.n75 56.0773
R473 commonsourceibias.n57 commonsourceibias.n56 56.0773
R474 commonsourceibias.n169 commonsourceibias.n168 56.0773
R475 commonsourceibias.n150 commonsourceibias.n149 56.0773
R476 commonsourceibias.n329 commonsourceibias.n328 56.0773
R477 commonsourceibias.n348 commonsourceibias.n347 56.0773
R478 commonsourceibias.n258 commonsourceibias.n257 56.0773
R479 commonsourceibias.n239 commonsourceibias.n238 56.0773
R480 commonsourceibias.n476 commonsourceibias.n475 56.0773
R481 commonsourceibias.n496 commonsourceibias.n495 56.0773
R482 commonsourceibias.n542 commonsourceibias.n541 56.0773
R483 commonsourceibias.n417 commonsourceibias.n416 56.0773
R484 commonsourceibias.n701 commonsourceibias.n700 56.0773
R485 commonsourceibias.n721 commonsourceibias.n720 56.0773
R486 commonsourceibias.n611 commonsourceibias.n610 56.0773
R487 commonsourceibias.n631 commonsourceibias.n630 56.0773
R488 commonsourceibias.n99 commonsourceibias.n98 55.3321
R489 commonsourceibias.n192 commonsourceibias.n191 55.3321
R490 commonsourceibias.n371 commonsourceibias.n370 55.3321
R491 commonsourceibias.n281 commonsourceibias.n280 55.3321
R492 commonsourceibias.n520 commonsourceibias.n519 55.3321
R493 commonsourceibias.n566 commonsourceibias.n565 55.3321
R494 commonsourceibias.n745 commonsourceibias.n744 55.3321
R495 commonsourceibias.n655 commonsourceibias.n654 55.3321
R496 commonsourceibias.n90 commonsourceibias.n89 55.1086
R497 commonsourceibias.n41 commonsourceibias.n31 55.1086
R498 commonsourceibias.n183 commonsourceibias.n182 55.1086
R499 commonsourceibias.n134 commonsourceibias.n124 55.1086
R500 commonsourceibias.n313 commonsourceibias.n303 55.1086
R501 commonsourceibias.n362 commonsourceibias.n361 55.1086
R502 commonsourceibias.n272 commonsourceibias.n271 55.1086
R503 commonsourceibias.n223 commonsourceibias.n213 55.1086
R504 commonsourceibias.n460 commonsourceibias.n450 55.1086
R505 commonsourceibias.n511 commonsourceibias.n510 55.1086
R506 commonsourceibias.n557 commonsourceibias.n556 55.1086
R507 commonsourceibias.n401 commonsourceibias.n391 55.1086
R508 commonsourceibias.n685 commonsourceibias.n675 55.1086
R509 commonsourceibias.n736 commonsourceibias.n735 55.1086
R510 commonsourceibias.n595 commonsourceibias.n585 55.1086
R511 commonsourceibias.n646 commonsourceibias.n645 55.1086
R512 commonsourceibias.n35 commonsourceibias.n34 47.4592
R513 commonsourceibias.n128 commonsourceibias.n127 47.4592
R514 commonsourceibias.n307 commonsourceibias.n306 47.4592
R515 commonsourceibias.n217 commonsourceibias.n216 47.4592
R516 commonsourceibias.n454 commonsourceibias.n453 47.4592
R517 commonsourceibias.n395 commonsourceibias.n394 47.4592
R518 commonsourceibias.n679 commonsourceibias.n678 47.4592
R519 commonsourceibias.n589 commonsourceibias.n588 47.4592
R520 commonsourceibias.n308 commonsourceibias.n307 44.0436
R521 commonsourceibias.n455 commonsourceibias.n454 44.0436
R522 commonsourceibias.n396 commonsourceibias.n395 44.0436
R523 commonsourceibias.n680 commonsourceibias.n679 44.0436
R524 commonsourceibias.n590 commonsourceibias.n589 44.0436
R525 commonsourceibias.n36 commonsourceibias.n35 44.0436
R526 commonsourceibias.n129 commonsourceibias.n128 44.0436
R527 commonsourceibias.n218 commonsourceibias.n217 44.0436
R528 commonsourceibias.n92 commonsourceibias.n13 42.5146
R529 commonsourceibias.n39 commonsourceibias.n38 42.5146
R530 commonsourceibias.n185 commonsourceibias.n1 42.5146
R531 commonsourceibias.n132 commonsourceibias.n131 42.5146
R532 commonsourceibias.n311 commonsourceibias.n310 42.5146
R533 commonsourceibias.n364 commonsourceibias.n285 42.5146
R534 commonsourceibias.n274 commonsourceibias.n195 42.5146
R535 commonsourceibias.n221 commonsourceibias.n220 42.5146
R536 commonsourceibias.n458 commonsourceibias.n457 42.5146
R537 commonsourceibias.n513 commonsourceibias.n434 42.5146
R538 commonsourceibias.n559 commonsourceibias.n375 42.5146
R539 commonsourceibias.n399 commonsourceibias.n398 42.5146
R540 commonsourceibias.n683 commonsourceibias.n682 42.5146
R541 commonsourceibias.n738 commonsourceibias.n659 42.5146
R542 commonsourceibias.n593 commonsourceibias.n592 42.5146
R543 commonsourceibias.n648 commonsourceibias.n569 42.5146
R544 commonsourceibias.n78 commonsourceibias.n18 41.5458
R545 commonsourceibias.n53 commonsourceibias.n52 41.5458
R546 commonsourceibias.n171 commonsourceibias.n6 41.5458
R547 commonsourceibias.n146 commonsourceibias.n145 41.5458
R548 commonsourceibias.n325 commonsourceibias.n324 41.5458
R549 commonsourceibias.n350 commonsourceibias.n290 41.5458
R550 commonsourceibias.n260 commonsourceibias.n200 41.5458
R551 commonsourceibias.n235 commonsourceibias.n234 41.5458
R552 commonsourceibias.n472 commonsourceibias.n471 41.5458
R553 commonsourceibias.n498 commonsourceibias.n438 41.5458
R554 commonsourceibias.n544 commonsourceibias.n379 41.5458
R555 commonsourceibias.n413 commonsourceibias.n412 41.5458
R556 commonsourceibias.n697 commonsourceibias.n696 41.5458
R557 commonsourceibias.n723 commonsourceibias.n663 41.5458
R558 commonsourceibias.n607 commonsourceibias.n606 41.5458
R559 commonsourceibias.n633 commonsourceibias.n573 41.5458
R560 commonsourceibias.n68 commonsourceibias.n23 40.577
R561 commonsourceibias.n64 commonsourceibias.n23 40.577
R562 commonsourceibias.n161 commonsourceibias.n11 40.577
R563 commonsourceibias.n157 commonsourceibias.n11 40.577
R564 commonsourceibias.n336 commonsourceibias.n295 40.577
R565 commonsourceibias.n340 commonsourceibias.n295 40.577
R566 commonsourceibias.n250 commonsourceibias.n205 40.577
R567 commonsourceibias.n246 commonsourceibias.n205 40.577
R568 commonsourceibias.n483 commonsourceibias.n442 40.577
R569 commonsourceibias.n487 commonsourceibias.n442 40.577
R570 commonsourceibias.n533 commonsourceibias.n383 40.577
R571 commonsourceibias.n424 commonsourceibias.n383 40.577
R572 commonsourceibias.n708 commonsourceibias.n667 40.577
R573 commonsourceibias.n712 commonsourceibias.n667 40.577
R574 commonsourceibias.n618 commonsourceibias.n577 40.577
R575 commonsourceibias.n622 commonsourceibias.n577 40.577
R576 commonsourceibias.n82 commonsourceibias.n18 39.6083
R577 commonsourceibias.n52 commonsourceibias.n51 39.6083
R578 commonsourceibias.n175 commonsourceibias.n6 39.6083
R579 commonsourceibias.n145 commonsourceibias.n144 39.6083
R580 commonsourceibias.n324 commonsourceibias.n323 39.6083
R581 commonsourceibias.n354 commonsourceibias.n290 39.6083
R582 commonsourceibias.n264 commonsourceibias.n200 39.6083
R583 commonsourceibias.n234 commonsourceibias.n233 39.6083
R584 commonsourceibias.n471 commonsourceibias.n470 39.6083
R585 commonsourceibias.n502 commonsourceibias.n438 39.6083
R586 commonsourceibias.n548 commonsourceibias.n379 39.6083
R587 commonsourceibias.n412 commonsourceibias.n411 39.6083
R588 commonsourceibias.n696 commonsourceibias.n695 39.6083
R589 commonsourceibias.n727 commonsourceibias.n663 39.6083
R590 commonsourceibias.n606 commonsourceibias.n605 39.6083
R591 commonsourceibias.n637 commonsourceibias.n573 39.6083
R592 commonsourceibias.n96 commonsourceibias.n13 38.6395
R593 commonsourceibias.n38 commonsourceibias.n33 38.6395
R594 commonsourceibias.n189 commonsourceibias.n1 38.6395
R595 commonsourceibias.n131 commonsourceibias.n126 38.6395
R596 commonsourceibias.n310 commonsourceibias.n305 38.6395
R597 commonsourceibias.n368 commonsourceibias.n285 38.6395
R598 commonsourceibias.n278 commonsourceibias.n195 38.6395
R599 commonsourceibias.n220 commonsourceibias.n215 38.6395
R600 commonsourceibias.n457 commonsourceibias.n452 38.6395
R601 commonsourceibias.n517 commonsourceibias.n434 38.6395
R602 commonsourceibias.n563 commonsourceibias.n375 38.6395
R603 commonsourceibias.n398 commonsourceibias.n393 38.6395
R604 commonsourceibias.n682 commonsourceibias.n677 38.6395
R605 commonsourceibias.n742 commonsourceibias.n659 38.6395
R606 commonsourceibias.n592 commonsourceibias.n587 38.6395
R607 commonsourceibias.n652 commonsourceibias.n569 38.6395
R608 commonsourceibias.n89 commonsourceibias.n15 26.0455
R609 commonsourceibias.n45 commonsourceibias.n31 26.0455
R610 commonsourceibias.n182 commonsourceibias.n3 26.0455
R611 commonsourceibias.n138 commonsourceibias.n124 26.0455
R612 commonsourceibias.n317 commonsourceibias.n303 26.0455
R613 commonsourceibias.n361 commonsourceibias.n287 26.0455
R614 commonsourceibias.n271 commonsourceibias.n197 26.0455
R615 commonsourceibias.n227 commonsourceibias.n213 26.0455
R616 commonsourceibias.n464 commonsourceibias.n450 26.0455
R617 commonsourceibias.n510 commonsourceibias.n436 26.0455
R618 commonsourceibias.n556 commonsourceibias.n377 26.0455
R619 commonsourceibias.n405 commonsourceibias.n391 26.0455
R620 commonsourceibias.n689 commonsourceibias.n675 26.0455
R621 commonsourceibias.n735 commonsourceibias.n661 26.0455
R622 commonsourceibias.n599 commonsourceibias.n585 26.0455
R623 commonsourceibias.n645 commonsourceibias.n571 26.0455
R624 commonsourceibias.n75 commonsourceibias.n20 25.0767
R625 commonsourceibias.n58 commonsourceibias.n57 25.0767
R626 commonsourceibias.n168 commonsourceibias.n8 25.0767
R627 commonsourceibias.n151 commonsourceibias.n150 25.0767
R628 commonsourceibias.n330 commonsourceibias.n329 25.0767
R629 commonsourceibias.n347 commonsourceibias.n292 25.0767
R630 commonsourceibias.n257 commonsourceibias.n202 25.0767
R631 commonsourceibias.n240 commonsourceibias.n239 25.0767
R632 commonsourceibias.n477 commonsourceibias.n476 25.0767
R633 commonsourceibias.n495 commonsourceibias.n440 25.0767
R634 commonsourceibias.n541 commonsourceibias.n381 25.0767
R635 commonsourceibias.n418 commonsourceibias.n417 25.0767
R636 commonsourceibias.n702 commonsourceibias.n701 25.0767
R637 commonsourceibias.n720 commonsourceibias.n665 25.0767
R638 commonsourceibias.n612 commonsourceibias.n611 25.0767
R639 commonsourceibias.n630 commonsourceibias.n575 25.0767
R640 commonsourceibias.n71 commonsourceibias.n22 24.3464
R641 commonsourceibias.n61 commonsourceibias.n25 24.3464
R642 commonsourceibias.n164 commonsourceibias.n10 24.3464
R643 commonsourceibias.n154 commonsourceibias.n118 24.3464
R644 commonsourceibias.n333 commonsourceibias.n297 24.3464
R645 commonsourceibias.n343 commonsourceibias.n294 24.3464
R646 commonsourceibias.n253 commonsourceibias.n204 24.3464
R647 commonsourceibias.n243 commonsourceibias.n207 24.3464
R648 commonsourceibias.n480 commonsourceibias.n444 24.3464
R649 commonsourceibias.n491 commonsourceibias.n490 24.3464
R650 commonsourceibias.n537 commonsourceibias.n536 24.3464
R651 commonsourceibias.n421 commonsourceibias.n385 24.3464
R652 commonsourceibias.n705 commonsourceibias.n669 24.3464
R653 commonsourceibias.n716 commonsourceibias.n715 24.3464
R654 commonsourceibias.n615 commonsourceibias.n579 24.3464
R655 commonsourceibias.n626 commonsourceibias.n625 24.3464
R656 commonsourceibias.n85 commonsourceibias.n17 23.8546
R657 commonsourceibias.n47 commonsourceibias.n46 23.8546
R658 commonsourceibias.n178 commonsourceibias.n5 23.8546
R659 commonsourceibias.n140 commonsourceibias.n139 23.8546
R660 commonsourceibias.n319 commonsourceibias.n318 23.8546
R661 commonsourceibias.n357 commonsourceibias.n289 23.8546
R662 commonsourceibias.n267 commonsourceibias.n199 23.8546
R663 commonsourceibias.n229 commonsourceibias.n228 23.8546
R664 commonsourceibias.n466 commonsourceibias.n465 23.8546
R665 commonsourceibias.n506 commonsourceibias.n505 23.8546
R666 commonsourceibias.n552 commonsourceibias.n551 23.8546
R667 commonsourceibias.n407 commonsourceibias.n406 23.8546
R668 commonsourceibias.n691 commonsourceibias.n690 23.8546
R669 commonsourceibias.n731 commonsourceibias.n730 23.8546
R670 commonsourceibias.n601 commonsourceibias.n600 23.8546
R671 commonsourceibias.n641 commonsourceibias.n640 23.8546
R672 commonsourceibias.n98 commonsourceibias.n97 17.4607
R673 commonsourceibias.n191 commonsourceibias.n190 17.4607
R674 commonsourceibias.n370 commonsourceibias.n369 17.4607
R675 commonsourceibias.n280 commonsourceibias.n279 17.4607
R676 commonsourceibias.n519 commonsourceibias.n518 17.4607
R677 commonsourceibias.n565 commonsourceibias.n564 17.4607
R678 commonsourceibias.n744 commonsourceibias.n743 17.4607
R679 commonsourceibias.n654 commonsourceibias.n653 17.4607
R680 commonsourceibias.n84 commonsourceibias.n83 16.9689
R681 commonsourceibias.n48 commonsourceibias.n29 16.9689
R682 commonsourceibias.n177 commonsourceibias.n176 16.9689
R683 commonsourceibias.n141 commonsourceibias.n122 16.9689
R684 commonsourceibias.n320 commonsourceibias.n301 16.9689
R685 commonsourceibias.n356 commonsourceibias.n355 16.9689
R686 commonsourceibias.n266 commonsourceibias.n265 16.9689
R687 commonsourceibias.n230 commonsourceibias.n211 16.9689
R688 commonsourceibias.n467 commonsourceibias.n448 16.9689
R689 commonsourceibias.n504 commonsourceibias.n503 16.9689
R690 commonsourceibias.n550 commonsourceibias.n549 16.9689
R691 commonsourceibias.n408 commonsourceibias.n389 16.9689
R692 commonsourceibias.n692 commonsourceibias.n673 16.9689
R693 commonsourceibias.n729 commonsourceibias.n728 16.9689
R694 commonsourceibias.n602 commonsourceibias.n583 16.9689
R695 commonsourceibias.n639 commonsourceibias.n638 16.9689
R696 commonsourceibias.n70 commonsourceibias.n69 16.477
R697 commonsourceibias.n63 commonsourceibias.n62 16.477
R698 commonsourceibias.n163 commonsourceibias.n162 16.477
R699 commonsourceibias.n156 commonsourceibias.n155 16.477
R700 commonsourceibias.n335 commonsourceibias.n334 16.477
R701 commonsourceibias.n342 commonsourceibias.n341 16.477
R702 commonsourceibias.n252 commonsourceibias.n251 16.477
R703 commonsourceibias.n245 commonsourceibias.n244 16.477
R704 commonsourceibias.n482 commonsourceibias.n481 16.477
R705 commonsourceibias.n489 commonsourceibias.n488 16.477
R706 commonsourceibias.n535 commonsourceibias.n534 16.477
R707 commonsourceibias.n423 commonsourceibias.n422 16.477
R708 commonsourceibias.n707 commonsourceibias.n706 16.477
R709 commonsourceibias.n714 commonsourceibias.n713 16.477
R710 commonsourceibias.n617 commonsourceibias.n616 16.477
R711 commonsourceibias.n624 commonsourceibias.n623 16.477
R712 commonsourceibias.n77 commonsourceibias.n76 15.9852
R713 commonsourceibias.n56 commonsourceibias.n27 15.9852
R714 commonsourceibias.n170 commonsourceibias.n169 15.9852
R715 commonsourceibias.n149 commonsourceibias.n120 15.9852
R716 commonsourceibias.n328 commonsourceibias.n299 15.9852
R717 commonsourceibias.n349 commonsourceibias.n348 15.9852
R718 commonsourceibias.n259 commonsourceibias.n258 15.9852
R719 commonsourceibias.n238 commonsourceibias.n209 15.9852
R720 commonsourceibias.n475 commonsourceibias.n446 15.9852
R721 commonsourceibias.n497 commonsourceibias.n496 15.9852
R722 commonsourceibias.n543 commonsourceibias.n542 15.9852
R723 commonsourceibias.n416 commonsourceibias.n387 15.9852
R724 commonsourceibias.n700 commonsourceibias.n671 15.9852
R725 commonsourceibias.n722 commonsourceibias.n721 15.9852
R726 commonsourceibias.n610 commonsourceibias.n581 15.9852
R727 commonsourceibias.n632 commonsourceibias.n631 15.9852
R728 commonsourceibias.n91 commonsourceibias.n90 15.4934
R729 commonsourceibias.n41 commonsourceibias.n40 15.4934
R730 commonsourceibias.n184 commonsourceibias.n183 15.4934
R731 commonsourceibias.n134 commonsourceibias.n133 15.4934
R732 commonsourceibias.n313 commonsourceibias.n312 15.4934
R733 commonsourceibias.n363 commonsourceibias.n362 15.4934
R734 commonsourceibias.n273 commonsourceibias.n272 15.4934
R735 commonsourceibias.n223 commonsourceibias.n222 15.4934
R736 commonsourceibias.n460 commonsourceibias.n459 15.4934
R737 commonsourceibias.n512 commonsourceibias.n511 15.4934
R738 commonsourceibias.n558 commonsourceibias.n557 15.4934
R739 commonsourceibias.n401 commonsourceibias.n400 15.4934
R740 commonsourceibias.n685 commonsourceibias.n684 15.4934
R741 commonsourceibias.n737 commonsourceibias.n736 15.4934
R742 commonsourceibias.n595 commonsourceibias.n594 15.4934
R743 commonsourceibias.n647 commonsourceibias.n646 15.4934
R744 commonsourceibias.n102 commonsourceibias.n100 13.2663
R745 commonsourceibias.n523 commonsourceibias.n521 13.2663
R746 commonsourceibias.n748 commonsourceibias.n373 10.122
R747 commonsourceibias.n159 commonsourceibias.n116 9.50363
R748 commonsourceibias.n531 commonsourceibias.n530 9.50363
R749 commonsourceibias.n92 commonsourceibias.n91 9.09948
R750 commonsourceibias.n40 commonsourceibias.n39 9.09948
R751 commonsourceibias.n185 commonsourceibias.n184 9.09948
R752 commonsourceibias.n133 commonsourceibias.n132 9.09948
R753 commonsourceibias.n312 commonsourceibias.n311 9.09948
R754 commonsourceibias.n364 commonsourceibias.n363 9.09948
R755 commonsourceibias.n274 commonsourceibias.n273 9.09948
R756 commonsourceibias.n222 commonsourceibias.n221 9.09948
R757 commonsourceibias.n459 commonsourceibias.n458 9.09948
R758 commonsourceibias.n513 commonsourceibias.n512 9.09948
R759 commonsourceibias.n559 commonsourceibias.n558 9.09948
R760 commonsourceibias.n400 commonsourceibias.n399 9.09948
R761 commonsourceibias.n684 commonsourceibias.n683 9.09948
R762 commonsourceibias.n738 commonsourceibias.n737 9.09948
R763 commonsourceibias.n594 commonsourceibias.n593 9.09948
R764 commonsourceibias.n648 commonsourceibias.n647 9.09948
R765 commonsourceibias.n283 commonsourceibias.n193 8.79451
R766 commonsourceibias.n657 commonsourceibias.n567 8.79451
R767 commonsourceibias.n78 commonsourceibias.n77 8.60764
R768 commonsourceibias.n53 commonsourceibias.n27 8.60764
R769 commonsourceibias.n171 commonsourceibias.n170 8.60764
R770 commonsourceibias.n146 commonsourceibias.n120 8.60764
R771 commonsourceibias.n325 commonsourceibias.n299 8.60764
R772 commonsourceibias.n350 commonsourceibias.n349 8.60764
R773 commonsourceibias.n260 commonsourceibias.n259 8.60764
R774 commonsourceibias.n235 commonsourceibias.n209 8.60764
R775 commonsourceibias.n472 commonsourceibias.n446 8.60764
R776 commonsourceibias.n498 commonsourceibias.n497 8.60764
R777 commonsourceibias.n544 commonsourceibias.n543 8.60764
R778 commonsourceibias.n413 commonsourceibias.n387 8.60764
R779 commonsourceibias.n697 commonsourceibias.n671 8.60764
R780 commonsourceibias.n723 commonsourceibias.n722 8.60764
R781 commonsourceibias.n607 commonsourceibias.n581 8.60764
R782 commonsourceibias.n633 commonsourceibias.n632 8.60764
R783 commonsourceibias.n748 commonsourceibias.n747 8.46921
R784 commonsourceibias.n69 commonsourceibias.n68 8.11581
R785 commonsourceibias.n64 commonsourceibias.n63 8.11581
R786 commonsourceibias.n162 commonsourceibias.n161 8.11581
R787 commonsourceibias.n157 commonsourceibias.n156 8.11581
R788 commonsourceibias.n336 commonsourceibias.n335 8.11581
R789 commonsourceibias.n341 commonsourceibias.n340 8.11581
R790 commonsourceibias.n251 commonsourceibias.n250 8.11581
R791 commonsourceibias.n246 commonsourceibias.n245 8.11581
R792 commonsourceibias.n483 commonsourceibias.n482 8.11581
R793 commonsourceibias.n488 commonsourceibias.n487 8.11581
R794 commonsourceibias.n534 commonsourceibias.n533 8.11581
R795 commonsourceibias.n424 commonsourceibias.n423 8.11581
R796 commonsourceibias.n708 commonsourceibias.n707 8.11581
R797 commonsourceibias.n713 commonsourceibias.n712 8.11581
R798 commonsourceibias.n618 commonsourceibias.n617 8.11581
R799 commonsourceibias.n623 commonsourceibias.n622 8.11581
R800 commonsourceibias.n83 commonsourceibias.n82 7.62397
R801 commonsourceibias.n51 commonsourceibias.n29 7.62397
R802 commonsourceibias.n176 commonsourceibias.n175 7.62397
R803 commonsourceibias.n144 commonsourceibias.n122 7.62397
R804 commonsourceibias.n323 commonsourceibias.n301 7.62397
R805 commonsourceibias.n355 commonsourceibias.n354 7.62397
R806 commonsourceibias.n265 commonsourceibias.n264 7.62397
R807 commonsourceibias.n233 commonsourceibias.n211 7.62397
R808 commonsourceibias.n470 commonsourceibias.n448 7.62397
R809 commonsourceibias.n503 commonsourceibias.n502 7.62397
R810 commonsourceibias.n549 commonsourceibias.n548 7.62397
R811 commonsourceibias.n411 commonsourceibias.n389 7.62397
R812 commonsourceibias.n695 commonsourceibias.n673 7.62397
R813 commonsourceibias.n728 commonsourceibias.n727 7.62397
R814 commonsourceibias.n605 commonsourceibias.n583 7.62397
R815 commonsourceibias.n638 commonsourceibias.n637 7.62397
R816 commonsourceibias.n97 commonsourceibias.n96 7.13213
R817 commonsourceibias.n34 commonsourceibias.n33 7.13213
R818 commonsourceibias.n190 commonsourceibias.n189 7.13213
R819 commonsourceibias.n127 commonsourceibias.n126 7.13213
R820 commonsourceibias.n306 commonsourceibias.n305 7.13213
R821 commonsourceibias.n369 commonsourceibias.n368 7.13213
R822 commonsourceibias.n279 commonsourceibias.n278 7.13213
R823 commonsourceibias.n216 commonsourceibias.n215 7.13213
R824 commonsourceibias.n453 commonsourceibias.n452 7.13213
R825 commonsourceibias.n518 commonsourceibias.n517 7.13213
R826 commonsourceibias.n564 commonsourceibias.n563 7.13213
R827 commonsourceibias.n394 commonsourceibias.n393 7.13213
R828 commonsourceibias.n678 commonsourceibias.n677 7.13213
R829 commonsourceibias.n743 commonsourceibias.n742 7.13213
R830 commonsourceibias.n588 commonsourceibias.n587 7.13213
R831 commonsourceibias.n653 commonsourceibias.n652 7.13213
R832 commonsourceibias.n373 commonsourceibias.n372 5.06534
R833 commonsourceibias.n283 commonsourceibias.n282 5.06534
R834 commonsourceibias.n747 commonsourceibias.n746 5.06534
R835 commonsourceibias.n657 commonsourceibias.n656 5.06534
R836 commonsourceibias commonsourceibias.n748 4.04308
R837 commonsourceibias.n373 commonsourceibias.n283 3.72967
R838 commonsourceibias.n747 commonsourceibias.n657 3.72967
R839 commonsourceibias.n109 commonsourceibias.t23 2.82907
R840 commonsourceibias.n109 commonsourceibias.t63 2.82907
R841 commonsourceibias.n110 commonsourceibias.t19 2.82907
R842 commonsourceibias.n110 commonsourceibias.t61 2.82907
R843 commonsourceibias.n112 commonsourceibias.t49 2.82907
R844 commonsourceibias.n112 commonsourceibias.t35 2.82907
R845 commonsourceibias.n114 commonsourceibias.t57 2.82907
R846 commonsourceibias.n114 commonsourceibias.t29 2.82907
R847 commonsourceibias.n107 commonsourceibias.t33 2.82907
R848 commonsourceibias.n107 commonsourceibias.t7 2.82907
R849 commonsourceibias.n105 commonsourceibias.t15 2.82907
R850 commonsourceibias.n105 commonsourceibias.t59 2.82907
R851 commonsourceibias.n103 commonsourceibias.t5 2.82907
R852 commonsourceibias.n103 commonsourceibias.t53 2.82907
R853 commonsourceibias.n101 commonsourceibias.t55 2.82907
R854 commonsourceibias.n101 commonsourceibias.t21 2.82907
R855 commonsourceibias.n522 commonsourceibias.t11 2.82907
R856 commonsourceibias.n522 commonsourceibias.t39 2.82907
R857 commonsourceibias.n524 commonsourceibias.t37 2.82907
R858 commonsourceibias.n524 commonsourceibias.t45 2.82907
R859 commonsourceibias.n526 commonsourceibias.t43 2.82907
R860 commonsourceibias.n526 commonsourceibias.t1 2.82907
R861 commonsourceibias.n528 commonsourceibias.t51 2.82907
R862 commonsourceibias.n528 commonsourceibias.t31 2.82907
R863 commonsourceibias.n431 commonsourceibias.t13 2.82907
R864 commonsourceibias.n431 commonsourceibias.t41 2.82907
R865 commonsourceibias.n429 commonsourceibias.t17 2.82907
R866 commonsourceibias.n429 commonsourceibias.t27 2.82907
R867 commonsourceibias.n427 commonsourceibias.t25 2.82907
R868 commonsourceibias.n427 commonsourceibias.t3 2.82907
R869 commonsourceibias.n426 commonsourceibias.t47 2.82907
R870 commonsourceibias.n426 commonsourceibias.t9 2.82907
R871 commonsourceibias.n17 commonsourceibias.n15 0.738255
R872 commonsourceibias.n46 commonsourceibias.n45 0.738255
R873 commonsourceibias.n5 commonsourceibias.n3 0.738255
R874 commonsourceibias.n139 commonsourceibias.n138 0.738255
R875 commonsourceibias.n318 commonsourceibias.n317 0.738255
R876 commonsourceibias.n289 commonsourceibias.n287 0.738255
R877 commonsourceibias.n199 commonsourceibias.n197 0.738255
R878 commonsourceibias.n228 commonsourceibias.n227 0.738255
R879 commonsourceibias.n465 commonsourceibias.n464 0.738255
R880 commonsourceibias.n505 commonsourceibias.n436 0.738255
R881 commonsourceibias.n551 commonsourceibias.n377 0.738255
R882 commonsourceibias.n406 commonsourceibias.n405 0.738255
R883 commonsourceibias.n690 commonsourceibias.n689 0.738255
R884 commonsourceibias.n730 commonsourceibias.n661 0.738255
R885 commonsourceibias.n600 commonsourceibias.n599 0.738255
R886 commonsourceibias.n640 commonsourceibias.n571 0.738255
R887 commonsourceibias.n104 commonsourceibias.n102 0.573776
R888 commonsourceibias.n106 commonsourceibias.n104 0.573776
R889 commonsourceibias.n108 commonsourceibias.n106 0.573776
R890 commonsourceibias.n115 commonsourceibias.n113 0.573776
R891 commonsourceibias.n113 commonsourceibias.n111 0.573776
R892 commonsourceibias.n430 commonsourceibias.n428 0.573776
R893 commonsourceibias.n432 commonsourceibias.n430 0.573776
R894 commonsourceibias.n529 commonsourceibias.n527 0.573776
R895 commonsourceibias.n527 commonsourceibias.n525 0.573776
R896 commonsourceibias.n525 commonsourceibias.n523 0.573776
R897 commonsourceibias.n116 commonsourceibias.n108 0.287138
R898 commonsourceibias.n116 commonsourceibias.n115 0.287138
R899 commonsourceibias.n530 commonsourceibias.n432 0.287138
R900 commonsourceibias.n530 commonsourceibias.n529 0.287138
R901 commonsourceibias.n100 commonsourceibias.n12 0.285035
R902 commonsourceibias.n193 commonsourceibias.n0 0.285035
R903 commonsourceibias.n372 commonsourceibias.n284 0.285035
R904 commonsourceibias.n282 commonsourceibias.n194 0.285035
R905 commonsourceibias.n521 commonsourceibias.n433 0.285035
R906 commonsourceibias.n567 commonsourceibias.n374 0.285035
R907 commonsourceibias.n746 commonsourceibias.n658 0.285035
R908 commonsourceibias.n656 commonsourceibias.n568 0.285035
R909 commonsourceibias.n22 commonsourceibias.n20 0.246418
R910 commonsourceibias.n58 commonsourceibias.n25 0.246418
R911 commonsourceibias.n10 commonsourceibias.n8 0.246418
R912 commonsourceibias.n151 commonsourceibias.n118 0.246418
R913 commonsourceibias.n330 commonsourceibias.n297 0.246418
R914 commonsourceibias.n294 commonsourceibias.n292 0.246418
R915 commonsourceibias.n204 commonsourceibias.n202 0.246418
R916 commonsourceibias.n240 commonsourceibias.n207 0.246418
R917 commonsourceibias.n477 commonsourceibias.n444 0.246418
R918 commonsourceibias.n490 commonsourceibias.n440 0.246418
R919 commonsourceibias.n536 commonsourceibias.n381 0.246418
R920 commonsourceibias.n418 commonsourceibias.n385 0.246418
R921 commonsourceibias.n702 commonsourceibias.n669 0.246418
R922 commonsourceibias.n715 commonsourceibias.n665 0.246418
R923 commonsourceibias.n612 commonsourceibias.n579 0.246418
R924 commonsourceibias.n625 commonsourceibias.n575 0.246418
R925 commonsourceibias.n95 commonsourceibias.n12 0.189894
R926 commonsourceibias.n95 commonsourceibias.n94 0.189894
R927 commonsourceibias.n94 commonsourceibias.n93 0.189894
R928 commonsourceibias.n93 commonsourceibias.n14 0.189894
R929 commonsourceibias.n88 commonsourceibias.n14 0.189894
R930 commonsourceibias.n88 commonsourceibias.n87 0.189894
R931 commonsourceibias.n87 commonsourceibias.n86 0.189894
R932 commonsourceibias.n86 commonsourceibias.n16 0.189894
R933 commonsourceibias.n81 commonsourceibias.n16 0.189894
R934 commonsourceibias.n81 commonsourceibias.n80 0.189894
R935 commonsourceibias.n80 commonsourceibias.n79 0.189894
R936 commonsourceibias.n79 commonsourceibias.n19 0.189894
R937 commonsourceibias.n74 commonsourceibias.n19 0.189894
R938 commonsourceibias.n74 commonsourceibias.n73 0.189894
R939 commonsourceibias.n73 commonsourceibias.n72 0.189894
R940 commonsourceibias.n72 commonsourceibias.n21 0.189894
R941 commonsourceibias.n67 commonsourceibias.n21 0.189894
R942 commonsourceibias.n67 commonsourceibias.n66 0.189894
R943 commonsourceibias.n66 commonsourceibias.n65 0.189894
R944 commonsourceibias.n65 commonsourceibias.n24 0.189894
R945 commonsourceibias.n60 commonsourceibias.n24 0.189894
R946 commonsourceibias.n60 commonsourceibias.n59 0.189894
R947 commonsourceibias.n59 commonsourceibias.n26 0.189894
R948 commonsourceibias.n55 commonsourceibias.n26 0.189894
R949 commonsourceibias.n55 commonsourceibias.n54 0.189894
R950 commonsourceibias.n54 commonsourceibias.n28 0.189894
R951 commonsourceibias.n50 commonsourceibias.n28 0.189894
R952 commonsourceibias.n50 commonsourceibias.n49 0.189894
R953 commonsourceibias.n49 commonsourceibias.n30 0.189894
R954 commonsourceibias.n44 commonsourceibias.n30 0.189894
R955 commonsourceibias.n44 commonsourceibias.n43 0.189894
R956 commonsourceibias.n43 commonsourceibias.n42 0.189894
R957 commonsourceibias.n42 commonsourceibias.n32 0.189894
R958 commonsourceibias.n37 commonsourceibias.n32 0.189894
R959 commonsourceibias.n37 commonsourceibias.n36 0.189894
R960 commonsourceibias.n158 commonsourceibias.n117 0.189894
R961 commonsourceibias.n153 commonsourceibias.n117 0.189894
R962 commonsourceibias.n153 commonsourceibias.n152 0.189894
R963 commonsourceibias.n152 commonsourceibias.n119 0.189894
R964 commonsourceibias.n148 commonsourceibias.n119 0.189894
R965 commonsourceibias.n148 commonsourceibias.n147 0.189894
R966 commonsourceibias.n147 commonsourceibias.n121 0.189894
R967 commonsourceibias.n143 commonsourceibias.n121 0.189894
R968 commonsourceibias.n143 commonsourceibias.n142 0.189894
R969 commonsourceibias.n142 commonsourceibias.n123 0.189894
R970 commonsourceibias.n137 commonsourceibias.n123 0.189894
R971 commonsourceibias.n137 commonsourceibias.n136 0.189894
R972 commonsourceibias.n136 commonsourceibias.n135 0.189894
R973 commonsourceibias.n135 commonsourceibias.n125 0.189894
R974 commonsourceibias.n130 commonsourceibias.n125 0.189894
R975 commonsourceibias.n130 commonsourceibias.n129 0.189894
R976 commonsourceibias.n188 commonsourceibias.n0 0.189894
R977 commonsourceibias.n188 commonsourceibias.n187 0.189894
R978 commonsourceibias.n187 commonsourceibias.n186 0.189894
R979 commonsourceibias.n186 commonsourceibias.n2 0.189894
R980 commonsourceibias.n181 commonsourceibias.n2 0.189894
R981 commonsourceibias.n181 commonsourceibias.n180 0.189894
R982 commonsourceibias.n180 commonsourceibias.n179 0.189894
R983 commonsourceibias.n179 commonsourceibias.n4 0.189894
R984 commonsourceibias.n174 commonsourceibias.n4 0.189894
R985 commonsourceibias.n174 commonsourceibias.n173 0.189894
R986 commonsourceibias.n173 commonsourceibias.n172 0.189894
R987 commonsourceibias.n172 commonsourceibias.n7 0.189894
R988 commonsourceibias.n167 commonsourceibias.n7 0.189894
R989 commonsourceibias.n167 commonsourceibias.n166 0.189894
R990 commonsourceibias.n166 commonsourceibias.n165 0.189894
R991 commonsourceibias.n165 commonsourceibias.n9 0.189894
R992 commonsourceibias.n160 commonsourceibias.n9 0.189894
R993 commonsourceibias.n367 commonsourceibias.n284 0.189894
R994 commonsourceibias.n367 commonsourceibias.n366 0.189894
R995 commonsourceibias.n366 commonsourceibias.n365 0.189894
R996 commonsourceibias.n365 commonsourceibias.n286 0.189894
R997 commonsourceibias.n360 commonsourceibias.n286 0.189894
R998 commonsourceibias.n360 commonsourceibias.n359 0.189894
R999 commonsourceibias.n359 commonsourceibias.n358 0.189894
R1000 commonsourceibias.n358 commonsourceibias.n288 0.189894
R1001 commonsourceibias.n353 commonsourceibias.n288 0.189894
R1002 commonsourceibias.n353 commonsourceibias.n352 0.189894
R1003 commonsourceibias.n352 commonsourceibias.n351 0.189894
R1004 commonsourceibias.n351 commonsourceibias.n291 0.189894
R1005 commonsourceibias.n346 commonsourceibias.n291 0.189894
R1006 commonsourceibias.n346 commonsourceibias.n345 0.189894
R1007 commonsourceibias.n345 commonsourceibias.n344 0.189894
R1008 commonsourceibias.n344 commonsourceibias.n293 0.189894
R1009 commonsourceibias.n339 commonsourceibias.n293 0.189894
R1010 commonsourceibias.n339 commonsourceibias.n338 0.189894
R1011 commonsourceibias.n338 commonsourceibias.n337 0.189894
R1012 commonsourceibias.n337 commonsourceibias.n296 0.189894
R1013 commonsourceibias.n332 commonsourceibias.n296 0.189894
R1014 commonsourceibias.n332 commonsourceibias.n331 0.189894
R1015 commonsourceibias.n331 commonsourceibias.n298 0.189894
R1016 commonsourceibias.n327 commonsourceibias.n298 0.189894
R1017 commonsourceibias.n327 commonsourceibias.n326 0.189894
R1018 commonsourceibias.n326 commonsourceibias.n300 0.189894
R1019 commonsourceibias.n322 commonsourceibias.n300 0.189894
R1020 commonsourceibias.n322 commonsourceibias.n321 0.189894
R1021 commonsourceibias.n321 commonsourceibias.n302 0.189894
R1022 commonsourceibias.n316 commonsourceibias.n302 0.189894
R1023 commonsourceibias.n316 commonsourceibias.n315 0.189894
R1024 commonsourceibias.n315 commonsourceibias.n314 0.189894
R1025 commonsourceibias.n314 commonsourceibias.n304 0.189894
R1026 commonsourceibias.n309 commonsourceibias.n304 0.189894
R1027 commonsourceibias.n309 commonsourceibias.n308 0.189894
R1028 commonsourceibias.n277 commonsourceibias.n194 0.189894
R1029 commonsourceibias.n277 commonsourceibias.n276 0.189894
R1030 commonsourceibias.n276 commonsourceibias.n275 0.189894
R1031 commonsourceibias.n275 commonsourceibias.n196 0.189894
R1032 commonsourceibias.n270 commonsourceibias.n196 0.189894
R1033 commonsourceibias.n270 commonsourceibias.n269 0.189894
R1034 commonsourceibias.n269 commonsourceibias.n268 0.189894
R1035 commonsourceibias.n268 commonsourceibias.n198 0.189894
R1036 commonsourceibias.n263 commonsourceibias.n198 0.189894
R1037 commonsourceibias.n263 commonsourceibias.n262 0.189894
R1038 commonsourceibias.n262 commonsourceibias.n261 0.189894
R1039 commonsourceibias.n261 commonsourceibias.n201 0.189894
R1040 commonsourceibias.n256 commonsourceibias.n201 0.189894
R1041 commonsourceibias.n256 commonsourceibias.n255 0.189894
R1042 commonsourceibias.n255 commonsourceibias.n254 0.189894
R1043 commonsourceibias.n254 commonsourceibias.n203 0.189894
R1044 commonsourceibias.n249 commonsourceibias.n203 0.189894
R1045 commonsourceibias.n249 commonsourceibias.n248 0.189894
R1046 commonsourceibias.n248 commonsourceibias.n247 0.189894
R1047 commonsourceibias.n247 commonsourceibias.n206 0.189894
R1048 commonsourceibias.n242 commonsourceibias.n206 0.189894
R1049 commonsourceibias.n242 commonsourceibias.n241 0.189894
R1050 commonsourceibias.n241 commonsourceibias.n208 0.189894
R1051 commonsourceibias.n237 commonsourceibias.n208 0.189894
R1052 commonsourceibias.n237 commonsourceibias.n236 0.189894
R1053 commonsourceibias.n236 commonsourceibias.n210 0.189894
R1054 commonsourceibias.n232 commonsourceibias.n210 0.189894
R1055 commonsourceibias.n232 commonsourceibias.n231 0.189894
R1056 commonsourceibias.n231 commonsourceibias.n212 0.189894
R1057 commonsourceibias.n226 commonsourceibias.n212 0.189894
R1058 commonsourceibias.n226 commonsourceibias.n225 0.189894
R1059 commonsourceibias.n225 commonsourceibias.n224 0.189894
R1060 commonsourceibias.n224 commonsourceibias.n214 0.189894
R1061 commonsourceibias.n219 commonsourceibias.n214 0.189894
R1062 commonsourceibias.n219 commonsourceibias.n218 0.189894
R1063 commonsourceibias.n456 commonsourceibias.n455 0.189894
R1064 commonsourceibias.n456 commonsourceibias.n451 0.189894
R1065 commonsourceibias.n461 commonsourceibias.n451 0.189894
R1066 commonsourceibias.n462 commonsourceibias.n461 0.189894
R1067 commonsourceibias.n463 commonsourceibias.n462 0.189894
R1068 commonsourceibias.n463 commonsourceibias.n449 0.189894
R1069 commonsourceibias.n468 commonsourceibias.n449 0.189894
R1070 commonsourceibias.n469 commonsourceibias.n468 0.189894
R1071 commonsourceibias.n469 commonsourceibias.n447 0.189894
R1072 commonsourceibias.n473 commonsourceibias.n447 0.189894
R1073 commonsourceibias.n474 commonsourceibias.n473 0.189894
R1074 commonsourceibias.n474 commonsourceibias.n445 0.189894
R1075 commonsourceibias.n478 commonsourceibias.n445 0.189894
R1076 commonsourceibias.n479 commonsourceibias.n478 0.189894
R1077 commonsourceibias.n479 commonsourceibias.n443 0.189894
R1078 commonsourceibias.n484 commonsourceibias.n443 0.189894
R1079 commonsourceibias.n485 commonsourceibias.n484 0.189894
R1080 commonsourceibias.n486 commonsourceibias.n485 0.189894
R1081 commonsourceibias.n486 commonsourceibias.n441 0.189894
R1082 commonsourceibias.n492 commonsourceibias.n441 0.189894
R1083 commonsourceibias.n493 commonsourceibias.n492 0.189894
R1084 commonsourceibias.n494 commonsourceibias.n493 0.189894
R1085 commonsourceibias.n494 commonsourceibias.n439 0.189894
R1086 commonsourceibias.n499 commonsourceibias.n439 0.189894
R1087 commonsourceibias.n500 commonsourceibias.n499 0.189894
R1088 commonsourceibias.n501 commonsourceibias.n500 0.189894
R1089 commonsourceibias.n501 commonsourceibias.n437 0.189894
R1090 commonsourceibias.n507 commonsourceibias.n437 0.189894
R1091 commonsourceibias.n508 commonsourceibias.n507 0.189894
R1092 commonsourceibias.n509 commonsourceibias.n508 0.189894
R1093 commonsourceibias.n509 commonsourceibias.n435 0.189894
R1094 commonsourceibias.n514 commonsourceibias.n435 0.189894
R1095 commonsourceibias.n515 commonsourceibias.n514 0.189894
R1096 commonsourceibias.n516 commonsourceibias.n515 0.189894
R1097 commonsourceibias.n516 commonsourceibias.n433 0.189894
R1098 commonsourceibias.n397 commonsourceibias.n396 0.189894
R1099 commonsourceibias.n397 commonsourceibias.n392 0.189894
R1100 commonsourceibias.n402 commonsourceibias.n392 0.189894
R1101 commonsourceibias.n403 commonsourceibias.n402 0.189894
R1102 commonsourceibias.n404 commonsourceibias.n403 0.189894
R1103 commonsourceibias.n404 commonsourceibias.n390 0.189894
R1104 commonsourceibias.n409 commonsourceibias.n390 0.189894
R1105 commonsourceibias.n410 commonsourceibias.n409 0.189894
R1106 commonsourceibias.n410 commonsourceibias.n388 0.189894
R1107 commonsourceibias.n414 commonsourceibias.n388 0.189894
R1108 commonsourceibias.n415 commonsourceibias.n414 0.189894
R1109 commonsourceibias.n415 commonsourceibias.n386 0.189894
R1110 commonsourceibias.n419 commonsourceibias.n386 0.189894
R1111 commonsourceibias.n420 commonsourceibias.n419 0.189894
R1112 commonsourceibias.n420 commonsourceibias.n384 0.189894
R1113 commonsourceibias.n425 commonsourceibias.n384 0.189894
R1114 commonsourceibias.n532 commonsourceibias.n382 0.189894
R1115 commonsourceibias.n538 commonsourceibias.n382 0.189894
R1116 commonsourceibias.n539 commonsourceibias.n538 0.189894
R1117 commonsourceibias.n540 commonsourceibias.n539 0.189894
R1118 commonsourceibias.n540 commonsourceibias.n380 0.189894
R1119 commonsourceibias.n545 commonsourceibias.n380 0.189894
R1120 commonsourceibias.n546 commonsourceibias.n545 0.189894
R1121 commonsourceibias.n547 commonsourceibias.n546 0.189894
R1122 commonsourceibias.n547 commonsourceibias.n378 0.189894
R1123 commonsourceibias.n553 commonsourceibias.n378 0.189894
R1124 commonsourceibias.n554 commonsourceibias.n553 0.189894
R1125 commonsourceibias.n555 commonsourceibias.n554 0.189894
R1126 commonsourceibias.n555 commonsourceibias.n376 0.189894
R1127 commonsourceibias.n560 commonsourceibias.n376 0.189894
R1128 commonsourceibias.n561 commonsourceibias.n560 0.189894
R1129 commonsourceibias.n562 commonsourceibias.n561 0.189894
R1130 commonsourceibias.n562 commonsourceibias.n374 0.189894
R1131 commonsourceibias.n681 commonsourceibias.n680 0.189894
R1132 commonsourceibias.n681 commonsourceibias.n676 0.189894
R1133 commonsourceibias.n686 commonsourceibias.n676 0.189894
R1134 commonsourceibias.n687 commonsourceibias.n686 0.189894
R1135 commonsourceibias.n688 commonsourceibias.n687 0.189894
R1136 commonsourceibias.n688 commonsourceibias.n674 0.189894
R1137 commonsourceibias.n693 commonsourceibias.n674 0.189894
R1138 commonsourceibias.n694 commonsourceibias.n693 0.189894
R1139 commonsourceibias.n694 commonsourceibias.n672 0.189894
R1140 commonsourceibias.n698 commonsourceibias.n672 0.189894
R1141 commonsourceibias.n699 commonsourceibias.n698 0.189894
R1142 commonsourceibias.n699 commonsourceibias.n670 0.189894
R1143 commonsourceibias.n703 commonsourceibias.n670 0.189894
R1144 commonsourceibias.n704 commonsourceibias.n703 0.189894
R1145 commonsourceibias.n704 commonsourceibias.n668 0.189894
R1146 commonsourceibias.n709 commonsourceibias.n668 0.189894
R1147 commonsourceibias.n710 commonsourceibias.n709 0.189894
R1148 commonsourceibias.n711 commonsourceibias.n710 0.189894
R1149 commonsourceibias.n711 commonsourceibias.n666 0.189894
R1150 commonsourceibias.n717 commonsourceibias.n666 0.189894
R1151 commonsourceibias.n718 commonsourceibias.n717 0.189894
R1152 commonsourceibias.n719 commonsourceibias.n718 0.189894
R1153 commonsourceibias.n719 commonsourceibias.n664 0.189894
R1154 commonsourceibias.n724 commonsourceibias.n664 0.189894
R1155 commonsourceibias.n725 commonsourceibias.n724 0.189894
R1156 commonsourceibias.n726 commonsourceibias.n725 0.189894
R1157 commonsourceibias.n726 commonsourceibias.n662 0.189894
R1158 commonsourceibias.n732 commonsourceibias.n662 0.189894
R1159 commonsourceibias.n733 commonsourceibias.n732 0.189894
R1160 commonsourceibias.n734 commonsourceibias.n733 0.189894
R1161 commonsourceibias.n734 commonsourceibias.n660 0.189894
R1162 commonsourceibias.n739 commonsourceibias.n660 0.189894
R1163 commonsourceibias.n740 commonsourceibias.n739 0.189894
R1164 commonsourceibias.n741 commonsourceibias.n740 0.189894
R1165 commonsourceibias.n741 commonsourceibias.n658 0.189894
R1166 commonsourceibias.n591 commonsourceibias.n590 0.189894
R1167 commonsourceibias.n591 commonsourceibias.n586 0.189894
R1168 commonsourceibias.n596 commonsourceibias.n586 0.189894
R1169 commonsourceibias.n597 commonsourceibias.n596 0.189894
R1170 commonsourceibias.n598 commonsourceibias.n597 0.189894
R1171 commonsourceibias.n598 commonsourceibias.n584 0.189894
R1172 commonsourceibias.n603 commonsourceibias.n584 0.189894
R1173 commonsourceibias.n604 commonsourceibias.n603 0.189894
R1174 commonsourceibias.n604 commonsourceibias.n582 0.189894
R1175 commonsourceibias.n608 commonsourceibias.n582 0.189894
R1176 commonsourceibias.n609 commonsourceibias.n608 0.189894
R1177 commonsourceibias.n609 commonsourceibias.n580 0.189894
R1178 commonsourceibias.n613 commonsourceibias.n580 0.189894
R1179 commonsourceibias.n614 commonsourceibias.n613 0.189894
R1180 commonsourceibias.n614 commonsourceibias.n578 0.189894
R1181 commonsourceibias.n619 commonsourceibias.n578 0.189894
R1182 commonsourceibias.n620 commonsourceibias.n619 0.189894
R1183 commonsourceibias.n621 commonsourceibias.n620 0.189894
R1184 commonsourceibias.n621 commonsourceibias.n576 0.189894
R1185 commonsourceibias.n627 commonsourceibias.n576 0.189894
R1186 commonsourceibias.n628 commonsourceibias.n627 0.189894
R1187 commonsourceibias.n629 commonsourceibias.n628 0.189894
R1188 commonsourceibias.n629 commonsourceibias.n574 0.189894
R1189 commonsourceibias.n634 commonsourceibias.n574 0.189894
R1190 commonsourceibias.n635 commonsourceibias.n634 0.189894
R1191 commonsourceibias.n636 commonsourceibias.n635 0.189894
R1192 commonsourceibias.n636 commonsourceibias.n572 0.189894
R1193 commonsourceibias.n642 commonsourceibias.n572 0.189894
R1194 commonsourceibias.n643 commonsourceibias.n642 0.189894
R1195 commonsourceibias.n644 commonsourceibias.n643 0.189894
R1196 commonsourceibias.n644 commonsourceibias.n570 0.189894
R1197 commonsourceibias.n649 commonsourceibias.n570 0.189894
R1198 commonsourceibias.n650 commonsourceibias.n649 0.189894
R1199 commonsourceibias.n651 commonsourceibias.n650 0.189894
R1200 commonsourceibias.n651 commonsourceibias.n568 0.189894
R1201 commonsourceibias.n159 commonsourceibias.n158 0.170955
R1202 commonsourceibias.n160 commonsourceibias.n159 0.170955
R1203 commonsourceibias.n531 commonsourceibias.n425 0.170955
R1204 commonsourceibias.n532 commonsourceibias.n531 0.170955
R1205 gnd.n4036 gnd.n3722 939.716
R1206 gnd.n6577 gnd.n520 870.29
R1207 gnd.n211 gnd.n201 795.207
R1208 gnd.n7024 gnd.n7023 795.207
R1209 gnd.n1399 gnd.n1287 795.207
R1210 gnd.n5591 gnd.n1401 795.207
R1211 gnd.n979 gnd.n967 795.207
R1212 gnd.n4625 gnd.n4624 795.207
R1213 gnd.n3876 gnd.n3759 795.207
R1214 gnd.n3915 gnd.n2237 795.207
R1215 gnd.n4352 gnd.n4351 771.183
R1216 gnd.n5780 gnd.n1223 771.183
R1217 gnd.n4632 gnd.n2007 771.183
R1218 gnd.n5782 gnd.n1218 771.183
R1219 gnd.n3630 gnd.n2245 766.379
R1220 gnd.n3633 gnd.n3632 766.379
R1221 gnd.n2872 gnd.n2775 766.379
R1222 gnd.n2868 gnd.n2773 766.379
R1223 gnd.n3721 gnd.n2267 756.769
R1224 gnd.n3624 gnd.n3623 756.769
R1225 gnd.n2965 gnd.n2682 756.769
R1226 gnd.n2963 gnd.n2685 756.769
R1227 gnd.n7184 gnd.n205 739.952
R1228 gnd.n7060 gnd.n7059 739.952
R1229 gnd.n5594 gnd.n5593 739.952
R1230 gnd.n5711 gnd.n1333 739.952
R1231 gnd.n6024 gnd.n972 739.952
R1232 gnd.n4574 gnd.n2038 739.952
R1233 gnd.n4039 gnd.n4038 739.952
R1234 gnd.n4034 gnd.n2233 739.952
R1235 gnd.n6249 gnd.n712 655.866
R1236 gnd.n6576 gnd.n521 655.866
R1237 gnd.n6788 gnd.n6787 655.866
R1238 gnd.n6081 gnd.n882 655.866
R1239 gnd.n6250 gnd.n6249 585
R1240 gnd.n6249 gnd.n6248 585
R1241 gnd.n716 gnd.n715 585
R1242 gnd.n6247 gnd.n716 585
R1243 gnd.n6245 gnd.n6244 585
R1244 gnd.n6246 gnd.n6245 585
R1245 gnd.n6243 gnd.n718 585
R1246 gnd.n718 gnd.n717 585
R1247 gnd.n6242 gnd.n6241 585
R1248 gnd.n6241 gnd.n6240 585
R1249 gnd.n723 gnd.n722 585
R1250 gnd.n6239 gnd.n723 585
R1251 gnd.n6237 gnd.n6236 585
R1252 gnd.n6238 gnd.n6237 585
R1253 gnd.n6235 gnd.n725 585
R1254 gnd.n725 gnd.n724 585
R1255 gnd.n6234 gnd.n6233 585
R1256 gnd.n6233 gnd.n6232 585
R1257 gnd.n731 gnd.n730 585
R1258 gnd.n6231 gnd.n731 585
R1259 gnd.n6229 gnd.n6228 585
R1260 gnd.n6230 gnd.n6229 585
R1261 gnd.n6227 gnd.n733 585
R1262 gnd.n733 gnd.n732 585
R1263 gnd.n6226 gnd.n6225 585
R1264 gnd.n6225 gnd.n6224 585
R1265 gnd.n739 gnd.n738 585
R1266 gnd.n6223 gnd.n739 585
R1267 gnd.n6221 gnd.n6220 585
R1268 gnd.n6222 gnd.n6221 585
R1269 gnd.n6219 gnd.n741 585
R1270 gnd.n741 gnd.n740 585
R1271 gnd.n6218 gnd.n6217 585
R1272 gnd.n6217 gnd.n6216 585
R1273 gnd.n747 gnd.n746 585
R1274 gnd.n6215 gnd.n747 585
R1275 gnd.n6213 gnd.n6212 585
R1276 gnd.n6214 gnd.n6213 585
R1277 gnd.n6211 gnd.n749 585
R1278 gnd.n749 gnd.n748 585
R1279 gnd.n6210 gnd.n6209 585
R1280 gnd.n6209 gnd.n6208 585
R1281 gnd.n755 gnd.n754 585
R1282 gnd.n6207 gnd.n755 585
R1283 gnd.n6205 gnd.n6204 585
R1284 gnd.n6206 gnd.n6205 585
R1285 gnd.n6203 gnd.n757 585
R1286 gnd.n757 gnd.n756 585
R1287 gnd.n6202 gnd.n6201 585
R1288 gnd.n6201 gnd.n6200 585
R1289 gnd.n763 gnd.n762 585
R1290 gnd.n6199 gnd.n763 585
R1291 gnd.n6197 gnd.n6196 585
R1292 gnd.n6198 gnd.n6197 585
R1293 gnd.n6195 gnd.n765 585
R1294 gnd.n765 gnd.n764 585
R1295 gnd.n6194 gnd.n6193 585
R1296 gnd.n6193 gnd.n6192 585
R1297 gnd.n771 gnd.n770 585
R1298 gnd.n6191 gnd.n771 585
R1299 gnd.n6189 gnd.n6188 585
R1300 gnd.n6190 gnd.n6189 585
R1301 gnd.n6187 gnd.n773 585
R1302 gnd.n773 gnd.n772 585
R1303 gnd.n6186 gnd.n6185 585
R1304 gnd.n6185 gnd.n6184 585
R1305 gnd.n779 gnd.n778 585
R1306 gnd.n6183 gnd.n779 585
R1307 gnd.n6181 gnd.n6180 585
R1308 gnd.n6182 gnd.n6181 585
R1309 gnd.n6179 gnd.n781 585
R1310 gnd.n781 gnd.n780 585
R1311 gnd.n6178 gnd.n6177 585
R1312 gnd.n6177 gnd.n6176 585
R1313 gnd.n787 gnd.n786 585
R1314 gnd.n6175 gnd.n787 585
R1315 gnd.n6173 gnd.n6172 585
R1316 gnd.n6174 gnd.n6173 585
R1317 gnd.n6171 gnd.n789 585
R1318 gnd.n789 gnd.n788 585
R1319 gnd.n6170 gnd.n6169 585
R1320 gnd.n6169 gnd.n6168 585
R1321 gnd.n795 gnd.n794 585
R1322 gnd.n6167 gnd.n795 585
R1323 gnd.n6165 gnd.n6164 585
R1324 gnd.n6166 gnd.n6165 585
R1325 gnd.n6163 gnd.n797 585
R1326 gnd.n797 gnd.n796 585
R1327 gnd.n6162 gnd.n6161 585
R1328 gnd.n6161 gnd.n6160 585
R1329 gnd.n803 gnd.n802 585
R1330 gnd.n6159 gnd.n803 585
R1331 gnd.n6157 gnd.n6156 585
R1332 gnd.n6158 gnd.n6157 585
R1333 gnd.n6155 gnd.n805 585
R1334 gnd.n805 gnd.n804 585
R1335 gnd.n6154 gnd.n6153 585
R1336 gnd.n6153 gnd.n6152 585
R1337 gnd.n811 gnd.n810 585
R1338 gnd.n6151 gnd.n811 585
R1339 gnd.n6149 gnd.n6148 585
R1340 gnd.n6150 gnd.n6149 585
R1341 gnd.n6147 gnd.n813 585
R1342 gnd.n813 gnd.n812 585
R1343 gnd.n6146 gnd.n6145 585
R1344 gnd.n6145 gnd.n6144 585
R1345 gnd.n819 gnd.n818 585
R1346 gnd.n6143 gnd.n819 585
R1347 gnd.n6141 gnd.n6140 585
R1348 gnd.n6142 gnd.n6141 585
R1349 gnd.n6139 gnd.n821 585
R1350 gnd.n821 gnd.n820 585
R1351 gnd.n6138 gnd.n6137 585
R1352 gnd.n6137 gnd.n6136 585
R1353 gnd.n827 gnd.n826 585
R1354 gnd.n6135 gnd.n827 585
R1355 gnd.n6133 gnd.n6132 585
R1356 gnd.n6134 gnd.n6133 585
R1357 gnd.n6131 gnd.n829 585
R1358 gnd.n829 gnd.n828 585
R1359 gnd.n6130 gnd.n6129 585
R1360 gnd.n6129 gnd.n6128 585
R1361 gnd.n835 gnd.n834 585
R1362 gnd.n6127 gnd.n835 585
R1363 gnd.n6125 gnd.n6124 585
R1364 gnd.n6126 gnd.n6125 585
R1365 gnd.n6123 gnd.n837 585
R1366 gnd.n837 gnd.n836 585
R1367 gnd.n6122 gnd.n6121 585
R1368 gnd.n6121 gnd.n6120 585
R1369 gnd.n843 gnd.n842 585
R1370 gnd.n6119 gnd.n843 585
R1371 gnd.n6117 gnd.n6116 585
R1372 gnd.n6118 gnd.n6117 585
R1373 gnd.n6115 gnd.n845 585
R1374 gnd.n845 gnd.n844 585
R1375 gnd.n6114 gnd.n6113 585
R1376 gnd.n6113 gnd.n6112 585
R1377 gnd.n851 gnd.n850 585
R1378 gnd.n6111 gnd.n851 585
R1379 gnd.n6109 gnd.n6108 585
R1380 gnd.n6110 gnd.n6109 585
R1381 gnd.n6107 gnd.n853 585
R1382 gnd.n853 gnd.n852 585
R1383 gnd.n6106 gnd.n6105 585
R1384 gnd.n6105 gnd.n6104 585
R1385 gnd.n859 gnd.n858 585
R1386 gnd.n6103 gnd.n859 585
R1387 gnd.n6101 gnd.n6100 585
R1388 gnd.n6102 gnd.n6101 585
R1389 gnd.n6099 gnd.n861 585
R1390 gnd.n861 gnd.n860 585
R1391 gnd.n6098 gnd.n6097 585
R1392 gnd.n6097 gnd.n6096 585
R1393 gnd.n867 gnd.n866 585
R1394 gnd.n6095 gnd.n867 585
R1395 gnd.n6093 gnd.n6092 585
R1396 gnd.n6094 gnd.n6093 585
R1397 gnd.n6091 gnd.n869 585
R1398 gnd.n869 gnd.n868 585
R1399 gnd.n6090 gnd.n6089 585
R1400 gnd.n6089 gnd.n6088 585
R1401 gnd.n875 gnd.n874 585
R1402 gnd.n6087 gnd.n875 585
R1403 gnd.n6085 gnd.n6084 585
R1404 gnd.n6086 gnd.n6085 585
R1405 gnd.n6083 gnd.n877 585
R1406 gnd.n877 gnd.n876 585
R1407 gnd.n713 gnd.n712 585
R1408 gnd.n712 gnd.n711 585
R1409 gnd.n6255 gnd.n6254 585
R1410 gnd.n6256 gnd.n6255 585
R1411 gnd.n710 gnd.n709 585
R1412 gnd.n6257 gnd.n710 585
R1413 gnd.n6260 gnd.n6259 585
R1414 gnd.n6259 gnd.n6258 585
R1415 gnd.n707 gnd.n706 585
R1416 gnd.n706 gnd.n705 585
R1417 gnd.n6265 gnd.n6264 585
R1418 gnd.n6266 gnd.n6265 585
R1419 gnd.n704 gnd.n703 585
R1420 gnd.n6267 gnd.n704 585
R1421 gnd.n6270 gnd.n6269 585
R1422 gnd.n6269 gnd.n6268 585
R1423 gnd.n701 gnd.n700 585
R1424 gnd.n700 gnd.n699 585
R1425 gnd.n6275 gnd.n6274 585
R1426 gnd.n6276 gnd.n6275 585
R1427 gnd.n698 gnd.n697 585
R1428 gnd.n6277 gnd.n698 585
R1429 gnd.n6280 gnd.n6279 585
R1430 gnd.n6279 gnd.n6278 585
R1431 gnd.n695 gnd.n694 585
R1432 gnd.n694 gnd.n693 585
R1433 gnd.n6285 gnd.n6284 585
R1434 gnd.n6286 gnd.n6285 585
R1435 gnd.n692 gnd.n691 585
R1436 gnd.n6287 gnd.n692 585
R1437 gnd.n6290 gnd.n6289 585
R1438 gnd.n6289 gnd.n6288 585
R1439 gnd.n689 gnd.n688 585
R1440 gnd.n688 gnd.n687 585
R1441 gnd.n6295 gnd.n6294 585
R1442 gnd.n6296 gnd.n6295 585
R1443 gnd.n686 gnd.n685 585
R1444 gnd.n6297 gnd.n686 585
R1445 gnd.n6300 gnd.n6299 585
R1446 gnd.n6299 gnd.n6298 585
R1447 gnd.n683 gnd.n682 585
R1448 gnd.n682 gnd.n681 585
R1449 gnd.n6305 gnd.n6304 585
R1450 gnd.n6306 gnd.n6305 585
R1451 gnd.n680 gnd.n679 585
R1452 gnd.n6307 gnd.n680 585
R1453 gnd.n6310 gnd.n6309 585
R1454 gnd.n6309 gnd.n6308 585
R1455 gnd.n677 gnd.n676 585
R1456 gnd.n676 gnd.n675 585
R1457 gnd.n6315 gnd.n6314 585
R1458 gnd.n6316 gnd.n6315 585
R1459 gnd.n674 gnd.n673 585
R1460 gnd.n6317 gnd.n674 585
R1461 gnd.n6320 gnd.n6319 585
R1462 gnd.n6319 gnd.n6318 585
R1463 gnd.n671 gnd.n670 585
R1464 gnd.n670 gnd.n669 585
R1465 gnd.n6325 gnd.n6324 585
R1466 gnd.n6326 gnd.n6325 585
R1467 gnd.n668 gnd.n667 585
R1468 gnd.n6327 gnd.n668 585
R1469 gnd.n6330 gnd.n6329 585
R1470 gnd.n6329 gnd.n6328 585
R1471 gnd.n665 gnd.n664 585
R1472 gnd.n664 gnd.n663 585
R1473 gnd.n6335 gnd.n6334 585
R1474 gnd.n6336 gnd.n6335 585
R1475 gnd.n662 gnd.n661 585
R1476 gnd.n6337 gnd.n662 585
R1477 gnd.n6340 gnd.n6339 585
R1478 gnd.n6339 gnd.n6338 585
R1479 gnd.n659 gnd.n658 585
R1480 gnd.n658 gnd.n657 585
R1481 gnd.n6345 gnd.n6344 585
R1482 gnd.n6346 gnd.n6345 585
R1483 gnd.n656 gnd.n655 585
R1484 gnd.n6347 gnd.n656 585
R1485 gnd.n6350 gnd.n6349 585
R1486 gnd.n6349 gnd.n6348 585
R1487 gnd.n653 gnd.n652 585
R1488 gnd.n652 gnd.n651 585
R1489 gnd.n6355 gnd.n6354 585
R1490 gnd.n6356 gnd.n6355 585
R1491 gnd.n650 gnd.n649 585
R1492 gnd.n6357 gnd.n650 585
R1493 gnd.n6360 gnd.n6359 585
R1494 gnd.n6359 gnd.n6358 585
R1495 gnd.n647 gnd.n646 585
R1496 gnd.n646 gnd.n645 585
R1497 gnd.n6365 gnd.n6364 585
R1498 gnd.n6366 gnd.n6365 585
R1499 gnd.n644 gnd.n643 585
R1500 gnd.n6367 gnd.n644 585
R1501 gnd.n6370 gnd.n6369 585
R1502 gnd.n6369 gnd.n6368 585
R1503 gnd.n641 gnd.n640 585
R1504 gnd.n640 gnd.n639 585
R1505 gnd.n6375 gnd.n6374 585
R1506 gnd.n6376 gnd.n6375 585
R1507 gnd.n638 gnd.n637 585
R1508 gnd.n6377 gnd.n638 585
R1509 gnd.n6380 gnd.n6379 585
R1510 gnd.n6379 gnd.n6378 585
R1511 gnd.n635 gnd.n634 585
R1512 gnd.n634 gnd.n633 585
R1513 gnd.n6385 gnd.n6384 585
R1514 gnd.n6386 gnd.n6385 585
R1515 gnd.n632 gnd.n631 585
R1516 gnd.n6387 gnd.n632 585
R1517 gnd.n6390 gnd.n6389 585
R1518 gnd.n6389 gnd.n6388 585
R1519 gnd.n629 gnd.n628 585
R1520 gnd.n628 gnd.n627 585
R1521 gnd.n6395 gnd.n6394 585
R1522 gnd.n6396 gnd.n6395 585
R1523 gnd.n626 gnd.n625 585
R1524 gnd.n6397 gnd.n626 585
R1525 gnd.n6400 gnd.n6399 585
R1526 gnd.n6399 gnd.n6398 585
R1527 gnd.n623 gnd.n622 585
R1528 gnd.n622 gnd.n621 585
R1529 gnd.n6405 gnd.n6404 585
R1530 gnd.n6406 gnd.n6405 585
R1531 gnd.n620 gnd.n619 585
R1532 gnd.n6407 gnd.n620 585
R1533 gnd.n6410 gnd.n6409 585
R1534 gnd.n6409 gnd.n6408 585
R1535 gnd.n617 gnd.n616 585
R1536 gnd.n616 gnd.n615 585
R1537 gnd.n6415 gnd.n6414 585
R1538 gnd.n6416 gnd.n6415 585
R1539 gnd.n614 gnd.n613 585
R1540 gnd.n6417 gnd.n614 585
R1541 gnd.n6420 gnd.n6419 585
R1542 gnd.n6419 gnd.n6418 585
R1543 gnd.n611 gnd.n610 585
R1544 gnd.n610 gnd.n609 585
R1545 gnd.n6425 gnd.n6424 585
R1546 gnd.n6426 gnd.n6425 585
R1547 gnd.n608 gnd.n607 585
R1548 gnd.n6427 gnd.n608 585
R1549 gnd.n6430 gnd.n6429 585
R1550 gnd.n6429 gnd.n6428 585
R1551 gnd.n605 gnd.n604 585
R1552 gnd.n604 gnd.n603 585
R1553 gnd.n6435 gnd.n6434 585
R1554 gnd.n6436 gnd.n6435 585
R1555 gnd.n602 gnd.n601 585
R1556 gnd.n6437 gnd.n602 585
R1557 gnd.n6440 gnd.n6439 585
R1558 gnd.n6439 gnd.n6438 585
R1559 gnd.n599 gnd.n598 585
R1560 gnd.n598 gnd.n597 585
R1561 gnd.n6445 gnd.n6444 585
R1562 gnd.n6446 gnd.n6445 585
R1563 gnd.n596 gnd.n595 585
R1564 gnd.n6447 gnd.n596 585
R1565 gnd.n6450 gnd.n6449 585
R1566 gnd.n6449 gnd.n6448 585
R1567 gnd.n593 gnd.n592 585
R1568 gnd.n592 gnd.n591 585
R1569 gnd.n6455 gnd.n6454 585
R1570 gnd.n6456 gnd.n6455 585
R1571 gnd.n590 gnd.n589 585
R1572 gnd.n6457 gnd.n590 585
R1573 gnd.n6460 gnd.n6459 585
R1574 gnd.n6459 gnd.n6458 585
R1575 gnd.n587 gnd.n586 585
R1576 gnd.n586 gnd.n585 585
R1577 gnd.n6465 gnd.n6464 585
R1578 gnd.n6466 gnd.n6465 585
R1579 gnd.n584 gnd.n583 585
R1580 gnd.n6467 gnd.n584 585
R1581 gnd.n6470 gnd.n6469 585
R1582 gnd.n6469 gnd.n6468 585
R1583 gnd.n581 gnd.n580 585
R1584 gnd.n580 gnd.n579 585
R1585 gnd.n6475 gnd.n6474 585
R1586 gnd.n6476 gnd.n6475 585
R1587 gnd.n578 gnd.n577 585
R1588 gnd.n6477 gnd.n578 585
R1589 gnd.n6480 gnd.n6479 585
R1590 gnd.n6479 gnd.n6478 585
R1591 gnd.n575 gnd.n574 585
R1592 gnd.n574 gnd.n573 585
R1593 gnd.n6485 gnd.n6484 585
R1594 gnd.n6486 gnd.n6485 585
R1595 gnd.n572 gnd.n571 585
R1596 gnd.n6487 gnd.n572 585
R1597 gnd.n6490 gnd.n6489 585
R1598 gnd.n6489 gnd.n6488 585
R1599 gnd.n569 gnd.n568 585
R1600 gnd.n568 gnd.n567 585
R1601 gnd.n6495 gnd.n6494 585
R1602 gnd.n6496 gnd.n6495 585
R1603 gnd.n566 gnd.n565 585
R1604 gnd.n6497 gnd.n566 585
R1605 gnd.n6500 gnd.n6499 585
R1606 gnd.n6499 gnd.n6498 585
R1607 gnd.n563 gnd.n562 585
R1608 gnd.n562 gnd.n561 585
R1609 gnd.n6505 gnd.n6504 585
R1610 gnd.n6506 gnd.n6505 585
R1611 gnd.n560 gnd.n559 585
R1612 gnd.n6507 gnd.n560 585
R1613 gnd.n6510 gnd.n6509 585
R1614 gnd.n6509 gnd.n6508 585
R1615 gnd.n557 gnd.n556 585
R1616 gnd.n556 gnd.n555 585
R1617 gnd.n6515 gnd.n6514 585
R1618 gnd.n6516 gnd.n6515 585
R1619 gnd.n554 gnd.n553 585
R1620 gnd.n6517 gnd.n554 585
R1621 gnd.n6520 gnd.n6519 585
R1622 gnd.n6519 gnd.n6518 585
R1623 gnd.n551 gnd.n550 585
R1624 gnd.n550 gnd.n549 585
R1625 gnd.n6525 gnd.n6524 585
R1626 gnd.n6526 gnd.n6525 585
R1627 gnd.n548 gnd.n547 585
R1628 gnd.n6527 gnd.n548 585
R1629 gnd.n6530 gnd.n6529 585
R1630 gnd.n6529 gnd.n6528 585
R1631 gnd.n545 gnd.n544 585
R1632 gnd.n544 gnd.n543 585
R1633 gnd.n6535 gnd.n6534 585
R1634 gnd.n6536 gnd.n6535 585
R1635 gnd.n542 gnd.n541 585
R1636 gnd.n6537 gnd.n542 585
R1637 gnd.n6540 gnd.n6539 585
R1638 gnd.n6539 gnd.n6538 585
R1639 gnd.n539 gnd.n538 585
R1640 gnd.n538 gnd.n537 585
R1641 gnd.n6545 gnd.n6544 585
R1642 gnd.n6546 gnd.n6545 585
R1643 gnd.n536 gnd.n535 585
R1644 gnd.n6547 gnd.n536 585
R1645 gnd.n6550 gnd.n6549 585
R1646 gnd.n6549 gnd.n6548 585
R1647 gnd.n533 gnd.n532 585
R1648 gnd.n532 gnd.n531 585
R1649 gnd.n6555 gnd.n6554 585
R1650 gnd.n6556 gnd.n6555 585
R1651 gnd.n530 gnd.n529 585
R1652 gnd.n6557 gnd.n530 585
R1653 gnd.n6560 gnd.n6559 585
R1654 gnd.n6559 gnd.n6558 585
R1655 gnd.n527 gnd.n526 585
R1656 gnd.n526 gnd.n525 585
R1657 gnd.n6566 gnd.n6565 585
R1658 gnd.n6567 gnd.n6566 585
R1659 gnd.n524 gnd.n523 585
R1660 gnd.n6568 gnd.n524 585
R1661 gnd.n6571 gnd.n6570 585
R1662 gnd.n6570 gnd.n6569 585
R1663 gnd.n6572 gnd.n521 585
R1664 gnd.n521 gnd.n520 585
R1665 gnd.n396 gnd.n395 585
R1666 gnd.n6779 gnd.n395 585
R1667 gnd.n6782 gnd.n6781 585
R1668 gnd.n6781 gnd.n6780 585
R1669 gnd.n399 gnd.n398 585
R1670 gnd.n6778 gnd.n399 585
R1671 gnd.n6776 gnd.n6775 585
R1672 gnd.n6777 gnd.n6776 585
R1673 gnd.n402 gnd.n401 585
R1674 gnd.n401 gnd.n400 585
R1675 gnd.n6771 gnd.n6770 585
R1676 gnd.n6770 gnd.n6769 585
R1677 gnd.n405 gnd.n404 585
R1678 gnd.n6768 gnd.n405 585
R1679 gnd.n6766 gnd.n6765 585
R1680 gnd.n6767 gnd.n6766 585
R1681 gnd.n408 gnd.n407 585
R1682 gnd.n407 gnd.n406 585
R1683 gnd.n6761 gnd.n6760 585
R1684 gnd.n6760 gnd.n6759 585
R1685 gnd.n411 gnd.n410 585
R1686 gnd.n6758 gnd.n411 585
R1687 gnd.n6756 gnd.n6755 585
R1688 gnd.n6757 gnd.n6756 585
R1689 gnd.n414 gnd.n413 585
R1690 gnd.n413 gnd.n412 585
R1691 gnd.n6751 gnd.n6750 585
R1692 gnd.n6750 gnd.n6749 585
R1693 gnd.n417 gnd.n416 585
R1694 gnd.n6748 gnd.n417 585
R1695 gnd.n6746 gnd.n6745 585
R1696 gnd.n6747 gnd.n6746 585
R1697 gnd.n420 gnd.n419 585
R1698 gnd.n419 gnd.n418 585
R1699 gnd.n6741 gnd.n6740 585
R1700 gnd.n6740 gnd.n6739 585
R1701 gnd.n423 gnd.n422 585
R1702 gnd.n6738 gnd.n423 585
R1703 gnd.n6736 gnd.n6735 585
R1704 gnd.n6737 gnd.n6736 585
R1705 gnd.n426 gnd.n425 585
R1706 gnd.n425 gnd.n424 585
R1707 gnd.n6731 gnd.n6730 585
R1708 gnd.n6730 gnd.n6729 585
R1709 gnd.n429 gnd.n428 585
R1710 gnd.n6728 gnd.n429 585
R1711 gnd.n6726 gnd.n6725 585
R1712 gnd.n6727 gnd.n6726 585
R1713 gnd.n432 gnd.n431 585
R1714 gnd.n431 gnd.n430 585
R1715 gnd.n6721 gnd.n6720 585
R1716 gnd.n6720 gnd.n6719 585
R1717 gnd.n435 gnd.n434 585
R1718 gnd.n6718 gnd.n435 585
R1719 gnd.n6716 gnd.n6715 585
R1720 gnd.n6717 gnd.n6716 585
R1721 gnd.n438 gnd.n437 585
R1722 gnd.n437 gnd.n436 585
R1723 gnd.n6711 gnd.n6710 585
R1724 gnd.n6710 gnd.n6709 585
R1725 gnd.n441 gnd.n440 585
R1726 gnd.n6708 gnd.n441 585
R1727 gnd.n6706 gnd.n6705 585
R1728 gnd.n6707 gnd.n6706 585
R1729 gnd.n444 gnd.n443 585
R1730 gnd.n443 gnd.n442 585
R1731 gnd.n6701 gnd.n6700 585
R1732 gnd.n6700 gnd.n6699 585
R1733 gnd.n447 gnd.n446 585
R1734 gnd.n6698 gnd.n447 585
R1735 gnd.n6696 gnd.n6695 585
R1736 gnd.n6697 gnd.n6696 585
R1737 gnd.n450 gnd.n449 585
R1738 gnd.n449 gnd.n448 585
R1739 gnd.n6691 gnd.n6690 585
R1740 gnd.n6690 gnd.n6689 585
R1741 gnd.n453 gnd.n452 585
R1742 gnd.n6688 gnd.n453 585
R1743 gnd.n6686 gnd.n6685 585
R1744 gnd.n6687 gnd.n6686 585
R1745 gnd.n456 gnd.n455 585
R1746 gnd.n455 gnd.n454 585
R1747 gnd.n6681 gnd.n6680 585
R1748 gnd.n6680 gnd.n6679 585
R1749 gnd.n459 gnd.n458 585
R1750 gnd.n6678 gnd.n459 585
R1751 gnd.n6676 gnd.n6675 585
R1752 gnd.n6677 gnd.n6676 585
R1753 gnd.n462 gnd.n461 585
R1754 gnd.n461 gnd.n460 585
R1755 gnd.n6671 gnd.n6670 585
R1756 gnd.n6670 gnd.n6669 585
R1757 gnd.n465 gnd.n464 585
R1758 gnd.n6668 gnd.n465 585
R1759 gnd.n6666 gnd.n6665 585
R1760 gnd.n6667 gnd.n6666 585
R1761 gnd.n468 gnd.n467 585
R1762 gnd.n467 gnd.n466 585
R1763 gnd.n6661 gnd.n6660 585
R1764 gnd.n6660 gnd.n6659 585
R1765 gnd.n471 gnd.n470 585
R1766 gnd.n6658 gnd.n471 585
R1767 gnd.n6656 gnd.n6655 585
R1768 gnd.n6657 gnd.n6656 585
R1769 gnd.n474 gnd.n473 585
R1770 gnd.n473 gnd.n472 585
R1771 gnd.n6651 gnd.n6650 585
R1772 gnd.n6650 gnd.n6649 585
R1773 gnd.n477 gnd.n476 585
R1774 gnd.n6648 gnd.n477 585
R1775 gnd.n6646 gnd.n6645 585
R1776 gnd.n6647 gnd.n6646 585
R1777 gnd.n480 gnd.n479 585
R1778 gnd.n479 gnd.n478 585
R1779 gnd.n6641 gnd.n6640 585
R1780 gnd.n6640 gnd.n6639 585
R1781 gnd.n483 gnd.n482 585
R1782 gnd.n6638 gnd.n483 585
R1783 gnd.n6636 gnd.n6635 585
R1784 gnd.n6637 gnd.n6636 585
R1785 gnd.n486 gnd.n485 585
R1786 gnd.n485 gnd.n484 585
R1787 gnd.n6631 gnd.n6630 585
R1788 gnd.n6630 gnd.n6629 585
R1789 gnd.n489 gnd.n488 585
R1790 gnd.n6628 gnd.n489 585
R1791 gnd.n6626 gnd.n6625 585
R1792 gnd.n6627 gnd.n6626 585
R1793 gnd.n492 gnd.n491 585
R1794 gnd.n491 gnd.n490 585
R1795 gnd.n6621 gnd.n6620 585
R1796 gnd.n6620 gnd.n6619 585
R1797 gnd.n495 gnd.n494 585
R1798 gnd.n6618 gnd.n495 585
R1799 gnd.n6616 gnd.n6615 585
R1800 gnd.n6617 gnd.n6616 585
R1801 gnd.n498 gnd.n497 585
R1802 gnd.n497 gnd.n496 585
R1803 gnd.n6611 gnd.n6610 585
R1804 gnd.n6610 gnd.n6609 585
R1805 gnd.n501 gnd.n500 585
R1806 gnd.n6608 gnd.n501 585
R1807 gnd.n6606 gnd.n6605 585
R1808 gnd.n6607 gnd.n6606 585
R1809 gnd.n504 gnd.n503 585
R1810 gnd.n503 gnd.n502 585
R1811 gnd.n6601 gnd.n6600 585
R1812 gnd.n6600 gnd.n6599 585
R1813 gnd.n507 gnd.n506 585
R1814 gnd.n6598 gnd.n507 585
R1815 gnd.n6596 gnd.n6595 585
R1816 gnd.n6597 gnd.n6596 585
R1817 gnd.n510 gnd.n509 585
R1818 gnd.n509 gnd.n508 585
R1819 gnd.n6591 gnd.n6590 585
R1820 gnd.n6590 gnd.n6589 585
R1821 gnd.n513 gnd.n512 585
R1822 gnd.n6588 gnd.n513 585
R1823 gnd.n6586 gnd.n6585 585
R1824 gnd.n6587 gnd.n6586 585
R1825 gnd.n516 gnd.n515 585
R1826 gnd.n515 gnd.n514 585
R1827 gnd.n6581 gnd.n6580 585
R1828 gnd.n6580 gnd.n6579 585
R1829 gnd.n519 gnd.n518 585
R1830 gnd.n6578 gnd.n519 585
R1831 gnd.n6576 gnd.n6575 585
R1832 gnd.n6577 gnd.n6576 585
R1833 gnd.n967 gnd.n966 585
R1834 gnd.n4623 gnd.n967 585
R1835 gnd.n6033 gnd.n6032 585
R1836 gnd.n6032 gnd.n6031 585
R1837 gnd.n6034 gnd.n962 585
R1838 gnd.n4583 gnd.n962 585
R1839 gnd.n6036 gnd.n6035 585
R1840 gnd.n6037 gnd.n6036 585
R1841 gnd.n946 gnd.n945 585
R1842 gnd.n4331 gnd.n946 585
R1843 gnd.n6045 gnd.n6044 585
R1844 gnd.n6044 gnd.n6043 585
R1845 gnd.n6046 gnd.n941 585
R1846 gnd.n4596 gnd.n941 585
R1847 gnd.n6048 gnd.n6047 585
R1848 gnd.n6049 gnd.n6048 585
R1849 gnd.n927 gnd.n926 585
R1850 gnd.n4324 gnd.n927 585
R1851 gnd.n6057 gnd.n6056 585
R1852 gnd.n6056 gnd.n6055 585
R1853 gnd.n6058 gnd.n922 585
R1854 gnd.n4316 gnd.n922 585
R1855 gnd.n6060 gnd.n6059 585
R1856 gnd.n6061 gnd.n6060 585
R1857 gnd.n906 gnd.n905 585
R1858 gnd.n4282 gnd.n906 585
R1859 gnd.n6069 gnd.n6068 585
R1860 gnd.n6068 gnd.n6067 585
R1861 gnd.n6070 gnd.n900 585
R1862 gnd.n4290 gnd.n900 585
R1863 gnd.n6072 gnd.n6071 585
R1864 gnd.n6073 gnd.n6072 585
R1865 gnd.n901 gnd.n899 585
R1866 gnd.n4271 gnd.n899 585
R1867 gnd.n4246 gnd.n887 585
R1868 gnd.n6079 gnd.n887 585
R1869 gnd.n4248 gnd.n4247 585
R1870 gnd.n4247 gnd.n883 585
R1871 gnd.n4249 gnd.n2077 585
R1872 gnd.n4262 gnd.n2077 585
R1873 gnd.n4250 gnd.n2088 585
R1874 gnd.n2088 gnd.n2086 585
R1875 gnd.n4252 gnd.n4251 585
R1876 gnd.n4253 gnd.n4252 585
R1877 gnd.n2089 gnd.n2087 585
R1878 gnd.n2087 gnd.n2083 585
R1879 gnd.n4222 gnd.n2098 585
R1880 gnd.n4234 gnd.n2098 585
R1881 gnd.n4223 gnd.n2107 585
R1882 gnd.n2107 gnd.n2096 585
R1883 gnd.n4225 gnd.n4224 585
R1884 gnd.n4226 gnd.n4225 585
R1885 gnd.n2108 gnd.n2106 585
R1886 gnd.n4215 gnd.n2106 585
R1887 gnd.n4178 gnd.n4177 585
R1888 gnd.n4177 gnd.n2113 585
R1889 gnd.n4179 gnd.n2122 585
R1890 gnd.n4193 gnd.n2122 585
R1891 gnd.n4180 gnd.n2132 585
R1892 gnd.n2132 gnd.n2120 585
R1893 gnd.n4182 gnd.n4181 585
R1894 gnd.n4183 gnd.n4182 585
R1895 gnd.n2133 gnd.n2131 585
R1896 gnd.n4168 gnd.n2131 585
R1897 gnd.n4143 gnd.n4142 585
R1898 gnd.n4142 gnd.n2139 585
R1899 gnd.n4144 gnd.n2146 585
R1900 gnd.n4158 gnd.n2146 585
R1901 gnd.n4145 gnd.n2157 585
R1902 gnd.n2157 gnd.n2155 585
R1903 gnd.n4147 gnd.n4146 585
R1904 gnd.n4148 gnd.n4147 585
R1905 gnd.n2158 gnd.n2156 585
R1906 gnd.n4133 gnd.n2156 585
R1907 gnd.n4108 gnd.n4107 585
R1908 gnd.n4107 gnd.n2164 585
R1909 gnd.n4109 gnd.n2171 585
R1910 gnd.n4123 gnd.n2171 585
R1911 gnd.n4110 gnd.n2183 585
R1912 gnd.n2183 gnd.n2181 585
R1913 gnd.n4112 gnd.n4111 585
R1914 gnd.n4113 gnd.n4112 585
R1915 gnd.n2184 gnd.n2182 585
R1916 gnd.n2182 gnd.n2178 585
R1917 gnd.n4085 gnd.n2192 585
R1918 gnd.n4097 gnd.n2192 585
R1919 gnd.n4086 gnd.n2202 585
R1920 gnd.n2202 gnd.n2190 585
R1921 gnd.n4088 gnd.n4087 585
R1922 gnd.n4089 gnd.n4088 585
R1923 gnd.n2203 gnd.n2201 585
R1924 gnd.n2201 gnd.n2198 585
R1925 gnd.n4065 gnd.n2209 585
R1926 gnd.n4077 gnd.n2209 585
R1927 gnd.n4066 gnd.n2220 585
R1928 gnd.n2220 gnd.n2218 585
R1929 gnd.n4068 gnd.n4067 585
R1930 gnd.n4069 gnd.n4068 585
R1931 gnd.n2221 gnd.n2219 585
R1932 gnd.n2219 gnd.n2215 585
R1933 gnd.n4045 gnd.n2228 585
R1934 gnd.n4057 gnd.n2228 585
R1935 gnd.n4046 gnd.n2238 585
R1936 gnd.n2238 gnd.n2226 585
R1937 gnd.n4048 gnd.n4047 585
R1938 gnd.n4049 gnd.n4048 585
R1939 gnd.n2239 gnd.n2237 585
R1940 gnd.n2237 gnd.n2234 585
R1941 gnd.n3916 gnd.n3915 585
R1942 gnd.n3914 gnd.n3913 585
R1943 gnd.n3912 gnd.n3911 585
R1944 gnd.n3910 gnd.n3909 585
R1945 gnd.n3908 gnd.n3907 585
R1946 gnd.n3906 gnd.n3905 585
R1947 gnd.n3904 gnd.n3903 585
R1948 gnd.n3902 gnd.n3901 585
R1949 gnd.n3900 gnd.n3899 585
R1950 gnd.n3898 gnd.n3897 585
R1951 gnd.n3896 gnd.n3895 585
R1952 gnd.n3894 gnd.n3893 585
R1953 gnd.n3892 gnd.n3891 585
R1954 gnd.n3890 gnd.n3889 585
R1955 gnd.n3888 gnd.n3887 585
R1956 gnd.n3886 gnd.n3885 585
R1957 gnd.n3884 gnd.n3883 585
R1958 gnd.n3843 gnd.n3840 585
R1959 gnd.n3879 gnd.n3759 585
R1960 gnd.n4036 gnd.n3759 585
R1961 gnd.n4626 gnd.n4625 585
R1962 gnd.n4420 gnd.n2036 585
R1963 gnd.n4432 gnd.n4421 585
R1964 gnd.n4433 gnd.n4419 585
R1965 gnd.n4418 gnd.n4410 585
R1966 gnd.n4440 gnd.n4409 585
R1967 gnd.n4441 gnd.n4408 585
R1968 gnd.n4402 gnd.n4401 585
R1969 gnd.n4448 gnd.n4400 585
R1970 gnd.n4449 gnd.n4399 585
R1971 gnd.n4398 gnd.n4390 585
R1972 gnd.n4456 gnd.n4389 585
R1973 gnd.n4457 gnd.n4388 585
R1974 gnd.n4382 gnd.n4381 585
R1975 gnd.n4464 gnd.n4380 585
R1976 gnd.n4465 gnd.n4379 585
R1977 gnd.n4378 gnd.n4370 585
R1978 gnd.n4472 gnd.n4369 585
R1979 gnd.n4473 gnd.n979 585
R1980 gnd.n6023 gnd.n979 585
R1981 gnd.n4624 gnd.n2037 585
R1982 gnd.n4624 gnd.n4623 585
R1983 gnd.n4585 gnd.n970 585
R1984 gnd.n6031 gnd.n970 585
R1985 gnd.n4588 gnd.n4584 585
R1986 gnd.n4584 gnd.n4583 585
R1987 gnd.n4589 gnd.n960 585
R1988 gnd.n6037 gnd.n960 585
R1989 gnd.n4590 gnd.n2054 585
R1990 gnd.n4331 gnd.n2054 585
R1991 gnd.n2051 gnd.n949 585
R1992 gnd.n6043 gnd.n949 585
R1993 gnd.n4595 gnd.n4594 585
R1994 gnd.n4596 gnd.n4595 585
R1995 gnd.n2050 gnd.n940 585
R1996 gnd.n6049 gnd.n940 585
R1997 gnd.n4323 gnd.n4322 585
R1998 gnd.n4324 gnd.n4323 585
R1999 gnd.n2057 gnd.n929 585
R2000 gnd.n6055 gnd.n929 585
R2001 gnd.n4318 gnd.n4317 585
R2002 gnd.n4317 gnd.n4316 585
R2003 gnd.n2059 gnd.n920 585
R2004 gnd.n6061 gnd.n920 585
R2005 gnd.n4284 gnd.n4283 585
R2006 gnd.n4283 gnd.n4282 585
R2007 gnd.n2068 gnd.n909 585
R2008 gnd.n6067 gnd.n909 585
R2009 gnd.n4289 gnd.n4288 585
R2010 gnd.n4290 gnd.n4289 585
R2011 gnd.n2067 gnd.n898 585
R2012 gnd.n6073 gnd.n898 585
R2013 gnd.n4270 gnd.n4269 585
R2014 gnd.n4271 gnd.n4270 585
R2015 gnd.n2072 gnd.n885 585
R2016 gnd.n6079 gnd.n885 585
R2017 gnd.n4265 gnd.n4264 585
R2018 gnd.n4264 gnd.n883 585
R2019 gnd.n4263 gnd.n2074 585
R2020 gnd.n4263 gnd.n4262 585
R2021 gnd.n4203 gnd.n2075 585
R2022 gnd.n2086 gnd.n2075 585
R2023 gnd.n4202 gnd.n2085 585
R2024 gnd.n4253 gnd.n2085 585
R2025 gnd.n4207 gnd.n4201 585
R2026 gnd.n4201 gnd.n2083 585
R2027 gnd.n4208 gnd.n2097 585
R2028 gnd.n4234 gnd.n2097 585
R2029 gnd.n4209 gnd.n4200 585
R2030 gnd.n4200 gnd.n2096 585
R2031 gnd.n2116 gnd.n2105 585
R2032 gnd.n4226 gnd.n2105 585
R2033 gnd.n4214 gnd.n4213 585
R2034 gnd.n4215 gnd.n4214 585
R2035 gnd.n2115 gnd.n2114 585
R2036 gnd.n2114 gnd.n2113 585
R2037 gnd.n4195 gnd.n4194 585
R2038 gnd.n4194 gnd.n4193 585
R2039 gnd.n2119 gnd.n2118 585
R2040 gnd.n2120 gnd.n2119 585
R2041 gnd.n4165 gnd.n2130 585
R2042 gnd.n4183 gnd.n2130 585
R2043 gnd.n4167 gnd.n4166 585
R2044 gnd.n4168 gnd.n4167 585
R2045 gnd.n2141 gnd.n2140 585
R2046 gnd.n2140 gnd.n2139 585
R2047 gnd.n4160 gnd.n4159 585
R2048 gnd.n4159 gnd.n4158 585
R2049 gnd.n2144 gnd.n2143 585
R2050 gnd.n2155 gnd.n2144 585
R2051 gnd.n4130 gnd.n2154 585
R2052 gnd.n4148 gnd.n2154 585
R2053 gnd.n4132 gnd.n4131 585
R2054 gnd.n4133 gnd.n4132 585
R2055 gnd.n2166 gnd.n2165 585
R2056 gnd.n2165 gnd.n2164 585
R2057 gnd.n4125 gnd.n4124 585
R2058 gnd.n4124 gnd.n4123 585
R2059 gnd.n2169 gnd.n2168 585
R2060 gnd.n2181 gnd.n2169 585
R2061 gnd.n3857 gnd.n2180 585
R2062 gnd.n4113 gnd.n2180 585
R2063 gnd.n3859 gnd.n3858 585
R2064 gnd.n3858 gnd.n2178 585
R2065 gnd.n3860 gnd.n2191 585
R2066 gnd.n4097 gnd.n2191 585
R2067 gnd.n3862 gnd.n3861 585
R2068 gnd.n3861 gnd.n2190 585
R2069 gnd.n3863 gnd.n2200 585
R2070 gnd.n4089 gnd.n2200 585
R2071 gnd.n3865 gnd.n3864 585
R2072 gnd.n3864 gnd.n2198 585
R2073 gnd.n3866 gnd.n2208 585
R2074 gnd.n4077 gnd.n2208 585
R2075 gnd.n3868 gnd.n3867 585
R2076 gnd.n3867 gnd.n2218 585
R2077 gnd.n3869 gnd.n2217 585
R2078 gnd.n4069 gnd.n2217 585
R2079 gnd.n3871 gnd.n3870 585
R2080 gnd.n3870 gnd.n2215 585
R2081 gnd.n3872 gnd.n2227 585
R2082 gnd.n4057 gnd.n2227 585
R2083 gnd.n3874 gnd.n3873 585
R2084 gnd.n3873 gnd.n2226 585
R2085 gnd.n3875 gnd.n2236 585
R2086 gnd.n4049 gnd.n2236 585
R2087 gnd.n3877 gnd.n3876 585
R2088 gnd.n3876 gnd.n2234 585
R2089 gnd.n3630 gnd.n3629 585
R2090 gnd.n3631 gnd.n3630 585
R2091 gnd.n2321 gnd.n2320 585
R2092 gnd.n2327 gnd.n2320 585
R2093 gnd.n3605 gnd.n2339 585
R2094 gnd.n2339 gnd.n2326 585
R2095 gnd.n3607 gnd.n3606 585
R2096 gnd.n3608 gnd.n3607 585
R2097 gnd.n2340 gnd.n2338 585
R2098 gnd.n2338 gnd.n2334 585
R2099 gnd.n3339 gnd.n3338 585
R2100 gnd.n3338 gnd.n3337 585
R2101 gnd.n2345 gnd.n2344 585
R2102 gnd.n3308 gnd.n2345 585
R2103 gnd.n3328 gnd.n3327 585
R2104 gnd.n3327 gnd.n3326 585
R2105 gnd.n2352 gnd.n2351 585
R2106 gnd.n3314 gnd.n2352 585
R2107 gnd.n3284 gnd.n2372 585
R2108 gnd.n2372 gnd.n2371 585
R2109 gnd.n3286 gnd.n3285 585
R2110 gnd.n3287 gnd.n3286 585
R2111 gnd.n2373 gnd.n2370 585
R2112 gnd.n2381 gnd.n2370 585
R2113 gnd.n3262 gnd.n2393 585
R2114 gnd.n2393 gnd.n2380 585
R2115 gnd.n3264 gnd.n3263 585
R2116 gnd.n3265 gnd.n3264 585
R2117 gnd.n2394 gnd.n2392 585
R2118 gnd.n2392 gnd.n2388 585
R2119 gnd.n3250 gnd.n3249 585
R2120 gnd.n3249 gnd.n3248 585
R2121 gnd.n2399 gnd.n2398 585
R2122 gnd.n2409 gnd.n2399 585
R2123 gnd.n3239 gnd.n3238 585
R2124 gnd.n3238 gnd.n3237 585
R2125 gnd.n2406 gnd.n2405 585
R2126 gnd.n3225 gnd.n2406 585
R2127 gnd.n3199 gnd.n2427 585
R2128 gnd.n2427 gnd.n2416 585
R2129 gnd.n3201 gnd.n3200 585
R2130 gnd.n3202 gnd.n3201 585
R2131 gnd.n2428 gnd.n2426 585
R2132 gnd.n2436 gnd.n2426 585
R2133 gnd.n3177 gnd.n2448 585
R2134 gnd.n2448 gnd.n2435 585
R2135 gnd.n3179 gnd.n3178 585
R2136 gnd.n3180 gnd.n3179 585
R2137 gnd.n2449 gnd.n2447 585
R2138 gnd.n2447 gnd.n2443 585
R2139 gnd.n3165 gnd.n3164 585
R2140 gnd.n3164 gnd.n3163 585
R2141 gnd.n2454 gnd.n2453 585
R2142 gnd.n2463 gnd.n2454 585
R2143 gnd.n3154 gnd.n3153 585
R2144 gnd.n3153 gnd.n3152 585
R2145 gnd.n2461 gnd.n2460 585
R2146 gnd.n3140 gnd.n2461 585
R2147 gnd.n2578 gnd.n2577 585
R2148 gnd.n2578 gnd.n2470 585
R2149 gnd.n3097 gnd.n3096 585
R2150 gnd.n3096 gnd.n3095 585
R2151 gnd.n3098 gnd.n2572 585
R2152 gnd.n2583 gnd.n2572 585
R2153 gnd.n3100 gnd.n3099 585
R2154 gnd.n3101 gnd.n3100 585
R2155 gnd.n2573 gnd.n2571 585
R2156 gnd.n2596 gnd.n2571 585
R2157 gnd.n2556 gnd.n2555 585
R2158 gnd.n2559 gnd.n2556 585
R2159 gnd.n3111 gnd.n3110 585
R2160 gnd.n3110 gnd.n3109 585
R2161 gnd.n3112 gnd.n2550 585
R2162 gnd.n3071 gnd.n2550 585
R2163 gnd.n3114 gnd.n3113 585
R2164 gnd.n3115 gnd.n3114 585
R2165 gnd.n2551 gnd.n2549 585
R2166 gnd.n2610 gnd.n2549 585
R2167 gnd.n3063 gnd.n3062 585
R2168 gnd.n3062 gnd.n3061 585
R2169 gnd.n2607 gnd.n2606 585
R2170 gnd.n3045 gnd.n2607 585
R2171 gnd.n3032 gnd.n2626 585
R2172 gnd.n2626 gnd.n2625 585
R2173 gnd.n3034 gnd.n3033 585
R2174 gnd.n3035 gnd.n3034 585
R2175 gnd.n2627 gnd.n2624 585
R2176 gnd.n2633 gnd.n2624 585
R2177 gnd.n3013 gnd.n3012 585
R2178 gnd.n3014 gnd.n3013 585
R2179 gnd.n2644 gnd.n2643 585
R2180 gnd.n2643 gnd.n2639 585
R2181 gnd.n3003 gnd.n3002 585
R2182 gnd.n3004 gnd.n3003 585
R2183 gnd.n2654 gnd.n2653 585
R2184 gnd.n2659 gnd.n2653 585
R2185 gnd.n2981 gnd.n2672 585
R2186 gnd.n2672 gnd.n2658 585
R2187 gnd.n2983 gnd.n2982 585
R2188 gnd.n2984 gnd.n2983 585
R2189 gnd.n2673 gnd.n2671 585
R2190 gnd.n2671 gnd.n2667 585
R2191 gnd.n2972 gnd.n2971 585
R2192 gnd.n2973 gnd.n2972 585
R2193 gnd.n2680 gnd.n2679 585
R2194 gnd.n2684 gnd.n2679 585
R2195 gnd.n2949 gnd.n2701 585
R2196 gnd.n2701 gnd.n2683 585
R2197 gnd.n2951 gnd.n2950 585
R2198 gnd.n2952 gnd.n2951 585
R2199 gnd.n2702 gnd.n2700 585
R2200 gnd.n2700 gnd.n2691 585
R2201 gnd.n2944 gnd.n2943 585
R2202 gnd.n2943 gnd.n2942 585
R2203 gnd.n2749 gnd.n2748 585
R2204 gnd.n2750 gnd.n2749 585
R2205 gnd.n2903 gnd.n2902 585
R2206 gnd.n2904 gnd.n2903 585
R2207 gnd.n2759 gnd.n2758 585
R2208 gnd.n2758 gnd.n2757 585
R2209 gnd.n2898 gnd.n2897 585
R2210 gnd.n2897 gnd.n2896 585
R2211 gnd.n2762 gnd.n2761 585
R2212 gnd.n2763 gnd.n2762 585
R2213 gnd.n2887 gnd.n2886 585
R2214 gnd.n2888 gnd.n2887 585
R2215 gnd.n2770 gnd.n2769 585
R2216 gnd.n2879 gnd.n2769 585
R2217 gnd.n2882 gnd.n2881 585
R2218 gnd.n2881 gnd.n2880 585
R2219 gnd.n2773 gnd.n2772 585
R2220 gnd.n2774 gnd.n2773 585
R2221 gnd.n2868 gnd.n2867 585
R2222 gnd.n2866 gnd.n2792 585
R2223 gnd.n2865 gnd.n2791 585
R2224 gnd.n2870 gnd.n2791 585
R2225 gnd.n2864 gnd.n2863 585
R2226 gnd.n2862 gnd.n2861 585
R2227 gnd.n2860 gnd.n2859 585
R2228 gnd.n2858 gnd.n2857 585
R2229 gnd.n2856 gnd.n2855 585
R2230 gnd.n2854 gnd.n2853 585
R2231 gnd.n2852 gnd.n2851 585
R2232 gnd.n2850 gnd.n2849 585
R2233 gnd.n2848 gnd.n2847 585
R2234 gnd.n2846 gnd.n2845 585
R2235 gnd.n2844 gnd.n2843 585
R2236 gnd.n2842 gnd.n2841 585
R2237 gnd.n2840 gnd.n2839 585
R2238 gnd.n2838 gnd.n2837 585
R2239 gnd.n2836 gnd.n2835 585
R2240 gnd.n2834 gnd.n2833 585
R2241 gnd.n2832 gnd.n2831 585
R2242 gnd.n2830 gnd.n2829 585
R2243 gnd.n2828 gnd.n2827 585
R2244 gnd.n2826 gnd.n2825 585
R2245 gnd.n2824 gnd.n2823 585
R2246 gnd.n2822 gnd.n2821 585
R2247 gnd.n2779 gnd.n2778 585
R2248 gnd.n2873 gnd.n2872 585
R2249 gnd.n3634 gnd.n3633 585
R2250 gnd.n3636 gnd.n3635 585
R2251 gnd.n3638 gnd.n3637 585
R2252 gnd.n3640 gnd.n3639 585
R2253 gnd.n3642 gnd.n3641 585
R2254 gnd.n3644 gnd.n3643 585
R2255 gnd.n3646 gnd.n3645 585
R2256 gnd.n3648 gnd.n3647 585
R2257 gnd.n3650 gnd.n3649 585
R2258 gnd.n3652 gnd.n3651 585
R2259 gnd.n3654 gnd.n3653 585
R2260 gnd.n3656 gnd.n3655 585
R2261 gnd.n3658 gnd.n3657 585
R2262 gnd.n3660 gnd.n3659 585
R2263 gnd.n3662 gnd.n3661 585
R2264 gnd.n3664 gnd.n3663 585
R2265 gnd.n3666 gnd.n3665 585
R2266 gnd.n3668 gnd.n3667 585
R2267 gnd.n3670 gnd.n3669 585
R2268 gnd.n3672 gnd.n3671 585
R2269 gnd.n3674 gnd.n3673 585
R2270 gnd.n3676 gnd.n3675 585
R2271 gnd.n3678 gnd.n3677 585
R2272 gnd.n3680 gnd.n3679 585
R2273 gnd.n3682 gnd.n3681 585
R2274 gnd.n3683 gnd.n2287 585
R2275 gnd.n3684 gnd.n2245 585
R2276 gnd.n3722 gnd.n2245 585
R2277 gnd.n3632 gnd.n2317 585
R2278 gnd.n3632 gnd.n3631 585
R2279 gnd.n3301 gnd.n2316 585
R2280 gnd.n2327 gnd.n2316 585
R2281 gnd.n3303 gnd.n3302 585
R2282 gnd.n3302 gnd.n2326 585
R2283 gnd.n3304 gnd.n2336 585
R2284 gnd.n3608 gnd.n2336 585
R2285 gnd.n3306 gnd.n3305 585
R2286 gnd.n3305 gnd.n2334 585
R2287 gnd.n3307 gnd.n2347 585
R2288 gnd.n3337 gnd.n2347 585
R2289 gnd.n3310 gnd.n3309 585
R2290 gnd.n3309 gnd.n3308 585
R2291 gnd.n3311 gnd.n2354 585
R2292 gnd.n3326 gnd.n2354 585
R2293 gnd.n3313 gnd.n3312 585
R2294 gnd.n3314 gnd.n3313 585
R2295 gnd.n2364 gnd.n2363 585
R2296 gnd.n2371 gnd.n2363 585
R2297 gnd.n3289 gnd.n3288 585
R2298 gnd.n3288 gnd.n3287 585
R2299 gnd.n2367 gnd.n2366 585
R2300 gnd.n2381 gnd.n2367 585
R2301 gnd.n3215 gnd.n3214 585
R2302 gnd.n3214 gnd.n2380 585
R2303 gnd.n3216 gnd.n2390 585
R2304 gnd.n3265 gnd.n2390 585
R2305 gnd.n3218 gnd.n3217 585
R2306 gnd.n3217 gnd.n2388 585
R2307 gnd.n3219 gnd.n2401 585
R2308 gnd.n3248 gnd.n2401 585
R2309 gnd.n3221 gnd.n3220 585
R2310 gnd.n3220 gnd.n2409 585
R2311 gnd.n3222 gnd.n2408 585
R2312 gnd.n3237 gnd.n2408 585
R2313 gnd.n3224 gnd.n3223 585
R2314 gnd.n3225 gnd.n3224 585
R2315 gnd.n2420 gnd.n2419 585
R2316 gnd.n2419 gnd.n2416 585
R2317 gnd.n3204 gnd.n3203 585
R2318 gnd.n3203 gnd.n3202 585
R2319 gnd.n2423 gnd.n2422 585
R2320 gnd.n2436 gnd.n2423 585
R2321 gnd.n3128 gnd.n3127 585
R2322 gnd.n3127 gnd.n2435 585
R2323 gnd.n3129 gnd.n2445 585
R2324 gnd.n3180 gnd.n2445 585
R2325 gnd.n3131 gnd.n3130 585
R2326 gnd.n3130 gnd.n2443 585
R2327 gnd.n3132 gnd.n2456 585
R2328 gnd.n3163 gnd.n2456 585
R2329 gnd.n3134 gnd.n3133 585
R2330 gnd.n3133 gnd.n2463 585
R2331 gnd.n3135 gnd.n2462 585
R2332 gnd.n3152 gnd.n2462 585
R2333 gnd.n3137 gnd.n3136 585
R2334 gnd.n3140 gnd.n3137 585
R2335 gnd.n2473 gnd.n2472 585
R2336 gnd.n2472 gnd.n2470 585
R2337 gnd.n2580 gnd.n2579 585
R2338 gnd.n3095 gnd.n2579 585
R2339 gnd.n2582 gnd.n2581 585
R2340 gnd.n2583 gnd.n2582 585
R2341 gnd.n2593 gnd.n2569 585
R2342 gnd.n3101 gnd.n2569 585
R2343 gnd.n2595 gnd.n2594 585
R2344 gnd.n2596 gnd.n2595 585
R2345 gnd.n2592 gnd.n2591 585
R2346 gnd.n2592 gnd.n2559 585
R2347 gnd.n2590 gnd.n2557 585
R2348 gnd.n3109 gnd.n2557 585
R2349 gnd.n2546 gnd.n2544 585
R2350 gnd.n3071 gnd.n2546 585
R2351 gnd.n3117 gnd.n3116 585
R2352 gnd.n3116 gnd.n3115 585
R2353 gnd.n2545 gnd.n2543 585
R2354 gnd.n2610 gnd.n2545 585
R2355 gnd.n3042 gnd.n2609 585
R2356 gnd.n3061 gnd.n2609 585
R2357 gnd.n3044 gnd.n3043 585
R2358 gnd.n3045 gnd.n3044 585
R2359 gnd.n2619 gnd.n2618 585
R2360 gnd.n2625 gnd.n2618 585
R2361 gnd.n3037 gnd.n3036 585
R2362 gnd.n3036 gnd.n3035 585
R2363 gnd.n2622 gnd.n2621 585
R2364 gnd.n2633 gnd.n2622 585
R2365 gnd.n2922 gnd.n2641 585
R2366 gnd.n3014 gnd.n2641 585
R2367 gnd.n2924 gnd.n2923 585
R2368 gnd.n2923 gnd.n2639 585
R2369 gnd.n2925 gnd.n2652 585
R2370 gnd.n3004 gnd.n2652 585
R2371 gnd.n2927 gnd.n2926 585
R2372 gnd.n2927 gnd.n2659 585
R2373 gnd.n2929 gnd.n2928 585
R2374 gnd.n2928 gnd.n2658 585
R2375 gnd.n2930 gnd.n2669 585
R2376 gnd.n2984 gnd.n2669 585
R2377 gnd.n2932 gnd.n2931 585
R2378 gnd.n2931 gnd.n2667 585
R2379 gnd.n2933 gnd.n2678 585
R2380 gnd.n2973 gnd.n2678 585
R2381 gnd.n2935 gnd.n2934 585
R2382 gnd.n2935 gnd.n2684 585
R2383 gnd.n2937 gnd.n2936 585
R2384 gnd.n2936 gnd.n2683 585
R2385 gnd.n2938 gnd.n2699 585
R2386 gnd.n2952 gnd.n2699 585
R2387 gnd.n2939 gnd.n2752 585
R2388 gnd.n2752 gnd.n2691 585
R2389 gnd.n2941 gnd.n2940 585
R2390 gnd.n2942 gnd.n2941 585
R2391 gnd.n2753 gnd.n2751 585
R2392 gnd.n2751 gnd.n2750 585
R2393 gnd.n2906 gnd.n2905 585
R2394 gnd.n2905 gnd.n2904 585
R2395 gnd.n2756 gnd.n2755 585
R2396 gnd.n2757 gnd.n2756 585
R2397 gnd.n2895 gnd.n2894 585
R2398 gnd.n2896 gnd.n2895 585
R2399 gnd.n2765 gnd.n2764 585
R2400 gnd.n2764 gnd.n2763 585
R2401 gnd.n2890 gnd.n2889 585
R2402 gnd.n2889 gnd.n2888 585
R2403 gnd.n2768 gnd.n2767 585
R2404 gnd.n2879 gnd.n2768 585
R2405 gnd.n2878 gnd.n2877 585
R2406 gnd.n2880 gnd.n2878 585
R2407 gnd.n2776 gnd.n2775 585
R2408 gnd.n2775 gnd.n2774 585
R2409 gnd.n201 gnd.n200 585
R2410 gnd.n204 gnd.n201 585
R2411 gnd.n7193 gnd.n7192 585
R2412 gnd.n7192 gnd.n7191 585
R2413 gnd.n7194 gnd.n196 585
R2414 gnd.n196 gnd.n195 585
R2415 gnd.n7196 gnd.n7195 585
R2416 gnd.n7197 gnd.n7196 585
R2417 gnd.n181 gnd.n180 585
R2418 gnd.n185 gnd.n181 585
R2419 gnd.n7205 gnd.n7204 585
R2420 gnd.n7204 gnd.n7203 585
R2421 gnd.n7206 gnd.n176 585
R2422 gnd.n182 gnd.n176 585
R2423 gnd.n7208 gnd.n7207 585
R2424 gnd.n7209 gnd.n7208 585
R2425 gnd.n163 gnd.n162 585
R2426 gnd.n166 gnd.n163 585
R2427 gnd.n7217 gnd.n7216 585
R2428 gnd.n7216 gnd.n7215 585
R2429 gnd.n7218 gnd.n158 585
R2430 gnd.n7041 gnd.n158 585
R2431 gnd.n7220 gnd.n7219 585
R2432 gnd.n7221 gnd.n7220 585
R2433 gnd.n143 gnd.n142 585
R2434 gnd.n147 gnd.n143 585
R2435 gnd.n7229 gnd.n7228 585
R2436 gnd.n7228 gnd.n7227 585
R2437 gnd.n7230 gnd.n138 585
R2438 gnd.n144 gnd.n138 585
R2439 gnd.n7232 gnd.n7231 585
R2440 gnd.n7233 gnd.n7232 585
R2441 gnd.n125 gnd.n124 585
R2442 gnd.n128 gnd.n125 585
R2443 gnd.n7241 gnd.n7240 585
R2444 gnd.n7240 gnd.n7239 585
R2445 gnd.n7242 gnd.n120 585
R2446 gnd.n120 gnd.n119 585
R2447 gnd.n7244 gnd.n7243 585
R2448 gnd.n7245 gnd.n7244 585
R2449 gnd.n105 gnd.n104 585
R2450 gnd.n109 gnd.n105 585
R2451 gnd.n7253 gnd.n7252 585
R2452 gnd.n7252 gnd.n7251 585
R2453 gnd.n7254 gnd.n99 585
R2454 gnd.n106 gnd.n99 585
R2455 gnd.n7256 gnd.n7255 585
R2456 gnd.n7257 gnd.n7256 585
R2457 gnd.n100 gnd.n98 585
R2458 gnd.n98 gnd.n86 585
R2459 gnd.n6896 gnd.n87 585
R2460 gnd.n7263 gnd.n87 585
R2461 gnd.n6895 gnd.n6894 585
R2462 gnd.n6894 gnd.n6893 585
R2463 gnd.n312 gnd.n311 585
R2464 gnd.n313 gnd.n312 585
R2465 gnd.n6887 gnd.n6886 585
R2466 gnd.n6886 gnd.n6885 585
R2467 gnd.n318 gnd.n317 585
R2468 gnd.n319 gnd.n318 585
R2469 gnd.n6873 gnd.n6872 585
R2470 gnd.n6874 gnd.n6873 585
R2471 gnd.n332 gnd.n331 585
R2472 gnd.n6865 gnd.n331 585
R2473 gnd.n6836 gnd.n6835 585
R2474 gnd.n6835 gnd.n336 585
R2475 gnd.n6837 gnd.n344 585
R2476 gnd.n6851 gnd.n344 585
R2477 gnd.n6838 gnd.n356 585
R2478 gnd.n356 gnd.n354 585
R2479 gnd.n6840 gnd.n6839 585
R2480 gnd.n6841 gnd.n6840 585
R2481 gnd.n357 gnd.n355 585
R2482 gnd.n6826 gnd.n355 585
R2483 gnd.n6802 gnd.n6801 585
R2484 gnd.n6801 gnd.n6800 585
R2485 gnd.n6803 gnd.n372 585
R2486 gnd.n6817 gnd.n372 585
R2487 gnd.n6804 gnd.n384 585
R2488 gnd.n6794 gnd.n384 585
R2489 gnd.n6806 gnd.n6805 585
R2490 gnd.n6807 gnd.n6806 585
R2491 gnd.n385 gnd.n383 585
R2492 gnd.n5502 gnd.n383 585
R2493 gnd.n1452 gnd.n1451 585
R2494 gnd.n5554 gnd.n1452 585
R2495 gnd.n5564 gnd.n5563 585
R2496 gnd.n5563 gnd.n5562 585
R2497 gnd.n5565 gnd.n1447 585
R2498 gnd.n5493 gnd.n1447 585
R2499 gnd.n5567 gnd.n5566 585
R2500 gnd.n5568 gnd.n5567 585
R2501 gnd.n1431 gnd.n1430 585
R2502 gnd.n5489 gnd.n1431 585
R2503 gnd.n5576 gnd.n5575 585
R2504 gnd.n5575 gnd.n5574 585
R2505 gnd.n5577 gnd.n1426 585
R2506 gnd.n5484 gnd.n1426 585
R2507 gnd.n5579 gnd.n5578 585
R2508 gnd.n5580 gnd.n5579 585
R2509 gnd.n1407 gnd.n1406 585
R2510 gnd.n5480 gnd.n1407 585
R2511 gnd.n5588 gnd.n5587 585
R2512 gnd.n5587 gnd.n5586 585
R2513 gnd.n5589 gnd.n1402 585
R2514 gnd.n5525 gnd.n1402 585
R2515 gnd.n5591 gnd.n5590 585
R2516 gnd.n5592 gnd.n5591 585
R2517 gnd.n1401 gnd.n1241 585
R2518 gnd.n5759 gnd.n1242 585
R2519 gnd.n5758 gnd.n1243 585
R2520 gnd.n1318 gnd.n1244 585
R2521 gnd.n5751 gnd.n1250 585
R2522 gnd.n5750 gnd.n1251 585
R2523 gnd.n1321 gnd.n1252 585
R2524 gnd.n5743 gnd.n1258 585
R2525 gnd.n5742 gnd.n1259 585
R2526 gnd.n1323 gnd.n1260 585
R2527 gnd.n5735 gnd.n1266 585
R2528 gnd.n5734 gnd.n1267 585
R2529 gnd.n1326 gnd.n1268 585
R2530 gnd.n5727 gnd.n1274 585
R2531 gnd.n5726 gnd.n1275 585
R2532 gnd.n1328 gnd.n1276 585
R2533 gnd.n5719 gnd.n1284 585
R2534 gnd.n5718 gnd.n5715 585
R2535 gnd.n1287 gnd.n1285 585
R2536 gnd.n5713 gnd.n1287 585
R2537 gnd.n7023 gnd.n7022 585
R2538 gnd.n7016 gnd.n6969 585
R2539 gnd.n7018 gnd.n7017 585
R2540 gnd.n7015 gnd.n7014 585
R2541 gnd.n7013 gnd.n7012 585
R2542 gnd.n7006 gnd.n6971 585
R2543 gnd.n7008 gnd.n7007 585
R2544 gnd.n7005 gnd.n7004 585
R2545 gnd.n7003 gnd.n7002 585
R2546 gnd.n6996 gnd.n6973 585
R2547 gnd.n6998 gnd.n6997 585
R2548 gnd.n6995 gnd.n6994 585
R2549 gnd.n6993 gnd.n6992 585
R2550 gnd.n6986 gnd.n6975 585
R2551 gnd.n6988 gnd.n6987 585
R2552 gnd.n6985 gnd.n6984 585
R2553 gnd.n6983 gnd.n6982 585
R2554 gnd.n6979 gnd.n6978 585
R2555 gnd.n6977 gnd.n211 585
R2556 gnd.n7183 gnd.n211 585
R2557 gnd.n7025 gnd.n7024 585
R2558 gnd.n7024 gnd.n204 585
R2559 gnd.n7026 gnd.n203 585
R2560 gnd.n7191 gnd.n203 585
R2561 gnd.n7028 gnd.n7027 585
R2562 gnd.n7027 gnd.n195 585
R2563 gnd.n7029 gnd.n194 585
R2564 gnd.n7197 gnd.n194 585
R2565 gnd.n7031 gnd.n7030 585
R2566 gnd.n7030 gnd.n185 585
R2567 gnd.n7032 gnd.n184 585
R2568 gnd.n7203 gnd.n184 585
R2569 gnd.n7034 gnd.n7033 585
R2570 gnd.n7033 gnd.n182 585
R2571 gnd.n7035 gnd.n175 585
R2572 gnd.n7209 gnd.n175 585
R2573 gnd.n7037 gnd.n7036 585
R2574 gnd.n7036 gnd.n166 585
R2575 gnd.n7038 gnd.n165 585
R2576 gnd.n7215 gnd.n165 585
R2577 gnd.n7040 gnd.n7039 585
R2578 gnd.n7041 gnd.n7040 585
R2579 gnd.n6923 gnd.n156 585
R2580 gnd.n7221 gnd.n156 585
R2581 gnd.n6953 gnd.n6952 585
R2582 gnd.n6952 gnd.n147 585
R2583 gnd.n6951 gnd.n146 585
R2584 gnd.n7227 gnd.n146 585
R2585 gnd.n6950 gnd.n6949 585
R2586 gnd.n6949 gnd.n144 585
R2587 gnd.n6925 gnd.n137 585
R2588 gnd.n7233 gnd.n137 585
R2589 gnd.n6945 gnd.n6944 585
R2590 gnd.n6944 gnd.n128 585
R2591 gnd.n6943 gnd.n127 585
R2592 gnd.n7239 gnd.n127 585
R2593 gnd.n6942 gnd.n6941 585
R2594 gnd.n6941 gnd.n119 585
R2595 gnd.n6927 gnd.n118 585
R2596 gnd.n7245 gnd.n118 585
R2597 gnd.n6937 gnd.n6936 585
R2598 gnd.n6936 gnd.n109 585
R2599 gnd.n6935 gnd.n108 585
R2600 gnd.n7251 gnd.n108 585
R2601 gnd.n6934 gnd.n6933 585
R2602 gnd.n6933 gnd.n106 585
R2603 gnd.n6929 gnd.n97 585
R2604 gnd.n7257 gnd.n97 585
R2605 gnd.n84 gnd.n83 585
R2606 gnd.n86 gnd.n84 585
R2607 gnd.n7265 gnd.n7264 585
R2608 gnd.n7264 gnd.n7263 585
R2609 gnd.n7266 gnd.n82 585
R2610 gnd.n6893 gnd.n82 585
R2611 gnd.n321 gnd.n81 585
R2612 gnd.n321 gnd.n313 585
R2613 gnd.n6858 gnd.n322 585
R2614 gnd.n6885 gnd.n322 585
R2615 gnd.n6859 gnd.n6857 585
R2616 gnd.n6857 gnd.n319 585
R2617 gnd.n339 gnd.n330 585
R2618 gnd.n6874 gnd.n330 585
R2619 gnd.n6864 gnd.n6863 585
R2620 gnd.n6865 gnd.n6864 585
R2621 gnd.n338 gnd.n337 585
R2622 gnd.n337 gnd.n336 585
R2623 gnd.n6853 gnd.n6852 585
R2624 gnd.n6852 gnd.n6851 585
R2625 gnd.n342 gnd.n341 585
R2626 gnd.n354 gnd.n342 585
R2627 gnd.n366 gnd.n353 585
R2628 gnd.n6841 gnd.n353 585
R2629 gnd.n6825 gnd.n6824 585
R2630 gnd.n6826 gnd.n6825 585
R2631 gnd.n365 gnd.n364 585
R2632 gnd.n6800 gnd.n364 585
R2633 gnd.n6819 gnd.n6818 585
R2634 gnd.n6818 gnd.n6817 585
R2635 gnd.n369 gnd.n368 585
R2636 gnd.n6794 gnd.n369 585
R2637 gnd.n5505 gnd.n381 585
R2638 gnd.n6807 gnd.n381 585
R2639 gnd.n5506 gnd.n5503 585
R2640 gnd.n5503 gnd.n5502 585
R2641 gnd.n5507 gnd.n1458 585
R2642 gnd.n5554 gnd.n1458 585
R2643 gnd.n5475 gnd.n1455 585
R2644 gnd.n5562 gnd.n1455 585
R2645 gnd.n5511 gnd.n5474 585
R2646 gnd.n5493 gnd.n5474 585
R2647 gnd.n5512 gnd.n1445 585
R2648 gnd.n5568 gnd.n1445 585
R2649 gnd.n5513 gnd.n5473 585
R2650 gnd.n5489 gnd.n5473 585
R2651 gnd.n5471 gnd.n1434 585
R2652 gnd.n5574 gnd.n1434 585
R2653 gnd.n5517 gnd.n5470 585
R2654 gnd.n5484 gnd.n5470 585
R2655 gnd.n5518 gnd.n1424 585
R2656 gnd.n5580 gnd.n1424 585
R2657 gnd.n5519 gnd.n5469 585
R2658 gnd.n5480 gnd.n5469 585
R2659 gnd.n1474 gnd.n1409 585
R2660 gnd.n5586 gnd.n1409 585
R2661 gnd.n5524 gnd.n5523 585
R2662 gnd.n5525 gnd.n5524 585
R2663 gnd.n1473 gnd.n1399 585
R2664 gnd.n5592 gnd.n1399 585
R2665 gnd.n3617 gnd.n2267 585
R2666 gnd.n2319 gnd.n2267 585
R2667 gnd.n3618 gnd.n2329 585
R2668 gnd.n2329 gnd.n2318 585
R2669 gnd.n3620 gnd.n3619 585
R2670 gnd.n3621 gnd.n3620 585
R2671 gnd.n2330 gnd.n2328 585
R2672 gnd.n2337 gnd.n2328 585
R2673 gnd.n3611 gnd.n3610 585
R2674 gnd.n3610 gnd.n3609 585
R2675 gnd.n2333 gnd.n2332 585
R2676 gnd.n3336 gnd.n2333 585
R2677 gnd.n3322 gnd.n2356 585
R2678 gnd.n2356 gnd.n2346 585
R2679 gnd.n3324 gnd.n3323 585
R2680 gnd.n3325 gnd.n3324 585
R2681 gnd.n2357 gnd.n2355 585
R2682 gnd.n2355 gnd.n2353 585
R2683 gnd.n3317 gnd.n3316 585
R2684 gnd.n3316 gnd.n3315 585
R2685 gnd.n2360 gnd.n2359 585
R2686 gnd.n2369 gnd.n2360 585
R2687 gnd.n3273 gnd.n2383 585
R2688 gnd.n2383 gnd.n2368 585
R2689 gnd.n3275 gnd.n3274 585
R2690 gnd.n3276 gnd.n3275 585
R2691 gnd.n2384 gnd.n2382 585
R2692 gnd.n2391 gnd.n2382 585
R2693 gnd.n3268 gnd.n3267 585
R2694 gnd.n3267 gnd.n3266 585
R2695 gnd.n2387 gnd.n2386 585
R2696 gnd.n3247 gnd.n2387 585
R2697 gnd.n3233 gnd.n2411 585
R2698 gnd.n2411 gnd.n2400 585
R2699 gnd.n3235 gnd.n3234 585
R2700 gnd.n3236 gnd.n3235 585
R2701 gnd.n2412 gnd.n2410 585
R2702 gnd.n2410 gnd.n2407 585
R2703 gnd.n3228 gnd.n3227 585
R2704 gnd.n3227 gnd.n3226 585
R2705 gnd.n2415 gnd.n2414 585
R2706 gnd.n2425 gnd.n2415 585
R2707 gnd.n3188 gnd.n2438 585
R2708 gnd.n2438 gnd.n2424 585
R2709 gnd.n3190 gnd.n3189 585
R2710 gnd.n3191 gnd.n3190 585
R2711 gnd.n2439 gnd.n2437 585
R2712 gnd.n2446 gnd.n2437 585
R2713 gnd.n3183 gnd.n3182 585
R2714 gnd.n3182 gnd.n3181 585
R2715 gnd.n2442 gnd.n2441 585
R2716 gnd.n3162 gnd.n2442 585
R2717 gnd.n3148 gnd.n2465 585
R2718 gnd.n2465 gnd.n2455 585
R2719 gnd.n3150 gnd.n3149 585
R2720 gnd.n3151 gnd.n3150 585
R2721 gnd.n2466 gnd.n2464 585
R2722 gnd.n3139 gnd.n2464 585
R2723 gnd.n3143 gnd.n3142 585
R2724 gnd.n3142 gnd.n3141 585
R2725 gnd.n2469 gnd.n2468 585
R2726 gnd.n3094 gnd.n2469 585
R2727 gnd.n2587 gnd.n2586 585
R2728 gnd.n2588 gnd.n2587 585
R2729 gnd.n2567 gnd.n2566 585
R2730 gnd.n2570 gnd.n2567 585
R2731 gnd.n3104 gnd.n3103 585
R2732 gnd.n3103 gnd.n3102 585
R2733 gnd.n3105 gnd.n2561 585
R2734 gnd.n2597 gnd.n2561 585
R2735 gnd.n3107 gnd.n3106 585
R2736 gnd.n3108 gnd.n3107 585
R2737 gnd.n2562 gnd.n2560 585
R2738 gnd.n3072 gnd.n2560 585
R2739 gnd.n3056 gnd.n3055 585
R2740 gnd.n3055 gnd.n2548 585
R2741 gnd.n3057 gnd.n2612 585
R2742 gnd.n2612 gnd.n2547 585
R2743 gnd.n3059 gnd.n3058 585
R2744 gnd.n3060 gnd.n3059 585
R2745 gnd.n2613 gnd.n2611 585
R2746 gnd.n2611 gnd.n2608 585
R2747 gnd.n3048 gnd.n3047 585
R2748 gnd.n3047 gnd.n3046 585
R2749 gnd.n2616 gnd.n2615 585
R2750 gnd.n2623 gnd.n2616 585
R2751 gnd.n3022 gnd.n3021 585
R2752 gnd.n3023 gnd.n3022 585
R2753 gnd.n2635 gnd.n2634 585
R2754 gnd.n2642 gnd.n2634 585
R2755 gnd.n3017 gnd.n3016 585
R2756 gnd.n3016 gnd.n3015 585
R2757 gnd.n2638 gnd.n2637 585
R2758 gnd.n3005 gnd.n2638 585
R2759 gnd.n2992 gnd.n2662 585
R2760 gnd.n2662 gnd.n2661 585
R2761 gnd.n2994 gnd.n2993 585
R2762 gnd.n2995 gnd.n2994 585
R2763 gnd.n2663 gnd.n2660 585
R2764 gnd.n2670 gnd.n2660 585
R2765 gnd.n2987 gnd.n2986 585
R2766 gnd.n2986 gnd.n2985 585
R2767 gnd.n2666 gnd.n2665 585
R2768 gnd.n2974 gnd.n2666 585
R2769 gnd.n2961 gnd.n2687 585
R2770 gnd.n2687 gnd.n2686 585
R2771 gnd.n2963 gnd.n2962 585
R2772 gnd.n2964 gnd.n2963 585
R2773 gnd.n2957 gnd.n2685 585
R2774 gnd.n2956 gnd.n2955 585
R2775 gnd.n2690 gnd.n2689 585
R2776 gnd.n2953 gnd.n2690 585
R2777 gnd.n2712 gnd.n2711 585
R2778 gnd.n2715 gnd.n2714 585
R2779 gnd.n2713 gnd.n2708 585
R2780 gnd.n2720 gnd.n2719 585
R2781 gnd.n2722 gnd.n2721 585
R2782 gnd.n2725 gnd.n2724 585
R2783 gnd.n2723 gnd.n2706 585
R2784 gnd.n2730 gnd.n2729 585
R2785 gnd.n2732 gnd.n2731 585
R2786 gnd.n2735 gnd.n2734 585
R2787 gnd.n2733 gnd.n2704 585
R2788 gnd.n2740 gnd.n2739 585
R2789 gnd.n2744 gnd.n2741 585
R2790 gnd.n2745 gnd.n2682 585
R2791 gnd.n3623 gnd.n2282 585
R2792 gnd.n3690 gnd.n3689 585
R2793 gnd.n3692 gnd.n3691 585
R2794 gnd.n3694 gnd.n3693 585
R2795 gnd.n3696 gnd.n3695 585
R2796 gnd.n3698 gnd.n3697 585
R2797 gnd.n3700 gnd.n3699 585
R2798 gnd.n3702 gnd.n3701 585
R2799 gnd.n3704 gnd.n3703 585
R2800 gnd.n3706 gnd.n3705 585
R2801 gnd.n3708 gnd.n3707 585
R2802 gnd.n3710 gnd.n3709 585
R2803 gnd.n3712 gnd.n3711 585
R2804 gnd.n3715 gnd.n3714 585
R2805 gnd.n3713 gnd.n2270 585
R2806 gnd.n3719 gnd.n2268 585
R2807 gnd.n3721 gnd.n3720 585
R2808 gnd.n3722 gnd.n3721 585
R2809 gnd.n3624 gnd.n2324 585
R2810 gnd.n3624 gnd.n2319 585
R2811 gnd.n3626 gnd.n3625 585
R2812 gnd.n3625 gnd.n2318 585
R2813 gnd.n3622 gnd.n2323 585
R2814 gnd.n3622 gnd.n3621 585
R2815 gnd.n3601 gnd.n2325 585
R2816 gnd.n2337 gnd.n2325 585
R2817 gnd.n3600 gnd.n2335 585
R2818 gnd.n3609 gnd.n2335 585
R2819 gnd.n3335 gnd.n2342 585
R2820 gnd.n3336 gnd.n3335 585
R2821 gnd.n3334 gnd.n3333 585
R2822 gnd.n3334 gnd.n2346 585
R2823 gnd.n3332 gnd.n2348 585
R2824 gnd.n3325 gnd.n2348 585
R2825 gnd.n2361 gnd.n2349 585
R2826 gnd.n2361 gnd.n2353 585
R2827 gnd.n3281 gnd.n2362 585
R2828 gnd.n3315 gnd.n2362 585
R2829 gnd.n3280 gnd.n3279 585
R2830 gnd.n3279 gnd.n2369 585
R2831 gnd.n3278 gnd.n2377 585
R2832 gnd.n3278 gnd.n2368 585
R2833 gnd.n3277 gnd.n2379 585
R2834 gnd.n3277 gnd.n3276 585
R2835 gnd.n3256 gnd.n2378 585
R2836 gnd.n2391 gnd.n2378 585
R2837 gnd.n3255 gnd.n2389 585
R2838 gnd.n3266 gnd.n2389 585
R2839 gnd.n3246 gnd.n2396 585
R2840 gnd.n3247 gnd.n3246 585
R2841 gnd.n3245 gnd.n3244 585
R2842 gnd.n3245 gnd.n2400 585
R2843 gnd.n3243 gnd.n2402 585
R2844 gnd.n3236 gnd.n2402 585
R2845 gnd.n2417 gnd.n2403 585
R2846 gnd.n2417 gnd.n2407 585
R2847 gnd.n3196 gnd.n2418 585
R2848 gnd.n3226 gnd.n2418 585
R2849 gnd.n3195 gnd.n3194 585
R2850 gnd.n3194 gnd.n2425 585
R2851 gnd.n3193 gnd.n2432 585
R2852 gnd.n3193 gnd.n2424 585
R2853 gnd.n3192 gnd.n2434 585
R2854 gnd.n3192 gnd.n3191 585
R2855 gnd.n3171 gnd.n2433 585
R2856 gnd.n2446 gnd.n2433 585
R2857 gnd.n3170 gnd.n2444 585
R2858 gnd.n3181 gnd.n2444 585
R2859 gnd.n3161 gnd.n2451 585
R2860 gnd.n3162 gnd.n3161 585
R2861 gnd.n3160 gnd.n3159 585
R2862 gnd.n3160 gnd.n2455 585
R2863 gnd.n3158 gnd.n2457 585
R2864 gnd.n3151 gnd.n2457 585
R2865 gnd.n3138 gnd.n2458 585
R2866 gnd.n3139 gnd.n3138 585
R2867 gnd.n3091 gnd.n2471 585
R2868 gnd.n3141 gnd.n2471 585
R2869 gnd.n3093 gnd.n3092 585
R2870 gnd.n3094 gnd.n3093 585
R2871 gnd.n3086 gnd.n2589 585
R2872 gnd.n2589 gnd.n2588 585
R2873 gnd.n3084 gnd.n3083 585
R2874 gnd.n3083 gnd.n2570 585
R2875 gnd.n3081 gnd.n2568 585
R2876 gnd.n3102 gnd.n2568 585
R2877 gnd.n2599 gnd.n2598 585
R2878 gnd.n2598 gnd.n2597 585
R2879 gnd.n3075 gnd.n2558 585
R2880 gnd.n3108 gnd.n2558 585
R2881 gnd.n3074 gnd.n3073 585
R2882 gnd.n3073 gnd.n3072 585
R2883 gnd.n3070 gnd.n2601 585
R2884 gnd.n3070 gnd.n2548 585
R2885 gnd.n3069 gnd.n3068 585
R2886 gnd.n3069 gnd.n2547 585
R2887 gnd.n2604 gnd.n2603 585
R2888 gnd.n3060 gnd.n2603 585
R2889 gnd.n3028 gnd.n3027 585
R2890 gnd.n3027 gnd.n2608 585
R2891 gnd.n3029 gnd.n2617 585
R2892 gnd.n3046 gnd.n2617 585
R2893 gnd.n3026 gnd.n3025 585
R2894 gnd.n3025 gnd.n2623 585
R2895 gnd.n3024 gnd.n2631 585
R2896 gnd.n3024 gnd.n3023 585
R2897 gnd.n3009 gnd.n2632 585
R2898 gnd.n2642 gnd.n2632 585
R2899 gnd.n3008 gnd.n2640 585
R2900 gnd.n3015 gnd.n2640 585
R2901 gnd.n3007 gnd.n3006 585
R2902 gnd.n3006 gnd.n3005 585
R2903 gnd.n2651 gnd.n2648 585
R2904 gnd.n2661 gnd.n2651 585
R2905 gnd.n2997 gnd.n2996 585
R2906 gnd.n2996 gnd.n2995 585
R2907 gnd.n2657 gnd.n2656 585
R2908 gnd.n2670 gnd.n2657 585
R2909 gnd.n2977 gnd.n2668 585
R2910 gnd.n2985 gnd.n2668 585
R2911 gnd.n2976 gnd.n2975 585
R2912 gnd.n2975 gnd.n2974 585
R2913 gnd.n2677 gnd.n2675 585
R2914 gnd.n2686 gnd.n2677 585
R2915 gnd.n2966 gnd.n2965 585
R2916 gnd.n2965 gnd.n2964 585
R2917 gnd.n5399 gnd.n5398 585
R2918 gnd.n5398 gnd.n1526 585
R2919 gnd.n5400 gnd.n1540 585
R2920 gnd.n1540 gnd.n1538 585
R2921 gnd.n5402 gnd.n5401 585
R2922 gnd.n5403 gnd.n5402 585
R2923 gnd.n1541 gnd.n1539 585
R2924 gnd.n5274 gnd.n1539 585
R2925 gnd.n1643 gnd.n1642 585
R2926 gnd.n1642 gnd.n1618 585
R2927 gnd.n5246 gnd.n1644 585
R2928 gnd.n5246 gnd.n5245 585
R2929 gnd.n5247 gnd.n1641 585
R2930 gnd.n5247 gnd.n1626 585
R2931 gnd.n5249 gnd.n5248 585
R2932 gnd.n5248 gnd.n1625 585
R2933 gnd.n5250 gnd.n1639 585
R2934 gnd.n5238 gnd.n1639 585
R2935 gnd.n5252 gnd.n5251 585
R2936 gnd.n5253 gnd.n5252 585
R2937 gnd.n1640 gnd.n1638 585
R2938 gnd.n1638 gnd.n1634 585
R2939 gnd.n5231 gnd.n5230 585
R2940 gnd.n5232 gnd.n5231 585
R2941 gnd.n5229 gnd.n1650 585
R2942 gnd.n1656 gnd.n1650 585
R2943 gnd.n5228 gnd.n5227 585
R2944 gnd.n5227 gnd.n5226 585
R2945 gnd.n1652 gnd.n1651 585
R2946 gnd.n1653 gnd.n1652 585
R2947 gnd.n5216 gnd.n5215 585
R2948 gnd.n5217 gnd.n5216 585
R2949 gnd.n5214 gnd.n1667 585
R2950 gnd.n1667 gnd.n1663 585
R2951 gnd.n5213 gnd.n5212 585
R2952 gnd.n5212 gnd.n5211 585
R2953 gnd.n1669 gnd.n1668 585
R2954 gnd.n1675 gnd.n1669 585
R2955 gnd.n5198 gnd.n5197 585
R2956 gnd.n5199 gnd.n5198 585
R2957 gnd.n5196 gnd.n1678 585
R2958 gnd.n1684 gnd.n1678 585
R2959 gnd.n5195 gnd.n5194 585
R2960 gnd.n5194 gnd.n5193 585
R2961 gnd.n1680 gnd.n1679 585
R2962 gnd.n1695 gnd.n1680 585
R2963 gnd.n5170 gnd.n1692 585
R2964 gnd.n5182 gnd.n1692 585
R2965 gnd.n5171 gnd.n1703 585
R2966 gnd.n1703 gnd.n1691 585
R2967 gnd.n5173 gnd.n5172 585
R2968 gnd.n5174 gnd.n5173 585
R2969 gnd.n5169 gnd.n1702 585
R2970 gnd.n5165 gnd.n1702 585
R2971 gnd.n5168 gnd.n5167 585
R2972 gnd.n5167 gnd.n5166 585
R2973 gnd.n1705 gnd.n1704 585
R2974 gnd.n1711 gnd.n1705 585
R2975 gnd.n5158 gnd.n5157 585
R2976 gnd.n5159 gnd.n5158 585
R2977 gnd.n5156 gnd.n1713 585
R2978 gnd.n1713 gnd.n1710 585
R2979 gnd.n5155 gnd.n5154 585
R2980 gnd.n5154 gnd.n5153 585
R2981 gnd.n1715 gnd.n1714 585
R2982 gnd.n1727 gnd.n1715 585
R2983 gnd.n5134 gnd.n5133 585
R2984 gnd.n5135 gnd.n5134 585
R2985 gnd.n5132 gnd.n1728 585
R2986 gnd.n5127 gnd.n1728 585
R2987 gnd.n5131 gnd.n5130 585
R2988 gnd.n5130 gnd.n5129 585
R2989 gnd.n1730 gnd.n1729 585
R2990 gnd.n1731 gnd.n1730 585
R2991 gnd.n5115 gnd.n5114 585
R2992 gnd.n5116 gnd.n5115 585
R2993 gnd.n5113 gnd.n1738 585
R2994 gnd.n5109 gnd.n1738 585
R2995 gnd.n5112 gnd.n5111 585
R2996 gnd.n5111 gnd.n5110 585
R2997 gnd.n1740 gnd.n1739 585
R2998 gnd.n5097 gnd.n1740 585
R2999 gnd.n5086 gnd.n1758 585
R3000 gnd.n1758 gnd.n1756 585
R3001 gnd.n5088 gnd.n5087 585
R3002 gnd.n5089 gnd.n5088 585
R3003 gnd.n5085 gnd.n1757 585
R3004 gnd.n1763 gnd.n1757 585
R3005 gnd.n5084 gnd.n5083 585
R3006 gnd.n5083 gnd.n5082 585
R3007 gnd.n1760 gnd.n1759 585
R3008 gnd.n5059 gnd.n1760 585
R3009 gnd.n5071 gnd.n5070 585
R3010 gnd.n5072 gnd.n5071 585
R3011 gnd.n5069 gnd.n1773 585
R3012 gnd.n1773 gnd.n1769 585
R3013 gnd.n5068 gnd.n5067 585
R3014 gnd.n5067 gnd.n5066 585
R3015 gnd.n1775 gnd.n1774 585
R3016 gnd.n1776 gnd.n1775 585
R3017 gnd.n5053 gnd.n5052 585
R3018 gnd.n5054 gnd.n5053 585
R3019 gnd.n5051 gnd.n1785 585
R3020 gnd.n5047 gnd.n1785 585
R3021 gnd.n5050 gnd.n5049 585
R3022 gnd.n5049 gnd.n5048 585
R3023 gnd.n1787 gnd.n1786 585
R3024 gnd.n1793 gnd.n1787 585
R3025 gnd.n5040 gnd.n5039 585
R3026 gnd.n5041 gnd.n5040 585
R3027 gnd.n5038 gnd.n1796 585
R3028 gnd.n1796 gnd.n1792 585
R3029 gnd.n5037 gnd.n5036 585
R3030 gnd.n5036 gnd.n5035 585
R3031 gnd.n1798 gnd.n1797 585
R3032 gnd.n1810 gnd.n1798 585
R3033 gnd.n5013 gnd.n5012 585
R3034 gnd.n5014 gnd.n5013 585
R3035 gnd.n5011 gnd.n1811 585
R3036 gnd.n5005 gnd.n1811 585
R3037 gnd.n5010 gnd.n5009 585
R3038 gnd.n5009 gnd.n5008 585
R3039 gnd.n1813 gnd.n1812 585
R3040 gnd.n1814 gnd.n1813 585
R3041 gnd.n4993 gnd.n4992 585
R3042 gnd.n4994 gnd.n4993 585
R3043 gnd.n4991 gnd.n1820 585
R3044 gnd.n4987 gnd.n1820 585
R3045 gnd.n4990 gnd.n4989 585
R3046 gnd.n4989 gnd.n4988 585
R3047 gnd.n1822 gnd.n1821 585
R3048 gnd.n4974 gnd.n1822 585
R3049 gnd.n4963 gnd.n1839 585
R3050 gnd.n1839 gnd.n1837 585
R3051 gnd.n4965 gnd.n4964 585
R3052 gnd.n4966 gnd.n4965 585
R3053 gnd.n4962 gnd.n1838 585
R3054 gnd.n1844 gnd.n1838 585
R3055 gnd.n4961 gnd.n4960 585
R3056 gnd.n4960 gnd.n4959 585
R3057 gnd.n1841 gnd.n1840 585
R3058 gnd.n4935 gnd.n1841 585
R3059 gnd.n4947 gnd.n4946 585
R3060 gnd.n4948 gnd.n4947 585
R3061 gnd.n4945 gnd.n1853 585
R3062 gnd.n1857 gnd.n1853 585
R3063 gnd.n4944 gnd.n4943 585
R3064 gnd.n4943 gnd.n4942 585
R3065 gnd.n1855 gnd.n1854 585
R3066 gnd.n1863 gnd.n1855 585
R3067 gnd.n4929 gnd.n4928 585
R3068 gnd.n4930 gnd.n4929 585
R3069 gnd.n4927 gnd.n1865 585
R3070 gnd.n4923 gnd.n1865 585
R3071 gnd.n4926 gnd.n4925 585
R3072 gnd.n4925 gnd.n4924 585
R3073 gnd.n1867 gnd.n1866 585
R3074 gnd.n1874 gnd.n1867 585
R3075 gnd.n4916 gnd.n4915 585
R3076 gnd.n4917 gnd.n4916 585
R3077 gnd.n4914 gnd.n1876 585
R3078 gnd.n1876 gnd.n1873 585
R3079 gnd.n4913 gnd.n4912 585
R3080 gnd.n4912 gnd.n4911 585
R3081 gnd.n1878 gnd.n1877 585
R3082 gnd.n1890 gnd.n1878 585
R3083 gnd.n4889 gnd.n4888 585
R3084 gnd.n4890 gnd.n4889 585
R3085 gnd.n4887 gnd.n1891 585
R3086 gnd.n4882 gnd.n1891 585
R3087 gnd.n4886 gnd.n4885 585
R3088 gnd.n4885 gnd.n4884 585
R3089 gnd.n1893 gnd.n1892 585
R3090 gnd.n4872 gnd.n1893 585
R3091 gnd.n4861 gnd.n4860 585
R3092 gnd.n4862 gnd.n4861 585
R3093 gnd.n4859 gnd.n1901 585
R3094 gnd.n1901 gnd.n1899 585
R3095 gnd.n4858 gnd.n4857 585
R3096 gnd.n4857 gnd.n4856 585
R3097 gnd.n1903 gnd.n1902 585
R3098 gnd.n1903 gnd.n1125 585
R3099 gnd.n4848 gnd.n4847 585
R3100 gnd.n4849 gnd.n4848 585
R3101 gnd.n4846 gnd.n4843 585
R3102 gnd.n4843 gnd.n4842 585
R3103 gnd.n4845 gnd.n4844 585
R3104 gnd.n4844 gnd.n1114 585
R3105 gnd.n1109 gnd.n1108 585
R3106 gnd.n5898 gnd.n1109 585
R3107 gnd.n5901 gnd.n5900 585
R3108 gnd.n5900 gnd.n5899 585
R3109 gnd.n5902 gnd.n1087 585
R3110 gnd.n1973 gnd.n1087 585
R3111 gnd.n5967 gnd.n5966 585
R3112 gnd.n5965 gnd.n1086 585
R3113 gnd.n5964 gnd.n1085 585
R3114 gnd.n5969 gnd.n1085 585
R3115 gnd.n5963 gnd.n5962 585
R3116 gnd.n5961 gnd.n5960 585
R3117 gnd.n5959 gnd.n5958 585
R3118 gnd.n5957 gnd.n5956 585
R3119 gnd.n5955 gnd.n5954 585
R3120 gnd.n5953 gnd.n5952 585
R3121 gnd.n5951 gnd.n5950 585
R3122 gnd.n5949 gnd.n5948 585
R3123 gnd.n5947 gnd.n5946 585
R3124 gnd.n5945 gnd.n5944 585
R3125 gnd.n5943 gnd.n5942 585
R3126 gnd.n5941 gnd.n5940 585
R3127 gnd.n5939 gnd.n5938 585
R3128 gnd.n5937 gnd.n5936 585
R3129 gnd.n5935 gnd.n5934 585
R3130 gnd.n5933 gnd.n5932 585
R3131 gnd.n5931 gnd.n5930 585
R3132 gnd.n5929 gnd.n5928 585
R3133 gnd.n5927 gnd.n5926 585
R3134 gnd.n5925 gnd.n5924 585
R3135 gnd.n5923 gnd.n5922 585
R3136 gnd.n5921 gnd.n5920 585
R3137 gnd.n5919 gnd.n5918 585
R3138 gnd.n5917 gnd.n5916 585
R3139 gnd.n5915 gnd.n5914 585
R3140 gnd.n5913 gnd.n5912 585
R3141 gnd.n5911 gnd.n5910 585
R3142 gnd.n5909 gnd.n5908 585
R3143 gnd.n5907 gnd.n1049 585
R3144 gnd.n5972 gnd.n5971 585
R3145 gnd.n1051 gnd.n1048 585
R3146 gnd.n1911 gnd.n1910 585
R3147 gnd.n1913 gnd.n1912 585
R3148 gnd.n1916 gnd.n1915 585
R3149 gnd.n1918 gnd.n1917 585
R3150 gnd.n1920 gnd.n1919 585
R3151 gnd.n1922 gnd.n1921 585
R3152 gnd.n1924 gnd.n1923 585
R3153 gnd.n1926 gnd.n1925 585
R3154 gnd.n1928 gnd.n1927 585
R3155 gnd.n1930 gnd.n1929 585
R3156 gnd.n1932 gnd.n1931 585
R3157 gnd.n1934 gnd.n1933 585
R3158 gnd.n1936 gnd.n1935 585
R3159 gnd.n1938 gnd.n1937 585
R3160 gnd.n1940 gnd.n1939 585
R3161 gnd.n1942 gnd.n1941 585
R3162 gnd.n1944 gnd.n1943 585
R3163 gnd.n1946 gnd.n1945 585
R3164 gnd.n1948 gnd.n1947 585
R3165 gnd.n1950 gnd.n1949 585
R3166 gnd.n1952 gnd.n1951 585
R3167 gnd.n1954 gnd.n1953 585
R3168 gnd.n1956 gnd.n1955 585
R3169 gnd.n1958 gnd.n1957 585
R3170 gnd.n1960 gnd.n1959 585
R3171 gnd.n1962 gnd.n1961 585
R3172 gnd.n1964 gnd.n1963 585
R3173 gnd.n1966 gnd.n1965 585
R3174 gnd.n1968 gnd.n1967 585
R3175 gnd.n1970 gnd.n1969 585
R3176 gnd.n1972 gnd.n1971 585
R3177 gnd.n5282 gnd.n5281 585
R3178 gnd.n5283 gnd.n1613 585
R3179 gnd.n5285 gnd.n5284 585
R3180 gnd.n5287 gnd.n1611 585
R3181 gnd.n5289 gnd.n5288 585
R3182 gnd.n5290 gnd.n1610 585
R3183 gnd.n5292 gnd.n5291 585
R3184 gnd.n5294 gnd.n1608 585
R3185 gnd.n5296 gnd.n5295 585
R3186 gnd.n5297 gnd.n1607 585
R3187 gnd.n5299 gnd.n5298 585
R3188 gnd.n5301 gnd.n1605 585
R3189 gnd.n5303 gnd.n5302 585
R3190 gnd.n5304 gnd.n1604 585
R3191 gnd.n5306 gnd.n5305 585
R3192 gnd.n5308 gnd.n1602 585
R3193 gnd.n5310 gnd.n5309 585
R3194 gnd.n5311 gnd.n1601 585
R3195 gnd.n5313 gnd.n5312 585
R3196 gnd.n5315 gnd.n1599 585
R3197 gnd.n5317 gnd.n5316 585
R3198 gnd.n5318 gnd.n1598 585
R3199 gnd.n5320 gnd.n5319 585
R3200 gnd.n5322 gnd.n1596 585
R3201 gnd.n5324 gnd.n5323 585
R3202 gnd.n5325 gnd.n1595 585
R3203 gnd.n5327 gnd.n5326 585
R3204 gnd.n5329 gnd.n1593 585
R3205 gnd.n5331 gnd.n5330 585
R3206 gnd.n5333 gnd.n1590 585
R3207 gnd.n5335 gnd.n5334 585
R3208 gnd.n5337 gnd.n1589 585
R3209 gnd.n5338 gnd.n1528 585
R3210 gnd.n5341 gnd.n1362 585
R3211 gnd.n5343 gnd.n5342 585
R3212 gnd.n5344 gnd.n1584 585
R3213 gnd.n5346 gnd.n5345 585
R3214 gnd.n5348 gnd.n1582 585
R3215 gnd.n5350 gnd.n5349 585
R3216 gnd.n5351 gnd.n1581 585
R3217 gnd.n5353 gnd.n5352 585
R3218 gnd.n5355 gnd.n1579 585
R3219 gnd.n5357 gnd.n5356 585
R3220 gnd.n5358 gnd.n1578 585
R3221 gnd.n5360 gnd.n5359 585
R3222 gnd.n5362 gnd.n1576 585
R3223 gnd.n5364 gnd.n5363 585
R3224 gnd.n5365 gnd.n1575 585
R3225 gnd.n5367 gnd.n5366 585
R3226 gnd.n5369 gnd.n1573 585
R3227 gnd.n5371 gnd.n5370 585
R3228 gnd.n5372 gnd.n1572 585
R3229 gnd.n5374 gnd.n5373 585
R3230 gnd.n5376 gnd.n1570 585
R3231 gnd.n5378 gnd.n5377 585
R3232 gnd.n5379 gnd.n1569 585
R3233 gnd.n5381 gnd.n5380 585
R3234 gnd.n5383 gnd.n1567 585
R3235 gnd.n5385 gnd.n5384 585
R3236 gnd.n5386 gnd.n1566 585
R3237 gnd.n5388 gnd.n5387 585
R3238 gnd.n5390 gnd.n1564 585
R3239 gnd.n5392 gnd.n5391 585
R3240 gnd.n5393 gnd.n1563 585
R3241 gnd.n5395 gnd.n5394 585
R3242 gnd.n5397 gnd.n1562 585
R3243 gnd.n5280 gnd.n1614 585
R3244 gnd.n5280 gnd.n1526 585
R3245 gnd.n5279 gnd.n5278 585
R3246 gnd.n5279 gnd.n1538 585
R3247 gnd.n5277 gnd.n1535 585
R3248 gnd.n5403 gnd.n1535 585
R3249 gnd.n5276 gnd.n5275 585
R3250 gnd.n5275 gnd.n5274 585
R3251 gnd.n1617 gnd.n1616 585
R3252 gnd.n1618 gnd.n1617 585
R3253 gnd.n5244 gnd.n5243 585
R3254 gnd.n5245 gnd.n5244 585
R3255 gnd.n5242 gnd.n1646 585
R3256 gnd.n1646 gnd.n1626 585
R3257 gnd.n5241 gnd.n5240 585
R3258 gnd.n5240 gnd.n1625 585
R3259 gnd.n5239 gnd.n5237 585
R3260 gnd.n5239 gnd.n5238 585
R3261 gnd.n5236 gnd.n1636 585
R3262 gnd.n5253 gnd.n1636 585
R3263 gnd.n5235 gnd.n5234 585
R3264 gnd.n5234 gnd.n1634 585
R3265 gnd.n5233 gnd.n1647 585
R3266 gnd.n5233 gnd.n5232 585
R3267 gnd.n5203 gnd.n1648 585
R3268 gnd.n1656 gnd.n1648 585
R3269 gnd.n5204 gnd.n1654 585
R3270 gnd.n5226 gnd.n1654 585
R3271 gnd.n5206 gnd.n5205 585
R3272 gnd.n5205 gnd.n1653 585
R3273 gnd.n5207 gnd.n1665 585
R3274 gnd.n5217 gnd.n1665 585
R3275 gnd.n5208 gnd.n1672 585
R3276 gnd.n1672 gnd.n1663 585
R3277 gnd.n5210 gnd.n5209 585
R3278 gnd.n5211 gnd.n5210 585
R3279 gnd.n5202 gnd.n1671 585
R3280 gnd.n1675 gnd.n1671 585
R3281 gnd.n5201 gnd.n5200 585
R3282 gnd.n5200 gnd.n5199 585
R3283 gnd.n1674 gnd.n1673 585
R3284 gnd.n1684 gnd.n1674 585
R3285 gnd.n5178 gnd.n1682 585
R3286 gnd.n5193 gnd.n1682 585
R3287 gnd.n5179 gnd.n1696 585
R3288 gnd.n1696 gnd.n1695 585
R3289 gnd.n5181 gnd.n5180 585
R3290 gnd.n5182 gnd.n5181 585
R3291 gnd.n5177 gnd.n1694 585
R3292 gnd.n1694 gnd.n1691 585
R3293 gnd.n5176 gnd.n5175 585
R3294 gnd.n5175 gnd.n5174 585
R3295 gnd.n1698 gnd.n1697 585
R3296 gnd.n5165 gnd.n1698 585
R3297 gnd.n5164 gnd.n5163 585
R3298 gnd.n5166 gnd.n5164 585
R3299 gnd.n5162 gnd.n1707 585
R3300 gnd.n1711 gnd.n1707 585
R3301 gnd.n5161 gnd.n5160 585
R3302 gnd.n5160 gnd.n5159 585
R3303 gnd.n1709 gnd.n1708 585
R3304 gnd.n1710 gnd.n1709 585
R3305 gnd.n5121 gnd.n1716 585
R3306 gnd.n5153 gnd.n1716 585
R3307 gnd.n5123 gnd.n5122 585
R3308 gnd.n5122 gnd.n1727 585
R3309 gnd.n5124 gnd.n1726 585
R3310 gnd.n5135 gnd.n1726 585
R3311 gnd.n5126 gnd.n5125 585
R3312 gnd.n5127 gnd.n5126 585
R3313 gnd.n5120 gnd.n1732 585
R3314 gnd.n5129 gnd.n1732 585
R3315 gnd.n5119 gnd.n5118 585
R3316 gnd.n5118 gnd.n1731 585
R3317 gnd.n5117 gnd.n1734 585
R3318 gnd.n5117 gnd.n5116 585
R3319 gnd.n5093 gnd.n1735 585
R3320 gnd.n5109 gnd.n1735 585
R3321 gnd.n5094 gnd.n1742 585
R3322 gnd.n5110 gnd.n1742 585
R3323 gnd.n5096 gnd.n5095 585
R3324 gnd.n5097 gnd.n5096 585
R3325 gnd.n5092 gnd.n1751 585
R3326 gnd.n1756 gnd.n1751 585
R3327 gnd.n5091 gnd.n5090 585
R3328 gnd.n5090 gnd.n5089 585
R3329 gnd.n1753 gnd.n1752 585
R3330 gnd.n1763 gnd.n1753 585
R3331 gnd.n5058 gnd.n1761 585
R3332 gnd.n5082 gnd.n1761 585
R3333 gnd.n5061 gnd.n5060 585
R3334 gnd.n5060 gnd.n5059 585
R3335 gnd.n5062 gnd.n1771 585
R3336 gnd.n5072 gnd.n1771 585
R3337 gnd.n5063 gnd.n1780 585
R3338 gnd.n1780 gnd.n1769 585
R3339 gnd.n5065 gnd.n5064 585
R3340 gnd.n5066 gnd.n5065 585
R3341 gnd.n5057 gnd.n1779 585
R3342 gnd.n1779 gnd.n1776 585
R3343 gnd.n5056 gnd.n5055 585
R3344 gnd.n5055 gnd.n5054 585
R3345 gnd.n1782 gnd.n1781 585
R3346 gnd.n5047 gnd.n1782 585
R3347 gnd.n5046 gnd.n5045 585
R3348 gnd.n5048 gnd.n5046 585
R3349 gnd.n5044 gnd.n1789 585
R3350 gnd.n1793 gnd.n1789 585
R3351 gnd.n5043 gnd.n5042 585
R3352 gnd.n5042 gnd.n5041 585
R3353 gnd.n1791 gnd.n1790 585
R3354 gnd.n1792 gnd.n1791 585
R3355 gnd.n4999 gnd.n1800 585
R3356 gnd.n5035 gnd.n1800 585
R3357 gnd.n5001 gnd.n5000 585
R3358 gnd.n5000 gnd.n1810 585
R3359 gnd.n5002 gnd.n1809 585
R3360 gnd.n5014 gnd.n1809 585
R3361 gnd.n5004 gnd.n5003 585
R3362 gnd.n5005 gnd.n5004 585
R3363 gnd.n4998 gnd.n1815 585
R3364 gnd.n5008 gnd.n1815 585
R3365 gnd.n4997 gnd.n4996 585
R3366 gnd.n4996 gnd.n1814 585
R3367 gnd.n4995 gnd.n1817 585
R3368 gnd.n4995 gnd.n4994 585
R3369 gnd.n4970 gnd.n1818 585
R3370 gnd.n4987 gnd.n1818 585
R3371 gnd.n4971 gnd.n1824 585
R3372 gnd.n4988 gnd.n1824 585
R3373 gnd.n4973 gnd.n4972 585
R3374 gnd.n4974 gnd.n4973 585
R3375 gnd.n4969 gnd.n1833 585
R3376 gnd.n1837 gnd.n1833 585
R3377 gnd.n4968 gnd.n4967 585
R3378 gnd.n4967 gnd.n4966 585
R3379 gnd.n1835 gnd.n1834 585
R3380 gnd.n1844 gnd.n1835 585
R3381 gnd.n4934 gnd.n1842 585
R3382 gnd.n4959 gnd.n1842 585
R3383 gnd.n4937 gnd.n4936 585
R3384 gnd.n4936 gnd.n4935 585
R3385 gnd.n4938 gnd.n1851 585
R3386 gnd.n4948 gnd.n1851 585
R3387 gnd.n4939 gnd.n1859 585
R3388 gnd.n1859 gnd.n1857 585
R3389 gnd.n4941 gnd.n4940 585
R3390 gnd.n4942 gnd.n4941 585
R3391 gnd.n4933 gnd.n1858 585
R3392 gnd.n1863 gnd.n1858 585
R3393 gnd.n4932 gnd.n4931 585
R3394 gnd.n4931 gnd.n4930 585
R3395 gnd.n1861 gnd.n1860 585
R3396 gnd.n4923 gnd.n1861 585
R3397 gnd.n4922 gnd.n4921 585
R3398 gnd.n4924 gnd.n4922 585
R3399 gnd.n4920 gnd.n1870 585
R3400 gnd.n1874 gnd.n1870 585
R3401 gnd.n4919 gnd.n4918 585
R3402 gnd.n4918 gnd.n4917 585
R3403 gnd.n1872 gnd.n1871 585
R3404 gnd.n1873 gnd.n1872 585
R3405 gnd.n4876 gnd.n1880 585
R3406 gnd.n4911 gnd.n1880 585
R3407 gnd.n4878 gnd.n4877 585
R3408 gnd.n4877 gnd.n1890 585
R3409 gnd.n4879 gnd.n1889 585
R3410 gnd.n4890 gnd.n1889 585
R3411 gnd.n4881 gnd.n4880 585
R3412 gnd.n4882 gnd.n4881 585
R3413 gnd.n4875 gnd.n1894 585
R3414 gnd.n4884 gnd.n1894 585
R3415 gnd.n4874 gnd.n4873 585
R3416 gnd.n4873 gnd.n4872 585
R3417 gnd.n1897 gnd.n1896 585
R3418 gnd.n4862 gnd.n1897 585
R3419 gnd.n4853 gnd.n1906 585
R3420 gnd.n1906 gnd.n1899 585
R3421 gnd.n4855 gnd.n4854 585
R3422 gnd.n4856 gnd.n4855 585
R3423 gnd.n4852 gnd.n1905 585
R3424 gnd.n1905 gnd.n1125 585
R3425 gnd.n4851 gnd.n4850 585
R3426 gnd.n4850 gnd.n4849 585
R3427 gnd.n1980 gnd.n1907 585
R3428 gnd.n4842 gnd.n1980 585
R3429 gnd.n1979 gnd.n1978 585
R3430 gnd.n1979 gnd.n1114 585
R3431 gnd.n1977 gnd.n1112 585
R3432 gnd.n5898 gnd.n1112 585
R3433 gnd.n1976 gnd.n1111 585
R3434 gnd.n5899 gnd.n1111 585
R3435 gnd.n1975 gnd.n1974 585
R3436 gnd.n1974 gnd.n1973 585
R3437 gnd.n6028 gnd.n972 585
R3438 gnd.n4623 gnd.n972 585
R3439 gnd.n6030 gnd.n6029 585
R3440 gnd.n6031 gnd.n6030 585
R3441 gnd.n957 gnd.n956 585
R3442 gnd.n4583 gnd.n957 585
R3443 gnd.n6039 gnd.n6038 585
R3444 gnd.n6038 gnd.n6037 585
R3445 gnd.n6040 gnd.n951 585
R3446 gnd.n4331 gnd.n951 585
R3447 gnd.n6042 gnd.n6041 585
R3448 gnd.n6043 gnd.n6042 585
R3449 gnd.n937 gnd.n936 585
R3450 gnd.n4596 gnd.n937 585
R3451 gnd.n6051 gnd.n6050 585
R3452 gnd.n6050 gnd.n6049 585
R3453 gnd.n6052 gnd.n931 585
R3454 gnd.n4324 gnd.n931 585
R3455 gnd.n6054 gnd.n6053 585
R3456 gnd.n6055 gnd.n6054 585
R3457 gnd.n917 gnd.n916 585
R3458 gnd.n4316 gnd.n917 585
R3459 gnd.n6063 gnd.n6062 585
R3460 gnd.n6062 gnd.n6061 585
R3461 gnd.n6064 gnd.n911 585
R3462 gnd.n4282 gnd.n911 585
R3463 gnd.n6066 gnd.n6065 585
R3464 gnd.n6067 gnd.n6066 585
R3465 gnd.n895 gnd.n894 585
R3466 gnd.n4290 gnd.n895 585
R3467 gnd.n6075 gnd.n6074 585
R3468 gnd.n6074 gnd.n6073 585
R3469 gnd.n6076 gnd.n889 585
R3470 gnd.n4271 gnd.n889 585
R3471 gnd.n6078 gnd.n6077 585
R3472 gnd.n6079 gnd.n6078 585
R3473 gnd.n890 gnd.n888 585
R3474 gnd.n888 gnd.n883 585
R3475 gnd.n4261 gnd.n4260 585
R3476 gnd.n4262 gnd.n4261 585
R3477 gnd.n2079 gnd.n2078 585
R3478 gnd.n2086 gnd.n2078 585
R3479 gnd.n4255 gnd.n4254 585
R3480 gnd.n4254 gnd.n4253 585
R3481 gnd.n2082 gnd.n2081 585
R3482 gnd.n2083 gnd.n2082 585
R3483 gnd.n4233 gnd.n4232 585
R3484 gnd.n4234 gnd.n4233 585
R3485 gnd.n2100 gnd.n2099 585
R3486 gnd.n2099 gnd.n2096 585
R3487 gnd.n4228 gnd.n4227 585
R3488 gnd.n4227 gnd.n4226 585
R3489 gnd.n2103 gnd.n2102 585
R3490 gnd.n4215 gnd.n2103 585
R3491 gnd.n4190 gnd.n2124 585
R3492 gnd.n2124 gnd.n2113 585
R3493 gnd.n4192 gnd.n4191 585
R3494 gnd.n4193 gnd.n4192 585
R3495 gnd.n2125 gnd.n2123 585
R3496 gnd.n2123 gnd.n2120 585
R3497 gnd.n4185 gnd.n4184 585
R3498 gnd.n4184 gnd.n4183 585
R3499 gnd.n2128 gnd.n2127 585
R3500 gnd.n4168 gnd.n2128 585
R3501 gnd.n4155 gnd.n2148 585
R3502 gnd.n2148 gnd.n2139 585
R3503 gnd.n4157 gnd.n4156 585
R3504 gnd.n4158 gnd.n4157 585
R3505 gnd.n2149 gnd.n2147 585
R3506 gnd.n2155 gnd.n2147 585
R3507 gnd.n4150 gnd.n4149 585
R3508 gnd.n4149 gnd.n4148 585
R3509 gnd.n2152 gnd.n2151 585
R3510 gnd.n4133 gnd.n2152 585
R3511 gnd.n4120 gnd.n2173 585
R3512 gnd.n2173 gnd.n2164 585
R3513 gnd.n4122 gnd.n4121 585
R3514 gnd.n4123 gnd.n4122 585
R3515 gnd.n2174 gnd.n2172 585
R3516 gnd.n2181 gnd.n2172 585
R3517 gnd.n4115 gnd.n4114 585
R3518 gnd.n4114 gnd.n4113 585
R3519 gnd.n2177 gnd.n2176 585
R3520 gnd.n2178 gnd.n2177 585
R3521 gnd.n4096 gnd.n4095 585
R3522 gnd.n4097 gnd.n4096 585
R3523 gnd.n2194 gnd.n2193 585
R3524 gnd.n2193 gnd.n2190 585
R3525 gnd.n4091 gnd.n4090 585
R3526 gnd.n4090 gnd.n4089 585
R3527 gnd.n2197 gnd.n2196 585
R3528 gnd.n2198 gnd.n2197 585
R3529 gnd.n4076 gnd.n4075 585
R3530 gnd.n4077 gnd.n4076 585
R3531 gnd.n2211 gnd.n2210 585
R3532 gnd.n2218 gnd.n2210 585
R3533 gnd.n4071 gnd.n4070 585
R3534 gnd.n4070 gnd.n4069 585
R3535 gnd.n2214 gnd.n2213 585
R3536 gnd.n2215 gnd.n2214 585
R3537 gnd.n4056 gnd.n4055 585
R3538 gnd.n4057 gnd.n4056 585
R3539 gnd.n2230 gnd.n2229 585
R3540 gnd.n2229 gnd.n2226 585
R3541 gnd.n4051 gnd.n4050 585
R3542 gnd.n4050 gnd.n4049 585
R3543 gnd.n2233 gnd.n2232 585
R3544 gnd.n2234 gnd.n2233 585
R3545 gnd.n4034 gnd.n4033 585
R3546 gnd.n4032 gnd.n3761 585
R3547 gnd.n4031 gnd.n3760 585
R3548 gnd.n4036 gnd.n3760 585
R3549 gnd.n4030 gnd.n4029 585
R3550 gnd.n4028 gnd.n4027 585
R3551 gnd.n4026 gnd.n4025 585
R3552 gnd.n4024 gnd.n4023 585
R3553 gnd.n4022 gnd.n4021 585
R3554 gnd.n4020 gnd.n4019 585
R3555 gnd.n4018 gnd.n4017 585
R3556 gnd.n4016 gnd.n4015 585
R3557 gnd.n4014 gnd.n4013 585
R3558 gnd.n4012 gnd.n4011 585
R3559 gnd.n4010 gnd.n4009 585
R3560 gnd.n4008 gnd.n4007 585
R3561 gnd.n4006 gnd.n4005 585
R3562 gnd.n4004 gnd.n4003 585
R3563 gnd.n4002 gnd.n4001 585
R3564 gnd.n3999 gnd.n3998 585
R3565 gnd.n3997 gnd.n3996 585
R3566 gnd.n3995 gnd.n3994 585
R3567 gnd.n3993 gnd.n3992 585
R3568 gnd.n3991 gnd.n3990 585
R3569 gnd.n3989 gnd.n3988 585
R3570 gnd.n3987 gnd.n3986 585
R3571 gnd.n3985 gnd.n3984 585
R3572 gnd.n3983 gnd.n3982 585
R3573 gnd.n3981 gnd.n3980 585
R3574 gnd.n3979 gnd.n3978 585
R3575 gnd.n3977 gnd.n3976 585
R3576 gnd.n3975 gnd.n3974 585
R3577 gnd.n3973 gnd.n3972 585
R3578 gnd.n3971 gnd.n3970 585
R3579 gnd.n3969 gnd.n3968 585
R3580 gnd.n3967 gnd.n3966 585
R3581 gnd.n3965 gnd.n3964 585
R3582 gnd.n3963 gnd.n3962 585
R3583 gnd.n3961 gnd.n3960 585
R3584 gnd.n3959 gnd.n3958 585
R3585 gnd.n3957 gnd.n3956 585
R3586 gnd.n3955 gnd.n3954 585
R3587 gnd.n3953 gnd.n3952 585
R3588 gnd.n3951 gnd.n3950 585
R3589 gnd.n3949 gnd.n3948 585
R3590 gnd.n3947 gnd.n3946 585
R3591 gnd.n3945 gnd.n3944 585
R3592 gnd.n3943 gnd.n3942 585
R3593 gnd.n3941 gnd.n3940 585
R3594 gnd.n3939 gnd.n3938 585
R3595 gnd.n3937 gnd.n3936 585
R3596 gnd.n3935 gnd.n3934 585
R3597 gnd.n3933 gnd.n3932 585
R3598 gnd.n3931 gnd.n3930 585
R3599 gnd.n3929 gnd.n3928 585
R3600 gnd.n3927 gnd.n3926 585
R3601 gnd.n3925 gnd.n3924 585
R3602 gnd.n3923 gnd.n3922 585
R3603 gnd.n3921 gnd.n2243 585
R3604 gnd.n4038 gnd.n2242 585
R3605 gnd.n4575 gnd.n4574 585
R3606 gnd.n4573 gnd.n4484 585
R3607 gnd.n4572 gnd.n4571 585
R3608 gnd.n4565 gnd.n4485 585
R3609 gnd.n4567 gnd.n4566 585
R3610 gnd.n4564 gnd.n4563 585
R3611 gnd.n4562 gnd.n4561 585
R3612 gnd.n4555 gnd.n4487 585
R3613 gnd.n4557 gnd.n4556 585
R3614 gnd.n4554 gnd.n4553 585
R3615 gnd.n4552 gnd.n4551 585
R3616 gnd.n4545 gnd.n4489 585
R3617 gnd.n4547 gnd.n4546 585
R3618 gnd.n4544 gnd.n4543 585
R3619 gnd.n4542 gnd.n4541 585
R3620 gnd.n4535 gnd.n4491 585
R3621 gnd.n4537 gnd.n4536 585
R3622 gnd.n4534 gnd.n4533 585
R3623 gnd.n4532 gnd.n4531 585
R3624 gnd.n4525 gnd.n4493 585
R3625 gnd.n4527 gnd.n4526 585
R3626 gnd.n4524 gnd.n4497 585
R3627 gnd.n4523 gnd.n4522 585
R3628 gnd.n4516 gnd.n4498 585
R3629 gnd.n4518 gnd.n4517 585
R3630 gnd.n4515 gnd.n4514 585
R3631 gnd.n4513 gnd.n4512 585
R3632 gnd.n4506 gnd.n4500 585
R3633 gnd.n4508 gnd.n4507 585
R3634 gnd.n4505 gnd.n4504 585
R3635 gnd.n4503 gnd.n1045 585
R3636 gnd.n5975 gnd.n5974 585
R3637 gnd.n5977 gnd.n5976 585
R3638 gnd.n5979 gnd.n5978 585
R3639 gnd.n5981 gnd.n5980 585
R3640 gnd.n5983 gnd.n5982 585
R3641 gnd.n5985 gnd.n5984 585
R3642 gnd.n5987 gnd.n5986 585
R3643 gnd.n5989 gnd.n5988 585
R3644 gnd.n5992 gnd.n5991 585
R3645 gnd.n5994 gnd.n5993 585
R3646 gnd.n5996 gnd.n5995 585
R3647 gnd.n5998 gnd.n5997 585
R3648 gnd.n6000 gnd.n5999 585
R3649 gnd.n6002 gnd.n6001 585
R3650 gnd.n6004 gnd.n6003 585
R3651 gnd.n6006 gnd.n6005 585
R3652 gnd.n6008 gnd.n6007 585
R3653 gnd.n6010 gnd.n6009 585
R3654 gnd.n6012 gnd.n6011 585
R3655 gnd.n6014 gnd.n6013 585
R3656 gnd.n6016 gnd.n6015 585
R3657 gnd.n6018 gnd.n6017 585
R3658 gnd.n6019 gnd.n1018 585
R3659 gnd.n6021 gnd.n6020 585
R3660 gnd.n977 gnd.n976 585
R3661 gnd.n6025 gnd.n6024 585
R3662 gnd.n6024 gnd.n6023 585
R3663 gnd.n4579 gnd.n2038 585
R3664 gnd.n4623 gnd.n2038 585
R3665 gnd.n4580 gnd.n969 585
R3666 gnd.n6031 gnd.n969 585
R3667 gnd.n4582 gnd.n4581 585
R3668 gnd.n4583 gnd.n4582 585
R3669 gnd.n4334 gnd.n959 585
R3670 gnd.n6037 gnd.n959 585
R3671 gnd.n4333 gnd.n4332 585
R3672 gnd.n4332 gnd.n4331 585
R3673 gnd.n4329 gnd.n948 585
R3674 gnd.n6043 gnd.n948 585
R3675 gnd.n4328 gnd.n2049 585
R3676 gnd.n4596 gnd.n2049 585
R3677 gnd.n4327 gnd.n939 585
R3678 gnd.n6049 gnd.n939 585
R3679 gnd.n4326 gnd.n4325 585
R3680 gnd.n4325 gnd.n4324 585
R3681 gnd.n2055 gnd.n928 585
R3682 gnd.n6055 gnd.n928 585
R3683 gnd.n4278 gnd.n2060 585
R3684 gnd.n4316 gnd.n2060 585
R3685 gnd.n4279 gnd.n919 585
R3686 gnd.n6061 gnd.n919 585
R3687 gnd.n4281 gnd.n4280 585
R3688 gnd.n4282 gnd.n4281 585
R3689 gnd.n4276 gnd.n908 585
R3690 gnd.n6067 gnd.n908 585
R3691 gnd.n4275 gnd.n2066 585
R3692 gnd.n4290 gnd.n2066 585
R3693 gnd.n4274 gnd.n897 585
R3694 gnd.n6073 gnd.n897 585
R3695 gnd.n4273 gnd.n4272 585
R3696 gnd.n4272 gnd.n4271 585
R3697 gnd.n2070 gnd.n884 585
R3698 gnd.n6079 gnd.n884 585
R3699 gnd.n4243 gnd.n4242 585
R3700 gnd.n4242 gnd.n883 585
R3701 gnd.n4241 gnd.n2076 585
R3702 gnd.n4262 gnd.n2076 585
R3703 gnd.n4240 gnd.n4239 585
R3704 gnd.n4239 gnd.n2086 585
R3705 gnd.n4238 gnd.n2084 585
R3706 gnd.n4253 gnd.n2084 585
R3707 gnd.n4237 gnd.n4236 585
R3708 gnd.n4236 gnd.n2083 585
R3709 gnd.n4235 gnd.n2093 585
R3710 gnd.n4235 gnd.n4234 585
R3711 gnd.n4219 gnd.n2095 585
R3712 gnd.n2096 gnd.n2095 585
R3713 gnd.n4218 gnd.n2104 585
R3714 gnd.n4226 gnd.n2104 585
R3715 gnd.n4217 gnd.n4216 585
R3716 gnd.n4216 gnd.n4215 585
R3717 gnd.n2112 gnd.n2110 585
R3718 gnd.n2113 gnd.n2112 585
R3719 gnd.n4174 gnd.n2121 585
R3720 gnd.n4193 gnd.n2121 585
R3721 gnd.n4173 gnd.n4172 585
R3722 gnd.n4172 gnd.n2120 585
R3723 gnd.n4171 gnd.n2129 585
R3724 gnd.n4183 gnd.n2129 585
R3725 gnd.n4170 gnd.n4169 585
R3726 gnd.n4169 gnd.n4168 585
R3727 gnd.n2138 gnd.n2136 585
R3728 gnd.n2139 gnd.n2138 585
R3729 gnd.n4139 gnd.n2145 585
R3730 gnd.n4158 gnd.n2145 585
R3731 gnd.n4138 gnd.n4137 585
R3732 gnd.n4137 gnd.n2155 585
R3733 gnd.n4136 gnd.n2153 585
R3734 gnd.n4148 gnd.n2153 585
R3735 gnd.n4135 gnd.n4134 585
R3736 gnd.n4134 gnd.n4133 585
R3737 gnd.n2163 gnd.n2161 585
R3738 gnd.n2164 gnd.n2163 585
R3739 gnd.n4104 gnd.n2170 585
R3740 gnd.n4123 gnd.n2170 585
R3741 gnd.n4103 gnd.n4102 585
R3742 gnd.n4102 gnd.n2181 585
R3743 gnd.n4101 gnd.n2179 585
R3744 gnd.n4113 gnd.n2179 585
R3745 gnd.n4100 gnd.n4099 585
R3746 gnd.n4099 gnd.n2178 585
R3747 gnd.n4098 gnd.n2187 585
R3748 gnd.n4098 gnd.n4097 585
R3749 gnd.n4082 gnd.n2189 585
R3750 gnd.n2190 gnd.n2189 585
R3751 gnd.n4081 gnd.n2199 585
R3752 gnd.n4089 gnd.n2199 585
R3753 gnd.n4080 gnd.n4079 585
R3754 gnd.n4079 gnd.n2198 585
R3755 gnd.n4078 gnd.n2205 585
R3756 gnd.n4078 gnd.n4077 585
R3757 gnd.n4062 gnd.n2207 585
R3758 gnd.n2218 gnd.n2207 585
R3759 gnd.n4061 gnd.n2216 585
R3760 gnd.n4069 gnd.n2216 585
R3761 gnd.n4060 gnd.n4059 585
R3762 gnd.n4059 gnd.n2215 585
R3763 gnd.n4058 gnd.n2223 585
R3764 gnd.n4058 gnd.n4057 585
R3765 gnd.n4042 gnd.n2225 585
R3766 gnd.n2226 gnd.n2225 585
R3767 gnd.n4041 gnd.n2235 585
R3768 gnd.n4049 gnd.n2235 585
R3769 gnd.n4040 gnd.n4039 585
R3770 gnd.n4039 gnd.n2234 585
R3771 gnd.n7188 gnd.n205 585
R3772 gnd.n205 gnd.n204 585
R3773 gnd.n7190 gnd.n7189 585
R3774 gnd.n7191 gnd.n7190 585
R3775 gnd.n192 gnd.n191 585
R3776 gnd.n195 gnd.n192 585
R3777 gnd.n7199 gnd.n7198 585
R3778 gnd.n7198 gnd.n7197 585
R3779 gnd.n7200 gnd.n186 585
R3780 gnd.n186 gnd.n185 585
R3781 gnd.n7202 gnd.n7201 585
R3782 gnd.n7203 gnd.n7202 585
R3783 gnd.n173 gnd.n172 585
R3784 gnd.n182 gnd.n173 585
R3785 gnd.n7211 gnd.n7210 585
R3786 gnd.n7210 gnd.n7209 585
R3787 gnd.n7212 gnd.n167 585
R3788 gnd.n167 gnd.n166 585
R3789 gnd.n7214 gnd.n7213 585
R3790 gnd.n7215 gnd.n7214 585
R3791 gnd.n154 gnd.n153 585
R3792 gnd.n7041 gnd.n154 585
R3793 gnd.n7223 gnd.n7222 585
R3794 gnd.n7222 gnd.n7221 585
R3795 gnd.n7224 gnd.n148 585
R3796 gnd.n148 gnd.n147 585
R3797 gnd.n7226 gnd.n7225 585
R3798 gnd.n7227 gnd.n7226 585
R3799 gnd.n135 gnd.n134 585
R3800 gnd.n144 gnd.n135 585
R3801 gnd.n7235 gnd.n7234 585
R3802 gnd.n7234 gnd.n7233 585
R3803 gnd.n7236 gnd.n129 585
R3804 gnd.n129 gnd.n128 585
R3805 gnd.n7238 gnd.n7237 585
R3806 gnd.n7239 gnd.n7238 585
R3807 gnd.n116 gnd.n115 585
R3808 gnd.n119 gnd.n116 585
R3809 gnd.n7247 gnd.n7246 585
R3810 gnd.n7246 gnd.n7245 585
R3811 gnd.n7248 gnd.n110 585
R3812 gnd.n110 gnd.n109 585
R3813 gnd.n7250 gnd.n7249 585
R3814 gnd.n7251 gnd.n7250 585
R3815 gnd.n95 gnd.n94 585
R3816 gnd.n106 gnd.n95 585
R3817 gnd.n7259 gnd.n7258 585
R3818 gnd.n7258 gnd.n7257 585
R3819 gnd.n7260 gnd.n89 585
R3820 gnd.n89 gnd.n86 585
R3821 gnd.n7262 gnd.n7261 585
R3822 gnd.n7263 gnd.n7262 585
R3823 gnd.n90 gnd.n88 585
R3824 gnd.n6893 gnd.n88 585
R3825 gnd.n6882 gnd.n324 585
R3826 gnd.n324 gnd.n313 585
R3827 gnd.n6884 gnd.n6883 585
R3828 gnd.n6885 gnd.n6884 585
R3829 gnd.n325 gnd.n323 585
R3830 gnd.n323 gnd.n319 585
R3831 gnd.n6876 gnd.n6875 585
R3832 gnd.n6875 gnd.n6874 585
R3833 gnd.n328 gnd.n327 585
R3834 gnd.n6865 gnd.n328 585
R3835 gnd.n6848 gnd.n346 585
R3836 gnd.n346 gnd.n336 585
R3837 gnd.n6850 gnd.n6849 585
R3838 gnd.n6851 gnd.n6850 585
R3839 gnd.n347 gnd.n345 585
R3840 gnd.n354 gnd.n345 585
R3841 gnd.n6843 gnd.n6842 585
R3842 gnd.n6842 gnd.n6841 585
R3843 gnd.n350 gnd.n349 585
R3844 gnd.n6826 gnd.n350 585
R3845 gnd.n6814 gnd.n374 585
R3846 gnd.n6800 gnd.n374 585
R3847 gnd.n6816 gnd.n6815 585
R3848 gnd.n6817 gnd.n6816 585
R3849 gnd.n375 gnd.n373 585
R3850 gnd.n6794 gnd.n373 585
R3851 gnd.n6809 gnd.n6808 585
R3852 gnd.n6808 gnd.n6807 585
R3853 gnd.n378 gnd.n377 585
R3854 gnd.n5502 gnd.n378 585
R3855 gnd.n5559 gnd.n5555 585
R3856 gnd.n5555 gnd.n5554 585
R3857 gnd.n5561 gnd.n5560 585
R3858 gnd.n5562 gnd.n5561 585
R3859 gnd.n1442 gnd.n1441 585
R3860 gnd.n5493 gnd.n1442 585
R3861 gnd.n5570 gnd.n5569 585
R3862 gnd.n5569 gnd.n5568 585
R3863 gnd.n5571 gnd.n1436 585
R3864 gnd.n5489 gnd.n1436 585
R3865 gnd.n5573 gnd.n5572 585
R3866 gnd.n5574 gnd.n5573 585
R3867 gnd.n1421 gnd.n1420 585
R3868 gnd.n5484 gnd.n1421 585
R3869 gnd.n5582 gnd.n5581 585
R3870 gnd.n5581 gnd.n5580 585
R3871 gnd.n5583 gnd.n1412 585
R3872 gnd.n5480 gnd.n1412 585
R3873 gnd.n5585 gnd.n5584 585
R3874 gnd.n5586 gnd.n5585 585
R3875 gnd.n1413 gnd.n1411 585
R3876 gnd.n5525 gnd.n1411 585
R3877 gnd.n1414 gnd.n1333 585
R3878 gnd.n5592 gnd.n1333 585
R3879 gnd.n5711 gnd.n5710 585
R3880 gnd.n5709 gnd.n1332 585
R3881 gnd.n5708 gnd.n1331 585
R3882 gnd.n5713 gnd.n1331 585
R3883 gnd.n5707 gnd.n5706 585
R3884 gnd.n5705 gnd.n5704 585
R3885 gnd.n5703 gnd.n5702 585
R3886 gnd.n5701 gnd.n5700 585
R3887 gnd.n5699 gnd.n5698 585
R3888 gnd.n5697 gnd.n5696 585
R3889 gnd.n5695 gnd.n5694 585
R3890 gnd.n5693 gnd.n5692 585
R3891 gnd.n5691 gnd.n5690 585
R3892 gnd.n5689 gnd.n5688 585
R3893 gnd.n5687 gnd.n5686 585
R3894 gnd.n5685 gnd.n5684 585
R3895 gnd.n5683 gnd.n5682 585
R3896 gnd.n5681 gnd.n5680 585
R3897 gnd.n5679 gnd.n5678 585
R3898 gnd.n5676 gnd.n5675 585
R3899 gnd.n5674 gnd.n5673 585
R3900 gnd.n5672 gnd.n5671 585
R3901 gnd.n5670 gnd.n5669 585
R3902 gnd.n5668 gnd.n5667 585
R3903 gnd.n5666 gnd.n5665 585
R3904 gnd.n5664 gnd.n5663 585
R3905 gnd.n5662 gnd.n5661 585
R3906 gnd.n5659 gnd.n5658 585
R3907 gnd.n5657 gnd.n5656 585
R3908 gnd.n5655 gnd.n5654 585
R3909 gnd.n5653 gnd.n5652 585
R3910 gnd.n5651 gnd.n5650 585
R3911 gnd.n5649 gnd.n5648 585
R3912 gnd.n5647 gnd.n5646 585
R3913 gnd.n5645 gnd.n5644 585
R3914 gnd.n5643 gnd.n5642 585
R3915 gnd.n5641 gnd.n5640 585
R3916 gnd.n5639 gnd.n5638 585
R3917 gnd.n5637 gnd.n5636 585
R3918 gnd.n5635 gnd.n5634 585
R3919 gnd.n5633 gnd.n5632 585
R3920 gnd.n5631 gnd.n5630 585
R3921 gnd.n5629 gnd.n5628 585
R3922 gnd.n5627 gnd.n5626 585
R3923 gnd.n5625 gnd.n5624 585
R3924 gnd.n5623 gnd.n5622 585
R3925 gnd.n5621 gnd.n5620 585
R3926 gnd.n5619 gnd.n5618 585
R3927 gnd.n5617 gnd.n5616 585
R3928 gnd.n5615 gnd.n5614 585
R3929 gnd.n5613 gnd.n5612 585
R3930 gnd.n5611 gnd.n5610 585
R3931 gnd.n5609 gnd.n5608 585
R3932 gnd.n5607 gnd.n5606 585
R3933 gnd.n5605 gnd.n5604 585
R3934 gnd.n5603 gnd.n5602 585
R3935 gnd.n5601 gnd.n5600 585
R3936 gnd.n5595 gnd.n5594 585
R3937 gnd.n7059 gnd.n305 585
R3938 gnd.n7067 gnd.n7066 585
R3939 gnd.n7069 gnd.n7068 585
R3940 gnd.n7071 gnd.n7070 585
R3941 gnd.n7073 gnd.n7072 585
R3942 gnd.n7075 gnd.n7074 585
R3943 gnd.n7077 gnd.n7076 585
R3944 gnd.n7079 gnd.n7078 585
R3945 gnd.n7081 gnd.n7080 585
R3946 gnd.n7083 gnd.n7082 585
R3947 gnd.n7085 gnd.n7084 585
R3948 gnd.n7087 gnd.n7086 585
R3949 gnd.n7089 gnd.n7088 585
R3950 gnd.n7091 gnd.n7090 585
R3951 gnd.n7093 gnd.n7092 585
R3952 gnd.n7095 gnd.n7094 585
R3953 gnd.n7097 gnd.n7096 585
R3954 gnd.n7099 gnd.n7098 585
R3955 gnd.n7101 gnd.n7100 585
R3956 gnd.n7104 gnd.n7103 585
R3957 gnd.n7102 gnd.n285 585
R3958 gnd.n7109 gnd.n7108 585
R3959 gnd.n7111 gnd.n7110 585
R3960 gnd.n7113 gnd.n7112 585
R3961 gnd.n7115 gnd.n7114 585
R3962 gnd.n7117 gnd.n7116 585
R3963 gnd.n7119 gnd.n7118 585
R3964 gnd.n7121 gnd.n7120 585
R3965 gnd.n7123 gnd.n7122 585
R3966 gnd.n7125 gnd.n7124 585
R3967 gnd.n7127 gnd.n7126 585
R3968 gnd.n7129 gnd.n7128 585
R3969 gnd.n7131 gnd.n7130 585
R3970 gnd.n7133 gnd.n7132 585
R3971 gnd.n7135 gnd.n7134 585
R3972 gnd.n7137 gnd.n7136 585
R3973 gnd.n7139 gnd.n7138 585
R3974 gnd.n7141 gnd.n7140 585
R3975 gnd.n7143 gnd.n7142 585
R3976 gnd.n7145 gnd.n7144 585
R3977 gnd.n7147 gnd.n7146 585
R3978 gnd.n7152 gnd.n7151 585
R3979 gnd.n7154 gnd.n7153 585
R3980 gnd.n7156 gnd.n7155 585
R3981 gnd.n7158 gnd.n7157 585
R3982 gnd.n7160 gnd.n7159 585
R3983 gnd.n7162 gnd.n7161 585
R3984 gnd.n7164 gnd.n7163 585
R3985 gnd.n7166 gnd.n7165 585
R3986 gnd.n7168 gnd.n7167 585
R3987 gnd.n7170 gnd.n7169 585
R3988 gnd.n7172 gnd.n7171 585
R3989 gnd.n7174 gnd.n7173 585
R3990 gnd.n7176 gnd.n7175 585
R3991 gnd.n7178 gnd.n7177 585
R3992 gnd.n7179 gnd.n249 585
R3993 gnd.n7181 gnd.n7180 585
R3994 gnd.n210 gnd.n209 585
R3995 gnd.n7185 gnd.n7184 585
R3996 gnd.n7184 gnd.n7183 585
R3997 gnd.n7061 gnd.n7060 585
R3998 gnd.n7060 gnd.n204 585
R3999 gnd.n7058 gnd.n202 585
R4000 gnd.n7191 gnd.n202 585
R4001 gnd.n7057 gnd.n7056 585
R4002 gnd.n7056 gnd.n195 585
R4003 gnd.n7055 gnd.n193 585
R4004 gnd.n7197 gnd.n193 585
R4005 gnd.n7054 gnd.n7053 585
R4006 gnd.n7053 gnd.n185 585
R4007 gnd.n7051 gnd.n183 585
R4008 gnd.n7203 gnd.n183 585
R4009 gnd.n7050 gnd.n7049 585
R4010 gnd.n7049 gnd.n182 585
R4011 gnd.n7048 gnd.n174 585
R4012 gnd.n7209 gnd.n174 585
R4013 gnd.n7047 gnd.n7046 585
R4014 gnd.n7046 gnd.n166 585
R4015 gnd.n7044 gnd.n164 585
R4016 gnd.n7215 gnd.n164 585
R4017 gnd.n7043 gnd.n7042 585
R4018 gnd.n7042 gnd.n7041 585
R4019 gnd.n6922 gnd.n155 585
R4020 gnd.n7221 gnd.n155 585
R4021 gnd.n6921 gnd.n6920 585
R4022 gnd.n6920 gnd.n147 585
R4023 gnd.n6918 gnd.n145 585
R4024 gnd.n7227 gnd.n145 585
R4025 gnd.n6917 gnd.n6916 585
R4026 gnd.n6916 gnd.n144 585
R4027 gnd.n6915 gnd.n136 585
R4028 gnd.n7233 gnd.n136 585
R4029 gnd.n6914 gnd.n6913 585
R4030 gnd.n6913 gnd.n128 585
R4031 gnd.n6911 gnd.n126 585
R4032 gnd.n7239 gnd.n126 585
R4033 gnd.n6910 gnd.n6909 585
R4034 gnd.n6909 gnd.n119 585
R4035 gnd.n6908 gnd.n117 585
R4036 gnd.n7245 gnd.n117 585
R4037 gnd.n6907 gnd.n6906 585
R4038 gnd.n6906 gnd.n109 585
R4039 gnd.n6904 gnd.n107 585
R4040 gnd.n7251 gnd.n107 585
R4041 gnd.n6903 gnd.n6902 585
R4042 gnd.n6902 gnd.n106 585
R4043 gnd.n6901 gnd.n96 585
R4044 gnd.n7257 gnd.n96 585
R4045 gnd.n6900 gnd.n6899 585
R4046 gnd.n6899 gnd.n86 585
R4047 gnd.n309 gnd.n85 585
R4048 gnd.n7263 gnd.n85 585
R4049 gnd.n6892 gnd.n6891 585
R4050 gnd.n6893 gnd.n6892 585
R4051 gnd.n6890 gnd.n314 585
R4052 gnd.n314 gnd.n313 585
R4053 gnd.n320 gnd.n315 585
R4054 gnd.n6885 gnd.n320 585
R4055 gnd.n6869 gnd.n6868 585
R4056 gnd.n6868 gnd.n319 585
R4057 gnd.n6870 gnd.n329 585
R4058 gnd.n6874 gnd.n329 585
R4059 gnd.n6867 gnd.n6866 585
R4060 gnd.n6866 gnd.n6865 585
R4061 gnd.n335 gnd.n334 585
R4062 gnd.n336 gnd.n335 585
R4063 gnd.n6832 gnd.n343 585
R4064 gnd.n6851 gnd.n343 585
R4065 gnd.n6831 gnd.n6830 585
R4066 gnd.n6830 gnd.n354 585
R4067 gnd.n6829 gnd.n352 585
R4068 gnd.n6841 gnd.n352 585
R4069 gnd.n6828 gnd.n6827 585
R4070 gnd.n6827 gnd.n6826 585
R4071 gnd.n362 gnd.n360 585
R4072 gnd.n6800 gnd.n362 585
R4073 gnd.n6797 gnd.n370 585
R4074 gnd.n6817 gnd.n370 585
R4075 gnd.n6796 gnd.n6795 585
R4076 gnd.n6795 gnd.n6794 585
R4077 gnd.n388 gnd.n380 585
R4078 gnd.n6807 gnd.n380 585
R4079 gnd.n5501 gnd.n5500 585
R4080 gnd.n5502 gnd.n5501 585
R4081 gnd.n5497 gnd.n1457 585
R4082 gnd.n5554 gnd.n1457 585
R4083 gnd.n5496 gnd.n1454 585
R4084 gnd.n5562 gnd.n1454 585
R4085 gnd.n5495 gnd.n5494 585
R4086 gnd.n5494 gnd.n5493 585
R4087 gnd.n5492 gnd.n1444 585
R4088 gnd.n5568 gnd.n1444 585
R4089 gnd.n5491 gnd.n5490 585
R4090 gnd.n5490 gnd.n5489 585
R4091 gnd.n5487 gnd.n1433 585
R4092 gnd.n5574 gnd.n1433 585
R4093 gnd.n5486 gnd.n5485 585
R4094 gnd.n5485 gnd.n5484 585
R4095 gnd.n5483 gnd.n1423 585
R4096 gnd.n5580 gnd.n1423 585
R4097 gnd.n5482 gnd.n5481 585
R4098 gnd.n5481 gnd.n5480 585
R4099 gnd.n5478 gnd.n1408 585
R4100 gnd.n5586 gnd.n1408 585
R4101 gnd.n5477 gnd.n1396 585
R4102 gnd.n5525 gnd.n1396 585
R4103 gnd.n5593 gnd.n1397 585
R4104 gnd.n5593 gnd.n5592 585
R4105 gnd.n6082 gnd.n6081 585
R4106 gnd.n6081 gnd.n6080 585
R4107 gnd.n6787 gnd.n6786 585
R4108 gnd.n6787 gnd.n351 585
R4109 gnd.n6789 gnd.n6788 585
R4110 gnd.n6788 gnd.n363 585
R4111 gnd.n6790 gnd.n390 585
R4112 gnd.n390 gnd.n371 585
R4113 gnd.n6792 gnd.n6791 585
R4114 gnd.n6793 gnd.n6792 585
R4115 gnd.n391 gnd.n389 585
R4116 gnd.n389 gnd.n382 585
R4117 gnd.n5550 gnd.n1460 585
R4118 gnd.n1460 gnd.n379 585
R4119 gnd.n5552 gnd.n5551 585
R4120 gnd.n5553 gnd.n5552 585
R4121 gnd.n1461 gnd.n1459 585
R4122 gnd.n1459 gnd.n1456 585
R4123 gnd.n5544 gnd.n5543 585
R4124 gnd.n5543 gnd.n1453 585
R4125 gnd.n5542 gnd.n1463 585
R4126 gnd.n5542 gnd.n1446 585
R4127 gnd.n5541 gnd.n5540 585
R4128 gnd.n5541 gnd.n1443 585
R4129 gnd.n1465 gnd.n1464 585
R4130 gnd.n1464 gnd.n1435 585
R4131 gnd.n5536 gnd.n5535 585
R4132 gnd.n5535 gnd.n1432 585
R4133 gnd.n5534 gnd.n1467 585
R4134 gnd.n5534 gnd.n1425 585
R4135 gnd.n5533 gnd.n5532 585
R4136 gnd.n5533 gnd.n1422 585
R4137 gnd.n1469 gnd.n1468 585
R4138 gnd.n1468 gnd.n1410 585
R4139 gnd.n5528 gnd.n5527 585
R4140 gnd.n5527 gnd.n5526 585
R4141 gnd.n1472 gnd.n1471 585
R4142 gnd.n1472 gnd.n1400 585
R4143 gnd.n5453 gnd.n5452 585
R4144 gnd.n5453 gnd.n1398 585
R4145 gnd.n5454 gnd.n5449 585
R4146 gnd.n5454 gnd.n1330 585
R4147 gnd.n5456 gnd.n5455 585
R4148 gnd.n5455 gnd.n1288 585
R4149 gnd.n5457 gnd.n1503 585
R4150 gnd.n1503 gnd.n1501 585
R4151 gnd.n5459 gnd.n5458 585
R4152 gnd.n5460 gnd.n5459 585
R4153 gnd.n1504 gnd.n1502 585
R4154 gnd.n1502 gnd.n1221 585
R4155 gnd.n5443 gnd.n1220 585
R4156 gnd.n5781 gnd.n1220 585
R4157 gnd.n5442 gnd.n5441 585
R4158 gnd.n5441 gnd.n1219 585
R4159 gnd.n5440 gnd.n1506 585
R4160 gnd.n5440 gnd.n5439 585
R4161 gnd.n5428 gnd.n1507 585
R4162 gnd.n1508 gnd.n1507 585
R4163 gnd.n5430 gnd.n5429 585
R4164 gnd.n5431 gnd.n5430 585
R4165 gnd.n1517 gnd.n1516 585
R4166 gnd.n1516 gnd.n1515 585
R4167 gnd.n5422 gnd.n5421 585
R4168 gnd.n5421 gnd.n5420 585
R4169 gnd.n1520 gnd.n1519 585
R4170 gnd.n1527 gnd.n1520 585
R4171 gnd.n5411 gnd.n5410 585
R4172 gnd.n5412 gnd.n5411 585
R4173 gnd.n1530 gnd.n1529 585
R4174 gnd.n1537 gnd.n1529 585
R4175 gnd.n5406 gnd.n5405 585
R4176 gnd.n5405 gnd.n5404 585
R4177 gnd.n1533 gnd.n1532 585
R4178 gnd.n5273 gnd.n1533 585
R4179 gnd.n5261 gnd.n1629 585
R4180 gnd.n1645 gnd.n1629 585
R4181 gnd.n5263 gnd.n5262 585
R4182 gnd.n5264 gnd.n5263 585
R4183 gnd.n1630 gnd.n1628 585
R4184 gnd.n1637 gnd.n1628 585
R4185 gnd.n5256 gnd.n5255 585
R4186 gnd.n5255 gnd.n5254 585
R4187 gnd.n1633 gnd.n1632 585
R4188 gnd.n1649 gnd.n1633 585
R4189 gnd.n5224 gnd.n5223 585
R4190 gnd.n5225 gnd.n5224 585
R4191 gnd.n1659 gnd.n1658 585
R4192 gnd.n1666 gnd.n1658 585
R4193 gnd.n5219 gnd.n5218 585
R4194 gnd.n5218 gnd.t189 585
R4195 gnd.n1662 gnd.n1661 585
R4196 gnd.n1670 gnd.n1662 585
R4197 gnd.n5189 gnd.n1686 585
R4198 gnd.n1686 gnd.n1677 585
R4199 gnd.n5191 gnd.n5190 585
R4200 gnd.n5192 gnd.n5191 585
R4201 gnd.n1687 gnd.n1685 585
R4202 gnd.n1685 gnd.n1681 585
R4203 gnd.n5184 gnd.n5183 585
R4204 gnd.n5183 gnd.n5182 585
R4205 gnd.n1690 gnd.n1689 585
R4206 gnd.n1701 gnd.n1690 585
R4207 gnd.n5146 gnd.n5145 585
R4208 gnd.n5146 gnd.n1699 585
R4209 gnd.n5148 gnd.n5147 585
R4210 gnd.n5147 gnd.n1706 585
R4211 gnd.n5149 gnd.n1720 585
R4212 gnd.n1720 gnd.n1712 585
R4213 gnd.n5151 gnd.n5150 585
R4214 gnd.n5152 gnd.n5151 585
R4215 gnd.n1721 gnd.n1719 585
R4216 gnd.n4735 gnd.n1719 585
R4217 gnd.n5138 gnd.n5137 585
R4218 gnd.n5137 gnd.n5136 585
R4219 gnd.n1724 gnd.n1723 585
R4220 gnd.n5128 gnd.n1724 585
R4221 gnd.n5105 gnd.n1745 585
R4222 gnd.n1745 gnd.n1737 585
R4223 gnd.n5107 gnd.n5106 585
R4224 gnd.n5108 gnd.n5107 585
R4225 gnd.n1746 gnd.n1744 585
R4226 gnd.n1744 gnd.n1741 585
R4227 gnd.n5100 gnd.n5099 585
R4228 gnd.n5099 gnd.n5098 585
R4229 gnd.n1749 gnd.n1748 585
R4230 gnd.n1755 gnd.n1749 585
R4231 gnd.n5080 gnd.n5079 585
R4232 gnd.n5081 gnd.n5080 585
R4233 gnd.n1765 gnd.n1764 585
R4234 gnd.n1772 gnd.n1764 585
R4235 gnd.n5075 gnd.n5074 585
R4236 gnd.n5074 gnd.n5073 585
R4237 gnd.n1768 gnd.n1767 585
R4238 gnd.n5066 gnd.n1768 585
R4239 gnd.n5027 gnd.n5026 585
R4240 gnd.n5027 gnd.n1784 585
R4241 gnd.n5028 gnd.n5023 585
R4242 gnd.n5028 gnd.n1783 585
R4243 gnd.n5030 gnd.n5029 585
R4244 gnd.n5029 gnd.n1788 585
R4245 gnd.n5031 gnd.n1803 585
R4246 gnd.n1803 gnd.n1795 585
R4247 gnd.n5033 gnd.n5032 585
R4248 gnd.n5034 gnd.n5033 585
R4249 gnd.n1804 gnd.n1802 585
R4250 gnd.n1802 gnd.n1799 585
R4251 gnd.n5017 gnd.n5016 585
R4252 gnd.n5016 gnd.n5015 585
R4253 gnd.n1807 gnd.n1806 585
R4254 gnd.n5007 gnd.n1807 585
R4255 gnd.n4983 gnd.n1827 585
R4256 gnd.n1827 gnd.n1819 585
R4257 gnd.n4985 gnd.n4984 585
R4258 gnd.n4986 gnd.n4985 585
R4259 gnd.n1828 gnd.n1826 585
R4260 gnd.n1826 gnd.n1823 585
R4261 gnd.n4978 gnd.n4977 585
R4262 gnd.n4977 gnd.n4976 585
R4263 gnd.n1831 gnd.n1830 585
R4264 gnd.n1836 gnd.n1831 585
R4265 gnd.n4957 gnd.n4956 585
R4266 gnd.n4958 gnd.n4957 585
R4267 gnd.n1846 gnd.n1845 585
R4268 gnd.n1852 gnd.n1845 585
R4269 gnd.n4952 gnd.n4951 585
R4270 gnd.n4951 gnd.n4950 585
R4271 gnd.n1849 gnd.n1848 585
R4272 gnd.n4942 gnd.n1849 585
R4273 gnd.n4904 gnd.n4903 585
R4274 gnd.n4904 gnd.n1864 585
R4275 gnd.n4905 gnd.n4900 585
R4276 gnd.n4905 gnd.n1862 585
R4277 gnd.n4907 gnd.n4906 585
R4278 gnd.n4906 gnd.n1869 585
R4279 gnd.n4908 gnd.n1883 585
R4280 gnd.n1883 gnd.n1875 585
R4281 gnd.n4910 gnd.n4909 585
R4282 gnd.t5 gnd.n4910 585
R4283 gnd.n1884 gnd.n1882 585
R4284 gnd.n1882 gnd.n1879 585
R4285 gnd.n4894 gnd.n4893 585
R4286 gnd.n4893 gnd.n4892 585
R4287 gnd.n1887 gnd.n1886 585
R4288 gnd.n4883 gnd.n1887 585
R4289 gnd.n4870 gnd.n4869 585
R4290 gnd.n4871 gnd.n4870 585
R4291 gnd.n4865 gnd.n4864 585
R4292 gnd.n4864 gnd.n4863 585
R4293 gnd.n1123 gnd.n1122 585
R4294 gnd.n1904 gnd.n1123 585
R4295 gnd.n5893 gnd.n5892 585
R4296 gnd.n5892 gnd.n5891 585
R4297 gnd.n5894 gnd.n1117 585
R4298 gnd.n4841 gnd.n1117 585
R4299 gnd.n5896 gnd.n5895 585
R4300 gnd.n5897 gnd.n5896 585
R4301 gnd.n1118 gnd.n1116 585
R4302 gnd.n1116 gnd.n1110 585
R4303 gnd.n4678 gnd.n4677 585
R4304 gnd.n4678 gnd.n1084 585
R4305 gnd.n4680 gnd.n4679 585
R4306 gnd.n4679 gnd.n1052 585
R4307 gnd.n4681 gnd.n1994 585
R4308 gnd.n1994 gnd.n1991 585
R4309 gnd.n4683 gnd.n4682 585
R4310 gnd.n4684 gnd.n4683 585
R4311 gnd.n1995 gnd.n1993 585
R4312 gnd.n1993 gnd.n1990 585
R4313 gnd.n4669 gnd.n4668 585
R4314 gnd.n4668 gnd.n4667 585
R4315 gnd.n1998 gnd.n1997 585
R4316 gnd.n1999 gnd.n1998 585
R4317 gnd.n4641 gnd.n4640 585
R4318 gnd.n4642 gnd.n4641 585
R4319 gnd.n2011 gnd.n2010 585
R4320 gnd.n2010 gnd.n2008 585
R4321 gnd.n4636 gnd.n4635 585
R4322 gnd.n4635 gnd.n4634 585
R4323 gnd.n2014 gnd.n2013 585
R4324 gnd.n4633 gnd.n2014 585
R4325 gnd.n4616 gnd.n4615 585
R4326 gnd.n4616 gnd.n2015 585
R4327 gnd.n4618 gnd.n4617 585
R4328 gnd.n4617 gnd.n989 585
R4329 gnd.n4619 gnd.n2040 585
R4330 gnd.n2040 gnd.n978 585
R4331 gnd.n4621 gnd.n4620 585
R4332 gnd.n4622 gnd.n4621 585
R4333 gnd.n2041 gnd.n2039 585
R4334 gnd.n2039 gnd.n971 585
R4335 gnd.n4608 gnd.n4607 585
R4336 gnd.n4607 gnd.n968 585
R4337 gnd.n4606 gnd.n2043 585
R4338 gnd.n4606 gnd.n961 585
R4339 gnd.n4605 gnd.n4604 585
R4340 gnd.n4605 gnd.n958 585
R4341 gnd.n2045 gnd.n2044 585
R4342 gnd.n2044 gnd.n950 585
R4343 gnd.n4600 gnd.n4599 585
R4344 gnd.n4599 gnd.n947 585
R4345 gnd.n4598 gnd.n2047 585
R4346 gnd.n4598 gnd.n4597 585
R4347 gnd.n4311 gnd.n2048 585
R4348 gnd.n2048 gnd.n938 585
R4349 gnd.n4312 gnd.n2062 585
R4350 gnd.n2062 gnd.n930 585
R4351 gnd.n4314 gnd.n4313 585
R4352 gnd.n4315 gnd.n4314 585
R4353 gnd.n2063 gnd.n2061 585
R4354 gnd.n2061 gnd.n921 585
R4355 gnd.n4305 gnd.n4304 585
R4356 gnd.n4304 gnd.n918 585
R4357 gnd.n4303 gnd.n2065 585
R4358 gnd.n4303 gnd.n910 585
R4359 gnd.n4302 gnd.n4301 585
R4360 gnd.n4302 gnd.n907 585
R4361 gnd.n4293 gnd.n4292 585
R4362 gnd.n4292 gnd.n4291 585
R4363 gnd.n4297 gnd.n4296 585
R4364 gnd.n4296 gnd.n896 585
R4365 gnd.n4295 gnd.n882 585
R4366 gnd.n886 gnd.n882 585
R4367 gnd.n5780 gnd.n5779 585
R4368 gnd.n5781 gnd.n5780 585
R4369 gnd.n1224 gnd.n1222 585
R4370 gnd.n1222 gnd.n1219 585
R4371 gnd.n5438 gnd.n5437 585
R4372 gnd.n5439 gnd.n5438 585
R4373 gnd.n1510 gnd.n1509 585
R4374 gnd.n1509 gnd.n1508 585
R4375 gnd.n5433 gnd.n5432 585
R4376 gnd.n5432 gnd.n5431 585
R4377 gnd.n1513 gnd.n1512 585
R4378 gnd.n1515 gnd.n1513 585
R4379 gnd.n5419 gnd.n5418 585
R4380 gnd.n5420 gnd.n5419 585
R4381 gnd.n1522 gnd.n1521 585
R4382 gnd.n1527 gnd.n1521 585
R4383 gnd.n5414 gnd.n5413 585
R4384 gnd.n5413 gnd.n5412 585
R4385 gnd.n1525 gnd.n1524 585
R4386 gnd.n1537 gnd.n1525 585
R4387 gnd.n1621 gnd.n1534 585
R4388 gnd.n5404 gnd.n1534 585
R4389 gnd.n5272 gnd.n5271 585
R4390 gnd.n5273 gnd.n5272 585
R4391 gnd.n1620 gnd.n1619 585
R4392 gnd.n1645 gnd.n1619 585
R4393 gnd.n5266 gnd.n5265 585
R4394 gnd.n5265 gnd.n5264 585
R4395 gnd.n1624 gnd.n1623 585
R4396 gnd.n1637 gnd.n1624 585
R4397 gnd.n4755 gnd.n1635 585
R4398 gnd.n5254 gnd.n1635 585
R4399 gnd.n4756 gnd.n4753 585
R4400 gnd.n4753 gnd.n1649 585
R4401 gnd.n4757 gnd.n1655 585
R4402 gnd.n5225 gnd.n1655 585
R4403 gnd.n4751 gnd.n4750 585
R4404 gnd.n4750 gnd.n1666 585
R4405 gnd.n4761 gnd.n1664 585
R4406 gnd.t189 gnd.n1664 585
R4407 gnd.n4762 gnd.n4749 585
R4408 gnd.n4749 gnd.n1670 585
R4409 gnd.n4763 gnd.n4748 585
R4410 gnd.n4748 gnd.n1677 585
R4411 gnd.n4746 gnd.n1683 585
R4412 gnd.n5192 gnd.n1683 585
R4413 gnd.n4767 gnd.n4745 585
R4414 gnd.n4745 gnd.n1681 585
R4415 gnd.n4768 gnd.n1693 585
R4416 gnd.n5182 gnd.n1693 585
R4417 gnd.n4769 gnd.n4744 585
R4418 gnd.n4744 gnd.n1701 585
R4419 gnd.n4743 gnd.n4741 585
R4420 gnd.n4743 gnd.n1699 585
R4421 gnd.n4773 gnd.n4740 585
R4422 gnd.n4740 gnd.n1706 585
R4423 gnd.n4774 gnd.n4739 585
R4424 gnd.n4739 gnd.n1712 585
R4425 gnd.n4775 gnd.n1717 585
R4426 gnd.n5152 gnd.n1717 585
R4427 gnd.n4737 gnd.n4736 585
R4428 gnd.n4736 gnd.n4735 585
R4429 gnd.n4779 gnd.n1725 585
R4430 gnd.n5136 gnd.n1725 585
R4431 gnd.n4780 gnd.n1733 585
R4432 gnd.n5128 gnd.n1733 585
R4433 gnd.n4781 gnd.n4734 585
R4434 gnd.n4734 gnd.n1737 585
R4435 gnd.n4732 gnd.n1743 585
R4436 gnd.n5108 gnd.n1743 585
R4437 gnd.n4785 gnd.n4731 585
R4438 gnd.n4731 gnd.n1741 585
R4439 gnd.n4786 gnd.n1750 585
R4440 gnd.n5098 gnd.n1750 585
R4441 gnd.n4787 gnd.n4730 585
R4442 gnd.n4730 gnd.n1755 585
R4443 gnd.n4728 gnd.n1762 585
R4444 gnd.n5081 gnd.n1762 585
R4445 gnd.n4791 gnd.n4727 585
R4446 gnd.n4727 gnd.n1772 585
R4447 gnd.n4792 gnd.n1770 585
R4448 gnd.n5073 gnd.n1770 585
R4449 gnd.n4793 gnd.n1777 585
R4450 gnd.n5066 gnd.n1777 585
R4451 gnd.n4725 gnd.n4724 585
R4452 gnd.n4724 gnd.n1784 585
R4453 gnd.n4797 gnd.n4723 585
R4454 gnd.n4723 gnd.n1783 585
R4455 gnd.n4798 gnd.n4722 585
R4456 gnd.n4722 gnd.n1788 585
R4457 gnd.n4799 gnd.n4721 585
R4458 gnd.n4721 gnd.n1795 585
R4459 gnd.n4719 gnd.n1801 585
R4460 gnd.n5034 gnd.n1801 585
R4461 gnd.n4803 gnd.n4718 585
R4462 gnd.n4718 gnd.n1799 585
R4463 gnd.n4804 gnd.n1808 585
R4464 gnd.n5015 gnd.n1808 585
R4465 gnd.n4805 gnd.n1816 585
R4466 gnd.n5007 gnd.n1816 585
R4467 gnd.n4716 gnd.n4715 585
R4468 gnd.n4715 gnd.n1819 585
R4469 gnd.n4809 gnd.n1825 585
R4470 gnd.n4986 gnd.n1825 585
R4471 gnd.n4810 gnd.n4714 585
R4472 gnd.n4714 gnd.n1823 585
R4473 gnd.n4811 gnd.n1832 585
R4474 gnd.n4976 gnd.n1832 585
R4475 gnd.n4712 gnd.n4711 585
R4476 gnd.n4711 gnd.n1836 585
R4477 gnd.n4815 gnd.n1843 585
R4478 gnd.n4958 gnd.n1843 585
R4479 gnd.n4816 gnd.n4710 585
R4480 gnd.n4710 gnd.n1852 585
R4481 gnd.n4817 gnd.n1850 585
R4482 gnd.n4950 gnd.n1850 585
R4483 gnd.n4708 gnd.n1856 585
R4484 gnd.n4942 gnd.n1856 585
R4485 gnd.n4821 gnd.n4707 585
R4486 gnd.n4707 gnd.n1864 585
R4487 gnd.n4822 gnd.n4706 585
R4488 gnd.n4706 gnd.n1862 585
R4489 gnd.n4823 gnd.n4705 585
R4490 gnd.n4705 gnd.n1869 585
R4491 gnd.n4704 gnd.n4702 585
R4492 gnd.n4704 gnd.n1875 585
R4493 gnd.n4827 gnd.n1881 585
R4494 gnd.t5 gnd.n1881 585
R4495 gnd.n4828 gnd.n4701 585
R4496 gnd.n4701 gnd.n1879 585
R4497 gnd.n4829 gnd.n1888 585
R4498 gnd.n4892 gnd.n1888 585
R4499 gnd.n4699 gnd.n1895 585
R4500 gnd.n4883 gnd.n1895 585
R4501 gnd.n4833 gnd.n1898 585
R4502 gnd.n4871 gnd.n1898 585
R4503 gnd.n4834 gnd.n1900 585
R4504 gnd.n4863 gnd.n1900 585
R4505 gnd.n4835 gnd.n4698 585
R4506 gnd.n4698 gnd.n1904 585
R4507 gnd.n1982 gnd.n1124 585
R4508 gnd.n5891 gnd.n1124 585
R4509 gnd.n4840 gnd.n4839 585
R4510 gnd.n4841 gnd.n4840 585
R4511 gnd.n1981 gnd.n1113 585
R4512 gnd.n5897 gnd.n1113 585
R4513 gnd.n4694 gnd.n4693 585
R4514 gnd.n4693 gnd.n1110 585
R4515 gnd.n4692 gnd.n1984 585
R4516 gnd.n4692 gnd.n1084 585
R4517 gnd.n4691 gnd.n4690 585
R4518 gnd.n4691 gnd.n1052 585
R4519 gnd.n1986 gnd.n1985 585
R4520 gnd.n1991 gnd.n1985 585
R4521 gnd.n4686 gnd.n4685 585
R4522 gnd.n4685 gnd.n4684 585
R4523 gnd.n1989 gnd.n1988 585
R4524 gnd.n1990 gnd.n1989 585
R4525 gnd.n4345 gnd.n2000 585
R4526 gnd.n4667 gnd.n2000 585
R4527 gnd.n4346 gnd.n4344 585
R4528 gnd.n4344 gnd.n1999 585
R4529 gnd.n4342 gnd.n2009 585
R4530 gnd.n4642 gnd.n2009 585
R4531 gnd.n4351 gnd.n4350 585
R4532 gnd.n4351 gnd.n2008 585
R4533 gnd.n4353 gnd.n4352 585
R4534 gnd.n4355 gnd.n4354 585
R4535 gnd.n4357 gnd.n4356 585
R4536 gnd.n4338 gnd.n4337 585
R4537 gnd.n4361 gnd.n4339 585
R4538 gnd.n4363 gnd.n4362 585
R4539 gnd.n4478 gnd.n4364 585
R4540 gnd.n4477 gnd.n4365 585
R4541 gnd.n4476 gnd.n4366 585
R4542 gnd.n4372 gnd.n4367 585
R4543 gnd.n4469 gnd.n4373 585
R4544 gnd.n4468 gnd.n4374 585
R4545 gnd.n4376 gnd.n4375 585
R4546 gnd.n4461 gnd.n4384 585
R4547 gnd.n4460 gnd.n4385 585
R4548 gnd.n4392 gnd.n4386 585
R4549 gnd.n4453 gnd.n4393 585
R4550 gnd.n4452 gnd.n4394 585
R4551 gnd.n4396 gnd.n4395 585
R4552 gnd.n4445 gnd.n4404 585
R4553 gnd.n4444 gnd.n4405 585
R4554 gnd.n4412 gnd.n4406 585
R4555 gnd.n4437 gnd.n4413 585
R4556 gnd.n4436 gnd.n4414 585
R4557 gnd.n4416 gnd.n4415 585
R4558 gnd.n4429 gnd.n4426 585
R4559 gnd.n4428 gnd.n4427 585
R4560 gnd.n2031 gnd.n2030 585
R4561 gnd.n4632 gnd.n4631 585
R4562 gnd.n4633 gnd.n4632 585
R4563 gnd.n5783 gnd.n5782 585
R4564 gnd.n5782 gnd.n5781 585
R4565 gnd.n1217 gnd.n1215 585
R4566 gnd.n1219 gnd.n1217 585
R4567 gnd.n5787 gnd.n1214 585
R4568 gnd.n5439 gnd.n1214 585
R4569 gnd.n5788 gnd.n1213 585
R4570 gnd.n1508 gnd.n1213 585
R4571 gnd.n5789 gnd.n1212 585
R4572 gnd.n5431 gnd.n1212 585
R4573 gnd.n1514 gnd.n1210 585
R4574 gnd.n1515 gnd.n1514 585
R4575 gnd.n5793 gnd.n1209 585
R4576 gnd.n5420 gnd.n1209 585
R4577 gnd.n5794 gnd.n1208 585
R4578 gnd.n1527 gnd.n1208 585
R4579 gnd.n5795 gnd.n1207 585
R4580 gnd.n5412 gnd.n1207 585
R4581 gnd.n1536 gnd.n1205 585
R4582 gnd.n1537 gnd.n1536 585
R4583 gnd.n5799 gnd.n1204 585
R4584 gnd.n5404 gnd.n1204 585
R4585 gnd.n5800 gnd.n1203 585
R4586 gnd.n5273 gnd.n1203 585
R4587 gnd.n5801 gnd.n1202 585
R4588 gnd.n1645 gnd.n1202 585
R4589 gnd.n1627 gnd.n1200 585
R4590 gnd.n5264 gnd.n1627 585
R4591 gnd.n5805 gnd.n1199 585
R4592 gnd.n1637 gnd.n1199 585
R4593 gnd.n5806 gnd.n1198 585
R4594 gnd.n5254 gnd.n1198 585
R4595 gnd.n5807 gnd.n1197 585
R4596 gnd.n1649 gnd.n1197 585
R4597 gnd.n1657 gnd.n1195 585
R4598 gnd.n5225 gnd.n1657 585
R4599 gnd.n5811 gnd.n1194 585
R4600 gnd.n1666 gnd.n1194 585
R4601 gnd.n5812 gnd.n1193 585
R4602 gnd.t189 gnd.n1193 585
R4603 gnd.n5813 gnd.n1192 585
R4604 gnd.n1670 gnd.n1192 585
R4605 gnd.n1676 gnd.n1190 585
R4606 gnd.n1677 gnd.n1676 585
R4607 gnd.n5817 gnd.n1189 585
R4608 gnd.n5192 gnd.n1189 585
R4609 gnd.n5818 gnd.n1188 585
R4610 gnd.n1681 gnd.n1188 585
R4611 gnd.n5819 gnd.n1187 585
R4612 gnd.n5182 gnd.n1187 585
R4613 gnd.n1700 gnd.n1185 585
R4614 gnd.n1701 gnd.n1700 585
R4615 gnd.n5823 gnd.n1184 585
R4616 gnd.n1699 gnd.n1184 585
R4617 gnd.n5824 gnd.n1183 585
R4618 gnd.n1706 gnd.n1183 585
R4619 gnd.n5825 gnd.n1182 585
R4620 gnd.n1712 gnd.n1182 585
R4621 gnd.n1718 gnd.n1180 585
R4622 gnd.n5152 gnd.n1718 585
R4623 gnd.n5829 gnd.n1179 585
R4624 gnd.n4735 gnd.n1179 585
R4625 gnd.n5830 gnd.n1178 585
R4626 gnd.n5136 gnd.n1178 585
R4627 gnd.n5831 gnd.n1177 585
R4628 gnd.n5128 gnd.n1177 585
R4629 gnd.n1736 gnd.n1175 585
R4630 gnd.n1737 gnd.n1736 585
R4631 gnd.n5835 gnd.n1174 585
R4632 gnd.n5108 gnd.n1174 585
R4633 gnd.n5836 gnd.n1173 585
R4634 gnd.n1741 gnd.n1173 585
R4635 gnd.n5837 gnd.n1172 585
R4636 gnd.n5098 gnd.n1172 585
R4637 gnd.n1754 gnd.n1170 585
R4638 gnd.n1755 gnd.n1754 585
R4639 gnd.n5841 gnd.n1169 585
R4640 gnd.n5081 gnd.n1169 585
R4641 gnd.n5842 gnd.n1168 585
R4642 gnd.n1772 gnd.n1168 585
R4643 gnd.n5843 gnd.n1167 585
R4644 gnd.n5073 gnd.n1167 585
R4645 gnd.n1778 gnd.n1165 585
R4646 gnd.n5066 gnd.n1778 585
R4647 gnd.n5847 gnd.n1164 585
R4648 gnd.n1784 gnd.n1164 585
R4649 gnd.n5848 gnd.n1163 585
R4650 gnd.n1783 gnd.n1163 585
R4651 gnd.n5849 gnd.n1162 585
R4652 gnd.n1788 gnd.n1162 585
R4653 gnd.n1794 gnd.n1160 585
R4654 gnd.n1795 gnd.n1794 585
R4655 gnd.n5853 gnd.n1159 585
R4656 gnd.n5034 gnd.n1159 585
R4657 gnd.n5854 gnd.n1158 585
R4658 gnd.n1799 gnd.n1158 585
R4659 gnd.n5855 gnd.n1157 585
R4660 gnd.n5015 gnd.n1157 585
R4661 gnd.n5006 gnd.n1155 585
R4662 gnd.n5007 gnd.n5006 585
R4663 gnd.n5859 gnd.n1154 585
R4664 gnd.n1819 gnd.n1154 585
R4665 gnd.n5860 gnd.n1153 585
R4666 gnd.n4986 gnd.n1153 585
R4667 gnd.n5861 gnd.n1152 585
R4668 gnd.n1823 gnd.n1152 585
R4669 gnd.n4975 gnd.n1150 585
R4670 gnd.n4976 gnd.n4975 585
R4671 gnd.n5865 gnd.n1149 585
R4672 gnd.n1836 gnd.n1149 585
R4673 gnd.n5866 gnd.n1148 585
R4674 gnd.n4958 gnd.n1148 585
R4675 gnd.n5867 gnd.n1147 585
R4676 gnd.n1852 gnd.n1147 585
R4677 gnd.n4949 gnd.n1145 585
R4678 gnd.n4950 gnd.n4949 585
R4679 gnd.n5871 gnd.n1144 585
R4680 gnd.n4942 gnd.n1144 585
R4681 gnd.n5872 gnd.n1143 585
R4682 gnd.n1864 gnd.n1143 585
R4683 gnd.n5873 gnd.n1142 585
R4684 gnd.n1862 gnd.n1142 585
R4685 gnd.n1868 gnd.n1140 585
R4686 gnd.n1869 gnd.n1868 585
R4687 gnd.n5877 gnd.n1139 585
R4688 gnd.n1875 gnd.n1139 585
R4689 gnd.n5878 gnd.n1138 585
R4690 gnd.t5 gnd.n1138 585
R4691 gnd.n5879 gnd.n1137 585
R4692 gnd.n1879 gnd.n1137 585
R4693 gnd.n4891 gnd.n1135 585
R4694 gnd.n4892 gnd.n4891 585
R4695 gnd.n5883 gnd.n1134 585
R4696 gnd.n4883 gnd.n1134 585
R4697 gnd.n5884 gnd.n1133 585
R4698 gnd.n4871 gnd.n1133 585
R4699 gnd.n5885 gnd.n1132 585
R4700 gnd.n4863 gnd.n1132 585
R4701 gnd.n1129 gnd.n1127 585
R4702 gnd.n1904 gnd.n1127 585
R4703 gnd.n5890 gnd.n5889 585
R4704 gnd.n5891 gnd.n5890 585
R4705 gnd.n1128 gnd.n1126 585
R4706 gnd.n4841 gnd.n1126 585
R4707 gnd.n4654 gnd.n1115 585
R4708 gnd.n5897 gnd.n1115 585
R4709 gnd.n4655 gnd.n4653 585
R4710 gnd.n4653 gnd.n1110 585
R4711 gnd.n4652 gnd.n4650 585
R4712 gnd.n4652 gnd.n1084 585
R4713 gnd.n4659 gnd.n4649 585
R4714 gnd.n4649 gnd.n1052 585
R4715 gnd.n4660 gnd.n4648 585
R4716 gnd.n4648 gnd.n1991 585
R4717 gnd.n4661 gnd.n1992 585
R4718 gnd.n4684 gnd.n1992 585
R4719 gnd.n2004 gnd.n2002 585
R4720 gnd.n2002 gnd.n1990 585
R4721 gnd.n4666 gnd.n4665 585
R4722 gnd.n4667 gnd.n4666 585
R4723 gnd.n2003 gnd.n2001 585
R4724 gnd.n2001 gnd.n1999 585
R4725 gnd.n4644 gnd.n4643 585
R4726 gnd.n4643 gnd.n4642 585
R4727 gnd.n2007 gnd.n2006 585
R4728 gnd.n2008 gnd.n2007 585
R4729 gnd.n5722 gnd.n1279 585
R4730 gnd.n5723 gnd.n1278 585
R4731 gnd.n1496 gnd.n1272 585
R4732 gnd.n5730 gnd.n1271 585
R4733 gnd.n5731 gnd.n1270 585
R4734 gnd.n1493 gnd.n1264 585
R4735 gnd.n5738 gnd.n1263 585
R4736 gnd.n5739 gnd.n1262 585
R4737 gnd.n1491 gnd.n1256 585
R4738 gnd.n5746 gnd.n1255 585
R4739 gnd.n5747 gnd.n1254 585
R4740 gnd.n1488 gnd.n1248 585
R4741 gnd.n5754 gnd.n1247 585
R4742 gnd.n5755 gnd.n1246 585
R4743 gnd.n1486 gnd.n1239 585
R4744 gnd.n5762 gnd.n1238 585
R4745 gnd.n5763 gnd.n1237 585
R4746 gnd.n1483 gnd.n1234 585
R4747 gnd.n5768 gnd.n1233 585
R4748 gnd.n5769 gnd.n1232 585
R4749 gnd.n5770 gnd.n1231 585
R4750 gnd.n1480 gnd.n1229 585
R4751 gnd.n5774 gnd.n1228 585
R4752 gnd.n5775 gnd.n1227 585
R4753 gnd.n5776 gnd.n1223 585
R4754 gnd.n5463 gnd.n1218 585
R4755 gnd.n5460 gnd.n1218 585
R4756 gnd.n5464 gnd.n5462 585
R4757 gnd.n1478 gnd.n1477 585
R4758 gnd.n1499 gnd.n1498 585
R4759 gnd.n5398 gnd.n5397 468.476
R4760 gnd.n5281 gnd.n5280 468.476
R4761 gnd.n1974 gnd.n1972 468.476
R4762 gnd.n5967 gnd.n1087 468.476
R4763 gnd.n1908 gnd.t145 389.64
R4764 gnd.n1591 gnd.t110 389.64
R4765 gnd.n5904 gnd.t69 389.64
R4766 gnd.n1585 gnd.t154 389.64
R4767 gnd.n4423 gnd.t83 371.625
R4768 gnd.n5716 gnd.t142 371.625
R4769 gnd.n306 gnd.t163 371.625
R4770 gnd.n286 gnd.t73 371.625
R4771 gnd.n7148 gnd.t120 371.625
R4772 gnd.n1352 gnd.t139 371.625
R4773 gnd.n1375 gnd.t129 371.625
R4774 gnd.n5596 gnd.t61 371.625
R4775 gnd.n6967 gnd.t114 371.625
R4776 gnd.n2034 gnd.t166 371.625
R4777 gnd.n3841 gnd.t151 371.625
R4778 gnd.n3780 gnd.t97 371.625
R4779 gnd.n3802 gnd.t94 371.625
R4780 gnd.n3823 gnd.t65 371.625
R4781 gnd.n1035 gnd.t157 371.625
R4782 gnd.n4482 gnd.t90 371.625
R4783 gnd.n4495 gnd.t117 371.625
R4784 gnd.n1280 gnd.t100 371.625
R4785 gnd.n6248 gnd.n711 345.092
R4786 gnd.n2742 gnd.t135 323.425
R4787 gnd.n2283 gnd.t169 323.425
R4788 gnd.n3590 gnd.n3564 289.615
R4789 gnd.n3558 gnd.n3532 289.615
R4790 gnd.n3526 gnd.n3500 289.615
R4791 gnd.n3495 gnd.n3469 289.615
R4792 gnd.n3463 gnd.n3437 289.615
R4793 gnd.n3431 gnd.n3405 289.615
R4794 gnd.n3399 gnd.n3373 289.615
R4795 gnd.n3368 gnd.n3342 289.615
R4796 gnd.n2816 gnd.t57 279.217
R4797 gnd.n2309 gnd.t53 279.217
R4798 gnd.n1094 gnd.t79 260.649
R4799 gnd.n1553 gnd.t125 260.649
R4800 gnd.n5969 gnd.n5968 256.663
R4801 gnd.n5969 gnd.n1053 256.663
R4802 gnd.n5969 gnd.n1054 256.663
R4803 gnd.n5969 gnd.n1055 256.663
R4804 gnd.n5969 gnd.n1056 256.663
R4805 gnd.n5969 gnd.n1057 256.663
R4806 gnd.n5969 gnd.n1058 256.663
R4807 gnd.n5969 gnd.n1059 256.663
R4808 gnd.n5969 gnd.n1060 256.663
R4809 gnd.n5969 gnd.n1061 256.663
R4810 gnd.n5969 gnd.n1062 256.663
R4811 gnd.n5969 gnd.n1063 256.663
R4812 gnd.n5969 gnd.n1064 256.663
R4813 gnd.n5969 gnd.n1065 256.663
R4814 gnd.n5969 gnd.n1066 256.663
R4815 gnd.n5969 gnd.n1067 256.663
R4816 gnd.n5972 gnd.n1050 256.663
R4817 gnd.n5970 gnd.n5969 256.663
R4818 gnd.n5969 gnd.n1068 256.663
R4819 gnd.n5969 gnd.n1069 256.663
R4820 gnd.n5969 gnd.n1070 256.663
R4821 gnd.n5969 gnd.n1071 256.663
R4822 gnd.n5969 gnd.n1072 256.663
R4823 gnd.n5969 gnd.n1073 256.663
R4824 gnd.n5969 gnd.n1074 256.663
R4825 gnd.n5969 gnd.n1075 256.663
R4826 gnd.n5969 gnd.n1076 256.663
R4827 gnd.n5969 gnd.n1077 256.663
R4828 gnd.n5969 gnd.n1078 256.663
R4829 gnd.n5969 gnd.n1079 256.663
R4830 gnd.n5969 gnd.n1080 256.663
R4831 gnd.n5969 gnd.n1081 256.663
R4832 gnd.n5969 gnd.n1082 256.663
R4833 gnd.n5969 gnd.n1083 256.663
R4834 gnd.n1615 gnd.n1528 256.663
R4835 gnd.n5286 gnd.n1528 256.663
R4836 gnd.n1612 gnd.n1528 256.663
R4837 gnd.n5293 gnd.n1528 256.663
R4838 gnd.n1609 gnd.n1528 256.663
R4839 gnd.n5300 gnd.n1528 256.663
R4840 gnd.n1606 gnd.n1528 256.663
R4841 gnd.n5307 gnd.n1528 256.663
R4842 gnd.n1603 gnd.n1528 256.663
R4843 gnd.n5314 gnd.n1528 256.663
R4844 gnd.n1600 gnd.n1528 256.663
R4845 gnd.n5321 gnd.n1528 256.663
R4846 gnd.n1597 gnd.n1528 256.663
R4847 gnd.n5328 gnd.n1528 256.663
R4848 gnd.n1594 gnd.n1528 256.663
R4849 gnd.n5336 gnd.n1528 256.663
R4850 gnd.n5339 gnd.n1362 256.663
R4851 gnd.n5340 gnd.n1528 256.663
R4852 gnd.n1588 gnd.n1528 256.663
R4853 gnd.n5347 gnd.n1528 256.663
R4854 gnd.n1583 gnd.n1528 256.663
R4855 gnd.n5354 gnd.n1528 256.663
R4856 gnd.n1580 gnd.n1528 256.663
R4857 gnd.n5361 gnd.n1528 256.663
R4858 gnd.n1577 gnd.n1528 256.663
R4859 gnd.n5368 gnd.n1528 256.663
R4860 gnd.n1574 gnd.n1528 256.663
R4861 gnd.n5375 gnd.n1528 256.663
R4862 gnd.n1571 gnd.n1528 256.663
R4863 gnd.n5382 gnd.n1528 256.663
R4864 gnd.n1568 gnd.n1528 256.663
R4865 gnd.n5389 gnd.n1528 256.663
R4866 gnd.n1565 gnd.n1528 256.663
R4867 gnd.n5396 gnd.n1528 256.663
R4868 gnd.n4036 gnd.n3750 242.672
R4869 gnd.n4036 gnd.n3751 242.672
R4870 gnd.n4036 gnd.n3752 242.672
R4871 gnd.n4036 gnd.n3753 242.672
R4872 gnd.n4036 gnd.n3754 242.672
R4873 gnd.n4036 gnd.n3755 242.672
R4874 gnd.n4036 gnd.n3756 242.672
R4875 gnd.n4036 gnd.n3757 242.672
R4876 gnd.n4036 gnd.n3758 242.672
R4877 gnd.n6023 gnd.n988 242.672
R4878 gnd.n6023 gnd.n987 242.672
R4879 gnd.n6023 gnd.n986 242.672
R4880 gnd.n6023 gnd.n985 242.672
R4881 gnd.n6023 gnd.n984 242.672
R4882 gnd.n6023 gnd.n983 242.672
R4883 gnd.n6023 gnd.n982 242.672
R4884 gnd.n6023 gnd.n981 242.672
R4885 gnd.n6023 gnd.n980 242.672
R4886 gnd.n2870 gnd.n2869 242.672
R4887 gnd.n2870 gnd.n2780 242.672
R4888 gnd.n2870 gnd.n2781 242.672
R4889 gnd.n2870 gnd.n2782 242.672
R4890 gnd.n2870 gnd.n2783 242.672
R4891 gnd.n2870 gnd.n2784 242.672
R4892 gnd.n2870 gnd.n2785 242.672
R4893 gnd.n2870 gnd.n2786 242.672
R4894 gnd.n2870 gnd.n2787 242.672
R4895 gnd.n2870 gnd.n2788 242.672
R4896 gnd.n2870 gnd.n2789 242.672
R4897 gnd.n2870 gnd.n2790 242.672
R4898 gnd.n2871 gnd.n2870 242.672
R4899 gnd.n3722 gnd.n2258 242.672
R4900 gnd.n3722 gnd.n2257 242.672
R4901 gnd.n3722 gnd.n2256 242.672
R4902 gnd.n3722 gnd.n2255 242.672
R4903 gnd.n3722 gnd.n2254 242.672
R4904 gnd.n3722 gnd.n2253 242.672
R4905 gnd.n3722 gnd.n2252 242.672
R4906 gnd.n3722 gnd.n2251 242.672
R4907 gnd.n3722 gnd.n2250 242.672
R4908 gnd.n3722 gnd.n2249 242.672
R4909 gnd.n3722 gnd.n2248 242.672
R4910 gnd.n3722 gnd.n2247 242.672
R4911 gnd.n3722 gnd.n2246 242.672
R4912 gnd.n5713 gnd.n1317 242.672
R4913 gnd.n5713 gnd.n1319 242.672
R4914 gnd.n5713 gnd.n1320 242.672
R4915 gnd.n5713 gnd.n1322 242.672
R4916 gnd.n5713 gnd.n1324 242.672
R4917 gnd.n5713 gnd.n1325 242.672
R4918 gnd.n5713 gnd.n1327 242.672
R4919 gnd.n5713 gnd.n1329 242.672
R4920 gnd.n5714 gnd.n5713 242.672
R4921 gnd.n7183 gnd.n220 242.672
R4922 gnd.n7183 gnd.n219 242.672
R4923 gnd.n7183 gnd.n218 242.672
R4924 gnd.n7183 gnd.n217 242.672
R4925 gnd.n7183 gnd.n216 242.672
R4926 gnd.n7183 gnd.n215 242.672
R4927 gnd.n7183 gnd.n214 242.672
R4928 gnd.n7183 gnd.n213 242.672
R4929 gnd.n7183 gnd.n212 242.672
R4930 gnd.n2954 gnd.n2953 242.672
R4931 gnd.n2953 gnd.n2692 242.672
R4932 gnd.n2953 gnd.n2693 242.672
R4933 gnd.n2953 gnd.n2694 242.672
R4934 gnd.n2953 gnd.n2695 242.672
R4935 gnd.n2953 gnd.n2696 242.672
R4936 gnd.n2953 gnd.n2697 242.672
R4937 gnd.n2953 gnd.n2698 242.672
R4938 gnd.n3722 gnd.n2259 242.672
R4939 gnd.n3722 gnd.n2260 242.672
R4940 gnd.n3722 gnd.n2261 242.672
R4941 gnd.n3722 gnd.n2262 242.672
R4942 gnd.n3722 gnd.n2263 242.672
R4943 gnd.n3722 gnd.n2264 242.672
R4944 gnd.n3722 gnd.n2265 242.672
R4945 gnd.n3722 gnd.n2266 242.672
R4946 gnd.n4036 gnd.n4035 242.672
R4947 gnd.n4036 gnd.n3723 242.672
R4948 gnd.n4036 gnd.n3724 242.672
R4949 gnd.n4036 gnd.n3725 242.672
R4950 gnd.n4036 gnd.n3726 242.672
R4951 gnd.n4036 gnd.n3727 242.672
R4952 gnd.n4036 gnd.n3728 242.672
R4953 gnd.n4036 gnd.n3729 242.672
R4954 gnd.n4036 gnd.n3730 242.672
R4955 gnd.n4036 gnd.n3731 242.672
R4956 gnd.n4036 gnd.n3732 242.672
R4957 gnd.n4036 gnd.n3733 242.672
R4958 gnd.n4036 gnd.n3734 242.672
R4959 gnd.n4036 gnd.n3735 242.672
R4960 gnd.n4036 gnd.n3736 242.672
R4961 gnd.n4036 gnd.n3737 242.672
R4962 gnd.n4036 gnd.n3738 242.672
R4963 gnd.n4036 gnd.n3739 242.672
R4964 gnd.n4036 gnd.n3740 242.672
R4965 gnd.n4036 gnd.n3741 242.672
R4966 gnd.n4036 gnd.n3742 242.672
R4967 gnd.n4036 gnd.n3743 242.672
R4968 gnd.n4036 gnd.n3744 242.672
R4969 gnd.n4036 gnd.n3745 242.672
R4970 gnd.n4036 gnd.n3746 242.672
R4971 gnd.n4036 gnd.n3747 242.672
R4972 gnd.n4036 gnd.n3748 242.672
R4973 gnd.n4036 gnd.n3749 242.672
R4974 gnd.n4037 gnd.n4036 242.672
R4975 gnd.n6023 gnd.n990 242.672
R4976 gnd.n6023 gnd.n991 242.672
R4977 gnd.n6023 gnd.n992 242.672
R4978 gnd.n6023 gnd.n993 242.672
R4979 gnd.n6023 gnd.n994 242.672
R4980 gnd.n6023 gnd.n995 242.672
R4981 gnd.n6023 gnd.n996 242.672
R4982 gnd.n6023 gnd.n997 242.672
R4983 gnd.n6023 gnd.n998 242.672
R4984 gnd.n6023 gnd.n999 242.672
R4985 gnd.n6023 gnd.n1000 242.672
R4986 gnd.n6023 gnd.n1001 242.672
R4987 gnd.n6023 gnd.n1002 242.672
R4988 gnd.n6023 gnd.n1003 242.672
R4989 gnd.n6023 gnd.n1004 242.672
R4990 gnd.n6023 gnd.n1005 242.672
R4991 gnd.n5973 gnd.n1046 242.672
R4992 gnd.n6023 gnd.n1006 242.672
R4993 gnd.n6023 gnd.n1007 242.672
R4994 gnd.n6023 gnd.n1008 242.672
R4995 gnd.n6023 gnd.n1009 242.672
R4996 gnd.n6023 gnd.n1010 242.672
R4997 gnd.n6023 gnd.n1011 242.672
R4998 gnd.n6023 gnd.n1012 242.672
R4999 gnd.n6023 gnd.n1013 242.672
R5000 gnd.n6023 gnd.n1014 242.672
R5001 gnd.n6023 gnd.n1015 242.672
R5002 gnd.n6023 gnd.n1016 242.672
R5003 gnd.n6023 gnd.n1017 242.672
R5004 gnd.n6023 gnd.n6022 242.672
R5005 gnd.n5713 gnd.n5712 242.672
R5006 gnd.n5713 gnd.n1289 242.672
R5007 gnd.n5713 gnd.n1290 242.672
R5008 gnd.n5713 gnd.n1291 242.672
R5009 gnd.n5713 gnd.n1292 242.672
R5010 gnd.n5713 gnd.n1293 242.672
R5011 gnd.n5713 gnd.n1294 242.672
R5012 gnd.n5713 gnd.n1295 242.672
R5013 gnd.n5713 gnd.n1296 242.672
R5014 gnd.n5713 gnd.n1297 242.672
R5015 gnd.n5713 gnd.n1298 242.672
R5016 gnd.n5713 gnd.n1299 242.672
R5017 gnd.n5713 gnd.n1300 242.672
R5018 gnd.n5660 gnd.n1363 242.672
R5019 gnd.n5713 gnd.n1301 242.672
R5020 gnd.n5713 gnd.n1302 242.672
R5021 gnd.n5713 gnd.n1303 242.672
R5022 gnd.n5713 gnd.n1304 242.672
R5023 gnd.n5713 gnd.n1305 242.672
R5024 gnd.n5713 gnd.n1306 242.672
R5025 gnd.n5713 gnd.n1307 242.672
R5026 gnd.n5713 gnd.n1308 242.672
R5027 gnd.n5713 gnd.n1309 242.672
R5028 gnd.n5713 gnd.n1310 242.672
R5029 gnd.n5713 gnd.n1311 242.672
R5030 gnd.n5713 gnd.n1312 242.672
R5031 gnd.n5713 gnd.n1313 242.672
R5032 gnd.n5713 gnd.n1314 242.672
R5033 gnd.n5713 gnd.n1315 242.672
R5034 gnd.n5713 gnd.n1316 242.672
R5035 gnd.n7183 gnd.n221 242.672
R5036 gnd.n7183 gnd.n222 242.672
R5037 gnd.n7183 gnd.n223 242.672
R5038 gnd.n7183 gnd.n224 242.672
R5039 gnd.n7183 gnd.n225 242.672
R5040 gnd.n7183 gnd.n226 242.672
R5041 gnd.n7183 gnd.n227 242.672
R5042 gnd.n7183 gnd.n228 242.672
R5043 gnd.n7183 gnd.n229 242.672
R5044 gnd.n7183 gnd.n230 242.672
R5045 gnd.n7183 gnd.n231 242.672
R5046 gnd.n7183 gnd.n232 242.672
R5047 gnd.n7183 gnd.n233 242.672
R5048 gnd.n7183 gnd.n234 242.672
R5049 gnd.n7183 gnd.n235 242.672
R5050 gnd.n7183 gnd.n236 242.672
R5051 gnd.n7183 gnd.n237 242.672
R5052 gnd.n7183 gnd.n238 242.672
R5053 gnd.n7183 gnd.n239 242.672
R5054 gnd.n7183 gnd.n240 242.672
R5055 gnd.n7183 gnd.n241 242.672
R5056 gnd.n7183 gnd.n242 242.672
R5057 gnd.n7183 gnd.n243 242.672
R5058 gnd.n7183 gnd.n244 242.672
R5059 gnd.n7183 gnd.n245 242.672
R5060 gnd.n7183 gnd.n246 242.672
R5061 gnd.n7183 gnd.n247 242.672
R5062 gnd.n7183 gnd.n248 242.672
R5063 gnd.n7183 gnd.n7182 242.672
R5064 gnd.n4633 gnd.n2016 242.672
R5065 gnd.n4633 gnd.n2017 242.672
R5066 gnd.n4633 gnd.n2018 242.672
R5067 gnd.n4633 gnd.n2019 242.672
R5068 gnd.n4633 gnd.n2020 242.672
R5069 gnd.n4633 gnd.n2021 242.672
R5070 gnd.n4633 gnd.n2022 242.672
R5071 gnd.n4633 gnd.n2023 242.672
R5072 gnd.n4633 gnd.n2024 242.672
R5073 gnd.n4633 gnd.n2025 242.672
R5074 gnd.n4633 gnd.n2026 242.672
R5075 gnd.n4633 gnd.n2027 242.672
R5076 gnd.n4633 gnd.n2028 242.672
R5077 gnd.n4633 gnd.n2029 242.672
R5078 gnd.n5460 gnd.n1500 242.672
R5079 gnd.n5460 gnd.n1497 242.672
R5080 gnd.n5460 gnd.n1495 242.672
R5081 gnd.n5460 gnd.n1494 242.672
R5082 gnd.n5460 gnd.n1492 242.672
R5083 gnd.n5460 gnd.n1490 242.672
R5084 gnd.n5460 gnd.n1489 242.672
R5085 gnd.n5460 gnd.n1487 242.672
R5086 gnd.n5460 gnd.n1485 242.672
R5087 gnd.n5460 gnd.n1484 242.672
R5088 gnd.n5460 gnd.n1482 242.672
R5089 gnd.n5460 gnd.n1481 242.672
R5090 gnd.n5460 gnd.n1479 242.672
R5091 gnd.n5461 gnd.n5460 242.672
R5092 gnd.n7184 gnd.n210 240.244
R5093 gnd.n7181 gnd.n249 240.244
R5094 gnd.n7177 gnd.n7176 240.244
R5095 gnd.n7173 gnd.n7172 240.244
R5096 gnd.n7169 gnd.n7168 240.244
R5097 gnd.n7165 gnd.n7164 240.244
R5098 gnd.n7161 gnd.n7160 240.244
R5099 gnd.n7157 gnd.n7156 240.244
R5100 gnd.n7153 gnd.n7152 240.244
R5101 gnd.n7146 gnd.n7145 240.244
R5102 gnd.n7142 gnd.n7141 240.244
R5103 gnd.n7138 gnd.n7137 240.244
R5104 gnd.n7134 gnd.n7133 240.244
R5105 gnd.n7130 gnd.n7129 240.244
R5106 gnd.n7126 gnd.n7125 240.244
R5107 gnd.n7122 gnd.n7121 240.244
R5108 gnd.n7118 gnd.n7117 240.244
R5109 gnd.n7114 gnd.n7113 240.244
R5110 gnd.n7110 gnd.n7109 240.244
R5111 gnd.n7103 gnd.n7102 240.244
R5112 gnd.n7100 gnd.n7099 240.244
R5113 gnd.n7096 gnd.n7095 240.244
R5114 gnd.n7092 gnd.n7091 240.244
R5115 gnd.n7088 gnd.n7087 240.244
R5116 gnd.n7084 gnd.n7083 240.244
R5117 gnd.n7080 gnd.n7079 240.244
R5118 gnd.n7076 gnd.n7075 240.244
R5119 gnd.n7072 gnd.n7071 240.244
R5120 gnd.n7068 gnd.n7067 240.244
R5121 gnd.n5593 gnd.n1396 240.244
R5122 gnd.n1408 gnd.n1396 240.244
R5123 gnd.n5481 gnd.n1408 240.244
R5124 gnd.n5481 gnd.n1423 240.244
R5125 gnd.n5485 gnd.n1423 240.244
R5126 gnd.n5485 gnd.n1433 240.244
R5127 gnd.n5490 gnd.n1433 240.244
R5128 gnd.n5490 gnd.n1444 240.244
R5129 gnd.n5494 gnd.n1444 240.244
R5130 gnd.n5494 gnd.n1454 240.244
R5131 gnd.n1457 gnd.n1454 240.244
R5132 gnd.n5501 gnd.n1457 240.244
R5133 gnd.n5501 gnd.n380 240.244
R5134 gnd.n6795 gnd.n380 240.244
R5135 gnd.n6795 gnd.n370 240.244
R5136 gnd.n370 gnd.n362 240.244
R5137 gnd.n6827 gnd.n362 240.244
R5138 gnd.n6827 gnd.n352 240.244
R5139 gnd.n6830 gnd.n352 240.244
R5140 gnd.n6830 gnd.n343 240.244
R5141 gnd.n343 gnd.n335 240.244
R5142 gnd.n6866 gnd.n335 240.244
R5143 gnd.n6866 gnd.n329 240.244
R5144 gnd.n6868 gnd.n329 240.244
R5145 gnd.n6868 gnd.n320 240.244
R5146 gnd.n320 gnd.n314 240.244
R5147 gnd.n6892 gnd.n314 240.244
R5148 gnd.n6892 gnd.n85 240.244
R5149 gnd.n6899 gnd.n85 240.244
R5150 gnd.n6899 gnd.n96 240.244
R5151 gnd.n6902 gnd.n96 240.244
R5152 gnd.n6902 gnd.n107 240.244
R5153 gnd.n6906 gnd.n107 240.244
R5154 gnd.n6906 gnd.n117 240.244
R5155 gnd.n6909 gnd.n117 240.244
R5156 gnd.n6909 gnd.n126 240.244
R5157 gnd.n6913 gnd.n126 240.244
R5158 gnd.n6913 gnd.n136 240.244
R5159 gnd.n6916 gnd.n136 240.244
R5160 gnd.n6916 gnd.n145 240.244
R5161 gnd.n6920 gnd.n145 240.244
R5162 gnd.n6920 gnd.n155 240.244
R5163 gnd.n7042 gnd.n155 240.244
R5164 gnd.n7042 gnd.n164 240.244
R5165 gnd.n7046 gnd.n164 240.244
R5166 gnd.n7046 gnd.n174 240.244
R5167 gnd.n7049 gnd.n174 240.244
R5168 gnd.n7049 gnd.n183 240.244
R5169 gnd.n7053 gnd.n183 240.244
R5170 gnd.n7053 gnd.n193 240.244
R5171 gnd.n7056 gnd.n193 240.244
R5172 gnd.n7056 gnd.n202 240.244
R5173 gnd.n7060 gnd.n202 240.244
R5174 gnd.n1332 gnd.n1331 240.244
R5175 gnd.n5706 gnd.n1331 240.244
R5176 gnd.n5704 gnd.n5703 240.244
R5177 gnd.n5700 gnd.n5699 240.244
R5178 gnd.n5696 gnd.n5695 240.244
R5179 gnd.n5692 gnd.n5691 240.244
R5180 gnd.n5688 gnd.n5687 240.244
R5181 gnd.n5684 gnd.n5683 240.244
R5182 gnd.n5680 gnd.n5679 240.244
R5183 gnd.n5675 gnd.n5674 240.244
R5184 gnd.n5671 gnd.n5670 240.244
R5185 gnd.n5667 gnd.n5666 240.244
R5186 gnd.n5663 gnd.n5662 240.244
R5187 gnd.n5658 gnd.n5657 240.244
R5188 gnd.n5654 gnd.n5653 240.244
R5189 gnd.n5650 gnd.n5649 240.244
R5190 gnd.n5646 gnd.n5645 240.244
R5191 gnd.n5642 gnd.n5641 240.244
R5192 gnd.n5638 gnd.n5637 240.244
R5193 gnd.n5634 gnd.n5633 240.244
R5194 gnd.n5630 gnd.n5629 240.244
R5195 gnd.n5626 gnd.n5625 240.244
R5196 gnd.n5622 gnd.n5621 240.244
R5197 gnd.n5618 gnd.n5617 240.244
R5198 gnd.n5614 gnd.n5613 240.244
R5199 gnd.n5610 gnd.n5609 240.244
R5200 gnd.n5606 gnd.n5605 240.244
R5201 gnd.n5602 gnd.n5601 240.244
R5202 gnd.n1411 gnd.n1333 240.244
R5203 gnd.n5585 gnd.n1411 240.244
R5204 gnd.n5585 gnd.n1412 240.244
R5205 gnd.n5581 gnd.n1412 240.244
R5206 gnd.n5581 gnd.n1421 240.244
R5207 gnd.n5573 gnd.n1421 240.244
R5208 gnd.n5573 gnd.n1436 240.244
R5209 gnd.n5569 gnd.n1436 240.244
R5210 gnd.n5569 gnd.n1442 240.244
R5211 gnd.n5561 gnd.n1442 240.244
R5212 gnd.n5561 gnd.n5555 240.244
R5213 gnd.n5555 gnd.n378 240.244
R5214 gnd.n6808 gnd.n378 240.244
R5215 gnd.n6808 gnd.n373 240.244
R5216 gnd.n6816 gnd.n373 240.244
R5217 gnd.n6816 gnd.n374 240.244
R5218 gnd.n374 gnd.n350 240.244
R5219 gnd.n6842 gnd.n350 240.244
R5220 gnd.n6842 gnd.n345 240.244
R5221 gnd.n6850 gnd.n345 240.244
R5222 gnd.n6850 gnd.n346 240.244
R5223 gnd.n346 gnd.n328 240.244
R5224 gnd.n6875 gnd.n328 240.244
R5225 gnd.n6875 gnd.n323 240.244
R5226 gnd.n6884 gnd.n323 240.244
R5227 gnd.n6884 gnd.n324 240.244
R5228 gnd.n324 gnd.n88 240.244
R5229 gnd.n7262 gnd.n88 240.244
R5230 gnd.n7262 gnd.n89 240.244
R5231 gnd.n7258 gnd.n89 240.244
R5232 gnd.n7258 gnd.n95 240.244
R5233 gnd.n7250 gnd.n95 240.244
R5234 gnd.n7250 gnd.n110 240.244
R5235 gnd.n7246 gnd.n110 240.244
R5236 gnd.n7246 gnd.n116 240.244
R5237 gnd.n7238 gnd.n116 240.244
R5238 gnd.n7238 gnd.n129 240.244
R5239 gnd.n7234 gnd.n129 240.244
R5240 gnd.n7234 gnd.n135 240.244
R5241 gnd.n7226 gnd.n135 240.244
R5242 gnd.n7226 gnd.n148 240.244
R5243 gnd.n7222 gnd.n148 240.244
R5244 gnd.n7222 gnd.n154 240.244
R5245 gnd.n7214 gnd.n154 240.244
R5246 gnd.n7214 gnd.n167 240.244
R5247 gnd.n7210 gnd.n167 240.244
R5248 gnd.n7210 gnd.n173 240.244
R5249 gnd.n7202 gnd.n173 240.244
R5250 gnd.n7202 gnd.n186 240.244
R5251 gnd.n7198 gnd.n186 240.244
R5252 gnd.n7198 gnd.n192 240.244
R5253 gnd.n7190 gnd.n192 240.244
R5254 gnd.n7190 gnd.n205 240.244
R5255 gnd.n6024 gnd.n977 240.244
R5256 gnd.n6021 gnd.n1018 240.244
R5257 gnd.n6017 gnd.n6016 240.244
R5258 gnd.n6013 gnd.n6012 240.244
R5259 gnd.n6009 gnd.n6008 240.244
R5260 gnd.n6005 gnd.n6004 240.244
R5261 gnd.n6001 gnd.n6000 240.244
R5262 gnd.n5997 gnd.n5996 240.244
R5263 gnd.n5993 gnd.n5992 240.244
R5264 gnd.n5988 gnd.n5987 240.244
R5265 gnd.n5984 gnd.n5983 240.244
R5266 gnd.n5980 gnd.n5979 240.244
R5267 gnd.n5976 gnd.n5975 240.244
R5268 gnd.n4504 gnd.n4503 240.244
R5269 gnd.n4507 gnd.n4506 240.244
R5270 gnd.n4514 gnd.n4513 240.244
R5271 gnd.n4517 gnd.n4516 240.244
R5272 gnd.n4522 gnd.n4497 240.244
R5273 gnd.n4526 gnd.n4525 240.244
R5274 gnd.n4533 gnd.n4532 240.244
R5275 gnd.n4536 gnd.n4535 240.244
R5276 gnd.n4543 gnd.n4542 240.244
R5277 gnd.n4546 gnd.n4545 240.244
R5278 gnd.n4553 gnd.n4552 240.244
R5279 gnd.n4556 gnd.n4555 240.244
R5280 gnd.n4563 gnd.n4562 240.244
R5281 gnd.n4566 gnd.n4565 240.244
R5282 gnd.n4571 gnd.n4484 240.244
R5283 gnd.n4039 gnd.n2235 240.244
R5284 gnd.n2235 gnd.n2225 240.244
R5285 gnd.n4058 gnd.n2225 240.244
R5286 gnd.n4059 gnd.n4058 240.244
R5287 gnd.n4059 gnd.n2216 240.244
R5288 gnd.n2216 gnd.n2207 240.244
R5289 gnd.n4078 gnd.n2207 240.244
R5290 gnd.n4079 gnd.n4078 240.244
R5291 gnd.n4079 gnd.n2199 240.244
R5292 gnd.n2199 gnd.n2189 240.244
R5293 gnd.n4098 gnd.n2189 240.244
R5294 gnd.n4099 gnd.n4098 240.244
R5295 gnd.n4099 gnd.n2179 240.244
R5296 gnd.n4102 gnd.n2179 240.244
R5297 gnd.n4102 gnd.n2170 240.244
R5298 gnd.n2170 gnd.n2163 240.244
R5299 gnd.n4134 gnd.n2163 240.244
R5300 gnd.n4134 gnd.n2153 240.244
R5301 gnd.n4137 gnd.n2153 240.244
R5302 gnd.n4137 gnd.n2145 240.244
R5303 gnd.n2145 gnd.n2138 240.244
R5304 gnd.n4169 gnd.n2138 240.244
R5305 gnd.n4169 gnd.n2129 240.244
R5306 gnd.n4172 gnd.n2129 240.244
R5307 gnd.n4172 gnd.n2121 240.244
R5308 gnd.n2121 gnd.n2112 240.244
R5309 gnd.n4216 gnd.n2112 240.244
R5310 gnd.n4216 gnd.n2104 240.244
R5311 gnd.n2104 gnd.n2095 240.244
R5312 gnd.n4235 gnd.n2095 240.244
R5313 gnd.n4236 gnd.n4235 240.244
R5314 gnd.n4236 gnd.n2084 240.244
R5315 gnd.n4239 gnd.n2084 240.244
R5316 gnd.n4239 gnd.n2076 240.244
R5317 gnd.n4242 gnd.n2076 240.244
R5318 gnd.n4242 gnd.n884 240.244
R5319 gnd.n4272 gnd.n884 240.244
R5320 gnd.n4272 gnd.n897 240.244
R5321 gnd.n2066 gnd.n897 240.244
R5322 gnd.n2066 gnd.n908 240.244
R5323 gnd.n4281 gnd.n908 240.244
R5324 gnd.n4281 gnd.n919 240.244
R5325 gnd.n2060 gnd.n919 240.244
R5326 gnd.n2060 gnd.n928 240.244
R5327 gnd.n4325 gnd.n928 240.244
R5328 gnd.n4325 gnd.n939 240.244
R5329 gnd.n2049 gnd.n939 240.244
R5330 gnd.n2049 gnd.n948 240.244
R5331 gnd.n4332 gnd.n948 240.244
R5332 gnd.n4332 gnd.n959 240.244
R5333 gnd.n4582 gnd.n959 240.244
R5334 gnd.n4582 gnd.n969 240.244
R5335 gnd.n2038 gnd.n969 240.244
R5336 gnd.n3761 gnd.n3760 240.244
R5337 gnd.n4029 gnd.n3760 240.244
R5338 gnd.n4027 gnd.n4026 240.244
R5339 gnd.n4023 gnd.n4022 240.244
R5340 gnd.n4019 gnd.n4018 240.244
R5341 gnd.n4015 gnd.n4014 240.244
R5342 gnd.n4011 gnd.n4010 240.244
R5343 gnd.n4007 gnd.n4006 240.244
R5344 gnd.n4003 gnd.n4002 240.244
R5345 gnd.n3998 gnd.n3997 240.244
R5346 gnd.n3994 gnd.n3993 240.244
R5347 gnd.n3990 gnd.n3989 240.244
R5348 gnd.n3986 gnd.n3985 240.244
R5349 gnd.n3982 gnd.n3981 240.244
R5350 gnd.n3978 gnd.n3977 240.244
R5351 gnd.n3974 gnd.n3973 240.244
R5352 gnd.n3970 gnd.n3969 240.244
R5353 gnd.n3966 gnd.n3965 240.244
R5354 gnd.n3962 gnd.n3961 240.244
R5355 gnd.n3958 gnd.n3957 240.244
R5356 gnd.n3954 gnd.n3953 240.244
R5357 gnd.n3950 gnd.n3949 240.244
R5358 gnd.n3946 gnd.n3945 240.244
R5359 gnd.n3942 gnd.n3941 240.244
R5360 gnd.n3938 gnd.n3937 240.244
R5361 gnd.n3934 gnd.n3933 240.244
R5362 gnd.n3930 gnd.n3929 240.244
R5363 gnd.n3926 gnd.n3925 240.244
R5364 gnd.n3922 gnd.n2243 240.244
R5365 gnd.n4050 gnd.n2233 240.244
R5366 gnd.n4050 gnd.n2229 240.244
R5367 gnd.n4056 gnd.n2229 240.244
R5368 gnd.n4056 gnd.n2214 240.244
R5369 gnd.n4070 gnd.n2214 240.244
R5370 gnd.n4070 gnd.n2210 240.244
R5371 gnd.n4076 gnd.n2210 240.244
R5372 gnd.n4076 gnd.n2197 240.244
R5373 gnd.n4090 gnd.n2197 240.244
R5374 gnd.n4090 gnd.n2193 240.244
R5375 gnd.n4096 gnd.n2193 240.244
R5376 gnd.n4096 gnd.n2177 240.244
R5377 gnd.n4114 gnd.n2177 240.244
R5378 gnd.n4114 gnd.n2172 240.244
R5379 gnd.n4122 gnd.n2172 240.244
R5380 gnd.n4122 gnd.n2173 240.244
R5381 gnd.n2173 gnd.n2152 240.244
R5382 gnd.n4149 gnd.n2152 240.244
R5383 gnd.n4149 gnd.n2147 240.244
R5384 gnd.n4157 gnd.n2147 240.244
R5385 gnd.n4157 gnd.n2148 240.244
R5386 gnd.n2148 gnd.n2128 240.244
R5387 gnd.n4184 gnd.n2128 240.244
R5388 gnd.n4184 gnd.n2123 240.244
R5389 gnd.n4192 gnd.n2123 240.244
R5390 gnd.n4192 gnd.n2124 240.244
R5391 gnd.n2124 gnd.n2103 240.244
R5392 gnd.n4227 gnd.n2103 240.244
R5393 gnd.n4227 gnd.n2099 240.244
R5394 gnd.n4233 gnd.n2099 240.244
R5395 gnd.n4233 gnd.n2082 240.244
R5396 gnd.n4254 gnd.n2082 240.244
R5397 gnd.n4254 gnd.n2078 240.244
R5398 gnd.n4261 gnd.n2078 240.244
R5399 gnd.n4261 gnd.n888 240.244
R5400 gnd.n6078 gnd.n888 240.244
R5401 gnd.n6078 gnd.n889 240.244
R5402 gnd.n6074 gnd.n889 240.244
R5403 gnd.n6074 gnd.n895 240.244
R5404 gnd.n6066 gnd.n895 240.244
R5405 gnd.n6066 gnd.n911 240.244
R5406 gnd.n6062 gnd.n911 240.244
R5407 gnd.n6062 gnd.n917 240.244
R5408 gnd.n6054 gnd.n917 240.244
R5409 gnd.n6054 gnd.n931 240.244
R5410 gnd.n6050 gnd.n931 240.244
R5411 gnd.n6050 gnd.n937 240.244
R5412 gnd.n6042 gnd.n937 240.244
R5413 gnd.n6042 gnd.n951 240.244
R5414 gnd.n6038 gnd.n951 240.244
R5415 gnd.n6038 gnd.n957 240.244
R5416 gnd.n6030 gnd.n957 240.244
R5417 gnd.n6030 gnd.n972 240.244
R5418 gnd.n3721 gnd.n2268 240.244
R5419 gnd.n3714 gnd.n3713 240.244
R5420 gnd.n3711 gnd.n3710 240.244
R5421 gnd.n3707 gnd.n3706 240.244
R5422 gnd.n3703 gnd.n3702 240.244
R5423 gnd.n3699 gnd.n3698 240.244
R5424 gnd.n3695 gnd.n3694 240.244
R5425 gnd.n3691 gnd.n3690 240.244
R5426 gnd.n2965 gnd.n2677 240.244
R5427 gnd.n2975 gnd.n2677 240.244
R5428 gnd.n2975 gnd.n2668 240.244
R5429 gnd.n2668 gnd.n2657 240.244
R5430 gnd.n2996 gnd.n2657 240.244
R5431 gnd.n2996 gnd.n2651 240.244
R5432 gnd.n3006 gnd.n2651 240.244
R5433 gnd.n3006 gnd.n2640 240.244
R5434 gnd.n2640 gnd.n2632 240.244
R5435 gnd.n3024 gnd.n2632 240.244
R5436 gnd.n3025 gnd.n3024 240.244
R5437 gnd.n3025 gnd.n2617 240.244
R5438 gnd.n3027 gnd.n2617 240.244
R5439 gnd.n3027 gnd.n2603 240.244
R5440 gnd.n3069 gnd.n2603 240.244
R5441 gnd.n3070 gnd.n3069 240.244
R5442 gnd.n3073 gnd.n3070 240.244
R5443 gnd.n3073 gnd.n2558 240.244
R5444 gnd.n2598 gnd.n2558 240.244
R5445 gnd.n2598 gnd.n2568 240.244
R5446 gnd.n3083 gnd.n2568 240.244
R5447 gnd.n3083 gnd.n2589 240.244
R5448 gnd.n3093 gnd.n2589 240.244
R5449 gnd.n3093 gnd.n2471 240.244
R5450 gnd.n3138 gnd.n2471 240.244
R5451 gnd.n3138 gnd.n2457 240.244
R5452 gnd.n3160 gnd.n2457 240.244
R5453 gnd.n3161 gnd.n3160 240.244
R5454 gnd.n3161 gnd.n2444 240.244
R5455 gnd.n2444 gnd.n2433 240.244
R5456 gnd.n3192 gnd.n2433 240.244
R5457 gnd.n3193 gnd.n3192 240.244
R5458 gnd.n3194 gnd.n3193 240.244
R5459 gnd.n3194 gnd.n2418 240.244
R5460 gnd.n2418 gnd.n2417 240.244
R5461 gnd.n2417 gnd.n2402 240.244
R5462 gnd.n3245 gnd.n2402 240.244
R5463 gnd.n3246 gnd.n3245 240.244
R5464 gnd.n3246 gnd.n2389 240.244
R5465 gnd.n2389 gnd.n2378 240.244
R5466 gnd.n3277 gnd.n2378 240.244
R5467 gnd.n3278 gnd.n3277 240.244
R5468 gnd.n3279 gnd.n3278 240.244
R5469 gnd.n3279 gnd.n2362 240.244
R5470 gnd.n2362 gnd.n2361 240.244
R5471 gnd.n2361 gnd.n2348 240.244
R5472 gnd.n3334 gnd.n2348 240.244
R5473 gnd.n3335 gnd.n3334 240.244
R5474 gnd.n3335 gnd.n2335 240.244
R5475 gnd.n2335 gnd.n2325 240.244
R5476 gnd.n3622 gnd.n2325 240.244
R5477 gnd.n3625 gnd.n3622 240.244
R5478 gnd.n3625 gnd.n3624 240.244
R5479 gnd.n2955 gnd.n2690 240.244
R5480 gnd.n2711 gnd.n2690 240.244
R5481 gnd.n2714 gnd.n2713 240.244
R5482 gnd.n2721 gnd.n2720 240.244
R5483 gnd.n2724 gnd.n2723 240.244
R5484 gnd.n2731 gnd.n2730 240.244
R5485 gnd.n2734 gnd.n2733 240.244
R5486 gnd.n2741 gnd.n2740 240.244
R5487 gnd.n2963 gnd.n2687 240.244
R5488 gnd.n2687 gnd.n2666 240.244
R5489 gnd.n2986 gnd.n2666 240.244
R5490 gnd.n2986 gnd.n2660 240.244
R5491 gnd.n2994 gnd.n2660 240.244
R5492 gnd.n2994 gnd.n2662 240.244
R5493 gnd.n2662 gnd.n2638 240.244
R5494 gnd.n3016 gnd.n2638 240.244
R5495 gnd.n3016 gnd.n2634 240.244
R5496 gnd.n3022 gnd.n2634 240.244
R5497 gnd.n3022 gnd.n2616 240.244
R5498 gnd.n3047 gnd.n2616 240.244
R5499 gnd.n3047 gnd.n2611 240.244
R5500 gnd.n3059 gnd.n2611 240.244
R5501 gnd.n3059 gnd.n2612 240.244
R5502 gnd.n3055 gnd.n2612 240.244
R5503 gnd.n3055 gnd.n2560 240.244
R5504 gnd.n3107 gnd.n2560 240.244
R5505 gnd.n3107 gnd.n2561 240.244
R5506 gnd.n3103 gnd.n2561 240.244
R5507 gnd.n3103 gnd.n2567 240.244
R5508 gnd.n2587 gnd.n2567 240.244
R5509 gnd.n2587 gnd.n2469 240.244
R5510 gnd.n3142 gnd.n2469 240.244
R5511 gnd.n3142 gnd.n2464 240.244
R5512 gnd.n3150 gnd.n2464 240.244
R5513 gnd.n3150 gnd.n2465 240.244
R5514 gnd.n2465 gnd.n2442 240.244
R5515 gnd.n3182 gnd.n2442 240.244
R5516 gnd.n3182 gnd.n2437 240.244
R5517 gnd.n3190 gnd.n2437 240.244
R5518 gnd.n3190 gnd.n2438 240.244
R5519 gnd.n2438 gnd.n2415 240.244
R5520 gnd.n3227 gnd.n2415 240.244
R5521 gnd.n3227 gnd.n2410 240.244
R5522 gnd.n3235 gnd.n2410 240.244
R5523 gnd.n3235 gnd.n2411 240.244
R5524 gnd.n2411 gnd.n2387 240.244
R5525 gnd.n3267 gnd.n2387 240.244
R5526 gnd.n3267 gnd.n2382 240.244
R5527 gnd.n3275 gnd.n2382 240.244
R5528 gnd.n3275 gnd.n2383 240.244
R5529 gnd.n2383 gnd.n2360 240.244
R5530 gnd.n3316 gnd.n2360 240.244
R5531 gnd.n3316 gnd.n2355 240.244
R5532 gnd.n3324 gnd.n2355 240.244
R5533 gnd.n3324 gnd.n2356 240.244
R5534 gnd.n2356 gnd.n2333 240.244
R5535 gnd.n3610 gnd.n2333 240.244
R5536 gnd.n3610 gnd.n2328 240.244
R5537 gnd.n3620 gnd.n2328 240.244
R5538 gnd.n3620 gnd.n2329 240.244
R5539 gnd.n2329 gnd.n2267 240.244
R5540 gnd.n6978 gnd.n211 240.244
R5541 gnd.n6984 gnd.n6983 240.244
R5542 gnd.n6987 gnd.n6986 240.244
R5543 gnd.n6994 gnd.n6993 240.244
R5544 gnd.n6997 gnd.n6996 240.244
R5545 gnd.n7004 gnd.n7003 240.244
R5546 gnd.n7007 gnd.n7006 240.244
R5547 gnd.n7014 gnd.n7013 240.244
R5548 gnd.n7017 gnd.n7016 240.244
R5549 gnd.n5524 gnd.n1399 240.244
R5550 gnd.n5524 gnd.n1409 240.244
R5551 gnd.n5469 gnd.n1409 240.244
R5552 gnd.n5469 gnd.n1424 240.244
R5553 gnd.n5470 gnd.n1424 240.244
R5554 gnd.n5470 gnd.n1434 240.244
R5555 gnd.n5473 gnd.n1434 240.244
R5556 gnd.n5473 gnd.n1445 240.244
R5557 gnd.n5474 gnd.n1445 240.244
R5558 gnd.n5474 gnd.n1455 240.244
R5559 gnd.n1458 gnd.n1455 240.244
R5560 gnd.n5503 gnd.n1458 240.244
R5561 gnd.n5503 gnd.n381 240.244
R5562 gnd.n381 gnd.n369 240.244
R5563 gnd.n6818 gnd.n369 240.244
R5564 gnd.n6818 gnd.n364 240.244
R5565 gnd.n6825 gnd.n364 240.244
R5566 gnd.n6825 gnd.n353 240.244
R5567 gnd.n353 gnd.n342 240.244
R5568 gnd.n6852 gnd.n342 240.244
R5569 gnd.n6852 gnd.n337 240.244
R5570 gnd.n6864 gnd.n337 240.244
R5571 gnd.n6864 gnd.n330 240.244
R5572 gnd.n6857 gnd.n330 240.244
R5573 gnd.n6857 gnd.n322 240.244
R5574 gnd.n322 gnd.n321 240.244
R5575 gnd.n321 gnd.n82 240.244
R5576 gnd.n7264 gnd.n82 240.244
R5577 gnd.n7264 gnd.n84 240.244
R5578 gnd.n97 gnd.n84 240.244
R5579 gnd.n6933 gnd.n97 240.244
R5580 gnd.n6933 gnd.n108 240.244
R5581 gnd.n6936 gnd.n108 240.244
R5582 gnd.n6936 gnd.n118 240.244
R5583 gnd.n6941 gnd.n118 240.244
R5584 gnd.n6941 gnd.n127 240.244
R5585 gnd.n6944 gnd.n127 240.244
R5586 gnd.n6944 gnd.n137 240.244
R5587 gnd.n6949 gnd.n137 240.244
R5588 gnd.n6949 gnd.n146 240.244
R5589 gnd.n6952 gnd.n146 240.244
R5590 gnd.n6952 gnd.n156 240.244
R5591 gnd.n7040 gnd.n156 240.244
R5592 gnd.n7040 gnd.n165 240.244
R5593 gnd.n7036 gnd.n165 240.244
R5594 gnd.n7036 gnd.n175 240.244
R5595 gnd.n7033 gnd.n175 240.244
R5596 gnd.n7033 gnd.n184 240.244
R5597 gnd.n7030 gnd.n184 240.244
R5598 gnd.n7030 gnd.n194 240.244
R5599 gnd.n7027 gnd.n194 240.244
R5600 gnd.n7027 gnd.n203 240.244
R5601 gnd.n7024 gnd.n203 240.244
R5602 gnd.n1243 gnd.n1242 240.244
R5603 gnd.n1318 gnd.n1250 240.244
R5604 gnd.n1321 gnd.n1251 240.244
R5605 gnd.n1259 gnd.n1258 240.244
R5606 gnd.n1323 gnd.n1266 240.244
R5607 gnd.n1326 gnd.n1267 240.244
R5608 gnd.n1275 gnd.n1274 240.244
R5609 gnd.n1328 gnd.n1284 240.244
R5610 gnd.n5715 gnd.n1287 240.244
R5611 gnd.n5591 gnd.n1402 240.244
R5612 gnd.n5587 gnd.n1402 240.244
R5613 gnd.n5587 gnd.n1407 240.244
R5614 gnd.n5579 gnd.n1407 240.244
R5615 gnd.n5579 gnd.n1426 240.244
R5616 gnd.n5575 gnd.n1426 240.244
R5617 gnd.n5575 gnd.n1431 240.244
R5618 gnd.n5567 gnd.n1431 240.244
R5619 gnd.n5567 gnd.n1447 240.244
R5620 gnd.n5563 gnd.n1447 240.244
R5621 gnd.n5563 gnd.n1452 240.244
R5622 gnd.n1452 gnd.n383 240.244
R5623 gnd.n6806 gnd.n383 240.244
R5624 gnd.n6806 gnd.n384 240.244
R5625 gnd.n384 gnd.n372 240.244
R5626 gnd.n6801 gnd.n372 240.244
R5627 gnd.n6801 gnd.n355 240.244
R5628 gnd.n6840 gnd.n355 240.244
R5629 gnd.n6840 gnd.n356 240.244
R5630 gnd.n356 gnd.n344 240.244
R5631 gnd.n6835 gnd.n344 240.244
R5632 gnd.n6835 gnd.n331 240.244
R5633 gnd.n6873 gnd.n331 240.244
R5634 gnd.n6873 gnd.n318 240.244
R5635 gnd.n6886 gnd.n318 240.244
R5636 gnd.n6886 gnd.n312 240.244
R5637 gnd.n6894 gnd.n312 240.244
R5638 gnd.n6894 gnd.n87 240.244
R5639 gnd.n98 gnd.n87 240.244
R5640 gnd.n7256 gnd.n98 240.244
R5641 gnd.n7256 gnd.n99 240.244
R5642 gnd.n7252 gnd.n99 240.244
R5643 gnd.n7252 gnd.n105 240.244
R5644 gnd.n7244 gnd.n105 240.244
R5645 gnd.n7244 gnd.n120 240.244
R5646 gnd.n7240 gnd.n120 240.244
R5647 gnd.n7240 gnd.n125 240.244
R5648 gnd.n7232 gnd.n125 240.244
R5649 gnd.n7232 gnd.n138 240.244
R5650 gnd.n7228 gnd.n138 240.244
R5651 gnd.n7228 gnd.n143 240.244
R5652 gnd.n7220 gnd.n143 240.244
R5653 gnd.n7220 gnd.n158 240.244
R5654 gnd.n7216 gnd.n158 240.244
R5655 gnd.n7216 gnd.n163 240.244
R5656 gnd.n7208 gnd.n163 240.244
R5657 gnd.n7208 gnd.n176 240.244
R5658 gnd.n7204 gnd.n176 240.244
R5659 gnd.n7204 gnd.n181 240.244
R5660 gnd.n7196 gnd.n181 240.244
R5661 gnd.n7196 gnd.n196 240.244
R5662 gnd.n7192 gnd.n196 240.244
R5663 gnd.n7192 gnd.n201 240.244
R5664 gnd.n2287 gnd.n2245 240.244
R5665 gnd.n3681 gnd.n3680 240.244
R5666 gnd.n3677 gnd.n3676 240.244
R5667 gnd.n3673 gnd.n3672 240.244
R5668 gnd.n3669 gnd.n3668 240.244
R5669 gnd.n3665 gnd.n3664 240.244
R5670 gnd.n3661 gnd.n3660 240.244
R5671 gnd.n3657 gnd.n3656 240.244
R5672 gnd.n3653 gnd.n3652 240.244
R5673 gnd.n3649 gnd.n3648 240.244
R5674 gnd.n3645 gnd.n3644 240.244
R5675 gnd.n3641 gnd.n3640 240.244
R5676 gnd.n3637 gnd.n3636 240.244
R5677 gnd.n2878 gnd.n2775 240.244
R5678 gnd.n2878 gnd.n2768 240.244
R5679 gnd.n2889 gnd.n2768 240.244
R5680 gnd.n2889 gnd.n2764 240.244
R5681 gnd.n2895 gnd.n2764 240.244
R5682 gnd.n2895 gnd.n2756 240.244
R5683 gnd.n2905 gnd.n2756 240.244
R5684 gnd.n2905 gnd.n2751 240.244
R5685 gnd.n2941 gnd.n2751 240.244
R5686 gnd.n2941 gnd.n2752 240.244
R5687 gnd.n2752 gnd.n2699 240.244
R5688 gnd.n2936 gnd.n2699 240.244
R5689 gnd.n2936 gnd.n2935 240.244
R5690 gnd.n2935 gnd.n2678 240.244
R5691 gnd.n2931 gnd.n2678 240.244
R5692 gnd.n2931 gnd.n2669 240.244
R5693 gnd.n2928 gnd.n2669 240.244
R5694 gnd.n2928 gnd.n2927 240.244
R5695 gnd.n2927 gnd.n2652 240.244
R5696 gnd.n2923 gnd.n2652 240.244
R5697 gnd.n2923 gnd.n2641 240.244
R5698 gnd.n2641 gnd.n2622 240.244
R5699 gnd.n3036 gnd.n2622 240.244
R5700 gnd.n3036 gnd.n2618 240.244
R5701 gnd.n3044 gnd.n2618 240.244
R5702 gnd.n3044 gnd.n2609 240.244
R5703 gnd.n2609 gnd.n2545 240.244
R5704 gnd.n3116 gnd.n2545 240.244
R5705 gnd.n3116 gnd.n2546 240.244
R5706 gnd.n2557 gnd.n2546 240.244
R5707 gnd.n2592 gnd.n2557 240.244
R5708 gnd.n2595 gnd.n2592 240.244
R5709 gnd.n2595 gnd.n2569 240.244
R5710 gnd.n2582 gnd.n2569 240.244
R5711 gnd.n2582 gnd.n2579 240.244
R5712 gnd.n2579 gnd.n2472 240.244
R5713 gnd.n3137 gnd.n2472 240.244
R5714 gnd.n3137 gnd.n2462 240.244
R5715 gnd.n3133 gnd.n2462 240.244
R5716 gnd.n3133 gnd.n2456 240.244
R5717 gnd.n3130 gnd.n2456 240.244
R5718 gnd.n3130 gnd.n2445 240.244
R5719 gnd.n3127 gnd.n2445 240.244
R5720 gnd.n3127 gnd.n2423 240.244
R5721 gnd.n3203 gnd.n2423 240.244
R5722 gnd.n3203 gnd.n2419 240.244
R5723 gnd.n3224 gnd.n2419 240.244
R5724 gnd.n3224 gnd.n2408 240.244
R5725 gnd.n3220 gnd.n2408 240.244
R5726 gnd.n3220 gnd.n2401 240.244
R5727 gnd.n3217 gnd.n2401 240.244
R5728 gnd.n3217 gnd.n2390 240.244
R5729 gnd.n3214 gnd.n2390 240.244
R5730 gnd.n3214 gnd.n2367 240.244
R5731 gnd.n3288 gnd.n2367 240.244
R5732 gnd.n3288 gnd.n2363 240.244
R5733 gnd.n3313 gnd.n2363 240.244
R5734 gnd.n3313 gnd.n2354 240.244
R5735 gnd.n3309 gnd.n2354 240.244
R5736 gnd.n3309 gnd.n2347 240.244
R5737 gnd.n3305 gnd.n2347 240.244
R5738 gnd.n3305 gnd.n2336 240.244
R5739 gnd.n3302 gnd.n2336 240.244
R5740 gnd.n3302 gnd.n2316 240.244
R5741 gnd.n3632 gnd.n2316 240.244
R5742 gnd.n2792 gnd.n2791 240.244
R5743 gnd.n2863 gnd.n2791 240.244
R5744 gnd.n2861 gnd.n2860 240.244
R5745 gnd.n2857 gnd.n2856 240.244
R5746 gnd.n2853 gnd.n2852 240.244
R5747 gnd.n2849 gnd.n2848 240.244
R5748 gnd.n2845 gnd.n2844 240.244
R5749 gnd.n2841 gnd.n2840 240.244
R5750 gnd.n2837 gnd.n2836 240.244
R5751 gnd.n2833 gnd.n2832 240.244
R5752 gnd.n2829 gnd.n2828 240.244
R5753 gnd.n2825 gnd.n2824 240.244
R5754 gnd.n2821 gnd.n2779 240.244
R5755 gnd.n2881 gnd.n2773 240.244
R5756 gnd.n2881 gnd.n2769 240.244
R5757 gnd.n2887 gnd.n2769 240.244
R5758 gnd.n2887 gnd.n2762 240.244
R5759 gnd.n2897 gnd.n2762 240.244
R5760 gnd.n2897 gnd.n2758 240.244
R5761 gnd.n2903 gnd.n2758 240.244
R5762 gnd.n2903 gnd.n2749 240.244
R5763 gnd.n2943 gnd.n2749 240.244
R5764 gnd.n2943 gnd.n2700 240.244
R5765 gnd.n2951 gnd.n2700 240.244
R5766 gnd.n2951 gnd.n2701 240.244
R5767 gnd.n2701 gnd.n2679 240.244
R5768 gnd.n2972 gnd.n2679 240.244
R5769 gnd.n2972 gnd.n2671 240.244
R5770 gnd.n2983 gnd.n2671 240.244
R5771 gnd.n2983 gnd.n2672 240.244
R5772 gnd.n2672 gnd.n2653 240.244
R5773 gnd.n3003 gnd.n2653 240.244
R5774 gnd.n3003 gnd.n2643 240.244
R5775 gnd.n3013 gnd.n2643 240.244
R5776 gnd.n3013 gnd.n2624 240.244
R5777 gnd.n3034 gnd.n2624 240.244
R5778 gnd.n3034 gnd.n2626 240.244
R5779 gnd.n2626 gnd.n2607 240.244
R5780 gnd.n3062 gnd.n2607 240.244
R5781 gnd.n3062 gnd.n2549 240.244
R5782 gnd.n3114 gnd.n2549 240.244
R5783 gnd.n3114 gnd.n2550 240.244
R5784 gnd.n3110 gnd.n2550 240.244
R5785 gnd.n3110 gnd.n2556 240.244
R5786 gnd.n2571 gnd.n2556 240.244
R5787 gnd.n3100 gnd.n2571 240.244
R5788 gnd.n3100 gnd.n2572 240.244
R5789 gnd.n3096 gnd.n2572 240.244
R5790 gnd.n3096 gnd.n2578 240.244
R5791 gnd.n2578 gnd.n2461 240.244
R5792 gnd.n3153 gnd.n2461 240.244
R5793 gnd.n3153 gnd.n2454 240.244
R5794 gnd.n3164 gnd.n2454 240.244
R5795 gnd.n3164 gnd.n2447 240.244
R5796 gnd.n3179 gnd.n2447 240.244
R5797 gnd.n3179 gnd.n2448 240.244
R5798 gnd.n2448 gnd.n2426 240.244
R5799 gnd.n3201 gnd.n2426 240.244
R5800 gnd.n3201 gnd.n2427 240.244
R5801 gnd.n2427 gnd.n2406 240.244
R5802 gnd.n3238 gnd.n2406 240.244
R5803 gnd.n3238 gnd.n2399 240.244
R5804 gnd.n3249 gnd.n2399 240.244
R5805 gnd.n3249 gnd.n2392 240.244
R5806 gnd.n3264 gnd.n2392 240.244
R5807 gnd.n3264 gnd.n2393 240.244
R5808 gnd.n2393 gnd.n2370 240.244
R5809 gnd.n3286 gnd.n2370 240.244
R5810 gnd.n3286 gnd.n2372 240.244
R5811 gnd.n2372 gnd.n2352 240.244
R5812 gnd.n3327 gnd.n2352 240.244
R5813 gnd.n3327 gnd.n2345 240.244
R5814 gnd.n3338 gnd.n2345 240.244
R5815 gnd.n3338 gnd.n2338 240.244
R5816 gnd.n3607 gnd.n2338 240.244
R5817 gnd.n3607 gnd.n2339 240.244
R5818 gnd.n2339 gnd.n2320 240.244
R5819 gnd.n3630 gnd.n2320 240.244
R5820 gnd.n4369 gnd.n979 240.244
R5821 gnd.n4379 gnd.n4378 240.244
R5822 gnd.n4381 gnd.n4380 240.244
R5823 gnd.n4389 gnd.n4388 240.244
R5824 gnd.n4399 gnd.n4398 240.244
R5825 gnd.n4401 gnd.n4400 240.244
R5826 gnd.n4409 gnd.n4408 240.244
R5827 gnd.n4419 gnd.n4418 240.244
R5828 gnd.n4421 gnd.n4420 240.244
R5829 gnd.n3876 gnd.n2236 240.244
R5830 gnd.n3873 gnd.n2236 240.244
R5831 gnd.n3873 gnd.n2227 240.244
R5832 gnd.n3870 gnd.n2227 240.244
R5833 gnd.n3870 gnd.n2217 240.244
R5834 gnd.n3867 gnd.n2217 240.244
R5835 gnd.n3867 gnd.n2208 240.244
R5836 gnd.n3864 gnd.n2208 240.244
R5837 gnd.n3864 gnd.n2200 240.244
R5838 gnd.n3861 gnd.n2200 240.244
R5839 gnd.n3861 gnd.n2191 240.244
R5840 gnd.n3858 gnd.n2191 240.244
R5841 gnd.n3858 gnd.n2180 240.244
R5842 gnd.n2180 gnd.n2169 240.244
R5843 gnd.n4124 gnd.n2169 240.244
R5844 gnd.n4124 gnd.n2165 240.244
R5845 gnd.n4132 gnd.n2165 240.244
R5846 gnd.n4132 gnd.n2154 240.244
R5847 gnd.n2154 gnd.n2144 240.244
R5848 gnd.n4159 gnd.n2144 240.244
R5849 gnd.n4159 gnd.n2140 240.244
R5850 gnd.n4167 gnd.n2140 240.244
R5851 gnd.n4167 gnd.n2130 240.244
R5852 gnd.n2130 gnd.n2119 240.244
R5853 gnd.n4194 gnd.n2119 240.244
R5854 gnd.n4194 gnd.n2114 240.244
R5855 gnd.n4214 gnd.n2114 240.244
R5856 gnd.n4214 gnd.n2105 240.244
R5857 gnd.n4200 gnd.n2105 240.244
R5858 gnd.n4200 gnd.n2097 240.244
R5859 gnd.n4201 gnd.n2097 240.244
R5860 gnd.n4201 gnd.n2085 240.244
R5861 gnd.n2085 gnd.n2075 240.244
R5862 gnd.n4263 gnd.n2075 240.244
R5863 gnd.n4264 gnd.n4263 240.244
R5864 gnd.n4264 gnd.n885 240.244
R5865 gnd.n4270 gnd.n885 240.244
R5866 gnd.n4270 gnd.n898 240.244
R5867 gnd.n4289 gnd.n898 240.244
R5868 gnd.n4289 gnd.n909 240.244
R5869 gnd.n4283 gnd.n909 240.244
R5870 gnd.n4283 gnd.n920 240.244
R5871 gnd.n4317 gnd.n920 240.244
R5872 gnd.n4317 gnd.n929 240.244
R5873 gnd.n4323 gnd.n929 240.244
R5874 gnd.n4323 gnd.n940 240.244
R5875 gnd.n4595 gnd.n940 240.244
R5876 gnd.n4595 gnd.n949 240.244
R5877 gnd.n2054 gnd.n949 240.244
R5878 gnd.n2054 gnd.n960 240.244
R5879 gnd.n4584 gnd.n960 240.244
R5880 gnd.n4584 gnd.n970 240.244
R5881 gnd.n4624 gnd.n970 240.244
R5882 gnd.n3913 gnd.n3912 240.244
R5883 gnd.n3909 gnd.n3908 240.244
R5884 gnd.n3905 gnd.n3904 240.244
R5885 gnd.n3901 gnd.n3900 240.244
R5886 gnd.n3897 gnd.n3896 240.244
R5887 gnd.n3893 gnd.n3892 240.244
R5888 gnd.n3889 gnd.n3888 240.244
R5889 gnd.n3885 gnd.n3884 240.244
R5890 gnd.n3840 gnd.n3759 240.244
R5891 gnd.n4048 gnd.n2237 240.244
R5892 gnd.n4048 gnd.n2238 240.244
R5893 gnd.n2238 gnd.n2228 240.244
R5894 gnd.n2228 gnd.n2219 240.244
R5895 gnd.n4068 gnd.n2219 240.244
R5896 gnd.n4068 gnd.n2220 240.244
R5897 gnd.n2220 gnd.n2209 240.244
R5898 gnd.n2209 gnd.n2201 240.244
R5899 gnd.n4088 gnd.n2201 240.244
R5900 gnd.n4088 gnd.n2202 240.244
R5901 gnd.n2202 gnd.n2192 240.244
R5902 gnd.n2192 gnd.n2182 240.244
R5903 gnd.n4112 gnd.n2182 240.244
R5904 gnd.n4112 gnd.n2183 240.244
R5905 gnd.n2183 gnd.n2171 240.244
R5906 gnd.n4107 gnd.n2171 240.244
R5907 gnd.n4107 gnd.n2156 240.244
R5908 gnd.n4147 gnd.n2156 240.244
R5909 gnd.n4147 gnd.n2157 240.244
R5910 gnd.n2157 gnd.n2146 240.244
R5911 gnd.n4142 gnd.n2146 240.244
R5912 gnd.n4142 gnd.n2131 240.244
R5913 gnd.n4182 gnd.n2131 240.244
R5914 gnd.n4182 gnd.n2132 240.244
R5915 gnd.n2132 gnd.n2122 240.244
R5916 gnd.n4177 gnd.n2122 240.244
R5917 gnd.n4177 gnd.n2106 240.244
R5918 gnd.n4225 gnd.n2106 240.244
R5919 gnd.n4225 gnd.n2107 240.244
R5920 gnd.n2107 gnd.n2098 240.244
R5921 gnd.n2098 gnd.n2087 240.244
R5922 gnd.n4252 gnd.n2087 240.244
R5923 gnd.n4252 gnd.n2088 240.244
R5924 gnd.n2088 gnd.n2077 240.244
R5925 gnd.n4247 gnd.n2077 240.244
R5926 gnd.n4247 gnd.n887 240.244
R5927 gnd.n899 gnd.n887 240.244
R5928 gnd.n6072 gnd.n899 240.244
R5929 gnd.n6072 gnd.n900 240.244
R5930 gnd.n6068 gnd.n900 240.244
R5931 gnd.n6068 gnd.n906 240.244
R5932 gnd.n6060 gnd.n906 240.244
R5933 gnd.n6060 gnd.n922 240.244
R5934 gnd.n6056 gnd.n922 240.244
R5935 gnd.n6056 gnd.n927 240.244
R5936 gnd.n6048 gnd.n927 240.244
R5937 gnd.n6048 gnd.n941 240.244
R5938 gnd.n6044 gnd.n941 240.244
R5939 gnd.n6044 gnd.n946 240.244
R5940 gnd.n6036 gnd.n946 240.244
R5941 gnd.n6036 gnd.n962 240.244
R5942 gnd.n6032 gnd.n962 240.244
R5943 gnd.n6032 gnd.n967 240.244
R5944 gnd.n6255 gnd.n712 240.244
R5945 gnd.n6255 gnd.n710 240.244
R5946 gnd.n6259 gnd.n710 240.244
R5947 gnd.n6259 gnd.n706 240.244
R5948 gnd.n6265 gnd.n706 240.244
R5949 gnd.n6265 gnd.n704 240.244
R5950 gnd.n6269 gnd.n704 240.244
R5951 gnd.n6269 gnd.n700 240.244
R5952 gnd.n6275 gnd.n700 240.244
R5953 gnd.n6275 gnd.n698 240.244
R5954 gnd.n6279 gnd.n698 240.244
R5955 gnd.n6279 gnd.n694 240.244
R5956 gnd.n6285 gnd.n694 240.244
R5957 gnd.n6285 gnd.n692 240.244
R5958 gnd.n6289 gnd.n692 240.244
R5959 gnd.n6289 gnd.n688 240.244
R5960 gnd.n6295 gnd.n688 240.244
R5961 gnd.n6295 gnd.n686 240.244
R5962 gnd.n6299 gnd.n686 240.244
R5963 gnd.n6299 gnd.n682 240.244
R5964 gnd.n6305 gnd.n682 240.244
R5965 gnd.n6305 gnd.n680 240.244
R5966 gnd.n6309 gnd.n680 240.244
R5967 gnd.n6309 gnd.n676 240.244
R5968 gnd.n6315 gnd.n676 240.244
R5969 gnd.n6315 gnd.n674 240.244
R5970 gnd.n6319 gnd.n674 240.244
R5971 gnd.n6319 gnd.n670 240.244
R5972 gnd.n6325 gnd.n670 240.244
R5973 gnd.n6325 gnd.n668 240.244
R5974 gnd.n6329 gnd.n668 240.244
R5975 gnd.n6329 gnd.n664 240.244
R5976 gnd.n6335 gnd.n664 240.244
R5977 gnd.n6335 gnd.n662 240.244
R5978 gnd.n6339 gnd.n662 240.244
R5979 gnd.n6339 gnd.n658 240.244
R5980 gnd.n6345 gnd.n658 240.244
R5981 gnd.n6345 gnd.n656 240.244
R5982 gnd.n6349 gnd.n656 240.244
R5983 gnd.n6349 gnd.n652 240.244
R5984 gnd.n6355 gnd.n652 240.244
R5985 gnd.n6355 gnd.n650 240.244
R5986 gnd.n6359 gnd.n650 240.244
R5987 gnd.n6359 gnd.n646 240.244
R5988 gnd.n6365 gnd.n646 240.244
R5989 gnd.n6365 gnd.n644 240.244
R5990 gnd.n6369 gnd.n644 240.244
R5991 gnd.n6369 gnd.n640 240.244
R5992 gnd.n6375 gnd.n640 240.244
R5993 gnd.n6375 gnd.n638 240.244
R5994 gnd.n6379 gnd.n638 240.244
R5995 gnd.n6379 gnd.n634 240.244
R5996 gnd.n6385 gnd.n634 240.244
R5997 gnd.n6385 gnd.n632 240.244
R5998 gnd.n6389 gnd.n632 240.244
R5999 gnd.n6389 gnd.n628 240.244
R6000 gnd.n6395 gnd.n628 240.244
R6001 gnd.n6395 gnd.n626 240.244
R6002 gnd.n6399 gnd.n626 240.244
R6003 gnd.n6399 gnd.n622 240.244
R6004 gnd.n6405 gnd.n622 240.244
R6005 gnd.n6405 gnd.n620 240.244
R6006 gnd.n6409 gnd.n620 240.244
R6007 gnd.n6409 gnd.n616 240.244
R6008 gnd.n6415 gnd.n616 240.244
R6009 gnd.n6415 gnd.n614 240.244
R6010 gnd.n6419 gnd.n614 240.244
R6011 gnd.n6419 gnd.n610 240.244
R6012 gnd.n6425 gnd.n610 240.244
R6013 gnd.n6425 gnd.n608 240.244
R6014 gnd.n6429 gnd.n608 240.244
R6015 gnd.n6429 gnd.n604 240.244
R6016 gnd.n6435 gnd.n604 240.244
R6017 gnd.n6435 gnd.n602 240.244
R6018 gnd.n6439 gnd.n602 240.244
R6019 gnd.n6439 gnd.n598 240.244
R6020 gnd.n6445 gnd.n598 240.244
R6021 gnd.n6445 gnd.n596 240.244
R6022 gnd.n6449 gnd.n596 240.244
R6023 gnd.n6449 gnd.n592 240.244
R6024 gnd.n6455 gnd.n592 240.244
R6025 gnd.n6455 gnd.n590 240.244
R6026 gnd.n6459 gnd.n590 240.244
R6027 gnd.n6459 gnd.n586 240.244
R6028 gnd.n6465 gnd.n586 240.244
R6029 gnd.n6465 gnd.n584 240.244
R6030 gnd.n6469 gnd.n584 240.244
R6031 gnd.n6469 gnd.n580 240.244
R6032 gnd.n6475 gnd.n580 240.244
R6033 gnd.n6475 gnd.n578 240.244
R6034 gnd.n6479 gnd.n578 240.244
R6035 gnd.n6479 gnd.n574 240.244
R6036 gnd.n6485 gnd.n574 240.244
R6037 gnd.n6485 gnd.n572 240.244
R6038 gnd.n6489 gnd.n572 240.244
R6039 gnd.n6489 gnd.n568 240.244
R6040 gnd.n6495 gnd.n568 240.244
R6041 gnd.n6495 gnd.n566 240.244
R6042 gnd.n6499 gnd.n566 240.244
R6043 gnd.n6499 gnd.n562 240.244
R6044 gnd.n6505 gnd.n562 240.244
R6045 gnd.n6505 gnd.n560 240.244
R6046 gnd.n6509 gnd.n560 240.244
R6047 gnd.n6509 gnd.n556 240.244
R6048 gnd.n6515 gnd.n556 240.244
R6049 gnd.n6515 gnd.n554 240.244
R6050 gnd.n6519 gnd.n554 240.244
R6051 gnd.n6519 gnd.n550 240.244
R6052 gnd.n6525 gnd.n550 240.244
R6053 gnd.n6525 gnd.n548 240.244
R6054 gnd.n6529 gnd.n548 240.244
R6055 gnd.n6529 gnd.n544 240.244
R6056 gnd.n6535 gnd.n544 240.244
R6057 gnd.n6535 gnd.n542 240.244
R6058 gnd.n6539 gnd.n542 240.244
R6059 gnd.n6539 gnd.n538 240.244
R6060 gnd.n6545 gnd.n538 240.244
R6061 gnd.n6545 gnd.n536 240.244
R6062 gnd.n6549 gnd.n536 240.244
R6063 gnd.n6549 gnd.n532 240.244
R6064 gnd.n6555 gnd.n532 240.244
R6065 gnd.n6555 gnd.n530 240.244
R6066 gnd.n6559 gnd.n530 240.244
R6067 gnd.n6559 gnd.n526 240.244
R6068 gnd.n6566 gnd.n526 240.244
R6069 gnd.n6566 gnd.n524 240.244
R6070 gnd.n6570 gnd.n524 240.244
R6071 gnd.n6570 gnd.n521 240.244
R6072 gnd.n6576 gnd.n519 240.244
R6073 gnd.n6580 gnd.n519 240.244
R6074 gnd.n6580 gnd.n515 240.244
R6075 gnd.n6586 gnd.n515 240.244
R6076 gnd.n6586 gnd.n513 240.244
R6077 gnd.n6590 gnd.n513 240.244
R6078 gnd.n6590 gnd.n509 240.244
R6079 gnd.n6596 gnd.n509 240.244
R6080 gnd.n6596 gnd.n507 240.244
R6081 gnd.n6600 gnd.n507 240.244
R6082 gnd.n6600 gnd.n503 240.244
R6083 gnd.n6606 gnd.n503 240.244
R6084 gnd.n6606 gnd.n501 240.244
R6085 gnd.n6610 gnd.n501 240.244
R6086 gnd.n6610 gnd.n497 240.244
R6087 gnd.n6616 gnd.n497 240.244
R6088 gnd.n6616 gnd.n495 240.244
R6089 gnd.n6620 gnd.n495 240.244
R6090 gnd.n6620 gnd.n491 240.244
R6091 gnd.n6626 gnd.n491 240.244
R6092 gnd.n6626 gnd.n489 240.244
R6093 gnd.n6630 gnd.n489 240.244
R6094 gnd.n6630 gnd.n485 240.244
R6095 gnd.n6636 gnd.n485 240.244
R6096 gnd.n6636 gnd.n483 240.244
R6097 gnd.n6640 gnd.n483 240.244
R6098 gnd.n6640 gnd.n479 240.244
R6099 gnd.n6646 gnd.n479 240.244
R6100 gnd.n6646 gnd.n477 240.244
R6101 gnd.n6650 gnd.n477 240.244
R6102 gnd.n6650 gnd.n473 240.244
R6103 gnd.n6656 gnd.n473 240.244
R6104 gnd.n6656 gnd.n471 240.244
R6105 gnd.n6660 gnd.n471 240.244
R6106 gnd.n6660 gnd.n467 240.244
R6107 gnd.n6666 gnd.n467 240.244
R6108 gnd.n6666 gnd.n465 240.244
R6109 gnd.n6670 gnd.n465 240.244
R6110 gnd.n6670 gnd.n461 240.244
R6111 gnd.n6676 gnd.n461 240.244
R6112 gnd.n6676 gnd.n459 240.244
R6113 gnd.n6680 gnd.n459 240.244
R6114 gnd.n6680 gnd.n455 240.244
R6115 gnd.n6686 gnd.n455 240.244
R6116 gnd.n6686 gnd.n453 240.244
R6117 gnd.n6690 gnd.n453 240.244
R6118 gnd.n6690 gnd.n449 240.244
R6119 gnd.n6696 gnd.n449 240.244
R6120 gnd.n6696 gnd.n447 240.244
R6121 gnd.n6700 gnd.n447 240.244
R6122 gnd.n6700 gnd.n443 240.244
R6123 gnd.n6706 gnd.n443 240.244
R6124 gnd.n6706 gnd.n441 240.244
R6125 gnd.n6710 gnd.n441 240.244
R6126 gnd.n6710 gnd.n437 240.244
R6127 gnd.n6716 gnd.n437 240.244
R6128 gnd.n6716 gnd.n435 240.244
R6129 gnd.n6720 gnd.n435 240.244
R6130 gnd.n6720 gnd.n431 240.244
R6131 gnd.n6726 gnd.n431 240.244
R6132 gnd.n6726 gnd.n429 240.244
R6133 gnd.n6730 gnd.n429 240.244
R6134 gnd.n6730 gnd.n425 240.244
R6135 gnd.n6736 gnd.n425 240.244
R6136 gnd.n6736 gnd.n423 240.244
R6137 gnd.n6740 gnd.n423 240.244
R6138 gnd.n6740 gnd.n419 240.244
R6139 gnd.n6746 gnd.n419 240.244
R6140 gnd.n6746 gnd.n417 240.244
R6141 gnd.n6750 gnd.n417 240.244
R6142 gnd.n6750 gnd.n413 240.244
R6143 gnd.n6756 gnd.n413 240.244
R6144 gnd.n6756 gnd.n411 240.244
R6145 gnd.n6760 gnd.n411 240.244
R6146 gnd.n6760 gnd.n407 240.244
R6147 gnd.n6766 gnd.n407 240.244
R6148 gnd.n6766 gnd.n405 240.244
R6149 gnd.n6770 gnd.n405 240.244
R6150 gnd.n6770 gnd.n401 240.244
R6151 gnd.n6776 gnd.n401 240.244
R6152 gnd.n6776 gnd.n399 240.244
R6153 gnd.n6781 gnd.n399 240.244
R6154 gnd.n6781 gnd.n395 240.244
R6155 gnd.n6787 gnd.n395 240.244
R6156 gnd.n4296 gnd.n882 240.244
R6157 gnd.n4296 gnd.n4292 240.244
R6158 gnd.n4302 gnd.n4292 240.244
R6159 gnd.n4303 gnd.n4302 240.244
R6160 gnd.n4304 gnd.n4303 240.244
R6161 gnd.n4304 gnd.n2061 240.244
R6162 gnd.n4314 gnd.n2061 240.244
R6163 gnd.n4314 gnd.n2062 240.244
R6164 gnd.n2062 gnd.n2048 240.244
R6165 gnd.n4598 gnd.n2048 240.244
R6166 gnd.n4599 gnd.n4598 240.244
R6167 gnd.n4599 gnd.n2044 240.244
R6168 gnd.n4605 gnd.n2044 240.244
R6169 gnd.n4606 gnd.n4605 240.244
R6170 gnd.n4607 gnd.n4606 240.244
R6171 gnd.n4607 gnd.n2039 240.244
R6172 gnd.n4621 gnd.n2039 240.244
R6173 gnd.n4621 gnd.n2040 240.244
R6174 gnd.n4617 gnd.n2040 240.244
R6175 gnd.n4617 gnd.n4616 240.244
R6176 gnd.n4616 gnd.n2014 240.244
R6177 gnd.n4635 gnd.n2014 240.244
R6178 gnd.n4635 gnd.n2010 240.244
R6179 gnd.n4641 gnd.n2010 240.244
R6180 gnd.n4641 gnd.n1998 240.244
R6181 gnd.n4668 gnd.n1998 240.244
R6182 gnd.n4668 gnd.n1993 240.244
R6183 gnd.n4683 gnd.n1993 240.244
R6184 gnd.n4683 gnd.n1994 240.244
R6185 gnd.n4679 gnd.n1994 240.244
R6186 gnd.n4679 gnd.n4678 240.244
R6187 gnd.n4678 gnd.n1116 240.244
R6188 gnd.n5896 gnd.n1116 240.244
R6189 gnd.n5896 gnd.n1117 240.244
R6190 gnd.n5892 gnd.n1117 240.244
R6191 gnd.n5892 gnd.n1123 240.244
R6192 gnd.n4864 gnd.n1123 240.244
R6193 gnd.n4870 gnd.n4864 240.244
R6194 gnd.n4870 gnd.n1887 240.244
R6195 gnd.n4893 gnd.n1887 240.244
R6196 gnd.n4893 gnd.n1882 240.244
R6197 gnd.n4910 gnd.n1882 240.244
R6198 gnd.n4910 gnd.n1883 240.244
R6199 gnd.n4906 gnd.n1883 240.244
R6200 gnd.n4906 gnd.n4905 240.244
R6201 gnd.n4905 gnd.n4904 240.244
R6202 gnd.n4904 gnd.n1849 240.244
R6203 gnd.n4951 gnd.n1849 240.244
R6204 gnd.n4951 gnd.n1845 240.244
R6205 gnd.n4957 gnd.n1845 240.244
R6206 gnd.n4957 gnd.n1831 240.244
R6207 gnd.n4977 gnd.n1831 240.244
R6208 gnd.n4977 gnd.n1826 240.244
R6209 gnd.n4985 gnd.n1826 240.244
R6210 gnd.n4985 gnd.n1827 240.244
R6211 gnd.n1827 gnd.n1807 240.244
R6212 gnd.n5016 gnd.n1807 240.244
R6213 gnd.n5016 gnd.n1802 240.244
R6214 gnd.n5033 gnd.n1802 240.244
R6215 gnd.n5033 gnd.n1803 240.244
R6216 gnd.n5029 gnd.n1803 240.244
R6217 gnd.n5029 gnd.n5028 240.244
R6218 gnd.n5028 gnd.n5027 240.244
R6219 gnd.n5027 gnd.n1768 240.244
R6220 gnd.n5074 gnd.n1768 240.244
R6221 gnd.n5074 gnd.n1764 240.244
R6222 gnd.n5080 gnd.n1764 240.244
R6223 gnd.n5080 gnd.n1749 240.244
R6224 gnd.n5099 gnd.n1749 240.244
R6225 gnd.n5099 gnd.n1744 240.244
R6226 gnd.n5107 gnd.n1744 240.244
R6227 gnd.n5107 gnd.n1745 240.244
R6228 gnd.n1745 gnd.n1724 240.244
R6229 gnd.n5137 gnd.n1724 240.244
R6230 gnd.n5137 gnd.n1719 240.244
R6231 gnd.n5151 gnd.n1719 240.244
R6232 gnd.n5151 gnd.n1720 240.244
R6233 gnd.n5147 gnd.n1720 240.244
R6234 gnd.n5147 gnd.n5146 240.244
R6235 gnd.n5146 gnd.n1690 240.244
R6236 gnd.n5183 gnd.n1690 240.244
R6237 gnd.n5183 gnd.n1685 240.244
R6238 gnd.n5191 gnd.n1685 240.244
R6239 gnd.n5191 gnd.n1686 240.244
R6240 gnd.n1686 gnd.n1662 240.244
R6241 gnd.n5218 gnd.n1662 240.244
R6242 gnd.n5218 gnd.n1658 240.244
R6243 gnd.n5224 gnd.n1658 240.244
R6244 gnd.n5224 gnd.n1633 240.244
R6245 gnd.n5255 gnd.n1633 240.244
R6246 gnd.n5255 gnd.n1628 240.244
R6247 gnd.n5263 gnd.n1628 240.244
R6248 gnd.n5263 gnd.n1629 240.244
R6249 gnd.n1629 gnd.n1533 240.244
R6250 gnd.n5405 gnd.n1533 240.244
R6251 gnd.n5405 gnd.n1529 240.244
R6252 gnd.n5411 gnd.n1529 240.244
R6253 gnd.n5411 gnd.n1520 240.244
R6254 gnd.n5421 gnd.n1520 240.244
R6255 gnd.n5421 gnd.n1516 240.244
R6256 gnd.n5430 gnd.n1516 240.244
R6257 gnd.n5430 gnd.n1507 240.244
R6258 gnd.n5440 gnd.n1507 240.244
R6259 gnd.n5441 gnd.n5440 240.244
R6260 gnd.n5441 gnd.n1220 240.244
R6261 gnd.n1502 gnd.n1220 240.244
R6262 gnd.n5459 gnd.n1502 240.244
R6263 gnd.n5459 gnd.n1503 240.244
R6264 gnd.n5455 gnd.n1503 240.244
R6265 gnd.n5455 gnd.n5454 240.244
R6266 gnd.n5454 gnd.n5453 240.244
R6267 gnd.n5453 gnd.n1472 240.244
R6268 gnd.n5527 gnd.n1472 240.244
R6269 gnd.n5527 gnd.n1468 240.244
R6270 gnd.n5533 gnd.n1468 240.244
R6271 gnd.n5534 gnd.n5533 240.244
R6272 gnd.n5535 gnd.n5534 240.244
R6273 gnd.n5535 gnd.n1464 240.244
R6274 gnd.n5541 gnd.n1464 240.244
R6275 gnd.n5542 gnd.n5541 240.244
R6276 gnd.n5543 gnd.n5542 240.244
R6277 gnd.n5543 gnd.n1459 240.244
R6278 gnd.n5552 gnd.n1459 240.244
R6279 gnd.n5552 gnd.n1460 240.244
R6280 gnd.n1460 gnd.n389 240.244
R6281 gnd.n6792 gnd.n389 240.244
R6282 gnd.n6792 gnd.n390 240.244
R6283 gnd.n6788 gnd.n390 240.244
R6284 gnd.n6249 gnd.n716 240.244
R6285 gnd.n6245 gnd.n716 240.244
R6286 gnd.n6245 gnd.n718 240.244
R6287 gnd.n6241 gnd.n718 240.244
R6288 gnd.n6241 gnd.n723 240.244
R6289 gnd.n6237 gnd.n723 240.244
R6290 gnd.n6237 gnd.n725 240.244
R6291 gnd.n6233 gnd.n725 240.244
R6292 gnd.n6233 gnd.n731 240.244
R6293 gnd.n6229 gnd.n731 240.244
R6294 gnd.n6229 gnd.n733 240.244
R6295 gnd.n6225 gnd.n733 240.244
R6296 gnd.n6225 gnd.n739 240.244
R6297 gnd.n6221 gnd.n739 240.244
R6298 gnd.n6221 gnd.n741 240.244
R6299 gnd.n6217 gnd.n741 240.244
R6300 gnd.n6217 gnd.n747 240.244
R6301 gnd.n6213 gnd.n747 240.244
R6302 gnd.n6213 gnd.n749 240.244
R6303 gnd.n6209 gnd.n749 240.244
R6304 gnd.n6209 gnd.n755 240.244
R6305 gnd.n6205 gnd.n755 240.244
R6306 gnd.n6205 gnd.n757 240.244
R6307 gnd.n6201 gnd.n757 240.244
R6308 gnd.n6201 gnd.n763 240.244
R6309 gnd.n6197 gnd.n763 240.244
R6310 gnd.n6197 gnd.n765 240.244
R6311 gnd.n6193 gnd.n765 240.244
R6312 gnd.n6193 gnd.n771 240.244
R6313 gnd.n6189 gnd.n771 240.244
R6314 gnd.n6189 gnd.n773 240.244
R6315 gnd.n6185 gnd.n773 240.244
R6316 gnd.n6185 gnd.n779 240.244
R6317 gnd.n6181 gnd.n779 240.244
R6318 gnd.n6181 gnd.n781 240.244
R6319 gnd.n6177 gnd.n781 240.244
R6320 gnd.n6177 gnd.n787 240.244
R6321 gnd.n6173 gnd.n787 240.244
R6322 gnd.n6173 gnd.n789 240.244
R6323 gnd.n6169 gnd.n789 240.244
R6324 gnd.n6169 gnd.n795 240.244
R6325 gnd.n6165 gnd.n795 240.244
R6326 gnd.n6165 gnd.n797 240.244
R6327 gnd.n6161 gnd.n797 240.244
R6328 gnd.n6161 gnd.n803 240.244
R6329 gnd.n6157 gnd.n803 240.244
R6330 gnd.n6157 gnd.n805 240.244
R6331 gnd.n6153 gnd.n805 240.244
R6332 gnd.n6153 gnd.n811 240.244
R6333 gnd.n6149 gnd.n811 240.244
R6334 gnd.n6149 gnd.n813 240.244
R6335 gnd.n6145 gnd.n813 240.244
R6336 gnd.n6145 gnd.n819 240.244
R6337 gnd.n6141 gnd.n819 240.244
R6338 gnd.n6141 gnd.n821 240.244
R6339 gnd.n6137 gnd.n821 240.244
R6340 gnd.n6137 gnd.n827 240.244
R6341 gnd.n6133 gnd.n827 240.244
R6342 gnd.n6133 gnd.n829 240.244
R6343 gnd.n6129 gnd.n829 240.244
R6344 gnd.n6129 gnd.n835 240.244
R6345 gnd.n6125 gnd.n835 240.244
R6346 gnd.n6125 gnd.n837 240.244
R6347 gnd.n6121 gnd.n837 240.244
R6348 gnd.n6121 gnd.n843 240.244
R6349 gnd.n6117 gnd.n843 240.244
R6350 gnd.n6117 gnd.n845 240.244
R6351 gnd.n6113 gnd.n845 240.244
R6352 gnd.n6113 gnd.n851 240.244
R6353 gnd.n6109 gnd.n851 240.244
R6354 gnd.n6109 gnd.n853 240.244
R6355 gnd.n6105 gnd.n853 240.244
R6356 gnd.n6105 gnd.n859 240.244
R6357 gnd.n6101 gnd.n859 240.244
R6358 gnd.n6101 gnd.n861 240.244
R6359 gnd.n6097 gnd.n861 240.244
R6360 gnd.n6097 gnd.n867 240.244
R6361 gnd.n6093 gnd.n867 240.244
R6362 gnd.n6093 gnd.n869 240.244
R6363 gnd.n6089 gnd.n869 240.244
R6364 gnd.n6089 gnd.n875 240.244
R6365 gnd.n6085 gnd.n875 240.244
R6366 gnd.n6085 gnd.n877 240.244
R6367 gnd.n6081 gnd.n877 240.244
R6368 gnd.n4351 gnd.n2009 240.244
R6369 gnd.n4344 gnd.n2009 240.244
R6370 gnd.n4344 gnd.n2000 240.244
R6371 gnd.n2000 gnd.n1989 240.244
R6372 gnd.n4685 gnd.n1989 240.244
R6373 gnd.n4685 gnd.n1985 240.244
R6374 gnd.n4691 gnd.n1985 240.244
R6375 gnd.n4692 gnd.n4691 240.244
R6376 gnd.n4693 gnd.n4692 240.244
R6377 gnd.n4693 gnd.n1113 240.244
R6378 gnd.n4840 gnd.n1113 240.244
R6379 gnd.n4840 gnd.n1124 240.244
R6380 gnd.n4698 gnd.n1124 240.244
R6381 gnd.n4698 gnd.n1900 240.244
R6382 gnd.n1900 gnd.n1898 240.244
R6383 gnd.n1898 gnd.n1895 240.244
R6384 gnd.n1895 gnd.n1888 240.244
R6385 gnd.n4701 gnd.n1888 240.244
R6386 gnd.n4701 gnd.n1881 240.244
R6387 gnd.n4704 gnd.n1881 240.244
R6388 gnd.n4705 gnd.n4704 240.244
R6389 gnd.n4706 gnd.n4705 240.244
R6390 gnd.n4707 gnd.n4706 240.244
R6391 gnd.n4707 gnd.n1856 240.244
R6392 gnd.n1856 gnd.n1850 240.244
R6393 gnd.n4710 gnd.n1850 240.244
R6394 gnd.n4710 gnd.n1843 240.244
R6395 gnd.n4711 gnd.n1843 240.244
R6396 gnd.n4711 gnd.n1832 240.244
R6397 gnd.n4714 gnd.n1832 240.244
R6398 gnd.n4714 gnd.n1825 240.244
R6399 gnd.n4715 gnd.n1825 240.244
R6400 gnd.n4715 gnd.n1816 240.244
R6401 gnd.n1816 gnd.n1808 240.244
R6402 gnd.n4718 gnd.n1808 240.244
R6403 gnd.n4718 gnd.n1801 240.244
R6404 gnd.n4721 gnd.n1801 240.244
R6405 gnd.n4722 gnd.n4721 240.244
R6406 gnd.n4723 gnd.n4722 240.244
R6407 gnd.n4724 gnd.n4723 240.244
R6408 gnd.n4724 gnd.n1777 240.244
R6409 gnd.n1777 gnd.n1770 240.244
R6410 gnd.n4727 gnd.n1770 240.244
R6411 gnd.n4727 gnd.n1762 240.244
R6412 gnd.n4730 gnd.n1762 240.244
R6413 gnd.n4730 gnd.n1750 240.244
R6414 gnd.n4731 gnd.n1750 240.244
R6415 gnd.n4731 gnd.n1743 240.244
R6416 gnd.n4734 gnd.n1743 240.244
R6417 gnd.n4734 gnd.n1733 240.244
R6418 gnd.n1733 gnd.n1725 240.244
R6419 gnd.n4736 gnd.n1725 240.244
R6420 gnd.n4736 gnd.n1717 240.244
R6421 gnd.n4739 gnd.n1717 240.244
R6422 gnd.n4740 gnd.n4739 240.244
R6423 gnd.n4743 gnd.n4740 240.244
R6424 gnd.n4744 gnd.n4743 240.244
R6425 gnd.n4744 gnd.n1693 240.244
R6426 gnd.n4745 gnd.n1693 240.244
R6427 gnd.n4745 gnd.n1683 240.244
R6428 gnd.n4748 gnd.n1683 240.244
R6429 gnd.n4749 gnd.n4748 240.244
R6430 gnd.n4749 gnd.n1664 240.244
R6431 gnd.n4750 gnd.n1664 240.244
R6432 gnd.n4750 gnd.n1655 240.244
R6433 gnd.n4753 gnd.n1655 240.244
R6434 gnd.n4753 gnd.n1635 240.244
R6435 gnd.n1635 gnd.n1624 240.244
R6436 gnd.n5265 gnd.n1624 240.244
R6437 gnd.n5265 gnd.n1619 240.244
R6438 gnd.n5272 gnd.n1619 240.244
R6439 gnd.n5272 gnd.n1534 240.244
R6440 gnd.n1534 gnd.n1525 240.244
R6441 gnd.n5413 gnd.n1525 240.244
R6442 gnd.n5413 gnd.n1521 240.244
R6443 gnd.n5419 gnd.n1521 240.244
R6444 gnd.n5419 gnd.n1513 240.244
R6445 gnd.n5432 gnd.n1513 240.244
R6446 gnd.n5432 gnd.n1509 240.244
R6447 gnd.n5438 gnd.n1509 240.244
R6448 gnd.n5438 gnd.n1222 240.244
R6449 gnd.n5780 gnd.n1222 240.244
R6450 gnd.n4356 gnd.n4355 240.244
R6451 gnd.n4339 gnd.n4338 240.244
R6452 gnd.n4364 gnd.n4363 240.244
R6453 gnd.n4366 gnd.n4365 240.244
R6454 gnd.n4373 gnd.n4372 240.244
R6455 gnd.n4375 gnd.n4374 240.244
R6456 gnd.n4385 gnd.n4384 240.244
R6457 gnd.n4393 gnd.n4392 240.244
R6458 gnd.n4395 gnd.n4394 240.244
R6459 gnd.n4405 gnd.n4404 240.244
R6460 gnd.n4413 gnd.n4412 240.244
R6461 gnd.n4415 gnd.n4414 240.244
R6462 gnd.n4427 gnd.n4426 240.244
R6463 gnd.n4632 gnd.n2030 240.244
R6464 gnd.n4643 gnd.n2007 240.244
R6465 gnd.n4643 gnd.n2001 240.244
R6466 gnd.n4666 gnd.n2001 240.244
R6467 gnd.n4666 gnd.n2002 240.244
R6468 gnd.n2002 gnd.n1992 240.244
R6469 gnd.n4648 gnd.n1992 240.244
R6470 gnd.n4649 gnd.n4648 240.244
R6471 gnd.n4652 gnd.n4649 240.244
R6472 gnd.n4653 gnd.n4652 240.244
R6473 gnd.n4653 gnd.n1115 240.244
R6474 gnd.n1126 gnd.n1115 240.244
R6475 gnd.n5890 gnd.n1126 240.244
R6476 gnd.n5890 gnd.n1127 240.244
R6477 gnd.n1132 gnd.n1127 240.244
R6478 gnd.n1133 gnd.n1132 240.244
R6479 gnd.n1134 gnd.n1133 240.244
R6480 gnd.n4891 gnd.n1134 240.244
R6481 gnd.n4891 gnd.n1137 240.244
R6482 gnd.n1138 gnd.n1137 240.244
R6483 gnd.n1139 gnd.n1138 240.244
R6484 gnd.n1868 gnd.n1139 240.244
R6485 gnd.n1868 gnd.n1142 240.244
R6486 gnd.n1143 gnd.n1142 240.244
R6487 gnd.n1144 gnd.n1143 240.244
R6488 gnd.n4949 gnd.n1144 240.244
R6489 gnd.n4949 gnd.n1147 240.244
R6490 gnd.n1148 gnd.n1147 240.244
R6491 gnd.n1149 gnd.n1148 240.244
R6492 gnd.n4975 gnd.n1149 240.244
R6493 gnd.n4975 gnd.n1152 240.244
R6494 gnd.n1153 gnd.n1152 240.244
R6495 gnd.n1154 gnd.n1153 240.244
R6496 gnd.n5006 gnd.n1154 240.244
R6497 gnd.n5006 gnd.n1157 240.244
R6498 gnd.n1158 gnd.n1157 240.244
R6499 gnd.n1159 gnd.n1158 240.244
R6500 gnd.n1794 gnd.n1159 240.244
R6501 gnd.n1794 gnd.n1162 240.244
R6502 gnd.n1163 gnd.n1162 240.244
R6503 gnd.n1164 gnd.n1163 240.244
R6504 gnd.n1778 gnd.n1164 240.244
R6505 gnd.n1778 gnd.n1167 240.244
R6506 gnd.n1168 gnd.n1167 240.244
R6507 gnd.n1169 gnd.n1168 240.244
R6508 gnd.n1754 gnd.n1169 240.244
R6509 gnd.n1754 gnd.n1172 240.244
R6510 gnd.n1173 gnd.n1172 240.244
R6511 gnd.n1174 gnd.n1173 240.244
R6512 gnd.n1736 gnd.n1174 240.244
R6513 gnd.n1736 gnd.n1177 240.244
R6514 gnd.n1178 gnd.n1177 240.244
R6515 gnd.n1179 gnd.n1178 240.244
R6516 gnd.n1718 gnd.n1179 240.244
R6517 gnd.n1718 gnd.n1182 240.244
R6518 gnd.n1183 gnd.n1182 240.244
R6519 gnd.n1184 gnd.n1183 240.244
R6520 gnd.n1700 gnd.n1184 240.244
R6521 gnd.n1700 gnd.n1187 240.244
R6522 gnd.n1188 gnd.n1187 240.244
R6523 gnd.n1189 gnd.n1188 240.244
R6524 gnd.n1676 gnd.n1189 240.244
R6525 gnd.n1676 gnd.n1192 240.244
R6526 gnd.n1193 gnd.n1192 240.244
R6527 gnd.n1194 gnd.n1193 240.244
R6528 gnd.n1657 gnd.n1194 240.244
R6529 gnd.n1657 gnd.n1197 240.244
R6530 gnd.n1198 gnd.n1197 240.244
R6531 gnd.n1199 gnd.n1198 240.244
R6532 gnd.n1627 gnd.n1199 240.244
R6533 gnd.n1627 gnd.n1202 240.244
R6534 gnd.n1203 gnd.n1202 240.244
R6535 gnd.n1204 gnd.n1203 240.244
R6536 gnd.n1536 gnd.n1204 240.244
R6537 gnd.n1536 gnd.n1207 240.244
R6538 gnd.n1208 gnd.n1207 240.244
R6539 gnd.n1209 gnd.n1208 240.244
R6540 gnd.n1514 gnd.n1209 240.244
R6541 gnd.n1514 gnd.n1212 240.244
R6542 gnd.n1213 gnd.n1212 240.244
R6543 gnd.n1214 gnd.n1213 240.244
R6544 gnd.n1217 gnd.n1214 240.244
R6545 gnd.n5782 gnd.n1217 240.244
R6546 gnd.n1228 gnd.n1227 240.244
R6547 gnd.n1480 gnd.n1231 240.244
R6548 gnd.n1233 gnd.n1232 240.244
R6549 gnd.n1483 gnd.n1237 240.244
R6550 gnd.n1486 gnd.n1238 240.244
R6551 gnd.n1247 gnd.n1246 240.244
R6552 gnd.n1488 gnd.n1254 240.244
R6553 gnd.n1491 gnd.n1255 240.244
R6554 gnd.n1263 gnd.n1262 240.244
R6555 gnd.n1493 gnd.n1270 240.244
R6556 gnd.n1496 gnd.n1271 240.244
R6557 gnd.n1279 gnd.n1278 240.244
R6558 gnd.n1499 gnd.n1478 240.244
R6559 gnd.n5462 gnd.n1218 240.244
R6560 gnd.n1094 gnd.n1093 240.132
R6561 gnd.n1553 gnd.n1552 240.132
R6562 gnd.n6256 gnd.n711 225.874
R6563 gnd.n6257 gnd.n6256 225.874
R6564 gnd.n6258 gnd.n6257 225.874
R6565 gnd.n6258 gnd.n705 225.874
R6566 gnd.n6266 gnd.n705 225.874
R6567 gnd.n6267 gnd.n6266 225.874
R6568 gnd.n6268 gnd.n6267 225.874
R6569 gnd.n6268 gnd.n699 225.874
R6570 gnd.n6276 gnd.n699 225.874
R6571 gnd.n6277 gnd.n6276 225.874
R6572 gnd.n6278 gnd.n6277 225.874
R6573 gnd.n6278 gnd.n693 225.874
R6574 gnd.n6286 gnd.n693 225.874
R6575 gnd.n6287 gnd.n6286 225.874
R6576 gnd.n6288 gnd.n6287 225.874
R6577 gnd.n6288 gnd.n687 225.874
R6578 gnd.n6296 gnd.n687 225.874
R6579 gnd.n6297 gnd.n6296 225.874
R6580 gnd.n6298 gnd.n6297 225.874
R6581 gnd.n6298 gnd.n681 225.874
R6582 gnd.n6306 gnd.n681 225.874
R6583 gnd.n6307 gnd.n6306 225.874
R6584 gnd.n6308 gnd.n6307 225.874
R6585 gnd.n6308 gnd.n675 225.874
R6586 gnd.n6316 gnd.n675 225.874
R6587 gnd.n6317 gnd.n6316 225.874
R6588 gnd.n6318 gnd.n6317 225.874
R6589 gnd.n6318 gnd.n669 225.874
R6590 gnd.n6326 gnd.n669 225.874
R6591 gnd.n6327 gnd.n6326 225.874
R6592 gnd.n6328 gnd.n6327 225.874
R6593 gnd.n6328 gnd.n663 225.874
R6594 gnd.n6336 gnd.n663 225.874
R6595 gnd.n6337 gnd.n6336 225.874
R6596 gnd.n6338 gnd.n6337 225.874
R6597 gnd.n6338 gnd.n657 225.874
R6598 gnd.n6346 gnd.n657 225.874
R6599 gnd.n6347 gnd.n6346 225.874
R6600 gnd.n6348 gnd.n6347 225.874
R6601 gnd.n6348 gnd.n651 225.874
R6602 gnd.n6356 gnd.n651 225.874
R6603 gnd.n6357 gnd.n6356 225.874
R6604 gnd.n6358 gnd.n6357 225.874
R6605 gnd.n6358 gnd.n645 225.874
R6606 gnd.n6366 gnd.n645 225.874
R6607 gnd.n6367 gnd.n6366 225.874
R6608 gnd.n6368 gnd.n6367 225.874
R6609 gnd.n6368 gnd.n639 225.874
R6610 gnd.n6376 gnd.n639 225.874
R6611 gnd.n6377 gnd.n6376 225.874
R6612 gnd.n6378 gnd.n6377 225.874
R6613 gnd.n6378 gnd.n633 225.874
R6614 gnd.n6386 gnd.n633 225.874
R6615 gnd.n6387 gnd.n6386 225.874
R6616 gnd.n6388 gnd.n6387 225.874
R6617 gnd.n6388 gnd.n627 225.874
R6618 gnd.n6396 gnd.n627 225.874
R6619 gnd.n6397 gnd.n6396 225.874
R6620 gnd.n6398 gnd.n6397 225.874
R6621 gnd.n6398 gnd.n621 225.874
R6622 gnd.n6406 gnd.n621 225.874
R6623 gnd.n6407 gnd.n6406 225.874
R6624 gnd.n6408 gnd.n6407 225.874
R6625 gnd.n6408 gnd.n615 225.874
R6626 gnd.n6416 gnd.n615 225.874
R6627 gnd.n6417 gnd.n6416 225.874
R6628 gnd.n6418 gnd.n6417 225.874
R6629 gnd.n6418 gnd.n609 225.874
R6630 gnd.n6426 gnd.n609 225.874
R6631 gnd.n6427 gnd.n6426 225.874
R6632 gnd.n6428 gnd.n6427 225.874
R6633 gnd.n6428 gnd.n603 225.874
R6634 gnd.n6436 gnd.n603 225.874
R6635 gnd.n6437 gnd.n6436 225.874
R6636 gnd.n6438 gnd.n6437 225.874
R6637 gnd.n6438 gnd.n597 225.874
R6638 gnd.n6446 gnd.n597 225.874
R6639 gnd.n6447 gnd.n6446 225.874
R6640 gnd.n6448 gnd.n6447 225.874
R6641 gnd.n6448 gnd.n591 225.874
R6642 gnd.n6456 gnd.n591 225.874
R6643 gnd.n6457 gnd.n6456 225.874
R6644 gnd.n6458 gnd.n6457 225.874
R6645 gnd.n6458 gnd.n585 225.874
R6646 gnd.n6466 gnd.n585 225.874
R6647 gnd.n6467 gnd.n6466 225.874
R6648 gnd.n6468 gnd.n6467 225.874
R6649 gnd.n6468 gnd.n579 225.874
R6650 gnd.n6476 gnd.n579 225.874
R6651 gnd.n6477 gnd.n6476 225.874
R6652 gnd.n6478 gnd.n6477 225.874
R6653 gnd.n6478 gnd.n573 225.874
R6654 gnd.n6486 gnd.n573 225.874
R6655 gnd.n6487 gnd.n6486 225.874
R6656 gnd.n6488 gnd.n6487 225.874
R6657 gnd.n6488 gnd.n567 225.874
R6658 gnd.n6496 gnd.n567 225.874
R6659 gnd.n6497 gnd.n6496 225.874
R6660 gnd.n6498 gnd.n6497 225.874
R6661 gnd.n6498 gnd.n561 225.874
R6662 gnd.n6506 gnd.n561 225.874
R6663 gnd.n6507 gnd.n6506 225.874
R6664 gnd.n6508 gnd.n6507 225.874
R6665 gnd.n6508 gnd.n555 225.874
R6666 gnd.n6516 gnd.n555 225.874
R6667 gnd.n6517 gnd.n6516 225.874
R6668 gnd.n6518 gnd.n6517 225.874
R6669 gnd.n6518 gnd.n549 225.874
R6670 gnd.n6526 gnd.n549 225.874
R6671 gnd.n6527 gnd.n6526 225.874
R6672 gnd.n6528 gnd.n6527 225.874
R6673 gnd.n6528 gnd.n543 225.874
R6674 gnd.n6536 gnd.n543 225.874
R6675 gnd.n6537 gnd.n6536 225.874
R6676 gnd.n6538 gnd.n6537 225.874
R6677 gnd.n6538 gnd.n537 225.874
R6678 gnd.n6546 gnd.n537 225.874
R6679 gnd.n6547 gnd.n6546 225.874
R6680 gnd.n6548 gnd.n6547 225.874
R6681 gnd.n6548 gnd.n531 225.874
R6682 gnd.n6556 gnd.n531 225.874
R6683 gnd.n6557 gnd.n6556 225.874
R6684 gnd.n6558 gnd.n6557 225.874
R6685 gnd.n6558 gnd.n525 225.874
R6686 gnd.n6567 gnd.n525 225.874
R6687 gnd.n6568 gnd.n6567 225.874
R6688 gnd.n6569 gnd.n6568 225.874
R6689 gnd.n6569 gnd.n520 225.874
R6690 gnd.n2816 gnd.t60 224.174
R6691 gnd.n2309 gnd.t55 224.174
R6692 gnd.n1363 gnd.n1300 199.319
R6693 gnd.n1363 gnd.n1301 199.319
R6694 gnd.n1046 gnd.n1006 199.319
R6695 gnd.n1046 gnd.n1005 199.319
R6696 gnd.n1095 gnd.n1092 186.49
R6697 gnd.n1554 gnd.n1551 186.49
R6698 gnd.n3591 gnd.n3590 185
R6699 gnd.n3589 gnd.n3588 185
R6700 gnd.n3568 gnd.n3567 185
R6701 gnd.n3583 gnd.n3582 185
R6702 gnd.n3581 gnd.n3580 185
R6703 gnd.n3572 gnd.n3571 185
R6704 gnd.n3575 gnd.n3574 185
R6705 gnd.n3559 gnd.n3558 185
R6706 gnd.n3557 gnd.n3556 185
R6707 gnd.n3536 gnd.n3535 185
R6708 gnd.n3551 gnd.n3550 185
R6709 gnd.n3549 gnd.n3548 185
R6710 gnd.n3540 gnd.n3539 185
R6711 gnd.n3543 gnd.n3542 185
R6712 gnd.n3527 gnd.n3526 185
R6713 gnd.n3525 gnd.n3524 185
R6714 gnd.n3504 gnd.n3503 185
R6715 gnd.n3519 gnd.n3518 185
R6716 gnd.n3517 gnd.n3516 185
R6717 gnd.n3508 gnd.n3507 185
R6718 gnd.n3511 gnd.n3510 185
R6719 gnd.n3496 gnd.n3495 185
R6720 gnd.n3494 gnd.n3493 185
R6721 gnd.n3473 gnd.n3472 185
R6722 gnd.n3488 gnd.n3487 185
R6723 gnd.n3486 gnd.n3485 185
R6724 gnd.n3477 gnd.n3476 185
R6725 gnd.n3480 gnd.n3479 185
R6726 gnd.n3464 gnd.n3463 185
R6727 gnd.n3462 gnd.n3461 185
R6728 gnd.n3441 gnd.n3440 185
R6729 gnd.n3456 gnd.n3455 185
R6730 gnd.n3454 gnd.n3453 185
R6731 gnd.n3445 gnd.n3444 185
R6732 gnd.n3448 gnd.n3447 185
R6733 gnd.n3432 gnd.n3431 185
R6734 gnd.n3430 gnd.n3429 185
R6735 gnd.n3409 gnd.n3408 185
R6736 gnd.n3424 gnd.n3423 185
R6737 gnd.n3422 gnd.n3421 185
R6738 gnd.n3413 gnd.n3412 185
R6739 gnd.n3416 gnd.n3415 185
R6740 gnd.n3400 gnd.n3399 185
R6741 gnd.n3398 gnd.n3397 185
R6742 gnd.n3377 gnd.n3376 185
R6743 gnd.n3392 gnd.n3391 185
R6744 gnd.n3390 gnd.n3389 185
R6745 gnd.n3381 gnd.n3380 185
R6746 gnd.n3384 gnd.n3383 185
R6747 gnd.n3369 gnd.n3368 185
R6748 gnd.n3367 gnd.n3366 185
R6749 gnd.n3346 gnd.n3345 185
R6750 gnd.n3361 gnd.n3360 185
R6751 gnd.n3359 gnd.n3358 185
R6752 gnd.n3350 gnd.n3349 185
R6753 gnd.n3353 gnd.n3352 185
R6754 gnd.n2817 gnd.t59 178.987
R6755 gnd.n2310 gnd.t56 178.987
R6756 gnd.n1 gnd.t363 170.774
R6757 gnd.n7 gnd.t10 170.103
R6758 gnd.n6 gnd.t1 170.103
R6759 gnd.n5 gnd.t175 170.103
R6760 gnd.n4 gnd.t23 170.103
R6761 gnd.n3 gnd.t3 170.103
R6762 gnd.n2 gnd.t49 170.103
R6763 gnd.n1 gnd.t359 170.103
R6764 gnd.n5395 gnd.n1563 163.367
R6765 gnd.n5391 gnd.n5390 163.367
R6766 gnd.n5388 gnd.n1566 163.367
R6767 gnd.n5384 gnd.n5383 163.367
R6768 gnd.n5381 gnd.n1569 163.367
R6769 gnd.n5377 gnd.n5376 163.367
R6770 gnd.n5374 gnd.n1572 163.367
R6771 gnd.n5370 gnd.n5369 163.367
R6772 gnd.n5367 gnd.n1575 163.367
R6773 gnd.n5363 gnd.n5362 163.367
R6774 gnd.n5360 gnd.n1578 163.367
R6775 gnd.n5356 gnd.n5355 163.367
R6776 gnd.n5353 gnd.n1581 163.367
R6777 gnd.n5349 gnd.n5348 163.367
R6778 gnd.n5346 gnd.n1584 163.367
R6779 gnd.n5342 gnd.n5341 163.367
R6780 gnd.n5338 gnd.n5337 163.367
R6781 gnd.n5335 gnd.n1590 163.367
R6782 gnd.n5330 gnd.n5329 163.367
R6783 gnd.n5327 gnd.n1595 163.367
R6784 gnd.n5323 gnd.n5322 163.367
R6785 gnd.n5320 gnd.n1598 163.367
R6786 gnd.n5316 gnd.n5315 163.367
R6787 gnd.n5313 gnd.n1601 163.367
R6788 gnd.n5309 gnd.n5308 163.367
R6789 gnd.n5306 gnd.n1604 163.367
R6790 gnd.n5302 gnd.n5301 163.367
R6791 gnd.n5299 gnd.n1607 163.367
R6792 gnd.n5295 gnd.n5294 163.367
R6793 gnd.n5292 gnd.n1610 163.367
R6794 gnd.n5288 gnd.n5287 163.367
R6795 gnd.n5285 gnd.n1613 163.367
R6796 gnd.n1974 gnd.n1111 163.367
R6797 gnd.n1112 gnd.n1111 163.367
R6798 gnd.n1979 gnd.n1112 163.367
R6799 gnd.n1980 gnd.n1979 163.367
R6800 gnd.n4850 gnd.n1980 163.367
R6801 gnd.n4850 gnd.n1905 163.367
R6802 gnd.n4855 gnd.n1905 163.367
R6803 gnd.n4855 gnd.n1906 163.367
R6804 gnd.n1906 gnd.n1897 163.367
R6805 gnd.n4873 gnd.n1897 163.367
R6806 gnd.n4873 gnd.n1894 163.367
R6807 gnd.n4881 gnd.n1894 163.367
R6808 gnd.n4881 gnd.n1889 163.367
R6809 gnd.n4877 gnd.n1889 163.367
R6810 gnd.n4877 gnd.n1880 163.367
R6811 gnd.n1880 gnd.n1872 163.367
R6812 gnd.n4918 gnd.n1872 163.367
R6813 gnd.n4918 gnd.n1870 163.367
R6814 gnd.n4922 gnd.n1870 163.367
R6815 gnd.n4922 gnd.n1861 163.367
R6816 gnd.n4931 gnd.n1861 163.367
R6817 gnd.n4931 gnd.n1858 163.367
R6818 gnd.n4941 gnd.n1858 163.367
R6819 gnd.n4941 gnd.n1859 163.367
R6820 gnd.n1859 gnd.n1851 163.367
R6821 gnd.n4936 gnd.n1851 163.367
R6822 gnd.n4936 gnd.n1842 163.367
R6823 gnd.n1842 gnd.n1835 163.367
R6824 gnd.n4967 gnd.n1835 163.367
R6825 gnd.n4967 gnd.n1833 163.367
R6826 gnd.n4973 gnd.n1833 163.367
R6827 gnd.n4973 gnd.n1824 163.367
R6828 gnd.n1824 gnd.n1818 163.367
R6829 gnd.n4995 gnd.n1818 163.367
R6830 gnd.n4996 gnd.n4995 163.367
R6831 gnd.n4996 gnd.n1815 163.367
R6832 gnd.n5004 gnd.n1815 163.367
R6833 gnd.n5004 gnd.n1809 163.367
R6834 gnd.n5000 gnd.n1809 163.367
R6835 gnd.n5000 gnd.n1800 163.367
R6836 gnd.n1800 gnd.n1791 163.367
R6837 gnd.n5042 gnd.n1791 163.367
R6838 gnd.n5042 gnd.n1789 163.367
R6839 gnd.n5046 gnd.n1789 163.367
R6840 gnd.n5046 gnd.n1782 163.367
R6841 gnd.n5055 gnd.n1782 163.367
R6842 gnd.n5055 gnd.n1779 163.367
R6843 gnd.n5065 gnd.n1779 163.367
R6844 gnd.n5065 gnd.n1780 163.367
R6845 gnd.n1780 gnd.n1771 163.367
R6846 gnd.n5060 gnd.n1771 163.367
R6847 gnd.n5060 gnd.n1761 163.367
R6848 gnd.n1761 gnd.n1753 163.367
R6849 gnd.n5090 gnd.n1753 163.367
R6850 gnd.n5090 gnd.n1751 163.367
R6851 gnd.n5096 gnd.n1751 163.367
R6852 gnd.n5096 gnd.n1742 163.367
R6853 gnd.n1742 gnd.n1735 163.367
R6854 gnd.n5117 gnd.n1735 163.367
R6855 gnd.n5118 gnd.n5117 163.367
R6856 gnd.n5118 gnd.n1732 163.367
R6857 gnd.n5126 gnd.n1732 163.367
R6858 gnd.n5126 gnd.n1726 163.367
R6859 gnd.n5122 gnd.n1726 163.367
R6860 gnd.n5122 gnd.n1716 163.367
R6861 gnd.n1716 gnd.n1709 163.367
R6862 gnd.n5160 gnd.n1709 163.367
R6863 gnd.n5160 gnd.n1707 163.367
R6864 gnd.n5164 gnd.n1707 163.367
R6865 gnd.n5164 gnd.n1698 163.367
R6866 gnd.n5175 gnd.n1698 163.367
R6867 gnd.n5175 gnd.n1694 163.367
R6868 gnd.n5181 gnd.n1694 163.367
R6869 gnd.n5181 gnd.n1696 163.367
R6870 gnd.n1696 gnd.n1682 163.367
R6871 gnd.n1682 gnd.n1674 163.367
R6872 gnd.n5200 gnd.n1674 163.367
R6873 gnd.n5200 gnd.n1671 163.367
R6874 gnd.n5210 gnd.n1671 163.367
R6875 gnd.n5210 gnd.n1672 163.367
R6876 gnd.n1672 gnd.n1665 163.367
R6877 gnd.n5205 gnd.n1665 163.367
R6878 gnd.n5205 gnd.n1654 163.367
R6879 gnd.n1654 gnd.n1648 163.367
R6880 gnd.n5233 gnd.n1648 163.367
R6881 gnd.n5234 gnd.n5233 163.367
R6882 gnd.n5234 gnd.n1636 163.367
R6883 gnd.n5239 gnd.n1636 163.367
R6884 gnd.n5240 gnd.n5239 163.367
R6885 gnd.n5240 gnd.n1646 163.367
R6886 gnd.n5244 gnd.n1646 163.367
R6887 gnd.n5244 gnd.n1617 163.367
R6888 gnd.n5275 gnd.n1617 163.367
R6889 gnd.n5275 gnd.n1535 163.367
R6890 gnd.n5279 gnd.n1535 163.367
R6891 gnd.n5280 gnd.n5279 163.367
R6892 gnd.n1086 gnd.n1085 163.367
R6893 gnd.n5962 gnd.n1085 163.367
R6894 gnd.n5960 gnd.n5959 163.367
R6895 gnd.n5956 gnd.n5955 163.367
R6896 gnd.n5952 gnd.n5951 163.367
R6897 gnd.n5948 gnd.n5947 163.367
R6898 gnd.n5944 gnd.n5943 163.367
R6899 gnd.n5940 gnd.n5939 163.367
R6900 gnd.n5936 gnd.n5935 163.367
R6901 gnd.n5932 gnd.n5931 163.367
R6902 gnd.n5928 gnd.n5927 163.367
R6903 gnd.n5924 gnd.n5923 163.367
R6904 gnd.n5920 gnd.n5919 163.367
R6905 gnd.n5916 gnd.n5915 163.367
R6906 gnd.n5912 gnd.n5911 163.367
R6907 gnd.n5908 gnd.n5907 163.367
R6908 gnd.n5971 gnd.n1051 163.367
R6909 gnd.n1912 gnd.n1911 163.367
R6910 gnd.n1917 gnd.n1916 163.367
R6911 gnd.n1921 gnd.n1920 163.367
R6912 gnd.n1925 gnd.n1924 163.367
R6913 gnd.n1929 gnd.n1928 163.367
R6914 gnd.n1933 gnd.n1932 163.367
R6915 gnd.n1937 gnd.n1936 163.367
R6916 gnd.n1941 gnd.n1940 163.367
R6917 gnd.n1945 gnd.n1944 163.367
R6918 gnd.n1949 gnd.n1948 163.367
R6919 gnd.n1953 gnd.n1952 163.367
R6920 gnd.n1957 gnd.n1956 163.367
R6921 gnd.n1961 gnd.n1960 163.367
R6922 gnd.n1965 gnd.n1964 163.367
R6923 gnd.n1969 gnd.n1968 163.367
R6924 gnd.n5900 gnd.n1087 163.367
R6925 gnd.n5900 gnd.n1109 163.367
R6926 gnd.n4844 gnd.n1109 163.367
R6927 gnd.n4844 gnd.n4843 163.367
R6928 gnd.n4848 gnd.n4843 163.367
R6929 gnd.n4848 gnd.n1903 163.367
R6930 gnd.n4857 gnd.n1903 163.367
R6931 gnd.n4857 gnd.n1901 163.367
R6932 gnd.n4861 gnd.n1901 163.367
R6933 gnd.n4861 gnd.n1893 163.367
R6934 gnd.n4885 gnd.n1893 163.367
R6935 gnd.n4885 gnd.n1891 163.367
R6936 gnd.n4889 gnd.n1891 163.367
R6937 gnd.n4889 gnd.n1878 163.367
R6938 gnd.n4912 gnd.n1878 163.367
R6939 gnd.n4912 gnd.n1876 163.367
R6940 gnd.n4916 gnd.n1876 163.367
R6941 gnd.n4916 gnd.n1867 163.367
R6942 gnd.n4925 gnd.n1867 163.367
R6943 gnd.n4925 gnd.n1865 163.367
R6944 gnd.n4929 gnd.n1865 163.367
R6945 gnd.n4929 gnd.n1855 163.367
R6946 gnd.n4943 gnd.n1855 163.367
R6947 gnd.n4943 gnd.n1853 163.367
R6948 gnd.n4947 gnd.n1853 163.367
R6949 gnd.n4947 gnd.n1841 163.367
R6950 gnd.n4960 gnd.n1841 163.367
R6951 gnd.n4960 gnd.n1838 163.367
R6952 gnd.n4965 gnd.n1838 163.367
R6953 gnd.n4965 gnd.n1839 163.367
R6954 gnd.n1839 gnd.n1822 163.367
R6955 gnd.n4989 gnd.n1822 163.367
R6956 gnd.n4989 gnd.n1820 163.367
R6957 gnd.n4993 gnd.n1820 163.367
R6958 gnd.n4993 gnd.n1813 163.367
R6959 gnd.n5009 gnd.n1813 163.367
R6960 gnd.n5009 gnd.n1811 163.367
R6961 gnd.n5013 gnd.n1811 163.367
R6962 gnd.n5013 gnd.n1798 163.367
R6963 gnd.n5036 gnd.n1798 163.367
R6964 gnd.n5036 gnd.n1796 163.367
R6965 gnd.n5040 gnd.n1796 163.367
R6966 gnd.n5040 gnd.n1787 163.367
R6967 gnd.n5049 gnd.n1787 163.367
R6968 gnd.n5049 gnd.n1785 163.367
R6969 gnd.n5053 gnd.n1785 163.367
R6970 gnd.n5053 gnd.n1775 163.367
R6971 gnd.n5067 gnd.n1775 163.367
R6972 gnd.n5067 gnd.n1773 163.367
R6973 gnd.n5071 gnd.n1773 163.367
R6974 gnd.n5071 gnd.n1760 163.367
R6975 gnd.n5083 gnd.n1760 163.367
R6976 gnd.n5083 gnd.n1757 163.367
R6977 gnd.n5088 gnd.n1757 163.367
R6978 gnd.n5088 gnd.n1758 163.367
R6979 gnd.n1758 gnd.n1740 163.367
R6980 gnd.n5111 gnd.n1740 163.367
R6981 gnd.n5111 gnd.n1738 163.367
R6982 gnd.n5115 gnd.n1738 163.367
R6983 gnd.n5115 gnd.n1730 163.367
R6984 gnd.n5130 gnd.n1730 163.367
R6985 gnd.n5130 gnd.n1728 163.367
R6986 gnd.n5134 gnd.n1728 163.367
R6987 gnd.n5134 gnd.n1715 163.367
R6988 gnd.n5154 gnd.n1715 163.367
R6989 gnd.n5154 gnd.n1713 163.367
R6990 gnd.n5158 gnd.n1713 163.367
R6991 gnd.n5158 gnd.n1705 163.367
R6992 gnd.n5167 gnd.n1705 163.367
R6993 gnd.n5167 gnd.n1702 163.367
R6994 gnd.n5173 gnd.n1702 163.367
R6995 gnd.n5173 gnd.n1703 163.367
R6996 gnd.n1703 gnd.n1692 163.367
R6997 gnd.n1692 gnd.n1680 163.367
R6998 gnd.n5194 gnd.n1680 163.367
R6999 gnd.n5194 gnd.n1678 163.367
R7000 gnd.n5198 gnd.n1678 163.367
R7001 gnd.n5198 gnd.n1669 163.367
R7002 gnd.n5212 gnd.n1669 163.367
R7003 gnd.n5212 gnd.n1667 163.367
R7004 gnd.n5216 gnd.n1667 163.367
R7005 gnd.n5216 gnd.n1652 163.367
R7006 gnd.n5227 gnd.n1652 163.367
R7007 gnd.n5227 gnd.n1650 163.367
R7008 gnd.n5231 gnd.n1650 163.367
R7009 gnd.n5231 gnd.n1638 163.367
R7010 gnd.n5252 gnd.n1638 163.367
R7011 gnd.n5252 gnd.n1639 163.367
R7012 gnd.n5248 gnd.n1639 163.367
R7013 gnd.n5248 gnd.n5247 163.367
R7014 gnd.n5247 gnd.n5246 163.367
R7015 gnd.n5246 gnd.n1642 163.367
R7016 gnd.n1642 gnd.n1539 163.367
R7017 gnd.n5402 gnd.n1539 163.367
R7018 gnd.n5402 gnd.n1540 163.367
R7019 gnd.n5398 gnd.n1540 163.367
R7020 gnd.n1560 gnd.n1559 156.462
R7021 gnd.n3531 gnd.n3499 153.042
R7022 gnd.n3595 gnd.n3594 152.079
R7023 gnd.n3563 gnd.n3562 152.079
R7024 gnd.n3531 gnd.n3530 152.079
R7025 gnd.n1100 gnd.n1099 152
R7026 gnd.n1101 gnd.n1090 152
R7027 gnd.n1103 gnd.n1102 152
R7028 gnd.n1105 gnd.n1088 152
R7029 gnd.n1107 gnd.n1106 152
R7030 gnd.n1558 gnd.n1542 152
R7031 gnd.n1550 gnd.n1543 152
R7032 gnd.n1549 gnd.n1548 152
R7033 gnd.n1547 gnd.n1544 152
R7034 gnd.n1545 gnd.t123 150.546
R7035 gnd.t36 gnd.n3573 147.661
R7036 gnd.t42 gnd.n3541 147.661
R7037 gnd.t180 gnd.n3509 147.661
R7038 gnd.t30 gnd.n3478 147.661
R7039 gnd.t38 gnd.n3446 147.661
R7040 gnd.t191 gnd.n3414 147.661
R7041 gnd.t40 gnd.n3382 147.661
R7042 gnd.t44 gnd.n3351 147.661
R7043 gnd.n5340 gnd.n5339 143.351
R7044 gnd.n1067 gnd.n1050 143.351
R7045 gnd.n5970 gnd.n1050 143.351
R7046 gnd.n1097 gnd.t87 130.484
R7047 gnd.n1106 gnd.t77 126.766
R7048 gnd.n1104 gnd.t132 126.766
R7049 gnd.n1090 gnd.t104 126.766
R7050 gnd.n1098 gnd.t160 126.766
R7051 gnd.n1546 gnd.t107 126.766
R7052 gnd.n1548 gnd.t126 126.766
R7053 gnd.n1557 gnd.t80 126.766
R7054 gnd.n1559 gnd.t148 126.766
R7055 gnd.n3590 gnd.n3589 104.615
R7056 gnd.n3589 gnd.n3567 104.615
R7057 gnd.n3582 gnd.n3567 104.615
R7058 gnd.n3582 gnd.n3581 104.615
R7059 gnd.n3581 gnd.n3571 104.615
R7060 gnd.n3574 gnd.n3571 104.615
R7061 gnd.n3558 gnd.n3557 104.615
R7062 gnd.n3557 gnd.n3535 104.615
R7063 gnd.n3550 gnd.n3535 104.615
R7064 gnd.n3550 gnd.n3549 104.615
R7065 gnd.n3549 gnd.n3539 104.615
R7066 gnd.n3542 gnd.n3539 104.615
R7067 gnd.n3526 gnd.n3525 104.615
R7068 gnd.n3525 gnd.n3503 104.615
R7069 gnd.n3518 gnd.n3503 104.615
R7070 gnd.n3518 gnd.n3517 104.615
R7071 gnd.n3517 gnd.n3507 104.615
R7072 gnd.n3510 gnd.n3507 104.615
R7073 gnd.n3495 gnd.n3494 104.615
R7074 gnd.n3494 gnd.n3472 104.615
R7075 gnd.n3487 gnd.n3472 104.615
R7076 gnd.n3487 gnd.n3486 104.615
R7077 gnd.n3486 gnd.n3476 104.615
R7078 gnd.n3479 gnd.n3476 104.615
R7079 gnd.n3463 gnd.n3462 104.615
R7080 gnd.n3462 gnd.n3440 104.615
R7081 gnd.n3455 gnd.n3440 104.615
R7082 gnd.n3455 gnd.n3454 104.615
R7083 gnd.n3454 gnd.n3444 104.615
R7084 gnd.n3447 gnd.n3444 104.615
R7085 gnd.n3431 gnd.n3430 104.615
R7086 gnd.n3430 gnd.n3408 104.615
R7087 gnd.n3423 gnd.n3408 104.615
R7088 gnd.n3423 gnd.n3422 104.615
R7089 gnd.n3422 gnd.n3412 104.615
R7090 gnd.n3415 gnd.n3412 104.615
R7091 gnd.n3399 gnd.n3398 104.615
R7092 gnd.n3398 gnd.n3376 104.615
R7093 gnd.n3391 gnd.n3376 104.615
R7094 gnd.n3391 gnd.n3390 104.615
R7095 gnd.n3390 gnd.n3380 104.615
R7096 gnd.n3383 gnd.n3380 104.615
R7097 gnd.n3368 gnd.n3367 104.615
R7098 gnd.n3367 gnd.n3345 104.615
R7099 gnd.n3360 gnd.n3345 104.615
R7100 gnd.n3360 gnd.n3359 104.615
R7101 gnd.n3359 gnd.n3349 104.615
R7102 gnd.n3352 gnd.n3349 104.615
R7103 gnd.n2742 gnd.t138 100.632
R7104 gnd.n2283 gnd.t171 100.632
R7105 gnd.n7182 gnd.n7181 99.6594
R7106 gnd.n7177 gnd.n248 99.6594
R7107 gnd.n7173 gnd.n247 99.6594
R7108 gnd.n7169 gnd.n246 99.6594
R7109 gnd.n7165 gnd.n245 99.6594
R7110 gnd.n7161 gnd.n244 99.6594
R7111 gnd.n7157 gnd.n243 99.6594
R7112 gnd.n7153 gnd.n242 99.6594
R7113 gnd.n7146 gnd.n241 99.6594
R7114 gnd.n7142 gnd.n240 99.6594
R7115 gnd.n7138 gnd.n239 99.6594
R7116 gnd.n7134 gnd.n238 99.6594
R7117 gnd.n7130 gnd.n237 99.6594
R7118 gnd.n7126 gnd.n236 99.6594
R7119 gnd.n7122 gnd.n235 99.6594
R7120 gnd.n7118 gnd.n234 99.6594
R7121 gnd.n7114 gnd.n233 99.6594
R7122 gnd.n7110 gnd.n232 99.6594
R7123 gnd.n7102 gnd.n231 99.6594
R7124 gnd.n7100 gnd.n230 99.6594
R7125 gnd.n7096 gnd.n229 99.6594
R7126 gnd.n7092 gnd.n228 99.6594
R7127 gnd.n7088 gnd.n227 99.6594
R7128 gnd.n7084 gnd.n226 99.6594
R7129 gnd.n7080 gnd.n225 99.6594
R7130 gnd.n7076 gnd.n224 99.6594
R7131 gnd.n7072 gnd.n223 99.6594
R7132 gnd.n7068 gnd.n222 99.6594
R7133 gnd.n7059 gnd.n221 99.6594
R7134 gnd.n5712 gnd.n5711 99.6594
R7135 gnd.n5706 gnd.n1289 99.6594
R7136 gnd.n5703 gnd.n1290 99.6594
R7137 gnd.n5699 gnd.n1291 99.6594
R7138 gnd.n5695 gnd.n1292 99.6594
R7139 gnd.n5691 gnd.n1293 99.6594
R7140 gnd.n5687 gnd.n1294 99.6594
R7141 gnd.n5683 gnd.n1295 99.6594
R7142 gnd.n5679 gnd.n1296 99.6594
R7143 gnd.n5674 gnd.n1297 99.6594
R7144 gnd.n5670 gnd.n1298 99.6594
R7145 gnd.n5666 gnd.n1299 99.6594
R7146 gnd.n5662 gnd.n1300 99.6594
R7147 gnd.n5657 gnd.n1302 99.6594
R7148 gnd.n5653 gnd.n1303 99.6594
R7149 gnd.n5649 gnd.n1304 99.6594
R7150 gnd.n5645 gnd.n1305 99.6594
R7151 gnd.n5641 gnd.n1306 99.6594
R7152 gnd.n5637 gnd.n1307 99.6594
R7153 gnd.n5633 gnd.n1308 99.6594
R7154 gnd.n5629 gnd.n1309 99.6594
R7155 gnd.n5625 gnd.n1310 99.6594
R7156 gnd.n5621 gnd.n1311 99.6594
R7157 gnd.n5617 gnd.n1312 99.6594
R7158 gnd.n5613 gnd.n1313 99.6594
R7159 gnd.n5609 gnd.n1314 99.6594
R7160 gnd.n5605 gnd.n1315 99.6594
R7161 gnd.n5601 gnd.n1316 99.6594
R7162 gnd.n6022 gnd.n6021 99.6594
R7163 gnd.n6017 gnd.n1017 99.6594
R7164 gnd.n6013 gnd.n1016 99.6594
R7165 gnd.n6009 gnd.n1015 99.6594
R7166 gnd.n6005 gnd.n1014 99.6594
R7167 gnd.n6001 gnd.n1013 99.6594
R7168 gnd.n5997 gnd.n1012 99.6594
R7169 gnd.n5993 gnd.n1011 99.6594
R7170 gnd.n5988 gnd.n1010 99.6594
R7171 gnd.n5984 gnd.n1009 99.6594
R7172 gnd.n5980 gnd.n1008 99.6594
R7173 gnd.n5976 gnd.n1007 99.6594
R7174 gnd.n4503 gnd.n1005 99.6594
R7175 gnd.n4507 gnd.n1004 99.6594
R7176 gnd.n4513 gnd.n1003 99.6594
R7177 gnd.n4517 gnd.n1002 99.6594
R7178 gnd.n4522 gnd.n1001 99.6594
R7179 gnd.n4526 gnd.n1000 99.6594
R7180 gnd.n4532 gnd.n999 99.6594
R7181 gnd.n4536 gnd.n998 99.6594
R7182 gnd.n4542 gnd.n997 99.6594
R7183 gnd.n4546 gnd.n996 99.6594
R7184 gnd.n4552 gnd.n995 99.6594
R7185 gnd.n4556 gnd.n994 99.6594
R7186 gnd.n4562 gnd.n993 99.6594
R7187 gnd.n4566 gnd.n992 99.6594
R7188 gnd.n4571 gnd.n991 99.6594
R7189 gnd.n4574 gnd.n990 99.6594
R7190 gnd.n4035 gnd.n4034 99.6594
R7191 gnd.n4029 gnd.n3723 99.6594
R7192 gnd.n4026 gnd.n3724 99.6594
R7193 gnd.n4022 gnd.n3725 99.6594
R7194 gnd.n4018 gnd.n3726 99.6594
R7195 gnd.n4014 gnd.n3727 99.6594
R7196 gnd.n4010 gnd.n3728 99.6594
R7197 gnd.n4006 gnd.n3729 99.6594
R7198 gnd.n4002 gnd.n3730 99.6594
R7199 gnd.n3997 gnd.n3731 99.6594
R7200 gnd.n3993 gnd.n3732 99.6594
R7201 gnd.n3989 gnd.n3733 99.6594
R7202 gnd.n3985 gnd.n3734 99.6594
R7203 gnd.n3981 gnd.n3735 99.6594
R7204 gnd.n3977 gnd.n3736 99.6594
R7205 gnd.n3973 gnd.n3737 99.6594
R7206 gnd.n3969 gnd.n3738 99.6594
R7207 gnd.n3965 gnd.n3739 99.6594
R7208 gnd.n3961 gnd.n3740 99.6594
R7209 gnd.n3957 gnd.n3741 99.6594
R7210 gnd.n3953 gnd.n3742 99.6594
R7211 gnd.n3949 gnd.n3743 99.6594
R7212 gnd.n3945 gnd.n3744 99.6594
R7213 gnd.n3941 gnd.n3745 99.6594
R7214 gnd.n3937 gnd.n3746 99.6594
R7215 gnd.n3933 gnd.n3747 99.6594
R7216 gnd.n3929 gnd.n3748 99.6594
R7217 gnd.n3925 gnd.n3749 99.6594
R7218 gnd.n4037 gnd.n2243 99.6594
R7219 gnd.n3713 gnd.n2266 99.6594
R7220 gnd.n3711 gnd.n2265 99.6594
R7221 gnd.n3707 gnd.n2264 99.6594
R7222 gnd.n3703 gnd.n2263 99.6594
R7223 gnd.n3699 gnd.n2262 99.6594
R7224 gnd.n3695 gnd.n2261 99.6594
R7225 gnd.n3691 gnd.n2260 99.6594
R7226 gnd.n3623 gnd.n2259 99.6594
R7227 gnd.n2954 gnd.n2685 99.6594
R7228 gnd.n2711 gnd.n2692 99.6594
R7229 gnd.n2713 gnd.n2693 99.6594
R7230 gnd.n2721 gnd.n2694 99.6594
R7231 gnd.n2723 gnd.n2695 99.6594
R7232 gnd.n2731 gnd.n2696 99.6594
R7233 gnd.n2733 gnd.n2697 99.6594
R7234 gnd.n2741 gnd.n2698 99.6594
R7235 gnd.n6983 gnd.n212 99.6594
R7236 gnd.n6987 gnd.n213 99.6594
R7237 gnd.n6993 gnd.n214 99.6594
R7238 gnd.n6997 gnd.n215 99.6594
R7239 gnd.n7003 gnd.n216 99.6594
R7240 gnd.n7007 gnd.n217 99.6594
R7241 gnd.n7013 gnd.n218 99.6594
R7242 gnd.n7017 gnd.n219 99.6594
R7243 gnd.n7023 gnd.n220 99.6594
R7244 gnd.n1401 gnd.n1317 99.6594
R7245 gnd.n1319 gnd.n1243 99.6594
R7246 gnd.n1320 gnd.n1250 99.6594
R7247 gnd.n1322 gnd.n1321 99.6594
R7248 gnd.n1324 gnd.n1259 99.6594
R7249 gnd.n1325 gnd.n1266 99.6594
R7250 gnd.n1327 gnd.n1326 99.6594
R7251 gnd.n1329 gnd.n1275 99.6594
R7252 gnd.n5714 gnd.n1284 99.6594
R7253 gnd.n3681 gnd.n2246 99.6594
R7254 gnd.n3677 gnd.n2247 99.6594
R7255 gnd.n3673 gnd.n2248 99.6594
R7256 gnd.n3669 gnd.n2249 99.6594
R7257 gnd.n3665 gnd.n2250 99.6594
R7258 gnd.n3661 gnd.n2251 99.6594
R7259 gnd.n3657 gnd.n2252 99.6594
R7260 gnd.n3653 gnd.n2253 99.6594
R7261 gnd.n3649 gnd.n2254 99.6594
R7262 gnd.n3645 gnd.n2255 99.6594
R7263 gnd.n3641 gnd.n2256 99.6594
R7264 gnd.n3637 gnd.n2257 99.6594
R7265 gnd.n3633 gnd.n2258 99.6594
R7266 gnd.n2869 gnd.n2868 99.6594
R7267 gnd.n2863 gnd.n2780 99.6594
R7268 gnd.n2860 gnd.n2781 99.6594
R7269 gnd.n2856 gnd.n2782 99.6594
R7270 gnd.n2852 gnd.n2783 99.6594
R7271 gnd.n2848 gnd.n2784 99.6594
R7272 gnd.n2844 gnd.n2785 99.6594
R7273 gnd.n2840 gnd.n2786 99.6594
R7274 gnd.n2836 gnd.n2787 99.6594
R7275 gnd.n2832 gnd.n2788 99.6594
R7276 gnd.n2828 gnd.n2789 99.6594
R7277 gnd.n2824 gnd.n2790 99.6594
R7278 gnd.n2871 gnd.n2779 99.6594
R7279 gnd.n4378 gnd.n980 99.6594
R7280 gnd.n4380 gnd.n981 99.6594
R7281 gnd.n4388 gnd.n982 99.6594
R7282 gnd.n4398 gnd.n983 99.6594
R7283 gnd.n4400 gnd.n984 99.6594
R7284 gnd.n4408 gnd.n985 99.6594
R7285 gnd.n4418 gnd.n986 99.6594
R7286 gnd.n4421 gnd.n987 99.6594
R7287 gnd.n4625 gnd.n988 99.6594
R7288 gnd.n3915 gnd.n3750 99.6594
R7289 gnd.n3912 gnd.n3751 99.6594
R7290 gnd.n3908 gnd.n3752 99.6594
R7291 gnd.n3904 gnd.n3753 99.6594
R7292 gnd.n3900 gnd.n3754 99.6594
R7293 gnd.n3896 gnd.n3755 99.6594
R7294 gnd.n3892 gnd.n3756 99.6594
R7295 gnd.n3888 gnd.n3757 99.6594
R7296 gnd.n3884 gnd.n3758 99.6594
R7297 gnd.n3913 gnd.n3750 99.6594
R7298 gnd.n3909 gnd.n3751 99.6594
R7299 gnd.n3905 gnd.n3752 99.6594
R7300 gnd.n3901 gnd.n3753 99.6594
R7301 gnd.n3897 gnd.n3754 99.6594
R7302 gnd.n3893 gnd.n3755 99.6594
R7303 gnd.n3889 gnd.n3756 99.6594
R7304 gnd.n3885 gnd.n3757 99.6594
R7305 gnd.n3840 gnd.n3758 99.6594
R7306 gnd.n4420 gnd.n988 99.6594
R7307 gnd.n4419 gnd.n987 99.6594
R7308 gnd.n4409 gnd.n986 99.6594
R7309 gnd.n4401 gnd.n985 99.6594
R7310 gnd.n4399 gnd.n984 99.6594
R7311 gnd.n4389 gnd.n983 99.6594
R7312 gnd.n4381 gnd.n982 99.6594
R7313 gnd.n4379 gnd.n981 99.6594
R7314 gnd.n4369 gnd.n980 99.6594
R7315 gnd.n2869 gnd.n2792 99.6594
R7316 gnd.n2861 gnd.n2780 99.6594
R7317 gnd.n2857 gnd.n2781 99.6594
R7318 gnd.n2853 gnd.n2782 99.6594
R7319 gnd.n2849 gnd.n2783 99.6594
R7320 gnd.n2845 gnd.n2784 99.6594
R7321 gnd.n2841 gnd.n2785 99.6594
R7322 gnd.n2837 gnd.n2786 99.6594
R7323 gnd.n2833 gnd.n2787 99.6594
R7324 gnd.n2829 gnd.n2788 99.6594
R7325 gnd.n2825 gnd.n2789 99.6594
R7326 gnd.n2821 gnd.n2790 99.6594
R7327 gnd.n2872 gnd.n2871 99.6594
R7328 gnd.n3636 gnd.n2258 99.6594
R7329 gnd.n3640 gnd.n2257 99.6594
R7330 gnd.n3644 gnd.n2256 99.6594
R7331 gnd.n3648 gnd.n2255 99.6594
R7332 gnd.n3652 gnd.n2254 99.6594
R7333 gnd.n3656 gnd.n2253 99.6594
R7334 gnd.n3660 gnd.n2252 99.6594
R7335 gnd.n3664 gnd.n2251 99.6594
R7336 gnd.n3668 gnd.n2250 99.6594
R7337 gnd.n3672 gnd.n2249 99.6594
R7338 gnd.n3676 gnd.n2248 99.6594
R7339 gnd.n3680 gnd.n2247 99.6594
R7340 gnd.n2287 gnd.n2246 99.6594
R7341 gnd.n1317 gnd.n1242 99.6594
R7342 gnd.n1319 gnd.n1318 99.6594
R7343 gnd.n1320 gnd.n1251 99.6594
R7344 gnd.n1322 gnd.n1258 99.6594
R7345 gnd.n1324 gnd.n1323 99.6594
R7346 gnd.n1325 gnd.n1267 99.6594
R7347 gnd.n1327 gnd.n1274 99.6594
R7348 gnd.n1329 gnd.n1328 99.6594
R7349 gnd.n5715 gnd.n5714 99.6594
R7350 gnd.n7016 gnd.n220 99.6594
R7351 gnd.n7014 gnd.n219 99.6594
R7352 gnd.n7006 gnd.n218 99.6594
R7353 gnd.n7004 gnd.n217 99.6594
R7354 gnd.n6996 gnd.n216 99.6594
R7355 gnd.n6994 gnd.n215 99.6594
R7356 gnd.n6986 gnd.n214 99.6594
R7357 gnd.n6984 gnd.n213 99.6594
R7358 gnd.n6978 gnd.n212 99.6594
R7359 gnd.n2955 gnd.n2954 99.6594
R7360 gnd.n2714 gnd.n2692 99.6594
R7361 gnd.n2720 gnd.n2693 99.6594
R7362 gnd.n2724 gnd.n2694 99.6594
R7363 gnd.n2730 gnd.n2695 99.6594
R7364 gnd.n2734 gnd.n2696 99.6594
R7365 gnd.n2740 gnd.n2697 99.6594
R7366 gnd.n2698 gnd.n2682 99.6594
R7367 gnd.n3690 gnd.n2259 99.6594
R7368 gnd.n3694 gnd.n2260 99.6594
R7369 gnd.n3698 gnd.n2261 99.6594
R7370 gnd.n3702 gnd.n2262 99.6594
R7371 gnd.n3706 gnd.n2263 99.6594
R7372 gnd.n3710 gnd.n2264 99.6594
R7373 gnd.n3714 gnd.n2265 99.6594
R7374 gnd.n2268 gnd.n2266 99.6594
R7375 gnd.n4035 gnd.n3761 99.6594
R7376 gnd.n4027 gnd.n3723 99.6594
R7377 gnd.n4023 gnd.n3724 99.6594
R7378 gnd.n4019 gnd.n3725 99.6594
R7379 gnd.n4015 gnd.n3726 99.6594
R7380 gnd.n4011 gnd.n3727 99.6594
R7381 gnd.n4007 gnd.n3728 99.6594
R7382 gnd.n4003 gnd.n3729 99.6594
R7383 gnd.n3998 gnd.n3730 99.6594
R7384 gnd.n3994 gnd.n3731 99.6594
R7385 gnd.n3990 gnd.n3732 99.6594
R7386 gnd.n3986 gnd.n3733 99.6594
R7387 gnd.n3982 gnd.n3734 99.6594
R7388 gnd.n3978 gnd.n3735 99.6594
R7389 gnd.n3974 gnd.n3736 99.6594
R7390 gnd.n3970 gnd.n3737 99.6594
R7391 gnd.n3966 gnd.n3738 99.6594
R7392 gnd.n3962 gnd.n3739 99.6594
R7393 gnd.n3958 gnd.n3740 99.6594
R7394 gnd.n3954 gnd.n3741 99.6594
R7395 gnd.n3950 gnd.n3742 99.6594
R7396 gnd.n3946 gnd.n3743 99.6594
R7397 gnd.n3942 gnd.n3744 99.6594
R7398 gnd.n3938 gnd.n3745 99.6594
R7399 gnd.n3934 gnd.n3746 99.6594
R7400 gnd.n3930 gnd.n3747 99.6594
R7401 gnd.n3926 gnd.n3748 99.6594
R7402 gnd.n3922 gnd.n3749 99.6594
R7403 gnd.n4038 gnd.n4037 99.6594
R7404 gnd.n4484 gnd.n990 99.6594
R7405 gnd.n4565 gnd.n991 99.6594
R7406 gnd.n4563 gnd.n992 99.6594
R7407 gnd.n4555 gnd.n993 99.6594
R7408 gnd.n4553 gnd.n994 99.6594
R7409 gnd.n4545 gnd.n995 99.6594
R7410 gnd.n4543 gnd.n996 99.6594
R7411 gnd.n4535 gnd.n997 99.6594
R7412 gnd.n4533 gnd.n998 99.6594
R7413 gnd.n4525 gnd.n999 99.6594
R7414 gnd.n4497 gnd.n1000 99.6594
R7415 gnd.n4516 gnd.n1001 99.6594
R7416 gnd.n4514 gnd.n1002 99.6594
R7417 gnd.n4506 gnd.n1003 99.6594
R7418 gnd.n4504 gnd.n1004 99.6594
R7419 gnd.n5975 gnd.n1006 99.6594
R7420 gnd.n5979 gnd.n1007 99.6594
R7421 gnd.n5983 gnd.n1008 99.6594
R7422 gnd.n5987 gnd.n1009 99.6594
R7423 gnd.n5992 gnd.n1010 99.6594
R7424 gnd.n5996 gnd.n1011 99.6594
R7425 gnd.n6000 gnd.n1012 99.6594
R7426 gnd.n6004 gnd.n1013 99.6594
R7427 gnd.n6008 gnd.n1014 99.6594
R7428 gnd.n6012 gnd.n1015 99.6594
R7429 gnd.n6016 gnd.n1016 99.6594
R7430 gnd.n1018 gnd.n1017 99.6594
R7431 gnd.n6022 gnd.n977 99.6594
R7432 gnd.n5712 gnd.n1332 99.6594
R7433 gnd.n5704 gnd.n1289 99.6594
R7434 gnd.n5700 gnd.n1290 99.6594
R7435 gnd.n5696 gnd.n1291 99.6594
R7436 gnd.n5692 gnd.n1292 99.6594
R7437 gnd.n5688 gnd.n1293 99.6594
R7438 gnd.n5684 gnd.n1294 99.6594
R7439 gnd.n5680 gnd.n1295 99.6594
R7440 gnd.n5675 gnd.n1296 99.6594
R7441 gnd.n5671 gnd.n1297 99.6594
R7442 gnd.n5667 gnd.n1298 99.6594
R7443 gnd.n5663 gnd.n1299 99.6594
R7444 gnd.n5658 gnd.n1301 99.6594
R7445 gnd.n5654 gnd.n1302 99.6594
R7446 gnd.n5650 gnd.n1303 99.6594
R7447 gnd.n5646 gnd.n1304 99.6594
R7448 gnd.n5642 gnd.n1305 99.6594
R7449 gnd.n5638 gnd.n1306 99.6594
R7450 gnd.n5634 gnd.n1307 99.6594
R7451 gnd.n5630 gnd.n1308 99.6594
R7452 gnd.n5626 gnd.n1309 99.6594
R7453 gnd.n5622 gnd.n1310 99.6594
R7454 gnd.n5618 gnd.n1311 99.6594
R7455 gnd.n5614 gnd.n1312 99.6594
R7456 gnd.n5610 gnd.n1313 99.6594
R7457 gnd.n5606 gnd.n1314 99.6594
R7458 gnd.n5602 gnd.n1315 99.6594
R7459 gnd.n5594 gnd.n1316 99.6594
R7460 gnd.n7067 gnd.n221 99.6594
R7461 gnd.n7071 gnd.n222 99.6594
R7462 gnd.n7075 gnd.n223 99.6594
R7463 gnd.n7079 gnd.n224 99.6594
R7464 gnd.n7083 gnd.n225 99.6594
R7465 gnd.n7087 gnd.n226 99.6594
R7466 gnd.n7091 gnd.n227 99.6594
R7467 gnd.n7095 gnd.n228 99.6594
R7468 gnd.n7099 gnd.n229 99.6594
R7469 gnd.n7103 gnd.n230 99.6594
R7470 gnd.n7109 gnd.n231 99.6594
R7471 gnd.n7113 gnd.n232 99.6594
R7472 gnd.n7117 gnd.n233 99.6594
R7473 gnd.n7121 gnd.n234 99.6594
R7474 gnd.n7125 gnd.n235 99.6594
R7475 gnd.n7129 gnd.n236 99.6594
R7476 gnd.n7133 gnd.n237 99.6594
R7477 gnd.n7137 gnd.n238 99.6594
R7478 gnd.n7141 gnd.n239 99.6594
R7479 gnd.n7145 gnd.n240 99.6594
R7480 gnd.n7152 gnd.n241 99.6594
R7481 gnd.n7156 gnd.n242 99.6594
R7482 gnd.n7160 gnd.n243 99.6594
R7483 gnd.n7164 gnd.n244 99.6594
R7484 gnd.n7168 gnd.n245 99.6594
R7485 gnd.n7172 gnd.n246 99.6594
R7486 gnd.n7176 gnd.n247 99.6594
R7487 gnd.n249 gnd.n248 99.6594
R7488 gnd.n7182 gnd.n210 99.6594
R7489 gnd.n4352 gnd.n2016 99.6594
R7490 gnd.n4356 gnd.n2017 99.6594
R7491 gnd.n4339 gnd.n2018 99.6594
R7492 gnd.n4364 gnd.n2019 99.6594
R7493 gnd.n4366 gnd.n2020 99.6594
R7494 gnd.n4373 gnd.n2021 99.6594
R7495 gnd.n4375 gnd.n2022 99.6594
R7496 gnd.n4385 gnd.n2023 99.6594
R7497 gnd.n4393 gnd.n2024 99.6594
R7498 gnd.n4395 gnd.n2025 99.6594
R7499 gnd.n4405 gnd.n2026 99.6594
R7500 gnd.n4413 gnd.n2027 99.6594
R7501 gnd.n4415 gnd.n2028 99.6594
R7502 gnd.n4427 gnd.n2029 99.6594
R7503 gnd.n4355 gnd.n2016 99.6594
R7504 gnd.n4338 gnd.n2017 99.6594
R7505 gnd.n4363 gnd.n2018 99.6594
R7506 gnd.n4365 gnd.n2019 99.6594
R7507 gnd.n4372 gnd.n2020 99.6594
R7508 gnd.n4374 gnd.n2021 99.6594
R7509 gnd.n4384 gnd.n2022 99.6594
R7510 gnd.n4392 gnd.n2023 99.6594
R7511 gnd.n4394 gnd.n2024 99.6594
R7512 gnd.n4404 gnd.n2025 99.6594
R7513 gnd.n4412 gnd.n2026 99.6594
R7514 gnd.n4414 gnd.n2027 99.6594
R7515 gnd.n4426 gnd.n2028 99.6594
R7516 gnd.n2030 gnd.n2029 99.6594
R7517 gnd.n1479 gnd.n1223 99.6594
R7518 gnd.n1481 gnd.n1228 99.6594
R7519 gnd.n1482 gnd.n1231 99.6594
R7520 gnd.n1484 gnd.n1233 99.6594
R7521 gnd.n1485 gnd.n1237 99.6594
R7522 gnd.n1487 gnd.n1486 99.6594
R7523 gnd.n1489 gnd.n1247 99.6594
R7524 gnd.n1490 gnd.n1254 99.6594
R7525 gnd.n1492 gnd.n1491 99.6594
R7526 gnd.n1494 gnd.n1263 99.6594
R7527 gnd.n1495 gnd.n1270 99.6594
R7528 gnd.n1497 gnd.n1496 99.6594
R7529 gnd.n1500 gnd.n1279 99.6594
R7530 gnd.n5461 gnd.n1478 99.6594
R7531 gnd.n1497 gnd.n1278 99.6594
R7532 gnd.n1495 gnd.n1271 99.6594
R7533 gnd.n1494 gnd.n1493 99.6594
R7534 gnd.n1492 gnd.n1262 99.6594
R7535 gnd.n1490 gnd.n1255 99.6594
R7536 gnd.n1489 gnd.n1488 99.6594
R7537 gnd.n1487 gnd.n1246 99.6594
R7538 gnd.n1485 gnd.n1238 99.6594
R7539 gnd.n1484 gnd.n1483 99.6594
R7540 gnd.n1482 gnd.n1232 99.6594
R7541 gnd.n1481 gnd.n1480 99.6594
R7542 gnd.n1479 gnd.n1227 99.6594
R7543 gnd.n5462 gnd.n5461 99.6594
R7544 gnd.n1500 gnd.n1499 99.6594
R7545 gnd.n4423 gnd.t86 98.63
R7546 gnd.n5716 gnd.t144 98.63
R7547 gnd.n306 gnd.t164 98.63
R7548 gnd.n286 gnd.t75 98.63
R7549 gnd.n7148 gnd.t121 98.63
R7550 gnd.n1352 gnd.t141 98.63
R7551 gnd.n1375 gnd.t131 98.63
R7552 gnd.n5596 gnd.t64 98.63
R7553 gnd.n6967 gnd.t115 98.63
R7554 gnd.n2034 gnd.t167 98.63
R7555 gnd.n3841 gnd.t153 98.63
R7556 gnd.n3780 gnd.t99 98.63
R7557 gnd.n3802 gnd.t96 98.63
R7558 gnd.n3823 gnd.t68 98.63
R7559 gnd.n1035 gnd.t158 98.63
R7560 gnd.n4482 gnd.t92 98.63
R7561 gnd.n4495 gnd.t118 98.63
R7562 gnd.n1280 gnd.t102 98.63
R7563 gnd.n1908 gnd.t147 96.6984
R7564 gnd.n1591 gnd.t112 96.6984
R7565 gnd.n5904 gnd.t72 96.6906
R7566 gnd.n1585 gnd.t155 96.6906
R7567 gnd.n6578 gnd.n6577 84.828
R7568 gnd.n6579 gnd.n6578 84.828
R7569 gnd.n6579 gnd.n514 84.828
R7570 gnd.n6587 gnd.n514 84.828
R7571 gnd.n6588 gnd.n6587 84.828
R7572 gnd.n6589 gnd.n6588 84.828
R7573 gnd.n6589 gnd.n508 84.828
R7574 gnd.n6597 gnd.n508 84.828
R7575 gnd.n6598 gnd.n6597 84.828
R7576 gnd.n6599 gnd.n6598 84.828
R7577 gnd.n6599 gnd.n502 84.828
R7578 gnd.n6607 gnd.n502 84.828
R7579 gnd.n6608 gnd.n6607 84.828
R7580 gnd.n6609 gnd.n6608 84.828
R7581 gnd.n6609 gnd.n496 84.828
R7582 gnd.n6617 gnd.n496 84.828
R7583 gnd.n6618 gnd.n6617 84.828
R7584 gnd.n6619 gnd.n6618 84.828
R7585 gnd.n6619 gnd.n490 84.828
R7586 gnd.n6627 gnd.n490 84.828
R7587 gnd.n6628 gnd.n6627 84.828
R7588 gnd.n6629 gnd.n6628 84.828
R7589 gnd.n6629 gnd.n484 84.828
R7590 gnd.n6637 gnd.n484 84.828
R7591 gnd.n6638 gnd.n6637 84.828
R7592 gnd.n6639 gnd.n6638 84.828
R7593 gnd.n6639 gnd.n478 84.828
R7594 gnd.n6647 gnd.n478 84.828
R7595 gnd.n6648 gnd.n6647 84.828
R7596 gnd.n6649 gnd.n6648 84.828
R7597 gnd.n6649 gnd.n472 84.828
R7598 gnd.n6657 gnd.n472 84.828
R7599 gnd.n6658 gnd.n6657 84.828
R7600 gnd.n6659 gnd.n6658 84.828
R7601 gnd.n6659 gnd.n466 84.828
R7602 gnd.n6667 gnd.n466 84.828
R7603 gnd.n6668 gnd.n6667 84.828
R7604 gnd.n6669 gnd.n6668 84.828
R7605 gnd.n6669 gnd.n460 84.828
R7606 gnd.n6677 gnd.n460 84.828
R7607 gnd.n6678 gnd.n6677 84.828
R7608 gnd.n6679 gnd.n6678 84.828
R7609 gnd.n6679 gnd.n454 84.828
R7610 gnd.n6687 gnd.n454 84.828
R7611 gnd.n6688 gnd.n6687 84.828
R7612 gnd.n6689 gnd.n6688 84.828
R7613 gnd.n6689 gnd.n448 84.828
R7614 gnd.n6697 gnd.n448 84.828
R7615 gnd.n6698 gnd.n6697 84.828
R7616 gnd.n6699 gnd.n6698 84.828
R7617 gnd.n6699 gnd.n442 84.828
R7618 gnd.n6707 gnd.n442 84.828
R7619 gnd.n6708 gnd.n6707 84.828
R7620 gnd.n6709 gnd.n6708 84.828
R7621 gnd.n6709 gnd.n436 84.828
R7622 gnd.n6717 gnd.n436 84.828
R7623 gnd.n6718 gnd.n6717 84.828
R7624 gnd.n6719 gnd.n6718 84.828
R7625 gnd.n6719 gnd.n430 84.828
R7626 gnd.n6727 gnd.n430 84.828
R7627 gnd.n6728 gnd.n6727 84.828
R7628 gnd.n6729 gnd.n6728 84.828
R7629 gnd.n6729 gnd.n424 84.828
R7630 gnd.n6737 gnd.n424 84.828
R7631 gnd.n6738 gnd.n6737 84.828
R7632 gnd.n6739 gnd.n6738 84.828
R7633 gnd.n6739 gnd.n418 84.828
R7634 gnd.n6747 gnd.n418 84.828
R7635 gnd.n6748 gnd.n6747 84.828
R7636 gnd.n6749 gnd.n6748 84.828
R7637 gnd.n6749 gnd.n412 84.828
R7638 gnd.n6757 gnd.n412 84.828
R7639 gnd.n6758 gnd.n6757 84.828
R7640 gnd.n6759 gnd.n6758 84.828
R7641 gnd.n6759 gnd.n406 84.828
R7642 gnd.n6767 gnd.n406 84.828
R7643 gnd.n6768 gnd.n6767 84.828
R7644 gnd.n6769 gnd.n6768 84.828
R7645 gnd.n6769 gnd.n400 84.828
R7646 gnd.n6777 gnd.n400 84.828
R7647 gnd.n6778 gnd.n6777 84.828
R7648 gnd.n6780 gnd.n6778 84.828
R7649 gnd.n6780 gnd.n6779 84.828
R7650 gnd.n1097 gnd.n1096 81.8399
R7651 gnd.n5660 gnd.n1362 77.1205
R7652 gnd.n5973 gnd.n5972 77.1205
R7653 gnd.n2743 gnd.t137 74.8376
R7654 gnd.n2284 gnd.t172 74.8376
R7655 gnd.n1909 gnd.t146 72.8438
R7656 gnd.n1592 gnd.t113 72.8438
R7657 gnd.n1098 gnd.n1091 72.8411
R7658 gnd.n1104 gnd.n1089 72.8411
R7659 gnd.n1557 gnd.n1556 72.8411
R7660 gnd.n4424 gnd.t85 72.836
R7661 gnd.n5905 gnd.t71 72.836
R7662 gnd.n1586 gnd.t156 72.836
R7663 gnd.n5717 gnd.t143 72.836
R7664 gnd.n307 gnd.t165 72.836
R7665 gnd.n287 gnd.t76 72.836
R7666 gnd.n7149 gnd.t122 72.836
R7667 gnd.n1353 gnd.t140 72.836
R7668 gnd.n1376 gnd.t130 72.836
R7669 gnd.n5597 gnd.t63 72.836
R7670 gnd.n6968 gnd.t116 72.836
R7671 gnd.n2035 gnd.t168 72.836
R7672 gnd.n3842 gnd.t152 72.836
R7673 gnd.n3781 gnd.t98 72.836
R7674 gnd.n3803 gnd.t95 72.836
R7675 gnd.n3824 gnd.t67 72.836
R7676 gnd.n1036 gnd.t159 72.836
R7677 gnd.n4483 gnd.t93 72.836
R7678 gnd.n4496 gnd.t119 72.836
R7679 gnd.n1281 gnd.t103 72.836
R7680 gnd.n5396 gnd.n5395 71.676
R7681 gnd.n5391 gnd.n1565 71.676
R7682 gnd.n5389 gnd.n5388 71.676
R7683 gnd.n5384 gnd.n1568 71.676
R7684 gnd.n5382 gnd.n5381 71.676
R7685 gnd.n5377 gnd.n1571 71.676
R7686 gnd.n5375 gnd.n5374 71.676
R7687 gnd.n5370 gnd.n1574 71.676
R7688 gnd.n5368 gnd.n5367 71.676
R7689 gnd.n5363 gnd.n1577 71.676
R7690 gnd.n5361 gnd.n5360 71.676
R7691 gnd.n5356 gnd.n1580 71.676
R7692 gnd.n5354 gnd.n5353 71.676
R7693 gnd.n5349 gnd.n1583 71.676
R7694 gnd.n5347 gnd.n5346 71.676
R7695 gnd.n5342 gnd.n1588 71.676
R7696 gnd.n5339 gnd.n5338 71.676
R7697 gnd.n5336 gnd.n5335 71.676
R7698 gnd.n5330 gnd.n1594 71.676
R7699 gnd.n5328 gnd.n5327 71.676
R7700 gnd.n5323 gnd.n1597 71.676
R7701 gnd.n5321 gnd.n5320 71.676
R7702 gnd.n5316 gnd.n1600 71.676
R7703 gnd.n5314 gnd.n5313 71.676
R7704 gnd.n5309 gnd.n1603 71.676
R7705 gnd.n5307 gnd.n5306 71.676
R7706 gnd.n5302 gnd.n1606 71.676
R7707 gnd.n5300 gnd.n5299 71.676
R7708 gnd.n5295 gnd.n1609 71.676
R7709 gnd.n5293 gnd.n5292 71.676
R7710 gnd.n5288 gnd.n1612 71.676
R7711 gnd.n5286 gnd.n5285 71.676
R7712 gnd.n5281 gnd.n1615 71.676
R7713 gnd.n5968 gnd.n5967 71.676
R7714 gnd.n5962 gnd.n1053 71.676
R7715 gnd.n5959 gnd.n1054 71.676
R7716 gnd.n5955 gnd.n1055 71.676
R7717 gnd.n5951 gnd.n1056 71.676
R7718 gnd.n5947 gnd.n1057 71.676
R7719 gnd.n5943 gnd.n1058 71.676
R7720 gnd.n5939 gnd.n1059 71.676
R7721 gnd.n5935 gnd.n1060 71.676
R7722 gnd.n5931 gnd.n1061 71.676
R7723 gnd.n5927 gnd.n1062 71.676
R7724 gnd.n5923 gnd.n1063 71.676
R7725 gnd.n5919 gnd.n1064 71.676
R7726 gnd.n5915 gnd.n1065 71.676
R7727 gnd.n5911 gnd.n1066 71.676
R7728 gnd.n5907 gnd.n1067 71.676
R7729 gnd.n1068 gnd.n1051 71.676
R7730 gnd.n1912 gnd.n1069 71.676
R7731 gnd.n1917 gnd.n1070 71.676
R7732 gnd.n1921 gnd.n1071 71.676
R7733 gnd.n1925 gnd.n1072 71.676
R7734 gnd.n1929 gnd.n1073 71.676
R7735 gnd.n1933 gnd.n1074 71.676
R7736 gnd.n1937 gnd.n1075 71.676
R7737 gnd.n1941 gnd.n1076 71.676
R7738 gnd.n1945 gnd.n1077 71.676
R7739 gnd.n1949 gnd.n1078 71.676
R7740 gnd.n1953 gnd.n1079 71.676
R7741 gnd.n1957 gnd.n1080 71.676
R7742 gnd.n1961 gnd.n1081 71.676
R7743 gnd.n1965 gnd.n1082 71.676
R7744 gnd.n1969 gnd.n1083 71.676
R7745 gnd.n5968 gnd.n1086 71.676
R7746 gnd.n5960 gnd.n1053 71.676
R7747 gnd.n5956 gnd.n1054 71.676
R7748 gnd.n5952 gnd.n1055 71.676
R7749 gnd.n5948 gnd.n1056 71.676
R7750 gnd.n5944 gnd.n1057 71.676
R7751 gnd.n5940 gnd.n1058 71.676
R7752 gnd.n5936 gnd.n1059 71.676
R7753 gnd.n5932 gnd.n1060 71.676
R7754 gnd.n5928 gnd.n1061 71.676
R7755 gnd.n5924 gnd.n1062 71.676
R7756 gnd.n5920 gnd.n1063 71.676
R7757 gnd.n5916 gnd.n1064 71.676
R7758 gnd.n5912 gnd.n1065 71.676
R7759 gnd.n5908 gnd.n1066 71.676
R7760 gnd.n5971 gnd.n5970 71.676
R7761 gnd.n1911 gnd.n1068 71.676
R7762 gnd.n1916 gnd.n1069 71.676
R7763 gnd.n1920 gnd.n1070 71.676
R7764 gnd.n1924 gnd.n1071 71.676
R7765 gnd.n1928 gnd.n1072 71.676
R7766 gnd.n1932 gnd.n1073 71.676
R7767 gnd.n1936 gnd.n1074 71.676
R7768 gnd.n1940 gnd.n1075 71.676
R7769 gnd.n1944 gnd.n1076 71.676
R7770 gnd.n1948 gnd.n1077 71.676
R7771 gnd.n1952 gnd.n1078 71.676
R7772 gnd.n1956 gnd.n1079 71.676
R7773 gnd.n1960 gnd.n1080 71.676
R7774 gnd.n1964 gnd.n1081 71.676
R7775 gnd.n1968 gnd.n1082 71.676
R7776 gnd.n1972 gnd.n1083 71.676
R7777 gnd.n1615 gnd.n1613 71.676
R7778 gnd.n5287 gnd.n5286 71.676
R7779 gnd.n1612 gnd.n1610 71.676
R7780 gnd.n5294 gnd.n5293 71.676
R7781 gnd.n1609 gnd.n1607 71.676
R7782 gnd.n5301 gnd.n5300 71.676
R7783 gnd.n1606 gnd.n1604 71.676
R7784 gnd.n5308 gnd.n5307 71.676
R7785 gnd.n1603 gnd.n1601 71.676
R7786 gnd.n5315 gnd.n5314 71.676
R7787 gnd.n1600 gnd.n1598 71.676
R7788 gnd.n5322 gnd.n5321 71.676
R7789 gnd.n1597 gnd.n1595 71.676
R7790 gnd.n5329 gnd.n5328 71.676
R7791 gnd.n1594 gnd.n1590 71.676
R7792 gnd.n5337 gnd.n5336 71.676
R7793 gnd.n5341 gnd.n5340 71.676
R7794 gnd.n1588 gnd.n1584 71.676
R7795 gnd.n5348 gnd.n5347 71.676
R7796 gnd.n1583 gnd.n1581 71.676
R7797 gnd.n5355 gnd.n5354 71.676
R7798 gnd.n1580 gnd.n1578 71.676
R7799 gnd.n5362 gnd.n5361 71.676
R7800 gnd.n1577 gnd.n1575 71.676
R7801 gnd.n5369 gnd.n5368 71.676
R7802 gnd.n1574 gnd.n1572 71.676
R7803 gnd.n5376 gnd.n5375 71.676
R7804 gnd.n1571 gnd.n1569 71.676
R7805 gnd.n5383 gnd.n5382 71.676
R7806 gnd.n1568 gnd.n1566 71.676
R7807 gnd.n5390 gnd.n5389 71.676
R7808 gnd.n1565 gnd.n1563 71.676
R7809 gnd.n5397 gnd.n5396 71.676
R7810 gnd.n8 gnd.t12 69.1507
R7811 gnd.n14 gnd.t27 68.4792
R7812 gnd.n13 gnd.t16 68.4792
R7813 gnd.n12 gnd.t25 68.4792
R7814 gnd.n11 gnd.t177 68.4792
R7815 gnd.n10 gnd.t361 68.4792
R7816 gnd.n9 gnd.t32 68.4792
R7817 gnd.n8 gnd.t51 68.4792
R7818 gnd.n2870 gnd.n2774 64.369
R7819 gnd.n1914 gnd.n1909 59.5399
R7820 gnd.n5332 gnd.n1592 59.5399
R7821 gnd.n5906 gnd.n5905 59.5399
R7822 gnd.n1587 gnd.n1586 59.5399
R7823 gnd.n5903 gnd.n1107 59.1804
R7824 gnd.n4036 gnd.n2234 57.3586
R7825 gnd.n7183 gnd.n204 57.3586
R7826 gnd.n2525 gnd.t274 56.407
R7827 gnd.n2478 gnd.t336 56.407
R7828 gnd.n2493 gnd.t222 56.407
R7829 gnd.n2509 gnd.t323 56.407
R7830 gnd.n64 gnd.t239 56.407
R7831 gnd.n17 gnd.t229 56.407
R7832 gnd.n32 gnd.t352 56.407
R7833 gnd.n48 gnd.t289 56.407
R7834 gnd.n2538 gnd.t257 55.8337
R7835 gnd.n2491 gnd.t346 55.8337
R7836 gnd.n2506 gnd.t316 55.8337
R7837 gnd.n2522 gnd.t300 55.8337
R7838 gnd.n77 gnd.t197 55.8337
R7839 gnd.n30 gnd.t244 55.8337
R7840 gnd.n45 gnd.t305 55.8337
R7841 gnd.n61 gnd.t268 55.8337
R7842 gnd.n1095 gnd.n1094 54.358
R7843 gnd.n1554 gnd.n1553 54.358
R7844 gnd.n2525 gnd.n2524 53.0052
R7845 gnd.n2527 gnd.n2526 53.0052
R7846 gnd.n2529 gnd.n2528 53.0052
R7847 gnd.n2531 gnd.n2530 53.0052
R7848 gnd.n2533 gnd.n2532 53.0052
R7849 gnd.n2535 gnd.n2534 53.0052
R7850 gnd.n2537 gnd.n2536 53.0052
R7851 gnd.n2478 gnd.n2477 53.0052
R7852 gnd.n2480 gnd.n2479 53.0052
R7853 gnd.n2482 gnd.n2481 53.0052
R7854 gnd.n2484 gnd.n2483 53.0052
R7855 gnd.n2486 gnd.n2485 53.0052
R7856 gnd.n2488 gnd.n2487 53.0052
R7857 gnd.n2490 gnd.n2489 53.0052
R7858 gnd.n2493 gnd.n2492 53.0052
R7859 gnd.n2495 gnd.n2494 53.0052
R7860 gnd.n2497 gnd.n2496 53.0052
R7861 gnd.n2499 gnd.n2498 53.0052
R7862 gnd.n2501 gnd.n2500 53.0052
R7863 gnd.n2503 gnd.n2502 53.0052
R7864 gnd.n2505 gnd.n2504 53.0052
R7865 gnd.n2509 gnd.n2508 53.0052
R7866 gnd.n2511 gnd.n2510 53.0052
R7867 gnd.n2513 gnd.n2512 53.0052
R7868 gnd.n2515 gnd.n2514 53.0052
R7869 gnd.n2517 gnd.n2516 53.0052
R7870 gnd.n2519 gnd.n2518 53.0052
R7871 gnd.n2521 gnd.n2520 53.0052
R7872 gnd.n76 gnd.n75 53.0052
R7873 gnd.n74 gnd.n73 53.0052
R7874 gnd.n72 gnd.n71 53.0052
R7875 gnd.n70 gnd.n69 53.0052
R7876 gnd.n68 gnd.n67 53.0052
R7877 gnd.n66 gnd.n65 53.0052
R7878 gnd.n64 gnd.n63 53.0052
R7879 gnd.n29 gnd.n28 53.0052
R7880 gnd.n27 gnd.n26 53.0052
R7881 gnd.n25 gnd.n24 53.0052
R7882 gnd.n23 gnd.n22 53.0052
R7883 gnd.n21 gnd.n20 53.0052
R7884 gnd.n19 gnd.n18 53.0052
R7885 gnd.n17 gnd.n16 53.0052
R7886 gnd.n44 gnd.n43 53.0052
R7887 gnd.n42 gnd.n41 53.0052
R7888 gnd.n40 gnd.n39 53.0052
R7889 gnd.n38 gnd.n37 53.0052
R7890 gnd.n36 gnd.n35 53.0052
R7891 gnd.n34 gnd.n33 53.0052
R7892 gnd.n32 gnd.n31 53.0052
R7893 gnd.n60 gnd.n59 53.0052
R7894 gnd.n58 gnd.n57 53.0052
R7895 gnd.n56 gnd.n55 53.0052
R7896 gnd.n54 gnd.n53 53.0052
R7897 gnd.n52 gnd.n51 53.0052
R7898 gnd.n50 gnd.n49 53.0052
R7899 gnd.n48 gnd.n47 53.0052
R7900 gnd.n1545 gnd.n1544 52.4801
R7901 gnd.n3574 gnd.t36 52.3082
R7902 gnd.n3542 gnd.t42 52.3082
R7903 gnd.n3510 gnd.t180 52.3082
R7904 gnd.n3479 gnd.t30 52.3082
R7905 gnd.n3447 gnd.t38 52.3082
R7906 gnd.n3415 gnd.t191 52.3082
R7907 gnd.n3383 gnd.t40 52.3082
R7908 gnd.n3352 gnd.t44 52.3082
R7909 gnd.n3404 gnd.n3372 51.4173
R7910 gnd.n6779 gnd.n157 50.897
R7911 gnd.n3468 gnd.n3467 50.455
R7912 gnd.n3436 gnd.n3435 50.455
R7913 gnd.n3404 gnd.n3403 50.455
R7914 gnd.n2817 gnd.n2816 45.1884
R7915 gnd.n2310 gnd.n2309 45.1884
R7916 gnd.n1561 gnd.n1560 44.3322
R7917 gnd.n1098 gnd.n1097 44.3189
R7918 gnd.n4425 gnd.n4424 42.2793
R7919 gnd.n5718 gnd.n5717 42.2793
R7920 gnd.n7066 gnd.n307 42.2793
R7921 gnd.n7108 gnd.n287 42.2793
R7922 gnd.n7150 gnd.n7149 42.2793
R7923 gnd.n5677 gnd.n1353 42.2793
R7924 gnd.n5640 gnd.n1376 42.2793
R7925 gnd.n5600 gnd.n5597 42.2793
R7926 gnd.n6969 gnd.n6968 42.2793
R7927 gnd.n2818 gnd.n2817 42.2793
R7928 gnd.n2311 gnd.n2310 42.2793
R7929 gnd.n2744 gnd.n2743 42.2793
R7930 gnd.n3689 gnd.n2284 42.2793
R7931 gnd.n2036 gnd.n2035 42.2793
R7932 gnd.n3843 gnd.n3842 42.2793
R7933 gnd.n4000 gnd.n3781 42.2793
R7934 gnd.n3960 gnd.n3803 42.2793
R7935 gnd.n3921 gnd.n3824 42.2793
R7936 gnd.n5990 gnd.n1036 42.2793
R7937 gnd.n4573 gnd.n4483 42.2793
R7938 gnd.n4524 gnd.n4496 42.2793
R7939 gnd.n1282 gnd.n1281 42.2793
R7940 gnd.n1096 gnd.n1095 41.6274
R7941 gnd.n1555 gnd.n1554 41.6274
R7942 gnd.n1105 gnd.n1104 40.8975
R7943 gnd.n1558 gnd.n1557 40.8975
R7944 gnd.n1104 gnd.n1103 35.055
R7945 gnd.n1099 gnd.n1098 35.055
R7946 gnd.n1547 gnd.n1546 35.055
R7947 gnd.n1557 gnd.n1543 35.055
R7948 gnd.n6248 gnd.n6247 31.9912
R7949 gnd.n6247 gnd.n6246 31.9912
R7950 gnd.n6246 gnd.n717 31.9912
R7951 gnd.n6240 gnd.n717 31.9912
R7952 gnd.n6240 gnd.n6239 31.9912
R7953 gnd.n6239 gnd.n6238 31.9912
R7954 gnd.n6238 gnd.n724 31.9912
R7955 gnd.n6232 gnd.n724 31.9912
R7956 gnd.n6232 gnd.n6231 31.9912
R7957 gnd.n6231 gnd.n6230 31.9912
R7958 gnd.n6230 gnd.n732 31.9912
R7959 gnd.n6224 gnd.n732 31.9912
R7960 gnd.n6224 gnd.n6223 31.9912
R7961 gnd.n6223 gnd.n6222 31.9912
R7962 gnd.n6222 gnd.n740 31.9912
R7963 gnd.n6216 gnd.n740 31.9912
R7964 gnd.n6216 gnd.n6215 31.9912
R7965 gnd.n6215 gnd.n6214 31.9912
R7966 gnd.n6214 gnd.n748 31.9912
R7967 gnd.n6208 gnd.n748 31.9912
R7968 gnd.n6208 gnd.n6207 31.9912
R7969 gnd.n6207 gnd.n6206 31.9912
R7970 gnd.n6206 gnd.n756 31.9912
R7971 gnd.n6200 gnd.n756 31.9912
R7972 gnd.n6200 gnd.n6199 31.9912
R7973 gnd.n6199 gnd.n6198 31.9912
R7974 gnd.n6198 gnd.n764 31.9912
R7975 gnd.n6192 gnd.n764 31.9912
R7976 gnd.n6192 gnd.n6191 31.9912
R7977 gnd.n6191 gnd.n6190 31.9912
R7978 gnd.n6190 gnd.n772 31.9912
R7979 gnd.n6184 gnd.n772 31.9912
R7980 gnd.n6184 gnd.n6183 31.9912
R7981 gnd.n6183 gnd.n6182 31.9912
R7982 gnd.n6182 gnd.n780 31.9912
R7983 gnd.n6176 gnd.n780 31.9912
R7984 gnd.n6176 gnd.n6175 31.9912
R7985 gnd.n6175 gnd.n6174 31.9912
R7986 gnd.n6174 gnd.n788 31.9912
R7987 gnd.n6168 gnd.n788 31.9912
R7988 gnd.n6168 gnd.n6167 31.9912
R7989 gnd.n6167 gnd.n6166 31.9912
R7990 gnd.n6166 gnd.n796 31.9912
R7991 gnd.n6160 gnd.n796 31.9912
R7992 gnd.n6160 gnd.n6159 31.9912
R7993 gnd.n6159 gnd.n6158 31.9912
R7994 gnd.n6158 gnd.n804 31.9912
R7995 gnd.n6152 gnd.n804 31.9912
R7996 gnd.n6152 gnd.n6151 31.9912
R7997 gnd.n6151 gnd.n6150 31.9912
R7998 gnd.n6150 gnd.n812 31.9912
R7999 gnd.n6144 gnd.n812 31.9912
R8000 gnd.n6144 gnd.n6143 31.9912
R8001 gnd.n6143 gnd.n6142 31.9912
R8002 gnd.n6142 gnd.n820 31.9912
R8003 gnd.n6136 gnd.n820 31.9912
R8004 gnd.n6136 gnd.n6135 31.9912
R8005 gnd.n6135 gnd.n6134 31.9912
R8006 gnd.n6134 gnd.n828 31.9912
R8007 gnd.n6128 gnd.n828 31.9912
R8008 gnd.n6128 gnd.n6127 31.9912
R8009 gnd.n6127 gnd.n6126 31.9912
R8010 gnd.n6126 gnd.n836 31.9912
R8011 gnd.n6120 gnd.n836 31.9912
R8012 gnd.n6120 gnd.n6119 31.9912
R8013 gnd.n6119 gnd.n6118 31.9912
R8014 gnd.n6118 gnd.n844 31.9912
R8015 gnd.n6112 gnd.n844 31.9912
R8016 gnd.n6112 gnd.n6111 31.9912
R8017 gnd.n6111 gnd.n6110 31.9912
R8018 gnd.n6110 gnd.n852 31.9912
R8019 gnd.n6104 gnd.n852 31.9912
R8020 gnd.n6104 gnd.n6103 31.9912
R8021 gnd.n6103 gnd.n6102 31.9912
R8022 gnd.n6102 gnd.n860 31.9912
R8023 gnd.n6096 gnd.n860 31.9912
R8024 gnd.n6096 gnd.n6095 31.9912
R8025 gnd.n6095 gnd.n6094 31.9912
R8026 gnd.n6094 gnd.n868 31.9912
R8027 gnd.n6088 gnd.n868 31.9912
R8028 gnd.n6088 gnd.n6087 31.9912
R8029 gnd.n6087 gnd.n6086 31.9912
R8030 gnd.n6086 gnd.n876 31.9912
R8031 gnd.n2880 gnd.n2774 31.8661
R8032 gnd.n2880 gnd.n2879 31.8661
R8033 gnd.n2888 gnd.n2763 31.8661
R8034 gnd.n2896 gnd.n2763 31.8661
R8035 gnd.n2896 gnd.n2757 31.8661
R8036 gnd.n2904 gnd.n2757 31.8661
R8037 gnd.n2904 gnd.n2750 31.8661
R8038 gnd.n2942 gnd.n2750 31.8661
R8039 gnd.n2952 gnd.n2683 31.8661
R8040 gnd.n4049 gnd.n2234 31.8661
R8041 gnd.n4057 gnd.n2226 31.8661
R8042 gnd.n4057 gnd.n2215 31.8661
R8043 gnd.n4069 gnd.n2215 31.8661
R8044 gnd.n4069 gnd.n2218 31.8661
R8045 gnd.n4077 gnd.n2198 31.8661
R8046 gnd.n4089 gnd.n2198 31.8661
R8047 gnd.n4097 gnd.n2190 31.8661
R8048 gnd.n4113 gnd.n2178 31.8661
R8049 gnd.n4113 gnd.n2181 31.8661
R8050 gnd.n4123 gnd.n2164 31.8661
R8051 gnd.n4133 gnd.n2164 31.8661
R8052 gnd.n4148 gnd.n2155 31.8661
R8053 gnd.n4158 gnd.n2139 31.8661
R8054 gnd.n4168 gnd.n2139 31.8661
R8055 gnd.n4183 gnd.n2120 31.8661
R8056 gnd.n4193 gnd.n2120 31.8661
R8057 gnd.n4215 gnd.n2113 31.8661
R8058 gnd.n4226 gnd.n2096 31.8661
R8059 gnd.n4234 gnd.n2096 31.8661
R8060 gnd.n4253 gnd.n2083 31.8661
R8061 gnd.n4253 gnd.n2086 31.8661
R8062 gnd.n4262 gnd.n883 31.8661
R8063 gnd.n4622 gnd.n978 31.8661
R8064 gnd.n2015 gnd.n989 31.8661
R8065 gnd.n4633 gnd.n2015 31.8661
R8066 gnd.n4634 gnd.n4633 31.8661
R8067 gnd.n4634 gnd.n2008 31.8661
R8068 gnd.n4642 gnd.n2008 31.8661
R8069 gnd.n4667 gnd.n1999 31.8661
R8070 gnd.n4667 gnd.n1990 31.8661
R8071 gnd.n4684 gnd.n1990 31.8661
R8072 gnd.n4684 gnd.n1991 31.8661
R8073 gnd.n5420 gnd.n1515 31.8661
R8074 gnd.n5431 gnd.n1515 31.8661
R8075 gnd.n5431 gnd.n1508 31.8661
R8076 gnd.n5439 gnd.n1508 31.8661
R8077 gnd.n5781 gnd.n1219 31.8661
R8078 gnd.n5781 gnd.n1221 31.8661
R8079 gnd.n5460 gnd.n1221 31.8661
R8080 gnd.n5460 gnd.n1501 31.8661
R8081 gnd.n1501 gnd.n1288 31.8661
R8082 gnd.n1398 gnd.n1330 31.8661
R8083 gnd.n6841 gnd.n354 31.8661
R8084 gnd.n6851 gnd.n336 31.8661
R8085 gnd.n6865 gnd.n336 31.8661
R8086 gnd.n6874 gnd.n319 31.8661
R8087 gnd.n6885 gnd.n319 31.8661
R8088 gnd.n6893 gnd.n313 31.8661
R8089 gnd.n7263 gnd.n86 31.8661
R8090 gnd.n7257 gnd.n86 31.8661
R8091 gnd.n7251 gnd.n106 31.8661
R8092 gnd.n7251 gnd.n109 31.8661
R8093 gnd.n7245 gnd.n119 31.8661
R8094 gnd.n7239 gnd.n128 31.8661
R8095 gnd.n7233 gnd.n128 31.8661
R8096 gnd.n7227 gnd.n144 31.8661
R8097 gnd.n7227 gnd.n147 31.8661
R8098 gnd.n7215 gnd.n166 31.8661
R8099 gnd.n7209 gnd.n166 31.8661
R8100 gnd.n7203 gnd.n182 31.8661
R8101 gnd.n7203 gnd.n185 31.8661
R8102 gnd.n7197 gnd.n185 31.8661
R8103 gnd.n7197 gnd.n195 31.8661
R8104 gnd.n7191 gnd.n204 31.8661
R8105 gnd.n5282 gnd.n1614 30.4395
R8106 gnd.n1975 gnd.n1971 30.4395
R8107 gnd.n3722 gnd.n2244 29.9541
R8108 gnd.n4097 gnd.t282 27.7236
R8109 gnd.n7221 gnd.t248 27.7236
R8110 gnd.n2319 gnd.n2244 27.4049
R8111 gnd.n6023 gnd.n989 27.4049
R8112 gnd.n5713 gnd.n1288 27.4049
R8113 gnd.n2155 gnd.t260 27.0862
R8114 gnd.n4262 gnd.t277 27.0862
R8115 gnd.n354 gnd.t245 27.0862
R8116 gnd.n7245 gnd.t206 27.0862
R8117 gnd.t275 gnd.n2113 26.4489
R8118 gnd.n4215 gnd.t231 26.4489
R8119 gnd.t204 gnd.n313 26.4489
R8120 gnd.n6893 gnd.t240 26.4489
R8121 gnd.n4148 gnd.t213 25.8116
R8122 gnd.n5969 gnd.n1084 25.8116
R8123 gnd.n5412 gnd.n1528 25.8116
R8124 gnd.t258 gnd.n119 25.8116
R8125 gnd.n4424 gnd.n4423 25.7944
R8126 gnd.n5717 gnd.n5716 25.7944
R8127 gnd.n307 gnd.n306 25.7944
R8128 gnd.n287 gnd.n286 25.7944
R8129 gnd.n7149 gnd.n7148 25.7944
R8130 gnd.n1353 gnd.n1352 25.7944
R8131 gnd.n1376 gnd.n1375 25.7944
R8132 gnd.n5597 gnd.n5596 25.7944
R8133 gnd.n6968 gnd.n6967 25.7944
R8134 gnd.n2743 gnd.n2742 25.7944
R8135 gnd.n2284 gnd.n2283 25.7944
R8136 gnd.n2035 gnd.n2034 25.7944
R8137 gnd.n3842 gnd.n3841 25.7944
R8138 gnd.n3781 gnd.n3780 25.7944
R8139 gnd.n3803 gnd.n3802 25.7944
R8140 gnd.n3824 gnd.n3823 25.7944
R8141 gnd.n1036 gnd.n1035 25.7944
R8142 gnd.n4483 gnd.n4482 25.7944
R8143 gnd.n4496 gnd.n4495 25.7944
R8144 gnd.n1281 gnd.n1280 25.7944
R8145 gnd.t198 gnd.n2190 25.1743
R8146 gnd.n7041 gnd.t215 25.1743
R8147 gnd.n2964 gnd.n2684 24.8557
R8148 gnd.n2974 gnd.n2667 24.8557
R8149 gnd.n2670 gnd.n2658 24.8557
R8150 gnd.n2995 gnd.n2659 24.8557
R8151 gnd.n3005 gnd.n2639 24.8557
R8152 gnd.n3015 gnd.n3014 24.8557
R8153 gnd.n2625 gnd.n2623 24.8557
R8154 gnd.n3046 gnd.n3045 24.8557
R8155 gnd.n3061 gnd.n2608 24.8557
R8156 gnd.n3115 gnd.n2547 24.8557
R8157 gnd.n3071 gnd.n2548 24.8557
R8158 gnd.n3108 gnd.n2559 24.8557
R8159 gnd.n2597 gnd.n2596 24.8557
R8160 gnd.n3102 gnd.n3101 24.8557
R8161 gnd.n2583 gnd.n2570 24.8557
R8162 gnd.n3141 gnd.n3140 24.8557
R8163 gnd.n3151 gnd.n2463 24.8557
R8164 gnd.n3163 gnd.n2455 24.8557
R8165 gnd.n3162 gnd.n2443 24.8557
R8166 gnd.n3181 gnd.n3180 24.8557
R8167 gnd.n3191 gnd.n2436 24.8557
R8168 gnd.n3202 gnd.n2424 24.8557
R8169 gnd.n3226 gnd.n3225 24.8557
R8170 gnd.n3237 gnd.n2407 24.8557
R8171 gnd.n3236 gnd.n2409 24.8557
R8172 gnd.n3248 gnd.n2400 24.8557
R8173 gnd.n3266 gnd.n3265 24.8557
R8174 gnd.n2391 gnd.n2380 24.8557
R8175 gnd.n3287 gnd.n2368 24.8557
R8176 gnd.n3315 gnd.n3314 24.8557
R8177 gnd.n3326 gnd.n2353 24.8557
R8178 gnd.n3337 gnd.n2346 24.8557
R8179 gnd.n3336 gnd.n2334 24.8557
R8180 gnd.n3609 gnd.n3608 24.8557
R8181 gnd.n3631 gnd.n2318 24.8557
R8182 gnd.n1909 gnd.n1908 23.855
R8183 gnd.n1592 gnd.n1591 23.855
R8184 gnd.n5905 gnd.n5904 23.855
R8185 gnd.n1586 gnd.n1585 23.855
R8186 gnd.n2985 gnd.t43 23.2624
R8187 gnd.n2686 gnd.t136 22.6251
R8188 gnd.n4049 gnd.t66 22.6251
R8189 gnd.n7191 gnd.t74 22.6251
R8190 gnd.n6080 gnd.t226 21.6691
R8191 gnd.n5899 gnd.n5898 21.6691
R8192 gnd.n4890 gnd.n1890 21.6691
R8193 gnd.n4917 gnd.n1873 21.6691
R8194 gnd.n4942 gnd.n1857 21.6691
R8195 gnd.n4966 gnd.n1837 21.6691
R8196 gnd.n4988 gnd.n4987 21.6691
R8197 gnd.n5008 gnd.n1814 21.6691
R8198 gnd.n5014 gnd.n1810 21.6691
R8199 gnd.n5041 gnd.n1792 21.6691
R8200 gnd.n5066 gnd.n1776 21.6691
R8201 gnd.n5066 gnd.n1769 21.6691
R8202 gnd.n5089 gnd.n1756 21.6691
R8203 gnd.n5110 gnd.n5109 21.6691
R8204 gnd.n5129 gnd.n1731 21.6691
R8205 gnd.n5135 gnd.n1727 21.6691
R8206 gnd.n5159 gnd.n1710 21.6691
R8207 gnd.n5182 gnd.n1691 21.6691
R8208 gnd.n5211 gnd.n1663 21.6691
R8209 gnd.n5226 gnd.n1653 21.6691
R8210 gnd.n5245 gnd.n1618 21.6691
R8211 gnd.n5403 gnd.n1538 21.6691
R8212 gnd.t202 gnd.n351 21.6691
R8213 gnd.t29 gnd.n2691 21.3504
R8214 gnd.n6079 gnd.n886 21.0318
R8215 gnd.n4271 gnd.n896 21.0318
R8216 gnd.n4290 gnd.n907 21.0318
R8217 gnd.n6067 gnd.n910 21.0318
R8218 gnd.n6061 gnd.n921 21.0318
R8219 gnd.n4316 gnd.n4315 21.0318
R8220 gnd.n6055 gnd.n930 21.0318
R8221 gnd.n4324 gnd.n938 21.0318
R8222 gnd.n4596 gnd.n947 21.0318
R8223 gnd.n6043 gnd.n950 21.0318
R8224 gnd.n4331 gnd.n958 21.0318
R8225 gnd.n6037 gnd.n961 21.0318
R8226 gnd.n6031 gnd.n971 21.0318
R8227 gnd.n4623 gnd.n4622 21.0318
R8228 gnd.n5592 gnd.n1398 21.0318
R8229 gnd.n5525 gnd.n1400 21.0318
R8230 gnd.n5480 gnd.n1410 21.0318
R8231 gnd.n5580 gnd.n1422 21.0318
R8232 gnd.n5484 gnd.n1425 21.0318
R8233 gnd.n5574 gnd.n1432 21.0318
R8234 gnd.n5568 gnd.n1443 21.0318
R8235 gnd.n5493 gnd.n1446 21.0318
R8236 gnd.n5562 gnd.n1453 21.0318
R8237 gnd.n5554 gnd.n1456 21.0318
R8238 gnd.n6807 gnd.n379 21.0318
R8239 gnd.n6794 gnd.n382 21.0318
R8240 gnd.n6800 gnd.n371 21.0318
R8241 gnd.n6826 gnd.n363 21.0318
R8242 gnd.t19 gnd.n2381 20.7131
R8243 gnd.t362 gnd.n1052 20.7131
R8244 gnd.n1527 gnd.t26 20.7131
R8245 gnd.n1973 gnd.n1110 20.3945
R8246 gnd.t161 gnd.n1899 20.3945
R8247 gnd.n4930 gnd.n1862 20.3945
R8248 gnd.n4948 gnd.n1852 20.3945
R8249 gnd.n5054 gnd.n1783 20.3945
R8250 gnd.n5072 gnd.n1772 20.3945
R8251 gnd.n5174 gnd.n1699 20.3945
R8252 gnd.n5193 gnd.n5192 20.3945
R8253 gnd.t184 gnd.n2416 20.0758
R8254 gnd.n1093 gnd.t134 19.8005
R8255 gnd.n1093 gnd.t106 19.8005
R8256 gnd.n1092 gnd.t162 19.8005
R8257 gnd.n1092 gnd.t89 19.8005
R8258 gnd.n1552 gnd.t109 19.8005
R8259 gnd.n1552 gnd.t128 19.8005
R8260 gnd.n1551 gnd.t82 19.8005
R8261 gnd.n1551 gnd.t150 19.8005
R8262 gnd.n1089 gnd.n1088 19.5087
R8263 gnd.n1102 gnd.n1089 19.5087
R8264 gnd.n1100 gnd.n1091 19.5087
R8265 gnd.n1556 gnd.n1550 19.5087
R8266 gnd.n3152 gnd.t45 19.4385
R8267 gnd.n4644 gnd.n2006 19.3944
R8268 gnd.n4644 gnd.n2003 19.3944
R8269 gnd.n4665 gnd.n2003 19.3944
R8270 gnd.n4665 gnd.n2004 19.3944
R8271 gnd.n4661 gnd.n2004 19.3944
R8272 gnd.n4661 gnd.n4660 19.3944
R8273 gnd.n4660 gnd.n4659 19.3944
R8274 gnd.n4659 gnd.n4650 19.3944
R8275 gnd.n4655 gnd.n4650 19.3944
R8276 gnd.n4655 gnd.n4654 19.3944
R8277 gnd.n4654 gnd.n1128 19.3944
R8278 gnd.n5889 gnd.n1128 19.3944
R8279 gnd.n5889 gnd.n1129 19.3944
R8280 gnd.n5885 gnd.n1129 19.3944
R8281 gnd.n5885 gnd.n5884 19.3944
R8282 gnd.n5884 gnd.n5883 19.3944
R8283 gnd.n5883 gnd.n1135 19.3944
R8284 gnd.n5879 gnd.n1135 19.3944
R8285 gnd.n5879 gnd.n5878 19.3944
R8286 gnd.n5878 gnd.n5877 19.3944
R8287 gnd.n5877 gnd.n1140 19.3944
R8288 gnd.n5873 gnd.n1140 19.3944
R8289 gnd.n5873 gnd.n5872 19.3944
R8290 gnd.n5872 gnd.n5871 19.3944
R8291 gnd.n5871 gnd.n1145 19.3944
R8292 gnd.n5867 gnd.n1145 19.3944
R8293 gnd.n5867 gnd.n5866 19.3944
R8294 gnd.n5866 gnd.n5865 19.3944
R8295 gnd.n5865 gnd.n1150 19.3944
R8296 gnd.n5861 gnd.n1150 19.3944
R8297 gnd.n5861 gnd.n5860 19.3944
R8298 gnd.n5860 gnd.n5859 19.3944
R8299 gnd.n5859 gnd.n1155 19.3944
R8300 gnd.n5855 gnd.n1155 19.3944
R8301 gnd.n5855 gnd.n5854 19.3944
R8302 gnd.n5854 gnd.n5853 19.3944
R8303 gnd.n5853 gnd.n1160 19.3944
R8304 gnd.n5849 gnd.n1160 19.3944
R8305 gnd.n5849 gnd.n5848 19.3944
R8306 gnd.n5848 gnd.n5847 19.3944
R8307 gnd.n5847 gnd.n1165 19.3944
R8308 gnd.n5843 gnd.n1165 19.3944
R8309 gnd.n5843 gnd.n5842 19.3944
R8310 gnd.n5842 gnd.n5841 19.3944
R8311 gnd.n5841 gnd.n1170 19.3944
R8312 gnd.n5837 gnd.n1170 19.3944
R8313 gnd.n5837 gnd.n5836 19.3944
R8314 gnd.n5836 gnd.n5835 19.3944
R8315 gnd.n5835 gnd.n1175 19.3944
R8316 gnd.n5831 gnd.n1175 19.3944
R8317 gnd.n5831 gnd.n5830 19.3944
R8318 gnd.n5830 gnd.n5829 19.3944
R8319 gnd.n5829 gnd.n1180 19.3944
R8320 gnd.n5825 gnd.n1180 19.3944
R8321 gnd.n5825 gnd.n5824 19.3944
R8322 gnd.n5824 gnd.n5823 19.3944
R8323 gnd.n5823 gnd.n1185 19.3944
R8324 gnd.n5819 gnd.n1185 19.3944
R8325 gnd.n5819 gnd.n5818 19.3944
R8326 gnd.n5818 gnd.n5817 19.3944
R8327 gnd.n5817 gnd.n1190 19.3944
R8328 gnd.n5813 gnd.n1190 19.3944
R8329 gnd.n5813 gnd.n5812 19.3944
R8330 gnd.n5812 gnd.n5811 19.3944
R8331 gnd.n5811 gnd.n1195 19.3944
R8332 gnd.n5807 gnd.n1195 19.3944
R8333 gnd.n5807 gnd.n5806 19.3944
R8334 gnd.n5806 gnd.n5805 19.3944
R8335 gnd.n5805 gnd.n1200 19.3944
R8336 gnd.n5801 gnd.n1200 19.3944
R8337 gnd.n5801 gnd.n5800 19.3944
R8338 gnd.n5800 gnd.n5799 19.3944
R8339 gnd.n5799 gnd.n1205 19.3944
R8340 gnd.n5795 gnd.n1205 19.3944
R8341 gnd.n5795 gnd.n5794 19.3944
R8342 gnd.n5794 gnd.n5793 19.3944
R8343 gnd.n5793 gnd.n1210 19.3944
R8344 gnd.n5789 gnd.n1210 19.3944
R8345 gnd.n5789 gnd.n5788 19.3944
R8346 gnd.n5788 gnd.n5787 19.3944
R8347 gnd.n5787 gnd.n1215 19.3944
R8348 gnd.n5783 gnd.n1215 19.3944
R8349 gnd.n4429 gnd.n4428 19.3944
R8350 gnd.n4428 gnd.n2031 19.3944
R8351 gnd.n4631 gnd.n2031 19.3944
R8352 gnd.n4354 gnd.n4353 19.3944
R8353 gnd.n4357 gnd.n4354 19.3944
R8354 gnd.n4357 gnd.n4337 19.3944
R8355 gnd.n4361 gnd.n4337 19.3944
R8356 gnd.n4362 gnd.n4361 19.3944
R8357 gnd.n4478 gnd.n4362 19.3944
R8358 gnd.n4478 gnd.n4477 19.3944
R8359 gnd.n4477 gnd.n4476 19.3944
R8360 gnd.n4476 gnd.n4367 19.3944
R8361 gnd.n4469 gnd.n4367 19.3944
R8362 gnd.n4469 gnd.n4468 19.3944
R8363 gnd.n4468 gnd.n4376 19.3944
R8364 gnd.n4461 gnd.n4376 19.3944
R8365 gnd.n4461 gnd.n4460 19.3944
R8366 gnd.n4460 gnd.n4386 19.3944
R8367 gnd.n4453 gnd.n4386 19.3944
R8368 gnd.n4453 gnd.n4452 19.3944
R8369 gnd.n4452 gnd.n4396 19.3944
R8370 gnd.n4445 gnd.n4396 19.3944
R8371 gnd.n4445 gnd.n4444 19.3944
R8372 gnd.n4444 gnd.n4406 19.3944
R8373 gnd.n4437 gnd.n4406 19.3944
R8374 gnd.n4437 gnd.n4436 19.3944
R8375 gnd.n4436 gnd.n4416 19.3944
R8376 gnd.n5759 gnd.n1241 19.3944
R8377 gnd.n5759 gnd.n5758 19.3944
R8378 gnd.n5758 gnd.n1244 19.3944
R8379 gnd.n5751 gnd.n1244 19.3944
R8380 gnd.n5751 gnd.n5750 19.3944
R8381 gnd.n5750 gnd.n1252 19.3944
R8382 gnd.n5743 gnd.n1252 19.3944
R8383 gnd.n5743 gnd.n5742 19.3944
R8384 gnd.n5742 gnd.n1260 19.3944
R8385 gnd.n5735 gnd.n1260 19.3944
R8386 gnd.n5735 gnd.n5734 19.3944
R8387 gnd.n5734 gnd.n1268 19.3944
R8388 gnd.n5727 gnd.n1268 19.3944
R8389 gnd.n5727 gnd.n5726 19.3944
R8390 gnd.n5726 gnd.n1276 19.3944
R8391 gnd.n5719 gnd.n1276 19.3944
R8392 gnd.n5477 gnd.n1397 19.3944
R8393 gnd.n5478 gnd.n5477 19.3944
R8394 gnd.n5482 gnd.n5478 19.3944
R8395 gnd.n5483 gnd.n5482 19.3944
R8396 gnd.n5486 gnd.n5483 19.3944
R8397 gnd.n5487 gnd.n5486 19.3944
R8398 gnd.n5491 gnd.n5487 19.3944
R8399 gnd.n5492 gnd.n5491 19.3944
R8400 gnd.n5495 gnd.n5492 19.3944
R8401 gnd.n5496 gnd.n5495 19.3944
R8402 gnd.n5497 gnd.n5496 19.3944
R8403 gnd.n5500 gnd.n5497 19.3944
R8404 gnd.n5500 gnd.n388 19.3944
R8405 gnd.n6796 gnd.n388 19.3944
R8406 gnd.n6797 gnd.n6796 19.3944
R8407 gnd.n6797 gnd.n360 19.3944
R8408 gnd.n6828 gnd.n360 19.3944
R8409 gnd.n6829 gnd.n6828 19.3944
R8410 gnd.n6831 gnd.n6829 19.3944
R8411 gnd.n6832 gnd.n6831 19.3944
R8412 gnd.n6832 gnd.n334 19.3944
R8413 gnd.n6867 gnd.n334 19.3944
R8414 gnd.n6870 gnd.n6867 19.3944
R8415 gnd.n6870 gnd.n6869 19.3944
R8416 gnd.n6869 gnd.n315 19.3944
R8417 gnd.n6890 gnd.n315 19.3944
R8418 gnd.n6891 gnd.n6890 19.3944
R8419 gnd.n6891 gnd.n309 19.3944
R8420 gnd.n6900 gnd.n309 19.3944
R8421 gnd.n6901 gnd.n6900 19.3944
R8422 gnd.n6903 gnd.n6901 19.3944
R8423 gnd.n6904 gnd.n6903 19.3944
R8424 gnd.n6907 gnd.n6904 19.3944
R8425 gnd.n6908 gnd.n6907 19.3944
R8426 gnd.n6910 gnd.n6908 19.3944
R8427 gnd.n6911 gnd.n6910 19.3944
R8428 gnd.n6914 gnd.n6911 19.3944
R8429 gnd.n6915 gnd.n6914 19.3944
R8430 gnd.n6917 gnd.n6915 19.3944
R8431 gnd.n6918 gnd.n6917 19.3944
R8432 gnd.n6921 gnd.n6918 19.3944
R8433 gnd.n6922 gnd.n6921 19.3944
R8434 gnd.n7043 gnd.n6922 19.3944
R8435 gnd.n7044 gnd.n7043 19.3944
R8436 gnd.n7047 gnd.n7044 19.3944
R8437 gnd.n7048 gnd.n7047 19.3944
R8438 gnd.n7050 gnd.n7048 19.3944
R8439 gnd.n7051 gnd.n7050 19.3944
R8440 gnd.n7054 gnd.n7051 19.3944
R8441 gnd.n7055 gnd.n7054 19.3944
R8442 gnd.n7057 gnd.n7055 19.3944
R8443 gnd.n7058 gnd.n7057 19.3944
R8444 gnd.n7061 gnd.n7058 19.3944
R8445 gnd.n7104 gnd.n285 19.3944
R8446 gnd.n7104 gnd.n7101 19.3944
R8447 gnd.n7101 gnd.n7098 19.3944
R8448 gnd.n7098 gnd.n7097 19.3944
R8449 gnd.n7097 gnd.n7094 19.3944
R8450 gnd.n7094 gnd.n7093 19.3944
R8451 gnd.n7093 gnd.n7090 19.3944
R8452 gnd.n7090 gnd.n7089 19.3944
R8453 gnd.n7089 gnd.n7086 19.3944
R8454 gnd.n7086 gnd.n7085 19.3944
R8455 gnd.n7085 gnd.n7082 19.3944
R8456 gnd.n7082 gnd.n7081 19.3944
R8457 gnd.n7081 gnd.n7078 19.3944
R8458 gnd.n7078 gnd.n7077 19.3944
R8459 gnd.n7077 gnd.n7074 19.3944
R8460 gnd.n7074 gnd.n7073 19.3944
R8461 gnd.n7073 gnd.n7070 19.3944
R8462 gnd.n7070 gnd.n7069 19.3944
R8463 gnd.n7147 gnd.n7144 19.3944
R8464 gnd.n7144 gnd.n7143 19.3944
R8465 gnd.n7143 gnd.n7140 19.3944
R8466 gnd.n7140 gnd.n7139 19.3944
R8467 gnd.n7139 gnd.n7136 19.3944
R8468 gnd.n7136 gnd.n7135 19.3944
R8469 gnd.n7135 gnd.n7132 19.3944
R8470 gnd.n7132 gnd.n7131 19.3944
R8471 gnd.n7131 gnd.n7128 19.3944
R8472 gnd.n7128 gnd.n7127 19.3944
R8473 gnd.n7127 gnd.n7124 19.3944
R8474 gnd.n7124 gnd.n7123 19.3944
R8475 gnd.n7123 gnd.n7120 19.3944
R8476 gnd.n7120 gnd.n7119 19.3944
R8477 gnd.n7119 gnd.n7116 19.3944
R8478 gnd.n7116 gnd.n7115 19.3944
R8479 gnd.n7115 gnd.n7112 19.3944
R8480 gnd.n7112 gnd.n7111 19.3944
R8481 gnd.n7185 gnd.n209 19.3944
R8482 gnd.n7180 gnd.n209 19.3944
R8483 gnd.n7180 gnd.n7179 19.3944
R8484 gnd.n7179 gnd.n7178 19.3944
R8485 gnd.n7178 gnd.n7175 19.3944
R8486 gnd.n7175 gnd.n7174 19.3944
R8487 gnd.n7174 gnd.n7171 19.3944
R8488 gnd.n7171 gnd.n7170 19.3944
R8489 gnd.n7170 gnd.n7167 19.3944
R8490 gnd.n7167 gnd.n7166 19.3944
R8491 gnd.n7166 gnd.n7163 19.3944
R8492 gnd.n7163 gnd.n7162 19.3944
R8493 gnd.n7162 gnd.n7159 19.3944
R8494 gnd.n7159 gnd.n7158 19.3944
R8495 gnd.n7158 gnd.n7155 19.3944
R8496 gnd.n7155 gnd.n7154 19.3944
R8497 gnd.n7154 gnd.n7151 19.3944
R8498 gnd.n1414 gnd.n1413 19.3944
R8499 gnd.n5584 gnd.n1413 19.3944
R8500 gnd.n5584 gnd.n5583 19.3944
R8501 gnd.n5583 gnd.n5582 19.3944
R8502 gnd.n5582 gnd.n1420 19.3944
R8503 gnd.n5572 gnd.n1420 19.3944
R8504 gnd.n5572 gnd.n5571 19.3944
R8505 gnd.n5571 gnd.n5570 19.3944
R8506 gnd.n5570 gnd.n1441 19.3944
R8507 gnd.n5560 gnd.n1441 19.3944
R8508 gnd.n5560 gnd.n5559 19.3944
R8509 gnd.n5559 gnd.n377 19.3944
R8510 gnd.n6809 gnd.n377 19.3944
R8511 gnd.n6809 gnd.n375 19.3944
R8512 gnd.n6815 gnd.n375 19.3944
R8513 gnd.n6815 gnd.n6814 19.3944
R8514 gnd.n6814 gnd.n349 19.3944
R8515 gnd.n6843 gnd.n349 19.3944
R8516 gnd.n6843 gnd.n347 19.3944
R8517 gnd.n6849 gnd.n347 19.3944
R8518 gnd.n6849 gnd.n6848 19.3944
R8519 gnd.n6848 gnd.n327 19.3944
R8520 gnd.n6876 gnd.n327 19.3944
R8521 gnd.n6876 gnd.n325 19.3944
R8522 gnd.n6883 gnd.n325 19.3944
R8523 gnd.n6883 gnd.n6882 19.3944
R8524 gnd.n6882 gnd.n90 19.3944
R8525 gnd.n7261 gnd.n90 19.3944
R8526 gnd.n7261 gnd.n7260 19.3944
R8527 gnd.n7260 gnd.n7259 19.3944
R8528 gnd.n7259 gnd.n94 19.3944
R8529 gnd.n7249 gnd.n94 19.3944
R8530 gnd.n7249 gnd.n7248 19.3944
R8531 gnd.n7248 gnd.n7247 19.3944
R8532 gnd.n7247 gnd.n115 19.3944
R8533 gnd.n7237 gnd.n115 19.3944
R8534 gnd.n7237 gnd.n7236 19.3944
R8535 gnd.n7236 gnd.n7235 19.3944
R8536 gnd.n7235 gnd.n134 19.3944
R8537 gnd.n7225 gnd.n134 19.3944
R8538 gnd.n7225 gnd.n7224 19.3944
R8539 gnd.n7224 gnd.n7223 19.3944
R8540 gnd.n7223 gnd.n153 19.3944
R8541 gnd.n7213 gnd.n153 19.3944
R8542 gnd.n7213 gnd.n7212 19.3944
R8543 gnd.n7212 gnd.n7211 19.3944
R8544 gnd.n7211 gnd.n172 19.3944
R8545 gnd.n7201 gnd.n172 19.3944
R8546 gnd.n7201 gnd.n7200 19.3944
R8547 gnd.n7200 gnd.n7199 19.3944
R8548 gnd.n7199 gnd.n191 19.3944
R8549 gnd.n7189 gnd.n191 19.3944
R8550 gnd.n7189 gnd.n7188 19.3944
R8551 gnd.n5710 gnd.n5709 19.3944
R8552 gnd.n5709 gnd.n5708 19.3944
R8553 gnd.n5708 gnd.n5707 19.3944
R8554 gnd.n5707 gnd.n5705 19.3944
R8555 gnd.n5705 gnd.n5702 19.3944
R8556 gnd.n5702 gnd.n5701 19.3944
R8557 gnd.n5701 gnd.n5698 19.3944
R8558 gnd.n5698 gnd.n5697 19.3944
R8559 gnd.n5697 gnd.n5694 19.3944
R8560 gnd.n5694 gnd.n5693 19.3944
R8561 gnd.n5693 gnd.n5690 19.3944
R8562 gnd.n5690 gnd.n5689 19.3944
R8563 gnd.n5689 gnd.n5686 19.3944
R8564 gnd.n5686 gnd.n5685 19.3944
R8565 gnd.n5685 gnd.n5682 19.3944
R8566 gnd.n5682 gnd.n5681 19.3944
R8567 gnd.n5681 gnd.n5678 19.3944
R8568 gnd.n5676 gnd.n5673 19.3944
R8569 gnd.n5673 gnd.n5672 19.3944
R8570 gnd.n5672 gnd.n5669 19.3944
R8571 gnd.n5669 gnd.n5668 19.3944
R8572 gnd.n5668 gnd.n5665 19.3944
R8573 gnd.n5665 gnd.n5664 19.3944
R8574 gnd.n5664 gnd.n5661 19.3944
R8575 gnd.n5659 gnd.n5656 19.3944
R8576 gnd.n5656 gnd.n5655 19.3944
R8577 gnd.n5655 gnd.n5652 19.3944
R8578 gnd.n5652 gnd.n5651 19.3944
R8579 gnd.n5651 gnd.n5648 19.3944
R8580 gnd.n5648 gnd.n5647 19.3944
R8581 gnd.n5647 gnd.n5644 19.3944
R8582 gnd.n5644 gnd.n5643 19.3944
R8583 gnd.n5639 gnd.n5636 19.3944
R8584 gnd.n5636 gnd.n5635 19.3944
R8585 gnd.n5635 gnd.n5632 19.3944
R8586 gnd.n5632 gnd.n5631 19.3944
R8587 gnd.n5631 gnd.n5628 19.3944
R8588 gnd.n5628 gnd.n5627 19.3944
R8589 gnd.n5627 gnd.n5624 19.3944
R8590 gnd.n5624 gnd.n5623 19.3944
R8591 gnd.n5623 gnd.n5620 19.3944
R8592 gnd.n5620 gnd.n5619 19.3944
R8593 gnd.n5619 gnd.n5616 19.3944
R8594 gnd.n5616 gnd.n5615 19.3944
R8595 gnd.n5615 gnd.n5612 19.3944
R8596 gnd.n5612 gnd.n5611 19.3944
R8597 gnd.n5611 gnd.n5608 19.3944
R8598 gnd.n5608 gnd.n5607 19.3944
R8599 gnd.n5607 gnd.n5604 19.3944
R8600 gnd.n5604 gnd.n5603 19.3944
R8601 gnd.n6979 gnd.n6977 19.3944
R8602 gnd.n6982 gnd.n6979 19.3944
R8603 gnd.n6985 gnd.n6982 19.3944
R8604 gnd.n6988 gnd.n6985 19.3944
R8605 gnd.n6988 gnd.n6975 19.3944
R8606 gnd.n6992 gnd.n6975 19.3944
R8607 gnd.n6995 gnd.n6992 19.3944
R8608 gnd.n6998 gnd.n6995 19.3944
R8609 gnd.n6998 gnd.n6973 19.3944
R8610 gnd.n7002 gnd.n6973 19.3944
R8611 gnd.n7005 gnd.n7002 19.3944
R8612 gnd.n7008 gnd.n7005 19.3944
R8613 gnd.n7008 gnd.n6971 19.3944
R8614 gnd.n7012 gnd.n6971 19.3944
R8615 gnd.n7015 gnd.n7012 19.3944
R8616 gnd.n7018 gnd.n7015 19.3944
R8617 gnd.n5523 gnd.n1473 19.3944
R8618 gnd.n5523 gnd.n1474 19.3944
R8619 gnd.n5519 gnd.n1474 19.3944
R8620 gnd.n5519 gnd.n5518 19.3944
R8621 gnd.n5518 gnd.n5517 19.3944
R8622 gnd.n5517 gnd.n5471 19.3944
R8623 gnd.n5513 gnd.n5471 19.3944
R8624 gnd.n5513 gnd.n5512 19.3944
R8625 gnd.n5512 gnd.n5511 19.3944
R8626 gnd.n5511 gnd.n5475 19.3944
R8627 gnd.n5507 gnd.n5475 19.3944
R8628 gnd.n5507 gnd.n5506 19.3944
R8629 gnd.n5506 gnd.n5505 19.3944
R8630 gnd.n5505 gnd.n368 19.3944
R8631 gnd.n6819 gnd.n368 19.3944
R8632 gnd.n6819 gnd.n365 19.3944
R8633 gnd.n6824 gnd.n365 19.3944
R8634 gnd.n6824 gnd.n366 19.3944
R8635 gnd.n366 gnd.n341 19.3944
R8636 gnd.n6853 gnd.n341 19.3944
R8637 gnd.n6853 gnd.n338 19.3944
R8638 gnd.n6863 gnd.n338 19.3944
R8639 gnd.n6863 gnd.n339 19.3944
R8640 gnd.n6859 gnd.n339 19.3944
R8641 gnd.n6859 gnd.n6858 19.3944
R8642 gnd.n6858 gnd.n81 19.3944
R8643 gnd.n7266 gnd.n81 19.3944
R8644 gnd.n7266 gnd.n7265 19.3944
R8645 gnd.n7265 gnd.n83 19.3944
R8646 gnd.n6929 gnd.n83 19.3944
R8647 gnd.n6934 gnd.n6929 19.3944
R8648 gnd.n6935 gnd.n6934 19.3944
R8649 gnd.n6937 gnd.n6935 19.3944
R8650 gnd.n6937 gnd.n6927 19.3944
R8651 gnd.n6942 gnd.n6927 19.3944
R8652 gnd.n6943 gnd.n6942 19.3944
R8653 gnd.n6945 gnd.n6943 19.3944
R8654 gnd.n6945 gnd.n6925 19.3944
R8655 gnd.n6950 gnd.n6925 19.3944
R8656 gnd.n6951 gnd.n6950 19.3944
R8657 gnd.n6953 gnd.n6951 19.3944
R8658 gnd.n6953 gnd.n6923 19.3944
R8659 gnd.n7039 gnd.n6923 19.3944
R8660 gnd.n7039 gnd.n7038 19.3944
R8661 gnd.n7038 gnd.n7037 19.3944
R8662 gnd.n7037 gnd.n7035 19.3944
R8663 gnd.n7035 gnd.n7034 19.3944
R8664 gnd.n7034 gnd.n7032 19.3944
R8665 gnd.n7032 gnd.n7031 19.3944
R8666 gnd.n7031 gnd.n7029 19.3944
R8667 gnd.n7029 gnd.n7028 19.3944
R8668 gnd.n7028 gnd.n7026 19.3944
R8669 gnd.n7026 gnd.n7025 19.3944
R8670 gnd.n5590 gnd.n5589 19.3944
R8671 gnd.n5589 gnd.n5588 19.3944
R8672 gnd.n5588 gnd.n1406 19.3944
R8673 gnd.n5578 gnd.n1406 19.3944
R8674 gnd.n5578 gnd.n5577 19.3944
R8675 gnd.n5577 gnd.n5576 19.3944
R8676 gnd.n5576 gnd.n1430 19.3944
R8677 gnd.n5566 gnd.n1430 19.3944
R8678 gnd.n5566 gnd.n5565 19.3944
R8679 gnd.n5565 gnd.n5564 19.3944
R8680 gnd.n5564 gnd.n1451 19.3944
R8681 gnd.n1451 gnd.n385 19.3944
R8682 gnd.n6805 gnd.n385 19.3944
R8683 gnd.n6805 gnd.n6804 19.3944
R8684 gnd.n6804 gnd.n6803 19.3944
R8685 gnd.n6803 gnd.n6802 19.3944
R8686 gnd.n6802 gnd.n357 19.3944
R8687 gnd.n6839 gnd.n357 19.3944
R8688 gnd.n6839 gnd.n6838 19.3944
R8689 gnd.n6838 gnd.n6837 19.3944
R8690 gnd.n6837 gnd.n6836 19.3944
R8691 gnd.n6836 gnd.n332 19.3944
R8692 gnd.n6872 gnd.n332 19.3944
R8693 gnd.n6872 gnd.n317 19.3944
R8694 gnd.n6887 gnd.n317 19.3944
R8695 gnd.n6887 gnd.n311 19.3944
R8696 gnd.n6895 gnd.n311 19.3944
R8697 gnd.n6896 gnd.n6895 19.3944
R8698 gnd.n6896 gnd.n100 19.3944
R8699 gnd.n7255 gnd.n100 19.3944
R8700 gnd.n7255 gnd.n7254 19.3944
R8701 gnd.n7254 gnd.n7253 19.3944
R8702 gnd.n7253 gnd.n104 19.3944
R8703 gnd.n7243 gnd.n104 19.3944
R8704 gnd.n7243 gnd.n7242 19.3944
R8705 gnd.n7242 gnd.n7241 19.3944
R8706 gnd.n7241 gnd.n124 19.3944
R8707 gnd.n7231 gnd.n124 19.3944
R8708 gnd.n7231 gnd.n7230 19.3944
R8709 gnd.n7230 gnd.n7229 19.3944
R8710 gnd.n7229 gnd.n142 19.3944
R8711 gnd.n7219 gnd.n142 19.3944
R8712 gnd.n7219 gnd.n7218 19.3944
R8713 gnd.n7218 gnd.n7217 19.3944
R8714 gnd.n7217 gnd.n162 19.3944
R8715 gnd.n7207 gnd.n162 19.3944
R8716 gnd.n7207 gnd.n7206 19.3944
R8717 gnd.n7206 gnd.n7205 19.3944
R8718 gnd.n7205 gnd.n180 19.3944
R8719 gnd.n7195 gnd.n180 19.3944
R8720 gnd.n7195 gnd.n7194 19.3944
R8721 gnd.n7194 gnd.n7193 19.3944
R8722 gnd.n7193 gnd.n200 19.3944
R8723 gnd.n2867 gnd.n2866 19.3944
R8724 gnd.n2866 gnd.n2865 19.3944
R8725 gnd.n2865 gnd.n2864 19.3944
R8726 gnd.n2864 gnd.n2862 19.3944
R8727 gnd.n2862 gnd.n2859 19.3944
R8728 gnd.n2859 gnd.n2858 19.3944
R8729 gnd.n2858 gnd.n2855 19.3944
R8730 gnd.n2855 gnd.n2854 19.3944
R8731 gnd.n2854 gnd.n2851 19.3944
R8732 gnd.n2851 gnd.n2850 19.3944
R8733 gnd.n2850 gnd.n2847 19.3944
R8734 gnd.n2847 gnd.n2846 19.3944
R8735 gnd.n2846 gnd.n2843 19.3944
R8736 gnd.n2843 gnd.n2842 19.3944
R8737 gnd.n2842 gnd.n2839 19.3944
R8738 gnd.n2839 gnd.n2838 19.3944
R8739 gnd.n2838 gnd.n2835 19.3944
R8740 gnd.n2835 gnd.n2834 19.3944
R8741 gnd.n2834 gnd.n2831 19.3944
R8742 gnd.n2831 gnd.n2830 19.3944
R8743 gnd.n2830 gnd.n2827 19.3944
R8744 gnd.n2827 gnd.n2826 19.3944
R8745 gnd.n2823 gnd.n2822 19.3944
R8746 gnd.n2822 gnd.n2778 19.3944
R8747 gnd.n2873 gnd.n2778 19.3944
R8748 gnd.n3639 gnd.n3638 19.3944
R8749 gnd.n3638 gnd.n3635 19.3944
R8750 gnd.n3635 gnd.n3634 19.3944
R8751 gnd.n3684 gnd.n3683 19.3944
R8752 gnd.n3683 gnd.n3682 19.3944
R8753 gnd.n3682 gnd.n3679 19.3944
R8754 gnd.n3679 gnd.n3678 19.3944
R8755 gnd.n3678 gnd.n3675 19.3944
R8756 gnd.n3675 gnd.n3674 19.3944
R8757 gnd.n3674 gnd.n3671 19.3944
R8758 gnd.n3671 gnd.n3670 19.3944
R8759 gnd.n3670 gnd.n3667 19.3944
R8760 gnd.n3667 gnd.n3666 19.3944
R8761 gnd.n3666 gnd.n3663 19.3944
R8762 gnd.n3663 gnd.n3662 19.3944
R8763 gnd.n3662 gnd.n3659 19.3944
R8764 gnd.n3659 gnd.n3658 19.3944
R8765 gnd.n3658 gnd.n3655 19.3944
R8766 gnd.n3655 gnd.n3654 19.3944
R8767 gnd.n3654 gnd.n3651 19.3944
R8768 gnd.n3651 gnd.n3650 19.3944
R8769 gnd.n3650 gnd.n3647 19.3944
R8770 gnd.n3647 gnd.n3646 19.3944
R8771 gnd.n3646 gnd.n3643 19.3944
R8772 gnd.n3643 gnd.n3642 19.3944
R8773 gnd.n2966 gnd.n2675 19.3944
R8774 gnd.n2976 gnd.n2675 19.3944
R8775 gnd.n2977 gnd.n2976 19.3944
R8776 gnd.n2977 gnd.n2656 19.3944
R8777 gnd.n2997 gnd.n2656 19.3944
R8778 gnd.n2997 gnd.n2648 19.3944
R8779 gnd.n3007 gnd.n2648 19.3944
R8780 gnd.n3008 gnd.n3007 19.3944
R8781 gnd.n3009 gnd.n3008 19.3944
R8782 gnd.n3009 gnd.n2631 19.3944
R8783 gnd.n3026 gnd.n2631 19.3944
R8784 gnd.n3029 gnd.n3026 19.3944
R8785 gnd.n3029 gnd.n3028 19.3944
R8786 gnd.n3028 gnd.n2604 19.3944
R8787 gnd.n3068 gnd.n2604 19.3944
R8788 gnd.n3068 gnd.n2601 19.3944
R8789 gnd.n3074 gnd.n2601 19.3944
R8790 gnd.n3075 gnd.n3074 19.3944
R8791 gnd.n3075 gnd.n2599 19.3944
R8792 gnd.n3081 gnd.n2599 19.3944
R8793 gnd.n3084 gnd.n3081 19.3944
R8794 gnd.n3086 gnd.n3084 19.3944
R8795 gnd.n3092 gnd.n3086 19.3944
R8796 gnd.n3092 gnd.n3091 19.3944
R8797 gnd.n3091 gnd.n2458 19.3944
R8798 gnd.n3158 gnd.n2458 19.3944
R8799 gnd.n3159 gnd.n3158 19.3944
R8800 gnd.n3159 gnd.n2451 19.3944
R8801 gnd.n3170 gnd.n2451 19.3944
R8802 gnd.n3171 gnd.n3170 19.3944
R8803 gnd.n3171 gnd.n2434 19.3944
R8804 gnd.n2434 gnd.n2432 19.3944
R8805 gnd.n3195 gnd.n2432 19.3944
R8806 gnd.n3196 gnd.n3195 19.3944
R8807 gnd.n3196 gnd.n2403 19.3944
R8808 gnd.n3243 gnd.n2403 19.3944
R8809 gnd.n3244 gnd.n3243 19.3944
R8810 gnd.n3244 gnd.n2396 19.3944
R8811 gnd.n3255 gnd.n2396 19.3944
R8812 gnd.n3256 gnd.n3255 19.3944
R8813 gnd.n3256 gnd.n2379 19.3944
R8814 gnd.n2379 gnd.n2377 19.3944
R8815 gnd.n3280 gnd.n2377 19.3944
R8816 gnd.n3281 gnd.n3280 19.3944
R8817 gnd.n3281 gnd.n2349 19.3944
R8818 gnd.n3332 gnd.n2349 19.3944
R8819 gnd.n3333 gnd.n3332 19.3944
R8820 gnd.n3333 gnd.n2342 19.3944
R8821 gnd.n3600 gnd.n2342 19.3944
R8822 gnd.n3601 gnd.n3600 19.3944
R8823 gnd.n3601 gnd.n2323 19.3944
R8824 gnd.n3626 gnd.n2323 19.3944
R8825 gnd.n3626 gnd.n2324 19.3944
R8826 gnd.n2957 gnd.n2956 19.3944
R8827 gnd.n2956 gnd.n2689 19.3944
R8828 gnd.n2712 gnd.n2689 19.3944
R8829 gnd.n2715 gnd.n2712 19.3944
R8830 gnd.n2715 gnd.n2708 19.3944
R8831 gnd.n2719 gnd.n2708 19.3944
R8832 gnd.n2722 gnd.n2719 19.3944
R8833 gnd.n2725 gnd.n2722 19.3944
R8834 gnd.n2725 gnd.n2706 19.3944
R8835 gnd.n2729 gnd.n2706 19.3944
R8836 gnd.n2732 gnd.n2729 19.3944
R8837 gnd.n2735 gnd.n2732 19.3944
R8838 gnd.n2735 gnd.n2704 19.3944
R8839 gnd.n2739 gnd.n2704 19.3944
R8840 gnd.n2962 gnd.n2961 19.3944
R8841 gnd.n2961 gnd.n2665 19.3944
R8842 gnd.n2987 gnd.n2665 19.3944
R8843 gnd.n2987 gnd.n2663 19.3944
R8844 gnd.n2993 gnd.n2663 19.3944
R8845 gnd.n2993 gnd.n2992 19.3944
R8846 gnd.n2992 gnd.n2637 19.3944
R8847 gnd.n3017 gnd.n2637 19.3944
R8848 gnd.n3017 gnd.n2635 19.3944
R8849 gnd.n3021 gnd.n2635 19.3944
R8850 gnd.n3021 gnd.n2615 19.3944
R8851 gnd.n3048 gnd.n2615 19.3944
R8852 gnd.n3048 gnd.n2613 19.3944
R8853 gnd.n3058 gnd.n2613 19.3944
R8854 gnd.n3058 gnd.n3057 19.3944
R8855 gnd.n3057 gnd.n3056 19.3944
R8856 gnd.n3056 gnd.n2562 19.3944
R8857 gnd.n3106 gnd.n2562 19.3944
R8858 gnd.n3106 gnd.n3105 19.3944
R8859 gnd.n3105 gnd.n3104 19.3944
R8860 gnd.n3104 gnd.n2566 19.3944
R8861 gnd.n2586 gnd.n2566 19.3944
R8862 gnd.n2586 gnd.n2468 19.3944
R8863 gnd.n3143 gnd.n2468 19.3944
R8864 gnd.n3143 gnd.n2466 19.3944
R8865 gnd.n3149 gnd.n2466 19.3944
R8866 gnd.n3149 gnd.n3148 19.3944
R8867 gnd.n3148 gnd.n2441 19.3944
R8868 gnd.n3183 gnd.n2441 19.3944
R8869 gnd.n3183 gnd.n2439 19.3944
R8870 gnd.n3189 gnd.n2439 19.3944
R8871 gnd.n3189 gnd.n3188 19.3944
R8872 gnd.n3188 gnd.n2414 19.3944
R8873 gnd.n3228 gnd.n2414 19.3944
R8874 gnd.n3228 gnd.n2412 19.3944
R8875 gnd.n3234 gnd.n2412 19.3944
R8876 gnd.n3234 gnd.n3233 19.3944
R8877 gnd.n3233 gnd.n2386 19.3944
R8878 gnd.n3268 gnd.n2386 19.3944
R8879 gnd.n3268 gnd.n2384 19.3944
R8880 gnd.n3274 gnd.n2384 19.3944
R8881 gnd.n3274 gnd.n3273 19.3944
R8882 gnd.n3273 gnd.n2359 19.3944
R8883 gnd.n3317 gnd.n2359 19.3944
R8884 gnd.n3317 gnd.n2357 19.3944
R8885 gnd.n3323 gnd.n2357 19.3944
R8886 gnd.n3323 gnd.n3322 19.3944
R8887 gnd.n3322 gnd.n2332 19.3944
R8888 gnd.n3611 gnd.n2332 19.3944
R8889 gnd.n3611 gnd.n2330 19.3944
R8890 gnd.n3619 gnd.n2330 19.3944
R8891 gnd.n3619 gnd.n3618 19.3944
R8892 gnd.n3618 gnd.n3617 19.3944
R8893 gnd.n3720 gnd.n3719 19.3944
R8894 gnd.n3719 gnd.n2270 19.3944
R8895 gnd.n3715 gnd.n2270 19.3944
R8896 gnd.n3715 gnd.n3712 19.3944
R8897 gnd.n3712 gnd.n3709 19.3944
R8898 gnd.n3709 gnd.n3708 19.3944
R8899 gnd.n3708 gnd.n3705 19.3944
R8900 gnd.n3705 gnd.n3704 19.3944
R8901 gnd.n3704 gnd.n3701 19.3944
R8902 gnd.n3701 gnd.n3700 19.3944
R8903 gnd.n3700 gnd.n3697 19.3944
R8904 gnd.n3697 gnd.n3696 19.3944
R8905 gnd.n3696 gnd.n3693 19.3944
R8906 gnd.n3693 gnd.n3692 19.3944
R8907 gnd.n2877 gnd.n2776 19.3944
R8908 gnd.n2877 gnd.n2767 19.3944
R8909 gnd.n2890 gnd.n2767 19.3944
R8910 gnd.n2890 gnd.n2765 19.3944
R8911 gnd.n2894 gnd.n2765 19.3944
R8912 gnd.n2894 gnd.n2755 19.3944
R8913 gnd.n2906 gnd.n2755 19.3944
R8914 gnd.n2906 gnd.n2753 19.3944
R8915 gnd.n2940 gnd.n2753 19.3944
R8916 gnd.n2940 gnd.n2939 19.3944
R8917 gnd.n2939 gnd.n2938 19.3944
R8918 gnd.n2938 gnd.n2937 19.3944
R8919 gnd.n2937 gnd.n2934 19.3944
R8920 gnd.n2934 gnd.n2933 19.3944
R8921 gnd.n2933 gnd.n2932 19.3944
R8922 gnd.n2932 gnd.n2930 19.3944
R8923 gnd.n2930 gnd.n2929 19.3944
R8924 gnd.n2929 gnd.n2926 19.3944
R8925 gnd.n2926 gnd.n2925 19.3944
R8926 gnd.n2925 gnd.n2924 19.3944
R8927 gnd.n2924 gnd.n2922 19.3944
R8928 gnd.n2922 gnd.n2621 19.3944
R8929 gnd.n3037 gnd.n2621 19.3944
R8930 gnd.n3037 gnd.n2619 19.3944
R8931 gnd.n3043 gnd.n2619 19.3944
R8932 gnd.n3043 gnd.n3042 19.3944
R8933 gnd.n3042 gnd.n2543 19.3944
R8934 gnd.n3117 gnd.n2543 19.3944
R8935 gnd.n3117 gnd.n2544 19.3944
R8936 gnd.n2591 gnd.n2590 19.3944
R8937 gnd.n2594 gnd.n2593 19.3944
R8938 gnd.n2581 gnd.n2580 19.3944
R8939 gnd.n3136 gnd.n2473 19.3944
R8940 gnd.n3136 gnd.n3135 19.3944
R8941 gnd.n3135 gnd.n3134 19.3944
R8942 gnd.n3134 gnd.n3132 19.3944
R8943 gnd.n3132 gnd.n3131 19.3944
R8944 gnd.n3131 gnd.n3129 19.3944
R8945 gnd.n3129 gnd.n3128 19.3944
R8946 gnd.n3128 gnd.n2422 19.3944
R8947 gnd.n3204 gnd.n2422 19.3944
R8948 gnd.n3204 gnd.n2420 19.3944
R8949 gnd.n3223 gnd.n2420 19.3944
R8950 gnd.n3223 gnd.n3222 19.3944
R8951 gnd.n3222 gnd.n3221 19.3944
R8952 gnd.n3221 gnd.n3219 19.3944
R8953 gnd.n3219 gnd.n3218 19.3944
R8954 gnd.n3218 gnd.n3216 19.3944
R8955 gnd.n3216 gnd.n3215 19.3944
R8956 gnd.n3215 gnd.n2366 19.3944
R8957 gnd.n3289 gnd.n2366 19.3944
R8958 gnd.n3289 gnd.n2364 19.3944
R8959 gnd.n3312 gnd.n2364 19.3944
R8960 gnd.n3312 gnd.n3311 19.3944
R8961 gnd.n3311 gnd.n3310 19.3944
R8962 gnd.n3310 gnd.n3307 19.3944
R8963 gnd.n3307 gnd.n3306 19.3944
R8964 gnd.n3306 gnd.n3304 19.3944
R8965 gnd.n3304 gnd.n3303 19.3944
R8966 gnd.n3303 gnd.n3301 19.3944
R8967 gnd.n3301 gnd.n2317 19.3944
R8968 gnd.n2882 gnd.n2772 19.3944
R8969 gnd.n2882 gnd.n2770 19.3944
R8970 gnd.n2886 gnd.n2770 19.3944
R8971 gnd.n2886 gnd.n2761 19.3944
R8972 gnd.n2898 gnd.n2761 19.3944
R8973 gnd.n2898 gnd.n2759 19.3944
R8974 gnd.n2902 gnd.n2759 19.3944
R8975 gnd.n2902 gnd.n2748 19.3944
R8976 gnd.n2944 gnd.n2748 19.3944
R8977 gnd.n2944 gnd.n2702 19.3944
R8978 gnd.n2950 gnd.n2702 19.3944
R8979 gnd.n2950 gnd.n2949 19.3944
R8980 gnd.n2949 gnd.n2680 19.3944
R8981 gnd.n2971 gnd.n2680 19.3944
R8982 gnd.n2971 gnd.n2673 19.3944
R8983 gnd.n2982 gnd.n2673 19.3944
R8984 gnd.n2982 gnd.n2981 19.3944
R8985 gnd.n2981 gnd.n2654 19.3944
R8986 gnd.n3002 gnd.n2654 19.3944
R8987 gnd.n3002 gnd.n2644 19.3944
R8988 gnd.n3012 gnd.n2644 19.3944
R8989 gnd.n3012 gnd.n2627 19.3944
R8990 gnd.n3033 gnd.n2627 19.3944
R8991 gnd.n3033 gnd.n3032 19.3944
R8992 gnd.n3032 gnd.n2606 19.3944
R8993 gnd.n3063 gnd.n2606 19.3944
R8994 gnd.n3063 gnd.n2551 19.3944
R8995 gnd.n3113 gnd.n2551 19.3944
R8996 gnd.n3113 gnd.n3112 19.3944
R8997 gnd.n3112 gnd.n3111 19.3944
R8998 gnd.n3111 gnd.n2555 19.3944
R8999 gnd.n2573 gnd.n2555 19.3944
R9000 gnd.n3099 gnd.n2573 19.3944
R9001 gnd.n3099 gnd.n3098 19.3944
R9002 gnd.n3098 gnd.n3097 19.3944
R9003 gnd.n3097 gnd.n2577 19.3944
R9004 gnd.n2577 gnd.n2460 19.3944
R9005 gnd.n3154 gnd.n2460 19.3944
R9006 gnd.n3154 gnd.n2453 19.3944
R9007 gnd.n3165 gnd.n2453 19.3944
R9008 gnd.n3165 gnd.n2449 19.3944
R9009 gnd.n3178 gnd.n2449 19.3944
R9010 gnd.n3178 gnd.n3177 19.3944
R9011 gnd.n3177 gnd.n2428 19.3944
R9012 gnd.n3200 gnd.n2428 19.3944
R9013 gnd.n3200 gnd.n3199 19.3944
R9014 gnd.n3199 gnd.n2405 19.3944
R9015 gnd.n3239 gnd.n2405 19.3944
R9016 gnd.n3239 gnd.n2398 19.3944
R9017 gnd.n3250 gnd.n2398 19.3944
R9018 gnd.n3250 gnd.n2394 19.3944
R9019 gnd.n3263 gnd.n2394 19.3944
R9020 gnd.n3263 gnd.n3262 19.3944
R9021 gnd.n3262 gnd.n2373 19.3944
R9022 gnd.n3285 gnd.n2373 19.3944
R9023 gnd.n3285 gnd.n3284 19.3944
R9024 gnd.n3284 gnd.n2351 19.3944
R9025 gnd.n3328 gnd.n2351 19.3944
R9026 gnd.n3328 gnd.n2344 19.3944
R9027 gnd.n3339 gnd.n2344 19.3944
R9028 gnd.n3339 gnd.n2340 19.3944
R9029 gnd.n3606 gnd.n2340 19.3944
R9030 gnd.n3606 gnd.n3605 19.3944
R9031 gnd.n3605 gnd.n2321 19.3944
R9032 gnd.n3629 gnd.n2321 19.3944
R9033 gnd.n4473 gnd.n4472 19.3944
R9034 gnd.n4472 gnd.n4370 19.3944
R9035 gnd.n4465 gnd.n4370 19.3944
R9036 gnd.n4465 gnd.n4464 19.3944
R9037 gnd.n4464 gnd.n4382 19.3944
R9038 gnd.n4457 gnd.n4382 19.3944
R9039 gnd.n4457 gnd.n4456 19.3944
R9040 gnd.n4456 gnd.n4390 19.3944
R9041 gnd.n4449 gnd.n4390 19.3944
R9042 gnd.n4449 gnd.n4448 19.3944
R9043 gnd.n4448 gnd.n4402 19.3944
R9044 gnd.n4441 gnd.n4402 19.3944
R9045 gnd.n4441 gnd.n4440 19.3944
R9046 gnd.n4440 gnd.n4410 19.3944
R9047 gnd.n4433 gnd.n4410 19.3944
R9048 gnd.n4433 gnd.n4432 19.3944
R9049 gnd.n4041 gnd.n4040 19.3944
R9050 gnd.n4042 gnd.n4041 19.3944
R9051 gnd.n4042 gnd.n2223 19.3944
R9052 gnd.n4060 gnd.n2223 19.3944
R9053 gnd.n4061 gnd.n4060 19.3944
R9054 gnd.n4062 gnd.n4061 19.3944
R9055 gnd.n4062 gnd.n2205 19.3944
R9056 gnd.n4080 gnd.n2205 19.3944
R9057 gnd.n4081 gnd.n4080 19.3944
R9058 gnd.n4082 gnd.n4081 19.3944
R9059 gnd.n4082 gnd.n2187 19.3944
R9060 gnd.n4100 gnd.n2187 19.3944
R9061 gnd.n4101 gnd.n4100 19.3944
R9062 gnd.n4103 gnd.n4101 19.3944
R9063 gnd.n4104 gnd.n4103 19.3944
R9064 gnd.n4104 gnd.n2161 19.3944
R9065 gnd.n4135 gnd.n2161 19.3944
R9066 gnd.n4136 gnd.n4135 19.3944
R9067 gnd.n4138 gnd.n4136 19.3944
R9068 gnd.n4139 gnd.n4138 19.3944
R9069 gnd.n4139 gnd.n2136 19.3944
R9070 gnd.n4170 gnd.n2136 19.3944
R9071 gnd.n4171 gnd.n4170 19.3944
R9072 gnd.n4173 gnd.n4171 19.3944
R9073 gnd.n4174 gnd.n4173 19.3944
R9074 gnd.n4174 gnd.n2110 19.3944
R9075 gnd.n4217 gnd.n2110 19.3944
R9076 gnd.n4218 gnd.n4217 19.3944
R9077 gnd.n4219 gnd.n4218 19.3944
R9078 gnd.n4219 gnd.n2093 19.3944
R9079 gnd.n4237 gnd.n2093 19.3944
R9080 gnd.n4238 gnd.n4237 19.3944
R9081 gnd.n4240 gnd.n4238 19.3944
R9082 gnd.n4241 gnd.n4240 19.3944
R9083 gnd.n4243 gnd.n4241 19.3944
R9084 gnd.n4243 gnd.n2070 19.3944
R9085 gnd.n4273 gnd.n2070 19.3944
R9086 gnd.n4274 gnd.n4273 19.3944
R9087 gnd.n4275 gnd.n4274 19.3944
R9088 gnd.n4276 gnd.n4275 19.3944
R9089 gnd.n4280 gnd.n4276 19.3944
R9090 gnd.n4280 gnd.n4279 19.3944
R9091 gnd.n4279 gnd.n4278 19.3944
R9092 gnd.n4278 gnd.n2055 19.3944
R9093 gnd.n4326 gnd.n2055 19.3944
R9094 gnd.n4327 gnd.n4326 19.3944
R9095 gnd.n4328 gnd.n4327 19.3944
R9096 gnd.n4329 gnd.n4328 19.3944
R9097 gnd.n4333 gnd.n4329 19.3944
R9098 gnd.n4334 gnd.n4333 19.3944
R9099 gnd.n4581 gnd.n4334 19.3944
R9100 gnd.n4581 gnd.n4580 19.3944
R9101 gnd.n4580 gnd.n4579 19.3944
R9102 gnd.n3916 gnd.n3914 19.3944
R9103 gnd.n3914 gnd.n3911 19.3944
R9104 gnd.n3911 gnd.n3910 19.3944
R9105 gnd.n3910 gnd.n3907 19.3944
R9106 gnd.n3907 gnd.n3906 19.3944
R9107 gnd.n3906 gnd.n3903 19.3944
R9108 gnd.n3903 gnd.n3902 19.3944
R9109 gnd.n3902 gnd.n3899 19.3944
R9110 gnd.n3899 gnd.n3898 19.3944
R9111 gnd.n3898 gnd.n3895 19.3944
R9112 gnd.n3895 gnd.n3894 19.3944
R9113 gnd.n3894 gnd.n3891 19.3944
R9114 gnd.n3891 gnd.n3890 19.3944
R9115 gnd.n3890 gnd.n3887 19.3944
R9116 gnd.n3887 gnd.n3886 19.3944
R9117 gnd.n3886 gnd.n3883 19.3944
R9118 gnd.n3877 gnd.n3875 19.3944
R9119 gnd.n3875 gnd.n3874 19.3944
R9120 gnd.n3874 gnd.n3872 19.3944
R9121 gnd.n3872 gnd.n3871 19.3944
R9122 gnd.n3871 gnd.n3869 19.3944
R9123 gnd.n3869 gnd.n3868 19.3944
R9124 gnd.n3868 gnd.n3866 19.3944
R9125 gnd.n3866 gnd.n3865 19.3944
R9126 gnd.n3865 gnd.n3863 19.3944
R9127 gnd.n3863 gnd.n3862 19.3944
R9128 gnd.n3862 gnd.n3860 19.3944
R9129 gnd.n3860 gnd.n3859 19.3944
R9130 gnd.n3859 gnd.n3857 19.3944
R9131 gnd.n3857 gnd.n2168 19.3944
R9132 gnd.n4125 gnd.n2168 19.3944
R9133 gnd.n4125 gnd.n2166 19.3944
R9134 gnd.n4131 gnd.n2166 19.3944
R9135 gnd.n4131 gnd.n4130 19.3944
R9136 gnd.n4130 gnd.n2143 19.3944
R9137 gnd.n4160 gnd.n2143 19.3944
R9138 gnd.n4160 gnd.n2141 19.3944
R9139 gnd.n4166 gnd.n2141 19.3944
R9140 gnd.n4166 gnd.n4165 19.3944
R9141 gnd.n4165 gnd.n2118 19.3944
R9142 gnd.n4195 gnd.n2118 19.3944
R9143 gnd.n4195 gnd.n2115 19.3944
R9144 gnd.n4213 gnd.n2115 19.3944
R9145 gnd.n4213 gnd.n2116 19.3944
R9146 gnd.n4209 gnd.n2116 19.3944
R9147 gnd.n4209 gnd.n4208 19.3944
R9148 gnd.n4208 gnd.n4207 19.3944
R9149 gnd.n4207 gnd.n4202 19.3944
R9150 gnd.n4203 gnd.n4202 19.3944
R9151 gnd.n4203 gnd.n2074 19.3944
R9152 gnd.n4265 gnd.n2074 19.3944
R9153 gnd.n4265 gnd.n2072 19.3944
R9154 gnd.n4269 gnd.n2072 19.3944
R9155 gnd.n4269 gnd.n2067 19.3944
R9156 gnd.n4288 gnd.n2067 19.3944
R9157 gnd.n4288 gnd.n2068 19.3944
R9158 gnd.n4284 gnd.n2068 19.3944
R9159 gnd.n4284 gnd.n2059 19.3944
R9160 gnd.n4318 gnd.n2059 19.3944
R9161 gnd.n4318 gnd.n2057 19.3944
R9162 gnd.n4322 gnd.n2057 19.3944
R9163 gnd.n4322 gnd.n2050 19.3944
R9164 gnd.n4594 gnd.n2050 19.3944
R9165 gnd.n4594 gnd.n2051 19.3944
R9166 gnd.n4590 gnd.n2051 19.3944
R9167 gnd.n4590 gnd.n4589 19.3944
R9168 gnd.n4589 gnd.n4588 19.3944
R9169 gnd.n4588 gnd.n4585 19.3944
R9170 gnd.n4585 gnd.n2037 19.3944
R9171 gnd.n4033 gnd.n4032 19.3944
R9172 gnd.n4032 gnd.n4031 19.3944
R9173 gnd.n4031 gnd.n4030 19.3944
R9174 gnd.n4030 gnd.n4028 19.3944
R9175 gnd.n4028 gnd.n4025 19.3944
R9176 gnd.n4025 gnd.n4024 19.3944
R9177 gnd.n4024 gnd.n4021 19.3944
R9178 gnd.n4021 gnd.n4020 19.3944
R9179 gnd.n4020 gnd.n4017 19.3944
R9180 gnd.n4017 gnd.n4016 19.3944
R9181 gnd.n4016 gnd.n4013 19.3944
R9182 gnd.n4013 gnd.n4012 19.3944
R9183 gnd.n4012 gnd.n4009 19.3944
R9184 gnd.n4009 gnd.n4008 19.3944
R9185 gnd.n4008 gnd.n4005 19.3944
R9186 gnd.n4005 gnd.n4004 19.3944
R9187 gnd.n4004 gnd.n4001 19.3944
R9188 gnd.n3999 gnd.n3996 19.3944
R9189 gnd.n3996 gnd.n3995 19.3944
R9190 gnd.n3995 gnd.n3992 19.3944
R9191 gnd.n3992 gnd.n3991 19.3944
R9192 gnd.n3991 gnd.n3988 19.3944
R9193 gnd.n3988 gnd.n3987 19.3944
R9194 gnd.n3987 gnd.n3984 19.3944
R9195 gnd.n3984 gnd.n3983 19.3944
R9196 gnd.n3983 gnd.n3980 19.3944
R9197 gnd.n3980 gnd.n3979 19.3944
R9198 gnd.n3979 gnd.n3976 19.3944
R9199 gnd.n3976 gnd.n3975 19.3944
R9200 gnd.n3975 gnd.n3972 19.3944
R9201 gnd.n3972 gnd.n3971 19.3944
R9202 gnd.n3971 gnd.n3968 19.3944
R9203 gnd.n3968 gnd.n3967 19.3944
R9204 gnd.n3967 gnd.n3964 19.3944
R9205 gnd.n3964 gnd.n3963 19.3944
R9206 gnd.n3959 gnd.n3956 19.3944
R9207 gnd.n3956 gnd.n3955 19.3944
R9208 gnd.n3955 gnd.n3952 19.3944
R9209 gnd.n3952 gnd.n3951 19.3944
R9210 gnd.n3951 gnd.n3948 19.3944
R9211 gnd.n3948 gnd.n3947 19.3944
R9212 gnd.n3947 gnd.n3944 19.3944
R9213 gnd.n3944 gnd.n3943 19.3944
R9214 gnd.n3943 gnd.n3940 19.3944
R9215 gnd.n3940 gnd.n3939 19.3944
R9216 gnd.n3939 gnd.n3936 19.3944
R9217 gnd.n3936 gnd.n3935 19.3944
R9218 gnd.n3935 gnd.n3932 19.3944
R9219 gnd.n3932 gnd.n3931 19.3944
R9220 gnd.n3931 gnd.n3928 19.3944
R9221 gnd.n3928 gnd.n3927 19.3944
R9222 gnd.n3927 gnd.n3924 19.3944
R9223 gnd.n3924 gnd.n3923 19.3944
R9224 gnd.n4051 gnd.n2232 19.3944
R9225 gnd.n4051 gnd.n2230 19.3944
R9226 gnd.n4055 gnd.n2230 19.3944
R9227 gnd.n4055 gnd.n2213 19.3944
R9228 gnd.n4071 gnd.n2213 19.3944
R9229 gnd.n4071 gnd.n2211 19.3944
R9230 gnd.n4075 gnd.n2211 19.3944
R9231 gnd.n4075 gnd.n2196 19.3944
R9232 gnd.n4091 gnd.n2196 19.3944
R9233 gnd.n4091 gnd.n2194 19.3944
R9234 gnd.n4095 gnd.n2194 19.3944
R9235 gnd.n4095 gnd.n2176 19.3944
R9236 gnd.n4115 gnd.n2176 19.3944
R9237 gnd.n4115 gnd.n2174 19.3944
R9238 gnd.n4121 gnd.n2174 19.3944
R9239 gnd.n4121 gnd.n4120 19.3944
R9240 gnd.n4120 gnd.n2151 19.3944
R9241 gnd.n4150 gnd.n2151 19.3944
R9242 gnd.n4150 gnd.n2149 19.3944
R9243 gnd.n4156 gnd.n2149 19.3944
R9244 gnd.n4156 gnd.n4155 19.3944
R9245 gnd.n4155 gnd.n2127 19.3944
R9246 gnd.n4185 gnd.n2127 19.3944
R9247 gnd.n4185 gnd.n2125 19.3944
R9248 gnd.n4191 gnd.n2125 19.3944
R9249 gnd.n4191 gnd.n4190 19.3944
R9250 gnd.n4190 gnd.n2102 19.3944
R9251 gnd.n4228 gnd.n2102 19.3944
R9252 gnd.n4228 gnd.n2100 19.3944
R9253 gnd.n4232 gnd.n2100 19.3944
R9254 gnd.n4232 gnd.n2081 19.3944
R9255 gnd.n4255 gnd.n2081 19.3944
R9256 gnd.n4255 gnd.n2079 19.3944
R9257 gnd.n4260 gnd.n2079 19.3944
R9258 gnd.n4260 gnd.n890 19.3944
R9259 gnd.n6077 gnd.n890 19.3944
R9260 gnd.n6077 gnd.n6076 19.3944
R9261 gnd.n6076 gnd.n6075 19.3944
R9262 gnd.n6075 gnd.n894 19.3944
R9263 gnd.n6065 gnd.n894 19.3944
R9264 gnd.n6065 gnd.n6064 19.3944
R9265 gnd.n6064 gnd.n6063 19.3944
R9266 gnd.n6063 gnd.n916 19.3944
R9267 gnd.n6053 gnd.n916 19.3944
R9268 gnd.n6053 gnd.n6052 19.3944
R9269 gnd.n6052 gnd.n6051 19.3944
R9270 gnd.n6051 gnd.n936 19.3944
R9271 gnd.n6041 gnd.n936 19.3944
R9272 gnd.n6041 gnd.n6040 19.3944
R9273 gnd.n6040 gnd.n6039 19.3944
R9274 gnd.n6039 gnd.n956 19.3944
R9275 gnd.n6029 gnd.n956 19.3944
R9276 gnd.n6029 gnd.n6028 19.3944
R9277 gnd.n6025 gnd.n976 19.3944
R9278 gnd.n6020 gnd.n976 19.3944
R9279 gnd.n6020 gnd.n6019 19.3944
R9280 gnd.n6019 gnd.n6018 19.3944
R9281 gnd.n6018 gnd.n6015 19.3944
R9282 gnd.n6015 gnd.n6014 19.3944
R9283 gnd.n6014 gnd.n6011 19.3944
R9284 gnd.n6011 gnd.n6010 19.3944
R9285 gnd.n6010 gnd.n6007 19.3944
R9286 gnd.n6007 gnd.n6006 19.3944
R9287 gnd.n6006 gnd.n6003 19.3944
R9288 gnd.n6003 gnd.n6002 19.3944
R9289 gnd.n6002 gnd.n5999 19.3944
R9290 gnd.n5999 gnd.n5998 19.3944
R9291 gnd.n5998 gnd.n5995 19.3944
R9292 gnd.n5995 gnd.n5994 19.3944
R9293 gnd.n5994 gnd.n5991 19.3944
R9294 gnd.n4527 gnd.n4493 19.3944
R9295 gnd.n4531 gnd.n4493 19.3944
R9296 gnd.n4534 gnd.n4531 19.3944
R9297 gnd.n4537 gnd.n4534 19.3944
R9298 gnd.n4537 gnd.n4491 19.3944
R9299 gnd.n4541 gnd.n4491 19.3944
R9300 gnd.n4544 gnd.n4541 19.3944
R9301 gnd.n4547 gnd.n4544 19.3944
R9302 gnd.n4547 gnd.n4489 19.3944
R9303 gnd.n4551 gnd.n4489 19.3944
R9304 gnd.n4554 gnd.n4551 19.3944
R9305 gnd.n4557 gnd.n4554 19.3944
R9306 gnd.n4557 gnd.n4487 19.3944
R9307 gnd.n4561 gnd.n4487 19.3944
R9308 gnd.n4564 gnd.n4561 19.3944
R9309 gnd.n4567 gnd.n4564 19.3944
R9310 gnd.n4567 gnd.n4485 19.3944
R9311 gnd.n4572 gnd.n4485 19.3944
R9312 gnd.n4505 gnd.n1045 19.3944
R9313 gnd.n4508 gnd.n4505 19.3944
R9314 gnd.n4508 gnd.n4500 19.3944
R9315 gnd.n4512 gnd.n4500 19.3944
R9316 gnd.n4515 gnd.n4512 19.3944
R9317 gnd.n4518 gnd.n4515 19.3944
R9318 gnd.n4518 gnd.n4498 19.3944
R9319 gnd.n4523 gnd.n4498 19.3944
R9320 gnd.n5989 gnd.n5986 19.3944
R9321 gnd.n5986 gnd.n5985 19.3944
R9322 gnd.n5985 gnd.n5982 19.3944
R9323 gnd.n5982 gnd.n5981 19.3944
R9324 gnd.n5981 gnd.n5978 19.3944
R9325 gnd.n5978 gnd.n5977 19.3944
R9326 gnd.n5977 gnd.n5974 19.3944
R9327 gnd.n4047 gnd.n2239 19.3944
R9328 gnd.n4047 gnd.n4046 19.3944
R9329 gnd.n4046 gnd.n4045 19.3944
R9330 gnd.n4045 gnd.n2221 19.3944
R9331 gnd.n4067 gnd.n2221 19.3944
R9332 gnd.n4067 gnd.n4066 19.3944
R9333 gnd.n4066 gnd.n4065 19.3944
R9334 gnd.n4065 gnd.n2203 19.3944
R9335 gnd.n4087 gnd.n2203 19.3944
R9336 gnd.n4087 gnd.n4086 19.3944
R9337 gnd.n4086 gnd.n4085 19.3944
R9338 gnd.n4085 gnd.n2184 19.3944
R9339 gnd.n4111 gnd.n2184 19.3944
R9340 gnd.n4111 gnd.n4110 19.3944
R9341 gnd.n4110 gnd.n4109 19.3944
R9342 gnd.n4109 gnd.n4108 19.3944
R9343 gnd.n4108 gnd.n2158 19.3944
R9344 gnd.n4146 gnd.n2158 19.3944
R9345 gnd.n4146 gnd.n4145 19.3944
R9346 gnd.n4145 gnd.n4144 19.3944
R9347 gnd.n4144 gnd.n4143 19.3944
R9348 gnd.n4143 gnd.n2133 19.3944
R9349 gnd.n4181 gnd.n2133 19.3944
R9350 gnd.n4181 gnd.n4180 19.3944
R9351 gnd.n4180 gnd.n4179 19.3944
R9352 gnd.n4179 gnd.n4178 19.3944
R9353 gnd.n4178 gnd.n2108 19.3944
R9354 gnd.n4224 gnd.n2108 19.3944
R9355 gnd.n4224 gnd.n4223 19.3944
R9356 gnd.n4223 gnd.n4222 19.3944
R9357 gnd.n4222 gnd.n2089 19.3944
R9358 gnd.n4251 gnd.n2089 19.3944
R9359 gnd.n4251 gnd.n4250 19.3944
R9360 gnd.n4250 gnd.n4249 19.3944
R9361 gnd.n4249 gnd.n4248 19.3944
R9362 gnd.n4248 gnd.n4246 19.3944
R9363 gnd.n4246 gnd.n901 19.3944
R9364 gnd.n6071 gnd.n901 19.3944
R9365 gnd.n6071 gnd.n6070 19.3944
R9366 gnd.n6070 gnd.n6069 19.3944
R9367 gnd.n6069 gnd.n905 19.3944
R9368 gnd.n6059 gnd.n905 19.3944
R9369 gnd.n6059 gnd.n6058 19.3944
R9370 gnd.n6058 gnd.n6057 19.3944
R9371 gnd.n6057 gnd.n926 19.3944
R9372 gnd.n6047 gnd.n926 19.3944
R9373 gnd.n6047 gnd.n6046 19.3944
R9374 gnd.n6046 gnd.n6045 19.3944
R9375 gnd.n6045 gnd.n945 19.3944
R9376 gnd.n6035 gnd.n945 19.3944
R9377 gnd.n6035 gnd.n6034 19.3944
R9378 gnd.n6034 gnd.n6033 19.3944
R9379 gnd.n6033 gnd.n966 19.3944
R9380 gnd.n4297 gnd.n4295 19.3944
R9381 gnd.n4297 gnd.n4293 19.3944
R9382 gnd.n4301 gnd.n4293 19.3944
R9383 gnd.n4301 gnd.n2065 19.3944
R9384 gnd.n4305 gnd.n2065 19.3944
R9385 gnd.n4305 gnd.n2063 19.3944
R9386 gnd.n4313 gnd.n2063 19.3944
R9387 gnd.n4313 gnd.n4312 19.3944
R9388 gnd.n4312 gnd.n4311 19.3944
R9389 gnd.n4311 gnd.n2047 19.3944
R9390 gnd.n4600 gnd.n2047 19.3944
R9391 gnd.n4600 gnd.n2045 19.3944
R9392 gnd.n4604 gnd.n2045 19.3944
R9393 gnd.n4604 gnd.n2043 19.3944
R9394 gnd.n4608 gnd.n2043 19.3944
R9395 gnd.n4608 gnd.n2041 19.3944
R9396 gnd.n4620 gnd.n2041 19.3944
R9397 gnd.n4620 gnd.n4619 19.3944
R9398 gnd.n4619 gnd.n4618 19.3944
R9399 gnd.n4618 gnd.n4615 19.3944
R9400 gnd.n4615 gnd.n2013 19.3944
R9401 gnd.n4636 gnd.n2013 19.3944
R9402 gnd.n4636 gnd.n2011 19.3944
R9403 gnd.n4640 gnd.n2011 19.3944
R9404 gnd.n4640 gnd.n1997 19.3944
R9405 gnd.n4669 gnd.n1997 19.3944
R9406 gnd.n4669 gnd.n1995 19.3944
R9407 gnd.n4682 gnd.n1995 19.3944
R9408 gnd.n4682 gnd.n4681 19.3944
R9409 gnd.n4681 gnd.n4680 19.3944
R9410 gnd.n4680 gnd.n4677 19.3944
R9411 gnd.n4677 gnd.n1118 19.3944
R9412 gnd.n5895 gnd.n1118 19.3944
R9413 gnd.n5895 gnd.n5894 19.3944
R9414 gnd.n5894 gnd.n5893 19.3944
R9415 gnd.n5893 gnd.n1122 19.3944
R9416 gnd.n4865 gnd.n1122 19.3944
R9417 gnd.n4869 gnd.n4865 19.3944
R9418 gnd.n4869 gnd.n1886 19.3944
R9419 gnd.n4894 gnd.n1886 19.3944
R9420 gnd.n4894 gnd.n1884 19.3944
R9421 gnd.n4909 gnd.n1884 19.3944
R9422 gnd.n4909 gnd.n4908 19.3944
R9423 gnd.n4908 gnd.n4907 19.3944
R9424 gnd.n4907 gnd.n4900 19.3944
R9425 gnd.n4903 gnd.n4900 19.3944
R9426 gnd.n4903 gnd.n1848 19.3944
R9427 gnd.n4952 gnd.n1848 19.3944
R9428 gnd.n4952 gnd.n1846 19.3944
R9429 gnd.n4956 gnd.n1846 19.3944
R9430 gnd.n4956 gnd.n1830 19.3944
R9431 gnd.n4978 gnd.n1830 19.3944
R9432 gnd.n4978 gnd.n1828 19.3944
R9433 gnd.n4984 gnd.n1828 19.3944
R9434 gnd.n4984 gnd.n4983 19.3944
R9435 gnd.n4983 gnd.n1806 19.3944
R9436 gnd.n5017 gnd.n1806 19.3944
R9437 gnd.n5017 gnd.n1804 19.3944
R9438 gnd.n5032 gnd.n1804 19.3944
R9439 gnd.n5032 gnd.n5031 19.3944
R9440 gnd.n5031 gnd.n5030 19.3944
R9441 gnd.n5030 gnd.n5023 19.3944
R9442 gnd.n5026 gnd.n5023 19.3944
R9443 gnd.n5026 gnd.n1767 19.3944
R9444 gnd.n5075 gnd.n1767 19.3944
R9445 gnd.n5075 gnd.n1765 19.3944
R9446 gnd.n5079 gnd.n1765 19.3944
R9447 gnd.n5079 gnd.n1748 19.3944
R9448 gnd.n5100 gnd.n1748 19.3944
R9449 gnd.n5100 gnd.n1746 19.3944
R9450 gnd.n5106 gnd.n1746 19.3944
R9451 gnd.n5106 gnd.n5105 19.3944
R9452 gnd.n5105 gnd.n1723 19.3944
R9453 gnd.n5138 gnd.n1723 19.3944
R9454 gnd.n5138 gnd.n1721 19.3944
R9455 gnd.n5150 gnd.n1721 19.3944
R9456 gnd.n5150 gnd.n5149 19.3944
R9457 gnd.n5149 gnd.n5148 19.3944
R9458 gnd.n5148 gnd.n5145 19.3944
R9459 gnd.n5145 gnd.n1689 19.3944
R9460 gnd.n5184 gnd.n1689 19.3944
R9461 gnd.n5184 gnd.n1687 19.3944
R9462 gnd.n5190 gnd.n1687 19.3944
R9463 gnd.n5190 gnd.n5189 19.3944
R9464 gnd.n5189 gnd.n1661 19.3944
R9465 gnd.n5219 gnd.n1661 19.3944
R9466 gnd.n5219 gnd.n1659 19.3944
R9467 gnd.n5223 gnd.n1659 19.3944
R9468 gnd.n5223 gnd.n1632 19.3944
R9469 gnd.n5256 gnd.n1632 19.3944
R9470 gnd.n5256 gnd.n1630 19.3944
R9471 gnd.n5262 gnd.n1630 19.3944
R9472 gnd.n5262 gnd.n5261 19.3944
R9473 gnd.n5261 gnd.n1532 19.3944
R9474 gnd.n5406 gnd.n1532 19.3944
R9475 gnd.n5406 gnd.n1530 19.3944
R9476 gnd.n5410 gnd.n1530 19.3944
R9477 gnd.n5410 gnd.n1519 19.3944
R9478 gnd.n5422 gnd.n1519 19.3944
R9479 gnd.n5422 gnd.n1517 19.3944
R9480 gnd.n5429 gnd.n1517 19.3944
R9481 gnd.n5429 gnd.n5428 19.3944
R9482 gnd.n5428 gnd.n1506 19.3944
R9483 gnd.n5442 gnd.n1506 19.3944
R9484 gnd.n5443 gnd.n5442 19.3944
R9485 gnd.n5443 gnd.n1504 19.3944
R9486 gnd.n5458 gnd.n1504 19.3944
R9487 gnd.n5458 gnd.n5457 19.3944
R9488 gnd.n5457 gnd.n5456 19.3944
R9489 gnd.n5456 gnd.n5449 19.3944
R9490 gnd.n5452 gnd.n5449 19.3944
R9491 gnd.n5452 gnd.n1471 19.3944
R9492 gnd.n5528 gnd.n1471 19.3944
R9493 gnd.n5528 gnd.n1469 19.3944
R9494 gnd.n5532 gnd.n1469 19.3944
R9495 gnd.n5532 gnd.n1467 19.3944
R9496 gnd.n5536 gnd.n1467 19.3944
R9497 gnd.n5536 gnd.n1465 19.3944
R9498 gnd.n5540 gnd.n1465 19.3944
R9499 gnd.n5540 gnd.n1463 19.3944
R9500 gnd.n5544 gnd.n1463 19.3944
R9501 gnd.n5544 gnd.n1461 19.3944
R9502 gnd.n5551 gnd.n1461 19.3944
R9503 gnd.n5551 gnd.n5550 19.3944
R9504 gnd.n5550 gnd.n391 19.3944
R9505 gnd.n6791 gnd.n391 19.3944
R9506 gnd.n6791 gnd.n6790 19.3944
R9507 gnd.n6790 gnd.n6789 19.3944
R9508 gnd.n6575 gnd.n518 19.3944
R9509 gnd.n6581 gnd.n518 19.3944
R9510 gnd.n6581 gnd.n516 19.3944
R9511 gnd.n6585 gnd.n516 19.3944
R9512 gnd.n6585 gnd.n512 19.3944
R9513 gnd.n6591 gnd.n512 19.3944
R9514 gnd.n6591 gnd.n510 19.3944
R9515 gnd.n6595 gnd.n510 19.3944
R9516 gnd.n6595 gnd.n506 19.3944
R9517 gnd.n6601 gnd.n506 19.3944
R9518 gnd.n6601 gnd.n504 19.3944
R9519 gnd.n6605 gnd.n504 19.3944
R9520 gnd.n6605 gnd.n500 19.3944
R9521 gnd.n6611 gnd.n500 19.3944
R9522 gnd.n6611 gnd.n498 19.3944
R9523 gnd.n6615 gnd.n498 19.3944
R9524 gnd.n6615 gnd.n494 19.3944
R9525 gnd.n6621 gnd.n494 19.3944
R9526 gnd.n6621 gnd.n492 19.3944
R9527 gnd.n6625 gnd.n492 19.3944
R9528 gnd.n6625 gnd.n488 19.3944
R9529 gnd.n6631 gnd.n488 19.3944
R9530 gnd.n6631 gnd.n486 19.3944
R9531 gnd.n6635 gnd.n486 19.3944
R9532 gnd.n6635 gnd.n482 19.3944
R9533 gnd.n6641 gnd.n482 19.3944
R9534 gnd.n6641 gnd.n480 19.3944
R9535 gnd.n6645 gnd.n480 19.3944
R9536 gnd.n6645 gnd.n476 19.3944
R9537 gnd.n6651 gnd.n476 19.3944
R9538 gnd.n6651 gnd.n474 19.3944
R9539 gnd.n6655 gnd.n474 19.3944
R9540 gnd.n6655 gnd.n470 19.3944
R9541 gnd.n6661 gnd.n470 19.3944
R9542 gnd.n6661 gnd.n468 19.3944
R9543 gnd.n6665 gnd.n468 19.3944
R9544 gnd.n6665 gnd.n464 19.3944
R9545 gnd.n6671 gnd.n464 19.3944
R9546 gnd.n6671 gnd.n462 19.3944
R9547 gnd.n6675 gnd.n462 19.3944
R9548 gnd.n6675 gnd.n458 19.3944
R9549 gnd.n6681 gnd.n458 19.3944
R9550 gnd.n6681 gnd.n456 19.3944
R9551 gnd.n6685 gnd.n456 19.3944
R9552 gnd.n6685 gnd.n452 19.3944
R9553 gnd.n6691 gnd.n452 19.3944
R9554 gnd.n6691 gnd.n450 19.3944
R9555 gnd.n6695 gnd.n450 19.3944
R9556 gnd.n6695 gnd.n446 19.3944
R9557 gnd.n6701 gnd.n446 19.3944
R9558 gnd.n6701 gnd.n444 19.3944
R9559 gnd.n6705 gnd.n444 19.3944
R9560 gnd.n6705 gnd.n440 19.3944
R9561 gnd.n6711 gnd.n440 19.3944
R9562 gnd.n6711 gnd.n438 19.3944
R9563 gnd.n6715 gnd.n438 19.3944
R9564 gnd.n6715 gnd.n434 19.3944
R9565 gnd.n6721 gnd.n434 19.3944
R9566 gnd.n6721 gnd.n432 19.3944
R9567 gnd.n6725 gnd.n432 19.3944
R9568 gnd.n6725 gnd.n428 19.3944
R9569 gnd.n6731 gnd.n428 19.3944
R9570 gnd.n6731 gnd.n426 19.3944
R9571 gnd.n6735 gnd.n426 19.3944
R9572 gnd.n6735 gnd.n422 19.3944
R9573 gnd.n6741 gnd.n422 19.3944
R9574 gnd.n6741 gnd.n420 19.3944
R9575 gnd.n6745 gnd.n420 19.3944
R9576 gnd.n6745 gnd.n416 19.3944
R9577 gnd.n6751 gnd.n416 19.3944
R9578 gnd.n6751 gnd.n414 19.3944
R9579 gnd.n6755 gnd.n414 19.3944
R9580 gnd.n6755 gnd.n410 19.3944
R9581 gnd.n6761 gnd.n410 19.3944
R9582 gnd.n6761 gnd.n408 19.3944
R9583 gnd.n6765 gnd.n408 19.3944
R9584 gnd.n6765 gnd.n404 19.3944
R9585 gnd.n6771 gnd.n404 19.3944
R9586 gnd.n6771 gnd.n402 19.3944
R9587 gnd.n6775 gnd.n402 19.3944
R9588 gnd.n6775 gnd.n398 19.3944
R9589 gnd.n6782 gnd.n398 19.3944
R9590 gnd.n6782 gnd.n396 19.3944
R9591 gnd.n6786 gnd.n396 19.3944
R9592 gnd.n6254 gnd.n713 19.3944
R9593 gnd.n6254 gnd.n709 19.3944
R9594 gnd.n6260 gnd.n709 19.3944
R9595 gnd.n6260 gnd.n707 19.3944
R9596 gnd.n6264 gnd.n707 19.3944
R9597 gnd.n6264 gnd.n703 19.3944
R9598 gnd.n6270 gnd.n703 19.3944
R9599 gnd.n6270 gnd.n701 19.3944
R9600 gnd.n6274 gnd.n701 19.3944
R9601 gnd.n6274 gnd.n697 19.3944
R9602 gnd.n6280 gnd.n697 19.3944
R9603 gnd.n6280 gnd.n695 19.3944
R9604 gnd.n6284 gnd.n695 19.3944
R9605 gnd.n6284 gnd.n691 19.3944
R9606 gnd.n6290 gnd.n691 19.3944
R9607 gnd.n6290 gnd.n689 19.3944
R9608 gnd.n6294 gnd.n689 19.3944
R9609 gnd.n6294 gnd.n685 19.3944
R9610 gnd.n6300 gnd.n685 19.3944
R9611 gnd.n6300 gnd.n683 19.3944
R9612 gnd.n6304 gnd.n683 19.3944
R9613 gnd.n6304 gnd.n679 19.3944
R9614 gnd.n6310 gnd.n679 19.3944
R9615 gnd.n6310 gnd.n677 19.3944
R9616 gnd.n6314 gnd.n677 19.3944
R9617 gnd.n6314 gnd.n673 19.3944
R9618 gnd.n6320 gnd.n673 19.3944
R9619 gnd.n6320 gnd.n671 19.3944
R9620 gnd.n6324 gnd.n671 19.3944
R9621 gnd.n6324 gnd.n667 19.3944
R9622 gnd.n6330 gnd.n667 19.3944
R9623 gnd.n6330 gnd.n665 19.3944
R9624 gnd.n6334 gnd.n665 19.3944
R9625 gnd.n6334 gnd.n661 19.3944
R9626 gnd.n6340 gnd.n661 19.3944
R9627 gnd.n6340 gnd.n659 19.3944
R9628 gnd.n6344 gnd.n659 19.3944
R9629 gnd.n6344 gnd.n655 19.3944
R9630 gnd.n6350 gnd.n655 19.3944
R9631 gnd.n6350 gnd.n653 19.3944
R9632 gnd.n6354 gnd.n653 19.3944
R9633 gnd.n6354 gnd.n649 19.3944
R9634 gnd.n6360 gnd.n649 19.3944
R9635 gnd.n6360 gnd.n647 19.3944
R9636 gnd.n6364 gnd.n647 19.3944
R9637 gnd.n6364 gnd.n643 19.3944
R9638 gnd.n6370 gnd.n643 19.3944
R9639 gnd.n6370 gnd.n641 19.3944
R9640 gnd.n6374 gnd.n641 19.3944
R9641 gnd.n6374 gnd.n637 19.3944
R9642 gnd.n6380 gnd.n637 19.3944
R9643 gnd.n6380 gnd.n635 19.3944
R9644 gnd.n6384 gnd.n635 19.3944
R9645 gnd.n6384 gnd.n631 19.3944
R9646 gnd.n6390 gnd.n631 19.3944
R9647 gnd.n6390 gnd.n629 19.3944
R9648 gnd.n6394 gnd.n629 19.3944
R9649 gnd.n6394 gnd.n625 19.3944
R9650 gnd.n6400 gnd.n625 19.3944
R9651 gnd.n6400 gnd.n623 19.3944
R9652 gnd.n6404 gnd.n623 19.3944
R9653 gnd.n6404 gnd.n619 19.3944
R9654 gnd.n6410 gnd.n619 19.3944
R9655 gnd.n6410 gnd.n617 19.3944
R9656 gnd.n6414 gnd.n617 19.3944
R9657 gnd.n6414 gnd.n613 19.3944
R9658 gnd.n6420 gnd.n613 19.3944
R9659 gnd.n6420 gnd.n611 19.3944
R9660 gnd.n6424 gnd.n611 19.3944
R9661 gnd.n6424 gnd.n607 19.3944
R9662 gnd.n6430 gnd.n607 19.3944
R9663 gnd.n6430 gnd.n605 19.3944
R9664 gnd.n6434 gnd.n605 19.3944
R9665 gnd.n6434 gnd.n601 19.3944
R9666 gnd.n6440 gnd.n601 19.3944
R9667 gnd.n6440 gnd.n599 19.3944
R9668 gnd.n6444 gnd.n599 19.3944
R9669 gnd.n6444 gnd.n595 19.3944
R9670 gnd.n6450 gnd.n595 19.3944
R9671 gnd.n6450 gnd.n593 19.3944
R9672 gnd.n6454 gnd.n593 19.3944
R9673 gnd.n6454 gnd.n589 19.3944
R9674 gnd.n6460 gnd.n589 19.3944
R9675 gnd.n6460 gnd.n587 19.3944
R9676 gnd.n6464 gnd.n587 19.3944
R9677 gnd.n6464 gnd.n583 19.3944
R9678 gnd.n6470 gnd.n583 19.3944
R9679 gnd.n6470 gnd.n581 19.3944
R9680 gnd.n6474 gnd.n581 19.3944
R9681 gnd.n6474 gnd.n577 19.3944
R9682 gnd.n6480 gnd.n577 19.3944
R9683 gnd.n6480 gnd.n575 19.3944
R9684 gnd.n6484 gnd.n575 19.3944
R9685 gnd.n6484 gnd.n571 19.3944
R9686 gnd.n6490 gnd.n571 19.3944
R9687 gnd.n6490 gnd.n569 19.3944
R9688 gnd.n6494 gnd.n569 19.3944
R9689 gnd.n6494 gnd.n565 19.3944
R9690 gnd.n6500 gnd.n565 19.3944
R9691 gnd.n6500 gnd.n563 19.3944
R9692 gnd.n6504 gnd.n563 19.3944
R9693 gnd.n6504 gnd.n559 19.3944
R9694 gnd.n6510 gnd.n559 19.3944
R9695 gnd.n6510 gnd.n557 19.3944
R9696 gnd.n6514 gnd.n557 19.3944
R9697 gnd.n6514 gnd.n553 19.3944
R9698 gnd.n6520 gnd.n553 19.3944
R9699 gnd.n6520 gnd.n551 19.3944
R9700 gnd.n6524 gnd.n551 19.3944
R9701 gnd.n6524 gnd.n547 19.3944
R9702 gnd.n6530 gnd.n547 19.3944
R9703 gnd.n6530 gnd.n545 19.3944
R9704 gnd.n6534 gnd.n545 19.3944
R9705 gnd.n6534 gnd.n541 19.3944
R9706 gnd.n6540 gnd.n541 19.3944
R9707 gnd.n6540 gnd.n539 19.3944
R9708 gnd.n6544 gnd.n539 19.3944
R9709 gnd.n6544 gnd.n535 19.3944
R9710 gnd.n6550 gnd.n535 19.3944
R9711 gnd.n6550 gnd.n533 19.3944
R9712 gnd.n6554 gnd.n533 19.3944
R9713 gnd.n6554 gnd.n529 19.3944
R9714 gnd.n6560 gnd.n529 19.3944
R9715 gnd.n6560 gnd.n527 19.3944
R9716 gnd.n6565 gnd.n527 19.3944
R9717 gnd.n6565 gnd.n523 19.3944
R9718 gnd.n6571 gnd.n523 19.3944
R9719 gnd.n6572 gnd.n6571 19.3944
R9720 gnd.n6250 gnd.n715 19.3944
R9721 gnd.n6244 gnd.n715 19.3944
R9722 gnd.n6244 gnd.n6243 19.3944
R9723 gnd.n6243 gnd.n6242 19.3944
R9724 gnd.n6242 gnd.n722 19.3944
R9725 gnd.n6236 gnd.n722 19.3944
R9726 gnd.n6236 gnd.n6235 19.3944
R9727 gnd.n6235 gnd.n6234 19.3944
R9728 gnd.n6234 gnd.n730 19.3944
R9729 gnd.n6228 gnd.n730 19.3944
R9730 gnd.n6228 gnd.n6227 19.3944
R9731 gnd.n6227 gnd.n6226 19.3944
R9732 gnd.n6226 gnd.n738 19.3944
R9733 gnd.n6220 gnd.n738 19.3944
R9734 gnd.n6220 gnd.n6219 19.3944
R9735 gnd.n6219 gnd.n6218 19.3944
R9736 gnd.n6218 gnd.n746 19.3944
R9737 gnd.n6212 gnd.n746 19.3944
R9738 gnd.n6212 gnd.n6211 19.3944
R9739 gnd.n6211 gnd.n6210 19.3944
R9740 gnd.n6210 gnd.n754 19.3944
R9741 gnd.n6204 gnd.n754 19.3944
R9742 gnd.n6204 gnd.n6203 19.3944
R9743 gnd.n6203 gnd.n6202 19.3944
R9744 gnd.n6202 gnd.n762 19.3944
R9745 gnd.n6196 gnd.n762 19.3944
R9746 gnd.n6196 gnd.n6195 19.3944
R9747 gnd.n6195 gnd.n6194 19.3944
R9748 gnd.n6194 gnd.n770 19.3944
R9749 gnd.n6188 gnd.n770 19.3944
R9750 gnd.n6188 gnd.n6187 19.3944
R9751 gnd.n6187 gnd.n6186 19.3944
R9752 gnd.n6186 gnd.n778 19.3944
R9753 gnd.n6180 gnd.n778 19.3944
R9754 gnd.n6180 gnd.n6179 19.3944
R9755 gnd.n6179 gnd.n6178 19.3944
R9756 gnd.n6178 gnd.n786 19.3944
R9757 gnd.n6172 gnd.n786 19.3944
R9758 gnd.n6172 gnd.n6171 19.3944
R9759 gnd.n6171 gnd.n6170 19.3944
R9760 gnd.n6170 gnd.n794 19.3944
R9761 gnd.n6164 gnd.n794 19.3944
R9762 gnd.n6164 gnd.n6163 19.3944
R9763 gnd.n6163 gnd.n6162 19.3944
R9764 gnd.n6162 gnd.n802 19.3944
R9765 gnd.n6156 gnd.n802 19.3944
R9766 gnd.n6156 gnd.n6155 19.3944
R9767 gnd.n6155 gnd.n6154 19.3944
R9768 gnd.n6154 gnd.n810 19.3944
R9769 gnd.n6148 gnd.n810 19.3944
R9770 gnd.n6148 gnd.n6147 19.3944
R9771 gnd.n6147 gnd.n6146 19.3944
R9772 gnd.n6146 gnd.n818 19.3944
R9773 gnd.n6140 gnd.n818 19.3944
R9774 gnd.n6140 gnd.n6139 19.3944
R9775 gnd.n6139 gnd.n6138 19.3944
R9776 gnd.n6138 gnd.n826 19.3944
R9777 gnd.n6132 gnd.n826 19.3944
R9778 gnd.n6132 gnd.n6131 19.3944
R9779 gnd.n6131 gnd.n6130 19.3944
R9780 gnd.n6130 gnd.n834 19.3944
R9781 gnd.n6124 gnd.n834 19.3944
R9782 gnd.n6124 gnd.n6123 19.3944
R9783 gnd.n6123 gnd.n6122 19.3944
R9784 gnd.n6122 gnd.n842 19.3944
R9785 gnd.n6116 gnd.n842 19.3944
R9786 gnd.n6116 gnd.n6115 19.3944
R9787 gnd.n6115 gnd.n6114 19.3944
R9788 gnd.n6114 gnd.n850 19.3944
R9789 gnd.n6108 gnd.n850 19.3944
R9790 gnd.n6108 gnd.n6107 19.3944
R9791 gnd.n6107 gnd.n6106 19.3944
R9792 gnd.n6106 gnd.n858 19.3944
R9793 gnd.n6100 gnd.n858 19.3944
R9794 gnd.n6100 gnd.n6099 19.3944
R9795 gnd.n6099 gnd.n6098 19.3944
R9796 gnd.n6098 gnd.n866 19.3944
R9797 gnd.n6092 gnd.n866 19.3944
R9798 gnd.n6092 gnd.n6091 19.3944
R9799 gnd.n6091 gnd.n6090 19.3944
R9800 gnd.n6090 gnd.n874 19.3944
R9801 gnd.n6084 gnd.n874 19.3944
R9802 gnd.n6084 gnd.n6083 19.3944
R9803 gnd.n6083 gnd.n6082 19.3944
R9804 gnd.n4350 gnd.n4342 19.3944
R9805 gnd.n4346 gnd.n4342 19.3944
R9806 gnd.n4346 gnd.n4345 19.3944
R9807 gnd.n4345 gnd.n1988 19.3944
R9808 gnd.n4686 gnd.n1988 19.3944
R9809 gnd.n4686 gnd.n1986 19.3944
R9810 gnd.n4690 gnd.n1986 19.3944
R9811 gnd.n4690 gnd.n1984 19.3944
R9812 gnd.n4694 gnd.n1984 19.3944
R9813 gnd.n4694 gnd.n1981 19.3944
R9814 gnd.n4839 gnd.n1981 19.3944
R9815 gnd.n4839 gnd.n1982 19.3944
R9816 gnd.n4835 gnd.n1982 19.3944
R9817 gnd.n4835 gnd.n4834 19.3944
R9818 gnd.n4834 gnd.n4833 19.3944
R9819 gnd.n4833 gnd.n4699 19.3944
R9820 gnd.n4829 gnd.n4699 19.3944
R9821 gnd.n4829 gnd.n4828 19.3944
R9822 gnd.n4828 gnd.n4827 19.3944
R9823 gnd.n4827 gnd.n4702 19.3944
R9824 gnd.n4823 gnd.n4702 19.3944
R9825 gnd.n4823 gnd.n4822 19.3944
R9826 gnd.n4822 gnd.n4821 19.3944
R9827 gnd.n4821 gnd.n4708 19.3944
R9828 gnd.n4817 gnd.n4708 19.3944
R9829 gnd.n4817 gnd.n4816 19.3944
R9830 gnd.n4816 gnd.n4815 19.3944
R9831 gnd.n4815 gnd.n4712 19.3944
R9832 gnd.n4811 gnd.n4712 19.3944
R9833 gnd.n4811 gnd.n4810 19.3944
R9834 gnd.n4810 gnd.n4809 19.3944
R9835 gnd.n4809 gnd.n4716 19.3944
R9836 gnd.n4805 gnd.n4716 19.3944
R9837 gnd.n4805 gnd.n4804 19.3944
R9838 gnd.n4804 gnd.n4803 19.3944
R9839 gnd.n4803 gnd.n4719 19.3944
R9840 gnd.n4799 gnd.n4719 19.3944
R9841 gnd.n4799 gnd.n4798 19.3944
R9842 gnd.n4798 gnd.n4797 19.3944
R9843 gnd.n4797 gnd.n4725 19.3944
R9844 gnd.n4793 gnd.n4725 19.3944
R9845 gnd.n4793 gnd.n4792 19.3944
R9846 gnd.n4792 gnd.n4791 19.3944
R9847 gnd.n4791 gnd.n4728 19.3944
R9848 gnd.n4787 gnd.n4728 19.3944
R9849 gnd.n4787 gnd.n4786 19.3944
R9850 gnd.n4786 gnd.n4785 19.3944
R9851 gnd.n4785 gnd.n4732 19.3944
R9852 gnd.n4781 gnd.n4732 19.3944
R9853 gnd.n4781 gnd.n4780 19.3944
R9854 gnd.n4780 gnd.n4779 19.3944
R9855 gnd.n4779 gnd.n4737 19.3944
R9856 gnd.n4775 gnd.n4737 19.3944
R9857 gnd.n4775 gnd.n4774 19.3944
R9858 gnd.n4774 gnd.n4773 19.3944
R9859 gnd.n4773 gnd.n4741 19.3944
R9860 gnd.n4769 gnd.n4741 19.3944
R9861 gnd.n4769 gnd.n4768 19.3944
R9862 gnd.n4768 gnd.n4767 19.3944
R9863 gnd.n4767 gnd.n4746 19.3944
R9864 gnd.n4763 gnd.n4746 19.3944
R9865 gnd.n4763 gnd.n4762 19.3944
R9866 gnd.n4762 gnd.n4761 19.3944
R9867 gnd.n4761 gnd.n4751 19.3944
R9868 gnd.n4757 gnd.n4751 19.3944
R9869 gnd.n4757 gnd.n4756 19.3944
R9870 gnd.n4756 gnd.n4755 19.3944
R9871 gnd.n4755 gnd.n1623 19.3944
R9872 gnd.n5266 gnd.n1623 19.3944
R9873 gnd.n5266 gnd.n1620 19.3944
R9874 gnd.n5271 gnd.n1620 19.3944
R9875 gnd.n5271 gnd.n1621 19.3944
R9876 gnd.n1621 gnd.n1524 19.3944
R9877 gnd.n5414 gnd.n1524 19.3944
R9878 gnd.n5414 gnd.n1522 19.3944
R9879 gnd.n5418 gnd.n1522 19.3944
R9880 gnd.n5418 gnd.n1512 19.3944
R9881 gnd.n5433 gnd.n1512 19.3944
R9882 gnd.n5433 gnd.n1510 19.3944
R9883 gnd.n5437 gnd.n1510 19.3944
R9884 gnd.n5437 gnd.n1224 19.3944
R9885 gnd.n5779 gnd.n1224 19.3944
R9886 gnd.n5776 gnd.n5775 19.3944
R9887 gnd.n5775 gnd.n5774 19.3944
R9888 gnd.n5774 gnd.n1229 19.3944
R9889 gnd.n5770 gnd.n1229 19.3944
R9890 gnd.n5770 gnd.n5769 19.3944
R9891 gnd.n5769 gnd.n5768 19.3944
R9892 gnd.n5768 gnd.n1234 19.3944
R9893 gnd.n5763 gnd.n1234 19.3944
R9894 gnd.n5763 gnd.n5762 19.3944
R9895 gnd.n5762 gnd.n1239 19.3944
R9896 gnd.n5755 gnd.n1239 19.3944
R9897 gnd.n5755 gnd.n5754 19.3944
R9898 gnd.n5754 gnd.n1248 19.3944
R9899 gnd.n5747 gnd.n1248 19.3944
R9900 gnd.n5747 gnd.n5746 19.3944
R9901 gnd.n5746 gnd.n1256 19.3944
R9902 gnd.n5739 gnd.n1256 19.3944
R9903 gnd.n5739 gnd.n5738 19.3944
R9904 gnd.n5738 gnd.n1264 19.3944
R9905 gnd.n5731 gnd.n1264 19.3944
R9906 gnd.n5731 gnd.n5730 19.3944
R9907 gnd.n5730 gnd.n1272 19.3944
R9908 gnd.n5723 gnd.n1272 19.3944
R9909 gnd.n5723 gnd.n5722 19.3944
R9910 gnd.n1498 gnd.n1477 19.3944
R9911 gnd.n5464 gnd.n1477 19.3944
R9912 gnd.n5464 gnd.n5463 19.3944
R9913 gnd.n2244 gnd.n876 19.1949
R9914 gnd.n1863 gnd.t4 19.1199
R9915 gnd.n1844 gnd.n1836 19.1199
R9916 gnd.n1795 gnd.n1793 19.1199
R9917 gnd.n1763 gnd.n1755 19.1199
R9918 gnd.n1712 gnd.n1711 19.1199
R9919 gnd.n1695 gnd.t52 19.1199
R9920 gnd.n7041 gnd.n157 19.1199
R9921 gnd.n3109 gnd.t21 18.8012
R9922 gnd.n3094 gnd.t41 18.8012
R9923 gnd.n2953 gnd.n2952 18.4825
R9924 gnd.n5661 gnd.n5660 18.4247
R9925 gnd.n5974 gnd.n5973 18.4247
R9926 gnd.n5903 gnd.n5902 18.2639
R9927 gnd.n5399 gnd.n1561 18.2639
R9928 gnd.n5719 gnd.n5718 18.2308
R9929 gnd.n7018 gnd.n6969 18.2308
R9930 gnd.n4432 gnd.n2036 18.2308
R9931 gnd.n3883 gnd.n3843 18.2308
R9932 gnd.t20 gnd.n2633 18.1639
R9933 gnd.t11 gnd.n1114 18.1639
R9934 gnd.n5274 gnd.t9 18.1639
R9935 gnd.n1904 gnd.n1125 17.8452
R9936 gnd.n4911 gnd.n1879 17.8452
R9937 gnd.n5035 gnd.n1799 17.8452
R9938 gnd.n5097 gnd.n1741 17.8452
R9939 gnd.n5217 gnd.n1666 17.8452
R9940 gnd.t124 gnd.n1625 17.8452
R9941 gnd.n5264 gnd.n1626 17.8452
R9942 gnd.n2661 gnd.t7 17.5266
R9943 gnd.n2218 gnd.t256 17.5266
R9944 gnd.t31 gnd.n1823 17.5266
R9945 gnd.n4735 gnd.t174 17.5266
R9946 gnd.n182 gnd.t196 17.5266
R9947 gnd.n3060 gnd.t181 16.8893
R9948 gnd.n2181 gnd.t209 16.8893
R9949 gnd.t251 gnd.n918 16.8893
R9950 gnd.n5553 gnd.t217 16.8893
R9951 gnd.n144 gnd.t223 16.8893
R9952 gnd.n7111 gnd.n7108 16.6793
R9953 gnd.n5643 gnd.n5640 16.6793
R9954 gnd.n3963 gnd.n3960 16.6793
R9955 gnd.n4524 gnd.n4523 16.6793
R9956 gnd.n4883 gnd.n4882 16.5706
R9957 gnd.n4994 gnd.n1819 16.5706
R9958 gnd.n5007 gnd.n5005 16.5706
R9959 gnd.n5116 gnd.n1737 16.5706
R9960 gnd.n5128 gnd.n5127 16.5706
R9961 gnd.n1656 gnd.n1649 16.5706
R9962 gnd.n5254 gnd.n5253 16.5706
R9963 gnd.n2888 gnd.t58 16.2519
R9964 gnd.n2588 gnd.t194 16.2519
R9965 gnd.n4168 gnd.t242 16.2519
R9966 gnd.t290 gnd.n2083 16.2519
R9967 gnd.n4642 gnd.t84 16.2519
R9968 gnd.t101 gnd.n1219 16.2519
R9969 gnd.n6865 gnd.t266 16.2519
R9970 gnd.n106 gnd.t286 16.2519
R9971 gnd.t357 gnd.n4923 15.9333
R9972 gnd.n1684 gnd.t173 15.9333
R9973 gnd.n3575 gnd.n3573 15.6674
R9974 gnd.n3543 gnd.n3541 15.6674
R9975 gnd.n3511 gnd.n3509 15.6674
R9976 gnd.n3480 gnd.n3478 15.6674
R9977 gnd.n3448 gnd.n3446 15.6674
R9978 gnd.n3416 gnd.n3414 15.6674
R9979 gnd.n3384 gnd.n3382 15.6674
R9980 gnd.n3353 gnd.n3351 15.6674
R9981 gnd.n2879 gnd.t58 15.6146
R9982 gnd.t54 gnd.n2326 15.6146
R9983 gnd.t170 gnd.n2327 15.6146
R9984 gnd.n4183 gnd.t242 15.6146
R9985 gnd.n4234 gnd.t290 15.6146
R9986 gnd.t84 gnd.n1999 15.6146
R9987 gnd.n5439 gnd.t101 15.6146
R9988 gnd.n6874 gnd.t266 15.6146
R9989 gnd.n7257 gnd.t286 15.6146
R9990 gnd.n7066 gnd.n305 15.3217
R9991 gnd.n5600 gnd.n5595 15.3217
R9992 gnd.n3921 gnd.n2242 15.3217
R9993 gnd.n4575 gnd.n4573 15.3217
R9994 gnd.n4863 gnd.n4862 15.296
R9995 gnd.n5253 gnd.n1637 15.296
R9996 gnd.n1546 gnd.n1545 15.0827
R9997 gnd.n1096 gnd.n1091 15.0481
R9998 gnd.n1556 gnd.n1555 15.0481
R9999 gnd.n3247 gnd.t185 14.9773
R10000 gnd.n4123 gnd.t209 14.9773
R10001 gnd.n6073 gnd.t211 14.9773
R10002 gnd.n6817 gnd.t237 14.9773
R10003 gnd.n7233 gnd.t223 14.9773
R10004 gnd.n4892 gnd.t193 14.6587
R10005 gnd.n5225 gnd.t47 14.6587
R10006 gnd.t37 gnd.n2369 14.34
R10007 gnd.n3325 gnd.t8 14.34
R10008 gnd.n4077 gnd.t256 14.34
R10009 gnd.n6049 gnd.t221 14.34
R10010 gnd.n5489 gnd.t228 14.34
R10011 gnd.n7209 gnd.t196 14.34
R10012 gnd.n5891 gnd.n1125 14.0214
R10013 gnd.n4911 gnd.t5 14.0214
R10014 gnd.n4976 gnd.n4974 14.0214
R10015 gnd.n5035 gnd.n5034 14.0214
R10016 gnd.n5098 gnd.n5097 14.0214
R10017 gnd.n5153 gnd.n5152 14.0214
R10018 gnd.t189 gnd.n5217 14.0214
R10019 gnd.n3035 gnd.t179 13.7027
R10020 gnd.n4872 gnd.t358 13.7027
R10021 gnd.t15 gnd.n1634 13.7027
R10022 gnd.n2745 gnd.n2744 13.5763
R10023 gnd.n3689 gnd.n2282 13.5763
R10024 gnd.n2953 gnd.n2691 13.384
R10025 gnd.n4842 gnd.t105 13.384
R10026 gnd.t108 gnd.n1626 13.384
R10027 gnd.n1107 gnd.n1088 13.1884
R10028 gnd.n1102 gnd.n1101 13.1884
R10029 gnd.n1101 gnd.n1100 13.1884
R10030 gnd.n1549 gnd.n1544 13.1884
R10031 gnd.n1550 gnd.n1549 13.1884
R10032 gnd.n1103 gnd.n1090 13.146
R10033 gnd.n1099 gnd.n1090 13.146
R10034 gnd.n1548 gnd.n1547 13.146
R10035 gnd.n1548 gnd.n1543 13.146
R10036 gnd.n3576 gnd.n3572 12.8005
R10037 gnd.n3544 gnd.n3540 12.8005
R10038 gnd.n3512 gnd.n3508 12.8005
R10039 gnd.n3481 gnd.n3477 12.8005
R10040 gnd.n3449 gnd.n3445 12.8005
R10041 gnd.n3417 gnd.n3413 12.8005
R10042 gnd.n3385 gnd.n3381 12.8005
R10043 gnd.n3354 gnd.n3350 12.8005
R10044 gnd.n5897 gnd.n1114 12.7467
R10045 gnd.n1874 gnd.n1869 12.7467
R10046 gnd.n4958 gnd.n1844 12.7467
R10047 gnd.n1793 gnd.n1788 12.7467
R10048 gnd.n5048 gnd.t28 12.7467
R10049 gnd.n5082 gnd.t13 12.7467
R10050 gnd.n5081 gnd.n1763 12.7467
R10051 gnd.n1711 gnd.n1706 12.7467
R10052 gnd.n1677 gnd.n1675 12.7467
R10053 gnd.n7221 gnd.n157 12.7467
R10054 gnd.t50 gnd.n1874 12.4281
R10055 gnd.n1675 gnd.t0 12.4281
R10056 gnd.n2744 gnd.n2739 12.4126
R10057 gnd.n3692 gnd.n3689 12.4126
R10058 gnd.n5966 gnd.n5903 12.1761
R10059 gnd.n1562 gnd.n1561 12.1761
R10060 gnd.n3580 gnd.n3579 12.0247
R10061 gnd.n3548 gnd.n3547 12.0247
R10062 gnd.n3516 gnd.n3515 12.0247
R10063 gnd.n3485 gnd.n3484 12.0247
R10064 gnd.n3453 gnd.n3452 12.0247
R10065 gnd.n3421 gnd.n3420 12.0247
R10066 gnd.n3389 gnd.n3388 12.0247
R10067 gnd.n3358 gnd.n3357 12.0247
R10068 gnd.t91 gnd.n968 11.7908
R10069 gnd.n5526 gnd.t62 11.7908
R10070 gnd.n4930 gnd.n1864 11.4721
R10071 gnd.n4950 gnd.n4948 11.4721
R10072 gnd.n5054 gnd.n1784 11.4721
R10073 gnd.n5073 gnd.n5072 11.4721
R10074 gnd.n5174 gnd.n1701 11.4721
R10075 gnd.n5193 gnd.n1681 11.4721
R10076 gnd.n5404 gnd.t127 11.4721
R10077 gnd.n5412 gnd.n1526 11.4721
R10078 gnd.n3583 gnd.n3570 11.249
R10079 gnd.n3551 gnd.n3538 11.249
R10080 gnd.n3519 gnd.n3506 11.249
R10081 gnd.n3488 gnd.n3475 11.249
R10082 gnd.n3456 gnd.n3443 11.249
R10083 gnd.n3424 gnd.n3411 11.249
R10084 gnd.n3392 gnd.n3379 11.249
R10085 gnd.n3361 gnd.n3348 11.249
R10086 gnd.n3023 gnd.t179 11.1535
R10087 gnd.n1991 gnd.t362 11.1535
R10088 gnd.n5420 gnd.t26 11.1535
R10089 gnd.n4271 gnd.n886 10.8348
R10090 gnd.n6073 gnd.n896 10.8348
R10091 gnd.n4291 gnd.n4290 10.8348
R10092 gnd.n6067 gnd.n907 10.8348
R10093 gnd.n4282 gnd.n910 10.8348
R10094 gnd.n6061 gnd.n918 10.8348
R10095 gnd.n4316 gnd.n921 10.8348
R10096 gnd.n4324 gnd.n930 10.8348
R10097 gnd.n6049 gnd.n938 10.8348
R10098 gnd.n4597 gnd.n4596 10.8348
R10099 gnd.n6043 gnd.n947 10.8348
R10100 gnd.n4331 gnd.n950 10.8348
R10101 gnd.n6037 gnd.n958 10.8348
R10102 gnd.n4583 gnd.n961 10.8348
R10103 gnd.n6031 gnd.n968 10.8348
R10104 gnd.n4623 gnd.n971 10.8348
R10105 gnd.n4862 gnd.t88 10.8348
R10106 gnd.n4935 gnd.t18 10.8348
R10107 gnd.n4959 gnd.t18 10.8348
R10108 gnd.n5166 gnd.t14 10.8348
R10109 gnd.t14 gnd.n5165 10.8348
R10110 gnd.t81 gnd.n1526 10.8348
R10111 gnd.n5592 gnd.n1400 10.8348
R10112 gnd.n5526 gnd.n5525 10.8348
R10113 gnd.n5586 gnd.n1410 10.8348
R10114 gnd.n5480 gnd.n1422 10.8348
R10115 gnd.n5580 gnd.n1425 10.8348
R10116 gnd.n5484 gnd.n1432 10.8348
R10117 gnd.n5574 gnd.n1435 10.8348
R10118 gnd.n5489 gnd.n1443 10.8348
R10119 gnd.n5568 gnd.n1446 10.8348
R10120 gnd.n5562 gnd.n1456 10.8348
R10121 gnd.n5554 gnd.n5553 10.8348
R10122 gnd.n5502 gnd.n379 10.8348
R10123 gnd.n6807 gnd.n382 10.8348
R10124 gnd.n6794 gnd.n6793 10.8348
R10125 gnd.n6817 gnd.n371 10.8348
R10126 gnd.n6800 gnd.n363 10.8348
R10127 gnd.n7069 gnd.n7066 10.6672
R10128 gnd.n5603 gnd.n5600 10.6672
R10129 gnd.n3923 gnd.n3921 10.6672
R10130 gnd.n4573 gnd.n4572 10.6672
R10131 gnd.n5334 gnd.n1589 10.6151
R10132 gnd.n5334 gnd.n5333 10.6151
R10133 gnd.n5331 gnd.n1593 10.6151
R10134 gnd.n5326 gnd.n1593 10.6151
R10135 gnd.n5326 gnd.n5325 10.6151
R10136 gnd.n5325 gnd.n5324 10.6151
R10137 gnd.n5324 gnd.n1596 10.6151
R10138 gnd.n5319 gnd.n1596 10.6151
R10139 gnd.n5319 gnd.n5318 10.6151
R10140 gnd.n5318 gnd.n5317 10.6151
R10141 gnd.n5317 gnd.n1599 10.6151
R10142 gnd.n5312 gnd.n1599 10.6151
R10143 gnd.n5312 gnd.n5311 10.6151
R10144 gnd.n5311 gnd.n5310 10.6151
R10145 gnd.n5310 gnd.n1602 10.6151
R10146 gnd.n5305 gnd.n1602 10.6151
R10147 gnd.n5305 gnd.n5304 10.6151
R10148 gnd.n5304 gnd.n5303 10.6151
R10149 gnd.n5303 gnd.n1605 10.6151
R10150 gnd.n5298 gnd.n1605 10.6151
R10151 gnd.n5298 gnd.n5297 10.6151
R10152 gnd.n5297 gnd.n5296 10.6151
R10153 gnd.n5296 gnd.n1608 10.6151
R10154 gnd.n5291 gnd.n1608 10.6151
R10155 gnd.n5291 gnd.n5290 10.6151
R10156 gnd.n5290 gnd.n5289 10.6151
R10157 gnd.n5289 gnd.n1611 10.6151
R10158 gnd.n5284 gnd.n1611 10.6151
R10159 gnd.n5284 gnd.n5283 10.6151
R10160 gnd.n5283 gnd.n5282 10.6151
R10161 gnd.n1976 gnd.n1975 10.6151
R10162 gnd.n1977 gnd.n1976 10.6151
R10163 gnd.n1978 gnd.n1977 10.6151
R10164 gnd.n1978 gnd.n1907 10.6151
R10165 gnd.n4851 gnd.n1907 10.6151
R10166 gnd.n4852 gnd.n4851 10.6151
R10167 gnd.n4854 gnd.n4852 10.6151
R10168 gnd.n4854 gnd.n4853 10.6151
R10169 gnd.n4853 gnd.n1896 10.6151
R10170 gnd.n4874 gnd.n1896 10.6151
R10171 gnd.n4875 gnd.n4874 10.6151
R10172 gnd.n4880 gnd.n4875 10.6151
R10173 gnd.n4880 gnd.n4879 10.6151
R10174 gnd.n4879 gnd.n4878 10.6151
R10175 gnd.n4878 gnd.n4876 10.6151
R10176 gnd.n4876 gnd.n1871 10.6151
R10177 gnd.n4919 gnd.n1871 10.6151
R10178 gnd.n4920 gnd.n4919 10.6151
R10179 gnd.n4921 gnd.n4920 10.6151
R10180 gnd.n4921 gnd.n1860 10.6151
R10181 gnd.n4932 gnd.n1860 10.6151
R10182 gnd.n4933 gnd.n4932 10.6151
R10183 gnd.n4940 gnd.n4933 10.6151
R10184 gnd.n4940 gnd.n4939 10.6151
R10185 gnd.n4939 gnd.n4938 10.6151
R10186 gnd.n4938 gnd.n4937 10.6151
R10187 gnd.n4937 gnd.n4934 10.6151
R10188 gnd.n4934 gnd.n1834 10.6151
R10189 gnd.n4968 gnd.n1834 10.6151
R10190 gnd.n4969 gnd.n4968 10.6151
R10191 gnd.n4972 gnd.n4969 10.6151
R10192 gnd.n4972 gnd.n4971 10.6151
R10193 gnd.n4971 gnd.n4970 10.6151
R10194 gnd.n4970 gnd.n1817 10.6151
R10195 gnd.n4997 gnd.n1817 10.6151
R10196 gnd.n4998 gnd.n4997 10.6151
R10197 gnd.n5003 gnd.n4998 10.6151
R10198 gnd.n5003 gnd.n5002 10.6151
R10199 gnd.n5002 gnd.n5001 10.6151
R10200 gnd.n5001 gnd.n4999 10.6151
R10201 gnd.n4999 gnd.n1790 10.6151
R10202 gnd.n5043 gnd.n1790 10.6151
R10203 gnd.n5044 gnd.n5043 10.6151
R10204 gnd.n5045 gnd.n5044 10.6151
R10205 gnd.n5045 gnd.n1781 10.6151
R10206 gnd.n5056 gnd.n1781 10.6151
R10207 gnd.n5057 gnd.n5056 10.6151
R10208 gnd.n5064 gnd.n5057 10.6151
R10209 gnd.n5064 gnd.n5063 10.6151
R10210 gnd.n5063 gnd.n5062 10.6151
R10211 gnd.n5062 gnd.n5061 10.6151
R10212 gnd.n5061 gnd.n5058 10.6151
R10213 gnd.n5058 gnd.n1752 10.6151
R10214 gnd.n5091 gnd.n1752 10.6151
R10215 gnd.n5092 gnd.n5091 10.6151
R10216 gnd.n5095 gnd.n5092 10.6151
R10217 gnd.n5095 gnd.n5094 10.6151
R10218 gnd.n5094 gnd.n5093 10.6151
R10219 gnd.n5093 gnd.n1734 10.6151
R10220 gnd.n5119 gnd.n1734 10.6151
R10221 gnd.n5120 gnd.n5119 10.6151
R10222 gnd.n5125 gnd.n5120 10.6151
R10223 gnd.n5125 gnd.n5124 10.6151
R10224 gnd.n5124 gnd.n5123 10.6151
R10225 gnd.n5123 gnd.n5121 10.6151
R10226 gnd.n5121 gnd.n1708 10.6151
R10227 gnd.n5161 gnd.n1708 10.6151
R10228 gnd.n5162 gnd.n5161 10.6151
R10229 gnd.n5163 gnd.n5162 10.6151
R10230 gnd.n5163 gnd.n1697 10.6151
R10231 gnd.n5176 gnd.n1697 10.6151
R10232 gnd.n5177 gnd.n5176 10.6151
R10233 gnd.n5180 gnd.n5177 10.6151
R10234 gnd.n5180 gnd.n5179 10.6151
R10235 gnd.n5179 gnd.n5178 10.6151
R10236 gnd.n5178 gnd.n1673 10.6151
R10237 gnd.n5201 gnd.n1673 10.6151
R10238 gnd.n5202 gnd.n5201 10.6151
R10239 gnd.n5209 gnd.n5202 10.6151
R10240 gnd.n5209 gnd.n5208 10.6151
R10241 gnd.n5208 gnd.n5207 10.6151
R10242 gnd.n5207 gnd.n5206 10.6151
R10243 gnd.n5206 gnd.n5204 10.6151
R10244 gnd.n5204 gnd.n5203 10.6151
R10245 gnd.n5203 gnd.n1647 10.6151
R10246 gnd.n5235 gnd.n1647 10.6151
R10247 gnd.n5236 gnd.n5235 10.6151
R10248 gnd.n5237 gnd.n5236 10.6151
R10249 gnd.n5241 gnd.n5237 10.6151
R10250 gnd.n5242 gnd.n5241 10.6151
R10251 gnd.n5243 gnd.n5242 10.6151
R10252 gnd.n5243 gnd.n1616 10.6151
R10253 gnd.n5276 gnd.n1616 10.6151
R10254 gnd.n5277 gnd.n5276 10.6151
R10255 gnd.n5278 gnd.n5277 10.6151
R10256 gnd.n5278 gnd.n1614 10.6151
R10257 gnd.n1910 gnd.n1048 10.6151
R10258 gnd.n1913 gnd.n1910 10.6151
R10259 gnd.n1918 gnd.n1915 10.6151
R10260 gnd.n1919 gnd.n1918 10.6151
R10261 gnd.n1922 gnd.n1919 10.6151
R10262 gnd.n1923 gnd.n1922 10.6151
R10263 gnd.n1926 gnd.n1923 10.6151
R10264 gnd.n1927 gnd.n1926 10.6151
R10265 gnd.n1930 gnd.n1927 10.6151
R10266 gnd.n1931 gnd.n1930 10.6151
R10267 gnd.n1934 gnd.n1931 10.6151
R10268 gnd.n1935 gnd.n1934 10.6151
R10269 gnd.n1938 gnd.n1935 10.6151
R10270 gnd.n1939 gnd.n1938 10.6151
R10271 gnd.n1942 gnd.n1939 10.6151
R10272 gnd.n1943 gnd.n1942 10.6151
R10273 gnd.n1946 gnd.n1943 10.6151
R10274 gnd.n1947 gnd.n1946 10.6151
R10275 gnd.n1950 gnd.n1947 10.6151
R10276 gnd.n1951 gnd.n1950 10.6151
R10277 gnd.n1954 gnd.n1951 10.6151
R10278 gnd.n1955 gnd.n1954 10.6151
R10279 gnd.n1958 gnd.n1955 10.6151
R10280 gnd.n1959 gnd.n1958 10.6151
R10281 gnd.n1962 gnd.n1959 10.6151
R10282 gnd.n1963 gnd.n1962 10.6151
R10283 gnd.n1966 gnd.n1963 10.6151
R10284 gnd.n1967 gnd.n1966 10.6151
R10285 gnd.n1970 gnd.n1967 10.6151
R10286 gnd.n1971 gnd.n1970 10.6151
R10287 gnd.n5966 gnd.n5965 10.6151
R10288 gnd.n5965 gnd.n5964 10.6151
R10289 gnd.n5964 gnd.n5963 10.6151
R10290 gnd.n5963 gnd.n5961 10.6151
R10291 gnd.n5961 gnd.n5958 10.6151
R10292 gnd.n5958 gnd.n5957 10.6151
R10293 gnd.n5957 gnd.n5954 10.6151
R10294 gnd.n5954 gnd.n5953 10.6151
R10295 gnd.n5953 gnd.n5950 10.6151
R10296 gnd.n5950 gnd.n5949 10.6151
R10297 gnd.n5949 gnd.n5946 10.6151
R10298 gnd.n5946 gnd.n5945 10.6151
R10299 gnd.n5945 gnd.n5942 10.6151
R10300 gnd.n5942 gnd.n5941 10.6151
R10301 gnd.n5941 gnd.n5938 10.6151
R10302 gnd.n5938 gnd.n5937 10.6151
R10303 gnd.n5937 gnd.n5934 10.6151
R10304 gnd.n5934 gnd.n5933 10.6151
R10305 gnd.n5933 gnd.n5930 10.6151
R10306 gnd.n5930 gnd.n5929 10.6151
R10307 gnd.n5929 gnd.n5926 10.6151
R10308 gnd.n5926 gnd.n5925 10.6151
R10309 gnd.n5925 gnd.n5922 10.6151
R10310 gnd.n5922 gnd.n5921 10.6151
R10311 gnd.n5921 gnd.n5918 10.6151
R10312 gnd.n5918 gnd.n5917 10.6151
R10313 gnd.n5917 gnd.n5914 10.6151
R10314 gnd.n5914 gnd.n5913 10.6151
R10315 gnd.n5910 gnd.n5909 10.6151
R10316 gnd.n5909 gnd.n1049 10.6151
R10317 gnd.n5394 gnd.n1562 10.6151
R10318 gnd.n5394 gnd.n5393 10.6151
R10319 gnd.n5393 gnd.n5392 10.6151
R10320 gnd.n5392 gnd.n1564 10.6151
R10321 gnd.n5387 gnd.n1564 10.6151
R10322 gnd.n5387 gnd.n5386 10.6151
R10323 gnd.n5386 gnd.n5385 10.6151
R10324 gnd.n5385 gnd.n1567 10.6151
R10325 gnd.n5380 gnd.n1567 10.6151
R10326 gnd.n5380 gnd.n5379 10.6151
R10327 gnd.n5379 gnd.n5378 10.6151
R10328 gnd.n5378 gnd.n1570 10.6151
R10329 gnd.n5373 gnd.n1570 10.6151
R10330 gnd.n5373 gnd.n5372 10.6151
R10331 gnd.n5372 gnd.n5371 10.6151
R10332 gnd.n5371 gnd.n1573 10.6151
R10333 gnd.n5366 gnd.n1573 10.6151
R10334 gnd.n5366 gnd.n5365 10.6151
R10335 gnd.n5365 gnd.n5364 10.6151
R10336 gnd.n5364 gnd.n1576 10.6151
R10337 gnd.n5359 gnd.n1576 10.6151
R10338 gnd.n5359 gnd.n5358 10.6151
R10339 gnd.n5358 gnd.n5357 10.6151
R10340 gnd.n5357 gnd.n1579 10.6151
R10341 gnd.n5352 gnd.n1579 10.6151
R10342 gnd.n5352 gnd.n5351 10.6151
R10343 gnd.n5351 gnd.n5350 10.6151
R10344 gnd.n5350 gnd.n1582 10.6151
R10345 gnd.n5345 gnd.n5344 10.6151
R10346 gnd.n5344 gnd.n5343 10.6151
R10347 gnd.n5902 gnd.n5901 10.6151
R10348 gnd.n5901 gnd.n1108 10.6151
R10349 gnd.n4845 gnd.n1108 10.6151
R10350 gnd.n4846 gnd.n4845 10.6151
R10351 gnd.n4847 gnd.n4846 10.6151
R10352 gnd.n4847 gnd.n1902 10.6151
R10353 gnd.n4858 gnd.n1902 10.6151
R10354 gnd.n4859 gnd.n4858 10.6151
R10355 gnd.n4860 gnd.n4859 10.6151
R10356 gnd.n4860 gnd.n1892 10.6151
R10357 gnd.n4886 gnd.n1892 10.6151
R10358 gnd.n4887 gnd.n4886 10.6151
R10359 gnd.n4888 gnd.n4887 10.6151
R10360 gnd.n4888 gnd.n1877 10.6151
R10361 gnd.n4913 gnd.n1877 10.6151
R10362 gnd.n4914 gnd.n4913 10.6151
R10363 gnd.n4915 gnd.n4914 10.6151
R10364 gnd.n4915 gnd.n1866 10.6151
R10365 gnd.n4926 gnd.n1866 10.6151
R10366 gnd.n4927 gnd.n4926 10.6151
R10367 gnd.n4928 gnd.n4927 10.6151
R10368 gnd.n4928 gnd.n1854 10.6151
R10369 gnd.n4944 gnd.n1854 10.6151
R10370 gnd.n4945 gnd.n4944 10.6151
R10371 gnd.n4946 gnd.n4945 10.6151
R10372 gnd.n4946 gnd.n1840 10.6151
R10373 gnd.n4961 gnd.n1840 10.6151
R10374 gnd.n4962 gnd.n4961 10.6151
R10375 gnd.n4964 gnd.n4962 10.6151
R10376 gnd.n4964 gnd.n4963 10.6151
R10377 gnd.n4963 gnd.n1821 10.6151
R10378 gnd.n4990 gnd.n1821 10.6151
R10379 gnd.n4991 gnd.n4990 10.6151
R10380 gnd.n4992 gnd.n4991 10.6151
R10381 gnd.n4992 gnd.n1812 10.6151
R10382 gnd.n5010 gnd.n1812 10.6151
R10383 gnd.n5011 gnd.n5010 10.6151
R10384 gnd.n5012 gnd.n5011 10.6151
R10385 gnd.n5012 gnd.n1797 10.6151
R10386 gnd.n5037 gnd.n1797 10.6151
R10387 gnd.n5038 gnd.n5037 10.6151
R10388 gnd.n5039 gnd.n5038 10.6151
R10389 gnd.n5039 gnd.n1786 10.6151
R10390 gnd.n5050 gnd.n1786 10.6151
R10391 gnd.n5051 gnd.n5050 10.6151
R10392 gnd.n5052 gnd.n5051 10.6151
R10393 gnd.n5052 gnd.n1774 10.6151
R10394 gnd.n5068 gnd.n1774 10.6151
R10395 gnd.n5069 gnd.n5068 10.6151
R10396 gnd.n5070 gnd.n5069 10.6151
R10397 gnd.n5070 gnd.n1759 10.6151
R10398 gnd.n5084 gnd.n1759 10.6151
R10399 gnd.n5085 gnd.n5084 10.6151
R10400 gnd.n5087 gnd.n5085 10.6151
R10401 gnd.n5087 gnd.n5086 10.6151
R10402 gnd.n5086 gnd.n1739 10.6151
R10403 gnd.n5112 gnd.n1739 10.6151
R10404 gnd.n5113 gnd.n5112 10.6151
R10405 gnd.n5114 gnd.n5113 10.6151
R10406 gnd.n5114 gnd.n1729 10.6151
R10407 gnd.n5131 gnd.n1729 10.6151
R10408 gnd.n5132 gnd.n5131 10.6151
R10409 gnd.n5133 gnd.n5132 10.6151
R10410 gnd.n5133 gnd.n1714 10.6151
R10411 gnd.n5155 gnd.n1714 10.6151
R10412 gnd.n5156 gnd.n5155 10.6151
R10413 gnd.n5157 gnd.n5156 10.6151
R10414 gnd.n5157 gnd.n1704 10.6151
R10415 gnd.n5168 gnd.n1704 10.6151
R10416 gnd.n5169 gnd.n5168 10.6151
R10417 gnd.n5172 gnd.n5169 10.6151
R10418 gnd.n5172 gnd.n5171 10.6151
R10419 gnd.n5171 gnd.n5170 10.6151
R10420 gnd.n5170 gnd.n1679 10.6151
R10421 gnd.n5195 gnd.n1679 10.6151
R10422 gnd.n5196 gnd.n5195 10.6151
R10423 gnd.n5197 gnd.n5196 10.6151
R10424 gnd.n5197 gnd.n1668 10.6151
R10425 gnd.n5213 gnd.n1668 10.6151
R10426 gnd.n5214 gnd.n5213 10.6151
R10427 gnd.n5215 gnd.n5214 10.6151
R10428 gnd.n5215 gnd.n1651 10.6151
R10429 gnd.n5228 gnd.n1651 10.6151
R10430 gnd.n5229 gnd.n5228 10.6151
R10431 gnd.n5230 gnd.n5229 10.6151
R10432 gnd.n5230 gnd.n1640 10.6151
R10433 gnd.n5251 gnd.n1640 10.6151
R10434 gnd.n5251 gnd.n5250 10.6151
R10435 gnd.n5250 gnd.n5249 10.6151
R10436 gnd.n5249 gnd.n1641 10.6151
R10437 gnd.n1644 gnd.n1641 10.6151
R10438 gnd.n1644 gnd.n1643 10.6151
R10439 gnd.n1643 gnd.n1541 10.6151
R10440 gnd.n5401 gnd.n1541 10.6151
R10441 gnd.n5401 gnd.n5400 10.6151
R10442 gnd.n5400 gnd.n5399 10.6151
R10443 gnd.n2942 gnd.t29 10.5161
R10444 gnd.n2371 gnd.t37 10.5161
R10445 gnd.n3308 gnd.t8 10.5161
R10446 gnd.n3584 gnd.n3568 10.4732
R10447 gnd.n3552 gnd.n3536 10.4732
R10448 gnd.n3520 gnd.n3504 10.4732
R10449 gnd.n3489 gnd.n3473 10.4732
R10450 gnd.n3457 gnd.n3441 10.4732
R10451 gnd.n3425 gnd.n3409 10.4732
R10452 gnd.n3393 gnd.n3377 10.4732
R10453 gnd.n3362 gnd.n3346 10.4732
R10454 gnd.n1864 gnd.n1863 10.1975
R10455 gnd.n1784 gnd.n1776 10.1975
R10456 gnd.n5073 gnd.n1769 10.1975
R10457 gnd.n1695 gnd.n1681 10.1975
R10458 gnd.t185 gnd.n2388 9.87883
R10459 gnd.n3588 gnd.n3587 9.69747
R10460 gnd.n3556 gnd.n3555 9.69747
R10461 gnd.n3524 gnd.n3523 9.69747
R10462 gnd.n3493 gnd.n3492 9.69747
R10463 gnd.n3461 gnd.n3460 9.69747
R10464 gnd.n3429 gnd.n3428 9.69747
R10465 gnd.n3397 gnd.n3396 9.69747
R10466 gnd.n3366 gnd.n3365 9.69747
R10467 gnd.n4986 gnd.t356 9.56018
R10468 gnd.n5136 gnd.t178 9.56018
R10469 gnd.n1537 gnd.t81 9.56018
R10470 gnd.n3594 gnd.n3593 9.45567
R10471 gnd.n3562 gnd.n3561 9.45567
R10472 gnd.n3530 gnd.n3529 9.45567
R10473 gnd.n3499 gnd.n3498 9.45567
R10474 gnd.n3467 gnd.n3466 9.45567
R10475 gnd.n3435 gnd.n3434 9.45567
R10476 gnd.n3403 gnd.n3402 9.45567
R10477 gnd.n3372 gnd.n3371 9.45567
R10478 gnd.n7108 gnd.n285 9.30959
R10479 gnd.n5640 gnd.n5639 9.30959
R10480 gnd.n3960 gnd.n3959 9.30959
R10481 gnd.n4527 gnd.n4524 9.30959
R10482 gnd.n5600 gnd.n5599 9.3005
R10483 gnd.n5603 gnd.n1395 9.3005
R10484 gnd.n5604 gnd.n1394 9.3005
R10485 gnd.n5607 gnd.n1393 9.3005
R10486 gnd.n5608 gnd.n1392 9.3005
R10487 gnd.n5611 gnd.n1391 9.3005
R10488 gnd.n5612 gnd.n1390 9.3005
R10489 gnd.n5615 gnd.n1389 9.3005
R10490 gnd.n5616 gnd.n1388 9.3005
R10491 gnd.n5619 gnd.n1387 9.3005
R10492 gnd.n5620 gnd.n1386 9.3005
R10493 gnd.n5623 gnd.n1385 9.3005
R10494 gnd.n5624 gnd.n1384 9.3005
R10495 gnd.n5627 gnd.n1383 9.3005
R10496 gnd.n5628 gnd.n1382 9.3005
R10497 gnd.n5631 gnd.n1381 9.3005
R10498 gnd.n5632 gnd.n1380 9.3005
R10499 gnd.n5635 gnd.n1379 9.3005
R10500 gnd.n5636 gnd.n1378 9.3005
R10501 gnd.n5639 gnd.n1377 9.3005
R10502 gnd.n5643 gnd.n1373 9.3005
R10503 gnd.n5644 gnd.n1372 9.3005
R10504 gnd.n5647 gnd.n1371 9.3005
R10505 gnd.n5648 gnd.n1370 9.3005
R10506 gnd.n5651 gnd.n1369 9.3005
R10507 gnd.n5652 gnd.n1368 9.3005
R10508 gnd.n5655 gnd.n1367 9.3005
R10509 gnd.n5656 gnd.n1366 9.3005
R10510 gnd.n5659 gnd.n1365 9.3005
R10511 gnd.n5661 gnd.n1361 9.3005
R10512 gnd.n5664 gnd.n1360 9.3005
R10513 gnd.n5665 gnd.n1359 9.3005
R10514 gnd.n5668 gnd.n1358 9.3005
R10515 gnd.n5669 gnd.n1357 9.3005
R10516 gnd.n5672 gnd.n1356 9.3005
R10517 gnd.n5673 gnd.n1355 9.3005
R10518 gnd.n5676 gnd.n1354 9.3005
R10519 gnd.n5678 gnd.n1351 9.3005
R10520 gnd.n5681 gnd.n1350 9.3005
R10521 gnd.n5682 gnd.n1349 9.3005
R10522 gnd.n5685 gnd.n1348 9.3005
R10523 gnd.n5686 gnd.n1347 9.3005
R10524 gnd.n5689 gnd.n1346 9.3005
R10525 gnd.n5690 gnd.n1345 9.3005
R10526 gnd.n5693 gnd.n1344 9.3005
R10527 gnd.n5694 gnd.n1343 9.3005
R10528 gnd.n5697 gnd.n1342 9.3005
R10529 gnd.n5698 gnd.n1341 9.3005
R10530 gnd.n5701 gnd.n1340 9.3005
R10531 gnd.n5702 gnd.n1339 9.3005
R10532 gnd.n5705 gnd.n1338 9.3005
R10533 gnd.n5707 gnd.n1337 9.3005
R10534 gnd.n5708 gnd.n1336 9.3005
R10535 gnd.n5709 gnd.n1335 9.3005
R10536 gnd.n5710 gnd.n1334 9.3005
R10537 gnd.n5640 gnd.n1374 9.3005
R10538 gnd.n5598 gnd.n5595 9.3005
R10539 gnd.n1416 gnd.n1413 9.3005
R10540 gnd.n5584 gnd.n1417 9.3005
R10541 gnd.n5583 gnd.n1418 9.3005
R10542 gnd.n5582 gnd.n1419 9.3005
R10543 gnd.n1437 gnd.n1420 9.3005
R10544 gnd.n5572 gnd.n1438 9.3005
R10545 gnd.n5571 gnd.n1439 9.3005
R10546 gnd.n5570 gnd.n1440 9.3005
R10547 gnd.n5556 gnd.n1441 9.3005
R10548 gnd.n5560 gnd.n5557 9.3005
R10549 gnd.n5559 gnd.n5558 9.3005
R10550 gnd.n377 gnd.n376 9.3005
R10551 gnd.n6810 gnd.n6809 9.3005
R10552 gnd.n6811 gnd.n375 9.3005
R10553 gnd.n6815 gnd.n6812 9.3005
R10554 gnd.n6814 gnd.n6813 9.3005
R10555 gnd.n349 gnd.n348 9.3005
R10556 gnd.n6844 gnd.n6843 9.3005
R10557 gnd.n6845 gnd.n347 9.3005
R10558 gnd.n6849 gnd.n6846 9.3005
R10559 gnd.n6848 gnd.n6847 9.3005
R10560 gnd.n1415 gnd.n1414 9.3005
R10561 gnd.n327 gnd.n326 9.3005
R10562 gnd.n6877 gnd.n6876 9.3005
R10563 gnd.n6878 gnd.n325 9.3005
R10564 gnd.n6883 gnd.n6879 9.3005
R10565 gnd.n6882 gnd.n6881 9.3005
R10566 gnd.n6880 gnd.n90 9.3005
R10567 gnd.n7261 gnd.n91 9.3005
R10568 gnd.n7260 gnd.n92 9.3005
R10569 gnd.n7259 gnd.n93 9.3005
R10570 gnd.n111 gnd.n94 9.3005
R10571 gnd.n7249 gnd.n112 9.3005
R10572 gnd.n7248 gnd.n113 9.3005
R10573 gnd.n7247 gnd.n114 9.3005
R10574 gnd.n130 gnd.n115 9.3005
R10575 gnd.n7237 gnd.n131 9.3005
R10576 gnd.n7236 gnd.n132 9.3005
R10577 gnd.n7235 gnd.n133 9.3005
R10578 gnd.n149 gnd.n134 9.3005
R10579 gnd.n7225 gnd.n150 9.3005
R10580 gnd.n7224 gnd.n151 9.3005
R10581 gnd.n7223 gnd.n152 9.3005
R10582 gnd.n168 gnd.n153 9.3005
R10583 gnd.n7213 gnd.n169 9.3005
R10584 gnd.n7212 gnd.n170 9.3005
R10585 gnd.n7211 gnd.n171 9.3005
R10586 gnd.n187 gnd.n172 9.3005
R10587 gnd.n7201 gnd.n188 9.3005
R10588 gnd.n7200 gnd.n189 9.3005
R10589 gnd.n7199 gnd.n190 9.3005
R10590 gnd.n206 gnd.n191 9.3005
R10591 gnd.n7189 gnd.n207 9.3005
R10592 gnd.n7188 gnd.n7187 9.3005
R10593 gnd.n7267 gnd.n7266 9.3005
R10594 gnd.n7265 gnd.n80 9.3005
R10595 gnd.n6930 gnd.n83 9.3005
R10596 gnd.n6931 gnd.n6929 9.3005
R10597 gnd.n6934 gnd.n6932 9.3005
R10598 gnd.n6935 gnd.n6928 9.3005
R10599 gnd.n6938 gnd.n6937 9.3005
R10600 gnd.n6939 gnd.n6927 9.3005
R10601 gnd.n6942 gnd.n6940 9.3005
R10602 gnd.n6943 gnd.n6926 9.3005
R10603 gnd.n6946 gnd.n6945 9.3005
R10604 gnd.n6947 gnd.n6925 9.3005
R10605 gnd.n6950 gnd.n6948 9.3005
R10606 gnd.n6951 gnd.n6924 9.3005
R10607 gnd.n6954 gnd.n6953 9.3005
R10608 gnd.n6955 gnd.n6923 9.3005
R10609 gnd.n7039 gnd.n6956 9.3005
R10610 gnd.n7038 gnd.n6957 9.3005
R10611 gnd.n7037 gnd.n6958 9.3005
R10612 gnd.n7035 gnd.n6959 9.3005
R10613 gnd.n7034 gnd.n6960 9.3005
R10614 gnd.n7032 gnd.n6961 9.3005
R10615 gnd.n7031 gnd.n6962 9.3005
R10616 gnd.n7029 gnd.n6963 9.3005
R10617 gnd.n7028 gnd.n6964 9.3005
R10618 gnd.n7026 gnd.n6965 9.3005
R10619 gnd.n7025 gnd.n6966 9.3005
R10620 gnd.n6980 gnd.n6979 9.3005
R10621 gnd.n6982 gnd.n6981 9.3005
R10622 gnd.n6985 gnd.n6976 9.3005
R10623 gnd.n6989 gnd.n6988 9.3005
R10624 gnd.n6990 gnd.n6975 9.3005
R10625 gnd.n6992 gnd.n6991 9.3005
R10626 gnd.n6995 gnd.n6974 9.3005
R10627 gnd.n6999 gnd.n6998 9.3005
R10628 gnd.n7000 gnd.n6973 9.3005
R10629 gnd.n7002 gnd.n7001 9.3005
R10630 gnd.n7005 gnd.n6972 9.3005
R10631 gnd.n7009 gnd.n7008 9.3005
R10632 gnd.n7010 gnd.n6971 9.3005
R10633 gnd.n7012 gnd.n7011 9.3005
R10634 gnd.n7015 gnd.n6970 9.3005
R10635 gnd.n7019 gnd.n7018 9.3005
R10636 gnd.n7020 gnd.n6969 9.3005
R10637 gnd.n7022 gnd.n7021 9.3005
R10638 gnd.n6977 gnd.n308 9.3005
R10639 gnd.n209 gnd.n208 9.3005
R10640 gnd.n7180 gnd.n250 9.3005
R10641 gnd.n7179 gnd.n251 9.3005
R10642 gnd.n7178 gnd.n252 9.3005
R10643 gnd.n7175 gnd.n253 9.3005
R10644 gnd.n7174 gnd.n254 9.3005
R10645 gnd.n7171 gnd.n255 9.3005
R10646 gnd.n7170 gnd.n256 9.3005
R10647 gnd.n7167 gnd.n257 9.3005
R10648 gnd.n7166 gnd.n258 9.3005
R10649 gnd.n7163 gnd.n259 9.3005
R10650 gnd.n7162 gnd.n260 9.3005
R10651 gnd.n7159 gnd.n261 9.3005
R10652 gnd.n7158 gnd.n262 9.3005
R10653 gnd.n7155 gnd.n263 9.3005
R10654 gnd.n7154 gnd.n264 9.3005
R10655 gnd.n7151 gnd.n265 9.3005
R10656 gnd.n7147 gnd.n266 9.3005
R10657 gnd.n7144 gnd.n267 9.3005
R10658 gnd.n7143 gnd.n268 9.3005
R10659 gnd.n7140 gnd.n269 9.3005
R10660 gnd.n7139 gnd.n270 9.3005
R10661 gnd.n7136 gnd.n271 9.3005
R10662 gnd.n7135 gnd.n272 9.3005
R10663 gnd.n7132 gnd.n273 9.3005
R10664 gnd.n7131 gnd.n274 9.3005
R10665 gnd.n7128 gnd.n275 9.3005
R10666 gnd.n7127 gnd.n276 9.3005
R10667 gnd.n7124 gnd.n277 9.3005
R10668 gnd.n7123 gnd.n278 9.3005
R10669 gnd.n7120 gnd.n279 9.3005
R10670 gnd.n7119 gnd.n280 9.3005
R10671 gnd.n7116 gnd.n281 9.3005
R10672 gnd.n7115 gnd.n282 9.3005
R10673 gnd.n7112 gnd.n283 9.3005
R10674 gnd.n7111 gnd.n284 9.3005
R10675 gnd.n7108 gnd.n7107 9.3005
R10676 gnd.n7106 gnd.n285 9.3005
R10677 gnd.n7105 gnd.n7104 9.3005
R10678 gnd.n7101 gnd.n288 9.3005
R10679 gnd.n7098 gnd.n289 9.3005
R10680 gnd.n7097 gnd.n290 9.3005
R10681 gnd.n7094 gnd.n291 9.3005
R10682 gnd.n7093 gnd.n292 9.3005
R10683 gnd.n7090 gnd.n293 9.3005
R10684 gnd.n7089 gnd.n294 9.3005
R10685 gnd.n7086 gnd.n295 9.3005
R10686 gnd.n7085 gnd.n296 9.3005
R10687 gnd.n7082 gnd.n297 9.3005
R10688 gnd.n7081 gnd.n298 9.3005
R10689 gnd.n7078 gnd.n299 9.3005
R10690 gnd.n7077 gnd.n300 9.3005
R10691 gnd.n7074 gnd.n301 9.3005
R10692 gnd.n7073 gnd.n302 9.3005
R10693 gnd.n7070 gnd.n303 9.3005
R10694 gnd.n7069 gnd.n304 9.3005
R10695 gnd.n7066 gnd.n7065 9.3005
R10696 gnd.n7064 gnd.n305 9.3005
R10697 gnd.n7186 gnd.n7185 9.3005
R10698 gnd.n5477 gnd.n1404 9.3005
R10699 gnd.n5478 gnd.n1405 9.3005
R10700 gnd.n5482 gnd.n5479 9.3005
R10701 gnd.n5483 gnd.n1427 9.3005
R10702 gnd.n5486 gnd.n1428 9.3005
R10703 gnd.n5487 gnd.n1429 9.3005
R10704 gnd.n5491 gnd.n5488 9.3005
R10705 gnd.n5492 gnd.n1448 9.3005
R10706 gnd.n5495 gnd.n1449 9.3005
R10707 gnd.n5496 gnd.n1450 9.3005
R10708 gnd.n5498 gnd.n5497 9.3005
R10709 gnd.n5500 gnd.n5499 9.3005
R10710 gnd.n388 gnd.n386 9.3005
R10711 gnd.n6796 gnd.n387 9.3005
R10712 gnd.n6798 gnd.n6797 9.3005
R10713 gnd.n6799 gnd.n360 9.3005
R10714 gnd.n6828 gnd.n361 9.3005
R10715 gnd.n6829 gnd.n358 9.3005
R10716 gnd.n6831 gnd.n359 9.3005
R10717 gnd.n6833 gnd.n6832 9.3005
R10718 gnd.n6834 gnd.n334 9.3005
R10719 gnd.n6867 gnd.n333 9.3005
R10720 gnd.n6871 gnd.n6870 9.3005
R10721 gnd.n6869 gnd.n316 9.3005
R10722 gnd.n6888 gnd.n315 9.3005
R10723 gnd.n6890 gnd.n6889 9.3005
R10724 gnd.n6891 gnd.n310 9.3005
R10725 gnd.n6897 gnd.n309 9.3005
R10726 gnd.n6900 gnd.n6898 9.3005
R10727 gnd.n6901 gnd.n101 9.3005
R10728 gnd.n6903 gnd.n102 9.3005
R10729 gnd.n6904 gnd.n103 9.3005
R10730 gnd.n6907 gnd.n6905 9.3005
R10731 gnd.n6908 gnd.n121 9.3005
R10732 gnd.n6910 gnd.n122 9.3005
R10733 gnd.n6911 gnd.n123 9.3005
R10734 gnd.n6914 gnd.n6912 9.3005
R10735 gnd.n6915 gnd.n139 9.3005
R10736 gnd.n6917 gnd.n140 9.3005
R10737 gnd.n6918 gnd.n141 9.3005
R10738 gnd.n6921 gnd.n6919 9.3005
R10739 gnd.n6922 gnd.n159 9.3005
R10740 gnd.n7043 gnd.n160 9.3005
R10741 gnd.n7044 gnd.n161 9.3005
R10742 gnd.n7047 gnd.n7045 9.3005
R10743 gnd.n7048 gnd.n177 9.3005
R10744 gnd.n7050 gnd.n178 9.3005
R10745 gnd.n7051 gnd.n179 9.3005
R10746 gnd.n7054 gnd.n7052 9.3005
R10747 gnd.n7055 gnd.n197 9.3005
R10748 gnd.n7057 gnd.n198 9.3005
R10749 gnd.n7058 gnd.n199 9.3005
R10750 gnd.n7062 gnd.n7061 9.3005
R10751 gnd.n1403 gnd.n1397 9.3005
R10752 gnd.n5589 gnd.n1404 9.3005
R10753 gnd.n5588 gnd.n1405 9.3005
R10754 gnd.n5479 gnd.n1406 9.3005
R10755 gnd.n5578 gnd.n1427 9.3005
R10756 gnd.n5577 gnd.n1428 9.3005
R10757 gnd.n5576 gnd.n1429 9.3005
R10758 gnd.n5488 gnd.n1430 9.3005
R10759 gnd.n5566 gnd.n1448 9.3005
R10760 gnd.n5565 gnd.n1449 9.3005
R10761 gnd.n5564 gnd.n1450 9.3005
R10762 gnd.n5498 gnd.n1451 9.3005
R10763 gnd.n5499 gnd.n385 9.3005
R10764 gnd.n6805 gnd.n386 9.3005
R10765 gnd.n6804 gnd.n387 9.3005
R10766 gnd.n6803 gnd.n6798 9.3005
R10767 gnd.n6802 gnd.n6799 9.3005
R10768 gnd.n361 gnd.n357 9.3005
R10769 gnd.n6839 gnd.n358 9.3005
R10770 gnd.n6838 gnd.n359 9.3005
R10771 gnd.n6837 gnd.n6833 9.3005
R10772 gnd.n6836 gnd.n6834 9.3005
R10773 gnd.n333 gnd.n332 9.3005
R10774 gnd.n6872 gnd.n6871 9.3005
R10775 gnd.n317 gnd.n316 9.3005
R10776 gnd.n6888 gnd.n6887 9.3005
R10777 gnd.n6889 gnd.n311 9.3005
R10778 gnd.n6895 gnd.n310 9.3005
R10779 gnd.n6897 gnd.n6896 9.3005
R10780 gnd.n6898 gnd.n100 9.3005
R10781 gnd.n7255 gnd.n101 9.3005
R10782 gnd.n7254 gnd.n102 9.3005
R10783 gnd.n7253 gnd.n103 9.3005
R10784 gnd.n6905 gnd.n104 9.3005
R10785 gnd.n7243 gnd.n121 9.3005
R10786 gnd.n7242 gnd.n122 9.3005
R10787 gnd.n7241 gnd.n123 9.3005
R10788 gnd.n6912 gnd.n124 9.3005
R10789 gnd.n7231 gnd.n139 9.3005
R10790 gnd.n7230 gnd.n140 9.3005
R10791 gnd.n7229 gnd.n141 9.3005
R10792 gnd.n6919 gnd.n142 9.3005
R10793 gnd.n7219 gnd.n159 9.3005
R10794 gnd.n7218 gnd.n160 9.3005
R10795 gnd.n7217 gnd.n161 9.3005
R10796 gnd.n7045 gnd.n162 9.3005
R10797 gnd.n7207 gnd.n177 9.3005
R10798 gnd.n7206 gnd.n178 9.3005
R10799 gnd.n7205 gnd.n179 9.3005
R10800 gnd.n7052 gnd.n180 9.3005
R10801 gnd.n7195 gnd.n197 9.3005
R10802 gnd.n7194 gnd.n198 9.3005
R10803 gnd.n7193 gnd.n199 9.3005
R10804 gnd.n7062 gnd.n200 9.3005
R10805 gnd.n5590 gnd.n1403 9.3005
R10806 gnd.n3593 gnd.n3592 9.3005
R10807 gnd.n3566 gnd.n3565 9.3005
R10808 gnd.n3587 gnd.n3586 9.3005
R10809 gnd.n3585 gnd.n3584 9.3005
R10810 gnd.n3570 gnd.n3569 9.3005
R10811 gnd.n3579 gnd.n3578 9.3005
R10812 gnd.n3577 gnd.n3576 9.3005
R10813 gnd.n3561 gnd.n3560 9.3005
R10814 gnd.n3534 gnd.n3533 9.3005
R10815 gnd.n3555 gnd.n3554 9.3005
R10816 gnd.n3553 gnd.n3552 9.3005
R10817 gnd.n3538 gnd.n3537 9.3005
R10818 gnd.n3547 gnd.n3546 9.3005
R10819 gnd.n3545 gnd.n3544 9.3005
R10820 gnd.n3529 gnd.n3528 9.3005
R10821 gnd.n3502 gnd.n3501 9.3005
R10822 gnd.n3523 gnd.n3522 9.3005
R10823 gnd.n3521 gnd.n3520 9.3005
R10824 gnd.n3506 gnd.n3505 9.3005
R10825 gnd.n3515 gnd.n3514 9.3005
R10826 gnd.n3513 gnd.n3512 9.3005
R10827 gnd.n3498 gnd.n3497 9.3005
R10828 gnd.n3471 gnd.n3470 9.3005
R10829 gnd.n3492 gnd.n3491 9.3005
R10830 gnd.n3490 gnd.n3489 9.3005
R10831 gnd.n3475 gnd.n3474 9.3005
R10832 gnd.n3484 gnd.n3483 9.3005
R10833 gnd.n3482 gnd.n3481 9.3005
R10834 gnd.n3466 gnd.n3465 9.3005
R10835 gnd.n3439 gnd.n3438 9.3005
R10836 gnd.n3460 gnd.n3459 9.3005
R10837 gnd.n3458 gnd.n3457 9.3005
R10838 gnd.n3443 gnd.n3442 9.3005
R10839 gnd.n3452 gnd.n3451 9.3005
R10840 gnd.n3450 gnd.n3449 9.3005
R10841 gnd.n3434 gnd.n3433 9.3005
R10842 gnd.n3407 gnd.n3406 9.3005
R10843 gnd.n3428 gnd.n3427 9.3005
R10844 gnd.n3426 gnd.n3425 9.3005
R10845 gnd.n3411 gnd.n3410 9.3005
R10846 gnd.n3420 gnd.n3419 9.3005
R10847 gnd.n3418 gnd.n3417 9.3005
R10848 gnd.n3402 gnd.n3401 9.3005
R10849 gnd.n3375 gnd.n3374 9.3005
R10850 gnd.n3396 gnd.n3395 9.3005
R10851 gnd.n3394 gnd.n3393 9.3005
R10852 gnd.n3379 gnd.n3378 9.3005
R10853 gnd.n3388 gnd.n3387 9.3005
R10854 gnd.n3386 gnd.n3385 9.3005
R10855 gnd.n3371 gnd.n3370 9.3005
R10856 gnd.n3344 gnd.n3343 9.3005
R10857 gnd.n3365 gnd.n3364 9.3005
R10858 gnd.n3363 gnd.n3362 9.3005
R10859 gnd.n3348 gnd.n3347 9.3005
R10860 gnd.n3357 gnd.n3356 9.3005
R10861 gnd.n3355 gnd.n3354 9.3005
R10862 gnd.n3719 gnd.n3718 9.3005
R10863 gnd.n3717 gnd.n2270 9.3005
R10864 gnd.n3716 gnd.n3715 9.3005
R10865 gnd.n3712 gnd.n2271 9.3005
R10866 gnd.n3709 gnd.n2272 9.3005
R10867 gnd.n3708 gnd.n2273 9.3005
R10868 gnd.n3705 gnd.n2274 9.3005
R10869 gnd.n3704 gnd.n2275 9.3005
R10870 gnd.n3701 gnd.n2276 9.3005
R10871 gnd.n3700 gnd.n2277 9.3005
R10872 gnd.n3697 gnd.n2278 9.3005
R10873 gnd.n3696 gnd.n2279 9.3005
R10874 gnd.n3693 gnd.n2280 9.3005
R10875 gnd.n3692 gnd.n2281 9.3005
R10876 gnd.n3689 gnd.n3688 9.3005
R10877 gnd.n3687 gnd.n2282 9.3005
R10878 gnd.n3720 gnd.n2269 9.3005
R10879 gnd.n2961 gnd.n2960 9.3005
R10880 gnd.n2665 gnd.n2664 9.3005
R10881 gnd.n2988 gnd.n2987 9.3005
R10882 gnd.n2989 gnd.n2663 9.3005
R10883 gnd.n2993 gnd.n2990 9.3005
R10884 gnd.n2992 gnd.n2991 9.3005
R10885 gnd.n2637 gnd.n2636 9.3005
R10886 gnd.n3018 gnd.n3017 9.3005
R10887 gnd.n3019 gnd.n2635 9.3005
R10888 gnd.n3021 gnd.n3020 9.3005
R10889 gnd.n2615 gnd.n2614 9.3005
R10890 gnd.n3049 gnd.n3048 9.3005
R10891 gnd.n3050 gnd.n2613 9.3005
R10892 gnd.n3058 gnd.n3051 9.3005
R10893 gnd.n3057 gnd.n3052 9.3005
R10894 gnd.n3056 gnd.n3054 9.3005
R10895 gnd.n3053 gnd.n2562 9.3005
R10896 gnd.n3106 gnd.n2563 9.3005
R10897 gnd.n3105 gnd.n2564 9.3005
R10898 gnd.n3104 gnd.n2565 9.3005
R10899 gnd.n2584 gnd.n2566 9.3005
R10900 gnd.n2586 gnd.n2585 9.3005
R10901 gnd.n2468 gnd.n2467 9.3005
R10902 gnd.n3144 gnd.n3143 9.3005
R10903 gnd.n3145 gnd.n2466 9.3005
R10904 gnd.n3149 gnd.n3146 9.3005
R10905 gnd.n3148 gnd.n3147 9.3005
R10906 gnd.n2441 gnd.n2440 9.3005
R10907 gnd.n3184 gnd.n3183 9.3005
R10908 gnd.n3185 gnd.n2439 9.3005
R10909 gnd.n3189 gnd.n3186 9.3005
R10910 gnd.n3188 gnd.n3187 9.3005
R10911 gnd.n2414 gnd.n2413 9.3005
R10912 gnd.n3229 gnd.n3228 9.3005
R10913 gnd.n3230 gnd.n2412 9.3005
R10914 gnd.n3234 gnd.n3231 9.3005
R10915 gnd.n3233 gnd.n3232 9.3005
R10916 gnd.n2386 gnd.n2385 9.3005
R10917 gnd.n3269 gnd.n3268 9.3005
R10918 gnd.n3270 gnd.n2384 9.3005
R10919 gnd.n3274 gnd.n3271 9.3005
R10920 gnd.n3273 gnd.n3272 9.3005
R10921 gnd.n2359 gnd.n2358 9.3005
R10922 gnd.n3318 gnd.n3317 9.3005
R10923 gnd.n3319 gnd.n2357 9.3005
R10924 gnd.n3323 gnd.n3320 9.3005
R10925 gnd.n3322 gnd.n3321 9.3005
R10926 gnd.n2332 gnd.n2331 9.3005
R10927 gnd.n3612 gnd.n3611 9.3005
R10928 gnd.n3613 gnd.n2330 9.3005
R10929 gnd.n3619 gnd.n3614 9.3005
R10930 gnd.n3618 gnd.n3615 9.3005
R10931 gnd.n3617 gnd.n3616 9.3005
R10932 gnd.n2962 gnd.n2959 9.3005
R10933 gnd.n2744 gnd.n2703 9.3005
R10934 gnd.n2739 gnd.n2738 9.3005
R10935 gnd.n2737 gnd.n2704 9.3005
R10936 gnd.n2736 gnd.n2735 9.3005
R10937 gnd.n2732 gnd.n2705 9.3005
R10938 gnd.n2729 gnd.n2728 9.3005
R10939 gnd.n2727 gnd.n2706 9.3005
R10940 gnd.n2726 gnd.n2725 9.3005
R10941 gnd.n2722 gnd.n2707 9.3005
R10942 gnd.n2719 gnd.n2718 9.3005
R10943 gnd.n2717 gnd.n2708 9.3005
R10944 gnd.n2716 gnd.n2715 9.3005
R10945 gnd.n2712 gnd.n2710 9.3005
R10946 gnd.n2709 gnd.n2689 9.3005
R10947 gnd.n2956 gnd.n2688 9.3005
R10948 gnd.n2958 gnd.n2957 9.3005
R10949 gnd.n2746 gnd.n2745 9.3005
R10950 gnd.n2969 gnd.n2675 9.3005
R10951 gnd.n2976 gnd.n2676 9.3005
R10952 gnd.n2978 gnd.n2977 9.3005
R10953 gnd.n2979 gnd.n2656 9.3005
R10954 gnd.n2998 gnd.n2997 9.3005
R10955 gnd.n3000 gnd.n2648 9.3005
R10956 gnd.n3007 gnd.n2650 9.3005
R10957 gnd.n3008 gnd.n2645 9.3005
R10958 gnd.n3010 gnd.n3009 9.3005
R10959 gnd.n2646 gnd.n2631 9.3005
R10960 gnd.n3026 gnd.n2629 9.3005
R10961 gnd.n3030 gnd.n3029 9.3005
R10962 gnd.n3028 gnd.n2605 9.3005
R10963 gnd.n3065 gnd.n2604 9.3005
R10964 gnd.n3068 gnd.n3067 9.3005
R10965 gnd.n2601 gnd.n2600 9.3005
R10966 gnd.n3074 gnd.n2602 9.3005
R10967 gnd.n3076 gnd.n3075 9.3005
R10968 gnd.n3078 gnd.n2599 9.3005
R10969 gnd.n3081 gnd.n3080 9.3005
R10970 gnd.n3084 gnd.n3082 9.3005
R10971 gnd.n3086 gnd.n3085 9.3005
R10972 gnd.n3092 gnd.n3087 9.3005
R10973 gnd.n3091 gnd.n3090 9.3005
R10974 gnd.n2459 gnd.n2458 9.3005
R10975 gnd.n3158 gnd.n3157 9.3005
R10976 gnd.n3159 gnd.n2452 9.3005
R10977 gnd.n3167 gnd.n2451 9.3005
R10978 gnd.n3170 gnd.n3169 9.3005
R10979 gnd.n3172 gnd.n3171 9.3005
R10980 gnd.n3175 gnd.n2434 9.3005
R10981 gnd.n3173 gnd.n2432 9.3005
R10982 gnd.n3195 gnd.n2430 9.3005
R10983 gnd.n3197 gnd.n3196 9.3005
R10984 gnd.n2404 gnd.n2403 9.3005
R10985 gnd.n3243 gnd.n3242 9.3005
R10986 gnd.n3244 gnd.n2397 9.3005
R10987 gnd.n3252 gnd.n2396 9.3005
R10988 gnd.n3255 gnd.n3254 9.3005
R10989 gnd.n3257 gnd.n3256 9.3005
R10990 gnd.n3260 gnd.n2379 9.3005
R10991 gnd.n3258 gnd.n2377 9.3005
R10992 gnd.n3280 gnd.n2375 9.3005
R10993 gnd.n3282 gnd.n3281 9.3005
R10994 gnd.n2350 gnd.n2349 9.3005
R10995 gnd.n3332 gnd.n3331 9.3005
R10996 gnd.n3333 gnd.n2343 9.3005
R10997 gnd.n3341 gnd.n2342 9.3005
R10998 gnd.n3600 gnd.n3599 9.3005
R10999 gnd.n3602 gnd.n3601 9.3005
R11000 gnd.n3603 gnd.n2323 9.3005
R11001 gnd.n3627 gnd.n3626 9.3005
R11002 gnd.n2324 gnd.n2285 9.3005
R11003 gnd.n2967 gnd.n2966 9.3005
R11004 gnd.n3683 gnd.n2286 9.3005
R11005 gnd.n3682 gnd.n2288 9.3005
R11006 gnd.n3679 gnd.n2289 9.3005
R11007 gnd.n3678 gnd.n2290 9.3005
R11008 gnd.n3675 gnd.n2291 9.3005
R11009 gnd.n3674 gnd.n2292 9.3005
R11010 gnd.n3671 gnd.n2293 9.3005
R11011 gnd.n3670 gnd.n2294 9.3005
R11012 gnd.n3667 gnd.n2295 9.3005
R11013 gnd.n3666 gnd.n2296 9.3005
R11014 gnd.n3663 gnd.n2297 9.3005
R11015 gnd.n3662 gnd.n2298 9.3005
R11016 gnd.n3659 gnd.n2299 9.3005
R11017 gnd.n3658 gnd.n2300 9.3005
R11018 gnd.n3655 gnd.n2301 9.3005
R11019 gnd.n3654 gnd.n2302 9.3005
R11020 gnd.n3651 gnd.n2303 9.3005
R11021 gnd.n3650 gnd.n2304 9.3005
R11022 gnd.n3647 gnd.n2305 9.3005
R11023 gnd.n3646 gnd.n2306 9.3005
R11024 gnd.n3643 gnd.n2307 9.3005
R11025 gnd.n3642 gnd.n2308 9.3005
R11026 gnd.n3639 gnd.n2312 9.3005
R11027 gnd.n3638 gnd.n2313 9.3005
R11028 gnd.n3635 gnd.n2314 9.3005
R11029 gnd.n3634 gnd.n2315 9.3005
R11030 gnd.n3685 gnd.n3684 9.3005
R11031 gnd.n3136 gnd.n3120 9.3005
R11032 gnd.n3135 gnd.n3121 9.3005
R11033 gnd.n3134 gnd.n3122 9.3005
R11034 gnd.n3132 gnd.n3123 9.3005
R11035 gnd.n3131 gnd.n3124 9.3005
R11036 gnd.n3129 gnd.n3125 9.3005
R11037 gnd.n3128 gnd.n3126 9.3005
R11038 gnd.n2422 gnd.n2421 9.3005
R11039 gnd.n3205 gnd.n3204 9.3005
R11040 gnd.n3206 gnd.n2420 9.3005
R11041 gnd.n3223 gnd.n3207 9.3005
R11042 gnd.n3222 gnd.n3208 9.3005
R11043 gnd.n3221 gnd.n3209 9.3005
R11044 gnd.n3219 gnd.n3210 9.3005
R11045 gnd.n3218 gnd.n3211 9.3005
R11046 gnd.n3216 gnd.n3212 9.3005
R11047 gnd.n3215 gnd.n3213 9.3005
R11048 gnd.n2366 gnd.n2365 9.3005
R11049 gnd.n3290 gnd.n3289 9.3005
R11050 gnd.n3291 gnd.n2364 9.3005
R11051 gnd.n3312 gnd.n3292 9.3005
R11052 gnd.n3311 gnd.n3293 9.3005
R11053 gnd.n3310 gnd.n3294 9.3005
R11054 gnd.n3307 gnd.n3295 9.3005
R11055 gnd.n3306 gnd.n3296 9.3005
R11056 gnd.n3304 gnd.n3297 9.3005
R11057 gnd.n3303 gnd.n3298 9.3005
R11058 gnd.n3301 gnd.n3300 9.3005
R11059 gnd.n3299 gnd.n2317 9.3005
R11060 gnd.n2877 gnd.n2876 9.3005
R11061 gnd.n2767 gnd.n2766 9.3005
R11062 gnd.n2891 gnd.n2890 9.3005
R11063 gnd.n2892 gnd.n2765 9.3005
R11064 gnd.n2894 gnd.n2893 9.3005
R11065 gnd.n2755 gnd.n2754 9.3005
R11066 gnd.n2907 gnd.n2906 9.3005
R11067 gnd.n2908 gnd.n2753 9.3005
R11068 gnd.n2940 gnd.n2909 9.3005
R11069 gnd.n2939 gnd.n2910 9.3005
R11070 gnd.n2938 gnd.n2911 9.3005
R11071 gnd.n2937 gnd.n2912 9.3005
R11072 gnd.n2934 gnd.n2913 9.3005
R11073 gnd.n2933 gnd.n2914 9.3005
R11074 gnd.n2932 gnd.n2915 9.3005
R11075 gnd.n2930 gnd.n2916 9.3005
R11076 gnd.n2929 gnd.n2917 9.3005
R11077 gnd.n2926 gnd.n2918 9.3005
R11078 gnd.n2925 gnd.n2919 9.3005
R11079 gnd.n2924 gnd.n2920 9.3005
R11080 gnd.n2922 gnd.n2921 9.3005
R11081 gnd.n2621 gnd.n2620 9.3005
R11082 gnd.n3038 gnd.n3037 9.3005
R11083 gnd.n3039 gnd.n2619 9.3005
R11084 gnd.n3043 gnd.n3040 9.3005
R11085 gnd.n3042 gnd.n3041 9.3005
R11086 gnd.n2543 gnd.n2542 9.3005
R11087 gnd.n3118 gnd.n3117 9.3005
R11088 gnd.n2875 gnd.n2776 9.3005
R11089 gnd.n2778 gnd.n2777 9.3005
R11090 gnd.n2822 gnd.n2820 9.3005
R11091 gnd.n2823 gnd.n2819 9.3005
R11092 gnd.n2826 gnd.n2815 9.3005
R11093 gnd.n2827 gnd.n2814 9.3005
R11094 gnd.n2830 gnd.n2813 9.3005
R11095 gnd.n2831 gnd.n2812 9.3005
R11096 gnd.n2834 gnd.n2811 9.3005
R11097 gnd.n2835 gnd.n2810 9.3005
R11098 gnd.n2838 gnd.n2809 9.3005
R11099 gnd.n2839 gnd.n2808 9.3005
R11100 gnd.n2842 gnd.n2807 9.3005
R11101 gnd.n2843 gnd.n2806 9.3005
R11102 gnd.n2846 gnd.n2805 9.3005
R11103 gnd.n2847 gnd.n2804 9.3005
R11104 gnd.n2850 gnd.n2803 9.3005
R11105 gnd.n2851 gnd.n2802 9.3005
R11106 gnd.n2854 gnd.n2801 9.3005
R11107 gnd.n2855 gnd.n2800 9.3005
R11108 gnd.n2858 gnd.n2799 9.3005
R11109 gnd.n2859 gnd.n2798 9.3005
R11110 gnd.n2862 gnd.n2797 9.3005
R11111 gnd.n2864 gnd.n2796 9.3005
R11112 gnd.n2865 gnd.n2795 9.3005
R11113 gnd.n2866 gnd.n2794 9.3005
R11114 gnd.n2867 gnd.n2793 9.3005
R11115 gnd.n2874 gnd.n2873 9.3005
R11116 gnd.n2883 gnd.n2882 9.3005
R11117 gnd.n2884 gnd.n2770 9.3005
R11118 gnd.n2886 gnd.n2885 9.3005
R11119 gnd.n2761 gnd.n2760 9.3005
R11120 gnd.n2899 gnd.n2898 9.3005
R11121 gnd.n2900 gnd.n2759 9.3005
R11122 gnd.n2902 gnd.n2901 9.3005
R11123 gnd.n2748 gnd.n2747 9.3005
R11124 gnd.n2945 gnd.n2944 9.3005
R11125 gnd.n2946 gnd.n2702 9.3005
R11126 gnd.n2950 gnd.n2948 9.3005
R11127 gnd.n2949 gnd.n2681 9.3005
R11128 gnd.n2968 gnd.n2680 9.3005
R11129 gnd.n2971 gnd.n2970 9.3005
R11130 gnd.n2674 gnd.n2673 9.3005
R11131 gnd.n2982 gnd.n2980 9.3005
R11132 gnd.n2981 gnd.n2655 9.3005
R11133 gnd.n2999 gnd.n2654 9.3005
R11134 gnd.n3002 gnd.n3001 9.3005
R11135 gnd.n2649 gnd.n2644 9.3005
R11136 gnd.n3012 gnd.n3011 9.3005
R11137 gnd.n2647 gnd.n2627 9.3005
R11138 gnd.n3033 gnd.n2628 9.3005
R11139 gnd.n3032 gnd.n3031 9.3005
R11140 gnd.n2630 gnd.n2606 9.3005
R11141 gnd.n3064 gnd.n3063 9.3005
R11142 gnd.n3066 gnd.n2551 9.3005
R11143 gnd.n3113 gnd.n2552 9.3005
R11144 gnd.n3112 gnd.n2553 9.3005
R11145 gnd.n3111 gnd.n2554 9.3005
R11146 gnd.n3077 gnd.n2555 9.3005
R11147 gnd.n3079 gnd.n2573 9.3005
R11148 gnd.n3099 gnd.n2574 9.3005
R11149 gnd.n3098 gnd.n2575 9.3005
R11150 gnd.n3097 gnd.n2576 9.3005
R11151 gnd.n3088 gnd.n2577 9.3005
R11152 gnd.n3089 gnd.n2460 9.3005
R11153 gnd.n3155 gnd.n3154 9.3005
R11154 gnd.n3156 gnd.n2453 9.3005
R11155 gnd.n3166 gnd.n3165 9.3005
R11156 gnd.n3168 gnd.n2449 9.3005
R11157 gnd.n3178 gnd.n2450 9.3005
R11158 gnd.n3177 gnd.n3176 9.3005
R11159 gnd.n3174 gnd.n2428 9.3005
R11160 gnd.n3200 gnd.n2429 9.3005
R11161 gnd.n3199 gnd.n3198 9.3005
R11162 gnd.n2431 gnd.n2405 9.3005
R11163 gnd.n3240 gnd.n3239 9.3005
R11164 gnd.n3241 gnd.n2398 9.3005
R11165 gnd.n3251 gnd.n3250 9.3005
R11166 gnd.n3253 gnd.n2394 9.3005
R11167 gnd.n3263 gnd.n2395 9.3005
R11168 gnd.n3262 gnd.n3261 9.3005
R11169 gnd.n3259 gnd.n2373 9.3005
R11170 gnd.n3285 gnd.n2374 9.3005
R11171 gnd.n3284 gnd.n3283 9.3005
R11172 gnd.n2376 gnd.n2351 9.3005
R11173 gnd.n3329 gnd.n3328 9.3005
R11174 gnd.n3330 gnd.n2344 9.3005
R11175 gnd.n3340 gnd.n3339 9.3005
R11176 gnd.n3598 gnd.n2340 9.3005
R11177 gnd.n3606 gnd.n2341 9.3005
R11178 gnd.n3605 gnd.n3604 9.3005
R11179 gnd.n2322 gnd.n2321 9.3005
R11180 gnd.n3629 gnd.n3628 9.3005
R11181 gnd.n2772 gnd.n2771 9.3005
R11182 gnd.n3875 gnd.n3844 9.3005
R11183 gnd.n3874 gnd.n3845 9.3005
R11184 gnd.n3872 gnd.n3846 9.3005
R11185 gnd.n3871 gnd.n3847 9.3005
R11186 gnd.n3869 gnd.n3848 9.3005
R11187 gnd.n3868 gnd.n3849 9.3005
R11188 gnd.n3866 gnd.n3850 9.3005
R11189 gnd.n3865 gnd.n3851 9.3005
R11190 gnd.n3863 gnd.n3852 9.3005
R11191 gnd.n3862 gnd.n3853 9.3005
R11192 gnd.n3860 gnd.n3854 9.3005
R11193 gnd.n3859 gnd.n3855 9.3005
R11194 gnd.n3857 gnd.n3856 9.3005
R11195 gnd.n2168 gnd.n2167 9.3005
R11196 gnd.n4126 gnd.n4125 9.3005
R11197 gnd.n4127 gnd.n2166 9.3005
R11198 gnd.n4131 gnd.n4128 9.3005
R11199 gnd.n4130 gnd.n4129 9.3005
R11200 gnd.n2143 gnd.n2142 9.3005
R11201 gnd.n4161 gnd.n4160 9.3005
R11202 gnd.n4162 gnd.n2141 9.3005
R11203 gnd.n4166 gnd.n4163 9.3005
R11204 gnd.n4165 gnd.n4164 9.3005
R11205 gnd.n2118 gnd.n2117 9.3005
R11206 gnd.n4196 gnd.n4195 9.3005
R11207 gnd.n4197 gnd.n2115 9.3005
R11208 gnd.n3878 gnd.n3877 9.3005
R11209 gnd.n5974 gnd.n1044 9.3005
R11210 gnd.n5977 gnd.n1043 9.3005
R11211 gnd.n5978 gnd.n1042 9.3005
R11212 gnd.n5981 gnd.n1041 9.3005
R11213 gnd.n5982 gnd.n1040 9.3005
R11214 gnd.n5985 gnd.n1039 9.3005
R11215 gnd.n5986 gnd.n1038 9.3005
R11216 gnd.n5989 gnd.n1037 9.3005
R11217 gnd.n5991 gnd.n1034 9.3005
R11218 gnd.n5994 gnd.n1033 9.3005
R11219 gnd.n5995 gnd.n1032 9.3005
R11220 gnd.n5998 gnd.n1031 9.3005
R11221 gnd.n5999 gnd.n1030 9.3005
R11222 gnd.n6002 gnd.n1029 9.3005
R11223 gnd.n6003 gnd.n1028 9.3005
R11224 gnd.n6006 gnd.n1027 9.3005
R11225 gnd.n6007 gnd.n1026 9.3005
R11226 gnd.n6010 gnd.n1025 9.3005
R11227 gnd.n6011 gnd.n1024 9.3005
R11228 gnd.n6014 gnd.n1023 9.3005
R11229 gnd.n6015 gnd.n1022 9.3005
R11230 gnd.n6018 gnd.n1021 9.3005
R11231 gnd.n6019 gnd.n1020 9.3005
R11232 gnd.n6020 gnd.n1019 9.3005
R11233 gnd.n976 gnd.n975 9.3005
R11234 gnd.n6026 gnd.n6025 9.3005
R11235 gnd.n4505 gnd.n4502 9.3005
R11236 gnd.n4509 gnd.n4508 9.3005
R11237 gnd.n4510 gnd.n4500 9.3005
R11238 gnd.n4512 gnd.n4511 9.3005
R11239 gnd.n4515 gnd.n4499 9.3005
R11240 gnd.n4519 gnd.n4518 9.3005
R11241 gnd.n4520 gnd.n4498 9.3005
R11242 gnd.n4523 gnd.n4521 9.3005
R11243 gnd.n4524 gnd.n4494 9.3005
R11244 gnd.n4528 gnd.n4527 9.3005
R11245 gnd.n4529 gnd.n4493 9.3005
R11246 gnd.n4531 gnd.n4530 9.3005
R11247 gnd.n4534 gnd.n4492 9.3005
R11248 gnd.n4538 gnd.n4537 9.3005
R11249 gnd.n4539 gnd.n4491 9.3005
R11250 gnd.n4541 gnd.n4540 9.3005
R11251 gnd.n4544 gnd.n4490 9.3005
R11252 gnd.n4548 gnd.n4547 9.3005
R11253 gnd.n4549 gnd.n4489 9.3005
R11254 gnd.n4551 gnd.n4550 9.3005
R11255 gnd.n4554 gnd.n4488 9.3005
R11256 gnd.n4558 gnd.n4557 9.3005
R11257 gnd.n4559 gnd.n4487 9.3005
R11258 gnd.n4561 gnd.n4560 9.3005
R11259 gnd.n4564 gnd.n4486 9.3005
R11260 gnd.n4568 gnd.n4567 9.3005
R11261 gnd.n4569 gnd.n4485 9.3005
R11262 gnd.n4572 gnd.n4570 9.3005
R11263 gnd.n4573 gnd.n4481 9.3005
R11264 gnd.n4576 gnd.n4575 9.3005
R11265 gnd.n4501 gnd.n1045 9.3005
R11266 gnd.n4256 gnd.n4255 9.3005
R11267 gnd.n4257 gnd.n2079 9.3005
R11268 gnd.n4260 gnd.n4259 9.3005
R11269 gnd.n4258 gnd.n890 9.3005
R11270 gnd.n6077 gnd.n891 9.3005
R11271 gnd.n6076 gnd.n892 9.3005
R11272 gnd.n6075 gnd.n893 9.3005
R11273 gnd.n912 gnd.n894 9.3005
R11274 gnd.n6065 gnd.n913 9.3005
R11275 gnd.n6064 gnd.n914 9.3005
R11276 gnd.n6063 gnd.n915 9.3005
R11277 gnd.n932 gnd.n916 9.3005
R11278 gnd.n6053 gnd.n933 9.3005
R11279 gnd.n6052 gnd.n934 9.3005
R11280 gnd.n6051 gnd.n935 9.3005
R11281 gnd.n952 gnd.n936 9.3005
R11282 gnd.n6041 gnd.n953 9.3005
R11283 gnd.n6040 gnd.n954 9.3005
R11284 gnd.n6039 gnd.n955 9.3005
R11285 gnd.n973 gnd.n956 9.3005
R11286 gnd.n6029 gnd.n974 9.3005
R11287 gnd.n6028 gnd.n6027 9.3005
R11288 gnd.n2127 gnd.n2126 9.3005
R11289 gnd.n4186 gnd.n4185 9.3005
R11290 gnd.n4187 gnd.n2125 9.3005
R11291 gnd.n4191 gnd.n4188 9.3005
R11292 gnd.n4190 gnd.n4189 9.3005
R11293 gnd.n2102 gnd.n2101 9.3005
R11294 gnd.n4229 gnd.n4228 9.3005
R11295 gnd.n4230 gnd.n2100 9.3005
R11296 gnd.n4232 gnd.n4231 9.3005
R11297 gnd.n2081 gnd.n2080 9.3005
R11298 gnd.n4052 gnd.n4051 9.3005
R11299 gnd.n4053 gnd.n2230 9.3005
R11300 gnd.n4055 gnd.n4054 9.3005
R11301 gnd.n2213 gnd.n2212 9.3005
R11302 gnd.n4072 gnd.n4071 9.3005
R11303 gnd.n4073 gnd.n2211 9.3005
R11304 gnd.n4075 gnd.n4074 9.3005
R11305 gnd.n2196 gnd.n2195 9.3005
R11306 gnd.n4092 gnd.n4091 9.3005
R11307 gnd.n4093 gnd.n2194 9.3005
R11308 gnd.n4095 gnd.n4094 9.3005
R11309 gnd.n2176 gnd.n2175 9.3005
R11310 gnd.n4116 gnd.n4115 9.3005
R11311 gnd.n4117 gnd.n2174 9.3005
R11312 gnd.n4121 gnd.n4118 9.3005
R11313 gnd.n4120 gnd.n4119 9.3005
R11314 gnd.n2151 gnd.n2150 9.3005
R11315 gnd.n4151 gnd.n4150 9.3005
R11316 gnd.n4152 gnd.n2149 9.3005
R11317 gnd.n4156 gnd.n4153 9.3005
R11318 gnd.n4155 gnd.n4154 9.3005
R11319 gnd.n2232 gnd.n2231 9.3005
R11320 gnd.n3921 gnd.n3920 9.3005
R11321 gnd.n3923 gnd.n3822 9.3005
R11322 gnd.n3924 gnd.n3821 9.3005
R11323 gnd.n3927 gnd.n3820 9.3005
R11324 gnd.n3928 gnd.n3819 9.3005
R11325 gnd.n3931 gnd.n3818 9.3005
R11326 gnd.n3932 gnd.n3817 9.3005
R11327 gnd.n3935 gnd.n3816 9.3005
R11328 gnd.n3936 gnd.n3815 9.3005
R11329 gnd.n3939 gnd.n3814 9.3005
R11330 gnd.n3940 gnd.n3813 9.3005
R11331 gnd.n3943 gnd.n3812 9.3005
R11332 gnd.n3944 gnd.n3811 9.3005
R11333 gnd.n3947 gnd.n3810 9.3005
R11334 gnd.n3948 gnd.n3809 9.3005
R11335 gnd.n3951 gnd.n3808 9.3005
R11336 gnd.n3952 gnd.n3807 9.3005
R11337 gnd.n3955 gnd.n3806 9.3005
R11338 gnd.n3956 gnd.n3805 9.3005
R11339 gnd.n3959 gnd.n3804 9.3005
R11340 gnd.n3963 gnd.n3800 9.3005
R11341 gnd.n3964 gnd.n3799 9.3005
R11342 gnd.n3967 gnd.n3798 9.3005
R11343 gnd.n3968 gnd.n3797 9.3005
R11344 gnd.n3971 gnd.n3796 9.3005
R11345 gnd.n3972 gnd.n3795 9.3005
R11346 gnd.n3975 gnd.n3794 9.3005
R11347 gnd.n3976 gnd.n3793 9.3005
R11348 gnd.n3979 gnd.n3792 9.3005
R11349 gnd.n3980 gnd.n3791 9.3005
R11350 gnd.n3983 gnd.n3790 9.3005
R11351 gnd.n3984 gnd.n3789 9.3005
R11352 gnd.n3987 gnd.n3788 9.3005
R11353 gnd.n3988 gnd.n3787 9.3005
R11354 gnd.n3991 gnd.n3786 9.3005
R11355 gnd.n3992 gnd.n3785 9.3005
R11356 gnd.n3995 gnd.n3784 9.3005
R11357 gnd.n3996 gnd.n3783 9.3005
R11358 gnd.n3999 gnd.n3782 9.3005
R11359 gnd.n4001 gnd.n3779 9.3005
R11360 gnd.n4004 gnd.n3778 9.3005
R11361 gnd.n4005 gnd.n3777 9.3005
R11362 gnd.n4008 gnd.n3776 9.3005
R11363 gnd.n4009 gnd.n3775 9.3005
R11364 gnd.n4012 gnd.n3774 9.3005
R11365 gnd.n4013 gnd.n3773 9.3005
R11366 gnd.n4016 gnd.n3772 9.3005
R11367 gnd.n4017 gnd.n3771 9.3005
R11368 gnd.n4020 gnd.n3770 9.3005
R11369 gnd.n4021 gnd.n3769 9.3005
R11370 gnd.n4024 gnd.n3768 9.3005
R11371 gnd.n4025 gnd.n3767 9.3005
R11372 gnd.n4028 gnd.n3766 9.3005
R11373 gnd.n4030 gnd.n3765 9.3005
R11374 gnd.n4031 gnd.n3764 9.3005
R11375 gnd.n4032 gnd.n3763 9.3005
R11376 gnd.n4033 gnd.n3762 9.3005
R11377 gnd.n3960 gnd.n3801 9.3005
R11378 gnd.n3919 gnd.n2242 9.3005
R11379 gnd.n3883 gnd.n3882 9.3005
R11380 gnd.n3886 gnd.n3839 9.3005
R11381 gnd.n3887 gnd.n3838 9.3005
R11382 gnd.n3890 gnd.n3837 9.3005
R11383 gnd.n3891 gnd.n3836 9.3005
R11384 gnd.n3894 gnd.n3835 9.3005
R11385 gnd.n3895 gnd.n3834 9.3005
R11386 gnd.n3898 gnd.n3833 9.3005
R11387 gnd.n3899 gnd.n3832 9.3005
R11388 gnd.n3902 gnd.n3831 9.3005
R11389 gnd.n3903 gnd.n3830 9.3005
R11390 gnd.n3906 gnd.n3829 9.3005
R11391 gnd.n3907 gnd.n3828 9.3005
R11392 gnd.n3910 gnd.n3827 9.3005
R11393 gnd.n3911 gnd.n3826 9.3005
R11394 gnd.n3914 gnd.n3825 9.3005
R11395 gnd.n3917 gnd.n3916 9.3005
R11396 gnd.n3881 gnd.n3843 9.3005
R11397 gnd.n3880 gnd.n3879 9.3005
R11398 gnd.n4041 gnd.n2240 9.3005
R11399 gnd.n4043 gnd.n4042 9.3005
R11400 gnd.n4044 gnd.n2223 9.3005
R11401 gnd.n4060 gnd.n2224 9.3005
R11402 gnd.n4061 gnd.n2222 9.3005
R11403 gnd.n4063 gnd.n4062 9.3005
R11404 gnd.n4064 gnd.n2205 9.3005
R11405 gnd.n4080 gnd.n2206 9.3005
R11406 gnd.n4081 gnd.n2204 9.3005
R11407 gnd.n4083 gnd.n4082 9.3005
R11408 gnd.n4084 gnd.n2187 9.3005
R11409 gnd.n4100 gnd.n2188 9.3005
R11410 gnd.n4101 gnd.n2185 9.3005
R11411 gnd.n4103 gnd.n2186 9.3005
R11412 gnd.n4105 gnd.n4104 9.3005
R11413 gnd.n4106 gnd.n2161 9.3005
R11414 gnd.n4135 gnd.n2162 9.3005
R11415 gnd.n4136 gnd.n2159 9.3005
R11416 gnd.n4138 gnd.n2160 9.3005
R11417 gnd.n4140 gnd.n4139 9.3005
R11418 gnd.n4141 gnd.n2136 9.3005
R11419 gnd.n4170 gnd.n2137 9.3005
R11420 gnd.n4171 gnd.n2134 9.3005
R11421 gnd.n4173 gnd.n2135 9.3005
R11422 gnd.n4175 gnd.n4174 9.3005
R11423 gnd.n4176 gnd.n2110 9.3005
R11424 gnd.n4217 gnd.n2111 9.3005
R11425 gnd.n4218 gnd.n2109 9.3005
R11426 gnd.n4220 gnd.n4219 9.3005
R11427 gnd.n4221 gnd.n2093 9.3005
R11428 gnd.n4237 gnd.n2094 9.3005
R11429 gnd.n4238 gnd.n2090 9.3005
R11430 gnd.n4240 gnd.n2091 9.3005
R11431 gnd.n4241 gnd.n2092 9.3005
R11432 gnd.n4244 gnd.n4243 9.3005
R11433 gnd.n4245 gnd.n2070 9.3005
R11434 gnd.n4273 gnd.n2071 9.3005
R11435 gnd.n4274 gnd.n902 9.3005
R11436 gnd.n4275 gnd.n903 9.3005
R11437 gnd.n4276 gnd.n904 9.3005
R11438 gnd.n4280 gnd.n4277 9.3005
R11439 gnd.n4279 gnd.n923 9.3005
R11440 gnd.n4278 gnd.n924 9.3005
R11441 gnd.n2055 gnd.n925 9.3005
R11442 gnd.n4326 gnd.n2056 9.3005
R11443 gnd.n4327 gnd.n942 9.3005
R11444 gnd.n4328 gnd.n943 9.3005
R11445 gnd.n4329 gnd.n944 9.3005
R11446 gnd.n4333 gnd.n4330 9.3005
R11447 gnd.n4334 gnd.n963 9.3005
R11448 gnd.n4581 gnd.n964 9.3005
R11449 gnd.n4580 gnd.n965 9.3005
R11450 gnd.n4579 gnd.n4578 9.3005
R11451 gnd.n4040 gnd.n2241 9.3005
R11452 gnd.n4047 gnd.n2240 9.3005
R11453 gnd.n4046 gnd.n4043 9.3005
R11454 gnd.n4045 gnd.n4044 9.3005
R11455 gnd.n2224 gnd.n2221 9.3005
R11456 gnd.n4067 gnd.n2222 9.3005
R11457 gnd.n4066 gnd.n4063 9.3005
R11458 gnd.n4065 gnd.n4064 9.3005
R11459 gnd.n2206 gnd.n2203 9.3005
R11460 gnd.n4087 gnd.n2204 9.3005
R11461 gnd.n4086 gnd.n4083 9.3005
R11462 gnd.n4085 gnd.n4084 9.3005
R11463 gnd.n2188 gnd.n2184 9.3005
R11464 gnd.n4111 gnd.n2185 9.3005
R11465 gnd.n4110 gnd.n2186 9.3005
R11466 gnd.n4109 gnd.n4105 9.3005
R11467 gnd.n4108 gnd.n4106 9.3005
R11468 gnd.n2162 gnd.n2158 9.3005
R11469 gnd.n4146 gnd.n2159 9.3005
R11470 gnd.n4145 gnd.n2160 9.3005
R11471 gnd.n4144 gnd.n4140 9.3005
R11472 gnd.n4143 gnd.n4141 9.3005
R11473 gnd.n2137 gnd.n2133 9.3005
R11474 gnd.n4181 gnd.n2134 9.3005
R11475 gnd.n4180 gnd.n2135 9.3005
R11476 gnd.n4179 gnd.n4175 9.3005
R11477 gnd.n4178 gnd.n4176 9.3005
R11478 gnd.n2111 gnd.n2108 9.3005
R11479 gnd.n4224 gnd.n2109 9.3005
R11480 gnd.n4223 gnd.n4220 9.3005
R11481 gnd.n4222 gnd.n4221 9.3005
R11482 gnd.n2094 gnd.n2089 9.3005
R11483 gnd.n4251 gnd.n2090 9.3005
R11484 gnd.n4250 gnd.n2091 9.3005
R11485 gnd.n4249 gnd.n2092 9.3005
R11486 gnd.n4248 gnd.n4244 9.3005
R11487 gnd.n4246 gnd.n4245 9.3005
R11488 gnd.n2071 gnd.n901 9.3005
R11489 gnd.n6071 gnd.n902 9.3005
R11490 gnd.n6070 gnd.n903 9.3005
R11491 gnd.n6069 gnd.n904 9.3005
R11492 gnd.n4277 gnd.n905 9.3005
R11493 gnd.n6059 gnd.n923 9.3005
R11494 gnd.n6058 gnd.n924 9.3005
R11495 gnd.n6057 gnd.n925 9.3005
R11496 gnd.n2056 gnd.n926 9.3005
R11497 gnd.n6047 gnd.n942 9.3005
R11498 gnd.n6046 gnd.n943 9.3005
R11499 gnd.n6045 gnd.n944 9.3005
R11500 gnd.n4330 gnd.n945 9.3005
R11501 gnd.n6035 gnd.n963 9.3005
R11502 gnd.n6034 gnd.n964 9.3005
R11503 gnd.n6033 gnd.n965 9.3005
R11504 gnd.n4578 gnd.n966 9.3005
R11505 gnd.n2241 gnd.n2239 9.3005
R11506 gnd.n6252 gnd.n713 9.3005
R11507 gnd.n6254 gnd.n6253 9.3005
R11508 gnd.n709 gnd.n708 9.3005
R11509 gnd.n6261 gnd.n6260 9.3005
R11510 gnd.n6262 gnd.n707 9.3005
R11511 gnd.n6264 gnd.n6263 9.3005
R11512 gnd.n703 gnd.n702 9.3005
R11513 gnd.n6271 gnd.n6270 9.3005
R11514 gnd.n6272 gnd.n701 9.3005
R11515 gnd.n6274 gnd.n6273 9.3005
R11516 gnd.n697 gnd.n696 9.3005
R11517 gnd.n6281 gnd.n6280 9.3005
R11518 gnd.n6282 gnd.n695 9.3005
R11519 gnd.n6284 gnd.n6283 9.3005
R11520 gnd.n691 gnd.n690 9.3005
R11521 gnd.n6291 gnd.n6290 9.3005
R11522 gnd.n6292 gnd.n689 9.3005
R11523 gnd.n6294 gnd.n6293 9.3005
R11524 gnd.n685 gnd.n684 9.3005
R11525 gnd.n6301 gnd.n6300 9.3005
R11526 gnd.n6302 gnd.n683 9.3005
R11527 gnd.n6304 gnd.n6303 9.3005
R11528 gnd.n679 gnd.n678 9.3005
R11529 gnd.n6311 gnd.n6310 9.3005
R11530 gnd.n6312 gnd.n677 9.3005
R11531 gnd.n6314 gnd.n6313 9.3005
R11532 gnd.n673 gnd.n672 9.3005
R11533 gnd.n6321 gnd.n6320 9.3005
R11534 gnd.n6322 gnd.n671 9.3005
R11535 gnd.n6324 gnd.n6323 9.3005
R11536 gnd.n667 gnd.n666 9.3005
R11537 gnd.n6331 gnd.n6330 9.3005
R11538 gnd.n6332 gnd.n665 9.3005
R11539 gnd.n6334 gnd.n6333 9.3005
R11540 gnd.n661 gnd.n660 9.3005
R11541 gnd.n6341 gnd.n6340 9.3005
R11542 gnd.n6342 gnd.n659 9.3005
R11543 gnd.n6344 gnd.n6343 9.3005
R11544 gnd.n655 gnd.n654 9.3005
R11545 gnd.n6351 gnd.n6350 9.3005
R11546 gnd.n6352 gnd.n653 9.3005
R11547 gnd.n6354 gnd.n6353 9.3005
R11548 gnd.n649 gnd.n648 9.3005
R11549 gnd.n6361 gnd.n6360 9.3005
R11550 gnd.n6362 gnd.n647 9.3005
R11551 gnd.n6364 gnd.n6363 9.3005
R11552 gnd.n643 gnd.n642 9.3005
R11553 gnd.n6371 gnd.n6370 9.3005
R11554 gnd.n6372 gnd.n641 9.3005
R11555 gnd.n6374 gnd.n6373 9.3005
R11556 gnd.n637 gnd.n636 9.3005
R11557 gnd.n6381 gnd.n6380 9.3005
R11558 gnd.n6382 gnd.n635 9.3005
R11559 gnd.n6384 gnd.n6383 9.3005
R11560 gnd.n631 gnd.n630 9.3005
R11561 gnd.n6391 gnd.n6390 9.3005
R11562 gnd.n6392 gnd.n629 9.3005
R11563 gnd.n6394 gnd.n6393 9.3005
R11564 gnd.n625 gnd.n624 9.3005
R11565 gnd.n6401 gnd.n6400 9.3005
R11566 gnd.n6402 gnd.n623 9.3005
R11567 gnd.n6404 gnd.n6403 9.3005
R11568 gnd.n619 gnd.n618 9.3005
R11569 gnd.n6411 gnd.n6410 9.3005
R11570 gnd.n6412 gnd.n617 9.3005
R11571 gnd.n6414 gnd.n6413 9.3005
R11572 gnd.n613 gnd.n612 9.3005
R11573 gnd.n6421 gnd.n6420 9.3005
R11574 gnd.n6422 gnd.n611 9.3005
R11575 gnd.n6424 gnd.n6423 9.3005
R11576 gnd.n607 gnd.n606 9.3005
R11577 gnd.n6431 gnd.n6430 9.3005
R11578 gnd.n6432 gnd.n605 9.3005
R11579 gnd.n6434 gnd.n6433 9.3005
R11580 gnd.n601 gnd.n600 9.3005
R11581 gnd.n6441 gnd.n6440 9.3005
R11582 gnd.n6442 gnd.n599 9.3005
R11583 gnd.n6444 gnd.n6443 9.3005
R11584 gnd.n595 gnd.n594 9.3005
R11585 gnd.n6451 gnd.n6450 9.3005
R11586 gnd.n6452 gnd.n593 9.3005
R11587 gnd.n6454 gnd.n6453 9.3005
R11588 gnd.n589 gnd.n588 9.3005
R11589 gnd.n6461 gnd.n6460 9.3005
R11590 gnd.n6462 gnd.n587 9.3005
R11591 gnd.n6464 gnd.n6463 9.3005
R11592 gnd.n583 gnd.n582 9.3005
R11593 gnd.n6471 gnd.n6470 9.3005
R11594 gnd.n6472 gnd.n581 9.3005
R11595 gnd.n6474 gnd.n6473 9.3005
R11596 gnd.n577 gnd.n576 9.3005
R11597 gnd.n6481 gnd.n6480 9.3005
R11598 gnd.n6482 gnd.n575 9.3005
R11599 gnd.n6484 gnd.n6483 9.3005
R11600 gnd.n571 gnd.n570 9.3005
R11601 gnd.n6491 gnd.n6490 9.3005
R11602 gnd.n6492 gnd.n569 9.3005
R11603 gnd.n6494 gnd.n6493 9.3005
R11604 gnd.n565 gnd.n564 9.3005
R11605 gnd.n6501 gnd.n6500 9.3005
R11606 gnd.n6502 gnd.n563 9.3005
R11607 gnd.n6504 gnd.n6503 9.3005
R11608 gnd.n559 gnd.n558 9.3005
R11609 gnd.n6511 gnd.n6510 9.3005
R11610 gnd.n6512 gnd.n557 9.3005
R11611 gnd.n6514 gnd.n6513 9.3005
R11612 gnd.n553 gnd.n552 9.3005
R11613 gnd.n6521 gnd.n6520 9.3005
R11614 gnd.n6522 gnd.n551 9.3005
R11615 gnd.n6524 gnd.n6523 9.3005
R11616 gnd.n547 gnd.n546 9.3005
R11617 gnd.n6531 gnd.n6530 9.3005
R11618 gnd.n6532 gnd.n545 9.3005
R11619 gnd.n6534 gnd.n6533 9.3005
R11620 gnd.n541 gnd.n540 9.3005
R11621 gnd.n6541 gnd.n6540 9.3005
R11622 gnd.n6542 gnd.n539 9.3005
R11623 gnd.n6544 gnd.n6543 9.3005
R11624 gnd.n535 gnd.n534 9.3005
R11625 gnd.n6551 gnd.n6550 9.3005
R11626 gnd.n6552 gnd.n533 9.3005
R11627 gnd.n6554 gnd.n6553 9.3005
R11628 gnd.n529 gnd.n528 9.3005
R11629 gnd.n6561 gnd.n6560 9.3005
R11630 gnd.n6562 gnd.n527 9.3005
R11631 gnd.n6565 gnd.n6564 9.3005
R11632 gnd.n6563 gnd.n523 9.3005
R11633 gnd.n6571 gnd.n522 9.3005
R11634 gnd.n6573 gnd.n6572 9.3005
R11635 gnd.n518 gnd.n517 9.3005
R11636 gnd.n6582 gnd.n6581 9.3005
R11637 gnd.n6583 gnd.n516 9.3005
R11638 gnd.n6585 gnd.n6584 9.3005
R11639 gnd.n512 gnd.n511 9.3005
R11640 gnd.n6592 gnd.n6591 9.3005
R11641 gnd.n6593 gnd.n510 9.3005
R11642 gnd.n6595 gnd.n6594 9.3005
R11643 gnd.n506 gnd.n505 9.3005
R11644 gnd.n6602 gnd.n6601 9.3005
R11645 gnd.n6603 gnd.n504 9.3005
R11646 gnd.n6605 gnd.n6604 9.3005
R11647 gnd.n500 gnd.n499 9.3005
R11648 gnd.n6612 gnd.n6611 9.3005
R11649 gnd.n6613 gnd.n498 9.3005
R11650 gnd.n6615 gnd.n6614 9.3005
R11651 gnd.n494 gnd.n493 9.3005
R11652 gnd.n6622 gnd.n6621 9.3005
R11653 gnd.n6623 gnd.n492 9.3005
R11654 gnd.n6625 gnd.n6624 9.3005
R11655 gnd.n488 gnd.n487 9.3005
R11656 gnd.n6632 gnd.n6631 9.3005
R11657 gnd.n6633 gnd.n486 9.3005
R11658 gnd.n6635 gnd.n6634 9.3005
R11659 gnd.n482 gnd.n481 9.3005
R11660 gnd.n6642 gnd.n6641 9.3005
R11661 gnd.n6643 gnd.n480 9.3005
R11662 gnd.n6645 gnd.n6644 9.3005
R11663 gnd.n476 gnd.n475 9.3005
R11664 gnd.n6652 gnd.n6651 9.3005
R11665 gnd.n6653 gnd.n474 9.3005
R11666 gnd.n6655 gnd.n6654 9.3005
R11667 gnd.n470 gnd.n469 9.3005
R11668 gnd.n6662 gnd.n6661 9.3005
R11669 gnd.n6663 gnd.n468 9.3005
R11670 gnd.n6665 gnd.n6664 9.3005
R11671 gnd.n464 gnd.n463 9.3005
R11672 gnd.n6672 gnd.n6671 9.3005
R11673 gnd.n6673 gnd.n462 9.3005
R11674 gnd.n6675 gnd.n6674 9.3005
R11675 gnd.n458 gnd.n457 9.3005
R11676 gnd.n6682 gnd.n6681 9.3005
R11677 gnd.n6683 gnd.n456 9.3005
R11678 gnd.n6685 gnd.n6684 9.3005
R11679 gnd.n452 gnd.n451 9.3005
R11680 gnd.n6692 gnd.n6691 9.3005
R11681 gnd.n6693 gnd.n450 9.3005
R11682 gnd.n6695 gnd.n6694 9.3005
R11683 gnd.n446 gnd.n445 9.3005
R11684 gnd.n6702 gnd.n6701 9.3005
R11685 gnd.n6703 gnd.n444 9.3005
R11686 gnd.n6705 gnd.n6704 9.3005
R11687 gnd.n440 gnd.n439 9.3005
R11688 gnd.n6712 gnd.n6711 9.3005
R11689 gnd.n6713 gnd.n438 9.3005
R11690 gnd.n6715 gnd.n6714 9.3005
R11691 gnd.n434 gnd.n433 9.3005
R11692 gnd.n6722 gnd.n6721 9.3005
R11693 gnd.n6723 gnd.n432 9.3005
R11694 gnd.n6725 gnd.n6724 9.3005
R11695 gnd.n428 gnd.n427 9.3005
R11696 gnd.n6732 gnd.n6731 9.3005
R11697 gnd.n6733 gnd.n426 9.3005
R11698 gnd.n6735 gnd.n6734 9.3005
R11699 gnd.n422 gnd.n421 9.3005
R11700 gnd.n6742 gnd.n6741 9.3005
R11701 gnd.n6743 gnd.n420 9.3005
R11702 gnd.n6745 gnd.n6744 9.3005
R11703 gnd.n416 gnd.n415 9.3005
R11704 gnd.n6752 gnd.n6751 9.3005
R11705 gnd.n6753 gnd.n414 9.3005
R11706 gnd.n6755 gnd.n6754 9.3005
R11707 gnd.n410 gnd.n409 9.3005
R11708 gnd.n6762 gnd.n6761 9.3005
R11709 gnd.n6763 gnd.n408 9.3005
R11710 gnd.n6765 gnd.n6764 9.3005
R11711 gnd.n404 gnd.n403 9.3005
R11712 gnd.n6772 gnd.n6771 9.3005
R11713 gnd.n6773 gnd.n402 9.3005
R11714 gnd.n6775 gnd.n6774 9.3005
R11715 gnd.n398 gnd.n397 9.3005
R11716 gnd.n6783 gnd.n6782 9.3005
R11717 gnd.n6784 gnd.n396 9.3005
R11718 gnd.n6786 gnd.n6785 9.3005
R11719 gnd.n6575 gnd.n6574 9.3005
R11720 gnd.n4298 gnd.n4297 9.3005
R11721 gnd.n4299 gnd.n4293 9.3005
R11722 gnd.n4301 gnd.n4300 9.3005
R11723 gnd.n2065 gnd.n2064 9.3005
R11724 gnd.n4306 gnd.n4305 9.3005
R11725 gnd.n4307 gnd.n2063 9.3005
R11726 gnd.n4313 gnd.n4308 9.3005
R11727 gnd.n4312 gnd.n4309 9.3005
R11728 gnd.n4311 gnd.n4310 9.3005
R11729 gnd.n2047 gnd.n2046 9.3005
R11730 gnd.n4601 gnd.n4600 9.3005
R11731 gnd.n4602 gnd.n2045 9.3005
R11732 gnd.n4604 gnd.n4603 9.3005
R11733 gnd.n2043 gnd.n2042 9.3005
R11734 gnd.n4609 gnd.n4608 9.3005
R11735 gnd.n4610 gnd.n2041 9.3005
R11736 gnd.n4620 gnd.n4611 9.3005
R11737 gnd.n4619 gnd.n4612 9.3005
R11738 gnd.n4618 gnd.n4613 9.3005
R11739 gnd.n4615 gnd.n4614 9.3005
R11740 gnd.n2013 gnd.n2012 9.3005
R11741 gnd.n4637 gnd.n4636 9.3005
R11742 gnd.n4638 gnd.n2011 9.3005
R11743 gnd.n4640 gnd.n4639 9.3005
R11744 gnd.n1997 gnd.n1996 9.3005
R11745 gnd.n4670 gnd.n4669 9.3005
R11746 gnd.n4671 gnd.n1995 9.3005
R11747 gnd.n4682 gnd.n4672 9.3005
R11748 gnd.n4681 gnd.n4673 9.3005
R11749 gnd.n4680 gnd.n4674 9.3005
R11750 gnd.n4677 gnd.n4676 9.3005
R11751 gnd.n4675 gnd.n1118 9.3005
R11752 gnd.n5895 gnd.n1119 9.3005
R11753 gnd.n5894 gnd.n1120 9.3005
R11754 gnd.n5893 gnd.n1121 9.3005
R11755 gnd.n4866 gnd.n1122 9.3005
R11756 gnd.n4867 gnd.n4865 9.3005
R11757 gnd.n4869 gnd.n4868 9.3005
R11758 gnd.n1886 gnd.n1885 9.3005
R11759 gnd.n4895 gnd.n4894 9.3005
R11760 gnd.n4896 gnd.n1884 9.3005
R11761 gnd.n4909 gnd.n4897 9.3005
R11762 gnd.n4908 gnd.n4898 9.3005
R11763 gnd.n4907 gnd.n4899 9.3005
R11764 gnd.n4901 gnd.n4900 9.3005
R11765 gnd.n4903 gnd.n4902 9.3005
R11766 gnd.n1848 gnd.n1847 9.3005
R11767 gnd.n4953 gnd.n4952 9.3005
R11768 gnd.n4954 gnd.n1846 9.3005
R11769 gnd.n4956 gnd.n4955 9.3005
R11770 gnd.n1830 gnd.n1829 9.3005
R11771 gnd.n4979 gnd.n4978 9.3005
R11772 gnd.n4980 gnd.n1828 9.3005
R11773 gnd.n4984 gnd.n4981 9.3005
R11774 gnd.n4983 gnd.n4982 9.3005
R11775 gnd.n1806 gnd.n1805 9.3005
R11776 gnd.n5018 gnd.n5017 9.3005
R11777 gnd.n5019 gnd.n1804 9.3005
R11778 gnd.n5032 gnd.n5020 9.3005
R11779 gnd.n5031 gnd.n5021 9.3005
R11780 gnd.n5030 gnd.n5022 9.3005
R11781 gnd.n5024 gnd.n5023 9.3005
R11782 gnd.n5026 gnd.n5025 9.3005
R11783 gnd.n1767 gnd.n1766 9.3005
R11784 gnd.n5076 gnd.n5075 9.3005
R11785 gnd.n5077 gnd.n1765 9.3005
R11786 gnd.n5079 gnd.n5078 9.3005
R11787 gnd.n1748 gnd.n1747 9.3005
R11788 gnd.n5101 gnd.n5100 9.3005
R11789 gnd.n5102 gnd.n1746 9.3005
R11790 gnd.n5106 gnd.n5103 9.3005
R11791 gnd.n5105 gnd.n5104 9.3005
R11792 gnd.n1723 gnd.n1722 9.3005
R11793 gnd.n5139 gnd.n5138 9.3005
R11794 gnd.n5140 gnd.n1721 9.3005
R11795 gnd.n5150 gnd.n5141 9.3005
R11796 gnd.n5149 gnd.n5142 9.3005
R11797 gnd.n5148 gnd.n5143 9.3005
R11798 gnd.n5145 gnd.n5144 9.3005
R11799 gnd.n1689 gnd.n1688 9.3005
R11800 gnd.n5185 gnd.n5184 9.3005
R11801 gnd.n5186 gnd.n1687 9.3005
R11802 gnd.n5190 gnd.n5187 9.3005
R11803 gnd.n5189 gnd.n5188 9.3005
R11804 gnd.n1661 gnd.n1660 9.3005
R11805 gnd.n5220 gnd.n5219 9.3005
R11806 gnd.n5221 gnd.n1659 9.3005
R11807 gnd.n5223 gnd.n5222 9.3005
R11808 gnd.n1632 gnd.n1631 9.3005
R11809 gnd.n5257 gnd.n5256 9.3005
R11810 gnd.n5258 gnd.n1630 9.3005
R11811 gnd.n5262 gnd.n5259 9.3005
R11812 gnd.n5261 gnd.n5260 9.3005
R11813 gnd.n1532 gnd.n1531 9.3005
R11814 gnd.n5407 gnd.n5406 9.3005
R11815 gnd.n5408 gnd.n1530 9.3005
R11816 gnd.n5410 gnd.n5409 9.3005
R11817 gnd.n1519 gnd.n1518 9.3005
R11818 gnd.n5423 gnd.n5422 9.3005
R11819 gnd.n5424 gnd.n1517 9.3005
R11820 gnd.n5429 gnd.n5425 9.3005
R11821 gnd.n5428 gnd.n5427 9.3005
R11822 gnd.n5426 gnd.n1506 9.3005
R11823 gnd.n5442 gnd.n1505 9.3005
R11824 gnd.n5444 gnd.n5443 9.3005
R11825 gnd.n5445 gnd.n1504 9.3005
R11826 gnd.n5458 gnd.n5446 9.3005
R11827 gnd.n5457 gnd.n5447 9.3005
R11828 gnd.n5456 gnd.n5448 9.3005
R11829 gnd.n5450 gnd.n5449 9.3005
R11830 gnd.n5452 gnd.n5451 9.3005
R11831 gnd.n1471 gnd.n1470 9.3005
R11832 gnd.n5529 gnd.n5528 9.3005
R11833 gnd.n5530 gnd.n1469 9.3005
R11834 gnd.n5532 gnd.n5531 9.3005
R11835 gnd.n1467 gnd.n1466 9.3005
R11836 gnd.n5537 gnd.n5536 9.3005
R11837 gnd.n5538 gnd.n1465 9.3005
R11838 gnd.n5540 gnd.n5539 9.3005
R11839 gnd.n1463 gnd.n1462 9.3005
R11840 gnd.n5545 gnd.n5544 9.3005
R11841 gnd.n5546 gnd.n1461 9.3005
R11842 gnd.n5551 gnd.n5547 9.3005
R11843 gnd.n5550 gnd.n5549 9.3005
R11844 gnd.n5548 gnd.n391 9.3005
R11845 gnd.n6791 gnd.n392 9.3005
R11846 gnd.n6790 gnd.n393 9.3005
R11847 gnd.n6789 gnd.n394 9.3005
R11848 gnd.n4295 gnd.n4294 9.3005
R11849 gnd.n6083 gnd.n880 9.3005
R11850 gnd.n6084 gnd.n879 9.3005
R11851 gnd.n878 gnd.n874 9.3005
R11852 gnd.n6090 gnd.n873 9.3005
R11853 gnd.n6091 gnd.n872 9.3005
R11854 gnd.n6092 gnd.n871 9.3005
R11855 gnd.n870 gnd.n866 9.3005
R11856 gnd.n6098 gnd.n865 9.3005
R11857 gnd.n6099 gnd.n864 9.3005
R11858 gnd.n6100 gnd.n863 9.3005
R11859 gnd.n862 gnd.n858 9.3005
R11860 gnd.n6106 gnd.n857 9.3005
R11861 gnd.n6107 gnd.n856 9.3005
R11862 gnd.n6108 gnd.n855 9.3005
R11863 gnd.n854 gnd.n850 9.3005
R11864 gnd.n6114 gnd.n849 9.3005
R11865 gnd.n6115 gnd.n848 9.3005
R11866 gnd.n6116 gnd.n847 9.3005
R11867 gnd.n846 gnd.n842 9.3005
R11868 gnd.n6122 gnd.n841 9.3005
R11869 gnd.n6123 gnd.n840 9.3005
R11870 gnd.n6124 gnd.n839 9.3005
R11871 gnd.n838 gnd.n834 9.3005
R11872 gnd.n6130 gnd.n833 9.3005
R11873 gnd.n6131 gnd.n832 9.3005
R11874 gnd.n6132 gnd.n831 9.3005
R11875 gnd.n830 gnd.n826 9.3005
R11876 gnd.n6138 gnd.n825 9.3005
R11877 gnd.n6139 gnd.n824 9.3005
R11878 gnd.n6140 gnd.n823 9.3005
R11879 gnd.n822 gnd.n818 9.3005
R11880 gnd.n6146 gnd.n817 9.3005
R11881 gnd.n6147 gnd.n816 9.3005
R11882 gnd.n6148 gnd.n815 9.3005
R11883 gnd.n814 gnd.n810 9.3005
R11884 gnd.n6154 gnd.n809 9.3005
R11885 gnd.n6155 gnd.n808 9.3005
R11886 gnd.n6156 gnd.n807 9.3005
R11887 gnd.n806 gnd.n802 9.3005
R11888 gnd.n6162 gnd.n801 9.3005
R11889 gnd.n6163 gnd.n800 9.3005
R11890 gnd.n6164 gnd.n799 9.3005
R11891 gnd.n798 gnd.n794 9.3005
R11892 gnd.n6170 gnd.n793 9.3005
R11893 gnd.n6171 gnd.n792 9.3005
R11894 gnd.n6172 gnd.n791 9.3005
R11895 gnd.n790 gnd.n786 9.3005
R11896 gnd.n6178 gnd.n785 9.3005
R11897 gnd.n6179 gnd.n784 9.3005
R11898 gnd.n6180 gnd.n783 9.3005
R11899 gnd.n782 gnd.n778 9.3005
R11900 gnd.n6186 gnd.n777 9.3005
R11901 gnd.n6187 gnd.n776 9.3005
R11902 gnd.n6188 gnd.n775 9.3005
R11903 gnd.n774 gnd.n770 9.3005
R11904 gnd.n6194 gnd.n769 9.3005
R11905 gnd.n6195 gnd.n768 9.3005
R11906 gnd.n6196 gnd.n767 9.3005
R11907 gnd.n766 gnd.n762 9.3005
R11908 gnd.n6202 gnd.n761 9.3005
R11909 gnd.n6203 gnd.n760 9.3005
R11910 gnd.n6204 gnd.n759 9.3005
R11911 gnd.n758 gnd.n754 9.3005
R11912 gnd.n6210 gnd.n753 9.3005
R11913 gnd.n6211 gnd.n752 9.3005
R11914 gnd.n6212 gnd.n751 9.3005
R11915 gnd.n750 gnd.n746 9.3005
R11916 gnd.n6218 gnd.n745 9.3005
R11917 gnd.n6219 gnd.n744 9.3005
R11918 gnd.n6220 gnd.n743 9.3005
R11919 gnd.n742 gnd.n738 9.3005
R11920 gnd.n6226 gnd.n737 9.3005
R11921 gnd.n6227 gnd.n736 9.3005
R11922 gnd.n6228 gnd.n735 9.3005
R11923 gnd.n734 gnd.n730 9.3005
R11924 gnd.n6234 gnd.n729 9.3005
R11925 gnd.n6235 gnd.n728 9.3005
R11926 gnd.n6236 gnd.n727 9.3005
R11927 gnd.n726 gnd.n722 9.3005
R11928 gnd.n6242 gnd.n721 9.3005
R11929 gnd.n6243 gnd.n720 9.3005
R11930 gnd.n6244 gnd.n719 9.3005
R11931 gnd.n715 gnd.n714 9.3005
R11932 gnd.n6251 gnd.n6250 9.3005
R11933 gnd.n6082 gnd.n881 9.3005
R11934 gnd.n5463 gnd.n1216 9.3005
R11935 gnd.n4645 gnd.n4644 9.3005
R11936 gnd.n4646 gnd.n2003 9.3005
R11937 gnd.n4665 gnd.n4664 9.3005
R11938 gnd.n4663 gnd.n2004 9.3005
R11939 gnd.n4662 gnd.n4661 9.3005
R11940 gnd.n4660 gnd.n4647 9.3005
R11941 gnd.n4659 gnd.n4658 9.3005
R11942 gnd.n4657 gnd.n4650 9.3005
R11943 gnd.n4656 gnd.n4655 9.3005
R11944 gnd.n4654 gnd.n4651 9.3005
R11945 gnd.n1130 gnd.n1128 9.3005
R11946 gnd.n5889 gnd.n5888 9.3005
R11947 gnd.n5887 gnd.n1129 9.3005
R11948 gnd.n5886 gnd.n5885 9.3005
R11949 gnd.n5884 gnd.n1131 9.3005
R11950 gnd.n5883 gnd.n5882 9.3005
R11951 gnd.n5881 gnd.n1135 9.3005
R11952 gnd.n5880 gnd.n5879 9.3005
R11953 gnd.n5878 gnd.n1136 9.3005
R11954 gnd.n5877 gnd.n5876 9.3005
R11955 gnd.n5875 gnd.n1140 9.3005
R11956 gnd.n5874 gnd.n5873 9.3005
R11957 gnd.n5872 gnd.n1141 9.3005
R11958 gnd.n5871 gnd.n5870 9.3005
R11959 gnd.n5869 gnd.n1145 9.3005
R11960 gnd.n5868 gnd.n5867 9.3005
R11961 gnd.n5866 gnd.n1146 9.3005
R11962 gnd.n5865 gnd.n5864 9.3005
R11963 gnd.n5863 gnd.n1150 9.3005
R11964 gnd.n5862 gnd.n5861 9.3005
R11965 gnd.n5860 gnd.n1151 9.3005
R11966 gnd.n5859 gnd.n5858 9.3005
R11967 gnd.n5857 gnd.n1155 9.3005
R11968 gnd.n5856 gnd.n5855 9.3005
R11969 gnd.n5854 gnd.n1156 9.3005
R11970 gnd.n5853 gnd.n5852 9.3005
R11971 gnd.n5851 gnd.n1160 9.3005
R11972 gnd.n5850 gnd.n5849 9.3005
R11973 gnd.n5848 gnd.n1161 9.3005
R11974 gnd.n5847 gnd.n5846 9.3005
R11975 gnd.n5845 gnd.n1165 9.3005
R11976 gnd.n5844 gnd.n5843 9.3005
R11977 gnd.n5842 gnd.n1166 9.3005
R11978 gnd.n5841 gnd.n5840 9.3005
R11979 gnd.n5839 gnd.n1170 9.3005
R11980 gnd.n5838 gnd.n5837 9.3005
R11981 gnd.n5836 gnd.n1171 9.3005
R11982 gnd.n5835 gnd.n5834 9.3005
R11983 gnd.n5833 gnd.n1175 9.3005
R11984 gnd.n5832 gnd.n5831 9.3005
R11985 gnd.n5830 gnd.n1176 9.3005
R11986 gnd.n5829 gnd.n5828 9.3005
R11987 gnd.n5827 gnd.n1180 9.3005
R11988 gnd.n5826 gnd.n5825 9.3005
R11989 gnd.n5824 gnd.n1181 9.3005
R11990 gnd.n5823 gnd.n5822 9.3005
R11991 gnd.n5821 gnd.n1185 9.3005
R11992 gnd.n5820 gnd.n5819 9.3005
R11993 gnd.n5818 gnd.n1186 9.3005
R11994 gnd.n5817 gnd.n5816 9.3005
R11995 gnd.n5815 gnd.n1190 9.3005
R11996 gnd.n5814 gnd.n5813 9.3005
R11997 gnd.n5812 gnd.n1191 9.3005
R11998 gnd.n5811 gnd.n5810 9.3005
R11999 gnd.n5809 gnd.n1195 9.3005
R12000 gnd.n5808 gnd.n5807 9.3005
R12001 gnd.n5806 gnd.n1196 9.3005
R12002 gnd.n5805 gnd.n5804 9.3005
R12003 gnd.n5803 gnd.n1200 9.3005
R12004 gnd.n5802 gnd.n5801 9.3005
R12005 gnd.n5800 gnd.n1201 9.3005
R12006 gnd.n5799 gnd.n5798 9.3005
R12007 gnd.n5797 gnd.n1205 9.3005
R12008 gnd.n5796 gnd.n5795 9.3005
R12009 gnd.n5794 gnd.n1206 9.3005
R12010 gnd.n5793 gnd.n5792 9.3005
R12011 gnd.n5791 gnd.n1210 9.3005
R12012 gnd.n5790 gnd.n5789 9.3005
R12013 gnd.n5788 gnd.n1211 9.3005
R12014 gnd.n5787 gnd.n5786 9.3005
R12015 gnd.n5785 gnd.n1215 9.3005
R12016 gnd.n5784 gnd.n5783 9.3005
R12017 gnd.n2006 gnd.n2005 9.3005
R12018 gnd.n4631 gnd.n4630 9.3005
R12019 gnd.n4213 gnd.n4212 9.3005
R12020 gnd.n4211 gnd.n2116 9.3005
R12021 gnd.n4210 gnd.n4209 9.3005
R12022 gnd.n4208 gnd.n4199 9.3005
R12023 gnd.n4207 gnd.n4206 9.3005
R12024 gnd.n4205 gnd.n4202 9.3005
R12025 gnd.n4204 gnd.n4203 9.3005
R12026 gnd.n2074 gnd.n2073 9.3005
R12027 gnd.n4266 gnd.n4265 9.3005
R12028 gnd.n4267 gnd.n2072 9.3005
R12029 gnd.n4269 gnd.n4268 9.3005
R12030 gnd.n2069 gnd.n2067 9.3005
R12031 gnd.n4288 gnd.n4287 9.3005
R12032 gnd.n4286 gnd.n2068 9.3005
R12033 gnd.n4285 gnd.n4284 9.3005
R12034 gnd.n2059 gnd.n2058 9.3005
R12035 gnd.n4319 gnd.n4318 9.3005
R12036 gnd.n4320 gnd.n2057 9.3005
R12037 gnd.n4322 gnd.n4321 9.3005
R12038 gnd.n2052 gnd.n2050 9.3005
R12039 gnd.n4594 gnd.n4593 9.3005
R12040 gnd.n4592 gnd.n2051 9.3005
R12041 gnd.n4591 gnd.n4590 9.3005
R12042 gnd.n4589 gnd.n2053 9.3005
R12043 gnd.n4588 gnd.n4587 9.3005
R12044 gnd.n4586 gnd.n4585 9.3005
R12045 gnd.n2037 gnd.n2032 9.3005
R12046 gnd.n4472 gnd.n4471 9.3005
R12047 gnd.n4371 gnd.n4370 9.3005
R12048 gnd.n4466 gnd.n4465 9.3005
R12049 gnd.n4464 gnd.n4463 9.3005
R12050 gnd.n4383 gnd.n4382 9.3005
R12051 gnd.n4458 gnd.n4457 9.3005
R12052 gnd.n4456 gnd.n4455 9.3005
R12053 gnd.n4391 gnd.n4390 9.3005
R12054 gnd.n4450 gnd.n4449 9.3005
R12055 gnd.n4448 gnd.n4447 9.3005
R12056 gnd.n4403 gnd.n4402 9.3005
R12057 gnd.n4442 gnd.n4441 9.3005
R12058 gnd.n4440 gnd.n4439 9.3005
R12059 gnd.n4411 gnd.n4410 9.3005
R12060 gnd.n4434 gnd.n4433 9.3005
R12061 gnd.n4432 gnd.n4431 9.3005
R12062 gnd.n4422 gnd.n2036 9.3005
R12063 gnd.n4627 gnd.n4626 9.3005
R12064 gnd.n4474 gnd.n4473 9.3005
R12065 gnd.n4628 gnd.n2031 9.3005
R12066 gnd.n4428 gnd.n2033 9.3005
R12067 gnd.n4430 gnd.n4429 9.3005
R12068 gnd.n4417 gnd.n4416 9.3005
R12069 gnd.n4436 gnd.n4435 9.3005
R12070 gnd.n4438 gnd.n4437 9.3005
R12071 gnd.n4407 gnd.n4406 9.3005
R12072 gnd.n4444 gnd.n4443 9.3005
R12073 gnd.n4446 gnd.n4445 9.3005
R12074 gnd.n4397 gnd.n4396 9.3005
R12075 gnd.n4452 gnd.n4451 9.3005
R12076 gnd.n4454 gnd.n4453 9.3005
R12077 gnd.n4387 gnd.n4386 9.3005
R12078 gnd.n4460 gnd.n4459 9.3005
R12079 gnd.n4462 gnd.n4461 9.3005
R12080 gnd.n4377 gnd.n4376 9.3005
R12081 gnd.n4468 gnd.n4467 9.3005
R12082 gnd.n4470 gnd.n4469 9.3005
R12083 gnd.n4368 gnd.n4367 9.3005
R12084 gnd.n4476 gnd.n4475 9.3005
R12085 gnd.n4477 gnd.n4335 9.3005
R12086 gnd.n4479 gnd.n4478 9.3005
R12087 gnd.n4362 gnd.n4336 9.3005
R12088 gnd.n4361 gnd.n4360 9.3005
R12089 gnd.n4359 gnd.n4337 9.3005
R12090 gnd.n4358 gnd.n4357 9.3005
R12091 gnd.n4354 gnd.n4340 9.3005
R12092 gnd.n4353 gnd.n4341 9.3005
R12093 gnd.n4348 gnd.n4342 9.3005
R12094 gnd.n4347 gnd.n4346 9.3005
R12095 gnd.n4345 gnd.n4343 9.3005
R12096 gnd.n1988 gnd.n1987 9.3005
R12097 gnd.n4687 gnd.n4686 9.3005
R12098 gnd.n4688 gnd.n1986 9.3005
R12099 gnd.n4690 gnd.n4689 9.3005
R12100 gnd.n1984 gnd.n1983 9.3005
R12101 gnd.n4695 gnd.n4694 9.3005
R12102 gnd.n4696 gnd.n1981 9.3005
R12103 gnd.n4839 gnd.n4838 9.3005
R12104 gnd.n4837 gnd.n1982 9.3005
R12105 gnd.n4836 gnd.n4835 9.3005
R12106 gnd.n4834 gnd.n4697 9.3005
R12107 gnd.n4833 gnd.n4832 9.3005
R12108 gnd.n4831 gnd.n4699 9.3005
R12109 gnd.n4830 gnd.n4829 9.3005
R12110 gnd.n4828 gnd.n4700 9.3005
R12111 gnd.n4827 gnd.n4826 9.3005
R12112 gnd.n4825 gnd.n4702 9.3005
R12113 gnd.n4824 gnd.n4823 9.3005
R12114 gnd.n4822 gnd.n4703 9.3005
R12115 gnd.n4821 gnd.n4820 9.3005
R12116 gnd.n4819 gnd.n4708 9.3005
R12117 gnd.n4818 gnd.n4817 9.3005
R12118 gnd.n4816 gnd.n4709 9.3005
R12119 gnd.n4815 gnd.n4814 9.3005
R12120 gnd.n4813 gnd.n4712 9.3005
R12121 gnd.n4812 gnd.n4811 9.3005
R12122 gnd.n4810 gnd.n4713 9.3005
R12123 gnd.n4809 gnd.n4808 9.3005
R12124 gnd.n4807 gnd.n4716 9.3005
R12125 gnd.n4806 gnd.n4805 9.3005
R12126 gnd.n4804 gnd.n4717 9.3005
R12127 gnd.n4803 gnd.n4802 9.3005
R12128 gnd.n4801 gnd.n4719 9.3005
R12129 gnd.n4800 gnd.n4799 9.3005
R12130 gnd.n4798 gnd.n4720 9.3005
R12131 gnd.n4797 gnd.n4796 9.3005
R12132 gnd.n4795 gnd.n4725 9.3005
R12133 gnd.n4794 gnd.n4793 9.3005
R12134 gnd.n4792 gnd.n4726 9.3005
R12135 gnd.n4791 gnd.n4790 9.3005
R12136 gnd.n4789 gnd.n4728 9.3005
R12137 gnd.n4788 gnd.n4787 9.3005
R12138 gnd.n4786 gnd.n4729 9.3005
R12139 gnd.n4785 gnd.n4784 9.3005
R12140 gnd.n4783 gnd.n4732 9.3005
R12141 gnd.n4782 gnd.n4781 9.3005
R12142 gnd.n4780 gnd.n4733 9.3005
R12143 gnd.n4779 gnd.n4778 9.3005
R12144 gnd.n4777 gnd.n4737 9.3005
R12145 gnd.n4776 gnd.n4775 9.3005
R12146 gnd.n4774 gnd.n4738 9.3005
R12147 gnd.n4773 gnd.n4772 9.3005
R12148 gnd.n4771 gnd.n4741 9.3005
R12149 gnd.n4770 gnd.n4769 9.3005
R12150 gnd.n4768 gnd.n4742 9.3005
R12151 gnd.n4767 gnd.n4766 9.3005
R12152 gnd.n4765 gnd.n4746 9.3005
R12153 gnd.n4764 gnd.n4763 9.3005
R12154 gnd.n4762 gnd.n4747 9.3005
R12155 gnd.n4761 gnd.n4760 9.3005
R12156 gnd.n4759 gnd.n4751 9.3005
R12157 gnd.n4758 gnd.n4757 9.3005
R12158 gnd.n4756 gnd.n4752 9.3005
R12159 gnd.n4755 gnd.n4754 9.3005
R12160 gnd.n1623 gnd.n1622 9.3005
R12161 gnd.n5267 gnd.n5266 9.3005
R12162 gnd.n5268 gnd.n1620 9.3005
R12163 gnd.n5271 gnd.n5270 9.3005
R12164 gnd.n5269 gnd.n1621 9.3005
R12165 gnd.n1524 gnd.n1523 9.3005
R12166 gnd.n5415 gnd.n5414 9.3005
R12167 gnd.n5416 gnd.n1522 9.3005
R12168 gnd.n5418 gnd.n5417 9.3005
R12169 gnd.n1512 gnd.n1511 9.3005
R12170 gnd.n5434 gnd.n5433 9.3005
R12171 gnd.n5435 gnd.n1510 9.3005
R12172 gnd.n5437 gnd.n5436 9.3005
R12173 gnd.n1225 gnd.n1224 9.3005
R12174 gnd.n5779 gnd.n5778 9.3005
R12175 gnd.n4350 gnd.n4349 9.3005
R12176 gnd.n5775 gnd.n1226 9.3005
R12177 gnd.n5774 gnd.n5773 9.3005
R12178 gnd.n5772 gnd.n1229 9.3005
R12179 gnd.n5771 gnd.n5770 9.3005
R12180 gnd.n5769 gnd.n1230 9.3005
R12181 gnd.n5768 gnd.n5767 9.3005
R12182 gnd.n5777 gnd.n5776 9.3005
R12183 gnd.n5720 gnd.n5719 9.3005
R12184 gnd.n1277 gnd.n1276 9.3005
R12185 gnd.n5726 gnd.n5725 9.3005
R12186 gnd.n5728 gnd.n5727 9.3005
R12187 gnd.n1269 gnd.n1268 9.3005
R12188 gnd.n5734 gnd.n5733 9.3005
R12189 gnd.n5736 gnd.n5735 9.3005
R12190 gnd.n1261 gnd.n1260 9.3005
R12191 gnd.n5742 gnd.n5741 9.3005
R12192 gnd.n5744 gnd.n5743 9.3005
R12193 gnd.n1253 gnd.n1252 9.3005
R12194 gnd.n5750 gnd.n5749 9.3005
R12195 gnd.n5752 gnd.n5751 9.3005
R12196 gnd.n1245 gnd.n1244 9.3005
R12197 gnd.n5758 gnd.n5757 9.3005
R12198 gnd.n5760 gnd.n5759 9.3005
R12199 gnd.n1241 gnd.n1236 9.3005
R12200 gnd.n5718 gnd.n1286 9.3005
R12201 gnd.n1475 gnd.n1285 9.3005
R12202 gnd.n5765 gnd.n1234 9.3005
R12203 gnd.n5764 gnd.n5763 9.3005
R12204 gnd.n5762 gnd.n5761 9.3005
R12205 gnd.n1240 gnd.n1239 9.3005
R12206 gnd.n5756 gnd.n5755 9.3005
R12207 gnd.n5754 gnd.n5753 9.3005
R12208 gnd.n1249 gnd.n1248 9.3005
R12209 gnd.n5748 gnd.n5747 9.3005
R12210 gnd.n5746 gnd.n5745 9.3005
R12211 gnd.n1257 gnd.n1256 9.3005
R12212 gnd.n5740 gnd.n5739 9.3005
R12213 gnd.n5738 gnd.n5737 9.3005
R12214 gnd.n1265 gnd.n1264 9.3005
R12215 gnd.n5732 gnd.n5731 9.3005
R12216 gnd.n5730 gnd.n5729 9.3005
R12217 gnd.n1273 gnd.n1272 9.3005
R12218 gnd.n5724 gnd.n5723 9.3005
R12219 gnd.n5722 gnd.n5721 9.3005
R12220 gnd.n1498 gnd.n1283 9.3005
R12221 gnd.n1477 gnd.n1476 9.3005
R12222 gnd.n5465 gnd.n5464 9.3005
R12223 gnd.n5523 gnd.n5522 9.3005
R12224 gnd.n5521 gnd.n1474 9.3005
R12225 gnd.n5520 gnd.n5519 9.3005
R12226 gnd.n5518 gnd.n5468 9.3005
R12227 gnd.n5517 gnd.n5516 9.3005
R12228 gnd.n5515 gnd.n5471 9.3005
R12229 gnd.n5514 gnd.n5513 9.3005
R12230 gnd.n5512 gnd.n5472 9.3005
R12231 gnd.n5511 gnd.n5510 9.3005
R12232 gnd.n5509 gnd.n5475 9.3005
R12233 gnd.n5508 gnd.n5507 9.3005
R12234 gnd.n5506 gnd.n5476 9.3005
R12235 gnd.n5505 gnd.n5504 9.3005
R12236 gnd.n368 gnd.n367 9.3005
R12237 gnd.n6820 gnd.n6819 9.3005
R12238 gnd.n6821 gnd.n365 9.3005
R12239 gnd.n6824 gnd.n6823 9.3005
R12240 gnd.n6822 gnd.n366 9.3005
R12241 gnd.n341 gnd.n340 9.3005
R12242 gnd.n6854 gnd.n6853 9.3005
R12243 gnd.n6855 gnd.n338 9.3005
R12244 gnd.n6863 gnd.n6862 9.3005
R12245 gnd.n6861 gnd.n339 9.3005
R12246 gnd.n6860 gnd.n6859 9.3005
R12247 gnd.n6858 gnd.n6856 9.3005
R12248 gnd.n81 gnd.n79 9.3005
R12249 gnd.n5467 gnd.n1473 9.3005
R12250 gnd.t182 gnd.n2435 9.24152
R12251 gnd.n2337 gnd.t54 9.24152
R12252 gnd.n3621 gnd.t170 9.24152
R12253 gnd.t66 gnd.n2226 9.24152
R12254 gnd.n4583 gnd.t91 9.24152
R12255 gnd.n5586 gnd.t62 9.24152
R12256 gnd.t74 gnd.n195 9.24152
R12257 gnd.t190 gnd.t182 8.92286
R12258 gnd.n4924 gnd.n1869 8.92286
R12259 gnd.n4959 gnd.n4958 8.92286
R12260 gnd.n5048 gnd.n1788 8.92286
R12261 gnd.n5082 gnd.n5081 8.92286
R12262 gnd.n5166 gnd.n1706 8.92286
R12263 gnd.n5199 gnd.n1677 8.92286
R12264 gnd.n5404 gnd.n5403 8.92286
R12265 gnd.n3591 gnd.n3566 8.92171
R12266 gnd.n3559 gnd.n3534 8.92171
R12267 gnd.n3527 gnd.n3502 8.92171
R12268 gnd.n3496 gnd.n3471 8.92171
R12269 gnd.n3464 gnd.n3439 8.92171
R12270 gnd.n3432 gnd.n3407 8.92171
R12271 gnd.n3400 gnd.n3375 8.92171
R12272 gnd.n3369 gnd.n3344 8.92171
R12273 gnd.n1560 gnd.n1542 8.72777
R12274 gnd.n3095 gnd.t194 8.60421
R12275 gnd.t360 gnd.n5047 8.60421
R12276 gnd.n5059 gnd.t22 8.60421
R12277 gnd.n2507 gnd.n2491 8.43656
R12278 gnd.n46 gnd.n30 8.43656
R12279 gnd.n4849 gnd.t105 8.28555
R12280 gnd.n3592 gnd.n3564 8.14595
R12281 gnd.n3560 gnd.n3532 8.14595
R12282 gnd.n3528 gnd.n3500 8.14595
R12283 gnd.n3497 gnd.n3469 8.14595
R12284 gnd.n3465 gnd.n3437 8.14595
R12285 gnd.n3433 gnd.n3405 8.14595
R12286 gnd.n3401 gnd.n3373 8.14595
R12287 gnd.n3370 gnd.n3342 8.14595
R12288 gnd.n4198 gnd.n0 8.10675
R12289 gnd.n7269 gnd.n7268 8.10675
R12290 gnd.n3597 gnd.n3596 7.97301
R12291 gnd.t181 gnd.n2610 7.9669
R12292 gnd.n4884 gnd.t358 7.9669
R12293 gnd.n5232 gnd.t15 7.9669
R12294 gnd.n7269 gnd.n78 7.86902
R12295 gnd.n5718 gnd.n1285 7.75808
R12296 gnd.n7022 gnd.n6969 7.75808
R12297 gnd.n4626 gnd.n2036 7.75808
R12298 gnd.n3879 gnd.n3843 7.75808
R12299 gnd.t5 gnd.n1873 7.64824
R12300 gnd.n5005 gnd.t17 7.64824
R12301 gnd.n5015 gnd.t17 7.64824
R12302 gnd.n5108 gnd.t34 7.64824
R12303 gnd.n5116 gnd.t34 7.64824
R12304 gnd.t189 gnd.n1663 7.64824
R12305 gnd.n2540 gnd.n2539 7.53171
R12306 gnd.n3004 gnd.t7 7.32958
R12307 gnd.n1106 gnd.n1105 7.30353
R12308 gnd.n1559 gnd.n1558 7.30353
R12309 gnd.n2964 gnd.n2683 7.01093
R12310 gnd.n2686 gnd.n2684 7.01093
R12311 gnd.n2974 gnd.n2973 7.01093
R12312 gnd.n2985 gnd.n2667 7.01093
R12313 gnd.n2984 gnd.n2670 7.01093
R12314 gnd.n2995 gnd.n2658 7.01093
R12315 gnd.n2661 gnd.n2659 7.01093
R12316 gnd.n3005 gnd.n3004 7.01093
R12317 gnd.n3015 gnd.n2639 7.01093
R12318 gnd.n3014 gnd.n2642 7.01093
R12319 gnd.n3023 gnd.n2633 7.01093
R12320 gnd.n3035 gnd.n2623 7.01093
R12321 gnd.n3045 gnd.n2608 7.01093
R12322 gnd.n3061 gnd.n3060 7.01093
R12323 gnd.n2610 gnd.n2547 7.01093
R12324 gnd.n3115 gnd.n2548 7.01093
R12325 gnd.n3109 gnd.n3108 7.01093
R12326 gnd.n2597 gnd.n2559 7.01093
R12327 gnd.n3101 gnd.n2570 7.01093
R12328 gnd.n2588 gnd.n2583 7.01093
R12329 gnd.n3095 gnd.n3094 7.01093
R12330 gnd.n3141 gnd.n2470 7.01093
R12331 gnd.n3140 gnd.n3139 7.01093
R12332 gnd.n3152 gnd.n3151 7.01093
R12333 gnd.n2463 gnd.n2455 7.01093
R12334 gnd.n3181 gnd.n2443 7.01093
R12335 gnd.n3180 gnd.n2446 7.01093
R12336 gnd.n3191 gnd.n2435 7.01093
R12337 gnd.n2436 gnd.n2424 7.01093
R12338 gnd.n3202 gnd.n2425 7.01093
R12339 gnd.n3226 gnd.n2416 7.01093
R12340 gnd.n3225 gnd.n2407 7.01093
R12341 gnd.n3248 gnd.n3247 7.01093
R12342 gnd.n3266 gnd.n2388 7.01093
R12343 gnd.n3265 gnd.n2391 7.01093
R12344 gnd.n3276 gnd.n2380 7.01093
R12345 gnd.n2381 gnd.n2368 7.01093
R12346 gnd.n3287 gnd.n2369 7.01093
R12347 gnd.n3314 gnd.n2353 7.01093
R12348 gnd.n3326 gnd.n3325 7.01093
R12349 gnd.n3308 gnd.n2346 7.01093
R12350 gnd.n3337 gnd.n3336 7.01093
R12351 gnd.n3609 gnd.n2334 7.01093
R12352 gnd.n3608 gnd.n2337 7.01093
R12353 gnd.n3621 gnd.n2326 7.01093
R12354 gnd.n2327 gnd.n2318 7.01093
R12355 gnd.n3631 gnd.n2319 7.01093
R12356 gnd.n5034 gnd.t192 7.01093
R12357 gnd.n5098 gnd.t186 7.01093
R12358 gnd.n2642 gnd.t20 6.69227
R12359 gnd.n2446 gnd.t190 6.69227
R12360 gnd.n3315 gnd.t195 6.69227
R12361 gnd.n4089 gnd.t198 6.69227
R12362 gnd.n6055 gnd.t234 6.69227
R12363 gnd.n4597 gnd.t221 6.69227
R12364 gnd.n1875 gnd.t50 6.69227
R12365 gnd.t0 gnd.n1670 6.69227
R12366 gnd.t228 gnd.n1435 6.69227
R12367 gnd.n5493 gnd.t200 6.69227
R12368 gnd.n7215 gnd.t215 6.69227
R12369 gnd.n5333 gnd.n5332 6.5566
R12370 gnd.n1914 gnd.n1913 6.5566
R12371 gnd.n5910 gnd.n5906 6.5566
R12372 gnd.n5345 gnd.n1587 6.5566
R12373 gnd.n4863 gnd.n1899 6.37362
R12374 gnd.n4892 gnd.n4890 6.37362
R12375 gnd.n4987 gnd.n4986 6.37362
R12376 gnd.n5136 gnd.n5135 6.37362
R12377 gnd.n5226 gnd.n5225 6.37362
R12378 gnd.n5238 gnd.n1637 6.37362
R12379 gnd.n4429 gnd.n4425 6.20656
R12380 gnd.n1498 gnd.n1282 6.20656
R12381 gnd.t39 gnd.n3071 6.05496
R12382 gnd.n3072 gnd.t21 6.05496
R12383 gnd.t41 gnd.n2470 6.05496
R12384 gnd.t188 gnd.n3236 6.05496
R12385 gnd.n4133 gnd.t213 6.05496
R12386 gnd.t226 gnd.n6079 6.05496
R12387 gnd.n4291 gnd.t211 6.05496
R12388 gnd.n5969 gnd.n1052 6.05496
R12389 gnd.n6793 gnd.t237 6.05496
R12390 gnd.n6826 gnd.t202 6.05496
R12391 gnd.n7239 gnd.t258 6.05496
R12392 gnd.n3594 gnd.n3564 5.81868
R12393 gnd.n3562 gnd.n3532 5.81868
R12394 gnd.n3530 gnd.n3500 5.81868
R12395 gnd.n3499 gnd.n3469 5.81868
R12396 gnd.n3467 gnd.n3437 5.81868
R12397 gnd.n3435 gnd.n3405 5.81868
R12398 gnd.n3403 gnd.n3373 5.81868
R12399 gnd.n3372 gnd.n3342 5.81868
R12400 gnd.t78 gnd.n1084 5.73631
R12401 gnd.n1973 gnd.t78 5.73631
R12402 gnd.n4871 gnd.t88 5.73631
R12403 gnd.n4924 gnd.t357 5.73631
R12404 gnd.n4994 gnd.t356 5.73631
R12405 gnd.n5127 gnd.t178 5.73631
R12406 gnd.n5199 gnd.t173 5.73631
R12407 gnd.n1589 gnd.n1362 5.62001
R12408 gnd.n5972 gnd.n1048 5.62001
R12409 gnd.n5972 gnd.n1049 5.62001
R12410 gnd.n5343 gnd.n1362 5.62001
R12411 gnd.n2823 gnd.n2818 5.4308
R12412 gnd.n3639 gnd.n2311 5.4308
R12413 gnd.n3139 gnd.t45 5.41765
R12414 gnd.t187 gnd.n3162 5.41765
R12415 gnd.t35 gnd.n2400 5.41765
R12416 gnd.n4193 gnd.t275 5.41765
R12417 gnd.n4226 gnd.t231 5.41765
R12418 gnd.n4950 gnd.t48 5.41765
R12419 gnd.n1701 gnd.t24 5.41765
R12420 gnd.n6885 gnd.t204 5.41765
R12421 gnd.n7263 gnd.t240 5.41765
R12422 gnd.t133 gnd.n5897 5.09899
R12423 gnd.n4872 gnd.n4871 5.09899
R12424 gnd.n4884 gnd.n4883 5.09899
R12425 gnd.n4976 gnd.t46 5.09899
R12426 gnd.n1819 gnd.n1814 5.09899
R12427 gnd.n5008 gnd.n5007 5.09899
R12428 gnd.n1737 gnd.n1731 5.09899
R12429 gnd.n5129 gnd.n5128 5.09899
R12430 gnd.n5152 gnd.t33 5.09899
R12431 gnd.n5232 gnd.n1649 5.09899
R12432 gnd.n5254 gnd.n1634 5.09899
R12433 gnd.n3592 gnd.n3591 5.04292
R12434 gnd.n3560 gnd.n3559 5.04292
R12435 gnd.n3528 gnd.n3527 5.04292
R12436 gnd.n3497 gnd.n3496 5.04292
R12437 gnd.n3465 gnd.n3464 5.04292
R12438 gnd.n3433 gnd.n3432 5.04292
R12439 gnd.n3401 gnd.n3400 5.04292
R12440 gnd.n3370 gnd.n3369 5.04292
R12441 gnd.n3102 gnd.t6 4.78034
R12442 gnd.n2425 gnd.t184 4.78034
R12443 gnd.n4158 gnd.t260 4.78034
R12444 gnd.n2086 gnd.t277 4.78034
R12445 gnd.n1857 gnd.t48 4.78034
R12446 gnd.t24 gnd.n1691 4.78034
R12447 gnd.n1528 gnd.t149 4.78034
R12448 gnd.n6851 gnd.t245 4.78034
R12449 gnd.t206 gnd.n109 4.78034
R12450 gnd.n2544 gnd.n2541 4.74817
R12451 gnd.n2594 gnd.n2476 4.74817
R12452 gnd.n2581 gnd.n2475 4.74817
R12453 gnd.n2474 gnd.n2473 4.74817
R12454 gnd.n2590 gnd.n2541 4.74817
R12455 gnd.n2591 gnd.n2476 4.74817
R12456 gnd.n2593 gnd.n2475 4.74817
R12457 gnd.n2580 gnd.n2474 4.74817
R12458 gnd.n2539 gnd.n2538 4.74296
R12459 gnd.n78 gnd.n77 4.74296
R12460 gnd.n2507 gnd.n2506 4.7074
R12461 gnd.n2523 gnd.n2522 4.7074
R12462 gnd.n46 gnd.n45 4.7074
R12463 gnd.n62 gnd.n61 4.7074
R12464 gnd.n2539 gnd.n2523 4.65959
R12465 gnd.n78 gnd.n62 4.65959
R12466 gnd.n5660 gnd.n1364 4.6132
R12467 gnd.n5973 gnd.n1047 4.6132
R12468 gnd.n6023 gnd.n978 4.46168
R12469 gnd.n4849 gnd.t70 4.46168
R12470 gnd.n5245 gnd.t111 4.46168
R12471 gnd.n5713 gnd.n1330 4.46168
R12472 gnd.n1555 gnd.n1542 4.46111
R12473 gnd.n3577 gnd.n3573 4.38594
R12474 gnd.n3545 gnd.n3541 4.38594
R12475 gnd.n3513 gnd.n3509 4.38594
R12476 gnd.n3482 gnd.n3478 4.38594
R12477 gnd.n3450 gnd.n3446 4.38594
R12478 gnd.n3418 gnd.n3414 4.38594
R12479 gnd.n3386 gnd.n3382 4.38594
R12480 gnd.n3355 gnd.n3351 4.38594
R12481 gnd.n3588 gnd.n3566 4.26717
R12482 gnd.n3556 gnd.n3534 4.26717
R12483 gnd.n3524 gnd.n3502 4.26717
R12484 gnd.n3493 gnd.n3471 4.26717
R12485 gnd.n3461 gnd.n3439 4.26717
R12486 gnd.n3429 gnd.n3407 4.26717
R12487 gnd.n3397 gnd.n3375 4.26717
R12488 gnd.n3366 gnd.n3344 4.26717
R12489 gnd.n3046 gnd.t183 4.14303
R12490 gnd.n3276 gnd.t19 4.14303
R12491 gnd.t282 gnd.n2178 4.14303
R12492 gnd.n6080 gnd.n883 4.14303
R12493 gnd.n4282 gnd.t251 4.14303
R12494 gnd.n4315 gnd.t234 4.14303
R12495 gnd.t2 gnd.n5014 4.14303
R12496 gnd.n5109 gnd.t176 4.14303
R12497 gnd.t200 gnd.n1453 4.14303
R12498 gnd.n5502 gnd.t217 4.14303
R12499 gnd.n6841 gnd.n351 4.14303
R12500 gnd.t248 gnd.n147 4.14303
R12501 gnd.n3596 gnd.n3595 4.08274
R12502 gnd.n5332 gnd.n5331 4.05904
R12503 gnd.n1915 gnd.n1914 4.05904
R12504 gnd.n5913 gnd.n5906 4.05904
R12505 gnd.n1587 gnd.n1582 4.05904
R12506 gnd.n15 gnd.n7 3.99943
R12507 gnd.n5898 gnd.t133 3.82437
R12508 gnd.n4856 gnd.n1904 3.82437
R12509 gnd.n1890 gnd.n1879 3.82437
R12510 gnd.n4988 gnd.n1823 3.82437
R12511 gnd.n1810 gnd.n1799 3.82437
R12512 gnd.n5110 gnd.n1741 3.82437
R12513 gnd.n4735 gnd.n1727 3.82437
R12514 gnd.n1666 gnd.n1653 3.82437
R12515 gnd.n5238 gnd.t124 3.82437
R12516 gnd.n5264 gnd.n1625 3.82437
R12517 gnd.n3119 gnd.n2540 3.81325
R12518 gnd.n2523 gnd.n2507 3.72967
R12519 gnd.n62 gnd.n46 3.72967
R12520 gnd.n3596 gnd.n3468 3.70378
R12521 gnd.n15 gnd.n14 3.60163
R12522 gnd.n3587 gnd.n3568 3.49141
R12523 gnd.n3555 gnd.n3536 3.49141
R12524 gnd.n3523 gnd.n3504 3.49141
R12525 gnd.n3492 gnd.n3473 3.49141
R12526 gnd.n3460 gnd.n3441 3.49141
R12527 gnd.n3428 gnd.n3409 3.49141
R12528 gnd.n3396 gnd.n3377 3.49141
R12529 gnd.n3365 gnd.n3346 3.49141
R12530 gnd.n7150 gnd.n7147 3.29747
R12531 gnd.n7151 gnd.n7150 3.29747
R12532 gnd.n5678 gnd.n5677 3.29747
R12533 gnd.n5677 gnd.n5676 3.29747
R12534 gnd.n4001 gnd.n4000 3.29747
R12535 gnd.n4000 gnd.n3999 3.29747
R12536 gnd.n5991 gnd.n5990 3.29747
R12537 gnd.n5990 gnd.n5989 3.29747
R12538 gnd.n5891 gnd.t70 3.18706
R12539 gnd.t111 gnd.n1645 3.18706
R12540 gnd.n2625 gnd.t183 2.8684
R12541 gnd.n2524 gnd.t252 2.82907
R12542 gnd.n2524 gnd.t335 2.82907
R12543 gnd.n2526 gnd.t227 2.82907
R12544 gnd.n2526 gnd.t272 2.82907
R12545 gnd.n2528 gnd.t291 2.82907
R12546 gnd.n2528 gnd.t278 2.82907
R12547 gnd.n2530 gnd.t276 2.82907
R12548 gnd.n2530 gnd.t264 2.82907
R12549 gnd.n2532 gnd.t284 2.82907
R12550 gnd.n2532 gnd.t319 2.82907
R12551 gnd.n2534 gnd.t210 2.82907
R12552 gnd.n2534 gnd.t306 2.82907
R12553 gnd.n2536 gnd.t345 2.82907
R12554 gnd.n2536 gnd.t283 2.82907
R12555 gnd.n2477 gnd.t285 2.82907
R12556 gnd.n2477 gnd.t309 2.82907
R12557 gnd.n2479 gnd.t318 2.82907
R12558 gnd.n2479 gnd.t253 2.82907
R12559 gnd.n2481 gnd.t303 2.82907
R12560 gnd.n2481 gnd.t296 2.82907
R12561 gnd.n2483 gnd.t351 2.82907
R12562 gnd.n2483 gnd.t337 2.82907
R12563 gnd.n2485 gnd.t261 2.82907
R12564 gnd.n2485 gnd.t311 2.82907
R12565 gnd.n2487 gnd.t331 2.82907
R12566 gnd.n2487 gnd.t214 2.82907
R12567 gnd.n2489 gnd.t199 2.82907
R12568 gnd.n2489 gnd.t302 2.82907
R12569 gnd.n2492 gnd.t353 2.82907
R12570 gnd.n2492 gnd.t235 2.82907
R12571 gnd.n2494 gnd.t233 2.82907
R12572 gnd.n2494 gnd.t212 2.82907
R12573 gnd.n2496 gnd.t317 2.82907
R12574 gnd.n2496 gnd.t350 2.82907
R12575 gnd.n2498 gnd.t349 2.82907
R12576 gnd.n2498 gnd.t232 2.82907
R12577 gnd.n2500 gnd.t338 2.82907
R12578 gnd.n2500 gnd.t314 2.82907
R12579 gnd.n2502 gnd.t315 2.82907
R12580 gnd.n2502 gnd.t347 2.82907
R12581 gnd.n2504 gnd.t348 2.82907
R12582 gnd.n2504 gnd.t330 2.82907
R12583 gnd.n2508 gnd.t297 2.82907
R12584 gnd.n2508 gnd.t255 2.82907
R12585 gnd.n2510 gnd.t281 2.82907
R12586 gnd.n2510 gnd.t320 2.82907
R12587 gnd.n2512 gnd.t344 2.82907
R12588 gnd.n2512 gnd.t327 2.82907
R12589 gnd.n2514 gnd.t328 2.82907
R12590 gnd.n2514 gnd.t310 2.82907
R12591 gnd.n2516 gnd.t334 2.82907
R12592 gnd.n2516 gnd.t243 2.82907
R12593 gnd.n2518 gnd.t271 2.82907
R12594 gnd.n2518 gnd.t220 2.82907
R12595 gnd.n2520 gnd.t263 2.82907
R12596 gnd.n2520 gnd.t333 2.82907
R12597 gnd.n75 gnd.t249 2.82907
R12598 gnd.n75 gnd.t301 2.82907
R12599 gnd.n73 gnd.t270 2.82907
R12600 gnd.n73 gnd.t312 2.82907
R12601 gnd.n71 gnd.t287 2.82907
R12602 gnd.n71 gnd.t262 2.82907
R12603 gnd.n69 gnd.t219 2.82907
R12604 gnd.n69 gnd.t241 2.82907
R12605 gnd.n67 gnd.t246 2.82907
R12606 gnd.n67 gnd.t267 2.82907
R12607 gnd.n65 gnd.t238 2.82907
R12608 gnd.n65 gnd.t326 2.82907
R12609 gnd.n63 gnd.t298 2.82907
R12610 gnd.n63 gnd.t218 2.82907
R12611 gnd.n28 gnd.t340 2.82907
R12612 gnd.n28 gnd.t265 2.82907
R12613 gnd.n26 gnd.t259 2.82907
R12614 gnd.n26 gnd.t224 2.82907
R12615 gnd.n24 gnd.t355 2.82907
R12616 gnd.n24 gnd.t250 2.82907
R12617 gnd.n22 gnd.t230 2.82907
R12618 gnd.n22 gnd.t247 2.82907
R12619 gnd.n20 gnd.t329 2.82907
R12620 gnd.n20 gnd.t293 2.82907
R12621 gnd.n18 gnd.t280 2.82907
R12622 gnd.n18 gnd.t208 2.82907
R12623 gnd.n16 gnd.t343 2.82907
R12624 gnd.n16 gnd.t269 2.82907
R12625 gnd.n43 gnd.t308 2.82907
R12626 gnd.n43 gnd.t325 2.82907
R12627 gnd.n41 gnd.t324 2.82907
R12628 gnd.n41 gnd.t304 2.82907
R12629 gnd.n39 gnd.t299 2.82907
R12630 gnd.n39 gnd.t207 2.82907
R12631 gnd.n37 gnd.t205 2.82907
R12632 gnd.n37 gnd.t322 2.82907
R12633 gnd.n35 gnd.t332 2.82907
R12634 gnd.n35 gnd.t342 2.82907
R12635 gnd.n33 gnd.t341 2.82907
R12636 gnd.n33 gnd.t203 2.82907
R12637 gnd.n31 gnd.t201 2.82907
R12638 gnd.n31 gnd.t225 2.82907
R12639 gnd.n59 gnd.t295 2.82907
R12640 gnd.n59 gnd.t216 2.82907
R12641 gnd.n57 gnd.t321 2.82907
R12642 gnd.n57 gnd.t236 2.82907
R12643 gnd.n55 gnd.t339 2.82907
R12644 gnd.n55 gnd.t307 2.82907
R12645 gnd.n53 gnd.t279 2.82907
R12646 gnd.n53 gnd.t292 2.82907
R12647 gnd.n51 gnd.t294 2.82907
R12648 gnd.n51 gnd.t313 2.82907
R12649 gnd.n49 gnd.t288 2.82907
R12650 gnd.n49 gnd.t254 2.82907
R12651 gnd.n47 gnd.t354 2.82907
R12652 gnd.n47 gnd.t273 2.82907
R12653 gnd.n3584 gnd.n3583 2.71565
R12654 gnd.n3552 gnd.n3551 2.71565
R12655 gnd.n3520 gnd.n3519 2.71565
R12656 gnd.n3489 gnd.n3488 2.71565
R12657 gnd.n3457 gnd.n3456 2.71565
R12658 gnd.n3425 gnd.n3424 2.71565
R12659 gnd.n3393 gnd.n3392 2.71565
R12660 gnd.n3362 gnd.n3361 2.71565
R12661 gnd.n4842 gnd.n4841 2.54975
R12662 gnd.n4917 gnd.n1875 2.54975
R12663 gnd.n4942 gnd.t4 2.54975
R12664 gnd.n4966 gnd.n1836 2.54975
R12665 gnd.n1837 gnd.t46 2.54975
R12666 gnd.n5041 gnd.n1795 2.54975
R12667 gnd.n5089 gnd.n1755 2.54975
R12668 gnd.t33 gnd.n1710 2.54975
R12669 gnd.n5159 gnd.n1712 2.54975
R12670 gnd.n5182 gnd.t52 2.54975
R12671 gnd.n5211 gnd.n1670 2.54975
R12672 gnd.n5273 gnd.n1618 2.54975
R12673 gnd.n3119 gnd.n2541 2.27742
R12674 gnd.n3119 gnd.n2476 2.27742
R12675 gnd.n3119 gnd.n2475 2.27742
R12676 gnd.n3119 gnd.n2474 2.27742
R12677 gnd.n2973 gnd.t136 2.23109
R12678 gnd.n2596 gnd.t6 2.23109
R12679 gnd.n5015 gnd.t2 2.23109
R12680 gnd.t176 gnd.n5108 2.23109
R12681 gnd.n3580 gnd.n3570 1.93989
R12682 gnd.n3548 gnd.n3538 1.93989
R12683 gnd.n3516 gnd.n3506 1.93989
R12684 gnd.n3485 gnd.n3475 1.93989
R12685 gnd.n3453 gnd.n3443 1.93989
R12686 gnd.n3421 gnd.n3411 1.93989
R12687 gnd.n3389 gnd.n3379 1.93989
R12688 gnd.n3358 gnd.n3348 1.93989
R12689 gnd.t43 gnd.n2984 1.59378
R12690 gnd.n3163 gnd.t187 1.59378
R12691 gnd.n2409 gnd.t35 1.59378
R12692 gnd.n5899 gnd.n1110 1.27512
R12693 gnd.n4856 gnd.t161 1.27512
R12694 gnd.n4923 gnd.n1862 1.27512
R12695 gnd.n4935 gnd.n1852 1.27512
R12696 gnd.n5047 gnd.n1783 1.27512
R12697 gnd.n5059 gnd.n1772 1.27512
R12698 gnd.n5165 gnd.n1699 1.27512
R12699 gnd.n5192 gnd.n1684 1.27512
R12700 gnd.n5274 gnd.t127 1.27512
R12701 gnd.n1538 gnd.n1537 1.27512
R12702 gnd.t149 gnd.n1527 1.27512
R12703 gnd.n2826 gnd.n2818 1.16414
R12704 gnd.n3642 gnd.n2311 1.16414
R12705 gnd.n3579 gnd.n3572 1.16414
R12706 gnd.n3547 gnd.n3540 1.16414
R12707 gnd.n3515 gnd.n3508 1.16414
R12708 gnd.n3484 gnd.n3477 1.16414
R12709 gnd.n3452 gnd.n3445 1.16414
R12710 gnd.n3420 gnd.n3413 1.16414
R12711 gnd.n3388 gnd.n3381 1.16414
R12712 gnd.n3357 gnd.n3350 1.16414
R12713 gnd.n5660 gnd.n5659 0.970197
R12714 gnd.n5973 gnd.n1045 0.970197
R12715 gnd.n3563 gnd.n3531 0.962709
R12716 gnd.n3595 gnd.n3563 0.962709
R12717 gnd.n3436 gnd.n3404 0.962709
R12718 gnd.n3468 gnd.n3436 0.962709
R12719 gnd.n3072 gnd.t39 0.956468
R12720 gnd.n3237 gnd.t188 0.956468
R12721 gnd.n4841 gnd.t11 0.956468
R12722 gnd.t9 gnd.n5273 0.956468
R12723 gnd.n2 gnd.n1 0.672012
R12724 gnd.n3 gnd.n2 0.672012
R12725 gnd.n4 gnd.n3 0.672012
R12726 gnd.n5 gnd.n4 0.672012
R12727 gnd.n6 gnd.n5 0.672012
R12728 gnd.n7 gnd.n6 0.672012
R12729 gnd.n9 gnd.n8 0.672012
R12730 gnd.n10 gnd.n9 0.672012
R12731 gnd.n11 gnd.n10 0.672012
R12732 gnd.n12 gnd.n11 0.672012
R12733 gnd.n13 gnd.n12 0.672012
R12734 gnd.n14 gnd.n13 0.672012
R12735 gnd.n4882 gnd.t193 0.637812
R12736 gnd.t192 gnd.n1792 0.637812
R12737 gnd.n1756 gnd.t186 0.637812
R12738 gnd.t47 gnd.n1656 0.637812
R12739 gnd.n1645 gnd.t108 0.637812
R12740 gnd gnd.n0 0.59317
R12741 gnd.n2538 gnd.n2537 0.573776
R12742 gnd.n2537 gnd.n2535 0.573776
R12743 gnd.n2535 gnd.n2533 0.573776
R12744 gnd.n2533 gnd.n2531 0.573776
R12745 gnd.n2531 gnd.n2529 0.573776
R12746 gnd.n2529 gnd.n2527 0.573776
R12747 gnd.n2527 gnd.n2525 0.573776
R12748 gnd.n2491 gnd.n2490 0.573776
R12749 gnd.n2490 gnd.n2488 0.573776
R12750 gnd.n2488 gnd.n2486 0.573776
R12751 gnd.n2486 gnd.n2484 0.573776
R12752 gnd.n2484 gnd.n2482 0.573776
R12753 gnd.n2482 gnd.n2480 0.573776
R12754 gnd.n2480 gnd.n2478 0.573776
R12755 gnd.n2506 gnd.n2505 0.573776
R12756 gnd.n2505 gnd.n2503 0.573776
R12757 gnd.n2503 gnd.n2501 0.573776
R12758 gnd.n2501 gnd.n2499 0.573776
R12759 gnd.n2499 gnd.n2497 0.573776
R12760 gnd.n2497 gnd.n2495 0.573776
R12761 gnd.n2495 gnd.n2493 0.573776
R12762 gnd.n2522 gnd.n2521 0.573776
R12763 gnd.n2521 gnd.n2519 0.573776
R12764 gnd.n2519 gnd.n2517 0.573776
R12765 gnd.n2517 gnd.n2515 0.573776
R12766 gnd.n2515 gnd.n2513 0.573776
R12767 gnd.n2513 gnd.n2511 0.573776
R12768 gnd.n2511 gnd.n2509 0.573776
R12769 gnd.n66 gnd.n64 0.573776
R12770 gnd.n68 gnd.n66 0.573776
R12771 gnd.n70 gnd.n68 0.573776
R12772 gnd.n72 gnd.n70 0.573776
R12773 gnd.n74 gnd.n72 0.573776
R12774 gnd.n76 gnd.n74 0.573776
R12775 gnd.n77 gnd.n76 0.573776
R12776 gnd.n19 gnd.n17 0.573776
R12777 gnd.n21 gnd.n19 0.573776
R12778 gnd.n23 gnd.n21 0.573776
R12779 gnd.n25 gnd.n23 0.573776
R12780 gnd.n27 gnd.n25 0.573776
R12781 gnd.n29 gnd.n27 0.573776
R12782 gnd.n30 gnd.n29 0.573776
R12783 gnd.n34 gnd.n32 0.573776
R12784 gnd.n36 gnd.n34 0.573776
R12785 gnd.n38 gnd.n36 0.573776
R12786 gnd.n40 gnd.n38 0.573776
R12787 gnd.n42 gnd.n40 0.573776
R12788 gnd.n44 gnd.n42 0.573776
R12789 gnd.n45 gnd.n44 0.573776
R12790 gnd.n50 gnd.n48 0.573776
R12791 gnd.n52 gnd.n50 0.573776
R12792 gnd.n54 gnd.n52 0.573776
R12793 gnd.n56 gnd.n54 0.573776
R12794 gnd.n58 gnd.n56 0.573776
R12795 gnd.n60 gnd.n58 0.573776
R12796 gnd.n61 gnd.n60 0.573776
R12797 gnd.n7270 gnd.n7269 0.553533
R12798 gnd.n7021 gnd.n6966 0.505073
R12799 gnd.n3880 gnd.n3878 0.505073
R12800 gnd.n5784 gnd.n1216 0.489829
R12801 gnd.n4630 gnd.n2005 0.489829
R12802 gnd.n4349 gnd.n4341 0.489829
R12803 gnd.n5778 gnd.n5777 0.489829
R12804 gnd.n3299 gnd.n2315 0.486781
R12805 gnd.n2875 gnd.n2874 0.48678
R12806 gnd.n3616 gnd.n2269 0.480683
R12807 gnd.n2959 gnd.n2958 0.480683
R12808 gnd.n1415 gnd.n1334 0.470012
R12809 gnd.n7187 gnd.n7186 0.470012
R12810 gnd.n6027 gnd.n6026 0.470012
R12811 gnd.n3762 gnd.n2231 0.470012
R12812 gnd.n6252 gnd.n6251 0.416659
R12813 gnd.n6574 gnd.n6573 0.416659
R12814 gnd.n6785 gnd.n394 0.416659
R12815 gnd.n4294 gnd.n881 0.416659
R12816 gnd.n4425 gnd.n4416 0.388379
R12817 gnd.n3576 gnd.n3575 0.388379
R12818 gnd.n3544 gnd.n3543 0.388379
R12819 gnd.n3512 gnd.n3511 0.388379
R12820 gnd.n3481 gnd.n3480 0.388379
R12821 gnd.n3449 gnd.n3448 0.388379
R12822 gnd.n3417 gnd.n3416 0.388379
R12823 gnd.n3385 gnd.n3384 0.388379
R12824 gnd.n3354 gnd.n3353 0.388379
R12825 gnd.n5722 gnd.n1282 0.388379
R12826 gnd.n7270 gnd.n15 0.374463
R12827 gnd.n2371 gnd.t195 0.319156
R12828 gnd.n4974 gnd.t31 0.319156
R12829 gnd.t28 gnd.t360 0.319156
R12830 gnd.t22 gnd.t13 0.319156
R12831 gnd.n5153 gnd.t174 0.319156
R12832 gnd.n2793 gnd.n2771 0.311721
R12833 gnd gnd.n7270 0.295112
R12834 gnd.n7063 gnd.n308 0.293183
R12835 gnd.n3918 gnd.n3917 0.293183
R12836 gnd.n4629 gnd.n2032 0.27489
R12837 gnd.n5467 gnd.n5466 0.27489
R12838 gnd.n3687 gnd.n3686 0.268793
R12839 gnd.n5598 gnd.n1235 0.258122
R12840 gnd.n7064 gnd.n7063 0.258122
R12841 gnd.n4577 gnd.n4576 0.258122
R12842 gnd.n3919 gnd.n3918 0.258122
R12843 gnd.n3686 gnd.n3685 0.241354
R12844 gnd.n1364 gnd.n1361 0.229039
R12845 gnd.n1365 gnd.n1364 0.229039
R12846 gnd.n1047 gnd.n1044 0.229039
R12847 gnd.n4501 gnd.n1047 0.229039
R12848 gnd.n2947 gnd.n2746 0.206293
R12849 gnd.n2540 gnd.n0 0.169152
R12850 gnd.n3593 gnd.n3565 0.155672
R12851 gnd.n3586 gnd.n3565 0.155672
R12852 gnd.n3586 gnd.n3585 0.155672
R12853 gnd.n3585 gnd.n3569 0.155672
R12854 gnd.n3578 gnd.n3569 0.155672
R12855 gnd.n3578 gnd.n3577 0.155672
R12856 gnd.n3561 gnd.n3533 0.155672
R12857 gnd.n3554 gnd.n3533 0.155672
R12858 gnd.n3554 gnd.n3553 0.155672
R12859 gnd.n3553 gnd.n3537 0.155672
R12860 gnd.n3546 gnd.n3537 0.155672
R12861 gnd.n3546 gnd.n3545 0.155672
R12862 gnd.n3529 gnd.n3501 0.155672
R12863 gnd.n3522 gnd.n3501 0.155672
R12864 gnd.n3522 gnd.n3521 0.155672
R12865 gnd.n3521 gnd.n3505 0.155672
R12866 gnd.n3514 gnd.n3505 0.155672
R12867 gnd.n3514 gnd.n3513 0.155672
R12868 gnd.n3498 gnd.n3470 0.155672
R12869 gnd.n3491 gnd.n3470 0.155672
R12870 gnd.n3491 gnd.n3490 0.155672
R12871 gnd.n3490 gnd.n3474 0.155672
R12872 gnd.n3483 gnd.n3474 0.155672
R12873 gnd.n3483 gnd.n3482 0.155672
R12874 gnd.n3466 gnd.n3438 0.155672
R12875 gnd.n3459 gnd.n3438 0.155672
R12876 gnd.n3459 gnd.n3458 0.155672
R12877 gnd.n3458 gnd.n3442 0.155672
R12878 gnd.n3451 gnd.n3442 0.155672
R12879 gnd.n3451 gnd.n3450 0.155672
R12880 gnd.n3434 gnd.n3406 0.155672
R12881 gnd.n3427 gnd.n3406 0.155672
R12882 gnd.n3427 gnd.n3426 0.155672
R12883 gnd.n3426 gnd.n3410 0.155672
R12884 gnd.n3419 gnd.n3410 0.155672
R12885 gnd.n3419 gnd.n3418 0.155672
R12886 gnd.n3402 gnd.n3374 0.155672
R12887 gnd.n3395 gnd.n3374 0.155672
R12888 gnd.n3395 gnd.n3394 0.155672
R12889 gnd.n3394 gnd.n3378 0.155672
R12890 gnd.n3387 gnd.n3378 0.155672
R12891 gnd.n3387 gnd.n3386 0.155672
R12892 gnd.n3371 gnd.n3343 0.155672
R12893 gnd.n3364 gnd.n3343 0.155672
R12894 gnd.n3364 gnd.n3363 0.155672
R12895 gnd.n3363 gnd.n3347 0.155672
R12896 gnd.n3356 gnd.n3347 0.155672
R12897 gnd.n3356 gnd.n3355 0.155672
R12898 gnd.n1335 gnd.n1334 0.152939
R12899 gnd.n1336 gnd.n1335 0.152939
R12900 gnd.n1337 gnd.n1336 0.152939
R12901 gnd.n1338 gnd.n1337 0.152939
R12902 gnd.n1339 gnd.n1338 0.152939
R12903 gnd.n1340 gnd.n1339 0.152939
R12904 gnd.n1341 gnd.n1340 0.152939
R12905 gnd.n1342 gnd.n1341 0.152939
R12906 gnd.n1343 gnd.n1342 0.152939
R12907 gnd.n1344 gnd.n1343 0.152939
R12908 gnd.n1345 gnd.n1344 0.152939
R12909 gnd.n1346 gnd.n1345 0.152939
R12910 gnd.n1347 gnd.n1346 0.152939
R12911 gnd.n1348 gnd.n1347 0.152939
R12912 gnd.n1349 gnd.n1348 0.152939
R12913 gnd.n1350 gnd.n1349 0.152939
R12914 gnd.n1351 gnd.n1350 0.152939
R12915 gnd.n1354 gnd.n1351 0.152939
R12916 gnd.n1355 gnd.n1354 0.152939
R12917 gnd.n1356 gnd.n1355 0.152939
R12918 gnd.n1357 gnd.n1356 0.152939
R12919 gnd.n1358 gnd.n1357 0.152939
R12920 gnd.n1359 gnd.n1358 0.152939
R12921 gnd.n1360 gnd.n1359 0.152939
R12922 gnd.n1361 gnd.n1360 0.152939
R12923 gnd.n1366 gnd.n1365 0.152939
R12924 gnd.n1367 gnd.n1366 0.152939
R12925 gnd.n1368 gnd.n1367 0.152939
R12926 gnd.n1369 gnd.n1368 0.152939
R12927 gnd.n1370 gnd.n1369 0.152939
R12928 gnd.n1371 gnd.n1370 0.152939
R12929 gnd.n1372 gnd.n1371 0.152939
R12930 gnd.n1373 gnd.n1372 0.152939
R12931 gnd.n1374 gnd.n1373 0.152939
R12932 gnd.n1377 gnd.n1374 0.152939
R12933 gnd.n1378 gnd.n1377 0.152939
R12934 gnd.n1379 gnd.n1378 0.152939
R12935 gnd.n1380 gnd.n1379 0.152939
R12936 gnd.n1381 gnd.n1380 0.152939
R12937 gnd.n1382 gnd.n1381 0.152939
R12938 gnd.n1383 gnd.n1382 0.152939
R12939 gnd.n1384 gnd.n1383 0.152939
R12940 gnd.n1385 gnd.n1384 0.152939
R12941 gnd.n1386 gnd.n1385 0.152939
R12942 gnd.n1387 gnd.n1386 0.152939
R12943 gnd.n1388 gnd.n1387 0.152939
R12944 gnd.n1389 gnd.n1388 0.152939
R12945 gnd.n1390 gnd.n1389 0.152939
R12946 gnd.n1391 gnd.n1390 0.152939
R12947 gnd.n1392 gnd.n1391 0.152939
R12948 gnd.n1393 gnd.n1392 0.152939
R12949 gnd.n1394 gnd.n1393 0.152939
R12950 gnd.n1395 gnd.n1394 0.152939
R12951 gnd.n5599 gnd.n1395 0.152939
R12952 gnd.n5599 gnd.n5598 0.152939
R12953 gnd.n1416 gnd.n1415 0.152939
R12954 gnd.n1417 gnd.n1416 0.152939
R12955 gnd.n1418 gnd.n1417 0.152939
R12956 gnd.n1419 gnd.n1418 0.152939
R12957 gnd.n1437 gnd.n1419 0.152939
R12958 gnd.n1438 gnd.n1437 0.152939
R12959 gnd.n1439 gnd.n1438 0.152939
R12960 gnd.n1440 gnd.n1439 0.152939
R12961 gnd.n5556 gnd.n1440 0.152939
R12962 gnd.n5557 gnd.n5556 0.152939
R12963 gnd.n5558 gnd.n5557 0.152939
R12964 gnd.n5558 gnd.n376 0.152939
R12965 gnd.n6810 gnd.n376 0.152939
R12966 gnd.n6811 gnd.n6810 0.152939
R12967 gnd.n6812 gnd.n6811 0.152939
R12968 gnd.n6813 gnd.n6812 0.152939
R12969 gnd.n6813 gnd.n348 0.152939
R12970 gnd.n6844 gnd.n348 0.152939
R12971 gnd.n6845 gnd.n6844 0.152939
R12972 gnd.n6846 gnd.n6845 0.152939
R12973 gnd.n6847 gnd.n6846 0.152939
R12974 gnd.n113 gnd.n112 0.152939
R12975 gnd.n114 gnd.n113 0.152939
R12976 gnd.n130 gnd.n114 0.152939
R12977 gnd.n131 gnd.n130 0.152939
R12978 gnd.n132 gnd.n131 0.152939
R12979 gnd.n133 gnd.n132 0.152939
R12980 gnd.n149 gnd.n133 0.152939
R12981 gnd.n150 gnd.n149 0.152939
R12982 gnd.n151 gnd.n150 0.152939
R12983 gnd.n152 gnd.n151 0.152939
R12984 gnd.n168 gnd.n152 0.152939
R12985 gnd.n169 gnd.n168 0.152939
R12986 gnd.n170 gnd.n169 0.152939
R12987 gnd.n171 gnd.n170 0.152939
R12988 gnd.n187 gnd.n171 0.152939
R12989 gnd.n188 gnd.n187 0.152939
R12990 gnd.n189 gnd.n188 0.152939
R12991 gnd.n190 gnd.n189 0.152939
R12992 gnd.n206 gnd.n190 0.152939
R12993 gnd.n207 gnd.n206 0.152939
R12994 gnd.n7187 gnd.n207 0.152939
R12995 gnd.n7267 gnd.n80 0.152939
R12996 gnd.n6930 gnd.n80 0.152939
R12997 gnd.n6931 gnd.n6930 0.152939
R12998 gnd.n6932 gnd.n6931 0.152939
R12999 gnd.n6932 gnd.n6928 0.152939
R13000 gnd.n6938 gnd.n6928 0.152939
R13001 gnd.n6939 gnd.n6938 0.152939
R13002 gnd.n6940 gnd.n6939 0.152939
R13003 gnd.n6940 gnd.n6926 0.152939
R13004 gnd.n6946 gnd.n6926 0.152939
R13005 gnd.n6947 gnd.n6946 0.152939
R13006 gnd.n6948 gnd.n6947 0.152939
R13007 gnd.n6948 gnd.n6924 0.152939
R13008 gnd.n6954 gnd.n6924 0.152939
R13009 gnd.n6955 gnd.n6954 0.152939
R13010 gnd.n6956 gnd.n6955 0.152939
R13011 gnd.n6957 gnd.n6956 0.152939
R13012 gnd.n6958 gnd.n6957 0.152939
R13013 gnd.n6959 gnd.n6958 0.152939
R13014 gnd.n6960 gnd.n6959 0.152939
R13015 gnd.n6961 gnd.n6960 0.152939
R13016 gnd.n6962 gnd.n6961 0.152939
R13017 gnd.n6963 gnd.n6962 0.152939
R13018 gnd.n6964 gnd.n6963 0.152939
R13019 gnd.n6965 gnd.n6964 0.152939
R13020 gnd.n6966 gnd.n6965 0.152939
R13021 gnd.n6980 gnd.n308 0.152939
R13022 gnd.n6981 gnd.n6980 0.152939
R13023 gnd.n6981 gnd.n6976 0.152939
R13024 gnd.n6989 gnd.n6976 0.152939
R13025 gnd.n6990 gnd.n6989 0.152939
R13026 gnd.n6991 gnd.n6990 0.152939
R13027 gnd.n6991 gnd.n6974 0.152939
R13028 gnd.n6999 gnd.n6974 0.152939
R13029 gnd.n7000 gnd.n6999 0.152939
R13030 gnd.n7001 gnd.n7000 0.152939
R13031 gnd.n7001 gnd.n6972 0.152939
R13032 gnd.n7009 gnd.n6972 0.152939
R13033 gnd.n7010 gnd.n7009 0.152939
R13034 gnd.n7011 gnd.n7010 0.152939
R13035 gnd.n7011 gnd.n6970 0.152939
R13036 gnd.n7019 gnd.n6970 0.152939
R13037 gnd.n7020 gnd.n7019 0.152939
R13038 gnd.n7021 gnd.n7020 0.152939
R13039 gnd.n7186 gnd.n208 0.152939
R13040 gnd.n250 gnd.n208 0.152939
R13041 gnd.n251 gnd.n250 0.152939
R13042 gnd.n252 gnd.n251 0.152939
R13043 gnd.n253 gnd.n252 0.152939
R13044 gnd.n254 gnd.n253 0.152939
R13045 gnd.n255 gnd.n254 0.152939
R13046 gnd.n256 gnd.n255 0.152939
R13047 gnd.n257 gnd.n256 0.152939
R13048 gnd.n258 gnd.n257 0.152939
R13049 gnd.n259 gnd.n258 0.152939
R13050 gnd.n260 gnd.n259 0.152939
R13051 gnd.n261 gnd.n260 0.152939
R13052 gnd.n262 gnd.n261 0.152939
R13053 gnd.n263 gnd.n262 0.152939
R13054 gnd.n264 gnd.n263 0.152939
R13055 gnd.n265 gnd.n264 0.152939
R13056 gnd.n266 gnd.n265 0.152939
R13057 gnd.n267 gnd.n266 0.152939
R13058 gnd.n268 gnd.n267 0.152939
R13059 gnd.n269 gnd.n268 0.152939
R13060 gnd.n270 gnd.n269 0.152939
R13061 gnd.n271 gnd.n270 0.152939
R13062 gnd.n272 gnd.n271 0.152939
R13063 gnd.n273 gnd.n272 0.152939
R13064 gnd.n274 gnd.n273 0.152939
R13065 gnd.n275 gnd.n274 0.152939
R13066 gnd.n276 gnd.n275 0.152939
R13067 gnd.n277 gnd.n276 0.152939
R13068 gnd.n278 gnd.n277 0.152939
R13069 gnd.n279 gnd.n278 0.152939
R13070 gnd.n280 gnd.n279 0.152939
R13071 gnd.n281 gnd.n280 0.152939
R13072 gnd.n282 gnd.n281 0.152939
R13073 gnd.n283 gnd.n282 0.152939
R13074 gnd.n284 gnd.n283 0.152939
R13075 gnd.n7107 gnd.n284 0.152939
R13076 gnd.n7107 gnd.n7106 0.152939
R13077 gnd.n7106 gnd.n7105 0.152939
R13078 gnd.n7105 gnd.n288 0.152939
R13079 gnd.n289 gnd.n288 0.152939
R13080 gnd.n290 gnd.n289 0.152939
R13081 gnd.n291 gnd.n290 0.152939
R13082 gnd.n292 gnd.n291 0.152939
R13083 gnd.n293 gnd.n292 0.152939
R13084 gnd.n294 gnd.n293 0.152939
R13085 gnd.n295 gnd.n294 0.152939
R13086 gnd.n296 gnd.n295 0.152939
R13087 gnd.n297 gnd.n296 0.152939
R13088 gnd.n298 gnd.n297 0.152939
R13089 gnd.n299 gnd.n298 0.152939
R13090 gnd.n300 gnd.n299 0.152939
R13091 gnd.n301 gnd.n300 0.152939
R13092 gnd.n302 gnd.n301 0.152939
R13093 gnd.n303 gnd.n302 0.152939
R13094 gnd.n304 gnd.n303 0.152939
R13095 gnd.n7065 gnd.n304 0.152939
R13096 gnd.n7065 gnd.n7064 0.152939
R13097 gnd.n3718 gnd.n2269 0.152939
R13098 gnd.n3718 gnd.n3717 0.152939
R13099 gnd.n3717 gnd.n3716 0.152939
R13100 gnd.n3716 gnd.n2271 0.152939
R13101 gnd.n2272 gnd.n2271 0.152939
R13102 gnd.n2273 gnd.n2272 0.152939
R13103 gnd.n2274 gnd.n2273 0.152939
R13104 gnd.n2275 gnd.n2274 0.152939
R13105 gnd.n2276 gnd.n2275 0.152939
R13106 gnd.n2277 gnd.n2276 0.152939
R13107 gnd.n2278 gnd.n2277 0.152939
R13108 gnd.n2279 gnd.n2278 0.152939
R13109 gnd.n2280 gnd.n2279 0.152939
R13110 gnd.n2281 gnd.n2280 0.152939
R13111 gnd.n3688 gnd.n2281 0.152939
R13112 gnd.n3688 gnd.n3687 0.152939
R13113 gnd.n2960 gnd.n2959 0.152939
R13114 gnd.n2960 gnd.n2664 0.152939
R13115 gnd.n2988 gnd.n2664 0.152939
R13116 gnd.n2989 gnd.n2988 0.152939
R13117 gnd.n2990 gnd.n2989 0.152939
R13118 gnd.n2991 gnd.n2990 0.152939
R13119 gnd.n2991 gnd.n2636 0.152939
R13120 gnd.n3018 gnd.n2636 0.152939
R13121 gnd.n3019 gnd.n3018 0.152939
R13122 gnd.n3020 gnd.n3019 0.152939
R13123 gnd.n3020 gnd.n2614 0.152939
R13124 gnd.n3049 gnd.n2614 0.152939
R13125 gnd.n3050 gnd.n3049 0.152939
R13126 gnd.n3051 gnd.n3050 0.152939
R13127 gnd.n3052 gnd.n3051 0.152939
R13128 gnd.n3054 gnd.n3052 0.152939
R13129 gnd.n3054 gnd.n3053 0.152939
R13130 gnd.n3053 gnd.n2563 0.152939
R13131 gnd.n2564 gnd.n2563 0.152939
R13132 gnd.n2565 gnd.n2564 0.152939
R13133 gnd.n2584 gnd.n2565 0.152939
R13134 gnd.n2585 gnd.n2584 0.152939
R13135 gnd.n2585 gnd.n2467 0.152939
R13136 gnd.n3144 gnd.n2467 0.152939
R13137 gnd.n3145 gnd.n3144 0.152939
R13138 gnd.n3146 gnd.n3145 0.152939
R13139 gnd.n3147 gnd.n3146 0.152939
R13140 gnd.n3147 gnd.n2440 0.152939
R13141 gnd.n3184 gnd.n2440 0.152939
R13142 gnd.n3185 gnd.n3184 0.152939
R13143 gnd.n3186 gnd.n3185 0.152939
R13144 gnd.n3187 gnd.n3186 0.152939
R13145 gnd.n3187 gnd.n2413 0.152939
R13146 gnd.n3229 gnd.n2413 0.152939
R13147 gnd.n3230 gnd.n3229 0.152939
R13148 gnd.n3231 gnd.n3230 0.152939
R13149 gnd.n3232 gnd.n3231 0.152939
R13150 gnd.n3232 gnd.n2385 0.152939
R13151 gnd.n3269 gnd.n2385 0.152939
R13152 gnd.n3270 gnd.n3269 0.152939
R13153 gnd.n3271 gnd.n3270 0.152939
R13154 gnd.n3272 gnd.n3271 0.152939
R13155 gnd.n3272 gnd.n2358 0.152939
R13156 gnd.n3318 gnd.n2358 0.152939
R13157 gnd.n3319 gnd.n3318 0.152939
R13158 gnd.n3320 gnd.n3319 0.152939
R13159 gnd.n3321 gnd.n3320 0.152939
R13160 gnd.n3321 gnd.n2331 0.152939
R13161 gnd.n3612 gnd.n2331 0.152939
R13162 gnd.n3613 gnd.n3612 0.152939
R13163 gnd.n3614 gnd.n3613 0.152939
R13164 gnd.n3615 gnd.n3614 0.152939
R13165 gnd.n3616 gnd.n3615 0.152939
R13166 gnd.n2958 gnd.n2688 0.152939
R13167 gnd.n2709 gnd.n2688 0.152939
R13168 gnd.n2710 gnd.n2709 0.152939
R13169 gnd.n2716 gnd.n2710 0.152939
R13170 gnd.n2717 gnd.n2716 0.152939
R13171 gnd.n2718 gnd.n2717 0.152939
R13172 gnd.n2718 gnd.n2707 0.152939
R13173 gnd.n2726 gnd.n2707 0.152939
R13174 gnd.n2727 gnd.n2726 0.152939
R13175 gnd.n2728 gnd.n2727 0.152939
R13176 gnd.n2728 gnd.n2705 0.152939
R13177 gnd.n2736 gnd.n2705 0.152939
R13178 gnd.n2737 gnd.n2736 0.152939
R13179 gnd.n2738 gnd.n2737 0.152939
R13180 gnd.n2738 gnd.n2703 0.152939
R13181 gnd.n2746 gnd.n2703 0.152939
R13182 gnd.n3685 gnd.n2286 0.152939
R13183 gnd.n2288 gnd.n2286 0.152939
R13184 gnd.n2289 gnd.n2288 0.152939
R13185 gnd.n2290 gnd.n2289 0.152939
R13186 gnd.n2291 gnd.n2290 0.152939
R13187 gnd.n2292 gnd.n2291 0.152939
R13188 gnd.n2293 gnd.n2292 0.152939
R13189 gnd.n2294 gnd.n2293 0.152939
R13190 gnd.n2295 gnd.n2294 0.152939
R13191 gnd.n2296 gnd.n2295 0.152939
R13192 gnd.n2297 gnd.n2296 0.152939
R13193 gnd.n2298 gnd.n2297 0.152939
R13194 gnd.n2299 gnd.n2298 0.152939
R13195 gnd.n2300 gnd.n2299 0.152939
R13196 gnd.n2301 gnd.n2300 0.152939
R13197 gnd.n2302 gnd.n2301 0.152939
R13198 gnd.n2303 gnd.n2302 0.152939
R13199 gnd.n2304 gnd.n2303 0.152939
R13200 gnd.n2305 gnd.n2304 0.152939
R13201 gnd.n2306 gnd.n2305 0.152939
R13202 gnd.n2307 gnd.n2306 0.152939
R13203 gnd.n2308 gnd.n2307 0.152939
R13204 gnd.n2312 gnd.n2308 0.152939
R13205 gnd.n2313 gnd.n2312 0.152939
R13206 gnd.n2314 gnd.n2313 0.152939
R13207 gnd.n2315 gnd.n2314 0.152939
R13208 gnd.n3121 gnd.n3120 0.152939
R13209 gnd.n3122 gnd.n3121 0.152939
R13210 gnd.n3123 gnd.n3122 0.152939
R13211 gnd.n3124 gnd.n3123 0.152939
R13212 gnd.n3125 gnd.n3124 0.152939
R13213 gnd.n3126 gnd.n3125 0.152939
R13214 gnd.n3126 gnd.n2421 0.152939
R13215 gnd.n3205 gnd.n2421 0.152939
R13216 gnd.n3206 gnd.n3205 0.152939
R13217 gnd.n3207 gnd.n3206 0.152939
R13218 gnd.n3208 gnd.n3207 0.152939
R13219 gnd.n3209 gnd.n3208 0.152939
R13220 gnd.n3210 gnd.n3209 0.152939
R13221 gnd.n3211 gnd.n3210 0.152939
R13222 gnd.n3212 gnd.n3211 0.152939
R13223 gnd.n3213 gnd.n3212 0.152939
R13224 gnd.n3213 gnd.n2365 0.152939
R13225 gnd.n3290 gnd.n2365 0.152939
R13226 gnd.n3291 gnd.n3290 0.152939
R13227 gnd.n3292 gnd.n3291 0.152939
R13228 gnd.n3293 gnd.n3292 0.152939
R13229 gnd.n3294 gnd.n3293 0.152939
R13230 gnd.n3295 gnd.n3294 0.152939
R13231 gnd.n3296 gnd.n3295 0.152939
R13232 gnd.n3297 gnd.n3296 0.152939
R13233 gnd.n3298 gnd.n3297 0.152939
R13234 gnd.n3300 gnd.n3298 0.152939
R13235 gnd.n3300 gnd.n3299 0.152939
R13236 gnd.n2876 gnd.n2875 0.152939
R13237 gnd.n2876 gnd.n2766 0.152939
R13238 gnd.n2891 gnd.n2766 0.152939
R13239 gnd.n2892 gnd.n2891 0.152939
R13240 gnd.n2893 gnd.n2892 0.152939
R13241 gnd.n2893 gnd.n2754 0.152939
R13242 gnd.n2907 gnd.n2754 0.152939
R13243 gnd.n2908 gnd.n2907 0.152939
R13244 gnd.n2909 gnd.n2908 0.152939
R13245 gnd.n2910 gnd.n2909 0.152939
R13246 gnd.n2911 gnd.n2910 0.152939
R13247 gnd.n2912 gnd.n2911 0.152939
R13248 gnd.n2913 gnd.n2912 0.152939
R13249 gnd.n2914 gnd.n2913 0.152939
R13250 gnd.n2915 gnd.n2914 0.152939
R13251 gnd.n2916 gnd.n2915 0.152939
R13252 gnd.n2917 gnd.n2916 0.152939
R13253 gnd.n2918 gnd.n2917 0.152939
R13254 gnd.n2919 gnd.n2918 0.152939
R13255 gnd.n2920 gnd.n2919 0.152939
R13256 gnd.n2921 gnd.n2920 0.152939
R13257 gnd.n2921 gnd.n2620 0.152939
R13258 gnd.n3038 gnd.n2620 0.152939
R13259 gnd.n3039 gnd.n3038 0.152939
R13260 gnd.n3040 gnd.n3039 0.152939
R13261 gnd.n3041 gnd.n3040 0.152939
R13262 gnd.n3041 gnd.n2542 0.152939
R13263 gnd.n3118 gnd.n2542 0.152939
R13264 gnd.n2794 gnd.n2793 0.152939
R13265 gnd.n2795 gnd.n2794 0.152939
R13266 gnd.n2796 gnd.n2795 0.152939
R13267 gnd.n2797 gnd.n2796 0.152939
R13268 gnd.n2798 gnd.n2797 0.152939
R13269 gnd.n2799 gnd.n2798 0.152939
R13270 gnd.n2800 gnd.n2799 0.152939
R13271 gnd.n2801 gnd.n2800 0.152939
R13272 gnd.n2802 gnd.n2801 0.152939
R13273 gnd.n2803 gnd.n2802 0.152939
R13274 gnd.n2804 gnd.n2803 0.152939
R13275 gnd.n2805 gnd.n2804 0.152939
R13276 gnd.n2806 gnd.n2805 0.152939
R13277 gnd.n2807 gnd.n2806 0.152939
R13278 gnd.n2808 gnd.n2807 0.152939
R13279 gnd.n2809 gnd.n2808 0.152939
R13280 gnd.n2810 gnd.n2809 0.152939
R13281 gnd.n2811 gnd.n2810 0.152939
R13282 gnd.n2812 gnd.n2811 0.152939
R13283 gnd.n2813 gnd.n2812 0.152939
R13284 gnd.n2814 gnd.n2813 0.152939
R13285 gnd.n2815 gnd.n2814 0.152939
R13286 gnd.n2819 gnd.n2815 0.152939
R13287 gnd.n2820 gnd.n2819 0.152939
R13288 gnd.n2820 gnd.n2777 0.152939
R13289 gnd.n2874 gnd.n2777 0.152939
R13290 gnd.n3878 gnd.n3844 0.152939
R13291 gnd.n3845 gnd.n3844 0.152939
R13292 gnd.n3846 gnd.n3845 0.152939
R13293 gnd.n3847 gnd.n3846 0.152939
R13294 gnd.n3848 gnd.n3847 0.152939
R13295 gnd.n3849 gnd.n3848 0.152939
R13296 gnd.n3850 gnd.n3849 0.152939
R13297 gnd.n3851 gnd.n3850 0.152939
R13298 gnd.n3852 gnd.n3851 0.152939
R13299 gnd.n3853 gnd.n3852 0.152939
R13300 gnd.n3854 gnd.n3853 0.152939
R13301 gnd.n3855 gnd.n3854 0.152939
R13302 gnd.n3856 gnd.n3855 0.152939
R13303 gnd.n3856 gnd.n2167 0.152939
R13304 gnd.n4126 gnd.n2167 0.152939
R13305 gnd.n4127 gnd.n4126 0.152939
R13306 gnd.n4128 gnd.n4127 0.152939
R13307 gnd.n4129 gnd.n4128 0.152939
R13308 gnd.n4129 gnd.n2142 0.152939
R13309 gnd.n4161 gnd.n2142 0.152939
R13310 gnd.n4162 gnd.n4161 0.152939
R13311 gnd.n4163 gnd.n4162 0.152939
R13312 gnd.n4164 gnd.n4163 0.152939
R13313 gnd.n4164 gnd.n2117 0.152939
R13314 gnd.n4196 gnd.n2117 0.152939
R13315 gnd.n4197 gnd.n4196 0.152939
R13316 gnd.n6026 gnd.n975 0.152939
R13317 gnd.n1019 gnd.n975 0.152939
R13318 gnd.n1020 gnd.n1019 0.152939
R13319 gnd.n1021 gnd.n1020 0.152939
R13320 gnd.n1022 gnd.n1021 0.152939
R13321 gnd.n1023 gnd.n1022 0.152939
R13322 gnd.n1024 gnd.n1023 0.152939
R13323 gnd.n1025 gnd.n1024 0.152939
R13324 gnd.n1026 gnd.n1025 0.152939
R13325 gnd.n1027 gnd.n1026 0.152939
R13326 gnd.n1028 gnd.n1027 0.152939
R13327 gnd.n1029 gnd.n1028 0.152939
R13328 gnd.n1030 gnd.n1029 0.152939
R13329 gnd.n1031 gnd.n1030 0.152939
R13330 gnd.n1032 gnd.n1031 0.152939
R13331 gnd.n1033 gnd.n1032 0.152939
R13332 gnd.n1034 gnd.n1033 0.152939
R13333 gnd.n1037 gnd.n1034 0.152939
R13334 gnd.n1038 gnd.n1037 0.152939
R13335 gnd.n1039 gnd.n1038 0.152939
R13336 gnd.n1040 gnd.n1039 0.152939
R13337 gnd.n1041 gnd.n1040 0.152939
R13338 gnd.n1042 gnd.n1041 0.152939
R13339 gnd.n1043 gnd.n1042 0.152939
R13340 gnd.n1044 gnd.n1043 0.152939
R13341 gnd.n4502 gnd.n4501 0.152939
R13342 gnd.n4509 gnd.n4502 0.152939
R13343 gnd.n4510 gnd.n4509 0.152939
R13344 gnd.n4511 gnd.n4510 0.152939
R13345 gnd.n4511 gnd.n4499 0.152939
R13346 gnd.n4519 gnd.n4499 0.152939
R13347 gnd.n4520 gnd.n4519 0.152939
R13348 gnd.n4521 gnd.n4520 0.152939
R13349 gnd.n4521 gnd.n4494 0.152939
R13350 gnd.n4528 gnd.n4494 0.152939
R13351 gnd.n4529 gnd.n4528 0.152939
R13352 gnd.n4530 gnd.n4529 0.152939
R13353 gnd.n4530 gnd.n4492 0.152939
R13354 gnd.n4538 gnd.n4492 0.152939
R13355 gnd.n4539 gnd.n4538 0.152939
R13356 gnd.n4540 gnd.n4539 0.152939
R13357 gnd.n4540 gnd.n4490 0.152939
R13358 gnd.n4548 gnd.n4490 0.152939
R13359 gnd.n4549 gnd.n4548 0.152939
R13360 gnd.n4550 gnd.n4549 0.152939
R13361 gnd.n4550 gnd.n4488 0.152939
R13362 gnd.n4558 gnd.n4488 0.152939
R13363 gnd.n4559 gnd.n4558 0.152939
R13364 gnd.n4560 gnd.n4559 0.152939
R13365 gnd.n4560 gnd.n4486 0.152939
R13366 gnd.n4568 gnd.n4486 0.152939
R13367 gnd.n4569 gnd.n4568 0.152939
R13368 gnd.n4570 gnd.n4569 0.152939
R13369 gnd.n4570 gnd.n4481 0.152939
R13370 gnd.n4576 gnd.n4481 0.152939
R13371 gnd.n4257 gnd.n4256 0.152939
R13372 gnd.n4259 gnd.n4257 0.152939
R13373 gnd.n4259 gnd.n4258 0.152939
R13374 gnd.n4258 gnd.n891 0.152939
R13375 gnd.n892 gnd.n891 0.152939
R13376 gnd.n893 gnd.n892 0.152939
R13377 gnd.n912 gnd.n893 0.152939
R13378 gnd.n913 gnd.n912 0.152939
R13379 gnd.n914 gnd.n913 0.152939
R13380 gnd.n915 gnd.n914 0.152939
R13381 gnd.n932 gnd.n915 0.152939
R13382 gnd.n933 gnd.n932 0.152939
R13383 gnd.n934 gnd.n933 0.152939
R13384 gnd.n935 gnd.n934 0.152939
R13385 gnd.n952 gnd.n935 0.152939
R13386 gnd.n953 gnd.n952 0.152939
R13387 gnd.n954 gnd.n953 0.152939
R13388 gnd.n955 gnd.n954 0.152939
R13389 gnd.n973 gnd.n955 0.152939
R13390 gnd.n974 gnd.n973 0.152939
R13391 gnd.n6027 gnd.n974 0.152939
R13392 gnd.n4052 gnd.n2231 0.152939
R13393 gnd.n4053 gnd.n4052 0.152939
R13394 gnd.n4054 gnd.n4053 0.152939
R13395 gnd.n4054 gnd.n2212 0.152939
R13396 gnd.n4072 gnd.n2212 0.152939
R13397 gnd.n4073 gnd.n4072 0.152939
R13398 gnd.n4074 gnd.n4073 0.152939
R13399 gnd.n4074 gnd.n2195 0.152939
R13400 gnd.n4092 gnd.n2195 0.152939
R13401 gnd.n4093 gnd.n4092 0.152939
R13402 gnd.n4094 gnd.n4093 0.152939
R13403 gnd.n4094 gnd.n2175 0.152939
R13404 gnd.n4116 gnd.n2175 0.152939
R13405 gnd.n4117 gnd.n4116 0.152939
R13406 gnd.n4118 gnd.n4117 0.152939
R13407 gnd.n4119 gnd.n4118 0.152939
R13408 gnd.n4119 gnd.n2150 0.152939
R13409 gnd.n4151 gnd.n2150 0.152939
R13410 gnd.n4152 gnd.n4151 0.152939
R13411 gnd.n4153 gnd.n4152 0.152939
R13412 gnd.n4154 gnd.n4153 0.152939
R13413 gnd.n3763 gnd.n3762 0.152939
R13414 gnd.n3764 gnd.n3763 0.152939
R13415 gnd.n3765 gnd.n3764 0.152939
R13416 gnd.n3766 gnd.n3765 0.152939
R13417 gnd.n3767 gnd.n3766 0.152939
R13418 gnd.n3768 gnd.n3767 0.152939
R13419 gnd.n3769 gnd.n3768 0.152939
R13420 gnd.n3770 gnd.n3769 0.152939
R13421 gnd.n3771 gnd.n3770 0.152939
R13422 gnd.n3772 gnd.n3771 0.152939
R13423 gnd.n3773 gnd.n3772 0.152939
R13424 gnd.n3774 gnd.n3773 0.152939
R13425 gnd.n3775 gnd.n3774 0.152939
R13426 gnd.n3776 gnd.n3775 0.152939
R13427 gnd.n3777 gnd.n3776 0.152939
R13428 gnd.n3778 gnd.n3777 0.152939
R13429 gnd.n3779 gnd.n3778 0.152939
R13430 gnd.n3782 gnd.n3779 0.152939
R13431 gnd.n3783 gnd.n3782 0.152939
R13432 gnd.n3784 gnd.n3783 0.152939
R13433 gnd.n3785 gnd.n3784 0.152939
R13434 gnd.n3786 gnd.n3785 0.152939
R13435 gnd.n3787 gnd.n3786 0.152939
R13436 gnd.n3788 gnd.n3787 0.152939
R13437 gnd.n3789 gnd.n3788 0.152939
R13438 gnd.n3790 gnd.n3789 0.152939
R13439 gnd.n3791 gnd.n3790 0.152939
R13440 gnd.n3792 gnd.n3791 0.152939
R13441 gnd.n3793 gnd.n3792 0.152939
R13442 gnd.n3794 gnd.n3793 0.152939
R13443 gnd.n3795 gnd.n3794 0.152939
R13444 gnd.n3796 gnd.n3795 0.152939
R13445 gnd.n3797 gnd.n3796 0.152939
R13446 gnd.n3798 gnd.n3797 0.152939
R13447 gnd.n3799 gnd.n3798 0.152939
R13448 gnd.n3800 gnd.n3799 0.152939
R13449 gnd.n3801 gnd.n3800 0.152939
R13450 gnd.n3804 gnd.n3801 0.152939
R13451 gnd.n3805 gnd.n3804 0.152939
R13452 gnd.n3806 gnd.n3805 0.152939
R13453 gnd.n3807 gnd.n3806 0.152939
R13454 gnd.n3808 gnd.n3807 0.152939
R13455 gnd.n3809 gnd.n3808 0.152939
R13456 gnd.n3810 gnd.n3809 0.152939
R13457 gnd.n3811 gnd.n3810 0.152939
R13458 gnd.n3812 gnd.n3811 0.152939
R13459 gnd.n3813 gnd.n3812 0.152939
R13460 gnd.n3814 gnd.n3813 0.152939
R13461 gnd.n3815 gnd.n3814 0.152939
R13462 gnd.n3816 gnd.n3815 0.152939
R13463 gnd.n3817 gnd.n3816 0.152939
R13464 gnd.n3818 gnd.n3817 0.152939
R13465 gnd.n3819 gnd.n3818 0.152939
R13466 gnd.n3820 gnd.n3819 0.152939
R13467 gnd.n3821 gnd.n3820 0.152939
R13468 gnd.n3822 gnd.n3821 0.152939
R13469 gnd.n3920 gnd.n3822 0.152939
R13470 gnd.n3920 gnd.n3919 0.152939
R13471 gnd.n3917 gnd.n3825 0.152939
R13472 gnd.n3826 gnd.n3825 0.152939
R13473 gnd.n3827 gnd.n3826 0.152939
R13474 gnd.n3828 gnd.n3827 0.152939
R13475 gnd.n3829 gnd.n3828 0.152939
R13476 gnd.n3830 gnd.n3829 0.152939
R13477 gnd.n3831 gnd.n3830 0.152939
R13478 gnd.n3832 gnd.n3831 0.152939
R13479 gnd.n3833 gnd.n3832 0.152939
R13480 gnd.n3834 gnd.n3833 0.152939
R13481 gnd.n3835 gnd.n3834 0.152939
R13482 gnd.n3836 gnd.n3835 0.152939
R13483 gnd.n3837 gnd.n3836 0.152939
R13484 gnd.n3838 gnd.n3837 0.152939
R13485 gnd.n3839 gnd.n3838 0.152939
R13486 gnd.n3882 gnd.n3839 0.152939
R13487 gnd.n3882 gnd.n3881 0.152939
R13488 gnd.n3881 gnd.n3880 0.152939
R13489 gnd.n6253 gnd.n6252 0.152939
R13490 gnd.n6253 gnd.n708 0.152939
R13491 gnd.n6261 gnd.n708 0.152939
R13492 gnd.n6262 gnd.n6261 0.152939
R13493 gnd.n6263 gnd.n6262 0.152939
R13494 gnd.n6263 gnd.n702 0.152939
R13495 gnd.n6271 gnd.n702 0.152939
R13496 gnd.n6272 gnd.n6271 0.152939
R13497 gnd.n6273 gnd.n6272 0.152939
R13498 gnd.n6273 gnd.n696 0.152939
R13499 gnd.n6281 gnd.n696 0.152939
R13500 gnd.n6282 gnd.n6281 0.152939
R13501 gnd.n6283 gnd.n6282 0.152939
R13502 gnd.n6283 gnd.n690 0.152939
R13503 gnd.n6291 gnd.n690 0.152939
R13504 gnd.n6292 gnd.n6291 0.152939
R13505 gnd.n6293 gnd.n6292 0.152939
R13506 gnd.n6293 gnd.n684 0.152939
R13507 gnd.n6301 gnd.n684 0.152939
R13508 gnd.n6302 gnd.n6301 0.152939
R13509 gnd.n6303 gnd.n6302 0.152939
R13510 gnd.n6303 gnd.n678 0.152939
R13511 gnd.n6311 gnd.n678 0.152939
R13512 gnd.n6312 gnd.n6311 0.152939
R13513 gnd.n6313 gnd.n6312 0.152939
R13514 gnd.n6313 gnd.n672 0.152939
R13515 gnd.n6321 gnd.n672 0.152939
R13516 gnd.n6322 gnd.n6321 0.152939
R13517 gnd.n6323 gnd.n6322 0.152939
R13518 gnd.n6323 gnd.n666 0.152939
R13519 gnd.n6331 gnd.n666 0.152939
R13520 gnd.n6332 gnd.n6331 0.152939
R13521 gnd.n6333 gnd.n6332 0.152939
R13522 gnd.n6333 gnd.n660 0.152939
R13523 gnd.n6341 gnd.n660 0.152939
R13524 gnd.n6342 gnd.n6341 0.152939
R13525 gnd.n6343 gnd.n6342 0.152939
R13526 gnd.n6343 gnd.n654 0.152939
R13527 gnd.n6351 gnd.n654 0.152939
R13528 gnd.n6352 gnd.n6351 0.152939
R13529 gnd.n6353 gnd.n6352 0.152939
R13530 gnd.n6353 gnd.n648 0.152939
R13531 gnd.n6361 gnd.n648 0.152939
R13532 gnd.n6362 gnd.n6361 0.152939
R13533 gnd.n6363 gnd.n6362 0.152939
R13534 gnd.n6363 gnd.n642 0.152939
R13535 gnd.n6371 gnd.n642 0.152939
R13536 gnd.n6372 gnd.n6371 0.152939
R13537 gnd.n6373 gnd.n6372 0.152939
R13538 gnd.n6373 gnd.n636 0.152939
R13539 gnd.n6381 gnd.n636 0.152939
R13540 gnd.n6382 gnd.n6381 0.152939
R13541 gnd.n6383 gnd.n6382 0.152939
R13542 gnd.n6383 gnd.n630 0.152939
R13543 gnd.n6391 gnd.n630 0.152939
R13544 gnd.n6392 gnd.n6391 0.152939
R13545 gnd.n6393 gnd.n6392 0.152939
R13546 gnd.n6393 gnd.n624 0.152939
R13547 gnd.n6401 gnd.n624 0.152939
R13548 gnd.n6402 gnd.n6401 0.152939
R13549 gnd.n6403 gnd.n6402 0.152939
R13550 gnd.n6403 gnd.n618 0.152939
R13551 gnd.n6411 gnd.n618 0.152939
R13552 gnd.n6412 gnd.n6411 0.152939
R13553 gnd.n6413 gnd.n6412 0.152939
R13554 gnd.n6413 gnd.n612 0.152939
R13555 gnd.n6421 gnd.n612 0.152939
R13556 gnd.n6422 gnd.n6421 0.152939
R13557 gnd.n6423 gnd.n6422 0.152939
R13558 gnd.n6423 gnd.n606 0.152939
R13559 gnd.n6431 gnd.n606 0.152939
R13560 gnd.n6432 gnd.n6431 0.152939
R13561 gnd.n6433 gnd.n6432 0.152939
R13562 gnd.n6433 gnd.n600 0.152939
R13563 gnd.n6441 gnd.n600 0.152939
R13564 gnd.n6442 gnd.n6441 0.152939
R13565 gnd.n6443 gnd.n6442 0.152939
R13566 gnd.n6443 gnd.n594 0.152939
R13567 gnd.n6451 gnd.n594 0.152939
R13568 gnd.n6452 gnd.n6451 0.152939
R13569 gnd.n6453 gnd.n6452 0.152939
R13570 gnd.n6453 gnd.n588 0.152939
R13571 gnd.n6461 gnd.n588 0.152939
R13572 gnd.n6462 gnd.n6461 0.152939
R13573 gnd.n6463 gnd.n6462 0.152939
R13574 gnd.n6463 gnd.n582 0.152939
R13575 gnd.n6471 gnd.n582 0.152939
R13576 gnd.n6472 gnd.n6471 0.152939
R13577 gnd.n6473 gnd.n6472 0.152939
R13578 gnd.n6473 gnd.n576 0.152939
R13579 gnd.n6481 gnd.n576 0.152939
R13580 gnd.n6482 gnd.n6481 0.152939
R13581 gnd.n6483 gnd.n6482 0.152939
R13582 gnd.n6483 gnd.n570 0.152939
R13583 gnd.n6491 gnd.n570 0.152939
R13584 gnd.n6492 gnd.n6491 0.152939
R13585 gnd.n6493 gnd.n6492 0.152939
R13586 gnd.n6493 gnd.n564 0.152939
R13587 gnd.n6501 gnd.n564 0.152939
R13588 gnd.n6502 gnd.n6501 0.152939
R13589 gnd.n6503 gnd.n6502 0.152939
R13590 gnd.n6503 gnd.n558 0.152939
R13591 gnd.n6511 gnd.n558 0.152939
R13592 gnd.n6512 gnd.n6511 0.152939
R13593 gnd.n6513 gnd.n6512 0.152939
R13594 gnd.n6513 gnd.n552 0.152939
R13595 gnd.n6521 gnd.n552 0.152939
R13596 gnd.n6522 gnd.n6521 0.152939
R13597 gnd.n6523 gnd.n6522 0.152939
R13598 gnd.n6523 gnd.n546 0.152939
R13599 gnd.n6531 gnd.n546 0.152939
R13600 gnd.n6532 gnd.n6531 0.152939
R13601 gnd.n6533 gnd.n6532 0.152939
R13602 gnd.n6533 gnd.n540 0.152939
R13603 gnd.n6541 gnd.n540 0.152939
R13604 gnd.n6542 gnd.n6541 0.152939
R13605 gnd.n6543 gnd.n6542 0.152939
R13606 gnd.n6543 gnd.n534 0.152939
R13607 gnd.n6551 gnd.n534 0.152939
R13608 gnd.n6552 gnd.n6551 0.152939
R13609 gnd.n6553 gnd.n6552 0.152939
R13610 gnd.n6553 gnd.n528 0.152939
R13611 gnd.n6561 gnd.n528 0.152939
R13612 gnd.n6562 gnd.n6561 0.152939
R13613 gnd.n6564 gnd.n6562 0.152939
R13614 gnd.n6564 gnd.n6563 0.152939
R13615 gnd.n6563 gnd.n522 0.152939
R13616 gnd.n6573 gnd.n522 0.152939
R13617 gnd.n6574 gnd.n517 0.152939
R13618 gnd.n6582 gnd.n517 0.152939
R13619 gnd.n6583 gnd.n6582 0.152939
R13620 gnd.n6584 gnd.n6583 0.152939
R13621 gnd.n6584 gnd.n511 0.152939
R13622 gnd.n6592 gnd.n511 0.152939
R13623 gnd.n6593 gnd.n6592 0.152939
R13624 gnd.n6594 gnd.n6593 0.152939
R13625 gnd.n6594 gnd.n505 0.152939
R13626 gnd.n6602 gnd.n505 0.152939
R13627 gnd.n6603 gnd.n6602 0.152939
R13628 gnd.n6604 gnd.n6603 0.152939
R13629 gnd.n6604 gnd.n499 0.152939
R13630 gnd.n6612 gnd.n499 0.152939
R13631 gnd.n6613 gnd.n6612 0.152939
R13632 gnd.n6614 gnd.n6613 0.152939
R13633 gnd.n6614 gnd.n493 0.152939
R13634 gnd.n6622 gnd.n493 0.152939
R13635 gnd.n6623 gnd.n6622 0.152939
R13636 gnd.n6624 gnd.n6623 0.152939
R13637 gnd.n6624 gnd.n487 0.152939
R13638 gnd.n6632 gnd.n487 0.152939
R13639 gnd.n6633 gnd.n6632 0.152939
R13640 gnd.n6634 gnd.n6633 0.152939
R13641 gnd.n6634 gnd.n481 0.152939
R13642 gnd.n6642 gnd.n481 0.152939
R13643 gnd.n6643 gnd.n6642 0.152939
R13644 gnd.n6644 gnd.n6643 0.152939
R13645 gnd.n6644 gnd.n475 0.152939
R13646 gnd.n6652 gnd.n475 0.152939
R13647 gnd.n6653 gnd.n6652 0.152939
R13648 gnd.n6654 gnd.n6653 0.152939
R13649 gnd.n6654 gnd.n469 0.152939
R13650 gnd.n6662 gnd.n469 0.152939
R13651 gnd.n6663 gnd.n6662 0.152939
R13652 gnd.n6664 gnd.n6663 0.152939
R13653 gnd.n6664 gnd.n463 0.152939
R13654 gnd.n6672 gnd.n463 0.152939
R13655 gnd.n6673 gnd.n6672 0.152939
R13656 gnd.n6674 gnd.n6673 0.152939
R13657 gnd.n6674 gnd.n457 0.152939
R13658 gnd.n6682 gnd.n457 0.152939
R13659 gnd.n6683 gnd.n6682 0.152939
R13660 gnd.n6684 gnd.n6683 0.152939
R13661 gnd.n6684 gnd.n451 0.152939
R13662 gnd.n6692 gnd.n451 0.152939
R13663 gnd.n6693 gnd.n6692 0.152939
R13664 gnd.n6694 gnd.n6693 0.152939
R13665 gnd.n6694 gnd.n445 0.152939
R13666 gnd.n6702 gnd.n445 0.152939
R13667 gnd.n6703 gnd.n6702 0.152939
R13668 gnd.n6704 gnd.n6703 0.152939
R13669 gnd.n6704 gnd.n439 0.152939
R13670 gnd.n6712 gnd.n439 0.152939
R13671 gnd.n6713 gnd.n6712 0.152939
R13672 gnd.n6714 gnd.n6713 0.152939
R13673 gnd.n6714 gnd.n433 0.152939
R13674 gnd.n6722 gnd.n433 0.152939
R13675 gnd.n6723 gnd.n6722 0.152939
R13676 gnd.n6724 gnd.n6723 0.152939
R13677 gnd.n6724 gnd.n427 0.152939
R13678 gnd.n6732 gnd.n427 0.152939
R13679 gnd.n6733 gnd.n6732 0.152939
R13680 gnd.n6734 gnd.n6733 0.152939
R13681 gnd.n6734 gnd.n421 0.152939
R13682 gnd.n6742 gnd.n421 0.152939
R13683 gnd.n6743 gnd.n6742 0.152939
R13684 gnd.n6744 gnd.n6743 0.152939
R13685 gnd.n6744 gnd.n415 0.152939
R13686 gnd.n6752 gnd.n415 0.152939
R13687 gnd.n6753 gnd.n6752 0.152939
R13688 gnd.n6754 gnd.n6753 0.152939
R13689 gnd.n6754 gnd.n409 0.152939
R13690 gnd.n6762 gnd.n409 0.152939
R13691 gnd.n6763 gnd.n6762 0.152939
R13692 gnd.n6764 gnd.n6763 0.152939
R13693 gnd.n6764 gnd.n403 0.152939
R13694 gnd.n6772 gnd.n403 0.152939
R13695 gnd.n6773 gnd.n6772 0.152939
R13696 gnd.n6774 gnd.n6773 0.152939
R13697 gnd.n6774 gnd.n397 0.152939
R13698 gnd.n6783 gnd.n397 0.152939
R13699 gnd.n6784 gnd.n6783 0.152939
R13700 gnd.n6785 gnd.n6784 0.152939
R13701 gnd.n4298 gnd.n4294 0.152939
R13702 gnd.n4299 gnd.n4298 0.152939
R13703 gnd.n4300 gnd.n4299 0.152939
R13704 gnd.n4300 gnd.n2064 0.152939
R13705 gnd.n4306 gnd.n2064 0.152939
R13706 gnd.n4307 gnd.n4306 0.152939
R13707 gnd.n4308 gnd.n4307 0.152939
R13708 gnd.n4309 gnd.n4308 0.152939
R13709 gnd.n4310 gnd.n4309 0.152939
R13710 gnd.n4310 gnd.n2046 0.152939
R13711 gnd.n4601 gnd.n2046 0.152939
R13712 gnd.n4602 gnd.n4601 0.152939
R13713 gnd.n4603 gnd.n4602 0.152939
R13714 gnd.n4603 gnd.n2042 0.152939
R13715 gnd.n4609 gnd.n2042 0.152939
R13716 gnd.n4610 gnd.n4609 0.152939
R13717 gnd.n4611 gnd.n4610 0.152939
R13718 gnd.n4612 gnd.n4611 0.152939
R13719 gnd.n4613 gnd.n4612 0.152939
R13720 gnd.n4614 gnd.n4613 0.152939
R13721 gnd.n4614 gnd.n2012 0.152939
R13722 gnd.n4637 gnd.n2012 0.152939
R13723 gnd.n4638 gnd.n4637 0.152939
R13724 gnd.n4639 gnd.n4638 0.152939
R13725 gnd.n4639 gnd.n1996 0.152939
R13726 gnd.n4670 gnd.n1996 0.152939
R13727 gnd.n4671 gnd.n4670 0.152939
R13728 gnd.n4672 gnd.n4671 0.152939
R13729 gnd.n4673 gnd.n4672 0.152939
R13730 gnd.n4674 gnd.n4673 0.152939
R13731 gnd.n4676 gnd.n4674 0.152939
R13732 gnd.n4676 gnd.n4675 0.152939
R13733 gnd.n4675 gnd.n1119 0.152939
R13734 gnd.n1120 gnd.n1119 0.152939
R13735 gnd.n1121 gnd.n1120 0.152939
R13736 gnd.n4866 gnd.n1121 0.152939
R13737 gnd.n4867 gnd.n4866 0.152939
R13738 gnd.n4868 gnd.n4867 0.152939
R13739 gnd.n4868 gnd.n1885 0.152939
R13740 gnd.n4895 gnd.n1885 0.152939
R13741 gnd.n4896 gnd.n4895 0.152939
R13742 gnd.n4897 gnd.n4896 0.152939
R13743 gnd.n4898 gnd.n4897 0.152939
R13744 gnd.n4899 gnd.n4898 0.152939
R13745 gnd.n4901 gnd.n4899 0.152939
R13746 gnd.n4902 gnd.n4901 0.152939
R13747 gnd.n4902 gnd.n1847 0.152939
R13748 gnd.n4953 gnd.n1847 0.152939
R13749 gnd.n4954 gnd.n4953 0.152939
R13750 gnd.n4955 gnd.n4954 0.152939
R13751 gnd.n4955 gnd.n1829 0.152939
R13752 gnd.n4979 gnd.n1829 0.152939
R13753 gnd.n4980 gnd.n4979 0.152939
R13754 gnd.n4981 gnd.n4980 0.152939
R13755 gnd.n4982 gnd.n4981 0.152939
R13756 gnd.n4982 gnd.n1805 0.152939
R13757 gnd.n5018 gnd.n1805 0.152939
R13758 gnd.n5019 gnd.n5018 0.152939
R13759 gnd.n5020 gnd.n5019 0.152939
R13760 gnd.n5021 gnd.n5020 0.152939
R13761 gnd.n5022 gnd.n5021 0.152939
R13762 gnd.n5024 gnd.n5022 0.152939
R13763 gnd.n5025 gnd.n5024 0.152939
R13764 gnd.n5025 gnd.n1766 0.152939
R13765 gnd.n5076 gnd.n1766 0.152939
R13766 gnd.n5077 gnd.n5076 0.152939
R13767 gnd.n5078 gnd.n5077 0.152939
R13768 gnd.n5078 gnd.n1747 0.152939
R13769 gnd.n5101 gnd.n1747 0.152939
R13770 gnd.n5102 gnd.n5101 0.152939
R13771 gnd.n5103 gnd.n5102 0.152939
R13772 gnd.n5104 gnd.n5103 0.152939
R13773 gnd.n5104 gnd.n1722 0.152939
R13774 gnd.n5139 gnd.n1722 0.152939
R13775 gnd.n5140 gnd.n5139 0.152939
R13776 gnd.n5141 gnd.n5140 0.152939
R13777 gnd.n5142 gnd.n5141 0.152939
R13778 gnd.n5143 gnd.n5142 0.152939
R13779 gnd.n5144 gnd.n5143 0.152939
R13780 gnd.n5144 gnd.n1688 0.152939
R13781 gnd.n5185 gnd.n1688 0.152939
R13782 gnd.n5186 gnd.n5185 0.152939
R13783 gnd.n5187 gnd.n5186 0.152939
R13784 gnd.n5188 gnd.n5187 0.152939
R13785 gnd.n5188 gnd.n1660 0.152939
R13786 gnd.n5220 gnd.n1660 0.152939
R13787 gnd.n5221 gnd.n5220 0.152939
R13788 gnd.n5222 gnd.n5221 0.152939
R13789 gnd.n5222 gnd.n1631 0.152939
R13790 gnd.n5257 gnd.n1631 0.152939
R13791 gnd.n5258 gnd.n5257 0.152939
R13792 gnd.n5259 gnd.n5258 0.152939
R13793 gnd.n5260 gnd.n5259 0.152939
R13794 gnd.n5260 gnd.n1531 0.152939
R13795 gnd.n5407 gnd.n1531 0.152939
R13796 gnd.n5408 gnd.n5407 0.152939
R13797 gnd.n5409 gnd.n5408 0.152939
R13798 gnd.n5409 gnd.n1518 0.152939
R13799 gnd.n5423 gnd.n1518 0.152939
R13800 gnd.n5424 gnd.n5423 0.152939
R13801 gnd.n5425 gnd.n5424 0.152939
R13802 gnd.n5427 gnd.n5425 0.152939
R13803 gnd.n5427 gnd.n5426 0.152939
R13804 gnd.n5426 gnd.n1505 0.152939
R13805 gnd.n5444 gnd.n1505 0.152939
R13806 gnd.n5445 gnd.n5444 0.152939
R13807 gnd.n5446 gnd.n5445 0.152939
R13808 gnd.n5447 gnd.n5446 0.152939
R13809 gnd.n5448 gnd.n5447 0.152939
R13810 gnd.n5450 gnd.n5448 0.152939
R13811 gnd.n5451 gnd.n5450 0.152939
R13812 gnd.n5451 gnd.n1470 0.152939
R13813 gnd.n5529 gnd.n1470 0.152939
R13814 gnd.n5530 gnd.n5529 0.152939
R13815 gnd.n5531 gnd.n5530 0.152939
R13816 gnd.n5531 gnd.n1466 0.152939
R13817 gnd.n5537 gnd.n1466 0.152939
R13818 gnd.n5538 gnd.n5537 0.152939
R13819 gnd.n5539 gnd.n5538 0.152939
R13820 gnd.n5539 gnd.n1462 0.152939
R13821 gnd.n5545 gnd.n1462 0.152939
R13822 gnd.n5546 gnd.n5545 0.152939
R13823 gnd.n5547 gnd.n5546 0.152939
R13824 gnd.n5549 gnd.n5547 0.152939
R13825 gnd.n5549 gnd.n5548 0.152939
R13826 gnd.n5548 gnd.n392 0.152939
R13827 gnd.n393 gnd.n392 0.152939
R13828 gnd.n394 gnd.n393 0.152939
R13829 gnd.n6251 gnd.n714 0.152939
R13830 gnd.n719 gnd.n714 0.152939
R13831 gnd.n720 gnd.n719 0.152939
R13832 gnd.n721 gnd.n720 0.152939
R13833 gnd.n726 gnd.n721 0.152939
R13834 gnd.n727 gnd.n726 0.152939
R13835 gnd.n728 gnd.n727 0.152939
R13836 gnd.n729 gnd.n728 0.152939
R13837 gnd.n734 gnd.n729 0.152939
R13838 gnd.n735 gnd.n734 0.152939
R13839 gnd.n736 gnd.n735 0.152939
R13840 gnd.n737 gnd.n736 0.152939
R13841 gnd.n742 gnd.n737 0.152939
R13842 gnd.n743 gnd.n742 0.152939
R13843 gnd.n744 gnd.n743 0.152939
R13844 gnd.n745 gnd.n744 0.152939
R13845 gnd.n750 gnd.n745 0.152939
R13846 gnd.n751 gnd.n750 0.152939
R13847 gnd.n752 gnd.n751 0.152939
R13848 gnd.n753 gnd.n752 0.152939
R13849 gnd.n758 gnd.n753 0.152939
R13850 gnd.n759 gnd.n758 0.152939
R13851 gnd.n760 gnd.n759 0.152939
R13852 gnd.n761 gnd.n760 0.152939
R13853 gnd.n766 gnd.n761 0.152939
R13854 gnd.n767 gnd.n766 0.152939
R13855 gnd.n768 gnd.n767 0.152939
R13856 gnd.n769 gnd.n768 0.152939
R13857 gnd.n774 gnd.n769 0.152939
R13858 gnd.n775 gnd.n774 0.152939
R13859 gnd.n776 gnd.n775 0.152939
R13860 gnd.n777 gnd.n776 0.152939
R13861 gnd.n782 gnd.n777 0.152939
R13862 gnd.n783 gnd.n782 0.152939
R13863 gnd.n784 gnd.n783 0.152939
R13864 gnd.n785 gnd.n784 0.152939
R13865 gnd.n790 gnd.n785 0.152939
R13866 gnd.n791 gnd.n790 0.152939
R13867 gnd.n792 gnd.n791 0.152939
R13868 gnd.n793 gnd.n792 0.152939
R13869 gnd.n798 gnd.n793 0.152939
R13870 gnd.n799 gnd.n798 0.152939
R13871 gnd.n800 gnd.n799 0.152939
R13872 gnd.n801 gnd.n800 0.152939
R13873 gnd.n806 gnd.n801 0.152939
R13874 gnd.n807 gnd.n806 0.152939
R13875 gnd.n808 gnd.n807 0.152939
R13876 gnd.n809 gnd.n808 0.152939
R13877 gnd.n814 gnd.n809 0.152939
R13878 gnd.n815 gnd.n814 0.152939
R13879 gnd.n816 gnd.n815 0.152939
R13880 gnd.n817 gnd.n816 0.152939
R13881 gnd.n822 gnd.n817 0.152939
R13882 gnd.n823 gnd.n822 0.152939
R13883 gnd.n824 gnd.n823 0.152939
R13884 gnd.n825 gnd.n824 0.152939
R13885 gnd.n830 gnd.n825 0.152939
R13886 gnd.n831 gnd.n830 0.152939
R13887 gnd.n832 gnd.n831 0.152939
R13888 gnd.n833 gnd.n832 0.152939
R13889 gnd.n838 gnd.n833 0.152939
R13890 gnd.n839 gnd.n838 0.152939
R13891 gnd.n840 gnd.n839 0.152939
R13892 gnd.n841 gnd.n840 0.152939
R13893 gnd.n846 gnd.n841 0.152939
R13894 gnd.n847 gnd.n846 0.152939
R13895 gnd.n848 gnd.n847 0.152939
R13896 gnd.n849 gnd.n848 0.152939
R13897 gnd.n854 gnd.n849 0.152939
R13898 gnd.n855 gnd.n854 0.152939
R13899 gnd.n856 gnd.n855 0.152939
R13900 gnd.n857 gnd.n856 0.152939
R13901 gnd.n862 gnd.n857 0.152939
R13902 gnd.n863 gnd.n862 0.152939
R13903 gnd.n864 gnd.n863 0.152939
R13904 gnd.n865 gnd.n864 0.152939
R13905 gnd.n870 gnd.n865 0.152939
R13906 gnd.n871 gnd.n870 0.152939
R13907 gnd.n872 gnd.n871 0.152939
R13908 gnd.n873 gnd.n872 0.152939
R13909 gnd.n878 gnd.n873 0.152939
R13910 gnd.n879 gnd.n878 0.152939
R13911 gnd.n880 gnd.n879 0.152939
R13912 gnd.n881 gnd.n880 0.152939
R13913 gnd.n4645 gnd.n2005 0.152939
R13914 gnd.n4646 gnd.n4645 0.152939
R13915 gnd.n4664 gnd.n4646 0.152939
R13916 gnd.n4664 gnd.n4663 0.152939
R13917 gnd.n4663 gnd.n4662 0.152939
R13918 gnd.n4662 gnd.n4647 0.152939
R13919 gnd.n4658 gnd.n4647 0.152939
R13920 gnd.n4658 gnd.n4657 0.152939
R13921 gnd.n4657 gnd.n4656 0.152939
R13922 gnd.n4656 gnd.n4651 0.152939
R13923 gnd.n4651 gnd.n1130 0.152939
R13924 gnd.n5888 gnd.n1130 0.152939
R13925 gnd.n5888 gnd.n5887 0.152939
R13926 gnd.n5887 gnd.n5886 0.152939
R13927 gnd.n5886 gnd.n1131 0.152939
R13928 gnd.n5882 gnd.n1131 0.152939
R13929 gnd.n5882 gnd.n5881 0.152939
R13930 gnd.n5881 gnd.n5880 0.152939
R13931 gnd.n5880 gnd.n1136 0.152939
R13932 gnd.n5876 gnd.n1136 0.152939
R13933 gnd.n5876 gnd.n5875 0.152939
R13934 gnd.n5875 gnd.n5874 0.152939
R13935 gnd.n5874 gnd.n1141 0.152939
R13936 gnd.n5870 gnd.n1141 0.152939
R13937 gnd.n5870 gnd.n5869 0.152939
R13938 gnd.n5869 gnd.n5868 0.152939
R13939 gnd.n5868 gnd.n1146 0.152939
R13940 gnd.n5864 gnd.n1146 0.152939
R13941 gnd.n5864 gnd.n5863 0.152939
R13942 gnd.n5863 gnd.n5862 0.152939
R13943 gnd.n5862 gnd.n1151 0.152939
R13944 gnd.n5858 gnd.n1151 0.152939
R13945 gnd.n5858 gnd.n5857 0.152939
R13946 gnd.n5857 gnd.n5856 0.152939
R13947 gnd.n5856 gnd.n1156 0.152939
R13948 gnd.n5852 gnd.n1156 0.152939
R13949 gnd.n5852 gnd.n5851 0.152939
R13950 gnd.n5851 gnd.n5850 0.152939
R13951 gnd.n5850 gnd.n1161 0.152939
R13952 gnd.n5846 gnd.n1161 0.152939
R13953 gnd.n5846 gnd.n5845 0.152939
R13954 gnd.n5845 gnd.n5844 0.152939
R13955 gnd.n5844 gnd.n1166 0.152939
R13956 gnd.n5840 gnd.n1166 0.152939
R13957 gnd.n5840 gnd.n5839 0.152939
R13958 gnd.n5839 gnd.n5838 0.152939
R13959 gnd.n5838 gnd.n1171 0.152939
R13960 gnd.n5834 gnd.n1171 0.152939
R13961 gnd.n5834 gnd.n5833 0.152939
R13962 gnd.n5833 gnd.n5832 0.152939
R13963 gnd.n5832 gnd.n1176 0.152939
R13964 gnd.n5828 gnd.n1176 0.152939
R13965 gnd.n5828 gnd.n5827 0.152939
R13966 gnd.n5827 gnd.n5826 0.152939
R13967 gnd.n5826 gnd.n1181 0.152939
R13968 gnd.n5822 gnd.n1181 0.152939
R13969 gnd.n5822 gnd.n5821 0.152939
R13970 gnd.n5821 gnd.n5820 0.152939
R13971 gnd.n5820 gnd.n1186 0.152939
R13972 gnd.n5816 gnd.n1186 0.152939
R13973 gnd.n5816 gnd.n5815 0.152939
R13974 gnd.n5815 gnd.n5814 0.152939
R13975 gnd.n5814 gnd.n1191 0.152939
R13976 gnd.n5810 gnd.n1191 0.152939
R13977 gnd.n5810 gnd.n5809 0.152939
R13978 gnd.n5809 gnd.n5808 0.152939
R13979 gnd.n5808 gnd.n1196 0.152939
R13980 gnd.n5804 gnd.n1196 0.152939
R13981 gnd.n5804 gnd.n5803 0.152939
R13982 gnd.n5803 gnd.n5802 0.152939
R13983 gnd.n5802 gnd.n1201 0.152939
R13984 gnd.n5798 gnd.n1201 0.152939
R13985 gnd.n5798 gnd.n5797 0.152939
R13986 gnd.n5797 gnd.n5796 0.152939
R13987 gnd.n5796 gnd.n1206 0.152939
R13988 gnd.n5792 gnd.n1206 0.152939
R13989 gnd.n5792 gnd.n5791 0.152939
R13990 gnd.n5791 gnd.n5790 0.152939
R13991 gnd.n5790 gnd.n1211 0.152939
R13992 gnd.n5786 gnd.n1211 0.152939
R13993 gnd.n5786 gnd.n5785 0.152939
R13994 gnd.n5785 gnd.n5784 0.152939
R13995 gnd.n4212 gnd.n4211 0.152939
R13996 gnd.n4211 gnd.n4210 0.152939
R13997 gnd.n4210 gnd.n4199 0.152939
R13998 gnd.n4206 gnd.n4199 0.152939
R13999 gnd.n4206 gnd.n4205 0.152939
R14000 gnd.n4205 gnd.n4204 0.152939
R14001 gnd.n4204 gnd.n2073 0.152939
R14002 gnd.n4266 gnd.n2073 0.152939
R14003 gnd.n4267 gnd.n4266 0.152939
R14004 gnd.n4268 gnd.n4267 0.152939
R14005 gnd.n4268 gnd.n2069 0.152939
R14006 gnd.n4287 gnd.n2069 0.152939
R14007 gnd.n4287 gnd.n4286 0.152939
R14008 gnd.n4286 gnd.n4285 0.152939
R14009 gnd.n4285 gnd.n2058 0.152939
R14010 gnd.n4319 gnd.n2058 0.152939
R14011 gnd.n4320 gnd.n4319 0.152939
R14012 gnd.n4321 gnd.n4320 0.152939
R14013 gnd.n4321 gnd.n2052 0.152939
R14014 gnd.n4593 gnd.n2052 0.152939
R14015 gnd.n4593 gnd.n4592 0.152939
R14016 gnd.n4592 gnd.n4591 0.152939
R14017 gnd.n4591 gnd.n2053 0.152939
R14018 gnd.n4587 gnd.n2053 0.152939
R14019 gnd.n4587 gnd.n4586 0.152939
R14020 gnd.n4586 gnd.n2032 0.152939
R14021 gnd.n4341 gnd.n4340 0.152939
R14022 gnd.n4358 gnd.n4340 0.152939
R14023 gnd.n4359 gnd.n4358 0.152939
R14024 gnd.n4360 gnd.n4359 0.152939
R14025 gnd.n4360 gnd.n4336 0.152939
R14026 gnd.n4479 gnd.n4336 0.152939
R14027 gnd.n4349 gnd.n4348 0.152939
R14028 gnd.n4348 gnd.n4347 0.152939
R14029 gnd.n4347 gnd.n4343 0.152939
R14030 gnd.n4343 gnd.n1987 0.152939
R14031 gnd.n4687 gnd.n1987 0.152939
R14032 gnd.n4688 gnd.n4687 0.152939
R14033 gnd.n4689 gnd.n4688 0.152939
R14034 gnd.n4689 gnd.n1983 0.152939
R14035 gnd.n4695 gnd.n1983 0.152939
R14036 gnd.n4696 gnd.n4695 0.152939
R14037 gnd.n4838 gnd.n4696 0.152939
R14038 gnd.n4838 gnd.n4837 0.152939
R14039 gnd.n4837 gnd.n4836 0.152939
R14040 gnd.n4836 gnd.n4697 0.152939
R14041 gnd.n4832 gnd.n4697 0.152939
R14042 gnd.n4832 gnd.n4831 0.152939
R14043 gnd.n4831 gnd.n4830 0.152939
R14044 gnd.n4830 gnd.n4700 0.152939
R14045 gnd.n4826 gnd.n4700 0.152939
R14046 gnd.n4826 gnd.n4825 0.152939
R14047 gnd.n4825 gnd.n4824 0.152939
R14048 gnd.n4824 gnd.n4703 0.152939
R14049 gnd.n4820 gnd.n4703 0.152939
R14050 gnd.n4820 gnd.n4819 0.152939
R14051 gnd.n4819 gnd.n4818 0.152939
R14052 gnd.n4818 gnd.n4709 0.152939
R14053 gnd.n4814 gnd.n4709 0.152939
R14054 gnd.n4814 gnd.n4813 0.152939
R14055 gnd.n4813 gnd.n4812 0.152939
R14056 gnd.n4812 gnd.n4713 0.152939
R14057 gnd.n4808 gnd.n4713 0.152939
R14058 gnd.n4808 gnd.n4807 0.152939
R14059 gnd.n4807 gnd.n4806 0.152939
R14060 gnd.n4806 gnd.n4717 0.152939
R14061 gnd.n4802 gnd.n4717 0.152939
R14062 gnd.n4802 gnd.n4801 0.152939
R14063 gnd.n4801 gnd.n4800 0.152939
R14064 gnd.n4800 gnd.n4720 0.152939
R14065 gnd.n4796 gnd.n4720 0.152939
R14066 gnd.n4796 gnd.n4795 0.152939
R14067 gnd.n4795 gnd.n4794 0.152939
R14068 gnd.n4794 gnd.n4726 0.152939
R14069 gnd.n4790 gnd.n4726 0.152939
R14070 gnd.n4790 gnd.n4789 0.152939
R14071 gnd.n4789 gnd.n4788 0.152939
R14072 gnd.n4788 gnd.n4729 0.152939
R14073 gnd.n4784 gnd.n4729 0.152939
R14074 gnd.n4784 gnd.n4783 0.152939
R14075 gnd.n4783 gnd.n4782 0.152939
R14076 gnd.n4782 gnd.n4733 0.152939
R14077 gnd.n4778 gnd.n4733 0.152939
R14078 gnd.n4778 gnd.n4777 0.152939
R14079 gnd.n4777 gnd.n4776 0.152939
R14080 gnd.n4776 gnd.n4738 0.152939
R14081 gnd.n4772 gnd.n4738 0.152939
R14082 gnd.n4772 gnd.n4771 0.152939
R14083 gnd.n4771 gnd.n4770 0.152939
R14084 gnd.n4770 gnd.n4742 0.152939
R14085 gnd.n4766 gnd.n4742 0.152939
R14086 gnd.n4766 gnd.n4765 0.152939
R14087 gnd.n4765 gnd.n4764 0.152939
R14088 gnd.n4764 gnd.n4747 0.152939
R14089 gnd.n4760 gnd.n4747 0.152939
R14090 gnd.n4760 gnd.n4759 0.152939
R14091 gnd.n4759 gnd.n4758 0.152939
R14092 gnd.n4758 gnd.n4752 0.152939
R14093 gnd.n4754 gnd.n4752 0.152939
R14094 gnd.n4754 gnd.n1622 0.152939
R14095 gnd.n5267 gnd.n1622 0.152939
R14096 gnd.n5268 gnd.n5267 0.152939
R14097 gnd.n5270 gnd.n5268 0.152939
R14098 gnd.n5270 gnd.n5269 0.152939
R14099 gnd.n5269 gnd.n1523 0.152939
R14100 gnd.n5415 gnd.n1523 0.152939
R14101 gnd.n5416 gnd.n5415 0.152939
R14102 gnd.n5417 gnd.n5416 0.152939
R14103 gnd.n5417 gnd.n1511 0.152939
R14104 gnd.n5434 gnd.n1511 0.152939
R14105 gnd.n5435 gnd.n5434 0.152939
R14106 gnd.n5436 gnd.n5435 0.152939
R14107 gnd.n5436 gnd.n1225 0.152939
R14108 gnd.n5778 gnd.n1225 0.152939
R14109 gnd.n5777 gnd.n1226 0.152939
R14110 gnd.n5773 gnd.n1226 0.152939
R14111 gnd.n5773 gnd.n5772 0.152939
R14112 gnd.n5772 gnd.n5771 0.152939
R14113 gnd.n5771 gnd.n1230 0.152939
R14114 gnd.n5767 gnd.n1230 0.152939
R14115 gnd.n5522 gnd.n5467 0.152939
R14116 gnd.n5522 gnd.n5521 0.152939
R14117 gnd.n5521 gnd.n5520 0.152939
R14118 gnd.n5520 gnd.n5468 0.152939
R14119 gnd.n5516 gnd.n5468 0.152939
R14120 gnd.n5516 gnd.n5515 0.152939
R14121 gnd.n5515 gnd.n5514 0.152939
R14122 gnd.n5514 gnd.n5472 0.152939
R14123 gnd.n5510 gnd.n5472 0.152939
R14124 gnd.n5510 gnd.n5509 0.152939
R14125 gnd.n5509 gnd.n5508 0.152939
R14126 gnd.n5508 gnd.n5476 0.152939
R14127 gnd.n5504 gnd.n5476 0.152939
R14128 gnd.n5504 gnd.n367 0.152939
R14129 gnd.n6820 gnd.n367 0.152939
R14130 gnd.n6821 gnd.n6820 0.152939
R14131 gnd.n6823 gnd.n6821 0.152939
R14132 gnd.n6823 gnd.n6822 0.152939
R14133 gnd.n6822 gnd.n340 0.152939
R14134 gnd.n6854 gnd.n340 0.152939
R14135 gnd.n6855 gnd.n6854 0.152939
R14136 gnd.n6862 gnd.n6855 0.152939
R14137 gnd.n6862 gnd.n6861 0.152939
R14138 gnd.n6861 gnd.n6860 0.152939
R14139 gnd.n6860 gnd.n6856 0.152939
R14140 gnd.n6856 gnd.n79 0.152939
R14141 gnd.n4480 gnd.n4479 0.128549
R14142 gnd.n5767 gnd.n5766 0.128549
R14143 gnd.n6847 gnd.n326 0.0785577
R14144 gnd.n112 gnd.n111 0.0785577
R14145 gnd.n4256 gnd.n2080 0.0785577
R14146 gnd.n4154 gnd.n2126 0.0785577
R14147 gnd.n3120 gnd.n3119 0.0767195
R14148 gnd.n3119 gnd.n3118 0.0767195
R14149 gnd.n7268 gnd.n7267 0.0695946
R14150 gnd.n4198 gnd.n4197 0.0695946
R14151 gnd.n4212 gnd.n4198 0.0695946
R14152 gnd.n7268 gnd.n79 0.0695946
R14153 gnd.n4577 gnd.n4480 0.063
R14154 gnd.n5766 gnd.n1235 0.063
R14155 gnd.n1403 gnd.n1235 0.0477147
R14156 gnd.n7063 gnd.n7062 0.0477147
R14157 gnd.n3686 gnd.n2285 0.0477147
R14158 gnd.n3918 gnd.n2241 0.0477147
R14159 gnd.n4578 gnd.n4577 0.0477147
R14160 gnd.n2883 gnd.n2771 0.0442063
R14161 gnd.n2884 gnd.n2883 0.0442063
R14162 gnd.n2885 gnd.n2884 0.0442063
R14163 gnd.n2885 gnd.n2760 0.0442063
R14164 gnd.n2899 gnd.n2760 0.0442063
R14165 gnd.n2900 gnd.n2899 0.0442063
R14166 gnd.n2901 gnd.n2900 0.0442063
R14167 gnd.n2901 gnd.n2747 0.0442063
R14168 gnd.n2945 gnd.n2747 0.0442063
R14169 gnd.n2946 gnd.n2945 0.0442063
R14170 gnd.n1404 gnd.n1403 0.0344674
R14171 gnd.n1405 gnd.n1404 0.0344674
R14172 gnd.n5479 gnd.n1405 0.0344674
R14173 gnd.n5479 gnd.n1427 0.0344674
R14174 gnd.n1428 gnd.n1427 0.0344674
R14175 gnd.n1429 gnd.n1428 0.0344674
R14176 gnd.n5488 gnd.n1429 0.0344674
R14177 gnd.n5488 gnd.n1448 0.0344674
R14178 gnd.n1449 gnd.n1448 0.0344674
R14179 gnd.n1450 gnd.n1449 0.0344674
R14180 gnd.n5498 gnd.n1450 0.0344674
R14181 gnd.n5499 gnd.n5498 0.0344674
R14182 gnd.n5499 gnd.n386 0.0344674
R14183 gnd.n387 gnd.n386 0.0344674
R14184 gnd.n6798 gnd.n387 0.0344674
R14185 gnd.n6799 gnd.n6798 0.0344674
R14186 gnd.n6799 gnd.n361 0.0344674
R14187 gnd.n361 gnd.n358 0.0344674
R14188 gnd.n359 gnd.n358 0.0344674
R14189 gnd.n6833 gnd.n359 0.0344674
R14190 gnd.n6834 gnd.n6833 0.0344674
R14191 gnd.n6834 gnd.n333 0.0344674
R14192 gnd.n6871 gnd.n333 0.0344674
R14193 gnd.n6871 gnd.n316 0.0344674
R14194 gnd.n6888 gnd.n316 0.0344674
R14195 gnd.n6889 gnd.n6888 0.0344674
R14196 gnd.n6889 gnd.n310 0.0344674
R14197 gnd.n6897 gnd.n310 0.0344674
R14198 gnd.n6898 gnd.n6897 0.0344674
R14199 gnd.n6898 gnd.n101 0.0344674
R14200 gnd.n102 gnd.n101 0.0344674
R14201 gnd.n103 gnd.n102 0.0344674
R14202 gnd.n6905 gnd.n103 0.0344674
R14203 gnd.n6905 gnd.n121 0.0344674
R14204 gnd.n122 gnd.n121 0.0344674
R14205 gnd.n123 gnd.n122 0.0344674
R14206 gnd.n6912 gnd.n123 0.0344674
R14207 gnd.n6912 gnd.n139 0.0344674
R14208 gnd.n140 gnd.n139 0.0344674
R14209 gnd.n141 gnd.n140 0.0344674
R14210 gnd.n6919 gnd.n141 0.0344674
R14211 gnd.n6919 gnd.n159 0.0344674
R14212 gnd.n160 gnd.n159 0.0344674
R14213 gnd.n161 gnd.n160 0.0344674
R14214 gnd.n7045 gnd.n161 0.0344674
R14215 gnd.n7045 gnd.n177 0.0344674
R14216 gnd.n178 gnd.n177 0.0344674
R14217 gnd.n179 gnd.n178 0.0344674
R14218 gnd.n7052 gnd.n179 0.0344674
R14219 gnd.n7052 gnd.n197 0.0344674
R14220 gnd.n198 gnd.n197 0.0344674
R14221 gnd.n199 gnd.n198 0.0344674
R14222 gnd.n7062 gnd.n199 0.0344674
R14223 gnd.n2948 gnd.n2681 0.0344674
R14224 gnd.n2241 gnd.n2240 0.0344674
R14225 gnd.n4043 gnd.n2240 0.0344674
R14226 gnd.n4044 gnd.n4043 0.0344674
R14227 gnd.n4044 gnd.n2224 0.0344674
R14228 gnd.n2224 gnd.n2222 0.0344674
R14229 gnd.n4063 gnd.n2222 0.0344674
R14230 gnd.n4064 gnd.n4063 0.0344674
R14231 gnd.n4064 gnd.n2206 0.0344674
R14232 gnd.n2206 gnd.n2204 0.0344674
R14233 gnd.n4083 gnd.n2204 0.0344674
R14234 gnd.n4084 gnd.n4083 0.0344674
R14235 gnd.n4084 gnd.n2188 0.0344674
R14236 gnd.n2188 gnd.n2185 0.0344674
R14237 gnd.n2186 gnd.n2185 0.0344674
R14238 gnd.n4105 gnd.n2186 0.0344674
R14239 gnd.n4106 gnd.n4105 0.0344674
R14240 gnd.n4106 gnd.n2162 0.0344674
R14241 gnd.n2162 gnd.n2159 0.0344674
R14242 gnd.n2160 gnd.n2159 0.0344674
R14243 gnd.n4140 gnd.n2160 0.0344674
R14244 gnd.n4141 gnd.n4140 0.0344674
R14245 gnd.n4141 gnd.n2137 0.0344674
R14246 gnd.n2137 gnd.n2134 0.0344674
R14247 gnd.n2135 gnd.n2134 0.0344674
R14248 gnd.n4175 gnd.n2135 0.0344674
R14249 gnd.n4176 gnd.n4175 0.0344674
R14250 gnd.n4176 gnd.n2111 0.0344674
R14251 gnd.n2111 gnd.n2109 0.0344674
R14252 gnd.n4220 gnd.n2109 0.0344674
R14253 gnd.n4221 gnd.n4220 0.0344674
R14254 gnd.n4221 gnd.n2094 0.0344674
R14255 gnd.n2094 gnd.n2090 0.0344674
R14256 gnd.n2091 gnd.n2090 0.0344674
R14257 gnd.n2092 gnd.n2091 0.0344674
R14258 gnd.n4244 gnd.n2092 0.0344674
R14259 gnd.n4245 gnd.n4244 0.0344674
R14260 gnd.n4245 gnd.n2071 0.0344674
R14261 gnd.n2071 gnd.n902 0.0344674
R14262 gnd.n903 gnd.n902 0.0344674
R14263 gnd.n904 gnd.n903 0.0344674
R14264 gnd.n4277 gnd.n904 0.0344674
R14265 gnd.n4277 gnd.n923 0.0344674
R14266 gnd.n924 gnd.n923 0.0344674
R14267 gnd.n925 gnd.n924 0.0344674
R14268 gnd.n2056 gnd.n925 0.0344674
R14269 gnd.n2056 gnd.n942 0.0344674
R14270 gnd.n943 gnd.n942 0.0344674
R14271 gnd.n944 gnd.n943 0.0344674
R14272 gnd.n4330 gnd.n944 0.0344674
R14273 gnd.n4330 gnd.n963 0.0344674
R14274 gnd.n964 gnd.n963 0.0344674
R14275 gnd.n965 gnd.n964 0.0344674
R14276 gnd.n4578 gnd.n965 0.0344674
R14277 gnd.n4475 gnd.n4335 0.0344674
R14278 gnd.n5765 gnd.n5764 0.0344674
R14279 gnd.n4629 gnd.n4628 0.029712
R14280 gnd.n5466 gnd.n5465 0.029712
R14281 gnd.n2968 gnd.n2967 0.0269946
R14282 gnd.n2970 gnd.n2969 0.0269946
R14283 gnd.n2676 gnd.n2674 0.0269946
R14284 gnd.n2980 gnd.n2978 0.0269946
R14285 gnd.n2979 gnd.n2655 0.0269946
R14286 gnd.n2999 gnd.n2998 0.0269946
R14287 gnd.n3001 gnd.n3000 0.0269946
R14288 gnd.n2650 gnd.n2649 0.0269946
R14289 gnd.n3011 gnd.n2645 0.0269946
R14290 gnd.n3010 gnd.n2647 0.0269946
R14291 gnd.n2646 gnd.n2628 0.0269946
R14292 gnd.n3031 gnd.n2629 0.0269946
R14293 gnd.n3030 gnd.n2630 0.0269946
R14294 gnd.n3064 gnd.n2605 0.0269946
R14295 gnd.n3066 gnd.n3065 0.0269946
R14296 gnd.n3067 gnd.n2552 0.0269946
R14297 gnd.n2600 gnd.n2553 0.0269946
R14298 gnd.n2602 gnd.n2554 0.0269946
R14299 gnd.n3077 gnd.n3076 0.0269946
R14300 gnd.n3079 gnd.n3078 0.0269946
R14301 gnd.n3080 gnd.n2574 0.0269946
R14302 gnd.n3082 gnd.n2575 0.0269946
R14303 gnd.n3085 gnd.n2576 0.0269946
R14304 gnd.n3088 gnd.n3087 0.0269946
R14305 gnd.n3090 gnd.n3089 0.0269946
R14306 gnd.n3155 gnd.n2459 0.0269946
R14307 gnd.n3157 gnd.n3156 0.0269946
R14308 gnd.n3166 gnd.n2452 0.0269946
R14309 gnd.n3168 gnd.n3167 0.0269946
R14310 gnd.n3169 gnd.n2450 0.0269946
R14311 gnd.n3176 gnd.n3172 0.0269946
R14312 gnd.n3175 gnd.n3174 0.0269946
R14313 gnd.n3173 gnd.n2429 0.0269946
R14314 gnd.n3198 gnd.n2430 0.0269946
R14315 gnd.n3197 gnd.n2431 0.0269946
R14316 gnd.n3240 gnd.n2404 0.0269946
R14317 gnd.n3242 gnd.n3241 0.0269946
R14318 gnd.n3251 gnd.n2397 0.0269946
R14319 gnd.n3253 gnd.n3252 0.0269946
R14320 gnd.n3254 gnd.n2395 0.0269946
R14321 gnd.n3261 gnd.n3257 0.0269946
R14322 gnd.n3260 gnd.n3259 0.0269946
R14323 gnd.n3258 gnd.n2374 0.0269946
R14324 gnd.n3283 gnd.n2375 0.0269946
R14325 gnd.n3282 gnd.n2376 0.0269946
R14326 gnd.n3329 gnd.n2350 0.0269946
R14327 gnd.n3331 gnd.n3330 0.0269946
R14328 gnd.n3340 gnd.n2343 0.0269946
R14329 gnd.n3599 gnd.n2341 0.0269946
R14330 gnd.n3604 gnd.n3602 0.0269946
R14331 gnd.n3603 gnd.n2322 0.0269946
R14332 gnd.n3628 gnd.n3627 0.0269946
R14333 gnd.n4474 gnd.n4368 0.0225788
R14334 gnd.n4471 gnd.n4470 0.0225788
R14335 gnd.n4467 gnd.n4371 0.0225788
R14336 gnd.n4466 gnd.n4377 0.0225788
R14337 gnd.n4463 gnd.n4462 0.0225788
R14338 gnd.n4459 gnd.n4383 0.0225788
R14339 gnd.n4458 gnd.n4387 0.0225788
R14340 gnd.n4455 gnd.n4454 0.0225788
R14341 gnd.n4451 gnd.n4391 0.0225788
R14342 gnd.n4450 gnd.n4397 0.0225788
R14343 gnd.n4447 gnd.n4446 0.0225788
R14344 gnd.n4443 gnd.n4403 0.0225788
R14345 gnd.n4442 gnd.n4407 0.0225788
R14346 gnd.n4439 gnd.n4438 0.0225788
R14347 gnd.n4435 gnd.n4411 0.0225788
R14348 gnd.n4434 gnd.n4417 0.0225788
R14349 gnd.n4431 gnd.n4430 0.0225788
R14350 gnd.n4422 gnd.n2033 0.0225788
R14351 gnd.n4628 gnd.n4627 0.0225788
R14352 gnd.n5761 gnd.n1236 0.0225788
R14353 gnd.n5760 gnd.n1240 0.0225788
R14354 gnd.n5757 gnd.n5756 0.0225788
R14355 gnd.n5753 gnd.n1245 0.0225788
R14356 gnd.n5752 gnd.n1249 0.0225788
R14357 gnd.n5749 gnd.n5748 0.0225788
R14358 gnd.n5745 gnd.n1253 0.0225788
R14359 gnd.n5744 gnd.n1257 0.0225788
R14360 gnd.n5741 gnd.n5740 0.0225788
R14361 gnd.n5737 gnd.n1261 0.0225788
R14362 gnd.n5736 gnd.n1265 0.0225788
R14363 gnd.n5733 gnd.n5732 0.0225788
R14364 gnd.n5729 gnd.n1269 0.0225788
R14365 gnd.n5728 gnd.n1273 0.0225788
R14366 gnd.n5725 gnd.n5724 0.0225788
R14367 gnd.n5721 gnd.n1277 0.0225788
R14368 gnd.n5720 gnd.n1283 0.0225788
R14369 gnd.n1476 gnd.n1286 0.0225788
R14370 gnd.n5465 gnd.n1475 0.0225788
R14371 gnd.n5466 gnd.n1216 0.0218415
R14372 gnd.n4630 gnd.n4629 0.0218415
R14373 gnd.n2948 gnd.n2947 0.0202011
R14374 gnd.n2947 gnd.n2946 0.0148637
R14375 gnd.n3597 gnd.n3341 0.0144266
R14376 gnd.n3598 gnd.n3597 0.0130679
R14377 gnd.n4475 gnd.n4474 0.0123886
R14378 gnd.n4471 gnd.n4368 0.0123886
R14379 gnd.n4470 gnd.n4371 0.0123886
R14380 gnd.n4467 gnd.n4466 0.0123886
R14381 gnd.n4463 gnd.n4377 0.0123886
R14382 gnd.n4462 gnd.n4383 0.0123886
R14383 gnd.n4459 gnd.n4458 0.0123886
R14384 gnd.n4455 gnd.n4387 0.0123886
R14385 gnd.n4454 gnd.n4391 0.0123886
R14386 gnd.n4451 gnd.n4450 0.0123886
R14387 gnd.n4447 gnd.n4397 0.0123886
R14388 gnd.n4446 gnd.n4403 0.0123886
R14389 gnd.n4443 gnd.n4442 0.0123886
R14390 gnd.n4439 gnd.n4407 0.0123886
R14391 gnd.n4438 gnd.n4411 0.0123886
R14392 gnd.n4435 gnd.n4434 0.0123886
R14393 gnd.n4431 gnd.n4417 0.0123886
R14394 gnd.n4430 gnd.n4422 0.0123886
R14395 gnd.n4627 gnd.n2033 0.0123886
R14396 gnd.n5764 gnd.n1236 0.0123886
R14397 gnd.n5761 gnd.n5760 0.0123886
R14398 gnd.n5757 gnd.n1240 0.0123886
R14399 gnd.n5756 gnd.n1245 0.0123886
R14400 gnd.n5753 gnd.n5752 0.0123886
R14401 gnd.n5749 gnd.n1249 0.0123886
R14402 gnd.n5748 gnd.n1253 0.0123886
R14403 gnd.n5745 gnd.n5744 0.0123886
R14404 gnd.n5741 gnd.n1257 0.0123886
R14405 gnd.n5740 gnd.n1261 0.0123886
R14406 gnd.n5737 gnd.n5736 0.0123886
R14407 gnd.n5733 gnd.n1265 0.0123886
R14408 gnd.n5732 gnd.n1269 0.0123886
R14409 gnd.n5729 gnd.n5728 0.0123886
R14410 gnd.n5725 gnd.n1273 0.0123886
R14411 gnd.n5724 gnd.n1277 0.0123886
R14412 gnd.n5721 gnd.n5720 0.0123886
R14413 gnd.n1286 gnd.n1283 0.0123886
R14414 gnd.n1476 gnd.n1475 0.0123886
R14415 gnd.n2967 gnd.n2681 0.00797283
R14416 gnd.n2969 gnd.n2968 0.00797283
R14417 gnd.n2970 gnd.n2676 0.00797283
R14418 gnd.n2978 gnd.n2674 0.00797283
R14419 gnd.n2980 gnd.n2979 0.00797283
R14420 gnd.n2998 gnd.n2655 0.00797283
R14421 gnd.n3000 gnd.n2999 0.00797283
R14422 gnd.n3001 gnd.n2650 0.00797283
R14423 gnd.n2649 gnd.n2645 0.00797283
R14424 gnd.n3011 gnd.n3010 0.00797283
R14425 gnd.n2647 gnd.n2646 0.00797283
R14426 gnd.n2629 gnd.n2628 0.00797283
R14427 gnd.n3031 gnd.n3030 0.00797283
R14428 gnd.n2630 gnd.n2605 0.00797283
R14429 gnd.n3065 gnd.n3064 0.00797283
R14430 gnd.n3067 gnd.n3066 0.00797283
R14431 gnd.n2600 gnd.n2552 0.00797283
R14432 gnd.n2602 gnd.n2553 0.00797283
R14433 gnd.n3076 gnd.n2554 0.00797283
R14434 gnd.n3078 gnd.n3077 0.00797283
R14435 gnd.n3080 gnd.n3079 0.00797283
R14436 gnd.n3082 gnd.n2574 0.00797283
R14437 gnd.n3085 gnd.n2575 0.00797283
R14438 gnd.n3087 gnd.n2576 0.00797283
R14439 gnd.n3090 gnd.n3088 0.00797283
R14440 gnd.n3089 gnd.n2459 0.00797283
R14441 gnd.n3157 gnd.n3155 0.00797283
R14442 gnd.n3156 gnd.n2452 0.00797283
R14443 gnd.n3167 gnd.n3166 0.00797283
R14444 gnd.n3169 gnd.n3168 0.00797283
R14445 gnd.n3172 gnd.n2450 0.00797283
R14446 gnd.n3176 gnd.n3175 0.00797283
R14447 gnd.n3174 gnd.n3173 0.00797283
R14448 gnd.n2430 gnd.n2429 0.00797283
R14449 gnd.n3198 gnd.n3197 0.00797283
R14450 gnd.n2431 gnd.n2404 0.00797283
R14451 gnd.n3242 gnd.n3240 0.00797283
R14452 gnd.n3241 gnd.n2397 0.00797283
R14453 gnd.n3252 gnd.n3251 0.00797283
R14454 gnd.n3254 gnd.n3253 0.00797283
R14455 gnd.n3257 gnd.n2395 0.00797283
R14456 gnd.n3261 gnd.n3260 0.00797283
R14457 gnd.n3259 gnd.n3258 0.00797283
R14458 gnd.n2375 gnd.n2374 0.00797283
R14459 gnd.n3283 gnd.n3282 0.00797283
R14460 gnd.n2376 gnd.n2350 0.00797283
R14461 gnd.n3331 gnd.n3329 0.00797283
R14462 gnd.n3330 gnd.n2343 0.00797283
R14463 gnd.n3341 gnd.n3340 0.00797283
R14464 gnd.n3599 gnd.n3598 0.00797283
R14465 gnd.n3602 gnd.n2341 0.00797283
R14466 gnd.n3604 gnd.n3603 0.00797283
R14467 gnd.n3627 gnd.n2322 0.00797283
R14468 gnd.n3628 gnd.n2285 0.00797283
R14469 gnd.n4480 gnd.n4335 0.00593478
R14470 gnd.n5766 gnd.n5765 0.00593478
R14471 gnd.n6877 gnd.n326 0.00417647
R14472 gnd.n6878 gnd.n6877 0.00417647
R14473 gnd.n6879 gnd.n6878 0.00417647
R14474 gnd.n6881 gnd.n6879 0.00417647
R14475 gnd.n6881 gnd.n6880 0.00417647
R14476 gnd.n6880 gnd.n91 0.00417647
R14477 gnd.n92 gnd.n91 0.00417647
R14478 gnd.n93 gnd.n92 0.00417647
R14479 gnd.n111 gnd.n93 0.00417647
R14480 gnd.n4186 gnd.n2126 0.00417647
R14481 gnd.n4187 gnd.n4186 0.00417647
R14482 gnd.n4188 gnd.n4187 0.00417647
R14483 gnd.n4189 gnd.n4188 0.00417647
R14484 gnd.n4189 gnd.n2101 0.00417647
R14485 gnd.n4229 gnd.n2101 0.00417647
R14486 gnd.n4230 gnd.n4229 0.00417647
R14487 gnd.n4231 gnd.n4230 0.00417647
R14488 gnd.n4231 gnd.n2080 0.00417647
R14489 CSoutput.n19 CSoutput.t160 184.661
R14490 CSoutput.n78 CSoutput.n77 165.8
R14491 CSoutput.n76 CSoutput.n0 165.8
R14492 CSoutput.n75 CSoutput.n74 165.8
R14493 CSoutput.n73 CSoutput.n72 165.8
R14494 CSoutput.n71 CSoutput.n2 165.8
R14495 CSoutput.n69 CSoutput.n68 165.8
R14496 CSoutput.n67 CSoutput.n3 165.8
R14497 CSoutput.n66 CSoutput.n65 165.8
R14498 CSoutput.n63 CSoutput.n4 165.8
R14499 CSoutput.n61 CSoutput.n60 165.8
R14500 CSoutput.n59 CSoutput.n5 165.8
R14501 CSoutput.n58 CSoutput.n57 165.8
R14502 CSoutput.n55 CSoutput.n6 165.8
R14503 CSoutput.n54 CSoutput.n53 165.8
R14504 CSoutput.n52 CSoutput.n51 165.8
R14505 CSoutput.n50 CSoutput.n8 165.8
R14506 CSoutput.n48 CSoutput.n47 165.8
R14507 CSoutput.n46 CSoutput.n9 165.8
R14508 CSoutput.n45 CSoutput.n44 165.8
R14509 CSoutput.n42 CSoutput.n10 165.8
R14510 CSoutput.n41 CSoutput.n40 165.8
R14511 CSoutput.n39 CSoutput.n38 165.8
R14512 CSoutput.n37 CSoutput.n12 165.8
R14513 CSoutput.n35 CSoutput.n34 165.8
R14514 CSoutput.n33 CSoutput.n13 165.8
R14515 CSoutput.n32 CSoutput.n31 165.8
R14516 CSoutput.n29 CSoutput.n14 165.8
R14517 CSoutput.n28 CSoutput.n27 165.8
R14518 CSoutput.n26 CSoutput.n25 165.8
R14519 CSoutput.n24 CSoutput.n16 165.8
R14520 CSoutput.n22 CSoutput.n21 165.8
R14521 CSoutput.n20 CSoutput.n17 165.8
R14522 CSoutput.n77 CSoutput.t161 162.194
R14523 CSoutput.n18 CSoutput.t157 120.501
R14524 CSoutput.n23 CSoutput.t151 120.501
R14525 CSoutput.n15 CSoutput.t145 120.501
R14526 CSoutput.n30 CSoutput.t158 120.501
R14527 CSoutput.n36 CSoutput.t159 120.501
R14528 CSoutput.n11 CSoutput.t147 120.501
R14529 CSoutput.n43 CSoutput.t165 120.501
R14530 CSoutput.n49 CSoutput.t162 120.501
R14531 CSoutput.n7 CSoutput.t150 120.501
R14532 CSoutput.n56 CSoutput.t152 120.501
R14533 CSoutput.n62 CSoutput.t163 120.501
R14534 CSoutput.n64 CSoutput.t154 120.501
R14535 CSoutput.n70 CSoutput.t156 120.501
R14536 CSoutput.n1 CSoutput.t148 120.501
R14537 CSoutput.n270 CSoutput.n268 103.469
R14538 CSoutput.n262 CSoutput.n260 103.469
R14539 CSoutput.n255 CSoutput.n253 103.469
R14540 CSoutput.n96 CSoutput.n94 103.469
R14541 CSoutput.n88 CSoutput.n86 103.469
R14542 CSoutput.n81 CSoutput.n79 103.469
R14543 CSoutput.n272 CSoutput.n271 103.111
R14544 CSoutput.n270 CSoutput.n269 103.111
R14545 CSoutput.n266 CSoutput.n265 103.111
R14546 CSoutput.n264 CSoutput.n263 103.111
R14547 CSoutput.n262 CSoutput.n261 103.111
R14548 CSoutput.n259 CSoutput.n258 103.111
R14549 CSoutput.n257 CSoutput.n256 103.111
R14550 CSoutput.n255 CSoutput.n254 103.111
R14551 CSoutput.n96 CSoutput.n95 103.111
R14552 CSoutput.n98 CSoutput.n97 103.111
R14553 CSoutput.n100 CSoutput.n99 103.111
R14554 CSoutput.n88 CSoutput.n87 103.111
R14555 CSoutput.n90 CSoutput.n89 103.111
R14556 CSoutput.n92 CSoutput.n91 103.111
R14557 CSoutput.n81 CSoutput.n80 103.111
R14558 CSoutput.n83 CSoutput.n82 103.111
R14559 CSoutput.n85 CSoutput.n84 103.111
R14560 CSoutput.n274 CSoutput.n273 103.111
R14561 CSoutput.n310 CSoutput.n308 81.5057
R14562 CSoutput.n294 CSoutput.n292 81.5057
R14563 CSoutput.n279 CSoutput.n277 81.5057
R14564 CSoutput.n358 CSoutput.n356 81.5057
R14565 CSoutput.n342 CSoutput.n340 81.5057
R14566 CSoutput.n327 CSoutput.n325 81.5057
R14567 CSoutput.n322 CSoutput.n321 80.9324
R14568 CSoutput.n320 CSoutput.n319 80.9324
R14569 CSoutput.n318 CSoutput.n317 80.9324
R14570 CSoutput.n316 CSoutput.n315 80.9324
R14571 CSoutput.n314 CSoutput.n313 80.9324
R14572 CSoutput.n312 CSoutput.n311 80.9324
R14573 CSoutput.n310 CSoutput.n309 80.9324
R14574 CSoutput.n306 CSoutput.n305 80.9324
R14575 CSoutput.n304 CSoutput.n303 80.9324
R14576 CSoutput.n302 CSoutput.n301 80.9324
R14577 CSoutput.n300 CSoutput.n299 80.9324
R14578 CSoutput.n298 CSoutput.n297 80.9324
R14579 CSoutput.n296 CSoutput.n295 80.9324
R14580 CSoutput.n294 CSoutput.n293 80.9324
R14581 CSoutput.n291 CSoutput.n290 80.9324
R14582 CSoutput.n289 CSoutput.n288 80.9324
R14583 CSoutput.n287 CSoutput.n286 80.9324
R14584 CSoutput.n285 CSoutput.n284 80.9324
R14585 CSoutput.n283 CSoutput.n282 80.9324
R14586 CSoutput.n281 CSoutput.n280 80.9324
R14587 CSoutput.n279 CSoutput.n278 80.9324
R14588 CSoutput.n358 CSoutput.n357 80.9324
R14589 CSoutput.n360 CSoutput.n359 80.9324
R14590 CSoutput.n362 CSoutput.n361 80.9324
R14591 CSoutput.n364 CSoutput.n363 80.9324
R14592 CSoutput.n366 CSoutput.n365 80.9324
R14593 CSoutput.n368 CSoutput.n367 80.9324
R14594 CSoutput.n370 CSoutput.n369 80.9324
R14595 CSoutput.n342 CSoutput.n341 80.9324
R14596 CSoutput.n344 CSoutput.n343 80.9324
R14597 CSoutput.n346 CSoutput.n345 80.9324
R14598 CSoutput.n348 CSoutput.n347 80.9324
R14599 CSoutput.n350 CSoutput.n349 80.9324
R14600 CSoutput.n352 CSoutput.n351 80.9324
R14601 CSoutput.n354 CSoutput.n353 80.9324
R14602 CSoutput.n327 CSoutput.n326 80.9324
R14603 CSoutput.n329 CSoutput.n328 80.9324
R14604 CSoutput.n331 CSoutput.n330 80.9324
R14605 CSoutput.n333 CSoutput.n332 80.9324
R14606 CSoutput.n335 CSoutput.n334 80.9324
R14607 CSoutput.n337 CSoutput.n336 80.9324
R14608 CSoutput.n339 CSoutput.n338 80.9324
R14609 CSoutput.n25 CSoutput.n24 48.1486
R14610 CSoutput.n69 CSoutput.n3 48.1486
R14611 CSoutput.n38 CSoutput.n37 48.1486
R14612 CSoutput.n42 CSoutput.n41 48.1486
R14613 CSoutput.n51 CSoutput.n50 48.1486
R14614 CSoutput.n55 CSoutput.n54 48.1486
R14615 CSoutput.n22 CSoutput.n17 46.462
R14616 CSoutput.n72 CSoutput.n71 46.462
R14617 CSoutput.n20 CSoutput.n19 44.9055
R14618 CSoutput.n29 CSoutput.n28 43.7635
R14619 CSoutput.n65 CSoutput.n63 43.7635
R14620 CSoutput.n35 CSoutput.n13 41.7396
R14621 CSoutput.n57 CSoutput.n5 41.7396
R14622 CSoutput.n44 CSoutput.n9 37.0171
R14623 CSoutput.n48 CSoutput.n9 37.0171
R14624 CSoutput.n76 CSoutput.n75 34.9932
R14625 CSoutput.n31 CSoutput.n13 32.2947
R14626 CSoutput.n61 CSoutput.n5 32.2947
R14627 CSoutput.n30 CSoutput.n29 29.6014
R14628 CSoutput.n63 CSoutput.n62 29.6014
R14629 CSoutput.n19 CSoutput.n18 28.4085
R14630 CSoutput.n18 CSoutput.n17 25.1176
R14631 CSoutput.n72 CSoutput.n1 25.1176
R14632 CSoutput.n43 CSoutput.n42 22.0922
R14633 CSoutput.n50 CSoutput.n49 22.0922
R14634 CSoutput.n77 CSoutput.n76 21.8586
R14635 CSoutput.n37 CSoutput.n36 18.9681
R14636 CSoutput.n56 CSoutput.n55 18.9681
R14637 CSoutput.n25 CSoutput.n15 17.6292
R14638 CSoutput.n64 CSoutput.n3 17.6292
R14639 CSoutput.n24 CSoutput.n23 15.844
R14640 CSoutput.n70 CSoutput.n69 15.844
R14641 CSoutput.n38 CSoutput.n11 14.5051
R14642 CSoutput.n54 CSoutput.n7 14.5051
R14643 CSoutput.n373 CSoutput.n78 11.4982
R14644 CSoutput.n41 CSoutput.n11 11.3811
R14645 CSoutput.n51 CSoutput.n7 11.3811
R14646 CSoutput.n23 CSoutput.n22 10.0422
R14647 CSoutput.n71 CSoutput.n70 10.0422
R14648 CSoutput.n267 CSoutput.n259 9.25285
R14649 CSoutput.n93 CSoutput.n85 9.25285
R14650 CSoutput.n324 CSoutput.n276 9.09499
R14651 CSoutput.n307 CSoutput.n291 8.98182
R14652 CSoutput.n355 CSoutput.n339 8.98182
R14653 CSoutput.n28 CSoutput.n15 8.25698
R14654 CSoutput.n65 CSoutput.n64 8.25698
R14655 CSoutput.n276 CSoutput.n275 7.12641
R14656 CSoutput.n102 CSoutput.n101 7.12641
R14657 CSoutput.n36 CSoutput.n35 6.91809
R14658 CSoutput.n57 CSoutput.n56 6.91809
R14659 CSoutput.n324 CSoutput.n323 6.02792
R14660 CSoutput.n372 CSoutput.n371 6.02792
R14661 CSoutput.n373 CSoutput.n102 5.50255
R14662 CSoutput.n323 CSoutput.n322 5.25266
R14663 CSoutput.n307 CSoutput.n306 5.25266
R14664 CSoutput.n371 CSoutput.n370 5.25266
R14665 CSoutput.n355 CSoutput.n354 5.25266
R14666 CSoutput.n275 CSoutput.n274 5.1449
R14667 CSoutput.n267 CSoutput.n266 5.1449
R14668 CSoutput.n101 CSoutput.n100 5.1449
R14669 CSoutput.n93 CSoutput.n92 5.1449
R14670 CSoutput.n193 CSoutput.n146 4.5005
R14671 CSoutput.n162 CSoutput.n146 4.5005
R14672 CSoutput.n157 CSoutput.n141 4.5005
R14673 CSoutput.n157 CSoutput.n143 4.5005
R14674 CSoutput.n157 CSoutput.n140 4.5005
R14675 CSoutput.n157 CSoutput.n144 4.5005
R14676 CSoutput.n157 CSoutput.n139 4.5005
R14677 CSoutput.n157 CSoutput.t164 4.5005
R14678 CSoutput.n157 CSoutput.n138 4.5005
R14679 CSoutput.n157 CSoutput.n145 4.5005
R14680 CSoutput.n157 CSoutput.n146 4.5005
R14681 CSoutput.n155 CSoutput.n141 4.5005
R14682 CSoutput.n155 CSoutput.n143 4.5005
R14683 CSoutput.n155 CSoutput.n140 4.5005
R14684 CSoutput.n155 CSoutput.n144 4.5005
R14685 CSoutput.n155 CSoutput.n139 4.5005
R14686 CSoutput.n155 CSoutput.t164 4.5005
R14687 CSoutput.n155 CSoutput.n138 4.5005
R14688 CSoutput.n155 CSoutput.n145 4.5005
R14689 CSoutput.n155 CSoutput.n146 4.5005
R14690 CSoutput.n154 CSoutput.n141 4.5005
R14691 CSoutput.n154 CSoutput.n143 4.5005
R14692 CSoutput.n154 CSoutput.n140 4.5005
R14693 CSoutput.n154 CSoutput.n144 4.5005
R14694 CSoutput.n154 CSoutput.n139 4.5005
R14695 CSoutput.n154 CSoutput.t164 4.5005
R14696 CSoutput.n154 CSoutput.n138 4.5005
R14697 CSoutput.n154 CSoutput.n145 4.5005
R14698 CSoutput.n154 CSoutput.n146 4.5005
R14699 CSoutput.n239 CSoutput.n141 4.5005
R14700 CSoutput.n239 CSoutput.n143 4.5005
R14701 CSoutput.n239 CSoutput.n140 4.5005
R14702 CSoutput.n239 CSoutput.n144 4.5005
R14703 CSoutput.n239 CSoutput.n139 4.5005
R14704 CSoutput.n239 CSoutput.t164 4.5005
R14705 CSoutput.n239 CSoutput.n138 4.5005
R14706 CSoutput.n239 CSoutput.n145 4.5005
R14707 CSoutput.n239 CSoutput.n146 4.5005
R14708 CSoutput.n237 CSoutput.n141 4.5005
R14709 CSoutput.n237 CSoutput.n143 4.5005
R14710 CSoutput.n237 CSoutput.n140 4.5005
R14711 CSoutput.n237 CSoutput.n144 4.5005
R14712 CSoutput.n237 CSoutput.n139 4.5005
R14713 CSoutput.n237 CSoutput.t164 4.5005
R14714 CSoutput.n237 CSoutput.n138 4.5005
R14715 CSoutput.n237 CSoutput.n145 4.5005
R14716 CSoutput.n235 CSoutput.n141 4.5005
R14717 CSoutput.n235 CSoutput.n143 4.5005
R14718 CSoutput.n235 CSoutput.n140 4.5005
R14719 CSoutput.n235 CSoutput.n144 4.5005
R14720 CSoutput.n235 CSoutput.n139 4.5005
R14721 CSoutput.n235 CSoutput.t164 4.5005
R14722 CSoutput.n235 CSoutput.n138 4.5005
R14723 CSoutput.n235 CSoutput.n145 4.5005
R14724 CSoutput.n165 CSoutput.n141 4.5005
R14725 CSoutput.n165 CSoutput.n143 4.5005
R14726 CSoutput.n165 CSoutput.n140 4.5005
R14727 CSoutput.n165 CSoutput.n144 4.5005
R14728 CSoutput.n165 CSoutput.n139 4.5005
R14729 CSoutput.n165 CSoutput.t164 4.5005
R14730 CSoutput.n165 CSoutput.n138 4.5005
R14731 CSoutput.n165 CSoutput.n145 4.5005
R14732 CSoutput.n165 CSoutput.n146 4.5005
R14733 CSoutput.n164 CSoutput.n141 4.5005
R14734 CSoutput.n164 CSoutput.n143 4.5005
R14735 CSoutput.n164 CSoutput.n140 4.5005
R14736 CSoutput.n164 CSoutput.n144 4.5005
R14737 CSoutput.n164 CSoutput.n139 4.5005
R14738 CSoutput.n164 CSoutput.t164 4.5005
R14739 CSoutput.n164 CSoutput.n138 4.5005
R14740 CSoutput.n164 CSoutput.n145 4.5005
R14741 CSoutput.n164 CSoutput.n146 4.5005
R14742 CSoutput.n168 CSoutput.n141 4.5005
R14743 CSoutput.n168 CSoutput.n143 4.5005
R14744 CSoutput.n168 CSoutput.n140 4.5005
R14745 CSoutput.n168 CSoutput.n144 4.5005
R14746 CSoutput.n168 CSoutput.n139 4.5005
R14747 CSoutput.n168 CSoutput.t164 4.5005
R14748 CSoutput.n168 CSoutput.n138 4.5005
R14749 CSoutput.n168 CSoutput.n145 4.5005
R14750 CSoutput.n168 CSoutput.n146 4.5005
R14751 CSoutput.n167 CSoutput.n141 4.5005
R14752 CSoutput.n167 CSoutput.n143 4.5005
R14753 CSoutput.n167 CSoutput.n140 4.5005
R14754 CSoutput.n167 CSoutput.n144 4.5005
R14755 CSoutput.n167 CSoutput.n139 4.5005
R14756 CSoutput.n167 CSoutput.t164 4.5005
R14757 CSoutput.n167 CSoutput.n138 4.5005
R14758 CSoutput.n167 CSoutput.n145 4.5005
R14759 CSoutput.n167 CSoutput.n146 4.5005
R14760 CSoutput.n150 CSoutput.n141 4.5005
R14761 CSoutput.n150 CSoutput.n143 4.5005
R14762 CSoutput.n150 CSoutput.n140 4.5005
R14763 CSoutput.n150 CSoutput.n144 4.5005
R14764 CSoutput.n150 CSoutput.n139 4.5005
R14765 CSoutput.n150 CSoutput.t164 4.5005
R14766 CSoutput.n150 CSoutput.n138 4.5005
R14767 CSoutput.n150 CSoutput.n145 4.5005
R14768 CSoutput.n150 CSoutput.n146 4.5005
R14769 CSoutput.n242 CSoutput.n141 4.5005
R14770 CSoutput.n242 CSoutput.n143 4.5005
R14771 CSoutput.n242 CSoutput.n140 4.5005
R14772 CSoutput.n242 CSoutput.n144 4.5005
R14773 CSoutput.n242 CSoutput.n139 4.5005
R14774 CSoutput.n242 CSoutput.t164 4.5005
R14775 CSoutput.n242 CSoutput.n138 4.5005
R14776 CSoutput.n242 CSoutput.n145 4.5005
R14777 CSoutput.n242 CSoutput.n146 4.5005
R14778 CSoutput.n229 CSoutput.n200 4.5005
R14779 CSoutput.n229 CSoutput.n206 4.5005
R14780 CSoutput.n187 CSoutput.n176 4.5005
R14781 CSoutput.n187 CSoutput.n178 4.5005
R14782 CSoutput.n187 CSoutput.n175 4.5005
R14783 CSoutput.n187 CSoutput.n179 4.5005
R14784 CSoutput.n187 CSoutput.n174 4.5005
R14785 CSoutput.n187 CSoutput.t144 4.5005
R14786 CSoutput.n187 CSoutput.n173 4.5005
R14787 CSoutput.n187 CSoutput.n180 4.5005
R14788 CSoutput.n229 CSoutput.n187 4.5005
R14789 CSoutput.n208 CSoutput.n176 4.5005
R14790 CSoutput.n208 CSoutput.n178 4.5005
R14791 CSoutput.n208 CSoutput.n175 4.5005
R14792 CSoutput.n208 CSoutput.n179 4.5005
R14793 CSoutput.n208 CSoutput.n174 4.5005
R14794 CSoutput.n208 CSoutput.t144 4.5005
R14795 CSoutput.n208 CSoutput.n173 4.5005
R14796 CSoutput.n208 CSoutput.n180 4.5005
R14797 CSoutput.n229 CSoutput.n208 4.5005
R14798 CSoutput.n186 CSoutput.n176 4.5005
R14799 CSoutput.n186 CSoutput.n178 4.5005
R14800 CSoutput.n186 CSoutput.n175 4.5005
R14801 CSoutput.n186 CSoutput.n179 4.5005
R14802 CSoutput.n186 CSoutput.n174 4.5005
R14803 CSoutput.n186 CSoutput.t144 4.5005
R14804 CSoutput.n186 CSoutput.n173 4.5005
R14805 CSoutput.n186 CSoutput.n180 4.5005
R14806 CSoutput.n229 CSoutput.n186 4.5005
R14807 CSoutput.n210 CSoutput.n176 4.5005
R14808 CSoutput.n210 CSoutput.n178 4.5005
R14809 CSoutput.n210 CSoutput.n175 4.5005
R14810 CSoutput.n210 CSoutput.n179 4.5005
R14811 CSoutput.n210 CSoutput.n174 4.5005
R14812 CSoutput.n210 CSoutput.t144 4.5005
R14813 CSoutput.n210 CSoutput.n173 4.5005
R14814 CSoutput.n210 CSoutput.n180 4.5005
R14815 CSoutput.n229 CSoutput.n210 4.5005
R14816 CSoutput.n176 CSoutput.n171 4.5005
R14817 CSoutput.n178 CSoutput.n171 4.5005
R14818 CSoutput.n175 CSoutput.n171 4.5005
R14819 CSoutput.n179 CSoutput.n171 4.5005
R14820 CSoutput.n174 CSoutput.n171 4.5005
R14821 CSoutput.t144 CSoutput.n171 4.5005
R14822 CSoutput.n173 CSoutput.n171 4.5005
R14823 CSoutput.n180 CSoutput.n171 4.5005
R14824 CSoutput.n232 CSoutput.n176 4.5005
R14825 CSoutput.n232 CSoutput.n178 4.5005
R14826 CSoutput.n232 CSoutput.n175 4.5005
R14827 CSoutput.n232 CSoutput.n179 4.5005
R14828 CSoutput.n232 CSoutput.n174 4.5005
R14829 CSoutput.n232 CSoutput.t144 4.5005
R14830 CSoutput.n232 CSoutput.n173 4.5005
R14831 CSoutput.n232 CSoutput.n180 4.5005
R14832 CSoutput.n230 CSoutput.n176 4.5005
R14833 CSoutput.n230 CSoutput.n178 4.5005
R14834 CSoutput.n230 CSoutput.n175 4.5005
R14835 CSoutput.n230 CSoutput.n179 4.5005
R14836 CSoutput.n230 CSoutput.n174 4.5005
R14837 CSoutput.n230 CSoutput.t144 4.5005
R14838 CSoutput.n230 CSoutput.n173 4.5005
R14839 CSoutput.n230 CSoutput.n180 4.5005
R14840 CSoutput.n230 CSoutput.n229 4.5005
R14841 CSoutput.n212 CSoutput.n176 4.5005
R14842 CSoutput.n212 CSoutput.n178 4.5005
R14843 CSoutput.n212 CSoutput.n175 4.5005
R14844 CSoutput.n212 CSoutput.n179 4.5005
R14845 CSoutput.n212 CSoutput.n174 4.5005
R14846 CSoutput.n212 CSoutput.t144 4.5005
R14847 CSoutput.n212 CSoutput.n173 4.5005
R14848 CSoutput.n212 CSoutput.n180 4.5005
R14849 CSoutput.n229 CSoutput.n212 4.5005
R14850 CSoutput.n184 CSoutput.n176 4.5005
R14851 CSoutput.n184 CSoutput.n178 4.5005
R14852 CSoutput.n184 CSoutput.n175 4.5005
R14853 CSoutput.n184 CSoutput.n179 4.5005
R14854 CSoutput.n184 CSoutput.n174 4.5005
R14855 CSoutput.n184 CSoutput.t144 4.5005
R14856 CSoutput.n184 CSoutput.n173 4.5005
R14857 CSoutput.n184 CSoutput.n180 4.5005
R14858 CSoutput.n229 CSoutput.n184 4.5005
R14859 CSoutput.n214 CSoutput.n176 4.5005
R14860 CSoutput.n214 CSoutput.n178 4.5005
R14861 CSoutput.n214 CSoutput.n175 4.5005
R14862 CSoutput.n214 CSoutput.n179 4.5005
R14863 CSoutput.n214 CSoutput.n174 4.5005
R14864 CSoutput.n214 CSoutput.t144 4.5005
R14865 CSoutput.n214 CSoutput.n173 4.5005
R14866 CSoutput.n214 CSoutput.n180 4.5005
R14867 CSoutput.n229 CSoutput.n214 4.5005
R14868 CSoutput.n183 CSoutput.n176 4.5005
R14869 CSoutput.n183 CSoutput.n178 4.5005
R14870 CSoutput.n183 CSoutput.n175 4.5005
R14871 CSoutput.n183 CSoutput.n179 4.5005
R14872 CSoutput.n183 CSoutput.n174 4.5005
R14873 CSoutput.n183 CSoutput.t144 4.5005
R14874 CSoutput.n183 CSoutput.n173 4.5005
R14875 CSoutput.n183 CSoutput.n180 4.5005
R14876 CSoutput.n229 CSoutput.n183 4.5005
R14877 CSoutput.n228 CSoutput.n176 4.5005
R14878 CSoutput.n228 CSoutput.n178 4.5005
R14879 CSoutput.n228 CSoutput.n175 4.5005
R14880 CSoutput.n228 CSoutput.n179 4.5005
R14881 CSoutput.n228 CSoutput.n174 4.5005
R14882 CSoutput.n228 CSoutput.t144 4.5005
R14883 CSoutput.n228 CSoutput.n173 4.5005
R14884 CSoutput.n228 CSoutput.n180 4.5005
R14885 CSoutput.n229 CSoutput.n228 4.5005
R14886 CSoutput.n227 CSoutput.n112 4.5005
R14887 CSoutput.n128 CSoutput.n112 4.5005
R14888 CSoutput.n123 CSoutput.n107 4.5005
R14889 CSoutput.n123 CSoutput.n109 4.5005
R14890 CSoutput.n123 CSoutput.n106 4.5005
R14891 CSoutput.n123 CSoutput.n110 4.5005
R14892 CSoutput.n123 CSoutput.n105 4.5005
R14893 CSoutput.n123 CSoutput.t153 4.5005
R14894 CSoutput.n123 CSoutput.n104 4.5005
R14895 CSoutput.n123 CSoutput.n111 4.5005
R14896 CSoutput.n123 CSoutput.n112 4.5005
R14897 CSoutput.n121 CSoutput.n107 4.5005
R14898 CSoutput.n121 CSoutput.n109 4.5005
R14899 CSoutput.n121 CSoutput.n106 4.5005
R14900 CSoutput.n121 CSoutput.n110 4.5005
R14901 CSoutput.n121 CSoutput.n105 4.5005
R14902 CSoutput.n121 CSoutput.t153 4.5005
R14903 CSoutput.n121 CSoutput.n104 4.5005
R14904 CSoutput.n121 CSoutput.n111 4.5005
R14905 CSoutput.n121 CSoutput.n112 4.5005
R14906 CSoutput.n120 CSoutput.n107 4.5005
R14907 CSoutput.n120 CSoutput.n109 4.5005
R14908 CSoutput.n120 CSoutput.n106 4.5005
R14909 CSoutput.n120 CSoutput.n110 4.5005
R14910 CSoutput.n120 CSoutput.n105 4.5005
R14911 CSoutput.n120 CSoutput.t153 4.5005
R14912 CSoutput.n120 CSoutput.n104 4.5005
R14913 CSoutput.n120 CSoutput.n111 4.5005
R14914 CSoutput.n120 CSoutput.n112 4.5005
R14915 CSoutput.n249 CSoutput.n107 4.5005
R14916 CSoutput.n249 CSoutput.n109 4.5005
R14917 CSoutput.n249 CSoutput.n106 4.5005
R14918 CSoutput.n249 CSoutput.n110 4.5005
R14919 CSoutput.n249 CSoutput.n105 4.5005
R14920 CSoutput.n249 CSoutput.t153 4.5005
R14921 CSoutput.n249 CSoutput.n104 4.5005
R14922 CSoutput.n249 CSoutput.n111 4.5005
R14923 CSoutput.n249 CSoutput.n112 4.5005
R14924 CSoutput.n247 CSoutput.n107 4.5005
R14925 CSoutput.n247 CSoutput.n109 4.5005
R14926 CSoutput.n247 CSoutput.n106 4.5005
R14927 CSoutput.n247 CSoutput.n110 4.5005
R14928 CSoutput.n247 CSoutput.n105 4.5005
R14929 CSoutput.n247 CSoutput.t153 4.5005
R14930 CSoutput.n247 CSoutput.n104 4.5005
R14931 CSoutput.n247 CSoutput.n111 4.5005
R14932 CSoutput.n245 CSoutput.n107 4.5005
R14933 CSoutput.n245 CSoutput.n109 4.5005
R14934 CSoutput.n245 CSoutput.n106 4.5005
R14935 CSoutput.n245 CSoutput.n110 4.5005
R14936 CSoutput.n245 CSoutput.n105 4.5005
R14937 CSoutput.n245 CSoutput.t153 4.5005
R14938 CSoutput.n245 CSoutput.n104 4.5005
R14939 CSoutput.n245 CSoutput.n111 4.5005
R14940 CSoutput.n131 CSoutput.n107 4.5005
R14941 CSoutput.n131 CSoutput.n109 4.5005
R14942 CSoutput.n131 CSoutput.n106 4.5005
R14943 CSoutput.n131 CSoutput.n110 4.5005
R14944 CSoutput.n131 CSoutput.n105 4.5005
R14945 CSoutput.n131 CSoutput.t153 4.5005
R14946 CSoutput.n131 CSoutput.n104 4.5005
R14947 CSoutput.n131 CSoutput.n111 4.5005
R14948 CSoutput.n131 CSoutput.n112 4.5005
R14949 CSoutput.n130 CSoutput.n107 4.5005
R14950 CSoutput.n130 CSoutput.n109 4.5005
R14951 CSoutput.n130 CSoutput.n106 4.5005
R14952 CSoutput.n130 CSoutput.n110 4.5005
R14953 CSoutput.n130 CSoutput.n105 4.5005
R14954 CSoutput.n130 CSoutput.t153 4.5005
R14955 CSoutput.n130 CSoutput.n104 4.5005
R14956 CSoutput.n130 CSoutput.n111 4.5005
R14957 CSoutput.n130 CSoutput.n112 4.5005
R14958 CSoutput.n134 CSoutput.n107 4.5005
R14959 CSoutput.n134 CSoutput.n109 4.5005
R14960 CSoutput.n134 CSoutput.n106 4.5005
R14961 CSoutput.n134 CSoutput.n110 4.5005
R14962 CSoutput.n134 CSoutput.n105 4.5005
R14963 CSoutput.n134 CSoutput.t153 4.5005
R14964 CSoutput.n134 CSoutput.n104 4.5005
R14965 CSoutput.n134 CSoutput.n111 4.5005
R14966 CSoutput.n134 CSoutput.n112 4.5005
R14967 CSoutput.n133 CSoutput.n107 4.5005
R14968 CSoutput.n133 CSoutput.n109 4.5005
R14969 CSoutput.n133 CSoutput.n106 4.5005
R14970 CSoutput.n133 CSoutput.n110 4.5005
R14971 CSoutput.n133 CSoutput.n105 4.5005
R14972 CSoutput.n133 CSoutput.t153 4.5005
R14973 CSoutput.n133 CSoutput.n104 4.5005
R14974 CSoutput.n133 CSoutput.n111 4.5005
R14975 CSoutput.n133 CSoutput.n112 4.5005
R14976 CSoutput.n116 CSoutput.n107 4.5005
R14977 CSoutput.n116 CSoutput.n109 4.5005
R14978 CSoutput.n116 CSoutput.n106 4.5005
R14979 CSoutput.n116 CSoutput.n110 4.5005
R14980 CSoutput.n116 CSoutput.n105 4.5005
R14981 CSoutput.n116 CSoutput.t153 4.5005
R14982 CSoutput.n116 CSoutput.n104 4.5005
R14983 CSoutput.n116 CSoutput.n111 4.5005
R14984 CSoutput.n116 CSoutput.n112 4.5005
R14985 CSoutput.n252 CSoutput.n107 4.5005
R14986 CSoutput.n252 CSoutput.n109 4.5005
R14987 CSoutput.n252 CSoutput.n106 4.5005
R14988 CSoutput.n252 CSoutput.n110 4.5005
R14989 CSoutput.n252 CSoutput.n105 4.5005
R14990 CSoutput.n252 CSoutput.t153 4.5005
R14991 CSoutput.n252 CSoutput.n104 4.5005
R14992 CSoutput.n252 CSoutput.n111 4.5005
R14993 CSoutput.n252 CSoutput.n112 4.5005
R14994 CSoutput.n275 CSoutput.n267 4.10845
R14995 CSoutput.n101 CSoutput.n93 4.10845
R14996 CSoutput.n273 CSoutput.t33 4.06363
R14997 CSoutput.n273 CSoutput.t0 4.06363
R14998 CSoutput.n271 CSoutput.t37 4.06363
R14999 CSoutput.n271 CSoutput.t140 4.06363
R15000 CSoutput.n269 CSoutput.t12 4.06363
R15001 CSoutput.n269 CSoutput.t2 4.06363
R15002 CSoutput.n268 CSoutput.t24 4.06363
R15003 CSoutput.n268 CSoutput.t141 4.06363
R15004 CSoutput.n265 CSoutput.t139 4.06363
R15005 CSoutput.n265 CSoutput.t17 4.06363
R15006 CSoutput.n263 CSoutput.t25 4.06363
R15007 CSoutput.n263 CSoutput.t14 4.06363
R15008 CSoutput.n261 CSoutput.t6 4.06363
R15009 CSoutput.n261 CSoutput.t4 4.06363
R15010 CSoutput.n260 CSoutput.t32 4.06363
R15011 CSoutput.n260 CSoutput.t36 4.06363
R15012 CSoutput.n258 CSoutput.t39 4.06363
R15013 CSoutput.n258 CSoutput.t22 4.06363
R15014 CSoutput.n256 CSoutput.t5 4.06363
R15015 CSoutput.n256 CSoutput.t26 4.06363
R15016 CSoutput.n254 CSoutput.t23 4.06363
R15017 CSoutput.n254 CSoutput.t30 4.06363
R15018 CSoutput.n253 CSoutput.t10 4.06363
R15019 CSoutput.n253 CSoutput.t31 4.06363
R15020 CSoutput.n94 CSoutput.t9 4.06363
R15021 CSoutput.n94 CSoutput.t11 4.06363
R15022 CSoutput.n95 CSoutput.t143 4.06363
R15023 CSoutput.n95 CSoutput.t21 4.06363
R15024 CSoutput.n97 CSoutput.t138 4.06363
R15025 CSoutput.n97 CSoutput.t19 4.06363
R15026 CSoutput.n99 CSoutput.t3 4.06363
R15027 CSoutput.n99 CSoutput.t137 4.06363
R15028 CSoutput.n86 CSoutput.t142 4.06363
R15029 CSoutput.n86 CSoutput.t27 4.06363
R15030 CSoutput.n87 CSoutput.t28 4.06363
R15031 CSoutput.n87 CSoutput.t18 4.06363
R15032 CSoutput.n89 CSoutput.t13 4.06363
R15033 CSoutput.n89 CSoutput.t34 4.06363
R15034 CSoutput.n91 CSoutput.t1 4.06363
R15035 CSoutput.n91 CSoutput.t35 4.06363
R15036 CSoutput.n79 CSoutput.t7 4.06363
R15037 CSoutput.n79 CSoutput.t16 4.06363
R15038 CSoutput.n80 CSoutput.t136 4.06363
R15039 CSoutput.n80 CSoutput.t38 4.06363
R15040 CSoutput.n82 CSoutput.t29 4.06363
R15041 CSoutput.n82 CSoutput.t8 4.06363
R15042 CSoutput.n84 CSoutput.t20 4.06363
R15043 CSoutput.n84 CSoutput.t15 4.06363
R15044 CSoutput.n44 CSoutput.n43 3.79402
R15045 CSoutput.n49 CSoutput.n48 3.79402
R15046 CSoutput.n323 CSoutput.n307 3.72967
R15047 CSoutput.n371 CSoutput.n355 3.72967
R15048 CSoutput.n373 CSoutput.n372 3.57343
R15049 CSoutput.n372 CSoutput.n324 3.08965
R15050 CSoutput.n321 CSoutput.t69 2.82907
R15051 CSoutput.n321 CSoutput.t60 2.82907
R15052 CSoutput.n319 CSoutput.t50 2.82907
R15053 CSoutput.n319 CSoutput.t123 2.82907
R15054 CSoutput.n317 CSoutput.t62 2.82907
R15055 CSoutput.n317 CSoutput.t66 2.82907
R15056 CSoutput.n315 CSoutput.t61 2.82907
R15057 CSoutput.n315 CSoutput.t135 2.82907
R15058 CSoutput.n313 CSoutput.t81 2.82907
R15059 CSoutput.n313 CSoutput.t53 2.82907
R15060 CSoutput.n311 CSoutput.t44 2.82907
R15061 CSoutput.n311 CSoutput.t110 2.82907
R15062 CSoutput.n309 CSoutput.t71 2.82907
R15063 CSoutput.n309 CSoutput.t75 2.82907
R15064 CSoutput.n308 CSoutput.t52 2.82907
R15065 CSoutput.n308 CSoutput.t124 2.82907
R15066 CSoutput.n305 CSoutput.t108 2.82907
R15067 CSoutput.n305 CSoutput.t91 2.82907
R15068 CSoutput.n303 CSoutput.t90 2.82907
R15069 CSoutput.n303 CSoutput.t94 2.82907
R15070 CSoutput.n301 CSoutput.t43 2.82907
R15071 CSoutput.n301 CSoutput.t107 2.82907
R15072 CSoutput.n299 CSoutput.t105 2.82907
R15073 CSoutput.n299 CSoutput.t86 2.82907
R15074 CSoutput.n297 CSoutput.t122 2.82907
R15075 CSoutput.n297 CSoutput.t42 2.82907
R15076 CSoutput.n295 CSoutput.t41 2.82907
R15077 CSoutput.n295 CSoutput.t114 2.82907
R15078 CSoutput.n293 CSoutput.t51 2.82907
R15079 CSoutput.n293 CSoutput.t121 2.82907
R15080 CSoutput.n292 CSoutput.t131 2.82907
R15081 CSoutput.n292 CSoutput.t40 2.82907
R15082 CSoutput.n290 CSoutput.t47 2.82907
R15083 CSoutput.n290 CSoutput.t70 2.82907
R15084 CSoutput.n288 CSoutput.t58 2.82907
R15085 CSoutput.n288 CSoutput.t83 2.82907
R15086 CSoutput.n286 CSoutput.t93 2.82907
R15087 CSoutput.n286 CSoutput.t103 2.82907
R15088 CSoutput.n284 CSoutput.t80 2.82907
R15089 CSoutput.n284 CSoutput.t120 2.82907
R15090 CSoutput.n282 CSoutput.t97 2.82907
R15091 CSoutput.n282 CSoutput.t74 2.82907
R15092 CSoutput.n280 CSoutput.t64 2.82907
R15093 CSoutput.n280 CSoutput.t82 2.82907
R15094 CSoutput.n278 CSoutput.t73 2.82907
R15095 CSoutput.n278 CSoutput.t78 2.82907
R15096 CSoutput.n277 CSoutput.t79 2.82907
R15097 CSoutput.n277 CSoutput.t134 2.82907
R15098 CSoutput.n356 CSoutput.t92 2.82907
R15099 CSoutput.n356 CSoutput.t117 2.82907
R15100 CSoutput.n357 CSoutput.t63 2.82907
R15101 CSoutput.n357 CSoutput.t77 2.82907
R15102 CSoutput.n359 CSoutput.t84 2.82907
R15103 CSoutput.n359 CSoutput.t102 2.82907
R15104 CSoutput.n361 CSoutput.t118 2.82907
R15105 CSoutput.n361 CSoutput.t89 2.82907
R15106 CSoutput.n363 CSoutput.t96 2.82907
R15107 CSoutput.n363 CSoutput.t130 2.82907
R15108 CSoutput.n365 CSoutput.t46 2.82907
R15109 CSoutput.n365 CSoutput.t67 2.82907
R15110 CSoutput.n367 CSoutput.t88 2.82907
R15111 CSoutput.n367 CSoutput.t113 2.82907
R15112 CSoutput.n369 CSoutput.t126 2.82907
R15113 CSoutput.n369 CSoutput.t54 2.82907
R15114 CSoutput.n340 CSoutput.t57 2.82907
R15115 CSoutput.n340 CSoutput.t49 2.82907
R15116 CSoutput.n341 CSoutput.t45 2.82907
R15117 CSoutput.n341 CSoutput.t133 2.82907
R15118 CSoutput.n343 CSoutput.t132 2.82907
R15119 CSoutput.n343 CSoutput.t56 2.82907
R15120 CSoutput.n345 CSoutput.t55 2.82907
R15121 CSoutput.n345 CSoutput.t101 2.82907
R15122 CSoutput.n347 CSoutput.t98 2.82907
R15123 CSoutput.n347 CSoutput.t129 2.82907
R15124 CSoutput.n349 CSoutput.t127 2.82907
R15125 CSoutput.n349 CSoutput.t119 2.82907
R15126 CSoutput.n351 CSoutput.t112 2.82907
R15127 CSoutput.n351 CSoutput.t99 2.82907
R15128 CSoutput.n353 CSoutput.t100 2.82907
R15129 CSoutput.n353 CSoutput.t128 2.82907
R15130 CSoutput.n325 CSoutput.t65 2.82907
R15131 CSoutput.n325 CSoutput.t106 2.82907
R15132 CSoutput.n326 CSoutput.t104 2.82907
R15133 CSoutput.n326 CSoutput.t85 2.82907
R15134 CSoutput.n328 CSoutput.t111 2.82907
R15135 CSoutput.n328 CSoutput.t76 2.82907
R15136 CSoutput.n330 CSoutput.t95 2.82907
R15137 CSoutput.n330 CSoutput.t125 2.82907
R15138 CSoutput.n332 CSoutput.t59 2.82907
R15139 CSoutput.n332 CSoutput.t109 2.82907
R15140 CSoutput.n334 CSoutput.t48 2.82907
R15141 CSoutput.n334 CSoutput.t116 2.82907
R15142 CSoutput.n336 CSoutput.t115 2.82907
R15143 CSoutput.n336 CSoutput.t72 2.82907
R15144 CSoutput.n338 CSoutput.t87 2.82907
R15145 CSoutput.n338 CSoutput.t68 2.82907
R15146 CSoutput.n75 CSoutput.n1 2.45513
R15147 CSoutput.n193 CSoutput.n191 2.251
R15148 CSoutput.n193 CSoutput.n190 2.251
R15149 CSoutput.n193 CSoutput.n189 2.251
R15150 CSoutput.n193 CSoutput.n188 2.251
R15151 CSoutput.n162 CSoutput.n161 2.251
R15152 CSoutput.n162 CSoutput.n160 2.251
R15153 CSoutput.n162 CSoutput.n159 2.251
R15154 CSoutput.n162 CSoutput.n158 2.251
R15155 CSoutput.n235 CSoutput.n234 2.251
R15156 CSoutput.n200 CSoutput.n198 2.251
R15157 CSoutput.n200 CSoutput.n197 2.251
R15158 CSoutput.n200 CSoutput.n196 2.251
R15159 CSoutput.n218 CSoutput.n200 2.251
R15160 CSoutput.n206 CSoutput.n205 2.251
R15161 CSoutput.n206 CSoutput.n204 2.251
R15162 CSoutput.n206 CSoutput.n203 2.251
R15163 CSoutput.n206 CSoutput.n202 2.251
R15164 CSoutput.n232 CSoutput.n172 2.251
R15165 CSoutput.n227 CSoutput.n225 2.251
R15166 CSoutput.n227 CSoutput.n224 2.251
R15167 CSoutput.n227 CSoutput.n223 2.251
R15168 CSoutput.n227 CSoutput.n222 2.251
R15169 CSoutput.n128 CSoutput.n127 2.251
R15170 CSoutput.n128 CSoutput.n126 2.251
R15171 CSoutput.n128 CSoutput.n125 2.251
R15172 CSoutput.n128 CSoutput.n124 2.251
R15173 CSoutput.n245 CSoutput.n244 2.251
R15174 CSoutput.n162 CSoutput.n142 2.2505
R15175 CSoutput.n157 CSoutput.n142 2.2505
R15176 CSoutput.n155 CSoutput.n142 2.2505
R15177 CSoutput.n154 CSoutput.n142 2.2505
R15178 CSoutput.n239 CSoutput.n142 2.2505
R15179 CSoutput.n237 CSoutput.n142 2.2505
R15180 CSoutput.n235 CSoutput.n142 2.2505
R15181 CSoutput.n165 CSoutput.n142 2.2505
R15182 CSoutput.n164 CSoutput.n142 2.2505
R15183 CSoutput.n168 CSoutput.n142 2.2505
R15184 CSoutput.n167 CSoutput.n142 2.2505
R15185 CSoutput.n150 CSoutput.n142 2.2505
R15186 CSoutput.n242 CSoutput.n142 2.2505
R15187 CSoutput.n242 CSoutput.n241 2.2505
R15188 CSoutput.n206 CSoutput.n177 2.2505
R15189 CSoutput.n187 CSoutput.n177 2.2505
R15190 CSoutput.n208 CSoutput.n177 2.2505
R15191 CSoutput.n186 CSoutput.n177 2.2505
R15192 CSoutput.n210 CSoutput.n177 2.2505
R15193 CSoutput.n177 CSoutput.n171 2.2505
R15194 CSoutput.n232 CSoutput.n177 2.2505
R15195 CSoutput.n230 CSoutput.n177 2.2505
R15196 CSoutput.n212 CSoutput.n177 2.2505
R15197 CSoutput.n184 CSoutput.n177 2.2505
R15198 CSoutput.n214 CSoutput.n177 2.2505
R15199 CSoutput.n183 CSoutput.n177 2.2505
R15200 CSoutput.n228 CSoutput.n177 2.2505
R15201 CSoutput.n228 CSoutput.n181 2.2505
R15202 CSoutput.n128 CSoutput.n108 2.2505
R15203 CSoutput.n123 CSoutput.n108 2.2505
R15204 CSoutput.n121 CSoutput.n108 2.2505
R15205 CSoutput.n120 CSoutput.n108 2.2505
R15206 CSoutput.n249 CSoutput.n108 2.2505
R15207 CSoutput.n247 CSoutput.n108 2.2505
R15208 CSoutput.n245 CSoutput.n108 2.2505
R15209 CSoutput.n131 CSoutput.n108 2.2505
R15210 CSoutput.n130 CSoutput.n108 2.2505
R15211 CSoutput.n134 CSoutput.n108 2.2505
R15212 CSoutput.n133 CSoutput.n108 2.2505
R15213 CSoutput.n116 CSoutput.n108 2.2505
R15214 CSoutput.n252 CSoutput.n108 2.2505
R15215 CSoutput.n252 CSoutput.n251 2.2505
R15216 CSoutput.n170 CSoutput.n163 2.25024
R15217 CSoutput.n170 CSoutput.n156 2.25024
R15218 CSoutput.n238 CSoutput.n170 2.25024
R15219 CSoutput.n170 CSoutput.n166 2.25024
R15220 CSoutput.n170 CSoutput.n169 2.25024
R15221 CSoutput.n170 CSoutput.n137 2.25024
R15222 CSoutput.n220 CSoutput.n217 2.25024
R15223 CSoutput.n220 CSoutput.n216 2.25024
R15224 CSoutput.n220 CSoutput.n215 2.25024
R15225 CSoutput.n220 CSoutput.n182 2.25024
R15226 CSoutput.n220 CSoutput.n219 2.25024
R15227 CSoutput.n221 CSoutput.n220 2.25024
R15228 CSoutput.n136 CSoutput.n129 2.25024
R15229 CSoutput.n136 CSoutput.n122 2.25024
R15230 CSoutput.n248 CSoutput.n136 2.25024
R15231 CSoutput.n136 CSoutput.n132 2.25024
R15232 CSoutput.n136 CSoutput.n135 2.25024
R15233 CSoutput.n136 CSoutput.n103 2.25024
R15234 CSoutput.n276 CSoutput.n102 1.95131
R15235 CSoutput.n237 CSoutput.n147 1.50111
R15236 CSoutput.n185 CSoutput.n171 1.50111
R15237 CSoutput.n247 CSoutput.n113 1.50111
R15238 CSoutput.n193 CSoutput.n192 1.501
R15239 CSoutput.n200 CSoutput.n199 1.501
R15240 CSoutput.n227 CSoutput.n226 1.501
R15241 CSoutput.n241 CSoutput.n152 1.12536
R15242 CSoutput.n241 CSoutput.n153 1.12536
R15243 CSoutput.n241 CSoutput.n240 1.12536
R15244 CSoutput.n201 CSoutput.n181 1.12536
R15245 CSoutput.n207 CSoutput.n181 1.12536
R15246 CSoutput.n209 CSoutput.n181 1.12536
R15247 CSoutput.n251 CSoutput.n118 1.12536
R15248 CSoutput.n251 CSoutput.n119 1.12536
R15249 CSoutput.n251 CSoutput.n250 1.12536
R15250 CSoutput.n241 CSoutput.n148 1.12536
R15251 CSoutput.n241 CSoutput.n149 1.12536
R15252 CSoutput.n241 CSoutput.n151 1.12536
R15253 CSoutput.n231 CSoutput.n181 1.12536
R15254 CSoutput.n211 CSoutput.n181 1.12536
R15255 CSoutput.n213 CSoutput.n181 1.12536
R15256 CSoutput.n251 CSoutput.n114 1.12536
R15257 CSoutput.n251 CSoutput.n115 1.12536
R15258 CSoutput.n251 CSoutput.n117 1.12536
R15259 CSoutput.n31 CSoutput.n30 0.669944
R15260 CSoutput.n62 CSoutput.n61 0.669944
R15261 CSoutput.n312 CSoutput.n310 0.573776
R15262 CSoutput.n314 CSoutput.n312 0.573776
R15263 CSoutput.n316 CSoutput.n314 0.573776
R15264 CSoutput.n318 CSoutput.n316 0.573776
R15265 CSoutput.n320 CSoutput.n318 0.573776
R15266 CSoutput.n322 CSoutput.n320 0.573776
R15267 CSoutput.n296 CSoutput.n294 0.573776
R15268 CSoutput.n298 CSoutput.n296 0.573776
R15269 CSoutput.n300 CSoutput.n298 0.573776
R15270 CSoutput.n302 CSoutput.n300 0.573776
R15271 CSoutput.n304 CSoutput.n302 0.573776
R15272 CSoutput.n306 CSoutput.n304 0.573776
R15273 CSoutput.n281 CSoutput.n279 0.573776
R15274 CSoutput.n283 CSoutput.n281 0.573776
R15275 CSoutput.n285 CSoutput.n283 0.573776
R15276 CSoutput.n287 CSoutput.n285 0.573776
R15277 CSoutput.n289 CSoutput.n287 0.573776
R15278 CSoutput.n291 CSoutput.n289 0.573776
R15279 CSoutput.n370 CSoutput.n368 0.573776
R15280 CSoutput.n368 CSoutput.n366 0.573776
R15281 CSoutput.n366 CSoutput.n364 0.573776
R15282 CSoutput.n364 CSoutput.n362 0.573776
R15283 CSoutput.n362 CSoutput.n360 0.573776
R15284 CSoutput.n360 CSoutput.n358 0.573776
R15285 CSoutput.n354 CSoutput.n352 0.573776
R15286 CSoutput.n352 CSoutput.n350 0.573776
R15287 CSoutput.n350 CSoutput.n348 0.573776
R15288 CSoutput.n348 CSoutput.n346 0.573776
R15289 CSoutput.n346 CSoutput.n344 0.573776
R15290 CSoutput.n344 CSoutput.n342 0.573776
R15291 CSoutput.n339 CSoutput.n337 0.573776
R15292 CSoutput.n337 CSoutput.n335 0.573776
R15293 CSoutput.n335 CSoutput.n333 0.573776
R15294 CSoutput.n333 CSoutput.n331 0.573776
R15295 CSoutput.n331 CSoutput.n329 0.573776
R15296 CSoutput.n329 CSoutput.n327 0.573776
R15297 CSoutput.n373 CSoutput.n252 0.53442
R15298 CSoutput.n272 CSoutput.n270 0.358259
R15299 CSoutput.n274 CSoutput.n272 0.358259
R15300 CSoutput.n264 CSoutput.n262 0.358259
R15301 CSoutput.n266 CSoutput.n264 0.358259
R15302 CSoutput.n257 CSoutput.n255 0.358259
R15303 CSoutput.n259 CSoutput.n257 0.358259
R15304 CSoutput.n100 CSoutput.n98 0.358259
R15305 CSoutput.n98 CSoutput.n96 0.358259
R15306 CSoutput.n92 CSoutput.n90 0.358259
R15307 CSoutput.n90 CSoutput.n88 0.358259
R15308 CSoutput.n85 CSoutput.n83 0.358259
R15309 CSoutput.n83 CSoutput.n81 0.358259
R15310 CSoutput.n21 CSoutput.n20 0.169105
R15311 CSoutput.n21 CSoutput.n16 0.169105
R15312 CSoutput.n26 CSoutput.n16 0.169105
R15313 CSoutput.n27 CSoutput.n26 0.169105
R15314 CSoutput.n27 CSoutput.n14 0.169105
R15315 CSoutput.n32 CSoutput.n14 0.169105
R15316 CSoutput.n33 CSoutput.n32 0.169105
R15317 CSoutput.n34 CSoutput.n33 0.169105
R15318 CSoutput.n34 CSoutput.n12 0.169105
R15319 CSoutput.n39 CSoutput.n12 0.169105
R15320 CSoutput.n40 CSoutput.n39 0.169105
R15321 CSoutput.n40 CSoutput.n10 0.169105
R15322 CSoutput.n45 CSoutput.n10 0.169105
R15323 CSoutput.n46 CSoutput.n45 0.169105
R15324 CSoutput.n47 CSoutput.n46 0.169105
R15325 CSoutput.n47 CSoutput.n8 0.169105
R15326 CSoutput.n52 CSoutput.n8 0.169105
R15327 CSoutput.n53 CSoutput.n52 0.169105
R15328 CSoutput.n53 CSoutput.n6 0.169105
R15329 CSoutput.n58 CSoutput.n6 0.169105
R15330 CSoutput.n59 CSoutput.n58 0.169105
R15331 CSoutput.n60 CSoutput.n59 0.169105
R15332 CSoutput.n60 CSoutput.n4 0.169105
R15333 CSoutput.n66 CSoutput.n4 0.169105
R15334 CSoutput.n67 CSoutput.n66 0.169105
R15335 CSoutput.n68 CSoutput.n67 0.169105
R15336 CSoutput.n68 CSoutput.n2 0.169105
R15337 CSoutput.n73 CSoutput.n2 0.169105
R15338 CSoutput.n74 CSoutput.n73 0.169105
R15339 CSoutput.n74 CSoutput.n0 0.169105
R15340 CSoutput.n78 CSoutput.n0 0.169105
R15341 CSoutput.n195 CSoutput.n194 0.0910737
R15342 CSoutput.n246 CSoutput.n243 0.0723685
R15343 CSoutput.n200 CSoutput.n195 0.0522944
R15344 CSoutput.n243 CSoutput.n242 0.0499135
R15345 CSoutput.n194 CSoutput.n193 0.0499135
R15346 CSoutput.n228 CSoutput.n227 0.0464294
R15347 CSoutput.n236 CSoutput.n233 0.0391444
R15348 CSoutput.n195 CSoutput.t155 0.023435
R15349 CSoutput.n243 CSoutput.t146 0.02262
R15350 CSoutput.n194 CSoutput.t149 0.02262
R15351 CSoutput CSoutput.n373 0.0052
R15352 CSoutput.n165 CSoutput.n148 0.00365111
R15353 CSoutput.n168 CSoutput.n149 0.00365111
R15354 CSoutput.n151 CSoutput.n150 0.00365111
R15355 CSoutput.n193 CSoutput.n152 0.00365111
R15356 CSoutput.n157 CSoutput.n153 0.00365111
R15357 CSoutput.n240 CSoutput.n154 0.00365111
R15358 CSoutput.n231 CSoutput.n230 0.00365111
R15359 CSoutput.n211 CSoutput.n184 0.00365111
R15360 CSoutput.n213 CSoutput.n183 0.00365111
R15361 CSoutput.n201 CSoutput.n200 0.00365111
R15362 CSoutput.n207 CSoutput.n187 0.00365111
R15363 CSoutput.n209 CSoutput.n186 0.00365111
R15364 CSoutput.n131 CSoutput.n114 0.00365111
R15365 CSoutput.n134 CSoutput.n115 0.00365111
R15366 CSoutput.n117 CSoutput.n116 0.00365111
R15367 CSoutput.n227 CSoutput.n118 0.00365111
R15368 CSoutput.n123 CSoutput.n119 0.00365111
R15369 CSoutput.n250 CSoutput.n120 0.00365111
R15370 CSoutput.n162 CSoutput.n152 0.00340054
R15371 CSoutput.n155 CSoutput.n153 0.00340054
R15372 CSoutput.n240 CSoutput.n239 0.00340054
R15373 CSoutput.n235 CSoutput.n148 0.00340054
R15374 CSoutput.n164 CSoutput.n149 0.00340054
R15375 CSoutput.n167 CSoutput.n151 0.00340054
R15376 CSoutput.n206 CSoutput.n201 0.00340054
R15377 CSoutput.n208 CSoutput.n207 0.00340054
R15378 CSoutput.n210 CSoutput.n209 0.00340054
R15379 CSoutput.n232 CSoutput.n231 0.00340054
R15380 CSoutput.n212 CSoutput.n211 0.00340054
R15381 CSoutput.n214 CSoutput.n213 0.00340054
R15382 CSoutput.n128 CSoutput.n118 0.00340054
R15383 CSoutput.n121 CSoutput.n119 0.00340054
R15384 CSoutput.n250 CSoutput.n249 0.00340054
R15385 CSoutput.n245 CSoutput.n114 0.00340054
R15386 CSoutput.n130 CSoutput.n115 0.00340054
R15387 CSoutput.n133 CSoutput.n117 0.00340054
R15388 CSoutput.n163 CSoutput.n157 0.00252698
R15389 CSoutput.n156 CSoutput.n154 0.00252698
R15390 CSoutput.n238 CSoutput.n237 0.00252698
R15391 CSoutput.n166 CSoutput.n164 0.00252698
R15392 CSoutput.n169 CSoutput.n167 0.00252698
R15393 CSoutput.n242 CSoutput.n137 0.00252698
R15394 CSoutput.n163 CSoutput.n162 0.00252698
R15395 CSoutput.n156 CSoutput.n155 0.00252698
R15396 CSoutput.n239 CSoutput.n238 0.00252698
R15397 CSoutput.n166 CSoutput.n165 0.00252698
R15398 CSoutput.n169 CSoutput.n168 0.00252698
R15399 CSoutput.n150 CSoutput.n137 0.00252698
R15400 CSoutput.n217 CSoutput.n187 0.00252698
R15401 CSoutput.n216 CSoutput.n186 0.00252698
R15402 CSoutput.n215 CSoutput.n171 0.00252698
R15403 CSoutput.n212 CSoutput.n182 0.00252698
R15404 CSoutput.n219 CSoutput.n214 0.00252698
R15405 CSoutput.n228 CSoutput.n221 0.00252698
R15406 CSoutput.n217 CSoutput.n206 0.00252698
R15407 CSoutput.n216 CSoutput.n208 0.00252698
R15408 CSoutput.n215 CSoutput.n210 0.00252698
R15409 CSoutput.n230 CSoutput.n182 0.00252698
R15410 CSoutput.n219 CSoutput.n184 0.00252698
R15411 CSoutput.n221 CSoutput.n183 0.00252698
R15412 CSoutput.n129 CSoutput.n123 0.00252698
R15413 CSoutput.n122 CSoutput.n120 0.00252698
R15414 CSoutput.n248 CSoutput.n247 0.00252698
R15415 CSoutput.n132 CSoutput.n130 0.00252698
R15416 CSoutput.n135 CSoutput.n133 0.00252698
R15417 CSoutput.n252 CSoutput.n103 0.00252698
R15418 CSoutput.n129 CSoutput.n128 0.00252698
R15419 CSoutput.n122 CSoutput.n121 0.00252698
R15420 CSoutput.n249 CSoutput.n248 0.00252698
R15421 CSoutput.n132 CSoutput.n131 0.00252698
R15422 CSoutput.n135 CSoutput.n134 0.00252698
R15423 CSoutput.n116 CSoutput.n103 0.00252698
R15424 CSoutput.n237 CSoutput.n236 0.0020275
R15425 CSoutput.n236 CSoutput.n235 0.0020275
R15426 CSoutput.n233 CSoutput.n171 0.0020275
R15427 CSoutput.n233 CSoutput.n232 0.0020275
R15428 CSoutput.n247 CSoutput.n246 0.0020275
R15429 CSoutput.n246 CSoutput.n245 0.0020275
R15430 CSoutput.n147 CSoutput.n146 0.00166668
R15431 CSoutput.n229 CSoutput.n185 0.00166668
R15432 CSoutput.n113 CSoutput.n112 0.00166668
R15433 CSoutput.n251 CSoutput.n113 0.00133328
R15434 CSoutput.n185 CSoutput.n181 0.00133328
R15435 CSoutput.n241 CSoutput.n147 0.00133328
R15436 CSoutput.n244 CSoutput.n136 0.001
R15437 CSoutput.n222 CSoutput.n136 0.001
R15438 CSoutput.n124 CSoutput.n104 0.001
R15439 CSoutput.n223 CSoutput.n104 0.001
R15440 CSoutput.n125 CSoutput.n105 0.001
R15441 CSoutput.n224 CSoutput.n105 0.001
R15442 CSoutput.n126 CSoutput.n106 0.001
R15443 CSoutput.n225 CSoutput.n106 0.001
R15444 CSoutput.n127 CSoutput.n107 0.001
R15445 CSoutput.n226 CSoutput.n107 0.001
R15446 CSoutput.n220 CSoutput.n172 0.001
R15447 CSoutput.n220 CSoutput.n218 0.001
R15448 CSoutput.n202 CSoutput.n173 0.001
R15449 CSoutput.n196 CSoutput.n173 0.001
R15450 CSoutput.n203 CSoutput.n174 0.001
R15451 CSoutput.n197 CSoutput.n174 0.001
R15452 CSoutput.n204 CSoutput.n175 0.001
R15453 CSoutput.n198 CSoutput.n175 0.001
R15454 CSoutput.n205 CSoutput.n176 0.001
R15455 CSoutput.n199 CSoutput.n176 0.001
R15456 CSoutput.n234 CSoutput.n170 0.001
R15457 CSoutput.n188 CSoutput.n170 0.001
R15458 CSoutput.n158 CSoutput.n138 0.001
R15459 CSoutput.n189 CSoutput.n138 0.001
R15460 CSoutput.n159 CSoutput.n139 0.001
R15461 CSoutput.n190 CSoutput.n139 0.001
R15462 CSoutput.n160 CSoutput.n140 0.001
R15463 CSoutput.n191 CSoutput.n140 0.001
R15464 CSoutput.n161 CSoutput.n141 0.001
R15465 CSoutput.n192 CSoutput.n141 0.001
R15466 CSoutput.n192 CSoutput.n142 0.001
R15467 CSoutput.n191 CSoutput.n143 0.001
R15468 CSoutput.n190 CSoutput.n144 0.001
R15469 CSoutput.n189 CSoutput.t164 0.001
R15470 CSoutput.n188 CSoutput.n145 0.001
R15471 CSoutput.n161 CSoutput.n143 0.001
R15472 CSoutput.n160 CSoutput.n144 0.001
R15473 CSoutput.n159 CSoutput.t164 0.001
R15474 CSoutput.n158 CSoutput.n145 0.001
R15475 CSoutput.n234 CSoutput.n146 0.001
R15476 CSoutput.n199 CSoutput.n177 0.001
R15477 CSoutput.n198 CSoutput.n178 0.001
R15478 CSoutput.n197 CSoutput.n179 0.001
R15479 CSoutput.n196 CSoutput.t144 0.001
R15480 CSoutput.n218 CSoutput.n180 0.001
R15481 CSoutput.n205 CSoutput.n178 0.001
R15482 CSoutput.n204 CSoutput.n179 0.001
R15483 CSoutput.n203 CSoutput.t144 0.001
R15484 CSoutput.n202 CSoutput.n180 0.001
R15485 CSoutput.n229 CSoutput.n172 0.001
R15486 CSoutput.n226 CSoutput.n108 0.001
R15487 CSoutput.n225 CSoutput.n109 0.001
R15488 CSoutput.n224 CSoutput.n110 0.001
R15489 CSoutput.n223 CSoutput.t153 0.001
R15490 CSoutput.n222 CSoutput.n111 0.001
R15491 CSoutput.n127 CSoutput.n109 0.001
R15492 CSoutput.n126 CSoutput.n110 0.001
R15493 CSoutput.n125 CSoutput.t153 0.001
R15494 CSoutput.n124 CSoutput.n111 0.001
R15495 CSoutput.n244 CSoutput.n112 0.001
R15496 a_n1986_8322.n2 a_n1986_8322.t10 74.6477
R15497 a_n1986_8322.t0 a_n1986_8322.n0 74.6477
R15498 a_n1986_8322.n1 a_n1986_8322.t18 74.6474
R15499 a_n1986_8322.n0 a_n1986_8322.t12 74.2899
R15500 a_n1986_8322.n0 a_n1986_8322.t17 74.2899
R15501 a_n1986_8322.n3 a_n1986_8322.t4 74.2899
R15502 a_n1986_8322.n6 a_n1986_8322.t14 74.2899
R15503 a_n1986_8322.n10 a_n1986_8322.t13 74.2899
R15504 a_n1986_8322.n0 a_n1986_8322.n13 70.6783
R15505 a_n1986_8322.n0 a_n1986_8322.n12 70.6783
R15506 a_n1986_8322.n1 a_n1986_8322.n4 70.6783
R15507 a_n1986_8322.n1 a_n1986_8322.n5 70.6783
R15508 a_n1986_8322.n2 a_n1986_8322.n8 70.6783
R15509 a_n1986_8322.n2 a_n1986_8322.n9 70.6783
R15510 a_n1986_8322.n11 a_n1986_8322.n10 22.7556
R15511 a_n1986_8322.n7 a_n1986_8322.t8 9.96389
R15512 a_n1986_8322.n3 a_n1986_8322.n11 6.2408
R15513 a_n1986_8322.n7 a_n1986_8322.n6 5.83671
R15514 a_n1986_8322.n11 a_n1986_8322.n7 5.3452
R15515 a_n1986_8322.n13 a_n1986_8322.t15 3.61217
R15516 a_n1986_8322.n13 a_n1986_8322.t16 3.61217
R15517 a_n1986_8322.n12 a_n1986_8322.t3 3.61217
R15518 a_n1986_8322.n12 a_n1986_8322.t9 3.61217
R15519 a_n1986_8322.n4 a_n1986_8322.t7 3.61217
R15520 a_n1986_8322.n4 a_n1986_8322.t2 3.61217
R15521 a_n1986_8322.n5 a_n1986_8322.t1 3.61217
R15522 a_n1986_8322.n5 a_n1986_8322.t20 3.61217
R15523 a_n1986_8322.n8 a_n1986_8322.t19 3.61217
R15524 a_n1986_8322.n8 a_n1986_8322.t11 3.61217
R15525 a_n1986_8322.n9 a_n1986_8322.t5 3.61217
R15526 a_n1986_8322.n9 a_n1986_8322.t6 3.61217
R15527 a_n1986_8322.n0 a_n1986_8322.n3 1.17507
R15528 a_n1986_8322.n10 a_n1986_8322.n2 0.716017
R15529 a_n1986_8322.n6 a_n1986_8322.n1 0.716017
R15530 a_n5644_8799.n95 a_n5644_8799.t65 485.149
R15531 a_n5644_8799.n102 a_n5644_8799.t68 485.149
R15532 a_n5644_8799.n110 a_n5644_8799.t34 485.149
R15533 a_n5644_8799.n71 a_n5644_8799.t49 485.149
R15534 a_n5644_8799.n78 a_n5644_8799.t54 485.149
R15535 a_n5644_8799.n86 a_n5644_8799.t35 485.149
R15536 a_n5644_8799.n20 a_n5644_8799.t56 485.135
R15537 a_n5644_8799.n99 a_n5644_8799.t55 464.166
R15538 a_n5644_8799.n93 a_n5644_8799.t42 464.166
R15539 a_n5644_8799.n98 a_n5644_8799.t72 464.166
R15540 a_n5644_8799.n97 a_n5644_8799.t57 464.166
R15541 a_n5644_8799.n94 a_n5644_8799.t47 464.166
R15542 a_n5644_8799.n96 a_n5644_8799.t74 464.166
R15543 a_n5644_8799.n25 a_n5644_8799.t60 485.135
R15544 a_n5644_8799.n106 a_n5644_8799.t59 464.166
R15545 a_n5644_8799.n100 a_n5644_8799.t51 464.166
R15546 a_n5644_8799.n105 a_n5644_8799.t76 464.166
R15547 a_n5644_8799.n104 a_n5644_8799.t63 464.166
R15548 a_n5644_8799.n101 a_n5644_8799.t52 464.166
R15549 a_n5644_8799.n103 a_n5644_8799.t32 464.166
R15550 a_n5644_8799.n30 a_n5644_8799.t78 485.135
R15551 a_n5644_8799.n114 a_n5644_8799.t40 464.166
R15552 a_n5644_8799.n108 a_n5644_8799.t61 464.166
R15553 a_n5644_8799.n113 a_n5644_8799.t33 464.166
R15554 a_n5644_8799.n112 a_n5644_8799.t69 464.166
R15555 a_n5644_8799.n109 a_n5644_8799.t46 464.166
R15556 a_n5644_8799.n111 a_n5644_8799.t66 464.166
R15557 a_n5644_8799.n72 a_n5644_8799.t58 464.166
R15558 a_n5644_8799.n73 a_n5644_8799.t73 464.166
R15559 a_n5644_8799.n74 a_n5644_8799.t38 464.166
R15560 a_n5644_8799.n75 a_n5644_8799.t48 464.166
R15561 a_n5644_8799.n70 a_n5644_8799.t71 464.166
R15562 a_n5644_8799.n76 a_n5644_8799.t37 464.166
R15563 a_n5644_8799.n79 a_n5644_8799.t64 464.166
R15564 a_n5644_8799.n80 a_n5644_8799.t77 464.166
R15565 a_n5644_8799.n81 a_n5644_8799.t45 464.166
R15566 a_n5644_8799.n82 a_n5644_8799.t53 464.166
R15567 a_n5644_8799.n77 a_n5644_8799.t75 464.166
R15568 a_n5644_8799.n83 a_n5644_8799.t41 464.166
R15569 a_n5644_8799.n87 a_n5644_8799.t67 464.166
R15570 a_n5644_8799.n88 a_n5644_8799.t44 464.166
R15571 a_n5644_8799.n89 a_n5644_8799.t70 464.166
R15572 a_n5644_8799.n90 a_n5644_8799.t50 464.166
R15573 a_n5644_8799.n85 a_n5644_8799.t62 464.166
R15574 a_n5644_8799.n91 a_n5644_8799.t39 464.166
R15575 a_n5644_8799.n16 a_n5644_8799.n24 72.3034
R15576 a_n5644_8799.n24 a_n5644_8799.n94 16.6962
R15577 a_n5644_8799.n23 a_n5644_8799.n16 77.6622
R15578 a_n5644_8799.n97 a_n5644_8799.n23 5.97853
R15579 a_n5644_8799.n22 a_n5644_8799.n15 77.6622
R15580 a_n5644_8799.n15 a_n5644_8799.n21 72.3034
R15581 a_n5644_8799.n99 a_n5644_8799.n20 20.9683
R15582 a_n5644_8799.n17 a_n5644_8799.n20 70.1674
R15583 a_n5644_8799.n13 a_n5644_8799.n29 72.3034
R15584 a_n5644_8799.n29 a_n5644_8799.n101 16.6962
R15585 a_n5644_8799.n28 a_n5644_8799.n13 77.6622
R15586 a_n5644_8799.n104 a_n5644_8799.n28 5.97853
R15587 a_n5644_8799.n27 a_n5644_8799.n12 77.6622
R15588 a_n5644_8799.n12 a_n5644_8799.n26 72.3034
R15589 a_n5644_8799.n106 a_n5644_8799.n25 20.9683
R15590 a_n5644_8799.n14 a_n5644_8799.n25 70.1674
R15591 a_n5644_8799.n10 a_n5644_8799.n34 72.3034
R15592 a_n5644_8799.n34 a_n5644_8799.n109 16.6962
R15593 a_n5644_8799.n33 a_n5644_8799.n10 77.6622
R15594 a_n5644_8799.n112 a_n5644_8799.n33 5.97853
R15595 a_n5644_8799.n32 a_n5644_8799.n9 77.6622
R15596 a_n5644_8799.n9 a_n5644_8799.n31 72.3034
R15597 a_n5644_8799.n114 a_n5644_8799.n30 20.9683
R15598 a_n5644_8799.n11 a_n5644_8799.n30 70.1674
R15599 a_n5644_8799.n7 a_n5644_8799.n39 70.1674
R15600 a_n5644_8799.n76 a_n5644_8799.n39 20.9683
R15601 a_n5644_8799.n38 a_n5644_8799.n7 72.3034
R15602 a_n5644_8799.n38 a_n5644_8799.n70 16.6962
R15603 a_n5644_8799.n6 a_n5644_8799.n37 77.6622
R15604 a_n5644_8799.n75 a_n5644_8799.n37 5.97853
R15605 a_n5644_8799.n36 a_n5644_8799.n6 77.6622
R15606 a_n5644_8799.n35 a_n5644_8799.n73 16.6962
R15607 a_n5644_8799.n35 a_n5644_8799.n8 72.3034
R15608 a_n5644_8799.n4 a_n5644_8799.n44 70.1674
R15609 a_n5644_8799.n83 a_n5644_8799.n44 20.9683
R15610 a_n5644_8799.n43 a_n5644_8799.n4 72.3034
R15611 a_n5644_8799.n43 a_n5644_8799.n77 16.6962
R15612 a_n5644_8799.n3 a_n5644_8799.n42 77.6622
R15613 a_n5644_8799.n82 a_n5644_8799.n42 5.97853
R15614 a_n5644_8799.n41 a_n5644_8799.n3 77.6622
R15615 a_n5644_8799.n40 a_n5644_8799.n80 16.6962
R15616 a_n5644_8799.n40 a_n5644_8799.n5 72.3034
R15617 a_n5644_8799.n1 a_n5644_8799.n49 70.1674
R15618 a_n5644_8799.n91 a_n5644_8799.n49 20.9683
R15619 a_n5644_8799.n48 a_n5644_8799.n1 72.3034
R15620 a_n5644_8799.n48 a_n5644_8799.n85 16.6962
R15621 a_n5644_8799.n0 a_n5644_8799.n47 77.6622
R15622 a_n5644_8799.n90 a_n5644_8799.n47 5.97853
R15623 a_n5644_8799.n46 a_n5644_8799.n0 77.6622
R15624 a_n5644_8799.n45 a_n5644_8799.n88 16.6962
R15625 a_n5644_8799.n45 a_n5644_8799.n2 72.3034
R15626 a_n5644_8799.n18 a_n5644_8799.n50 98.9633
R15627 a_n5644_8799.n19 a_n5644_8799.n119 98.9631
R15628 a_n5644_8799.n19 a_n5644_8799.n120 98.6055
R15629 a_n5644_8799.n18 a_n5644_8799.n52 98.6055
R15630 a_n5644_8799.n18 a_n5644_8799.n51 98.6055
R15631 a_n5644_8799.n121 a_n5644_8799.n19 98.6054
R15632 a_n5644_8799.n55 a_n5644_8799.n53 81.4626
R15633 a_n5644_8799.n63 a_n5644_8799.n61 81.4626
R15634 a_n5644_8799.n59 a_n5644_8799.n57 81.4626
R15635 a_n5644_8799.n66 a_n5644_8799.n65 80.9324
R15636 a_n5644_8799.n68 a_n5644_8799.n67 80.9324
R15637 a_n5644_8799.n69 a_n5644_8799.n56 80.9324
R15638 a_n5644_8799.n55 a_n5644_8799.n54 80.9324
R15639 a_n5644_8799.n63 a_n5644_8799.n62 80.9324
R15640 a_n5644_8799.n64 a_n5644_8799.n60 80.9324
R15641 a_n5644_8799.n59 a_n5644_8799.n58 80.9324
R15642 a_n5644_8799.n16 a_n5644_8799.n95 70.4033
R15643 a_n5644_8799.n13 a_n5644_8799.n102 70.4033
R15644 a_n5644_8799.n10 a_n5644_8799.n110 70.4033
R15645 a_n5644_8799.n71 a_n5644_8799.n8 70.4033
R15646 a_n5644_8799.n78 a_n5644_8799.n5 70.4033
R15647 a_n5644_8799.n86 a_n5644_8799.n2 70.4033
R15648 a_n5644_8799.n98 a_n5644_8799.n97 48.2005
R15649 a_n5644_8799.n105 a_n5644_8799.n104 48.2005
R15650 a_n5644_8799.n113 a_n5644_8799.n112 48.2005
R15651 a_n5644_8799.n75 a_n5644_8799.n74 48.2005
R15652 a_n5644_8799.t36 a_n5644_8799.n39 485.135
R15653 a_n5644_8799.n82 a_n5644_8799.n81 48.2005
R15654 a_n5644_8799.t43 a_n5644_8799.n44 485.135
R15655 a_n5644_8799.n90 a_n5644_8799.n89 48.2005
R15656 a_n5644_8799.t79 a_n5644_8799.n49 485.135
R15657 a_n5644_8799.n21 a_n5644_8799.n93 16.6962
R15658 a_n5644_8799.n96 a_n5644_8799.n24 27.6507
R15659 a_n5644_8799.n26 a_n5644_8799.n100 16.6962
R15660 a_n5644_8799.n103 a_n5644_8799.n29 27.6507
R15661 a_n5644_8799.n31 a_n5644_8799.n108 16.6962
R15662 a_n5644_8799.n111 a_n5644_8799.n34 27.6507
R15663 a_n5644_8799.n76 a_n5644_8799.n38 27.6507
R15664 a_n5644_8799.n83 a_n5644_8799.n43 27.6507
R15665 a_n5644_8799.n91 a_n5644_8799.n48 27.6507
R15666 a_n5644_8799.n22 a_n5644_8799.n93 41.7634
R15667 a_n5644_8799.n27 a_n5644_8799.n100 41.7634
R15668 a_n5644_8799.n32 a_n5644_8799.n108 41.7634
R15669 a_n5644_8799.n73 a_n5644_8799.n36 41.7634
R15670 a_n5644_8799.n80 a_n5644_8799.n41 41.7634
R15671 a_n5644_8799.n88 a_n5644_8799.n46 41.7634
R15672 a_n5644_8799.n66 a_n5644_8799.n64 33.5285
R15673 a_n5644_8799.n96 a_n5644_8799.n95 20.9576
R15674 a_n5644_8799.n103 a_n5644_8799.n102 20.9576
R15675 a_n5644_8799.n111 a_n5644_8799.n110 20.9576
R15676 a_n5644_8799.n72 a_n5644_8799.n71 20.9576
R15677 a_n5644_8799.n79 a_n5644_8799.n78 20.9576
R15678 a_n5644_8799.n87 a_n5644_8799.n86 20.9576
R15679 a_n5644_8799.n22 a_n5644_8799.n98 5.97853
R15680 a_n5644_8799.n23 a_n5644_8799.n94 41.7634
R15681 a_n5644_8799.n27 a_n5644_8799.n105 5.97853
R15682 a_n5644_8799.n28 a_n5644_8799.n101 41.7634
R15683 a_n5644_8799.n32 a_n5644_8799.n113 5.97853
R15684 a_n5644_8799.n33 a_n5644_8799.n109 41.7634
R15685 a_n5644_8799.n74 a_n5644_8799.n36 5.97853
R15686 a_n5644_8799.n70 a_n5644_8799.n37 41.7634
R15687 a_n5644_8799.n81 a_n5644_8799.n41 5.97853
R15688 a_n5644_8799.n77 a_n5644_8799.n42 41.7634
R15689 a_n5644_8799.n89 a_n5644_8799.n46 5.97853
R15690 a_n5644_8799.n85 a_n5644_8799.n47 41.7634
R15691 a_n5644_8799.n19 a_n5644_8799.n118 31.2868
R15692 a_n5644_8799.n117 a_n5644_8799.n69 12.3339
R15693 a_n5644_8799.n118 a_n5644_8799.n117 11.4887
R15694 a_n5644_8799.n99 a_n5644_8799.n21 27.6507
R15695 a_n5644_8799.n106 a_n5644_8799.n26 27.6507
R15696 a_n5644_8799.n114 a_n5644_8799.n31 27.6507
R15697 a_n5644_8799.n35 a_n5644_8799.n72 27.6507
R15698 a_n5644_8799.n40 a_n5644_8799.n79 27.6507
R15699 a_n5644_8799.n45 a_n5644_8799.n87 27.6507
R15700 a_n5644_8799.n118 a_n5644_8799.n18 17.8783
R15701 a_n5644_8799.n107 a_n5644_8799.n17 9.05164
R15702 a_n5644_8799.n84 a_n5644_8799.n7 9.05164
R15703 a_n5644_8799.n116 a_n5644_8799.n92 6.90118
R15704 a_n5644_8799.n116 a_n5644_8799.n115 6.48163
R15705 a_n5644_8799.n107 a_n5644_8799.n14 4.94368
R15706 a_n5644_8799.n115 a_n5644_8799.n11 4.94368
R15707 a_n5644_8799.n84 a_n5644_8799.n4 4.94368
R15708 a_n5644_8799.n92 a_n5644_8799.n1 4.94368
R15709 a_n5644_8799.n115 a_n5644_8799.n107 4.10845
R15710 a_n5644_8799.n92 a_n5644_8799.n84 4.10845
R15711 a_n5644_8799.n119 a_n5644_8799.t1 3.61217
R15712 a_n5644_8799.n119 a_n5644_8799.t25 3.61217
R15713 a_n5644_8799.n120 a_n5644_8799.t30 3.61217
R15714 a_n5644_8799.n120 a_n5644_8799.t6 3.61217
R15715 a_n5644_8799.n52 a_n5644_8799.t13 3.61217
R15716 a_n5644_8799.n52 a_n5644_8799.t12 3.61217
R15717 a_n5644_8799.n51 a_n5644_8799.t5 3.61217
R15718 a_n5644_8799.n51 a_n5644_8799.t26 3.61217
R15719 a_n5644_8799.n50 a_n5644_8799.t16 3.61217
R15720 a_n5644_8799.n50 a_n5644_8799.t2 3.61217
R15721 a_n5644_8799.n121 a_n5644_8799.t17 3.61217
R15722 a_n5644_8799.t0 a_n5644_8799.n121 3.61217
R15723 a_n5644_8799.n117 a_n5644_8799.n116 3.4105
R15724 a_n5644_8799.n65 a_n5644_8799.t24 2.82907
R15725 a_n5644_8799.n65 a_n5644_8799.t10 2.82907
R15726 a_n5644_8799.n67 a_n5644_8799.t11 2.82907
R15727 a_n5644_8799.n67 a_n5644_8799.t14 2.82907
R15728 a_n5644_8799.n56 a_n5644_8799.t7 2.82907
R15729 a_n5644_8799.n56 a_n5644_8799.t31 2.82907
R15730 a_n5644_8799.n54 a_n5644_8799.t8 2.82907
R15731 a_n5644_8799.n54 a_n5644_8799.t19 2.82907
R15732 a_n5644_8799.n53 a_n5644_8799.t22 2.82907
R15733 a_n5644_8799.n53 a_n5644_8799.t15 2.82907
R15734 a_n5644_8799.n61 a_n5644_8799.t18 2.82907
R15735 a_n5644_8799.n61 a_n5644_8799.t4 2.82907
R15736 a_n5644_8799.n62 a_n5644_8799.t20 2.82907
R15737 a_n5644_8799.n62 a_n5644_8799.t23 2.82907
R15738 a_n5644_8799.n60 a_n5644_8799.t28 2.82907
R15739 a_n5644_8799.n60 a_n5644_8799.t9 2.82907
R15740 a_n5644_8799.n58 a_n5644_8799.t27 2.82907
R15741 a_n5644_8799.n58 a_n5644_8799.t3 2.82907
R15742 a_n5644_8799.n57 a_n5644_8799.t21 2.82907
R15743 a_n5644_8799.n57 a_n5644_8799.t29 2.82907
R15744 a_n5644_8799.n16 a_n5644_8799.n15 1.13686
R15745 a_n5644_8799.n13 a_n5644_8799.n12 1.13686
R15746 a_n5644_8799.n10 a_n5644_8799.n9 1.13686
R15747 a_n5644_8799.n7 a_n5644_8799.n6 1.13686
R15748 a_n5644_8799.n4 a_n5644_8799.n3 1.13686
R15749 a_n5644_8799.n1 a_n5644_8799.n0 1.13686
R15750 a_n5644_8799.n0 a_n5644_8799.n2 0.568682
R15751 a_n5644_8799.n3 a_n5644_8799.n5 0.568682
R15752 a_n5644_8799.n6 a_n5644_8799.n8 0.568682
R15753 a_n5644_8799.n9 a_n5644_8799.n11 0.568682
R15754 a_n5644_8799.n12 a_n5644_8799.n14 0.568682
R15755 a_n5644_8799.n15 a_n5644_8799.n17 0.568682
R15756 a_n5644_8799.n64 a_n5644_8799.n59 0.530672
R15757 a_n5644_8799.n64 a_n5644_8799.n63 0.530672
R15758 a_n5644_8799.n69 a_n5644_8799.n55 0.530672
R15759 a_n5644_8799.n69 a_n5644_8799.n68 0.530672
R15760 a_n5644_8799.n68 a_n5644_8799.n66 0.530672
R15761 vdd.n291 vdd.n255 756.745
R15762 vdd.n244 vdd.n208 756.745
R15763 vdd.n201 vdd.n165 756.745
R15764 vdd.n154 vdd.n118 756.745
R15765 vdd.n112 vdd.n76 756.745
R15766 vdd.n65 vdd.n29 756.745
R15767 vdd.n1106 vdd.n1070 756.745
R15768 vdd.n1153 vdd.n1117 756.745
R15769 vdd.n1016 vdd.n980 756.745
R15770 vdd.n1063 vdd.n1027 756.745
R15771 vdd.n927 vdd.n891 756.745
R15772 vdd.n974 vdd.n938 756.745
R15773 vdd.n1791 vdd.t112 640.208
R15774 vdd.n755 vdd.t97 640.208
R15775 vdd.n1765 vdd.t138 640.208
R15776 vdd.n747 vdd.t129 640.208
R15777 vdd.n2536 vdd.t80 640.208
R15778 vdd.n2256 vdd.t120 640.208
R15779 vdd.n622 vdd.t101 640.208
R15780 vdd.n2253 vdd.t105 640.208
R15781 vdd.n589 vdd.t109 640.208
R15782 vdd.n817 vdd.t116 640.208
R15783 vdd.n1320 vdd.t76 592.009
R15784 vdd.n1358 vdd.t123 592.009
R15785 vdd.n1254 vdd.t126 592.009
R15786 vdd.n1947 vdd.t72 592.009
R15787 vdd.n1584 vdd.t84 592.009
R15788 vdd.n1544 vdd.t91 592.009
R15789 vdd.n2908 vdd.t135 592.009
R15790 vdd.n405 vdd.t87 592.009
R15791 vdd.n365 vdd.t94 592.009
R15792 vdd.n557 vdd.t65 592.009
R15793 vdd.n2804 vdd.t69 592.009
R15794 vdd.n2711 vdd.t132 592.009
R15795 vdd.n292 vdd.n291 585
R15796 vdd.n290 vdd.n257 585
R15797 vdd.n289 vdd.n288 585
R15798 vdd.n260 vdd.n258 585
R15799 vdd.n283 vdd.n282 585
R15800 vdd.n281 vdd.n280 585
R15801 vdd.n264 vdd.n263 585
R15802 vdd.n275 vdd.n274 585
R15803 vdd.n273 vdd.n272 585
R15804 vdd.n268 vdd.n267 585
R15805 vdd.n245 vdd.n244 585
R15806 vdd.n243 vdd.n210 585
R15807 vdd.n242 vdd.n241 585
R15808 vdd.n213 vdd.n211 585
R15809 vdd.n236 vdd.n235 585
R15810 vdd.n234 vdd.n233 585
R15811 vdd.n217 vdd.n216 585
R15812 vdd.n228 vdd.n227 585
R15813 vdd.n226 vdd.n225 585
R15814 vdd.n221 vdd.n220 585
R15815 vdd.n202 vdd.n201 585
R15816 vdd.n200 vdd.n167 585
R15817 vdd.n199 vdd.n198 585
R15818 vdd.n170 vdd.n168 585
R15819 vdd.n193 vdd.n192 585
R15820 vdd.n191 vdd.n190 585
R15821 vdd.n174 vdd.n173 585
R15822 vdd.n185 vdd.n184 585
R15823 vdd.n183 vdd.n182 585
R15824 vdd.n178 vdd.n177 585
R15825 vdd.n155 vdd.n154 585
R15826 vdd.n153 vdd.n120 585
R15827 vdd.n152 vdd.n151 585
R15828 vdd.n123 vdd.n121 585
R15829 vdd.n146 vdd.n145 585
R15830 vdd.n144 vdd.n143 585
R15831 vdd.n127 vdd.n126 585
R15832 vdd.n138 vdd.n137 585
R15833 vdd.n136 vdd.n135 585
R15834 vdd.n131 vdd.n130 585
R15835 vdd.n113 vdd.n112 585
R15836 vdd.n111 vdd.n78 585
R15837 vdd.n110 vdd.n109 585
R15838 vdd.n81 vdd.n79 585
R15839 vdd.n104 vdd.n103 585
R15840 vdd.n102 vdd.n101 585
R15841 vdd.n85 vdd.n84 585
R15842 vdd.n96 vdd.n95 585
R15843 vdd.n94 vdd.n93 585
R15844 vdd.n89 vdd.n88 585
R15845 vdd.n66 vdd.n65 585
R15846 vdd.n64 vdd.n31 585
R15847 vdd.n63 vdd.n62 585
R15848 vdd.n34 vdd.n32 585
R15849 vdd.n57 vdd.n56 585
R15850 vdd.n55 vdd.n54 585
R15851 vdd.n38 vdd.n37 585
R15852 vdd.n49 vdd.n48 585
R15853 vdd.n47 vdd.n46 585
R15854 vdd.n42 vdd.n41 585
R15855 vdd.n1107 vdd.n1106 585
R15856 vdd.n1105 vdd.n1072 585
R15857 vdd.n1104 vdd.n1103 585
R15858 vdd.n1075 vdd.n1073 585
R15859 vdd.n1098 vdd.n1097 585
R15860 vdd.n1096 vdd.n1095 585
R15861 vdd.n1079 vdd.n1078 585
R15862 vdd.n1090 vdd.n1089 585
R15863 vdd.n1088 vdd.n1087 585
R15864 vdd.n1083 vdd.n1082 585
R15865 vdd.n1154 vdd.n1153 585
R15866 vdd.n1152 vdd.n1119 585
R15867 vdd.n1151 vdd.n1150 585
R15868 vdd.n1122 vdd.n1120 585
R15869 vdd.n1145 vdd.n1144 585
R15870 vdd.n1143 vdd.n1142 585
R15871 vdd.n1126 vdd.n1125 585
R15872 vdd.n1137 vdd.n1136 585
R15873 vdd.n1135 vdd.n1134 585
R15874 vdd.n1130 vdd.n1129 585
R15875 vdd.n1017 vdd.n1016 585
R15876 vdd.n1015 vdd.n982 585
R15877 vdd.n1014 vdd.n1013 585
R15878 vdd.n985 vdd.n983 585
R15879 vdd.n1008 vdd.n1007 585
R15880 vdd.n1006 vdd.n1005 585
R15881 vdd.n989 vdd.n988 585
R15882 vdd.n1000 vdd.n999 585
R15883 vdd.n998 vdd.n997 585
R15884 vdd.n993 vdd.n992 585
R15885 vdd.n1064 vdd.n1063 585
R15886 vdd.n1062 vdd.n1029 585
R15887 vdd.n1061 vdd.n1060 585
R15888 vdd.n1032 vdd.n1030 585
R15889 vdd.n1055 vdd.n1054 585
R15890 vdd.n1053 vdd.n1052 585
R15891 vdd.n1036 vdd.n1035 585
R15892 vdd.n1047 vdd.n1046 585
R15893 vdd.n1045 vdd.n1044 585
R15894 vdd.n1040 vdd.n1039 585
R15895 vdd.n928 vdd.n927 585
R15896 vdd.n926 vdd.n893 585
R15897 vdd.n925 vdd.n924 585
R15898 vdd.n896 vdd.n894 585
R15899 vdd.n919 vdd.n918 585
R15900 vdd.n917 vdd.n916 585
R15901 vdd.n900 vdd.n899 585
R15902 vdd.n911 vdd.n910 585
R15903 vdd.n909 vdd.n908 585
R15904 vdd.n904 vdd.n903 585
R15905 vdd.n975 vdd.n974 585
R15906 vdd.n973 vdd.n940 585
R15907 vdd.n972 vdd.n971 585
R15908 vdd.n943 vdd.n941 585
R15909 vdd.n966 vdd.n965 585
R15910 vdd.n964 vdd.n963 585
R15911 vdd.n947 vdd.n946 585
R15912 vdd.n958 vdd.n957 585
R15913 vdd.n956 vdd.n955 585
R15914 vdd.n951 vdd.n950 585
R15915 vdd.n3024 vdd.n330 515.122
R15916 vdd.n2906 vdd.n328 515.122
R15917 vdd.n515 vdd.n478 515.122
R15918 vdd.n2842 vdd.n479 515.122
R15919 vdd.n1942 vdd.n865 515.122
R15920 vdd.n1945 vdd.n1944 515.122
R15921 vdd.n1227 vdd.n1191 515.122
R15922 vdd.n1423 vdd.n1192 515.122
R15923 vdd.n269 vdd.t25 329.043
R15924 vdd.n222 vdd.t36 329.043
R15925 vdd.n179 vdd.t21 329.043
R15926 vdd.n132 vdd.t31 329.043
R15927 vdd.n90 vdd.t62 329.043
R15928 vdd.n43 vdd.t4 329.043
R15929 vdd.n1084 vdd.t60 329.043
R15930 vdd.n1131 vdd.t46 329.043
R15931 vdd.n994 vdd.t52 329.043
R15932 vdd.n1041 vdd.t39 329.043
R15933 vdd.n905 vdd.t2 329.043
R15934 vdd.n952 vdd.t61 329.043
R15935 vdd.n1320 vdd.t79 319.788
R15936 vdd.n1358 vdd.t125 319.788
R15937 vdd.n1254 vdd.t128 319.788
R15938 vdd.n1947 vdd.t74 319.788
R15939 vdd.n1584 vdd.t85 319.788
R15940 vdd.n1544 vdd.t92 319.788
R15941 vdd.n2908 vdd.t136 319.788
R15942 vdd.n405 vdd.t89 319.788
R15943 vdd.n365 vdd.t95 319.788
R15944 vdd.n557 vdd.t68 319.788
R15945 vdd.n2804 vdd.t71 319.788
R15946 vdd.n2711 vdd.t134 319.788
R15947 vdd.n1321 vdd.t78 303.69
R15948 vdd.n1359 vdd.t124 303.69
R15949 vdd.n1255 vdd.t127 303.69
R15950 vdd.n1948 vdd.t75 303.69
R15951 vdd.n1585 vdd.t86 303.69
R15952 vdd.n1545 vdd.t93 303.69
R15953 vdd.n2909 vdd.t137 303.69
R15954 vdd.n406 vdd.t90 303.69
R15955 vdd.n366 vdd.t96 303.69
R15956 vdd.n558 vdd.t67 303.69
R15957 vdd.n2805 vdd.t70 303.69
R15958 vdd.n2712 vdd.t133 303.69
R15959 vdd.n2479 vdd.n703 297.074
R15960 vdd.n2672 vdd.n599 297.074
R15961 vdd.n2609 vdd.n596 297.074
R15962 vdd.n2402 vdd.n704 297.074
R15963 vdd.n2217 vdd.n744 297.074
R15964 vdd.n2148 vdd.n2147 297.074
R15965 vdd.n1894 vdd.n840 297.074
R15966 vdd.n1990 vdd.n838 297.074
R15967 vdd.n2588 vdd.n597 297.074
R15968 vdd.n2675 vdd.n2674 297.074
R15969 vdd.n2251 vdd.n705 297.074
R15970 vdd.n2477 vdd.n706 297.074
R15971 vdd.n2145 vdd.n753 297.074
R15972 vdd.n751 vdd.n726 297.074
R15973 vdd.n1831 vdd.n841 297.074
R15974 vdd.n1988 vdd.n842 297.074
R15975 vdd.n2590 vdd.n597 185
R15976 vdd.n2673 vdd.n597 185
R15977 vdd.n2592 vdd.n2591 185
R15978 vdd.n2591 vdd.n595 185
R15979 vdd.n2593 vdd.n629 185
R15980 vdd.n2603 vdd.n629 185
R15981 vdd.n2594 vdd.n638 185
R15982 vdd.n638 vdd.n636 185
R15983 vdd.n2596 vdd.n2595 185
R15984 vdd.n2597 vdd.n2596 185
R15985 vdd.n2549 vdd.n637 185
R15986 vdd.n637 vdd.n633 185
R15987 vdd.n2548 vdd.n2547 185
R15988 vdd.n2547 vdd.n2546 185
R15989 vdd.n640 vdd.n639 185
R15990 vdd.n641 vdd.n640 185
R15991 vdd.n2539 vdd.n2538 185
R15992 vdd.n2540 vdd.n2539 185
R15993 vdd.n2535 vdd.n650 185
R15994 vdd.n650 vdd.n647 185
R15995 vdd.n2534 vdd.n2533 185
R15996 vdd.n2533 vdd.n2532 185
R15997 vdd.n652 vdd.n651 185
R15998 vdd.n660 vdd.n652 185
R15999 vdd.n2525 vdd.n2524 185
R16000 vdd.n2526 vdd.n2525 185
R16001 vdd.n2523 vdd.n661 185
R16002 vdd.n2374 vdd.n661 185
R16003 vdd.n2522 vdd.n2521 185
R16004 vdd.n2521 vdd.n2520 185
R16005 vdd.n663 vdd.n662 185
R16006 vdd.n664 vdd.n663 185
R16007 vdd.n2513 vdd.n2512 185
R16008 vdd.n2514 vdd.n2513 185
R16009 vdd.n2511 vdd.n673 185
R16010 vdd.n673 vdd.n670 185
R16011 vdd.n2510 vdd.n2509 185
R16012 vdd.n2509 vdd.n2508 185
R16013 vdd.n675 vdd.n674 185
R16014 vdd.n683 vdd.n675 185
R16015 vdd.n2501 vdd.n2500 185
R16016 vdd.n2502 vdd.n2501 185
R16017 vdd.n2499 vdd.n684 185
R16018 vdd.n690 vdd.n684 185
R16019 vdd.n2498 vdd.n2497 185
R16020 vdd.n2497 vdd.n2496 185
R16021 vdd.n686 vdd.n685 185
R16022 vdd.n687 vdd.n686 185
R16023 vdd.n2489 vdd.n2488 185
R16024 vdd.n2490 vdd.n2489 185
R16025 vdd.n2487 vdd.n696 185
R16026 vdd.n2395 vdd.n696 185
R16027 vdd.n2486 vdd.n2485 185
R16028 vdd.n2485 vdd.n2484 185
R16029 vdd.n698 vdd.n697 185
R16030 vdd.t195 vdd.n698 185
R16031 vdd.n2477 vdd.n2476 185
R16032 vdd.n2478 vdd.n2477 185
R16033 vdd.n2475 vdd.n706 185
R16034 vdd.n2474 vdd.n2473 185
R16035 vdd.n708 vdd.n707 185
R16036 vdd.n2260 vdd.n2259 185
R16037 vdd.n2262 vdd.n2261 185
R16038 vdd.n2264 vdd.n2263 185
R16039 vdd.n2266 vdd.n2265 185
R16040 vdd.n2268 vdd.n2267 185
R16041 vdd.n2270 vdd.n2269 185
R16042 vdd.n2272 vdd.n2271 185
R16043 vdd.n2274 vdd.n2273 185
R16044 vdd.n2276 vdd.n2275 185
R16045 vdd.n2278 vdd.n2277 185
R16046 vdd.n2280 vdd.n2279 185
R16047 vdd.n2282 vdd.n2281 185
R16048 vdd.n2284 vdd.n2283 185
R16049 vdd.n2286 vdd.n2285 185
R16050 vdd.n2288 vdd.n2287 185
R16051 vdd.n2290 vdd.n2289 185
R16052 vdd.n2292 vdd.n2291 185
R16053 vdd.n2294 vdd.n2293 185
R16054 vdd.n2296 vdd.n2295 185
R16055 vdd.n2298 vdd.n2297 185
R16056 vdd.n2300 vdd.n2299 185
R16057 vdd.n2302 vdd.n2301 185
R16058 vdd.n2304 vdd.n2303 185
R16059 vdd.n2306 vdd.n2305 185
R16060 vdd.n2308 vdd.n2307 185
R16061 vdd.n2310 vdd.n2309 185
R16062 vdd.n2312 vdd.n2311 185
R16063 vdd.n2314 vdd.n2313 185
R16064 vdd.n2316 vdd.n2315 185
R16065 vdd.n2318 vdd.n2317 185
R16066 vdd.n2320 vdd.n2319 185
R16067 vdd.n2321 vdd.n2251 185
R16068 vdd.n2471 vdd.n2251 185
R16069 vdd.n2676 vdd.n2675 185
R16070 vdd.n2677 vdd.n588 185
R16071 vdd.n2679 vdd.n2678 185
R16072 vdd.n2681 vdd.n586 185
R16073 vdd.n2683 vdd.n2682 185
R16074 vdd.n2684 vdd.n585 185
R16075 vdd.n2686 vdd.n2685 185
R16076 vdd.n2688 vdd.n583 185
R16077 vdd.n2690 vdd.n2689 185
R16078 vdd.n2691 vdd.n582 185
R16079 vdd.n2693 vdd.n2692 185
R16080 vdd.n2695 vdd.n580 185
R16081 vdd.n2697 vdd.n2696 185
R16082 vdd.n2698 vdd.n579 185
R16083 vdd.n2700 vdd.n2699 185
R16084 vdd.n2702 vdd.n578 185
R16085 vdd.n2703 vdd.n576 185
R16086 vdd.n2706 vdd.n2705 185
R16087 vdd.n577 vdd.n575 185
R16088 vdd.n2562 vdd.n2561 185
R16089 vdd.n2564 vdd.n2563 185
R16090 vdd.n2566 vdd.n2558 185
R16091 vdd.n2568 vdd.n2567 185
R16092 vdd.n2569 vdd.n2557 185
R16093 vdd.n2571 vdd.n2570 185
R16094 vdd.n2573 vdd.n2555 185
R16095 vdd.n2575 vdd.n2574 185
R16096 vdd.n2576 vdd.n2554 185
R16097 vdd.n2578 vdd.n2577 185
R16098 vdd.n2580 vdd.n2552 185
R16099 vdd.n2582 vdd.n2581 185
R16100 vdd.n2583 vdd.n2551 185
R16101 vdd.n2585 vdd.n2584 185
R16102 vdd.n2587 vdd.n2550 185
R16103 vdd.n2589 vdd.n2588 185
R16104 vdd.n2588 vdd.n484 185
R16105 vdd.n2674 vdd.n592 185
R16106 vdd.n2674 vdd.n2673 185
R16107 vdd.n2326 vdd.n594 185
R16108 vdd.n595 vdd.n594 185
R16109 vdd.n2327 vdd.n628 185
R16110 vdd.n2603 vdd.n628 185
R16111 vdd.n2329 vdd.n2328 185
R16112 vdd.n2328 vdd.n636 185
R16113 vdd.n2330 vdd.n635 185
R16114 vdd.n2597 vdd.n635 185
R16115 vdd.n2332 vdd.n2331 185
R16116 vdd.n2331 vdd.n633 185
R16117 vdd.n2333 vdd.n643 185
R16118 vdd.n2546 vdd.n643 185
R16119 vdd.n2335 vdd.n2334 185
R16120 vdd.n2334 vdd.n641 185
R16121 vdd.n2336 vdd.n649 185
R16122 vdd.n2540 vdd.n649 185
R16123 vdd.n2338 vdd.n2337 185
R16124 vdd.n2337 vdd.n647 185
R16125 vdd.n2339 vdd.n654 185
R16126 vdd.n2532 vdd.n654 185
R16127 vdd.n2341 vdd.n2340 185
R16128 vdd.n2340 vdd.n660 185
R16129 vdd.n2342 vdd.n659 185
R16130 vdd.n2526 vdd.n659 185
R16131 vdd.n2376 vdd.n2375 185
R16132 vdd.n2375 vdd.n2374 185
R16133 vdd.n2377 vdd.n666 185
R16134 vdd.n2520 vdd.n666 185
R16135 vdd.n2379 vdd.n2378 185
R16136 vdd.n2378 vdd.n664 185
R16137 vdd.n2380 vdd.n672 185
R16138 vdd.n2514 vdd.n672 185
R16139 vdd.n2382 vdd.n2381 185
R16140 vdd.n2381 vdd.n670 185
R16141 vdd.n2383 vdd.n677 185
R16142 vdd.n2508 vdd.n677 185
R16143 vdd.n2385 vdd.n2384 185
R16144 vdd.n2384 vdd.n683 185
R16145 vdd.n2386 vdd.n682 185
R16146 vdd.n2502 vdd.n682 185
R16147 vdd.n2388 vdd.n2387 185
R16148 vdd.n2387 vdd.n690 185
R16149 vdd.n2389 vdd.n689 185
R16150 vdd.n2496 vdd.n689 185
R16151 vdd.n2391 vdd.n2390 185
R16152 vdd.n2390 vdd.n687 185
R16153 vdd.n2392 vdd.n695 185
R16154 vdd.n2490 vdd.n695 185
R16155 vdd.n2394 vdd.n2393 185
R16156 vdd.n2395 vdd.n2394 185
R16157 vdd.n2325 vdd.n700 185
R16158 vdd.n2484 vdd.n700 185
R16159 vdd.n2324 vdd.n2323 185
R16160 vdd.n2323 vdd.t195 185
R16161 vdd.n2322 vdd.n705 185
R16162 vdd.n2478 vdd.n705 185
R16163 vdd.n1942 vdd.n1941 185
R16164 vdd.n1943 vdd.n1942 185
R16165 vdd.n866 vdd.n864 185
R16166 vdd.n1508 vdd.n864 185
R16167 vdd.n1511 vdd.n1510 185
R16168 vdd.n1510 vdd.n1509 185
R16169 vdd.n869 vdd.n868 185
R16170 vdd.n870 vdd.n869 185
R16171 vdd.n1497 vdd.n1496 185
R16172 vdd.n1498 vdd.n1497 185
R16173 vdd.n878 vdd.n877 185
R16174 vdd.n1489 vdd.n877 185
R16175 vdd.n1492 vdd.n1491 185
R16176 vdd.n1491 vdd.n1490 185
R16177 vdd.n881 vdd.n880 185
R16178 vdd.n888 vdd.n881 185
R16179 vdd.n1480 vdd.n1479 185
R16180 vdd.n1481 vdd.n1480 185
R16181 vdd.n890 vdd.n889 185
R16182 vdd.n889 vdd.n887 185
R16183 vdd.n1475 vdd.n1474 185
R16184 vdd.n1474 vdd.n1473 185
R16185 vdd.n1163 vdd.n1162 185
R16186 vdd.n1164 vdd.n1163 185
R16187 vdd.n1464 vdd.n1463 185
R16188 vdd.n1465 vdd.n1464 185
R16189 vdd.n1171 vdd.n1170 185
R16190 vdd.n1455 vdd.n1170 185
R16191 vdd.n1458 vdd.n1457 185
R16192 vdd.n1457 vdd.n1456 185
R16193 vdd.n1174 vdd.n1173 185
R16194 vdd.n1180 vdd.n1174 185
R16195 vdd.n1446 vdd.n1445 185
R16196 vdd.n1447 vdd.n1446 185
R16197 vdd.n1182 vdd.n1181 185
R16198 vdd.n1438 vdd.n1181 185
R16199 vdd.n1441 vdd.n1440 185
R16200 vdd.n1440 vdd.n1439 185
R16201 vdd.n1185 vdd.n1184 185
R16202 vdd.n1186 vdd.n1185 185
R16203 vdd.n1429 vdd.n1428 185
R16204 vdd.n1430 vdd.n1429 185
R16205 vdd.n1193 vdd.n1192 185
R16206 vdd.n1228 vdd.n1192 185
R16207 vdd.n1424 vdd.n1423 185
R16208 vdd.n1196 vdd.n1195 185
R16209 vdd.n1420 vdd.n1419 185
R16210 vdd.n1421 vdd.n1420 185
R16211 vdd.n1230 vdd.n1229 185
R16212 vdd.n1415 vdd.n1232 185
R16213 vdd.n1414 vdd.n1233 185
R16214 vdd.n1413 vdd.n1234 185
R16215 vdd.n1236 vdd.n1235 185
R16216 vdd.n1409 vdd.n1238 185
R16217 vdd.n1408 vdd.n1239 185
R16218 vdd.n1407 vdd.n1240 185
R16219 vdd.n1242 vdd.n1241 185
R16220 vdd.n1403 vdd.n1244 185
R16221 vdd.n1402 vdd.n1245 185
R16222 vdd.n1401 vdd.n1246 185
R16223 vdd.n1248 vdd.n1247 185
R16224 vdd.n1397 vdd.n1250 185
R16225 vdd.n1396 vdd.n1251 185
R16226 vdd.n1395 vdd.n1252 185
R16227 vdd.n1256 vdd.n1253 185
R16228 vdd.n1391 vdd.n1258 185
R16229 vdd.n1390 vdd.n1259 185
R16230 vdd.n1389 vdd.n1260 185
R16231 vdd.n1262 vdd.n1261 185
R16232 vdd.n1385 vdd.n1264 185
R16233 vdd.n1384 vdd.n1265 185
R16234 vdd.n1383 vdd.n1266 185
R16235 vdd.n1268 vdd.n1267 185
R16236 vdd.n1379 vdd.n1270 185
R16237 vdd.n1378 vdd.n1271 185
R16238 vdd.n1377 vdd.n1272 185
R16239 vdd.n1274 vdd.n1273 185
R16240 vdd.n1373 vdd.n1276 185
R16241 vdd.n1372 vdd.n1277 185
R16242 vdd.n1371 vdd.n1278 185
R16243 vdd.n1280 vdd.n1279 185
R16244 vdd.n1367 vdd.n1282 185
R16245 vdd.n1366 vdd.n1283 185
R16246 vdd.n1365 vdd.n1284 185
R16247 vdd.n1286 vdd.n1285 185
R16248 vdd.n1361 vdd.n1288 185
R16249 vdd.n1360 vdd.n1357 185
R16250 vdd.n1356 vdd.n1289 185
R16251 vdd.n1291 vdd.n1290 185
R16252 vdd.n1352 vdd.n1293 185
R16253 vdd.n1351 vdd.n1294 185
R16254 vdd.n1350 vdd.n1295 185
R16255 vdd.n1297 vdd.n1296 185
R16256 vdd.n1346 vdd.n1299 185
R16257 vdd.n1345 vdd.n1300 185
R16258 vdd.n1344 vdd.n1301 185
R16259 vdd.n1303 vdd.n1302 185
R16260 vdd.n1340 vdd.n1305 185
R16261 vdd.n1339 vdd.n1306 185
R16262 vdd.n1338 vdd.n1307 185
R16263 vdd.n1309 vdd.n1308 185
R16264 vdd.n1334 vdd.n1311 185
R16265 vdd.n1333 vdd.n1312 185
R16266 vdd.n1332 vdd.n1313 185
R16267 vdd.n1315 vdd.n1314 185
R16268 vdd.n1328 vdd.n1317 185
R16269 vdd.n1327 vdd.n1318 185
R16270 vdd.n1326 vdd.n1319 185
R16271 vdd.n1323 vdd.n1227 185
R16272 vdd.n1421 vdd.n1227 185
R16273 vdd.n1946 vdd.n1945 185
R16274 vdd.n1950 vdd.n859 185
R16275 vdd.n1613 vdd.n858 185
R16276 vdd.n1616 vdd.n1615 185
R16277 vdd.n1618 vdd.n1617 185
R16278 vdd.n1621 vdd.n1620 185
R16279 vdd.n1623 vdd.n1622 185
R16280 vdd.n1625 vdd.n1611 185
R16281 vdd.n1627 vdd.n1626 185
R16282 vdd.n1628 vdd.n1605 185
R16283 vdd.n1630 vdd.n1629 185
R16284 vdd.n1632 vdd.n1603 185
R16285 vdd.n1634 vdd.n1633 185
R16286 vdd.n1635 vdd.n1598 185
R16287 vdd.n1637 vdd.n1636 185
R16288 vdd.n1639 vdd.n1596 185
R16289 vdd.n1641 vdd.n1640 185
R16290 vdd.n1642 vdd.n1592 185
R16291 vdd.n1644 vdd.n1643 185
R16292 vdd.n1646 vdd.n1589 185
R16293 vdd.n1648 vdd.n1647 185
R16294 vdd.n1590 vdd.n1583 185
R16295 vdd.n1652 vdd.n1587 185
R16296 vdd.n1653 vdd.n1579 185
R16297 vdd.n1655 vdd.n1654 185
R16298 vdd.n1657 vdd.n1577 185
R16299 vdd.n1659 vdd.n1658 185
R16300 vdd.n1660 vdd.n1572 185
R16301 vdd.n1662 vdd.n1661 185
R16302 vdd.n1664 vdd.n1570 185
R16303 vdd.n1666 vdd.n1665 185
R16304 vdd.n1667 vdd.n1565 185
R16305 vdd.n1669 vdd.n1668 185
R16306 vdd.n1671 vdd.n1563 185
R16307 vdd.n1673 vdd.n1672 185
R16308 vdd.n1674 vdd.n1558 185
R16309 vdd.n1676 vdd.n1675 185
R16310 vdd.n1678 vdd.n1556 185
R16311 vdd.n1680 vdd.n1679 185
R16312 vdd.n1681 vdd.n1552 185
R16313 vdd.n1683 vdd.n1682 185
R16314 vdd.n1685 vdd.n1549 185
R16315 vdd.n1687 vdd.n1686 185
R16316 vdd.n1550 vdd.n1543 185
R16317 vdd.n1691 vdd.n1547 185
R16318 vdd.n1692 vdd.n1539 185
R16319 vdd.n1694 vdd.n1693 185
R16320 vdd.n1696 vdd.n1537 185
R16321 vdd.n1698 vdd.n1697 185
R16322 vdd.n1699 vdd.n1532 185
R16323 vdd.n1701 vdd.n1700 185
R16324 vdd.n1703 vdd.n1530 185
R16325 vdd.n1705 vdd.n1704 185
R16326 vdd.n1706 vdd.n1525 185
R16327 vdd.n1708 vdd.n1707 185
R16328 vdd.n1710 vdd.n1524 185
R16329 vdd.n1711 vdd.n1521 185
R16330 vdd.n1714 vdd.n1713 185
R16331 vdd.n1523 vdd.n1519 185
R16332 vdd.n1931 vdd.n1517 185
R16333 vdd.n1933 vdd.n1932 185
R16334 vdd.n1935 vdd.n1515 185
R16335 vdd.n1937 vdd.n1936 185
R16336 vdd.n1938 vdd.n865 185
R16337 vdd.n1944 vdd.n862 185
R16338 vdd.n1944 vdd.n1943 185
R16339 vdd.n873 vdd.n861 185
R16340 vdd.n1508 vdd.n861 185
R16341 vdd.n1507 vdd.n1506 185
R16342 vdd.n1509 vdd.n1507 185
R16343 vdd.n872 vdd.n871 185
R16344 vdd.n871 vdd.n870 185
R16345 vdd.n1500 vdd.n1499 185
R16346 vdd.n1499 vdd.n1498 185
R16347 vdd.n876 vdd.n875 185
R16348 vdd.n1489 vdd.n876 185
R16349 vdd.n1488 vdd.n1487 185
R16350 vdd.n1490 vdd.n1488 185
R16351 vdd.n883 vdd.n882 185
R16352 vdd.n888 vdd.n882 185
R16353 vdd.n1483 vdd.n1482 185
R16354 vdd.n1482 vdd.n1481 185
R16355 vdd.n886 vdd.n885 185
R16356 vdd.n887 vdd.n886 185
R16357 vdd.n1472 vdd.n1471 185
R16358 vdd.n1473 vdd.n1472 185
R16359 vdd.n1166 vdd.n1165 185
R16360 vdd.n1165 vdd.n1164 185
R16361 vdd.n1467 vdd.n1466 185
R16362 vdd.n1466 vdd.n1465 185
R16363 vdd.n1169 vdd.n1168 185
R16364 vdd.n1455 vdd.n1169 185
R16365 vdd.n1454 vdd.n1453 185
R16366 vdd.n1456 vdd.n1454 185
R16367 vdd.n1176 vdd.n1175 185
R16368 vdd.n1180 vdd.n1175 185
R16369 vdd.n1449 vdd.n1448 185
R16370 vdd.n1448 vdd.n1447 185
R16371 vdd.n1179 vdd.n1178 185
R16372 vdd.n1438 vdd.n1179 185
R16373 vdd.n1437 vdd.n1436 185
R16374 vdd.n1439 vdd.n1437 185
R16375 vdd.n1188 vdd.n1187 185
R16376 vdd.n1187 vdd.n1186 185
R16377 vdd.n1432 vdd.n1431 185
R16378 vdd.n1431 vdd.n1430 185
R16379 vdd.n1191 vdd.n1190 185
R16380 vdd.n1228 vdd.n1191 185
R16381 vdd.n746 vdd.n744 185
R16382 vdd.n2146 vdd.n744 185
R16383 vdd.n2068 vdd.n763 185
R16384 vdd.n763 vdd.t189 185
R16385 vdd.n2070 vdd.n2069 185
R16386 vdd.n2071 vdd.n2070 185
R16387 vdd.n2067 vdd.n762 185
R16388 vdd.n1770 vdd.n762 185
R16389 vdd.n2066 vdd.n2065 185
R16390 vdd.n2065 vdd.n2064 185
R16391 vdd.n765 vdd.n764 185
R16392 vdd.n766 vdd.n765 185
R16393 vdd.n2055 vdd.n2054 185
R16394 vdd.n2056 vdd.n2055 185
R16395 vdd.n2053 vdd.n776 185
R16396 vdd.n776 vdd.n773 185
R16397 vdd.n2052 vdd.n2051 185
R16398 vdd.n2051 vdd.n2050 185
R16399 vdd.n778 vdd.n777 185
R16400 vdd.n779 vdd.n778 185
R16401 vdd.n2043 vdd.n2042 185
R16402 vdd.n2044 vdd.n2043 185
R16403 vdd.n2041 vdd.n787 185
R16404 vdd.n792 vdd.n787 185
R16405 vdd.n2040 vdd.n2039 185
R16406 vdd.n2039 vdd.n2038 185
R16407 vdd.n789 vdd.n788 185
R16408 vdd.n798 vdd.n789 185
R16409 vdd.n2031 vdd.n2030 185
R16410 vdd.n2032 vdd.n2031 185
R16411 vdd.n2029 vdd.n799 185
R16412 vdd.n1871 vdd.n799 185
R16413 vdd.n2028 vdd.n2027 185
R16414 vdd.n2027 vdd.n2026 185
R16415 vdd.n801 vdd.n800 185
R16416 vdd.n802 vdd.n801 185
R16417 vdd.n2019 vdd.n2018 185
R16418 vdd.n2020 vdd.n2019 185
R16419 vdd.n2017 vdd.n811 185
R16420 vdd.n811 vdd.n808 185
R16421 vdd.n2016 vdd.n2015 185
R16422 vdd.n2015 vdd.n2014 185
R16423 vdd.n813 vdd.n812 185
R16424 vdd.n823 vdd.n813 185
R16425 vdd.n2006 vdd.n2005 185
R16426 vdd.n2007 vdd.n2006 185
R16427 vdd.n2004 vdd.n824 185
R16428 vdd.n824 vdd.n820 185
R16429 vdd.n2003 vdd.n2002 185
R16430 vdd.n2002 vdd.n2001 185
R16431 vdd.n826 vdd.n825 185
R16432 vdd.n827 vdd.n826 185
R16433 vdd.n1994 vdd.n1993 185
R16434 vdd.n1995 vdd.n1994 185
R16435 vdd.n1992 vdd.n836 185
R16436 vdd.n836 vdd.n833 185
R16437 vdd.n1991 vdd.n1990 185
R16438 vdd.n1990 vdd.n1989 185
R16439 vdd.n838 vdd.n837 185
R16440 vdd.n1726 vdd.n1725 185
R16441 vdd.n1727 vdd.n1723 185
R16442 vdd.n1723 vdd.n839 185
R16443 vdd.n1729 vdd.n1728 185
R16444 vdd.n1731 vdd.n1722 185
R16445 vdd.n1734 vdd.n1733 185
R16446 vdd.n1735 vdd.n1721 185
R16447 vdd.n1737 vdd.n1736 185
R16448 vdd.n1739 vdd.n1720 185
R16449 vdd.n1742 vdd.n1741 185
R16450 vdd.n1743 vdd.n1719 185
R16451 vdd.n1745 vdd.n1744 185
R16452 vdd.n1747 vdd.n1718 185
R16453 vdd.n1750 vdd.n1749 185
R16454 vdd.n1751 vdd.n1717 185
R16455 vdd.n1753 vdd.n1752 185
R16456 vdd.n1755 vdd.n1716 185
R16457 vdd.n1928 vdd.n1756 185
R16458 vdd.n1927 vdd.n1926 185
R16459 vdd.n1924 vdd.n1757 185
R16460 vdd.n1922 vdd.n1921 185
R16461 vdd.n1920 vdd.n1758 185
R16462 vdd.n1919 vdd.n1918 185
R16463 vdd.n1916 vdd.n1759 185
R16464 vdd.n1914 vdd.n1913 185
R16465 vdd.n1912 vdd.n1760 185
R16466 vdd.n1911 vdd.n1910 185
R16467 vdd.n1908 vdd.n1761 185
R16468 vdd.n1906 vdd.n1905 185
R16469 vdd.n1904 vdd.n1762 185
R16470 vdd.n1903 vdd.n1902 185
R16471 vdd.n1900 vdd.n1763 185
R16472 vdd.n1898 vdd.n1897 185
R16473 vdd.n1896 vdd.n1764 185
R16474 vdd.n1895 vdd.n1894 185
R16475 vdd.n2149 vdd.n2148 185
R16476 vdd.n2151 vdd.n2150 185
R16477 vdd.n2153 vdd.n2152 185
R16478 vdd.n2156 vdd.n2155 185
R16479 vdd.n2158 vdd.n2157 185
R16480 vdd.n2160 vdd.n2159 185
R16481 vdd.n2162 vdd.n2161 185
R16482 vdd.n2164 vdd.n2163 185
R16483 vdd.n2166 vdd.n2165 185
R16484 vdd.n2168 vdd.n2167 185
R16485 vdd.n2170 vdd.n2169 185
R16486 vdd.n2172 vdd.n2171 185
R16487 vdd.n2174 vdd.n2173 185
R16488 vdd.n2176 vdd.n2175 185
R16489 vdd.n2178 vdd.n2177 185
R16490 vdd.n2180 vdd.n2179 185
R16491 vdd.n2182 vdd.n2181 185
R16492 vdd.n2184 vdd.n2183 185
R16493 vdd.n2186 vdd.n2185 185
R16494 vdd.n2188 vdd.n2187 185
R16495 vdd.n2190 vdd.n2189 185
R16496 vdd.n2192 vdd.n2191 185
R16497 vdd.n2194 vdd.n2193 185
R16498 vdd.n2196 vdd.n2195 185
R16499 vdd.n2198 vdd.n2197 185
R16500 vdd.n2200 vdd.n2199 185
R16501 vdd.n2202 vdd.n2201 185
R16502 vdd.n2204 vdd.n2203 185
R16503 vdd.n2206 vdd.n2205 185
R16504 vdd.n2208 vdd.n2207 185
R16505 vdd.n2210 vdd.n2209 185
R16506 vdd.n2212 vdd.n2211 185
R16507 vdd.n2214 vdd.n2213 185
R16508 vdd.n2215 vdd.n745 185
R16509 vdd.n2217 vdd.n2216 185
R16510 vdd.n2218 vdd.n2217 185
R16511 vdd.n2147 vdd.n749 185
R16512 vdd.n2147 vdd.n2146 185
R16513 vdd.n1768 vdd.n750 185
R16514 vdd.t189 vdd.n750 185
R16515 vdd.n1769 vdd.n760 185
R16516 vdd.n2071 vdd.n760 185
R16517 vdd.n1772 vdd.n1771 185
R16518 vdd.n1771 vdd.n1770 185
R16519 vdd.n1773 vdd.n767 185
R16520 vdd.n2064 vdd.n767 185
R16521 vdd.n1775 vdd.n1774 185
R16522 vdd.n1774 vdd.n766 185
R16523 vdd.n1776 vdd.n774 185
R16524 vdd.n2056 vdd.n774 185
R16525 vdd.n1778 vdd.n1777 185
R16526 vdd.n1777 vdd.n773 185
R16527 vdd.n1779 vdd.n780 185
R16528 vdd.n2050 vdd.n780 185
R16529 vdd.n1781 vdd.n1780 185
R16530 vdd.n1780 vdd.n779 185
R16531 vdd.n1782 vdd.n785 185
R16532 vdd.n2044 vdd.n785 185
R16533 vdd.n1784 vdd.n1783 185
R16534 vdd.n1783 vdd.n792 185
R16535 vdd.n1785 vdd.n790 185
R16536 vdd.n2038 vdd.n790 185
R16537 vdd.n1787 vdd.n1786 185
R16538 vdd.n1786 vdd.n798 185
R16539 vdd.n1788 vdd.n796 185
R16540 vdd.n2032 vdd.n796 185
R16541 vdd.n1873 vdd.n1872 185
R16542 vdd.n1872 vdd.n1871 185
R16543 vdd.n1874 vdd.n803 185
R16544 vdd.n2026 vdd.n803 185
R16545 vdd.n1876 vdd.n1875 185
R16546 vdd.n1875 vdd.n802 185
R16547 vdd.n1877 vdd.n809 185
R16548 vdd.n2020 vdd.n809 185
R16549 vdd.n1879 vdd.n1878 185
R16550 vdd.n1878 vdd.n808 185
R16551 vdd.n1880 vdd.n814 185
R16552 vdd.n2014 vdd.n814 185
R16553 vdd.n1882 vdd.n1881 185
R16554 vdd.n1881 vdd.n823 185
R16555 vdd.n1883 vdd.n821 185
R16556 vdd.n2007 vdd.n821 185
R16557 vdd.n1885 vdd.n1884 185
R16558 vdd.n1884 vdd.n820 185
R16559 vdd.n1886 vdd.n828 185
R16560 vdd.n2001 vdd.n828 185
R16561 vdd.n1888 vdd.n1887 185
R16562 vdd.n1887 vdd.n827 185
R16563 vdd.n1889 vdd.n834 185
R16564 vdd.n1995 vdd.n834 185
R16565 vdd.n1891 vdd.n1890 185
R16566 vdd.n1890 vdd.n833 185
R16567 vdd.n1892 vdd.n840 185
R16568 vdd.n1989 vdd.n840 185
R16569 vdd.n3024 vdd.n3023 185
R16570 vdd.n3025 vdd.n3024 185
R16571 vdd.n325 vdd.n324 185
R16572 vdd.n3026 vdd.n325 185
R16573 vdd.n3029 vdd.n3028 185
R16574 vdd.n3028 vdd.n3027 185
R16575 vdd.n3030 vdd.n319 185
R16576 vdd.n319 vdd.n318 185
R16577 vdd.n3032 vdd.n3031 185
R16578 vdd.n3033 vdd.n3032 185
R16579 vdd.n314 vdd.n313 185
R16580 vdd.n3034 vdd.n314 185
R16581 vdd.n3037 vdd.n3036 185
R16582 vdd.n3036 vdd.n3035 185
R16583 vdd.n3038 vdd.n309 185
R16584 vdd.n309 vdd.n308 185
R16585 vdd.n3040 vdd.n3039 185
R16586 vdd.n3041 vdd.n3040 185
R16587 vdd.n303 vdd.n301 185
R16588 vdd.n3042 vdd.n303 185
R16589 vdd.n3045 vdd.n3044 185
R16590 vdd.n3044 vdd.n3043 185
R16591 vdd.n302 vdd.n300 185
R16592 vdd.n304 vdd.n302 185
R16593 vdd.n2881 vdd.n2880 185
R16594 vdd.n2882 vdd.n2881 185
R16595 vdd.n458 vdd.n457 185
R16596 vdd.n457 vdd.n456 185
R16597 vdd.n2876 vdd.n2875 185
R16598 vdd.n2875 vdd.n2874 185
R16599 vdd.n461 vdd.n460 185
R16600 vdd.n467 vdd.n461 185
R16601 vdd.n2865 vdd.n2864 185
R16602 vdd.n2866 vdd.n2865 185
R16603 vdd.n469 vdd.n468 185
R16604 vdd.n2857 vdd.n468 185
R16605 vdd.n2860 vdd.n2859 185
R16606 vdd.n2859 vdd.n2858 185
R16607 vdd.n472 vdd.n471 185
R16608 vdd.n473 vdd.n472 185
R16609 vdd.n2848 vdd.n2847 185
R16610 vdd.n2849 vdd.n2848 185
R16611 vdd.n480 vdd.n479 185
R16612 vdd.n516 vdd.n479 185
R16613 vdd.n2843 vdd.n2842 185
R16614 vdd.n483 vdd.n482 185
R16615 vdd.n2839 vdd.n2838 185
R16616 vdd.n2840 vdd.n2839 185
R16617 vdd.n518 vdd.n517 185
R16618 vdd.n522 vdd.n521 185
R16619 vdd.n2834 vdd.n523 185
R16620 vdd.n2833 vdd.n2832 185
R16621 vdd.n2831 vdd.n2830 185
R16622 vdd.n2829 vdd.n2828 185
R16623 vdd.n2827 vdd.n2826 185
R16624 vdd.n2825 vdd.n2824 185
R16625 vdd.n2823 vdd.n2822 185
R16626 vdd.n2821 vdd.n2820 185
R16627 vdd.n2819 vdd.n2818 185
R16628 vdd.n2817 vdd.n2816 185
R16629 vdd.n2815 vdd.n2814 185
R16630 vdd.n2813 vdd.n2812 185
R16631 vdd.n2811 vdd.n2810 185
R16632 vdd.n2809 vdd.n2808 185
R16633 vdd.n2807 vdd.n2806 185
R16634 vdd.n2798 vdd.n536 185
R16635 vdd.n2800 vdd.n2799 185
R16636 vdd.n2797 vdd.n2796 185
R16637 vdd.n2795 vdd.n2794 185
R16638 vdd.n2793 vdd.n2792 185
R16639 vdd.n2791 vdd.n2790 185
R16640 vdd.n2789 vdd.n2788 185
R16641 vdd.n2787 vdd.n2786 185
R16642 vdd.n2785 vdd.n2784 185
R16643 vdd.n2783 vdd.n2782 185
R16644 vdd.n2781 vdd.n2780 185
R16645 vdd.n2779 vdd.n2778 185
R16646 vdd.n2777 vdd.n2776 185
R16647 vdd.n2775 vdd.n2774 185
R16648 vdd.n2773 vdd.n2772 185
R16649 vdd.n2771 vdd.n2770 185
R16650 vdd.n2769 vdd.n2768 185
R16651 vdd.n2767 vdd.n2766 185
R16652 vdd.n2765 vdd.n2764 185
R16653 vdd.n2763 vdd.n2762 185
R16654 vdd.n2761 vdd.n2760 185
R16655 vdd.n2759 vdd.n2758 185
R16656 vdd.n2752 vdd.n556 185
R16657 vdd.n2754 vdd.n2753 185
R16658 vdd.n2751 vdd.n2750 185
R16659 vdd.n2749 vdd.n2748 185
R16660 vdd.n2747 vdd.n2746 185
R16661 vdd.n2745 vdd.n2744 185
R16662 vdd.n2743 vdd.n2742 185
R16663 vdd.n2741 vdd.n2740 185
R16664 vdd.n2739 vdd.n2738 185
R16665 vdd.n2737 vdd.n2736 185
R16666 vdd.n2735 vdd.n2734 185
R16667 vdd.n2733 vdd.n2732 185
R16668 vdd.n2731 vdd.n2730 185
R16669 vdd.n2729 vdd.n2728 185
R16670 vdd.n2727 vdd.n2726 185
R16671 vdd.n2725 vdd.n2724 185
R16672 vdd.n2723 vdd.n2722 185
R16673 vdd.n2721 vdd.n2720 185
R16674 vdd.n2719 vdd.n2718 185
R16675 vdd.n2717 vdd.n2716 185
R16676 vdd.n2715 vdd.n2714 185
R16677 vdd.n2710 vdd.n515 185
R16678 vdd.n2840 vdd.n515 185
R16679 vdd.n2907 vdd.n2906 185
R16680 vdd.n2911 vdd.n440 185
R16681 vdd.n2913 vdd.n2912 185
R16682 vdd.n2915 vdd.n438 185
R16683 vdd.n2917 vdd.n2916 185
R16684 vdd.n2918 vdd.n433 185
R16685 vdd.n2920 vdd.n2919 185
R16686 vdd.n2922 vdd.n431 185
R16687 vdd.n2924 vdd.n2923 185
R16688 vdd.n2925 vdd.n426 185
R16689 vdd.n2927 vdd.n2926 185
R16690 vdd.n2929 vdd.n424 185
R16691 vdd.n2931 vdd.n2930 185
R16692 vdd.n2932 vdd.n419 185
R16693 vdd.n2934 vdd.n2933 185
R16694 vdd.n2936 vdd.n417 185
R16695 vdd.n2938 vdd.n2937 185
R16696 vdd.n2939 vdd.n413 185
R16697 vdd.n2941 vdd.n2940 185
R16698 vdd.n2943 vdd.n410 185
R16699 vdd.n2945 vdd.n2944 185
R16700 vdd.n411 vdd.n404 185
R16701 vdd.n2949 vdd.n408 185
R16702 vdd.n2950 vdd.n400 185
R16703 vdd.n2952 vdd.n2951 185
R16704 vdd.n2954 vdd.n398 185
R16705 vdd.n2956 vdd.n2955 185
R16706 vdd.n2957 vdd.n393 185
R16707 vdd.n2959 vdd.n2958 185
R16708 vdd.n2961 vdd.n391 185
R16709 vdd.n2963 vdd.n2962 185
R16710 vdd.n2964 vdd.n386 185
R16711 vdd.n2966 vdd.n2965 185
R16712 vdd.n2968 vdd.n384 185
R16713 vdd.n2970 vdd.n2969 185
R16714 vdd.n2971 vdd.n379 185
R16715 vdd.n2973 vdd.n2972 185
R16716 vdd.n2975 vdd.n377 185
R16717 vdd.n2977 vdd.n2976 185
R16718 vdd.n2978 vdd.n373 185
R16719 vdd.n2980 vdd.n2979 185
R16720 vdd.n2982 vdd.n370 185
R16721 vdd.n2984 vdd.n2983 185
R16722 vdd.n371 vdd.n364 185
R16723 vdd.n2988 vdd.n368 185
R16724 vdd.n2989 vdd.n360 185
R16725 vdd.n2991 vdd.n2990 185
R16726 vdd.n2993 vdd.n358 185
R16727 vdd.n2995 vdd.n2994 185
R16728 vdd.n2996 vdd.n353 185
R16729 vdd.n2998 vdd.n2997 185
R16730 vdd.n3000 vdd.n351 185
R16731 vdd.n3002 vdd.n3001 185
R16732 vdd.n3003 vdd.n346 185
R16733 vdd.n3005 vdd.n3004 185
R16734 vdd.n3007 vdd.n344 185
R16735 vdd.n3009 vdd.n3008 185
R16736 vdd.n3010 vdd.n338 185
R16737 vdd.n3012 vdd.n3011 185
R16738 vdd.n3014 vdd.n337 185
R16739 vdd.n3015 vdd.n336 185
R16740 vdd.n3018 vdd.n3017 185
R16741 vdd.n3019 vdd.n334 185
R16742 vdd.n3020 vdd.n330 185
R16743 vdd.n2902 vdd.n328 185
R16744 vdd.n3025 vdd.n328 185
R16745 vdd.n2901 vdd.n327 185
R16746 vdd.n3026 vdd.n327 185
R16747 vdd.n2900 vdd.n326 185
R16748 vdd.n3027 vdd.n326 185
R16749 vdd.n446 vdd.n445 185
R16750 vdd.n445 vdd.n318 185
R16751 vdd.n2896 vdd.n317 185
R16752 vdd.n3033 vdd.n317 185
R16753 vdd.n2895 vdd.n316 185
R16754 vdd.n3034 vdd.n316 185
R16755 vdd.n2894 vdd.n315 185
R16756 vdd.n3035 vdd.n315 185
R16757 vdd.n449 vdd.n448 185
R16758 vdd.n448 vdd.n308 185
R16759 vdd.n2890 vdd.n307 185
R16760 vdd.n3041 vdd.n307 185
R16761 vdd.n2889 vdd.n306 185
R16762 vdd.n3042 vdd.n306 185
R16763 vdd.n2888 vdd.n305 185
R16764 vdd.n3043 vdd.n305 185
R16765 vdd.n455 vdd.n451 185
R16766 vdd.n455 vdd.n304 185
R16767 vdd.n2884 vdd.n2883 185
R16768 vdd.n2883 vdd.n2882 185
R16769 vdd.n454 vdd.n453 185
R16770 vdd.n456 vdd.n454 185
R16771 vdd.n2873 vdd.n2872 185
R16772 vdd.n2874 vdd.n2873 185
R16773 vdd.n463 vdd.n462 185
R16774 vdd.n467 vdd.n462 185
R16775 vdd.n2868 vdd.n2867 185
R16776 vdd.n2867 vdd.n2866 185
R16777 vdd.n466 vdd.n465 185
R16778 vdd.n2857 vdd.n466 185
R16779 vdd.n2856 vdd.n2855 185
R16780 vdd.n2858 vdd.n2856 185
R16781 vdd.n475 vdd.n474 185
R16782 vdd.n474 vdd.n473 185
R16783 vdd.n2851 vdd.n2850 185
R16784 vdd.n2850 vdd.n2849 185
R16785 vdd.n478 vdd.n477 185
R16786 vdd.n516 vdd.n478 185
R16787 vdd.n703 vdd.n702 185
R16788 vdd.n2469 vdd.n2468 185
R16789 vdd.n2467 vdd.n2252 185
R16790 vdd.n2471 vdd.n2252 185
R16791 vdd.n2466 vdd.n2465 185
R16792 vdd.n2464 vdd.n2463 185
R16793 vdd.n2462 vdd.n2461 185
R16794 vdd.n2460 vdd.n2459 185
R16795 vdd.n2458 vdd.n2457 185
R16796 vdd.n2456 vdd.n2455 185
R16797 vdd.n2454 vdd.n2453 185
R16798 vdd.n2452 vdd.n2451 185
R16799 vdd.n2450 vdd.n2449 185
R16800 vdd.n2448 vdd.n2447 185
R16801 vdd.n2446 vdd.n2445 185
R16802 vdd.n2444 vdd.n2443 185
R16803 vdd.n2442 vdd.n2441 185
R16804 vdd.n2440 vdd.n2439 185
R16805 vdd.n2438 vdd.n2437 185
R16806 vdd.n2436 vdd.n2435 185
R16807 vdd.n2434 vdd.n2433 185
R16808 vdd.n2432 vdd.n2431 185
R16809 vdd.n2430 vdd.n2429 185
R16810 vdd.n2428 vdd.n2427 185
R16811 vdd.n2426 vdd.n2425 185
R16812 vdd.n2424 vdd.n2423 185
R16813 vdd.n2422 vdd.n2421 185
R16814 vdd.n2420 vdd.n2419 185
R16815 vdd.n2418 vdd.n2417 185
R16816 vdd.n2416 vdd.n2415 185
R16817 vdd.n2414 vdd.n2413 185
R16818 vdd.n2412 vdd.n2411 185
R16819 vdd.n2410 vdd.n2409 185
R16820 vdd.n2407 vdd.n2406 185
R16821 vdd.n2405 vdd.n2404 185
R16822 vdd.n2403 vdd.n2402 185
R16823 vdd.n2609 vdd.n2608 185
R16824 vdd.n2611 vdd.n624 185
R16825 vdd.n2613 vdd.n2612 185
R16826 vdd.n2615 vdd.n621 185
R16827 vdd.n2617 vdd.n2616 185
R16828 vdd.n2619 vdd.n619 185
R16829 vdd.n2621 vdd.n2620 185
R16830 vdd.n2622 vdd.n618 185
R16831 vdd.n2624 vdd.n2623 185
R16832 vdd.n2626 vdd.n616 185
R16833 vdd.n2628 vdd.n2627 185
R16834 vdd.n2629 vdd.n615 185
R16835 vdd.n2631 vdd.n2630 185
R16836 vdd.n2633 vdd.n613 185
R16837 vdd.n2635 vdd.n2634 185
R16838 vdd.n2636 vdd.n612 185
R16839 vdd.n2638 vdd.n2637 185
R16840 vdd.n2640 vdd.n520 185
R16841 vdd.n2642 vdd.n2641 185
R16842 vdd.n2644 vdd.n610 185
R16843 vdd.n2646 vdd.n2645 185
R16844 vdd.n2647 vdd.n609 185
R16845 vdd.n2649 vdd.n2648 185
R16846 vdd.n2651 vdd.n607 185
R16847 vdd.n2653 vdd.n2652 185
R16848 vdd.n2654 vdd.n606 185
R16849 vdd.n2656 vdd.n2655 185
R16850 vdd.n2658 vdd.n604 185
R16851 vdd.n2660 vdd.n2659 185
R16852 vdd.n2661 vdd.n603 185
R16853 vdd.n2663 vdd.n2662 185
R16854 vdd.n2665 vdd.n602 185
R16855 vdd.n2666 vdd.n601 185
R16856 vdd.n2669 vdd.n2668 185
R16857 vdd.n2670 vdd.n599 185
R16858 vdd.n599 vdd.n484 185
R16859 vdd.n2607 vdd.n596 185
R16860 vdd.n2673 vdd.n596 185
R16861 vdd.n2606 vdd.n2605 185
R16862 vdd.n2605 vdd.n595 185
R16863 vdd.n2604 vdd.n626 185
R16864 vdd.n2604 vdd.n2603 185
R16865 vdd.n2358 vdd.n627 185
R16866 vdd.n636 vdd.n627 185
R16867 vdd.n2359 vdd.n634 185
R16868 vdd.n2597 vdd.n634 185
R16869 vdd.n2361 vdd.n2360 185
R16870 vdd.n2360 vdd.n633 185
R16871 vdd.n2362 vdd.n642 185
R16872 vdd.n2546 vdd.n642 185
R16873 vdd.n2364 vdd.n2363 185
R16874 vdd.n2363 vdd.n641 185
R16875 vdd.n2365 vdd.n648 185
R16876 vdd.n2540 vdd.n648 185
R16877 vdd.n2367 vdd.n2366 185
R16878 vdd.n2366 vdd.n647 185
R16879 vdd.n2368 vdd.n653 185
R16880 vdd.n2532 vdd.n653 185
R16881 vdd.n2370 vdd.n2369 185
R16882 vdd.n2369 vdd.n660 185
R16883 vdd.n2371 vdd.n658 185
R16884 vdd.n2526 vdd.n658 185
R16885 vdd.n2373 vdd.n2372 185
R16886 vdd.n2374 vdd.n2373 185
R16887 vdd.n2357 vdd.n665 185
R16888 vdd.n2520 vdd.n665 185
R16889 vdd.n2356 vdd.n2355 185
R16890 vdd.n2355 vdd.n664 185
R16891 vdd.n2354 vdd.n671 185
R16892 vdd.n2514 vdd.n671 185
R16893 vdd.n2353 vdd.n2352 185
R16894 vdd.n2352 vdd.n670 185
R16895 vdd.n2351 vdd.n676 185
R16896 vdd.n2508 vdd.n676 185
R16897 vdd.n2350 vdd.n2349 185
R16898 vdd.n2349 vdd.n683 185
R16899 vdd.n2348 vdd.n681 185
R16900 vdd.n2502 vdd.n681 185
R16901 vdd.n2347 vdd.n2346 185
R16902 vdd.n2346 vdd.n690 185
R16903 vdd.n2345 vdd.n688 185
R16904 vdd.n2496 vdd.n688 185
R16905 vdd.n2344 vdd.n2343 185
R16906 vdd.n2343 vdd.n687 185
R16907 vdd.n2255 vdd.n694 185
R16908 vdd.n2490 vdd.n694 185
R16909 vdd.n2397 vdd.n2396 185
R16910 vdd.n2396 vdd.n2395 185
R16911 vdd.n2398 vdd.n699 185
R16912 vdd.n2484 vdd.n699 185
R16913 vdd.n2400 vdd.n2399 185
R16914 vdd.n2399 vdd.t195 185
R16915 vdd.n2401 vdd.n704 185
R16916 vdd.n2478 vdd.n704 185
R16917 vdd.n2480 vdd.n2479 185
R16918 vdd.n2479 vdd.n2478 185
R16919 vdd.n2481 vdd.n701 185
R16920 vdd.n701 vdd.t195 185
R16921 vdd.n2483 vdd.n2482 185
R16922 vdd.n2484 vdd.n2483 185
R16923 vdd.n693 vdd.n692 185
R16924 vdd.n2395 vdd.n693 185
R16925 vdd.n2492 vdd.n2491 185
R16926 vdd.n2491 vdd.n2490 185
R16927 vdd.n2493 vdd.n691 185
R16928 vdd.n691 vdd.n687 185
R16929 vdd.n2495 vdd.n2494 185
R16930 vdd.n2496 vdd.n2495 185
R16931 vdd.n680 vdd.n679 185
R16932 vdd.n690 vdd.n680 185
R16933 vdd.n2504 vdd.n2503 185
R16934 vdd.n2503 vdd.n2502 185
R16935 vdd.n2505 vdd.n678 185
R16936 vdd.n683 vdd.n678 185
R16937 vdd.n2507 vdd.n2506 185
R16938 vdd.n2508 vdd.n2507 185
R16939 vdd.n669 vdd.n668 185
R16940 vdd.n670 vdd.n669 185
R16941 vdd.n2516 vdd.n2515 185
R16942 vdd.n2515 vdd.n2514 185
R16943 vdd.n2517 vdd.n667 185
R16944 vdd.n667 vdd.n664 185
R16945 vdd.n2519 vdd.n2518 185
R16946 vdd.n2520 vdd.n2519 185
R16947 vdd.n657 vdd.n656 185
R16948 vdd.n2374 vdd.n657 185
R16949 vdd.n2528 vdd.n2527 185
R16950 vdd.n2527 vdd.n2526 185
R16951 vdd.n2529 vdd.n655 185
R16952 vdd.n660 vdd.n655 185
R16953 vdd.n2531 vdd.n2530 185
R16954 vdd.n2532 vdd.n2531 185
R16955 vdd.n646 vdd.n645 185
R16956 vdd.n647 vdd.n646 185
R16957 vdd.n2542 vdd.n2541 185
R16958 vdd.n2541 vdd.n2540 185
R16959 vdd.n2543 vdd.n644 185
R16960 vdd.n644 vdd.n641 185
R16961 vdd.n2545 vdd.n2544 185
R16962 vdd.n2546 vdd.n2545 185
R16963 vdd.n632 vdd.n631 185
R16964 vdd.n633 vdd.n632 185
R16965 vdd.n2599 vdd.n2598 185
R16966 vdd.n2598 vdd.n2597 185
R16967 vdd.n2600 vdd.n630 185
R16968 vdd.n636 vdd.n630 185
R16969 vdd.n2602 vdd.n2601 185
R16970 vdd.n2603 vdd.n2602 185
R16971 vdd.n600 vdd.n598 185
R16972 vdd.n598 vdd.n595 185
R16973 vdd.n2672 vdd.n2671 185
R16974 vdd.n2673 vdd.n2672 185
R16975 vdd.n2145 vdd.n2144 185
R16976 vdd.n2146 vdd.n2145 185
R16977 vdd.n754 vdd.n752 185
R16978 vdd.n752 vdd.t189 185
R16979 vdd.n2060 vdd.n761 185
R16980 vdd.n2071 vdd.n761 185
R16981 vdd.n2061 vdd.n770 185
R16982 vdd.n1770 vdd.n770 185
R16983 vdd.n2063 vdd.n2062 185
R16984 vdd.n2064 vdd.n2063 185
R16985 vdd.n2059 vdd.n769 185
R16986 vdd.n769 vdd.n766 185
R16987 vdd.n2058 vdd.n2057 185
R16988 vdd.n2057 vdd.n2056 185
R16989 vdd.n772 vdd.n771 185
R16990 vdd.n773 vdd.n772 185
R16991 vdd.n2049 vdd.n2048 185
R16992 vdd.n2050 vdd.n2049 185
R16993 vdd.n2047 vdd.n782 185
R16994 vdd.n782 vdd.n779 185
R16995 vdd.n2046 vdd.n2045 185
R16996 vdd.n2045 vdd.n2044 185
R16997 vdd.n784 vdd.n783 185
R16998 vdd.n792 vdd.n784 185
R16999 vdd.n2037 vdd.n2036 185
R17000 vdd.n2038 vdd.n2037 185
R17001 vdd.n2035 vdd.n793 185
R17002 vdd.n798 vdd.n793 185
R17003 vdd.n2034 vdd.n2033 185
R17004 vdd.n2033 vdd.n2032 185
R17005 vdd.n795 vdd.n794 185
R17006 vdd.n1871 vdd.n795 185
R17007 vdd.n2025 vdd.n2024 185
R17008 vdd.n2026 vdd.n2025 185
R17009 vdd.n2023 vdd.n805 185
R17010 vdd.n805 vdd.n802 185
R17011 vdd.n2022 vdd.n2021 185
R17012 vdd.n2021 vdd.n2020 185
R17013 vdd.n807 vdd.n806 185
R17014 vdd.n808 vdd.n807 185
R17015 vdd.n2013 vdd.n2012 185
R17016 vdd.n2014 vdd.n2013 185
R17017 vdd.n2010 vdd.n816 185
R17018 vdd.n823 vdd.n816 185
R17019 vdd.n2009 vdd.n2008 185
R17020 vdd.n2008 vdd.n2007 185
R17021 vdd.n819 vdd.n818 185
R17022 vdd.n820 vdd.n819 185
R17023 vdd.n2000 vdd.n1999 185
R17024 vdd.n2001 vdd.n2000 185
R17025 vdd.n1998 vdd.n830 185
R17026 vdd.n830 vdd.n827 185
R17027 vdd.n1997 vdd.n1996 185
R17028 vdd.n1996 vdd.n1995 185
R17029 vdd.n832 vdd.n831 185
R17030 vdd.n833 vdd.n832 185
R17031 vdd.n1988 vdd.n1987 185
R17032 vdd.n1989 vdd.n1988 185
R17033 vdd.n2076 vdd.n726 185
R17034 vdd.n2218 vdd.n726 185
R17035 vdd.n2078 vdd.n2077 185
R17036 vdd.n2080 vdd.n2079 185
R17037 vdd.n2082 vdd.n2081 185
R17038 vdd.n2084 vdd.n2083 185
R17039 vdd.n2086 vdd.n2085 185
R17040 vdd.n2088 vdd.n2087 185
R17041 vdd.n2090 vdd.n2089 185
R17042 vdd.n2092 vdd.n2091 185
R17043 vdd.n2094 vdd.n2093 185
R17044 vdd.n2096 vdd.n2095 185
R17045 vdd.n2098 vdd.n2097 185
R17046 vdd.n2100 vdd.n2099 185
R17047 vdd.n2102 vdd.n2101 185
R17048 vdd.n2104 vdd.n2103 185
R17049 vdd.n2106 vdd.n2105 185
R17050 vdd.n2108 vdd.n2107 185
R17051 vdd.n2110 vdd.n2109 185
R17052 vdd.n2112 vdd.n2111 185
R17053 vdd.n2114 vdd.n2113 185
R17054 vdd.n2116 vdd.n2115 185
R17055 vdd.n2118 vdd.n2117 185
R17056 vdd.n2120 vdd.n2119 185
R17057 vdd.n2122 vdd.n2121 185
R17058 vdd.n2124 vdd.n2123 185
R17059 vdd.n2126 vdd.n2125 185
R17060 vdd.n2128 vdd.n2127 185
R17061 vdd.n2130 vdd.n2129 185
R17062 vdd.n2132 vdd.n2131 185
R17063 vdd.n2134 vdd.n2133 185
R17064 vdd.n2136 vdd.n2135 185
R17065 vdd.n2138 vdd.n2137 185
R17066 vdd.n2140 vdd.n2139 185
R17067 vdd.n2142 vdd.n2141 185
R17068 vdd.n2143 vdd.n753 185
R17069 vdd.n2075 vdd.n751 185
R17070 vdd.n2146 vdd.n751 185
R17071 vdd.n2074 vdd.n2073 185
R17072 vdd.n2073 vdd.t189 185
R17073 vdd.n2072 vdd.n758 185
R17074 vdd.n2072 vdd.n2071 185
R17075 vdd.n1852 vdd.n759 185
R17076 vdd.n1770 vdd.n759 185
R17077 vdd.n1853 vdd.n768 185
R17078 vdd.n2064 vdd.n768 185
R17079 vdd.n1855 vdd.n1854 185
R17080 vdd.n1854 vdd.n766 185
R17081 vdd.n1856 vdd.n775 185
R17082 vdd.n2056 vdd.n775 185
R17083 vdd.n1858 vdd.n1857 185
R17084 vdd.n1857 vdd.n773 185
R17085 vdd.n1859 vdd.n781 185
R17086 vdd.n2050 vdd.n781 185
R17087 vdd.n1861 vdd.n1860 185
R17088 vdd.n1860 vdd.n779 185
R17089 vdd.n1862 vdd.n786 185
R17090 vdd.n2044 vdd.n786 185
R17091 vdd.n1864 vdd.n1863 185
R17092 vdd.n1863 vdd.n792 185
R17093 vdd.n1865 vdd.n791 185
R17094 vdd.n2038 vdd.n791 185
R17095 vdd.n1867 vdd.n1866 185
R17096 vdd.n1866 vdd.n798 185
R17097 vdd.n1868 vdd.n797 185
R17098 vdd.n2032 vdd.n797 185
R17099 vdd.n1870 vdd.n1869 185
R17100 vdd.n1871 vdd.n1870 185
R17101 vdd.n1851 vdd.n804 185
R17102 vdd.n2026 vdd.n804 185
R17103 vdd.n1850 vdd.n1849 185
R17104 vdd.n1849 vdd.n802 185
R17105 vdd.n1848 vdd.n810 185
R17106 vdd.n2020 vdd.n810 185
R17107 vdd.n1847 vdd.n1846 185
R17108 vdd.n1846 vdd.n808 185
R17109 vdd.n1845 vdd.n815 185
R17110 vdd.n2014 vdd.n815 185
R17111 vdd.n1844 vdd.n1843 185
R17112 vdd.n1843 vdd.n823 185
R17113 vdd.n1842 vdd.n822 185
R17114 vdd.n2007 vdd.n822 185
R17115 vdd.n1841 vdd.n1840 185
R17116 vdd.n1840 vdd.n820 185
R17117 vdd.n1839 vdd.n829 185
R17118 vdd.n2001 vdd.n829 185
R17119 vdd.n1838 vdd.n1837 185
R17120 vdd.n1837 vdd.n827 185
R17121 vdd.n1836 vdd.n835 185
R17122 vdd.n1995 vdd.n835 185
R17123 vdd.n1835 vdd.n1834 185
R17124 vdd.n1834 vdd.n833 185
R17125 vdd.n1833 vdd.n841 185
R17126 vdd.n1989 vdd.n841 185
R17127 vdd.n1986 vdd.n842 185
R17128 vdd.n1985 vdd.n1984 185
R17129 vdd.n1982 vdd.n843 185
R17130 vdd.n1980 vdd.n1979 185
R17131 vdd.n1978 vdd.n844 185
R17132 vdd.n1977 vdd.n1976 185
R17133 vdd.n1974 vdd.n845 185
R17134 vdd.n1972 vdd.n1971 185
R17135 vdd.n1970 vdd.n846 185
R17136 vdd.n1969 vdd.n1968 185
R17137 vdd.n1966 vdd.n847 185
R17138 vdd.n1964 vdd.n1963 185
R17139 vdd.n1962 vdd.n848 185
R17140 vdd.n1961 vdd.n1960 185
R17141 vdd.n1958 vdd.n849 185
R17142 vdd.n1956 vdd.n1955 185
R17143 vdd.n1954 vdd.n850 185
R17144 vdd.n1953 vdd.n852 185
R17145 vdd.n1798 vdd.n853 185
R17146 vdd.n1801 vdd.n1800 185
R17147 vdd.n1803 vdd.n1802 185
R17148 vdd.n1805 vdd.n1797 185
R17149 vdd.n1808 vdd.n1807 185
R17150 vdd.n1809 vdd.n1796 185
R17151 vdd.n1811 vdd.n1810 185
R17152 vdd.n1813 vdd.n1795 185
R17153 vdd.n1816 vdd.n1815 185
R17154 vdd.n1817 vdd.n1794 185
R17155 vdd.n1819 vdd.n1818 185
R17156 vdd.n1821 vdd.n1793 185
R17157 vdd.n1824 vdd.n1823 185
R17158 vdd.n1825 vdd.n1790 185
R17159 vdd.n1828 vdd.n1827 185
R17160 vdd.n1830 vdd.n1789 185
R17161 vdd.n1832 vdd.n1831 185
R17162 vdd.n1831 vdd.n839 185
R17163 vdd.n291 vdd.n290 171.744
R17164 vdd.n290 vdd.n289 171.744
R17165 vdd.n289 vdd.n258 171.744
R17166 vdd.n282 vdd.n258 171.744
R17167 vdd.n282 vdd.n281 171.744
R17168 vdd.n281 vdd.n263 171.744
R17169 vdd.n274 vdd.n263 171.744
R17170 vdd.n274 vdd.n273 171.744
R17171 vdd.n273 vdd.n267 171.744
R17172 vdd.n244 vdd.n243 171.744
R17173 vdd.n243 vdd.n242 171.744
R17174 vdd.n242 vdd.n211 171.744
R17175 vdd.n235 vdd.n211 171.744
R17176 vdd.n235 vdd.n234 171.744
R17177 vdd.n234 vdd.n216 171.744
R17178 vdd.n227 vdd.n216 171.744
R17179 vdd.n227 vdd.n226 171.744
R17180 vdd.n226 vdd.n220 171.744
R17181 vdd.n201 vdd.n200 171.744
R17182 vdd.n200 vdd.n199 171.744
R17183 vdd.n199 vdd.n168 171.744
R17184 vdd.n192 vdd.n168 171.744
R17185 vdd.n192 vdd.n191 171.744
R17186 vdd.n191 vdd.n173 171.744
R17187 vdd.n184 vdd.n173 171.744
R17188 vdd.n184 vdd.n183 171.744
R17189 vdd.n183 vdd.n177 171.744
R17190 vdd.n154 vdd.n153 171.744
R17191 vdd.n153 vdd.n152 171.744
R17192 vdd.n152 vdd.n121 171.744
R17193 vdd.n145 vdd.n121 171.744
R17194 vdd.n145 vdd.n144 171.744
R17195 vdd.n144 vdd.n126 171.744
R17196 vdd.n137 vdd.n126 171.744
R17197 vdd.n137 vdd.n136 171.744
R17198 vdd.n136 vdd.n130 171.744
R17199 vdd.n112 vdd.n111 171.744
R17200 vdd.n111 vdd.n110 171.744
R17201 vdd.n110 vdd.n79 171.744
R17202 vdd.n103 vdd.n79 171.744
R17203 vdd.n103 vdd.n102 171.744
R17204 vdd.n102 vdd.n84 171.744
R17205 vdd.n95 vdd.n84 171.744
R17206 vdd.n95 vdd.n94 171.744
R17207 vdd.n94 vdd.n88 171.744
R17208 vdd.n65 vdd.n64 171.744
R17209 vdd.n64 vdd.n63 171.744
R17210 vdd.n63 vdd.n32 171.744
R17211 vdd.n56 vdd.n32 171.744
R17212 vdd.n56 vdd.n55 171.744
R17213 vdd.n55 vdd.n37 171.744
R17214 vdd.n48 vdd.n37 171.744
R17215 vdd.n48 vdd.n47 171.744
R17216 vdd.n47 vdd.n41 171.744
R17217 vdd.n1106 vdd.n1105 171.744
R17218 vdd.n1105 vdd.n1104 171.744
R17219 vdd.n1104 vdd.n1073 171.744
R17220 vdd.n1097 vdd.n1073 171.744
R17221 vdd.n1097 vdd.n1096 171.744
R17222 vdd.n1096 vdd.n1078 171.744
R17223 vdd.n1089 vdd.n1078 171.744
R17224 vdd.n1089 vdd.n1088 171.744
R17225 vdd.n1088 vdd.n1082 171.744
R17226 vdd.n1153 vdd.n1152 171.744
R17227 vdd.n1152 vdd.n1151 171.744
R17228 vdd.n1151 vdd.n1120 171.744
R17229 vdd.n1144 vdd.n1120 171.744
R17230 vdd.n1144 vdd.n1143 171.744
R17231 vdd.n1143 vdd.n1125 171.744
R17232 vdd.n1136 vdd.n1125 171.744
R17233 vdd.n1136 vdd.n1135 171.744
R17234 vdd.n1135 vdd.n1129 171.744
R17235 vdd.n1016 vdd.n1015 171.744
R17236 vdd.n1015 vdd.n1014 171.744
R17237 vdd.n1014 vdd.n983 171.744
R17238 vdd.n1007 vdd.n983 171.744
R17239 vdd.n1007 vdd.n1006 171.744
R17240 vdd.n1006 vdd.n988 171.744
R17241 vdd.n999 vdd.n988 171.744
R17242 vdd.n999 vdd.n998 171.744
R17243 vdd.n998 vdd.n992 171.744
R17244 vdd.n1063 vdd.n1062 171.744
R17245 vdd.n1062 vdd.n1061 171.744
R17246 vdd.n1061 vdd.n1030 171.744
R17247 vdd.n1054 vdd.n1030 171.744
R17248 vdd.n1054 vdd.n1053 171.744
R17249 vdd.n1053 vdd.n1035 171.744
R17250 vdd.n1046 vdd.n1035 171.744
R17251 vdd.n1046 vdd.n1045 171.744
R17252 vdd.n1045 vdd.n1039 171.744
R17253 vdd.n927 vdd.n926 171.744
R17254 vdd.n926 vdd.n925 171.744
R17255 vdd.n925 vdd.n894 171.744
R17256 vdd.n918 vdd.n894 171.744
R17257 vdd.n918 vdd.n917 171.744
R17258 vdd.n917 vdd.n899 171.744
R17259 vdd.n910 vdd.n899 171.744
R17260 vdd.n910 vdd.n909 171.744
R17261 vdd.n909 vdd.n903 171.744
R17262 vdd.n974 vdd.n973 171.744
R17263 vdd.n973 vdd.n972 171.744
R17264 vdd.n972 vdd.n941 171.744
R17265 vdd.n965 vdd.n941 171.744
R17266 vdd.n965 vdd.n964 171.744
R17267 vdd.n964 vdd.n946 171.744
R17268 vdd.n957 vdd.n946 171.744
R17269 vdd.n957 vdd.n956 171.744
R17270 vdd.n956 vdd.n950 171.744
R17271 vdd.n3017 vdd.n334 146.341
R17272 vdd.n3015 vdd.n3014 146.341
R17273 vdd.n3012 vdd.n338 146.341
R17274 vdd.n3008 vdd.n3007 146.341
R17275 vdd.n3005 vdd.n346 146.341
R17276 vdd.n3001 vdd.n3000 146.341
R17277 vdd.n2998 vdd.n353 146.341
R17278 vdd.n2994 vdd.n2993 146.341
R17279 vdd.n2991 vdd.n360 146.341
R17280 vdd.n371 vdd.n368 146.341
R17281 vdd.n2983 vdd.n2982 146.341
R17282 vdd.n2980 vdd.n373 146.341
R17283 vdd.n2976 vdd.n2975 146.341
R17284 vdd.n2973 vdd.n379 146.341
R17285 vdd.n2969 vdd.n2968 146.341
R17286 vdd.n2966 vdd.n386 146.341
R17287 vdd.n2962 vdd.n2961 146.341
R17288 vdd.n2959 vdd.n393 146.341
R17289 vdd.n2955 vdd.n2954 146.341
R17290 vdd.n2952 vdd.n400 146.341
R17291 vdd.n411 vdd.n408 146.341
R17292 vdd.n2944 vdd.n2943 146.341
R17293 vdd.n2941 vdd.n413 146.341
R17294 vdd.n2937 vdd.n2936 146.341
R17295 vdd.n2934 vdd.n419 146.341
R17296 vdd.n2930 vdd.n2929 146.341
R17297 vdd.n2927 vdd.n426 146.341
R17298 vdd.n2923 vdd.n2922 146.341
R17299 vdd.n2920 vdd.n433 146.341
R17300 vdd.n2916 vdd.n2915 146.341
R17301 vdd.n2913 vdd.n440 146.341
R17302 vdd.n2850 vdd.n478 146.341
R17303 vdd.n2850 vdd.n474 146.341
R17304 vdd.n2856 vdd.n474 146.341
R17305 vdd.n2856 vdd.n466 146.341
R17306 vdd.n2867 vdd.n466 146.341
R17307 vdd.n2867 vdd.n462 146.341
R17308 vdd.n2873 vdd.n462 146.341
R17309 vdd.n2873 vdd.n454 146.341
R17310 vdd.n2883 vdd.n454 146.341
R17311 vdd.n2883 vdd.n455 146.341
R17312 vdd.n455 vdd.n305 146.341
R17313 vdd.n306 vdd.n305 146.341
R17314 vdd.n307 vdd.n306 146.341
R17315 vdd.n448 vdd.n307 146.341
R17316 vdd.n448 vdd.n315 146.341
R17317 vdd.n316 vdd.n315 146.341
R17318 vdd.n317 vdd.n316 146.341
R17319 vdd.n445 vdd.n317 146.341
R17320 vdd.n445 vdd.n326 146.341
R17321 vdd.n327 vdd.n326 146.341
R17322 vdd.n328 vdd.n327 146.341
R17323 vdd.n2839 vdd.n483 146.341
R17324 vdd.n2839 vdd.n517 146.341
R17325 vdd.n523 vdd.n522 146.341
R17326 vdd.n2832 vdd.n2831 146.341
R17327 vdd.n2828 vdd.n2827 146.341
R17328 vdd.n2824 vdd.n2823 146.341
R17329 vdd.n2820 vdd.n2819 146.341
R17330 vdd.n2816 vdd.n2815 146.341
R17331 vdd.n2812 vdd.n2811 146.341
R17332 vdd.n2808 vdd.n2807 146.341
R17333 vdd.n2799 vdd.n2798 146.341
R17334 vdd.n2796 vdd.n2795 146.341
R17335 vdd.n2792 vdd.n2791 146.341
R17336 vdd.n2788 vdd.n2787 146.341
R17337 vdd.n2784 vdd.n2783 146.341
R17338 vdd.n2780 vdd.n2779 146.341
R17339 vdd.n2776 vdd.n2775 146.341
R17340 vdd.n2772 vdd.n2771 146.341
R17341 vdd.n2768 vdd.n2767 146.341
R17342 vdd.n2764 vdd.n2763 146.341
R17343 vdd.n2760 vdd.n2759 146.341
R17344 vdd.n2753 vdd.n2752 146.341
R17345 vdd.n2750 vdd.n2749 146.341
R17346 vdd.n2746 vdd.n2745 146.341
R17347 vdd.n2742 vdd.n2741 146.341
R17348 vdd.n2738 vdd.n2737 146.341
R17349 vdd.n2734 vdd.n2733 146.341
R17350 vdd.n2730 vdd.n2729 146.341
R17351 vdd.n2726 vdd.n2725 146.341
R17352 vdd.n2722 vdd.n2721 146.341
R17353 vdd.n2718 vdd.n2717 146.341
R17354 vdd.n2714 vdd.n515 146.341
R17355 vdd.n2848 vdd.n479 146.341
R17356 vdd.n2848 vdd.n472 146.341
R17357 vdd.n2859 vdd.n472 146.341
R17358 vdd.n2859 vdd.n468 146.341
R17359 vdd.n2865 vdd.n468 146.341
R17360 vdd.n2865 vdd.n461 146.341
R17361 vdd.n2875 vdd.n461 146.341
R17362 vdd.n2875 vdd.n457 146.341
R17363 vdd.n2881 vdd.n457 146.341
R17364 vdd.n2881 vdd.n302 146.341
R17365 vdd.n3044 vdd.n302 146.341
R17366 vdd.n3044 vdd.n303 146.341
R17367 vdd.n3040 vdd.n303 146.341
R17368 vdd.n3040 vdd.n309 146.341
R17369 vdd.n3036 vdd.n309 146.341
R17370 vdd.n3036 vdd.n314 146.341
R17371 vdd.n3032 vdd.n314 146.341
R17372 vdd.n3032 vdd.n319 146.341
R17373 vdd.n3028 vdd.n319 146.341
R17374 vdd.n3028 vdd.n325 146.341
R17375 vdd.n3024 vdd.n325 146.341
R17376 vdd.n1936 vdd.n1935 146.341
R17377 vdd.n1933 vdd.n1517 146.341
R17378 vdd.n1713 vdd.n1523 146.341
R17379 vdd.n1711 vdd.n1710 146.341
R17380 vdd.n1708 vdd.n1525 146.341
R17381 vdd.n1704 vdd.n1703 146.341
R17382 vdd.n1701 vdd.n1532 146.341
R17383 vdd.n1697 vdd.n1696 146.341
R17384 vdd.n1694 vdd.n1539 146.341
R17385 vdd.n1550 vdd.n1547 146.341
R17386 vdd.n1686 vdd.n1685 146.341
R17387 vdd.n1683 vdd.n1552 146.341
R17388 vdd.n1679 vdd.n1678 146.341
R17389 vdd.n1676 vdd.n1558 146.341
R17390 vdd.n1672 vdd.n1671 146.341
R17391 vdd.n1669 vdd.n1565 146.341
R17392 vdd.n1665 vdd.n1664 146.341
R17393 vdd.n1662 vdd.n1572 146.341
R17394 vdd.n1658 vdd.n1657 146.341
R17395 vdd.n1655 vdd.n1579 146.341
R17396 vdd.n1590 vdd.n1587 146.341
R17397 vdd.n1647 vdd.n1646 146.341
R17398 vdd.n1644 vdd.n1592 146.341
R17399 vdd.n1640 vdd.n1639 146.341
R17400 vdd.n1637 vdd.n1598 146.341
R17401 vdd.n1633 vdd.n1632 146.341
R17402 vdd.n1630 vdd.n1605 146.341
R17403 vdd.n1626 vdd.n1625 146.341
R17404 vdd.n1623 vdd.n1620 146.341
R17405 vdd.n1618 vdd.n1615 146.341
R17406 vdd.n1613 vdd.n859 146.341
R17407 vdd.n1431 vdd.n1191 146.341
R17408 vdd.n1431 vdd.n1187 146.341
R17409 vdd.n1437 vdd.n1187 146.341
R17410 vdd.n1437 vdd.n1179 146.341
R17411 vdd.n1448 vdd.n1179 146.341
R17412 vdd.n1448 vdd.n1175 146.341
R17413 vdd.n1454 vdd.n1175 146.341
R17414 vdd.n1454 vdd.n1169 146.341
R17415 vdd.n1466 vdd.n1169 146.341
R17416 vdd.n1466 vdd.n1165 146.341
R17417 vdd.n1472 vdd.n1165 146.341
R17418 vdd.n1472 vdd.n886 146.341
R17419 vdd.n1482 vdd.n886 146.341
R17420 vdd.n1482 vdd.n882 146.341
R17421 vdd.n1488 vdd.n882 146.341
R17422 vdd.n1488 vdd.n876 146.341
R17423 vdd.n1499 vdd.n876 146.341
R17424 vdd.n1499 vdd.n871 146.341
R17425 vdd.n1507 vdd.n871 146.341
R17426 vdd.n1507 vdd.n861 146.341
R17427 vdd.n1944 vdd.n861 146.341
R17428 vdd.n1420 vdd.n1196 146.341
R17429 vdd.n1420 vdd.n1229 146.341
R17430 vdd.n1233 vdd.n1232 146.341
R17431 vdd.n1235 vdd.n1234 146.341
R17432 vdd.n1239 vdd.n1238 146.341
R17433 vdd.n1241 vdd.n1240 146.341
R17434 vdd.n1245 vdd.n1244 146.341
R17435 vdd.n1247 vdd.n1246 146.341
R17436 vdd.n1251 vdd.n1250 146.341
R17437 vdd.n1253 vdd.n1252 146.341
R17438 vdd.n1259 vdd.n1258 146.341
R17439 vdd.n1261 vdd.n1260 146.341
R17440 vdd.n1265 vdd.n1264 146.341
R17441 vdd.n1267 vdd.n1266 146.341
R17442 vdd.n1271 vdd.n1270 146.341
R17443 vdd.n1273 vdd.n1272 146.341
R17444 vdd.n1277 vdd.n1276 146.341
R17445 vdd.n1279 vdd.n1278 146.341
R17446 vdd.n1283 vdd.n1282 146.341
R17447 vdd.n1285 vdd.n1284 146.341
R17448 vdd.n1357 vdd.n1288 146.341
R17449 vdd.n1290 vdd.n1289 146.341
R17450 vdd.n1294 vdd.n1293 146.341
R17451 vdd.n1296 vdd.n1295 146.341
R17452 vdd.n1300 vdd.n1299 146.341
R17453 vdd.n1302 vdd.n1301 146.341
R17454 vdd.n1306 vdd.n1305 146.341
R17455 vdd.n1308 vdd.n1307 146.341
R17456 vdd.n1312 vdd.n1311 146.341
R17457 vdd.n1314 vdd.n1313 146.341
R17458 vdd.n1318 vdd.n1317 146.341
R17459 vdd.n1319 vdd.n1227 146.341
R17460 vdd.n1429 vdd.n1192 146.341
R17461 vdd.n1429 vdd.n1185 146.341
R17462 vdd.n1440 vdd.n1185 146.341
R17463 vdd.n1440 vdd.n1181 146.341
R17464 vdd.n1446 vdd.n1181 146.341
R17465 vdd.n1446 vdd.n1174 146.341
R17466 vdd.n1457 vdd.n1174 146.341
R17467 vdd.n1457 vdd.n1170 146.341
R17468 vdd.n1464 vdd.n1170 146.341
R17469 vdd.n1464 vdd.n1163 146.341
R17470 vdd.n1474 vdd.n1163 146.341
R17471 vdd.n1474 vdd.n889 146.341
R17472 vdd.n1480 vdd.n889 146.341
R17473 vdd.n1480 vdd.n881 146.341
R17474 vdd.n1491 vdd.n881 146.341
R17475 vdd.n1491 vdd.n877 146.341
R17476 vdd.n1497 vdd.n877 146.341
R17477 vdd.n1497 vdd.n869 146.341
R17478 vdd.n1510 vdd.n869 146.341
R17479 vdd.n1510 vdd.n864 146.341
R17480 vdd.n1942 vdd.n864 146.341
R17481 vdd.n863 vdd.n839 141.707
R17482 vdd.n2840 vdd.n484 141.707
R17483 vdd.n1791 vdd.t115 127.284
R17484 vdd.n755 vdd.t99 127.284
R17485 vdd.n1765 vdd.t140 127.284
R17486 vdd.n747 vdd.t130 127.284
R17487 vdd.n2536 vdd.t82 127.284
R17488 vdd.n2536 vdd.t83 127.284
R17489 vdd.n2256 vdd.t122 127.284
R17490 vdd.n622 vdd.t103 127.284
R17491 vdd.n2253 vdd.t108 127.284
R17492 vdd.n589 vdd.t110 127.284
R17493 vdd.n817 vdd.t118 127.284
R17494 vdd.n817 vdd.t119 127.284
R17495 vdd.n22 vdd.n20 117.314
R17496 vdd.n17 vdd.n15 117.314
R17497 vdd.n27 vdd.n26 116.927
R17498 vdd.n24 vdd.n23 116.927
R17499 vdd.n22 vdd.n21 116.927
R17500 vdd.n17 vdd.n16 116.927
R17501 vdd.n19 vdd.n18 116.927
R17502 vdd.n27 vdd.n25 116.927
R17503 vdd.n1792 vdd.t114 111.188
R17504 vdd.n756 vdd.t100 111.188
R17505 vdd.n1766 vdd.t139 111.188
R17506 vdd.n748 vdd.t131 111.188
R17507 vdd.n2257 vdd.t121 111.188
R17508 vdd.n623 vdd.t104 111.188
R17509 vdd.n2254 vdd.t107 111.188
R17510 vdd.n590 vdd.t111 111.188
R17511 vdd.n2479 vdd.n701 99.5127
R17512 vdd.n2483 vdd.n701 99.5127
R17513 vdd.n2483 vdd.n693 99.5127
R17514 vdd.n2491 vdd.n693 99.5127
R17515 vdd.n2491 vdd.n691 99.5127
R17516 vdd.n2495 vdd.n691 99.5127
R17517 vdd.n2495 vdd.n680 99.5127
R17518 vdd.n2503 vdd.n680 99.5127
R17519 vdd.n2503 vdd.n678 99.5127
R17520 vdd.n2507 vdd.n678 99.5127
R17521 vdd.n2507 vdd.n669 99.5127
R17522 vdd.n2515 vdd.n669 99.5127
R17523 vdd.n2515 vdd.n667 99.5127
R17524 vdd.n2519 vdd.n667 99.5127
R17525 vdd.n2519 vdd.n657 99.5127
R17526 vdd.n2527 vdd.n657 99.5127
R17527 vdd.n2527 vdd.n655 99.5127
R17528 vdd.n2531 vdd.n655 99.5127
R17529 vdd.n2531 vdd.n646 99.5127
R17530 vdd.n2541 vdd.n646 99.5127
R17531 vdd.n2541 vdd.n644 99.5127
R17532 vdd.n2545 vdd.n644 99.5127
R17533 vdd.n2545 vdd.n632 99.5127
R17534 vdd.n2598 vdd.n632 99.5127
R17535 vdd.n2598 vdd.n630 99.5127
R17536 vdd.n2602 vdd.n630 99.5127
R17537 vdd.n2602 vdd.n598 99.5127
R17538 vdd.n2672 vdd.n598 99.5127
R17539 vdd.n2668 vdd.n599 99.5127
R17540 vdd.n2666 vdd.n2665 99.5127
R17541 vdd.n2663 vdd.n603 99.5127
R17542 vdd.n2659 vdd.n2658 99.5127
R17543 vdd.n2656 vdd.n606 99.5127
R17544 vdd.n2652 vdd.n2651 99.5127
R17545 vdd.n2649 vdd.n609 99.5127
R17546 vdd.n2645 vdd.n2644 99.5127
R17547 vdd.n2642 vdd.n2640 99.5127
R17548 vdd.n2638 vdd.n612 99.5127
R17549 vdd.n2634 vdd.n2633 99.5127
R17550 vdd.n2631 vdd.n615 99.5127
R17551 vdd.n2627 vdd.n2626 99.5127
R17552 vdd.n2624 vdd.n618 99.5127
R17553 vdd.n2620 vdd.n2619 99.5127
R17554 vdd.n2617 vdd.n621 99.5127
R17555 vdd.n2612 vdd.n2611 99.5127
R17556 vdd.n2399 vdd.n704 99.5127
R17557 vdd.n2399 vdd.n699 99.5127
R17558 vdd.n2396 vdd.n699 99.5127
R17559 vdd.n2396 vdd.n694 99.5127
R17560 vdd.n2343 vdd.n694 99.5127
R17561 vdd.n2343 vdd.n688 99.5127
R17562 vdd.n2346 vdd.n688 99.5127
R17563 vdd.n2346 vdd.n681 99.5127
R17564 vdd.n2349 vdd.n681 99.5127
R17565 vdd.n2349 vdd.n676 99.5127
R17566 vdd.n2352 vdd.n676 99.5127
R17567 vdd.n2352 vdd.n671 99.5127
R17568 vdd.n2355 vdd.n671 99.5127
R17569 vdd.n2355 vdd.n665 99.5127
R17570 vdd.n2373 vdd.n665 99.5127
R17571 vdd.n2373 vdd.n658 99.5127
R17572 vdd.n2369 vdd.n658 99.5127
R17573 vdd.n2369 vdd.n653 99.5127
R17574 vdd.n2366 vdd.n653 99.5127
R17575 vdd.n2366 vdd.n648 99.5127
R17576 vdd.n2363 vdd.n648 99.5127
R17577 vdd.n2363 vdd.n642 99.5127
R17578 vdd.n2360 vdd.n642 99.5127
R17579 vdd.n2360 vdd.n634 99.5127
R17580 vdd.n634 vdd.n627 99.5127
R17581 vdd.n2604 vdd.n627 99.5127
R17582 vdd.n2605 vdd.n2604 99.5127
R17583 vdd.n2605 vdd.n596 99.5127
R17584 vdd.n2469 vdd.n2252 99.5127
R17585 vdd.n2465 vdd.n2252 99.5127
R17586 vdd.n2463 vdd.n2462 99.5127
R17587 vdd.n2459 vdd.n2458 99.5127
R17588 vdd.n2455 vdd.n2454 99.5127
R17589 vdd.n2451 vdd.n2450 99.5127
R17590 vdd.n2447 vdd.n2446 99.5127
R17591 vdd.n2443 vdd.n2442 99.5127
R17592 vdd.n2439 vdd.n2438 99.5127
R17593 vdd.n2435 vdd.n2434 99.5127
R17594 vdd.n2431 vdd.n2430 99.5127
R17595 vdd.n2427 vdd.n2426 99.5127
R17596 vdd.n2423 vdd.n2422 99.5127
R17597 vdd.n2419 vdd.n2418 99.5127
R17598 vdd.n2415 vdd.n2414 99.5127
R17599 vdd.n2411 vdd.n2410 99.5127
R17600 vdd.n2406 vdd.n2405 99.5127
R17601 vdd.n2217 vdd.n745 99.5127
R17602 vdd.n2213 vdd.n2212 99.5127
R17603 vdd.n2209 vdd.n2208 99.5127
R17604 vdd.n2205 vdd.n2204 99.5127
R17605 vdd.n2201 vdd.n2200 99.5127
R17606 vdd.n2197 vdd.n2196 99.5127
R17607 vdd.n2193 vdd.n2192 99.5127
R17608 vdd.n2189 vdd.n2188 99.5127
R17609 vdd.n2185 vdd.n2184 99.5127
R17610 vdd.n2181 vdd.n2180 99.5127
R17611 vdd.n2177 vdd.n2176 99.5127
R17612 vdd.n2173 vdd.n2172 99.5127
R17613 vdd.n2169 vdd.n2168 99.5127
R17614 vdd.n2165 vdd.n2164 99.5127
R17615 vdd.n2161 vdd.n2160 99.5127
R17616 vdd.n2157 vdd.n2156 99.5127
R17617 vdd.n2152 vdd.n2151 99.5127
R17618 vdd.n1890 vdd.n840 99.5127
R17619 vdd.n1890 vdd.n834 99.5127
R17620 vdd.n1887 vdd.n834 99.5127
R17621 vdd.n1887 vdd.n828 99.5127
R17622 vdd.n1884 vdd.n828 99.5127
R17623 vdd.n1884 vdd.n821 99.5127
R17624 vdd.n1881 vdd.n821 99.5127
R17625 vdd.n1881 vdd.n814 99.5127
R17626 vdd.n1878 vdd.n814 99.5127
R17627 vdd.n1878 vdd.n809 99.5127
R17628 vdd.n1875 vdd.n809 99.5127
R17629 vdd.n1875 vdd.n803 99.5127
R17630 vdd.n1872 vdd.n803 99.5127
R17631 vdd.n1872 vdd.n796 99.5127
R17632 vdd.n1786 vdd.n796 99.5127
R17633 vdd.n1786 vdd.n790 99.5127
R17634 vdd.n1783 vdd.n790 99.5127
R17635 vdd.n1783 vdd.n785 99.5127
R17636 vdd.n1780 vdd.n785 99.5127
R17637 vdd.n1780 vdd.n780 99.5127
R17638 vdd.n1777 vdd.n780 99.5127
R17639 vdd.n1777 vdd.n774 99.5127
R17640 vdd.n1774 vdd.n774 99.5127
R17641 vdd.n1774 vdd.n767 99.5127
R17642 vdd.n1771 vdd.n767 99.5127
R17643 vdd.n1771 vdd.n760 99.5127
R17644 vdd.n760 vdd.n750 99.5127
R17645 vdd.n2147 vdd.n750 99.5127
R17646 vdd.n1725 vdd.n1723 99.5127
R17647 vdd.n1729 vdd.n1723 99.5127
R17648 vdd.n1733 vdd.n1731 99.5127
R17649 vdd.n1737 vdd.n1721 99.5127
R17650 vdd.n1741 vdd.n1739 99.5127
R17651 vdd.n1745 vdd.n1719 99.5127
R17652 vdd.n1749 vdd.n1747 99.5127
R17653 vdd.n1753 vdd.n1717 99.5127
R17654 vdd.n1756 vdd.n1755 99.5127
R17655 vdd.n1926 vdd.n1924 99.5127
R17656 vdd.n1922 vdd.n1758 99.5127
R17657 vdd.n1918 vdd.n1916 99.5127
R17658 vdd.n1914 vdd.n1760 99.5127
R17659 vdd.n1910 vdd.n1908 99.5127
R17660 vdd.n1906 vdd.n1762 99.5127
R17661 vdd.n1902 vdd.n1900 99.5127
R17662 vdd.n1898 vdd.n1764 99.5127
R17663 vdd.n1990 vdd.n836 99.5127
R17664 vdd.n1994 vdd.n836 99.5127
R17665 vdd.n1994 vdd.n826 99.5127
R17666 vdd.n2002 vdd.n826 99.5127
R17667 vdd.n2002 vdd.n824 99.5127
R17668 vdd.n2006 vdd.n824 99.5127
R17669 vdd.n2006 vdd.n813 99.5127
R17670 vdd.n2015 vdd.n813 99.5127
R17671 vdd.n2015 vdd.n811 99.5127
R17672 vdd.n2019 vdd.n811 99.5127
R17673 vdd.n2019 vdd.n801 99.5127
R17674 vdd.n2027 vdd.n801 99.5127
R17675 vdd.n2027 vdd.n799 99.5127
R17676 vdd.n2031 vdd.n799 99.5127
R17677 vdd.n2031 vdd.n789 99.5127
R17678 vdd.n2039 vdd.n789 99.5127
R17679 vdd.n2039 vdd.n787 99.5127
R17680 vdd.n2043 vdd.n787 99.5127
R17681 vdd.n2043 vdd.n778 99.5127
R17682 vdd.n2051 vdd.n778 99.5127
R17683 vdd.n2051 vdd.n776 99.5127
R17684 vdd.n2055 vdd.n776 99.5127
R17685 vdd.n2055 vdd.n765 99.5127
R17686 vdd.n2065 vdd.n765 99.5127
R17687 vdd.n2065 vdd.n762 99.5127
R17688 vdd.n2070 vdd.n762 99.5127
R17689 vdd.n2070 vdd.n763 99.5127
R17690 vdd.n763 vdd.n744 99.5127
R17691 vdd.n2588 vdd.n2587 99.5127
R17692 vdd.n2585 vdd.n2551 99.5127
R17693 vdd.n2581 vdd.n2580 99.5127
R17694 vdd.n2578 vdd.n2554 99.5127
R17695 vdd.n2574 vdd.n2573 99.5127
R17696 vdd.n2571 vdd.n2557 99.5127
R17697 vdd.n2567 vdd.n2566 99.5127
R17698 vdd.n2564 vdd.n2561 99.5127
R17699 vdd.n2705 vdd.n577 99.5127
R17700 vdd.n2703 vdd.n2702 99.5127
R17701 vdd.n2700 vdd.n579 99.5127
R17702 vdd.n2696 vdd.n2695 99.5127
R17703 vdd.n2693 vdd.n582 99.5127
R17704 vdd.n2689 vdd.n2688 99.5127
R17705 vdd.n2686 vdd.n585 99.5127
R17706 vdd.n2682 vdd.n2681 99.5127
R17707 vdd.n2679 vdd.n588 99.5127
R17708 vdd.n2323 vdd.n705 99.5127
R17709 vdd.n2323 vdd.n700 99.5127
R17710 vdd.n2394 vdd.n700 99.5127
R17711 vdd.n2394 vdd.n695 99.5127
R17712 vdd.n2390 vdd.n695 99.5127
R17713 vdd.n2390 vdd.n689 99.5127
R17714 vdd.n2387 vdd.n689 99.5127
R17715 vdd.n2387 vdd.n682 99.5127
R17716 vdd.n2384 vdd.n682 99.5127
R17717 vdd.n2384 vdd.n677 99.5127
R17718 vdd.n2381 vdd.n677 99.5127
R17719 vdd.n2381 vdd.n672 99.5127
R17720 vdd.n2378 vdd.n672 99.5127
R17721 vdd.n2378 vdd.n666 99.5127
R17722 vdd.n2375 vdd.n666 99.5127
R17723 vdd.n2375 vdd.n659 99.5127
R17724 vdd.n2340 vdd.n659 99.5127
R17725 vdd.n2340 vdd.n654 99.5127
R17726 vdd.n2337 vdd.n654 99.5127
R17727 vdd.n2337 vdd.n649 99.5127
R17728 vdd.n2334 vdd.n649 99.5127
R17729 vdd.n2334 vdd.n643 99.5127
R17730 vdd.n2331 vdd.n643 99.5127
R17731 vdd.n2331 vdd.n635 99.5127
R17732 vdd.n2328 vdd.n635 99.5127
R17733 vdd.n2328 vdd.n628 99.5127
R17734 vdd.n628 vdd.n594 99.5127
R17735 vdd.n2674 vdd.n594 99.5127
R17736 vdd.n2473 vdd.n708 99.5127
R17737 vdd.n2261 vdd.n2260 99.5127
R17738 vdd.n2265 vdd.n2264 99.5127
R17739 vdd.n2269 vdd.n2268 99.5127
R17740 vdd.n2273 vdd.n2272 99.5127
R17741 vdd.n2277 vdd.n2276 99.5127
R17742 vdd.n2281 vdd.n2280 99.5127
R17743 vdd.n2285 vdd.n2284 99.5127
R17744 vdd.n2289 vdd.n2288 99.5127
R17745 vdd.n2293 vdd.n2292 99.5127
R17746 vdd.n2297 vdd.n2296 99.5127
R17747 vdd.n2301 vdd.n2300 99.5127
R17748 vdd.n2305 vdd.n2304 99.5127
R17749 vdd.n2309 vdd.n2308 99.5127
R17750 vdd.n2313 vdd.n2312 99.5127
R17751 vdd.n2317 vdd.n2316 99.5127
R17752 vdd.n2319 vdd.n2251 99.5127
R17753 vdd.n2477 vdd.n698 99.5127
R17754 vdd.n2485 vdd.n698 99.5127
R17755 vdd.n2485 vdd.n696 99.5127
R17756 vdd.n2489 vdd.n696 99.5127
R17757 vdd.n2489 vdd.n686 99.5127
R17758 vdd.n2497 vdd.n686 99.5127
R17759 vdd.n2497 vdd.n684 99.5127
R17760 vdd.n2501 vdd.n684 99.5127
R17761 vdd.n2501 vdd.n675 99.5127
R17762 vdd.n2509 vdd.n675 99.5127
R17763 vdd.n2509 vdd.n673 99.5127
R17764 vdd.n2513 vdd.n673 99.5127
R17765 vdd.n2513 vdd.n663 99.5127
R17766 vdd.n2521 vdd.n663 99.5127
R17767 vdd.n2521 vdd.n661 99.5127
R17768 vdd.n2525 vdd.n661 99.5127
R17769 vdd.n2525 vdd.n652 99.5127
R17770 vdd.n2533 vdd.n652 99.5127
R17771 vdd.n2533 vdd.n650 99.5127
R17772 vdd.n2539 vdd.n650 99.5127
R17773 vdd.n2539 vdd.n640 99.5127
R17774 vdd.n2547 vdd.n640 99.5127
R17775 vdd.n2547 vdd.n637 99.5127
R17776 vdd.n2596 vdd.n637 99.5127
R17777 vdd.n2596 vdd.n638 99.5127
R17778 vdd.n638 vdd.n629 99.5127
R17779 vdd.n2591 vdd.n629 99.5127
R17780 vdd.n2591 vdd.n597 99.5127
R17781 vdd.n2141 vdd.n2140 99.5127
R17782 vdd.n2137 vdd.n2136 99.5127
R17783 vdd.n2133 vdd.n2132 99.5127
R17784 vdd.n2129 vdd.n2128 99.5127
R17785 vdd.n2125 vdd.n2124 99.5127
R17786 vdd.n2121 vdd.n2120 99.5127
R17787 vdd.n2117 vdd.n2116 99.5127
R17788 vdd.n2113 vdd.n2112 99.5127
R17789 vdd.n2109 vdd.n2108 99.5127
R17790 vdd.n2105 vdd.n2104 99.5127
R17791 vdd.n2101 vdd.n2100 99.5127
R17792 vdd.n2097 vdd.n2096 99.5127
R17793 vdd.n2093 vdd.n2092 99.5127
R17794 vdd.n2089 vdd.n2088 99.5127
R17795 vdd.n2085 vdd.n2084 99.5127
R17796 vdd.n2081 vdd.n2080 99.5127
R17797 vdd.n2077 vdd.n726 99.5127
R17798 vdd.n1834 vdd.n841 99.5127
R17799 vdd.n1834 vdd.n835 99.5127
R17800 vdd.n1837 vdd.n835 99.5127
R17801 vdd.n1837 vdd.n829 99.5127
R17802 vdd.n1840 vdd.n829 99.5127
R17803 vdd.n1840 vdd.n822 99.5127
R17804 vdd.n1843 vdd.n822 99.5127
R17805 vdd.n1843 vdd.n815 99.5127
R17806 vdd.n1846 vdd.n815 99.5127
R17807 vdd.n1846 vdd.n810 99.5127
R17808 vdd.n1849 vdd.n810 99.5127
R17809 vdd.n1849 vdd.n804 99.5127
R17810 vdd.n1870 vdd.n804 99.5127
R17811 vdd.n1870 vdd.n797 99.5127
R17812 vdd.n1866 vdd.n797 99.5127
R17813 vdd.n1866 vdd.n791 99.5127
R17814 vdd.n1863 vdd.n791 99.5127
R17815 vdd.n1863 vdd.n786 99.5127
R17816 vdd.n1860 vdd.n786 99.5127
R17817 vdd.n1860 vdd.n781 99.5127
R17818 vdd.n1857 vdd.n781 99.5127
R17819 vdd.n1857 vdd.n775 99.5127
R17820 vdd.n1854 vdd.n775 99.5127
R17821 vdd.n1854 vdd.n768 99.5127
R17822 vdd.n768 vdd.n759 99.5127
R17823 vdd.n2072 vdd.n759 99.5127
R17824 vdd.n2073 vdd.n2072 99.5127
R17825 vdd.n2073 vdd.n751 99.5127
R17826 vdd.n1984 vdd.n1982 99.5127
R17827 vdd.n1980 vdd.n844 99.5127
R17828 vdd.n1976 vdd.n1974 99.5127
R17829 vdd.n1972 vdd.n846 99.5127
R17830 vdd.n1968 vdd.n1966 99.5127
R17831 vdd.n1964 vdd.n848 99.5127
R17832 vdd.n1960 vdd.n1958 99.5127
R17833 vdd.n1956 vdd.n850 99.5127
R17834 vdd.n1798 vdd.n852 99.5127
R17835 vdd.n1803 vdd.n1800 99.5127
R17836 vdd.n1807 vdd.n1805 99.5127
R17837 vdd.n1811 vdd.n1796 99.5127
R17838 vdd.n1815 vdd.n1813 99.5127
R17839 vdd.n1819 vdd.n1794 99.5127
R17840 vdd.n1823 vdd.n1821 99.5127
R17841 vdd.n1828 vdd.n1790 99.5127
R17842 vdd.n1831 vdd.n1830 99.5127
R17843 vdd.n1988 vdd.n832 99.5127
R17844 vdd.n1996 vdd.n832 99.5127
R17845 vdd.n1996 vdd.n830 99.5127
R17846 vdd.n2000 vdd.n830 99.5127
R17847 vdd.n2000 vdd.n819 99.5127
R17848 vdd.n2008 vdd.n819 99.5127
R17849 vdd.n2008 vdd.n816 99.5127
R17850 vdd.n2013 vdd.n816 99.5127
R17851 vdd.n2013 vdd.n807 99.5127
R17852 vdd.n2021 vdd.n807 99.5127
R17853 vdd.n2021 vdd.n805 99.5127
R17854 vdd.n2025 vdd.n805 99.5127
R17855 vdd.n2025 vdd.n795 99.5127
R17856 vdd.n2033 vdd.n795 99.5127
R17857 vdd.n2033 vdd.n793 99.5127
R17858 vdd.n2037 vdd.n793 99.5127
R17859 vdd.n2037 vdd.n784 99.5127
R17860 vdd.n2045 vdd.n784 99.5127
R17861 vdd.n2045 vdd.n782 99.5127
R17862 vdd.n2049 vdd.n782 99.5127
R17863 vdd.n2049 vdd.n772 99.5127
R17864 vdd.n2057 vdd.n772 99.5127
R17865 vdd.n2057 vdd.n769 99.5127
R17866 vdd.n2063 vdd.n769 99.5127
R17867 vdd.n2063 vdd.n770 99.5127
R17868 vdd.n770 vdd.n761 99.5127
R17869 vdd.n761 vdd.n752 99.5127
R17870 vdd.n2145 vdd.n752 99.5127
R17871 vdd.n9 vdd.n7 98.9633
R17872 vdd.n2 vdd.n0 98.9633
R17873 vdd.n9 vdd.n8 98.6055
R17874 vdd.n11 vdd.n10 98.6055
R17875 vdd.n13 vdd.n12 98.6055
R17876 vdd.n6 vdd.n5 98.6055
R17877 vdd.n4 vdd.n3 98.6055
R17878 vdd.n2 vdd.n1 98.6055
R17879 vdd.t25 vdd.n267 85.8723
R17880 vdd.t36 vdd.n220 85.8723
R17881 vdd.t21 vdd.n177 85.8723
R17882 vdd.t31 vdd.n130 85.8723
R17883 vdd.t62 vdd.n88 85.8723
R17884 vdd.t4 vdd.n41 85.8723
R17885 vdd.t60 vdd.n1082 85.8723
R17886 vdd.t46 vdd.n1129 85.8723
R17887 vdd.t52 vdd.n992 85.8723
R17888 vdd.t39 vdd.n1039 85.8723
R17889 vdd.t2 vdd.n903 85.8723
R17890 vdd.t61 vdd.n950 85.8723
R17891 vdd.n2537 vdd.n2536 78.546
R17892 vdd.n2011 vdd.n817 78.546
R17893 vdd.n254 vdd.n253 75.1835
R17894 vdd.n252 vdd.n251 75.1835
R17895 vdd.n250 vdd.n249 75.1835
R17896 vdd.n164 vdd.n163 75.1835
R17897 vdd.n162 vdd.n161 75.1835
R17898 vdd.n160 vdd.n159 75.1835
R17899 vdd.n75 vdd.n74 75.1835
R17900 vdd.n73 vdd.n72 75.1835
R17901 vdd.n71 vdd.n70 75.1835
R17902 vdd.n1112 vdd.n1111 75.1835
R17903 vdd.n1114 vdd.n1113 75.1835
R17904 vdd.n1116 vdd.n1115 75.1835
R17905 vdd.n1022 vdd.n1021 75.1835
R17906 vdd.n1024 vdd.n1023 75.1835
R17907 vdd.n1026 vdd.n1025 75.1835
R17908 vdd.n933 vdd.n932 75.1835
R17909 vdd.n935 vdd.n934 75.1835
R17910 vdd.n937 vdd.n936 75.1835
R17911 vdd.n2472 vdd.n2471 72.8958
R17912 vdd.n2471 vdd.n2235 72.8958
R17913 vdd.n2471 vdd.n2236 72.8958
R17914 vdd.n2471 vdd.n2237 72.8958
R17915 vdd.n2471 vdd.n2238 72.8958
R17916 vdd.n2471 vdd.n2239 72.8958
R17917 vdd.n2471 vdd.n2240 72.8958
R17918 vdd.n2471 vdd.n2241 72.8958
R17919 vdd.n2471 vdd.n2242 72.8958
R17920 vdd.n2471 vdd.n2243 72.8958
R17921 vdd.n2471 vdd.n2244 72.8958
R17922 vdd.n2471 vdd.n2245 72.8958
R17923 vdd.n2471 vdd.n2246 72.8958
R17924 vdd.n2471 vdd.n2247 72.8958
R17925 vdd.n2471 vdd.n2248 72.8958
R17926 vdd.n2471 vdd.n2249 72.8958
R17927 vdd.n2471 vdd.n2250 72.8958
R17928 vdd.n593 vdd.n484 72.8958
R17929 vdd.n2680 vdd.n484 72.8958
R17930 vdd.n587 vdd.n484 72.8958
R17931 vdd.n2687 vdd.n484 72.8958
R17932 vdd.n584 vdd.n484 72.8958
R17933 vdd.n2694 vdd.n484 72.8958
R17934 vdd.n581 vdd.n484 72.8958
R17935 vdd.n2701 vdd.n484 72.8958
R17936 vdd.n2704 vdd.n484 72.8958
R17937 vdd.n2560 vdd.n484 72.8958
R17938 vdd.n2565 vdd.n484 72.8958
R17939 vdd.n2559 vdd.n484 72.8958
R17940 vdd.n2572 vdd.n484 72.8958
R17941 vdd.n2556 vdd.n484 72.8958
R17942 vdd.n2579 vdd.n484 72.8958
R17943 vdd.n2553 vdd.n484 72.8958
R17944 vdd.n2586 vdd.n484 72.8958
R17945 vdd.n1724 vdd.n839 72.8958
R17946 vdd.n1730 vdd.n839 72.8958
R17947 vdd.n1732 vdd.n839 72.8958
R17948 vdd.n1738 vdd.n839 72.8958
R17949 vdd.n1740 vdd.n839 72.8958
R17950 vdd.n1746 vdd.n839 72.8958
R17951 vdd.n1748 vdd.n839 72.8958
R17952 vdd.n1754 vdd.n839 72.8958
R17953 vdd.n1925 vdd.n839 72.8958
R17954 vdd.n1923 vdd.n839 72.8958
R17955 vdd.n1917 vdd.n839 72.8958
R17956 vdd.n1915 vdd.n839 72.8958
R17957 vdd.n1909 vdd.n839 72.8958
R17958 vdd.n1907 vdd.n839 72.8958
R17959 vdd.n1901 vdd.n839 72.8958
R17960 vdd.n1899 vdd.n839 72.8958
R17961 vdd.n1893 vdd.n839 72.8958
R17962 vdd.n2218 vdd.n727 72.8958
R17963 vdd.n2218 vdd.n728 72.8958
R17964 vdd.n2218 vdd.n729 72.8958
R17965 vdd.n2218 vdd.n730 72.8958
R17966 vdd.n2218 vdd.n731 72.8958
R17967 vdd.n2218 vdd.n732 72.8958
R17968 vdd.n2218 vdd.n733 72.8958
R17969 vdd.n2218 vdd.n734 72.8958
R17970 vdd.n2218 vdd.n735 72.8958
R17971 vdd.n2218 vdd.n736 72.8958
R17972 vdd.n2218 vdd.n737 72.8958
R17973 vdd.n2218 vdd.n738 72.8958
R17974 vdd.n2218 vdd.n739 72.8958
R17975 vdd.n2218 vdd.n740 72.8958
R17976 vdd.n2218 vdd.n741 72.8958
R17977 vdd.n2218 vdd.n742 72.8958
R17978 vdd.n2218 vdd.n743 72.8958
R17979 vdd.n2471 vdd.n2470 72.8958
R17980 vdd.n2471 vdd.n2219 72.8958
R17981 vdd.n2471 vdd.n2220 72.8958
R17982 vdd.n2471 vdd.n2221 72.8958
R17983 vdd.n2471 vdd.n2222 72.8958
R17984 vdd.n2471 vdd.n2223 72.8958
R17985 vdd.n2471 vdd.n2224 72.8958
R17986 vdd.n2471 vdd.n2225 72.8958
R17987 vdd.n2471 vdd.n2226 72.8958
R17988 vdd.n2471 vdd.n2227 72.8958
R17989 vdd.n2471 vdd.n2228 72.8958
R17990 vdd.n2471 vdd.n2229 72.8958
R17991 vdd.n2471 vdd.n2230 72.8958
R17992 vdd.n2471 vdd.n2231 72.8958
R17993 vdd.n2471 vdd.n2232 72.8958
R17994 vdd.n2471 vdd.n2233 72.8958
R17995 vdd.n2471 vdd.n2234 72.8958
R17996 vdd.n2610 vdd.n484 72.8958
R17997 vdd.n625 vdd.n484 72.8958
R17998 vdd.n2618 vdd.n484 72.8958
R17999 vdd.n620 vdd.n484 72.8958
R18000 vdd.n2625 vdd.n484 72.8958
R18001 vdd.n617 vdd.n484 72.8958
R18002 vdd.n2632 vdd.n484 72.8958
R18003 vdd.n614 vdd.n484 72.8958
R18004 vdd.n2639 vdd.n484 72.8958
R18005 vdd.n2643 vdd.n484 72.8958
R18006 vdd.n611 vdd.n484 72.8958
R18007 vdd.n2650 vdd.n484 72.8958
R18008 vdd.n608 vdd.n484 72.8958
R18009 vdd.n2657 vdd.n484 72.8958
R18010 vdd.n605 vdd.n484 72.8958
R18011 vdd.n2664 vdd.n484 72.8958
R18012 vdd.n2667 vdd.n484 72.8958
R18013 vdd.n2218 vdd.n725 72.8958
R18014 vdd.n2218 vdd.n724 72.8958
R18015 vdd.n2218 vdd.n723 72.8958
R18016 vdd.n2218 vdd.n722 72.8958
R18017 vdd.n2218 vdd.n721 72.8958
R18018 vdd.n2218 vdd.n720 72.8958
R18019 vdd.n2218 vdd.n719 72.8958
R18020 vdd.n2218 vdd.n718 72.8958
R18021 vdd.n2218 vdd.n717 72.8958
R18022 vdd.n2218 vdd.n716 72.8958
R18023 vdd.n2218 vdd.n715 72.8958
R18024 vdd.n2218 vdd.n714 72.8958
R18025 vdd.n2218 vdd.n713 72.8958
R18026 vdd.n2218 vdd.n712 72.8958
R18027 vdd.n2218 vdd.n711 72.8958
R18028 vdd.n2218 vdd.n710 72.8958
R18029 vdd.n2218 vdd.n709 72.8958
R18030 vdd.n1983 vdd.n839 72.8958
R18031 vdd.n1981 vdd.n839 72.8958
R18032 vdd.n1975 vdd.n839 72.8958
R18033 vdd.n1973 vdd.n839 72.8958
R18034 vdd.n1967 vdd.n839 72.8958
R18035 vdd.n1965 vdd.n839 72.8958
R18036 vdd.n1959 vdd.n839 72.8958
R18037 vdd.n1957 vdd.n839 72.8958
R18038 vdd.n851 vdd.n839 72.8958
R18039 vdd.n1799 vdd.n839 72.8958
R18040 vdd.n1804 vdd.n839 72.8958
R18041 vdd.n1806 vdd.n839 72.8958
R18042 vdd.n1812 vdd.n839 72.8958
R18043 vdd.n1814 vdd.n839 72.8958
R18044 vdd.n1820 vdd.n839 72.8958
R18045 vdd.n1822 vdd.n839 72.8958
R18046 vdd.n1829 vdd.n839 72.8958
R18047 vdd.n1422 vdd.n1421 66.2847
R18048 vdd.n1421 vdd.n1197 66.2847
R18049 vdd.n1421 vdd.n1198 66.2847
R18050 vdd.n1421 vdd.n1199 66.2847
R18051 vdd.n1421 vdd.n1200 66.2847
R18052 vdd.n1421 vdd.n1201 66.2847
R18053 vdd.n1421 vdd.n1202 66.2847
R18054 vdd.n1421 vdd.n1203 66.2847
R18055 vdd.n1421 vdd.n1204 66.2847
R18056 vdd.n1421 vdd.n1205 66.2847
R18057 vdd.n1421 vdd.n1206 66.2847
R18058 vdd.n1421 vdd.n1207 66.2847
R18059 vdd.n1421 vdd.n1208 66.2847
R18060 vdd.n1421 vdd.n1209 66.2847
R18061 vdd.n1421 vdd.n1210 66.2847
R18062 vdd.n1421 vdd.n1211 66.2847
R18063 vdd.n1421 vdd.n1212 66.2847
R18064 vdd.n1421 vdd.n1213 66.2847
R18065 vdd.n1421 vdd.n1214 66.2847
R18066 vdd.n1421 vdd.n1215 66.2847
R18067 vdd.n1421 vdd.n1216 66.2847
R18068 vdd.n1421 vdd.n1217 66.2847
R18069 vdd.n1421 vdd.n1218 66.2847
R18070 vdd.n1421 vdd.n1219 66.2847
R18071 vdd.n1421 vdd.n1220 66.2847
R18072 vdd.n1421 vdd.n1221 66.2847
R18073 vdd.n1421 vdd.n1222 66.2847
R18074 vdd.n1421 vdd.n1223 66.2847
R18075 vdd.n1421 vdd.n1224 66.2847
R18076 vdd.n1421 vdd.n1225 66.2847
R18077 vdd.n1421 vdd.n1226 66.2847
R18078 vdd.n863 vdd.n860 66.2847
R18079 vdd.n1614 vdd.n863 66.2847
R18080 vdd.n1619 vdd.n863 66.2847
R18081 vdd.n1624 vdd.n863 66.2847
R18082 vdd.n1612 vdd.n863 66.2847
R18083 vdd.n1631 vdd.n863 66.2847
R18084 vdd.n1604 vdd.n863 66.2847
R18085 vdd.n1638 vdd.n863 66.2847
R18086 vdd.n1597 vdd.n863 66.2847
R18087 vdd.n1645 vdd.n863 66.2847
R18088 vdd.n1591 vdd.n863 66.2847
R18089 vdd.n1586 vdd.n863 66.2847
R18090 vdd.n1656 vdd.n863 66.2847
R18091 vdd.n1578 vdd.n863 66.2847
R18092 vdd.n1663 vdd.n863 66.2847
R18093 vdd.n1571 vdd.n863 66.2847
R18094 vdd.n1670 vdd.n863 66.2847
R18095 vdd.n1564 vdd.n863 66.2847
R18096 vdd.n1677 vdd.n863 66.2847
R18097 vdd.n1557 vdd.n863 66.2847
R18098 vdd.n1684 vdd.n863 66.2847
R18099 vdd.n1551 vdd.n863 66.2847
R18100 vdd.n1546 vdd.n863 66.2847
R18101 vdd.n1695 vdd.n863 66.2847
R18102 vdd.n1538 vdd.n863 66.2847
R18103 vdd.n1702 vdd.n863 66.2847
R18104 vdd.n1531 vdd.n863 66.2847
R18105 vdd.n1709 vdd.n863 66.2847
R18106 vdd.n1712 vdd.n863 66.2847
R18107 vdd.n1522 vdd.n863 66.2847
R18108 vdd.n1934 vdd.n863 66.2847
R18109 vdd.n1516 vdd.n863 66.2847
R18110 vdd.n2841 vdd.n2840 66.2847
R18111 vdd.n2840 vdd.n485 66.2847
R18112 vdd.n2840 vdd.n486 66.2847
R18113 vdd.n2840 vdd.n487 66.2847
R18114 vdd.n2840 vdd.n488 66.2847
R18115 vdd.n2840 vdd.n489 66.2847
R18116 vdd.n2840 vdd.n490 66.2847
R18117 vdd.n2840 vdd.n491 66.2847
R18118 vdd.n2840 vdd.n492 66.2847
R18119 vdd.n2840 vdd.n493 66.2847
R18120 vdd.n2840 vdd.n494 66.2847
R18121 vdd.n2840 vdd.n495 66.2847
R18122 vdd.n2840 vdd.n496 66.2847
R18123 vdd.n2840 vdd.n497 66.2847
R18124 vdd.n2840 vdd.n498 66.2847
R18125 vdd.n2840 vdd.n499 66.2847
R18126 vdd.n2840 vdd.n500 66.2847
R18127 vdd.n2840 vdd.n501 66.2847
R18128 vdd.n2840 vdd.n502 66.2847
R18129 vdd.n2840 vdd.n503 66.2847
R18130 vdd.n2840 vdd.n504 66.2847
R18131 vdd.n2840 vdd.n505 66.2847
R18132 vdd.n2840 vdd.n506 66.2847
R18133 vdd.n2840 vdd.n507 66.2847
R18134 vdd.n2840 vdd.n508 66.2847
R18135 vdd.n2840 vdd.n509 66.2847
R18136 vdd.n2840 vdd.n510 66.2847
R18137 vdd.n2840 vdd.n511 66.2847
R18138 vdd.n2840 vdd.n512 66.2847
R18139 vdd.n2840 vdd.n513 66.2847
R18140 vdd.n2840 vdd.n514 66.2847
R18141 vdd.n2905 vdd.n329 66.2847
R18142 vdd.n2914 vdd.n329 66.2847
R18143 vdd.n439 vdd.n329 66.2847
R18144 vdd.n2921 vdd.n329 66.2847
R18145 vdd.n432 vdd.n329 66.2847
R18146 vdd.n2928 vdd.n329 66.2847
R18147 vdd.n425 vdd.n329 66.2847
R18148 vdd.n2935 vdd.n329 66.2847
R18149 vdd.n418 vdd.n329 66.2847
R18150 vdd.n2942 vdd.n329 66.2847
R18151 vdd.n412 vdd.n329 66.2847
R18152 vdd.n407 vdd.n329 66.2847
R18153 vdd.n2953 vdd.n329 66.2847
R18154 vdd.n399 vdd.n329 66.2847
R18155 vdd.n2960 vdd.n329 66.2847
R18156 vdd.n392 vdd.n329 66.2847
R18157 vdd.n2967 vdd.n329 66.2847
R18158 vdd.n385 vdd.n329 66.2847
R18159 vdd.n2974 vdd.n329 66.2847
R18160 vdd.n378 vdd.n329 66.2847
R18161 vdd.n2981 vdd.n329 66.2847
R18162 vdd.n372 vdd.n329 66.2847
R18163 vdd.n367 vdd.n329 66.2847
R18164 vdd.n2992 vdd.n329 66.2847
R18165 vdd.n359 vdd.n329 66.2847
R18166 vdd.n2999 vdd.n329 66.2847
R18167 vdd.n352 vdd.n329 66.2847
R18168 vdd.n3006 vdd.n329 66.2847
R18169 vdd.n345 vdd.n329 66.2847
R18170 vdd.n3013 vdd.n329 66.2847
R18171 vdd.n3016 vdd.n329 66.2847
R18172 vdd.n333 vdd.n329 66.2847
R18173 vdd.n334 vdd.n333 52.4337
R18174 vdd.n3016 vdd.n3015 52.4337
R18175 vdd.n3013 vdd.n3012 52.4337
R18176 vdd.n3008 vdd.n345 52.4337
R18177 vdd.n3006 vdd.n3005 52.4337
R18178 vdd.n3001 vdd.n352 52.4337
R18179 vdd.n2999 vdd.n2998 52.4337
R18180 vdd.n2994 vdd.n359 52.4337
R18181 vdd.n2992 vdd.n2991 52.4337
R18182 vdd.n368 vdd.n367 52.4337
R18183 vdd.n2983 vdd.n372 52.4337
R18184 vdd.n2981 vdd.n2980 52.4337
R18185 vdd.n2976 vdd.n378 52.4337
R18186 vdd.n2974 vdd.n2973 52.4337
R18187 vdd.n2969 vdd.n385 52.4337
R18188 vdd.n2967 vdd.n2966 52.4337
R18189 vdd.n2962 vdd.n392 52.4337
R18190 vdd.n2960 vdd.n2959 52.4337
R18191 vdd.n2955 vdd.n399 52.4337
R18192 vdd.n2953 vdd.n2952 52.4337
R18193 vdd.n408 vdd.n407 52.4337
R18194 vdd.n2944 vdd.n412 52.4337
R18195 vdd.n2942 vdd.n2941 52.4337
R18196 vdd.n2937 vdd.n418 52.4337
R18197 vdd.n2935 vdd.n2934 52.4337
R18198 vdd.n2930 vdd.n425 52.4337
R18199 vdd.n2928 vdd.n2927 52.4337
R18200 vdd.n2923 vdd.n432 52.4337
R18201 vdd.n2921 vdd.n2920 52.4337
R18202 vdd.n2916 vdd.n439 52.4337
R18203 vdd.n2914 vdd.n2913 52.4337
R18204 vdd.n2906 vdd.n2905 52.4337
R18205 vdd.n2842 vdd.n2841 52.4337
R18206 vdd.n517 vdd.n485 52.4337
R18207 vdd.n523 vdd.n486 52.4337
R18208 vdd.n2831 vdd.n487 52.4337
R18209 vdd.n2827 vdd.n488 52.4337
R18210 vdd.n2823 vdd.n489 52.4337
R18211 vdd.n2819 vdd.n490 52.4337
R18212 vdd.n2815 vdd.n491 52.4337
R18213 vdd.n2811 vdd.n492 52.4337
R18214 vdd.n2807 vdd.n493 52.4337
R18215 vdd.n2799 vdd.n494 52.4337
R18216 vdd.n2795 vdd.n495 52.4337
R18217 vdd.n2791 vdd.n496 52.4337
R18218 vdd.n2787 vdd.n497 52.4337
R18219 vdd.n2783 vdd.n498 52.4337
R18220 vdd.n2779 vdd.n499 52.4337
R18221 vdd.n2775 vdd.n500 52.4337
R18222 vdd.n2771 vdd.n501 52.4337
R18223 vdd.n2767 vdd.n502 52.4337
R18224 vdd.n2763 vdd.n503 52.4337
R18225 vdd.n2759 vdd.n504 52.4337
R18226 vdd.n2753 vdd.n505 52.4337
R18227 vdd.n2749 vdd.n506 52.4337
R18228 vdd.n2745 vdd.n507 52.4337
R18229 vdd.n2741 vdd.n508 52.4337
R18230 vdd.n2737 vdd.n509 52.4337
R18231 vdd.n2733 vdd.n510 52.4337
R18232 vdd.n2729 vdd.n511 52.4337
R18233 vdd.n2725 vdd.n512 52.4337
R18234 vdd.n2721 vdd.n513 52.4337
R18235 vdd.n2717 vdd.n514 52.4337
R18236 vdd.n1936 vdd.n1516 52.4337
R18237 vdd.n1934 vdd.n1933 52.4337
R18238 vdd.n1523 vdd.n1522 52.4337
R18239 vdd.n1712 vdd.n1711 52.4337
R18240 vdd.n1709 vdd.n1708 52.4337
R18241 vdd.n1704 vdd.n1531 52.4337
R18242 vdd.n1702 vdd.n1701 52.4337
R18243 vdd.n1697 vdd.n1538 52.4337
R18244 vdd.n1695 vdd.n1694 52.4337
R18245 vdd.n1547 vdd.n1546 52.4337
R18246 vdd.n1686 vdd.n1551 52.4337
R18247 vdd.n1684 vdd.n1683 52.4337
R18248 vdd.n1679 vdd.n1557 52.4337
R18249 vdd.n1677 vdd.n1676 52.4337
R18250 vdd.n1672 vdd.n1564 52.4337
R18251 vdd.n1670 vdd.n1669 52.4337
R18252 vdd.n1665 vdd.n1571 52.4337
R18253 vdd.n1663 vdd.n1662 52.4337
R18254 vdd.n1658 vdd.n1578 52.4337
R18255 vdd.n1656 vdd.n1655 52.4337
R18256 vdd.n1587 vdd.n1586 52.4337
R18257 vdd.n1647 vdd.n1591 52.4337
R18258 vdd.n1645 vdd.n1644 52.4337
R18259 vdd.n1640 vdd.n1597 52.4337
R18260 vdd.n1638 vdd.n1637 52.4337
R18261 vdd.n1633 vdd.n1604 52.4337
R18262 vdd.n1631 vdd.n1630 52.4337
R18263 vdd.n1626 vdd.n1612 52.4337
R18264 vdd.n1624 vdd.n1623 52.4337
R18265 vdd.n1619 vdd.n1618 52.4337
R18266 vdd.n1614 vdd.n1613 52.4337
R18267 vdd.n1945 vdd.n860 52.4337
R18268 vdd.n1423 vdd.n1422 52.4337
R18269 vdd.n1229 vdd.n1197 52.4337
R18270 vdd.n1233 vdd.n1198 52.4337
R18271 vdd.n1235 vdd.n1199 52.4337
R18272 vdd.n1239 vdd.n1200 52.4337
R18273 vdd.n1241 vdd.n1201 52.4337
R18274 vdd.n1245 vdd.n1202 52.4337
R18275 vdd.n1247 vdd.n1203 52.4337
R18276 vdd.n1251 vdd.n1204 52.4337
R18277 vdd.n1253 vdd.n1205 52.4337
R18278 vdd.n1259 vdd.n1206 52.4337
R18279 vdd.n1261 vdd.n1207 52.4337
R18280 vdd.n1265 vdd.n1208 52.4337
R18281 vdd.n1267 vdd.n1209 52.4337
R18282 vdd.n1271 vdd.n1210 52.4337
R18283 vdd.n1273 vdd.n1211 52.4337
R18284 vdd.n1277 vdd.n1212 52.4337
R18285 vdd.n1279 vdd.n1213 52.4337
R18286 vdd.n1283 vdd.n1214 52.4337
R18287 vdd.n1285 vdd.n1215 52.4337
R18288 vdd.n1357 vdd.n1216 52.4337
R18289 vdd.n1290 vdd.n1217 52.4337
R18290 vdd.n1294 vdd.n1218 52.4337
R18291 vdd.n1296 vdd.n1219 52.4337
R18292 vdd.n1300 vdd.n1220 52.4337
R18293 vdd.n1302 vdd.n1221 52.4337
R18294 vdd.n1306 vdd.n1222 52.4337
R18295 vdd.n1308 vdd.n1223 52.4337
R18296 vdd.n1312 vdd.n1224 52.4337
R18297 vdd.n1314 vdd.n1225 52.4337
R18298 vdd.n1318 vdd.n1226 52.4337
R18299 vdd.n1422 vdd.n1196 52.4337
R18300 vdd.n1232 vdd.n1197 52.4337
R18301 vdd.n1234 vdd.n1198 52.4337
R18302 vdd.n1238 vdd.n1199 52.4337
R18303 vdd.n1240 vdd.n1200 52.4337
R18304 vdd.n1244 vdd.n1201 52.4337
R18305 vdd.n1246 vdd.n1202 52.4337
R18306 vdd.n1250 vdd.n1203 52.4337
R18307 vdd.n1252 vdd.n1204 52.4337
R18308 vdd.n1258 vdd.n1205 52.4337
R18309 vdd.n1260 vdd.n1206 52.4337
R18310 vdd.n1264 vdd.n1207 52.4337
R18311 vdd.n1266 vdd.n1208 52.4337
R18312 vdd.n1270 vdd.n1209 52.4337
R18313 vdd.n1272 vdd.n1210 52.4337
R18314 vdd.n1276 vdd.n1211 52.4337
R18315 vdd.n1278 vdd.n1212 52.4337
R18316 vdd.n1282 vdd.n1213 52.4337
R18317 vdd.n1284 vdd.n1214 52.4337
R18318 vdd.n1288 vdd.n1215 52.4337
R18319 vdd.n1289 vdd.n1216 52.4337
R18320 vdd.n1293 vdd.n1217 52.4337
R18321 vdd.n1295 vdd.n1218 52.4337
R18322 vdd.n1299 vdd.n1219 52.4337
R18323 vdd.n1301 vdd.n1220 52.4337
R18324 vdd.n1305 vdd.n1221 52.4337
R18325 vdd.n1307 vdd.n1222 52.4337
R18326 vdd.n1311 vdd.n1223 52.4337
R18327 vdd.n1313 vdd.n1224 52.4337
R18328 vdd.n1317 vdd.n1225 52.4337
R18329 vdd.n1319 vdd.n1226 52.4337
R18330 vdd.n860 vdd.n859 52.4337
R18331 vdd.n1615 vdd.n1614 52.4337
R18332 vdd.n1620 vdd.n1619 52.4337
R18333 vdd.n1625 vdd.n1624 52.4337
R18334 vdd.n1612 vdd.n1605 52.4337
R18335 vdd.n1632 vdd.n1631 52.4337
R18336 vdd.n1604 vdd.n1598 52.4337
R18337 vdd.n1639 vdd.n1638 52.4337
R18338 vdd.n1597 vdd.n1592 52.4337
R18339 vdd.n1646 vdd.n1645 52.4337
R18340 vdd.n1591 vdd.n1590 52.4337
R18341 vdd.n1586 vdd.n1579 52.4337
R18342 vdd.n1657 vdd.n1656 52.4337
R18343 vdd.n1578 vdd.n1572 52.4337
R18344 vdd.n1664 vdd.n1663 52.4337
R18345 vdd.n1571 vdd.n1565 52.4337
R18346 vdd.n1671 vdd.n1670 52.4337
R18347 vdd.n1564 vdd.n1558 52.4337
R18348 vdd.n1678 vdd.n1677 52.4337
R18349 vdd.n1557 vdd.n1552 52.4337
R18350 vdd.n1685 vdd.n1684 52.4337
R18351 vdd.n1551 vdd.n1550 52.4337
R18352 vdd.n1546 vdd.n1539 52.4337
R18353 vdd.n1696 vdd.n1695 52.4337
R18354 vdd.n1538 vdd.n1532 52.4337
R18355 vdd.n1703 vdd.n1702 52.4337
R18356 vdd.n1531 vdd.n1525 52.4337
R18357 vdd.n1710 vdd.n1709 52.4337
R18358 vdd.n1713 vdd.n1712 52.4337
R18359 vdd.n1522 vdd.n1517 52.4337
R18360 vdd.n1935 vdd.n1934 52.4337
R18361 vdd.n1516 vdd.n865 52.4337
R18362 vdd.n2841 vdd.n483 52.4337
R18363 vdd.n522 vdd.n485 52.4337
R18364 vdd.n2832 vdd.n486 52.4337
R18365 vdd.n2828 vdd.n487 52.4337
R18366 vdd.n2824 vdd.n488 52.4337
R18367 vdd.n2820 vdd.n489 52.4337
R18368 vdd.n2816 vdd.n490 52.4337
R18369 vdd.n2812 vdd.n491 52.4337
R18370 vdd.n2808 vdd.n492 52.4337
R18371 vdd.n2798 vdd.n493 52.4337
R18372 vdd.n2796 vdd.n494 52.4337
R18373 vdd.n2792 vdd.n495 52.4337
R18374 vdd.n2788 vdd.n496 52.4337
R18375 vdd.n2784 vdd.n497 52.4337
R18376 vdd.n2780 vdd.n498 52.4337
R18377 vdd.n2776 vdd.n499 52.4337
R18378 vdd.n2772 vdd.n500 52.4337
R18379 vdd.n2768 vdd.n501 52.4337
R18380 vdd.n2764 vdd.n502 52.4337
R18381 vdd.n2760 vdd.n503 52.4337
R18382 vdd.n2752 vdd.n504 52.4337
R18383 vdd.n2750 vdd.n505 52.4337
R18384 vdd.n2746 vdd.n506 52.4337
R18385 vdd.n2742 vdd.n507 52.4337
R18386 vdd.n2738 vdd.n508 52.4337
R18387 vdd.n2734 vdd.n509 52.4337
R18388 vdd.n2730 vdd.n510 52.4337
R18389 vdd.n2726 vdd.n511 52.4337
R18390 vdd.n2722 vdd.n512 52.4337
R18391 vdd.n2718 vdd.n513 52.4337
R18392 vdd.n2714 vdd.n514 52.4337
R18393 vdd.n2905 vdd.n440 52.4337
R18394 vdd.n2915 vdd.n2914 52.4337
R18395 vdd.n439 vdd.n433 52.4337
R18396 vdd.n2922 vdd.n2921 52.4337
R18397 vdd.n432 vdd.n426 52.4337
R18398 vdd.n2929 vdd.n2928 52.4337
R18399 vdd.n425 vdd.n419 52.4337
R18400 vdd.n2936 vdd.n2935 52.4337
R18401 vdd.n418 vdd.n413 52.4337
R18402 vdd.n2943 vdd.n2942 52.4337
R18403 vdd.n412 vdd.n411 52.4337
R18404 vdd.n407 vdd.n400 52.4337
R18405 vdd.n2954 vdd.n2953 52.4337
R18406 vdd.n399 vdd.n393 52.4337
R18407 vdd.n2961 vdd.n2960 52.4337
R18408 vdd.n392 vdd.n386 52.4337
R18409 vdd.n2968 vdd.n2967 52.4337
R18410 vdd.n385 vdd.n379 52.4337
R18411 vdd.n2975 vdd.n2974 52.4337
R18412 vdd.n378 vdd.n373 52.4337
R18413 vdd.n2982 vdd.n2981 52.4337
R18414 vdd.n372 vdd.n371 52.4337
R18415 vdd.n367 vdd.n360 52.4337
R18416 vdd.n2993 vdd.n2992 52.4337
R18417 vdd.n359 vdd.n353 52.4337
R18418 vdd.n3000 vdd.n2999 52.4337
R18419 vdd.n352 vdd.n346 52.4337
R18420 vdd.n3007 vdd.n3006 52.4337
R18421 vdd.n345 vdd.n338 52.4337
R18422 vdd.n3014 vdd.n3013 52.4337
R18423 vdd.n3017 vdd.n3016 52.4337
R18424 vdd.n333 vdd.n330 52.4337
R18425 vdd.t147 vdd.t141 51.4683
R18426 vdd.n250 vdd.n248 42.0461
R18427 vdd.n160 vdd.n158 42.0461
R18428 vdd.n71 vdd.n69 42.0461
R18429 vdd.n1112 vdd.n1110 42.0461
R18430 vdd.n1022 vdd.n1020 42.0461
R18431 vdd.n933 vdd.n931 42.0461
R18432 vdd.n296 vdd.n295 41.6884
R18433 vdd.n206 vdd.n205 41.6884
R18434 vdd.n117 vdd.n116 41.6884
R18435 vdd.n1158 vdd.n1157 41.6884
R18436 vdd.n1068 vdd.n1067 41.6884
R18437 vdd.n979 vdd.n978 41.6884
R18438 vdd.n1322 vdd.n1321 41.1157
R18439 vdd.n1360 vdd.n1359 41.1157
R18440 vdd.n1256 vdd.n1255 41.1157
R18441 vdd.n2910 vdd.n2909 41.1157
R18442 vdd.n2949 vdd.n406 41.1157
R18443 vdd.n2988 vdd.n366 41.1157
R18444 vdd.n2667 vdd.n2666 39.2114
R18445 vdd.n2664 vdd.n2663 39.2114
R18446 vdd.n2659 vdd.n605 39.2114
R18447 vdd.n2657 vdd.n2656 39.2114
R18448 vdd.n2652 vdd.n608 39.2114
R18449 vdd.n2650 vdd.n2649 39.2114
R18450 vdd.n2645 vdd.n611 39.2114
R18451 vdd.n2643 vdd.n2642 39.2114
R18452 vdd.n2639 vdd.n2638 39.2114
R18453 vdd.n2634 vdd.n614 39.2114
R18454 vdd.n2632 vdd.n2631 39.2114
R18455 vdd.n2627 vdd.n617 39.2114
R18456 vdd.n2625 vdd.n2624 39.2114
R18457 vdd.n2620 vdd.n620 39.2114
R18458 vdd.n2618 vdd.n2617 39.2114
R18459 vdd.n2612 vdd.n625 39.2114
R18460 vdd.n2610 vdd.n2609 39.2114
R18461 vdd.n2470 vdd.n703 39.2114
R18462 vdd.n2465 vdd.n2219 39.2114
R18463 vdd.n2462 vdd.n2220 39.2114
R18464 vdd.n2458 vdd.n2221 39.2114
R18465 vdd.n2454 vdd.n2222 39.2114
R18466 vdd.n2450 vdd.n2223 39.2114
R18467 vdd.n2446 vdd.n2224 39.2114
R18468 vdd.n2442 vdd.n2225 39.2114
R18469 vdd.n2438 vdd.n2226 39.2114
R18470 vdd.n2434 vdd.n2227 39.2114
R18471 vdd.n2430 vdd.n2228 39.2114
R18472 vdd.n2426 vdd.n2229 39.2114
R18473 vdd.n2422 vdd.n2230 39.2114
R18474 vdd.n2418 vdd.n2231 39.2114
R18475 vdd.n2414 vdd.n2232 39.2114
R18476 vdd.n2410 vdd.n2233 39.2114
R18477 vdd.n2405 vdd.n2234 39.2114
R18478 vdd.n2213 vdd.n743 39.2114
R18479 vdd.n2209 vdd.n742 39.2114
R18480 vdd.n2205 vdd.n741 39.2114
R18481 vdd.n2201 vdd.n740 39.2114
R18482 vdd.n2197 vdd.n739 39.2114
R18483 vdd.n2193 vdd.n738 39.2114
R18484 vdd.n2189 vdd.n737 39.2114
R18485 vdd.n2185 vdd.n736 39.2114
R18486 vdd.n2181 vdd.n735 39.2114
R18487 vdd.n2177 vdd.n734 39.2114
R18488 vdd.n2173 vdd.n733 39.2114
R18489 vdd.n2169 vdd.n732 39.2114
R18490 vdd.n2165 vdd.n731 39.2114
R18491 vdd.n2161 vdd.n730 39.2114
R18492 vdd.n2157 vdd.n729 39.2114
R18493 vdd.n2152 vdd.n728 39.2114
R18494 vdd.n2148 vdd.n727 39.2114
R18495 vdd.n1724 vdd.n838 39.2114
R18496 vdd.n1730 vdd.n1729 39.2114
R18497 vdd.n1733 vdd.n1732 39.2114
R18498 vdd.n1738 vdd.n1737 39.2114
R18499 vdd.n1741 vdd.n1740 39.2114
R18500 vdd.n1746 vdd.n1745 39.2114
R18501 vdd.n1749 vdd.n1748 39.2114
R18502 vdd.n1754 vdd.n1753 39.2114
R18503 vdd.n1925 vdd.n1756 39.2114
R18504 vdd.n1924 vdd.n1923 39.2114
R18505 vdd.n1917 vdd.n1758 39.2114
R18506 vdd.n1916 vdd.n1915 39.2114
R18507 vdd.n1909 vdd.n1760 39.2114
R18508 vdd.n1908 vdd.n1907 39.2114
R18509 vdd.n1901 vdd.n1762 39.2114
R18510 vdd.n1900 vdd.n1899 39.2114
R18511 vdd.n1893 vdd.n1764 39.2114
R18512 vdd.n2586 vdd.n2585 39.2114
R18513 vdd.n2581 vdd.n2553 39.2114
R18514 vdd.n2579 vdd.n2578 39.2114
R18515 vdd.n2574 vdd.n2556 39.2114
R18516 vdd.n2572 vdd.n2571 39.2114
R18517 vdd.n2567 vdd.n2559 39.2114
R18518 vdd.n2565 vdd.n2564 39.2114
R18519 vdd.n2560 vdd.n577 39.2114
R18520 vdd.n2704 vdd.n2703 39.2114
R18521 vdd.n2701 vdd.n2700 39.2114
R18522 vdd.n2696 vdd.n581 39.2114
R18523 vdd.n2694 vdd.n2693 39.2114
R18524 vdd.n2689 vdd.n584 39.2114
R18525 vdd.n2687 vdd.n2686 39.2114
R18526 vdd.n2682 vdd.n587 39.2114
R18527 vdd.n2680 vdd.n2679 39.2114
R18528 vdd.n2675 vdd.n593 39.2114
R18529 vdd.n2472 vdd.n706 39.2114
R18530 vdd.n2235 vdd.n708 39.2114
R18531 vdd.n2261 vdd.n2236 39.2114
R18532 vdd.n2265 vdd.n2237 39.2114
R18533 vdd.n2269 vdd.n2238 39.2114
R18534 vdd.n2273 vdd.n2239 39.2114
R18535 vdd.n2277 vdd.n2240 39.2114
R18536 vdd.n2281 vdd.n2241 39.2114
R18537 vdd.n2285 vdd.n2242 39.2114
R18538 vdd.n2289 vdd.n2243 39.2114
R18539 vdd.n2293 vdd.n2244 39.2114
R18540 vdd.n2297 vdd.n2245 39.2114
R18541 vdd.n2301 vdd.n2246 39.2114
R18542 vdd.n2305 vdd.n2247 39.2114
R18543 vdd.n2309 vdd.n2248 39.2114
R18544 vdd.n2313 vdd.n2249 39.2114
R18545 vdd.n2317 vdd.n2250 39.2114
R18546 vdd.n2473 vdd.n2472 39.2114
R18547 vdd.n2260 vdd.n2235 39.2114
R18548 vdd.n2264 vdd.n2236 39.2114
R18549 vdd.n2268 vdd.n2237 39.2114
R18550 vdd.n2272 vdd.n2238 39.2114
R18551 vdd.n2276 vdd.n2239 39.2114
R18552 vdd.n2280 vdd.n2240 39.2114
R18553 vdd.n2284 vdd.n2241 39.2114
R18554 vdd.n2288 vdd.n2242 39.2114
R18555 vdd.n2292 vdd.n2243 39.2114
R18556 vdd.n2296 vdd.n2244 39.2114
R18557 vdd.n2300 vdd.n2245 39.2114
R18558 vdd.n2304 vdd.n2246 39.2114
R18559 vdd.n2308 vdd.n2247 39.2114
R18560 vdd.n2312 vdd.n2248 39.2114
R18561 vdd.n2316 vdd.n2249 39.2114
R18562 vdd.n2319 vdd.n2250 39.2114
R18563 vdd.n593 vdd.n588 39.2114
R18564 vdd.n2681 vdd.n2680 39.2114
R18565 vdd.n587 vdd.n585 39.2114
R18566 vdd.n2688 vdd.n2687 39.2114
R18567 vdd.n584 vdd.n582 39.2114
R18568 vdd.n2695 vdd.n2694 39.2114
R18569 vdd.n581 vdd.n579 39.2114
R18570 vdd.n2702 vdd.n2701 39.2114
R18571 vdd.n2705 vdd.n2704 39.2114
R18572 vdd.n2561 vdd.n2560 39.2114
R18573 vdd.n2566 vdd.n2565 39.2114
R18574 vdd.n2559 vdd.n2557 39.2114
R18575 vdd.n2573 vdd.n2572 39.2114
R18576 vdd.n2556 vdd.n2554 39.2114
R18577 vdd.n2580 vdd.n2579 39.2114
R18578 vdd.n2553 vdd.n2551 39.2114
R18579 vdd.n2587 vdd.n2586 39.2114
R18580 vdd.n1725 vdd.n1724 39.2114
R18581 vdd.n1731 vdd.n1730 39.2114
R18582 vdd.n1732 vdd.n1721 39.2114
R18583 vdd.n1739 vdd.n1738 39.2114
R18584 vdd.n1740 vdd.n1719 39.2114
R18585 vdd.n1747 vdd.n1746 39.2114
R18586 vdd.n1748 vdd.n1717 39.2114
R18587 vdd.n1755 vdd.n1754 39.2114
R18588 vdd.n1926 vdd.n1925 39.2114
R18589 vdd.n1923 vdd.n1922 39.2114
R18590 vdd.n1918 vdd.n1917 39.2114
R18591 vdd.n1915 vdd.n1914 39.2114
R18592 vdd.n1910 vdd.n1909 39.2114
R18593 vdd.n1907 vdd.n1906 39.2114
R18594 vdd.n1902 vdd.n1901 39.2114
R18595 vdd.n1899 vdd.n1898 39.2114
R18596 vdd.n1894 vdd.n1893 39.2114
R18597 vdd.n2151 vdd.n727 39.2114
R18598 vdd.n2156 vdd.n728 39.2114
R18599 vdd.n2160 vdd.n729 39.2114
R18600 vdd.n2164 vdd.n730 39.2114
R18601 vdd.n2168 vdd.n731 39.2114
R18602 vdd.n2172 vdd.n732 39.2114
R18603 vdd.n2176 vdd.n733 39.2114
R18604 vdd.n2180 vdd.n734 39.2114
R18605 vdd.n2184 vdd.n735 39.2114
R18606 vdd.n2188 vdd.n736 39.2114
R18607 vdd.n2192 vdd.n737 39.2114
R18608 vdd.n2196 vdd.n738 39.2114
R18609 vdd.n2200 vdd.n739 39.2114
R18610 vdd.n2204 vdd.n740 39.2114
R18611 vdd.n2208 vdd.n741 39.2114
R18612 vdd.n2212 vdd.n742 39.2114
R18613 vdd.n745 vdd.n743 39.2114
R18614 vdd.n2470 vdd.n2469 39.2114
R18615 vdd.n2463 vdd.n2219 39.2114
R18616 vdd.n2459 vdd.n2220 39.2114
R18617 vdd.n2455 vdd.n2221 39.2114
R18618 vdd.n2451 vdd.n2222 39.2114
R18619 vdd.n2447 vdd.n2223 39.2114
R18620 vdd.n2443 vdd.n2224 39.2114
R18621 vdd.n2439 vdd.n2225 39.2114
R18622 vdd.n2435 vdd.n2226 39.2114
R18623 vdd.n2431 vdd.n2227 39.2114
R18624 vdd.n2427 vdd.n2228 39.2114
R18625 vdd.n2423 vdd.n2229 39.2114
R18626 vdd.n2419 vdd.n2230 39.2114
R18627 vdd.n2415 vdd.n2231 39.2114
R18628 vdd.n2411 vdd.n2232 39.2114
R18629 vdd.n2406 vdd.n2233 39.2114
R18630 vdd.n2402 vdd.n2234 39.2114
R18631 vdd.n2611 vdd.n2610 39.2114
R18632 vdd.n625 vdd.n621 39.2114
R18633 vdd.n2619 vdd.n2618 39.2114
R18634 vdd.n620 vdd.n618 39.2114
R18635 vdd.n2626 vdd.n2625 39.2114
R18636 vdd.n617 vdd.n615 39.2114
R18637 vdd.n2633 vdd.n2632 39.2114
R18638 vdd.n614 vdd.n612 39.2114
R18639 vdd.n2640 vdd.n2639 39.2114
R18640 vdd.n2644 vdd.n2643 39.2114
R18641 vdd.n611 vdd.n609 39.2114
R18642 vdd.n2651 vdd.n2650 39.2114
R18643 vdd.n608 vdd.n606 39.2114
R18644 vdd.n2658 vdd.n2657 39.2114
R18645 vdd.n605 vdd.n603 39.2114
R18646 vdd.n2665 vdd.n2664 39.2114
R18647 vdd.n2668 vdd.n2667 39.2114
R18648 vdd.n753 vdd.n709 39.2114
R18649 vdd.n2140 vdd.n710 39.2114
R18650 vdd.n2136 vdd.n711 39.2114
R18651 vdd.n2132 vdd.n712 39.2114
R18652 vdd.n2128 vdd.n713 39.2114
R18653 vdd.n2124 vdd.n714 39.2114
R18654 vdd.n2120 vdd.n715 39.2114
R18655 vdd.n2116 vdd.n716 39.2114
R18656 vdd.n2112 vdd.n717 39.2114
R18657 vdd.n2108 vdd.n718 39.2114
R18658 vdd.n2104 vdd.n719 39.2114
R18659 vdd.n2100 vdd.n720 39.2114
R18660 vdd.n2096 vdd.n721 39.2114
R18661 vdd.n2092 vdd.n722 39.2114
R18662 vdd.n2088 vdd.n723 39.2114
R18663 vdd.n2084 vdd.n724 39.2114
R18664 vdd.n2080 vdd.n725 39.2114
R18665 vdd.n1983 vdd.n842 39.2114
R18666 vdd.n1982 vdd.n1981 39.2114
R18667 vdd.n1975 vdd.n844 39.2114
R18668 vdd.n1974 vdd.n1973 39.2114
R18669 vdd.n1967 vdd.n846 39.2114
R18670 vdd.n1966 vdd.n1965 39.2114
R18671 vdd.n1959 vdd.n848 39.2114
R18672 vdd.n1958 vdd.n1957 39.2114
R18673 vdd.n851 vdd.n850 39.2114
R18674 vdd.n1799 vdd.n1798 39.2114
R18675 vdd.n1804 vdd.n1803 39.2114
R18676 vdd.n1807 vdd.n1806 39.2114
R18677 vdd.n1812 vdd.n1811 39.2114
R18678 vdd.n1815 vdd.n1814 39.2114
R18679 vdd.n1820 vdd.n1819 39.2114
R18680 vdd.n1823 vdd.n1822 39.2114
R18681 vdd.n1829 vdd.n1828 39.2114
R18682 vdd.n2077 vdd.n725 39.2114
R18683 vdd.n2081 vdd.n724 39.2114
R18684 vdd.n2085 vdd.n723 39.2114
R18685 vdd.n2089 vdd.n722 39.2114
R18686 vdd.n2093 vdd.n721 39.2114
R18687 vdd.n2097 vdd.n720 39.2114
R18688 vdd.n2101 vdd.n719 39.2114
R18689 vdd.n2105 vdd.n718 39.2114
R18690 vdd.n2109 vdd.n717 39.2114
R18691 vdd.n2113 vdd.n716 39.2114
R18692 vdd.n2117 vdd.n715 39.2114
R18693 vdd.n2121 vdd.n714 39.2114
R18694 vdd.n2125 vdd.n713 39.2114
R18695 vdd.n2129 vdd.n712 39.2114
R18696 vdd.n2133 vdd.n711 39.2114
R18697 vdd.n2137 vdd.n710 39.2114
R18698 vdd.n2141 vdd.n709 39.2114
R18699 vdd.n1984 vdd.n1983 39.2114
R18700 vdd.n1981 vdd.n1980 39.2114
R18701 vdd.n1976 vdd.n1975 39.2114
R18702 vdd.n1973 vdd.n1972 39.2114
R18703 vdd.n1968 vdd.n1967 39.2114
R18704 vdd.n1965 vdd.n1964 39.2114
R18705 vdd.n1960 vdd.n1959 39.2114
R18706 vdd.n1957 vdd.n1956 39.2114
R18707 vdd.n852 vdd.n851 39.2114
R18708 vdd.n1800 vdd.n1799 39.2114
R18709 vdd.n1805 vdd.n1804 39.2114
R18710 vdd.n1806 vdd.n1796 39.2114
R18711 vdd.n1813 vdd.n1812 39.2114
R18712 vdd.n1814 vdd.n1794 39.2114
R18713 vdd.n1821 vdd.n1820 39.2114
R18714 vdd.n1822 vdd.n1790 39.2114
R18715 vdd.n1830 vdd.n1829 39.2114
R18716 vdd.n1949 vdd.n1948 37.2369
R18717 vdd.n1652 vdd.n1585 37.2369
R18718 vdd.n1691 vdd.n1545 37.2369
R18719 vdd.n2758 vdd.n558 37.2369
R18720 vdd.n2806 vdd.n2805 37.2369
R18721 vdd.n2713 vdd.n2712 37.2369
R18722 vdd.n1991 vdd.n837 31.6883
R18723 vdd.n2216 vdd.n746 31.6883
R18724 vdd.n2149 vdd.n749 31.6883
R18725 vdd.n1895 vdd.n1892 31.6883
R18726 vdd.n2403 vdd.n2401 31.6883
R18727 vdd.n2608 vdd.n2607 31.6883
R18728 vdd.n2480 vdd.n702 31.6883
R18729 vdd.n2671 vdd.n2670 31.6883
R18730 vdd.n2590 vdd.n2589 31.6883
R18731 vdd.n2676 vdd.n592 31.6883
R18732 vdd.n2322 vdd.n2321 31.6883
R18733 vdd.n2476 vdd.n2475 31.6883
R18734 vdd.n1987 vdd.n1986 31.6883
R18735 vdd.n2144 vdd.n2143 31.6883
R18736 vdd.n2076 vdd.n2075 31.6883
R18737 vdd.n1833 vdd.n1832 31.6883
R18738 vdd.n1826 vdd.n1792 30.449
R18739 vdd.n757 vdd.n756 30.449
R18740 vdd.n1767 vdd.n1766 30.449
R18741 vdd.n2154 vdd.n748 30.449
R18742 vdd.n2258 vdd.n2257 30.449
R18743 vdd.n2614 vdd.n623 30.449
R18744 vdd.n2408 vdd.n2254 30.449
R18745 vdd.n591 vdd.n590 30.449
R18746 vdd.n1421 vdd.n1228 22.6735
R18747 vdd.n1943 vdd.n863 22.6735
R18748 vdd.n2840 vdd.n516 22.6735
R18749 vdd.n3025 vdd.n329 22.6735
R18750 vdd.n1432 vdd.n1190 19.3944
R18751 vdd.n1432 vdd.n1188 19.3944
R18752 vdd.n1436 vdd.n1188 19.3944
R18753 vdd.n1436 vdd.n1178 19.3944
R18754 vdd.n1449 vdd.n1178 19.3944
R18755 vdd.n1449 vdd.n1176 19.3944
R18756 vdd.n1453 vdd.n1176 19.3944
R18757 vdd.n1453 vdd.n1168 19.3944
R18758 vdd.n1467 vdd.n1168 19.3944
R18759 vdd.n1467 vdd.n1166 19.3944
R18760 vdd.n1471 vdd.n1166 19.3944
R18761 vdd.n1471 vdd.n885 19.3944
R18762 vdd.n1483 vdd.n885 19.3944
R18763 vdd.n1483 vdd.n883 19.3944
R18764 vdd.n1487 vdd.n883 19.3944
R18765 vdd.n1487 vdd.n875 19.3944
R18766 vdd.n1500 vdd.n875 19.3944
R18767 vdd.n1500 vdd.n872 19.3944
R18768 vdd.n1506 vdd.n872 19.3944
R18769 vdd.n1506 vdd.n873 19.3944
R18770 vdd.n873 vdd.n862 19.3944
R18771 vdd.n1356 vdd.n1291 19.3944
R18772 vdd.n1352 vdd.n1291 19.3944
R18773 vdd.n1352 vdd.n1351 19.3944
R18774 vdd.n1351 vdd.n1350 19.3944
R18775 vdd.n1350 vdd.n1297 19.3944
R18776 vdd.n1346 vdd.n1297 19.3944
R18777 vdd.n1346 vdd.n1345 19.3944
R18778 vdd.n1345 vdd.n1344 19.3944
R18779 vdd.n1344 vdd.n1303 19.3944
R18780 vdd.n1340 vdd.n1303 19.3944
R18781 vdd.n1340 vdd.n1339 19.3944
R18782 vdd.n1339 vdd.n1338 19.3944
R18783 vdd.n1338 vdd.n1309 19.3944
R18784 vdd.n1334 vdd.n1309 19.3944
R18785 vdd.n1334 vdd.n1333 19.3944
R18786 vdd.n1333 vdd.n1332 19.3944
R18787 vdd.n1332 vdd.n1315 19.3944
R18788 vdd.n1328 vdd.n1315 19.3944
R18789 vdd.n1328 vdd.n1327 19.3944
R18790 vdd.n1327 vdd.n1326 19.3944
R18791 vdd.n1391 vdd.n1390 19.3944
R18792 vdd.n1390 vdd.n1389 19.3944
R18793 vdd.n1389 vdd.n1262 19.3944
R18794 vdd.n1385 vdd.n1262 19.3944
R18795 vdd.n1385 vdd.n1384 19.3944
R18796 vdd.n1384 vdd.n1383 19.3944
R18797 vdd.n1383 vdd.n1268 19.3944
R18798 vdd.n1379 vdd.n1268 19.3944
R18799 vdd.n1379 vdd.n1378 19.3944
R18800 vdd.n1378 vdd.n1377 19.3944
R18801 vdd.n1377 vdd.n1274 19.3944
R18802 vdd.n1373 vdd.n1274 19.3944
R18803 vdd.n1373 vdd.n1372 19.3944
R18804 vdd.n1372 vdd.n1371 19.3944
R18805 vdd.n1371 vdd.n1280 19.3944
R18806 vdd.n1367 vdd.n1280 19.3944
R18807 vdd.n1367 vdd.n1366 19.3944
R18808 vdd.n1366 vdd.n1365 19.3944
R18809 vdd.n1365 vdd.n1286 19.3944
R18810 vdd.n1361 vdd.n1286 19.3944
R18811 vdd.n1424 vdd.n1195 19.3944
R18812 vdd.n1419 vdd.n1195 19.3944
R18813 vdd.n1419 vdd.n1230 19.3944
R18814 vdd.n1415 vdd.n1230 19.3944
R18815 vdd.n1415 vdd.n1414 19.3944
R18816 vdd.n1414 vdd.n1413 19.3944
R18817 vdd.n1413 vdd.n1236 19.3944
R18818 vdd.n1409 vdd.n1236 19.3944
R18819 vdd.n1409 vdd.n1408 19.3944
R18820 vdd.n1408 vdd.n1407 19.3944
R18821 vdd.n1407 vdd.n1242 19.3944
R18822 vdd.n1403 vdd.n1242 19.3944
R18823 vdd.n1403 vdd.n1402 19.3944
R18824 vdd.n1402 vdd.n1401 19.3944
R18825 vdd.n1401 vdd.n1248 19.3944
R18826 vdd.n1397 vdd.n1248 19.3944
R18827 vdd.n1397 vdd.n1396 19.3944
R18828 vdd.n1396 vdd.n1395 19.3944
R18829 vdd.n1648 vdd.n1583 19.3944
R18830 vdd.n1648 vdd.n1589 19.3944
R18831 vdd.n1643 vdd.n1589 19.3944
R18832 vdd.n1643 vdd.n1642 19.3944
R18833 vdd.n1642 vdd.n1641 19.3944
R18834 vdd.n1641 vdd.n1596 19.3944
R18835 vdd.n1636 vdd.n1596 19.3944
R18836 vdd.n1636 vdd.n1635 19.3944
R18837 vdd.n1635 vdd.n1634 19.3944
R18838 vdd.n1634 vdd.n1603 19.3944
R18839 vdd.n1629 vdd.n1603 19.3944
R18840 vdd.n1629 vdd.n1628 19.3944
R18841 vdd.n1628 vdd.n1627 19.3944
R18842 vdd.n1627 vdd.n1611 19.3944
R18843 vdd.n1622 vdd.n1611 19.3944
R18844 vdd.n1622 vdd.n1621 19.3944
R18845 vdd.n1617 vdd.n1616 19.3944
R18846 vdd.n1950 vdd.n858 19.3944
R18847 vdd.n1687 vdd.n1543 19.3944
R18848 vdd.n1687 vdd.n1549 19.3944
R18849 vdd.n1682 vdd.n1549 19.3944
R18850 vdd.n1682 vdd.n1681 19.3944
R18851 vdd.n1681 vdd.n1680 19.3944
R18852 vdd.n1680 vdd.n1556 19.3944
R18853 vdd.n1675 vdd.n1556 19.3944
R18854 vdd.n1675 vdd.n1674 19.3944
R18855 vdd.n1674 vdd.n1673 19.3944
R18856 vdd.n1673 vdd.n1563 19.3944
R18857 vdd.n1668 vdd.n1563 19.3944
R18858 vdd.n1668 vdd.n1667 19.3944
R18859 vdd.n1667 vdd.n1666 19.3944
R18860 vdd.n1666 vdd.n1570 19.3944
R18861 vdd.n1661 vdd.n1570 19.3944
R18862 vdd.n1661 vdd.n1660 19.3944
R18863 vdd.n1660 vdd.n1659 19.3944
R18864 vdd.n1659 vdd.n1577 19.3944
R18865 vdd.n1654 vdd.n1577 19.3944
R18866 vdd.n1654 vdd.n1653 19.3944
R18867 vdd.n1938 vdd.n1937 19.3944
R18868 vdd.n1937 vdd.n1515 19.3944
R18869 vdd.n1932 vdd.n1931 19.3944
R18870 vdd.n1714 vdd.n1519 19.3944
R18871 vdd.n1714 vdd.n1521 19.3944
R18872 vdd.n1524 vdd.n1521 19.3944
R18873 vdd.n1707 vdd.n1524 19.3944
R18874 vdd.n1707 vdd.n1706 19.3944
R18875 vdd.n1706 vdd.n1705 19.3944
R18876 vdd.n1705 vdd.n1530 19.3944
R18877 vdd.n1700 vdd.n1530 19.3944
R18878 vdd.n1700 vdd.n1699 19.3944
R18879 vdd.n1699 vdd.n1698 19.3944
R18880 vdd.n1698 vdd.n1537 19.3944
R18881 vdd.n1693 vdd.n1537 19.3944
R18882 vdd.n1693 vdd.n1692 19.3944
R18883 vdd.n1428 vdd.n1193 19.3944
R18884 vdd.n1428 vdd.n1184 19.3944
R18885 vdd.n1441 vdd.n1184 19.3944
R18886 vdd.n1441 vdd.n1182 19.3944
R18887 vdd.n1445 vdd.n1182 19.3944
R18888 vdd.n1445 vdd.n1173 19.3944
R18889 vdd.n1458 vdd.n1173 19.3944
R18890 vdd.n1458 vdd.n1171 19.3944
R18891 vdd.n1463 vdd.n1171 19.3944
R18892 vdd.n1463 vdd.n1162 19.3944
R18893 vdd.n1475 vdd.n1162 19.3944
R18894 vdd.n1475 vdd.n890 19.3944
R18895 vdd.n1479 vdd.n890 19.3944
R18896 vdd.n1479 vdd.n880 19.3944
R18897 vdd.n1492 vdd.n880 19.3944
R18898 vdd.n1492 vdd.n878 19.3944
R18899 vdd.n1496 vdd.n878 19.3944
R18900 vdd.n1496 vdd.n868 19.3944
R18901 vdd.n1511 vdd.n868 19.3944
R18902 vdd.n1511 vdd.n866 19.3944
R18903 vdd.n1941 vdd.n866 19.3944
R18904 vdd.n2851 vdd.n477 19.3944
R18905 vdd.n2851 vdd.n475 19.3944
R18906 vdd.n2855 vdd.n475 19.3944
R18907 vdd.n2855 vdd.n465 19.3944
R18908 vdd.n2868 vdd.n465 19.3944
R18909 vdd.n2868 vdd.n463 19.3944
R18910 vdd.n2872 vdd.n463 19.3944
R18911 vdd.n2872 vdd.n453 19.3944
R18912 vdd.n2884 vdd.n453 19.3944
R18913 vdd.n2884 vdd.n451 19.3944
R18914 vdd.n2888 vdd.n451 19.3944
R18915 vdd.n2889 vdd.n2888 19.3944
R18916 vdd.n2890 vdd.n2889 19.3944
R18917 vdd.n2890 vdd.n449 19.3944
R18918 vdd.n2894 vdd.n449 19.3944
R18919 vdd.n2895 vdd.n2894 19.3944
R18920 vdd.n2896 vdd.n2895 19.3944
R18921 vdd.n2896 vdd.n446 19.3944
R18922 vdd.n2900 vdd.n446 19.3944
R18923 vdd.n2901 vdd.n2900 19.3944
R18924 vdd.n2902 vdd.n2901 19.3944
R18925 vdd.n2945 vdd.n404 19.3944
R18926 vdd.n2945 vdd.n410 19.3944
R18927 vdd.n2940 vdd.n410 19.3944
R18928 vdd.n2940 vdd.n2939 19.3944
R18929 vdd.n2939 vdd.n2938 19.3944
R18930 vdd.n2938 vdd.n417 19.3944
R18931 vdd.n2933 vdd.n417 19.3944
R18932 vdd.n2933 vdd.n2932 19.3944
R18933 vdd.n2932 vdd.n2931 19.3944
R18934 vdd.n2931 vdd.n424 19.3944
R18935 vdd.n2926 vdd.n424 19.3944
R18936 vdd.n2926 vdd.n2925 19.3944
R18937 vdd.n2925 vdd.n2924 19.3944
R18938 vdd.n2924 vdd.n431 19.3944
R18939 vdd.n2919 vdd.n431 19.3944
R18940 vdd.n2919 vdd.n2918 19.3944
R18941 vdd.n2918 vdd.n2917 19.3944
R18942 vdd.n2917 vdd.n438 19.3944
R18943 vdd.n2912 vdd.n438 19.3944
R18944 vdd.n2912 vdd.n2911 19.3944
R18945 vdd.n2984 vdd.n364 19.3944
R18946 vdd.n2984 vdd.n370 19.3944
R18947 vdd.n2979 vdd.n370 19.3944
R18948 vdd.n2979 vdd.n2978 19.3944
R18949 vdd.n2978 vdd.n2977 19.3944
R18950 vdd.n2977 vdd.n377 19.3944
R18951 vdd.n2972 vdd.n377 19.3944
R18952 vdd.n2972 vdd.n2971 19.3944
R18953 vdd.n2971 vdd.n2970 19.3944
R18954 vdd.n2970 vdd.n384 19.3944
R18955 vdd.n2965 vdd.n384 19.3944
R18956 vdd.n2965 vdd.n2964 19.3944
R18957 vdd.n2964 vdd.n2963 19.3944
R18958 vdd.n2963 vdd.n391 19.3944
R18959 vdd.n2958 vdd.n391 19.3944
R18960 vdd.n2958 vdd.n2957 19.3944
R18961 vdd.n2957 vdd.n2956 19.3944
R18962 vdd.n2956 vdd.n398 19.3944
R18963 vdd.n2951 vdd.n398 19.3944
R18964 vdd.n2951 vdd.n2950 19.3944
R18965 vdd.n3020 vdd.n3019 19.3944
R18966 vdd.n3019 vdd.n3018 19.3944
R18967 vdd.n3018 vdd.n336 19.3944
R18968 vdd.n337 vdd.n336 19.3944
R18969 vdd.n3011 vdd.n337 19.3944
R18970 vdd.n3011 vdd.n3010 19.3944
R18971 vdd.n3010 vdd.n3009 19.3944
R18972 vdd.n3009 vdd.n344 19.3944
R18973 vdd.n3004 vdd.n344 19.3944
R18974 vdd.n3004 vdd.n3003 19.3944
R18975 vdd.n3003 vdd.n3002 19.3944
R18976 vdd.n3002 vdd.n351 19.3944
R18977 vdd.n2997 vdd.n351 19.3944
R18978 vdd.n2997 vdd.n2996 19.3944
R18979 vdd.n2996 vdd.n2995 19.3944
R18980 vdd.n2995 vdd.n358 19.3944
R18981 vdd.n2990 vdd.n358 19.3944
R18982 vdd.n2990 vdd.n2989 19.3944
R18983 vdd.n2847 vdd.n480 19.3944
R18984 vdd.n2847 vdd.n471 19.3944
R18985 vdd.n2860 vdd.n471 19.3944
R18986 vdd.n2860 vdd.n469 19.3944
R18987 vdd.n2864 vdd.n469 19.3944
R18988 vdd.n2864 vdd.n460 19.3944
R18989 vdd.n2876 vdd.n460 19.3944
R18990 vdd.n2876 vdd.n458 19.3944
R18991 vdd.n2880 vdd.n458 19.3944
R18992 vdd.n2880 vdd.n300 19.3944
R18993 vdd.n3045 vdd.n300 19.3944
R18994 vdd.n3045 vdd.n301 19.3944
R18995 vdd.n3039 vdd.n301 19.3944
R18996 vdd.n3039 vdd.n3038 19.3944
R18997 vdd.n3038 vdd.n3037 19.3944
R18998 vdd.n3037 vdd.n313 19.3944
R18999 vdd.n3031 vdd.n313 19.3944
R19000 vdd.n3031 vdd.n3030 19.3944
R19001 vdd.n3030 vdd.n3029 19.3944
R19002 vdd.n3029 vdd.n324 19.3944
R19003 vdd.n3023 vdd.n324 19.3944
R19004 vdd.n2800 vdd.n536 19.3944
R19005 vdd.n2800 vdd.n2797 19.3944
R19006 vdd.n2797 vdd.n2794 19.3944
R19007 vdd.n2794 vdd.n2793 19.3944
R19008 vdd.n2793 vdd.n2790 19.3944
R19009 vdd.n2790 vdd.n2789 19.3944
R19010 vdd.n2789 vdd.n2786 19.3944
R19011 vdd.n2786 vdd.n2785 19.3944
R19012 vdd.n2785 vdd.n2782 19.3944
R19013 vdd.n2782 vdd.n2781 19.3944
R19014 vdd.n2781 vdd.n2778 19.3944
R19015 vdd.n2778 vdd.n2777 19.3944
R19016 vdd.n2777 vdd.n2774 19.3944
R19017 vdd.n2774 vdd.n2773 19.3944
R19018 vdd.n2773 vdd.n2770 19.3944
R19019 vdd.n2770 vdd.n2769 19.3944
R19020 vdd.n2769 vdd.n2766 19.3944
R19021 vdd.n2766 vdd.n2765 19.3944
R19022 vdd.n2765 vdd.n2762 19.3944
R19023 vdd.n2762 vdd.n2761 19.3944
R19024 vdd.n2843 vdd.n482 19.3944
R19025 vdd.n2838 vdd.n482 19.3944
R19026 vdd.n521 vdd.n518 19.3944
R19027 vdd.n2834 vdd.n2833 19.3944
R19028 vdd.n2833 vdd.n2830 19.3944
R19029 vdd.n2830 vdd.n2829 19.3944
R19030 vdd.n2829 vdd.n2826 19.3944
R19031 vdd.n2826 vdd.n2825 19.3944
R19032 vdd.n2825 vdd.n2822 19.3944
R19033 vdd.n2822 vdd.n2821 19.3944
R19034 vdd.n2821 vdd.n2818 19.3944
R19035 vdd.n2818 vdd.n2817 19.3944
R19036 vdd.n2817 vdd.n2814 19.3944
R19037 vdd.n2814 vdd.n2813 19.3944
R19038 vdd.n2813 vdd.n2810 19.3944
R19039 vdd.n2810 vdd.n2809 19.3944
R19040 vdd.n2754 vdd.n556 19.3944
R19041 vdd.n2754 vdd.n2751 19.3944
R19042 vdd.n2751 vdd.n2748 19.3944
R19043 vdd.n2748 vdd.n2747 19.3944
R19044 vdd.n2747 vdd.n2744 19.3944
R19045 vdd.n2744 vdd.n2743 19.3944
R19046 vdd.n2743 vdd.n2740 19.3944
R19047 vdd.n2740 vdd.n2739 19.3944
R19048 vdd.n2739 vdd.n2736 19.3944
R19049 vdd.n2736 vdd.n2735 19.3944
R19050 vdd.n2735 vdd.n2732 19.3944
R19051 vdd.n2732 vdd.n2731 19.3944
R19052 vdd.n2731 vdd.n2728 19.3944
R19053 vdd.n2728 vdd.n2727 19.3944
R19054 vdd.n2727 vdd.n2724 19.3944
R19055 vdd.n2724 vdd.n2723 19.3944
R19056 vdd.n2720 vdd.n2719 19.3944
R19057 vdd.n2716 vdd.n2715 19.3944
R19058 vdd.n1360 vdd.n1356 19.0066
R19059 vdd.n1652 vdd.n1583 19.0066
R19060 vdd.n2949 vdd.n404 19.0066
R19061 vdd.n2758 vdd.n556 19.0066
R19062 vdd.n1792 vdd.n1791 16.0975
R19063 vdd.n756 vdd.n755 16.0975
R19064 vdd.n1321 vdd.n1320 16.0975
R19065 vdd.n1359 vdd.n1358 16.0975
R19066 vdd.n1255 vdd.n1254 16.0975
R19067 vdd.n1948 vdd.n1947 16.0975
R19068 vdd.n1585 vdd.n1584 16.0975
R19069 vdd.n1545 vdd.n1544 16.0975
R19070 vdd.n1766 vdd.n1765 16.0975
R19071 vdd.n748 vdd.n747 16.0975
R19072 vdd.n2257 vdd.n2256 16.0975
R19073 vdd.n2909 vdd.n2908 16.0975
R19074 vdd.n406 vdd.n405 16.0975
R19075 vdd.n366 vdd.n365 16.0975
R19076 vdd.n558 vdd.n557 16.0975
R19077 vdd.n2805 vdd.n2804 16.0975
R19078 vdd.n623 vdd.n622 16.0975
R19079 vdd.n2254 vdd.n2253 16.0975
R19080 vdd.n2712 vdd.n2711 16.0975
R19081 vdd.n590 vdd.n589 16.0975
R19082 vdd.t141 vdd.n2218 15.4182
R19083 vdd.n2471 vdd.t147 15.4182
R19084 vdd.n28 vdd.n27 14.5674
R19085 vdd.n1989 vdd.n839 14.5112
R19086 vdd.n2673 vdd.n484 14.5112
R19087 vdd.n292 vdd.n257 13.1884
R19088 vdd.n245 vdd.n210 13.1884
R19089 vdd.n202 vdd.n167 13.1884
R19090 vdd.n155 vdd.n120 13.1884
R19091 vdd.n113 vdd.n78 13.1884
R19092 vdd.n66 vdd.n31 13.1884
R19093 vdd.n1107 vdd.n1072 13.1884
R19094 vdd.n1154 vdd.n1119 13.1884
R19095 vdd.n1017 vdd.n982 13.1884
R19096 vdd.n1064 vdd.n1029 13.1884
R19097 vdd.n928 vdd.n893 13.1884
R19098 vdd.n975 vdd.n940 13.1884
R19099 vdd.n1391 vdd.n1256 12.9944
R19100 vdd.n1395 vdd.n1256 12.9944
R19101 vdd.n1691 vdd.n1543 12.9944
R19102 vdd.n1692 vdd.n1691 12.9944
R19103 vdd.n2988 vdd.n364 12.9944
R19104 vdd.n2989 vdd.n2988 12.9944
R19105 vdd.n2806 vdd.n536 12.9944
R19106 vdd.n2809 vdd.n2806 12.9944
R19107 vdd.n293 vdd.n255 12.8005
R19108 vdd.n288 vdd.n259 12.8005
R19109 vdd.n246 vdd.n208 12.8005
R19110 vdd.n241 vdd.n212 12.8005
R19111 vdd.n203 vdd.n165 12.8005
R19112 vdd.n198 vdd.n169 12.8005
R19113 vdd.n156 vdd.n118 12.8005
R19114 vdd.n151 vdd.n122 12.8005
R19115 vdd.n114 vdd.n76 12.8005
R19116 vdd.n109 vdd.n80 12.8005
R19117 vdd.n67 vdd.n29 12.8005
R19118 vdd.n62 vdd.n33 12.8005
R19119 vdd.n1108 vdd.n1070 12.8005
R19120 vdd.n1103 vdd.n1074 12.8005
R19121 vdd.n1155 vdd.n1117 12.8005
R19122 vdd.n1150 vdd.n1121 12.8005
R19123 vdd.n1018 vdd.n980 12.8005
R19124 vdd.n1013 vdd.n984 12.8005
R19125 vdd.n1065 vdd.n1027 12.8005
R19126 vdd.n1060 vdd.n1031 12.8005
R19127 vdd.n929 vdd.n891 12.8005
R19128 vdd.n924 vdd.n895 12.8005
R19129 vdd.n976 vdd.n938 12.8005
R19130 vdd.n971 vdd.n942 12.8005
R19131 vdd.n287 vdd.n260 12.0247
R19132 vdd.n240 vdd.n213 12.0247
R19133 vdd.n197 vdd.n170 12.0247
R19134 vdd.n150 vdd.n123 12.0247
R19135 vdd.n108 vdd.n81 12.0247
R19136 vdd.n61 vdd.n34 12.0247
R19137 vdd.n1102 vdd.n1075 12.0247
R19138 vdd.n1149 vdd.n1122 12.0247
R19139 vdd.n1012 vdd.n985 12.0247
R19140 vdd.n1059 vdd.n1032 12.0247
R19141 vdd.n923 vdd.n896 12.0247
R19142 vdd.n970 vdd.n943 12.0247
R19143 vdd.n1430 vdd.n1186 11.337
R19144 vdd.n1439 vdd.n1186 11.337
R19145 vdd.n1439 vdd.n1438 11.337
R19146 vdd.n1447 vdd.n1180 11.337
R19147 vdd.n1456 vdd.n1455 11.337
R19148 vdd.n1473 vdd.n1164 11.337
R19149 vdd.n1481 vdd.n887 11.337
R19150 vdd.n1490 vdd.n1489 11.337
R19151 vdd.n1498 vdd.n870 11.337
R19152 vdd.n1509 vdd.n870 11.337
R19153 vdd.n1509 vdd.n1508 11.337
R19154 vdd.n2849 vdd.n473 11.337
R19155 vdd.n2858 vdd.n473 11.337
R19156 vdd.n2858 vdd.n2857 11.337
R19157 vdd.n2866 vdd.n467 11.337
R19158 vdd.n2882 vdd.n456 11.337
R19159 vdd.n3043 vdd.n304 11.337
R19160 vdd.n3041 vdd.n308 11.337
R19161 vdd.n3035 vdd.n3034 11.337
R19162 vdd.n3033 vdd.n318 11.337
R19163 vdd.n3027 vdd.n318 11.337
R19164 vdd.n3027 vdd.n3026 11.337
R19165 vdd.n284 vdd.n283 11.249
R19166 vdd.n237 vdd.n236 11.249
R19167 vdd.n194 vdd.n193 11.249
R19168 vdd.n147 vdd.n146 11.249
R19169 vdd.n105 vdd.n104 11.249
R19170 vdd.n58 vdd.n57 11.249
R19171 vdd.n1099 vdd.n1098 11.249
R19172 vdd.n1146 vdd.n1145 11.249
R19173 vdd.n1009 vdd.n1008 11.249
R19174 vdd.n1056 vdd.n1055 11.249
R19175 vdd.n920 vdd.n919 11.249
R19176 vdd.n967 vdd.n966 11.249
R19177 vdd.n2146 vdd.t191 11.1103
R19178 vdd.n2478 vdd.t154 11.1103
R19179 vdd.n1228 vdd.t77 10.7702
R19180 vdd.t88 vdd.n3025 10.7702
R19181 vdd.n269 vdd.n268 10.7238
R19182 vdd.n222 vdd.n221 10.7238
R19183 vdd.n179 vdd.n178 10.7238
R19184 vdd.n132 vdd.n131 10.7238
R19185 vdd.n90 vdd.n89 10.7238
R19186 vdd.n43 vdd.n42 10.7238
R19187 vdd.n1084 vdd.n1083 10.7238
R19188 vdd.n1131 vdd.n1130 10.7238
R19189 vdd.n994 vdd.n993 10.7238
R19190 vdd.n1041 vdd.n1040 10.7238
R19191 vdd.n905 vdd.n904 10.7238
R19192 vdd.n952 vdd.n951 10.7238
R19193 vdd.n1992 vdd.n1991 10.6151
R19194 vdd.n1993 vdd.n1992 10.6151
R19195 vdd.n1993 vdd.n825 10.6151
R19196 vdd.n2003 vdd.n825 10.6151
R19197 vdd.n2004 vdd.n2003 10.6151
R19198 vdd.n2005 vdd.n2004 10.6151
R19199 vdd.n2005 vdd.n812 10.6151
R19200 vdd.n2016 vdd.n812 10.6151
R19201 vdd.n2017 vdd.n2016 10.6151
R19202 vdd.n2018 vdd.n2017 10.6151
R19203 vdd.n2018 vdd.n800 10.6151
R19204 vdd.n2028 vdd.n800 10.6151
R19205 vdd.n2029 vdd.n2028 10.6151
R19206 vdd.n2030 vdd.n2029 10.6151
R19207 vdd.n2030 vdd.n788 10.6151
R19208 vdd.n2040 vdd.n788 10.6151
R19209 vdd.n2041 vdd.n2040 10.6151
R19210 vdd.n2042 vdd.n2041 10.6151
R19211 vdd.n2042 vdd.n777 10.6151
R19212 vdd.n2052 vdd.n777 10.6151
R19213 vdd.n2053 vdd.n2052 10.6151
R19214 vdd.n2054 vdd.n2053 10.6151
R19215 vdd.n2054 vdd.n764 10.6151
R19216 vdd.n2066 vdd.n764 10.6151
R19217 vdd.n2067 vdd.n2066 10.6151
R19218 vdd.n2069 vdd.n2067 10.6151
R19219 vdd.n2069 vdd.n2068 10.6151
R19220 vdd.n2068 vdd.n746 10.6151
R19221 vdd.n2216 vdd.n2215 10.6151
R19222 vdd.n2215 vdd.n2214 10.6151
R19223 vdd.n2214 vdd.n2211 10.6151
R19224 vdd.n2211 vdd.n2210 10.6151
R19225 vdd.n2210 vdd.n2207 10.6151
R19226 vdd.n2207 vdd.n2206 10.6151
R19227 vdd.n2206 vdd.n2203 10.6151
R19228 vdd.n2203 vdd.n2202 10.6151
R19229 vdd.n2202 vdd.n2199 10.6151
R19230 vdd.n2199 vdd.n2198 10.6151
R19231 vdd.n2198 vdd.n2195 10.6151
R19232 vdd.n2195 vdd.n2194 10.6151
R19233 vdd.n2194 vdd.n2191 10.6151
R19234 vdd.n2191 vdd.n2190 10.6151
R19235 vdd.n2190 vdd.n2187 10.6151
R19236 vdd.n2187 vdd.n2186 10.6151
R19237 vdd.n2186 vdd.n2183 10.6151
R19238 vdd.n2183 vdd.n2182 10.6151
R19239 vdd.n2182 vdd.n2179 10.6151
R19240 vdd.n2179 vdd.n2178 10.6151
R19241 vdd.n2178 vdd.n2175 10.6151
R19242 vdd.n2175 vdd.n2174 10.6151
R19243 vdd.n2174 vdd.n2171 10.6151
R19244 vdd.n2171 vdd.n2170 10.6151
R19245 vdd.n2170 vdd.n2167 10.6151
R19246 vdd.n2167 vdd.n2166 10.6151
R19247 vdd.n2166 vdd.n2163 10.6151
R19248 vdd.n2163 vdd.n2162 10.6151
R19249 vdd.n2162 vdd.n2159 10.6151
R19250 vdd.n2159 vdd.n2158 10.6151
R19251 vdd.n2158 vdd.n2155 10.6151
R19252 vdd.n2153 vdd.n2150 10.6151
R19253 vdd.n2150 vdd.n2149 10.6151
R19254 vdd.n1892 vdd.n1891 10.6151
R19255 vdd.n1891 vdd.n1889 10.6151
R19256 vdd.n1889 vdd.n1888 10.6151
R19257 vdd.n1888 vdd.n1886 10.6151
R19258 vdd.n1886 vdd.n1885 10.6151
R19259 vdd.n1885 vdd.n1883 10.6151
R19260 vdd.n1883 vdd.n1882 10.6151
R19261 vdd.n1882 vdd.n1880 10.6151
R19262 vdd.n1880 vdd.n1879 10.6151
R19263 vdd.n1879 vdd.n1877 10.6151
R19264 vdd.n1877 vdd.n1876 10.6151
R19265 vdd.n1876 vdd.n1874 10.6151
R19266 vdd.n1874 vdd.n1873 10.6151
R19267 vdd.n1873 vdd.n1788 10.6151
R19268 vdd.n1788 vdd.n1787 10.6151
R19269 vdd.n1787 vdd.n1785 10.6151
R19270 vdd.n1785 vdd.n1784 10.6151
R19271 vdd.n1784 vdd.n1782 10.6151
R19272 vdd.n1782 vdd.n1781 10.6151
R19273 vdd.n1781 vdd.n1779 10.6151
R19274 vdd.n1779 vdd.n1778 10.6151
R19275 vdd.n1778 vdd.n1776 10.6151
R19276 vdd.n1776 vdd.n1775 10.6151
R19277 vdd.n1775 vdd.n1773 10.6151
R19278 vdd.n1773 vdd.n1772 10.6151
R19279 vdd.n1772 vdd.n1769 10.6151
R19280 vdd.n1769 vdd.n1768 10.6151
R19281 vdd.n1768 vdd.n749 10.6151
R19282 vdd.n1726 vdd.n837 10.6151
R19283 vdd.n1727 vdd.n1726 10.6151
R19284 vdd.n1728 vdd.n1727 10.6151
R19285 vdd.n1728 vdd.n1722 10.6151
R19286 vdd.n1734 vdd.n1722 10.6151
R19287 vdd.n1735 vdd.n1734 10.6151
R19288 vdd.n1736 vdd.n1735 10.6151
R19289 vdd.n1736 vdd.n1720 10.6151
R19290 vdd.n1742 vdd.n1720 10.6151
R19291 vdd.n1743 vdd.n1742 10.6151
R19292 vdd.n1744 vdd.n1743 10.6151
R19293 vdd.n1744 vdd.n1718 10.6151
R19294 vdd.n1750 vdd.n1718 10.6151
R19295 vdd.n1751 vdd.n1750 10.6151
R19296 vdd.n1752 vdd.n1751 10.6151
R19297 vdd.n1752 vdd.n1716 10.6151
R19298 vdd.n1928 vdd.n1716 10.6151
R19299 vdd.n1928 vdd.n1927 10.6151
R19300 vdd.n1927 vdd.n1757 10.6151
R19301 vdd.n1921 vdd.n1757 10.6151
R19302 vdd.n1921 vdd.n1920 10.6151
R19303 vdd.n1920 vdd.n1919 10.6151
R19304 vdd.n1919 vdd.n1759 10.6151
R19305 vdd.n1913 vdd.n1759 10.6151
R19306 vdd.n1913 vdd.n1912 10.6151
R19307 vdd.n1912 vdd.n1911 10.6151
R19308 vdd.n1911 vdd.n1761 10.6151
R19309 vdd.n1905 vdd.n1761 10.6151
R19310 vdd.n1905 vdd.n1904 10.6151
R19311 vdd.n1904 vdd.n1903 10.6151
R19312 vdd.n1903 vdd.n1763 10.6151
R19313 vdd.n1897 vdd.n1896 10.6151
R19314 vdd.n1896 vdd.n1895 10.6151
R19315 vdd.n2401 vdd.n2400 10.6151
R19316 vdd.n2400 vdd.n2398 10.6151
R19317 vdd.n2398 vdd.n2397 10.6151
R19318 vdd.n2397 vdd.n2255 10.6151
R19319 vdd.n2344 vdd.n2255 10.6151
R19320 vdd.n2345 vdd.n2344 10.6151
R19321 vdd.n2347 vdd.n2345 10.6151
R19322 vdd.n2348 vdd.n2347 10.6151
R19323 vdd.n2350 vdd.n2348 10.6151
R19324 vdd.n2351 vdd.n2350 10.6151
R19325 vdd.n2353 vdd.n2351 10.6151
R19326 vdd.n2354 vdd.n2353 10.6151
R19327 vdd.n2356 vdd.n2354 10.6151
R19328 vdd.n2357 vdd.n2356 10.6151
R19329 vdd.n2372 vdd.n2357 10.6151
R19330 vdd.n2372 vdd.n2371 10.6151
R19331 vdd.n2371 vdd.n2370 10.6151
R19332 vdd.n2370 vdd.n2368 10.6151
R19333 vdd.n2368 vdd.n2367 10.6151
R19334 vdd.n2367 vdd.n2365 10.6151
R19335 vdd.n2365 vdd.n2364 10.6151
R19336 vdd.n2364 vdd.n2362 10.6151
R19337 vdd.n2362 vdd.n2361 10.6151
R19338 vdd.n2361 vdd.n2359 10.6151
R19339 vdd.n2359 vdd.n2358 10.6151
R19340 vdd.n2358 vdd.n626 10.6151
R19341 vdd.n2606 vdd.n626 10.6151
R19342 vdd.n2607 vdd.n2606 10.6151
R19343 vdd.n2468 vdd.n702 10.6151
R19344 vdd.n2468 vdd.n2467 10.6151
R19345 vdd.n2467 vdd.n2466 10.6151
R19346 vdd.n2466 vdd.n2464 10.6151
R19347 vdd.n2464 vdd.n2461 10.6151
R19348 vdd.n2461 vdd.n2460 10.6151
R19349 vdd.n2460 vdd.n2457 10.6151
R19350 vdd.n2457 vdd.n2456 10.6151
R19351 vdd.n2456 vdd.n2453 10.6151
R19352 vdd.n2453 vdd.n2452 10.6151
R19353 vdd.n2452 vdd.n2449 10.6151
R19354 vdd.n2449 vdd.n2448 10.6151
R19355 vdd.n2448 vdd.n2445 10.6151
R19356 vdd.n2445 vdd.n2444 10.6151
R19357 vdd.n2444 vdd.n2441 10.6151
R19358 vdd.n2441 vdd.n2440 10.6151
R19359 vdd.n2440 vdd.n2437 10.6151
R19360 vdd.n2437 vdd.n2436 10.6151
R19361 vdd.n2436 vdd.n2433 10.6151
R19362 vdd.n2433 vdd.n2432 10.6151
R19363 vdd.n2432 vdd.n2429 10.6151
R19364 vdd.n2429 vdd.n2428 10.6151
R19365 vdd.n2428 vdd.n2425 10.6151
R19366 vdd.n2425 vdd.n2424 10.6151
R19367 vdd.n2424 vdd.n2421 10.6151
R19368 vdd.n2421 vdd.n2420 10.6151
R19369 vdd.n2420 vdd.n2417 10.6151
R19370 vdd.n2417 vdd.n2416 10.6151
R19371 vdd.n2416 vdd.n2413 10.6151
R19372 vdd.n2413 vdd.n2412 10.6151
R19373 vdd.n2412 vdd.n2409 10.6151
R19374 vdd.n2407 vdd.n2404 10.6151
R19375 vdd.n2404 vdd.n2403 10.6151
R19376 vdd.n2481 vdd.n2480 10.6151
R19377 vdd.n2482 vdd.n2481 10.6151
R19378 vdd.n2482 vdd.n692 10.6151
R19379 vdd.n2492 vdd.n692 10.6151
R19380 vdd.n2493 vdd.n2492 10.6151
R19381 vdd.n2494 vdd.n2493 10.6151
R19382 vdd.n2494 vdd.n679 10.6151
R19383 vdd.n2504 vdd.n679 10.6151
R19384 vdd.n2505 vdd.n2504 10.6151
R19385 vdd.n2506 vdd.n2505 10.6151
R19386 vdd.n2506 vdd.n668 10.6151
R19387 vdd.n2516 vdd.n668 10.6151
R19388 vdd.n2517 vdd.n2516 10.6151
R19389 vdd.n2518 vdd.n2517 10.6151
R19390 vdd.n2518 vdd.n656 10.6151
R19391 vdd.n2528 vdd.n656 10.6151
R19392 vdd.n2529 vdd.n2528 10.6151
R19393 vdd.n2530 vdd.n2529 10.6151
R19394 vdd.n2530 vdd.n645 10.6151
R19395 vdd.n2542 vdd.n645 10.6151
R19396 vdd.n2543 vdd.n2542 10.6151
R19397 vdd.n2544 vdd.n2543 10.6151
R19398 vdd.n2544 vdd.n631 10.6151
R19399 vdd.n2599 vdd.n631 10.6151
R19400 vdd.n2600 vdd.n2599 10.6151
R19401 vdd.n2601 vdd.n2600 10.6151
R19402 vdd.n2601 vdd.n600 10.6151
R19403 vdd.n2671 vdd.n600 10.6151
R19404 vdd.n2670 vdd.n2669 10.6151
R19405 vdd.n2669 vdd.n601 10.6151
R19406 vdd.n602 vdd.n601 10.6151
R19407 vdd.n2662 vdd.n602 10.6151
R19408 vdd.n2662 vdd.n2661 10.6151
R19409 vdd.n2661 vdd.n2660 10.6151
R19410 vdd.n2660 vdd.n604 10.6151
R19411 vdd.n2655 vdd.n604 10.6151
R19412 vdd.n2655 vdd.n2654 10.6151
R19413 vdd.n2654 vdd.n2653 10.6151
R19414 vdd.n2653 vdd.n607 10.6151
R19415 vdd.n2648 vdd.n607 10.6151
R19416 vdd.n2648 vdd.n2647 10.6151
R19417 vdd.n2647 vdd.n2646 10.6151
R19418 vdd.n2646 vdd.n610 10.6151
R19419 vdd.n2641 vdd.n610 10.6151
R19420 vdd.n2641 vdd.n520 10.6151
R19421 vdd.n2637 vdd.n520 10.6151
R19422 vdd.n2637 vdd.n2636 10.6151
R19423 vdd.n2636 vdd.n2635 10.6151
R19424 vdd.n2635 vdd.n613 10.6151
R19425 vdd.n2630 vdd.n613 10.6151
R19426 vdd.n2630 vdd.n2629 10.6151
R19427 vdd.n2629 vdd.n2628 10.6151
R19428 vdd.n2628 vdd.n616 10.6151
R19429 vdd.n2623 vdd.n616 10.6151
R19430 vdd.n2623 vdd.n2622 10.6151
R19431 vdd.n2622 vdd.n2621 10.6151
R19432 vdd.n2621 vdd.n619 10.6151
R19433 vdd.n2616 vdd.n619 10.6151
R19434 vdd.n2616 vdd.n2615 10.6151
R19435 vdd.n2613 vdd.n624 10.6151
R19436 vdd.n2608 vdd.n624 10.6151
R19437 vdd.n2589 vdd.n2550 10.6151
R19438 vdd.n2584 vdd.n2550 10.6151
R19439 vdd.n2584 vdd.n2583 10.6151
R19440 vdd.n2583 vdd.n2582 10.6151
R19441 vdd.n2582 vdd.n2552 10.6151
R19442 vdd.n2577 vdd.n2552 10.6151
R19443 vdd.n2577 vdd.n2576 10.6151
R19444 vdd.n2576 vdd.n2575 10.6151
R19445 vdd.n2575 vdd.n2555 10.6151
R19446 vdd.n2570 vdd.n2555 10.6151
R19447 vdd.n2570 vdd.n2569 10.6151
R19448 vdd.n2569 vdd.n2568 10.6151
R19449 vdd.n2568 vdd.n2558 10.6151
R19450 vdd.n2563 vdd.n2558 10.6151
R19451 vdd.n2563 vdd.n2562 10.6151
R19452 vdd.n2562 vdd.n575 10.6151
R19453 vdd.n2706 vdd.n575 10.6151
R19454 vdd.n2706 vdd.n576 10.6151
R19455 vdd.n578 vdd.n576 10.6151
R19456 vdd.n2699 vdd.n578 10.6151
R19457 vdd.n2699 vdd.n2698 10.6151
R19458 vdd.n2698 vdd.n2697 10.6151
R19459 vdd.n2697 vdd.n580 10.6151
R19460 vdd.n2692 vdd.n580 10.6151
R19461 vdd.n2692 vdd.n2691 10.6151
R19462 vdd.n2691 vdd.n2690 10.6151
R19463 vdd.n2690 vdd.n583 10.6151
R19464 vdd.n2685 vdd.n583 10.6151
R19465 vdd.n2685 vdd.n2684 10.6151
R19466 vdd.n2684 vdd.n2683 10.6151
R19467 vdd.n2683 vdd.n586 10.6151
R19468 vdd.n2678 vdd.n2677 10.6151
R19469 vdd.n2677 vdd.n2676 10.6151
R19470 vdd.n2324 vdd.n2322 10.6151
R19471 vdd.n2325 vdd.n2324 10.6151
R19472 vdd.n2393 vdd.n2325 10.6151
R19473 vdd.n2393 vdd.n2392 10.6151
R19474 vdd.n2392 vdd.n2391 10.6151
R19475 vdd.n2391 vdd.n2389 10.6151
R19476 vdd.n2389 vdd.n2388 10.6151
R19477 vdd.n2388 vdd.n2386 10.6151
R19478 vdd.n2386 vdd.n2385 10.6151
R19479 vdd.n2385 vdd.n2383 10.6151
R19480 vdd.n2383 vdd.n2382 10.6151
R19481 vdd.n2382 vdd.n2380 10.6151
R19482 vdd.n2380 vdd.n2379 10.6151
R19483 vdd.n2379 vdd.n2377 10.6151
R19484 vdd.n2377 vdd.n2376 10.6151
R19485 vdd.n2376 vdd.n2342 10.6151
R19486 vdd.n2342 vdd.n2341 10.6151
R19487 vdd.n2341 vdd.n2339 10.6151
R19488 vdd.n2339 vdd.n2338 10.6151
R19489 vdd.n2338 vdd.n2336 10.6151
R19490 vdd.n2336 vdd.n2335 10.6151
R19491 vdd.n2335 vdd.n2333 10.6151
R19492 vdd.n2333 vdd.n2332 10.6151
R19493 vdd.n2332 vdd.n2330 10.6151
R19494 vdd.n2330 vdd.n2329 10.6151
R19495 vdd.n2329 vdd.n2327 10.6151
R19496 vdd.n2327 vdd.n2326 10.6151
R19497 vdd.n2326 vdd.n592 10.6151
R19498 vdd.n2475 vdd.n2474 10.6151
R19499 vdd.n2474 vdd.n707 10.6151
R19500 vdd.n2259 vdd.n707 10.6151
R19501 vdd.n2262 vdd.n2259 10.6151
R19502 vdd.n2263 vdd.n2262 10.6151
R19503 vdd.n2266 vdd.n2263 10.6151
R19504 vdd.n2267 vdd.n2266 10.6151
R19505 vdd.n2270 vdd.n2267 10.6151
R19506 vdd.n2271 vdd.n2270 10.6151
R19507 vdd.n2274 vdd.n2271 10.6151
R19508 vdd.n2275 vdd.n2274 10.6151
R19509 vdd.n2278 vdd.n2275 10.6151
R19510 vdd.n2279 vdd.n2278 10.6151
R19511 vdd.n2282 vdd.n2279 10.6151
R19512 vdd.n2283 vdd.n2282 10.6151
R19513 vdd.n2286 vdd.n2283 10.6151
R19514 vdd.n2287 vdd.n2286 10.6151
R19515 vdd.n2290 vdd.n2287 10.6151
R19516 vdd.n2291 vdd.n2290 10.6151
R19517 vdd.n2294 vdd.n2291 10.6151
R19518 vdd.n2295 vdd.n2294 10.6151
R19519 vdd.n2298 vdd.n2295 10.6151
R19520 vdd.n2299 vdd.n2298 10.6151
R19521 vdd.n2302 vdd.n2299 10.6151
R19522 vdd.n2303 vdd.n2302 10.6151
R19523 vdd.n2306 vdd.n2303 10.6151
R19524 vdd.n2307 vdd.n2306 10.6151
R19525 vdd.n2310 vdd.n2307 10.6151
R19526 vdd.n2311 vdd.n2310 10.6151
R19527 vdd.n2314 vdd.n2311 10.6151
R19528 vdd.n2315 vdd.n2314 10.6151
R19529 vdd.n2320 vdd.n2318 10.6151
R19530 vdd.n2321 vdd.n2320 10.6151
R19531 vdd.n2476 vdd.n697 10.6151
R19532 vdd.n2486 vdd.n697 10.6151
R19533 vdd.n2487 vdd.n2486 10.6151
R19534 vdd.n2488 vdd.n2487 10.6151
R19535 vdd.n2488 vdd.n685 10.6151
R19536 vdd.n2498 vdd.n685 10.6151
R19537 vdd.n2499 vdd.n2498 10.6151
R19538 vdd.n2500 vdd.n2499 10.6151
R19539 vdd.n2500 vdd.n674 10.6151
R19540 vdd.n2510 vdd.n674 10.6151
R19541 vdd.n2511 vdd.n2510 10.6151
R19542 vdd.n2512 vdd.n2511 10.6151
R19543 vdd.n2512 vdd.n662 10.6151
R19544 vdd.n2522 vdd.n662 10.6151
R19545 vdd.n2523 vdd.n2522 10.6151
R19546 vdd.n2524 vdd.n2523 10.6151
R19547 vdd.n2524 vdd.n651 10.6151
R19548 vdd.n2534 vdd.n651 10.6151
R19549 vdd.n2535 vdd.n2534 10.6151
R19550 vdd.n2538 vdd.n2535 10.6151
R19551 vdd.n2548 vdd.n639 10.6151
R19552 vdd.n2549 vdd.n2548 10.6151
R19553 vdd.n2595 vdd.n2549 10.6151
R19554 vdd.n2595 vdd.n2594 10.6151
R19555 vdd.n2594 vdd.n2593 10.6151
R19556 vdd.n2593 vdd.n2592 10.6151
R19557 vdd.n2592 vdd.n2590 10.6151
R19558 vdd.n1987 vdd.n831 10.6151
R19559 vdd.n1997 vdd.n831 10.6151
R19560 vdd.n1998 vdd.n1997 10.6151
R19561 vdd.n1999 vdd.n1998 10.6151
R19562 vdd.n1999 vdd.n818 10.6151
R19563 vdd.n2009 vdd.n818 10.6151
R19564 vdd.n2010 vdd.n2009 10.6151
R19565 vdd.n2012 vdd.n806 10.6151
R19566 vdd.n2022 vdd.n806 10.6151
R19567 vdd.n2023 vdd.n2022 10.6151
R19568 vdd.n2024 vdd.n2023 10.6151
R19569 vdd.n2024 vdd.n794 10.6151
R19570 vdd.n2034 vdd.n794 10.6151
R19571 vdd.n2035 vdd.n2034 10.6151
R19572 vdd.n2036 vdd.n2035 10.6151
R19573 vdd.n2036 vdd.n783 10.6151
R19574 vdd.n2046 vdd.n783 10.6151
R19575 vdd.n2047 vdd.n2046 10.6151
R19576 vdd.n2048 vdd.n2047 10.6151
R19577 vdd.n2048 vdd.n771 10.6151
R19578 vdd.n2058 vdd.n771 10.6151
R19579 vdd.n2059 vdd.n2058 10.6151
R19580 vdd.n2062 vdd.n2059 10.6151
R19581 vdd.n2062 vdd.n2061 10.6151
R19582 vdd.n2061 vdd.n2060 10.6151
R19583 vdd.n2060 vdd.n754 10.6151
R19584 vdd.n2144 vdd.n754 10.6151
R19585 vdd.n2143 vdd.n2142 10.6151
R19586 vdd.n2142 vdd.n2139 10.6151
R19587 vdd.n2139 vdd.n2138 10.6151
R19588 vdd.n2138 vdd.n2135 10.6151
R19589 vdd.n2135 vdd.n2134 10.6151
R19590 vdd.n2134 vdd.n2131 10.6151
R19591 vdd.n2131 vdd.n2130 10.6151
R19592 vdd.n2130 vdd.n2127 10.6151
R19593 vdd.n2127 vdd.n2126 10.6151
R19594 vdd.n2126 vdd.n2123 10.6151
R19595 vdd.n2123 vdd.n2122 10.6151
R19596 vdd.n2122 vdd.n2119 10.6151
R19597 vdd.n2119 vdd.n2118 10.6151
R19598 vdd.n2118 vdd.n2115 10.6151
R19599 vdd.n2115 vdd.n2114 10.6151
R19600 vdd.n2114 vdd.n2111 10.6151
R19601 vdd.n2111 vdd.n2110 10.6151
R19602 vdd.n2110 vdd.n2107 10.6151
R19603 vdd.n2107 vdd.n2106 10.6151
R19604 vdd.n2106 vdd.n2103 10.6151
R19605 vdd.n2103 vdd.n2102 10.6151
R19606 vdd.n2102 vdd.n2099 10.6151
R19607 vdd.n2099 vdd.n2098 10.6151
R19608 vdd.n2098 vdd.n2095 10.6151
R19609 vdd.n2095 vdd.n2094 10.6151
R19610 vdd.n2094 vdd.n2091 10.6151
R19611 vdd.n2091 vdd.n2090 10.6151
R19612 vdd.n2090 vdd.n2087 10.6151
R19613 vdd.n2087 vdd.n2086 10.6151
R19614 vdd.n2086 vdd.n2083 10.6151
R19615 vdd.n2083 vdd.n2082 10.6151
R19616 vdd.n2079 vdd.n2078 10.6151
R19617 vdd.n2078 vdd.n2076 10.6151
R19618 vdd.n1835 vdd.n1833 10.6151
R19619 vdd.n1836 vdd.n1835 10.6151
R19620 vdd.n1838 vdd.n1836 10.6151
R19621 vdd.n1839 vdd.n1838 10.6151
R19622 vdd.n1841 vdd.n1839 10.6151
R19623 vdd.n1842 vdd.n1841 10.6151
R19624 vdd.n1844 vdd.n1842 10.6151
R19625 vdd.n1845 vdd.n1844 10.6151
R19626 vdd.n1847 vdd.n1845 10.6151
R19627 vdd.n1848 vdd.n1847 10.6151
R19628 vdd.n1850 vdd.n1848 10.6151
R19629 vdd.n1851 vdd.n1850 10.6151
R19630 vdd.n1869 vdd.n1851 10.6151
R19631 vdd.n1869 vdd.n1868 10.6151
R19632 vdd.n1868 vdd.n1867 10.6151
R19633 vdd.n1867 vdd.n1865 10.6151
R19634 vdd.n1865 vdd.n1864 10.6151
R19635 vdd.n1864 vdd.n1862 10.6151
R19636 vdd.n1862 vdd.n1861 10.6151
R19637 vdd.n1861 vdd.n1859 10.6151
R19638 vdd.n1859 vdd.n1858 10.6151
R19639 vdd.n1858 vdd.n1856 10.6151
R19640 vdd.n1856 vdd.n1855 10.6151
R19641 vdd.n1855 vdd.n1853 10.6151
R19642 vdd.n1853 vdd.n1852 10.6151
R19643 vdd.n1852 vdd.n758 10.6151
R19644 vdd.n2074 vdd.n758 10.6151
R19645 vdd.n2075 vdd.n2074 10.6151
R19646 vdd.n1986 vdd.n1985 10.6151
R19647 vdd.n1985 vdd.n843 10.6151
R19648 vdd.n1979 vdd.n843 10.6151
R19649 vdd.n1979 vdd.n1978 10.6151
R19650 vdd.n1978 vdd.n1977 10.6151
R19651 vdd.n1977 vdd.n845 10.6151
R19652 vdd.n1971 vdd.n845 10.6151
R19653 vdd.n1971 vdd.n1970 10.6151
R19654 vdd.n1970 vdd.n1969 10.6151
R19655 vdd.n1969 vdd.n847 10.6151
R19656 vdd.n1963 vdd.n847 10.6151
R19657 vdd.n1963 vdd.n1962 10.6151
R19658 vdd.n1962 vdd.n1961 10.6151
R19659 vdd.n1961 vdd.n849 10.6151
R19660 vdd.n1955 vdd.n849 10.6151
R19661 vdd.n1955 vdd.n1954 10.6151
R19662 vdd.n1954 vdd.n1953 10.6151
R19663 vdd.n1953 vdd.n853 10.6151
R19664 vdd.n1801 vdd.n853 10.6151
R19665 vdd.n1802 vdd.n1801 10.6151
R19666 vdd.n1802 vdd.n1797 10.6151
R19667 vdd.n1808 vdd.n1797 10.6151
R19668 vdd.n1809 vdd.n1808 10.6151
R19669 vdd.n1810 vdd.n1809 10.6151
R19670 vdd.n1810 vdd.n1795 10.6151
R19671 vdd.n1816 vdd.n1795 10.6151
R19672 vdd.n1817 vdd.n1816 10.6151
R19673 vdd.n1818 vdd.n1817 10.6151
R19674 vdd.n1818 vdd.n1793 10.6151
R19675 vdd.n1824 vdd.n1793 10.6151
R19676 vdd.n1825 vdd.n1824 10.6151
R19677 vdd.n1827 vdd.n1789 10.6151
R19678 vdd.n1832 vdd.n1789 10.6151
R19679 vdd.n280 vdd.n262 10.4732
R19680 vdd.n233 vdd.n215 10.4732
R19681 vdd.n190 vdd.n172 10.4732
R19682 vdd.n143 vdd.n125 10.4732
R19683 vdd.n101 vdd.n83 10.4732
R19684 vdd.n54 vdd.n36 10.4732
R19685 vdd.n1095 vdd.n1077 10.4732
R19686 vdd.n1142 vdd.n1124 10.4732
R19687 vdd.n1005 vdd.n987 10.4732
R19688 vdd.n1052 vdd.n1034 10.4732
R19689 vdd.n916 vdd.n898 10.4732
R19690 vdd.n963 vdd.n945 10.4732
R19691 vdd.t9 vdd.n888 10.3167
R19692 vdd.n2874 vdd.t29 10.3167
R19693 vdd.n1465 vdd.t5 10.09
R19694 vdd.n3042 vdd.t42 10.09
R19695 vdd.n279 vdd.n264 9.69747
R19696 vdd.n232 vdd.n217 9.69747
R19697 vdd.n189 vdd.n174 9.69747
R19698 vdd.n142 vdd.n127 9.69747
R19699 vdd.n100 vdd.n85 9.69747
R19700 vdd.n53 vdd.n38 9.69747
R19701 vdd.n1094 vdd.n1079 9.69747
R19702 vdd.n1141 vdd.n1126 9.69747
R19703 vdd.n1004 vdd.n989 9.69747
R19704 vdd.n1051 vdd.n1036 9.69747
R19705 vdd.n915 vdd.n900 9.69747
R19706 vdd.n962 vdd.n947 9.69747
R19707 vdd.n1929 vdd.n1928 9.67831
R19708 vdd.n2836 vdd.n520 9.67831
R19709 vdd.n2707 vdd.n2706 9.67831
R19710 vdd.n1953 vdd.n1952 9.67831
R19711 vdd.n295 vdd.n294 9.45567
R19712 vdd.n248 vdd.n247 9.45567
R19713 vdd.n205 vdd.n204 9.45567
R19714 vdd.n158 vdd.n157 9.45567
R19715 vdd.n116 vdd.n115 9.45567
R19716 vdd.n69 vdd.n68 9.45567
R19717 vdd.n1110 vdd.n1109 9.45567
R19718 vdd.n1157 vdd.n1156 9.45567
R19719 vdd.n1020 vdd.n1019 9.45567
R19720 vdd.n1067 vdd.n1066 9.45567
R19721 vdd.n931 vdd.n930 9.45567
R19722 vdd.n978 vdd.n977 9.45567
R19723 vdd.n1689 vdd.n1543 9.3005
R19724 vdd.n1688 vdd.n1687 9.3005
R19725 vdd.n1549 vdd.n1548 9.3005
R19726 vdd.n1682 vdd.n1553 9.3005
R19727 vdd.n1681 vdd.n1554 9.3005
R19728 vdd.n1680 vdd.n1555 9.3005
R19729 vdd.n1559 vdd.n1556 9.3005
R19730 vdd.n1675 vdd.n1560 9.3005
R19731 vdd.n1674 vdd.n1561 9.3005
R19732 vdd.n1673 vdd.n1562 9.3005
R19733 vdd.n1566 vdd.n1563 9.3005
R19734 vdd.n1668 vdd.n1567 9.3005
R19735 vdd.n1667 vdd.n1568 9.3005
R19736 vdd.n1666 vdd.n1569 9.3005
R19737 vdd.n1573 vdd.n1570 9.3005
R19738 vdd.n1661 vdd.n1574 9.3005
R19739 vdd.n1660 vdd.n1575 9.3005
R19740 vdd.n1659 vdd.n1576 9.3005
R19741 vdd.n1580 vdd.n1577 9.3005
R19742 vdd.n1654 vdd.n1581 9.3005
R19743 vdd.n1653 vdd.n1582 9.3005
R19744 vdd.n1652 vdd.n1651 9.3005
R19745 vdd.n1650 vdd.n1583 9.3005
R19746 vdd.n1649 vdd.n1648 9.3005
R19747 vdd.n1589 vdd.n1588 9.3005
R19748 vdd.n1643 vdd.n1593 9.3005
R19749 vdd.n1642 vdd.n1594 9.3005
R19750 vdd.n1641 vdd.n1595 9.3005
R19751 vdd.n1599 vdd.n1596 9.3005
R19752 vdd.n1636 vdd.n1600 9.3005
R19753 vdd.n1635 vdd.n1601 9.3005
R19754 vdd.n1634 vdd.n1602 9.3005
R19755 vdd.n1606 vdd.n1603 9.3005
R19756 vdd.n1629 vdd.n1607 9.3005
R19757 vdd.n1628 vdd.n1608 9.3005
R19758 vdd.n1627 vdd.n1609 9.3005
R19759 vdd.n1611 vdd.n1610 9.3005
R19760 vdd.n1622 vdd.n854 9.3005
R19761 vdd.n1691 vdd.n1690 9.3005
R19762 vdd.n1715 vdd.n1714 9.3005
R19763 vdd.n1521 vdd.n1520 9.3005
R19764 vdd.n1526 vdd.n1524 9.3005
R19765 vdd.n1707 vdd.n1527 9.3005
R19766 vdd.n1706 vdd.n1528 9.3005
R19767 vdd.n1705 vdd.n1529 9.3005
R19768 vdd.n1533 vdd.n1530 9.3005
R19769 vdd.n1700 vdd.n1534 9.3005
R19770 vdd.n1699 vdd.n1535 9.3005
R19771 vdd.n1698 vdd.n1536 9.3005
R19772 vdd.n1540 vdd.n1537 9.3005
R19773 vdd.n1693 vdd.n1541 9.3005
R19774 vdd.n1692 vdd.n1542 9.3005
R19775 vdd.n1937 vdd.n1514 9.3005
R19776 vdd.n1939 vdd.n1938 9.3005
R19777 vdd.n1476 vdd.n1475 9.3005
R19778 vdd.n1477 vdd.n890 9.3005
R19779 vdd.n1479 vdd.n1478 9.3005
R19780 vdd.n880 vdd.n879 9.3005
R19781 vdd.n1493 vdd.n1492 9.3005
R19782 vdd.n1494 vdd.n878 9.3005
R19783 vdd.n1496 vdd.n1495 9.3005
R19784 vdd.n868 vdd.n867 9.3005
R19785 vdd.n1512 vdd.n1511 9.3005
R19786 vdd.n1513 vdd.n866 9.3005
R19787 vdd.n1941 vdd.n1940 9.3005
R19788 vdd.n271 vdd.n270 9.3005
R19789 vdd.n266 vdd.n265 9.3005
R19790 vdd.n277 vdd.n276 9.3005
R19791 vdd.n279 vdd.n278 9.3005
R19792 vdd.n262 vdd.n261 9.3005
R19793 vdd.n285 vdd.n284 9.3005
R19794 vdd.n287 vdd.n286 9.3005
R19795 vdd.n259 vdd.n256 9.3005
R19796 vdd.n294 vdd.n293 9.3005
R19797 vdd.n224 vdd.n223 9.3005
R19798 vdd.n219 vdd.n218 9.3005
R19799 vdd.n230 vdd.n229 9.3005
R19800 vdd.n232 vdd.n231 9.3005
R19801 vdd.n215 vdd.n214 9.3005
R19802 vdd.n238 vdd.n237 9.3005
R19803 vdd.n240 vdd.n239 9.3005
R19804 vdd.n212 vdd.n209 9.3005
R19805 vdd.n247 vdd.n246 9.3005
R19806 vdd.n181 vdd.n180 9.3005
R19807 vdd.n176 vdd.n175 9.3005
R19808 vdd.n187 vdd.n186 9.3005
R19809 vdd.n189 vdd.n188 9.3005
R19810 vdd.n172 vdd.n171 9.3005
R19811 vdd.n195 vdd.n194 9.3005
R19812 vdd.n197 vdd.n196 9.3005
R19813 vdd.n169 vdd.n166 9.3005
R19814 vdd.n204 vdd.n203 9.3005
R19815 vdd.n134 vdd.n133 9.3005
R19816 vdd.n129 vdd.n128 9.3005
R19817 vdd.n140 vdd.n139 9.3005
R19818 vdd.n142 vdd.n141 9.3005
R19819 vdd.n125 vdd.n124 9.3005
R19820 vdd.n148 vdd.n147 9.3005
R19821 vdd.n150 vdd.n149 9.3005
R19822 vdd.n122 vdd.n119 9.3005
R19823 vdd.n157 vdd.n156 9.3005
R19824 vdd.n92 vdd.n91 9.3005
R19825 vdd.n87 vdd.n86 9.3005
R19826 vdd.n98 vdd.n97 9.3005
R19827 vdd.n100 vdd.n99 9.3005
R19828 vdd.n83 vdd.n82 9.3005
R19829 vdd.n106 vdd.n105 9.3005
R19830 vdd.n108 vdd.n107 9.3005
R19831 vdd.n80 vdd.n77 9.3005
R19832 vdd.n115 vdd.n114 9.3005
R19833 vdd.n45 vdd.n44 9.3005
R19834 vdd.n40 vdd.n39 9.3005
R19835 vdd.n51 vdd.n50 9.3005
R19836 vdd.n53 vdd.n52 9.3005
R19837 vdd.n36 vdd.n35 9.3005
R19838 vdd.n59 vdd.n58 9.3005
R19839 vdd.n61 vdd.n60 9.3005
R19840 vdd.n33 vdd.n30 9.3005
R19841 vdd.n68 vdd.n67 9.3005
R19842 vdd.n2758 vdd.n2757 9.3005
R19843 vdd.n2761 vdd.n555 9.3005
R19844 vdd.n2762 vdd.n554 9.3005
R19845 vdd.n2765 vdd.n553 9.3005
R19846 vdd.n2766 vdd.n552 9.3005
R19847 vdd.n2769 vdd.n551 9.3005
R19848 vdd.n2770 vdd.n550 9.3005
R19849 vdd.n2773 vdd.n549 9.3005
R19850 vdd.n2774 vdd.n548 9.3005
R19851 vdd.n2777 vdd.n547 9.3005
R19852 vdd.n2778 vdd.n546 9.3005
R19853 vdd.n2781 vdd.n545 9.3005
R19854 vdd.n2782 vdd.n544 9.3005
R19855 vdd.n2785 vdd.n543 9.3005
R19856 vdd.n2786 vdd.n542 9.3005
R19857 vdd.n2789 vdd.n541 9.3005
R19858 vdd.n2790 vdd.n540 9.3005
R19859 vdd.n2793 vdd.n539 9.3005
R19860 vdd.n2794 vdd.n538 9.3005
R19861 vdd.n2797 vdd.n537 9.3005
R19862 vdd.n2801 vdd.n2800 9.3005
R19863 vdd.n2802 vdd.n536 9.3005
R19864 vdd.n2806 vdd.n2803 9.3005
R19865 vdd.n2809 vdd.n535 9.3005
R19866 vdd.n2810 vdd.n534 9.3005
R19867 vdd.n2813 vdd.n533 9.3005
R19868 vdd.n2814 vdd.n532 9.3005
R19869 vdd.n2817 vdd.n531 9.3005
R19870 vdd.n2818 vdd.n530 9.3005
R19871 vdd.n2821 vdd.n529 9.3005
R19872 vdd.n2822 vdd.n528 9.3005
R19873 vdd.n2825 vdd.n527 9.3005
R19874 vdd.n2826 vdd.n526 9.3005
R19875 vdd.n2829 vdd.n525 9.3005
R19876 vdd.n2830 vdd.n524 9.3005
R19877 vdd.n2833 vdd.n519 9.3005
R19878 vdd.n482 vdd.n481 9.3005
R19879 vdd.n2844 vdd.n2843 9.3005
R19880 vdd.n2847 vdd.n2846 9.3005
R19881 vdd.n471 vdd.n470 9.3005
R19882 vdd.n2861 vdd.n2860 9.3005
R19883 vdd.n2862 vdd.n469 9.3005
R19884 vdd.n2864 vdd.n2863 9.3005
R19885 vdd.n460 vdd.n459 9.3005
R19886 vdd.n2877 vdd.n2876 9.3005
R19887 vdd.n2878 vdd.n458 9.3005
R19888 vdd.n2880 vdd.n2879 9.3005
R19889 vdd.n300 vdd.n298 9.3005
R19890 vdd.n2845 vdd.n480 9.3005
R19891 vdd.n3046 vdd.n3045 9.3005
R19892 vdd.n301 vdd.n299 9.3005
R19893 vdd.n3039 vdd.n310 9.3005
R19894 vdd.n3038 vdd.n311 9.3005
R19895 vdd.n3037 vdd.n312 9.3005
R19896 vdd.n320 vdd.n313 9.3005
R19897 vdd.n3031 vdd.n321 9.3005
R19898 vdd.n3030 vdd.n322 9.3005
R19899 vdd.n3029 vdd.n323 9.3005
R19900 vdd.n331 vdd.n324 9.3005
R19901 vdd.n3023 vdd.n3022 9.3005
R19902 vdd.n3019 vdd.n332 9.3005
R19903 vdd.n3018 vdd.n335 9.3005
R19904 vdd.n339 vdd.n336 9.3005
R19905 vdd.n340 vdd.n337 9.3005
R19906 vdd.n3011 vdd.n341 9.3005
R19907 vdd.n3010 vdd.n342 9.3005
R19908 vdd.n3009 vdd.n343 9.3005
R19909 vdd.n347 vdd.n344 9.3005
R19910 vdd.n3004 vdd.n348 9.3005
R19911 vdd.n3003 vdd.n349 9.3005
R19912 vdd.n3002 vdd.n350 9.3005
R19913 vdd.n354 vdd.n351 9.3005
R19914 vdd.n2997 vdd.n355 9.3005
R19915 vdd.n2996 vdd.n356 9.3005
R19916 vdd.n2995 vdd.n357 9.3005
R19917 vdd.n361 vdd.n358 9.3005
R19918 vdd.n2990 vdd.n362 9.3005
R19919 vdd.n2989 vdd.n363 9.3005
R19920 vdd.n2988 vdd.n2987 9.3005
R19921 vdd.n2986 vdd.n364 9.3005
R19922 vdd.n2985 vdd.n2984 9.3005
R19923 vdd.n370 vdd.n369 9.3005
R19924 vdd.n2979 vdd.n374 9.3005
R19925 vdd.n2978 vdd.n375 9.3005
R19926 vdd.n2977 vdd.n376 9.3005
R19927 vdd.n380 vdd.n377 9.3005
R19928 vdd.n2972 vdd.n381 9.3005
R19929 vdd.n2971 vdd.n382 9.3005
R19930 vdd.n2970 vdd.n383 9.3005
R19931 vdd.n387 vdd.n384 9.3005
R19932 vdd.n2965 vdd.n388 9.3005
R19933 vdd.n2964 vdd.n389 9.3005
R19934 vdd.n2963 vdd.n390 9.3005
R19935 vdd.n394 vdd.n391 9.3005
R19936 vdd.n2958 vdd.n395 9.3005
R19937 vdd.n2957 vdd.n396 9.3005
R19938 vdd.n2956 vdd.n397 9.3005
R19939 vdd.n401 vdd.n398 9.3005
R19940 vdd.n2951 vdd.n402 9.3005
R19941 vdd.n2950 vdd.n403 9.3005
R19942 vdd.n2949 vdd.n2948 9.3005
R19943 vdd.n2947 vdd.n404 9.3005
R19944 vdd.n2946 vdd.n2945 9.3005
R19945 vdd.n410 vdd.n409 9.3005
R19946 vdd.n2940 vdd.n414 9.3005
R19947 vdd.n2939 vdd.n415 9.3005
R19948 vdd.n2938 vdd.n416 9.3005
R19949 vdd.n420 vdd.n417 9.3005
R19950 vdd.n2933 vdd.n421 9.3005
R19951 vdd.n2932 vdd.n422 9.3005
R19952 vdd.n2931 vdd.n423 9.3005
R19953 vdd.n427 vdd.n424 9.3005
R19954 vdd.n2926 vdd.n428 9.3005
R19955 vdd.n2925 vdd.n429 9.3005
R19956 vdd.n2924 vdd.n430 9.3005
R19957 vdd.n434 vdd.n431 9.3005
R19958 vdd.n2919 vdd.n435 9.3005
R19959 vdd.n2918 vdd.n436 9.3005
R19960 vdd.n2917 vdd.n437 9.3005
R19961 vdd.n441 vdd.n438 9.3005
R19962 vdd.n2912 vdd.n442 9.3005
R19963 vdd.n2911 vdd.n443 9.3005
R19964 vdd.n2907 vdd.n2904 9.3005
R19965 vdd.n3021 vdd.n3020 9.3005
R19966 vdd.n2852 vdd.n2851 9.3005
R19967 vdd.n2853 vdd.n475 9.3005
R19968 vdd.n2855 vdd.n2854 9.3005
R19969 vdd.n465 vdd.n464 9.3005
R19970 vdd.n2869 vdd.n2868 9.3005
R19971 vdd.n2870 vdd.n463 9.3005
R19972 vdd.n2872 vdd.n2871 9.3005
R19973 vdd.n453 vdd.n452 9.3005
R19974 vdd.n2885 vdd.n2884 9.3005
R19975 vdd.n2886 vdd.n451 9.3005
R19976 vdd.n2888 vdd.n2887 9.3005
R19977 vdd.n2889 vdd.n450 9.3005
R19978 vdd.n2891 vdd.n2890 9.3005
R19979 vdd.n2892 vdd.n449 9.3005
R19980 vdd.n2894 vdd.n2893 9.3005
R19981 vdd.n2895 vdd.n447 9.3005
R19982 vdd.n2897 vdd.n2896 9.3005
R19983 vdd.n2898 vdd.n446 9.3005
R19984 vdd.n2900 vdd.n2899 9.3005
R19985 vdd.n2901 vdd.n444 9.3005
R19986 vdd.n2903 vdd.n2902 9.3005
R19987 vdd.n477 vdd.n476 9.3005
R19988 vdd.n2710 vdd.n2709 9.3005
R19989 vdd.n2715 vdd.n2708 9.3005
R19990 vdd.n2724 vdd.n572 9.3005
R19991 vdd.n2727 vdd.n571 9.3005
R19992 vdd.n2728 vdd.n570 9.3005
R19993 vdd.n2731 vdd.n569 9.3005
R19994 vdd.n2732 vdd.n568 9.3005
R19995 vdd.n2735 vdd.n567 9.3005
R19996 vdd.n2736 vdd.n566 9.3005
R19997 vdd.n2739 vdd.n565 9.3005
R19998 vdd.n2740 vdd.n564 9.3005
R19999 vdd.n2743 vdd.n563 9.3005
R20000 vdd.n2744 vdd.n562 9.3005
R20001 vdd.n2747 vdd.n561 9.3005
R20002 vdd.n2748 vdd.n560 9.3005
R20003 vdd.n2751 vdd.n559 9.3005
R20004 vdd.n2755 vdd.n2754 9.3005
R20005 vdd.n2756 vdd.n556 9.3005
R20006 vdd.n1951 vdd.n1950 9.3005
R20007 vdd.n1946 vdd.n857 9.3005
R20008 vdd.n1433 vdd.n1432 9.3005
R20009 vdd.n1434 vdd.n1188 9.3005
R20010 vdd.n1436 vdd.n1435 9.3005
R20011 vdd.n1178 vdd.n1177 9.3005
R20012 vdd.n1450 vdd.n1449 9.3005
R20013 vdd.n1451 vdd.n1176 9.3005
R20014 vdd.n1453 vdd.n1452 9.3005
R20015 vdd.n1168 vdd.n1167 9.3005
R20016 vdd.n1468 vdd.n1467 9.3005
R20017 vdd.n1469 vdd.n1166 9.3005
R20018 vdd.n1471 vdd.n1470 9.3005
R20019 vdd.n885 vdd.n884 9.3005
R20020 vdd.n1484 vdd.n1483 9.3005
R20021 vdd.n1485 vdd.n883 9.3005
R20022 vdd.n1487 vdd.n1486 9.3005
R20023 vdd.n875 vdd.n874 9.3005
R20024 vdd.n1501 vdd.n1500 9.3005
R20025 vdd.n1502 vdd.n872 9.3005
R20026 vdd.n1506 vdd.n1505 9.3005
R20027 vdd.n1504 vdd.n873 9.3005
R20028 vdd.n1503 vdd.n862 9.3005
R20029 vdd.n1190 vdd.n1189 9.3005
R20030 vdd.n1326 vdd.n1325 9.3005
R20031 vdd.n1327 vdd.n1316 9.3005
R20032 vdd.n1329 vdd.n1328 9.3005
R20033 vdd.n1330 vdd.n1315 9.3005
R20034 vdd.n1332 vdd.n1331 9.3005
R20035 vdd.n1333 vdd.n1310 9.3005
R20036 vdd.n1335 vdd.n1334 9.3005
R20037 vdd.n1336 vdd.n1309 9.3005
R20038 vdd.n1338 vdd.n1337 9.3005
R20039 vdd.n1339 vdd.n1304 9.3005
R20040 vdd.n1341 vdd.n1340 9.3005
R20041 vdd.n1342 vdd.n1303 9.3005
R20042 vdd.n1344 vdd.n1343 9.3005
R20043 vdd.n1345 vdd.n1298 9.3005
R20044 vdd.n1347 vdd.n1346 9.3005
R20045 vdd.n1348 vdd.n1297 9.3005
R20046 vdd.n1350 vdd.n1349 9.3005
R20047 vdd.n1351 vdd.n1292 9.3005
R20048 vdd.n1353 vdd.n1352 9.3005
R20049 vdd.n1354 vdd.n1291 9.3005
R20050 vdd.n1356 vdd.n1355 9.3005
R20051 vdd.n1360 vdd.n1287 9.3005
R20052 vdd.n1362 vdd.n1361 9.3005
R20053 vdd.n1363 vdd.n1286 9.3005
R20054 vdd.n1365 vdd.n1364 9.3005
R20055 vdd.n1366 vdd.n1281 9.3005
R20056 vdd.n1368 vdd.n1367 9.3005
R20057 vdd.n1369 vdd.n1280 9.3005
R20058 vdd.n1371 vdd.n1370 9.3005
R20059 vdd.n1372 vdd.n1275 9.3005
R20060 vdd.n1374 vdd.n1373 9.3005
R20061 vdd.n1375 vdd.n1274 9.3005
R20062 vdd.n1377 vdd.n1376 9.3005
R20063 vdd.n1378 vdd.n1269 9.3005
R20064 vdd.n1380 vdd.n1379 9.3005
R20065 vdd.n1381 vdd.n1268 9.3005
R20066 vdd.n1383 vdd.n1382 9.3005
R20067 vdd.n1384 vdd.n1263 9.3005
R20068 vdd.n1386 vdd.n1385 9.3005
R20069 vdd.n1387 vdd.n1262 9.3005
R20070 vdd.n1389 vdd.n1388 9.3005
R20071 vdd.n1390 vdd.n1257 9.3005
R20072 vdd.n1392 vdd.n1391 9.3005
R20073 vdd.n1393 vdd.n1256 9.3005
R20074 vdd.n1395 vdd.n1394 9.3005
R20075 vdd.n1396 vdd.n1249 9.3005
R20076 vdd.n1398 vdd.n1397 9.3005
R20077 vdd.n1399 vdd.n1248 9.3005
R20078 vdd.n1401 vdd.n1400 9.3005
R20079 vdd.n1402 vdd.n1243 9.3005
R20080 vdd.n1404 vdd.n1403 9.3005
R20081 vdd.n1405 vdd.n1242 9.3005
R20082 vdd.n1407 vdd.n1406 9.3005
R20083 vdd.n1408 vdd.n1237 9.3005
R20084 vdd.n1410 vdd.n1409 9.3005
R20085 vdd.n1411 vdd.n1236 9.3005
R20086 vdd.n1413 vdd.n1412 9.3005
R20087 vdd.n1414 vdd.n1231 9.3005
R20088 vdd.n1416 vdd.n1415 9.3005
R20089 vdd.n1417 vdd.n1230 9.3005
R20090 vdd.n1419 vdd.n1418 9.3005
R20091 vdd.n1195 vdd.n1194 9.3005
R20092 vdd.n1425 vdd.n1424 9.3005
R20093 vdd.n1324 vdd.n1323 9.3005
R20094 vdd.n1428 vdd.n1427 9.3005
R20095 vdd.n1184 vdd.n1183 9.3005
R20096 vdd.n1442 vdd.n1441 9.3005
R20097 vdd.n1443 vdd.n1182 9.3005
R20098 vdd.n1445 vdd.n1444 9.3005
R20099 vdd.n1173 vdd.n1172 9.3005
R20100 vdd.n1459 vdd.n1458 9.3005
R20101 vdd.n1460 vdd.n1171 9.3005
R20102 vdd.n1463 vdd.n1462 9.3005
R20103 vdd.n1461 vdd.n1162 9.3005
R20104 vdd.n1426 vdd.n1193 9.3005
R20105 vdd.n1086 vdd.n1085 9.3005
R20106 vdd.n1081 vdd.n1080 9.3005
R20107 vdd.n1092 vdd.n1091 9.3005
R20108 vdd.n1094 vdd.n1093 9.3005
R20109 vdd.n1077 vdd.n1076 9.3005
R20110 vdd.n1100 vdd.n1099 9.3005
R20111 vdd.n1102 vdd.n1101 9.3005
R20112 vdd.n1074 vdd.n1071 9.3005
R20113 vdd.n1109 vdd.n1108 9.3005
R20114 vdd.n1133 vdd.n1132 9.3005
R20115 vdd.n1128 vdd.n1127 9.3005
R20116 vdd.n1139 vdd.n1138 9.3005
R20117 vdd.n1141 vdd.n1140 9.3005
R20118 vdd.n1124 vdd.n1123 9.3005
R20119 vdd.n1147 vdd.n1146 9.3005
R20120 vdd.n1149 vdd.n1148 9.3005
R20121 vdd.n1121 vdd.n1118 9.3005
R20122 vdd.n1156 vdd.n1155 9.3005
R20123 vdd.n996 vdd.n995 9.3005
R20124 vdd.n991 vdd.n990 9.3005
R20125 vdd.n1002 vdd.n1001 9.3005
R20126 vdd.n1004 vdd.n1003 9.3005
R20127 vdd.n987 vdd.n986 9.3005
R20128 vdd.n1010 vdd.n1009 9.3005
R20129 vdd.n1012 vdd.n1011 9.3005
R20130 vdd.n984 vdd.n981 9.3005
R20131 vdd.n1019 vdd.n1018 9.3005
R20132 vdd.n1043 vdd.n1042 9.3005
R20133 vdd.n1038 vdd.n1037 9.3005
R20134 vdd.n1049 vdd.n1048 9.3005
R20135 vdd.n1051 vdd.n1050 9.3005
R20136 vdd.n1034 vdd.n1033 9.3005
R20137 vdd.n1057 vdd.n1056 9.3005
R20138 vdd.n1059 vdd.n1058 9.3005
R20139 vdd.n1031 vdd.n1028 9.3005
R20140 vdd.n1066 vdd.n1065 9.3005
R20141 vdd.n907 vdd.n906 9.3005
R20142 vdd.n902 vdd.n901 9.3005
R20143 vdd.n913 vdd.n912 9.3005
R20144 vdd.n915 vdd.n914 9.3005
R20145 vdd.n898 vdd.n897 9.3005
R20146 vdd.n921 vdd.n920 9.3005
R20147 vdd.n923 vdd.n922 9.3005
R20148 vdd.n895 vdd.n892 9.3005
R20149 vdd.n930 vdd.n929 9.3005
R20150 vdd.n954 vdd.n953 9.3005
R20151 vdd.n949 vdd.n948 9.3005
R20152 vdd.n960 vdd.n959 9.3005
R20153 vdd.n962 vdd.n961 9.3005
R20154 vdd.n945 vdd.n944 9.3005
R20155 vdd.n968 vdd.n967 9.3005
R20156 vdd.n970 vdd.n969 9.3005
R20157 vdd.n942 vdd.n939 9.3005
R20158 vdd.n977 vdd.n976 9.3005
R20159 vdd.n1438 vdd.t38 8.95635
R20160 vdd.t20 vdd.n3033 8.95635
R20161 vdd.n276 vdd.n275 8.92171
R20162 vdd.n229 vdd.n228 8.92171
R20163 vdd.n186 vdd.n185 8.92171
R20164 vdd.n139 vdd.n138 8.92171
R20165 vdd.n97 vdd.n96 8.92171
R20166 vdd.n50 vdd.n49 8.92171
R20167 vdd.n1091 vdd.n1090 8.92171
R20168 vdd.n1138 vdd.n1137 8.92171
R20169 vdd.n1001 vdd.n1000 8.92171
R20170 vdd.n1048 vdd.n1047 8.92171
R20171 vdd.n912 vdd.n911 8.92171
R20172 vdd.n959 vdd.n958 8.92171
R20173 vdd.n207 vdd.n117 8.81535
R20174 vdd.n1069 vdd.n979 8.81535
R20175 vdd.n1465 vdd.t16 8.72962
R20176 vdd.t18 vdd.n3042 8.72962
R20177 vdd.n888 vdd.t54 8.50289
R20178 vdd.n1943 vdd.t73 8.50289
R20179 vdd.n516 vdd.t66 8.50289
R20180 vdd.n2874 vdd.t32 8.50289
R20181 vdd.n28 vdd.n14 8.42249
R20182 vdd.n3048 vdd.n3047 8.16225
R20183 vdd.n1161 vdd.n1160 8.16225
R20184 vdd.n272 vdd.n266 8.14595
R20185 vdd.n225 vdd.n219 8.14595
R20186 vdd.n182 vdd.n176 8.14595
R20187 vdd.n135 vdd.n129 8.14595
R20188 vdd.n93 vdd.n87 8.14595
R20189 vdd.n46 vdd.n40 8.14595
R20190 vdd.n1087 vdd.n1081 8.14595
R20191 vdd.n1134 vdd.n1128 8.14595
R20192 vdd.n997 vdd.n991 8.14595
R20193 vdd.n1044 vdd.n1038 8.14595
R20194 vdd.n908 vdd.n902 8.14595
R20195 vdd.n955 vdd.n949 8.14595
R20196 vdd.n2537 vdd.n639 8.11757
R20197 vdd.n2011 vdd.n2010 8.11757
R20198 vdd.n1989 vdd.n833 7.70933
R20199 vdd.n1995 vdd.n833 7.70933
R20200 vdd.n2001 vdd.n827 7.70933
R20201 vdd.n2001 vdd.n820 7.70933
R20202 vdd.n2007 vdd.n820 7.70933
R20203 vdd.n2007 vdd.n823 7.70933
R20204 vdd.n2014 vdd.n808 7.70933
R20205 vdd.n2020 vdd.n808 7.70933
R20206 vdd.n2026 vdd.n802 7.70933
R20207 vdd.n2032 vdd.n798 7.70933
R20208 vdd.n2038 vdd.n792 7.70933
R20209 vdd.n2050 vdd.n779 7.70933
R20210 vdd.n2056 vdd.n773 7.70933
R20211 vdd.n2056 vdd.n766 7.70933
R20212 vdd.n2064 vdd.n766 7.70933
R20213 vdd.n2071 vdd.t189 7.70933
R20214 vdd.n2146 vdd.t189 7.70933
R20215 vdd.n2478 vdd.t195 7.70933
R20216 vdd.n2484 vdd.t195 7.70933
R20217 vdd.n2490 vdd.n687 7.70933
R20218 vdd.n2496 vdd.n687 7.70933
R20219 vdd.n2496 vdd.n690 7.70933
R20220 vdd.n2502 vdd.n683 7.70933
R20221 vdd.n2514 vdd.n670 7.70933
R20222 vdd.n2520 vdd.n664 7.70933
R20223 vdd.n2526 vdd.n660 7.70933
R20224 vdd.n2532 vdd.n647 7.70933
R20225 vdd.n2540 vdd.n647 7.70933
R20226 vdd.n2546 vdd.n641 7.70933
R20227 vdd.n2546 vdd.n633 7.70933
R20228 vdd.n2597 vdd.n633 7.70933
R20229 vdd.n2597 vdd.n636 7.70933
R20230 vdd.n2603 vdd.n595 7.70933
R20231 vdd.n2673 vdd.n595 7.70933
R20232 vdd.n271 vdd.n268 7.3702
R20233 vdd.n224 vdd.n221 7.3702
R20234 vdd.n181 vdd.n178 7.3702
R20235 vdd.n134 vdd.n131 7.3702
R20236 vdd.n92 vdd.n89 7.3702
R20237 vdd.n45 vdd.n42 7.3702
R20238 vdd.n1086 vdd.n1083 7.3702
R20239 vdd.n1133 vdd.n1130 7.3702
R20240 vdd.n996 vdd.n993 7.3702
R20241 vdd.n1043 vdd.n1040 7.3702
R20242 vdd.n907 vdd.n904 7.3702
R20243 vdd.n954 vdd.n951 7.3702
R20244 vdd.n1361 vdd.n1360 6.98232
R20245 vdd.n1653 vdd.n1652 6.98232
R20246 vdd.n2950 vdd.n2949 6.98232
R20247 vdd.n2761 vdd.n2758 6.98232
R20248 vdd.n1498 vdd.t1 6.68904
R20249 vdd.n2857 vdd.t3 6.68904
R20250 vdd.t40 vdd.n887 6.46231
R20251 vdd.n2882 vdd.t7 6.46231
R20252 vdd.n1456 vdd.t22 6.23558
R20253 vdd.t11 vdd.n308 6.23558
R20254 vdd.n3048 vdd.n297 6.22547
R20255 vdd.n1160 vdd.n1159 6.22547
R20256 vdd.n2026 vdd.t145 6.00885
R20257 vdd.n2526 vdd.t185 6.00885
R20258 vdd.n823 vdd.t117 5.89549
R20259 vdd.t81 vdd.n641 5.89549
R20260 vdd.n272 vdd.n271 5.81868
R20261 vdd.n225 vdd.n224 5.81868
R20262 vdd.n182 vdd.n181 5.81868
R20263 vdd.n135 vdd.n134 5.81868
R20264 vdd.n93 vdd.n92 5.81868
R20265 vdd.n46 vdd.n45 5.81868
R20266 vdd.n1087 vdd.n1086 5.81868
R20267 vdd.n1134 vdd.n1133 5.81868
R20268 vdd.n997 vdd.n996 5.81868
R20269 vdd.n1044 vdd.n1043 5.81868
R20270 vdd.n908 vdd.n907 5.81868
R20271 vdd.n955 vdd.n954 5.81868
R20272 vdd.t113 vdd.n827 5.78212
R20273 vdd.n1770 vdd.t98 5.78212
R20274 vdd.n2395 vdd.t106 5.78212
R20275 vdd.n636 vdd.t102 5.78212
R20276 vdd.n2154 vdd.n2153 5.77611
R20277 vdd.n1897 vdd.n1767 5.77611
R20278 vdd.n2408 vdd.n2407 5.77611
R20279 vdd.n2614 vdd.n2613 5.77611
R20280 vdd.n2678 vdd.n591 5.77611
R20281 vdd.n2318 vdd.n2258 5.77611
R20282 vdd.n2079 vdd.n757 5.77611
R20283 vdd.n1827 vdd.n1826 5.77611
R20284 vdd.n1323 vdd.n1322 5.62474
R20285 vdd.n1949 vdd.n1946 5.62474
R20286 vdd.n2910 vdd.n2907 5.62474
R20287 vdd.n2713 vdd.n2710 5.62474
R20288 vdd.t177 vdd.n779 5.44203
R20289 vdd.n683 vdd.t157 5.44203
R20290 vdd.n1180 vdd.t22 5.10193
R20291 vdd.t146 vdd.n802 5.10193
R20292 vdd.n792 vdd.t0 5.10193
R20293 vdd.t153 vdd.n670 5.10193
R20294 vdd.n660 vdd.t182 5.10193
R20295 vdd.n3035 vdd.t11 5.10193
R20296 vdd.n275 vdd.n266 5.04292
R20297 vdd.n228 vdd.n219 5.04292
R20298 vdd.n185 vdd.n176 5.04292
R20299 vdd.n138 vdd.n129 5.04292
R20300 vdd.n96 vdd.n87 5.04292
R20301 vdd.n49 vdd.n40 5.04292
R20302 vdd.n1090 vdd.n1081 5.04292
R20303 vdd.n1137 vdd.n1128 5.04292
R20304 vdd.n1000 vdd.n991 5.04292
R20305 vdd.n1047 vdd.n1038 5.04292
R20306 vdd.n911 vdd.n902 5.04292
R20307 vdd.n958 vdd.n949 5.04292
R20308 vdd.n1473 vdd.t40 4.8752
R20309 vdd.t159 vdd.t149 4.8752
R20310 vdd.t197 vdd.t193 4.8752
R20311 vdd.t143 vdd.t186 4.8752
R20312 vdd.t198 vdd.t156 4.8752
R20313 vdd.t7 vdd.n304 4.8752
R20314 vdd.n2155 vdd.n2154 4.83952
R20315 vdd.n1767 vdd.n1763 4.83952
R20316 vdd.n2409 vdd.n2408 4.83952
R20317 vdd.n2615 vdd.n2614 4.83952
R20318 vdd.n591 vdd.n586 4.83952
R20319 vdd.n2315 vdd.n2258 4.83952
R20320 vdd.n2082 vdd.n757 4.83952
R20321 vdd.n1826 vdd.n1825 4.83952
R20322 vdd.n1621 vdd.n855 4.74817
R20323 vdd.n1616 vdd.n856 4.74817
R20324 vdd.n1518 vdd.n1515 4.74817
R20325 vdd.n1930 vdd.n1519 4.74817
R20326 vdd.n1932 vdd.n1518 4.74817
R20327 vdd.n1931 vdd.n1930 4.74817
R20328 vdd.n2838 vdd.n2837 4.74817
R20329 vdd.n2835 vdd.n2834 4.74817
R20330 vdd.n2835 vdd.n521 4.74817
R20331 vdd.n2837 vdd.n518 4.74817
R20332 vdd.n2720 vdd.n573 4.74817
R20333 vdd.n2716 vdd.n574 4.74817
R20334 vdd.n2719 vdd.n574 4.74817
R20335 vdd.n2723 vdd.n573 4.74817
R20336 vdd.n1617 vdd.n855 4.74817
R20337 vdd.n858 vdd.n856 4.74817
R20338 vdd.n297 vdd.n296 4.7074
R20339 vdd.n207 vdd.n206 4.7074
R20340 vdd.n1159 vdd.n1158 4.7074
R20341 vdd.n1069 vdd.n1068 4.7074
R20342 vdd.n1489 vdd.t1 4.64847
R20343 vdd.n2866 vdd.t3 4.64847
R20344 vdd.n2032 vdd.t151 4.53511
R20345 vdd.n2520 vdd.t187 4.53511
R20346 vdd.n2064 vdd.t183 4.30838
R20347 vdd.n2490 vdd.t180 4.30838
R20348 vdd.n276 vdd.n264 4.26717
R20349 vdd.n229 vdd.n217 4.26717
R20350 vdd.n186 vdd.n174 4.26717
R20351 vdd.n139 vdd.n127 4.26717
R20352 vdd.n97 vdd.n85 4.26717
R20353 vdd.n50 vdd.n38 4.26717
R20354 vdd.n1091 vdd.n1079 4.26717
R20355 vdd.n1138 vdd.n1126 4.26717
R20356 vdd.n1001 vdd.n989 4.26717
R20357 vdd.n1048 vdd.n1036 4.26717
R20358 vdd.n912 vdd.n900 4.26717
R20359 vdd.n959 vdd.n947 4.26717
R20360 vdd.n297 vdd.n207 4.10845
R20361 vdd.n1159 vdd.n1069 4.10845
R20362 vdd.n253 vdd.t48 4.06363
R20363 vdd.n253 vdd.t12 4.06363
R20364 vdd.n251 vdd.t14 4.06363
R20365 vdd.n251 vdd.t35 4.06363
R20366 vdd.n249 vdd.t37 4.06363
R20367 vdd.n249 vdd.t53 4.06363
R20368 vdd.n163 vdd.t43 4.06363
R20369 vdd.n163 vdd.t64 4.06363
R20370 vdd.n161 vdd.t8 4.06363
R20371 vdd.n161 vdd.t27 4.06363
R20372 vdd.n159 vdd.t33 4.06363
R20373 vdd.n159 vdd.t44 4.06363
R20374 vdd.n74 vdd.t49 4.06363
R20375 vdd.n74 vdd.t24 4.06363
R20376 vdd.n72 vdd.t63 4.06363
R20377 vdd.n72 vdd.t19 4.06363
R20378 vdd.n70 vdd.t56 4.06363
R20379 vdd.n70 vdd.t30 4.06363
R20380 vdd.n1111 vdd.t15 4.06363
R20381 vdd.n1111 vdd.t59 4.06363
R20382 vdd.n1113 vdd.t58 4.06363
R20383 vdd.n1113 vdd.t47 4.06363
R20384 vdd.n1115 vdd.t34 4.06363
R20385 vdd.n1115 vdd.t13 4.06363
R20386 vdd.n1021 vdd.t10 4.06363
R20387 vdd.n1021 vdd.t55 4.06363
R20388 vdd.n1023 vdd.t50 4.06363
R20389 vdd.n1023 vdd.t41 4.06363
R20390 vdd.n1025 vdd.t26 4.06363
R20391 vdd.n1025 vdd.t6 4.06363
R20392 vdd.n932 vdd.t28 4.06363
R20393 vdd.n932 vdd.t57 4.06363
R20394 vdd.n934 vdd.t17 4.06363
R20395 vdd.n934 vdd.t45 4.06363
R20396 vdd.n936 vdd.t23 4.06363
R20397 vdd.n936 vdd.t51 4.06363
R20398 vdd.n26 vdd.t164 3.9605
R20399 vdd.n26 vdd.t174 3.9605
R20400 vdd.n23 vdd.t163 3.9605
R20401 vdd.n23 vdd.t165 3.9605
R20402 vdd.n21 vdd.t173 3.9605
R20403 vdd.n21 vdd.t160 3.9605
R20404 vdd.n20 vdd.t167 3.9605
R20405 vdd.n20 vdd.t175 3.9605
R20406 vdd.n15 vdd.t170 3.9605
R20407 vdd.n15 vdd.t171 3.9605
R20408 vdd.n16 vdd.t168 3.9605
R20409 vdd.n16 vdd.t169 3.9605
R20410 vdd.n18 vdd.t172 3.9605
R20411 vdd.n18 vdd.t166 3.9605
R20412 vdd.n25 vdd.t161 3.9605
R20413 vdd.n25 vdd.t162 3.9605
R20414 vdd.n7 vdd.t199 3.61217
R20415 vdd.n7 vdd.t188 3.61217
R20416 vdd.n8 vdd.t144 3.61217
R20417 vdd.n8 vdd.t158 3.61217
R20418 vdd.n10 vdd.t196 3.61217
R20419 vdd.n10 vdd.t181 3.61217
R20420 vdd.n12 vdd.t148 3.61217
R20421 vdd.n12 vdd.t155 3.61217
R20422 vdd.n5 vdd.t192 3.61217
R20423 vdd.n5 vdd.t142 3.61217
R20424 vdd.n3 vdd.t184 3.61217
R20425 vdd.n3 vdd.t190 3.61217
R20426 vdd.n1 vdd.t178 3.61217
R20427 vdd.n1 vdd.t194 3.61217
R20428 vdd.n0 vdd.t152 3.61217
R20429 vdd.n0 vdd.t150 3.61217
R20430 vdd.n280 vdd.n279 3.49141
R20431 vdd.n233 vdd.n232 3.49141
R20432 vdd.n190 vdd.n189 3.49141
R20433 vdd.n143 vdd.n142 3.49141
R20434 vdd.n101 vdd.n100 3.49141
R20435 vdd.n54 vdd.n53 3.49141
R20436 vdd.n1095 vdd.n1094 3.49141
R20437 vdd.n1142 vdd.n1141 3.49141
R20438 vdd.n1005 vdd.n1004 3.49141
R20439 vdd.n1052 vdd.n1051 3.49141
R20440 vdd.n916 vdd.n915 3.49141
R20441 vdd.n963 vdd.n962 3.49141
R20442 vdd.n1770 vdd.t183 3.40145
R20443 vdd.n2218 vdd.t191 3.40145
R20444 vdd.n2471 vdd.t154 3.40145
R20445 vdd.n2395 vdd.t180 3.40145
R20446 vdd.n1871 vdd.t151 3.17472
R20447 vdd.n2374 vdd.t187 3.17472
R20448 vdd.n1490 vdd.t54 2.83463
R20449 vdd.n1508 vdd.t73 2.83463
R20450 vdd.n2849 vdd.t66 2.83463
R20451 vdd.n467 vdd.t32 2.83463
R20452 vdd.n283 vdd.n262 2.71565
R20453 vdd.n236 vdd.n215 2.71565
R20454 vdd.n193 vdd.n172 2.71565
R20455 vdd.n146 vdd.n125 2.71565
R20456 vdd.n104 vdd.n83 2.71565
R20457 vdd.n57 vdd.n36 2.71565
R20458 vdd.n1098 vdd.n1077 2.71565
R20459 vdd.n1145 vdd.n1124 2.71565
R20460 vdd.n1008 vdd.n987 2.71565
R20461 vdd.n1055 vdd.n1034 2.71565
R20462 vdd.n919 vdd.n898 2.71565
R20463 vdd.n966 vdd.n945 2.71565
R20464 vdd.t16 vdd.n1164 2.6079
R20465 vdd.n2020 vdd.t146 2.6079
R20466 vdd.n2044 vdd.t0 2.6079
R20467 vdd.n2508 vdd.t153 2.6079
R20468 vdd.n2532 vdd.t182 2.6079
R20469 vdd.n3043 vdd.t18 2.6079
R20470 vdd.n2538 vdd.n2537 2.49806
R20471 vdd.n2012 vdd.n2011 2.49806
R20472 vdd.n270 vdd.n269 2.4129
R20473 vdd.n223 vdd.n222 2.4129
R20474 vdd.n180 vdd.n179 2.4129
R20475 vdd.n133 vdd.n132 2.4129
R20476 vdd.n91 vdd.n90 2.4129
R20477 vdd.n44 vdd.n43 2.4129
R20478 vdd.n1085 vdd.n1084 2.4129
R20479 vdd.n1132 vdd.n1131 2.4129
R20480 vdd.n995 vdd.n994 2.4129
R20481 vdd.n1042 vdd.n1041 2.4129
R20482 vdd.n906 vdd.n905 2.4129
R20483 vdd.n953 vdd.n952 2.4129
R20484 vdd.n1447 vdd.t38 2.38117
R20485 vdd.n3034 vdd.t20 2.38117
R20486 vdd.n1929 vdd.n1518 2.27742
R20487 vdd.n1930 vdd.n1929 2.27742
R20488 vdd.n2836 vdd.n2835 2.27742
R20489 vdd.n2837 vdd.n2836 2.27742
R20490 vdd.n2707 vdd.n574 2.27742
R20491 vdd.n2707 vdd.n573 2.27742
R20492 vdd.n1952 vdd.n855 2.27742
R20493 vdd.n1952 vdd.n856 2.27742
R20494 vdd.n2044 vdd.t177 2.2678
R20495 vdd.n2508 vdd.t157 2.2678
R20496 vdd.t193 vdd.n773 2.04107
R20497 vdd.n690 vdd.t143 2.04107
R20498 vdd.n284 vdd.n260 1.93989
R20499 vdd.n237 vdd.n213 1.93989
R20500 vdd.n194 vdd.n170 1.93989
R20501 vdd.n147 vdd.n123 1.93989
R20502 vdd.n105 vdd.n81 1.93989
R20503 vdd.n58 vdd.n34 1.93989
R20504 vdd.n1099 vdd.n1075 1.93989
R20505 vdd.n1146 vdd.n1122 1.93989
R20506 vdd.n1009 vdd.n985 1.93989
R20507 vdd.n1056 vdd.n1032 1.93989
R20508 vdd.n920 vdd.n896 1.93989
R20509 vdd.n967 vdd.n943 1.93989
R20510 vdd.n1995 vdd.t113 1.92771
R20511 vdd.n2071 vdd.t98 1.92771
R20512 vdd.n2484 vdd.t106 1.92771
R20513 vdd.n2603 vdd.t102 1.92771
R20514 vdd.n1871 vdd.t145 1.70098
R20515 vdd.n798 vdd.t159 1.70098
R20516 vdd.t156 vdd.n664 1.70098
R20517 vdd.n2374 vdd.t185 1.70098
R20518 vdd.n1455 vdd.t5 1.24752
R20519 vdd.t42 vdd.n3041 1.24752
R20520 vdd.n295 vdd.n255 1.16414
R20521 vdd.n288 vdd.n287 1.16414
R20522 vdd.n248 vdd.n208 1.16414
R20523 vdd.n241 vdd.n240 1.16414
R20524 vdd.n205 vdd.n165 1.16414
R20525 vdd.n198 vdd.n197 1.16414
R20526 vdd.n158 vdd.n118 1.16414
R20527 vdd.n151 vdd.n150 1.16414
R20528 vdd.n116 vdd.n76 1.16414
R20529 vdd.n109 vdd.n108 1.16414
R20530 vdd.n69 vdd.n29 1.16414
R20531 vdd.n62 vdd.n61 1.16414
R20532 vdd.n1110 vdd.n1070 1.16414
R20533 vdd.n1103 vdd.n1102 1.16414
R20534 vdd.n1157 vdd.n1117 1.16414
R20535 vdd.n1150 vdd.n1149 1.16414
R20536 vdd.n1020 vdd.n980 1.16414
R20537 vdd.n1013 vdd.n1012 1.16414
R20538 vdd.n1067 vdd.n1027 1.16414
R20539 vdd.n1060 vdd.n1059 1.16414
R20540 vdd.n931 vdd.n891 1.16414
R20541 vdd.n924 vdd.n923 1.16414
R20542 vdd.n978 vdd.n938 1.16414
R20543 vdd.n971 vdd.n970 1.16414
R20544 vdd.n2038 vdd.t149 1.13415
R20545 vdd.n2514 vdd.t198 1.13415
R20546 vdd.n1481 vdd.t9 1.02079
R20547 vdd.t117 vdd.t176 1.02079
R20548 vdd.t179 vdd.t81 1.02079
R20549 vdd.t29 vdd.n456 1.02079
R20550 vdd.n1326 vdd.n1322 0.970197
R20551 vdd.n1950 vdd.n1949 0.970197
R20552 vdd.n2911 vdd.n2910 0.970197
R20553 vdd.n2715 vdd.n2713 0.970197
R20554 vdd.n2014 vdd.t176 0.794056
R20555 vdd.n2050 vdd.t197 0.794056
R20556 vdd.n2502 vdd.t186 0.794056
R20557 vdd.n2540 vdd.t179 0.794056
R20558 vdd.n1160 vdd.n28 0.74827
R20559 vdd vdd.n3048 0.740437
R20560 vdd.n1430 vdd.t77 0.567326
R20561 vdd.n3026 vdd.t88 0.567326
R20562 vdd.n1940 vdd.n1939 0.537085
R20563 vdd.n2845 vdd.n2844 0.537085
R20564 vdd.n3022 vdd.n3021 0.537085
R20565 vdd.n2904 vdd.n2903 0.537085
R20566 vdd.n2709 vdd.n476 0.537085
R20567 vdd.n1503 vdd.n857 0.537085
R20568 vdd.n1324 vdd.n1189 0.537085
R20569 vdd.n1426 vdd.n1425 0.537085
R20570 vdd.n4 vdd.n2 0.459552
R20571 vdd.n11 vdd.n9 0.459552
R20572 vdd.n293 vdd.n292 0.388379
R20573 vdd.n259 vdd.n257 0.388379
R20574 vdd.n246 vdd.n245 0.388379
R20575 vdd.n212 vdd.n210 0.388379
R20576 vdd.n203 vdd.n202 0.388379
R20577 vdd.n169 vdd.n167 0.388379
R20578 vdd.n156 vdd.n155 0.388379
R20579 vdd.n122 vdd.n120 0.388379
R20580 vdd.n114 vdd.n113 0.388379
R20581 vdd.n80 vdd.n78 0.388379
R20582 vdd.n67 vdd.n66 0.388379
R20583 vdd.n33 vdd.n31 0.388379
R20584 vdd.n1108 vdd.n1107 0.388379
R20585 vdd.n1074 vdd.n1072 0.388379
R20586 vdd.n1155 vdd.n1154 0.388379
R20587 vdd.n1121 vdd.n1119 0.388379
R20588 vdd.n1018 vdd.n1017 0.388379
R20589 vdd.n984 vdd.n982 0.388379
R20590 vdd.n1065 vdd.n1064 0.388379
R20591 vdd.n1031 vdd.n1029 0.388379
R20592 vdd.n929 vdd.n928 0.388379
R20593 vdd.n895 vdd.n893 0.388379
R20594 vdd.n976 vdd.n975 0.388379
R20595 vdd.n942 vdd.n940 0.388379
R20596 vdd.n19 vdd.n17 0.387128
R20597 vdd.n24 vdd.n22 0.387128
R20598 vdd.n6 vdd.n4 0.358259
R20599 vdd.n13 vdd.n11 0.358259
R20600 vdd.n252 vdd.n250 0.358259
R20601 vdd.n254 vdd.n252 0.358259
R20602 vdd.n296 vdd.n254 0.358259
R20603 vdd.n162 vdd.n160 0.358259
R20604 vdd.n164 vdd.n162 0.358259
R20605 vdd.n206 vdd.n164 0.358259
R20606 vdd.n73 vdd.n71 0.358259
R20607 vdd.n75 vdd.n73 0.358259
R20608 vdd.n117 vdd.n75 0.358259
R20609 vdd.n1158 vdd.n1116 0.358259
R20610 vdd.n1116 vdd.n1114 0.358259
R20611 vdd.n1114 vdd.n1112 0.358259
R20612 vdd.n1068 vdd.n1026 0.358259
R20613 vdd.n1026 vdd.n1024 0.358259
R20614 vdd.n1024 vdd.n1022 0.358259
R20615 vdd.n979 vdd.n937 0.358259
R20616 vdd.n937 vdd.n935 0.358259
R20617 vdd.n935 vdd.n933 0.358259
R20618 vdd.n14 vdd.n6 0.334552
R20619 vdd.n14 vdd.n13 0.334552
R20620 vdd.n27 vdd.n19 0.21707
R20621 vdd.n27 vdd.n24 0.21707
R20622 vdd.n294 vdd.n256 0.155672
R20623 vdd.n286 vdd.n256 0.155672
R20624 vdd.n286 vdd.n285 0.155672
R20625 vdd.n285 vdd.n261 0.155672
R20626 vdd.n278 vdd.n261 0.155672
R20627 vdd.n278 vdd.n277 0.155672
R20628 vdd.n277 vdd.n265 0.155672
R20629 vdd.n270 vdd.n265 0.155672
R20630 vdd.n247 vdd.n209 0.155672
R20631 vdd.n239 vdd.n209 0.155672
R20632 vdd.n239 vdd.n238 0.155672
R20633 vdd.n238 vdd.n214 0.155672
R20634 vdd.n231 vdd.n214 0.155672
R20635 vdd.n231 vdd.n230 0.155672
R20636 vdd.n230 vdd.n218 0.155672
R20637 vdd.n223 vdd.n218 0.155672
R20638 vdd.n204 vdd.n166 0.155672
R20639 vdd.n196 vdd.n166 0.155672
R20640 vdd.n196 vdd.n195 0.155672
R20641 vdd.n195 vdd.n171 0.155672
R20642 vdd.n188 vdd.n171 0.155672
R20643 vdd.n188 vdd.n187 0.155672
R20644 vdd.n187 vdd.n175 0.155672
R20645 vdd.n180 vdd.n175 0.155672
R20646 vdd.n157 vdd.n119 0.155672
R20647 vdd.n149 vdd.n119 0.155672
R20648 vdd.n149 vdd.n148 0.155672
R20649 vdd.n148 vdd.n124 0.155672
R20650 vdd.n141 vdd.n124 0.155672
R20651 vdd.n141 vdd.n140 0.155672
R20652 vdd.n140 vdd.n128 0.155672
R20653 vdd.n133 vdd.n128 0.155672
R20654 vdd.n115 vdd.n77 0.155672
R20655 vdd.n107 vdd.n77 0.155672
R20656 vdd.n107 vdd.n106 0.155672
R20657 vdd.n106 vdd.n82 0.155672
R20658 vdd.n99 vdd.n82 0.155672
R20659 vdd.n99 vdd.n98 0.155672
R20660 vdd.n98 vdd.n86 0.155672
R20661 vdd.n91 vdd.n86 0.155672
R20662 vdd.n68 vdd.n30 0.155672
R20663 vdd.n60 vdd.n30 0.155672
R20664 vdd.n60 vdd.n59 0.155672
R20665 vdd.n59 vdd.n35 0.155672
R20666 vdd.n52 vdd.n35 0.155672
R20667 vdd.n52 vdd.n51 0.155672
R20668 vdd.n51 vdd.n39 0.155672
R20669 vdd.n44 vdd.n39 0.155672
R20670 vdd.n1109 vdd.n1071 0.155672
R20671 vdd.n1101 vdd.n1071 0.155672
R20672 vdd.n1101 vdd.n1100 0.155672
R20673 vdd.n1100 vdd.n1076 0.155672
R20674 vdd.n1093 vdd.n1076 0.155672
R20675 vdd.n1093 vdd.n1092 0.155672
R20676 vdd.n1092 vdd.n1080 0.155672
R20677 vdd.n1085 vdd.n1080 0.155672
R20678 vdd.n1156 vdd.n1118 0.155672
R20679 vdd.n1148 vdd.n1118 0.155672
R20680 vdd.n1148 vdd.n1147 0.155672
R20681 vdd.n1147 vdd.n1123 0.155672
R20682 vdd.n1140 vdd.n1123 0.155672
R20683 vdd.n1140 vdd.n1139 0.155672
R20684 vdd.n1139 vdd.n1127 0.155672
R20685 vdd.n1132 vdd.n1127 0.155672
R20686 vdd.n1019 vdd.n981 0.155672
R20687 vdd.n1011 vdd.n981 0.155672
R20688 vdd.n1011 vdd.n1010 0.155672
R20689 vdd.n1010 vdd.n986 0.155672
R20690 vdd.n1003 vdd.n986 0.155672
R20691 vdd.n1003 vdd.n1002 0.155672
R20692 vdd.n1002 vdd.n990 0.155672
R20693 vdd.n995 vdd.n990 0.155672
R20694 vdd.n1066 vdd.n1028 0.155672
R20695 vdd.n1058 vdd.n1028 0.155672
R20696 vdd.n1058 vdd.n1057 0.155672
R20697 vdd.n1057 vdd.n1033 0.155672
R20698 vdd.n1050 vdd.n1033 0.155672
R20699 vdd.n1050 vdd.n1049 0.155672
R20700 vdd.n1049 vdd.n1037 0.155672
R20701 vdd.n1042 vdd.n1037 0.155672
R20702 vdd.n930 vdd.n892 0.155672
R20703 vdd.n922 vdd.n892 0.155672
R20704 vdd.n922 vdd.n921 0.155672
R20705 vdd.n921 vdd.n897 0.155672
R20706 vdd.n914 vdd.n897 0.155672
R20707 vdd.n914 vdd.n913 0.155672
R20708 vdd.n913 vdd.n901 0.155672
R20709 vdd.n906 vdd.n901 0.155672
R20710 vdd.n977 vdd.n939 0.155672
R20711 vdd.n969 vdd.n939 0.155672
R20712 vdd.n969 vdd.n968 0.155672
R20713 vdd.n968 vdd.n944 0.155672
R20714 vdd.n961 vdd.n944 0.155672
R20715 vdd.n961 vdd.n960 0.155672
R20716 vdd.n960 vdd.n948 0.155672
R20717 vdd.n953 vdd.n948 0.155672
R20718 vdd.n1715 vdd.n1520 0.152939
R20719 vdd.n1526 vdd.n1520 0.152939
R20720 vdd.n1527 vdd.n1526 0.152939
R20721 vdd.n1528 vdd.n1527 0.152939
R20722 vdd.n1529 vdd.n1528 0.152939
R20723 vdd.n1533 vdd.n1529 0.152939
R20724 vdd.n1534 vdd.n1533 0.152939
R20725 vdd.n1535 vdd.n1534 0.152939
R20726 vdd.n1536 vdd.n1535 0.152939
R20727 vdd.n1540 vdd.n1536 0.152939
R20728 vdd.n1541 vdd.n1540 0.152939
R20729 vdd.n1542 vdd.n1541 0.152939
R20730 vdd.n1690 vdd.n1542 0.152939
R20731 vdd.n1690 vdd.n1689 0.152939
R20732 vdd.n1689 vdd.n1688 0.152939
R20733 vdd.n1688 vdd.n1548 0.152939
R20734 vdd.n1553 vdd.n1548 0.152939
R20735 vdd.n1554 vdd.n1553 0.152939
R20736 vdd.n1555 vdd.n1554 0.152939
R20737 vdd.n1559 vdd.n1555 0.152939
R20738 vdd.n1560 vdd.n1559 0.152939
R20739 vdd.n1561 vdd.n1560 0.152939
R20740 vdd.n1562 vdd.n1561 0.152939
R20741 vdd.n1566 vdd.n1562 0.152939
R20742 vdd.n1567 vdd.n1566 0.152939
R20743 vdd.n1568 vdd.n1567 0.152939
R20744 vdd.n1569 vdd.n1568 0.152939
R20745 vdd.n1573 vdd.n1569 0.152939
R20746 vdd.n1574 vdd.n1573 0.152939
R20747 vdd.n1575 vdd.n1574 0.152939
R20748 vdd.n1576 vdd.n1575 0.152939
R20749 vdd.n1580 vdd.n1576 0.152939
R20750 vdd.n1581 vdd.n1580 0.152939
R20751 vdd.n1582 vdd.n1581 0.152939
R20752 vdd.n1651 vdd.n1582 0.152939
R20753 vdd.n1651 vdd.n1650 0.152939
R20754 vdd.n1650 vdd.n1649 0.152939
R20755 vdd.n1649 vdd.n1588 0.152939
R20756 vdd.n1593 vdd.n1588 0.152939
R20757 vdd.n1594 vdd.n1593 0.152939
R20758 vdd.n1595 vdd.n1594 0.152939
R20759 vdd.n1599 vdd.n1595 0.152939
R20760 vdd.n1600 vdd.n1599 0.152939
R20761 vdd.n1601 vdd.n1600 0.152939
R20762 vdd.n1602 vdd.n1601 0.152939
R20763 vdd.n1606 vdd.n1602 0.152939
R20764 vdd.n1607 vdd.n1606 0.152939
R20765 vdd.n1608 vdd.n1607 0.152939
R20766 vdd.n1609 vdd.n1608 0.152939
R20767 vdd.n1610 vdd.n1609 0.152939
R20768 vdd.n1610 vdd.n854 0.152939
R20769 vdd.n1939 vdd.n1514 0.152939
R20770 vdd.n1477 vdd.n1476 0.152939
R20771 vdd.n1478 vdd.n1477 0.152939
R20772 vdd.n1478 vdd.n879 0.152939
R20773 vdd.n1493 vdd.n879 0.152939
R20774 vdd.n1494 vdd.n1493 0.152939
R20775 vdd.n1495 vdd.n1494 0.152939
R20776 vdd.n1495 vdd.n867 0.152939
R20777 vdd.n1512 vdd.n867 0.152939
R20778 vdd.n1513 vdd.n1512 0.152939
R20779 vdd.n1940 vdd.n1513 0.152939
R20780 vdd.n524 vdd.n519 0.152939
R20781 vdd.n525 vdd.n524 0.152939
R20782 vdd.n526 vdd.n525 0.152939
R20783 vdd.n527 vdd.n526 0.152939
R20784 vdd.n528 vdd.n527 0.152939
R20785 vdd.n529 vdd.n528 0.152939
R20786 vdd.n530 vdd.n529 0.152939
R20787 vdd.n531 vdd.n530 0.152939
R20788 vdd.n532 vdd.n531 0.152939
R20789 vdd.n533 vdd.n532 0.152939
R20790 vdd.n534 vdd.n533 0.152939
R20791 vdd.n535 vdd.n534 0.152939
R20792 vdd.n2803 vdd.n535 0.152939
R20793 vdd.n2803 vdd.n2802 0.152939
R20794 vdd.n2802 vdd.n2801 0.152939
R20795 vdd.n2801 vdd.n537 0.152939
R20796 vdd.n538 vdd.n537 0.152939
R20797 vdd.n539 vdd.n538 0.152939
R20798 vdd.n540 vdd.n539 0.152939
R20799 vdd.n541 vdd.n540 0.152939
R20800 vdd.n542 vdd.n541 0.152939
R20801 vdd.n543 vdd.n542 0.152939
R20802 vdd.n544 vdd.n543 0.152939
R20803 vdd.n545 vdd.n544 0.152939
R20804 vdd.n546 vdd.n545 0.152939
R20805 vdd.n547 vdd.n546 0.152939
R20806 vdd.n548 vdd.n547 0.152939
R20807 vdd.n549 vdd.n548 0.152939
R20808 vdd.n550 vdd.n549 0.152939
R20809 vdd.n551 vdd.n550 0.152939
R20810 vdd.n552 vdd.n551 0.152939
R20811 vdd.n553 vdd.n552 0.152939
R20812 vdd.n554 vdd.n553 0.152939
R20813 vdd.n555 vdd.n554 0.152939
R20814 vdd.n2757 vdd.n555 0.152939
R20815 vdd.n2757 vdd.n2756 0.152939
R20816 vdd.n2756 vdd.n2755 0.152939
R20817 vdd.n2755 vdd.n559 0.152939
R20818 vdd.n560 vdd.n559 0.152939
R20819 vdd.n561 vdd.n560 0.152939
R20820 vdd.n562 vdd.n561 0.152939
R20821 vdd.n563 vdd.n562 0.152939
R20822 vdd.n564 vdd.n563 0.152939
R20823 vdd.n565 vdd.n564 0.152939
R20824 vdd.n566 vdd.n565 0.152939
R20825 vdd.n567 vdd.n566 0.152939
R20826 vdd.n568 vdd.n567 0.152939
R20827 vdd.n569 vdd.n568 0.152939
R20828 vdd.n570 vdd.n569 0.152939
R20829 vdd.n571 vdd.n570 0.152939
R20830 vdd.n572 vdd.n571 0.152939
R20831 vdd.n2844 vdd.n481 0.152939
R20832 vdd.n2846 vdd.n2845 0.152939
R20833 vdd.n2846 vdd.n470 0.152939
R20834 vdd.n2861 vdd.n470 0.152939
R20835 vdd.n2862 vdd.n2861 0.152939
R20836 vdd.n2863 vdd.n2862 0.152939
R20837 vdd.n2863 vdd.n459 0.152939
R20838 vdd.n2877 vdd.n459 0.152939
R20839 vdd.n2878 vdd.n2877 0.152939
R20840 vdd.n2879 vdd.n2878 0.152939
R20841 vdd.n2879 vdd.n298 0.152939
R20842 vdd.n3046 vdd.n299 0.152939
R20843 vdd.n310 vdd.n299 0.152939
R20844 vdd.n311 vdd.n310 0.152939
R20845 vdd.n312 vdd.n311 0.152939
R20846 vdd.n320 vdd.n312 0.152939
R20847 vdd.n321 vdd.n320 0.152939
R20848 vdd.n322 vdd.n321 0.152939
R20849 vdd.n323 vdd.n322 0.152939
R20850 vdd.n331 vdd.n323 0.152939
R20851 vdd.n3022 vdd.n331 0.152939
R20852 vdd.n3021 vdd.n332 0.152939
R20853 vdd.n335 vdd.n332 0.152939
R20854 vdd.n339 vdd.n335 0.152939
R20855 vdd.n340 vdd.n339 0.152939
R20856 vdd.n341 vdd.n340 0.152939
R20857 vdd.n342 vdd.n341 0.152939
R20858 vdd.n343 vdd.n342 0.152939
R20859 vdd.n347 vdd.n343 0.152939
R20860 vdd.n348 vdd.n347 0.152939
R20861 vdd.n349 vdd.n348 0.152939
R20862 vdd.n350 vdd.n349 0.152939
R20863 vdd.n354 vdd.n350 0.152939
R20864 vdd.n355 vdd.n354 0.152939
R20865 vdd.n356 vdd.n355 0.152939
R20866 vdd.n357 vdd.n356 0.152939
R20867 vdd.n361 vdd.n357 0.152939
R20868 vdd.n362 vdd.n361 0.152939
R20869 vdd.n363 vdd.n362 0.152939
R20870 vdd.n2987 vdd.n363 0.152939
R20871 vdd.n2987 vdd.n2986 0.152939
R20872 vdd.n2986 vdd.n2985 0.152939
R20873 vdd.n2985 vdd.n369 0.152939
R20874 vdd.n374 vdd.n369 0.152939
R20875 vdd.n375 vdd.n374 0.152939
R20876 vdd.n376 vdd.n375 0.152939
R20877 vdd.n380 vdd.n376 0.152939
R20878 vdd.n381 vdd.n380 0.152939
R20879 vdd.n382 vdd.n381 0.152939
R20880 vdd.n383 vdd.n382 0.152939
R20881 vdd.n387 vdd.n383 0.152939
R20882 vdd.n388 vdd.n387 0.152939
R20883 vdd.n389 vdd.n388 0.152939
R20884 vdd.n390 vdd.n389 0.152939
R20885 vdd.n394 vdd.n390 0.152939
R20886 vdd.n395 vdd.n394 0.152939
R20887 vdd.n396 vdd.n395 0.152939
R20888 vdd.n397 vdd.n396 0.152939
R20889 vdd.n401 vdd.n397 0.152939
R20890 vdd.n402 vdd.n401 0.152939
R20891 vdd.n403 vdd.n402 0.152939
R20892 vdd.n2948 vdd.n403 0.152939
R20893 vdd.n2948 vdd.n2947 0.152939
R20894 vdd.n2947 vdd.n2946 0.152939
R20895 vdd.n2946 vdd.n409 0.152939
R20896 vdd.n414 vdd.n409 0.152939
R20897 vdd.n415 vdd.n414 0.152939
R20898 vdd.n416 vdd.n415 0.152939
R20899 vdd.n420 vdd.n416 0.152939
R20900 vdd.n421 vdd.n420 0.152939
R20901 vdd.n422 vdd.n421 0.152939
R20902 vdd.n423 vdd.n422 0.152939
R20903 vdd.n427 vdd.n423 0.152939
R20904 vdd.n428 vdd.n427 0.152939
R20905 vdd.n429 vdd.n428 0.152939
R20906 vdd.n430 vdd.n429 0.152939
R20907 vdd.n434 vdd.n430 0.152939
R20908 vdd.n435 vdd.n434 0.152939
R20909 vdd.n436 vdd.n435 0.152939
R20910 vdd.n437 vdd.n436 0.152939
R20911 vdd.n441 vdd.n437 0.152939
R20912 vdd.n442 vdd.n441 0.152939
R20913 vdd.n443 vdd.n442 0.152939
R20914 vdd.n2904 vdd.n443 0.152939
R20915 vdd.n2852 vdd.n476 0.152939
R20916 vdd.n2853 vdd.n2852 0.152939
R20917 vdd.n2854 vdd.n2853 0.152939
R20918 vdd.n2854 vdd.n464 0.152939
R20919 vdd.n2869 vdd.n464 0.152939
R20920 vdd.n2870 vdd.n2869 0.152939
R20921 vdd.n2871 vdd.n2870 0.152939
R20922 vdd.n2871 vdd.n452 0.152939
R20923 vdd.n2885 vdd.n452 0.152939
R20924 vdd.n2886 vdd.n2885 0.152939
R20925 vdd.n2887 vdd.n2886 0.152939
R20926 vdd.n2887 vdd.n450 0.152939
R20927 vdd.n2891 vdd.n450 0.152939
R20928 vdd.n2892 vdd.n2891 0.152939
R20929 vdd.n2893 vdd.n2892 0.152939
R20930 vdd.n2893 vdd.n447 0.152939
R20931 vdd.n2897 vdd.n447 0.152939
R20932 vdd.n2898 vdd.n2897 0.152939
R20933 vdd.n2899 vdd.n2898 0.152939
R20934 vdd.n2899 vdd.n444 0.152939
R20935 vdd.n2903 vdd.n444 0.152939
R20936 vdd.n2709 vdd.n2708 0.152939
R20937 vdd.n1951 vdd.n857 0.152939
R20938 vdd.n1433 vdd.n1189 0.152939
R20939 vdd.n1434 vdd.n1433 0.152939
R20940 vdd.n1435 vdd.n1434 0.152939
R20941 vdd.n1435 vdd.n1177 0.152939
R20942 vdd.n1450 vdd.n1177 0.152939
R20943 vdd.n1451 vdd.n1450 0.152939
R20944 vdd.n1452 vdd.n1451 0.152939
R20945 vdd.n1452 vdd.n1167 0.152939
R20946 vdd.n1468 vdd.n1167 0.152939
R20947 vdd.n1469 vdd.n1468 0.152939
R20948 vdd.n1470 vdd.n1469 0.152939
R20949 vdd.n1470 vdd.n884 0.152939
R20950 vdd.n1484 vdd.n884 0.152939
R20951 vdd.n1485 vdd.n1484 0.152939
R20952 vdd.n1486 vdd.n1485 0.152939
R20953 vdd.n1486 vdd.n874 0.152939
R20954 vdd.n1501 vdd.n874 0.152939
R20955 vdd.n1502 vdd.n1501 0.152939
R20956 vdd.n1505 vdd.n1502 0.152939
R20957 vdd.n1505 vdd.n1504 0.152939
R20958 vdd.n1504 vdd.n1503 0.152939
R20959 vdd.n1425 vdd.n1194 0.152939
R20960 vdd.n1418 vdd.n1194 0.152939
R20961 vdd.n1418 vdd.n1417 0.152939
R20962 vdd.n1417 vdd.n1416 0.152939
R20963 vdd.n1416 vdd.n1231 0.152939
R20964 vdd.n1412 vdd.n1231 0.152939
R20965 vdd.n1412 vdd.n1411 0.152939
R20966 vdd.n1411 vdd.n1410 0.152939
R20967 vdd.n1410 vdd.n1237 0.152939
R20968 vdd.n1406 vdd.n1237 0.152939
R20969 vdd.n1406 vdd.n1405 0.152939
R20970 vdd.n1405 vdd.n1404 0.152939
R20971 vdd.n1404 vdd.n1243 0.152939
R20972 vdd.n1400 vdd.n1243 0.152939
R20973 vdd.n1400 vdd.n1399 0.152939
R20974 vdd.n1399 vdd.n1398 0.152939
R20975 vdd.n1398 vdd.n1249 0.152939
R20976 vdd.n1394 vdd.n1249 0.152939
R20977 vdd.n1394 vdd.n1393 0.152939
R20978 vdd.n1393 vdd.n1392 0.152939
R20979 vdd.n1392 vdd.n1257 0.152939
R20980 vdd.n1388 vdd.n1257 0.152939
R20981 vdd.n1388 vdd.n1387 0.152939
R20982 vdd.n1387 vdd.n1386 0.152939
R20983 vdd.n1386 vdd.n1263 0.152939
R20984 vdd.n1382 vdd.n1263 0.152939
R20985 vdd.n1382 vdd.n1381 0.152939
R20986 vdd.n1381 vdd.n1380 0.152939
R20987 vdd.n1380 vdd.n1269 0.152939
R20988 vdd.n1376 vdd.n1269 0.152939
R20989 vdd.n1376 vdd.n1375 0.152939
R20990 vdd.n1375 vdd.n1374 0.152939
R20991 vdd.n1374 vdd.n1275 0.152939
R20992 vdd.n1370 vdd.n1275 0.152939
R20993 vdd.n1370 vdd.n1369 0.152939
R20994 vdd.n1369 vdd.n1368 0.152939
R20995 vdd.n1368 vdd.n1281 0.152939
R20996 vdd.n1364 vdd.n1281 0.152939
R20997 vdd.n1364 vdd.n1363 0.152939
R20998 vdd.n1363 vdd.n1362 0.152939
R20999 vdd.n1362 vdd.n1287 0.152939
R21000 vdd.n1355 vdd.n1287 0.152939
R21001 vdd.n1355 vdd.n1354 0.152939
R21002 vdd.n1354 vdd.n1353 0.152939
R21003 vdd.n1353 vdd.n1292 0.152939
R21004 vdd.n1349 vdd.n1292 0.152939
R21005 vdd.n1349 vdd.n1348 0.152939
R21006 vdd.n1348 vdd.n1347 0.152939
R21007 vdd.n1347 vdd.n1298 0.152939
R21008 vdd.n1343 vdd.n1298 0.152939
R21009 vdd.n1343 vdd.n1342 0.152939
R21010 vdd.n1342 vdd.n1341 0.152939
R21011 vdd.n1341 vdd.n1304 0.152939
R21012 vdd.n1337 vdd.n1304 0.152939
R21013 vdd.n1337 vdd.n1336 0.152939
R21014 vdd.n1336 vdd.n1335 0.152939
R21015 vdd.n1335 vdd.n1310 0.152939
R21016 vdd.n1331 vdd.n1310 0.152939
R21017 vdd.n1331 vdd.n1330 0.152939
R21018 vdd.n1330 vdd.n1329 0.152939
R21019 vdd.n1329 vdd.n1316 0.152939
R21020 vdd.n1325 vdd.n1316 0.152939
R21021 vdd.n1325 vdd.n1324 0.152939
R21022 vdd.n1427 vdd.n1426 0.152939
R21023 vdd.n1427 vdd.n1183 0.152939
R21024 vdd.n1442 vdd.n1183 0.152939
R21025 vdd.n1443 vdd.n1442 0.152939
R21026 vdd.n1444 vdd.n1443 0.152939
R21027 vdd.n1444 vdd.n1172 0.152939
R21028 vdd.n1459 vdd.n1172 0.152939
R21029 vdd.n1460 vdd.n1459 0.152939
R21030 vdd.n1462 vdd.n1460 0.152939
R21031 vdd.n1462 vdd.n1461 0.152939
R21032 vdd.n1929 vdd.n1514 0.110256
R21033 vdd.n2836 vdd.n481 0.110256
R21034 vdd.n2708 vdd.n2707 0.110256
R21035 vdd.n1952 vdd.n1951 0.110256
R21036 vdd.n1476 vdd.n1161 0.0695946
R21037 vdd.n3047 vdd.n298 0.0695946
R21038 vdd.n3047 vdd.n3046 0.0695946
R21039 vdd.n1461 vdd.n1161 0.0695946
R21040 vdd.n1929 vdd.n1715 0.0431829
R21041 vdd.n1952 vdd.n854 0.0431829
R21042 vdd.n2836 vdd.n519 0.0431829
R21043 vdd.n2707 vdd.n572 0.0431829
R21044 vdd vdd.n28 0.00833333
R21045 a_n2356_n452.n84 a_n2356_n452.t60 512.366
R21046 a_n2356_n452.n83 a_n2356_n452.t51 512.366
R21047 a_n2356_n452.n82 a_n2356_n452.t45 512.366
R21048 a_n2356_n452.n86 a_n2356_n452.t68 512.366
R21049 a_n2356_n452.n85 a_n2356_n452.t57 512.366
R21050 a_n2356_n452.n81 a_n2356_n452.t56 512.366
R21051 a_n2356_n452.n88 a_n2356_n452.t64 512.366
R21052 a_n2356_n452.n87 a_n2356_n452.t49 512.366
R21053 a_n2356_n452.n80 a_n2356_n452.t50 512.366
R21054 a_n2356_n452.n90 a_n2356_n452.t53 512.366
R21055 a_n2356_n452.n89 a_n2356_n452.t62 512.366
R21056 a_n2356_n452.n79 a_n2356_n452.t44 512.366
R21057 a_n2356_n452.n21 a_n2356_n452.t71 539.01
R21058 a_n2356_n452.n54 a_n2356_n452.t54 512.366
R21059 a_n2356_n452.n53 a_n2356_n452.t58 512.366
R21060 a_n2356_n452.n51 a_n2356_n452.t48 512.366
R21061 a_n2356_n452.n52 a_n2356_n452.t63 512.366
R21062 a_n2356_n452.n17 a_n2356_n452.t8 539.01
R21063 a_n2356_n452.n74 a_n2356_n452.t12 512.366
R21064 a_n2356_n452.n73 a_n2356_n452.t6 512.366
R21065 a_n2356_n452.n47 a_n2356_n452.t4 512.366
R21066 a_n2356_n452.n55 a_n2356_n452.t16 512.366
R21067 a_n2356_n452.n11 a_n2356_n452.t22 539.01
R21068 a_n2356_n452.n95 a_n2356_n452.t14 512.366
R21069 a_n2356_n452.n96 a_n2356_n452.t20 512.366
R21070 a_n2356_n452.n49 a_n2356_n452.t2 512.366
R21071 a_n2356_n452.n97 a_n2356_n452.t10 512.366
R21072 a_n2356_n452.n15 a_n2356_n452.t66 539.01
R21073 a_n2356_n452.n92 a_n2356_n452.t67 512.366
R21074 a_n2356_n452.n93 a_n2356_n452.t46 512.366
R21075 a_n2356_n452.n50 a_n2356_n452.t52 512.366
R21076 a_n2356_n452.n94 a_n2356_n452.t61 512.366
R21077 a_n2356_n452.n0 a_n2356_n452.n45 70.1674
R21078 a_n2356_n452.n2 a_n2356_n452.n43 70.1674
R21079 a_n2356_n452.n4 a_n2356_n452.n41 70.1674
R21080 a_n2356_n452.n6 a_n2356_n452.n39 70.1674
R21081 a_n2356_n452.n30 a_n2356_n452.n19 70.3058
R21082 a_n2356_n452.n26 a_n2356_n452.n22 70.3058
R21083 a_n2356_n452.n22 a_n2356_n452.n46 70.1674
R21084 a_n2356_n452.n20 a_n2356_n452.n28 70.1674
R21085 a_n2356_n452.n28 a_n2356_n452.n51 20.9683
R21086 a_n2356_n452.n27 a_n2356_n452.n20 75.0448
R21087 a_n2356_n452.n53 a_n2356_n452.n27 11.2134
R21088 a_n2356_n452.n18 a_n2356_n452.n21 44.8194
R21089 a_n2356_n452.n46 a_n2356_n452.n47 20.9683
R21090 a_n2356_n452.n31 a_n2356_n452.n22 75.0448
R21091 a_n2356_n452.n73 a_n2356_n452.n31 11.2134
R21092 a_n2356_n452.n16 a_n2356_n452.n17 44.8194
R21093 a_n2356_n452.n8 a_n2356_n452.n37 70.3058
R21094 a_n2356_n452.n12 a_n2356_n452.n34 70.3058
R21095 a_n2356_n452.n33 a_n2356_n452.n13 70.1674
R21096 a_n2356_n452.n33 a_n2356_n452.n50 20.9683
R21097 a_n2356_n452.n13 a_n2356_n452.n32 75.0448
R21098 a_n2356_n452.n93 a_n2356_n452.n32 11.2134
R21099 a_n2356_n452.n14 a_n2356_n452.n15 44.8194
R21100 a_n2356_n452.n36 a_n2356_n452.n9 70.1674
R21101 a_n2356_n452.n36 a_n2356_n452.n49 20.9683
R21102 a_n2356_n452.n9 a_n2356_n452.n35 75.0448
R21103 a_n2356_n452.n96 a_n2356_n452.n35 11.2134
R21104 a_n2356_n452.n10 a_n2356_n452.n11 44.8194
R21105 a_n2356_n452.n39 a_n2356_n452.n79 20.9683
R21106 a_n2356_n452.n38 a_n2356_n452.n7 75.0448
R21107 a_n2356_n452.n89 a_n2356_n452.n38 11.2134
R21108 a_n2356_n452.n7 a_n2356_n452.n90 161.3
R21109 a_n2356_n452.n41 a_n2356_n452.n80 20.9683
R21110 a_n2356_n452.n40 a_n2356_n452.n5 75.0448
R21111 a_n2356_n452.n87 a_n2356_n452.n40 11.2134
R21112 a_n2356_n452.n5 a_n2356_n452.n88 161.3
R21113 a_n2356_n452.n43 a_n2356_n452.n81 20.9683
R21114 a_n2356_n452.n42 a_n2356_n452.n3 75.0448
R21115 a_n2356_n452.n85 a_n2356_n452.n42 11.2134
R21116 a_n2356_n452.n3 a_n2356_n452.n86 161.3
R21117 a_n2356_n452.n45 a_n2356_n452.n82 20.9683
R21118 a_n2356_n452.n44 a_n2356_n452.n1 75.0448
R21119 a_n2356_n452.n83 a_n2356_n452.n44 11.2134
R21120 a_n2356_n452.n1 a_n2356_n452.n84 161.3
R21121 a_n2356_n452.n71 a_n2356_n452.n69 81.4626
R21122 a_n2356_n452.n62 a_n2356_n452.n60 81.4626
R21123 a_n2356_n452.n58 a_n2356_n452.n56 81.4626
R21124 a_n2356_n452.n71 a_n2356_n452.n70 80.9324
R21125 a_n2356_n452.n72 a_n2356_n452.n68 80.9324
R21126 a_n2356_n452.n67 a_n2356_n452.n66 80.9324
R21127 a_n2356_n452.n65 a_n2356_n452.n64 80.9324
R21128 a_n2356_n452.n62 a_n2356_n452.n61 80.9324
R21129 a_n2356_n452.n63 a_n2356_n452.n59 80.9324
R21130 a_n2356_n452.n58 a_n2356_n452.n57 80.9324
R21131 a_n2356_n452.n24 a_n2356_n452.t23 74.6477
R21132 a_n2356_n452.n23 a_n2356_n452.t19 74.6477
R21133 a_n2356_n452.n77 a_n2356_n452.t9 74.2899
R21134 a_n2356_n452.n25 a_n2356_n452.t25 74.2897
R21135 a_n2356_n452.n24 a_n2356_n452.n48 70.6783
R21136 a_n2356_n452.n23 a_n2356_n452.n75 70.6783
R21137 a_n2356_n452.n23 a_n2356_n452.n76 70.6783
R21138 a_n2356_n452.n99 a_n2356_n452.n25 70.6782
R21139 a_n2356_n452.n84 a_n2356_n452.n83 48.2005
R21140 a_n2356_n452.t65 a_n2356_n452.n45 533.335
R21141 a_n2356_n452.n86 a_n2356_n452.n85 48.2005
R21142 a_n2356_n452.t70 a_n2356_n452.n43 533.335
R21143 a_n2356_n452.n88 a_n2356_n452.n87 48.2005
R21144 a_n2356_n452.t59 a_n2356_n452.n41 533.335
R21145 a_n2356_n452.n90 a_n2356_n452.n89 48.2005
R21146 a_n2356_n452.t55 a_n2356_n452.n39 533.335
R21147 a_n2356_n452.n54 a_n2356_n452.n53 48.2005
R21148 a_n2356_n452.n52 a_n2356_n452.n28 20.9683
R21149 a_n2356_n452.n74 a_n2356_n452.n73 48.2005
R21150 a_n2356_n452.n55 a_n2356_n452.n46 20.9683
R21151 a_n2356_n452.n96 a_n2356_n452.n95 48.2005
R21152 a_n2356_n452.n97 a_n2356_n452.n36 20.9683
R21153 a_n2356_n452.n93 a_n2356_n452.n92 48.2005
R21154 a_n2356_n452.n94 a_n2356_n452.n33 20.9683
R21155 a_n2356_n452.n30 a_n2356_n452.t69 533.058
R21156 a_n2356_n452.n26 a_n2356_n452.t18 533.058
R21157 a_n2356_n452.t24 a_n2356_n452.n37 533.058
R21158 a_n2356_n452.t47 a_n2356_n452.n34 533.058
R21159 a_n2356_n452.n65 a_n2356_n452.n63 32.7898
R21160 a_n2356_n452.n44 a_n2356_n452.n82 35.3134
R21161 a_n2356_n452.n42 a_n2356_n452.n81 35.3134
R21162 a_n2356_n452.n40 a_n2356_n452.n80 35.3134
R21163 a_n2356_n452.n38 a_n2356_n452.n79 35.3134
R21164 a_n2356_n452.n27 a_n2356_n452.n51 35.3134
R21165 a_n2356_n452.n31 a_n2356_n452.n47 35.3134
R21166 a_n2356_n452.n49 a_n2356_n452.n35 35.3134
R21167 a_n2356_n452.n50 a_n2356_n452.n32 35.3134
R21168 a_n2356_n452.n22 a_n2356_n452.n72 23.891
R21169 a_n2356_n452.n14 a_n2356_n452.n91 12.046
R21170 a_n2356_n452.n19 a_n2356_n452.n29 11.8414
R21171 a_n2356_n452.n78 a_n2356_n452.n16 10.5365
R21172 a_n2356_n452.n25 a_n2356_n452.n98 9.50122
R21173 a_n2356_n452.n91 a_n2356_n452.n7 7.47588
R21174 a_n2356_n452.n0 a_n2356_n452.n29 7.47588
R21175 a_n2356_n452.n98 a_n2356_n452.n8 6.70126
R21176 a_n2356_n452.n78 a_n2356_n452.n77 5.65783
R21177 a_n2356_n452.n98 a_n2356_n452.n29 5.3452
R21178 a_n2356_n452.n22 a_n2356_n452.n18 3.95126
R21179 a_n2356_n452.n10 a_n2356_n452.n12 3.95126
R21180 a_n2356_n452.n48 a_n2356_n452.t15 3.61217
R21181 a_n2356_n452.n48 a_n2356_n452.t21 3.61217
R21182 a_n2356_n452.n75 a_n2356_n452.t5 3.61217
R21183 a_n2356_n452.n75 a_n2356_n452.t17 3.61217
R21184 a_n2356_n452.n76 a_n2356_n452.t13 3.61217
R21185 a_n2356_n452.n76 a_n2356_n452.t7 3.61217
R21186 a_n2356_n452.t3 a_n2356_n452.n99 3.61217
R21187 a_n2356_n452.n99 a_n2356_n452.t11 3.61217
R21188 a_n2356_n452.n69 a_n2356_n452.t39 2.82907
R21189 a_n2356_n452.n69 a_n2356_n452.t38 2.82907
R21190 a_n2356_n452.n70 a_n2356_n452.t43 2.82907
R21191 a_n2356_n452.n70 a_n2356_n452.t28 2.82907
R21192 a_n2356_n452.n68 a_n2356_n452.t29 2.82907
R21193 a_n2356_n452.n68 a_n2356_n452.t35 2.82907
R21194 a_n2356_n452.n66 a_n2356_n452.t42 2.82907
R21195 a_n2356_n452.n66 a_n2356_n452.t0 2.82907
R21196 a_n2356_n452.n64 a_n2356_n452.t40 2.82907
R21197 a_n2356_n452.n64 a_n2356_n452.t1 2.82907
R21198 a_n2356_n452.n60 a_n2356_n452.t36 2.82907
R21199 a_n2356_n452.n60 a_n2356_n452.t34 2.82907
R21200 a_n2356_n452.n61 a_n2356_n452.t41 2.82907
R21201 a_n2356_n452.n61 a_n2356_n452.t30 2.82907
R21202 a_n2356_n452.n59 a_n2356_n452.t37 2.82907
R21203 a_n2356_n452.n59 a_n2356_n452.t27 2.82907
R21204 a_n2356_n452.n57 a_n2356_n452.t31 2.82907
R21205 a_n2356_n452.n57 a_n2356_n452.t32 2.82907
R21206 a_n2356_n452.n56 a_n2356_n452.t26 2.82907
R21207 a_n2356_n452.n56 a_n2356_n452.t33 2.82907
R21208 a_n2356_n452.n91 a_n2356_n452.n78 1.30542
R21209 a_n2356_n452.n4 a_n2356_n452.n3 1.04595
R21210 a_n2356_n452.n21 a_n2356_n452.n54 13.657
R21211 a_n2356_n452.n52 a_n2356_n452.n30 21.4216
R21212 a_n2356_n452.n17 a_n2356_n452.n74 13.657
R21213 a_n2356_n452.n55 a_n2356_n452.n26 21.4216
R21214 a_n2356_n452.n95 a_n2356_n452.n11 13.657
R21215 a_n2356_n452.n37 a_n2356_n452.n97 21.4216
R21216 a_n2356_n452.n92 a_n2356_n452.n15 13.657
R21217 a_n2356_n452.n34 a_n2356_n452.n94 21.4216
R21218 a_n2356_n452.n22 a_n2356_n452.n16 1.47777
R21219 a_n2356_n452.n20 a_n2356_n452.n18 0.758076
R21220 a_n2356_n452.n20 a_n2356_n452.n19 0.758076
R21221 a_n2356_n452.n14 a_n2356_n452.n13 0.758076
R21222 a_n2356_n452.n13 a_n2356_n452.n12 0.758076
R21223 a_n2356_n452.n10 a_n2356_n452.n9 0.758076
R21224 a_n2356_n452.n9 a_n2356_n452.n8 0.758076
R21225 a_n2356_n452.n7 a_n2356_n452.n6 0.758076
R21226 a_n2356_n452.n5 a_n2356_n452.n4 0.758076
R21227 a_n2356_n452.n3 a_n2356_n452.n2 0.758076
R21228 a_n2356_n452.n1 a_n2356_n452.n0 0.758076
R21229 a_n2356_n452.n25 a_n2356_n452.n24 0.716017
R21230 a_n2356_n452.n77 a_n2356_n452.n23 0.716017
R21231 a_n2356_n452.n6 a_n2356_n452.n5 0.67853
R21232 a_n2356_n452.n2 a_n2356_n452.n1 0.67853
R21233 a_n2356_n452.n63 a_n2356_n452.n58 0.530672
R21234 a_n2356_n452.n63 a_n2356_n452.n62 0.530672
R21235 a_n2356_n452.n67 a_n2356_n452.n65 0.530672
R21236 a_n2356_n452.n72 a_n2356_n452.n67 0.530672
R21237 a_n2356_n452.n72 a_n2356_n452.n71 0.530672
R21238 a_n1808_13878.n5 a_n1808_13878.n3 98.9633
R21239 a_n1808_13878.n2 a_n1808_13878.n0 98.7517
R21240 a_n1808_13878.n2 a_n1808_13878.n1 98.6055
R21241 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R21242 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R21243 a_n1808_13878.n7 a_n1808_13878.n6 98.6054
R21244 a_n1808_13878.n9 a_n1808_13878.t13 74.6477
R21245 a_n1808_13878.n14 a_n1808_13878.t14 74.2899
R21246 a_n1808_13878.n11 a_n1808_13878.t15 74.2899
R21247 a_n1808_13878.n10 a_n1808_13878.t12 74.2899
R21248 a_n1808_13878.n13 a_n1808_13878.n12 70.6783
R21249 a_n1808_13878.n9 a_n1808_13878.n8 70.6783
R21250 a_n1808_13878.n16 a_n1808_13878.n15 13.5694
R21251 a_n1808_13878.n15 a_n1808_13878.n7 11.5762
R21252 a_n1808_13878.n15 a_n1808_13878.n14 6.2408
R21253 a_n1808_13878.n1 a_n1808_13878.t6 3.61217
R21254 a_n1808_13878.n1 a_n1808_13878.t1 3.61217
R21255 a_n1808_13878.n0 a_n1808_13878.t0 3.61217
R21256 a_n1808_13878.n0 a_n1808_13878.t2 3.61217
R21257 a_n1808_13878.n6 a_n1808_13878.t7 3.61217
R21258 a_n1808_13878.n6 a_n1808_13878.t8 3.61217
R21259 a_n1808_13878.n4 a_n1808_13878.t10 3.61217
R21260 a_n1808_13878.n4 a_n1808_13878.t3 3.61217
R21261 a_n1808_13878.n3 a_n1808_13878.t5 3.61217
R21262 a_n1808_13878.n3 a_n1808_13878.t9 3.61217
R21263 a_n1808_13878.n12 a_n1808_13878.t18 3.61217
R21264 a_n1808_13878.n12 a_n1808_13878.t19 3.61217
R21265 a_n1808_13878.n8 a_n1808_13878.t16 3.61217
R21266 a_n1808_13878.n8 a_n1808_13878.t17 3.61217
R21267 a_n1808_13878.n17 a_n1808_13878.t4 3.61217
R21268 a_n1808_13878.t11 a_n1808_13878.n17 3.61217
R21269 a_n1808_13878.n7 a_n1808_13878.n5 0.358259
R21270 a_n1808_13878.n10 a_n1808_13878.n9 0.358259
R21271 a_n1808_13878.n13 a_n1808_13878.n11 0.358259
R21272 a_n1808_13878.n14 a_n1808_13878.n13 0.358259
R21273 a_n1808_13878.n16 a_n1808_13878.n2 0.146627
R21274 a_n1808_13878.n11 a_n1808_13878.n10 0.101793
R21275 plus.n61 plus.t11 251.488
R21276 plus.n12 plus.t14 251.488
R21277 plus.n100 plus.t1 243.97
R21278 plus.n96 plus.t23 231.093
R21279 plus.n47 plus.t6 231.093
R21280 plus.n100 plus.n99 223.454
R21281 plus.n102 plus.n101 223.454
R21282 plus.n60 plus.t5 187.445
R21283 plus.n65 plus.t21 187.445
R21284 plus.n71 plus.t20 187.445
R21285 plus.n56 plus.t16 187.445
R21286 plus.n54 plus.t17 187.445
R21287 plus.n83 plus.t13 187.445
R21288 plus.n89 plus.t15 187.445
R21289 plus.n50 plus.t10 187.445
R21290 plus.n1 plus.t12 187.445
R21291 plus.n40 plus.t8 187.445
R21292 plus.n34 plus.t7 187.445
R21293 plus.n5 plus.t19 187.445
R21294 plus.n7 plus.t18 187.445
R21295 plus.n22 plus.t24 187.445
R21296 plus.n16 plus.t22 187.445
R21297 plus.n11 plus.t9 187.445
R21298 plus.n97 plus.n96 161.3
R21299 plus.n95 plus.n49 161.3
R21300 plus.n94 plus.n93 161.3
R21301 plus.n92 plus.n91 161.3
R21302 plus.n90 plus.n51 161.3
R21303 plus.n88 plus.n87 161.3
R21304 plus.n86 plus.n52 161.3
R21305 plus.n85 plus.n84 161.3
R21306 plus.n82 plus.n53 161.3
R21307 plus.n81 plus.n80 161.3
R21308 plus.n79 plus.n78 161.3
R21309 plus.n77 plus.n55 161.3
R21310 plus.n76 plus.n75 161.3
R21311 plus.n74 plus.n73 161.3
R21312 plus.n72 plus.n57 161.3
R21313 plus.n70 plus.n69 161.3
R21314 plus.n68 plus.n58 161.3
R21315 plus.n67 plus.n66 161.3
R21316 plus.n64 plus.n59 161.3
R21317 plus.n63 plus.n62 161.3
R21318 plus.n14 plus.n13 161.3
R21319 plus.n15 plus.n10 161.3
R21320 plus.n18 plus.n17 161.3
R21321 plus.n19 plus.n9 161.3
R21322 plus.n21 plus.n20 161.3
R21323 plus.n23 plus.n8 161.3
R21324 plus.n25 plus.n24 161.3
R21325 plus.n27 plus.n26 161.3
R21326 plus.n28 plus.n6 161.3
R21327 plus.n30 plus.n29 161.3
R21328 plus.n32 plus.n31 161.3
R21329 plus.n33 plus.n4 161.3
R21330 plus.n36 plus.n35 161.3
R21331 plus.n37 plus.n3 161.3
R21332 plus.n39 plus.n38 161.3
R21333 plus.n41 plus.n2 161.3
R21334 plus.n43 plus.n42 161.3
R21335 plus.n45 plus.n44 161.3
R21336 plus.n46 plus.n0 161.3
R21337 plus.n48 plus.n47 161.3
R21338 plus.n64 plus.n63 56.5617
R21339 plus.n91 plus.n90 56.5617
R21340 plus.n42 plus.n41 56.5617
R21341 plus.n15 plus.n14 56.5617
R21342 plus.n73 plus.n72 56.5617
R21343 plus.n82 plus.n81 56.5617
R21344 plus.n33 plus.n32 56.5617
R21345 plus.n24 plus.n23 56.5617
R21346 plus.n95 plus.n94 48.3272
R21347 plus.n46 plus.n45 48.3272
R21348 plus.n70 plus.n58 44.4521
R21349 plus.n84 plus.n52 44.4521
R21350 plus.n35 plus.n3 44.4521
R21351 plus.n21 plus.n9 44.4521
R21352 plus.n62 plus.n61 43.0014
R21353 plus.n13 plus.n12 43.0014
R21354 plus.n77 plus.n76 40.577
R21355 plus.n78 plus.n77 40.577
R21356 plus.n29 plus.n28 40.577
R21357 plus.n28 plus.n27 40.577
R21358 plus.n61 plus.n60 39.4345
R21359 plus.n12 plus.n11 39.4345
R21360 plus.n66 plus.n58 36.702
R21361 plus.n88 plus.n52 36.702
R21362 plus.n39 plus.n3 36.702
R21363 plus.n17 plus.n9 36.702
R21364 plus.n98 plus.n97 33.3471
R21365 plus.n65 plus.n64 20.9036
R21366 plus.n90 plus.n89 20.9036
R21367 plus.n41 plus.n40 20.9036
R21368 plus.n16 plus.n15 20.9036
R21369 plus.n99 plus.t2 19.8005
R21370 plus.n99 plus.t4 19.8005
R21371 plus.n101 plus.t0 19.8005
R21372 plus.n101 plus.t3 19.8005
R21373 plus.n73 plus.n56 18.9362
R21374 plus.n81 plus.n54 18.9362
R21375 plus.n32 plus.n5 18.9362
R21376 plus.n24 plus.n7 18.9362
R21377 plus.n72 plus.n71 16.9689
R21378 plus.n83 plus.n82 16.9689
R21379 plus.n34 plus.n33 16.9689
R21380 plus.n23 plus.n22 16.9689
R21381 plus.n63 plus.n60 15.0015
R21382 plus.n91 plus.n50 15.0015
R21383 plus.n42 plus.n1 15.0015
R21384 plus.n14 plus.n11 15.0015
R21385 plus plus.n103 14.5821
R21386 plus.n96 plus.n95 12.4157
R21387 plus.n47 plus.n46 12.4157
R21388 plus.n98 plus.n48 11.9418
R21389 plus.n94 plus.n50 9.59132
R21390 plus.n45 plus.n1 9.59132
R21391 plus.n71 plus.n70 7.62397
R21392 plus.n84 plus.n83 7.62397
R21393 plus.n35 plus.n34 7.62397
R21394 plus.n22 plus.n21 7.62397
R21395 plus.n76 plus.n56 5.65662
R21396 plus.n78 plus.n54 5.65662
R21397 plus.n29 plus.n5 5.65662
R21398 plus.n27 plus.n7 5.65662
R21399 plus.n103 plus.n102 5.40567
R21400 plus.n66 plus.n65 3.68928
R21401 plus.n89 plus.n88 3.68928
R21402 plus.n40 plus.n39 3.68928
R21403 plus.n17 plus.n16 3.68928
R21404 plus.n103 plus.n98 1.188
R21405 plus.n102 plus.n100 0.716017
R21406 plus.n62 plus.n59 0.189894
R21407 plus.n67 plus.n59 0.189894
R21408 plus.n68 plus.n67 0.189894
R21409 plus.n69 plus.n68 0.189894
R21410 plus.n69 plus.n57 0.189894
R21411 plus.n74 plus.n57 0.189894
R21412 plus.n75 plus.n74 0.189894
R21413 plus.n75 plus.n55 0.189894
R21414 plus.n79 plus.n55 0.189894
R21415 plus.n80 plus.n79 0.189894
R21416 plus.n80 plus.n53 0.189894
R21417 plus.n85 plus.n53 0.189894
R21418 plus.n86 plus.n85 0.189894
R21419 plus.n87 plus.n86 0.189894
R21420 plus.n87 plus.n51 0.189894
R21421 plus.n92 plus.n51 0.189894
R21422 plus.n93 plus.n92 0.189894
R21423 plus.n93 plus.n49 0.189894
R21424 plus.n97 plus.n49 0.189894
R21425 plus.n48 plus.n0 0.189894
R21426 plus.n44 plus.n0 0.189894
R21427 plus.n44 plus.n43 0.189894
R21428 plus.n43 plus.n2 0.189894
R21429 plus.n38 plus.n2 0.189894
R21430 plus.n38 plus.n37 0.189894
R21431 plus.n37 plus.n36 0.189894
R21432 plus.n36 plus.n4 0.189894
R21433 plus.n31 plus.n4 0.189894
R21434 plus.n31 plus.n30 0.189894
R21435 plus.n30 plus.n6 0.189894
R21436 plus.n26 plus.n6 0.189894
R21437 plus.n26 plus.n25 0.189894
R21438 plus.n25 plus.n8 0.189894
R21439 plus.n20 plus.n8 0.189894
R21440 plus.n20 plus.n19 0.189894
R21441 plus.n19 plus.n18 0.189894
R21442 plus.n18 plus.n10 0.189894
R21443 plus.n13 plus.n10 0.189894
R21444 a_n2903_n3924.n18 a_n2903_n3924.t47 214.624
R21445 a_n2903_n3924.n1 a_n2903_n3924.t4 214.321
R21446 a_n2903_n3924.n12 a_n2903_n3924.t0 214.321
R21447 a_n2903_n3924.n13 a_n2903_n3924.t33 214.321
R21448 a_n2903_n3924.n14 a_n2903_n3924.t29 214.321
R21449 a_n2903_n3924.n15 a_n2903_n3924.t1 214.321
R21450 a_n2903_n3924.n16 a_n2903_n3924.t30 214.321
R21451 a_n2903_n3924.n17 a_n2903_n3924.t46 214.321
R21452 a_n2903_n3924.n0 a_n2903_n3924.t20 55.8337
R21453 a_n2903_n3924.n2 a_n2903_n3924.t40 55.8337
R21454 a_n2903_n3924.n11 a_n2903_n3924.t42 55.8337
R21455 a_n2903_n3924.n41 a_n2903_n3924.t8 55.8335
R21456 a_n2903_n3924.n39 a_n2903_n3924.t36 55.8335
R21457 a_n2903_n3924.n30 a_n2903_n3924.t5 55.8335
R21458 a_n2903_n3924.n29 a_n2903_n3924.t17 55.8335
R21459 a_n2903_n3924.n20 a_n2903_n3924.t25 55.8335
R21460 a_n2903_n3924.n43 a_n2903_n3924.n42 53.0052
R21461 a_n2903_n3924.n45 a_n2903_n3924.n44 53.0052
R21462 a_n2903_n3924.n47 a_n2903_n3924.n46 53.0052
R21463 a_n2903_n3924.n4 a_n2903_n3924.n3 53.0052
R21464 a_n2903_n3924.n6 a_n2903_n3924.n5 53.0052
R21465 a_n2903_n3924.n8 a_n2903_n3924.n7 53.0052
R21466 a_n2903_n3924.n10 a_n2903_n3924.n9 53.0052
R21467 a_n2903_n3924.n38 a_n2903_n3924.n37 53.0051
R21468 a_n2903_n3924.n36 a_n2903_n3924.n35 53.0051
R21469 a_n2903_n3924.n34 a_n2903_n3924.n33 53.0051
R21470 a_n2903_n3924.n32 a_n2903_n3924.n31 53.0051
R21471 a_n2903_n3924.n28 a_n2903_n3924.n27 53.0051
R21472 a_n2903_n3924.n26 a_n2903_n3924.n25 53.0051
R21473 a_n2903_n3924.n24 a_n2903_n3924.n23 53.0051
R21474 a_n2903_n3924.n22 a_n2903_n3924.n21 53.0051
R21475 a_n2903_n3924.n49 a_n2903_n3924.n48 53.0051
R21476 a_n2903_n3924.n19 a_n2903_n3924.n11 12.2417
R21477 a_n2903_n3924.n41 a_n2903_n3924.n40 12.2417
R21478 a_n2903_n3924.n20 a_n2903_n3924.n19 5.16214
R21479 a_n2903_n3924.n40 a_n2903_n3924.n39 5.16214
R21480 a_n2903_n3924.n42 a_n2903_n3924.t16 2.82907
R21481 a_n2903_n3924.n42 a_n2903_n3924.t21 2.82907
R21482 a_n2903_n3924.n44 a_n2903_n3924.t14 2.82907
R21483 a_n2903_n3924.n44 a_n2903_n3924.t18 2.82907
R21484 a_n2903_n3924.n46 a_n2903_n3924.t11 2.82907
R21485 a_n2903_n3924.n46 a_n2903_n3924.t15 2.82907
R21486 a_n2903_n3924.n3 a_n2903_n3924.t27 2.82907
R21487 a_n2903_n3924.n3 a_n2903_n3924.t41 2.82907
R21488 a_n2903_n3924.n5 a_n2903_n3924.t37 2.82907
R21489 a_n2903_n3924.n5 a_n2903_n3924.t45 2.82907
R21490 a_n2903_n3924.n7 a_n2903_n3924.t2 2.82907
R21491 a_n2903_n3924.n7 a_n2903_n3924.t28 2.82907
R21492 a_n2903_n3924.n9 a_n2903_n3924.t3 2.82907
R21493 a_n2903_n3924.n9 a_n2903_n3924.t44 2.82907
R21494 a_n2903_n3924.n37 a_n2903_n3924.t31 2.82907
R21495 a_n2903_n3924.n37 a_n2903_n3924.t38 2.82907
R21496 a_n2903_n3924.n35 a_n2903_n3924.t6 2.82907
R21497 a_n2903_n3924.n35 a_n2903_n3924.t43 2.82907
R21498 a_n2903_n3924.n33 a_n2903_n3924.t34 2.82907
R21499 a_n2903_n3924.n33 a_n2903_n3924.t39 2.82907
R21500 a_n2903_n3924.n31 a_n2903_n3924.t35 2.82907
R21501 a_n2903_n3924.n31 a_n2903_n3924.t32 2.82907
R21502 a_n2903_n3924.n27 a_n2903_n3924.t9 2.82907
R21503 a_n2903_n3924.n27 a_n2903_n3924.t22 2.82907
R21504 a_n2903_n3924.n25 a_n2903_n3924.t13 2.82907
R21505 a_n2903_n3924.n25 a_n2903_n3924.t7 2.82907
R21506 a_n2903_n3924.n23 a_n2903_n3924.t24 2.82907
R21507 a_n2903_n3924.n23 a_n2903_n3924.t12 2.82907
R21508 a_n2903_n3924.n21 a_n2903_n3924.t19 2.82907
R21509 a_n2903_n3924.n21 a_n2903_n3924.t23 2.82907
R21510 a_n2903_n3924.t26 a_n2903_n3924.n49 2.82907
R21511 a_n2903_n3924.n49 a_n2903_n3924.t10 2.82907
R21512 a_n2903_n3924.n40 a_n2903_n3924.n1 2.18441
R21513 a_n2903_n3924.n19 a_n2903_n3924.n18 1.95694
R21514 a_n2903_n3924.n17 a_n2903_n3924.n16 0.672012
R21515 a_n2903_n3924.n16 a_n2903_n3924.n15 0.672012
R21516 a_n2903_n3924.n15 a_n2903_n3924.n14 0.672012
R21517 a_n2903_n3924.n14 a_n2903_n3924.n13 0.672012
R21518 a_n2903_n3924.n13 a_n2903_n3924.n12 0.672012
R21519 a_n2903_n3924.n12 a_n2903_n3924.n1 0.672012
R21520 a_n2903_n3924.n22 a_n2903_n3924.n20 0.530672
R21521 a_n2903_n3924.n24 a_n2903_n3924.n22 0.530672
R21522 a_n2903_n3924.n26 a_n2903_n3924.n24 0.530672
R21523 a_n2903_n3924.n28 a_n2903_n3924.n26 0.530672
R21524 a_n2903_n3924.n29 a_n2903_n3924.n28 0.530672
R21525 a_n2903_n3924.n32 a_n2903_n3924.n30 0.530672
R21526 a_n2903_n3924.n34 a_n2903_n3924.n32 0.530672
R21527 a_n2903_n3924.n36 a_n2903_n3924.n34 0.530672
R21528 a_n2903_n3924.n38 a_n2903_n3924.n36 0.530672
R21529 a_n2903_n3924.n39 a_n2903_n3924.n38 0.530672
R21530 a_n2903_n3924.n11 a_n2903_n3924.n10 0.530672
R21531 a_n2903_n3924.n10 a_n2903_n3924.n8 0.530672
R21532 a_n2903_n3924.n8 a_n2903_n3924.n6 0.530672
R21533 a_n2903_n3924.n6 a_n2903_n3924.n4 0.530672
R21534 a_n2903_n3924.n4 a_n2903_n3924.n2 0.530672
R21535 a_n2903_n3924.n48 a_n2903_n3924.n0 0.530672
R21536 a_n2903_n3924.n48 a_n2903_n3924.n47 0.530672
R21537 a_n2903_n3924.n47 a_n2903_n3924.n45 0.530672
R21538 a_n2903_n3924.n45 a_n2903_n3924.n43 0.530672
R21539 a_n2903_n3924.n43 a_n2903_n3924.n41 0.530672
R21540 a_n2903_n3924.n18 a_n2903_n3924.n17 0.370413
R21541 a_n2903_n3924.n30 a_n2903_n3924.n29 0.235414
R21542 a_n2903_n3924.n2 a_n2903_n3924.n0 0.235414
R21543 output.n41 output.n15 289.615
R21544 output.n72 output.n46 289.615
R21545 output.n104 output.n78 289.615
R21546 output.n136 output.n110 289.615
R21547 output.n77 output.n45 197.26
R21548 output.n77 output.n76 196.298
R21549 output.n109 output.n108 196.298
R21550 output.n141 output.n140 196.298
R21551 output.n42 output.n41 185
R21552 output.n40 output.n39 185
R21553 output.n19 output.n18 185
R21554 output.n34 output.n33 185
R21555 output.n32 output.n31 185
R21556 output.n23 output.n22 185
R21557 output.n26 output.n25 185
R21558 output.n73 output.n72 185
R21559 output.n71 output.n70 185
R21560 output.n50 output.n49 185
R21561 output.n65 output.n64 185
R21562 output.n63 output.n62 185
R21563 output.n54 output.n53 185
R21564 output.n57 output.n56 185
R21565 output.n105 output.n104 185
R21566 output.n103 output.n102 185
R21567 output.n82 output.n81 185
R21568 output.n97 output.n96 185
R21569 output.n95 output.n94 185
R21570 output.n86 output.n85 185
R21571 output.n89 output.n88 185
R21572 output.n137 output.n136 185
R21573 output.n135 output.n134 185
R21574 output.n114 output.n113 185
R21575 output.n129 output.n128 185
R21576 output.n127 output.n126 185
R21577 output.n118 output.n117 185
R21578 output.n121 output.n120 185
R21579 output.t1 output.n24 147.661
R21580 output.t2 output.n55 147.661
R21581 output.t19 output.n87 147.661
R21582 output.t0 output.n119 147.661
R21583 output.n41 output.n40 104.615
R21584 output.n40 output.n18 104.615
R21585 output.n33 output.n18 104.615
R21586 output.n33 output.n32 104.615
R21587 output.n32 output.n22 104.615
R21588 output.n25 output.n22 104.615
R21589 output.n72 output.n71 104.615
R21590 output.n71 output.n49 104.615
R21591 output.n64 output.n49 104.615
R21592 output.n64 output.n63 104.615
R21593 output.n63 output.n53 104.615
R21594 output.n56 output.n53 104.615
R21595 output.n104 output.n103 104.615
R21596 output.n103 output.n81 104.615
R21597 output.n96 output.n81 104.615
R21598 output.n96 output.n95 104.615
R21599 output.n95 output.n85 104.615
R21600 output.n88 output.n85 104.615
R21601 output.n136 output.n135 104.615
R21602 output.n135 output.n113 104.615
R21603 output.n128 output.n113 104.615
R21604 output.n128 output.n127 104.615
R21605 output.n127 output.n117 104.615
R21606 output.n120 output.n117 104.615
R21607 output.n1 output.t6 77.056
R21608 output.n14 output.t7 76.6694
R21609 output.n1 output.n0 72.7095
R21610 output.n3 output.n2 72.7095
R21611 output.n5 output.n4 72.7095
R21612 output.n7 output.n6 72.7095
R21613 output.n9 output.n8 72.7095
R21614 output.n11 output.n10 72.7095
R21615 output.n13 output.n12 72.7095
R21616 output.n25 output.t1 52.3082
R21617 output.n56 output.t2 52.3082
R21618 output.n88 output.t19 52.3082
R21619 output.n120 output.t0 52.3082
R21620 output.n26 output.n24 15.6674
R21621 output.n57 output.n55 15.6674
R21622 output.n89 output.n87 15.6674
R21623 output.n121 output.n119 15.6674
R21624 output.n27 output.n23 12.8005
R21625 output.n58 output.n54 12.8005
R21626 output.n90 output.n86 12.8005
R21627 output.n122 output.n118 12.8005
R21628 output.n31 output.n30 12.0247
R21629 output.n62 output.n61 12.0247
R21630 output.n94 output.n93 12.0247
R21631 output.n126 output.n125 12.0247
R21632 output.n34 output.n21 11.249
R21633 output.n65 output.n52 11.249
R21634 output.n97 output.n84 11.249
R21635 output.n129 output.n116 11.249
R21636 output.n35 output.n19 10.4732
R21637 output.n66 output.n50 10.4732
R21638 output.n98 output.n82 10.4732
R21639 output.n130 output.n114 10.4732
R21640 output.n39 output.n38 9.69747
R21641 output.n70 output.n69 9.69747
R21642 output.n102 output.n101 9.69747
R21643 output.n134 output.n133 9.69747
R21644 output.n45 output.n44 9.45567
R21645 output.n76 output.n75 9.45567
R21646 output.n108 output.n107 9.45567
R21647 output.n140 output.n139 9.45567
R21648 output.n44 output.n43 9.3005
R21649 output.n17 output.n16 9.3005
R21650 output.n38 output.n37 9.3005
R21651 output.n36 output.n35 9.3005
R21652 output.n21 output.n20 9.3005
R21653 output.n30 output.n29 9.3005
R21654 output.n28 output.n27 9.3005
R21655 output.n75 output.n74 9.3005
R21656 output.n48 output.n47 9.3005
R21657 output.n69 output.n68 9.3005
R21658 output.n67 output.n66 9.3005
R21659 output.n52 output.n51 9.3005
R21660 output.n61 output.n60 9.3005
R21661 output.n59 output.n58 9.3005
R21662 output.n107 output.n106 9.3005
R21663 output.n80 output.n79 9.3005
R21664 output.n101 output.n100 9.3005
R21665 output.n99 output.n98 9.3005
R21666 output.n84 output.n83 9.3005
R21667 output.n93 output.n92 9.3005
R21668 output.n91 output.n90 9.3005
R21669 output.n139 output.n138 9.3005
R21670 output.n112 output.n111 9.3005
R21671 output.n133 output.n132 9.3005
R21672 output.n131 output.n130 9.3005
R21673 output.n116 output.n115 9.3005
R21674 output.n125 output.n124 9.3005
R21675 output.n123 output.n122 9.3005
R21676 output.n42 output.n17 8.92171
R21677 output.n73 output.n48 8.92171
R21678 output.n105 output.n80 8.92171
R21679 output.n137 output.n112 8.92171
R21680 output output.n141 8.15037
R21681 output.n43 output.n15 8.14595
R21682 output.n74 output.n46 8.14595
R21683 output.n106 output.n78 8.14595
R21684 output.n138 output.n110 8.14595
R21685 output.n45 output.n15 5.81868
R21686 output.n76 output.n46 5.81868
R21687 output.n108 output.n78 5.81868
R21688 output.n140 output.n110 5.81868
R21689 output.n43 output.n42 5.04292
R21690 output.n74 output.n73 5.04292
R21691 output.n106 output.n105 5.04292
R21692 output.n138 output.n137 5.04292
R21693 output.n28 output.n24 4.38594
R21694 output.n59 output.n55 4.38594
R21695 output.n91 output.n87 4.38594
R21696 output.n123 output.n119 4.38594
R21697 output.n39 output.n17 4.26717
R21698 output.n70 output.n48 4.26717
R21699 output.n102 output.n80 4.26717
R21700 output.n134 output.n112 4.26717
R21701 output.n0 output.t11 3.9605
R21702 output.n0 output.t16 3.9605
R21703 output.n2 output.t4 3.9605
R21704 output.n2 output.t12 3.9605
R21705 output.n4 output.t15 3.9605
R21706 output.n4 output.t13 3.9605
R21707 output.n6 output.t3 3.9605
R21708 output.n6 output.t5 3.9605
R21709 output.n8 output.t8 3.9605
R21710 output.n8 output.t17 3.9605
R21711 output.n10 output.t18 3.9605
R21712 output.n10 output.t9 3.9605
R21713 output.n12 output.t10 3.9605
R21714 output.n12 output.t14 3.9605
R21715 output.n38 output.n19 3.49141
R21716 output.n69 output.n50 3.49141
R21717 output.n101 output.n82 3.49141
R21718 output.n133 output.n114 3.49141
R21719 output.n35 output.n34 2.71565
R21720 output.n66 output.n65 2.71565
R21721 output.n98 output.n97 2.71565
R21722 output.n130 output.n129 2.71565
R21723 output.n31 output.n21 1.93989
R21724 output.n62 output.n52 1.93989
R21725 output.n94 output.n84 1.93989
R21726 output.n126 output.n116 1.93989
R21727 output.n30 output.n23 1.16414
R21728 output.n61 output.n54 1.16414
R21729 output.n93 output.n86 1.16414
R21730 output.n125 output.n118 1.16414
R21731 output.n141 output.n109 0.962709
R21732 output.n109 output.n77 0.962709
R21733 output.n27 output.n26 0.388379
R21734 output.n58 output.n57 0.388379
R21735 output.n90 output.n89 0.388379
R21736 output.n122 output.n121 0.388379
R21737 output.n14 output.n13 0.387128
R21738 output.n13 output.n11 0.387128
R21739 output.n11 output.n9 0.387128
R21740 output.n9 output.n7 0.387128
R21741 output.n7 output.n5 0.387128
R21742 output.n5 output.n3 0.387128
R21743 output.n3 output.n1 0.387128
R21744 output.n44 output.n16 0.155672
R21745 output.n37 output.n16 0.155672
R21746 output.n37 output.n36 0.155672
R21747 output.n36 output.n20 0.155672
R21748 output.n29 output.n20 0.155672
R21749 output.n29 output.n28 0.155672
R21750 output.n75 output.n47 0.155672
R21751 output.n68 output.n47 0.155672
R21752 output.n68 output.n67 0.155672
R21753 output.n67 output.n51 0.155672
R21754 output.n60 output.n51 0.155672
R21755 output.n60 output.n59 0.155672
R21756 output.n107 output.n79 0.155672
R21757 output.n100 output.n79 0.155672
R21758 output.n100 output.n99 0.155672
R21759 output.n99 output.n83 0.155672
R21760 output.n92 output.n83 0.155672
R21761 output.n92 output.n91 0.155672
R21762 output.n139 output.n111 0.155672
R21763 output.n132 output.n111 0.155672
R21764 output.n132 output.n131 0.155672
R21765 output.n131 output.n115 0.155672
R21766 output.n124 output.n115 0.155672
R21767 output.n124 output.n123 0.155672
R21768 output output.n14 0.126227
R21769 minus.n61 minus.t24 251.488
R21770 minus.n12 minus.t16 251.488
R21771 minus.n102 minus.t4 243.255
R21772 minus.n96 minus.t14 231.093
R21773 minus.n47 minus.t9 231.093
R21774 minus.n101 minus.n99 224.169
R21775 minus.n101 minus.n100 223.454
R21776 minus.n50 minus.t21 187.445
R21777 minus.n89 minus.t18 187.445
R21778 minus.n83 minus.t15 187.445
R21779 minus.n54 minus.t7 187.445
R21780 minus.n56 minus.t6 187.445
R21781 minus.n71 minus.t12 187.445
R21782 minus.n65 minus.t11 187.445
R21783 minus.n60 minus.t19 187.445
R21784 minus.n11 minus.t10 187.445
R21785 minus.n16 minus.t8 187.445
R21786 minus.n22 minus.t5 187.445
R21787 minus.n7 minus.t22 187.445
R21788 minus.n5 minus.t23 187.445
R21789 minus.n34 minus.t17 187.445
R21790 minus.n40 minus.t20 187.445
R21791 minus.n1 minus.t13 187.445
R21792 minus.n63 minus.n62 161.3
R21793 minus.n64 minus.n59 161.3
R21794 minus.n67 minus.n66 161.3
R21795 minus.n68 minus.n58 161.3
R21796 minus.n70 minus.n69 161.3
R21797 minus.n72 minus.n57 161.3
R21798 minus.n74 minus.n73 161.3
R21799 minus.n76 minus.n75 161.3
R21800 minus.n77 minus.n55 161.3
R21801 minus.n79 minus.n78 161.3
R21802 minus.n81 minus.n80 161.3
R21803 minus.n82 minus.n53 161.3
R21804 minus.n85 minus.n84 161.3
R21805 minus.n86 minus.n52 161.3
R21806 minus.n88 minus.n87 161.3
R21807 minus.n90 minus.n51 161.3
R21808 minus.n92 minus.n91 161.3
R21809 minus.n94 minus.n93 161.3
R21810 minus.n95 minus.n49 161.3
R21811 minus.n97 minus.n96 161.3
R21812 minus.n48 minus.n47 161.3
R21813 minus.n46 minus.n0 161.3
R21814 minus.n45 minus.n44 161.3
R21815 minus.n43 minus.n42 161.3
R21816 minus.n41 minus.n2 161.3
R21817 minus.n39 minus.n38 161.3
R21818 minus.n37 minus.n3 161.3
R21819 minus.n36 minus.n35 161.3
R21820 minus.n33 minus.n4 161.3
R21821 minus.n32 minus.n31 161.3
R21822 minus.n30 minus.n29 161.3
R21823 minus.n28 minus.n6 161.3
R21824 minus.n27 minus.n26 161.3
R21825 minus.n25 minus.n24 161.3
R21826 minus.n23 minus.n8 161.3
R21827 minus.n21 minus.n20 161.3
R21828 minus.n19 minus.n9 161.3
R21829 minus.n18 minus.n17 161.3
R21830 minus.n15 minus.n10 161.3
R21831 minus.n14 minus.n13 161.3
R21832 minus.n91 minus.n90 56.5617
R21833 minus.n64 minus.n63 56.5617
R21834 minus.n15 minus.n14 56.5617
R21835 minus.n42 minus.n41 56.5617
R21836 minus.n82 minus.n81 56.5617
R21837 minus.n73 minus.n72 56.5617
R21838 minus.n24 minus.n23 56.5617
R21839 minus.n33 minus.n32 56.5617
R21840 minus.n95 minus.n94 48.3272
R21841 minus.n46 minus.n45 48.3272
R21842 minus.n84 minus.n52 44.4521
R21843 minus.n70 minus.n58 44.4521
R21844 minus.n21 minus.n9 44.4521
R21845 minus.n35 minus.n3 44.4521
R21846 minus.n13 minus.n12 43.0014
R21847 minus.n62 minus.n61 43.0014
R21848 minus.n78 minus.n77 40.577
R21849 minus.n77 minus.n76 40.577
R21850 minus.n28 minus.n27 40.577
R21851 minus.n29 minus.n28 40.577
R21852 minus.n61 minus.n60 39.4345
R21853 minus.n12 minus.n11 39.4345
R21854 minus.n88 minus.n52 36.702
R21855 minus.n66 minus.n58 36.702
R21856 minus.n17 minus.n9 36.702
R21857 minus.n39 minus.n3 36.702
R21858 minus.n98 minus.n97 33.563
R21859 minus.n90 minus.n89 20.9036
R21860 minus.n65 minus.n64 20.9036
R21861 minus.n16 minus.n15 20.9036
R21862 minus.n41 minus.n40 20.9036
R21863 minus.n100 minus.t3 19.8005
R21864 minus.n100 minus.t0 19.8005
R21865 minus.n99 minus.t2 19.8005
R21866 minus.n99 minus.t1 19.8005
R21867 minus.n81 minus.n54 18.9362
R21868 minus.n73 minus.n56 18.9362
R21869 minus.n24 minus.n7 18.9362
R21870 minus.n32 minus.n5 18.9362
R21871 minus.n83 minus.n82 16.9689
R21872 minus.n72 minus.n71 16.9689
R21873 minus.n23 minus.n22 16.9689
R21874 minus.n34 minus.n33 16.9689
R21875 minus.n91 minus.n50 15.0015
R21876 minus.n63 minus.n60 15.0015
R21877 minus.n14 minus.n11 15.0015
R21878 minus.n42 minus.n1 15.0015
R21879 minus.n96 minus.n95 12.4157
R21880 minus.n47 minus.n46 12.4157
R21881 minus.n98 minus.n48 12.1577
R21882 minus minus.n103 11.4024
R21883 minus.n94 minus.n50 9.59132
R21884 minus.n45 minus.n1 9.59132
R21885 minus.n84 minus.n83 7.62397
R21886 minus.n71 minus.n70 7.62397
R21887 minus.n22 minus.n21 7.62397
R21888 minus.n35 minus.n34 7.62397
R21889 minus.n78 minus.n54 5.65662
R21890 minus.n76 minus.n56 5.65662
R21891 minus.n27 minus.n7 5.65662
R21892 minus.n29 minus.n5 5.65662
R21893 minus.n103 minus.n102 4.80222
R21894 minus.n89 minus.n88 3.68928
R21895 minus.n66 minus.n65 3.68928
R21896 minus.n17 minus.n16 3.68928
R21897 minus.n40 minus.n39 3.68928
R21898 minus.n103 minus.n98 0.972091
R21899 minus.n102 minus.n101 0.716017
R21900 minus.n97 minus.n49 0.189894
R21901 minus.n93 minus.n49 0.189894
R21902 minus.n93 minus.n92 0.189894
R21903 minus.n92 minus.n51 0.189894
R21904 minus.n87 minus.n51 0.189894
R21905 minus.n87 minus.n86 0.189894
R21906 minus.n86 minus.n85 0.189894
R21907 minus.n85 minus.n53 0.189894
R21908 minus.n80 minus.n53 0.189894
R21909 minus.n80 minus.n79 0.189894
R21910 minus.n79 minus.n55 0.189894
R21911 minus.n75 minus.n55 0.189894
R21912 minus.n75 minus.n74 0.189894
R21913 minus.n74 minus.n57 0.189894
R21914 minus.n69 minus.n57 0.189894
R21915 minus.n69 minus.n68 0.189894
R21916 minus.n68 minus.n67 0.189894
R21917 minus.n67 minus.n59 0.189894
R21918 minus.n62 minus.n59 0.189894
R21919 minus.n13 minus.n10 0.189894
R21920 minus.n18 minus.n10 0.189894
R21921 minus.n19 minus.n18 0.189894
R21922 minus.n20 minus.n19 0.189894
R21923 minus.n20 minus.n8 0.189894
R21924 minus.n25 minus.n8 0.189894
R21925 minus.n26 minus.n25 0.189894
R21926 minus.n26 minus.n6 0.189894
R21927 minus.n30 minus.n6 0.189894
R21928 minus.n31 minus.n30 0.189894
R21929 minus.n31 minus.n4 0.189894
R21930 minus.n36 minus.n4 0.189894
R21931 minus.n37 minus.n36 0.189894
R21932 minus.n38 minus.n37 0.189894
R21933 minus.n38 minus.n2 0.189894
R21934 minus.n43 minus.n2 0.189894
R21935 minus.n44 minus.n43 0.189894
R21936 minus.n44 minus.n0 0.189894
R21937 minus.n48 minus.n0 0.189894
R21938 diffpairibias.n0 diffpairibias.t18 436.822
R21939 diffpairibias.n21 diffpairibias.t19 435.479
R21940 diffpairibias.n20 diffpairibias.t16 435.479
R21941 diffpairibias.n19 diffpairibias.t17 435.479
R21942 diffpairibias.n18 diffpairibias.t21 435.479
R21943 diffpairibias.n0 diffpairibias.t22 435.479
R21944 diffpairibias.n1 diffpairibias.t20 435.479
R21945 diffpairibias.n2 diffpairibias.t23 435.479
R21946 diffpairibias.n10 diffpairibias.t0 377.536
R21947 diffpairibias.n10 diffpairibias.t8 376.193
R21948 diffpairibias.n11 diffpairibias.t10 376.193
R21949 diffpairibias.n12 diffpairibias.t6 376.193
R21950 diffpairibias.n13 diffpairibias.t2 376.193
R21951 diffpairibias.n14 diffpairibias.t12 376.193
R21952 diffpairibias.n15 diffpairibias.t4 376.193
R21953 diffpairibias.n16 diffpairibias.t14 376.193
R21954 diffpairibias.n3 diffpairibias.t1 113.368
R21955 diffpairibias.n3 diffpairibias.t9 112.698
R21956 diffpairibias.n4 diffpairibias.t11 112.698
R21957 diffpairibias.n5 diffpairibias.t7 112.698
R21958 diffpairibias.n6 diffpairibias.t3 112.698
R21959 diffpairibias.n7 diffpairibias.t13 112.698
R21960 diffpairibias.n8 diffpairibias.t5 112.698
R21961 diffpairibias.n9 diffpairibias.t15 112.698
R21962 diffpairibias.n17 diffpairibias.n16 4.77242
R21963 diffpairibias.n17 diffpairibias.n9 4.30807
R21964 diffpairibias.n18 diffpairibias.n17 4.13945
R21965 diffpairibias.n16 diffpairibias.n15 1.34352
R21966 diffpairibias.n15 diffpairibias.n14 1.34352
R21967 diffpairibias.n14 diffpairibias.n13 1.34352
R21968 diffpairibias.n13 diffpairibias.n12 1.34352
R21969 diffpairibias.n12 diffpairibias.n11 1.34352
R21970 diffpairibias.n11 diffpairibias.n10 1.34352
R21971 diffpairibias.n2 diffpairibias.n1 1.34352
R21972 diffpairibias.n1 diffpairibias.n0 1.34352
R21973 diffpairibias.n19 diffpairibias.n18 1.34352
R21974 diffpairibias.n20 diffpairibias.n19 1.34352
R21975 diffpairibias.n21 diffpairibias.n20 1.34352
R21976 diffpairibias.n22 diffpairibias.n21 0.862419
R21977 diffpairibias diffpairibias.n22 0.684875
R21978 diffpairibias.n9 diffpairibias.n8 0.672012
R21979 diffpairibias.n8 diffpairibias.n7 0.672012
R21980 diffpairibias.n7 diffpairibias.n6 0.672012
R21981 diffpairibias.n6 diffpairibias.n5 0.672012
R21982 diffpairibias.n5 diffpairibias.n4 0.672012
R21983 diffpairibias.n4 diffpairibias.n3 0.672012
R21984 diffpairibias.n22 diffpairibias.n2 0.190907
R21985 outputibias.n27 outputibias.n1 289.615
R21986 outputibias.n58 outputibias.n32 289.615
R21987 outputibias.n90 outputibias.n64 289.615
R21988 outputibias.n122 outputibias.n96 289.615
R21989 outputibias.n28 outputibias.n27 185
R21990 outputibias.n26 outputibias.n25 185
R21991 outputibias.n5 outputibias.n4 185
R21992 outputibias.n20 outputibias.n19 185
R21993 outputibias.n18 outputibias.n17 185
R21994 outputibias.n9 outputibias.n8 185
R21995 outputibias.n12 outputibias.n11 185
R21996 outputibias.n59 outputibias.n58 185
R21997 outputibias.n57 outputibias.n56 185
R21998 outputibias.n36 outputibias.n35 185
R21999 outputibias.n51 outputibias.n50 185
R22000 outputibias.n49 outputibias.n48 185
R22001 outputibias.n40 outputibias.n39 185
R22002 outputibias.n43 outputibias.n42 185
R22003 outputibias.n91 outputibias.n90 185
R22004 outputibias.n89 outputibias.n88 185
R22005 outputibias.n68 outputibias.n67 185
R22006 outputibias.n83 outputibias.n82 185
R22007 outputibias.n81 outputibias.n80 185
R22008 outputibias.n72 outputibias.n71 185
R22009 outputibias.n75 outputibias.n74 185
R22010 outputibias.n123 outputibias.n122 185
R22011 outputibias.n121 outputibias.n120 185
R22012 outputibias.n100 outputibias.n99 185
R22013 outputibias.n115 outputibias.n114 185
R22014 outputibias.n113 outputibias.n112 185
R22015 outputibias.n104 outputibias.n103 185
R22016 outputibias.n107 outputibias.n106 185
R22017 outputibias.n0 outputibias.t10 178.945
R22018 outputibias.n133 outputibias.t8 177.018
R22019 outputibias.n132 outputibias.t11 177.018
R22020 outputibias.n0 outputibias.t9 177.018
R22021 outputibias.t7 outputibias.n10 147.661
R22022 outputibias.t1 outputibias.n41 147.661
R22023 outputibias.t3 outputibias.n73 147.661
R22024 outputibias.t5 outputibias.n105 147.661
R22025 outputibias.n128 outputibias.t6 132.363
R22026 outputibias.n128 outputibias.t0 130.436
R22027 outputibias.n129 outputibias.t2 130.436
R22028 outputibias.n130 outputibias.t4 130.436
R22029 outputibias.n27 outputibias.n26 104.615
R22030 outputibias.n26 outputibias.n4 104.615
R22031 outputibias.n19 outputibias.n4 104.615
R22032 outputibias.n19 outputibias.n18 104.615
R22033 outputibias.n18 outputibias.n8 104.615
R22034 outputibias.n11 outputibias.n8 104.615
R22035 outputibias.n58 outputibias.n57 104.615
R22036 outputibias.n57 outputibias.n35 104.615
R22037 outputibias.n50 outputibias.n35 104.615
R22038 outputibias.n50 outputibias.n49 104.615
R22039 outputibias.n49 outputibias.n39 104.615
R22040 outputibias.n42 outputibias.n39 104.615
R22041 outputibias.n90 outputibias.n89 104.615
R22042 outputibias.n89 outputibias.n67 104.615
R22043 outputibias.n82 outputibias.n67 104.615
R22044 outputibias.n82 outputibias.n81 104.615
R22045 outputibias.n81 outputibias.n71 104.615
R22046 outputibias.n74 outputibias.n71 104.615
R22047 outputibias.n122 outputibias.n121 104.615
R22048 outputibias.n121 outputibias.n99 104.615
R22049 outputibias.n114 outputibias.n99 104.615
R22050 outputibias.n114 outputibias.n113 104.615
R22051 outputibias.n113 outputibias.n103 104.615
R22052 outputibias.n106 outputibias.n103 104.615
R22053 outputibias.n63 outputibias.n31 95.6354
R22054 outputibias.n63 outputibias.n62 94.6732
R22055 outputibias.n95 outputibias.n94 94.6732
R22056 outputibias.n127 outputibias.n126 94.6732
R22057 outputibias.n11 outputibias.t7 52.3082
R22058 outputibias.n42 outputibias.t1 52.3082
R22059 outputibias.n74 outputibias.t3 52.3082
R22060 outputibias.n106 outputibias.t5 52.3082
R22061 outputibias.n12 outputibias.n10 15.6674
R22062 outputibias.n43 outputibias.n41 15.6674
R22063 outputibias.n75 outputibias.n73 15.6674
R22064 outputibias.n107 outputibias.n105 15.6674
R22065 outputibias.n13 outputibias.n9 12.8005
R22066 outputibias.n44 outputibias.n40 12.8005
R22067 outputibias.n76 outputibias.n72 12.8005
R22068 outputibias.n108 outputibias.n104 12.8005
R22069 outputibias.n17 outputibias.n16 12.0247
R22070 outputibias.n48 outputibias.n47 12.0247
R22071 outputibias.n80 outputibias.n79 12.0247
R22072 outputibias.n112 outputibias.n111 12.0247
R22073 outputibias.n20 outputibias.n7 11.249
R22074 outputibias.n51 outputibias.n38 11.249
R22075 outputibias.n83 outputibias.n70 11.249
R22076 outputibias.n115 outputibias.n102 11.249
R22077 outputibias.n21 outputibias.n5 10.4732
R22078 outputibias.n52 outputibias.n36 10.4732
R22079 outputibias.n84 outputibias.n68 10.4732
R22080 outputibias.n116 outputibias.n100 10.4732
R22081 outputibias.n25 outputibias.n24 9.69747
R22082 outputibias.n56 outputibias.n55 9.69747
R22083 outputibias.n88 outputibias.n87 9.69747
R22084 outputibias.n120 outputibias.n119 9.69747
R22085 outputibias.n31 outputibias.n30 9.45567
R22086 outputibias.n62 outputibias.n61 9.45567
R22087 outputibias.n94 outputibias.n93 9.45567
R22088 outputibias.n126 outputibias.n125 9.45567
R22089 outputibias.n30 outputibias.n29 9.3005
R22090 outputibias.n3 outputibias.n2 9.3005
R22091 outputibias.n24 outputibias.n23 9.3005
R22092 outputibias.n22 outputibias.n21 9.3005
R22093 outputibias.n7 outputibias.n6 9.3005
R22094 outputibias.n16 outputibias.n15 9.3005
R22095 outputibias.n14 outputibias.n13 9.3005
R22096 outputibias.n61 outputibias.n60 9.3005
R22097 outputibias.n34 outputibias.n33 9.3005
R22098 outputibias.n55 outputibias.n54 9.3005
R22099 outputibias.n53 outputibias.n52 9.3005
R22100 outputibias.n38 outputibias.n37 9.3005
R22101 outputibias.n47 outputibias.n46 9.3005
R22102 outputibias.n45 outputibias.n44 9.3005
R22103 outputibias.n93 outputibias.n92 9.3005
R22104 outputibias.n66 outputibias.n65 9.3005
R22105 outputibias.n87 outputibias.n86 9.3005
R22106 outputibias.n85 outputibias.n84 9.3005
R22107 outputibias.n70 outputibias.n69 9.3005
R22108 outputibias.n79 outputibias.n78 9.3005
R22109 outputibias.n77 outputibias.n76 9.3005
R22110 outputibias.n125 outputibias.n124 9.3005
R22111 outputibias.n98 outputibias.n97 9.3005
R22112 outputibias.n119 outputibias.n118 9.3005
R22113 outputibias.n117 outputibias.n116 9.3005
R22114 outputibias.n102 outputibias.n101 9.3005
R22115 outputibias.n111 outputibias.n110 9.3005
R22116 outputibias.n109 outputibias.n108 9.3005
R22117 outputibias.n28 outputibias.n3 8.92171
R22118 outputibias.n59 outputibias.n34 8.92171
R22119 outputibias.n91 outputibias.n66 8.92171
R22120 outputibias.n123 outputibias.n98 8.92171
R22121 outputibias.n29 outputibias.n1 8.14595
R22122 outputibias.n60 outputibias.n32 8.14595
R22123 outputibias.n92 outputibias.n64 8.14595
R22124 outputibias.n124 outputibias.n96 8.14595
R22125 outputibias.n31 outputibias.n1 5.81868
R22126 outputibias.n62 outputibias.n32 5.81868
R22127 outputibias.n94 outputibias.n64 5.81868
R22128 outputibias.n126 outputibias.n96 5.81868
R22129 outputibias.n131 outputibias.n130 5.20947
R22130 outputibias.n29 outputibias.n28 5.04292
R22131 outputibias.n60 outputibias.n59 5.04292
R22132 outputibias.n92 outputibias.n91 5.04292
R22133 outputibias.n124 outputibias.n123 5.04292
R22134 outputibias.n131 outputibias.n127 4.42209
R22135 outputibias.n14 outputibias.n10 4.38594
R22136 outputibias.n45 outputibias.n41 4.38594
R22137 outputibias.n77 outputibias.n73 4.38594
R22138 outputibias.n109 outputibias.n105 4.38594
R22139 outputibias.n132 outputibias.n131 4.28454
R22140 outputibias.n25 outputibias.n3 4.26717
R22141 outputibias.n56 outputibias.n34 4.26717
R22142 outputibias.n88 outputibias.n66 4.26717
R22143 outputibias.n120 outputibias.n98 4.26717
R22144 outputibias.n24 outputibias.n5 3.49141
R22145 outputibias.n55 outputibias.n36 3.49141
R22146 outputibias.n87 outputibias.n68 3.49141
R22147 outputibias.n119 outputibias.n100 3.49141
R22148 outputibias.n21 outputibias.n20 2.71565
R22149 outputibias.n52 outputibias.n51 2.71565
R22150 outputibias.n84 outputibias.n83 2.71565
R22151 outputibias.n116 outputibias.n115 2.71565
R22152 outputibias.n17 outputibias.n7 1.93989
R22153 outputibias.n48 outputibias.n38 1.93989
R22154 outputibias.n80 outputibias.n70 1.93989
R22155 outputibias.n112 outputibias.n102 1.93989
R22156 outputibias.n130 outputibias.n129 1.9266
R22157 outputibias.n129 outputibias.n128 1.9266
R22158 outputibias.n133 outputibias.n132 1.92658
R22159 outputibias.n134 outputibias.n133 1.29913
R22160 outputibias.n16 outputibias.n9 1.16414
R22161 outputibias.n47 outputibias.n40 1.16414
R22162 outputibias.n79 outputibias.n72 1.16414
R22163 outputibias.n111 outputibias.n104 1.16414
R22164 outputibias.n127 outputibias.n95 0.962709
R22165 outputibias.n95 outputibias.n63 0.962709
R22166 outputibias.n13 outputibias.n12 0.388379
R22167 outputibias.n44 outputibias.n43 0.388379
R22168 outputibias.n76 outputibias.n75 0.388379
R22169 outputibias.n108 outputibias.n107 0.388379
R22170 outputibias.n134 outputibias.n0 0.337251
R22171 outputibias outputibias.n134 0.302375
R22172 outputibias.n30 outputibias.n2 0.155672
R22173 outputibias.n23 outputibias.n2 0.155672
R22174 outputibias.n23 outputibias.n22 0.155672
R22175 outputibias.n22 outputibias.n6 0.155672
R22176 outputibias.n15 outputibias.n6 0.155672
R22177 outputibias.n15 outputibias.n14 0.155672
R22178 outputibias.n61 outputibias.n33 0.155672
R22179 outputibias.n54 outputibias.n33 0.155672
R22180 outputibias.n54 outputibias.n53 0.155672
R22181 outputibias.n53 outputibias.n37 0.155672
R22182 outputibias.n46 outputibias.n37 0.155672
R22183 outputibias.n46 outputibias.n45 0.155672
R22184 outputibias.n93 outputibias.n65 0.155672
R22185 outputibias.n86 outputibias.n65 0.155672
R22186 outputibias.n86 outputibias.n85 0.155672
R22187 outputibias.n85 outputibias.n69 0.155672
R22188 outputibias.n78 outputibias.n69 0.155672
R22189 outputibias.n78 outputibias.n77 0.155672
R22190 outputibias.n125 outputibias.n97 0.155672
R22191 outputibias.n118 outputibias.n97 0.155672
R22192 outputibias.n118 outputibias.n117 0.155672
R22193 outputibias.n117 outputibias.n101 0.155672
R22194 outputibias.n110 outputibias.n101 0.155672
R22195 outputibias.n110 outputibias.n109 0.155672
C0 CSoutput output 6.13881f
C1 CSoutput outputibias 0.032386f
C2 vdd CSoutput 67.6707f
C3 minus diffpairibias 5.12e-19
C4 commonsourceibias output 0.006808f
C5 CSoutput minus 2.65135f
C6 vdd plus 0.070154f
C7 plus diffpairibias 4.13e-19
C8 commonsourceibias outputibias 0.003832f
C9 vdd commonsourceibias 0.004218f
C10 CSoutput plus 0.875866f
C11 commonsourceibias diffpairibias 0.06482f
C12 CSoutput commonsourceibias 54.0646f
C13 minus plus 9.61291f
C14 minus commonsourceibias 0.462932f
C15 plus commonsourceibias 0.417773f
C16 output outputibias 2.34152f
C17 vdd output 7.23429f
C18 diffpairibias gnd 48.98024f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.183165p
C22 plus gnd 35.556202f
C23 minus gnd 28.47191f
C24 CSoutput gnd 0.125529p
C25 vdd gnd 0.345104p
C26 outputibias.t9 gnd 0.11477f
C27 outputibias.t10 gnd 0.115567f
C28 outputibias.n0 gnd 0.130108f
C29 outputibias.n1 gnd 0.001372f
C30 outputibias.n2 gnd 9.76e-19
C31 outputibias.n3 gnd 5.24e-19
C32 outputibias.n4 gnd 0.001239f
C33 outputibias.n5 gnd 5.55e-19
C34 outputibias.n6 gnd 9.76e-19
C35 outputibias.n7 gnd 5.24e-19
C36 outputibias.n8 gnd 0.001239f
C37 outputibias.n9 gnd 5.55e-19
C38 outputibias.n10 gnd 0.004176f
C39 outputibias.t7 gnd 0.00202f
C40 outputibias.n11 gnd 9.3e-19
C41 outputibias.n12 gnd 7.32e-19
C42 outputibias.n13 gnd 5.24e-19
C43 outputibias.n14 gnd 0.02322f
C44 outputibias.n15 gnd 9.76e-19
C45 outputibias.n16 gnd 5.24e-19
C46 outputibias.n17 gnd 5.55e-19
C47 outputibias.n18 gnd 0.001239f
C48 outputibias.n19 gnd 0.001239f
C49 outputibias.n20 gnd 5.55e-19
C50 outputibias.n21 gnd 5.24e-19
C51 outputibias.n22 gnd 9.76e-19
C52 outputibias.n23 gnd 9.76e-19
C53 outputibias.n24 gnd 5.24e-19
C54 outputibias.n25 gnd 5.55e-19
C55 outputibias.n26 gnd 0.001239f
C56 outputibias.n27 gnd 0.002683f
C57 outputibias.n28 gnd 5.55e-19
C58 outputibias.n29 gnd 5.24e-19
C59 outputibias.n30 gnd 0.002256f
C60 outputibias.n31 gnd 0.005781f
C61 outputibias.n32 gnd 0.001372f
C62 outputibias.n33 gnd 9.76e-19
C63 outputibias.n34 gnd 5.24e-19
C64 outputibias.n35 gnd 0.001239f
C65 outputibias.n36 gnd 5.55e-19
C66 outputibias.n37 gnd 9.76e-19
C67 outputibias.n38 gnd 5.24e-19
C68 outputibias.n39 gnd 0.001239f
C69 outputibias.n40 gnd 5.55e-19
C70 outputibias.n41 gnd 0.004176f
C71 outputibias.t1 gnd 0.00202f
C72 outputibias.n42 gnd 9.3e-19
C73 outputibias.n43 gnd 7.32e-19
C74 outputibias.n44 gnd 5.24e-19
C75 outputibias.n45 gnd 0.02322f
C76 outputibias.n46 gnd 9.76e-19
C77 outputibias.n47 gnd 5.24e-19
C78 outputibias.n48 gnd 5.55e-19
C79 outputibias.n49 gnd 0.001239f
C80 outputibias.n50 gnd 0.001239f
C81 outputibias.n51 gnd 5.55e-19
C82 outputibias.n52 gnd 5.24e-19
C83 outputibias.n53 gnd 9.76e-19
C84 outputibias.n54 gnd 9.76e-19
C85 outputibias.n55 gnd 5.24e-19
C86 outputibias.n56 gnd 5.55e-19
C87 outputibias.n57 gnd 0.001239f
C88 outputibias.n58 gnd 0.002683f
C89 outputibias.n59 gnd 5.55e-19
C90 outputibias.n60 gnd 5.24e-19
C91 outputibias.n61 gnd 0.002256f
C92 outputibias.n62 gnd 0.005197f
C93 outputibias.n63 gnd 0.121892f
C94 outputibias.n64 gnd 0.001372f
C95 outputibias.n65 gnd 9.76e-19
C96 outputibias.n66 gnd 5.24e-19
C97 outputibias.n67 gnd 0.001239f
C98 outputibias.n68 gnd 5.55e-19
C99 outputibias.n69 gnd 9.76e-19
C100 outputibias.n70 gnd 5.24e-19
C101 outputibias.n71 gnd 0.001239f
C102 outputibias.n72 gnd 5.55e-19
C103 outputibias.n73 gnd 0.004176f
C104 outputibias.t3 gnd 0.00202f
C105 outputibias.n74 gnd 9.3e-19
C106 outputibias.n75 gnd 7.32e-19
C107 outputibias.n76 gnd 5.24e-19
C108 outputibias.n77 gnd 0.02322f
C109 outputibias.n78 gnd 9.76e-19
C110 outputibias.n79 gnd 5.24e-19
C111 outputibias.n80 gnd 5.55e-19
C112 outputibias.n81 gnd 0.001239f
C113 outputibias.n82 gnd 0.001239f
C114 outputibias.n83 gnd 5.55e-19
C115 outputibias.n84 gnd 5.24e-19
C116 outputibias.n85 gnd 9.76e-19
C117 outputibias.n86 gnd 9.76e-19
C118 outputibias.n87 gnd 5.24e-19
C119 outputibias.n88 gnd 5.55e-19
C120 outputibias.n89 gnd 0.001239f
C121 outputibias.n90 gnd 0.002683f
C122 outputibias.n91 gnd 5.55e-19
C123 outputibias.n92 gnd 5.24e-19
C124 outputibias.n93 gnd 0.002256f
C125 outputibias.n94 gnd 0.005197f
C126 outputibias.n95 gnd 0.064513f
C127 outputibias.n96 gnd 0.001372f
C128 outputibias.n97 gnd 9.76e-19
C129 outputibias.n98 gnd 5.24e-19
C130 outputibias.n99 gnd 0.001239f
C131 outputibias.n100 gnd 5.55e-19
C132 outputibias.n101 gnd 9.76e-19
C133 outputibias.n102 gnd 5.24e-19
C134 outputibias.n103 gnd 0.001239f
C135 outputibias.n104 gnd 5.55e-19
C136 outputibias.n105 gnd 0.004176f
C137 outputibias.t5 gnd 0.00202f
C138 outputibias.n106 gnd 9.3e-19
C139 outputibias.n107 gnd 7.32e-19
C140 outputibias.n108 gnd 5.24e-19
C141 outputibias.n109 gnd 0.02322f
C142 outputibias.n110 gnd 9.76e-19
C143 outputibias.n111 gnd 5.24e-19
C144 outputibias.n112 gnd 5.55e-19
C145 outputibias.n113 gnd 0.001239f
C146 outputibias.n114 gnd 0.001239f
C147 outputibias.n115 gnd 5.55e-19
C148 outputibias.n116 gnd 5.24e-19
C149 outputibias.n117 gnd 9.76e-19
C150 outputibias.n118 gnd 9.76e-19
C151 outputibias.n119 gnd 5.24e-19
C152 outputibias.n120 gnd 5.55e-19
C153 outputibias.n121 gnd 0.001239f
C154 outputibias.n122 gnd 0.002683f
C155 outputibias.n123 gnd 5.55e-19
C156 outputibias.n124 gnd 5.24e-19
C157 outputibias.n125 gnd 0.002256f
C158 outputibias.n126 gnd 0.005197f
C159 outputibias.n127 gnd 0.084814f
C160 outputibias.t4 gnd 0.108319f
C161 outputibias.t2 gnd 0.108319f
C162 outputibias.t0 gnd 0.108319f
C163 outputibias.t6 gnd 0.109238f
C164 outputibias.n128 gnd 0.134674f
C165 outputibias.n129 gnd 0.07244f
C166 outputibias.n130 gnd 0.079818f
C167 outputibias.n131 gnd 0.164901f
C168 outputibias.t11 gnd 0.11477f
C169 outputibias.n132 gnd 0.067481f
C170 outputibias.t8 gnd 0.11477f
C171 outputibias.n133 gnd 0.065115f
C172 outputibias.n134 gnd 0.029159f
C173 diffpairibias.t18 gnd 0.087401f
C174 diffpairibias.t22 gnd 0.087239f
C175 diffpairibias.n0 gnd 0.102784f
C176 diffpairibias.t20 gnd 0.087239f
C177 diffpairibias.n1 gnd 0.050171f
C178 diffpairibias.t23 gnd 0.087239f
C179 diffpairibias.n2 gnd 0.039841f
C180 diffpairibias.t1 gnd 0.083757f
C181 diffpairibias.t9 gnd 0.083392f
C182 diffpairibias.n3 gnd 0.131682f
C183 diffpairibias.t11 gnd 0.083392f
C184 diffpairibias.n4 gnd 0.07027f
C185 diffpairibias.t7 gnd 0.083392f
C186 diffpairibias.n5 gnd 0.07027f
C187 diffpairibias.t3 gnd 0.083392f
C188 diffpairibias.n6 gnd 0.07027f
C189 diffpairibias.t13 gnd 0.083392f
C190 diffpairibias.n7 gnd 0.07027f
C191 diffpairibias.t5 gnd 0.083392f
C192 diffpairibias.n8 gnd 0.07027f
C193 diffpairibias.t15 gnd 0.083392f
C194 diffpairibias.n9 gnd 0.099771f
C195 diffpairibias.t0 gnd 0.08427f
C196 diffpairibias.t8 gnd 0.084123f
C197 diffpairibias.n10 gnd 0.091784f
C198 diffpairibias.t10 gnd 0.084123f
C199 diffpairibias.n11 gnd 0.050681f
C200 diffpairibias.t6 gnd 0.084123f
C201 diffpairibias.n12 gnd 0.050681f
C202 diffpairibias.t2 gnd 0.084123f
C203 diffpairibias.n13 gnd 0.050681f
C204 diffpairibias.t12 gnd 0.084123f
C205 diffpairibias.n14 gnd 0.050681f
C206 diffpairibias.t4 gnd 0.084123f
C207 diffpairibias.n15 gnd 0.050681f
C208 diffpairibias.t14 gnd 0.084123f
C209 diffpairibias.n16 gnd 0.059977f
C210 diffpairibias.n17 gnd 0.226448f
C211 diffpairibias.t21 gnd 0.087239f
C212 diffpairibias.n18 gnd 0.050181f
C213 diffpairibias.t17 gnd 0.087239f
C214 diffpairibias.n19 gnd 0.050171f
C215 diffpairibias.t16 gnd 0.087239f
C216 diffpairibias.n20 gnd 0.050171f
C217 diffpairibias.t19 gnd 0.087239f
C218 diffpairibias.n21 gnd 0.045859f
C219 diffpairibias.n22 gnd 0.046268f
C220 minus.n0 gnd 0.030653f
C221 minus.t13 gnd 0.51542f
C222 minus.n1 gnd 0.208459f
C223 minus.n2 gnd 0.030653f
C224 minus.t20 gnd 0.51542f
C225 minus.n3 gnd 0.025388f
C226 minus.n4 gnd 0.030653f
C227 minus.t17 gnd 0.51542f
C228 minus.t23 gnd 0.51542f
C229 minus.n5 gnd 0.208459f
C230 minus.n6 gnd 0.030653f
C231 minus.t22 gnd 0.51542f
C232 minus.n7 gnd 0.208459f
C233 minus.n8 gnd 0.030653f
C234 minus.t5 gnd 0.51542f
C235 minus.n9 gnd 0.025388f
C236 minus.n10 gnd 0.030653f
C237 minus.t8 gnd 0.51542f
C238 minus.t10 gnd 0.51542f
C239 minus.n11 gnd 0.239719f
C240 minus.t16 gnd 0.57765f
C241 minus.n12 gnd 0.242787f
C242 minus.n13 gnd 0.130833f
C243 minus.n14 gnd 0.038703f
C244 minus.n15 gnd 0.035261f
C245 minus.n16 gnd 0.208459f
C246 minus.n17 gnd 0.03762f
C247 minus.n18 gnd 0.030653f
C248 minus.n19 gnd 0.030653f
C249 minus.n20 gnd 0.030653f
C250 minus.n21 gnd 0.039737f
C251 minus.n22 gnd 0.208459f
C252 minus.n23 gnd 0.037555f
C253 minus.n24 gnd 0.036408f
C254 minus.n25 gnd 0.030653f
C255 minus.n26 gnd 0.030653f
C256 minus.n27 gnd 0.038994f
C257 minus.n28 gnd 0.024757f
C258 minus.n29 gnd 0.038994f
C259 minus.n30 gnd 0.030653f
C260 minus.n31 gnd 0.030653f
C261 minus.n32 gnd 0.036408f
C262 minus.n33 gnd 0.037555f
C263 minus.n34 gnd 0.208459f
C264 minus.n35 gnd 0.039737f
C265 minus.n36 gnd 0.030653f
C266 minus.n37 gnd 0.030653f
C267 minus.n38 gnd 0.030653f
C268 minus.n39 gnd 0.03762f
C269 minus.n40 gnd 0.208459f
C270 minus.n41 gnd 0.035261f
C271 minus.n42 gnd 0.038703f
C272 minus.n43 gnd 0.030653f
C273 minus.n44 gnd 0.030653f
C274 minus.n45 gnd 0.040001f
C275 minus.n46 gnd 0.011871f
C276 minus.t9 gnd 0.557427f
C277 minus.n47 gnd 0.241738f
C278 minus.n48 gnd 0.359629f
C279 minus.n49 gnd 0.030653f
C280 minus.t14 gnd 0.557427f
C281 minus.t21 gnd 0.51542f
C282 minus.n50 gnd 0.208459f
C283 minus.n51 gnd 0.030653f
C284 minus.t18 gnd 0.51542f
C285 minus.n52 gnd 0.025388f
C286 minus.n53 gnd 0.030653f
C287 minus.t15 gnd 0.51542f
C288 minus.t7 gnd 0.51542f
C289 minus.n54 gnd 0.208459f
C290 minus.n55 gnd 0.030653f
C291 minus.t6 gnd 0.51542f
C292 minus.n56 gnd 0.208459f
C293 minus.n57 gnd 0.030653f
C294 minus.t12 gnd 0.51542f
C295 minus.n58 gnd 0.025388f
C296 minus.n59 gnd 0.030653f
C297 minus.t11 gnd 0.51542f
C298 minus.t19 gnd 0.51542f
C299 minus.n60 gnd 0.239719f
C300 minus.t24 gnd 0.57765f
C301 minus.n61 gnd 0.242787f
C302 minus.n62 gnd 0.130833f
C303 minus.n63 gnd 0.038703f
C304 minus.n64 gnd 0.035261f
C305 minus.n65 gnd 0.208459f
C306 minus.n66 gnd 0.03762f
C307 minus.n67 gnd 0.030653f
C308 minus.n68 gnd 0.030653f
C309 minus.n69 gnd 0.030653f
C310 minus.n70 gnd 0.039737f
C311 minus.n71 gnd 0.208459f
C312 minus.n72 gnd 0.037555f
C313 minus.n73 gnd 0.036408f
C314 minus.n74 gnd 0.030653f
C315 minus.n75 gnd 0.030653f
C316 minus.n76 gnd 0.038994f
C317 minus.n77 gnd 0.024757f
C318 minus.n78 gnd 0.038994f
C319 minus.n79 gnd 0.030653f
C320 minus.n80 gnd 0.030653f
C321 minus.n81 gnd 0.036408f
C322 minus.n82 gnd 0.037555f
C323 minus.n83 gnd 0.208459f
C324 minus.n84 gnd 0.039737f
C325 minus.n85 gnd 0.030653f
C326 minus.n86 gnd 0.030653f
C327 minus.n87 gnd 0.030653f
C328 minus.n88 gnd 0.03762f
C329 minus.n89 gnd 0.208459f
C330 minus.n90 gnd 0.035261f
C331 minus.n91 gnd 0.038703f
C332 minus.n92 gnd 0.030653f
C333 minus.n93 gnd 0.030653f
C334 minus.n94 gnd 0.040001f
C335 minus.n95 gnd 0.011871f
C336 minus.n96 gnd 0.241738f
C337 minus.n97 gnd 1.03605f
C338 minus.n98 gnd 1.5397f
C339 minus.t2 gnd 0.009449f
C340 minus.t1 gnd 0.009449f
C341 minus.n99 gnd 0.031072f
C342 minus.t3 gnd 0.009449f
C343 minus.t0 gnd 0.009449f
C344 minus.n100 gnd 0.030646f
C345 minus.n101 gnd 0.261548f
C346 minus.t4 gnd 0.052594f
C347 minus.n102 gnd 0.142724f
C348 minus.n103 gnd 1.83725f
C349 output.t6 gnd 0.464308f
C350 output.t11 gnd 0.044422f
C351 output.t16 gnd 0.044422f
C352 output.n0 gnd 0.364624f
C353 output.n1 gnd 0.614102f
C354 output.t4 gnd 0.044422f
C355 output.t12 gnd 0.044422f
C356 output.n2 gnd 0.364624f
C357 output.n3 gnd 0.350265f
C358 output.t15 gnd 0.044422f
C359 output.t13 gnd 0.044422f
C360 output.n4 gnd 0.364624f
C361 output.n5 gnd 0.350265f
C362 output.t3 gnd 0.044422f
C363 output.t5 gnd 0.044422f
C364 output.n6 gnd 0.364624f
C365 output.n7 gnd 0.350265f
C366 output.t8 gnd 0.044422f
C367 output.t17 gnd 0.044422f
C368 output.n8 gnd 0.364624f
C369 output.n9 gnd 0.350265f
C370 output.t18 gnd 0.044422f
C371 output.t9 gnd 0.044422f
C372 output.n10 gnd 0.364624f
C373 output.n11 gnd 0.350265f
C374 output.t10 gnd 0.044422f
C375 output.t14 gnd 0.044422f
C376 output.n12 gnd 0.364624f
C377 output.n13 gnd 0.350265f
C378 output.t7 gnd 0.462979f
C379 output.n14 gnd 0.28994f
C380 output.n15 gnd 0.015803f
C381 output.n16 gnd 0.011243f
C382 output.n17 gnd 0.006041f
C383 output.n18 gnd 0.01428f
C384 output.n19 gnd 0.006397f
C385 output.n20 gnd 0.011243f
C386 output.n21 gnd 0.006041f
C387 output.n22 gnd 0.01428f
C388 output.n23 gnd 0.006397f
C389 output.n24 gnd 0.048111f
C390 output.t1 gnd 0.023274f
C391 output.n25 gnd 0.01071f
C392 output.n26 gnd 0.008435f
C393 output.n27 gnd 0.006041f
C394 output.n28 gnd 0.267512f
C395 output.n29 gnd 0.011243f
C396 output.n30 gnd 0.006041f
C397 output.n31 gnd 0.006397f
C398 output.n32 gnd 0.01428f
C399 output.n33 gnd 0.01428f
C400 output.n34 gnd 0.006397f
C401 output.n35 gnd 0.006041f
C402 output.n36 gnd 0.011243f
C403 output.n37 gnd 0.011243f
C404 output.n38 gnd 0.006041f
C405 output.n39 gnd 0.006397f
C406 output.n40 gnd 0.01428f
C407 output.n41 gnd 0.030913f
C408 output.n42 gnd 0.006397f
C409 output.n43 gnd 0.006041f
C410 output.n44 gnd 0.025987f
C411 output.n45 gnd 0.097665f
C412 output.n46 gnd 0.015803f
C413 output.n47 gnd 0.011243f
C414 output.n48 gnd 0.006041f
C415 output.n49 gnd 0.01428f
C416 output.n50 gnd 0.006397f
C417 output.n51 gnd 0.011243f
C418 output.n52 gnd 0.006041f
C419 output.n53 gnd 0.01428f
C420 output.n54 gnd 0.006397f
C421 output.n55 gnd 0.048111f
C422 output.t2 gnd 0.023274f
C423 output.n56 gnd 0.01071f
C424 output.n57 gnd 0.008435f
C425 output.n58 gnd 0.006041f
C426 output.n59 gnd 0.267512f
C427 output.n60 gnd 0.011243f
C428 output.n61 gnd 0.006041f
C429 output.n62 gnd 0.006397f
C430 output.n63 gnd 0.01428f
C431 output.n64 gnd 0.01428f
C432 output.n65 gnd 0.006397f
C433 output.n66 gnd 0.006041f
C434 output.n67 gnd 0.011243f
C435 output.n68 gnd 0.011243f
C436 output.n69 gnd 0.006041f
C437 output.n70 gnd 0.006397f
C438 output.n71 gnd 0.01428f
C439 output.n72 gnd 0.030913f
C440 output.n73 gnd 0.006397f
C441 output.n74 gnd 0.006041f
C442 output.n75 gnd 0.025987f
C443 output.n76 gnd 0.09306f
C444 output.n77 gnd 1.65264f
C445 output.n78 gnd 0.015803f
C446 output.n79 gnd 0.011243f
C447 output.n80 gnd 0.006041f
C448 output.n81 gnd 0.01428f
C449 output.n82 gnd 0.006397f
C450 output.n83 gnd 0.011243f
C451 output.n84 gnd 0.006041f
C452 output.n85 gnd 0.01428f
C453 output.n86 gnd 0.006397f
C454 output.n87 gnd 0.048111f
C455 output.t19 gnd 0.023274f
C456 output.n88 gnd 0.01071f
C457 output.n89 gnd 0.008435f
C458 output.n90 gnd 0.006041f
C459 output.n91 gnd 0.267512f
C460 output.n92 gnd 0.011243f
C461 output.n93 gnd 0.006041f
C462 output.n94 gnd 0.006397f
C463 output.n95 gnd 0.01428f
C464 output.n96 gnd 0.01428f
C465 output.n97 gnd 0.006397f
C466 output.n98 gnd 0.006041f
C467 output.n99 gnd 0.011243f
C468 output.n100 gnd 0.011243f
C469 output.n101 gnd 0.006041f
C470 output.n102 gnd 0.006397f
C471 output.n103 gnd 0.01428f
C472 output.n104 gnd 0.030913f
C473 output.n105 gnd 0.006397f
C474 output.n106 gnd 0.006041f
C475 output.n107 gnd 0.025987f
C476 output.n108 gnd 0.09306f
C477 output.n109 gnd 0.713089f
C478 output.n110 gnd 0.015803f
C479 output.n111 gnd 0.011243f
C480 output.n112 gnd 0.006041f
C481 output.n113 gnd 0.01428f
C482 output.n114 gnd 0.006397f
C483 output.n115 gnd 0.011243f
C484 output.n116 gnd 0.006041f
C485 output.n117 gnd 0.01428f
C486 output.n118 gnd 0.006397f
C487 output.n119 gnd 0.048111f
C488 output.t0 gnd 0.023274f
C489 output.n120 gnd 0.01071f
C490 output.n121 gnd 0.008435f
C491 output.n122 gnd 0.006041f
C492 output.n123 gnd 0.267512f
C493 output.n124 gnd 0.011243f
C494 output.n125 gnd 0.006041f
C495 output.n126 gnd 0.006397f
C496 output.n127 gnd 0.01428f
C497 output.n128 gnd 0.01428f
C498 output.n129 gnd 0.006397f
C499 output.n130 gnd 0.006041f
C500 output.n131 gnd 0.011243f
C501 output.n132 gnd 0.011243f
C502 output.n133 gnd 0.006041f
C503 output.n134 gnd 0.006397f
C504 output.n135 gnd 0.01428f
C505 output.n136 gnd 0.030913f
C506 output.n137 gnd 0.006397f
C507 output.n138 gnd 0.006041f
C508 output.n139 gnd 0.025987f
C509 output.n140 gnd 0.09306f
C510 output.n141 gnd 1.67353f
C511 a_n2903_n3924.t10 gnd 0.094851f
C512 a_n2903_n3924.t20 gnd 0.985803f
C513 a_n2903_n3924.n0 gnd 0.372677f
C514 a_n2903_n3924.t4 gnd 1.22484f
C515 a_n2903_n3924.n1 gnd 1.15477f
C516 a_n2903_n3924.t40 gnd 0.985803f
C517 a_n2903_n3924.n2 gnd 0.372677f
C518 a_n2903_n3924.t27 gnd 0.094851f
C519 a_n2903_n3924.t41 gnd 0.094851f
C520 a_n2903_n3924.n3 gnd 0.774663f
C521 a_n2903_n3924.n4 gnd 0.390386f
C522 a_n2903_n3924.t37 gnd 0.094851f
C523 a_n2903_n3924.t45 gnd 0.094851f
C524 a_n2903_n3924.n5 gnd 0.774663f
C525 a_n2903_n3924.n6 gnd 0.390386f
C526 a_n2903_n3924.t2 gnd 0.094851f
C527 a_n2903_n3924.t28 gnd 0.094851f
C528 a_n2903_n3924.n7 gnd 0.774663f
C529 a_n2903_n3924.n8 gnd 0.390386f
C530 a_n2903_n3924.t3 gnd 0.094851f
C531 a_n2903_n3924.t44 gnd 0.094851f
C532 a_n2903_n3924.n9 gnd 0.774663f
C533 a_n2903_n3924.n10 gnd 0.390386f
C534 a_n2903_n3924.t42 gnd 0.985803f
C535 a_n2903_n3924.n11 gnd 0.922787f
C536 a_n2903_n3924.t47 gnd 1.22537f
C537 a_n2903_n3924.t0 gnd 1.22484f
C538 a_n2903_n3924.n12 gnd 0.862674f
C539 a_n2903_n3924.t33 gnd 1.22484f
C540 a_n2903_n3924.n13 gnd 0.862674f
C541 a_n2903_n3924.t29 gnd 1.22484f
C542 a_n2903_n3924.n14 gnd 0.862674f
C543 a_n2903_n3924.t1 gnd 1.22484f
C544 a_n2903_n3924.n15 gnd 0.862674f
C545 a_n2903_n3924.t30 gnd 1.22484f
C546 a_n2903_n3924.n16 gnd 0.862674f
C547 a_n2903_n3924.t46 gnd 1.22484f
C548 a_n2903_n3924.n17 gnd 0.716127f
C549 a_n2903_n3924.n18 gnd 0.845678f
C550 a_n2903_n3924.n19 gnd 0.894202f
C551 a_n2903_n3924.t25 gnd 0.985799f
C552 a_n2903_n3924.n20 gnd 0.612329f
C553 a_n2903_n3924.t19 gnd 0.094851f
C554 a_n2903_n3924.t23 gnd 0.094851f
C555 a_n2903_n3924.n21 gnd 0.774662f
C556 a_n2903_n3924.n22 gnd 0.390388f
C557 a_n2903_n3924.t24 gnd 0.094851f
C558 a_n2903_n3924.t12 gnd 0.094851f
C559 a_n2903_n3924.n23 gnd 0.774662f
C560 a_n2903_n3924.n24 gnd 0.390388f
C561 a_n2903_n3924.t13 gnd 0.094851f
C562 a_n2903_n3924.t7 gnd 0.094851f
C563 a_n2903_n3924.n25 gnd 0.774662f
C564 a_n2903_n3924.n26 gnd 0.390388f
C565 a_n2903_n3924.t9 gnd 0.094851f
C566 a_n2903_n3924.t22 gnd 0.094851f
C567 a_n2903_n3924.n27 gnd 0.774662f
C568 a_n2903_n3924.n28 gnd 0.390388f
C569 a_n2903_n3924.t17 gnd 0.985799f
C570 a_n2903_n3924.n29 gnd 0.372681f
C571 a_n2903_n3924.t5 gnd 0.985799f
C572 a_n2903_n3924.n30 gnd 0.372681f
C573 a_n2903_n3924.t35 gnd 0.094851f
C574 a_n2903_n3924.t32 gnd 0.094851f
C575 a_n2903_n3924.n31 gnd 0.774662f
C576 a_n2903_n3924.n32 gnd 0.390388f
C577 a_n2903_n3924.t34 gnd 0.094851f
C578 a_n2903_n3924.t39 gnd 0.094851f
C579 a_n2903_n3924.n33 gnd 0.774662f
C580 a_n2903_n3924.n34 gnd 0.390388f
C581 a_n2903_n3924.t6 gnd 0.094851f
C582 a_n2903_n3924.t43 gnd 0.094851f
C583 a_n2903_n3924.n35 gnd 0.774662f
C584 a_n2903_n3924.n36 gnd 0.390388f
C585 a_n2903_n3924.t31 gnd 0.094851f
C586 a_n2903_n3924.t38 gnd 0.094851f
C587 a_n2903_n3924.n37 gnd 0.774662f
C588 a_n2903_n3924.n38 gnd 0.390388f
C589 a_n2903_n3924.t36 gnd 0.985799f
C590 a_n2903_n3924.n39 gnd 0.612329f
C591 a_n2903_n3924.n40 gnd 0.953249f
C592 a_n2903_n3924.t8 gnd 0.985799f
C593 a_n2903_n3924.n41 gnd 0.922791f
C594 a_n2903_n3924.t16 gnd 0.094851f
C595 a_n2903_n3924.t21 gnd 0.094851f
C596 a_n2903_n3924.n42 gnd 0.774663f
C597 a_n2903_n3924.n43 gnd 0.390386f
C598 a_n2903_n3924.t14 gnd 0.094851f
C599 a_n2903_n3924.t18 gnd 0.094851f
C600 a_n2903_n3924.n44 gnd 0.774663f
C601 a_n2903_n3924.n45 gnd 0.390386f
C602 a_n2903_n3924.t11 gnd 0.094851f
C603 a_n2903_n3924.t15 gnd 0.094851f
C604 a_n2903_n3924.n46 gnd 0.774663f
C605 a_n2903_n3924.n47 gnd 0.390386f
C606 a_n2903_n3924.n48 gnd 0.390385f
C607 a_n2903_n3924.n49 gnd 0.774664f
C608 a_n2903_n3924.t26 gnd 0.094851f
C609 plus.n0 gnd 0.022688f
C610 plus.t6 gnd 0.412586f
C611 plus.t12 gnd 0.381494f
C612 plus.n1 gnd 0.154293f
C613 plus.n2 gnd 0.022688f
C614 plus.t8 gnd 0.381494f
C615 plus.n3 gnd 0.018791f
C616 plus.n4 gnd 0.022688f
C617 plus.t7 gnd 0.381494f
C618 plus.t19 gnd 0.381494f
C619 plus.n5 gnd 0.154293f
C620 plus.n6 gnd 0.022688f
C621 plus.t18 gnd 0.381494f
C622 plus.n7 gnd 0.154293f
C623 plus.n8 gnd 0.022688f
C624 plus.t24 gnd 0.381494f
C625 plus.n9 gnd 0.018791f
C626 plus.n10 gnd 0.022688f
C627 plus.t22 gnd 0.381494f
C628 plus.t9 gnd 0.381494f
C629 plus.n11 gnd 0.177431f
C630 plus.t14 gnd 0.427554f
C631 plus.n12 gnd 0.179702f
C632 plus.n13 gnd 0.096838f
C633 plus.n14 gnd 0.028646f
C634 plus.n15 gnd 0.026099f
C635 plus.n16 gnd 0.154293f
C636 plus.n17 gnd 0.027845f
C637 plus.n18 gnd 0.022688f
C638 plus.n19 gnd 0.022688f
C639 plus.n20 gnd 0.022688f
C640 plus.n21 gnd 0.029412f
C641 plus.n22 gnd 0.154293f
C642 plus.n23 gnd 0.027797f
C643 plus.n24 gnd 0.026948f
C644 plus.n25 gnd 0.022688f
C645 plus.n26 gnd 0.022688f
C646 plus.n27 gnd 0.028862f
C647 plus.n28 gnd 0.018324f
C648 plus.n29 gnd 0.028862f
C649 plus.n30 gnd 0.022688f
C650 plus.n31 gnd 0.022688f
C651 plus.n32 gnd 0.026948f
C652 plus.n33 gnd 0.027797f
C653 plus.n34 gnd 0.154293f
C654 plus.n35 gnd 0.029412f
C655 plus.n36 gnd 0.022688f
C656 plus.n37 gnd 0.022688f
C657 plus.n38 gnd 0.022688f
C658 plus.n39 gnd 0.027845f
C659 plus.n40 gnd 0.154293f
C660 plus.n41 gnd 0.026099f
C661 plus.n42 gnd 0.028646f
C662 plus.n43 gnd 0.022688f
C663 plus.n44 gnd 0.022688f
C664 plus.n45 gnd 0.029607f
C665 plus.n46 gnd 0.008787f
C666 plus.n47 gnd 0.178925f
C667 plus.n48 gnd 0.260348f
C668 plus.n49 gnd 0.022688f
C669 plus.t10 gnd 0.381494f
C670 plus.n50 gnd 0.154293f
C671 plus.n51 gnd 0.022688f
C672 plus.t15 gnd 0.381494f
C673 plus.n52 gnd 0.018791f
C674 plus.n53 gnd 0.022688f
C675 plus.t13 gnd 0.381494f
C676 plus.t17 gnd 0.381494f
C677 plus.n54 gnd 0.154293f
C678 plus.n55 gnd 0.022688f
C679 plus.t16 gnd 0.381494f
C680 plus.n56 gnd 0.154293f
C681 plus.n57 gnd 0.022688f
C682 plus.t20 gnd 0.381494f
C683 plus.n58 gnd 0.018791f
C684 plus.n59 gnd 0.022688f
C685 plus.t21 gnd 0.381494f
C686 plus.t5 gnd 0.381494f
C687 plus.n60 gnd 0.177431f
C688 plus.t11 gnd 0.427554f
C689 plus.n61 gnd 0.179702f
C690 plus.n62 gnd 0.096838f
C691 plus.n63 gnd 0.028646f
C692 plus.n64 gnd 0.026099f
C693 plus.n65 gnd 0.154293f
C694 plus.n66 gnd 0.027845f
C695 plus.n67 gnd 0.022688f
C696 plus.n68 gnd 0.022688f
C697 plus.n69 gnd 0.022688f
C698 plus.n70 gnd 0.029412f
C699 plus.n71 gnd 0.154293f
C700 plus.n72 gnd 0.027797f
C701 plus.n73 gnd 0.026948f
C702 plus.n74 gnd 0.022688f
C703 plus.n75 gnd 0.022688f
C704 plus.n76 gnd 0.028862f
C705 plus.n77 gnd 0.018324f
C706 plus.n78 gnd 0.028862f
C707 plus.n79 gnd 0.022688f
C708 plus.n80 gnd 0.022688f
C709 plus.n81 gnd 0.026948f
C710 plus.n82 gnd 0.027797f
C711 plus.n83 gnd 0.154293f
C712 plus.n84 gnd 0.029412f
C713 plus.n85 gnd 0.022688f
C714 plus.n86 gnd 0.022688f
C715 plus.n87 gnd 0.022688f
C716 plus.n88 gnd 0.027845f
C717 plus.n89 gnd 0.154293f
C718 plus.n90 gnd 0.026099f
C719 plus.n91 gnd 0.028646f
C720 plus.n92 gnd 0.022688f
C721 plus.n93 gnd 0.022688f
C722 plus.n94 gnd 0.029607f
C723 plus.n95 gnd 0.008787f
C724 plus.t23 gnd 0.412586f
C725 plus.n96 gnd 0.178925f
C726 plus.n97 gnd 0.757758f
C727 plus.n98 gnd 1.13063f
C728 plus.t1 gnd 0.039166f
C729 plus.t2 gnd 0.006994f
C730 plus.t4 gnd 0.006994f
C731 plus.n99 gnd 0.022683f
C732 plus.n100 gnd 0.176089f
C733 plus.t0 gnd 0.006994f
C734 plus.t3 gnd 0.006994f
C735 plus.n101 gnd 0.022683f
C736 plus.n102 gnd 0.132176f
C737 plus.n103 gnd 2.65938f
C738 a_n1808_13878.t4 gnd 0.185683f
C739 a_n1808_13878.t0 gnd 0.185683f
C740 a_n1808_13878.t2 gnd 0.185683f
C741 a_n1808_13878.n0 gnd 1.46364f
C742 a_n1808_13878.t6 gnd 0.185683f
C743 a_n1808_13878.t1 gnd 0.185683f
C744 a_n1808_13878.n1 gnd 1.46209f
C745 a_n1808_13878.n2 gnd 2.04299f
C746 a_n1808_13878.t5 gnd 0.185683f
C747 a_n1808_13878.t9 gnd 0.185683f
C748 a_n1808_13878.n3 gnd 1.46451f
C749 a_n1808_13878.t10 gnd 0.185683f
C750 a_n1808_13878.t3 gnd 0.185683f
C751 a_n1808_13878.n4 gnd 1.46209f
C752 a_n1808_13878.n5 gnd 1.31424f
C753 a_n1808_13878.t7 gnd 0.185683f
C754 a_n1808_13878.t8 gnd 0.185683f
C755 a_n1808_13878.n6 gnd 1.46209f
C756 a_n1808_13878.n7 gnd 1.80499f
C757 a_n1808_13878.t13 gnd 1.73864f
C758 a_n1808_13878.t16 gnd 0.185683f
C759 a_n1808_13878.t17 gnd 0.185683f
C760 a_n1808_13878.n8 gnd 1.30795f
C761 a_n1808_13878.n9 gnd 1.46144f
C762 a_n1808_13878.t12 gnd 1.73518f
C763 a_n1808_13878.n10 gnd 0.735417f
C764 a_n1808_13878.t15 gnd 1.73518f
C765 a_n1808_13878.n11 gnd 0.735417f
C766 a_n1808_13878.t18 gnd 0.185683f
C767 a_n1808_13878.t19 gnd 0.185683f
C768 a_n1808_13878.n12 gnd 1.30795f
C769 a_n1808_13878.n13 gnd 0.742539f
C770 a_n1808_13878.t14 gnd 1.73518f
C771 a_n1808_13878.n14 gnd 1.73174f
C772 a_n1808_13878.n15 gnd 2.52099f
C773 a_n1808_13878.n16 gnd 3.70273f
C774 a_n1808_13878.n17 gnd 1.46209f
C775 a_n1808_13878.t11 gnd 0.185683f
C776 a_n2356_n452.n0 gnd 0.521964f
C777 a_n2356_n452.n1 gnd 0.203307f
C778 a_n2356_n452.n2 gnd 0.149739f
C779 a_n2356_n452.n3 gnd 0.235343f
C780 a_n2356_n452.n4 gnd 0.181775f
C781 a_n2356_n452.n5 gnd 0.203307f
C782 a_n2356_n452.n6 gnd 0.149739f
C783 a_n2356_n452.n7 gnd 0.575531f
C784 a_n2356_n452.n8 gnd 0.428941f
C785 a_n2356_n452.n9 gnd 0.21427f
C786 a_n2356_n452.n10 gnd 0.488658f
C787 a_n2356_n452.n11 gnd 0.280324f
C788 a_n2356_n452.n12 gnd 0.43509f
C789 a_n2356_n452.n13 gnd 0.21427f
C790 a_n2356_n452.n14 gnd 0.725869f
C791 a_n2356_n452.n15 gnd 0.280324f
C792 a_n2356_n452.n16 gnd 0.634249f
C793 a_n2356_n452.n17 gnd 0.280324f
C794 a_n2356_n452.n18 gnd 0.488658f
C795 a_n2356_n452.n19 gnd 0.659289f
C796 a_n2356_n452.n20 gnd 0.21427f
C797 a_n2356_n452.n21 gnd 0.280324f
C798 a_n2356_n452.n22 gnd 3.29653f
C799 a_n2356_n452.n23 gnd 1.76406f
C800 a_n2356_n452.n24 gnd 1.16973f
C801 a_n2356_n452.n25 gnd 1.90084f
C802 a_n2356_n452.n26 gnd 0.283453f
C803 a_n2356_n452.n27 gnd 0.008296f
C804 a_n2356_n452.n29 gnd 1.32808f
C805 a_n2356_n452.n30 gnd 0.283453f
C806 a_n2356_n452.n31 gnd 0.008296f
C807 a_n2356_n452.n32 gnd 0.008296f
C808 a_n2356_n452.n34 gnd 0.283453f
C809 a_n2356_n452.n35 gnd 0.008296f
C810 a_n2356_n452.n37 gnd 0.283453f
C811 a_n2356_n452.n38 gnd 0.008296f
C812 a_n2356_n452.n39 gnd 0.28305f
C813 a_n2356_n452.n40 gnd 0.008296f
C814 a_n2356_n452.n41 gnd 0.28305f
C815 a_n2356_n452.n42 gnd 0.008296f
C816 a_n2356_n452.n43 gnd 0.28305f
C817 a_n2356_n452.n44 gnd 0.008296f
C818 a_n2356_n452.n45 gnd 0.28305f
C819 a_n2356_n452.n47 gnd 0.303943f
C820 a_n2356_n452.t11 gnd 0.14862f
C821 a_n2356_n452.t23 gnd 1.3916f
C822 a_n2356_n452.t15 gnd 0.14862f
C823 a_n2356_n452.t21 gnd 0.14862f
C824 a_n2356_n452.n48 gnd 1.04688f
C825 a_n2356_n452.t2 gnd 0.691309f
C826 a_n2356_n452.n49 gnd 0.303943f
C827 a_n2356_n452.t10 gnd 0.691309f
C828 a_n2356_n452.t14 gnd 0.691309f
C829 a_n2356_n452.t52 gnd 0.691309f
C830 a_n2356_n452.n50 gnd 0.303943f
C831 a_n2356_n452.t61 gnd 0.691309f
C832 a_n2356_n452.t67 gnd 0.691309f
C833 a_n2356_n452.t8 gnd 0.705869f
C834 a_n2356_n452.t12 gnd 0.691309f
C835 a_n2356_n452.t6 gnd 0.691309f
C836 a_n2356_n452.t4 gnd 0.691309f
C837 a_n2356_n452.t16 gnd 0.691309f
C838 a_n2356_n452.t18 gnd 0.702738f
C839 a_n2356_n452.t71 gnd 0.705869f
C840 a_n2356_n452.t54 gnd 0.691309f
C841 a_n2356_n452.t58 gnd 0.691309f
C842 a_n2356_n452.t48 gnd 0.691309f
C843 a_n2356_n452.n51 gnd 0.303943f
C844 a_n2356_n452.t63 gnd 0.691309f
C845 a_n2356_n452.t69 gnd 0.702738f
C846 a_n2356_n452.n52 gnd 0.30654f
C847 a_n2356_n452.n53 gnd 0.300083f
C848 a_n2356_n452.n54 gnd 0.30654f
C849 a_n2356_n452.n55 gnd 0.30654f
C850 a_n2356_n452.t26 gnd 0.115593f
C851 a_n2356_n452.t33 gnd 0.115593f
C852 a_n2356_n452.n56 gnd 1.02443f
C853 a_n2356_n452.t31 gnd 0.115593f
C854 a_n2356_n452.t32 gnd 0.115593f
C855 a_n2356_n452.n57 gnd 1.02142f
C856 a_n2356_n452.n58 gnd 0.905747f
C857 a_n2356_n452.t37 gnd 0.115593f
C858 a_n2356_n452.t27 gnd 0.115593f
C859 a_n2356_n452.n59 gnd 1.02142f
C860 a_n2356_n452.t36 gnd 0.115593f
C861 a_n2356_n452.t34 gnd 0.115593f
C862 a_n2356_n452.n60 gnd 1.02443f
C863 a_n2356_n452.t41 gnd 0.115593f
C864 a_n2356_n452.t30 gnd 0.115593f
C865 a_n2356_n452.n61 gnd 1.02142f
C866 a_n2356_n452.n62 gnd 0.905747f
C867 a_n2356_n452.n63 gnd 2.76749f
C868 a_n2356_n452.t40 gnd 0.115593f
C869 a_n2356_n452.t1 gnd 0.115593f
C870 a_n2356_n452.n64 gnd 1.02142f
C871 a_n2356_n452.n65 gnd 2.95023f
C872 a_n2356_n452.t42 gnd 0.115593f
C873 a_n2356_n452.t0 gnd 0.115593f
C874 a_n2356_n452.n66 gnd 1.02142f
C875 a_n2356_n452.n67 gnd 0.445962f
C876 a_n2356_n452.t29 gnd 0.115593f
C877 a_n2356_n452.t35 gnd 0.115593f
C878 a_n2356_n452.n68 gnd 1.02142f
C879 a_n2356_n452.t39 gnd 0.115593f
C880 a_n2356_n452.t38 gnd 0.115593f
C881 a_n2356_n452.n69 gnd 1.02444f
C882 a_n2356_n452.t43 gnd 0.115593f
C883 a_n2356_n452.t28 gnd 0.115593f
C884 a_n2356_n452.n70 gnd 1.02142f
C885 a_n2356_n452.n71 gnd 0.905745f
C886 a_n2356_n452.n72 gnd 3.10539f
C887 a_n2356_n452.n73 gnd 0.300083f
C888 a_n2356_n452.n74 gnd 0.30654f
C889 a_n2356_n452.t19 gnd 1.3916f
C890 a_n2356_n452.t5 gnd 0.14862f
C891 a_n2356_n452.t17 gnd 0.14862f
C892 a_n2356_n452.n75 gnd 1.04688f
C893 a_n2356_n452.t13 gnd 0.14862f
C894 a_n2356_n452.t7 gnd 0.14862f
C895 a_n2356_n452.n76 gnd 1.04688f
C896 a_n2356_n452.t9 gnd 1.38883f
C897 a_n2356_n452.n77 gnd 1.13572f
C898 a_n2356_n452.n78 gnd 0.78084f
C899 a_n2356_n452.t53 gnd 0.691309f
C900 a_n2356_n452.t62 gnd 0.691309f
C901 a_n2356_n452.t44 gnd 0.691309f
C902 a_n2356_n452.n79 gnd 0.303943f
C903 a_n2356_n452.t64 gnd 0.691309f
C904 a_n2356_n452.t49 gnd 0.691309f
C905 a_n2356_n452.t50 gnd 0.691309f
C906 a_n2356_n452.n80 gnd 0.303943f
C907 a_n2356_n452.t68 gnd 0.691309f
C908 a_n2356_n452.t57 gnd 0.691309f
C909 a_n2356_n452.t56 gnd 0.691309f
C910 a_n2356_n452.n81 gnd 0.303943f
C911 a_n2356_n452.t60 gnd 0.691309f
C912 a_n2356_n452.t51 gnd 0.691309f
C913 a_n2356_n452.t45 gnd 0.691309f
C914 a_n2356_n452.n82 gnd 0.303943f
C915 a_n2356_n452.t65 gnd 0.702892f
C916 a_n2356_n452.n83 gnd 0.300083f
C917 a_n2356_n452.n84 gnd 0.294634f
C918 a_n2356_n452.t70 gnd 0.702892f
C919 a_n2356_n452.n85 gnd 0.300083f
C920 a_n2356_n452.n86 gnd 0.294634f
C921 a_n2356_n452.t59 gnd 0.702892f
C922 a_n2356_n452.n87 gnd 0.300083f
C923 a_n2356_n452.n88 gnd 0.294634f
C924 a_n2356_n452.t55 gnd 0.702892f
C925 a_n2356_n452.n89 gnd 0.300083f
C926 a_n2356_n452.n90 gnd 0.294634f
C927 a_n2356_n452.n91 gnd 0.998508f
C928 a_n2356_n452.t66 gnd 0.705869f
C929 a_n2356_n452.n92 gnd 0.30654f
C930 a_n2356_n452.t46 gnd 0.691309f
C931 a_n2356_n452.n93 gnd 0.300083f
C932 a_n2356_n452.n94 gnd 0.30654f
C933 a_n2356_n452.t47 gnd 0.702738f
C934 a_n2356_n452.t22 gnd 0.705869f
C935 a_n2356_n452.n95 gnd 0.30654f
C936 a_n2356_n452.t20 gnd 0.691309f
C937 a_n2356_n452.n96 gnd 0.300083f
C938 a_n2356_n452.n97 gnd 0.30654f
C939 a_n2356_n452.t24 gnd 0.702738f
C940 a_n2356_n452.n98 gnd 1.12327f
C941 a_n2356_n452.t25 gnd 1.38883f
C942 a_n2356_n452.n99 gnd 1.04688f
C943 a_n2356_n452.t3 gnd 0.14862f
C944 vdd.t152 gnd 0.032956f
C945 vdd.t150 gnd 0.032956f
C946 vdd.n0 gnd 0.259932f
C947 vdd.t178 gnd 0.032956f
C948 vdd.t194 gnd 0.032956f
C949 vdd.n1 gnd 0.259503f
C950 vdd.n2 gnd 0.239312f
C951 vdd.t184 gnd 0.032956f
C952 vdd.t190 gnd 0.032956f
C953 vdd.n3 gnd 0.259503f
C954 vdd.n4 gnd 0.121029f
C955 vdd.t192 gnd 0.032956f
C956 vdd.t142 gnd 0.032956f
C957 vdd.n5 gnd 0.259503f
C958 vdd.n6 gnd 0.113563f
C959 vdd.t199 gnd 0.032956f
C960 vdd.t188 gnd 0.032956f
C961 vdd.n7 gnd 0.259932f
C962 vdd.t144 gnd 0.032956f
C963 vdd.t158 gnd 0.032956f
C964 vdd.n8 gnd 0.259503f
C965 vdd.n9 gnd 0.239312f
C966 vdd.t196 gnd 0.032956f
C967 vdd.t181 gnd 0.032956f
C968 vdd.n10 gnd 0.259503f
C969 vdd.n11 gnd 0.121029f
C970 vdd.t148 gnd 0.032956f
C971 vdd.t155 gnd 0.032956f
C972 vdd.n12 gnd 0.259503f
C973 vdd.n13 gnd 0.113563f
C974 vdd.n14 gnd 0.080287f
C975 vdd.t170 gnd 0.018309f
C976 vdd.t171 gnd 0.018309f
C977 vdd.n15 gnd 0.168528f
C978 vdd.t168 gnd 0.018309f
C979 vdd.t169 gnd 0.018309f
C980 vdd.n16 gnd 0.168034f
C981 vdd.n17 gnd 0.292432f
C982 vdd.t172 gnd 0.018309f
C983 vdd.t166 gnd 0.018309f
C984 vdd.n18 gnd 0.168034f
C985 vdd.n19 gnd 0.120983f
C986 vdd.t167 gnd 0.018309f
C987 vdd.t175 gnd 0.018309f
C988 vdd.n20 gnd 0.168528f
C989 vdd.t173 gnd 0.018309f
C990 vdd.t160 gnd 0.018309f
C991 vdd.n21 gnd 0.168034f
C992 vdd.n22 gnd 0.292432f
C993 vdd.t163 gnd 0.018309f
C994 vdd.t165 gnd 0.018309f
C995 vdd.n23 gnd 0.168034f
C996 vdd.n24 gnd 0.120983f
C997 vdd.t161 gnd 0.018309f
C998 vdd.t162 gnd 0.018309f
C999 vdd.n25 gnd 0.168034f
C1000 vdd.t164 gnd 0.018309f
C1001 vdd.t174 gnd 0.018309f
C1002 vdd.n26 gnd 0.168034f
C1003 vdd.n27 gnd 18.423f
C1004 vdd.n28 gnd 6.88036f
C1005 vdd.n29 gnd 0.004994f
C1006 vdd.n30 gnd 0.004634f
C1007 vdd.n31 gnd 0.002563f
C1008 vdd.n32 gnd 0.005886f
C1009 vdd.n33 gnd 0.00249f
C1010 vdd.n34 gnd 0.002637f
C1011 vdd.n35 gnd 0.004634f
C1012 vdd.n36 gnd 0.00249f
C1013 vdd.n37 gnd 0.005886f
C1014 vdd.n38 gnd 0.002637f
C1015 vdd.n39 gnd 0.004634f
C1016 vdd.n40 gnd 0.00249f
C1017 vdd.n41 gnd 0.004414f
C1018 vdd.n42 gnd 0.004427f
C1019 vdd.t4 gnd 0.012645f
C1020 vdd.n43 gnd 0.028134f
C1021 vdd.n44 gnd 0.146416f
C1022 vdd.n45 gnd 0.00249f
C1023 vdd.n46 gnd 0.002637f
C1024 vdd.n47 gnd 0.005886f
C1025 vdd.n48 gnd 0.005886f
C1026 vdd.n49 gnd 0.002637f
C1027 vdd.n50 gnd 0.00249f
C1028 vdd.n51 gnd 0.004634f
C1029 vdd.n52 gnd 0.004634f
C1030 vdd.n53 gnd 0.00249f
C1031 vdd.n54 gnd 0.002637f
C1032 vdd.n55 gnd 0.005886f
C1033 vdd.n56 gnd 0.005886f
C1034 vdd.n57 gnd 0.002637f
C1035 vdd.n58 gnd 0.00249f
C1036 vdd.n59 gnd 0.004634f
C1037 vdd.n60 gnd 0.004634f
C1038 vdd.n61 gnd 0.00249f
C1039 vdd.n62 gnd 0.002637f
C1040 vdd.n63 gnd 0.005886f
C1041 vdd.n64 gnd 0.005886f
C1042 vdd.n65 gnd 0.013915f
C1043 vdd.n66 gnd 0.002563f
C1044 vdd.n67 gnd 0.00249f
C1045 vdd.n68 gnd 0.011977f
C1046 vdd.n69 gnd 0.008362f
C1047 vdd.t56 gnd 0.029295f
C1048 vdd.t30 gnd 0.029295f
C1049 vdd.n70 gnd 0.201332f
C1050 vdd.n71 gnd 0.158317f
C1051 vdd.t63 gnd 0.029295f
C1052 vdd.t19 gnd 0.029295f
C1053 vdd.n72 gnd 0.201332f
C1054 vdd.n73 gnd 0.127761f
C1055 vdd.t49 gnd 0.029295f
C1056 vdd.t24 gnd 0.029295f
C1057 vdd.n74 gnd 0.201332f
C1058 vdd.n75 gnd 0.127761f
C1059 vdd.n76 gnd 0.004994f
C1060 vdd.n77 gnd 0.004634f
C1061 vdd.n78 gnd 0.002563f
C1062 vdd.n79 gnd 0.005886f
C1063 vdd.n80 gnd 0.00249f
C1064 vdd.n81 gnd 0.002637f
C1065 vdd.n82 gnd 0.004634f
C1066 vdd.n83 gnd 0.00249f
C1067 vdd.n84 gnd 0.005886f
C1068 vdd.n85 gnd 0.002637f
C1069 vdd.n86 gnd 0.004634f
C1070 vdd.n87 gnd 0.00249f
C1071 vdd.n88 gnd 0.004414f
C1072 vdd.n89 gnd 0.004427f
C1073 vdd.t62 gnd 0.012645f
C1074 vdd.n90 gnd 0.028134f
C1075 vdd.n91 gnd 0.146416f
C1076 vdd.n92 gnd 0.00249f
C1077 vdd.n93 gnd 0.002637f
C1078 vdd.n94 gnd 0.005886f
C1079 vdd.n95 gnd 0.005886f
C1080 vdd.n96 gnd 0.002637f
C1081 vdd.n97 gnd 0.00249f
C1082 vdd.n98 gnd 0.004634f
C1083 vdd.n99 gnd 0.004634f
C1084 vdd.n100 gnd 0.00249f
C1085 vdd.n101 gnd 0.002637f
C1086 vdd.n102 gnd 0.005886f
C1087 vdd.n103 gnd 0.005886f
C1088 vdd.n104 gnd 0.002637f
C1089 vdd.n105 gnd 0.00249f
C1090 vdd.n106 gnd 0.004634f
C1091 vdd.n107 gnd 0.004634f
C1092 vdd.n108 gnd 0.00249f
C1093 vdd.n109 gnd 0.002637f
C1094 vdd.n110 gnd 0.005886f
C1095 vdd.n111 gnd 0.005886f
C1096 vdd.n112 gnd 0.013915f
C1097 vdd.n113 gnd 0.002563f
C1098 vdd.n114 gnd 0.00249f
C1099 vdd.n115 gnd 0.011977f
C1100 vdd.n116 gnd 0.008099f
C1101 vdd.n117 gnd 0.095055f
C1102 vdd.n118 gnd 0.004994f
C1103 vdd.n119 gnd 0.004634f
C1104 vdd.n120 gnd 0.002563f
C1105 vdd.n121 gnd 0.005886f
C1106 vdd.n122 gnd 0.00249f
C1107 vdd.n123 gnd 0.002637f
C1108 vdd.n124 gnd 0.004634f
C1109 vdd.n125 gnd 0.00249f
C1110 vdd.n126 gnd 0.005886f
C1111 vdd.n127 gnd 0.002637f
C1112 vdd.n128 gnd 0.004634f
C1113 vdd.n129 gnd 0.00249f
C1114 vdd.n130 gnd 0.004414f
C1115 vdd.n131 gnd 0.004427f
C1116 vdd.t31 gnd 0.012645f
C1117 vdd.n132 gnd 0.028134f
C1118 vdd.n133 gnd 0.146416f
C1119 vdd.n134 gnd 0.00249f
C1120 vdd.n135 gnd 0.002637f
C1121 vdd.n136 gnd 0.005886f
C1122 vdd.n137 gnd 0.005886f
C1123 vdd.n138 gnd 0.002637f
C1124 vdd.n139 gnd 0.00249f
C1125 vdd.n140 gnd 0.004634f
C1126 vdd.n141 gnd 0.004634f
C1127 vdd.n142 gnd 0.00249f
C1128 vdd.n143 gnd 0.002637f
C1129 vdd.n144 gnd 0.005886f
C1130 vdd.n145 gnd 0.005886f
C1131 vdd.n146 gnd 0.002637f
C1132 vdd.n147 gnd 0.00249f
C1133 vdd.n148 gnd 0.004634f
C1134 vdd.n149 gnd 0.004634f
C1135 vdd.n150 gnd 0.00249f
C1136 vdd.n151 gnd 0.002637f
C1137 vdd.n152 gnd 0.005886f
C1138 vdd.n153 gnd 0.005886f
C1139 vdd.n154 gnd 0.013915f
C1140 vdd.n155 gnd 0.002563f
C1141 vdd.n156 gnd 0.00249f
C1142 vdd.n157 gnd 0.011977f
C1143 vdd.n158 gnd 0.008362f
C1144 vdd.t33 gnd 0.029295f
C1145 vdd.t44 gnd 0.029295f
C1146 vdd.n159 gnd 0.201332f
C1147 vdd.n160 gnd 0.158317f
C1148 vdd.t8 gnd 0.029295f
C1149 vdd.t27 gnd 0.029295f
C1150 vdd.n161 gnd 0.201332f
C1151 vdd.n162 gnd 0.127761f
C1152 vdd.t43 gnd 0.029295f
C1153 vdd.t64 gnd 0.029295f
C1154 vdd.n163 gnd 0.201332f
C1155 vdd.n164 gnd 0.127761f
C1156 vdd.n165 gnd 0.004994f
C1157 vdd.n166 gnd 0.004634f
C1158 vdd.n167 gnd 0.002563f
C1159 vdd.n168 gnd 0.005886f
C1160 vdd.n169 gnd 0.00249f
C1161 vdd.n170 gnd 0.002637f
C1162 vdd.n171 gnd 0.004634f
C1163 vdd.n172 gnd 0.00249f
C1164 vdd.n173 gnd 0.005886f
C1165 vdd.n174 gnd 0.002637f
C1166 vdd.n175 gnd 0.004634f
C1167 vdd.n176 gnd 0.00249f
C1168 vdd.n177 gnd 0.004414f
C1169 vdd.n178 gnd 0.004427f
C1170 vdd.t21 gnd 0.012645f
C1171 vdd.n179 gnd 0.028134f
C1172 vdd.n180 gnd 0.146416f
C1173 vdd.n181 gnd 0.00249f
C1174 vdd.n182 gnd 0.002637f
C1175 vdd.n183 gnd 0.005886f
C1176 vdd.n184 gnd 0.005886f
C1177 vdd.n185 gnd 0.002637f
C1178 vdd.n186 gnd 0.00249f
C1179 vdd.n187 gnd 0.004634f
C1180 vdd.n188 gnd 0.004634f
C1181 vdd.n189 gnd 0.00249f
C1182 vdd.n190 gnd 0.002637f
C1183 vdd.n191 gnd 0.005886f
C1184 vdd.n192 gnd 0.005886f
C1185 vdd.n193 gnd 0.002637f
C1186 vdd.n194 gnd 0.00249f
C1187 vdd.n195 gnd 0.004634f
C1188 vdd.n196 gnd 0.004634f
C1189 vdd.n197 gnd 0.00249f
C1190 vdd.n198 gnd 0.002637f
C1191 vdd.n199 gnd 0.005886f
C1192 vdd.n200 gnd 0.005886f
C1193 vdd.n201 gnd 0.013915f
C1194 vdd.n202 gnd 0.002563f
C1195 vdd.n203 gnd 0.00249f
C1196 vdd.n204 gnd 0.011977f
C1197 vdd.n205 gnd 0.008099f
C1198 vdd.n206 gnd 0.056548f
C1199 vdd.n207 gnd 0.203758f
C1200 vdd.n208 gnd 0.004994f
C1201 vdd.n209 gnd 0.004634f
C1202 vdd.n210 gnd 0.002563f
C1203 vdd.n211 gnd 0.005886f
C1204 vdd.n212 gnd 0.00249f
C1205 vdd.n213 gnd 0.002637f
C1206 vdd.n214 gnd 0.004634f
C1207 vdd.n215 gnd 0.00249f
C1208 vdd.n216 gnd 0.005886f
C1209 vdd.n217 gnd 0.002637f
C1210 vdd.n218 gnd 0.004634f
C1211 vdd.n219 gnd 0.00249f
C1212 vdd.n220 gnd 0.004414f
C1213 vdd.n221 gnd 0.004427f
C1214 vdd.t36 gnd 0.012645f
C1215 vdd.n222 gnd 0.028134f
C1216 vdd.n223 gnd 0.146416f
C1217 vdd.n224 gnd 0.00249f
C1218 vdd.n225 gnd 0.002637f
C1219 vdd.n226 gnd 0.005886f
C1220 vdd.n227 gnd 0.005886f
C1221 vdd.n228 gnd 0.002637f
C1222 vdd.n229 gnd 0.00249f
C1223 vdd.n230 gnd 0.004634f
C1224 vdd.n231 gnd 0.004634f
C1225 vdd.n232 gnd 0.00249f
C1226 vdd.n233 gnd 0.002637f
C1227 vdd.n234 gnd 0.005886f
C1228 vdd.n235 gnd 0.005886f
C1229 vdd.n236 gnd 0.002637f
C1230 vdd.n237 gnd 0.00249f
C1231 vdd.n238 gnd 0.004634f
C1232 vdd.n239 gnd 0.004634f
C1233 vdd.n240 gnd 0.00249f
C1234 vdd.n241 gnd 0.002637f
C1235 vdd.n242 gnd 0.005886f
C1236 vdd.n243 gnd 0.005886f
C1237 vdd.n244 gnd 0.013915f
C1238 vdd.n245 gnd 0.002563f
C1239 vdd.n246 gnd 0.00249f
C1240 vdd.n247 gnd 0.011977f
C1241 vdd.n248 gnd 0.008362f
C1242 vdd.t37 gnd 0.029295f
C1243 vdd.t53 gnd 0.029295f
C1244 vdd.n249 gnd 0.201332f
C1245 vdd.n250 gnd 0.158317f
C1246 vdd.t14 gnd 0.029295f
C1247 vdd.t35 gnd 0.029295f
C1248 vdd.n251 gnd 0.201332f
C1249 vdd.n252 gnd 0.127761f
C1250 vdd.t48 gnd 0.029295f
C1251 vdd.t12 gnd 0.029295f
C1252 vdd.n253 gnd 0.201332f
C1253 vdd.n254 gnd 0.127761f
C1254 vdd.n255 gnd 0.004994f
C1255 vdd.n256 gnd 0.004634f
C1256 vdd.n257 gnd 0.002563f
C1257 vdd.n258 gnd 0.005886f
C1258 vdd.n259 gnd 0.00249f
C1259 vdd.n260 gnd 0.002637f
C1260 vdd.n261 gnd 0.004634f
C1261 vdd.n262 gnd 0.00249f
C1262 vdd.n263 gnd 0.005886f
C1263 vdd.n264 gnd 0.002637f
C1264 vdd.n265 gnd 0.004634f
C1265 vdd.n266 gnd 0.00249f
C1266 vdd.n267 gnd 0.004414f
C1267 vdd.n268 gnd 0.004427f
C1268 vdd.t25 gnd 0.012645f
C1269 vdd.n269 gnd 0.028134f
C1270 vdd.n270 gnd 0.146416f
C1271 vdd.n271 gnd 0.00249f
C1272 vdd.n272 gnd 0.002637f
C1273 vdd.n273 gnd 0.005886f
C1274 vdd.n274 gnd 0.005886f
C1275 vdd.n275 gnd 0.002637f
C1276 vdd.n276 gnd 0.00249f
C1277 vdd.n277 gnd 0.004634f
C1278 vdd.n278 gnd 0.004634f
C1279 vdd.n279 gnd 0.00249f
C1280 vdd.n280 gnd 0.002637f
C1281 vdd.n281 gnd 0.005886f
C1282 vdd.n282 gnd 0.005886f
C1283 vdd.n283 gnd 0.002637f
C1284 vdd.n284 gnd 0.00249f
C1285 vdd.n285 gnd 0.004634f
C1286 vdd.n286 gnd 0.004634f
C1287 vdd.n287 gnd 0.00249f
C1288 vdd.n288 gnd 0.002637f
C1289 vdd.n289 gnd 0.005886f
C1290 vdd.n290 gnd 0.005886f
C1291 vdd.n291 gnd 0.013915f
C1292 vdd.n292 gnd 0.002563f
C1293 vdd.n293 gnd 0.00249f
C1294 vdd.n294 gnd 0.011977f
C1295 vdd.n295 gnd 0.008099f
C1296 vdd.n296 gnd 0.056548f
C1297 vdd.n297 gnd 0.220543f
C1298 vdd.n298 gnd 0.006993f
C1299 vdd.n299 gnd 0.009099f
C1300 vdd.n300 gnd 0.007324f
C1301 vdd.n301 gnd 0.007324f
C1302 vdd.n302 gnd 0.009099f
C1303 vdd.n303 gnd 0.009099f
C1304 vdd.n304 gnd 0.664865f
C1305 vdd.n305 gnd 0.009099f
C1306 vdd.n306 gnd 0.009099f
C1307 vdd.n307 gnd 0.009099f
C1308 vdd.n308 gnd 0.720658f
C1309 vdd.n309 gnd 0.009099f
C1310 vdd.n310 gnd 0.009099f
C1311 vdd.n311 gnd 0.009099f
C1312 vdd.n312 gnd 0.009099f
C1313 vdd.n313 gnd 0.007324f
C1314 vdd.n314 gnd 0.009099f
C1315 vdd.t11 gnd 0.46494f
C1316 vdd.n315 gnd 0.009099f
C1317 vdd.n316 gnd 0.009099f
C1318 vdd.n317 gnd 0.009099f
C1319 vdd.n318 gnd 0.929881f
C1320 vdd.n319 gnd 0.009099f
C1321 vdd.n320 gnd 0.009099f
C1322 vdd.n321 gnd 0.009099f
C1323 vdd.n322 gnd 0.009099f
C1324 vdd.n323 gnd 0.009099f
C1325 vdd.n324 gnd 0.007324f
C1326 vdd.n325 gnd 0.009099f
C1327 vdd.n326 gnd 0.009099f
C1328 vdd.n327 gnd 0.009099f
C1329 vdd.n328 gnd 0.022175f
C1330 vdd.n329 gnd 2.22242f
C1331 vdd.n330 gnd 0.022684f
C1332 vdd.n331 gnd 0.009099f
C1333 vdd.n332 gnd 0.009099f
C1334 vdd.n334 gnd 0.009099f
C1335 vdd.n335 gnd 0.009099f
C1336 vdd.n336 gnd 0.007324f
C1337 vdd.n337 gnd 0.007324f
C1338 vdd.n338 gnd 0.009099f
C1339 vdd.n339 gnd 0.009099f
C1340 vdd.n340 gnd 0.009099f
C1341 vdd.n341 gnd 0.009099f
C1342 vdd.n342 gnd 0.009099f
C1343 vdd.n343 gnd 0.009099f
C1344 vdd.n344 gnd 0.007324f
C1345 vdd.n346 gnd 0.009099f
C1346 vdd.n347 gnd 0.009099f
C1347 vdd.n348 gnd 0.009099f
C1348 vdd.n349 gnd 0.009099f
C1349 vdd.n350 gnd 0.009099f
C1350 vdd.n351 gnd 0.007324f
C1351 vdd.n353 gnd 0.009099f
C1352 vdd.n354 gnd 0.009099f
C1353 vdd.n355 gnd 0.009099f
C1354 vdd.n356 gnd 0.009099f
C1355 vdd.n357 gnd 0.009099f
C1356 vdd.n358 gnd 0.007324f
C1357 vdd.n360 gnd 0.009099f
C1358 vdd.n361 gnd 0.009099f
C1359 vdd.n362 gnd 0.009099f
C1360 vdd.n363 gnd 0.009099f
C1361 vdd.n364 gnd 0.006115f
C1362 vdd.t96 gnd 0.111942f
C1363 vdd.t95 gnd 0.119636f
C1364 vdd.t94 gnd 0.146195f
C1365 vdd.n365 gnd 0.187402f
C1366 vdd.n366 gnd 0.158184f
C1367 vdd.n368 gnd 0.009099f
C1368 vdd.n369 gnd 0.009099f
C1369 vdd.n370 gnd 0.007324f
C1370 vdd.n371 gnd 0.009099f
C1371 vdd.n373 gnd 0.009099f
C1372 vdd.n374 gnd 0.009099f
C1373 vdd.n375 gnd 0.009099f
C1374 vdd.n376 gnd 0.009099f
C1375 vdd.n377 gnd 0.007324f
C1376 vdd.n379 gnd 0.009099f
C1377 vdd.n380 gnd 0.009099f
C1378 vdd.n381 gnd 0.009099f
C1379 vdd.n382 gnd 0.009099f
C1380 vdd.n383 gnd 0.009099f
C1381 vdd.n384 gnd 0.007324f
C1382 vdd.n386 gnd 0.009099f
C1383 vdd.n387 gnd 0.009099f
C1384 vdd.n388 gnd 0.009099f
C1385 vdd.n389 gnd 0.009099f
C1386 vdd.n390 gnd 0.009099f
C1387 vdd.n391 gnd 0.007324f
C1388 vdd.n393 gnd 0.009099f
C1389 vdd.n394 gnd 0.009099f
C1390 vdd.n395 gnd 0.009099f
C1391 vdd.n396 gnd 0.009099f
C1392 vdd.n397 gnd 0.009099f
C1393 vdd.n398 gnd 0.007324f
C1394 vdd.n400 gnd 0.009099f
C1395 vdd.n401 gnd 0.009099f
C1396 vdd.n402 gnd 0.009099f
C1397 vdd.n403 gnd 0.009099f
C1398 vdd.n404 gnd 0.00725f
C1399 vdd.t90 gnd 0.111942f
C1400 vdd.t89 gnd 0.119636f
C1401 vdd.t87 gnd 0.146195f
C1402 vdd.n405 gnd 0.187402f
C1403 vdd.n406 gnd 0.158184f
C1404 vdd.n408 gnd 0.009099f
C1405 vdd.n409 gnd 0.009099f
C1406 vdd.n410 gnd 0.007324f
C1407 vdd.n411 gnd 0.009099f
C1408 vdd.n413 gnd 0.009099f
C1409 vdd.n414 gnd 0.009099f
C1410 vdd.n415 gnd 0.009099f
C1411 vdd.n416 gnd 0.009099f
C1412 vdd.n417 gnd 0.007324f
C1413 vdd.n419 gnd 0.009099f
C1414 vdd.n420 gnd 0.009099f
C1415 vdd.n421 gnd 0.009099f
C1416 vdd.n422 gnd 0.009099f
C1417 vdd.n423 gnd 0.009099f
C1418 vdd.n424 gnd 0.007324f
C1419 vdd.n426 gnd 0.009099f
C1420 vdd.n427 gnd 0.009099f
C1421 vdd.n428 gnd 0.009099f
C1422 vdd.n429 gnd 0.009099f
C1423 vdd.n430 gnd 0.009099f
C1424 vdd.n431 gnd 0.007324f
C1425 vdd.n433 gnd 0.009099f
C1426 vdd.n434 gnd 0.009099f
C1427 vdd.n435 gnd 0.009099f
C1428 vdd.n436 gnd 0.009099f
C1429 vdd.n437 gnd 0.009099f
C1430 vdd.n438 gnd 0.007324f
C1431 vdd.n440 gnd 0.009099f
C1432 vdd.n441 gnd 0.009099f
C1433 vdd.n442 gnd 0.009099f
C1434 vdd.n443 gnd 0.009099f
C1435 vdd.n444 gnd 0.009099f
C1436 vdd.n445 gnd 0.009099f
C1437 vdd.n446 gnd 0.007324f
C1438 vdd.n447 gnd 0.009099f
C1439 vdd.n448 gnd 0.009099f
C1440 vdd.n449 gnd 0.007324f
C1441 vdd.n450 gnd 0.009099f
C1442 vdd.n451 gnd 0.007324f
C1443 vdd.n452 gnd 0.009099f
C1444 vdd.n453 gnd 0.007324f
C1445 vdd.n454 gnd 0.009099f
C1446 vdd.n455 gnd 0.009099f
C1447 vdd.n456 gnd 0.506785f
C1448 vdd.t7 gnd 0.46494f
C1449 vdd.n457 gnd 0.009099f
C1450 vdd.n458 gnd 0.007324f
C1451 vdd.n459 gnd 0.009099f
C1452 vdd.n460 gnd 0.007324f
C1453 vdd.n461 gnd 0.009099f
C1454 vdd.t32 gnd 0.46494f
C1455 vdd.n462 gnd 0.009099f
C1456 vdd.n463 gnd 0.007324f
C1457 vdd.n464 gnd 0.009099f
C1458 vdd.n465 gnd 0.007324f
C1459 vdd.n466 gnd 0.009099f
C1460 vdd.t3 gnd 0.46494f
C1461 vdd.n467 gnd 0.581176f
C1462 vdd.n468 gnd 0.009099f
C1463 vdd.n469 gnd 0.007324f
C1464 vdd.n470 gnd 0.009099f
C1465 vdd.n471 gnd 0.007324f
C1466 vdd.n472 gnd 0.009099f
C1467 vdd.n473 gnd 0.929881f
C1468 vdd.n474 gnd 0.009099f
C1469 vdd.n475 gnd 0.007324f
C1470 vdd.n476 gnd 0.022175f
C1471 vdd.n477 gnd 0.006079f
C1472 vdd.n478 gnd 0.022175f
C1473 vdd.t66 gnd 0.46494f
C1474 vdd.n479 gnd 0.022175f
C1475 vdd.n480 gnd 0.006079f
C1476 vdd.n481 gnd 0.007825f
C1477 vdd.n482 gnd 0.007324f
C1478 vdd.n483 gnd 0.009099f
C1479 vdd.n484 gnd 6.40688f
C1480 vdd.n515 gnd 0.022684f
C1481 vdd.n516 gnd 1.27859f
C1482 vdd.n517 gnd 0.009099f
C1483 vdd.n518 gnd 0.007324f
C1484 vdd.n519 gnd 0.005823f
C1485 vdd.n520 gnd 0.014868f
C1486 vdd.n521 gnd 0.007324f
C1487 vdd.n522 gnd 0.009099f
C1488 vdd.n523 gnd 0.009099f
C1489 vdd.n524 gnd 0.009099f
C1490 vdd.n525 gnd 0.009099f
C1491 vdd.n526 gnd 0.009099f
C1492 vdd.n527 gnd 0.009099f
C1493 vdd.n528 gnd 0.009099f
C1494 vdd.n529 gnd 0.009099f
C1495 vdd.n530 gnd 0.009099f
C1496 vdd.n531 gnd 0.009099f
C1497 vdd.n532 gnd 0.009099f
C1498 vdd.n533 gnd 0.009099f
C1499 vdd.n534 gnd 0.009099f
C1500 vdd.n535 gnd 0.009099f
C1501 vdd.n536 gnd 0.006115f
C1502 vdd.n537 gnd 0.009099f
C1503 vdd.n538 gnd 0.009099f
C1504 vdd.n539 gnd 0.009099f
C1505 vdd.n540 gnd 0.009099f
C1506 vdd.n541 gnd 0.009099f
C1507 vdd.n542 gnd 0.009099f
C1508 vdd.n543 gnd 0.009099f
C1509 vdd.n544 gnd 0.009099f
C1510 vdd.n545 gnd 0.009099f
C1511 vdd.n546 gnd 0.009099f
C1512 vdd.n547 gnd 0.009099f
C1513 vdd.n548 gnd 0.009099f
C1514 vdd.n549 gnd 0.009099f
C1515 vdd.n550 gnd 0.009099f
C1516 vdd.n551 gnd 0.009099f
C1517 vdd.n552 gnd 0.009099f
C1518 vdd.n553 gnd 0.009099f
C1519 vdd.n554 gnd 0.009099f
C1520 vdd.n555 gnd 0.009099f
C1521 vdd.n556 gnd 0.00725f
C1522 vdd.t67 gnd 0.111942f
C1523 vdd.t68 gnd 0.119636f
C1524 vdd.t65 gnd 0.146195f
C1525 vdd.n557 gnd 0.187402f
C1526 vdd.n558 gnd 0.157451f
C1527 vdd.n559 gnd 0.009099f
C1528 vdd.n560 gnd 0.009099f
C1529 vdd.n561 gnd 0.009099f
C1530 vdd.n562 gnd 0.009099f
C1531 vdd.n563 gnd 0.009099f
C1532 vdd.n564 gnd 0.009099f
C1533 vdd.n565 gnd 0.009099f
C1534 vdd.n566 gnd 0.009099f
C1535 vdd.n567 gnd 0.009099f
C1536 vdd.n568 gnd 0.009099f
C1537 vdd.n569 gnd 0.009099f
C1538 vdd.n570 gnd 0.009099f
C1539 vdd.n571 gnd 0.009099f
C1540 vdd.n572 gnd 0.005823f
C1541 vdd.n575 gnd 0.006187f
C1542 vdd.n576 gnd 0.006187f
C1543 vdd.n577 gnd 0.006187f
C1544 vdd.n578 gnd 0.006187f
C1545 vdd.n579 gnd 0.006187f
C1546 vdd.n580 gnd 0.006187f
C1547 vdd.n582 gnd 0.006187f
C1548 vdd.n583 gnd 0.006187f
C1549 vdd.n585 gnd 0.006187f
C1550 vdd.n586 gnd 0.004504f
C1551 vdd.n588 gnd 0.006187f
C1552 vdd.t111 gnd 0.25003f
C1553 vdd.t110 gnd 0.255937f
C1554 vdd.t109 gnd 0.163229f
C1555 vdd.n589 gnd 0.088216f
C1556 vdd.n590 gnd 0.050039f
C1557 vdd.n591 gnd 0.008843f
C1558 vdd.n592 gnd 0.014461f
C1559 vdd.n594 gnd 0.006187f
C1560 vdd.n595 gnd 0.632319f
C1561 vdd.n596 gnd 0.013708f
C1562 vdd.n597 gnd 0.013708f
C1563 vdd.n598 gnd 0.006187f
C1564 vdd.n599 gnd 0.014682f
C1565 vdd.n600 gnd 0.006187f
C1566 vdd.n601 gnd 0.006187f
C1567 vdd.n602 gnd 0.006187f
C1568 vdd.n603 gnd 0.006187f
C1569 vdd.n604 gnd 0.006187f
C1570 vdd.n606 gnd 0.006187f
C1571 vdd.n607 gnd 0.006187f
C1572 vdd.n609 gnd 0.006187f
C1573 vdd.n610 gnd 0.006187f
C1574 vdd.n612 gnd 0.006187f
C1575 vdd.n613 gnd 0.006187f
C1576 vdd.n615 gnd 0.006187f
C1577 vdd.n616 gnd 0.006187f
C1578 vdd.n618 gnd 0.006187f
C1579 vdd.n619 gnd 0.006187f
C1580 vdd.n621 gnd 0.006187f
C1581 vdd.t104 gnd 0.25003f
C1582 vdd.t103 gnd 0.255937f
C1583 vdd.t101 gnd 0.163229f
C1584 vdd.n622 gnd 0.088216f
C1585 vdd.n623 gnd 0.050039f
C1586 vdd.n624 gnd 0.006187f
C1587 vdd.n626 gnd 0.006187f
C1588 vdd.n627 gnd 0.006187f
C1589 vdd.t102 gnd 0.316159f
C1590 vdd.n628 gnd 0.006187f
C1591 vdd.n629 gnd 0.006187f
C1592 vdd.n630 gnd 0.006187f
C1593 vdd.n631 gnd 0.006187f
C1594 vdd.n632 gnd 0.006187f
C1595 vdd.n633 gnd 0.632319f
C1596 vdd.n634 gnd 0.006187f
C1597 vdd.n635 gnd 0.006187f
C1598 vdd.n636 gnd 0.553279f
C1599 vdd.n637 gnd 0.006187f
C1600 vdd.n638 gnd 0.006187f
C1601 vdd.n639 gnd 0.005459f
C1602 vdd.n640 gnd 0.006187f
C1603 vdd.n641 gnd 0.557929f
C1604 vdd.n642 gnd 0.006187f
C1605 vdd.n643 gnd 0.006187f
C1606 vdd.n644 gnd 0.006187f
C1607 vdd.n645 gnd 0.006187f
C1608 vdd.n646 gnd 0.006187f
C1609 vdd.n647 gnd 0.632319f
C1610 vdd.n648 gnd 0.006187f
C1611 vdd.n649 gnd 0.006187f
C1612 vdd.t81 gnd 0.283614f
C1613 vdd.t179 gnd 0.074391f
C1614 vdd.n650 gnd 0.006187f
C1615 vdd.n651 gnd 0.006187f
C1616 vdd.n652 gnd 0.006187f
C1617 vdd.t182 gnd 0.316159f
C1618 vdd.n653 gnd 0.006187f
C1619 vdd.n654 gnd 0.006187f
C1620 vdd.n655 gnd 0.006187f
C1621 vdd.n656 gnd 0.006187f
C1622 vdd.n657 gnd 0.006187f
C1623 vdd.t185 gnd 0.316159f
C1624 vdd.n658 gnd 0.006187f
C1625 vdd.n659 gnd 0.006187f
C1626 vdd.n660 gnd 0.525383f
C1627 vdd.n661 gnd 0.006187f
C1628 vdd.n662 gnd 0.006187f
C1629 vdd.n663 gnd 0.006187f
C1630 vdd.n664 gnd 0.385901f
C1631 vdd.n665 gnd 0.006187f
C1632 vdd.n666 gnd 0.006187f
C1633 vdd.t187 gnd 0.316159f
C1634 vdd.n667 gnd 0.006187f
C1635 vdd.n668 gnd 0.006187f
C1636 vdd.n669 gnd 0.006187f
C1637 vdd.n670 gnd 0.525383f
C1638 vdd.n671 gnd 0.006187f
C1639 vdd.n672 gnd 0.006187f
C1640 vdd.t156 gnd 0.269665f
C1641 vdd.t198 gnd 0.246418f
C1642 vdd.n673 gnd 0.006187f
C1643 vdd.n674 gnd 0.006187f
C1644 vdd.n675 gnd 0.006187f
C1645 vdd.t157 gnd 0.316159f
C1646 vdd.n676 gnd 0.006187f
C1647 vdd.n677 gnd 0.006187f
C1648 vdd.t153 gnd 0.316159f
C1649 vdd.n678 gnd 0.006187f
C1650 vdd.n679 gnd 0.006187f
C1651 vdd.n680 gnd 0.006187f
C1652 vdd.t186 gnd 0.23247f
C1653 vdd.n681 gnd 0.006187f
C1654 vdd.n682 gnd 0.006187f
C1655 vdd.n683 gnd 0.539331f
C1656 vdd.n684 gnd 0.006187f
C1657 vdd.n685 gnd 0.006187f
C1658 vdd.n686 gnd 0.006187f
C1659 vdd.n687 gnd 0.632319f
C1660 vdd.n688 gnd 0.006187f
C1661 vdd.n689 gnd 0.006187f
C1662 vdd.t143 gnd 0.283614f
C1663 vdd.n690 gnd 0.399849f
C1664 vdd.n691 gnd 0.006187f
C1665 vdd.n692 gnd 0.006187f
C1666 vdd.n693 gnd 0.006187f
C1667 vdd.t180 gnd 0.316159f
C1668 vdd.n694 gnd 0.006187f
C1669 vdd.n695 gnd 0.006187f
C1670 vdd.n696 gnd 0.006187f
C1671 vdd.n697 gnd 0.006187f
C1672 vdd.n698 gnd 0.006187f
C1673 vdd.t195 gnd 0.632319f
C1674 vdd.n699 gnd 0.006187f
C1675 vdd.n700 gnd 0.006187f
C1676 vdd.t106 gnd 0.316159f
C1677 vdd.n701 gnd 0.006187f
C1678 vdd.n702 gnd 0.014682f
C1679 vdd.n703 gnd 0.014682f
C1680 vdd.t154 gnd 0.595124f
C1681 vdd.n704 gnd 0.013708f
C1682 vdd.n705 gnd 0.013708f
C1683 vdd.n706 gnd 0.014682f
C1684 vdd.n707 gnd 0.006187f
C1685 vdd.n708 gnd 0.006187f
C1686 vdd.t191 gnd 0.595124f
C1687 vdd.n726 gnd 0.014682f
C1688 vdd.n744 gnd 0.013708f
C1689 vdd.n745 gnd 0.006187f
C1690 vdd.n746 gnd 0.013708f
C1691 vdd.t131 gnd 0.25003f
C1692 vdd.t130 gnd 0.255937f
C1693 vdd.t129 gnd 0.163229f
C1694 vdd.n747 gnd 0.088216f
C1695 vdd.n748 gnd 0.050039f
C1696 vdd.n749 gnd 0.014461f
C1697 vdd.n750 gnd 0.006187f
C1698 vdd.t189 gnd 0.632319f
C1699 vdd.n751 gnd 0.013708f
C1700 vdd.n752 gnd 0.006187f
C1701 vdd.n753 gnd 0.014682f
C1702 vdd.n754 gnd 0.006187f
C1703 vdd.t100 gnd 0.25003f
C1704 vdd.t99 gnd 0.255937f
C1705 vdd.t97 gnd 0.163229f
C1706 vdd.n755 gnd 0.088216f
C1707 vdd.n756 gnd 0.050039f
C1708 vdd.n757 gnd 0.008843f
C1709 vdd.n758 gnd 0.006187f
C1710 vdd.n759 gnd 0.006187f
C1711 vdd.t98 gnd 0.316159f
C1712 vdd.n760 gnd 0.006187f
C1713 vdd.n761 gnd 0.006187f
C1714 vdd.n762 gnd 0.006187f
C1715 vdd.n763 gnd 0.006187f
C1716 vdd.n764 gnd 0.006187f
C1717 vdd.n765 gnd 0.006187f
C1718 vdd.n766 gnd 0.632319f
C1719 vdd.n767 gnd 0.006187f
C1720 vdd.n768 gnd 0.006187f
C1721 vdd.t183 gnd 0.316159f
C1722 vdd.n769 gnd 0.006187f
C1723 vdd.n770 gnd 0.006187f
C1724 vdd.n771 gnd 0.006187f
C1725 vdd.n772 gnd 0.006187f
C1726 vdd.n773 gnd 0.399849f
C1727 vdd.n774 gnd 0.006187f
C1728 vdd.n775 gnd 0.006187f
C1729 vdd.n776 gnd 0.006187f
C1730 vdd.n777 gnd 0.006187f
C1731 vdd.n778 gnd 0.006187f
C1732 vdd.n779 gnd 0.539331f
C1733 vdd.n780 gnd 0.006187f
C1734 vdd.n781 gnd 0.006187f
C1735 vdd.t193 gnd 0.283614f
C1736 vdd.t197 gnd 0.23247f
C1737 vdd.n782 gnd 0.006187f
C1738 vdd.n783 gnd 0.006187f
C1739 vdd.n784 gnd 0.006187f
C1740 vdd.t0 gnd 0.316159f
C1741 vdd.n785 gnd 0.006187f
C1742 vdd.n786 gnd 0.006187f
C1743 vdd.t177 gnd 0.316159f
C1744 vdd.n787 gnd 0.006187f
C1745 vdd.n788 gnd 0.006187f
C1746 vdd.n789 gnd 0.006187f
C1747 vdd.t149 gnd 0.246418f
C1748 vdd.n790 gnd 0.006187f
C1749 vdd.n791 gnd 0.006187f
C1750 vdd.n792 gnd 0.525383f
C1751 vdd.n793 gnd 0.006187f
C1752 vdd.n794 gnd 0.006187f
C1753 vdd.n795 gnd 0.006187f
C1754 vdd.t151 gnd 0.316159f
C1755 vdd.n796 gnd 0.006187f
C1756 vdd.n797 gnd 0.006187f
C1757 vdd.t159 gnd 0.269665f
C1758 vdd.n798 gnd 0.385901f
C1759 vdd.n799 gnd 0.006187f
C1760 vdd.n800 gnd 0.006187f
C1761 vdd.n801 gnd 0.006187f
C1762 vdd.n802 gnd 0.525383f
C1763 vdd.n803 gnd 0.006187f
C1764 vdd.n804 gnd 0.006187f
C1765 vdd.t145 gnd 0.316159f
C1766 vdd.n805 gnd 0.006187f
C1767 vdd.n806 gnd 0.006187f
C1768 vdd.n807 gnd 0.006187f
C1769 vdd.n808 gnd 0.632319f
C1770 vdd.n809 gnd 0.006187f
C1771 vdd.n810 gnd 0.006187f
C1772 vdd.t146 gnd 0.316159f
C1773 vdd.n811 gnd 0.006187f
C1774 vdd.n812 gnd 0.006187f
C1775 vdd.n813 gnd 0.006187f
C1776 vdd.t176 gnd 0.074391f
C1777 vdd.n814 gnd 0.006187f
C1778 vdd.n815 gnd 0.006187f
C1779 vdd.n816 gnd 0.006187f
C1780 vdd.t118 gnd 0.255937f
C1781 vdd.t116 gnd 0.163229f
C1782 vdd.t119 gnd 0.255937f
C1783 vdd.n817 gnd 0.143847f
C1784 vdd.n818 gnd 0.006187f
C1785 vdd.n819 gnd 0.006187f
C1786 vdd.n820 gnd 0.632319f
C1787 vdd.n821 gnd 0.006187f
C1788 vdd.n822 gnd 0.006187f
C1789 vdd.t117 gnd 0.283614f
C1790 vdd.n823 gnd 0.557929f
C1791 vdd.n824 gnd 0.006187f
C1792 vdd.n825 gnd 0.006187f
C1793 vdd.n826 gnd 0.006187f
C1794 vdd.n827 gnd 0.553279f
C1795 vdd.n828 gnd 0.006187f
C1796 vdd.n829 gnd 0.006187f
C1797 vdd.n830 gnd 0.006187f
C1798 vdd.n831 gnd 0.006187f
C1799 vdd.n832 gnd 0.006187f
C1800 vdd.n833 gnd 0.632319f
C1801 vdd.n834 gnd 0.006187f
C1802 vdd.n835 gnd 0.006187f
C1803 vdd.t113 gnd 0.316159f
C1804 vdd.n836 gnd 0.006187f
C1805 vdd.n837 gnd 0.014682f
C1806 vdd.n838 gnd 0.014682f
C1807 vdd.n839 gnd 6.40688f
C1808 vdd.n840 gnd 0.013708f
C1809 vdd.n841 gnd 0.013708f
C1810 vdd.n842 gnd 0.014682f
C1811 vdd.n843 gnd 0.006187f
C1812 vdd.n844 gnd 0.006187f
C1813 vdd.n845 gnd 0.006187f
C1814 vdd.n846 gnd 0.006187f
C1815 vdd.n847 gnd 0.006187f
C1816 vdd.n848 gnd 0.006187f
C1817 vdd.n849 gnd 0.006187f
C1818 vdd.n850 gnd 0.006187f
C1819 vdd.n852 gnd 0.006187f
C1820 vdd.n853 gnd 0.006187f
C1821 vdd.n854 gnd 0.005823f
C1822 vdd.n857 gnd 0.022684f
C1823 vdd.n858 gnd 0.007324f
C1824 vdd.n859 gnd 0.009099f
C1825 vdd.n861 gnd 0.009099f
C1826 vdd.n862 gnd 0.006079f
C1827 vdd.t73 gnd 0.46494f
C1828 vdd.n863 gnd 6.74164f
C1829 vdd.n864 gnd 0.009099f
C1830 vdd.n865 gnd 0.022684f
C1831 vdd.n866 gnd 0.007324f
C1832 vdd.n867 gnd 0.009099f
C1833 vdd.n868 gnd 0.007324f
C1834 vdd.n869 gnd 0.009099f
C1835 vdd.n870 gnd 0.929881f
C1836 vdd.n871 gnd 0.009099f
C1837 vdd.n872 gnd 0.007324f
C1838 vdd.n873 gnd 0.007324f
C1839 vdd.n874 gnd 0.009099f
C1840 vdd.n875 gnd 0.007324f
C1841 vdd.n876 gnd 0.009099f
C1842 vdd.t1 gnd 0.46494f
C1843 vdd.n877 gnd 0.009099f
C1844 vdd.n878 gnd 0.007324f
C1845 vdd.n879 gnd 0.009099f
C1846 vdd.n880 gnd 0.007324f
C1847 vdd.n881 gnd 0.009099f
C1848 vdd.t54 gnd 0.46494f
C1849 vdd.n882 gnd 0.009099f
C1850 vdd.n883 gnd 0.007324f
C1851 vdd.n884 gnd 0.009099f
C1852 vdd.n885 gnd 0.007324f
C1853 vdd.n886 gnd 0.009099f
C1854 vdd.n887 gnd 0.729956f
C1855 vdd.n888 gnd 0.771801f
C1856 vdd.t9 gnd 0.46494f
C1857 vdd.n889 gnd 0.009099f
C1858 vdd.n890 gnd 0.007324f
C1859 vdd.n891 gnd 0.004994f
C1860 vdd.n892 gnd 0.004634f
C1861 vdd.n893 gnd 0.002563f
C1862 vdd.n894 gnd 0.005886f
C1863 vdd.n895 gnd 0.00249f
C1864 vdd.n896 gnd 0.002637f
C1865 vdd.n897 gnd 0.004634f
C1866 vdd.n898 gnd 0.00249f
C1867 vdd.n899 gnd 0.005886f
C1868 vdd.n900 gnd 0.002637f
C1869 vdd.n901 gnd 0.004634f
C1870 vdd.n902 gnd 0.00249f
C1871 vdd.n903 gnd 0.004414f
C1872 vdd.n904 gnd 0.004427f
C1873 vdd.t2 gnd 0.012645f
C1874 vdd.n905 gnd 0.028134f
C1875 vdd.n906 gnd 0.146416f
C1876 vdd.n907 gnd 0.00249f
C1877 vdd.n908 gnd 0.002637f
C1878 vdd.n909 gnd 0.005886f
C1879 vdd.n910 gnd 0.005886f
C1880 vdd.n911 gnd 0.002637f
C1881 vdd.n912 gnd 0.00249f
C1882 vdd.n913 gnd 0.004634f
C1883 vdd.n914 gnd 0.004634f
C1884 vdd.n915 gnd 0.00249f
C1885 vdd.n916 gnd 0.002637f
C1886 vdd.n917 gnd 0.005886f
C1887 vdd.n918 gnd 0.005886f
C1888 vdd.n919 gnd 0.002637f
C1889 vdd.n920 gnd 0.00249f
C1890 vdd.n921 gnd 0.004634f
C1891 vdd.n922 gnd 0.004634f
C1892 vdd.n923 gnd 0.00249f
C1893 vdd.n924 gnd 0.002637f
C1894 vdd.n925 gnd 0.005886f
C1895 vdd.n926 gnd 0.005886f
C1896 vdd.n927 gnd 0.013915f
C1897 vdd.n928 gnd 0.002563f
C1898 vdd.n929 gnd 0.00249f
C1899 vdd.n930 gnd 0.011977f
C1900 vdd.n931 gnd 0.008362f
C1901 vdd.t28 gnd 0.029295f
C1902 vdd.t57 gnd 0.029295f
C1903 vdd.n932 gnd 0.201332f
C1904 vdd.n933 gnd 0.158317f
C1905 vdd.t17 gnd 0.029295f
C1906 vdd.t45 gnd 0.029295f
C1907 vdd.n934 gnd 0.201332f
C1908 vdd.n935 gnd 0.127761f
C1909 vdd.t23 gnd 0.029295f
C1910 vdd.t51 gnd 0.029295f
C1911 vdd.n936 gnd 0.201332f
C1912 vdd.n937 gnd 0.127761f
C1913 vdd.n938 gnd 0.004994f
C1914 vdd.n939 gnd 0.004634f
C1915 vdd.n940 gnd 0.002563f
C1916 vdd.n941 gnd 0.005886f
C1917 vdd.n942 gnd 0.00249f
C1918 vdd.n943 gnd 0.002637f
C1919 vdd.n944 gnd 0.004634f
C1920 vdd.n945 gnd 0.00249f
C1921 vdd.n946 gnd 0.005886f
C1922 vdd.n947 gnd 0.002637f
C1923 vdd.n948 gnd 0.004634f
C1924 vdd.n949 gnd 0.00249f
C1925 vdd.n950 gnd 0.004414f
C1926 vdd.n951 gnd 0.004427f
C1927 vdd.t61 gnd 0.012645f
C1928 vdd.n952 gnd 0.028134f
C1929 vdd.n953 gnd 0.146416f
C1930 vdd.n954 gnd 0.00249f
C1931 vdd.n955 gnd 0.002637f
C1932 vdd.n956 gnd 0.005886f
C1933 vdd.n957 gnd 0.005886f
C1934 vdd.n958 gnd 0.002637f
C1935 vdd.n959 gnd 0.00249f
C1936 vdd.n960 gnd 0.004634f
C1937 vdd.n961 gnd 0.004634f
C1938 vdd.n962 gnd 0.00249f
C1939 vdd.n963 gnd 0.002637f
C1940 vdd.n964 gnd 0.005886f
C1941 vdd.n965 gnd 0.005886f
C1942 vdd.n966 gnd 0.002637f
C1943 vdd.n967 gnd 0.00249f
C1944 vdd.n968 gnd 0.004634f
C1945 vdd.n969 gnd 0.004634f
C1946 vdd.n970 gnd 0.00249f
C1947 vdd.n971 gnd 0.002637f
C1948 vdd.n972 gnd 0.005886f
C1949 vdd.n973 gnd 0.005886f
C1950 vdd.n974 gnd 0.013915f
C1951 vdd.n975 gnd 0.002563f
C1952 vdd.n976 gnd 0.00249f
C1953 vdd.n977 gnd 0.011977f
C1954 vdd.n978 gnd 0.008099f
C1955 vdd.n979 gnd 0.095055f
C1956 vdd.n980 gnd 0.004994f
C1957 vdd.n981 gnd 0.004634f
C1958 vdd.n982 gnd 0.002563f
C1959 vdd.n983 gnd 0.005886f
C1960 vdd.n984 gnd 0.00249f
C1961 vdd.n985 gnd 0.002637f
C1962 vdd.n986 gnd 0.004634f
C1963 vdd.n987 gnd 0.00249f
C1964 vdd.n988 gnd 0.005886f
C1965 vdd.n989 gnd 0.002637f
C1966 vdd.n990 gnd 0.004634f
C1967 vdd.n991 gnd 0.00249f
C1968 vdd.n992 gnd 0.004414f
C1969 vdd.n993 gnd 0.004427f
C1970 vdd.t52 gnd 0.012645f
C1971 vdd.n994 gnd 0.028134f
C1972 vdd.n995 gnd 0.146416f
C1973 vdd.n996 gnd 0.00249f
C1974 vdd.n997 gnd 0.002637f
C1975 vdd.n998 gnd 0.005886f
C1976 vdd.n999 gnd 0.005886f
C1977 vdd.n1000 gnd 0.002637f
C1978 vdd.n1001 gnd 0.00249f
C1979 vdd.n1002 gnd 0.004634f
C1980 vdd.n1003 gnd 0.004634f
C1981 vdd.n1004 gnd 0.00249f
C1982 vdd.n1005 gnd 0.002637f
C1983 vdd.n1006 gnd 0.005886f
C1984 vdd.n1007 gnd 0.005886f
C1985 vdd.n1008 gnd 0.002637f
C1986 vdd.n1009 gnd 0.00249f
C1987 vdd.n1010 gnd 0.004634f
C1988 vdd.n1011 gnd 0.004634f
C1989 vdd.n1012 gnd 0.00249f
C1990 vdd.n1013 gnd 0.002637f
C1991 vdd.n1014 gnd 0.005886f
C1992 vdd.n1015 gnd 0.005886f
C1993 vdd.n1016 gnd 0.013915f
C1994 vdd.n1017 gnd 0.002563f
C1995 vdd.n1018 gnd 0.00249f
C1996 vdd.n1019 gnd 0.011977f
C1997 vdd.n1020 gnd 0.008362f
C1998 vdd.t10 gnd 0.029295f
C1999 vdd.t55 gnd 0.029295f
C2000 vdd.n1021 gnd 0.201332f
C2001 vdd.n1022 gnd 0.158317f
C2002 vdd.t50 gnd 0.029295f
C2003 vdd.t41 gnd 0.029295f
C2004 vdd.n1023 gnd 0.201332f
C2005 vdd.n1024 gnd 0.127761f
C2006 vdd.t26 gnd 0.029295f
C2007 vdd.t6 gnd 0.029295f
C2008 vdd.n1025 gnd 0.201332f
C2009 vdd.n1026 gnd 0.127761f
C2010 vdd.n1027 gnd 0.004994f
C2011 vdd.n1028 gnd 0.004634f
C2012 vdd.n1029 gnd 0.002563f
C2013 vdd.n1030 gnd 0.005886f
C2014 vdd.n1031 gnd 0.00249f
C2015 vdd.n1032 gnd 0.002637f
C2016 vdd.n1033 gnd 0.004634f
C2017 vdd.n1034 gnd 0.00249f
C2018 vdd.n1035 gnd 0.005886f
C2019 vdd.n1036 gnd 0.002637f
C2020 vdd.n1037 gnd 0.004634f
C2021 vdd.n1038 gnd 0.00249f
C2022 vdd.n1039 gnd 0.004414f
C2023 vdd.n1040 gnd 0.004427f
C2024 vdd.t39 gnd 0.012645f
C2025 vdd.n1041 gnd 0.028134f
C2026 vdd.n1042 gnd 0.146416f
C2027 vdd.n1043 gnd 0.00249f
C2028 vdd.n1044 gnd 0.002637f
C2029 vdd.n1045 gnd 0.005886f
C2030 vdd.n1046 gnd 0.005886f
C2031 vdd.n1047 gnd 0.002637f
C2032 vdd.n1048 gnd 0.00249f
C2033 vdd.n1049 gnd 0.004634f
C2034 vdd.n1050 gnd 0.004634f
C2035 vdd.n1051 gnd 0.00249f
C2036 vdd.n1052 gnd 0.002637f
C2037 vdd.n1053 gnd 0.005886f
C2038 vdd.n1054 gnd 0.005886f
C2039 vdd.n1055 gnd 0.002637f
C2040 vdd.n1056 gnd 0.00249f
C2041 vdd.n1057 gnd 0.004634f
C2042 vdd.n1058 gnd 0.004634f
C2043 vdd.n1059 gnd 0.00249f
C2044 vdd.n1060 gnd 0.002637f
C2045 vdd.n1061 gnd 0.005886f
C2046 vdd.n1062 gnd 0.005886f
C2047 vdd.n1063 gnd 0.013915f
C2048 vdd.n1064 gnd 0.002563f
C2049 vdd.n1065 gnd 0.00249f
C2050 vdd.n1066 gnd 0.011977f
C2051 vdd.n1067 gnd 0.008099f
C2052 vdd.n1068 gnd 0.056548f
C2053 vdd.n1069 gnd 0.203758f
C2054 vdd.n1070 gnd 0.004994f
C2055 vdd.n1071 gnd 0.004634f
C2056 vdd.n1072 gnd 0.002563f
C2057 vdd.n1073 gnd 0.005886f
C2058 vdd.n1074 gnd 0.00249f
C2059 vdd.n1075 gnd 0.002637f
C2060 vdd.n1076 gnd 0.004634f
C2061 vdd.n1077 gnd 0.00249f
C2062 vdd.n1078 gnd 0.005886f
C2063 vdd.n1079 gnd 0.002637f
C2064 vdd.n1080 gnd 0.004634f
C2065 vdd.n1081 gnd 0.00249f
C2066 vdd.n1082 gnd 0.004414f
C2067 vdd.n1083 gnd 0.004427f
C2068 vdd.t60 gnd 0.012645f
C2069 vdd.n1084 gnd 0.028134f
C2070 vdd.n1085 gnd 0.146416f
C2071 vdd.n1086 gnd 0.00249f
C2072 vdd.n1087 gnd 0.002637f
C2073 vdd.n1088 gnd 0.005886f
C2074 vdd.n1089 gnd 0.005886f
C2075 vdd.n1090 gnd 0.002637f
C2076 vdd.n1091 gnd 0.00249f
C2077 vdd.n1092 gnd 0.004634f
C2078 vdd.n1093 gnd 0.004634f
C2079 vdd.n1094 gnd 0.00249f
C2080 vdd.n1095 gnd 0.002637f
C2081 vdd.n1096 gnd 0.005886f
C2082 vdd.n1097 gnd 0.005886f
C2083 vdd.n1098 gnd 0.002637f
C2084 vdd.n1099 gnd 0.00249f
C2085 vdd.n1100 gnd 0.004634f
C2086 vdd.n1101 gnd 0.004634f
C2087 vdd.n1102 gnd 0.00249f
C2088 vdd.n1103 gnd 0.002637f
C2089 vdd.n1104 gnd 0.005886f
C2090 vdd.n1105 gnd 0.005886f
C2091 vdd.n1106 gnd 0.013915f
C2092 vdd.n1107 gnd 0.002563f
C2093 vdd.n1108 gnd 0.00249f
C2094 vdd.n1109 gnd 0.011977f
C2095 vdd.n1110 gnd 0.008362f
C2096 vdd.t15 gnd 0.029295f
C2097 vdd.t59 gnd 0.029295f
C2098 vdd.n1111 gnd 0.201332f
C2099 vdd.n1112 gnd 0.158317f
C2100 vdd.t58 gnd 0.029295f
C2101 vdd.t47 gnd 0.029295f
C2102 vdd.n1113 gnd 0.201332f
C2103 vdd.n1114 gnd 0.127761f
C2104 vdd.t34 gnd 0.029295f
C2105 vdd.t13 gnd 0.029295f
C2106 vdd.n1115 gnd 0.201332f
C2107 vdd.n1116 gnd 0.127761f
C2108 vdd.n1117 gnd 0.004994f
C2109 vdd.n1118 gnd 0.004634f
C2110 vdd.n1119 gnd 0.002563f
C2111 vdd.n1120 gnd 0.005886f
C2112 vdd.n1121 gnd 0.00249f
C2113 vdd.n1122 gnd 0.002637f
C2114 vdd.n1123 gnd 0.004634f
C2115 vdd.n1124 gnd 0.00249f
C2116 vdd.n1125 gnd 0.005886f
C2117 vdd.n1126 gnd 0.002637f
C2118 vdd.n1127 gnd 0.004634f
C2119 vdd.n1128 gnd 0.00249f
C2120 vdd.n1129 gnd 0.004414f
C2121 vdd.n1130 gnd 0.004427f
C2122 vdd.t46 gnd 0.012645f
C2123 vdd.n1131 gnd 0.028134f
C2124 vdd.n1132 gnd 0.146416f
C2125 vdd.n1133 gnd 0.00249f
C2126 vdd.n1134 gnd 0.002637f
C2127 vdd.n1135 gnd 0.005886f
C2128 vdd.n1136 gnd 0.005886f
C2129 vdd.n1137 gnd 0.002637f
C2130 vdd.n1138 gnd 0.00249f
C2131 vdd.n1139 gnd 0.004634f
C2132 vdd.n1140 gnd 0.004634f
C2133 vdd.n1141 gnd 0.00249f
C2134 vdd.n1142 gnd 0.002637f
C2135 vdd.n1143 gnd 0.005886f
C2136 vdd.n1144 gnd 0.005886f
C2137 vdd.n1145 gnd 0.002637f
C2138 vdd.n1146 gnd 0.00249f
C2139 vdd.n1147 gnd 0.004634f
C2140 vdd.n1148 gnd 0.004634f
C2141 vdd.n1149 gnd 0.00249f
C2142 vdd.n1150 gnd 0.002637f
C2143 vdd.n1151 gnd 0.005886f
C2144 vdd.n1152 gnd 0.005886f
C2145 vdd.n1153 gnd 0.013915f
C2146 vdd.n1154 gnd 0.002563f
C2147 vdd.n1155 gnd 0.00249f
C2148 vdd.n1156 gnd 0.011977f
C2149 vdd.n1157 gnd 0.008099f
C2150 vdd.n1158 gnd 0.056548f
C2151 vdd.n1159 gnd 0.220543f
C2152 vdd.n1160 gnd 1.8535f
C2153 vdd.n1161 gnd 0.536697f
C2154 vdd.n1162 gnd 0.007324f
C2155 vdd.n1163 gnd 0.009099f
C2156 vdd.n1164 gnd 0.571877f
C2157 vdd.n1165 gnd 0.009099f
C2158 vdd.n1166 gnd 0.007324f
C2159 vdd.n1167 gnd 0.009099f
C2160 vdd.n1168 gnd 0.007324f
C2161 vdd.n1169 gnd 0.009099f
C2162 vdd.t5 gnd 0.46494f
C2163 vdd.t16 gnd 0.46494f
C2164 vdd.n1170 gnd 0.009099f
C2165 vdd.n1171 gnd 0.007324f
C2166 vdd.n1172 gnd 0.009099f
C2167 vdd.n1173 gnd 0.007324f
C2168 vdd.n1174 gnd 0.009099f
C2169 vdd.t22 gnd 0.46494f
C2170 vdd.n1175 gnd 0.009099f
C2171 vdd.n1176 gnd 0.007324f
C2172 vdd.n1177 gnd 0.009099f
C2173 vdd.n1178 gnd 0.007324f
C2174 vdd.n1179 gnd 0.009099f
C2175 vdd.t38 gnd 0.46494f
C2176 vdd.n1180 gnd 0.674164f
C2177 vdd.n1181 gnd 0.009099f
C2178 vdd.n1182 gnd 0.007324f
C2179 vdd.n1183 gnd 0.009099f
C2180 vdd.n1184 gnd 0.007324f
C2181 vdd.n1185 gnd 0.009099f
C2182 vdd.n1186 gnd 0.929881f
C2183 vdd.n1187 gnd 0.009099f
C2184 vdd.n1188 gnd 0.007324f
C2185 vdd.n1189 gnd 0.022175f
C2186 vdd.n1190 gnd 0.006079f
C2187 vdd.n1191 gnd 0.022175f
C2188 vdd.t77 gnd 0.46494f
C2189 vdd.n1192 gnd 0.022175f
C2190 vdd.n1193 gnd 0.006079f
C2191 vdd.n1194 gnd 0.009099f
C2192 vdd.n1195 gnd 0.007324f
C2193 vdd.n1196 gnd 0.009099f
C2194 vdd.n1227 gnd 0.022684f
C2195 vdd.n1228 gnd 1.37157f
C2196 vdd.n1229 gnd 0.009099f
C2197 vdd.n1230 gnd 0.007324f
C2198 vdd.n1231 gnd 0.009099f
C2199 vdd.n1232 gnd 0.009099f
C2200 vdd.n1233 gnd 0.009099f
C2201 vdd.n1234 gnd 0.009099f
C2202 vdd.n1235 gnd 0.009099f
C2203 vdd.n1236 gnd 0.007324f
C2204 vdd.n1237 gnd 0.009099f
C2205 vdd.n1238 gnd 0.009099f
C2206 vdd.n1239 gnd 0.009099f
C2207 vdd.n1240 gnd 0.009099f
C2208 vdd.n1241 gnd 0.009099f
C2209 vdd.n1242 gnd 0.007324f
C2210 vdd.n1243 gnd 0.009099f
C2211 vdd.n1244 gnd 0.009099f
C2212 vdd.n1245 gnd 0.009099f
C2213 vdd.n1246 gnd 0.009099f
C2214 vdd.n1247 gnd 0.009099f
C2215 vdd.n1248 gnd 0.007324f
C2216 vdd.n1249 gnd 0.009099f
C2217 vdd.n1250 gnd 0.009099f
C2218 vdd.n1251 gnd 0.009099f
C2219 vdd.n1252 gnd 0.009099f
C2220 vdd.n1253 gnd 0.009099f
C2221 vdd.t127 gnd 0.111942f
C2222 vdd.t128 gnd 0.119636f
C2223 vdd.t126 gnd 0.146195f
C2224 vdd.n1254 gnd 0.187402f
C2225 vdd.n1255 gnd 0.158184f
C2226 vdd.n1256 gnd 0.015673f
C2227 vdd.n1257 gnd 0.009099f
C2228 vdd.n1258 gnd 0.009099f
C2229 vdd.n1259 gnd 0.009099f
C2230 vdd.n1260 gnd 0.009099f
C2231 vdd.n1261 gnd 0.009099f
C2232 vdd.n1262 gnd 0.007324f
C2233 vdd.n1263 gnd 0.009099f
C2234 vdd.n1264 gnd 0.009099f
C2235 vdd.n1265 gnd 0.009099f
C2236 vdd.n1266 gnd 0.009099f
C2237 vdd.n1267 gnd 0.009099f
C2238 vdd.n1268 gnd 0.007324f
C2239 vdd.n1269 gnd 0.009099f
C2240 vdd.n1270 gnd 0.009099f
C2241 vdd.n1271 gnd 0.009099f
C2242 vdd.n1272 gnd 0.009099f
C2243 vdd.n1273 gnd 0.009099f
C2244 vdd.n1274 gnd 0.007324f
C2245 vdd.n1275 gnd 0.009099f
C2246 vdd.n1276 gnd 0.009099f
C2247 vdd.n1277 gnd 0.009099f
C2248 vdd.n1278 gnd 0.009099f
C2249 vdd.n1279 gnd 0.009099f
C2250 vdd.n1280 gnd 0.007324f
C2251 vdd.n1281 gnd 0.009099f
C2252 vdd.n1282 gnd 0.009099f
C2253 vdd.n1283 gnd 0.009099f
C2254 vdd.n1284 gnd 0.009099f
C2255 vdd.n1285 gnd 0.009099f
C2256 vdd.n1286 gnd 0.007324f
C2257 vdd.n1287 gnd 0.009099f
C2258 vdd.n1288 gnd 0.009099f
C2259 vdd.n1289 gnd 0.009099f
C2260 vdd.n1290 gnd 0.009099f
C2261 vdd.n1291 gnd 0.007324f
C2262 vdd.n1292 gnd 0.009099f
C2263 vdd.n1293 gnd 0.009099f
C2264 vdd.n1294 gnd 0.009099f
C2265 vdd.n1295 gnd 0.009099f
C2266 vdd.n1296 gnd 0.009099f
C2267 vdd.n1297 gnd 0.007324f
C2268 vdd.n1298 gnd 0.009099f
C2269 vdd.n1299 gnd 0.009099f
C2270 vdd.n1300 gnd 0.009099f
C2271 vdd.n1301 gnd 0.009099f
C2272 vdd.n1302 gnd 0.009099f
C2273 vdd.n1303 gnd 0.007324f
C2274 vdd.n1304 gnd 0.009099f
C2275 vdd.n1305 gnd 0.009099f
C2276 vdd.n1306 gnd 0.009099f
C2277 vdd.n1307 gnd 0.009099f
C2278 vdd.n1308 gnd 0.009099f
C2279 vdd.n1309 gnd 0.007324f
C2280 vdd.n1310 gnd 0.009099f
C2281 vdd.n1311 gnd 0.009099f
C2282 vdd.n1312 gnd 0.009099f
C2283 vdd.n1313 gnd 0.009099f
C2284 vdd.n1314 gnd 0.009099f
C2285 vdd.n1315 gnd 0.007324f
C2286 vdd.n1316 gnd 0.009099f
C2287 vdd.n1317 gnd 0.009099f
C2288 vdd.n1318 gnd 0.009099f
C2289 vdd.n1319 gnd 0.009099f
C2290 vdd.t78 gnd 0.111942f
C2291 vdd.t79 gnd 0.119636f
C2292 vdd.t76 gnd 0.146195f
C2293 vdd.n1320 gnd 0.187402f
C2294 vdd.n1321 gnd 0.158184f
C2295 vdd.n1322 gnd 0.012011f
C2296 vdd.n1323 gnd 0.003479f
C2297 vdd.n1324 gnd 0.022684f
C2298 vdd.n1325 gnd 0.009099f
C2299 vdd.n1326 gnd 0.003845f
C2300 vdd.n1327 gnd 0.007324f
C2301 vdd.n1328 gnd 0.007324f
C2302 vdd.n1329 gnd 0.009099f
C2303 vdd.n1330 gnd 0.009099f
C2304 vdd.n1331 gnd 0.009099f
C2305 vdd.n1332 gnd 0.007324f
C2306 vdd.n1333 gnd 0.007324f
C2307 vdd.n1334 gnd 0.007324f
C2308 vdd.n1335 gnd 0.009099f
C2309 vdd.n1336 gnd 0.009099f
C2310 vdd.n1337 gnd 0.009099f
C2311 vdd.n1338 gnd 0.007324f
C2312 vdd.n1339 gnd 0.007324f
C2313 vdd.n1340 gnd 0.007324f
C2314 vdd.n1341 gnd 0.009099f
C2315 vdd.n1342 gnd 0.009099f
C2316 vdd.n1343 gnd 0.009099f
C2317 vdd.n1344 gnd 0.007324f
C2318 vdd.n1345 gnd 0.007324f
C2319 vdd.n1346 gnd 0.007324f
C2320 vdd.n1347 gnd 0.009099f
C2321 vdd.n1348 gnd 0.009099f
C2322 vdd.n1349 gnd 0.009099f
C2323 vdd.n1350 gnd 0.007324f
C2324 vdd.n1351 gnd 0.007324f
C2325 vdd.n1352 gnd 0.007324f
C2326 vdd.n1353 gnd 0.009099f
C2327 vdd.n1354 gnd 0.009099f
C2328 vdd.n1355 gnd 0.009099f
C2329 vdd.n1356 gnd 0.00725f
C2330 vdd.n1357 gnd 0.009099f
C2331 vdd.t124 gnd 0.111942f
C2332 vdd.t125 gnd 0.119636f
C2333 vdd.t123 gnd 0.146195f
C2334 vdd.n1358 gnd 0.187402f
C2335 vdd.n1359 gnd 0.158184f
C2336 vdd.n1360 gnd 0.015673f
C2337 vdd.n1361 gnd 0.00498f
C2338 vdd.n1362 gnd 0.009099f
C2339 vdd.n1363 gnd 0.009099f
C2340 vdd.n1364 gnd 0.009099f
C2341 vdd.n1365 gnd 0.007324f
C2342 vdd.n1366 gnd 0.007324f
C2343 vdd.n1367 gnd 0.007324f
C2344 vdd.n1368 gnd 0.009099f
C2345 vdd.n1369 gnd 0.009099f
C2346 vdd.n1370 gnd 0.009099f
C2347 vdd.n1371 gnd 0.007324f
C2348 vdd.n1372 gnd 0.007324f
C2349 vdd.n1373 gnd 0.007324f
C2350 vdd.n1374 gnd 0.009099f
C2351 vdd.n1375 gnd 0.009099f
C2352 vdd.n1376 gnd 0.009099f
C2353 vdd.n1377 gnd 0.007324f
C2354 vdd.n1378 gnd 0.007324f
C2355 vdd.n1379 gnd 0.007324f
C2356 vdd.n1380 gnd 0.009099f
C2357 vdd.n1381 gnd 0.009099f
C2358 vdd.n1382 gnd 0.009099f
C2359 vdd.n1383 gnd 0.007324f
C2360 vdd.n1384 gnd 0.007324f
C2361 vdd.n1385 gnd 0.007324f
C2362 vdd.n1386 gnd 0.009099f
C2363 vdd.n1387 gnd 0.009099f
C2364 vdd.n1388 gnd 0.009099f
C2365 vdd.n1389 gnd 0.007324f
C2366 vdd.n1390 gnd 0.007324f
C2367 vdd.n1391 gnd 0.006115f
C2368 vdd.n1392 gnd 0.009099f
C2369 vdd.n1393 gnd 0.009099f
C2370 vdd.n1394 gnd 0.009099f
C2371 vdd.n1395 gnd 0.006115f
C2372 vdd.n1396 gnd 0.007324f
C2373 vdd.n1397 gnd 0.007324f
C2374 vdd.n1398 gnd 0.009099f
C2375 vdd.n1399 gnd 0.009099f
C2376 vdd.n1400 gnd 0.009099f
C2377 vdd.n1401 gnd 0.007324f
C2378 vdd.n1402 gnd 0.007324f
C2379 vdd.n1403 gnd 0.007324f
C2380 vdd.n1404 gnd 0.009099f
C2381 vdd.n1405 gnd 0.009099f
C2382 vdd.n1406 gnd 0.009099f
C2383 vdd.n1407 gnd 0.007324f
C2384 vdd.n1408 gnd 0.007324f
C2385 vdd.n1409 gnd 0.007324f
C2386 vdd.n1410 gnd 0.009099f
C2387 vdd.n1411 gnd 0.009099f
C2388 vdd.n1412 gnd 0.009099f
C2389 vdd.n1413 gnd 0.007324f
C2390 vdd.n1414 gnd 0.007324f
C2391 vdd.n1415 gnd 0.007324f
C2392 vdd.n1416 gnd 0.009099f
C2393 vdd.n1417 gnd 0.009099f
C2394 vdd.n1418 gnd 0.009099f
C2395 vdd.n1419 gnd 0.007324f
C2396 vdd.n1420 gnd 0.009099f
C2397 vdd.n1421 gnd 2.22242f
C2398 vdd.n1423 gnd 0.022684f
C2399 vdd.n1424 gnd 0.006079f
C2400 vdd.n1425 gnd 0.022684f
C2401 vdd.n1426 gnd 0.022175f
C2402 vdd.n1427 gnd 0.009099f
C2403 vdd.n1428 gnd 0.007324f
C2404 vdd.n1429 gnd 0.009099f
C2405 vdd.n1430 gnd 0.488187f
C2406 vdd.n1431 gnd 0.009099f
C2407 vdd.n1432 gnd 0.007324f
C2408 vdd.n1433 gnd 0.009099f
C2409 vdd.n1434 gnd 0.009099f
C2410 vdd.n1435 gnd 0.009099f
C2411 vdd.n1436 gnd 0.007324f
C2412 vdd.n1437 gnd 0.009099f
C2413 vdd.n1438 gnd 0.832243f
C2414 vdd.n1439 gnd 0.929881f
C2415 vdd.n1440 gnd 0.009099f
C2416 vdd.n1441 gnd 0.007324f
C2417 vdd.n1442 gnd 0.009099f
C2418 vdd.n1443 gnd 0.009099f
C2419 vdd.n1444 gnd 0.009099f
C2420 vdd.n1445 gnd 0.007324f
C2421 vdd.n1446 gnd 0.009099f
C2422 vdd.n1447 gnd 0.562578f
C2423 vdd.n1448 gnd 0.009099f
C2424 vdd.n1449 gnd 0.007324f
C2425 vdd.n1450 gnd 0.009099f
C2426 vdd.n1451 gnd 0.009099f
C2427 vdd.n1452 gnd 0.009099f
C2428 vdd.n1453 gnd 0.007324f
C2429 vdd.n1454 gnd 0.009099f
C2430 vdd.n1455 gnd 0.516084f
C2431 vdd.n1456 gnd 0.720658f
C2432 vdd.n1457 gnd 0.009099f
C2433 vdd.n1458 gnd 0.007324f
C2434 vdd.n1459 gnd 0.009099f
C2435 vdd.n1460 gnd 0.009099f
C2436 vdd.n1461 gnd 0.006993f
C2437 vdd.n1462 gnd 0.009099f
C2438 vdd.n1463 gnd 0.007324f
C2439 vdd.n1464 gnd 0.009099f
C2440 vdd.n1465 gnd 0.771801f
C2441 vdd.n1466 gnd 0.009099f
C2442 vdd.n1467 gnd 0.007324f
C2443 vdd.n1468 gnd 0.009099f
C2444 vdd.n1469 gnd 0.009099f
C2445 vdd.n1470 gnd 0.009099f
C2446 vdd.n1471 gnd 0.007324f
C2447 vdd.n1472 gnd 0.009099f
C2448 vdd.t40 gnd 0.46494f
C2449 vdd.n1473 gnd 0.664865f
C2450 vdd.n1474 gnd 0.009099f
C2451 vdd.n1475 gnd 0.007324f
C2452 vdd.n1476 gnd 0.006993f
C2453 vdd.n1477 gnd 0.009099f
C2454 vdd.n1478 gnd 0.009099f
C2455 vdd.n1479 gnd 0.007324f
C2456 vdd.n1480 gnd 0.009099f
C2457 vdd.n1481 gnd 0.506785f
C2458 vdd.n1482 gnd 0.009099f
C2459 vdd.n1483 gnd 0.007324f
C2460 vdd.n1484 gnd 0.009099f
C2461 vdd.n1485 gnd 0.009099f
C2462 vdd.n1486 gnd 0.009099f
C2463 vdd.n1487 gnd 0.007324f
C2464 vdd.n1488 gnd 0.009099f
C2465 vdd.n1489 gnd 0.655566f
C2466 vdd.n1490 gnd 0.581176f
C2467 vdd.n1491 gnd 0.009099f
C2468 vdd.n1492 gnd 0.007324f
C2469 vdd.n1493 gnd 0.009099f
C2470 vdd.n1494 gnd 0.009099f
C2471 vdd.n1495 gnd 0.009099f
C2472 vdd.n1496 gnd 0.007324f
C2473 vdd.n1497 gnd 0.009099f
C2474 vdd.n1498 gnd 0.739255f
C2475 vdd.n1499 gnd 0.009099f
C2476 vdd.n1500 gnd 0.007324f
C2477 vdd.n1501 gnd 0.009099f
C2478 vdd.n1502 gnd 0.009099f
C2479 vdd.n1503 gnd 0.022175f
C2480 vdd.n1504 gnd 0.009099f
C2481 vdd.n1505 gnd 0.009099f
C2482 vdd.n1506 gnd 0.007324f
C2483 vdd.n1507 gnd 0.009099f
C2484 vdd.n1508 gnd 0.581176f
C2485 vdd.n1509 gnd 0.929881f
C2486 vdd.n1510 gnd 0.009099f
C2487 vdd.n1511 gnd 0.007324f
C2488 vdd.n1512 gnd 0.009099f
C2489 vdd.n1513 gnd 0.009099f
C2490 vdd.n1514 gnd 0.007825f
C2491 vdd.n1515 gnd 0.007324f
C2492 vdd.n1517 gnd 0.009099f
C2493 vdd.n1519 gnd 0.007324f
C2494 vdd.n1520 gnd 0.009099f
C2495 vdd.n1521 gnd 0.007324f
C2496 vdd.n1523 gnd 0.009099f
C2497 vdd.n1524 gnd 0.007324f
C2498 vdd.n1525 gnd 0.009099f
C2499 vdd.n1526 gnd 0.009099f
C2500 vdd.n1527 gnd 0.009099f
C2501 vdd.n1528 gnd 0.009099f
C2502 vdd.n1529 gnd 0.009099f
C2503 vdd.n1530 gnd 0.007324f
C2504 vdd.n1532 gnd 0.009099f
C2505 vdd.n1533 gnd 0.009099f
C2506 vdd.n1534 gnd 0.009099f
C2507 vdd.n1535 gnd 0.009099f
C2508 vdd.n1536 gnd 0.009099f
C2509 vdd.n1537 gnd 0.007324f
C2510 vdd.n1539 gnd 0.009099f
C2511 vdd.n1540 gnd 0.009099f
C2512 vdd.n1541 gnd 0.009099f
C2513 vdd.n1542 gnd 0.009099f
C2514 vdd.n1543 gnd 0.006115f
C2515 vdd.t93 gnd 0.111942f
C2516 vdd.t92 gnd 0.119636f
C2517 vdd.t91 gnd 0.146195f
C2518 vdd.n1544 gnd 0.187402f
C2519 vdd.n1545 gnd 0.157451f
C2520 vdd.n1547 gnd 0.009099f
C2521 vdd.n1548 gnd 0.009099f
C2522 vdd.n1549 gnd 0.007324f
C2523 vdd.n1550 gnd 0.009099f
C2524 vdd.n1552 gnd 0.009099f
C2525 vdd.n1553 gnd 0.009099f
C2526 vdd.n1554 gnd 0.009099f
C2527 vdd.n1555 gnd 0.009099f
C2528 vdd.n1556 gnd 0.007324f
C2529 vdd.n1558 gnd 0.009099f
C2530 vdd.n1559 gnd 0.009099f
C2531 vdd.n1560 gnd 0.009099f
C2532 vdd.n1561 gnd 0.009099f
C2533 vdd.n1562 gnd 0.009099f
C2534 vdd.n1563 gnd 0.007324f
C2535 vdd.n1565 gnd 0.009099f
C2536 vdd.n1566 gnd 0.009099f
C2537 vdd.n1567 gnd 0.009099f
C2538 vdd.n1568 gnd 0.009099f
C2539 vdd.n1569 gnd 0.009099f
C2540 vdd.n1570 gnd 0.007324f
C2541 vdd.n1572 gnd 0.009099f
C2542 vdd.n1573 gnd 0.009099f
C2543 vdd.n1574 gnd 0.009099f
C2544 vdd.n1575 gnd 0.009099f
C2545 vdd.n1576 gnd 0.009099f
C2546 vdd.n1577 gnd 0.007324f
C2547 vdd.n1579 gnd 0.009099f
C2548 vdd.n1580 gnd 0.009099f
C2549 vdd.n1581 gnd 0.009099f
C2550 vdd.n1582 gnd 0.009099f
C2551 vdd.n1583 gnd 0.00725f
C2552 vdd.t86 gnd 0.111942f
C2553 vdd.t85 gnd 0.119636f
C2554 vdd.t84 gnd 0.146195f
C2555 vdd.n1584 gnd 0.187402f
C2556 vdd.n1585 gnd 0.157451f
C2557 vdd.n1587 gnd 0.009099f
C2558 vdd.n1588 gnd 0.009099f
C2559 vdd.n1589 gnd 0.007324f
C2560 vdd.n1590 gnd 0.009099f
C2561 vdd.n1592 gnd 0.009099f
C2562 vdd.n1593 gnd 0.009099f
C2563 vdd.n1594 gnd 0.009099f
C2564 vdd.n1595 gnd 0.009099f
C2565 vdd.n1596 gnd 0.007324f
C2566 vdd.n1598 gnd 0.009099f
C2567 vdd.n1599 gnd 0.009099f
C2568 vdd.n1600 gnd 0.009099f
C2569 vdd.n1601 gnd 0.009099f
C2570 vdd.n1602 gnd 0.009099f
C2571 vdd.n1603 gnd 0.007324f
C2572 vdd.n1605 gnd 0.009099f
C2573 vdd.n1606 gnd 0.009099f
C2574 vdd.n1607 gnd 0.009099f
C2575 vdd.n1608 gnd 0.009099f
C2576 vdd.n1609 gnd 0.009099f
C2577 vdd.n1610 gnd 0.009099f
C2578 vdd.n1611 gnd 0.007324f
C2579 vdd.n1613 gnd 0.009099f
C2580 vdd.n1615 gnd 0.009099f
C2581 vdd.n1616 gnd 0.007324f
C2582 vdd.n1617 gnd 0.007324f
C2583 vdd.n1618 gnd 0.009099f
C2584 vdd.n1620 gnd 0.009099f
C2585 vdd.n1621 gnd 0.007324f
C2586 vdd.n1622 gnd 0.007324f
C2587 vdd.n1623 gnd 0.009099f
C2588 vdd.n1625 gnd 0.009099f
C2589 vdd.n1626 gnd 0.009099f
C2590 vdd.n1627 gnd 0.007324f
C2591 vdd.n1628 gnd 0.007324f
C2592 vdd.n1629 gnd 0.007324f
C2593 vdd.n1630 gnd 0.009099f
C2594 vdd.n1632 gnd 0.009099f
C2595 vdd.n1633 gnd 0.009099f
C2596 vdd.n1634 gnd 0.007324f
C2597 vdd.n1635 gnd 0.007324f
C2598 vdd.n1636 gnd 0.007324f
C2599 vdd.n1637 gnd 0.009099f
C2600 vdd.n1639 gnd 0.009099f
C2601 vdd.n1640 gnd 0.009099f
C2602 vdd.n1641 gnd 0.007324f
C2603 vdd.n1642 gnd 0.007324f
C2604 vdd.n1643 gnd 0.007324f
C2605 vdd.n1644 gnd 0.009099f
C2606 vdd.n1646 gnd 0.009099f
C2607 vdd.n1647 gnd 0.009099f
C2608 vdd.n1648 gnd 0.007324f
C2609 vdd.n1649 gnd 0.009099f
C2610 vdd.n1650 gnd 0.009099f
C2611 vdd.n1651 gnd 0.009099f
C2612 vdd.n1652 gnd 0.01494f
C2613 vdd.n1653 gnd 0.00498f
C2614 vdd.n1654 gnd 0.007324f
C2615 vdd.n1655 gnd 0.009099f
C2616 vdd.n1657 gnd 0.009099f
C2617 vdd.n1658 gnd 0.009099f
C2618 vdd.n1659 gnd 0.007324f
C2619 vdd.n1660 gnd 0.007324f
C2620 vdd.n1661 gnd 0.007324f
C2621 vdd.n1662 gnd 0.009099f
C2622 vdd.n1664 gnd 0.009099f
C2623 vdd.n1665 gnd 0.009099f
C2624 vdd.n1666 gnd 0.007324f
C2625 vdd.n1667 gnd 0.007324f
C2626 vdd.n1668 gnd 0.007324f
C2627 vdd.n1669 gnd 0.009099f
C2628 vdd.n1671 gnd 0.009099f
C2629 vdd.n1672 gnd 0.009099f
C2630 vdd.n1673 gnd 0.007324f
C2631 vdd.n1674 gnd 0.007324f
C2632 vdd.n1675 gnd 0.007324f
C2633 vdd.n1676 gnd 0.009099f
C2634 vdd.n1678 gnd 0.009099f
C2635 vdd.n1679 gnd 0.009099f
C2636 vdd.n1680 gnd 0.007324f
C2637 vdd.n1681 gnd 0.007324f
C2638 vdd.n1682 gnd 0.007324f
C2639 vdd.n1683 gnd 0.009099f
C2640 vdd.n1685 gnd 0.009099f
C2641 vdd.n1686 gnd 0.009099f
C2642 vdd.n1687 gnd 0.007324f
C2643 vdd.n1688 gnd 0.009099f
C2644 vdd.n1689 gnd 0.009099f
C2645 vdd.n1690 gnd 0.009099f
C2646 vdd.n1691 gnd 0.01494f
C2647 vdd.n1692 gnd 0.006115f
C2648 vdd.n1693 gnd 0.007324f
C2649 vdd.n1694 gnd 0.009099f
C2650 vdd.n1696 gnd 0.009099f
C2651 vdd.n1697 gnd 0.009099f
C2652 vdd.n1698 gnd 0.007324f
C2653 vdd.n1699 gnd 0.007324f
C2654 vdd.n1700 gnd 0.007324f
C2655 vdd.n1701 gnd 0.009099f
C2656 vdd.n1703 gnd 0.009099f
C2657 vdd.n1704 gnd 0.009099f
C2658 vdd.n1705 gnd 0.007324f
C2659 vdd.n1706 gnd 0.007324f
C2660 vdd.n1707 gnd 0.007324f
C2661 vdd.n1708 gnd 0.009099f
C2662 vdd.n1710 gnd 0.009099f
C2663 vdd.n1711 gnd 0.009099f
C2664 vdd.n1713 gnd 0.009099f
C2665 vdd.n1714 gnd 0.007324f
C2666 vdd.n1715 gnd 0.005823f
C2667 vdd.n1716 gnd 0.006187f
C2668 vdd.n1717 gnd 0.006187f
C2669 vdd.n1718 gnd 0.006187f
C2670 vdd.n1719 gnd 0.006187f
C2671 vdd.n1720 gnd 0.006187f
C2672 vdd.n1721 gnd 0.006187f
C2673 vdd.n1722 gnd 0.006187f
C2674 vdd.n1723 gnd 0.006187f
C2675 vdd.n1725 gnd 0.006187f
C2676 vdd.n1726 gnd 0.006187f
C2677 vdd.n1727 gnd 0.006187f
C2678 vdd.n1728 gnd 0.006187f
C2679 vdd.n1729 gnd 0.006187f
C2680 vdd.n1731 gnd 0.006187f
C2681 vdd.n1733 gnd 0.006187f
C2682 vdd.n1734 gnd 0.006187f
C2683 vdd.n1735 gnd 0.006187f
C2684 vdd.n1736 gnd 0.006187f
C2685 vdd.n1737 gnd 0.006187f
C2686 vdd.n1739 gnd 0.006187f
C2687 vdd.n1741 gnd 0.006187f
C2688 vdd.n1742 gnd 0.006187f
C2689 vdd.n1743 gnd 0.006187f
C2690 vdd.n1744 gnd 0.006187f
C2691 vdd.n1745 gnd 0.006187f
C2692 vdd.n1747 gnd 0.006187f
C2693 vdd.n1749 gnd 0.006187f
C2694 vdd.n1750 gnd 0.006187f
C2695 vdd.n1751 gnd 0.006187f
C2696 vdd.n1752 gnd 0.006187f
C2697 vdd.n1753 gnd 0.006187f
C2698 vdd.n1755 gnd 0.006187f
C2699 vdd.n1756 gnd 0.006187f
C2700 vdd.n1757 gnd 0.006187f
C2701 vdd.n1758 gnd 0.006187f
C2702 vdd.n1759 gnd 0.006187f
C2703 vdd.n1760 gnd 0.006187f
C2704 vdd.n1761 gnd 0.006187f
C2705 vdd.n1762 gnd 0.006187f
C2706 vdd.n1763 gnd 0.004504f
C2707 vdd.n1764 gnd 0.006187f
C2708 vdd.t139 gnd 0.25003f
C2709 vdd.t140 gnd 0.255937f
C2710 vdd.t138 gnd 0.163229f
C2711 vdd.n1765 gnd 0.088216f
C2712 vdd.n1766 gnd 0.050039f
C2713 vdd.n1767 gnd 0.008843f
C2714 vdd.n1768 gnd 0.006187f
C2715 vdd.n1769 gnd 0.006187f
C2716 vdd.n1770 gnd 0.376602f
C2717 vdd.n1771 gnd 0.006187f
C2718 vdd.n1772 gnd 0.006187f
C2719 vdd.n1773 gnd 0.006187f
C2720 vdd.n1774 gnd 0.006187f
C2721 vdd.n1775 gnd 0.006187f
C2722 vdd.n1776 gnd 0.006187f
C2723 vdd.n1777 gnd 0.006187f
C2724 vdd.n1778 gnd 0.006187f
C2725 vdd.n1779 gnd 0.006187f
C2726 vdd.n1780 gnd 0.006187f
C2727 vdd.n1781 gnd 0.006187f
C2728 vdd.n1782 gnd 0.006187f
C2729 vdd.n1783 gnd 0.006187f
C2730 vdd.n1784 gnd 0.006187f
C2731 vdd.n1785 gnd 0.006187f
C2732 vdd.n1786 gnd 0.006187f
C2733 vdd.n1787 gnd 0.006187f
C2734 vdd.n1788 gnd 0.006187f
C2735 vdd.n1789 gnd 0.006187f
C2736 vdd.n1790 gnd 0.006187f
C2737 vdd.t114 gnd 0.25003f
C2738 vdd.t115 gnd 0.255937f
C2739 vdd.t112 gnd 0.163229f
C2740 vdd.n1791 gnd 0.088216f
C2741 vdd.n1792 gnd 0.050039f
C2742 vdd.n1793 gnd 0.006187f
C2743 vdd.n1794 gnd 0.006187f
C2744 vdd.n1795 gnd 0.006187f
C2745 vdd.n1796 gnd 0.006187f
C2746 vdd.n1797 gnd 0.006187f
C2747 vdd.n1798 gnd 0.006187f
C2748 vdd.n1800 gnd 0.006187f
C2749 vdd.n1801 gnd 0.006187f
C2750 vdd.n1802 gnd 0.006187f
C2751 vdd.n1803 gnd 0.006187f
C2752 vdd.n1805 gnd 0.006187f
C2753 vdd.n1807 gnd 0.006187f
C2754 vdd.n1808 gnd 0.006187f
C2755 vdd.n1809 gnd 0.006187f
C2756 vdd.n1810 gnd 0.006187f
C2757 vdd.n1811 gnd 0.006187f
C2758 vdd.n1813 gnd 0.006187f
C2759 vdd.n1815 gnd 0.006187f
C2760 vdd.n1816 gnd 0.006187f
C2761 vdd.n1817 gnd 0.006187f
C2762 vdd.n1818 gnd 0.006187f
C2763 vdd.n1819 gnd 0.006187f
C2764 vdd.n1821 gnd 0.006187f
C2765 vdd.n1823 gnd 0.006187f
C2766 vdd.n1824 gnd 0.006187f
C2767 vdd.n1825 gnd 0.004504f
C2768 vdd.n1826 gnd 0.008843f
C2769 vdd.n1827 gnd 0.004777f
C2770 vdd.n1828 gnd 0.006187f
C2771 vdd.n1830 gnd 0.006187f
C2772 vdd.n1831 gnd 0.014682f
C2773 vdd.n1832 gnd 0.014682f
C2774 vdd.n1833 gnd 0.013708f
C2775 vdd.n1834 gnd 0.006187f
C2776 vdd.n1835 gnd 0.006187f
C2777 vdd.n1836 gnd 0.006187f
C2778 vdd.n1837 gnd 0.006187f
C2779 vdd.n1838 gnd 0.006187f
C2780 vdd.n1839 gnd 0.006187f
C2781 vdd.n1840 gnd 0.006187f
C2782 vdd.n1841 gnd 0.006187f
C2783 vdd.n1842 gnd 0.006187f
C2784 vdd.n1843 gnd 0.006187f
C2785 vdd.n1844 gnd 0.006187f
C2786 vdd.n1845 gnd 0.006187f
C2787 vdd.n1846 gnd 0.006187f
C2788 vdd.n1847 gnd 0.006187f
C2789 vdd.n1848 gnd 0.006187f
C2790 vdd.n1849 gnd 0.006187f
C2791 vdd.n1850 gnd 0.006187f
C2792 vdd.n1851 gnd 0.006187f
C2793 vdd.n1852 gnd 0.006187f
C2794 vdd.n1853 gnd 0.006187f
C2795 vdd.n1854 gnd 0.006187f
C2796 vdd.n1855 gnd 0.006187f
C2797 vdd.n1856 gnd 0.006187f
C2798 vdd.n1857 gnd 0.006187f
C2799 vdd.n1858 gnd 0.006187f
C2800 vdd.n1859 gnd 0.006187f
C2801 vdd.n1860 gnd 0.006187f
C2802 vdd.n1861 gnd 0.006187f
C2803 vdd.n1862 gnd 0.006187f
C2804 vdd.n1863 gnd 0.006187f
C2805 vdd.n1864 gnd 0.006187f
C2806 vdd.n1865 gnd 0.006187f
C2807 vdd.n1866 gnd 0.006187f
C2808 vdd.n1867 gnd 0.006187f
C2809 vdd.n1868 gnd 0.006187f
C2810 vdd.n1869 gnd 0.006187f
C2811 vdd.n1870 gnd 0.006187f
C2812 vdd.n1871 gnd 0.199924f
C2813 vdd.n1872 gnd 0.006187f
C2814 vdd.n1873 gnd 0.006187f
C2815 vdd.n1874 gnd 0.006187f
C2816 vdd.n1875 gnd 0.006187f
C2817 vdd.n1876 gnd 0.006187f
C2818 vdd.n1877 gnd 0.006187f
C2819 vdd.n1878 gnd 0.006187f
C2820 vdd.n1879 gnd 0.006187f
C2821 vdd.n1880 gnd 0.006187f
C2822 vdd.n1881 gnd 0.006187f
C2823 vdd.n1882 gnd 0.006187f
C2824 vdd.n1883 gnd 0.006187f
C2825 vdd.n1884 gnd 0.006187f
C2826 vdd.n1885 gnd 0.006187f
C2827 vdd.n1886 gnd 0.006187f
C2828 vdd.n1887 gnd 0.006187f
C2829 vdd.n1888 gnd 0.006187f
C2830 vdd.n1889 gnd 0.006187f
C2831 vdd.n1890 gnd 0.006187f
C2832 vdd.n1891 gnd 0.006187f
C2833 vdd.n1892 gnd 0.013708f
C2834 vdd.n1894 gnd 0.014682f
C2835 vdd.n1895 gnd 0.014682f
C2836 vdd.n1896 gnd 0.006187f
C2837 vdd.n1897 gnd 0.004777f
C2838 vdd.n1898 gnd 0.006187f
C2839 vdd.n1900 gnd 0.006187f
C2840 vdd.n1902 gnd 0.006187f
C2841 vdd.n1903 gnd 0.006187f
C2842 vdd.n1904 gnd 0.006187f
C2843 vdd.n1905 gnd 0.006187f
C2844 vdd.n1906 gnd 0.006187f
C2845 vdd.n1908 gnd 0.006187f
C2846 vdd.n1910 gnd 0.006187f
C2847 vdd.n1911 gnd 0.006187f
C2848 vdd.n1912 gnd 0.006187f
C2849 vdd.n1913 gnd 0.006187f
C2850 vdd.n1914 gnd 0.006187f
C2851 vdd.n1916 gnd 0.006187f
C2852 vdd.n1918 gnd 0.006187f
C2853 vdd.n1919 gnd 0.006187f
C2854 vdd.n1920 gnd 0.006187f
C2855 vdd.n1921 gnd 0.006187f
C2856 vdd.n1922 gnd 0.006187f
C2857 vdd.n1924 gnd 0.006187f
C2858 vdd.n1926 gnd 0.006187f
C2859 vdd.n1927 gnd 0.006187f
C2860 vdd.n1928 gnd 0.018456f
C2861 vdd.n1929 gnd 0.547103f
C2862 vdd.n1931 gnd 0.007324f
C2863 vdd.n1932 gnd 0.007324f
C2864 vdd.n1933 gnd 0.009099f
C2865 vdd.n1935 gnd 0.009099f
C2866 vdd.n1936 gnd 0.009099f
C2867 vdd.n1937 gnd 0.007324f
C2868 vdd.n1938 gnd 0.006079f
C2869 vdd.n1939 gnd 0.022684f
C2870 vdd.n1940 gnd 0.022175f
C2871 vdd.n1941 gnd 0.006079f
C2872 vdd.n1942 gnd 0.022175f
C2873 vdd.n1943 gnd 1.27859f
C2874 vdd.n1944 gnd 0.022175f
C2875 vdd.n1945 gnd 0.022684f
C2876 vdd.n1946 gnd 0.003479f
C2877 vdd.t75 gnd 0.111942f
C2878 vdd.t74 gnd 0.119636f
C2879 vdd.t72 gnd 0.146195f
C2880 vdd.n1947 gnd 0.187402f
C2881 vdd.n1948 gnd 0.157451f
C2882 vdd.n1949 gnd 0.011278f
C2883 vdd.n1950 gnd 0.003845f
C2884 vdd.n1951 gnd 0.007825f
C2885 vdd.n1952 gnd 0.547103f
C2886 vdd.n1953 gnd 0.018456f
C2887 vdd.n1954 gnd 0.006187f
C2888 vdd.n1955 gnd 0.006187f
C2889 vdd.n1956 gnd 0.006187f
C2890 vdd.n1958 gnd 0.006187f
C2891 vdd.n1960 gnd 0.006187f
C2892 vdd.n1961 gnd 0.006187f
C2893 vdd.n1962 gnd 0.006187f
C2894 vdd.n1963 gnd 0.006187f
C2895 vdd.n1964 gnd 0.006187f
C2896 vdd.n1966 gnd 0.006187f
C2897 vdd.n1968 gnd 0.006187f
C2898 vdd.n1969 gnd 0.006187f
C2899 vdd.n1970 gnd 0.006187f
C2900 vdd.n1971 gnd 0.006187f
C2901 vdd.n1972 gnd 0.006187f
C2902 vdd.n1974 gnd 0.006187f
C2903 vdd.n1976 gnd 0.006187f
C2904 vdd.n1977 gnd 0.006187f
C2905 vdd.n1978 gnd 0.006187f
C2906 vdd.n1979 gnd 0.006187f
C2907 vdd.n1980 gnd 0.006187f
C2908 vdd.n1982 gnd 0.006187f
C2909 vdd.n1984 gnd 0.006187f
C2910 vdd.n1985 gnd 0.006187f
C2911 vdd.n1986 gnd 0.014682f
C2912 vdd.n1987 gnd 0.013708f
C2913 vdd.n1988 gnd 0.013708f
C2914 vdd.n1989 gnd 0.911283f
C2915 vdd.n1990 gnd 0.013708f
C2916 vdd.n1991 gnd 0.013708f
C2917 vdd.n1992 gnd 0.006187f
C2918 vdd.n1993 gnd 0.006187f
C2919 vdd.n1994 gnd 0.006187f
C2920 vdd.n1995 gnd 0.395199f
C2921 vdd.n1996 gnd 0.006187f
C2922 vdd.n1997 gnd 0.006187f
C2923 vdd.n1998 gnd 0.006187f
C2924 vdd.n1999 gnd 0.006187f
C2925 vdd.n2000 gnd 0.006187f
C2926 vdd.n2001 gnd 0.632319f
C2927 vdd.n2002 gnd 0.006187f
C2928 vdd.n2003 gnd 0.006187f
C2929 vdd.n2004 gnd 0.006187f
C2930 vdd.n2005 gnd 0.006187f
C2931 vdd.n2006 gnd 0.006187f
C2932 vdd.n2007 gnd 0.632319f
C2933 vdd.n2008 gnd 0.006187f
C2934 vdd.n2009 gnd 0.006187f
C2935 vdd.n2010 gnd 0.005459f
C2936 vdd.n2011 gnd 0.017924f
C2937 vdd.n2012 gnd 0.003822f
C2938 vdd.n2013 gnd 0.006187f
C2939 vdd.n2014 gnd 0.348705f
C2940 vdd.n2015 gnd 0.006187f
C2941 vdd.n2016 gnd 0.006187f
C2942 vdd.n2017 gnd 0.006187f
C2943 vdd.n2018 gnd 0.006187f
C2944 vdd.n2019 gnd 0.006187f
C2945 vdd.n2020 gnd 0.423096f
C2946 vdd.n2021 gnd 0.006187f
C2947 vdd.n2022 gnd 0.006187f
C2948 vdd.n2023 gnd 0.006187f
C2949 vdd.n2024 gnd 0.006187f
C2950 vdd.n2025 gnd 0.006187f
C2951 vdd.n2026 gnd 0.562578f
C2952 vdd.n2027 gnd 0.006187f
C2953 vdd.n2028 gnd 0.006187f
C2954 vdd.n2029 gnd 0.006187f
C2955 vdd.n2030 gnd 0.006187f
C2956 vdd.n2031 gnd 0.006187f
C2957 vdd.n2032 gnd 0.502136f
C2958 vdd.n2033 gnd 0.006187f
C2959 vdd.n2034 gnd 0.006187f
C2960 vdd.n2035 gnd 0.006187f
C2961 vdd.n2036 gnd 0.006187f
C2962 vdd.n2037 gnd 0.006187f
C2963 vdd.n2038 gnd 0.362654f
C2964 vdd.n2039 gnd 0.006187f
C2965 vdd.n2040 gnd 0.006187f
C2966 vdd.n2041 gnd 0.006187f
C2967 vdd.n2042 gnd 0.006187f
C2968 vdd.n2043 gnd 0.006187f
C2969 vdd.n2044 gnd 0.199924f
C2970 vdd.n2045 gnd 0.006187f
C2971 vdd.n2046 gnd 0.006187f
C2972 vdd.n2047 gnd 0.006187f
C2973 vdd.n2048 gnd 0.006187f
C2974 vdd.n2049 gnd 0.006187f
C2975 vdd.n2050 gnd 0.348705f
C2976 vdd.n2051 gnd 0.006187f
C2977 vdd.n2052 gnd 0.006187f
C2978 vdd.n2053 gnd 0.006187f
C2979 vdd.n2054 gnd 0.006187f
C2980 vdd.n2055 gnd 0.006187f
C2981 vdd.n2056 gnd 0.632319f
C2982 vdd.n2057 gnd 0.006187f
C2983 vdd.n2058 gnd 0.006187f
C2984 vdd.n2059 gnd 0.006187f
C2985 vdd.n2060 gnd 0.006187f
C2986 vdd.n2061 gnd 0.006187f
C2987 vdd.n2062 gnd 0.006187f
C2988 vdd.n2063 gnd 0.006187f
C2989 vdd.n2064 gnd 0.492837f
C2990 vdd.n2065 gnd 0.006187f
C2991 vdd.n2066 gnd 0.006187f
C2992 vdd.n2067 gnd 0.006187f
C2993 vdd.n2068 gnd 0.006187f
C2994 vdd.n2069 gnd 0.006187f
C2995 vdd.n2070 gnd 0.006187f
C2996 vdd.n2071 gnd 0.395199f
C2997 vdd.n2072 gnd 0.006187f
C2998 vdd.n2073 gnd 0.006187f
C2999 vdd.n2074 gnd 0.006187f
C3000 vdd.n2075 gnd 0.014461f
C3001 vdd.n2076 gnd 0.013928f
C3002 vdd.n2077 gnd 0.006187f
C3003 vdd.n2078 gnd 0.006187f
C3004 vdd.n2079 gnd 0.004777f
C3005 vdd.n2080 gnd 0.006187f
C3006 vdd.n2081 gnd 0.006187f
C3007 vdd.n2082 gnd 0.004504f
C3008 vdd.n2083 gnd 0.006187f
C3009 vdd.n2084 gnd 0.006187f
C3010 vdd.n2085 gnd 0.006187f
C3011 vdd.n2086 gnd 0.006187f
C3012 vdd.n2087 gnd 0.006187f
C3013 vdd.n2088 gnd 0.006187f
C3014 vdd.n2089 gnd 0.006187f
C3015 vdd.n2090 gnd 0.006187f
C3016 vdd.n2091 gnd 0.006187f
C3017 vdd.n2092 gnd 0.006187f
C3018 vdd.n2093 gnd 0.006187f
C3019 vdd.n2094 gnd 0.006187f
C3020 vdd.n2095 gnd 0.006187f
C3021 vdd.n2096 gnd 0.006187f
C3022 vdd.n2097 gnd 0.006187f
C3023 vdd.n2098 gnd 0.006187f
C3024 vdd.n2099 gnd 0.006187f
C3025 vdd.n2100 gnd 0.006187f
C3026 vdd.n2101 gnd 0.006187f
C3027 vdd.n2102 gnd 0.006187f
C3028 vdd.n2103 gnd 0.006187f
C3029 vdd.n2104 gnd 0.006187f
C3030 vdd.n2105 gnd 0.006187f
C3031 vdd.n2106 gnd 0.006187f
C3032 vdd.n2107 gnd 0.006187f
C3033 vdd.n2108 gnd 0.006187f
C3034 vdd.n2109 gnd 0.006187f
C3035 vdd.n2110 gnd 0.006187f
C3036 vdd.n2111 gnd 0.006187f
C3037 vdd.n2112 gnd 0.006187f
C3038 vdd.n2113 gnd 0.006187f
C3039 vdd.n2114 gnd 0.006187f
C3040 vdd.n2115 gnd 0.006187f
C3041 vdd.n2116 gnd 0.006187f
C3042 vdd.n2117 gnd 0.006187f
C3043 vdd.n2118 gnd 0.006187f
C3044 vdd.n2119 gnd 0.006187f
C3045 vdd.n2120 gnd 0.006187f
C3046 vdd.n2121 gnd 0.006187f
C3047 vdd.n2122 gnd 0.006187f
C3048 vdd.n2123 gnd 0.006187f
C3049 vdd.n2124 gnd 0.006187f
C3050 vdd.n2125 gnd 0.006187f
C3051 vdd.n2126 gnd 0.006187f
C3052 vdd.n2127 gnd 0.006187f
C3053 vdd.n2128 gnd 0.006187f
C3054 vdd.n2129 gnd 0.006187f
C3055 vdd.n2130 gnd 0.006187f
C3056 vdd.n2131 gnd 0.006187f
C3057 vdd.n2132 gnd 0.006187f
C3058 vdd.n2133 gnd 0.006187f
C3059 vdd.n2134 gnd 0.006187f
C3060 vdd.n2135 gnd 0.006187f
C3061 vdd.n2136 gnd 0.006187f
C3062 vdd.n2137 gnd 0.006187f
C3063 vdd.n2138 gnd 0.006187f
C3064 vdd.n2139 gnd 0.006187f
C3065 vdd.n2140 gnd 0.006187f
C3066 vdd.n2141 gnd 0.006187f
C3067 vdd.n2142 gnd 0.006187f
C3068 vdd.n2143 gnd 0.014682f
C3069 vdd.n2144 gnd 0.013708f
C3070 vdd.n2145 gnd 0.013708f
C3071 vdd.n2146 gnd 0.771801f
C3072 vdd.n2147 gnd 0.013708f
C3073 vdd.n2148 gnd 0.014682f
C3074 vdd.n2149 gnd 0.013928f
C3075 vdd.n2150 gnd 0.006187f
C3076 vdd.n2151 gnd 0.006187f
C3077 vdd.n2152 gnd 0.006187f
C3078 vdd.n2153 gnd 0.004777f
C3079 vdd.n2154 gnd 0.008843f
C3080 vdd.n2155 gnd 0.004504f
C3081 vdd.n2156 gnd 0.006187f
C3082 vdd.n2157 gnd 0.006187f
C3083 vdd.n2158 gnd 0.006187f
C3084 vdd.n2159 gnd 0.006187f
C3085 vdd.n2160 gnd 0.006187f
C3086 vdd.n2161 gnd 0.006187f
C3087 vdd.n2162 gnd 0.006187f
C3088 vdd.n2163 gnd 0.006187f
C3089 vdd.n2164 gnd 0.006187f
C3090 vdd.n2165 gnd 0.006187f
C3091 vdd.n2166 gnd 0.006187f
C3092 vdd.n2167 gnd 0.006187f
C3093 vdd.n2168 gnd 0.006187f
C3094 vdd.n2169 gnd 0.006187f
C3095 vdd.n2170 gnd 0.006187f
C3096 vdd.n2171 gnd 0.006187f
C3097 vdd.n2172 gnd 0.006187f
C3098 vdd.n2173 gnd 0.006187f
C3099 vdd.n2174 gnd 0.006187f
C3100 vdd.n2175 gnd 0.006187f
C3101 vdd.n2176 gnd 0.006187f
C3102 vdd.n2177 gnd 0.006187f
C3103 vdd.n2178 gnd 0.006187f
C3104 vdd.n2179 gnd 0.006187f
C3105 vdd.n2180 gnd 0.006187f
C3106 vdd.n2181 gnd 0.006187f
C3107 vdd.n2182 gnd 0.006187f
C3108 vdd.n2183 gnd 0.006187f
C3109 vdd.n2184 gnd 0.006187f
C3110 vdd.n2185 gnd 0.006187f
C3111 vdd.n2186 gnd 0.006187f
C3112 vdd.n2187 gnd 0.006187f
C3113 vdd.n2188 gnd 0.006187f
C3114 vdd.n2189 gnd 0.006187f
C3115 vdd.n2190 gnd 0.006187f
C3116 vdd.n2191 gnd 0.006187f
C3117 vdd.n2192 gnd 0.006187f
C3118 vdd.n2193 gnd 0.006187f
C3119 vdd.n2194 gnd 0.006187f
C3120 vdd.n2195 gnd 0.006187f
C3121 vdd.n2196 gnd 0.006187f
C3122 vdd.n2197 gnd 0.006187f
C3123 vdd.n2198 gnd 0.006187f
C3124 vdd.n2199 gnd 0.006187f
C3125 vdd.n2200 gnd 0.006187f
C3126 vdd.n2201 gnd 0.006187f
C3127 vdd.n2202 gnd 0.006187f
C3128 vdd.n2203 gnd 0.006187f
C3129 vdd.n2204 gnd 0.006187f
C3130 vdd.n2205 gnd 0.006187f
C3131 vdd.n2206 gnd 0.006187f
C3132 vdd.n2207 gnd 0.006187f
C3133 vdd.n2208 gnd 0.006187f
C3134 vdd.n2209 gnd 0.006187f
C3135 vdd.n2210 gnd 0.006187f
C3136 vdd.n2211 gnd 0.006187f
C3137 vdd.n2212 gnd 0.006187f
C3138 vdd.n2213 gnd 0.006187f
C3139 vdd.n2214 gnd 0.006187f
C3140 vdd.n2215 gnd 0.006187f
C3141 vdd.n2216 gnd 0.014682f
C3142 vdd.n2217 gnd 0.014682f
C3143 vdd.n2218 gnd 0.771801f
C3144 vdd.t141 gnd 2.74315f
C3145 vdd.t147 gnd 2.74315f
C3146 vdd.n2251 gnd 0.014682f
C3147 vdd.n2252 gnd 0.006187f
C3148 vdd.t107 gnd 0.25003f
C3149 vdd.t108 gnd 0.255937f
C3150 vdd.t105 gnd 0.163229f
C3151 vdd.n2253 gnd 0.088216f
C3152 vdd.n2254 gnd 0.050039f
C3153 vdd.n2255 gnd 0.006187f
C3154 vdd.t121 gnd 0.25003f
C3155 vdd.t122 gnd 0.255937f
C3156 vdd.t120 gnd 0.163229f
C3157 vdd.n2256 gnd 0.088216f
C3158 vdd.n2257 gnd 0.050039f
C3159 vdd.n2258 gnd 0.008843f
C3160 vdd.n2259 gnd 0.006187f
C3161 vdd.n2260 gnd 0.006187f
C3162 vdd.n2261 gnd 0.006187f
C3163 vdd.n2262 gnd 0.006187f
C3164 vdd.n2263 gnd 0.006187f
C3165 vdd.n2264 gnd 0.006187f
C3166 vdd.n2265 gnd 0.006187f
C3167 vdd.n2266 gnd 0.006187f
C3168 vdd.n2267 gnd 0.006187f
C3169 vdd.n2268 gnd 0.006187f
C3170 vdd.n2269 gnd 0.006187f
C3171 vdd.n2270 gnd 0.006187f
C3172 vdd.n2271 gnd 0.006187f
C3173 vdd.n2272 gnd 0.006187f
C3174 vdd.n2273 gnd 0.006187f
C3175 vdd.n2274 gnd 0.006187f
C3176 vdd.n2275 gnd 0.006187f
C3177 vdd.n2276 gnd 0.006187f
C3178 vdd.n2277 gnd 0.006187f
C3179 vdd.n2278 gnd 0.006187f
C3180 vdd.n2279 gnd 0.006187f
C3181 vdd.n2280 gnd 0.006187f
C3182 vdd.n2281 gnd 0.006187f
C3183 vdd.n2282 gnd 0.006187f
C3184 vdd.n2283 gnd 0.006187f
C3185 vdd.n2284 gnd 0.006187f
C3186 vdd.n2285 gnd 0.006187f
C3187 vdd.n2286 gnd 0.006187f
C3188 vdd.n2287 gnd 0.006187f
C3189 vdd.n2288 gnd 0.006187f
C3190 vdd.n2289 gnd 0.006187f
C3191 vdd.n2290 gnd 0.006187f
C3192 vdd.n2291 gnd 0.006187f
C3193 vdd.n2292 gnd 0.006187f
C3194 vdd.n2293 gnd 0.006187f
C3195 vdd.n2294 gnd 0.006187f
C3196 vdd.n2295 gnd 0.006187f
C3197 vdd.n2296 gnd 0.006187f
C3198 vdd.n2297 gnd 0.006187f
C3199 vdd.n2298 gnd 0.006187f
C3200 vdd.n2299 gnd 0.006187f
C3201 vdd.n2300 gnd 0.006187f
C3202 vdd.n2301 gnd 0.006187f
C3203 vdd.n2302 gnd 0.006187f
C3204 vdd.n2303 gnd 0.006187f
C3205 vdd.n2304 gnd 0.006187f
C3206 vdd.n2305 gnd 0.006187f
C3207 vdd.n2306 gnd 0.006187f
C3208 vdd.n2307 gnd 0.006187f
C3209 vdd.n2308 gnd 0.006187f
C3210 vdd.n2309 gnd 0.006187f
C3211 vdd.n2310 gnd 0.006187f
C3212 vdd.n2311 gnd 0.006187f
C3213 vdd.n2312 gnd 0.006187f
C3214 vdd.n2313 gnd 0.006187f
C3215 vdd.n2314 gnd 0.006187f
C3216 vdd.n2315 gnd 0.004504f
C3217 vdd.n2316 gnd 0.006187f
C3218 vdd.n2317 gnd 0.006187f
C3219 vdd.n2318 gnd 0.004777f
C3220 vdd.n2319 gnd 0.006187f
C3221 vdd.n2320 gnd 0.006187f
C3222 vdd.n2321 gnd 0.014682f
C3223 vdd.n2322 gnd 0.013708f
C3224 vdd.n2323 gnd 0.006187f
C3225 vdd.n2324 gnd 0.006187f
C3226 vdd.n2325 gnd 0.006187f
C3227 vdd.n2326 gnd 0.006187f
C3228 vdd.n2327 gnd 0.006187f
C3229 vdd.n2328 gnd 0.006187f
C3230 vdd.n2329 gnd 0.006187f
C3231 vdd.n2330 gnd 0.006187f
C3232 vdd.n2331 gnd 0.006187f
C3233 vdd.n2332 gnd 0.006187f
C3234 vdd.n2333 gnd 0.006187f
C3235 vdd.n2334 gnd 0.006187f
C3236 vdd.n2335 gnd 0.006187f
C3237 vdd.n2336 gnd 0.006187f
C3238 vdd.n2337 gnd 0.006187f
C3239 vdd.n2338 gnd 0.006187f
C3240 vdd.n2339 gnd 0.006187f
C3241 vdd.n2340 gnd 0.006187f
C3242 vdd.n2341 gnd 0.006187f
C3243 vdd.n2342 gnd 0.006187f
C3244 vdd.n2343 gnd 0.006187f
C3245 vdd.n2344 gnd 0.006187f
C3246 vdd.n2345 gnd 0.006187f
C3247 vdd.n2346 gnd 0.006187f
C3248 vdd.n2347 gnd 0.006187f
C3249 vdd.n2348 gnd 0.006187f
C3250 vdd.n2349 gnd 0.006187f
C3251 vdd.n2350 gnd 0.006187f
C3252 vdd.n2351 gnd 0.006187f
C3253 vdd.n2352 gnd 0.006187f
C3254 vdd.n2353 gnd 0.006187f
C3255 vdd.n2354 gnd 0.006187f
C3256 vdd.n2355 gnd 0.006187f
C3257 vdd.n2356 gnd 0.006187f
C3258 vdd.n2357 gnd 0.006187f
C3259 vdd.n2358 gnd 0.006187f
C3260 vdd.n2359 gnd 0.006187f
C3261 vdd.n2360 gnd 0.006187f
C3262 vdd.n2361 gnd 0.006187f
C3263 vdd.n2362 gnd 0.006187f
C3264 vdd.n2363 gnd 0.006187f
C3265 vdd.n2364 gnd 0.006187f
C3266 vdd.n2365 gnd 0.006187f
C3267 vdd.n2366 gnd 0.006187f
C3268 vdd.n2367 gnd 0.006187f
C3269 vdd.n2368 gnd 0.006187f
C3270 vdd.n2369 gnd 0.006187f
C3271 vdd.n2370 gnd 0.006187f
C3272 vdd.n2371 gnd 0.006187f
C3273 vdd.n2372 gnd 0.006187f
C3274 vdd.n2373 gnd 0.006187f
C3275 vdd.n2374 gnd 0.199924f
C3276 vdd.n2375 gnd 0.006187f
C3277 vdd.n2376 gnd 0.006187f
C3278 vdd.n2377 gnd 0.006187f
C3279 vdd.n2378 gnd 0.006187f
C3280 vdd.n2379 gnd 0.006187f
C3281 vdd.n2380 gnd 0.006187f
C3282 vdd.n2381 gnd 0.006187f
C3283 vdd.n2382 gnd 0.006187f
C3284 vdd.n2383 gnd 0.006187f
C3285 vdd.n2384 gnd 0.006187f
C3286 vdd.n2385 gnd 0.006187f
C3287 vdd.n2386 gnd 0.006187f
C3288 vdd.n2387 gnd 0.006187f
C3289 vdd.n2388 gnd 0.006187f
C3290 vdd.n2389 gnd 0.006187f
C3291 vdd.n2390 gnd 0.006187f
C3292 vdd.n2391 gnd 0.006187f
C3293 vdd.n2392 gnd 0.006187f
C3294 vdd.n2393 gnd 0.006187f
C3295 vdd.n2394 gnd 0.006187f
C3296 vdd.n2395 gnd 0.376602f
C3297 vdd.n2396 gnd 0.006187f
C3298 vdd.n2397 gnd 0.006187f
C3299 vdd.n2398 gnd 0.006187f
C3300 vdd.n2399 gnd 0.006187f
C3301 vdd.n2400 gnd 0.006187f
C3302 vdd.n2401 gnd 0.013708f
C3303 vdd.n2402 gnd 0.014682f
C3304 vdd.n2403 gnd 0.014682f
C3305 vdd.n2404 gnd 0.006187f
C3306 vdd.n2405 gnd 0.006187f
C3307 vdd.n2406 gnd 0.006187f
C3308 vdd.n2407 gnd 0.004777f
C3309 vdd.n2408 gnd 0.008843f
C3310 vdd.n2409 gnd 0.004504f
C3311 vdd.n2410 gnd 0.006187f
C3312 vdd.n2411 gnd 0.006187f
C3313 vdd.n2412 gnd 0.006187f
C3314 vdd.n2413 gnd 0.006187f
C3315 vdd.n2414 gnd 0.006187f
C3316 vdd.n2415 gnd 0.006187f
C3317 vdd.n2416 gnd 0.006187f
C3318 vdd.n2417 gnd 0.006187f
C3319 vdd.n2418 gnd 0.006187f
C3320 vdd.n2419 gnd 0.006187f
C3321 vdd.n2420 gnd 0.006187f
C3322 vdd.n2421 gnd 0.006187f
C3323 vdd.n2422 gnd 0.006187f
C3324 vdd.n2423 gnd 0.006187f
C3325 vdd.n2424 gnd 0.006187f
C3326 vdd.n2425 gnd 0.006187f
C3327 vdd.n2426 gnd 0.006187f
C3328 vdd.n2427 gnd 0.006187f
C3329 vdd.n2428 gnd 0.006187f
C3330 vdd.n2429 gnd 0.006187f
C3331 vdd.n2430 gnd 0.006187f
C3332 vdd.n2431 gnd 0.006187f
C3333 vdd.n2432 gnd 0.006187f
C3334 vdd.n2433 gnd 0.006187f
C3335 vdd.n2434 gnd 0.006187f
C3336 vdd.n2435 gnd 0.006187f
C3337 vdd.n2436 gnd 0.006187f
C3338 vdd.n2437 gnd 0.006187f
C3339 vdd.n2438 gnd 0.006187f
C3340 vdd.n2439 gnd 0.006187f
C3341 vdd.n2440 gnd 0.006187f
C3342 vdd.n2441 gnd 0.006187f
C3343 vdd.n2442 gnd 0.006187f
C3344 vdd.n2443 gnd 0.006187f
C3345 vdd.n2444 gnd 0.006187f
C3346 vdd.n2445 gnd 0.006187f
C3347 vdd.n2446 gnd 0.006187f
C3348 vdd.n2447 gnd 0.006187f
C3349 vdd.n2448 gnd 0.006187f
C3350 vdd.n2449 gnd 0.006187f
C3351 vdd.n2450 gnd 0.006187f
C3352 vdd.n2451 gnd 0.006187f
C3353 vdd.n2452 gnd 0.006187f
C3354 vdd.n2453 gnd 0.006187f
C3355 vdd.n2454 gnd 0.006187f
C3356 vdd.n2455 gnd 0.006187f
C3357 vdd.n2456 gnd 0.006187f
C3358 vdd.n2457 gnd 0.006187f
C3359 vdd.n2458 gnd 0.006187f
C3360 vdd.n2459 gnd 0.006187f
C3361 vdd.n2460 gnd 0.006187f
C3362 vdd.n2461 gnd 0.006187f
C3363 vdd.n2462 gnd 0.006187f
C3364 vdd.n2463 gnd 0.006187f
C3365 vdd.n2464 gnd 0.006187f
C3366 vdd.n2465 gnd 0.006187f
C3367 vdd.n2466 gnd 0.006187f
C3368 vdd.n2467 gnd 0.006187f
C3369 vdd.n2468 gnd 0.006187f
C3370 vdd.n2469 gnd 0.006187f
C3371 vdd.n2471 gnd 0.771801f
C3372 vdd.n2473 gnd 0.006187f
C3373 vdd.n2474 gnd 0.006187f
C3374 vdd.n2475 gnd 0.014682f
C3375 vdd.n2476 gnd 0.013708f
C3376 vdd.n2477 gnd 0.013708f
C3377 vdd.n2478 gnd 0.771801f
C3378 vdd.n2479 gnd 0.013708f
C3379 vdd.n2480 gnd 0.013708f
C3380 vdd.n2481 gnd 0.006187f
C3381 vdd.n2482 gnd 0.006187f
C3382 vdd.n2483 gnd 0.006187f
C3383 vdd.n2484 gnd 0.395199f
C3384 vdd.n2485 gnd 0.006187f
C3385 vdd.n2486 gnd 0.006187f
C3386 vdd.n2487 gnd 0.006187f
C3387 vdd.n2488 gnd 0.006187f
C3388 vdd.n2489 gnd 0.006187f
C3389 vdd.n2490 gnd 0.492837f
C3390 vdd.n2491 gnd 0.006187f
C3391 vdd.n2492 gnd 0.006187f
C3392 vdd.n2493 gnd 0.006187f
C3393 vdd.n2494 gnd 0.006187f
C3394 vdd.n2495 gnd 0.006187f
C3395 vdd.n2496 gnd 0.632319f
C3396 vdd.n2497 gnd 0.006187f
C3397 vdd.n2498 gnd 0.006187f
C3398 vdd.n2499 gnd 0.006187f
C3399 vdd.n2500 gnd 0.006187f
C3400 vdd.n2501 gnd 0.006187f
C3401 vdd.n2502 gnd 0.348705f
C3402 vdd.n2503 gnd 0.006187f
C3403 vdd.n2504 gnd 0.006187f
C3404 vdd.n2505 gnd 0.006187f
C3405 vdd.n2506 gnd 0.006187f
C3406 vdd.n2507 gnd 0.006187f
C3407 vdd.n2508 gnd 0.199924f
C3408 vdd.n2509 gnd 0.006187f
C3409 vdd.n2510 gnd 0.006187f
C3410 vdd.n2511 gnd 0.006187f
C3411 vdd.n2512 gnd 0.006187f
C3412 vdd.n2513 gnd 0.006187f
C3413 vdd.n2514 gnd 0.362654f
C3414 vdd.n2515 gnd 0.006187f
C3415 vdd.n2516 gnd 0.006187f
C3416 vdd.n2517 gnd 0.006187f
C3417 vdd.n2518 gnd 0.006187f
C3418 vdd.n2519 gnd 0.006187f
C3419 vdd.n2520 gnd 0.502136f
C3420 vdd.n2521 gnd 0.006187f
C3421 vdd.n2522 gnd 0.006187f
C3422 vdd.n2523 gnd 0.006187f
C3423 vdd.n2524 gnd 0.006187f
C3424 vdd.n2525 gnd 0.006187f
C3425 vdd.n2526 gnd 0.562578f
C3426 vdd.n2527 gnd 0.006187f
C3427 vdd.n2528 gnd 0.006187f
C3428 vdd.n2529 gnd 0.006187f
C3429 vdd.n2530 gnd 0.006187f
C3430 vdd.n2531 gnd 0.006187f
C3431 vdd.n2532 gnd 0.423096f
C3432 vdd.n2533 gnd 0.006187f
C3433 vdd.n2534 gnd 0.006187f
C3434 vdd.n2535 gnd 0.006187f
C3435 vdd.t82 gnd 0.255937f
C3436 vdd.t80 gnd 0.163229f
C3437 vdd.t83 gnd 0.255937f
C3438 vdd.n2536 gnd 0.143847f
C3439 vdd.n2537 gnd 0.017924f
C3440 vdd.n2538 gnd 0.003822f
C3441 vdd.n2539 gnd 0.006187f
C3442 vdd.n2540 gnd 0.348705f
C3443 vdd.n2541 gnd 0.006187f
C3444 vdd.n2542 gnd 0.006187f
C3445 vdd.n2543 gnd 0.006187f
C3446 vdd.n2544 gnd 0.006187f
C3447 vdd.n2545 gnd 0.006187f
C3448 vdd.n2546 gnd 0.632319f
C3449 vdd.n2547 gnd 0.006187f
C3450 vdd.n2548 gnd 0.006187f
C3451 vdd.n2549 gnd 0.006187f
C3452 vdd.n2550 gnd 0.006187f
C3453 vdd.n2551 gnd 0.006187f
C3454 vdd.n2552 gnd 0.006187f
C3455 vdd.n2554 gnd 0.006187f
C3456 vdd.n2555 gnd 0.006187f
C3457 vdd.n2557 gnd 0.006187f
C3458 vdd.n2558 gnd 0.006187f
C3459 vdd.n2561 gnd 0.006187f
C3460 vdd.n2562 gnd 0.006187f
C3461 vdd.n2563 gnd 0.006187f
C3462 vdd.n2564 gnd 0.006187f
C3463 vdd.n2566 gnd 0.006187f
C3464 vdd.n2567 gnd 0.006187f
C3465 vdd.n2568 gnd 0.006187f
C3466 vdd.n2569 gnd 0.006187f
C3467 vdd.n2570 gnd 0.006187f
C3468 vdd.n2571 gnd 0.006187f
C3469 vdd.n2573 gnd 0.006187f
C3470 vdd.n2574 gnd 0.006187f
C3471 vdd.n2575 gnd 0.006187f
C3472 vdd.n2576 gnd 0.006187f
C3473 vdd.n2577 gnd 0.006187f
C3474 vdd.n2578 gnd 0.006187f
C3475 vdd.n2580 gnd 0.006187f
C3476 vdd.n2581 gnd 0.006187f
C3477 vdd.n2582 gnd 0.006187f
C3478 vdd.n2583 gnd 0.006187f
C3479 vdd.n2584 gnd 0.006187f
C3480 vdd.n2585 gnd 0.006187f
C3481 vdd.n2587 gnd 0.006187f
C3482 vdd.n2588 gnd 0.014682f
C3483 vdd.n2589 gnd 0.014682f
C3484 vdd.n2590 gnd 0.013708f
C3485 vdd.n2591 gnd 0.006187f
C3486 vdd.n2592 gnd 0.006187f
C3487 vdd.n2593 gnd 0.006187f
C3488 vdd.n2594 gnd 0.006187f
C3489 vdd.n2595 gnd 0.006187f
C3490 vdd.n2596 gnd 0.006187f
C3491 vdd.n2597 gnd 0.632319f
C3492 vdd.n2598 gnd 0.006187f
C3493 vdd.n2599 gnd 0.006187f
C3494 vdd.n2600 gnd 0.006187f
C3495 vdd.n2601 gnd 0.006187f
C3496 vdd.n2602 gnd 0.006187f
C3497 vdd.n2603 gnd 0.395199f
C3498 vdd.n2604 gnd 0.006187f
C3499 vdd.n2605 gnd 0.006187f
C3500 vdd.n2606 gnd 0.006187f
C3501 vdd.n2607 gnd 0.014461f
C3502 vdd.n2608 gnd 0.013928f
C3503 vdd.n2609 gnd 0.014682f
C3504 vdd.n2611 gnd 0.006187f
C3505 vdd.n2612 gnd 0.006187f
C3506 vdd.n2613 gnd 0.004777f
C3507 vdd.n2614 gnd 0.008843f
C3508 vdd.n2615 gnd 0.004504f
C3509 vdd.n2616 gnd 0.006187f
C3510 vdd.n2617 gnd 0.006187f
C3511 vdd.n2619 gnd 0.006187f
C3512 vdd.n2620 gnd 0.006187f
C3513 vdd.n2621 gnd 0.006187f
C3514 vdd.n2622 gnd 0.006187f
C3515 vdd.n2623 gnd 0.006187f
C3516 vdd.n2624 gnd 0.006187f
C3517 vdd.n2626 gnd 0.006187f
C3518 vdd.n2627 gnd 0.006187f
C3519 vdd.n2628 gnd 0.006187f
C3520 vdd.n2629 gnd 0.006187f
C3521 vdd.n2630 gnd 0.006187f
C3522 vdd.n2631 gnd 0.006187f
C3523 vdd.n2633 gnd 0.006187f
C3524 vdd.n2634 gnd 0.006187f
C3525 vdd.n2635 gnd 0.006187f
C3526 vdd.n2636 gnd 0.006187f
C3527 vdd.n2637 gnd 0.006187f
C3528 vdd.n2638 gnd 0.006187f
C3529 vdd.n2640 gnd 0.006187f
C3530 vdd.n2641 gnd 0.006187f
C3531 vdd.n2642 gnd 0.006187f
C3532 vdd.n2644 gnd 0.006187f
C3533 vdd.n2645 gnd 0.006187f
C3534 vdd.n2646 gnd 0.006187f
C3535 vdd.n2647 gnd 0.006187f
C3536 vdd.n2648 gnd 0.006187f
C3537 vdd.n2649 gnd 0.006187f
C3538 vdd.n2651 gnd 0.006187f
C3539 vdd.n2652 gnd 0.006187f
C3540 vdd.n2653 gnd 0.006187f
C3541 vdd.n2654 gnd 0.006187f
C3542 vdd.n2655 gnd 0.006187f
C3543 vdd.n2656 gnd 0.006187f
C3544 vdd.n2658 gnd 0.006187f
C3545 vdd.n2659 gnd 0.006187f
C3546 vdd.n2660 gnd 0.006187f
C3547 vdd.n2661 gnd 0.006187f
C3548 vdd.n2662 gnd 0.006187f
C3549 vdd.n2663 gnd 0.006187f
C3550 vdd.n2665 gnd 0.006187f
C3551 vdd.n2666 gnd 0.006187f
C3552 vdd.n2668 gnd 0.006187f
C3553 vdd.n2669 gnd 0.006187f
C3554 vdd.n2670 gnd 0.014682f
C3555 vdd.n2671 gnd 0.013708f
C3556 vdd.n2672 gnd 0.013708f
C3557 vdd.n2673 gnd 0.911283f
C3558 vdd.n2674 gnd 0.013708f
C3559 vdd.n2675 gnd 0.014682f
C3560 vdd.n2676 gnd 0.013928f
C3561 vdd.n2677 gnd 0.006187f
C3562 vdd.n2678 gnd 0.004777f
C3563 vdd.n2679 gnd 0.006187f
C3564 vdd.n2681 gnd 0.006187f
C3565 vdd.n2682 gnd 0.006187f
C3566 vdd.n2683 gnd 0.006187f
C3567 vdd.n2684 gnd 0.006187f
C3568 vdd.n2685 gnd 0.006187f
C3569 vdd.n2686 gnd 0.006187f
C3570 vdd.n2688 gnd 0.006187f
C3571 vdd.n2689 gnd 0.006187f
C3572 vdd.n2690 gnd 0.006187f
C3573 vdd.n2691 gnd 0.006187f
C3574 vdd.n2692 gnd 0.006187f
C3575 vdd.n2693 gnd 0.006187f
C3576 vdd.n2695 gnd 0.006187f
C3577 vdd.n2696 gnd 0.006187f
C3578 vdd.n2697 gnd 0.006187f
C3579 vdd.n2698 gnd 0.006187f
C3580 vdd.n2699 gnd 0.006187f
C3581 vdd.n2700 gnd 0.006187f
C3582 vdd.n2702 gnd 0.006187f
C3583 vdd.n2703 gnd 0.006187f
C3584 vdd.n2705 gnd 0.006187f
C3585 vdd.n2706 gnd 0.014868f
C3586 vdd.n2707 gnd 0.55069f
C3587 vdd.n2708 gnd 0.007825f
C3588 vdd.n2709 gnd 0.022684f
C3589 vdd.n2710 gnd 0.003479f
C3590 vdd.t133 gnd 0.111942f
C3591 vdd.t134 gnd 0.119636f
C3592 vdd.t132 gnd 0.146195f
C3593 vdd.n2711 gnd 0.187402f
C3594 vdd.n2712 gnd 0.157451f
C3595 vdd.n2713 gnd 0.011278f
C3596 vdd.n2714 gnd 0.009099f
C3597 vdd.n2715 gnd 0.003845f
C3598 vdd.n2716 gnd 0.007324f
C3599 vdd.n2717 gnd 0.009099f
C3600 vdd.n2718 gnd 0.009099f
C3601 vdd.n2719 gnd 0.007324f
C3602 vdd.n2720 gnd 0.007324f
C3603 vdd.n2721 gnd 0.009099f
C3604 vdd.n2722 gnd 0.009099f
C3605 vdd.n2723 gnd 0.007324f
C3606 vdd.n2724 gnd 0.007324f
C3607 vdd.n2725 gnd 0.009099f
C3608 vdd.n2726 gnd 0.009099f
C3609 vdd.n2727 gnd 0.007324f
C3610 vdd.n2728 gnd 0.007324f
C3611 vdd.n2729 gnd 0.009099f
C3612 vdd.n2730 gnd 0.009099f
C3613 vdd.n2731 gnd 0.007324f
C3614 vdd.n2732 gnd 0.007324f
C3615 vdd.n2733 gnd 0.009099f
C3616 vdd.n2734 gnd 0.009099f
C3617 vdd.n2735 gnd 0.007324f
C3618 vdd.n2736 gnd 0.007324f
C3619 vdd.n2737 gnd 0.009099f
C3620 vdd.n2738 gnd 0.009099f
C3621 vdd.n2739 gnd 0.007324f
C3622 vdd.n2740 gnd 0.007324f
C3623 vdd.n2741 gnd 0.009099f
C3624 vdd.n2742 gnd 0.009099f
C3625 vdd.n2743 gnd 0.007324f
C3626 vdd.n2744 gnd 0.007324f
C3627 vdd.n2745 gnd 0.009099f
C3628 vdd.n2746 gnd 0.009099f
C3629 vdd.n2747 gnd 0.007324f
C3630 vdd.n2748 gnd 0.007324f
C3631 vdd.n2749 gnd 0.009099f
C3632 vdd.n2750 gnd 0.009099f
C3633 vdd.n2751 gnd 0.007324f
C3634 vdd.n2752 gnd 0.009099f
C3635 vdd.n2753 gnd 0.009099f
C3636 vdd.n2754 gnd 0.007324f
C3637 vdd.n2755 gnd 0.009099f
C3638 vdd.n2756 gnd 0.009099f
C3639 vdd.n2757 gnd 0.009099f
C3640 vdd.n2758 gnd 0.01494f
C3641 vdd.n2759 gnd 0.009099f
C3642 vdd.n2760 gnd 0.009099f
C3643 vdd.n2761 gnd 0.00498f
C3644 vdd.n2762 gnd 0.007324f
C3645 vdd.n2763 gnd 0.009099f
C3646 vdd.n2764 gnd 0.009099f
C3647 vdd.n2765 gnd 0.007324f
C3648 vdd.n2766 gnd 0.007324f
C3649 vdd.n2767 gnd 0.009099f
C3650 vdd.n2768 gnd 0.009099f
C3651 vdd.n2769 gnd 0.007324f
C3652 vdd.n2770 gnd 0.007324f
C3653 vdd.n2771 gnd 0.009099f
C3654 vdd.n2772 gnd 0.009099f
C3655 vdd.n2773 gnd 0.007324f
C3656 vdd.n2774 gnd 0.007324f
C3657 vdd.n2775 gnd 0.009099f
C3658 vdd.n2776 gnd 0.009099f
C3659 vdd.n2777 gnd 0.007324f
C3660 vdd.n2778 gnd 0.007324f
C3661 vdd.n2779 gnd 0.009099f
C3662 vdd.n2780 gnd 0.009099f
C3663 vdd.n2781 gnd 0.007324f
C3664 vdd.n2782 gnd 0.007324f
C3665 vdd.n2783 gnd 0.009099f
C3666 vdd.n2784 gnd 0.009099f
C3667 vdd.n2785 gnd 0.007324f
C3668 vdd.n2786 gnd 0.007324f
C3669 vdd.n2787 gnd 0.009099f
C3670 vdd.n2788 gnd 0.009099f
C3671 vdd.n2789 gnd 0.007324f
C3672 vdd.n2790 gnd 0.007324f
C3673 vdd.n2791 gnd 0.009099f
C3674 vdd.n2792 gnd 0.009099f
C3675 vdd.n2793 gnd 0.007324f
C3676 vdd.n2794 gnd 0.007324f
C3677 vdd.n2795 gnd 0.009099f
C3678 vdd.n2796 gnd 0.009099f
C3679 vdd.n2797 gnd 0.007324f
C3680 vdd.n2798 gnd 0.009099f
C3681 vdd.n2799 gnd 0.009099f
C3682 vdd.n2800 gnd 0.007324f
C3683 vdd.n2801 gnd 0.009099f
C3684 vdd.n2802 gnd 0.009099f
C3685 vdd.n2803 gnd 0.009099f
C3686 vdd.t70 gnd 0.111942f
C3687 vdd.t71 gnd 0.119636f
C3688 vdd.t69 gnd 0.146195f
C3689 vdd.n2804 gnd 0.187402f
C3690 vdd.n2805 gnd 0.157451f
C3691 vdd.n2806 gnd 0.01494f
C3692 vdd.n2807 gnd 0.009099f
C3693 vdd.n2808 gnd 0.009099f
C3694 vdd.n2809 gnd 0.006115f
C3695 vdd.n2810 gnd 0.007324f
C3696 vdd.n2811 gnd 0.009099f
C3697 vdd.n2812 gnd 0.009099f
C3698 vdd.n2813 gnd 0.007324f
C3699 vdd.n2814 gnd 0.007324f
C3700 vdd.n2815 gnd 0.009099f
C3701 vdd.n2816 gnd 0.009099f
C3702 vdd.n2817 gnd 0.007324f
C3703 vdd.n2818 gnd 0.007324f
C3704 vdd.n2819 gnd 0.009099f
C3705 vdd.n2820 gnd 0.009099f
C3706 vdd.n2821 gnd 0.007324f
C3707 vdd.n2822 gnd 0.007324f
C3708 vdd.n2823 gnd 0.009099f
C3709 vdd.n2824 gnd 0.009099f
C3710 vdd.n2825 gnd 0.007324f
C3711 vdd.n2826 gnd 0.007324f
C3712 vdd.n2827 gnd 0.009099f
C3713 vdd.n2828 gnd 0.009099f
C3714 vdd.n2829 gnd 0.007324f
C3715 vdd.n2830 gnd 0.007324f
C3716 vdd.n2831 gnd 0.009099f
C3717 vdd.n2832 gnd 0.009099f
C3718 vdd.n2833 gnd 0.007324f
C3719 vdd.n2834 gnd 0.007324f
C3720 vdd.n2836 gnd 0.55069f
C3721 vdd.n2838 gnd 0.007324f
C3722 vdd.n2839 gnd 0.009099f
C3723 vdd.n2840 gnd 6.74164f
C3724 vdd.n2842 gnd 0.022684f
C3725 vdd.n2843 gnd 0.006079f
C3726 vdd.n2844 gnd 0.022684f
C3727 vdd.n2845 gnd 0.022175f
C3728 vdd.n2846 gnd 0.009099f
C3729 vdd.n2847 gnd 0.007324f
C3730 vdd.n2848 gnd 0.009099f
C3731 vdd.n2849 gnd 0.581176f
C3732 vdd.n2850 gnd 0.009099f
C3733 vdd.n2851 gnd 0.007324f
C3734 vdd.n2852 gnd 0.009099f
C3735 vdd.n2853 gnd 0.009099f
C3736 vdd.n2854 gnd 0.009099f
C3737 vdd.n2855 gnd 0.007324f
C3738 vdd.n2856 gnd 0.009099f
C3739 vdd.n2857 gnd 0.739255f
C3740 vdd.n2858 gnd 0.929881f
C3741 vdd.n2859 gnd 0.009099f
C3742 vdd.n2860 gnd 0.007324f
C3743 vdd.n2861 gnd 0.009099f
C3744 vdd.n2862 gnd 0.009099f
C3745 vdd.n2863 gnd 0.009099f
C3746 vdd.n2864 gnd 0.007324f
C3747 vdd.n2865 gnd 0.009099f
C3748 vdd.n2866 gnd 0.655566f
C3749 vdd.n2867 gnd 0.009099f
C3750 vdd.n2868 gnd 0.007324f
C3751 vdd.n2869 gnd 0.009099f
C3752 vdd.n2870 gnd 0.009099f
C3753 vdd.n2871 gnd 0.009099f
C3754 vdd.n2872 gnd 0.007324f
C3755 vdd.n2873 gnd 0.009099f
C3756 vdd.t29 gnd 0.46494f
C3757 vdd.n2874 gnd 0.771801f
C3758 vdd.n2875 gnd 0.009099f
C3759 vdd.n2876 gnd 0.007324f
C3760 vdd.n2877 gnd 0.009099f
C3761 vdd.n2878 gnd 0.009099f
C3762 vdd.n2879 gnd 0.009099f
C3763 vdd.n2880 gnd 0.007324f
C3764 vdd.n2881 gnd 0.009099f
C3765 vdd.n2882 gnd 0.729956f
C3766 vdd.n2883 gnd 0.009099f
C3767 vdd.n2884 gnd 0.007324f
C3768 vdd.n2885 gnd 0.009099f
C3769 vdd.n2886 gnd 0.009099f
C3770 vdd.n2887 gnd 0.009099f
C3771 vdd.n2888 gnd 0.007324f
C3772 vdd.n2889 gnd 0.007324f
C3773 vdd.n2890 gnd 0.007324f
C3774 vdd.n2891 gnd 0.009099f
C3775 vdd.n2892 gnd 0.009099f
C3776 vdd.n2893 gnd 0.009099f
C3777 vdd.n2894 gnd 0.007324f
C3778 vdd.n2895 gnd 0.007324f
C3779 vdd.n2896 gnd 0.007324f
C3780 vdd.n2897 gnd 0.009099f
C3781 vdd.n2898 gnd 0.009099f
C3782 vdd.n2899 gnd 0.009099f
C3783 vdd.n2900 gnd 0.007324f
C3784 vdd.n2901 gnd 0.007324f
C3785 vdd.n2902 gnd 0.006079f
C3786 vdd.n2903 gnd 0.022175f
C3787 vdd.n2904 gnd 0.022684f
C3788 vdd.n2906 gnd 0.022684f
C3789 vdd.n2907 gnd 0.003479f
C3790 vdd.t137 gnd 0.111942f
C3791 vdd.t136 gnd 0.119636f
C3792 vdd.t135 gnd 0.146195f
C3793 vdd.n2908 gnd 0.187402f
C3794 vdd.n2909 gnd 0.158184f
C3795 vdd.n2910 gnd 0.012011f
C3796 vdd.n2911 gnd 0.003845f
C3797 vdd.n2912 gnd 0.007324f
C3798 vdd.n2913 gnd 0.009099f
C3799 vdd.n2915 gnd 0.009099f
C3800 vdd.n2916 gnd 0.009099f
C3801 vdd.n2917 gnd 0.007324f
C3802 vdd.n2918 gnd 0.007324f
C3803 vdd.n2919 gnd 0.007324f
C3804 vdd.n2920 gnd 0.009099f
C3805 vdd.n2922 gnd 0.009099f
C3806 vdd.n2923 gnd 0.009099f
C3807 vdd.n2924 gnd 0.007324f
C3808 vdd.n2925 gnd 0.007324f
C3809 vdd.n2926 gnd 0.007324f
C3810 vdd.n2927 gnd 0.009099f
C3811 vdd.n2929 gnd 0.009099f
C3812 vdd.n2930 gnd 0.009099f
C3813 vdd.n2931 gnd 0.007324f
C3814 vdd.n2932 gnd 0.007324f
C3815 vdd.n2933 gnd 0.007324f
C3816 vdd.n2934 gnd 0.009099f
C3817 vdd.n2936 gnd 0.009099f
C3818 vdd.n2937 gnd 0.009099f
C3819 vdd.n2938 gnd 0.007324f
C3820 vdd.n2939 gnd 0.007324f
C3821 vdd.n2940 gnd 0.007324f
C3822 vdd.n2941 gnd 0.009099f
C3823 vdd.n2943 gnd 0.009099f
C3824 vdd.n2944 gnd 0.009099f
C3825 vdd.n2945 gnd 0.007324f
C3826 vdd.n2946 gnd 0.009099f
C3827 vdd.n2947 gnd 0.009099f
C3828 vdd.n2948 gnd 0.009099f
C3829 vdd.n2949 gnd 0.015673f
C3830 vdd.n2950 gnd 0.00498f
C3831 vdd.n2951 gnd 0.007324f
C3832 vdd.n2952 gnd 0.009099f
C3833 vdd.n2954 gnd 0.009099f
C3834 vdd.n2955 gnd 0.009099f
C3835 vdd.n2956 gnd 0.007324f
C3836 vdd.n2957 gnd 0.007324f
C3837 vdd.n2958 gnd 0.007324f
C3838 vdd.n2959 gnd 0.009099f
C3839 vdd.n2961 gnd 0.009099f
C3840 vdd.n2962 gnd 0.009099f
C3841 vdd.n2963 gnd 0.007324f
C3842 vdd.n2964 gnd 0.007324f
C3843 vdd.n2965 gnd 0.007324f
C3844 vdd.n2966 gnd 0.009099f
C3845 vdd.n2968 gnd 0.009099f
C3846 vdd.n2969 gnd 0.009099f
C3847 vdd.n2970 gnd 0.007324f
C3848 vdd.n2971 gnd 0.007324f
C3849 vdd.n2972 gnd 0.007324f
C3850 vdd.n2973 gnd 0.009099f
C3851 vdd.n2975 gnd 0.009099f
C3852 vdd.n2976 gnd 0.009099f
C3853 vdd.n2977 gnd 0.007324f
C3854 vdd.n2978 gnd 0.007324f
C3855 vdd.n2979 gnd 0.007324f
C3856 vdd.n2980 gnd 0.009099f
C3857 vdd.n2982 gnd 0.009099f
C3858 vdd.n2983 gnd 0.009099f
C3859 vdd.n2984 gnd 0.007324f
C3860 vdd.n2985 gnd 0.009099f
C3861 vdd.n2986 gnd 0.009099f
C3862 vdd.n2987 gnd 0.009099f
C3863 vdd.n2988 gnd 0.015673f
C3864 vdd.n2989 gnd 0.006115f
C3865 vdd.n2990 gnd 0.007324f
C3866 vdd.n2991 gnd 0.009099f
C3867 vdd.n2993 gnd 0.009099f
C3868 vdd.n2994 gnd 0.009099f
C3869 vdd.n2995 gnd 0.007324f
C3870 vdd.n2996 gnd 0.007324f
C3871 vdd.n2997 gnd 0.007324f
C3872 vdd.n2998 gnd 0.009099f
C3873 vdd.n3000 gnd 0.009099f
C3874 vdd.n3001 gnd 0.009099f
C3875 vdd.n3002 gnd 0.007324f
C3876 vdd.n3003 gnd 0.007324f
C3877 vdd.n3004 gnd 0.007324f
C3878 vdd.n3005 gnd 0.009099f
C3879 vdd.n3007 gnd 0.009099f
C3880 vdd.n3008 gnd 0.009099f
C3881 vdd.n3009 gnd 0.007324f
C3882 vdd.n3010 gnd 0.007324f
C3883 vdd.n3011 gnd 0.007324f
C3884 vdd.n3012 gnd 0.009099f
C3885 vdd.n3014 gnd 0.009099f
C3886 vdd.n3015 gnd 0.009099f
C3887 vdd.n3017 gnd 0.009099f
C3888 vdd.n3018 gnd 0.007324f
C3889 vdd.n3019 gnd 0.007324f
C3890 vdd.n3020 gnd 0.006079f
C3891 vdd.n3021 gnd 0.022684f
C3892 vdd.n3022 gnd 0.022175f
C3893 vdd.n3023 gnd 0.006079f
C3894 vdd.n3024 gnd 0.022175f
C3895 vdd.n3025 gnd 1.37157f
C3896 vdd.t88 gnd 0.46494f
C3897 vdd.n3026 gnd 0.488187f
C3898 vdd.n3027 gnd 0.929881f
C3899 vdd.n3028 gnd 0.009099f
C3900 vdd.n3029 gnd 0.007324f
C3901 vdd.n3030 gnd 0.007324f
C3902 vdd.n3031 gnd 0.007324f
C3903 vdd.n3032 gnd 0.009099f
C3904 vdd.n3033 gnd 0.832243f
C3905 vdd.t20 gnd 0.46494f
C3906 vdd.n3034 gnd 0.562578f
C3907 vdd.n3035 gnd 0.674164f
C3908 vdd.n3036 gnd 0.009099f
C3909 vdd.n3037 gnd 0.007324f
C3910 vdd.n3038 gnd 0.007324f
C3911 vdd.n3039 gnd 0.007324f
C3912 vdd.n3040 gnd 0.009099f
C3913 vdd.n3041 gnd 0.516084f
C3914 vdd.t42 gnd 0.46494f
C3915 vdd.n3042 gnd 0.771801f
C3916 vdd.t18 gnd 0.46494f
C3917 vdd.n3043 gnd 0.571877f
C3918 vdd.n3044 gnd 0.009099f
C3919 vdd.n3045 gnd 0.007324f
C3920 vdd.n3046 gnd 0.006993f
C3921 vdd.n3047 gnd 0.536697f
C3922 vdd.n3048 gnd 1.84287f
C3923 a_n5644_8799.n0 gnd 0.206002f
C3924 a_n5644_8799.n1 gnd 0.283995f
C3925 a_n5644_8799.n2 gnd 0.21547f
C3926 a_n5644_8799.n3 gnd 0.206002f
C3927 a_n5644_8799.n4 gnd 0.283995f
C3928 a_n5644_8799.n5 gnd 0.21547f
C3929 a_n5644_8799.n6 gnd 0.206002f
C3930 a_n5644_8799.n7 gnd 0.447551f
C3931 a_n5644_8799.n8 gnd 0.21547f
C3932 a_n5644_8799.n9 gnd 0.206002f
C3933 a_n5644_8799.n10 gnd 0.318471f
C3934 a_n5644_8799.n11 gnd 0.180994f
C3935 a_n5644_8799.n12 gnd 0.206002f
C3936 a_n5644_8799.n13 gnd 0.318471f
C3937 a_n5644_8799.n14 gnd 0.180994f
C3938 a_n5644_8799.n15 gnd 0.206002f
C3939 a_n5644_8799.n16 gnd 0.318471f
C3940 a_n5644_8799.n17 gnd 0.34455f
C3941 a_n5644_8799.n18 gnd 2.78901f
C3942 a_n5644_8799.n19 gnd 3.96341f
C3943 a_n5644_8799.n20 gnd 0.248007f
C3944 a_n5644_8799.n21 gnd 0.00463f
C3945 a_n5644_8799.n22 gnd 0.010014f
C3946 a_n5644_8799.n23 gnd 0.010014f
C3947 a_n5644_8799.n24 gnd 0.00463f
C3948 a_n5644_8799.n25 gnd 0.248007f
C3949 a_n5644_8799.n26 gnd 0.00463f
C3950 a_n5644_8799.n27 gnd 0.010014f
C3951 a_n5644_8799.n28 gnd 0.010014f
C3952 a_n5644_8799.n29 gnd 0.00463f
C3953 a_n5644_8799.n30 gnd 0.248007f
C3954 a_n5644_8799.n31 gnd 0.00463f
C3955 a_n5644_8799.n32 gnd 0.010014f
C3956 a_n5644_8799.n33 gnd 0.010014f
C3957 a_n5644_8799.n34 gnd 0.00463f
C3958 a_n5644_8799.n35 gnd 0.00463f
C3959 a_n5644_8799.n36 gnd 0.010014f
C3960 a_n5644_8799.n37 gnd 0.010014f
C3961 a_n5644_8799.n38 gnd 0.00463f
C3962 a_n5644_8799.n39 gnd 0.248007f
C3963 a_n5644_8799.n40 gnd 0.00463f
C3964 a_n5644_8799.n41 gnd 0.010014f
C3965 a_n5644_8799.n42 gnd 0.010014f
C3966 a_n5644_8799.n43 gnd 0.00463f
C3967 a_n5644_8799.n44 gnd 0.248007f
C3968 a_n5644_8799.n45 gnd 0.00463f
C3969 a_n5644_8799.n46 gnd 0.010014f
C3970 a_n5644_8799.n47 gnd 0.010014f
C3971 a_n5644_8799.n48 gnd 0.00463f
C3972 a_n5644_8799.n49 gnd 0.248007f
C3973 a_n5644_8799.t17 gnd 0.142885f
C3974 a_n5644_8799.t16 gnd 0.142885f
C3975 a_n5644_8799.t2 gnd 0.142885f
C3976 a_n5644_8799.n50 gnd 1.12696f
C3977 a_n5644_8799.t5 gnd 0.142885f
C3978 a_n5644_8799.t26 gnd 0.142885f
C3979 a_n5644_8799.n51 gnd 1.1251f
C3980 a_n5644_8799.t13 gnd 0.142885f
C3981 a_n5644_8799.t12 gnd 0.142885f
C3982 a_n5644_8799.n52 gnd 1.1251f
C3983 a_n5644_8799.t22 gnd 0.111133f
C3984 a_n5644_8799.t15 gnd 0.111133f
C3985 a_n5644_8799.n53 gnd 0.984906f
C3986 a_n5644_8799.t8 gnd 0.111133f
C3987 a_n5644_8799.t19 gnd 0.111133f
C3988 a_n5644_8799.n54 gnd 0.982011f
C3989 a_n5644_8799.n55 gnd 0.870796f
C3990 a_n5644_8799.t7 gnd 0.111133f
C3991 a_n5644_8799.t31 gnd 0.111133f
C3992 a_n5644_8799.n56 gnd 0.982011f
C3993 a_n5644_8799.t21 gnd 0.111133f
C3994 a_n5644_8799.t29 gnd 0.111133f
C3995 a_n5644_8799.n57 gnd 0.984906f
C3996 a_n5644_8799.t27 gnd 0.111133f
C3997 a_n5644_8799.t3 gnd 0.111133f
C3998 a_n5644_8799.n58 gnd 0.98201f
C3999 a_n5644_8799.n59 gnd 0.870798f
C4000 a_n5644_8799.t28 gnd 0.111133f
C4001 a_n5644_8799.t9 gnd 0.111133f
C4002 a_n5644_8799.n60 gnd 0.98201f
C4003 a_n5644_8799.t18 gnd 0.111133f
C4004 a_n5644_8799.t4 gnd 0.111133f
C4005 a_n5644_8799.n61 gnd 0.984906f
C4006 a_n5644_8799.t20 gnd 0.111133f
C4007 a_n5644_8799.t23 gnd 0.111133f
C4008 a_n5644_8799.n62 gnd 0.98201f
C4009 a_n5644_8799.n63 gnd 0.870798f
C4010 a_n5644_8799.n64 gnd 2.70771f
C4011 a_n5644_8799.t24 gnd 0.111133f
C4012 a_n5644_8799.t10 gnd 0.111133f
C4013 a_n5644_8799.n65 gnd 0.982011f
C4014 a_n5644_8799.n66 gnd 2.89323f
C4015 a_n5644_8799.t11 gnd 0.111133f
C4016 a_n5644_8799.t14 gnd 0.111133f
C4017 a_n5644_8799.n67 gnd 0.982011f
C4018 a_n5644_8799.n68 gnd 0.428754f
C4019 a_n5644_8799.n69 gnd 0.780109f
C4020 a_n5644_8799.t71 gnd 0.592469f
C4021 a_n5644_8799.n70 gnd 0.266281f
C4022 a_n5644_8799.t38 gnd 0.592469f
C4023 a_n5644_8799.t58 gnd 0.592469f
C4024 a_n5644_8799.t49 gnd 0.603683f
C4025 a_n5644_8799.n71 gnd 0.248372f
C4026 a_n5644_8799.n72 gnd 0.268648f
C4027 a_n5644_8799.t73 gnd 0.592469f
C4028 a_n5644_8799.n73 gnd 0.266281f
C4029 a_n5644_8799.n74 gnd 0.261909f
C4030 a_n5644_8799.t48 gnd 0.592469f
C4031 a_n5644_8799.n75 gnd 0.261909f
C4032 a_n5644_8799.t37 gnd 0.592469f
C4033 a_n5644_8799.n76 gnd 0.268648f
C4034 a_n5644_8799.t36 gnd 0.603672f
C4035 a_n5644_8799.t75 gnd 0.592469f
C4036 a_n5644_8799.n77 gnd 0.266281f
C4037 a_n5644_8799.t45 gnd 0.592469f
C4038 a_n5644_8799.t64 gnd 0.592469f
C4039 a_n5644_8799.t54 gnd 0.603683f
C4040 a_n5644_8799.n78 gnd 0.248372f
C4041 a_n5644_8799.n79 gnd 0.268648f
C4042 a_n5644_8799.t77 gnd 0.592469f
C4043 a_n5644_8799.n80 gnd 0.266281f
C4044 a_n5644_8799.n81 gnd 0.261909f
C4045 a_n5644_8799.t53 gnd 0.592469f
C4046 a_n5644_8799.n82 gnd 0.261909f
C4047 a_n5644_8799.t41 gnd 0.592469f
C4048 a_n5644_8799.n83 gnd 0.268648f
C4049 a_n5644_8799.t43 gnd 0.603672f
C4050 a_n5644_8799.n84 gnd 0.891053f
C4051 a_n5644_8799.t62 gnd 0.592469f
C4052 a_n5644_8799.n85 gnd 0.266281f
C4053 a_n5644_8799.t70 gnd 0.592469f
C4054 a_n5644_8799.t67 gnd 0.592469f
C4055 a_n5644_8799.t35 gnd 0.603683f
C4056 a_n5644_8799.n86 gnd 0.248372f
C4057 a_n5644_8799.n87 gnd 0.268648f
C4058 a_n5644_8799.t44 gnd 0.592469f
C4059 a_n5644_8799.n88 gnd 0.266281f
C4060 a_n5644_8799.n89 gnd 0.261909f
C4061 a_n5644_8799.t50 gnd 0.592469f
C4062 a_n5644_8799.n90 gnd 0.261909f
C4063 a_n5644_8799.t39 gnd 0.592469f
C4064 a_n5644_8799.n91 gnd 0.268648f
C4065 a_n5644_8799.t79 gnd 0.603672f
C4066 a_n5644_8799.n92 gnd 1.48132f
C4067 a_n5644_8799.t56 gnd 0.603672f
C4068 a_n5644_8799.t55 gnd 0.592469f
C4069 a_n5644_8799.t42 gnd 0.592469f
C4070 a_n5644_8799.n93 gnd 0.266281f
C4071 a_n5644_8799.t72 gnd 0.592469f
C4072 a_n5644_8799.t57 gnd 0.592469f
C4073 a_n5644_8799.t47 gnd 0.592469f
C4074 a_n5644_8799.n94 gnd 0.266281f
C4075 a_n5644_8799.t65 gnd 0.603683f
C4076 a_n5644_8799.n95 gnd 0.248372f
C4077 a_n5644_8799.t74 gnd 0.592469f
C4078 a_n5644_8799.n96 gnd 0.268648f
C4079 a_n5644_8799.n97 gnd 0.261909f
C4080 a_n5644_8799.n98 gnd 0.261909f
C4081 a_n5644_8799.n99 gnd 0.268648f
C4082 a_n5644_8799.t60 gnd 0.603672f
C4083 a_n5644_8799.t59 gnd 0.592469f
C4084 a_n5644_8799.t51 gnd 0.592469f
C4085 a_n5644_8799.n100 gnd 0.266281f
C4086 a_n5644_8799.t76 gnd 0.592469f
C4087 a_n5644_8799.t63 gnd 0.592469f
C4088 a_n5644_8799.t52 gnd 0.592469f
C4089 a_n5644_8799.n101 gnd 0.266281f
C4090 a_n5644_8799.t68 gnd 0.603683f
C4091 a_n5644_8799.n102 gnd 0.248372f
C4092 a_n5644_8799.t32 gnd 0.592469f
C4093 a_n5644_8799.n103 gnd 0.268648f
C4094 a_n5644_8799.n104 gnd 0.261909f
C4095 a_n5644_8799.n105 gnd 0.261909f
C4096 a_n5644_8799.n106 gnd 0.268648f
C4097 a_n5644_8799.n107 gnd 0.891053f
C4098 a_n5644_8799.t78 gnd 0.603672f
C4099 a_n5644_8799.t40 gnd 0.592469f
C4100 a_n5644_8799.t61 gnd 0.592469f
C4101 a_n5644_8799.n108 gnd 0.266281f
C4102 a_n5644_8799.t33 gnd 0.592469f
C4103 a_n5644_8799.t69 gnd 0.592469f
C4104 a_n5644_8799.t46 gnd 0.592469f
C4105 a_n5644_8799.n109 gnd 0.266281f
C4106 a_n5644_8799.t34 gnd 0.603683f
C4107 a_n5644_8799.n110 gnd 0.248372f
C4108 a_n5644_8799.t66 gnd 0.592469f
C4109 a_n5644_8799.n111 gnd 0.268648f
C4110 a_n5644_8799.n112 gnd 0.261909f
C4111 a_n5644_8799.n113 gnd 0.261909f
C4112 a_n5644_8799.n114 gnd 0.268648f
C4113 a_n5644_8799.n115 gnd 1.10132f
C4114 a_n5644_8799.n116 gnd 12.120501f
C4115 a_n5644_8799.n117 gnd 4.33602f
C4116 a_n5644_8799.n118 gnd 5.634759f
C4117 a_n5644_8799.t1 gnd 0.142885f
C4118 a_n5644_8799.t25 gnd 0.142885f
C4119 a_n5644_8799.n119 gnd 1.12696f
C4120 a_n5644_8799.t30 gnd 0.142885f
C4121 a_n5644_8799.t6 gnd 0.142885f
C4122 a_n5644_8799.n120 gnd 1.1251f
C4123 a_n5644_8799.n121 gnd 1.1251f
C4124 a_n5644_8799.t0 gnd 0.142885f
C4125 a_n1986_8322.n0 gnd 1.85102f
C4126 a_n1986_8322.n1 gnd 1.11016f
C4127 a_n1986_8322.n2 gnd 1.11016f
C4128 a_n1986_8322.n3 gnd 0.872286f
C4129 a_n1986_8322.t8 gnd 0.124841p
C4130 a_n1986_8322.t18 gnd 0.875759f
C4131 a_n1986_8322.t7 gnd 0.093529f
C4132 a_n1986_8322.t2 gnd 0.093529f
C4133 a_n1986_8322.n4 gnd 0.65882f
C4134 a_n1986_8322.t1 gnd 0.093529f
C4135 a_n1986_8322.t20 gnd 0.093529f
C4136 a_n1986_8322.n5 gnd 0.65882f
C4137 a_n1986_8322.t14 gnd 0.874017f
C4138 a_n1986_8322.n6 gnd 0.766493f
C4139 a_n1986_8322.n7 gnd 3.48702f
C4140 a_n1986_8322.t10 gnd 0.875761f
C4141 a_n1986_8322.t19 gnd 0.093529f
C4142 a_n1986_8322.t11 gnd 0.093529f
C4143 a_n1986_8322.n8 gnd 0.65882f
C4144 a_n1986_8322.t5 gnd 0.093529f
C4145 a_n1986_8322.t6 gnd 0.093529f
C4146 a_n1986_8322.n9 gnd 0.65882f
C4147 a_n1986_8322.t13 gnd 0.874017f
C4148 a_n1986_8322.n10 gnd 1.39891f
C4149 a_n1986_8322.n11 gnd 1.59065f
C4150 a_n1986_8322.t4 gnd 0.874017f
C4151 a_n1986_8322.t3 gnd 0.093529f
C4152 a_n1986_8322.t9 gnd 0.093529f
C4153 a_n1986_8322.n12 gnd 0.65882f
C4154 a_n1986_8322.t17 gnd 0.874017f
C4155 a_n1986_8322.t12 gnd 0.874017f
C4156 a_n1986_8322.t15 gnd 0.093529f
C4157 a_n1986_8322.t16 gnd 0.093529f
C4158 a_n1986_8322.n13 gnd 0.65882f
C4159 a_n1986_8322.t0 gnd 0.875761f
C4160 CSoutput.n0 gnd 0.037845f
C4161 CSoutput.t148 gnd 0.250336f
C4162 CSoutput.n1 gnd 0.113039f
C4163 CSoutput.n2 gnd 0.037845f
C4164 CSoutput.t156 gnd 0.250336f
C4165 CSoutput.n3 gnd 0.029995f
C4166 CSoutput.n4 gnd 0.037845f
C4167 CSoutput.t163 gnd 0.250336f
C4168 CSoutput.n5 gnd 0.025865f
C4169 CSoutput.n6 gnd 0.037845f
C4170 CSoutput.t152 gnd 0.250336f
C4171 CSoutput.t150 gnd 0.250336f
C4172 CSoutput.n7 gnd 0.111807f
C4173 CSoutput.n8 gnd 0.037845f
C4174 CSoutput.t162 gnd 0.250336f
C4175 CSoutput.n9 gnd 0.024661f
C4176 CSoutput.n10 gnd 0.037845f
C4177 CSoutput.t165 gnd 0.250336f
C4178 CSoutput.t147 gnd 0.250336f
C4179 CSoutput.n11 gnd 0.111807f
C4180 CSoutput.n12 gnd 0.037845f
C4181 CSoutput.t159 gnd 0.250336f
C4182 CSoutput.n13 gnd 0.025865f
C4183 CSoutput.n14 gnd 0.037845f
C4184 CSoutput.t158 gnd 0.250336f
C4185 CSoutput.t145 gnd 0.250336f
C4186 CSoutput.n15 gnd 0.111807f
C4187 CSoutput.n16 gnd 0.037845f
C4188 CSoutput.t151 gnd 0.250336f
C4189 CSoutput.n17 gnd 0.027625f
C4190 CSoutput.t160 gnd 0.299159f
C4191 CSoutput.t157 gnd 0.250336f
C4192 CSoutput.n18 gnd 0.142735f
C4193 CSoutput.n19 gnd 0.138502f
C4194 CSoutput.n20 gnd 0.160679f
C4195 CSoutput.n21 gnd 0.037845f
C4196 CSoutput.n22 gnd 0.031586f
C4197 CSoutput.n23 gnd 0.111807f
C4198 CSoutput.n24 gnd 0.030448f
C4199 CSoutput.n25 gnd 0.029995f
C4200 CSoutput.n26 gnd 0.037845f
C4201 CSoutput.n27 gnd 0.037845f
C4202 CSoutput.n28 gnd 0.031343f
C4203 CSoutput.n29 gnd 0.026611f
C4204 CSoutput.n30 gnd 0.114296f
C4205 CSoutput.n31 gnd 0.026978f
C4206 CSoutput.n32 gnd 0.037845f
C4207 CSoutput.n33 gnd 0.037845f
C4208 CSoutput.n34 gnd 0.037845f
C4209 CSoutput.n35 gnd 0.031009f
C4210 CSoutput.n36 gnd 0.111807f
C4211 CSoutput.n37 gnd 0.029656f
C4212 CSoutput.n38 gnd 0.030787f
C4213 CSoutput.n39 gnd 0.037845f
C4214 CSoutput.n40 gnd 0.037845f
C4215 CSoutput.n41 gnd 0.031579f
C4216 CSoutput.n42 gnd 0.028864f
C4217 CSoutput.n43 gnd 0.111807f
C4218 CSoutput.n44 gnd 0.029595f
C4219 CSoutput.n45 gnd 0.037845f
C4220 CSoutput.n46 gnd 0.037845f
C4221 CSoutput.n47 gnd 0.037845f
C4222 CSoutput.n48 gnd 0.029595f
C4223 CSoutput.n49 gnd 0.111807f
C4224 CSoutput.n50 gnd 0.028864f
C4225 CSoutput.n51 gnd 0.031579f
C4226 CSoutput.n52 gnd 0.037845f
C4227 CSoutput.n53 gnd 0.037845f
C4228 CSoutput.n54 gnd 0.030787f
C4229 CSoutput.n55 gnd 0.029656f
C4230 CSoutput.n56 gnd 0.111807f
C4231 CSoutput.n57 gnd 0.031009f
C4232 CSoutput.n58 gnd 0.037845f
C4233 CSoutput.n59 gnd 0.037845f
C4234 CSoutput.n60 gnd 0.037845f
C4235 CSoutput.n61 gnd 0.026978f
C4236 CSoutput.n62 gnd 0.114296f
C4237 CSoutput.n63 gnd 0.026611f
C4238 CSoutput.t154 gnd 0.250336f
C4239 CSoutput.n64 gnd 0.111807f
C4240 CSoutput.n65 gnd 0.031343f
C4241 CSoutput.n66 gnd 0.037845f
C4242 CSoutput.n67 gnd 0.037845f
C4243 CSoutput.n68 gnd 0.037845f
C4244 CSoutput.n69 gnd 0.030448f
C4245 CSoutput.n70 gnd 0.111807f
C4246 CSoutput.n71 gnd 0.031586f
C4247 CSoutput.n72 gnd 0.027625f
C4248 CSoutput.n73 gnd 0.037845f
C4249 CSoutput.n74 gnd 0.037845f
C4250 CSoutput.n75 gnd 0.028649f
C4251 CSoutput.n76 gnd 0.017015f
C4252 CSoutput.t161 gnd 0.281271f
C4253 CSoutput.n77 gnd 0.139724f
C4254 CSoutput.n78 gnd 0.571604f
C4255 CSoutput.t7 gnd 0.047206f
C4256 CSoutput.t16 gnd 0.047206f
C4257 CSoutput.n79 gnd 0.365487f
C4258 CSoutput.t136 gnd 0.047206f
C4259 CSoutput.t38 gnd 0.047206f
C4260 CSoutput.n80 gnd 0.364835f
C4261 CSoutput.n81 gnd 0.370307f
C4262 CSoutput.t29 gnd 0.047206f
C4263 CSoutput.t8 gnd 0.047206f
C4264 CSoutput.n82 gnd 0.364835f
C4265 CSoutput.n83 gnd 0.182472f
C4266 CSoutput.t20 gnd 0.047206f
C4267 CSoutput.t15 gnd 0.047206f
C4268 CSoutput.n84 gnd 0.364835f
C4269 CSoutput.n85 gnd 0.334611f
C4270 CSoutput.t142 gnd 0.047206f
C4271 CSoutput.t27 gnd 0.047206f
C4272 CSoutput.n86 gnd 0.365487f
C4273 CSoutput.t28 gnd 0.047206f
C4274 CSoutput.t18 gnd 0.047206f
C4275 CSoutput.n87 gnd 0.364835f
C4276 CSoutput.n88 gnd 0.370307f
C4277 CSoutput.t13 gnd 0.047206f
C4278 CSoutput.t34 gnd 0.047206f
C4279 CSoutput.n89 gnd 0.364835f
C4280 CSoutput.n90 gnd 0.182472f
C4281 CSoutput.t1 gnd 0.047206f
C4282 CSoutput.t35 gnd 0.047206f
C4283 CSoutput.n91 gnd 0.364835f
C4284 CSoutput.n92 gnd 0.272111f
C4285 CSoutput.n93 gnd 0.343131f
C4286 CSoutput.t9 gnd 0.047206f
C4287 CSoutput.t11 gnd 0.047206f
C4288 CSoutput.n94 gnd 0.365487f
C4289 CSoutput.t143 gnd 0.047206f
C4290 CSoutput.t21 gnd 0.047206f
C4291 CSoutput.n95 gnd 0.364835f
C4292 CSoutput.n96 gnd 0.370307f
C4293 CSoutput.t138 gnd 0.047206f
C4294 CSoutput.t19 gnd 0.047206f
C4295 CSoutput.n97 gnd 0.364835f
C4296 CSoutput.n98 gnd 0.182472f
C4297 CSoutput.t3 gnd 0.047206f
C4298 CSoutput.t137 gnd 0.047206f
C4299 CSoutput.n99 gnd 0.364835f
C4300 CSoutput.n100 gnd 0.272111f
C4301 CSoutput.n101 gnd 0.383532f
C4302 CSoutput.n102 gnd 6.9206f
C4303 CSoutput.n104 gnd 0.669471f
C4304 CSoutput.n105 gnd 0.502103f
C4305 CSoutput.n106 gnd 0.669471f
C4306 CSoutput.n107 gnd 0.669471f
C4307 CSoutput.n108 gnd 1.80242f
C4308 CSoutput.n109 gnd 0.669471f
C4309 CSoutput.n110 gnd 0.669471f
C4310 CSoutput.t153 gnd 0.836839f
C4311 CSoutput.n111 gnd 0.669471f
C4312 CSoutput.n112 gnd 0.669471f
C4313 CSoutput.n116 gnd 0.669471f
C4314 CSoutput.n120 gnd 0.669471f
C4315 CSoutput.n121 gnd 0.669471f
C4316 CSoutput.n123 gnd 0.669471f
C4317 CSoutput.n128 gnd 0.669471f
C4318 CSoutput.n130 gnd 0.669471f
C4319 CSoutput.n131 gnd 0.669471f
C4320 CSoutput.n133 gnd 0.669471f
C4321 CSoutput.n134 gnd 0.669471f
C4322 CSoutput.n136 gnd 0.669471f
C4323 CSoutput.t146 gnd 11.1868f
C4324 CSoutput.n138 gnd 0.669471f
C4325 CSoutput.n139 gnd 0.502103f
C4326 CSoutput.n140 gnd 0.669471f
C4327 CSoutput.n141 gnd 0.669471f
C4328 CSoutput.n142 gnd 1.80242f
C4329 CSoutput.n143 gnd 0.669471f
C4330 CSoutput.n144 gnd 0.669471f
C4331 CSoutput.t164 gnd 0.836839f
C4332 CSoutput.n145 gnd 0.669471f
C4333 CSoutput.n146 gnd 0.669471f
C4334 CSoutput.n150 gnd 0.669471f
C4335 CSoutput.n154 gnd 0.669471f
C4336 CSoutput.n155 gnd 0.669471f
C4337 CSoutput.n157 gnd 0.669471f
C4338 CSoutput.n162 gnd 0.669471f
C4339 CSoutput.n164 gnd 0.669471f
C4340 CSoutput.n165 gnd 0.669471f
C4341 CSoutput.n167 gnd 0.669471f
C4342 CSoutput.n168 gnd 0.669471f
C4343 CSoutput.n170 gnd 0.669471f
C4344 CSoutput.n171 gnd 0.502103f
C4345 CSoutput.n173 gnd 0.669471f
C4346 CSoutput.n174 gnd 0.502103f
C4347 CSoutput.n175 gnd 0.669471f
C4348 CSoutput.n176 gnd 0.669471f
C4349 CSoutput.n177 gnd 1.80242f
C4350 CSoutput.n178 gnd 0.669471f
C4351 CSoutput.n179 gnd 0.669471f
C4352 CSoutput.t144 gnd 0.836839f
C4353 CSoutput.n180 gnd 0.669471f
C4354 CSoutput.n181 gnd 1.80242f
C4355 CSoutput.n183 gnd 0.669471f
C4356 CSoutput.n184 gnd 0.669471f
C4357 CSoutput.n186 gnd 0.669471f
C4358 CSoutput.n187 gnd 0.669471f
C4359 CSoutput.t155 gnd 11.004499f
C4360 CSoutput.t149 gnd 11.1868f
C4361 CSoutput.n193 gnd 2.10023f
C4362 CSoutput.n194 gnd 8.555571f
C4363 CSoutput.n195 gnd 8.91357f
C4364 CSoutput.n200 gnd 2.27511f
C4365 CSoutput.n206 gnd 0.669471f
C4366 CSoutput.n208 gnd 0.669471f
C4367 CSoutput.n210 gnd 0.669471f
C4368 CSoutput.n212 gnd 0.669471f
C4369 CSoutput.n214 gnd 0.669471f
C4370 CSoutput.n220 gnd 0.669471f
C4371 CSoutput.n227 gnd 1.22822f
C4372 CSoutput.n228 gnd 1.22822f
C4373 CSoutput.n229 gnd 0.669471f
C4374 CSoutput.n230 gnd 0.669471f
C4375 CSoutput.n232 gnd 0.502103f
C4376 CSoutput.n233 gnd 0.430006f
C4377 CSoutput.n235 gnd 0.502103f
C4378 CSoutput.n236 gnd 0.430006f
C4379 CSoutput.n237 gnd 0.502103f
C4380 CSoutput.n239 gnd 0.669471f
C4381 CSoutput.n241 gnd 1.80242f
C4382 CSoutput.n242 gnd 2.10023f
C4383 CSoutput.n243 gnd 7.86892f
C4384 CSoutput.n245 gnd 0.502103f
C4385 CSoutput.n246 gnd 1.29194f
C4386 CSoutput.n247 gnd 0.502103f
C4387 CSoutput.n249 gnd 0.669471f
C4388 CSoutput.n251 gnd 1.80242f
C4389 CSoutput.n252 gnd 3.92597f
C4390 CSoutput.t10 gnd 0.047206f
C4391 CSoutput.t31 gnd 0.047206f
C4392 CSoutput.n253 gnd 0.365487f
C4393 CSoutput.t23 gnd 0.047206f
C4394 CSoutput.t30 gnd 0.047206f
C4395 CSoutput.n254 gnd 0.364835f
C4396 CSoutput.n255 gnd 0.370307f
C4397 CSoutput.t5 gnd 0.047206f
C4398 CSoutput.t26 gnd 0.047206f
C4399 CSoutput.n256 gnd 0.364835f
C4400 CSoutput.n257 gnd 0.182472f
C4401 CSoutput.t39 gnd 0.047206f
C4402 CSoutput.t22 gnd 0.047206f
C4403 CSoutput.n258 gnd 0.364835f
C4404 CSoutput.n259 gnd 0.334611f
C4405 CSoutput.t32 gnd 0.047206f
C4406 CSoutput.t36 gnd 0.047206f
C4407 CSoutput.n260 gnd 0.365487f
C4408 CSoutput.t6 gnd 0.047206f
C4409 CSoutput.t4 gnd 0.047206f
C4410 CSoutput.n261 gnd 0.364835f
C4411 CSoutput.n262 gnd 0.370307f
C4412 CSoutput.t25 gnd 0.047206f
C4413 CSoutput.t14 gnd 0.047206f
C4414 CSoutput.n263 gnd 0.364835f
C4415 CSoutput.n264 gnd 0.182472f
C4416 CSoutput.t139 gnd 0.047206f
C4417 CSoutput.t17 gnd 0.047206f
C4418 CSoutput.n265 gnd 0.364835f
C4419 CSoutput.n266 gnd 0.272111f
C4420 CSoutput.n267 gnd 0.343131f
C4421 CSoutput.t24 gnd 0.047206f
C4422 CSoutput.t141 gnd 0.047206f
C4423 CSoutput.n268 gnd 0.365487f
C4424 CSoutput.t12 gnd 0.047206f
C4425 CSoutput.t2 gnd 0.047206f
C4426 CSoutput.n269 gnd 0.364835f
C4427 CSoutput.n270 gnd 0.370307f
C4428 CSoutput.t37 gnd 0.047206f
C4429 CSoutput.t140 gnd 0.047206f
C4430 CSoutput.n271 gnd 0.364835f
C4431 CSoutput.n272 gnd 0.182472f
C4432 CSoutput.t33 gnd 0.047206f
C4433 CSoutput.t0 gnd 0.047206f
C4434 CSoutput.n273 gnd 0.364834f
C4435 CSoutput.n274 gnd 0.272113f
C4436 CSoutput.n275 gnd 0.383532f
C4437 CSoutput.n276 gnd 9.9266f
C4438 CSoutput.t79 gnd 0.041305f
C4439 CSoutput.t134 gnd 0.041305f
C4440 CSoutput.n277 gnd 0.366211f
C4441 CSoutput.t73 gnd 0.041305f
C4442 CSoutput.t78 gnd 0.041305f
C4443 CSoutput.n278 gnd 0.36499f
C4444 CSoutput.n279 gnd 0.340103f
C4445 CSoutput.t64 gnd 0.041305f
C4446 CSoutput.t82 gnd 0.041305f
C4447 CSoutput.n280 gnd 0.36499f
C4448 CSoutput.n281 gnd 0.167654f
C4449 CSoutput.t97 gnd 0.041305f
C4450 CSoutput.t74 gnd 0.041305f
C4451 CSoutput.n282 gnd 0.36499f
C4452 CSoutput.n283 gnd 0.167654f
C4453 CSoutput.t80 gnd 0.041305f
C4454 CSoutput.t120 gnd 0.041305f
C4455 CSoutput.n284 gnd 0.36499f
C4456 CSoutput.n285 gnd 0.167654f
C4457 CSoutput.t93 gnd 0.041305f
C4458 CSoutput.t103 gnd 0.041305f
C4459 CSoutput.n286 gnd 0.36499f
C4460 CSoutput.n287 gnd 0.167654f
C4461 CSoutput.t58 gnd 0.041305f
C4462 CSoutput.t83 gnd 0.041305f
C4463 CSoutput.n288 gnd 0.36499f
C4464 CSoutput.n289 gnd 0.167654f
C4465 CSoutput.t47 gnd 0.041305f
C4466 CSoutput.t70 gnd 0.041305f
C4467 CSoutput.n290 gnd 0.36499f
C4468 CSoutput.n291 gnd 0.30923f
C4469 CSoutput.t131 gnd 0.041305f
C4470 CSoutput.t40 gnd 0.041305f
C4471 CSoutput.n292 gnd 0.366211f
C4472 CSoutput.t51 gnd 0.041305f
C4473 CSoutput.t121 gnd 0.041305f
C4474 CSoutput.n293 gnd 0.36499f
C4475 CSoutput.n294 gnd 0.340103f
C4476 CSoutput.t41 gnd 0.041305f
C4477 CSoutput.t114 gnd 0.041305f
C4478 CSoutput.n295 gnd 0.36499f
C4479 CSoutput.n296 gnd 0.167654f
C4480 CSoutput.t122 gnd 0.041305f
C4481 CSoutput.t42 gnd 0.041305f
C4482 CSoutput.n297 gnd 0.36499f
C4483 CSoutput.n298 gnd 0.167654f
C4484 CSoutput.t105 gnd 0.041305f
C4485 CSoutput.t86 gnd 0.041305f
C4486 CSoutput.n299 gnd 0.36499f
C4487 CSoutput.n300 gnd 0.167654f
C4488 CSoutput.t43 gnd 0.041305f
C4489 CSoutput.t107 gnd 0.041305f
C4490 CSoutput.n301 gnd 0.36499f
C4491 CSoutput.n302 gnd 0.167654f
C4492 CSoutput.t90 gnd 0.041305f
C4493 CSoutput.t94 gnd 0.041305f
C4494 CSoutput.n303 gnd 0.36499f
C4495 CSoutput.n304 gnd 0.167654f
C4496 CSoutput.t108 gnd 0.041305f
C4497 CSoutput.t91 gnd 0.041305f
C4498 CSoutput.n305 gnd 0.36499f
C4499 CSoutput.n306 gnd 0.254535f
C4500 CSoutput.n307 gnd 0.321048f
C4501 CSoutput.t52 gnd 0.041305f
C4502 CSoutput.t124 gnd 0.041305f
C4503 CSoutput.n308 gnd 0.366211f
C4504 CSoutput.t71 gnd 0.041305f
C4505 CSoutput.t75 gnd 0.041305f
C4506 CSoutput.n309 gnd 0.36499f
C4507 CSoutput.n310 gnd 0.340103f
C4508 CSoutput.t44 gnd 0.041305f
C4509 CSoutput.t110 gnd 0.041305f
C4510 CSoutput.n311 gnd 0.36499f
C4511 CSoutput.n312 gnd 0.167654f
C4512 CSoutput.t81 gnd 0.041305f
C4513 CSoutput.t53 gnd 0.041305f
C4514 CSoutput.n313 gnd 0.36499f
C4515 CSoutput.n314 gnd 0.167654f
C4516 CSoutput.t61 gnd 0.041305f
C4517 CSoutput.t135 gnd 0.041305f
C4518 CSoutput.n315 gnd 0.36499f
C4519 CSoutput.n316 gnd 0.167654f
C4520 CSoutput.t62 gnd 0.041305f
C4521 CSoutput.t66 gnd 0.041305f
C4522 CSoutput.n317 gnd 0.36499f
C4523 CSoutput.n318 gnd 0.167654f
C4524 CSoutput.t50 gnd 0.041305f
C4525 CSoutput.t123 gnd 0.041305f
C4526 CSoutput.n319 gnd 0.36499f
C4527 CSoutput.n320 gnd 0.167654f
C4528 CSoutput.t69 gnd 0.041305f
C4529 CSoutput.t60 gnd 0.041305f
C4530 CSoutput.n321 gnd 0.36499f
C4531 CSoutput.n322 gnd 0.254535f
C4532 CSoutput.n323 gnd 0.344755f
C4533 CSoutput.n324 gnd 10.6183f
C4534 CSoutput.t65 gnd 0.041305f
C4535 CSoutput.t106 gnd 0.041305f
C4536 CSoutput.n325 gnd 0.366211f
C4537 CSoutput.t104 gnd 0.041305f
C4538 CSoutput.t85 gnd 0.041305f
C4539 CSoutput.n326 gnd 0.36499f
C4540 CSoutput.n327 gnd 0.340103f
C4541 CSoutput.t111 gnd 0.041305f
C4542 CSoutput.t76 gnd 0.041305f
C4543 CSoutput.n328 gnd 0.36499f
C4544 CSoutput.n329 gnd 0.167654f
C4545 CSoutput.t95 gnd 0.041305f
C4546 CSoutput.t125 gnd 0.041305f
C4547 CSoutput.n330 gnd 0.36499f
C4548 CSoutput.n331 gnd 0.167654f
C4549 CSoutput.t59 gnd 0.041305f
C4550 CSoutput.t109 gnd 0.041305f
C4551 CSoutput.n332 gnd 0.36499f
C4552 CSoutput.n333 gnd 0.167654f
C4553 CSoutput.t48 gnd 0.041305f
C4554 CSoutput.t116 gnd 0.041305f
C4555 CSoutput.n334 gnd 0.36499f
C4556 CSoutput.n335 gnd 0.167654f
C4557 CSoutput.t115 gnd 0.041305f
C4558 CSoutput.t72 gnd 0.041305f
C4559 CSoutput.n336 gnd 0.36499f
C4560 CSoutput.n337 gnd 0.167654f
C4561 CSoutput.t87 gnd 0.041305f
C4562 CSoutput.t68 gnd 0.041305f
C4563 CSoutput.n338 gnd 0.36499f
C4564 CSoutput.n339 gnd 0.30923f
C4565 CSoutput.t57 gnd 0.041305f
C4566 CSoutput.t49 gnd 0.041305f
C4567 CSoutput.n340 gnd 0.366211f
C4568 CSoutput.t45 gnd 0.041305f
C4569 CSoutput.t133 gnd 0.041305f
C4570 CSoutput.n341 gnd 0.36499f
C4571 CSoutput.n342 gnd 0.340103f
C4572 CSoutput.t132 gnd 0.041305f
C4573 CSoutput.t56 gnd 0.041305f
C4574 CSoutput.n343 gnd 0.36499f
C4575 CSoutput.n344 gnd 0.167654f
C4576 CSoutput.t55 gnd 0.041305f
C4577 CSoutput.t101 gnd 0.041305f
C4578 CSoutput.n345 gnd 0.36499f
C4579 CSoutput.n346 gnd 0.167654f
C4580 CSoutput.t98 gnd 0.041305f
C4581 CSoutput.t129 gnd 0.041305f
C4582 CSoutput.n347 gnd 0.36499f
C4583 CSoutput.n348 gnd 0.167654f
C4584 CSoutput.t127 gnd 0.041305f
C4585 CSoutput.t119 gnd 0.041305f
C4586 CSoutput.n349 gnd 0.36499f
C4587 CSoutput.n350 gnd 0.167654f
C4588 CSoutput.t112 gnd 0.041305f
C4589 CSoutput.t99 gnd 0.041305f
C4590 CSoutput.n351 gnd 0.36499f
C4591 CSoutput.n352 gnd 0.167654f
C4592 CSoutput.t100 gnd 0.041305f
C4593 CSoutput.t128 gnd 0.041305f
C4594 CSoutput.n353 gnd 0.36499f
C4595 CSoutput.n354 gnd 0.254535f
C4596 CSoutput.n355 gnd 0.321048f
C4597 CSoutput.t92 gnd 0.041305f
C4598 CSoutput.t117 gnd 0.041305f
C4599 CSoutput.n356 gnd 0.366211f
C4600 CSoutput.t63 gnd 0.041305f
C4601 CSoutput.t77 gnd 0.041305f
C4602 CSoutput.n357 gnd 0.36499f
C4603 CSoutput.n358 gnd 0.340103f
C4604 CSoutput.t84 gnd 0.041305f
C4605 CSoutput.t102 gnd 0.041305f
C4606 CSoutput.n359 gnd 0.36499f
C4607 CSoutput.n360 gnd 0.167654f
C4608 CSoutput.t118 gnd 0.041305f
C4609 CSoutput.t89 gnd 0.041305f
C4610 CSoutput.n361 gnd 0.36499f
C4611 CSoutput.n362 gnd 0.167654f
C4612 CSoutput.t96 gnd 0.041305f
C4613 CSoutput.t130 gnd 0.041305f
C4614 CSoutput.n363 gnd 0.36499f
C4615 CSoutput.n364 gnd 0.167654f
C4616 CSoutput.t46 gnd 0.041305f
C4617 CSoutput.t67 gnd 0.041305f
C4618 CSoutput.n365 gnd 0.36499f
C4619 CSoutput.n366 gnd 0.167654f
C4620 CSoutput.t88 gnd 0.041305f
C4621 CSoutput.t113 gnd 0.041305f
C4622 CSoutput.n367 gnd 0.36499f
C4623 CSoutput.n368 gnd 0.167654f
C4624 CSoutput.t126 gnd 0.041305f
C4625 CSoutput.t54 gnd 0.041305f
C4626 CSoutput.n369 gnd 0.36499f
C4627 CSoutput.n370 gnd 0.254535f
C4628 CSoutput.n371 gnd 0.344755f
C4629 CSoutput.n372 gnd 6.01389f
C4630 CSoutput.n373 gnd 11.6587f
C4631 commonsourceibias.n0 gnd 0.012624f
C4632 commonsourceibias.t120 gnd 0.191163f
C4633 commonsourceibias.t65 gnd 0.176757f
C4634 commonsourceibias.n1 gnd 0.00769f
C4635 commonsourceibias.n2 gnd 0.009461f
C4636 commonsourceibias.t126 gnd 0.176757f
C4637 commonsourceibias.n3 gnd 0.009597f
C4638 commonsourceibias.n4 gnd 0.009461f
C4639 commonsourceibias.t121 gnd 0.176757f
C4640 commonsourceibias.n5 gnd 0.070526f
C4641 commonsourceibias.t135 gnd 0.176757f
C4642 commonsourceibias.n6 gnd 0.007653f
C4643 commonsourceibias.n7 gnd 0.009461f
C4644 commonsourceibias.t117 gnd 0.176757f
C4645 commonsourceibias.n8 gnd 0.009134f
C4646 commonsourceibias.n9 gnd 0.009461f
C4647 commonsourceibias.t102 gnd 0.176757f
C4648 commonsourceibias.n10 gnd 0.070526f
C4649 commonsourceibias.t125 gnd 0.176757f
C4650 commonsourceibias.n11 gnd 0.007641f
C4651 commonsourceibias.n12 gnd 0.012624f
C4652 commonsourceibias.t54 gnd 0.191163f
C4653 commonsourceibias.t20 gnd 0.176757f
C4654 commonsourceibias.n13 gnd 0.00769f
C4655 commonsourceibias.n14 gnd 0.009461f
C4656 commonsourceibias.t4 gnd 0.176757f
C4657 commonsourceibias.n15 gnd 0.009597f
C4658 commonsourceibias.n16 gnd 0.009461f
C4659 commonsourceibias.t52 gnd 0.176757f
C4660 commonsourceibias.n17 gnd 0.070526f
C4661 commonsourceibias.t14 gnd 0.176757f
C4662 commonsourceibias.n18 gnd 0.007653f
C4663 commonsourceibias.n19 gnd 0.009461f
C4664 commonsourceibias.t58 gnd 0.176757f
C4665 commonsourceibias.n20 gnd 0.009134f
C4666 commonsourceibias.n21 gnd 0.009461f
C4667 commonsourceibias.t32 gnd 0.176757f
C4668 commonsourceibias.n22 gnd 0.070526f
C4669 commonsourceibias.t6 gnd 0.176757f
C4670 commonsourceibias.n23 gnd 0.007641f
C4671 commonsourceibias.n24 gnd 0.009461f
C4672 commonsourceibias.t56 gnd 0.176757f
C4673 commonsourceibias.t28 gnd 0.176757f
C4674 commonsourceibias.n25 gnd 0.070526f
C4675 commonsourceibias.n26 gnd 0.009461f
C4676 commonsourceibias.t48 gnd 0.176757f
C4677 commonsourceibias.n27 gnd 0.070526f
C4678 commonsourceibias.n28 gnd 0.009461f
C4679 commonsourceibias.t34 gnd 0.176757f
C4680 commonsourceibias.n29 gnd 0.070526f
C4681 commonsourceibias.n30 gnd 0.009461f
C4682 commonsourceibias.t18 gnd 0.176757f
C4683 commonsourceibias.n31 gnd 0.010754f
C4684 commonsourceibias.n32 gnd 0.009461f
C4685 commonsourceibias.t60 gnd 0.176757f
C4686 commonsourceibias.n33 gnd 0.012717f
C4687 commonsourceibias.t62 gnd 0.196904f
C4688 commonsourceibias.t22 gnd 0.176757f
C4689 commonsourceibias.n34 gnd 0.078584f
C4690 commonsourceibias.n35 gnd 0.084191f
C4691 commonsourceibias.n36 gnd 0.04027f
C4692 commonsourceibias.n37 gnd 0.009461f
C4693 commonsourceibias.n38 gnd 0.00769f
C4694 commonsourceibias.n39 gnd 0.013037f
C4695 commonsourceibias.n40 gnd 0.070526f
C4696 commonsourceibias.n41 gnd 0.013093f
C4697 commonsourceibias.n42 gnd 0.009461f
C4698 commonsourceibias.n43 gnd 0.009461f
C4699 commonsourceibias.n44 gnd 0.009461f
C4700 commonsourceibias.n45 gnd 0.009597f
C4701 commonsourceibias.n46 gnd 0.070526f
C4702 commonsourceibias.n47 gnd 0.011661f
C4703 commonsourceibias.n48 gnd 0.0129f
C4704 commonsourceibias.n49 gnd 0.009461f
C4705 commonsourceibias.n50 gnd 0.009461f
C4706 commonsourceibias.n51 gnd 0.012816f
C4707 commonsourceibias.n52 gnd 0.007653f
C4708 commonsourceibias.n53 gnd 0.012975f
C4709 commonsourceibias.n54 gnd 0.009461f
C4710 commonsourceibias.n55 gnd 0.009461f
C4711 commonsourceibias.n56 gnd 0.013054f
C4712 commonsourceibias.n57 gnd 0.011256f
C4713 commonsourceibias.n58 gnd 0.009134f
C4714 commonsourceibias.n59 gnd 0.009461f
C4715 commonsourceibias.n60 gnd 0.009461f
C4716 commonsourceibias.n61 gnd 0.011572f
C4717 commonsourceibias.n62 gnd 0.012989f
C4718 commonsourceibias.n63 gnd 0.070526f
C4719 commonsourceibias.n64 gnd 0.012901f
C4720 commonsourceibias.n65 gnd 0.009461f
C4721 commonsourceibias.n66 gnd 0.009461f
C4722 commonsourceibias.n67 gnd 0.009461f
C4723 commonsourceibias.n68 gnd 0.012901f
C4724 commonsourceibias.n69 gnd 0.070526f
C4725 commonsourceibias.n70 gnd 0.012989f
C4726 commonsourceibias.n71 gnd 0.011572f
C4727 commonsourceibias.n72 gnd 0.009461f
C4728 commonsourceibias.n73 gnd 0.009461f
C4729 commonsourceibias.n74 gnd 0.009461f
C4730 commonsourceibias.n75 gnd 0.011256f
C4731 commonsourceibias.n76 gnd 0.013054f
C4732 commonsourceibias.n77 gnd 0.070526f
C4733 commonsourceibias.n78 gnd 0.012975f
C4734 commonsourceibias.n79 gnd 0.009461f
C4735 commonsourceibias.n80 gnd 0.009461f
C4736 commonsourceibias.n81 gnd 0.009461f
C4737 commonsourceibias.n82 gnd 0.012816f
C4738 commonsourceibias.n83 gnd 0.070526f
C4739 commonsourceibias.n84 gnd 0.0129f
C4740 commonsourceibias.n85 gnd 0.011661f
C4741 commonsourceibias.n86 gnd 0.009461f
C4742 commonsourceibias.n87 gnd 0.009461f
C4743 commonsourceibias.n88 gnd 0.009461f
C4744 commonsourceibias.n89 gnd 0.010754f
C4745 commonsourceibias.n90 gnd 0.013093f
C4746 commonsourceibias.n91 gnd 0.070526f
C4747 commonsourceibias.n92 gnd 0.013037f
C4748 commonsourceibias.n93 gnd 0.009461f
C4749 commonsourceibias.n94 gnd 0.009461f
C4750 commonsourceibias.n95 gnd 0.009461f
C4751 commonsourceibias.n96 gnd 0.012717f
C4752 commonsourceibias.n97 gnd 0.070526f
C4753 commonsourceibias.n98 gnd 0.012748f
C4754 commonsourceibias.n99 gnd 0.085044f
C4755 commonsourceibias.n100 gnd 0.095092f
C4756 commonsourceibias.t55 gnd 0.020415f
C4757 commonsourceibias.t21 gnd 0.020415f
C4758 commonsourceibias.n101 gnd 0.180398f
C4759 commonsourceibias.n102 gnd 0.156264f
C4760 commonsourceibias.t5 gnd 0.020415f
C4761 commonsourceibias.t53 gnd 0.020415f
C4762 commonsourceibias.n103 gnd 0.180398f
C4763 commonsourceibias.n104 gnd 0.082864f
C4764 commonsourceibias.t15 gnd 0.020415f
C4765 commonsourceibias.t59 gnd 0.020415f
C4766 commonsourceibias.n105 gnd 0.180398f
C4767 commonsourceibias.n106 gnd 0.082864f
C4768 commonsourceibias.t33 gnd 0.020415f
C4769 commonsourceibias.t7 gnd 0.020415f
C4770 commonsourceibias.n107 gnd 0.180398f
C4771 commonsourceibias.n108 gnd 0.069229f
C4772 commonsourceibias.t23 gnd 0.020415f
C4773 commonsourceibias.t63 gnd 0.020415f
C4774 commonsourceibias.n109 gnd 0.181002f
C4775 commonsourceibias.t19 gnd 0.020415f
C4776 commonsourceibias.t61 gnd 0.020415f
C4777 commonsourceibias.n110 gnd 0.180398f
C4778 commonsourceibias.n111 gnd 0.168097f
C4779 commonsourceibias.t49 gnd 0.020415f
C4780 commonsourceibias.t35 gnd 0.020415f
C4781 commonsourceibias.n112 gnd 0.180398f
C4782 commonsourceibias.n113 gnd 0.082864f
C4783 commonsourceibias.t57 gnd 0.020415f
C4784 commonsourceibias.t29 gnd 0.020415f
C4785 commonsourceibias.n114 gnd 0.180398f
C4786 commonsourceibias.n115 gnd 0.069229f
C4787 commonsourceibias.n116 gnd 0.083829f
C4788 commonsourceibias.n117 gnd 0.009461f
C4789 commonsourceibias.t119 gnd 0.176757f
C4790 commonsourceibias.t79 gnd 0.176757f
C4791 commonsourceibias.n118 gnd 0.070526f
C4792 commonsourceibias.n119 gnd 0.009461f
C4793 commonsourceibias.t106 gnd 0.176757f
C4794 commonsourceibias.n120 gnd 0.070526f
C4795 commonsourceibias.n121 gnd 0.009461f
C4796 commonsourceibias.t96 gnd 0.176757f
C4797 commonsourceibias.n122 gnd 0.070526f
C4798 commonsourceibias.n123 gnd 0.009461f
C4799 commonsourceibias.t141 gnd 0.176757f
C4800 commonsourceibias.n124 gnd 0.010754f
C4801 commonsourceibias.n125 gnd 0.009461f
C4802 commonsourceibias.t116 gnd 0.176757f
C4803 commonsourceibias.n126 gnd 0.012717f
C4804 commonsourceibias.t129 gnd 0.196904f
C4805 commonsourceibias.t152 gnd 0.176757f
C4806 commonsourceibias.n127 gnd 0.078584f
C4807 commonsourceibias.n128 gnd 0.084191f
C4808 commonsourceibias.n129 gnd 0.04027f
C4809 commonsourceibias.n130 gnd 0.009461f
C4810 commonsourceibias.n131 gnd 0.00769f
C4811 commonsourceibias.n132 gnd 0.013037f
C4812 commonsourceibias.n133 gnd 0.070526f
C4813 commonsourceibias.n134 gnd 0.013093f
C4814 commonsourceibias.n135 gnd 0.009461f
C4815 commonsourceibias.n136 gnd 0.009461f
C4816 commonsourceibias.n137 gnd 0.009461f
C4817 commonsourceibias.n138 gnd 0.009597f
C4818 commonsourceibias.n139 gnd 0.070526f
C4819 commonsourceibias.n140 gnd 0.011661f
C4820 commonsourceibias.n141 gnd 0.0129f
C4821 commonsourceibias.n142 gnd 0.009461f
C4822 commonsourceibias.n143 gnd 0.009461f
C4823 commonsourceibias.n144 gnd 0.012816f
C4824 commonsourceibias.n145 gnd 0.007653f
C4825 commonsourceibias.n146 gnd 0.012975f
C4826 commonsourceibias.n147 gnd 0.009461f
C4827 commonsourceibias.n148 gnd 0.009461f
C4828 commonsourceibias.n149 gnd 0.013054f
C4829 commonsourceibias.n150 gnd 0.011256f
C4830 commonsourceibias.n151 gnd 0.009134f
C4831 commonsourceibias.n152 gnd 0.009461f
C4832 commonsourceibias.n153 gnd 0.009461f
C4833 commonsourceibias.n154 gnd 0.011572f
C4834 commonsourceibias.n155 gnd 0.012989f
C4835 commonsourceibias.n156 gnd 0.070526f
C4836 commonsourceibias.n157 gnd 0.012901f
C4837 commonsourceibias.n158 gnd 0.009415f
C4838 commonsourceibias.n159 gnd 0.06839f
C4839 commonsourceibias.n160 gnd 0.009415f
C4840 commonsourceibias.n161 gnd 0.012901f
C4841 commonsourceibias.n162 gnd 0.070526f
C4842 commonsourceibias.n163 gnd 0.012989f
C4843 commonsourceibias.n164 gnd 0.011572f
C4844 commonsourceibias.n165 gnd 0.009461f
C4845 commonsourceibias.n166 gnd 0.009461f
C4846 commonsourceibias.n167 gnd 0.009461f
C4847 commonsourceibias.n168 gnd 0.011256f
C4848 commonsourceibias.n169 gnd 0.013054f
C4849 commonsourceibias.n170 gnd 0.070526f
C4850 commonsourceibias.n171 gnd 0.012975f
C4851 commonsourceibias.n172 gnd 0.009461f
C4852 commonsourceibias.n173 gnd 0.009461f
C4853 commonsourceibias.n174 gnd 0.009461f
C4854 commonsourceibias.n175 gnd 0.012816f
C4855 commonsourceibias.n176 gnd 0.070526f
C4856 commonsourceibias.n177 gnd 0.0129f
C4857 commonsourceibias.n178 gnd 0.011661f
C4858 commonsourceibias.n179 gnd 0.009461f
C4859 commonsourceibias.n180 gnd 0.009461f
C4860 commonsourceibias.n181 gnd 0.009461f
C4861 commonsourceibias.n182 gnd 0.010754f
C4862 commonsourceibias.n183 gnd 0.013093f
C4863 commonsourceibias.n184 gnd 0.070526f
C4864 commonsourceibias.n185 gnd 0.013037f
C4865 commonsourceibias.n186 gnd 0.009461f
C4866 commonsourceibias.n187 gnd 0.009461f
C4867 commonsourceibias.n188 gnd 0.009461f
C4868 commonsourceibias.n189 gnd 0.012717f
C4869 commonsourceibias.n190 gnd 0.070526f
C4870 commonsourceibias.n191 gnd 0.012748f
C4871 commonsourceibias.n192 gnd 0.085044f
C4872 commonsourceibias.n193 gnd 0.056182f
C4873 commonsourceibias.n194 gnd 0.012624f
C4874 commonsourceibias.t68 gnd 0.191163f
C4875 commonsourceibias.t159 gnd 0.176757f
C4876 commonsourceibias.n195 gnd 0.00769f
C4877 commonsourceibias.n196 gnd 0.009461f
C4878 commonsourceibias.t148 gnd 0.176757f
C4879 commonsourceibias.n197 gnd 0.009597f
C4880 commonsourceibias.n198 gnd 0.009461f
C4881 commonsourceibias.t78 gnd 0.176757f
C4882 commonsourceibias.n199 gnd 0.070526f
C4883 commonsourceibias.t158 gnd 0.176757f
C4884 commonsourceibias.n200 gnd 0.007653f
C4885 commonsourceibias.n201 gnd 0.009461f
C4886 commonsourceibias.t85 gnd 0.176757f
C4887 commonsourceibias.n202 gnd 0.009134f
C4888 commonsourceibias.n203 gnd 0.009461f
C4889 commonsourceibias.t77 gnd 0.176757f
C4890 commonsourceibias.n204 gnd 0.070526f
C4891 commonsourceibias.t157 gnd 0.176757f
C4892 commonsourceibias.n205 gnd 0.007641f
C4893 commonsourceibias.n206 gnd 0.009461f
C4894 commonsourceibias.t94 gnd 0.176757f
C4895 commonsourceibias.t113 gnd 0.176757f
C4896 commonsourceibias.n207 gnd 0.070526f
C4897 commonsourceibias.n208 gnd 0.009461f
C4898 commonsourceibias.t156 gnd 0.176757f
C4899 commonsourceibias.n209 gnd 0.070526f
C4900 commonsourceibias.n210 gnd 0.009461f
C4901 commonsourceibias.t92 gnd 0.176757f
C4902 commonsourceibias.n211 gnd 0.070526f
C4903 commonsourceibias.n212 gnd 0.009461f
C4904 commonsourceibias.t109 gnd 0.176757f
C4905 commonsourceibias.n213 gnd 0.010754f
C4906 commonsourceibias.n214 gnd 0.009461f
C4907 commonsourceibias.t105 gnd 0.176757f
C4908 commonsourceibias.n215 gnd 0.012717f
C4909 commonsourceibias.t108 gnd 0.196904f
C4910 commonsourceibias.t91 gnd 0.176757f
C4911 commonsourceibias.n216 gnd 0.078584f
C4912 commonsourceibias.n217 gnd 0.084191f
C4913 commonsourceibias.n218 gnd 0.04027f
C4914 commonsourceibias.n219 gnd 0.009461f
C4915 commonsourceibias.n220 gnd 0.00769f
C4916 commonsourceibias.n221 gnd 0.013037f
C4917 commonsourceibias.n222 gnd 0.070526f
C4918 commonsourceibias.n223 gnd 0.013093f
C4919 commonsourceibias.n224 gnd 0.009461f
C4920 commonsourceibias.n225 gnd 0.009461f
C4921 commonsourceibias.n226 gnd 0.009461f
C4922 commonsourceibias.n227 gnd 0.009597f
C4923 commonsourceibias.n228 gnd 0.070526f
C4924 commonsourceibias.n229 gnd 0.011661f
C4925 commonsourceibias.n230 gnd 0.0129f
C4926 commonsourceibias.n231 gnd 0.009461f
C4927 commonsourceibias.n232 gnd 0.009461f
C4928 commonsourceibias.n233 gnd 0.012816f
C4929 commonsourceibias.n234 gnd 0.007653f
C4930 commonsourceibias.n235 gnd 0.012975f
C4931 commonsourceibias.n236 gnd 0.009461f
C4932 commonsourceibias.n237 gnd 0.009461f
C4933 commonsourceibias.n238 gnd 0.013054f
C4934 commonsourceibias.n239 gnd 0.011256f
C4935 commonsourceibias.n240 gnd 0.009134f
C4936 commonsourceibias.n241 gnd 0.009461f
C4937 commonsourceibias.n242 gnd 0.009461f
C4938 commonsourceibias.n243 gnd 0.011572f
C4939 commonsourceibias.n244 gnd 0.012989f
C4940 commonsourceibias.n245 gnd 0.070526f
C4941 commonsourceibias.n246 gnd 0.012901f
C4942 commonsourceibias.n247 gnd 0.009461f
C4943 commonsourceibias.n248 gnd 0.009461f
C4944 commonsourceibias.n249 gnd 0.009461f
C4945 commonsourceibias.n250 gnd 0.012901f
C4946 commonsourceibias.n251 gnd 0.070526f
C4947 commonsourceibias.n252 gnd 0.012989f
C4948 commonsourceibias.n253 gnd 0.011572f
C4949 commonsourceibias.n254 gnd 0.009461f
C4950 commonsourceibias.n255 gnd 0.009461f
C4951 commonsourceibias.n256 gnd 0.009461f
C4952 commonsourceibias.n257 gnd 0.011256f
C4953 commonsourceibias.n258 gnd 0.013054f
C4954 commonsourceibias.n259 gnd 0.070526f
C4955 commonsourceibias.n260 gnd 0.012975f
C4956 commonsourceibias.n261 gnd 0.009461f
C4957 commonsourceibias.n262 gnd 0.009461f
C4958 commonsourceibias.n263 gnd 0.009461f
C4959 commonsourceibias.n264 gnd 0.012816f
C4960 commonsourceibias.n265 gnd 0.070526f
C4961 commonsourceibias.n266 gnd 0.0129f
C4962 commonsourceibias.n267 gnd 0.011661f
C4963 commonsourceibias.n268 gnd 0.009461f
C4964 commonsourceibias.n269 gnd 0.009461f
C4965 commonsourceibias.n270 gnd 0.009461f
C4966 commonsourceibias.n271 gnd 0.010754f
C4967 commonsourceibias.n272 gnd 0.013093f
C4968 commonsourceibias.n273 gnd 0.070526f
C4969 commonsourceibias.n274 gnd 0.013037f
C4970 commonsourceibias.n275 gnd 0.009461f
C4971 commonsourceibias.n276 gnd 0.009461f
C4972 commonsourceibias.n277 gnd 0.009461f
C4973 commonsourceibias.n278 gnd 0.012717f
C4974 commonsourceibias.n279 gnd 0.070526f
C4975 commonsourceibias.n280 gnd 0.012748f
C4976 commonsourceibias.n281 gnd 0.085044f
C4977 commonsourceibias.n282 gnd 0.030348f
C4978 commonsourceibias.n283 gnd 0.15151f
C4979 commonsourceibias.n284 gnd 0.012624f
C4980 commonsourceibias.t75 gnd 0.176757f
C4981 commonsourceibias.n285 gnd 0.00769f
C4982 commonsourceibias.n286 gnd 0.009461f
C4983 commonsourceibias.t128 gnd 0.176757f
C4984 commonsourceibias.n287 gnd 0.009597f
C4985 commonsourceibias.n288 gnd 0.009461f
C4986 commonsourceibias.t124 gnd 0.176757f
C4987 commonsourceibias.n289 gnd 0.070526f
C4988 commonsourceibias.t155 gnd 0.176757f
C4989 commonsourceibias.n290 gnd 0.007653f
C4990 commonsourceibias.n291 gnd 0.009461f
C4991 commonsourceibias.t89 gnd 0.176757f
C4992 commonsourceibias.n292 gnd 0.009134f
C4993 commonsourceibias.n293 gnd 0.009461f
C4994 commonsourceibias.t118 gnd 0.176757f
C4995 commonsourceibias.n294 gnd 0.070526f
C4996 commonsourceibias.t146 gnd 0.176757f
C4997 commonsourceibias.n295 gnd 0.007641f
C4998 commonsourceibias.n296 gnd 0.009461f
C4999 commonsourceibias.t138 gnd 0.176757f
C5000 commonsourceibias.t64 gnd 0.176757f
C5001 commonsourceibias.n297 gnd 0.070526f
C5002 commonsourceibias.n298 gnd 0.009461f
C5003 commonsourceibias.t137 gnd 0.176757f
C5004 commonsourceibias.n299 gnd 0.070526f
C5005 commonsourceibias.n300 gnd 0.009461f
C5006 commonsourceibias.t133 gnd 0.176757f
C5007 commonsourceibias.n301 gnd 0.070526f
C5008 commonsourceibias.n302 gnd 0.009461f
C5009 commonsourceibias.t149 gnd 0.176757f
C5010 commonsourceibias.n303 gnd 0.010754f
C5011 commonsourceibias.n304 gnd 0.009461f
C5012 commonsourceibias.t76 gnd 0.176757f
C5013 commonsourceibias.n305 gnd 0.012717f
C5014 commonsourceibias.t139 gnd 0.196904f
C5015 commonsourceibias.t130 gnd 0.176757f
C5016 commonsourceibias.n306 gnd 0.078584f
C5017 commonsourceibias.n307 gnd 0.084191f
C5018 commonsourceibias.n308 gnd 0.04027f
C5019 commonsourceibias.n309 gnd 0.009461f
C5020 commonsourceibias.n310 gnd 0.00769f
C5021 commonsourceibias.n311 gnd 0.013037f
C5022 commonsourceibias.n312 gnd 0.070526f
C5023 commonsourceibias.n313 gnd 0.013093f
C5024 commonsourceibias.n314 gnd 0.009461f
C5025 commonsourceibias.n315 gnd 0.009461f
C5026 commonsourceibias.n316 gnd 0.009461f
C5027 commonsourceibias.n317 gnd 0.009597f
C5028 commonsourceibias.n318 gnd 0.070526f
C5029 commonsourceibias.n319 gnd 0.011661f
C5030 commonsourceibias.n320 gnd 0.0129f
C5031 commonsourceibias.n321 gnd 0.009461f
C5032 commonsourceibias.n322 gnd 0.009461f
C5033 commonsourceibias.n323 gnd 0.012816f
C5034 commonsourceibias.n324 gnd 0.007653f
C5035 commonsourceibias.n325 gnd 0.012975f
C5036 commonsourceibias.n326 gnd 0.009461f
C5037 commonsourceibias.n327 gnd 0.009461f
C5038 commonsourceibias.n328 gnd 0.013054f
C5039 commonsourceibias.n329 gnd 0.011256f
C5040 commonsourceibias.n330 gnd 0.009134f
C5041 commonsourceibias.n331 gnd 0.009461f
C5042 commonsourceibias.n332 gnd 0.009461f
C5043 commonsourceibias.n333 gnd 0.011572f
C5044 commonsourceibias.n334 gnd 0.012989f
C5045 commonsourceibias.n335 gnd 0.070526f
C5046 commonsourceibias.n336 gnd 0.012901f
C5047 commonsourceibias.n337 gnd 0.009461f
C5048 commonsourceibias.n338 gnd 0.009461f
C5049 commonsourceibias.n339 gnd 0.009461f
C5050 commonsourceibias.n340 gnd 0.012901f
C5051 commonsourceibias.n341 gnd 0.070526f
C5052 commonsourceibias.n342 gnd 0.012989f
C5053 commonsourceibias.n343 gnd 0.011572f
C5054 commonsourceibias.n344 gnd 0.009461f
C5055 commonsourceibias.n345 gnd 0.009461f
C5056 commonsourceibias.n346 gnd 0.009461f
C5057 commonsourceibias.n347 gnd 0.011256f
C5058 commonsourceibias.n348 gnd 0.013054f
C5059 commonsourceibias.n349 gnd 0.070526f
C5060 commonsourceibias.n350 gnd 0.012975f
C5061 commonsourceibias.n351 gnd 0.009461f
C5062 commonsourceibias.n352 gnd 0.009461f
C5063 commonsourceibias.n353 gnd 0.009461f
C5064 commonsourceibias.n354 gnd 0.012816f
C5065 commonsourceibias.n355 gnd 0.070526f
C5066 commonsourceibias.n356 gnd 0.0129f
C5067 commonsourceibias.n357 gnd 0.011661f
C5068 commonsourceibias.n358 gnd 0.009461f
C5069 commonsourceibias.n359 gnd 0.009461f
C5070 commonsourceibias.n360 gnd 0.009461f
C5071 commonsourceibias.n361 gnd 0.010754f
C5072 commonsourceibias.n362 gnd 0.013093f
C5073 commonsourceibias.n363 gnd 0.070526f
C5074 commonsourceibias.n364 gnd 0.013037f
C5075 commonsourceibias.n365 gnd 0.009461f
C5076 commonsourceibias.n366 gnd 0.009461f
C5077 commonsourceibias.n367 gnd 0.009461f
C5078 commonsourceibias.n368 gnd 0.012717f
C5079 commonsourceibias.n369 gnd 0.070526f
C5080 commonsourceibias.n370 gnd 0.012748f
C5081 commonsourceibias.t147 gnd 0.191163f
C5082 commonsourceibias.n371 gnd 0.085044f
C5083 commonsourceibias.n372 gnd 0.030348f
C5084 commonsourceibias.n373 gnd 0.449685f
C5085 commonsourceibias.n374 gnd 0.012624f
C5086 commonsourceibias.t93 gnd 0.191163f
C5087 commonsourceibias.t134 gnd 0.176757f
C5088 commonsourceibias.n375 gnd 0.00769f
C5089 commonsourceibias.n376 gnd 0.009461f
C5090 commonsourceibias.t114 gnd 0.176757f
C5091 commonsourceibias.n377 gnd 0.009597f
C5092 commonsourceibias.n378 gnd 0.009461f
C5093 commonsourceibias.t123 gnd 0.176757f
C5094 commonsourceibias.n379 gnd 0.007653f
C5095 commonsourceibias.n380 gnd 0.009461f
C5096 commonsourceibias.t88 gnd 0.176757f
C5097 commonsourceibias.n381 gnd 0.009134f
C5098 commonsourceibias.n382 gnd 0.009461f
C5099 commonsourceibias.t104 gnd 0.176757f
C5100 commonsourceibias.n383 gnd 0.007641f
C5101 commonsourceibias.n384 gnd 0.009461f
C5102 commonsourceibias.t90 gnd 0.176757f
C5103 commonsourceibias.t140 gnd 0.176757f
C5104 commonsourceibias.n385 gnd 0.070526f
C5105 commonsourceibias.n386 gnd 0.009461f
C5106 commonsourceibias.t83 gnd 0.176757f
C5107 commonsourceibias.n387 gnd 0.070526f
C5108 commonsourceibias.n388 gnd 0.009461f
C5109 commonsourceibias.t151 gnd 0.176757f
C5110 commonsourceibias.n389 gnd 0.070526f
C5111 commonsourceibias.n390 gnd 0.009461f
C5112 commonsourceibias.t127 gnd 0.176757f
C5113 commonsourceibias.n391 gnd 0.010754f
C5114 commonsourceibias.n392 gnd 0.009461f
C5115 commonsourceibias.t84 gnd 0.176757f
C5116 commonsourceibias.n393 gnd 0.012717f
C5117 commonsourceibias.t112 gnd 0.196904f
C5118 commonsourceibias.t131 gnd 0.176757f
C5119 commonsourceibias.n394 gnd 0.078584f
C5120 commonsourceibias.n395 gnd 0.084191f
C5121 commonsourceibias.n396 gnd 0.04027f
C5122 commonsourceibias.n397 gnd 0.009461f
C5123 commonsourceibias.n398 gnd 0.00769f
C5124 commonsourceibias.n399 gnd 0.013037f
C5125 commonsourceibias.n400 gnd 0.070526f
C5126 commonsourceibias.n401 gnd 0.013093f
C5127 commonsourceibias.n402 gnd 0.009461f
C5128 commonsourceibias.n403 gnd 0.009461f
C5129 commonsourceibias.n404 gnd 0.009461f
C5130 commonsourceibias.n405 gnd 0.009597f
C5131 commonsourceibias.n406 gnd 0.070526f
C5132 commonsourceibias.n407 gnd 0.011661f
C5133 commonsourceibias.n408 gnd 0.0129f
C5134 commonsourceibias.n409 gnd 0.009461f
C5135 commonsourceibias.n410 gnd 0.009461f
C5136 commonsourceibias.n411 gnd 0.012816f
C5137 commonsourceibias.n412 gnd 0.007653f
C5138 commonsourceibias.n413 gnd 0.012975f
C5139 commonsourceibias.n414 gnd 0.009461f
C5140 commonsourceibias.n415 gnd 0.009461f
C5141 commonsourceibias.n416 gnd 0.013054f
C5142 commonsourceibias.n417 gnd 0.011256f
C5143 commonsourceibias.n418 gnd 0.009134f
C5144 commonsourceibias.n419 gnd 0.009461f
C5145 commonsourceibias.n420 gnd 0.009461f
C5146 commonsourceibias.n421 gnd 0.011572f
C5147 commonsourceibias.n422 gnd 0.012989f
C5148 commonsourceibias.n423 gnd 0.070526f
C5149 commonsourceibias.n424 gnd 0.012901f
C5150 commonsourceibias.n425 gnd 0.009415f
C5151 commonsourceibias.t47 gnd 0.020415f
C5152 commonsourceibias.t9 gnd 0.020415f
C5153 commonsourceibias.n426 gnd 0.181002f
C5154 commonsourceibias.t25 gnd 0.020415f
C5155 commonsourceibias.t3 gnd 0.020415f
C5156 commonsourceibias.n427 gnd 0.180398f
C5157 commonsourceibias.n428 gnd 0.168097f
C5158 commonsourceibias.t17 gnd 0.020415f
C5159 commonsourceibias.t27 gnd 0.020415f
C5160 commonsourceibias.n429 gnd 0.180398f
C5161 commonsourceibias.n430 gnd 0.082864f
C5162 commonsourceibias.t13 gnd 0.020415f
C5163 commonsourceibias.t41 gnd 0.020415f
C5164 commonsourceibias.n431 gnd 0.180398f
C5165 commonsourceibias.n432 gnd 0.069229f
C5166 commonsourceibias.n433 gnd 0.012624f
C5167 commonsourceibias.t10 gnd 0.176757f
C5168 commonsourceibias.n434 gnd 0.00769f
C5169 commonsourceibias.n435 gnd 0.009461f
C5170 commonsourceibias.t44 gnd 0.176757f
C5171 commonsourceibias.n436 gnd 0.009597f
C5172 commonsourceibias.n437 gnd 0.009461f
C5173 commonsourceibias.t0 gnd 0.176757f
C5174 commonsourceibias.n438 gnd 0.007653f
C5175 commonsourceibias.n439 gnd 0.009461f
C5176 commonsourceibias.t42 gnd 0.176757f
C5177 commonsourceibias.n440 gnd 0.009134f
C5178 commonsourceibias.n441 gnd 0.009461f
C5179 commonsourceibias.t50 gnd 0.176757f
C5180 commonsourceibias.n442 gnd 0.007641f
C5181 commonsourceibias.n443 gnd 0.009461f
C5182 commonsourceibias.t40 gnd 0.176757f
C5183 commonsourceibias.t12 gnd 0.176757f
C5184 commonsourceibias.n444 gnd 0.070526f
C5185 commonsourceibias.n445 gnd 0.009461f
C5186 commonsourceibias.t26 gnd 0.176757f
C5187 commonsourceibias.n446 gnd 0.070526f
C5188 commonsourceibias.n447 gnd 0.009461f
C5189 commonsourceibias.t16 gnd 0.176757f
C5190 commonsourceibias.n448 gnd 0.070526f
C5191 commonsourceibias.n449 gnd 0.009461f
C5192 commonsourceibias.t2 gnd 0.176757f
C5193 commonsourceibias.n450 gnd 0.010754f
C5194 commonsourceibias.n451 gnd 0.009461f
C5195 commonsourceibias.t24 gnd 0.176757f
C5196 commonsourceibias.n452 gnd 0.012717f
C5197 commonsourceibias.t46 gnd 0.196904f
C5198 commonsourceibias.t8 gnd 0.176757f
C5199 commonsourceibias.n453 gnd 0.078584f
C5200 commonsourceibias.n454 gnd 0.084191f
C5201 commonsourceibias.n455 gnd 0.04027f
C5202 commonsourceibias.n456 gnd 0.009461f
C5203 commonsourceibias.n457 gnd 0.00769f
C5204 commonsourceibias.n458 gnd 0.013037f
C5205 commonsourceibias.n459 gnd 0.070526f
C5206 commonsourceibias.n460 gnd 0.013093f
C5207 commonsourceibias.n461 gnd 0.009461f
C5208 commonsourceibias.n462 gnd 0.009461f
C5209 commonsourceibias.n463 gnd 0.009461f
C5210 commonsourceibias.n464 gnd 0.009597f
C5211 commonsourceibias.n465 gnd 0.070526f
C5212 commonsourceibias.n466 gnd 0.011661f
C5213 commonsourceibias.n467 gnd 0.0129f
C5214 commonsourceibias.n468 gnd 0.009461f
C5215 commonsourceibias.n469 gnd 0.009461f
C5216 commonsourceibias.n470 gnd 0.012816f
C5217 commonsourceibias.n471 gnd 0.007653f
C5218 commonsourceibias.n472 gnd 0.012975f
C5219 commonsourceibias.n473 gnd 0.009461f
C5220 commonsourceibias.n474 gnd 0.009461f
C5221 commonsourceibias.n475 gnd 0.013054f
C5222 commonsourceibias.n476 gnd 0.011256f
C5223 commonsourceibias.n477 gnd 0.009134f
C5224 commonsourceibias.n478 gnd 0.009461f
C5225 commonsourceibias.n479 gnd 0.009461f
C5226 commonsourceibias.n480 gnd 0.011572f
C5227 commonsourceibias.n481 gnd 0.012989f
C5228 commonsourceibias.n482 gnd 0.070526f
C5229 commonsourceibias.n483 gnd 0.012901f
C5230 commonsourceibias.n484 gnd 0.009461f
C5231 commonsourceibias.n485 gnd 0.009461f
C5232 commonsourceibias.n486 gnd 0.009461f
C5233 commonsourceibias.n487 gnd 0.012901f
C5234 commonsourceibias.n488 gnd 0.070526f
C5235 commonsourceibias.n489 gnd 0.012989f
C5236 commonsourceibias.t30 gnd 0.176757f
C5237 commonsourceibias.n490 gnd 0.070526f
C5238 commonsourceibias.n491 gnd 0.011572f
C5239 commonsourceibias.n492 gnd 0.009461f
C5240 commonsourceibias.n493 gnd 0.009461f
C5241 commonsourceibias.n494 gnd 0.009461f
C5242 commonsourceibias.n495 gnd 0.011256f
C5243 commonsourceibias.n496 gnd 0.013054f
C5244 commonsourceibias.n497 gnd 0.070526f
C5245 commonsourceibias.n498 gnd 0.012975f
C5246 commonsourceibias.n499 gnd 0.009461f
C5247 commonsourceibias.n500 gnd 0.009461f
C5248 commonsourceibias.n501 gnd 0.009461f
C5249 commonsourceibias.n502 gnd 0.012816f
C5250 commonsourceibias.n503 gnd 0.070526f
C5251 commonsourceibias.n504 gnd 0.0129f
C5252 commonsourceibias.t36 gnd 0.176757f
C5253 commonsourceibias.n505 gnd 0.070526f
C5254 commonsourceibias.n506 gnd 0.011661f
C5255 commonsourceibias.n507 gnd 0.009461f
C5256 commonsourceibias.n508 gnd 0.009461f
C5257 commonsourceibias.n509 gnd 0.009461f
C5258 commonsourceibias.n510 gnd 0.010754f
C5259 commonsourceibias.n511 gnd 0.013093f
C5260 commonsourceibias.n512 gnd 0.070526f
C5261 commonsourceibias.n513 gnd 0.013037f
C5262 commonsourceibias.n514 gnd 0.009461f
C5263 commonsourceibias.n515 gnd 0.009461f
C5264 commonsourceibias.n516 gnd 0.009461f
C5265 commonsourceibias.n517 gnd 0.012717f
C5266 commonsourceibias.n518 gnd 0.070526f
C5267 commonsourceibias.n519 gnd 0.012748f
C5268 commonsourceibias.t38 gnd 0.191163f
C5269 commonsourceibias.n520 gnd 0.085044f
C5270 commonsourceibias.n521 gnd 0.095092f
C5271 commonsourceibias.t11 gnd 0.020415f
C5272 commonsourceibias.t39 gnd 0.020415f
C5273 commonsourceibias.n522 gnd 0.180398f
C5274 commonsourceibias.n523 gnd 0.156264f
C5275 commonsourceibias.t37 gnd 0.020415f
C5276 commonsourceibias.t45 gnd 0.020415f
C5277 commonsourceibias.n524 gnd 0.180398f
C5278 commonsourceibias.n525 gnd 0.082864f
C5279 commonsourceibias.t43 gnd 0.020415f
C5280 commonsourceibias.t1 gnd 0.020415f
C5281 commonsourceibias.n526 gnd 0.180398f
C5282 commonsourceibias.n527 gnd 0.082864f
C5283 commonsourceibias.t51 gnd 0.020415f
C5284 commonsourceibias.t31 gnd 0.020415f
C5285 commonsourceibias.n528 gnd 0.180398f
C5286 commonsourceibias.n529 gnd 0.069229f
C5287 commonsourceibias.n530 gnd 0.083829f
C5288 commonsourceibias.n531 gnd 0.06839f
C5289 commonsourceibias.n532 gnd 0.009415f
C5290 commonsourceibias.n533 gnd 0.012901f
C5291 commonsourceibias.n534 gnd 0.070526f
C5292 commonsourceibias.n535 gnd 0.012989f
C5293 commonsourceibias.t74 gnd 0.176757f
C5294 commonsourceibias.n536 gnd 0.070526f
C5295 commonsourceibias.n537 gnd 0.011572f
C5296 commonsourceibias.n538 gnd 0.009461f
C5297 commonsourceibias.n539 gnd 0.009461f
C5298 commonsourceibias.n540 gnd 0.009461f
C5299 commonsourceibias.n541 gnd 0.011256f
C5300 commonsourceibias.n542 gnd 0.013054f
C5301 commonsourceibias.n543 gnd 0.070526f
C5302 commonsourceibias.n544 gnd 0.012975f
C5303 commonsourceibias.n545 gnd 0.009461f
C5304 commonsourceibias.n546 gnd 0.009461f
C5305 commonsourceibias.n547 gnd 0.009461f
C5306 commonsourceibias.n548 gnd 0.012816f
C5307 commonsourceibias.n549 gnd 0.070526f
C5308 commonsourceibias.n550 gnd 0.0129f
C5309 commonsourceibias.t95 gnd 0.176757f
C5310 commonsourceibias.n551 gnd 0.070526f
C5311 commonsourceibias.n552 gnd 0.011661f
C5312 commonsourceibias.n553 gnd 0.009461f
C5313 commonsourceibias.n554 gnd 0.009461f
C5314 commonsourceibias.n555 gnd 0.009461f
C5315 commonsourceibias.n556 gnd 0.010754f
C5316 commonsourceibias.n557 gnd 0.013093f
C5317 commonsourceibias.n558 gnd 0.070526f
C5318 commonsourceibias.n559 gnd 0.013037f
C5319 commonsourceibias.n560 gnd 0.009461f
C5320 commonsourceibias.n561 gnd 0.009461f
C5321 commonsourceibias.n562 gnd 0.009461f
C5322 commonsourceibias.n563 gnd 0.012717f
C5323 commonsourceibias.n564 gnd 0.070526f
C5324 commonsourceibias.n565 gnd 0.012748f
C5325 commonsourceibias.n566 gnd 0.085044f
C5326 commonsourceibias.n567 gnd 0.056182f
C5327 commonsourceibias.n568 gnd 0.012624f
C5328 commonsourceibias.t142 gnd 0.176757f
C5329 commonsourceibias.n569 gnd 0.00769f
C5330 commonsourceibias.n570 gnd 0.009461f
C5331 commonsourceibias.t66 gnd 0.176757f
C5332 commonsourceibias.n571 gnd 0.009597f
C5333 commonsourceibias.n572 gnd 0.009461f
C5334 commonsourceibias.t143 gnd 0.176757f
C5335 commonsourceibias.n573 gnd 0.007653f
C5336 commonsourceibias.n574 gnd 0.009461f
C5337 commonsourceibias.t67 gnd 0.176757f
C5338 commonsourceibias.n575 gnd 0.009134f
C5339 commonsourceibias.n576 gnd 0.009461f
C5340 commonsourceibias.t144 gnd 0.176757f
C5341 commonsourceibias.n577 gnd 0.007641f
C5342 commonsourceibias.n578 gnd 0.009461f
C5343 commonsourceibias.t70 gnd 0.176757f
C5344 commonsourceibias.t101 gnd 0.176757f
C5345 commonsourceibias.n579 gnd 0.070526f
C5346 commonsourceibias.n580 gnd 0.009461f
C5347 commonsourceibias.t80 gnd 0.176757f
C5348 commonsourceibias.n581 gnd 0.070526f
C5349 commonsourceibias.n582 gnd 0.009461f
C5350 commonsourceibias.t72 gnd 0.176757f
C5351 commonsourceibias.n583 gnd 0.070526f
C5352 commonsourceibias.n584 gnd 0.009461f
C5353 commonsourceibias.t100 gnd 0.176757f
C5354 commonsourceibias.n585 gnd 0.010754f
C5355 commonsourceibias.n586 gnd 0.009461f
C5356 commonsourceibias.t87 gnd 0.176757f
C5357 commonsourceibias.n587 gnd 0.012717f
C5358 commonsourceibias.t99 gnd 0.196904f
C5359 commonsourceibias.t71 gnd 0.176757f
C5360 commonsourceibias.n588 gnd 0.078584f
C5361 commonsourceibias.n589 gnd 0.084191f
C5362 commonsourceibias.n590 gnd 0.04027f
C5363 commonsourceibias.n591 gnd 0.009461f
C5364 commonsourceibias.n592 gnd 0.00769f
C5365 commonsourceibias.n593 gnd 0.013037f
C5366 commonsourceibias.n594 gnd 0.070526f
C5367 commonsourceibias.n595 gnd 0.013093f
C5368 commonsourceibias.n596 gnd 0.009461f
C5369 commonsourceibias.n597 gnd 0.009461f
C5370 commonsourceibias.n598 gnd 0.009461f
C5371 commonsourceibias.n599 gnd 0.009597f
C5372 commonsourceibias.n600 gnd 0.070526f
C5373 commonsourceibias.n601 gnd 0.011661f
C5374 commonsourceibias.n602 gnd 0.0129f
C5375 commonsourceibias.n603 gnd 0.009461f
C5376 commonsourceibias.n604 gnd 0.009461f
C5377 commonsourceibias.n605 gnd 0.012816f
C5378 commonsourceibias.n606 gnd 0.007653f
C5379 commonsourceibias.n607 gnd 0.012975f
C5380 commonsourceibias.n608 gnd 0.009461f
C5381 commonsourceibias.n609 gnd 0.009461f
C5382 commonsourceibias.n610 gnd 0.013054f
C5383 commonsourceibias.n611 gnd 0.011256f
C5384 commonsourceibias.n612 gnd 0.009134f
C5385 commonsourceibias.n613 gnd 0.009461f
C5386 commonsourceibias.n614 gnd 0.009461f
C5387 commonsourceibias.n615 gnd 0.011572f
C5388 commonsourceibias.n616 gnd 0.012989f
C5389 commonsourceibias.n617 gnd 0.070526f
C5390 commonsourceibias.n618 gnd 0.012901f
C5391 commonsourceibias.n619 gnd 0.009461f
C5392 commonsourceibias.n620 gnd 0.009461f
C5393 commonsourceibias.n621 gnd 0.009461f
C5394 commonsourceibias.n622 gnd 0.012901f
C5395 commonsourceibias.n623 gnd 0.070526f
C5396 commonsourceibias.n624 gnd 0.012989f
C5397 commonsourceibias.t98 gnd 0.176757f
C5398 commonsourceibias.n625 gnd 0.070526f
C5399 commonsourceibias.n626 gnd 0.011572f
C5400 commonsourceibias.n627 gnd 0.009461f
C5401 commonsourceibias.n628 gnd 0.009461f
C5402 commonsourceibias.n629 gnd 0.009461f
C5403 commonsourceibias.n630 gnd 0.011256f
C5404 commonsourceibias.n631 gnd 0.013054f
C5405 commonsourceibias.n632 gnd 0.070526f
C5406 commonsourceibias.n633 gnd 0.012975f
C5407 commonsourceibias.n634 gnd 0.009461f
C5408 commonsourceibias.n635 gnd 0.009461f
C5409 commonsourceibias.n636 gnd 0.009461f
C5410 commonsourceibias.n637 gnd 0.012816f
C5411 commonsourceibias.n638 gnd 0.070526f
C5412 commonsourceibias.n639 gnd 0.0129f
C5413 commonsourceibias.t154 gnd 0.176757f
C5414 commonsourceibias.n640 gnd 0.070526f
C5415 commonsourceibias.n641 gnd 0.011661f
C5416 commonsourceibias.n642 gnd 0.009461f
C5417 commonsourceibias.n643 gnd 0.009461f
C5418 commonsourceibias.n644 gnd 0.009461f
C5419 commonsourceibias.n645 gnd 0.010754f
C5420 commonsourceibias.n646 gnd 0.013093f
C5421 commonsourceibias.n647 gnd 0.070526f
C5422 commonsourceibias.n648 gnd 0.013037f
C5423 commonsourceibias.n649 gnd 0.009461f
C5424 commonsourceibias.n650 gnd 0.009461f
C5425 commonsourceibias.n651 gnd 0.009461f
C5426 commonsourceibias.n652 gnd 0.012717f
C5427 commonsourceibias.n653 gnd 0.070526f
C5428 commonsourceibias.n654 gnd 0.012748f
C5429 commonsourceibias.t150 gnd 0.191163f
C5430 commonsourceibias.n655 gnd 0.085044f
C5431 commonsourceibias.n656 gnd 0.030348f
C5432 commonsourceibias.n657 gnd 0.15151f
C5433 commonsourceibias.n658 gnd 0.012624f
C5434 commonsourceibias.t107 gnd 0.176757f
C5435 commonsourceibias.n659 gnd 0.00769f
C5436 commonsourceibias.n660 gnd 0.009461f
C5437 commonsourceibias.t122 gnd 0.176757f
C5438 commonsourceibias.n661 gnd 0.009597f
C5439 commonsourceibias.n662 gnd 0.009461f
C5440 commonsourceibias.t97 gnd 0.176757f
C5441 commonsourceibias.n663 gnd 0.007653f
C5442 commonsourceibias.n664 gnd 0.009461f
C5443 commonsourceibias.t115 gnd 0.176757f
C5444 commonsourceibias.n665 gnd 0.009134f
C5445 commonsourceibias.n666 gnd 0.009461f
C5446 commonsourceibias.t81 gnd 0.176757f
C5447 commonsourceibias.n667 gnd 0.007641f
C5448 commonsourceibias.n668 gnd 0.009461f
C5449 commonsourceibias.t69 gnd 0.176757f
C5450 commonsourceibias.t103 gnd 0.176757f
C5451 commonsourceibias.n669 gnd 0.070526f
C5452 commonsourceibias.n670 gnd 0.009461f
C5453 commonsourceibias.t132 gnd 0.176757f
C5454 commonsourceibias.n671 gnd 0.070526f
C5455 commonsourceibias.n672 gnd 0.009461f
C5456 commonsourceibias.t153 gnd 0.176757f
C5457 commonsourceibias.n673 gnd 0.070526f
C5458 commonsourceibias.n674 gnd 0.009461f
C5459 commonsourceibias.t86 gnd 0.176757f
C5460 commonsourceibias.n675 gnd 0.010754f
C5461 commonsourceibias.n676 gnd 0.009461f
C5462 commonsourceibias.t111 gnd 0.176757f
C5463 commonsourceibias.n677 gnd 0.012717f
C5464 commonsourceibias.t73 gnd 0.196904f
C5465 commonsourceibias.t145 gnd 0.176757f
C5466 commonsourceibias.n678 gnd 0.078584f
C5467 commonsourceibias.n679 gnd 0.084191f
C5468 commonsourceibias.n680 gnd 0.04027f
C5469 commonsourceibias.n681 gnd 0.009461f
C5470 commonsourceibias.n682 gnd 0.00769f
C5471 commonsourceibias.n683 gnd 0.013037f
C5472 commonsourceibias.n684 gnd 0.070526f
C5473 commonsourceibias.n685 gnd 0.013093f
C5474 commonsourceibias.n686 gnd 0.009461f
C5475 commonsourceibias.n687 gnd 0.009461f
C5476 commonsourceibias.n688 gnd 0.009461f
C5477 commonsourceibias.n689 gnd 0.009597f
C5478 commonsourceibias.n690 gnd 0.070526f
C5479 commonsourceibias.n691 gnd 0.011661f
C5480 commonsourceibias.n692 gnd 0.0129f
C5481 commonsourceibias.n693 gnd 0.009461f
C5482 commonsourceibias.n694 gnd 0.009461f
C5483 commonsourceibias.n695 gnd 0.012816f
C5484 commonsourceibias.n696 gnd 0.007653f
C5485 commonsourceibias.n697 gnd 0.012975f
C5486 commonsourceibias.n698 gnd 0.009461f
C5487 commonsourceibias.n699 gnd 0.009461f
C5488 commonsourceibias.n700 gnd 0.013054f
C5489 commonsourceibias.n701 gnd 0.011256f
C5490 commonsourceibias.n702 gnd 0.009134f
C5491 commonsourceibias.n703 gnd 0.009461f
C5492 commonsourceibias.n704 gnd 0.009461f
C5493 commonsourceibias.n705 gnd 0.011572f
C5494 commonsourceibias.n706 gnd 0.012989f
C5495 commonsourceibias.n707 gnd 0.070526f
C5496 commonsourceibias.n708 gnd 0.012901f
C5497 commonsourceibias.n709 gnd 0.009461f
C5498 commonsourceibias.n710 gnd 0.009461f
C5499 commonsourceibias.n711 gnd 0.009461f
C5500 commonsourceibias.n712 gnd 0.012901f
C5501 commonsourceibias.n713 gnd 0.070526f
C5502 commonsourceibias.n714 gnd 0.012989f
C5503 commonsourceibias.t110 gnd 0.176757f
C5504 commonsourceibias.n715 gnd 0.070526f
C5505 commonsourceibias.n716 gnd 0.011572f
C5506 commonsourceibias.n717 gnd 0.009461f
C5507 commonsourceibias.n718 gnd 0.009461f
C5508 commonsourceibias.n719 gnd 0.009461f
C5509 commonsourceibias.n720 gnd 0.011256f
C5510 commonsourceibias.n721 gnd 0.013054f
C5511 commonsourceibias.n722 gnd 0.070526f
C5512 commonsourceibias.n723 gnd 0.012975f
C5513 commonsourceibias.n724 gnd 0.009461f
C5514 commonsourceibias.n725 gnd 0.009461f
C5515 commonsourceibias.n726 gnd 0.009461f
C5516 commonsourceibias.n727 gnd 0.012816f
C5517 commonsourceibias.n728 gnd 0.070526f
C5518 commonsourceibias.n729 gnd 0.0129f
C5519 commonsourceibias.t136 gnd 0.176757f
C5520 commonsourceibias.n730 gnd 0.070526f
C5521 commonsourceibias.n731 gnd 0.011661f
C5522 commonsourceibias.n732 gnd 0.009461f
C5523 commonsourceibias.n733 gnd 0.009461f
C5524 commonsourceibias.n734 gnd 0.009461f
C5525 commonsourceibias.n735 gnd 0.010754f
C5526 commonsourceibias.n736 gnd 0.013093f
C5527 commonsourceibias.n737 gnd 0.070526f
C5528 commonsourceibias.n738 gnd 0.013037f
C5529 commonsourceibias.n739 gnd 0.009461f
C5530 commonsourceibias.n740 gnd 0.009461f
C5531 commonsourceibias.n741 gnd 0.009461f
C5532 commonsourceibias.n742 gnd 0.012717f
C5533 commonsourceibias.n743 gnd 0.070526f
C5534 commonsourceibias.n744 gnd 0.012748f
C5535 commonsourceibias.t82 gnd 0.191163f
C5536 commonsourceibias.n745 gnd 0.085044f
C5537 commonsourceibias.n746 gnd 0.030348f
C5538 commonsourceibias.n747 gnd 0.199656f
C5539 commonsourceibias.n748 gnd 5.01419f
.ends

