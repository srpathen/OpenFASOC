* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t13 plus.t0 drain_left.t6 a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X1 source.t5 minus.t0 drain_right.t7 a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X2 drain_left.t4 plus.t1 source.t12 a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X3 drain_left.t3 plus.t2 source.t11 a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=1
X4 a_n2046_n2688# a_n2046_n2688# a_n2046_n2688# a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=1
X5 a_n2046_n2688# a_n2046_n2688# a_n2046_n2688# a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=1
X6 source.t10 plus.t3 drain_left.t2 a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=1
X7 source.t9 plus.t4 drain_left.t1 a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X8 drain_right.t6 minus.t1 source.t0 a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=1
X9 a_n2046_n2688# a_n2046_n2688# a_n2046_n2688# a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=1
X10 drain_left.t7 plus.t5 source.t8 a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=1
X11 drain_right.t5 minus.t2 source.t14 a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X12 drain_right.t4 minus.t3 source.t2 a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X13 a_n2046_n2688# a_n2046_n2688# a_n2046_n2688# a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=1
X14 source.t3 minus.t4 drain_right.t3 a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X15 source.t1 minus.t5 drain_right.t2 a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=1
X16 source.t4 minus.t6 drain_right.t1 a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=1
X17 source.t7 plus.t6 drain_left.t5 a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=1
X18 drain_right.t0 minus.t7 source.t15 a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=1
X19 drain_left.t0 plus.t7 source.t6 a_n2046_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
R0 plus.n2 plus.t6 271.445
R1 plus.n15 plus.t5 271.445
R2 plus.n11 plus.t2 256.183
R3 plus.n24 plus.t3 256.183
R4 plus.n9 plus.t0 216.9
R5 plus.n3 plus.t1 216.9
R6 plus.n22 plus.t7 216.9
R7 plus.n16 plus.t4 216.9
R8 plus.n5 plus.n4 161.3
R9 plus.n6 plus.n1 161.3
R10 plus.n8 plus.n7 161.3
R11 plus.n10 plus.n0 161.3
R12 plus.n18 plus.n17 161.3
R13 plus.n19 plus.n14 161.3
R14 plus.n21 plus.n20 161.3
R15 plus.n23 plus.n13 161.3
R16 plus.n12 plus.n11 80.6037
R17 plus.n25 plus.n24 80.6037
R18 plus.n11 plus.n10 56.3158
R19 plus.n24 plus.n23 56.3158
R20 plus.n3 plus.n2 46.9082
R21 plus.n16 plus.n15 46.9082
R22 plus.n5 plus.n2 43.8991
R23 plus.n18 plus.n15 43.8991
R24 plus.n8 plus.n1 40.577
R25 plus.n4 plus.n1 40.577
R26 plus.n21 plus.n14 40.577
R27 plus.n17 plus.n14 40.577
R28 plus plus.n25 29.9957
R29 plus.n10 plus.n9 16.477
R30 plus.n23 plus.n22 16.477
R31 plus plus.n12 11.3873
R32 plus.n9 plus.n8 8.11581
R33 plus.n4 plus.n3 8.11581
R34 plus.n22 plus.n21 8.11581
R35 plus.n17 plus.n16 8.11581
R36 plus.n12 plus.n0 0.285035
R37 plus.n25 plus.n13 0.285035
R38 plus.n6 plus.n5 0.189894
R39 plus.n7 plus.n6 0.189894
R40 plus.n7 plus.n0 0.189894
R41 plus.n20 plus.n13 0.189894
R42 plus.n20 plus.n19 0.189894
R43 plus.n19 plus.n18 0.189894
R44 drain_left.n5 drain_left.n3 66.6841
R45 drain_left.n2 drain_left.n1 66.0553
R46 drain_left.n2 drain_left.n0 66.0553
R47 drain_left.n5 drain_left.n4 65.5374
R48 drain_left drain_left.n2 29.1073
R49 drain_left drain_left.n5 6.79977
R50 drain_left.n1 drain_left.t1 2.2005
R51 drain_left.n1 drain_left.t7 2.2005
R52 drain_left.n0 drain_left.t2 2.2005
R53 drain_left.n0 drain_left.t0 2.2005
R54 drain_left.n4 drain_left.t6 2.2005
R55 drain_left.n4 drain_left.t3 2.2005
R56 drain_left.n3 drain_left.t5 2.2005
R57 drain_left.n3 drain_left.t4 2.2005
R58 source.n3 source.t7 51.0588
R59 source.n4 source.t0 51.0588
R60 source.n7 source.t4 51.0588
R61 source.n15 source.t15 51.0586
R62 source.n12 source.t1 51.0586
R63 source.n11 source.t8 51.0586
R64 source.n8 source.t10 51.0586
R65 source.n0 source.t11 51.0586
R66 source.n2 source.n1 48.8588
R67 source.n6 source.n5 48.8588
R68 source.n14 source.n13 48.8586
R69 source.n10 source.n9 48.8586
R70 source.n8 source.n7 20.1616
R71 source.n16 source.n0 14.3253
R72 source.n16 source.n15 5.83671
R73 source.n13 source.t2 2.2005
R74 source.n13 source.t5 2.2005
R75 source.n9 source.t6 2.2005
R76 source.n9 source.t9 2.2005
R77 source.n1 source.t12 2.2005
R78 source.n1 source.t13 2.2005
R79 source.n5 source.t14 2.2005
R80 source.n5 source.t3 2.2005
R81 source.n7 source.n6 1.14705
R82 source.n6 source.n4 1.14705
R83 source.n3 source.n2 1.14705
R84 source.n2 source.n0 1.14705
R85 source.n10 source.n8 1.14705
R86 source.n11 source.n10 1.14705
R87 source.n14 source.n12 1.14705
R88 source.n15 source.n14 1.14705
R89 source.n4 source.n3 0.470328
R90 source.n12 source.n11 0.470328
R91 source source.n16 0.188
R92 minus.n2 minus.t1 271.445
R93 minus.n15 minus.t5 271.445
R94 minus.n11 minus.t6 256.183
R95 minus.n24 minus.t7 256.183
R96 minus.n3 minus.t4 216.9
R97 minus.n9 minus.t2 216.9
R98 minus.n16 minus.t3 216.9
R99 minus.n22 minus.t0 216.9
R100 minus.n10 minus.n0 161.3
R101 minus.n8 minus.n7 161.3
R102 minus.n6 minus.n1 161.3
R103 minus.n5 minus.n4 161.3
R104 minus.n23 minus.n13 161.3
R105 minus.n21 minus.n20 161.3
R106 minus.n19 minus.n14 161.3
R107 minus.n18 minus.n17 161.3
R108 minus.n12 minus.n11 80.6037
R109 minus.n25 minus.n24 80.6037
R110 minus.n11 minus.n10 56.3158
R111 minus.n24 minus.n23 56.3158
R112 minus.n3 minus.n2 46.9082
R113 minus.n16 minus.n15 46.9082
R114 minus.n5 minus.n2 43.8991
R115 minus.n18 minus.n15 43.8991
R116 minus.n4 minus.n1 40.577
R117 minus.n8 minus.n1 40.577
R118 minus.n17 minus.n14 40.577
R119 minus.n21 minus.n14 40.577
R120 minus.n26 minus.n12 34.9782
R121 minus.n10 minus.n9 16.477
R122 minus.n23 minus.n22 16.477
R123 minus.n4 minus.n3 8.11581
R124 minus.n9 minus.n8 8.11581
R125 minus.n17 minus.n16 8.11581
R126 minus.n22 minus.n21 8.11581
R127 minus.n26 minus.n25 6.87973
R128 minus.n12 minus.n0 0.285035
R129 minus.n25 minus.n13 0.285035
R130 minus.n7 minus.n0 0.189894
R131 minus.n7 minus.n6 0.189894
R132 minus.n6 minus.n5 0.189894
R133 minus.n19 minus.n18 0.189894
R134 minus.n20 minus.n19 0.189894
R135 minus.n20 minus.n13 0.189894
R136 minus minus.n26 0.188
R137 drain_right.n5 drain_right.n3 66.684
R138 drain_right.n2 drain_right.n1 66.0553
R139 drain_right.n2 drain_right.n0 66.0553
R140 drain_right.n5 drain_right.n4 65.5376
R141 drain_right drain_right.n2 28.554
R142 drain_right drain_right.n5 6.79977
R143 drain_right.n1 drain_right.t7 2.2005
R144 drain_right.n1 drain_right.t0 2.2005
R145 drain_right.n0 drain_right.t2 2.2005
R146 drain_right.n0 drain_right.t4 2.2005
R147 drain_right.n3 drain_right.t3 2.2005
R148 drain_right.n3 drain_right.t6 2.2005
R149 drain_right.n4 drain_right.t1 2.2005
R150 drain_right.n4 drain_right.t5 2.2005
C0 minus plus 5.12721f
C1 minus source 4.99285f
C2 minus drain_left 0.172134f
C3 minus drain_right 4.99164f
C4 plus source 5.00689f
C5 plus drain_left 5.19171f
C6 source drain_left 7.90708f
C7 drain_right plus 0.355422f
C8 drain_right source 7.91064f
C9 drain_right drain_left 0.975109f
C10 drain_right a_n2046_n2688# 5.33224f
C11 drain_left a_n2046_n2688# 5.62594f
C12 source a_n2046_n2688# 7.508057f
C13 minus a_n2046_n2688# 7.729917f
C14 plus a_n2046_n2688# 9.13055f
C15 drain_right.t2 a_n2046_n2688# 0.181755f
C16 drain_right.t4 a_n2046_n2688# 0.181755f
C17 drain_right.n0 a_n2046_n2688# 1.59252f
C18 drain_right.t7 a_n2046_n2688# 0.181755f
C19 drain_right.t0 a_n2046_n2688# 0.181755f
C20 drain_right.n1 a_n2046_n2688# 1.59252f
C21 drain_right.n2 a_n2046_n2688# 1.82074f
C22 drain_right.t3 a_n2046_n2688# 0.181755f
C23 drain_right.t6 a_n2046_n2688# 0.181755f
C24 drain_right.n3 a_n2046_n2688# 1.59669f
C25 drain_right.t1 a_n2046_n2688# 0.181755f
C26 drain_right.t5 a_n2046_n2688# 0.181755f
C27 drain_right.n4 a_n2046_n2688# 1.58975f
C28 drain_right.n5 a_n2046_n2688# 1.02557f
C29 minus.n0 a_n2046_n2688# 0.051342f
C30 minus.t2 a_n2046_n2688# 0.93451f
C31 minus.n1 a_n2046_n2688# 0.031076f
C32 minus.t1 a_n2046_n2688# 1.01662f
C33 minus.n2 a_n2046_n2688# 0.414053f
C34 minus.t4 a_n2046_n2688# 0.93451f
C35 minus.n3 a_n2046_n2688# 0.392946f
C36 minus.n4 a_n2046_n2688# 0.052468f
C37 minus.n5 a_n2046_n2688# 0.164715f
C38 minus.n6 a_n2046_n2688# 0.038476f
C39 minus.n7 a_n2046_n2688# 0.038476f
C40 minus.n8 a_n2046_n2688# 0.052468f
C41 minus.n9 a_n2046_n2688# 0.358708f
C42 minus.n10 a_n2046_n2688# 0.052776f
C43 minus.t6 a_n2046_n2688# 0.993097f
C44 minus.n11 a_n2046_n2688# 0.41823f
C45 minus.n12 a_n2046_n2688# 1.31385f
C46 minus.n13 a_n2046_n2688# 0.051342f
C47 minus.t0 a_n2046_n2688# 0.93451f
C48 minus.n14 a_n2046_n2688# 0.031076f
C49 minus.t5 a_n2046_n2688# 1.01662f
C50 minus.n15 a_n2046_n2688# 0.414053f
C51 minus.t3 a_n2046_n2688# 0.93451f
C52 minus.n16 a_n2046_n2688# 0.392946f
C53 minus.n17 a_n2046_n2688# 0.052468f
C54 minus.n18 a_n2046_n2688# 0.164715f
C55 minus.n19 a_n2046_n2688# 0.038476f
C56 minus.n20 a_n2046_n2688# 0.038476f
C57 minus.n21 a_n2046_n2688# 0.052468f
C58 minus.n22 a_n2046_n2688# 0.358708f
C59 minus.n23 a_n2046_n2688# 0.052776f
C60 minus.t7 a_n2046_n2688# 0.993097f
C61 minus.n24 a_n2046_n2688# 0.41823f
C62 minus.n25 a_n2046_n2688# 0.298789f
C63 minus.n26 a_n2046_n2688# 1.57315f
C64 source.t11 a_n2046_n2688# 1.51726f
C65 source.n0 a_n2046_n2688# 0.937448f
C66 source.t12 a_n2046_n2688# 0.142286f
C67 source.t13 a_n2046_n2688# 0.142286f
C68 source.n1 a_n2046_n2688# 1.19112f
C69 source.n2 a_n2046_n2688# 0.334285f
C70 source.t7 a_n2046_n2688# 1.51726f
C71 source.n3 a_n2046_n2688# 0.352573f
C72 source.t0 a_n2046_n2688# 1.51726f
C73 source.n4 a_n2046_n2688# 0.352573f
C74 source.t14 a_n2046_n2688# 0.142286f
C75 source.t3 a_n2046_n2688# 0.142286f
C76 source.n5 a_n2046_n2688# 1.19112f
C77 source.n6 a_n2046_n2688# 0.334285f
C78 source.t4 a_n2046_n2688# 1.51726f
C79 source.n7 a_n2046_n2688# 1.24095f
C80 source.t10 a_n2046_n2688# 1.51726f
C81 source.n8 a_n2046_n2688# 1.24096f
C82 source.t6 a_n2046_n2688# 0.142286f
C83 source.t9 a_n2046_n2688# 0.142286f
C84 source.n9 a_n2046_n2688# 1.19112f
C85 source.n10 a_n2046_n2688# 0.334288f
C86 source.t8 a_n2046_n2688# 1.51726f
C87 source.n11 a_n2046_n2688# 0.352576f
C88 source.t1 a_n2046_n2688# 1.51726f
C89 source.n12 a_n2046_n2688# 0.352576f
C90 source.t2 a_n2046_n2688# 0.142286f
C91 source.t5 a_n2046_n2688# 0.142286f
C92 source.n13 a_n2046_n2688# 1.19112f
C93 source.n14 a_n2046_n2688# 0.334288f
C94 source.t15 a_n2046_n2688# 1.51726f
C95 source.n15 a_n2046_n2688# 0.496002f
C96 source.n16 a_n2046_n2688# 1.06269f
C97 drain_left.t2 a_n2046_n2688# 0.183153f
C98 drain_left.t0 a_n2046_n2688# 0.183153f
C99 drain_left.n0 a_n2046_n2688# 1.60477f
C100 drain_left.t1 a_n2046_n2688# 0.183153f
C101 drain_left.t7 a_n2046_n2688# 0.183153f
C102 drain_left.n1 a_n2046_n2688# 1.60477f
C103 drain_left.n2 a_n2046_n2688# 1.88761f
C104 drain_left.t5 a_n2046_n2688# 0.183153f
C105 drain_left.t4 a_n2046_n2688# 0.183153f
C106 drain_left.n3 a_n2046_n2688# 1.60898f
C107 drain_left.t6 a_n2046_n2688# 0.183153f
C108 drain_left.t3 a_n2046_n2688# 0.183153f
C109 drain_left.n4 a_n2046_n2688# 1.60197f
C110 drain_left.n5 a_n2046_n2688# 1.03346f
C111 plus.n0 a_n2046_n2688# 0.052291f
C112 plus.t2 a_n2046_n2688# 1.01146f
C113 plus.t0 a_n2046_n2688# 0.951792f
C114 plus.n1 a_n2046_n2688# 0.03165f
C115 plus.t6 a_n2046_n2688# 1.03543f
C116 plus.n2 a_n2046_n2688# 0.42171f
C117 plus.t1 a_n2046_n2688# 0.951792f
C118 plus.n3 a_n2046_n2688# 0.400213f
C119 plus.n4 a_n2046_n2688# 0.053439f
C120 plus.n5 a_n2046_n2688# 0.167761f
C121 plus.n6 a_n2046_n2688# 0.039188f
C122 plus.n7 a_n2046_n2688# 0.039188f
C123 plus.n8 a_n2046_n2688# 0.053439f
C124 plus.n9 a_n2046_n2688# 0.365342f
C125 plus.n10 a_n2046_n2688# 0.053752f
C126 plus.n11 a_n2046_n2688# 0.425964f
C127 plus.n12 a_n2046_n2688# 0.434412f
C128 plus.n13 a_n2046_n2688# 0.052291f
C129 plus.t3 a_n2046_n2688# 1.01146f
C130 plus.t7 a_n2046_n2688# 0.951792f
C131 plus.n14 a_n2046_n2688# 0.03165f
C132 plus.t5 a_n2046_n2688# 1.03543f
C133 plus.n15 a_n2046_n2688# 0.42171f
C134 plus.t4 a_n2046_n2688# 0.951792f
C135 plus.n16 a_n2046_n2688# 0.400213f
C136 plus.n17 a_n2046_n2688# 0.053439f
C137 plus.n18 a_n2046_n2688# 0.167761f
C138 plus.n19 a_n2046_n2688# 0.039188f
C139 plus.n20 a_n2046_n2688# 0.039188f
C140 plus.n21 a_n2046_n2688# 0.053439f
C141 plus.n22 a_n2046_n2688# 0.365342f
C142 plus.n23 a_n2046_n2688# 0.053752f
C143 plus.n24 a_n2046_n2688# 0.425964f
C144 plus.n25 a_n2046_n2688# 1.17407f
.ends

