* NGSPICE file created from opamp263.ext - technology: sky130A

.subckt opamp263 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 gnd.t337 commonsourceibias.t80 CSoutput.t84 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X1 CSoutput.t163 a_n6972_8799.t28 vdd.t237 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X2 commonsourceibias.t5 commonsourceibias.t4 gnd.t336 gnd.t300 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X3 a_n1808_13878.t7 a_n1986_13878.t40 vdd.t95 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 a_n1808_13878.t19 a_n1986_13878.t25 a_n1986_13878.t26 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X5 vdd.t236 a_n6972_8799.t29 CSoutput.t175 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X6 CSoutput.t160 a_n6972_8799.t30 vdd.t235 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X7 vdd.t75 vdd.t73 vdd.t74 vdd.t9 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X8 outputibias.t7 outputibias.t6 gnd.t143 gnd.t142 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X9 gnd.t141 gnd.t139 gnd.t140 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X10 a_n6972_8799.t6 plus.t5 a_n2903_n3924.t30 gnd.t144 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X11 gnd.t335 commonsourceibias.t81 CSoutput.t83 gnd.t294 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X12 CSoutput.t174 a_n6972_8799.t31 vdd.t234 vdd.t120 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X13 CSoutput.t176 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X14 gnd.t334 commonsourceibias.t82 CSoutput.t82 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X15 gnd.t333 commonsourceibias.t2 commonsourceibias.t3 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X16 minus.t4 gnd.t136 gnd.t138 gnd.t137 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X17 gnd.t332 commonsourceibias.t83 CSoutput.t81 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X18 a_n1986_8322.t21 a_n1986_13878.t41 a_n6972_8799.t2 vdd.t99 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X19 gnd.t331 commonsourceibias.t84 CSoutput.t80 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 output.t15 CSoutput.t177 vdd.t80 gnd.t25 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X21 CSoutput.t15 a_n6972_8799.t32 vdd.t233 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X22 outputibias.t5 outputibias.t4 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X23 gnd.t330 commonsourceibias.t85 CSoutput.t79 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X24 vdd.t232 a_n6972_8799.t33 CSoutput.t39 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X25 a_n1986_13878.t32 minus.t5 a_n2903_n3924.t9 gnd.t147 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X26 gnd.t329 commonsourceibias.t26 commonsourceibias.t27 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X27 a_n6972_8799.t0 plus.t6 a_n2903_n3924.t29 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X28 a_n1986_13878.t3 minus.t6 a_n2903_n3924.t3 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X29 vdd.t231 a_n6972_8799.t34 CSoutput.t24 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X30 CSoutput.t161 a_n6972_8799.t35 vdd.t230 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X31 vdd.t229 a_n6972_8799.t36 CSoutput.t32 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X32 a_n6972_8799.t3 a_n1986_13878.t42 a_n1986_8322.t20 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X33 CSoutput.t33 a_n6972_8799.t37 vdd.t228 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X34 CSoutput.t94 commonsourceibias.t86 gnd.t328 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 gnd.t327 commonsourceibias.t24 commonsourceibias.t25 gnd.t290 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X36 CSoutput.t93 commonsourceibias.t87 gnd.t326 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 CSoutput.t6 a_n6972_8799.t38 vdd.t227 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X38 vdd.t77 CSoutput.t178 output.t14 gnd.t24 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X39 a_n2903_n3924.t28 plus.t7 a_n6972_8799.t13 gnd.t28 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X40 vdd.t72 vdd.t70 vdd.t71 vdd.t5 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X41 CSoutput.t91 commonsourceibias.t88 gnd.t324 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X42 CSoutput.t92 commonsourceibias.t89 gnd.t325 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 a_n2903_n3924.t8 diffpairibias.t16 gnd.t146 gnd.t145 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X44 CSoutput.t49 a_n6972_8799.t39 vdd.t226 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X45 a_n2903_n3924.t4 minus.t7 a_n1986_13878.t4 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X46 vdd.t69 vdd.t67 vdd.t68 vdd.t9 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X47 CSoutput.t90 commonsourceibias.t90 gnd.t323 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X48 CSoutput.t60 a_n6972_8799.t40 vdd.t225 vdd.t120 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X49 gnd.t322 commonsourceibias.t22 commonsourceibias.t23 gnd.t250 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X50 outputibias.t3 outputibias.t2 gnd.t173 gnd.t172 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X51 output.t13 CSoutput.t179 vdd.t76 gnd.t23 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X52 vdd.t224 a_n6972_8799.t41 CSoutput.t167 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X53 a_n1808_13878.t18 a_n1986_13878.t23 a_n1986_13878.t24 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X54 CSoutput.t98 commonsourceibias.t91 gnd.t306 gnd.t300 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X55 CSoutput.t20 a_n6972_8799.t42 vdd.t223 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X56 commonsourceibias.t21 commonsourceibias.t20 gnd.t321 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X57 a_n1986_13878.t8 a_n1986_13878.t7 a_n1808_13878.t17 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X58 CSoutput.t180 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X59 gnd.t135 gnd.t133 plus.t4 gnd.t134 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X60 CSoutput.t10 a_n6972_8799.t43 vdd.t222 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X61 vdd.t66 vdd.t64 vdd.t65 vdd.t40 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X62 a_n2903_n3924.t27 plus.t8 a_n6972_8799.t9 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X63 vdd.t221 a_n6972_8799.t44 CSoutput.t76 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X64 diffpairibias.t15 diffpairibias.t14 gnd.t33 gnd.t32 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X65 gnd.t132 gnd.t130 gnd.t131 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X66 CSoutput.t71 a_n6972_8799.t45 vdd.t220 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X67 vdd.t219 a_n6972_8799.t46 CSoutput.t165 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X68 vdd.t218 a_n6972_8799.t47 CSoutput.t62 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X69 gnd.t320 commonsourceibias.t92 CSoutput.t89 gnd.t294 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X70 vdd.t216 a_n6972_8799.t48 CSoutput.t64 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X71 diffpairibias.t13 diffpairibias.t12 gnd.t159 gnd.t158 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X72 gnd.t319 commonsourceibias.t93 CSoutput.t88 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X73 CSoutput.t18 a_n6972_8799.t49 vdd.t215 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X74 CSoutput.t4 a_n6972_8799.t50 vdd.t214 vdd.t135 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X75 output.t12 CSoutput.t181 vdd.t83 gnd.t22 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X76 commonsourceibias.t19 commonsourceibias.t18 gnd.t318 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X77 gnd.t317 commonsourceibias.t94 CSoutput.t87 gnd.t290 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X78 vdd.t213 a_n6972_8799.t51 CSoutput.t38 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X79 CSoutput.t51 a_n6972_8799.t52 vdd.t212 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X80 CSoutput.t27 a_n6972_8799.t53 vdd.t211 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 commonsourceibias.t17 commonsourceibias.t16 gnd.t316 gnd.t241 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X82 gnd.t315 commonsourceibias.t95 CSoutput.t103 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X83 CSoutput.t22 a_n6972_8799.t54 vdd.t210 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X84 a_n2903_n3924.t2 minus.t8 a_n1986_13878.t2 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X85 output.t11 CSoutput.t182 vdd.t82 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X86 a_n2903_n3924.t26 plus.t9 a_n6972_8799.t15 gnd.t176 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X87 vdd.t209 a_n6972_8799.t55 CSoutput.t31 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X88 commonsourceibias.t37 commonsourceibias.t36 gnd.t314 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 gnd.t313 commonsourceibias.t96 CSoutput.t102 gnd.t286 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 CSoutput.t97 commonsourceibias.t97 gnd.t305 gnd.t282 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 gnd.t312 commonsourceibias.t34 commonsourceibias.t35 gnd.t286 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X92 a_n2903_n3924.t13 diffpairibias.t17 gnd.t168 gnd.t167 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X93 CSoutput.t183 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X94 a_n1986_13878.t14 a_n1986_13878.t13 a_n1808_13878.t16 vdd.t99 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X95 vdd.t208 a_n6972_8799.t56 CSoutput.t41 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X96 a_n2903_n3924.t25 plus.t10 a_n6972_8799.t4 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X97 a_n6972_8799.t27 a_n1986_13878.t43 a_n1986_8322.t19 vdd.t93 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X98 vdd.t207 a_n6972_8799.t57 CSoutput.t40 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X99 a_n1986_13878.t10 a_n1986_13878.t9 a_n1808_13878.t15 vdd.t104 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X100 gnd.t311 commonsourceibias.t32 commonsourceibias.t33 gnd.t274 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X101 vdd.t206 a_n6972_8799.t58 CSoutput.t63 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X102 commonsourceibias.t31 commonsourceibias.t30 gnd.t310 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X103 CSoutput.t101 commonsourceibias.t98 gnd.t309 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X104 vdd.t205 a_n6972_8799.t59 CSoutput.t17 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X105 CSoutput.t3 a_n6972_8799.t60 vdd.t204 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X106 CSoutput.t100 commonsourceibias.t99 gnd.t308 gnd.t269 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X107 vdd.t90 CSoutput.t184 output.t10 gnd.t20 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X108 vdd.t63 vdd.t61 vdd.t62 vdd.t48 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X109 vdd.t203 a_n6972_8799.t61 CSoutput.t57 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X110 CSoutput.t99 commonsourceibias.t100 gnd.t307 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X111 CSoutput.t35 a_n6972_8799.t62 vdd.t202 vdd.t135 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X112 vdd.t60 vdd.t57 vdd.t59 vdd.t58 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X113 gnd.t304 commonsourceibias.t101 CSoutput.t96 gnd.t274 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X114 commonsourceibias.t29 commonsourceibias.t28 gnd.t303 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X115 CSoutput.t95 commonsourceibias.t102 gnd.t302 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X116 CSoutput.t110 commonsourceibias.t103 gnd.t301 gnd.t300 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X117 vdd.t56 vdd.t54 vdd.t55 vdd.t1 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X118 vdd.t53 vdd.t51 vdd.t52 vdd.t44 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X119 vdd.t263 a_n1986_13878.t44 a_n1986_8322.t9 vdd.t262 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X120 gnd.t129 gnd.t127 minus.t3 gnd.t128 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X121 a_n1986_8322.t8 a_n1986_13878.t45 vdd.t259 vdd.t258 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X122 a_n2903_n3924.t12 diffpairibias.t18 gnd.t166 gnd.t165 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X123 CSoutput.t45 a_n6972_8799.t63 vdd.t201 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X124 gnd.t299 commonsourceibias.t104 CSoutput.t109 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X125 vdd.t199 a_n6972_8799.t64 CSoutput.t29 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X126 commonsourceibias.t47 commonsourceibias.t46 gnd.t298 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X127 gnd.t126 gnd.t124 gnd.t125 gnd.t68 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X128 commonsourceibias.t45 commonsourceibias.t44 gnd.t297 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X129 vdd.t261 a_n1986_13878.t46 a_n1808_13878.t6 vdd.t260 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X130 vdd.t50 vdd.t47 vdd.t49 vdd.t48 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X131 gnd.t296 commonsourceibias.t42 commonsourceibias.t43 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X132 gnd.t285 commonsourceibias.t105 CSoutput.t120 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X133 vdd.t197 a_n6972_8799.t65 CSoutput.t8 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X134 vdd.t46 vdd.t43 vdd.t45 vdd.t44 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X135 gnd.t295 commonsourceibias.t40 commonsourceibias.t41 gnd.t294 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X136 outputibias.t1 outputibias.t0 gnd.t175 gnd.t174 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X137 a_n6972_8799.t17 plus.t11 a_n2903_n3924.t24 gnd.t177 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X138 vdd.t42 vdd.t39 vdd.t41 vdd.t40 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X139 a_n1986_8322.t7 a_n1986_13878.t47 vdd.t257 vdd.t256 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X140 commonsourceibias.t39 commonsourceibias.t38 gnd.t293 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X141 gnd.t292 commonsourceibias.t106 CSoutput.t108 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X142 gnd.t291 commonsourceibias.t107 CSoutput.t107 gnd.t290 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X143 a_n6972_8799.t26 a_n1986_13878.t48 a_n1986_8322.t18 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X144 gnd.t289 commonsourceibias.t108 CSoutput.t106 gnd.t246 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X145 a_n6972_8799.t7 plus.t12 a_n2903_n3924.t23 gnd.t150 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X146 diffpairibias.t11 diffpairibias.t10 gnd.t149 gnd.t148 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X147 a_n1986_13878.t28 a_n1986_13878.t27 a_n1808_13878.t14 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X148 vdd.t195 a_n6972_8799.t66 CSoutput.t65 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X149 a_n6972_8799.t25 a_n1986_13878.t49 a_n1986_8322.t17 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X150 CSoutput.t74 a_n6972_8799.t67 vdd.t194 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X151 gnd.t288 commonsourceibias.t109 CSoutput.t105 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X152 output.t19 outputibias.t8 gnd.t31 gnd.t30 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X153 a_n1808_13878.t13 a_n1986_13878.t15 a_n1986_13878.t16 vdd.t93 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X154 gnd.t123 gnd.t121 gnd.t122 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X155 gnd.t287 commonsourceibias.t110 CSoutput.t104 gnd.t286 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X156 CSoutput.t119 commonsourceibias.t111 gnd.t284 gnd.t282 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X157 commonsourceibias.t49 commonsourceibias.t48 gnd.t283 gnd.t282 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X158 CSoutput.t69 a_n6972_8799.t68 vdd.t193 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X159 gnd.t281 commonsourceibias.t112 CSoutput.t118 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X160 vdd.t255 a_n1986_13878.t50 a_n1986_8322.t6 vdd.t254 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X161 CSoutput.t117 commonsourceibias.t113 gnd.t280 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X162 vdd.t192 a_n6972_8799.t69 CSoutput.t168 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X163 a_n1986_13878.t31 minus.t9 a_n2903_n3924.t7 gnd.t144 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X164 a_n2903_n3924.t22 plus.t13 a_n6972_8799.t12 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X165 CSoutput.t56 a_n6972_8799.t70 vdd.t191 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X166 plus.t3 gnd.t118 gnd.t120 gnd.t119 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X167 vdd.t190 a_n6972_8799.t71 CSoutput.t19 vdd.t112 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X168 CSoutput.t116 commonsourceibias.t114 gnd.t279 gnd.t269 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X169 a_n2903_n3924.t38 diffpairibias.t19 gnd.t347 gnd.t346 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X170 gnd.t117 gnd.t115 minus.t2 gnd.t116 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X171 gnd.t114 gnd.t111 gnd.t113 gnd.t112 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X172 a_n2903_n3924.t35 diffpairibias.t20 gnd.t339 gnd.t338 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X173 vdd.t81 CSoutput.t185 output.t9 gnd.t19 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X174 a_n6972_8799.t1 plus.t14 a_n2903_n3924.t21 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X175 CSoutput.t115 commonsourceibias.t115 gnd.t278 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X176 CSoutput.t114 commonsourceibias.t116 gnd.t277 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X177 vdd.t189 a_n6972_8799.t72 CSoutput.t70 vdd.t145 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X178 gnd.t275 commonsourceibias.t117 CSoutput.t113 gnd.t274 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X179 gnd.t273 commonsourceibias.t118 CSoutput.t112 gnd.t250 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X180 CSoutput.t111 commonsourceibias.t119 gnd.t272 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X181 commonsourceibias.t55 commonsourceibias.t54 gnd.t270 gnd.t269 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X182 CSoutput.t129 commonsourceibias.t120 gnd.t268 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X183 gnd.t110 gnd.t108 gnd.t109 gnd.t43 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X184 a_n6972_8799.t14 plus.t15 a_n2903_n3924.t20 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X185 gnd.t107 gnd.t104 gnd.t106 gnd.t105 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X186 gnd.t267 commonsourceibias.t121 CSoutput.t128 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X187 CSoutput.t73 a_n6972_8799.t73 vdd.t188 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X188 CSoutput.t47 a_n6972_8799.t74 vdd.t186 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X189 gnd.t103 gnd.t101 gnd.t102 gnd.t72 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X190 CSoutput.t127 commonsourceibias.t122 gnd.t266 gnd.t241 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X191 diffpairibias.t9 diffpairibias.t8 gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X192 a_n1808_13878.t5 a_n1986_13878.t51 vdd.t249 vdd.t248 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X193 a_n1986_13878.t0 minus.t10 a_n2903_n3924.t0 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X194 vdd.t251 a_n1986_13878.t52 a_n1808_13878.t4 vdd.t250 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X195 vdd.t38 vdd.t36 vdd.t37 vdd.t20 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X196 CSoutput.t30 a_n6972_8799.t75 vdd.t185 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X197 a_n2903_n3924.t19 plus.t16 a_n6972_8799.t19 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X198 vdd.t183 a_n6972_8799.t76 CSoutput.t46 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X199 gnd.t183 commonsourceibias.t123 CSoutput.t85 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X200 CSoutput.t126 commonsourceibias.t124 gnd.t265 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X201 gnd.t264 commonsourceibias.t52 commonsourceibias.t53 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X202 gnd.t263 commonsourceibias.t125 CSoutput.t125 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X203 gnd.t262 commonsourceibias.t126 CSoutput.t124 gnd.t246 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X204 CSoutput.t171 a_n6972_8799.t77 vdd.t181 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X205 vdd.t179 a_n6972_8799.t78 CSoutput.t162 vdd.t112 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X206 a_n2903_n3924.t31 minus.t11 a_n1986_13878.t35 gnd.t171 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X207 gnd.t261 commonsourceibias.t127 CSoutput.t123 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X208 a_n1986_8322.t16 a_n1986_13878.t53 a_n6972_8799.t22 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X209 vdd.t86 CSoutput.t186 output.t8 gnd.t18 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X210 CSoutput.t2 a_n6972_8799.t79 vdd.t178 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X211 diffpairibias.t7 diffpairibias.t6 gnd.t161 gnd.t160 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X212 CSoutput.t122 commonsourceibias.t128 gnd.t260 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X213 vdd.t177 a_n6972_8799.t80 CSoutput.t42 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X214 CSoutput.t14 a_n6972_8799.t81 vdd.t175 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X215 vdd.t174 a_n6972_8799.t82 CSoutput.t7 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X216 vdd.t253 a_n1986_13878.t54 a_n1986_8322.t5 vdd.t252 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X217 gnd.t259 commonsourceibias.t50 commonsourceibias.t51 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X218 vdd.t172 a_n6972_8799.t83 CSoutput.t170 vdd.t145 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X219 gnd.t100 gnd.t98 gnd.t99 gnd.t72 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X220 CSoutput.t121 commonsourceibias.t129 gnd.t257 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X221 plus.t2 gnd.t95 gnd.t97 gnd.t96 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X222 gnd.t94 gnd.t92 minus.t1 gnd.t93 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X223 gnd.t256 commonsourceibias.t130 CSoutput.t138 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X224 CSoutput.t137 commonsourceibias.t131 gnd.t255 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X225 a_n1808_13878.t3 a_n1986_13878.t55 vdd.t241 vdd.t240 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X226 vdd.t171 a_n6972_8799.t84 CSoutput.t169 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X227 CSoutput.t9 a_n6972_8799.t85 vdd.t170 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X228 CSoutput.t43 a_n6972_8799.t86 vdd.t169 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X229 gnd.t254 commonsourceibias.t60 commonsourceibias.t61 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X230 gnd.t91 gnd.t88 gnd.t90 gnd.t89 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X231 vdd.t35 vdd.t33 vdd.t34 vdd.t20 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X232 a_n2903_n3924.t36 diffpairibias.t21 gnd.t343 gnd.t342 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X233 CSoutput.t136 commonsourceibias.t132 gnd.t253 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X234 vdd.t243 a_n1986_13878.t56 a_n1986_8322.t4 vdd.t242 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X235 a_n1986_8322.t15 a_n1986_13878.t57 a_n6972_8799.t23 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X236 CSoutput.t187 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X237 CSoutput.t21 a_n6972_8799.t87 vdd.t168 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X238 a_n6972_8799.t10 plus.t17 a_n2903_n3924.t18 gnd.t147 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X239 vdd.t166 a_n6972_8799.t88 CSoutput.t36 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X240 vdd.t32 vdd.t30 vdd.t31 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X241 a_n1986_13878.t36 minus.t12 a_n2903_n3924.t32 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X242 CSoutput.t135 commonsourceibias.t133 gnd.t252 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X243 CSoutput.t12 a_n6972_8799.t89 vdd.t165 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X244 a_n2903_n3924.t33 minus.t13 a_n1986_13878.t37 gnd.t176 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X245 gnd.t251 commonsourceibias.t134 CSoutput.t134 gnd.t250 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X246 vdd.t164 a_n6972_8799.t90 CSoutput.t53 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X247 vdd.t163 a_n6972_8799.t91 CSoutput.t172 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X248 gnd.t249 commonsourceibias.t58 commonsourceibias.t59 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X249 gnd.t247 commonsourceibias.t56 commonsourceibias.t57 gnd.t246 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X250 vdd.t78 CSoutput.t188 output.t7 gnd.t17 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X251 CSoutput.t133 commonsourceibias.t135 gnd.t245 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X252 output.t6 CSoutput.t189 vdd.t84 gnd.t16 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X253 CSoutput.t132 commonsourceibias.t136 gnd.t244 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X254 gnd.t243 commonsourceibias.t137 CSoutput.t131 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X255 vdd.t29 vdd.t26 vdd.t28 vdd.t27 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X256 a_n2903_n3924.t34 minus.t14 a_n1986_13878.t38 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X257 gnd.t87 gnd.t85 gnd.t86 gnd.t57 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X258 gnd.t84 gnd.t81 gnd.t83 gnd.t82 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X259 a_n2903_n3924.t6 minus.t15 a_n1986_13878.t6 gnd.t28 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X260 a_n1808_13878.t12 a_n1986_13878.t17 a_n1986_13878.t18 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X261 CSoutput.t66 a_n6972_8799.t92 vdd.t162 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X262 gnd.t80 gnd.t78 gnd.t79 gnd.t57 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X263 CSoutput.t130 commonsourceibias.t138 gnd.t242 gnd.t241 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X264 a_n1986_8322.t14 a_n1986_13878.t58 a_n6972_8799.t24 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X265 diffpairibias.t5 diffpairibias.t4 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X266 CSoutput.t190 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X267 commonsourceibias.t79 commonsourceibias.t78 gnd.t240 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X268 CSoutput.t58 a_n6972_8799.t93 vdd.t161 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X269 vdd.t159 a_n6972_8799.t94 CSoutput.t37 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X270 gnd.t239 commonsourceibias.t139 CSoutput.t157 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X271 CSoutput.t156 commonsourceibias.t140 gnd.t238 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X272 vdd.t158 a_n6972_8799.t95 CSoutput.t75 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 a_n1986_8322.t3 a_n1986_13878.t59 vdd.t245 vdd.t244 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X274 gnd.t237 commonsourceibias.t76 commonsourceibias.t77 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 gnd.t235 commonsourceibias.t141 CSoutput.t155 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X276 CSoutput.t77 a_n6972_8799.t96 vdd.t156 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X277 a_n2903_n3924.t1 minus.t16 a_n1986_13878.t1 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X278 gnd.t77 gnd.t75 gnd.t76 gnd.t43 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X279 output.t18 outputibias.t9 gnd.t157 gnd.t156 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X280 CSoutput.t78 commonsourceibias.t142 gnd.t181 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X281 vdd.t247 a_n1986_13878.t60 a_n1808_13878.t2 vdd.t246 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X282 CSoutput.t23 a_n6972_8799.t97 vdd.t154 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X283 vdd.t25 vdd.t23 vdd.t24 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X284 output.t5 CSoutput.t191 vdd.t88 gnd.t15 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X285 CSoutput.t13 a_n6972_8799.t98 vdd.t152 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X286 gnd.t74 gnd.t71 gnd.t73 gnd.t72 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X287 vdd.t89 CSoutput.t192 output.t4 gnd.t14 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X288 gnd.t234 commonsourceibias.t143 CSoutput.t154 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X289 CSoutput.t153 commonsourceibias.t144 gnd.t233 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X290 CSoutput.t152 commonsourceibias.t145 gnd.t232 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X291 vdd.t151 a_n6972_8799.t99 CSoutput.t52 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X292 gnd.t230 commonsourceibias.t74 commonsourceibias.t75 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X293 vdd.t149 a_n6972_8799.t100 CSoutput.t11 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X294 output.t17 outputibias.t10 gnd.t155 gnd.t154 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X295 gnd.t70 gnd.t67 gnd.t69 gnd.t68 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X296 vdd.t22 vdd.t19 vdd.t21 vdd.t20 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X297 gnd.t66 gnd.t64 plus.t1 gnd.t65 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X298 a_n1986_8322.t13 a_n1986_13878.t61 a_n6972_8799.t20 vdd.t105 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X299 CSoutput.t61 a_n6972_8799.t101 vdd.t148 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X300 vdd.t18 vdd.t16 vdd.t17 vdd.t5 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X301 a_n6972_8799.t21 a_n1986_13878.t62 a_n1986_8322.t12 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X302 vdd.t146 a_n6972_8799.t102 CSoutput.t44 vdd.t145 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X303 a_n1808_13878.t1 a_n1986_13878.t63 vdd.t239 vdd.t238 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X304 output.t16 outputibias.t11 gnd.t170 gnd.t169 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X305 vdd.t85 CSoutput.t193 output.t3 gnd.t13 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X306 vdd.t144 a_n6972_8799.t103 CSoutput.t158 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X307 CSoutput.t0 a_n6972_8799.t104 vdd.t143 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X308 a_n2903_n3924.t17 plus.t18 a_n6972_8799.t8 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X309 a_n1986_13878.t33 minus.t17 a_n2903_n3924.t10 gnd.t150 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X310 CSoutput.t151 commonsourceibias.t146 gnd.t228 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X311 gnd.t63 gnd.t60 gnd.t62 gnd.t61 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X312 vdd.t15 vdd.t12 vdd.t14 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X313 vdd.t11 vdd.t8 vdd.t10 vdd.t9 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X314 output.t2 CSoutput.t194 vdd.t91 gnd.t12 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X315 a_n1808_13878.t11 a_n1986_13878.t29 a_n1986_13878.t30 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X316 CSoutput.t1 a_n6972_8799.t105 vdd.t141 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X317 commonsourceibias.t67 commonsourceibias.t66 gnd.t226 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X318 gnd.t224 commonsourceibias.t147 CSoutput.t144 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X319 vdd.t140 a_n6972_8799.t106 CSoutput.t166 vdd.t122 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X320 gnd.t223 commonsourceibias.t64 commonsourceibias.t65 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X321 CSoutput.t141 commonsourceibias.t148 gnd.t218 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X322 gnd.t222 commonsourceibias.t149 CSoutput.t143 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X323 CSoutput.t54 a_n6972_8799.t107 vdd.t139 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X324 a_n2903_n3924.t5 minus.t18 a_n1986_13878.t5 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X325 a_n2903_n3924.t37 diffpairibias.t22 gnd.t345 gnd.t344 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X326 output.t1 CSoutput.t195 vdd.t87 gnd.t11 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X327 gnd.t220 commonsourceibias.t150 CSoutput.t142 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X328 vdd.t138 a_n6972_8799.t108 CSoutput.t16 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X329 gnd.t59 gnd.t56 gnd.t58 gnd.t57 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X330 gnd.t216 commonsourceibias.t151 CSoutput.t140 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X331 a_n1986_13878.t12 a_n1986_13878.t11 a_n1808_13878.t10 vdd.t105 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X332 commonsourceibias.t63 commonsourceibias.t62 gnd.t214 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X333 a_n6972_8799.t16 a_n1986_13878.t64 a_n1986_8322.t11 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X334 gnd.t55 gnd.t52 gnd.t54 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X335 gnd.t213 commonsourceibias.t152 CSoutput.t139 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X336 vdd.t137 a_n6972_8799.t109 CSoutput.t48 vdd.t122 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X337 CSoutput.t55 a_n6972_8799.t110 vdd.t136 vdd.t135 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X338 vdd.t134 a_n6972_8799.t111 CSoutput.t26 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X339 diffpairibias.t3 diffpairibias.t2 gnd.t164 gnd.t163 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X340 vdd.t133 a_n6972_8799.t112 CSoutput.t50 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X341 vdd.t7 vdd.t4 vdd.t6 vdd.t5 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X342 gnd.t51 gnd.t49 plus.t0 gnd.t50 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X343 minus.t0 gnd.t46 gnd.t48 gnd.t47 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X344 CSoutput.t28 a_n6972_8799.t113 vdd.t131 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X345 a_n1986_13878.t34 minus.t19 a_n2903_n3924.t14 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X346 commonsourceibias.t73 commonsourceibias.t72 gnd.t211 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X347 vdd.t129 a_n6972_8799.t114 CSoutput.t59 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X348 gnd.t209 commonsourceibias.t153 CSoutput.t150 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X349 diffpairibias.t1 diffpairibias.t0 gnd.t341 gnd.t340 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X350 CSoutput.t196 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X351 gnd.t45 gnd.t42 gnd.t44 gnd.t43 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X352 CSoutput.t149 commonsourceibias.t154 gnd.t207 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X353 vdd.t103 a_n1986_13878.t65 a_n1808_13878.t0 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X354 commonsourceibias.t71 commonsourceibias.t70 gnd.t205 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X355 gnd.t41 gnd.t38 gnd.t40 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X356 gnd.t204 commonsourceibias.t155 CSoutput.t148 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X357 CSoutput.t147 commonsourceibias.t156 gnd.t203 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X358 CSoutput.t68 a_n6972_8799.t115 vdd.t127 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X359 CSoutput.t146 commonsourceibias.t157 gnd.t201 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X360 vdd.t125 a_n6972_8799.t116 CSoutput.t25 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X361 commonsourceibias.t69 commonsourceibias.t68 gnd.t199 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X362 vdd.t123 a_n6972_8799.t117 CSoutput.t164 vdd.t122 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X363 CSoutput.t145 commonsourceibias.t158 gnd.t197 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X364 CSoutput.t159 a_n6972_8799.t118 vdd.t121 vdd.t120 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X365 gnd.t195 commonsourceibias.t14 commonsourceibias.t15 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X366 vdd.t79 CSoutput.t197 output.t0 gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X367 a_n6972_8799.t11 plus.t19 a_n2903_n3924.t16 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X368 a_n1986_13878.t39 minus.t20 a_n2903_n3924.t39 gnd.t177 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X369 CSoutput.t86 commonsourceibias.t159 gnd.t193 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X370 CSoutput.t67 a_n6972_8799.t119 vdd.t119 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X371 a_n1986_8322.t10 a_n1986_13878.t66 a_n6972_8799.t5 vdd.t104 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X372 gnd.t191 commonsourceibias.t12 commonsourceibias.t13 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X373 vdd.t117 a_n6972_8799.t120 CSoutput.t34 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X374 CSoutput.t72 a_n6972_8799.t121 vdd.t115 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X375 vdd.t113 a_n6972_8799.t122 CSoutput.t173 vdd.t112 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X376 commonsourceibias.t11 commonsourceibias.t10 gnd.t189 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X377 gnd.t187 commonsourceibias.t8 commonsourceibias.t9 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X378 a_n1986_8322.t2 a_n1986_13878.t67 vdd.t101 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X379 gnd.t37 gnd.t34 gnd.t36 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X380 a_n1808_13878.t9 a_n1986_13878.t19 a_n1986_13878.t20 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X381 vdd.t111 a_n6972_8799.t123 CSoutput.t5 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X382 commonsourceibias.t7 commonsourceibias.t6 gnd.t185 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X383 a_n2903_n3924.t15 plus.t20 a_n6972_8799.t18 gnd.t171 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X384 a_n2903_n3924.t11 diffpairibias.t23 gnd.t153 gnd.t152 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X385 gnd.t179 commonsourceibias.t0 commonsourceibias.t1 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X386 a_n1986_13878.t22 a_n1986_13878.t21 a_n1808_13878.t8 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X387 vdd.t3 vdd.t0 vdd.t2 vdd.t1 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
R0 commonsourceibias.n281 commonsourceibias.t102 222.032
R1 commonsourceibias.n44 commonsourceibias.t20 222.032
R2 commonsourceibias.n166 commonsourceibias.t119 222.032
R3 commonsourceibias.n643 commonsourceibias.t108 222.032
R4 commonsourceibias.n413 commonsourceibias.t56 222.032
R5 commonsourceibias.n529 commonsourceibias.t126 222.032
R6 commonsourceibias.n364 commonsourceibias.t101 207.983
R7 commonsourceibias.n127 commonsourceibias.t32 207.983
R8 commonsourceibias.n249 commonsourceibias.t117 207.983
R9 commonsourceibias.n731 commonsourceibias.t124 207.983
R10 commonsourceibias.n501 commonsourceibias.t6 207.983
R11 commonsourceibias.n616 commonsourceibias.t140 207.983
R12 commonsourceibias.n280 commonsourceibias.t152 168.701
R13 commonsourceibias.n286 commonsourceibias.t157 168.701
R14 commonsourceibias.n292 commonsourceibias.t112 168.701
R15 commonsourceibias.n276 commonsourceibias.t97 168.701
R16 commonsourceibias.n300 commonsourceibias.t85 168.701
R17 commonsourceibias.n306 commonsourceibias.t122 168.701
R18 commonsourceibias.n271 commonsourceibias.t104 168.701
R19 commonsourceibias.n314 commonsourceibias.t91 168.701
R20 commonsourceibias.n320 commonsourceibias.t94 168.701
R21 commonsourceibias.n266 commonsourceibias.t113 168.701
R22 commonsourceibias.n328 commonsourceibias.t96 168.701
R23 commonsourceibias.n334 commonsourceibias.t100 168.701
R24 commonsourceibias.n261 commonsourceibias.t151 168.701
R25 commonsourceibias.n342 commonsourceibias.t129 168.701
R26 commonsourceibias.n348 commonsourceibias.t109 168.701
R27 commonsourceibias.n256 commonsourceibias.t159 168.701
R28 commonsourceibias.n356 commonsourceibias.t81 168.701
R29 commonsourceibias.n362 commonsourceibias.t120 168.701
R30 commonsourceibias.n125 commonsourceibias.t66 168.701
R31 commonsourceibias.n119 commonsourceibias.t40 168.701
R32 commonsourceibias.n19 commonsourceibias.t30 168.701
R33 commonsourceibias.n111 commonsourceibias.t50 168.701
R34 commonsourceibias.n105 commonsourceibias.t36 168.701
R35 commonsourceibias.n24 commonsourceibias.t2 168.701
R36 commonsourceibias.n97 commonsourceibias.t46 168.701
R37 commonsourceibias.n91 commonsourceibias.t34 168.701
R38 commonsourceibias.n29 commonsourceibias.t72 168.701
R39 commonsourceibias.n83 commonsourceibias.t24 168.701
R40 commonsourceibias.n77 commonsourceibias.t4 168.701
R41 commonsourceibias.n34 commonsourceibias.t58 168.701
R42 commonsourceibias.n69 commonsourceibias.t16 168.701
R43 commonsourceibias.n63 commonsourceibias.t74 168.701
R44 commonsourceibias.n39 commonsourceibias.t48 168.701
R45 commonsourceibias.n55 commonsourceibias.t8 168.701
R46 commonsourceibias.n49 commonsourceibias.t70 168.701
R47 commonsourceibias.n43 commonsourceibias.t64 168.701
R48 commonsourceibias.n247 commonsourceibias.t135 168.701
R49 commonsourceibias.n241 commonsourceibias.t92 168.701
R50 commonsourceibias.n5 commonsourceibias.t90 168.701
R51 commonsourceibias.n233 commonsourceibias.t127 168.701
R52 commonsourceibias.n227 commonsourceibias.t145 168.701
R53 commonsourceibias.n10 commonsourceibias.t83 168.701
R54 commonsourceibias.n219 commonsourceibias.t116 168.701
R55 commonsourceibias.n213 commonsourceibias.t110 168.701
R56 commonsourceibias.n150 commonsourceibias.t131 168.701
R57 commonsourceibias.n151 commonsourceibias.t107 168.701
R58 commonsourceibias.n153 commonsourceibias.t103 168.701
R59 commonsourceibias.n155 commonsourceibias.t121 168.701
R60 commonsourceibias.n191 commonsourceibias.t138 168.701
R61 commonsourceibias.n185 commonsourceibias.t95 168.701
R62 commonsourceibias.n161 commonsourceibias.t111 168.701
R63 commonsourceibias.n177 commonsourceibias.t130 168.701
R64 commonsourceibias.n171 commonsourceibias.t87 168.701
R65 commonsourceibias.n165 commonsourceibias.t84 168.701
R66 commonsourceibias.n642 commonsourceibias.t158 168.701
R67 commonsourceibias.n648 commonsourceibias.t150 168.701
R68 commonsourceibias.n654 commonsourceibias.t136 168.701
R69 commonsourceibias.n656 commonsourceibias.t118 168.701
R70 commonsourceibias.n663 commonsourceibias.t99 168.701
R71 commonsourceibias.n669 commonsourceibias.t143 168.701
R72 commonsourceibias.n671 commonsourceibias.t128 168.701
R73 commonsourceibias.n678 commonsourceibias.t106 168.701
R74 commonsourceibias.n684 commonsourceibias.t88 168.701
R75 commonsourceibias.n686 commonsourceibias.t137 168.701
R76 commonsourceibias.n693 commonsourceibias.t115 168.701
R77 commonsourceibias.n699 commonsourceibias.t123 168.701
R78 commonsourceibias.n701 commonsourceibias.t144 168.701
R79 commonsourceibias.n708 commonsourceibias.t147 168.701
R80 commonsourceibias.n714 commonsourceibias.t132 168.701
R81 commonsourceibias.n716 commonsourceibias.t93 168.701
R82 commonsourceibias.n723 commonsourceibias.t154 168.701
R83 commonsourceibias.n729 commonsourceibias.t141 168.701
R84 commonsourceibias.n412 commonsourceibias.t44 168.701
R85 commonsourceibias.n418 commonsourceibias.t42 168.701
R86 commonsourceibias.n424 commonsourceibias.t78 168.701
R87 commonsourceibias.n426 commonsourceibias.t22 168.701
R88 commonsourceibias.n433 commonsourceibias.t54 168.701
R89 commonsourceibias.n439 commonsourceibias.t14 168.701
R90 commonsourceibias.n441 commonsourceibias.t38 168.701
R91 commonsourceibias.n448 commonsourceibias.t76 168.701
R92 commonsourceibias.n454 commonsourceibias.t68 168.701
R93 commonsourceibias.n456 commonsourceibias.t60 168.701
R94 commonsourceibias.n463 commonsourceibias.t10 168.701
R95 commonsourceibias.n469 commonsourceibias.t26 168.701
R96 commonsourceibias.n471 commonsourceibias.t62 168.701
R97 commonsourceibias.n478 commonsourceibias.t12 168.701
R98 commonsourceibias.n484 commonsourceibias.t28 168.701
R99 commonsourceibias.n486 commonsourceibias.t0 168.701
R100 commonsourceibias.n493 commonsourceibias.t18 168.701
R101 commonsourceibias.n499 commonsourceibias.t52 168.701
R102 commonsourceibias.n614 commonsourceibias.t153 168.701
R103 commonsourceibias.n608 commonsourceibias.t86 168.701
R104 commonsourceibias.n601 commonsourceibias.t105 168.701
R105 commonsourceibias.n599 commonsourceibias.t146 168.701
R106 commonsourceibias.n593 commonsourceibias.t80 168.701
R107 commonsourceibias.n586 commonsourceibias.t156 168.701
R108 commonsourceibias.n584 commonsourceibias.t139 168.701
R109 commonsourceibias.n578 commonsourceibias.t133 168.701
R110 commonsourceibias.n571 commonsourceibias.t149 168.701
R111 commonsourceibias.n528 commonsourceibias.t89 168.701
R112 commonsourceibias.n534 commonsourceibias.t82 168.701
R113 commonsourceibias.n540 commonsourceibias.t148 168.701
R114 commonsourceibias.n542 commonsourceibias.t134 168.701
R115 commonsourceibias.n549 commonsourceibias.t114 168.701
R116 commonsourceibias.n555 commonsourceibias.t155 168.701
R117 commonsourceibias.n519 commonsourceibias.t142 168.701
R118 commonsourceibias.n517 commonsourceibias.t125 168.701
R119 commonsourceibias.n515 commonsourceibias.t98 168.701
R120 commonsourceibias.n363 commonsourceibias.n251 161.3
R121 commonsourceibias.n361 commonsourceibias.n360 161.3
R122 commonsourceibias.n359 commonsourceibias.n252 161.3
R123 commonsourceibias.n358 commonsourceibias.n357 161.3
R124 commonsourceibias.n355 commonsourceibias.n253 161.3
R125 commonsourceibias.n354 commonsourceibias.n353 161.3
R126 commonsourceibias.n352 commonsourceibias.n254 161.3
R127 commonsourceibias.n351 commonsourceibias.n350 161.3
R128 commonsourceibias.n349 commonsourceibias.n255 161.3
R129 commonsourceibias.n347 commonsourceibias.n346 161.3
R130 commonsourceibias.n345 commonsourceibias.n257 161.3
R131 commonsourceibias.n344 commonsourceibias.n343 161.3
R132 commonsourceibias.n341 commonsourceibias.n258 161.3
R133 commonsourceibias.n340 commonsourceibias.n339 161.3
R134 commonsourceibias.n338 commonsourceibias.n259 161.3
R135 commonsourceibias.n337 commonsourceibias.n336 161.3
R136 commonsourceibias.n335 commonsourceibias.n260 161.3
R137 commonsourceibias.n333 commonsourceibias.n332 161.3
R138 commonsourceibias.n331 commonsourceibias.n262 161.3
R139 commonsourceibias.n330 commonsourceibias.n329 161.3
R140 commonsourceibias.n327 commonsourceibias.n263 161.3
R141 commonsourceibias.n326 commonsourceibias.n325 161.3
R142 commonsourceibias.n324 commonsourceibias.n264 161.3
R143 commonsourceibias.n323 commonsourceibias.n322 161.3
R144 commonsourceibias.n321 commonsourceibias.n265 161.3
R145 commonsourceibias.n319 commonsourceibias.n318 161.3
R146 commonsourceibias.n317 commonsourceibias.n267 161.3
R147 commonsourceibias.n316 commonsourceibias.n315 161.3
R148 commonsourceibias.n313 commonsourceibias.n268 161.3
R149 commonsourceibias.n312 commonsourceibias.n311 161.3
R150 commonsourceibias.n310 commonsourceibias.n269 161.3
R151 commonsourceibias.n309 commonsourceibias.n308 161.3
R152 commonsourceibias.n307 commonsourceibias.n270 161.3
R153 commonsourceibias.n305 commonsourceibias.n304 161.3
R154 commonsourceibias.n303 commonsourceibias.n272 161.3
R155 commonsourceibias.n302 commonsourceibias.n301 161.3
R156 commonsourceibias.n299 commonsourceibias.n273 161.3
R157 commonsourceibias.n298 commonsourceibias.n297 161.3
R158 commonsourceibias.n296 commonsourceibias.n274 161.3
R159 commonsourceibias.n295 commonsourceibias.n294 161.3
R160 commonsourceibias.n293 commonsourceibias.n275 161.3
R161 commonsourceibias.n291 commonsourceibias.n290 161.3
R162 commonsourceibias.n289 commonsourceibias.n277 161.3
R163 commonsourceibias.n288 commonsourceibias.n287 161.3
R164 commonsourceibias.n285 commonsourceibias.n278 161.3
R165 commonsourceibias.n284 commonsourceibias.n283 161.3
R166 commonsourceibias.n282 commonsourceibias.n279 161.3
R167 commonsourceibias.n45 commonsourceibias.n42 161.3
R168 commonsourceibias.n47 commonsourceibias.n46 161.3
R169 commonsourceibias.n48 commonsourceibias.n41 161.3
R170 commonsourceibias.n51 commonsourceibias.n50 161.3
R171 commonsourceibias.n52 commonsourceibias.n40 161.3
R172 commonsourceibias.n54 commonsourceibias.n53 161.3
R173 commonsourceibias.n56 commonsourceibias.n38 161.3
R174 commonsourceibias.n58 commonsourceibias.n57 161.3
R175 commonsourceibias.n59 commonsourceibias.n37 161.3
R176 commonsourceibias.n61 commonsourceibias.n60 161.3
R177 commonsourceibias.n62 commonsourceibias.n36 161.3
R178 commonsourceibias.n65 commonsourceibias.n64 161.3
R179 commonsourceibias.n66 commonsourceibias.n35 161.3
R180 commonsourceibias.n68 commonsourceibias.n67 161.3
R181 commonsourceibias.n70 commonsourceibias.n33 161.3
R182 commonsourceibias.n72 commonsourceibias.n71 161.3
R183 commonsourceibias.n73 commonsourceibias.n32 161.3
R184 commonsourceibias.n75 commonsourceibias.n74 161.3
R185 commonsourceibias.n76 commonsourceibias.n31 161.3
R186 commonsourceibias.n79 commonsourceibias.n78 161.3
R187 commonsourceibias.n80 commonsourceibias.n30 161.3
R188 commonsourceibias.n82 commonsourceibias.n81 161.3
R189 commonsourceibias.n84 commonsourceibias.n28 161.3
R190 commonsourceibias.n86 commonsourceibias.n85 161.3
R191 commonsourceibias.n87 commonsourceibias.n27 161.3
R192 commonsourceibias.n89 commonsourceibias.n88 161.3
R193 commonsourceibias.n90 commonsourceibias.n26 161.3
R194 commonsourceibias.n93 commonsourceibias.n92 161.3
R195 commonsourceibias.n94 commonsourceibias.n25 161.3
R196 commonsourceibias.n96 commonsourceibias.n95 161.3
R197 commonsourceibias.n98 commonsourceibias.n23 161.3
R198 commonsourceibias.n100 commonsourceibias.n99 161.3
R199 commonsourceibias.n101 commonsourceibias.n22 161.3
R200 commonsourceibias.n103 commonsourceibias.n102 161.3
R201 commonsourceibias.n104 commonsourceibias.n21 161.3
R202 commonsourceibias.n107 commonsourceibias.n106 161.3
R203 commonsourceibias.n108 commonsourceibias.n20 161.3
R204 commonsourceibias.n110 commonsourceibias.n109 161.3
R205 commonsourceibias.n112 commonsourceibias.n18 161.3
R206 commonsourceibias.n114 commonsourceibias.n113 161.3
R207 commonsourceibias.n115 commonsourceibias.n17 161.3
R208 commonsourceibias.n117 commonsourceibias.n116 161.3
R209 commonsourceibias.n118 commonsourceibias.n16 161.3
R210 commonsourceibias.n121 commonsourceibias.n120 161.3
R211 commonsourceibias.n122 commonsourceibias.n15 161.3
R212 commonsourceibias.n124 commonsourceibias.n123 161.3
R213 commonsourceibias.n126 commonsourceibias.n14 161.3
R214 commonsourceibias.n167 commonsourceibias.n164 161.3
R215 commonsourceibias.n169 commonsourceibias.n168 161.3
R216 commonsourceibias.n170 commonsourceibias.n163 161.3
R217 commonsourceibias.n173 commonsourceibias.n172 161.3
R218 commonsourceibias.n174 commonsourceibias.n162 161.3
R219 commonsourceibias.n176 commonsourceibias.n175 161.3
R220 commonsourceibias.n178 commonsourceibias.n160 161.3
R221 commonsourceibias.n180 commonsourceibias.n179 161.3
R222 commonsourceibias.n181 commonsourceibias.n159 161.3
R223 commonsourceibias.n183 commonsourceibias.n182 161.3
R224 commonsourceibias.n184 commonsourceibias.n158 161.3
R225 commonsourceibias.n187 commonsourceibias.n186 161.3
R226 commonsourceibias.n188 commonsourceibias.n157 161.3
R227 commonsourceibias.n190 commonsourceibias.n189 161.3
R228 commonsourceibias.n192 commonsourceibias.n156 161.3
R229 commonsourceibias.n194 commonsourceibias.n193 161.3
R230 commonsourceibias.n196 commonsourceibias.n195 161.3
R231 commonsourceibias.n197 commonsourceibias.n154 161.3
R232 commonsourceibias.n199 commonsourceibias.n198 161.3
R233 commonsourceibias.n201 commonsourceibias.n200 161.3
R234 commonsourceibias.n202 commonsourceibias.n152 161.3
R235 commonsourceibias.n204 commonsourceibias.n203 161.3
R236 commonsourceibias.n206 commonsourceibias.n205 161.3
R237 commonsourceibias.n208 commonsourceibias.n207 161.3
R238 commonsourceibias.n209 commonsourceibias.n13 161.3
R239 commonsourceibias.n211 commonsourceibias.n210 161.3
R240 commonsourceibias.n212 commonsourceibias.n12 161.3
R241 commonsourceibias.n215 commonsourceibias.n214 161.3
R242 commonsourceibias.n216 commonsourceibias.n11 161.3
R243 commonsourceibias.n218 commonsourceibias.n217 161.3
R244 commonsourceibias.n220 commonsourceibias.n9 161.3
R245 commonsourceibias.n222 commonsourceibias.n221 161.3
R246 commonsourceibias.n223 commonsourceibias.n8 161.3
R247 commonsourceibias.n225 commonsourceibias.n224 161.3
R248 commonsourceibias.n226 commonsourceibias.n7 161.3
R249 commonsourceibias.n229 commonsourceibias.n228 161.3
R250 commonsourceibias.n230 commonsourceibias.n6 161.3
R251 commonsourceibias.n232 commonsourceibias.n231 161.3
R252 commonsourceibias.n234 commonsourceibias.n4 161.3
R253 commonsourceibias.n236 commonsourceibias.n235 161.3
R254 commonsourceibias.n237 commonsourceibias.n3 161.3
R255 commonsourceibias.n239 commonsourceibias.n238 161.3
R256 commonsourceibias.n240 commonsourceibias.n2 161.3
R257 commonsourceibias.n243 commonsourceibias.n242 161.3
R258 commonsourceibias.n244 commonsourceibias.n1 161.3
R259 commonsourceibias.n246 commonsourceibias.n245 161.3
R260 commonsourceibias.n248 commonsourceibias.n0 161.3
R261 commonsourceibias.n730 commonsourceibias.n618 161.3
R262 commonsourceibias.n728 commonsourceibias.n727 161.3
R263 commonsourceibias.n726 commonsourceibias.n619 161.3
R264 commonsourceibias.n725 commonsourceibias.n724 161.3
R265 commonsourceibias.n722 commonsourceibias.n620 161.3
R266 commonsourceibias.n721 commonsourceibias.n720 161.3
R267 commonsourceibias.n719 commonsourceibias.n621 161.3
R268 commonsourceibias.n718 commonsourceibias.n717 161.3
R269 commonsourceibias.n715 commonsourceibias.n622 161.3
R270 commonsourceibias.n713 commonsourceibias.n712 161.3
R271 commonsourceibias.n711 commonsourceibias.n623 161.3
R272 commonsourceibias.n710 commonsourceibias.n709 161.3
R273 commonsourceibias.n707 commonsourceibias.n624 161.3
R274 commonsourceibias.n706 commonsourceibias.n705 161.3
R275 commonsourceibias.n704 commonsourceibias.n625 161.3
R276 commonsourceibias.n703 commonsourceibias.n702 161.3
R277 commonsourceibias.n700 commonsourceibias.n626 161.3
R278 commonsourceibias.n698 commonsourceibias.n697 161.3
R279 commonsourceibias.n696 commonsourceibias.n627 161.3
R280 commonsourceibias.n695 commonsourceibias.n694 161.3
R281 commonsourceibias.n692 commonsourceibias.n628 161.3
R282 commonsourceibias.n691 commonsourceibias.n690 161.3
R283 commonsourceibias.n689 commonsourceibias.n629 161.3
R284 commonsourceibias.n688 commonsourceibias.n687 161.3
R285 commonsourceibias.n685 commonsourceibias.n630 161.3
R286 commonsourceibias.n683 commonsourceibias.n682 161.3
R287 commonsourceibias.n681 commonsourceibias.n631 161.3
R288 commonsourceibias.n680 commonsourceibias.n679 161.3
R289 commonsourceibias.n677 commonsourceibias.n632 161.3
R290 commonsourceibias.n676 commonsourceibias.n675 161.3
R291 commonsourceibias.n674 commonsourceibias.n633 161.3
R292 commonsourceibias.n673 commonsourceibias.n672 161.3
R293 commonsourceibias.n670 commonsourceibias.n634 161.3
R294 commonsourceibias.n668 commonsourceibias.n667 161.3
R295 commonsourceibias.n666 commonsourceibias.n635 161.3
R296 commonsourceibias.n665 commonsourceibias.n664 161.3
R297 commonsourceibias.n662 commonsourceibias.n636 161.3
R298 commonsourceibias.n661 commonsourceibias.n660 161.3
R299 commonsourceibias.n659 commonsourceibias.n637 161.3
R300 commonsourceibias.n658 commonsourceibias.n657 161.3
R301 commonsourceibias.n655 commonsourceibias.n638 161.3
R302 commonsourceibias.n653 commonsourceibias.n652 161.3
R303 commonsourceibias.n651 commonsourceibias.n639 161.3
R304 commonsourceibias.n650 commonsourceibias.n649 161.3
R305 commonsourceibias.n647 commonsourceibias.n640 161.3
R306 commonsourceibias.n646 commonsourceibias.n645 161.3
R307 commonsourceibias.n644 commonsourceibias.n641 161.3
R308 commonsourceibias.n500 commonsourceibias.n388 161.3
R309 commonsourceibias.n498 commonsourceibias.n497 161.3
R310 commonsourceibias.n496 commonsourceibias.n389 161.3
R311 commonsourceibias.n495 commonsourceibias.n494 161.3
R312 commonsourceibias.n492 commonsourceibias.n390 161.3
R313 commonsourceibias.n491 commonsourceibias.n490 161.3
R314 commonsourceibias.n489 commonsourceibias.n391 161.3
R315 commonsourceibias.n488 commonsourceibias.n487 161.3
R316 commonsourceibias.n485 commonsourceibias.n392 161.3
R317 commonsourceibias.n483 commonsourceibias.n482 161.3
R318 commonsourceibias.n481 commonsourceibias.n393 161.3
R319 commonsourceibias.n480 commonsourceibias.n479 161.3
R320 commonsourceibias.n477 commonsourceibias.n394 161.3
R321 commonsourceibias.n476 commonsourceibias.n475 161.3
R322 commonsourceibias.n474 commonsourceibias.n395 161.3
R323 commonsourceibias.n473 commonsourceibias.n472 161.3
R324 commonsourceibias.n470 commonsourceibias.n396 161.3
R325 commonsourceibias.n468 commonsourceibias.n467 161.3
R326 commonsourceibias.n466 commonsourceibias.n397 161.3
R327 commonsourceibias.n465 commonsourceibias.n464 161.3
R328 commonsourceibias.n462 commonsourceibias.n398 161.3
R329 commonsourceibias.n461 commonsourceibias.n460 161.3
R330 commonsourceibias.n459 commonsourceibias.n399 161.3
R331 commonsourceibias.n458 commonsourceibias.n457 161.3
R332 commonsourceibias.n455 commonsourceibias.n400 161.3
R333 commonsourceibias.n453 commonsourceibias.n452 161.3
R334 commonsourceibias.n451 commonsourceibias.n401 161.3
R335 commonsourceibias.n450 commonsourceibias.n449 161.3
R336 commonsourceibias.n447 commonsourceibias.n402 161.3
R337 commonsourceibias.n446 commonsourceibias.n445 161.3
R338 commonsourceibias.n444 commonsourceibias.n403 161.3
R339 commonsourceibias.n443 commonsourceibias.n442 161.3
R340 commonsourceibias.n440 commonsourceibias.n404 161.3
R341 commonsourceibias.n438 commonsourceibias.n437 161.3
R342 commonsourceibias.n436 commonsourceibias.n405 161.3
R343 commonsourceibias.n435 commonsourceibias.n434 161.3
R344 commonsourceibias.n432 commonsourceibias.n406 161.3
R345 commonsourceibias.n431 commonsourceibias.n430 161.3
R346 commonsourceibias.n429 commonsourceibias.n407 161.3
R347 commonsourceibias.n428 commonsourceibias.n427 161.3
R348 commonsourceibias.n425 commonsourceibias.n408 161.3
R349 commonsourceibias.n423 commonsourceibias.n422 161.3
R350 commonsourceibias.n421 commonsourceibias.n409 161.3
R351 commonsourceibias.n420 commonsourceibias.n419 161.3
R352 commonsourceibias.n417 commonsourceibias.n410 161.3
R353 commonsourceibias.n416 commonsourceibias.n415 161.3
R354 commonsourceibias.n414 commonsourceibias.n411 161.3
R355 commonsourceibias.n570 commonsourceibias.n569 161.3
R356 commonsourceibias.n568 commonsourceibias.n567 161.3
R357 commonsourceibias.n566 commonsourceibias.n516 161.3
R358 commonsourceibias.n565 commonsourceibias.n564 161.3
R359 commonsourceibias.n563 commonsourceibias.n562 161.3
R360 commonsourceibias.n561 commonsourceibias.n518 161.3
R361 commonsourceibias.n560 commonsourceibias.n559 161.3
R362 commonsourceibias.n558 commonsourceibias.n557 161.3
R363 commonsourceibias.n556 commonsourceibias.n520 161.3
R364 commonsourceibias.n554 commonsourceibias.n553 161.3
R365 commonsourceibias.n552 commonsourceibias.n521 161.3
R366 commonsourceibias.n551 commonsourceibias.n550 161.3
R367 commonsourceibias.n548 commonsourceibias.n522 161.3
R368 commonsourceibias.n547 commonsourceibias.n546 161.3
R369 commonsourceibias.n545 commonsourceibias.n523 161.3
R370 commonsourceibias.n544 commonsourceibias.n543 161.3
R371 commonsourceibias.n541 commonsourceibias.n524 161.3
R372 commonsourceibias.n539 commonsourceibias.n538 161.3
R373 commonsourceibias.n537 commonsourceibias.n525 161.3
R374 commonsourceibias.n536 commonsourceibias.n535 161.3
R375 commonsourceibias.n533 commonsourceibias.n526 161.3
R376 commonsourceibias.n532 commonsourceibias.n531 161.3
R377 commonsourceibias.n530 commonsourceibias.n527 161.3
R378 commonsourceibias.n615 commonsourceibias.n367 161.3
R379 commonsourceibias.n613 commonsourceibias.n612 161.3
R380 commonsourceibias.n611 commonsourceibias.n368 161.3
R381 commonsourceibias.n610 commonsourceibias.n609 161.3
R382 commonsourceibias.n607 commonsourceibias.n369 161.3
R383 commonsourceibias.n606 commonsourceibias.n605 161.3
R384 commonsourceibias.n604 commonsourceibias.n370 161.3
R385 commonsourceibias.n603 commonsourceibias.n602 161.3
R386 commonsourceibias.n600 commonsourceibias.n371 161.3
R387 commonsourceibias.n598 commonsourceibias.n597 161.3
R388 commonsourceibias.n596 commonsourceibias.n372 161.3
R389 commonsourceibias.n595 commonsourceibias.n594 161.3
R390 commonsourceibias.n592 commonsourceibias.n373 161.3
R391 commonsourceibias.n591 commonsourceibias.n590 161.3
R392 commonsourceibias.n589 commonsourceibias.n374 161.3
R393 commonsourceibias.n588 commonsourceibias.n587 161.3
R394 commonsourceibias.n585 commonsourceibias.n375 161.3
R395 commonsourceibias.n583 commonsourceibias.n582 161.3
R396 commonsourceibias.n581 commonsourceibias.n376 161.3
R397 commonsourceibias.n580 commonsourceibias.n579 161.3
R398 commonsourceibias.n577 commonsourceibias.n377 161.3
R399 commonsourceibias.n576 commonsourceibias.n575 161.3
R400 commonsourceibias.n574 commonsourceibias.n378 161.3
R401 commonsourceibias.n573 commonsourceibias.n572 161.3
R402 commonsourceibias.n141 commonsourceibias.n139 81.5057
R403 commonsourceibias.n381 commonsourceibias.n379 81.5057
R404 commonsourceibias.n141 commonsourceibias.n140 80.9324
R405 commonsourceibias.n143 commonsourceibias.n142 80.9324
R406 commonsourceibias.n145 commonsourceibias.n144 80.9324
R407 commonsourceibias.n147 commonsourceibias.n146 80.9324
R408 commonsourceibias.n138 commonsourceibias.n137 80.9324
R409 commonsourceibias.n136 commonsourceibias.n135 80.9324
R410 commonsourceibias.n134 commonsourceibias.n133 80.9324
R411 commonsourceibias.n132 commonsourceibias.n131 80.9324
R412 commonsourceibias.n130 commonsourceibias.n129 80.9324
R413 commonsourceibias.n504 commonsourceibias.n503 80.9324
R414 commonsourceibias.n506 commonsourceibias.n505 80.9324
R415 commonsourceibias.n508 commonsourceibias.n507 80.9324
R416 commonsourceibias.n510 commonsourceibias.n509 80.9324
R417 commonsourceibias.n512 commonsourceibias.n511 80.9324
R418 commonsourceibias.n387 commonsourceibias.n386 80.9324
R419 commonsourceibias.n385 commonsourceibias.n384 80.9324
R420 commonsourceibias.n383 commonsourceibias.n382 80.9324
R421 commonsourceibias.n381 commonsourceibias.n380 80.9324
R422 commonsourceibias.n365 commonsourceibias.n364 80.6037
R423 commonsourceibias.n128 commonsourceibias.n127 80.6037
R424 commonsourceibias.n250 commonsourceibias.n249 80.6037
R425 commonsourceibias.n732 commonsourceibias.n731 80.6037
R426 commonsourceibias.n502 commonsourceibias.n501 80.6037
R427 commonsourceibias.n617 commonsourceibias.n616 80.6037
R428 commonsourceibias.n322 commonsourceibias.n321 56.5617
R429 commonsourceibias.n336 commonsourceibias.n335 56.5617
R430 commonsourceibias.n85 commonsourceibias.n84 56.5617
R431 commonsourceibias.n71 commonsourceibias.n70 56.5617
R432 commonsourceibias.n207 commonsourceibias.n206 56.5617
R433 commonsourceibias.n193 commonsourceibias.n192 56.5617
R434 commonsourceibias.n687 commonsourceibias.n685 56.5617
R435 commonsourceibias.n702 commonsourceibias.n700 56.5617
R436 commonsourceibias.n457 commonsourceibias.n455 56.5617
R437 commonsourceibias.n472 commonsourceibias.n470 56.5617
R438 commonsourceibias.n572 commonsourceibias.n570 56.5617
R439 commonsourceibias.n294 commonsourceibias.n293 56.5617
R440 commonsourceibias.n308 commonsourceibias.n307 56.5617
R441 commonsourceibias.n350 commonsourceibias.n349 56.5617
R442 commonsourceibias.n113 commonsourceibias.n112 56.5617
R443 commonsourceibias.n99 commonsourceibias.n98 56.5617
R444 commonsourceibias.n57 commonsourceibias.n56 56.5617
R445 commonsourceibias.n235 commonsourceibias.n234 56.5617
R446 commonsourceibias.n221 commonsourceibias.n220 56.5617
R447 commonsourceibias.n179 commonsourceibias.n178 56.5617
R448 commonsourceibias.n657 commonsourceibias.n655 56.5617
R449 commonsourceibias.n672 commonsourceibias.n670 56.5617
R450 commonsourceibias.n717 commonsourceibias.n715 56.5617
R451 commonsourceibias.n427 commonsourceibias.n425 56.5617
R452 commonsourceibias.n442 commonsourceibias.n440 56.5617
R453 commonsourceibias.n487 commonsourceibias.n485 56.5617
R454 commonsourceibias.n602 commonsourceibias.n600 56.5617
R455 commonsourceibias.n587 commonsourceibias.n585 56.5617
R456 commonsourceibias.n543 commonsourceibias.n541 56.5617
R457 commonsourceibias.n557 commonsourceibias.n556 56.5617
R458 commonsourceibias.n285 commonsourceibias.n284 51.2335
R459 commonsourceibias.n357 commonsourceibias.n252 51.2335
R460 commonsourceibias.n120 commonsourceibias.n15 51.2335
R461 commonsourceibias.n48 commonsourceibias.n47 51.2335
R462 commonsourceibias.n242 commonsourceibias.n1 51.2335
R463 commonsourceibias.n170 commonsourceibias.n169 51.2335
R464 commonsourceibias.n647 commonsourceibias.n646 51.2335
R465 commonsourceibias.n724 commonsourceibias.n619 51.2335
R466 commonsourceibias.n417 commonsourceibias.n416 51.2335
R467 commonsourceibias.n494 commonsourceibias.n389 51.2335
R468 commonsourceibias.n609 commonsourceibias.n368 51.2335
R469 commonsourceibias.n533 commonsourceibias.n532 51.2335
R470 commonsourceibias.n364 commonsourceibias.n363 50.9056
R471 commonsourceibias.n127 commonsourceibias.n126 50.9056
R472 commonsourceibias.n249 commonsourceibias.n248 50.9056
R473 commonsourceibias.n731 commonsourceibias.n730 50.9056
R474 commonsourceibias.n501 commonsourceibias.n500 50.9056
R475 commonsourceibias.n616 commonsourceibias.n615 50.9056
R476 commonsourceibias.n299 commonsourceibias.n298 50.2647
R477 commonsourceibias.n343 commonsourceibias.n257 50.2647
R478 commonsourceibias.n106 commonsourceibias.n20 50.2647
R479 commonsourceibias.n62 commonsourceibias.n61 50.2647
R480 commonsourceibias.n228 commonsourceibias.n6 50.2647
R481 commonsourceibias.n184 commonsourceibias.n183 50.2647
R482 commonsourceibias.n662 commonsourceibias.n661 50.2647
R483 commonsourceibias.n709 commonsourceibias.n623 50.2647
R484 commonsourceibias.n432 commonsourceibias.n431 50.2647
R485 commonsourceibias.n479 commonsourceibias.n393 50.2647
R486 commonsourceibias.n594 commonsourceibias.n372 50.2647
R487 commonsourceibias.n548 commonsourceibias.n547 50.2647
R488 commonsourceibias.n281 commonsourceibias.n280 49.9027
R489 commonsourceibias.n44 commonsourceibias.n43 49.9027
R490 commonsourceibias.n166 commonsourceibias.n165 49.9027
R491 commonsourceibias.n643 commonsourceibias.n642 49.9027
R492 commonsourceibias.n413 commonsourceibias.n412 49.9027
R493 commonsourceibias.n529 commonsourceibias.n528 49.9027
R494 commonsourceibias.n313 commonsourceibias.n312 49.296
R495 commonsourceibias.n329 commonsourceibias.n262 49.296
R496 commonsourceibias.n92 commonsourceibias.n25 49.296
R497 commonsourceibias.n76 commonsourceibias.n75 49.296
R498 commonsourceibias.n214 commonsourceibias.n11 49.296
R499 commonsourceibias.n198 commonsourceibias.n197 49.296
R500 commonsourceibias.n677 commonsourceibias.n676 49.296
R501 commonsourceibias.n694 commonsourceibias.n627 49.296
R502 commonsourceibias.n447 commonsourceibias.n446 49.296
R503 commonsourceibias.n464 commonsourceibias.n397 49.296
R504 commonsourceibias.n579 commonsourceibias.n376 49.296
R505 commonsourceibias.n562 commonsourceibias.n561 49.296
R506 commonsourceibias.n315 commonsourceibias.n267 48.3272
R507 commonsourceibias.n327 commonsourceibias.n326 48.3272
R508 commonsourceibias.n90 commonsourceibias.n89 48.3272
R509 commonsourceibias.n78 commonsourceibias.n30 48.3272
R510 commonsourceibias.n212 commonsourceibias.n211 48.3272
R511 commonsourceibias.n202 commonsourceibias.n201 48.3272
R512 commonsourceibias.n679 commonsourceibias.n631 48.3272
R513 commonsourceibias.n692 commonsourceibias.n691 48.3272
R514 commonsourceibias.n449 commonsourceibias.n401 48.3272
R515 commonsourceibias.n462 commonsourceibias.n461 48.3272
R516 commonsourceibias.n577 commonsourceibias.n576 48.3272
R517 commonsourceibias.n566 commonsourceibias.n565 48.3272
R518 commonsourceibias.n301 commonsourceibias.n272 47.3584
R519 commonsourceibias.n341 commonsourceibias.n340 47.3584
R520 commonsourceibias.n104 commonsourceibias.n103 47.3584
R521 commonsourceibias.n64 commonsourceibias.n35 47.3584
R522 commonsourceibias.n226 commonsourceibias.n225 47.3584
R523 commonsourceibias.n186 commonsourceibias.n157 47.3584
R524 commonsourceibias.n664 commonsourceibias.n635 47.3584
R525 commonsourceibias.n707 commonsourceibias.n706 47.3584
R526 commonsourceibias.n434 commonsourceibias.n405 47.3584
R527 commonsourceibias.n477 commonsourceibias.n476 47.3584
R528 commonsourceibias.n592 commonsourceibias.n591 47.3584
R529 commonsourceibias.n550 commonsourceibias.n521 47.3584
R530 commonsourceibias.n287 commonsourceibias.n277 46.3896
R531 commonsourceibias.n355 commonsourceibias.n354 46.3896
R532 commonsourceibias.n118 commonsourceibias.n117 46.3896
R533 commonsourceibias.n50 commonsourceibias.n40 46.3896
R534 commonsourceibias.n240 commonsourceibias.n239 46.3896
R535 commonsourceibias.n172 commonsourceibias.n162 46.3896
R536 commonsourceibias.n649 commonsourceibias.n639 46.3896
R537 commonsourceibias.n722 commonsourceibias.n721 46.3896
R538 commonsourceibias.n419 commonsourceibias.n409 46.3896
R539 commonsourceibias.n492 commonsourceibias.n491 46.3896
R540 commonsourceibias.n607 commonsourceibias.n606 46.3896
R541 commonsourceibias.n535 commonsourceibias.n525 46.3896
R542 commonsourceibias.n282 commonsourceibias.n281 44.7059
R543 commonsourceibias.n644 commonsourceibias.n643 44.7059
R544 commonsourceibias.n414 commonsourceibias.n413 44.7059
R545 commonsourceibias.n530 commonsourceibias.n529 44.7059
R546 commonsourceibias.n45 commonsourceibias.n44 44.7059
R547 commonsourceibias.n167 commonsourceibias.n166 44.7059
R548 commonsourceibias.n291 commonsourceibias.n277 34.7644
R549 commonsourceibias.n354 commonsourceibias.n254 34.7644
R550 commonsourceibias.n117 commonsourceibias.n17 34.7644
R551 commonsourceibias.n54 commonsourceibias.n40 34.7644
R552 commonsourceibias.n239 commonsourceibias.n3 34.7644
R553 commonsourceibias.n176 commonsourceibias.n162 34.7644
R554 commonsourceibias.n653 commonsourceibias.n639 34.7644
R555 commonsourceibias.n721 commonsourceibias.n621 34.7644
R556 commonsourceibias.n423 commonsourceibias.n409 34.7644
R557 commonsourceibias.n491 commonsourceibias.n391 34.7644
R558 commonsourceibias.n606 commonsourceibias.n370 34.7644
R559 commonsourceibias.n539 commonsourceibias.n525 34.7644
R560 commonsourceibias.n305 commonsourceibias.n272 33.7956
R561 commonsourceibias.n340 commonsourceibias.n259 33.7956
R562 commonsourceibias.n103 commonsourceibias.n22 33.7956
R563 commonsourceibias.n68 commonsourceibias.n35 33.7956
R564 commonsourceibias.n225 commonsourceibias.n8 33.7956
R565 commonsourceibias.n190 commonsourceibias.n157 33.7956
R566 commonsourceibias.n668 commonsourceibias.n635 33.7956
R567 commonsourceibias.n706 commonsourceibias.n625 33.7956
R568 commonsourceibias.n438 commonsourceibias.n405 33.7956
R569 commonsourceibias.n476 commonsourceibias.n395 33.7956
R570 commonsourceibias.n591 commonsourceibias.n374 33.7956
R571 commonsourceibias.n554 commonsourceibias.n521 33.7956
R572 commonsourceibias.n319 commonsourceibias.n267 32.8269
R573 commonsourceibias.n326 commonsourceibias.n264 32.8269
R574 commonsourceibias.n89 commonsourceibias.n27 32.8269
R575 commonsourceibias.n82 commonsourceibias.n30 32.8269
R576 commonsourceibias.n211 commonsourceibias.n13 32.8269
R577 commonsourceibias.n203 commonsourceibias.n202 32.8269
R578 commonsourceibias.n683 commonsourceibias.n631 32.8269
R579 commonsourceibias.n691 commonsourceibias.n629 32.8269
R580 commonsourceibias.n453 commonsourceibias.n401 32.8269
R581 commonsourceibias.n461 commonsourceibias.n399 32.8269
R582 commonsourceibias.n576 commonsourceibias.n378 32.8269
R583 commonsourceibias.n567 commonsourceibias.n566 32.8269
R584 commonsourceibias.n312 commonsourceibias.n269 31.8581
R585 commonsourceibias.n333 commonsourceibias.n262 31.8581
R586 commonsourceibias.n96 commonsourceibias.n25 31.8581
R587 commonsourceibias.n75 commonsourceibias.n32 31.8581
R588 commonsourceibias.n218 commonsourceibias.n11 31.8581
R589 commonsourceibias.n197 commonsourceibias.n196 31.8581
R590 commonsourceibias.n676 commonsourceibias.n633 31.8581
R591 commonsourceibias.n698 commonsourceibias.n627 31.8581
R592 commonsourceibias.n446 commonsourceibias.n403 31.8581
R593 commonsourceibias.n468 commonsourceibias.n397 31.8581
R594 commonsourceibias.n583 commonsourceibias.n376 31.8581
R595 commonsourceibias.n561 commonsourceibias.n560 31.8581
R596 commonsourceibias.n298 commonsourceibias.n274 30.8893
R597 commonsourceibias.n347 commonsourceibias.n257 30.8893
R598 commonsourceibias.n110 commonsourceibias.n20 30.8893
R599 commonsourceibias.n61 commonsourceibias.n37 30.8893
R600 commonsourceibias.n232 commonsourceibias.n6 30.8893
R601 commonsourceibias.n183 commonsourceibias.n159 30.8893
R602 commonsourceibias.n661 commonsourceibias.n637 30.8893
R603 commonsourceibias.n713 commonsourceibias.n623 30.8893
R604 commonsourceibias.n431 commonsourceibias.n407 30.8893
R605 commonsourceibias.n483 commonsourceibias.n393 30.8893
R606 commonsourceibias.n598 commonsourceibias.n372 30.8893
R607 commonsourceibias.n547 commonsourceibias.n523 30.8893
R608 commonsourceibias.n284 commonsourceibias.n279 29.9206
R609 commonsourceibias.n361 commonsourceibias.n252 29.9206
R610 commonsourceibias.n124 commonsourceibias.n15 29.9206
R611 commonsourceibias.n47 commonsourceibias.n42 29.9206
R612 commonsourceibias.n246 commonsourceibias.n1 29.9206
R613 commonsourceibias.n169 commonsourceibias.n164 29.9206
R614 commonsourceibias.n646 commonsourceibias.n641 29.9206
R615 commonsourceibias.n728 commonsourceibias.n619 29.9206
R616 commonsourceibias.n416 commonsourceibias.n411 29.9206
R617 commonsourceibias.n498 commonsourceibias.n389 29.9206
R618 commonsourceibias.n613 commonsourceibias.n368 29.9206
R619 commonsourceibias.n532 commonsourceibias.n527 29.9206
R620 commonsourceibias.n363 commonsourceibias.n362 21.8872
R621 commonsourceibias.n126 commonsourceibias.n125 21.8872
R622 commonsourceibias.n248 commonsourceibias.n247 21.8872
R623 commonsourceibias.n730 commonsourceibias.n729 21.8872
R624 commonsourceibias.n500 commonsourceibias.n499 21.8872
R625 commonsourceibias.n615 commonsourceibias.n614 21.8872
R626 commonsourceibias.n294 commonsourceibias.n276 21.3954
R627 commonsourceibias.n349 commonsourceibias.n348 21.3954
R628 commonsourceibias.n112 commonsourceibias.n111 21.3954
R629 commonsourceibias.n57 commonsourceibias.n39 21.3954
R630 commonsourceibias.n234 commonsourceibias.n233 21.3954
R631 commonsourceibias.n179 commonsourceibias.n161 21.3954
R632 commonsourceibias.n657 commonsourceibias.n656 21.3954
R633 commonsourceibias.n715 commonsourceibias.n714 21.3954
R634 commonsourceibias.n427 commonsourceibias.n426 21.3954
R635 commonsourceibias.n485 commonsourceibias.n484 21.3954
R636 commonsourceibias.n600 commonsourceibias.n599 21.3954
R637 commonsourceibias.n543 commonsourceibias.n542 21.3954
R638 commonsourceibias.n308 commonsourceibias.n271 20.9036
R639 commonsourceibias.n335 commonsourceibias.n334 20.9036
R640 commonsourceibias.n98 commonsourceibias.n97 20.9036
R641 commonsourceibias.n71 commonsourceibias.n34 20.9036
R642 commonsourceibias.n220 commonsourceibias.n219 20.9036
R643 commonsourceibias.n193 commonsourceibias.n155 20.9036
R644 commonsourceibias.n672 commonsourceibias.n671 20.9036
R645 commonsourceibias.n700 commonsourceibias.n699 20.9036
R646 commonsourceibias.n442 commonsourceibias.n441 20.9036
R647 commonsourceibias.n470 commonsourceibias.n469 20.9036
R648 commonsourceibias.n585 commonsourceibias.n584 20.9036
R649 commonsourceibias.n557 commonsourceibias.n519 20.9036
R650 commonsourceibias.n321 commonsourceibias.n320 20.4117
R651 commonsourceibias.n322 commonsourceibias.n266 20.4117
R652 commonsourceibias.n85 commonsourceibias.n29 20.4117
R653 commonsourceibias.n84 commonsourceibias.n83 20.4117
R654 commonsourceibias.n207 commonsourceibias.n150 20.4117
R655 commonsourceibias.n206 commonsourceibias.n151 20.4117
R656 commonsourceibias.n685 commonsourceibias.n684 20.4117
R657 commonsourceibias.n687 commonsourceibias.n686 20.4117
R658 commonsourceibias.n455 commonsourceibias.n454 20.4117
R659 commonsourceibias.n457 commonsourceibias.n456 20.4117
R660 commonsourceibias.n572 commonsourceibias.n571 20.4117
R661 commonsourceibias.n570 commonsourceibias.n515 20.4117
R662 commonsourceibias.n307 commonsourceibias.n306 19.9199
R663 commonsourceibias.n336 commonsourceibias.n261 19.9199
R664 commonsourceibias.n99 commonsourceibias.n24 19.9199
R665 commonsourceibias.n70 commonsourceibias.n69 19.9199
R666 commonsourceibias.n221 commonsourceibias.n10 19.9199
R667 commonsourceibias.n192 commonsourceibias.n191 19.9199
R668 commonsourceibias.n670 commonsourceibias.n669 19.9199
R669 commonsourceibias.n702 commonsourceibias.n701 19.9199
R670 commonsourceibias.n440 commonsourceibias.n439 19.9199
R671 commonsourceibias.n472 commonsourceibias.n471 19.9199
R672 commonsourceibias.n587 commonsourceibias.n586 19.9199
R673 commonsourceibias.n556 commonsourceibias.n555 19.9199
R674 commonsourceibias.n293 commonsourceibias.n292 19.4281
R675 commonsourceibias.n350 commonsourceibias.n256 19.4281
R676 commonsourceibias.n113 commonsourceibias.n19 19.4281
R677 commonsourceibias.n56 commonsourceibias.n55 19.4281
R678 commonsourceibias.n235 commonsourceibias.n5 19.4281
R679 commonsourceibias.n178 commonsourceibias.n177 19.4281
R680 commonsourceibias.n655 commonsourceibias.n654 19.4281
R681 commonsourceibias.n717 commonsourceibias.n716 19.4281
R682 commonsourceibias.n425 commonsourceibias.n424 19.4281
R683 commonsourceibias.n487 commonsourceibias.n486 19.4281
R684 commonsourceibias.n602 commonsourceibias.n601 19.4281
R685 commonsourceibias.n541 commonsourceibias.n540 19.4281
R686 commonsourceibias.n286 commonsourceibias.n285 13.526
R687 commonsourceibias.n357 commonsourceibias.n356 13.526
R688 commonsourceibias.n120 commonsourceibias.n119 13.526
R689 commonsourceibias.n49 commonsourceibias.n48 13.526
R690 commonsourceibias.n242 commonsourceibias.n241 13.526
R691 commonsourceibias.n171 commonsourceibias.n170 13.526
R692 commonsourceibias.n648 commonsourceibias.n647 13.526
R693 commonsourceibias.n724 commonsourceibias.n723 13.526
R694 commonsourceibias.n418 commonsourceibias.n417 13.526
R695 commonsourceibias.n494 commonsourceibias.n493 13.526
R696 commonsourceibias.n609 commonsourceibias.n608 13.526
R697 commonsourceibias.n534 commonsourceibias.n533 13.526
R698 commonsourceibias.n130 commonsourceibias.n128 13.2322
R699 commonsourceibias.n504 commonsourceibias.n502 13.2322
R700 commonsourceibias.n300 commonsourceibias.n299 13.0342
R701 commonsourceibias.n343 commonsourceibias.n342 13.0342
R702 commonsourceibias.n106 commonsourceibias.n105 13.0342
R703 commonsourceibias.n63 commonsourceibias.n62 13.0342
R704 commonsourceibias.n228 commonsourceibias.n227 13.0342
R705 commonsourceibias.n185 commonsourceibias.n184 13.0342
R706 commonsourceibias.n663 commonsourceibias.n662 13.0342
R707 commonsourceibias.n709 commonsourceibias.n708 13.0342
R708 commonsourceibias.n433 commonsourceibias.n432 13.0342
R709 commonsourceibias.n479 commonsourceibias.n478 13.0342
R710 commonsourceibias.n594 commonsourceibias.n593 13.0342
R711 commonsourceibias.n549 commonsourceibias.n548 13.0342
R712 commonsourceibias.n314 commonsourceibias.n313 12.5423
R713 commonsourceibias.n329 commonsourceibias.n328 12.5423
R714 commonsourceibias.n92 commonsourceibias.n91 12.5423
R715 commonsourceibias.n77 commonsourceibias.n76 12.5423
R716 commonsourceibias.n214 commonsourceibias.n213 12.5423
R717 commonsourceibias.n198 commonsourceibias.n153 12.5423
R718 commonsourceibias.n678 commonsourceibias.n677 12.5423
R719 commonsourceibias.n694 commonsourceibias.n693 12.5423
R720 commonsourceibias.n448 commonsourceibias.n447 12.5423
R721 commonsourceibias.n464 commonsourceibias.n463 12.5423
R722 commonsourceibias.n579 commonsourceibias.n578 12.5423
R723 commonsourceibias.n562 commonsourceibias.n517 12.5423
R724 commonsourceibias.n315 commonsourceibias.n314 12.0505
R725 commonsourceibias.n328 commonsourceibias.n327 12.0505
R726 commonsourceibias.n91 commonsourceibias.n90 12.0505
R727 commonsourceibias.n78 commonsourceibias.n77 12.0505
R728 commonsourceibias.n213 commonsourceibias.n212 12.0505
R729 commonsourceibias.n201 commonsourceibias.n153 12.0505
R730 commonsourceibias.n679 commonsourceibias.n678 12.0505
R731 commonsourceibias.n693 commonsourceibias.n692 12.0505
R732 commonsourceibias.n449 commonsourceibias.n448 12.0505
R733 commonsourceibias.n463 commonsourceibias.n462 12.0505
R734 commonsourceibias.n578 commonsourceibias.n577 12.0505
R735 commonsourceibias.n565 commonsourceibias.n517 12.0505
R736 commonsourceibias.n734 commonsourceibias.n366 11.9876
R737 commonsourceibias.n301 commonsourceibias.n300 11.5587
R738 commonsourceibias.n342 commonsourceibias.n341 11.5587
R739 commonsourceibias.n105 commonsourceibias.n104 11.5587
R740 commonsourceibias.n64 commonsourceibias.n63 11.5587
R741 commonsourceibias.n227 commonsourceibias.n226 11.5587
R742 commonsourceibias.n186 commonsourceibias.n185 11.5587
R743 commonsourceibias.n664 commonsourceibias.n663 11.5587
R744 commonsourceibias.n708 commonsourceibias.n707 11.5587
R745 commonsourceibias.n434 commonsourceibias.n433 11.5587
R746 commonsourceibias.n478 commonsourceibias.n477 11.5587
R747 commonsourceibias.n593 commonsourceibias.n592 11.5587
R748 commonsourceibias.n550 commonsourceibias.n549 11.5587
R749 commonsourceibias.n287 commonsourceibias.n286 11.0668
R750 commonsourceibias.n356 commonsourceibias.n355 11.0668
R751 commonsourceibias.n119 commonsourceibias.n118 11.0668
R752 commonsourceibias.n50 commonsourceibias.n49 11.0668
R753 commonsourceibias.n241 commonsourceibias.n240 11.0668
R754 commonsourceibias.n172 commonsourceibias.n171 11.0668
R755 commonsourceibias.n649 commonsourceibias.n648 11.0668
R756 commonsourceibias.n723 commonsourceibias.n722 11.0668
R757 commonsourceibias.n419 commonsourceibias.n418 11.0668
R758 commonsourceibias.n493 commonsourceibias.n492 11.0668
R759 commonsourceibias.n608 commonsourceibias.n607 11.0668
R760 commonsourceibias.n535 commonsourceibias.n534 11.0668
R761 commonsourceibias.n734 commonsourceibias.n733 10.3347
R762 commonsourceibias.n149 commonsourceibias.n148 9.50363
R763 commonsourceibias.n514 commonsourceibias.n513 9.50363
R764 commonsourceibias.n366 commonsourceibias.n250 8.75852
R765 commonsourceibias.n733 commonsourceibias.n617 8.75852
R766 commonsourceibias.n292 commonsourceibias.n291 5.16479
R767 commonsourceibias.n256 commonsourceibias.n254 5.16479
R768 commonsourceibias.n19 commonsourceibias.n17 5.16479
R769 commonsourceibias.n55 commonsourceibias.n54 5.16479
R770 commonsourceibias.n5 commonsourceibias.n3 5.16479
R771 commonsourceibias.n177 commonsourceibias.n176 5.16479
R772 commonsourceibias.n654 commonsourceibias.n653 5.16479
R773 commonsourceibias.n716 commonsourceibias.n621 5.16479
R774 commonsourceibias.n424 commonsourceibias.n423 5.16479
R775 commonsourceibias.n486 commonsourceibias.n391 5.16479
R776 commonsourceibias.n601 commonsourceibias.n370 5.16479
R777 commonsourceibias.n540 commonsourceibias.n539 5.16479
R778 commonsourceibias.n366 commonsourceibias.n365 5.03125
R779 commonsourceibias.n733 commonsourceibias.n732 5.03125
R780 commonsourceibias.n306 commonsourceibias.n305 4.67295
R781 commonsourceibias.n261 commonsourceibias.n259 4.67295
R782 commonsourceibias.n24 commonsourceibias.n22 4.67295
R783 commonsourceibias.n69 commonsourceibias.n68 4.67295
R784 commonsourceibias.n10 commonsourceibias.n8 4.67295
R785 commonsourceibias.n191 commonsourceibias.n190 4.67295
R786 commonsourceibias.n669 commonsourceibias.n668 4.67295
R787 commonsourceibias.n701 commonsourceibias.n625 4.67295
R788 commonsourceibias.n439 commonsourceibias.n438 4.67295
R789 commonsourceibias.n471 commonsourceibias.n395 4.67295
R790 commonsourceibias.n586 commonsourceibias.n374 4.67295
R791 commonsourceibias.n555 commonsourceibias.n554 4.67295
R792 commonsourceibias commonsourceibias.n734 4.20978
R793 commonsourceibias.n320 commonsourceibias.n319 4.18111
R794 commonsourceibias.n266 commonsourceibias.n264 4.18111
R795 commonsourceibias.n29 commonsourceibias.n27 4.18111
R796 commonsourceibias.n83 commonsourceibias.n82 4.18111
R797 commonsourceibias.n150 commonsourceibias.n13 4.18111
R798 commonsourceibias.n203 commonsourceibias.n151 4.18111
R799 commonsourceibias.n684 commonsourceibias.n683 4.18111
R800 commonsourceibias.n686 commonsourceibias.n629 4.18111
R801 commonsourceibias.n454 commonsourceibias.n453 4.18111
R802 commonsourceibias.n456 commonsourceibias.n399 4.18111
R803 commonsourceibias.n571 commonsourceibias.n378 4.18111
R804 commonsourceibias.n567 commonsourceibias.n515 4.18111
R805 commonsourceibias.n271 commonsourceibias.n269 3.68928
R806 commonsourceibias.n334 commonsourceibias.n333 3.68928
R807 commonsourceibias.n97 commonsourceibias.n96 3.68928
R808 commonsourceibias.n34 commonsourceibias.n32 3.68928
R809 commonsourceibias.n219 commonsourceibias.n218 3.68928
R810 commonsourceibias.n196 commonsourceibias.n155 3.68928
R811 commonsourceibias.n671 commonsourceibias.n633 3.68928
R812 commonsourceibias.n699 commonsourceibias.n698 3.68928
R813 commonsourceibias.n441 commonsourceibias.n403 3.68928
R814 commonsourceibias.n469 commonsourceibias.n468 3.68928
R815 commonsourceibias.n584 commonsourceibias.n583 3.68928
R816 commonsourceibias.n560 commonsourceibias.n519 3.68928
R817 commonsourceibias.n276 commonsourceibias.n274 3.19744
R818 commonsourceibias.n348 commonsourceibias.n347 3.19744
R819 commonsourceibias.n111 commonsourceibias.n110 3.19744
R820 commonsourceibias.n39 commonsourceibias.n37 3.19744
R821 commonsourceibias.n233 commonsourceibias.n232 3.19744
R822 commonsourceibias.n161 commonsourceibias.n159 3.19744
R823 commonsourceibias.n656 commonsourceibias.n637 3.19744
R824 commonsourceibias.n714 commonsourceibias.n713 3.19744
R825 commonsourceibias.n426 commonsourceibias.n407 3.19744
R826 commonsourceibias.n484 commonsourceibias.n483 3.19744
R827 commonsourceibias.n599 commonsourceibias.n598 3.19744
R828 commonsourceibias.n542 commonsourceibias.n523 3.19744
R829 commonsourceibias.n139 commonsourceibias.t65 2.82907
R830 commonsourceibias.n139 commonsourceibias.t21 2.82907
R831 commonsourceibias.n140 commonsourceibias.t9 2.82907
R832 commonsourceibias.n140 commonsourceibias.t71 2.82907
R833 commonsourceibias.n142 commonsourceibias.t75 2.82907
R834 commonsourceibias.n142 commonsourceibias.t49 2.82907
R835 commonsourceibias.n144 commonsourceibias.t59 2.82907
R836 commonsourceibias.n144 commonsourceibias.t17 2.82907
R837 commonsourceibias.n146 commonsourceibias.t25 2.82907
R838 commonsourceibias.n146 commonsourceibias.t5 2.82907
R839 commonsourceibias.n137 commonsourceibias.t35 2.82907
R840 commonsourceibias.n137 commonsourceibias.t73 2.82907
R841 commonsourceibias.n135 commonsourceibias.t3 2.82907
R842 commonsourceibias.n135 commonsourceibias.t47 2.82907
R843 commonsourceibias.n133 commonsourceibias.t51 2.82907
R844 commonsourceibias.n133 commonsourceibias.t37 2.82907
R845 commonsourceibias.n131 commonsourceibias.t41 2.82907
R846 commonsourceibias.n131 commonsourceibias.t31 2.82907
R847 commonsourceibias.n129 commonsourceibias.t33 2.82907
R848 commonsourceibias.n129 commonsourceibias.t67 2.82907
R849 commonsourceibias.n503 commonsourceibias.t53 2.82907
R850 commonsourceibias.n503 commonsourceibias.t7 2.82907
R851 commonsourceibias.n505 commonsourceibias.t1 2.82907
R852 commonsourceibias.n505 commonsourceibias.t19 2.82907
R853 commonsourceibias.n507 commonsourceibias.t13 2.82907
R854 commonsourceibias.n507 commonsourceibias.t29 2.82907
R855 commonsourceibias.n509 commonsourceibias.t27 2.82907
R856 commonsourceibias.n509 commonsourceibias.t63 2.82907
R857 commonsourceibias.n511 commonsourceibias.t61 2.82907
R858 commonsourceibias.n511 commonsourceibias.t11 2.82907
R859 commonsourceibias.n386 commonsourceibias.t77 2.82907
R860 commonsourceibias.n386 commonsourceibias.t69 2.82907
R861 commonsourceibias.n384 commonsourceibias.t15 2.82907
R862 commonsourceibias.n384 commonsourceibias.t39 2.82907
R863 commonsourceibias.n382 commonsourceibias.t23 2.82907
R864 commonsourceibias.n382 commonsourceibias.t55 2.82907
R865 commonsourceibias.n380 commonsourceibias.t43 2.82907
R866 commonsourceibias.n380 commonsourceibias.t79 2.82907
R867 commonsourceibias.n379 commonsourceibias.t57 2.82907
R868 commonsourceibias.n379 commonsourceibias.t45 2.82907
R869 commonsourceibias.n280 commonsourceibias.n279 2.7056
R870 commonsourceibias.n362 commonsourceibias.n361 2.7056
R871 commonsourceibias.n125 commonsourceibias.n124 2.7056
R872 commonsourceibias.n43 commonsourceibias.n42 2.7056
R873 commonsourceibias.n247 commonsourceibias.n246 2.7056
R874 commonsourceibias.n165 commonsourceibias.n164 2.7056
R875 commonsourceibias.n642 commonsourceibias.n641 2.7056
R876 commonsourceibias.n729 commonsourceibias.n728 2.7056
R877 commonsourceibias.n412 commonsourceibias.n411 2.7056
R878 commonsourceibias.n499 commonsourceibias.n498 2.7056
R879 commonsourceibias.n614 commonsourceibias.n613 2.7056
R880 commonsourceibias.n528 commonsourceibias.n527 2.7056
R881 commonsourceibias.n132 commonsourceibias.n130 0.573776
R882 commonsourceibias.n134 commonsourceibias.n132 0.573776
R883 commonsourceibias.n136 commonsourceibias.n134 0.573776
R884 commonsourceibias.n138 commonsourceibias.n136 0.573776
R885 commonsourceibias.n147 commonsourceibias.n145 0.573776
R886 commonsourceibias.n145 commonsourceibias.n143 0.573776
R887 commonsourceibias.n143 commonsourceibias.n141 0.573776
R888 commonsourceibias.n383 commonsourceibias.n381 0.573776
R889 commonsourceibias.n385 commonsourceibias.n383 0.573776
R890 commonsourceibias.n387 commonsourceibias.n385 0.573776
R891 commonsourceibias.n512 commonsourceibias.n510 0.573776
R892 commonsourceibias.n510 commonsourceibias.n508 0.573776
R893 commonsourceibias.n508 commonsourceibias.n506 0.573776
R894 commonsourceibias.n506 commonsourceibias.n504 0.573776
R895 commonsourceibias.n148 commonsourceibias.n138 0.287138
R896 commonsourceibias.n148 commonsourceibias.n147 0.287138
R897 commonsourceibias.n513 commonsourceibias.n387 0.287138
R898 commonsourceibias.n513 commonsourceibias.n512 0.287138
R899 commonsourceibias.n365 commonsourceibias.n251 0.285035
R900 commonsourceibias.n128 commonsourceibias.n14 0.285035
R901 commonsourceibias.n250 commonsourceibias.n0 0.285035
R902 commonsourceibias.n732 commonsourceibias.n618 0.285035
R903 commonsourceibias.n502 commonsourceibias.n388 0.285035
R904 commonsourceibias.n617 commonsourceibias.n367 0.285035
R905 commonsourceibias.n360 commonsourceibias.n251 0.189894
R906 commonsourceibias.n360 commonsourceibias.n359 0.189894
R907 commonsourceibias.n359 commonsourceibias.n358 0.189894
R908 commonsourceibias.n358 commonsourceibias.n253 0.189894
R909 commonsourceibias.n353 commonsourceibias.n253 0.189894
R910 commonsourceibias.n353 commonsourceibias.n352 0.189894
R911 commonsourceibias.n352 commonsourceibias.n351 0.189894
R912 commonsourceibias.n351 commonsourceibias.n255 0.189894
R913 commonsourceibias.n346 commonsourceibias.n255 0.189894
R914 commonsourceibias.n346 commonsourceibias.n345 0.189894
R915 commonsourceibias.n345 commonsourceibias.n344 0.189894
R916 commonsourceibias.n344 commonsourceibias.n258 0.189894
R917 commonsourceibias.n339 commonsourceibias.n258 0.189894
R918 commonsourceibias.n339 commonsourceibias.n338 0.189894
R919 commonsourceibias.n338 commonsourceibias.n337 0.189894
R920 commonsourceibias.n337 commonsourceibias.n260 0.189894
R921 commonsourceibias.n332 commonsourceibias.n260 0.189894
R922 commonsourceibias.n332 commonsourceibias.n331 0.189894
R923 commonsourceibias.n331 commonsourceibias.n330 0.189894
R924 commonsourceibias.n330 commonsourceibias.n263 0.189894
R925 commonsourceibias.n325 commonsourceibias.n263 0.189894
R926 commonsourceibias.n325 commonsourceibias.n324 0.189894
R927 commonsourceibias.n324 commonsourceibias.n323 0.189894
R928 commonsourceibias.n323 commonsourceibias.n265 0.189894
R929 commonsourceibias.n318 commonsourceibias.n265 0.189894
R930 commonsourceibias.n318 commonsourceibias.n317 0.189894
R931 commonsourceibias.n317 commonsourceibias.n316 0.189894
R932 commonsourceibias.n316 commonsourceibias.n268 0.189894
R933 commonsourceibias.n311 commonsourceibias.n268 0.189894
R934 commonsourceibias.n311 commonsourceibias.n310 0.189894
R935 commonsourceibias.n310 commonsourceibias.n309 0.189894
R936 commonsourceibias.n309 commonsourceibias.n270 0.189894
R937 commonsourceibias.n304 commonsourceibias.n270 0.189894
R938 commonsourceibias.n304 commonsourceibias.n303 0.189894
R939 commonsourceibias.n303 commonsourceibias.n302 0.189894
R940 commonsourceibias.n302 commonsourceibias.n273 0.189894
R941 commonsourceibias.n297 commonsourceibias.n273 0.189894
R942 commonsourceibias.n297 commonsourceibias.n296 0.189894
R943 commonsourceibias.n296 commonsourceibias.n295 0.189894
R944 commonsourceibias.n295 commonsourceibias.n275 0.189894
R945 commonsourceibias.n290 commonsourceibias.n275 0.189894
R946 commonsourceibias.n290 commonsourceibias.n289 0.189894
R947 commonsourceibias.n289 commonsourceibias.n288 0.189894
R948 commonsourceibias.n288 commonsourceibias.n278 0.189894
R949 commonsourceibias.n283 commonsourceibias.n278 0.189894
R950 commonsourceibias.n283 commonsourceibias.n282 0.189894
R951 commonsourceibias.n123 commonsourceibias.n14 0.189894
R952 commonsourceibias.n123 commonsourceibias.n122 0.189894
R953 commonsourceibias.n122 commonsourceibias.n121 0.189894
R954 commonsourceibias.n121 commonsourceibias.n16 0.189894
R955 commonsourceibias.n116 commonsourceibias.n16 0.189894
R956 commonsourceibias.n116 commonsourceibias.n115 0.189894
R957 commonsourceibias.n115 commonsourceibias.n114 0.189894
R958 commonsourceibias.n114 commonsourceibias.n18 0.189894
R959 commonsourceibias.n109 commonsourceibias.n18 0.189894
R960 commonsourceibias.n109 commonsourceibias.n108 0.189894
R961 commonsourceibias.n108 commonsourceibias.n107 0.189894
R962 commonsourceibias.n107 commonsourceibias.n21 0.189894
R963 commonsourceibias.n102 commonsourceibias.n21 0.189894
R964 commonsourceibias.n102 commonsourceibias.n101 0.189894
R965 commonsourceibias.n101 commonsourceibias.n100 0.189894
R966 commonsourceibias.n100 commonsourceibias.n23 0.189894
R967 commonsourceibias.n95 commonsourceibias.n23 0.189894
R968 commonsourceibias.n95 commonsourceibias.n94 0.189894
R969 commonsourceibias.n94 commonsourceibias.n93 0.189894
R970 commonsourceibias.n93 commonsourceibias.n26 0.189894
R971 commonsourceibias.n88 commonsourceibias.n26 0.189894
R972 commonsourceibias.n88 commonsourceibias.n87 0.189894
R973 commonsourceibias.n87 commonsourceibias.n86 0.189894
R974 commonsourceibias.n86 commonsourceibias.n28 0.189894
R975 commonsourceibias.n81 commonsourceibias.n28 0.189894
R976 commonsourceibias.n81 commonsourceibias.n80 0.189894
R977 commonsourceibias.n80 commonsourceibias.n79 0.189894
R978 commonsourceibias.n79 commonsourceibias.n31 0.189894
R979 commonsourceibias.n74 commonsourceibias.n31 0.189894
R980 commonsourceibias.n74 commonsourceibias.n73 0.189894
R981 commonsourceibias.n73 commonsourceibias.n72 0.189894
R982 commonsourceibias.n72 commonsourceibias.n33 0.189894
R983 commonsourceibias.n67 commonsourceibias.n33 0.189894
R984 commonsourceibias.n67 commonsourceibias.n66 0.189894
R985 commonsourceibias.n66 commonsourceibias.n65 0.189894
R986 commonsourceibias.n65 commonsourceibias.n36 0.189894
R987 commonsourceibias.n60 commonsourceibias.n36 0.189894
R988 commonsourceibias.n60 commonsourceibias.n59 0.189894
R989 commonsourceibias.n59 commonsourceibias.n58 0.189894
R990 commonsourceibias.n58 commonsourceibias.n38 0.189894
R991 commonsourceibias.n53 commonsourceibias.n38 0.189894
R992 commonsourceibias.n53 commonsourceibias.n52 0.189894
R993 commonsourceibias.n52 commonsourceibias.n51 0.189894
R994 commonsourceibias.n51 commonsourceibias.n41 0.189894
R995 commonsourceibias.n46 commonsourceibias.n41 0.189894
R996 commonsourceibias.n46 commonsourceibias.n45 0.189894
R997 commonsourceibias.n205 commonsourceibias.n204 0.189894
R998 commonsourceibias.n204 commonsourceibias.n152 0.189894
R999 commonsourceibias.n200 commonsourceibias.n152 0.189894
R1000 commonsourceibias.n200 commonsourceibias.n199 0.189894
R1001 commonsourceibias.n199 commonsourceibias.n154 0.189894
R1002 commonsourceibias.n195 commonsourceibias.n154 0.189894
R1003 commonsourceibias.n195 commonsourceibias.n194 0.189894
R1004 commonsourceibias.n194 commonsourceibias.n156 0.189894
R1005 commonsourceibias.n189 commonsourceibias.n156 0.189894
R1006 commonsourceibias.n189 commonsourceibias.n188 0.189894
R1007 commonsourceibias.n188 commonsourceibias.n187 0.189894
R1008 commonsourceibias.n187 commonsourceibias.n158 0.189894
R1009 commonsourceibias.n182 commonsourceibias.n158 0.189894
R1010 commonsourceibias.n182 commonsourceibias.n181 0.189894
R1011 commonsourceibias.n181 commonsourceibias.n180 0.189894
R1012 commonsourceibias.n180 commonsourceibias.n160 0.189894
R1013 commonsourceibias.n175 commonsourceibias.n160 0.189894
R1014 commonsourceibias.n175 commonsourceibias.n174 0.189894
R1015 commonsourceibias.n174 commonsourceibias.n173 0.189894
R1016 commonsourceibias.n173 commonsourceibias.n163 0.189894
R1017 commonsourceibias.n168 commonsourceibias.n163 0.189894
R1018 commonsourceibias.n168 commonsourceibias.n167 0.189894
R1019 commonsourceibias.n245 commonsourceibias.n0 0.189894
R1020 commonsourceibias.n245 commonsourceibias.n244 0.189894
R1021 commonsourceibias.n244 commonsourceibias.n243 0.189894
R1022 commonsourceibias.n243 commonsourceibias.n2 0.189894
R1023 commonsourceibias.n238 commonsourceibias.n2 0.189894
R1024 commonsourceibias.n238 commonsourceibias.n237 0.189894
R1025 commonsourceibias.n237 commonsourceibias.n236 0.189894
R1026 commonsourceibias.n236 commonsourceibias.n4 0.189894
R1027 commonsourceibias.n231 commonsourceibias.n4 0.189894
R1028 commonsourceibias.n231 commonsourceibias.n230 0.189894
R1029 commonsourceibias.n230 commonsourceibias.n229 0.189894
R1030 commonsourceibias.n229 commonsourceibias.n7 0.189894
R1031 commonsourceibias.n224 commonsourceibias.n7 0.189894
R1032 commonsourceibias.n224 commonsourceibias.n223 0.189894
R1033 commonsourceibias.n223 commonsourceibias.n222 0.189894
R1034 commonsourceibias.n222 commonsourceibias.n9 0.189894
R1035 commonsourceibias.n217 commonsourceibias.n9 0.189894
R1036 commonsourceibias.n217 commonsourceibias.n216 0.189894
R1037 commonsourceibias.n216 commonsourceibias.n215 0.189894
R1038 commonsourceibias.n215 commonsourceibias.n12 0.189894
R1039 commonsourceibias.n210 commonsourceibias.n12 0.189894
R1040 commonsourceibias.n210 commonsourceibias.n209 0.189894
R1041 commonsourceibias.n209 commonsourceibias.n208 0.189894
R1042 commonsourceibias.n645 commonsourceibias.n644 0.189894
R1043 commonsourceibias.n645 commonsourceibias.n640 0.189894
R1044 commonsourceibias.n650 commonsourceibias.n640 0.189894
R1045 commonsourceibias.n651 commonsourceibias.n650 0.189894
R1046 commonsourceibias.n652 commonsourceibias.n651 0.189894
R1047 commonsourceibias.n652 commonsourceibias.n638 0.189894
R1048 commonsourceibias.n658 commonsourceibias.n638 0.189894
R1049 commonsourceibias.n659 commonsourceibias.n658 0.189894
R1050 commonsourceibias.n660 commonsourceibias.n659 0.189894
R1051 commonsourceibias.n660 commonsourceibias.n636 0.189894
R1052 commonsourceibias.n665 commonsourceibias.n636 0.189894
R1053 commonsourceibias.n666 commonsourceibias.n665 0.189894
R1054 commonsourceibias.n667 commonsourceibias.n666 0.189894
R1055 commonsourceibias.n667 commonsourceibias.n634 0.189894
R1056 commonsourceibias.n673 commonsourceibias.n634 0.189894
R1057 commonsourceibias.n674 commonsourceibias.n673 0.189894
R1058 commonsourceibias.n675 commonsourceibias.n674 0.189894
R1059 commonsourceibias.n675 commonsourceibias.n632 0.189894
R1060 commonsourceibias.n680 commonsourceibias.n632 0.189894
R1061 commonsourceibias.n681 commonsourceibias.n680 0.189894
R1062 commonsourceibias.n682 commonsourceibias.n681 0.189894
R1063 commonsourceibias.n682 commonsourceibias.n630 0.189894
R1064 commonsourceibias.n688 commonsourceibias.n630 0.189894
R1065 commonsourceibias.n689 commonsourceibias.n688 0.189894
R1066 commonsourceibias.n690 commonsourceibias.n689 0.189894
R1067 commonsourceibias.n690 commonsourceibias.n628 0.189894
R1068 commonsourceibias.n695 commonsourceibias.n628 0.189894
R1069 commonsourceibias.n696 commonsourceibias.n695 0.189894
R1070 commonsourceibias.n697 commonsourceibias.n696 0.189894
R1071 commonsourceibias.n697 commonsourceibias.n626 0.189894
R1072 commonsourceibias.n703 commonsourceibias.n626 0.189894
R1073 commonsourceibias.n704 commonsourceibias.n703 0.189894
R1074 commonsourceibias.n705 commonsourceibias.n704 0.189894
R1075 commonsourceibias.n705 commonsourceibias.n624 0.189894
R1076 commonsourceibias.n710 commonsourceibias.n624 0.189894
R1077 commonsourceibias.n711 commonsourceibias.n710 0.189894
R1078 commonsourceibias.n712 commonsourceibias.n711 0.189894
R1079 commonsourceibias.n712 commonsourceibias.n622 0.189894
R1080 commonsourceibias.n718 commonsourceibias.n622 0.189894
R1081 commonsourceibias.n719 commonsourceibias.n718 0.189894
R1082 commonsourceibias.n720 commonsourceibias.n719 0.189894
R1083 commonsourceibias.n720 commonsourceibias.n620 0.189894
R1084 commonsourceibias.n725 commonsourceibias.n620 0.189894
R1085 commonsourceibias.n726 commonsourceibias.n725 0.189894
R1086 commonsourceibias.n727 commonsourceibias.n726 0.189894
R1087 commonsourceibias.n727 commonsourceibias.n618 0.189894
R1088 commonsourceibias.n415 commonsourceibias.n414 0.189894
R1089 commonsourceibias.n415 commonsourceibias.n410 0.189894
R1090 commonsourceibias.n420 commonsourceibias.n410 0.189894
R1091 commonsourceibias.n421 commonsourceibias.n420 0.189894
R1092 commonsourceibias.n422 commonsourceibias.n421 0.189894
R1093 commonsourceibias.n422 commonsourceibias.n408 0.189894
R1094 commonsourceibias.n428 commonsourceibias.n408 0.189894
R1095 commonsourceibias.n429 commonsourceibias.n428 0.189894
R1096 commonsourceibias.n430 commonsourceibias.n429 0.189894
R1097 commonsourceibias.n430 commonsourceibias.n406 0.189894
R1098 commonsourceibias.n435 commonsourceibias.n406 0.189894
R1099 commonsourceibias.n436 commonsourceibias.n435 0.189894
R1100 commonsourceibias.n437 commonsourceibias.n436 0.189894
R1101 commonsourceibias.n437 commonsourceibias.n404 0.189894
R1102 commonsourceibias.n443 commonsourceibias.n404 0.189894
R1103 commonsourceibias.n444 commonsourceibias.n443 0.189894
R1104 commonsourceibias.n445 commonsourceibias.n444 0.189894
R1105 commonsourceibias.n445 commonsourceibias.n402 0.189894
R1106 commonsourceibias.n450 commonsourceibias.n402 0.189894
R1107 commonsourceibias.n451 commonsourceibias.n450 0.189894
R1108 commonsourceibias.n452 commonsourceibias.n451 0.189894
R1109 commonsourceibias.n452 commonsourceibias.n400 0.189894
R1110 commonsourceibias.n458 commonsourceibias.n400 0.189894
R1111 commonsourceibias.n459 commonsourceibias.n458 0.189894
R1112 commonsourceibias.n460 commonsourceibias.n459 0.189894
R1113 commonsourceibias.n460 commonsourceibias.n398 0.189894
R1114 commonsourceibias.n465 commonsourceibias.n398 0.189894
R1115 commonsourceibias.n466 commonsourceibias.n465 0.189894
R1116 commonsourceibias.n467 commonsourceibias.n466 0.189894
R1117 commonsourceibias.n467 commonsourceibias.n396 0.189894
R1118 commonsourceibias.n473 commonsourceibias.n396 0.189894
R1119 commonsourceibias.n474 commonsourceibias.n473 0.189894
R1120 commonsourceibias.n475 commonsourceibias.n474 0.189894
R1121 commonsourceibias.n475 commonsourceibias.n394 0.189894
R1122 commonsourceibias.n480 commonsourceibias.n394 0.189894
R1123 commonsourceibias.n481 commonsourceibias.n480 0.189894
R1124 commonsourceibias.n482 commonsourceibias.n481 0.189894
R1125 commonsourceibias.n482 commonsourceibias.n392 0.189894
R1126 commonsourceibias.n488 commonsourceibias.n392 0.189894
R1127 commonsourceibias.n489 commonsourceibias.n488 0.189894
R1128 commonsourceibias.n490 commonsourceibias.n489 0.189894
R1129 commonsourceibias.n490 commonsourceibias.n390 0.189894
R1130 commonsourceibias.n495 commonsourceibias.n390 0.189894
R1131 commonsourceibias.n496 commonsourceibias.n495 0.189894
R1132 commonsourceibias.n497 commonsourceibias.n496 0.189894
R1133 commonsourceibias.n497 commonsourceibias.n388 0.189894
R1134 commonsourceibias.n531 commonsourceibias.n530 0.189894
R1135 commonsourceibias.n531 commonsourceibias.n526 0.189894
R1136 commonsourceibias.n536 commonsourceibias.n526 0.189894
R1137 commonsourceibias.n537 commonsourceibias.n536 0.189894
R1138 commonsourceibias.n538 commonsourceibias.n537 0.189894
R1139 commonsourceibias.n538 commonsourceibias.n524 0.189894
R1140 commonsourceibias.n544 commonsourceibias.n524 0.189894
R1141 commonsourceibias.n545 commonsourceibias.n544 0.189894
R1142 commonsourceibias.n546 commonsourceibias.n545 0.189894
R1143 commonsourceibias.n546 commonsourceibias.n522 0.189894
R1144 commonsourceibias.n551 commonsourceibias.n522 0.189894
R1145 commonsourceibias.n552 commonsourceibias.n551 0.189894
R1146 commonsourceibias.n553 commonsourceibias.n552 0.189894
R1147 commonsourceibias.n553 commonsourceibias.n520 0.189894
R1148 commonsourceibias.n558 commonsourceibias.n520 0.189894
R1149 commonsourceibias.n559 commonsourceibias.n558 0.189894
R1150 commonsourceibias.n559 commonsourceibias.n518 0.189894
R1151 commonsourceibias.n563 commonsourceibias.n518 0.189894
R1152 commonsourceibias.n564 commonsourceibias.n563 0.189894
R1153 commonsourceibias.n564 commonsourceibias.n516 0.189894
R1154 commonsourceibias.n568 commonsourceibias.n516 0.189894
R1155 commonsourceibias.n569 commonsourceibias.n568 0.189894
R1156 commonsourceibias.n574 commonsourceibias.n573 0.189894
R1157 commonsourceibias.n575 commonsourceibias.n574 0.189894
R1158 commonsourceibias.n575 commonsourceibias.n377 0.189894
R1159 commonsourceibias.n580 commonsourceibias.n377 0.189894
R1160 commonsourceibias.n581 commonsourceibias.n580 0.189894
R1161 commonsourceibias.n582 commonsourceibias.n581 0.189894
R1162 commonsourceibias.n582 commonsourceibias.n375 0.189894
R1163 commonsourceibias.n588 commonsourceibias.n375 0.189894
R1164 commonsourceibias.n589 commonsourceibias.n588 0.189894
R1165 commonsourceibias.n590 commonsourceibias.n589 0.189894
R1166 commonsourceibias.n590 commonsourceibias.n373 0.189894
R1167 commonsourceibias.n595 commonsourceibias.n373 0.189894
R1168 commonsourceibias.n596 commonsourceibias.n595 0.189894
R1169 commonsourceibias.n597 commonsourceibias.n596 0.189894
R1170 commonsourceibias.n597 commonsourceibias.n371 0.189894
R1171 commonsourceibias.n603 commonsourceibias.n371 0.189894
R1172 commonsourceibias.n604 commonsourceibias.n603 0.189894
R1173 commonsourceibias.n605 commonsourceibias.n604 0.189894
R1174 commonsourceibias.n605 commonsourceibias.n369 0.189894
R1175 commonsourceibias.n610 commonsourceibias.n369 0.189894
R1176 commonsourceibias.n611 commonsourceibias.n610 0.189894
R1177 commonsourceibias.n612 commonsourceibias.n611 0.189894
R1178 commonsourceibias.n612 commonsourceibias.n367 0.189894
R1179 commonsourceibias.n205 commonsourceibias.n149 0.0762576
R1180 commonsourceibias.n208 commonsourceibias.n149 0.0762576
R1181 commonsourceibias.n569 commonsourceibias.n514 0.0762576
R1182 commonsourceibias.n573 commonsourceibias.n514 0.0762576
R1183 CSoutput.n19 CSoutput.t182 184.661
R1184 CSoutput.n78 CSoutput.n77 165.8
R1185 CSoutput.n76 CSoutput.n0 165.8
R1186 CSoutput.n75 CSoutput.n74 165.8
R1187 CSoutput.n73 CSoutput.n72 165.8
R1188 CSoutput.n71 CSoutput.n2 165.8
R1189 CSoutput.n69 CSoutput.n68 165.8
R1190 CSoutput.n67 CSoutput.n3 165.8
R1191 CSoutput.n66 CSoutput.n65 165.8
R1192 CSoutput.n63 CSoutput.n4 165.8
R1193 CSoutput.n61 CSoutput.n60 165.8
R1194 CSoutput.n59 CSoutput.n5 165.8
R1195 CSoutput.n58 CSoutput.n57 165.8
R1196 CSoutput.n55 CSoutput.n6 165.8
R1197 CSoutput.n54 CSoutput.n53 165.8
R1198 CSoutput.n52 CSoutput.n51 165.8
R1199 CSoutput.n50 CSoutput.n8 165.8
R1200 CSoutput.n48 CSoutput.n47 165.8
R1201 CSoutput.n46 CSoutput.n9 165.8
R1202 CSoutput.n45 CSoutput.n44 165.8
R1203 CSoutput.n42 CSoutput.n10 165.8
R1204 CSoutput.n41 CSoutput.n40 165.8
R1205 CSoutput.n39 CSoutput.n38 165.8
R1206 CSoutput.n37 CSoutput.n12 165.8
R1207 CSoutput.n35 CSoutput.n34 165.8
R1208 CSoutput.n33 CSoutput.n13 165.8
R1209 CSoutput.n32 CSoutput.n31 165.8
R1210 CSoutput.n29 CSoutput.n14 165.8
R1211 CSoutput.n28 CSoutput.n27 165.8
R1212 CSoutput.n26 CSoutput.n25 165.8
R1213 CSoutput.n24 CSoutput.n16 165.8
R1214 CSoutput.n22 CSoutput.n21 165.8
R1215 CSoutput.n20 CSoutput.n17 165.8
R1216 CSoutput.n77 CSoutput.t184 162.194
R1217 CSoutput.n18 CSoutput.t193 120.501
R1218 CSoutput.n23 CSoutput.t195 120.501
R1219 CSoutput.n15 CSoutput.t188 120.501
R1220 CSoutput.n30 CSoutput.t179 120.501
R1221 CSoutput.n36 CSoutput.t197 120.501
R1222 CSoutput.n11 CSoutput.t191 120.501
R1223 CSoutput.n43 CSoutput.t186 120.501
R1224 CSoutput.n49 CSoutput.t177 120.501
R1225 CSoutput.n7 CSoutput.t178 120.501
R1226 CSoutput.n56 CSoutput.t189 120.501
R1227 CSoutput.n62 CSoutput.t185 120.501
R1228 CSoutput.n64 CSoutput.t181 120.501
R1229 CSoutput.n70 CSoutput.t192 120.501
R1230 CSoutput.n1 CSoutput.t194 120.501
R1231 CSoutput.n310 CSoutput.n308 103.469
R1232 CSoutput.n294 CSoutput.n292 103.469
R1233 CSoutput.n279 CSoutput.n277 103.469
R1234 CSoutput.n112 CSoutput.n110 103.469
R1235 CSoutput.n96 CSoutput.n94 103.469
R1236 CSoutput.n81 CSoutput.n79 103.469
R1237 CSoutput.n320 CSoutput.n319 103.111
R1238 CSoutput.n318 CSoutput.n317 103.111
R1239 CSoutput.n316 CSoutput.n315 103.111
R1240 CSoutput.n314 CSoutput.n313 103.111
R1241 CSoutput.n312 CSoutput.n311 103.111
R1242 CSoutput.n310 CSoutput.n309 103.111
R1243 CSoutput.n306 CSoutput.n305 103.111
R1244 CSoutput.n304 CSoutput.n303 103.111
R1245 CSoutput.n302 CSoutput.n301 103.111
R1246 CSoutput.n300 CSoutput.n299 103.111
R1247 CSoutput.n298 CSoutput.n297 103.111
R1248 CSoutput.n296 CSoutput.n295 103.111
R1249 CSoutput.n294 CSoutput.n293 103.111
R1250 CSoutput.n291 CSoutput.n290 103.111
R1251 CSoutput.n289 CSoutput.n288 103.111
R1252 CSoutput.n287 CSoutput.n286 103.111
R1253 CSoutput.n285 CSoutput.n284 103.111
R1254 CSoutput.n283 CSoutput.n282 103.111
R1255 CSoutput.n281 CSoutput.n280 103.111
R1256 CSoutput.n279 CSoutput.n278 103.111
R1257 CSoutput.n112 CSoutput.n111 103.111
R1258 CSoutput.n114 CSoutput.n113 103.111
R1259 CSoutput.n116 CSoutput.n115 103.111
R1260 CSoutput.n118 CSoutput.n117 103.111
R1261 CSoutput.n120 CSoutput.n119 103.111
R1262 CSoutput.n122 CSoutput.n121 103.111
R1263 CSoutput.n124 CSoutput.n123 103.111
R1264 CSoutput.n96 CSoutput.n95 103.111
R1265 CSoutput.n98 CSoutput.n97 103.111
R1266 CSoutput.n100 CSoutput.n99 103.111
R1267 CSoutput.n102 CSoutput.n101 103.111
R1268 CSoutput.n104 CSoutput.n103 103.111
R1269 CSoutput.n106 CSoutput.n105 103.111
R1270 CSoutput.n108 CSoutput.n107 103.111
R1271 CSoutput.n81 CSoutput.n80 103.111
R1272 CSoutput.n83 CSoutput.n82 103.111
R1273 CSoutput.n85 CSoutput.n84 103.111
R1274 CSoutput.n87 CSoutput.n86 103.111
R1275 CSoutput.n89 CSoutput.n88 103.111
R1276 CSoutput.n91 CSoutput.n90 103.111
R1277 CSoutput.n93 CSoutput.n92 103.111
R1278 CSoutput.n322 CSoutput.n321 103.111
R1279 CSoutput.n346 CSoutput.n344 81.5057
R1280 CSoutput.n327 CSoutput.n325 81.5057
R1281 CSoutput.n386 CSoutput.n384 81.5057
R1282 CSoutput.n367 CSoutput.n365 81.5057
R1283 CSoutput.n362 CSoutput.n361 80.9324
R1284 CSoutput.n360 CSoutput.n359 80.9324
R1285 CSoutput.n358 CSoutput.n357 80.9324
R1286 CSoutput.n356 CSoutput.n355 80.9324
R1287 CSoutput.n354 CSoutput.n353 80.9324
R1288 CSoutput.n352 CSoutput.n351 80.9324
R1289 CSoutput.n350 CSoutput.n349 80.9324
R1290 CSoutput.n348 CSoutput.n347 80.9324
R1291 CSoutput.n346 CSoutput.n345 80.9324
R1292 CSoutput.n343 CSoutput.n342 80.9324
R1293 CSoutput.n341 CSoutput.n340 80.9324
R1294 CSoutput.n339 CSoutput.n338 80.9324
R1295 CSoutput.n337 CSoutput.n336 80.9324
R1296 CSoutput.n335 CSoutput.n334 80.9324
R1297 CSoutput.n333 CSoutput.n332 80.9324
R1298 CSoutput.n331 CSoutput.n330 80.9324
R1299 CSoutput.n329 CSoutput.n328 80.9324
R1300 CSoutput.n327 CSoutput.n326 80.9324
R1301 CSoutput.n386 CSoutput.n385 80.9324
R1302 CSoutput.n388 CSoutput.n387 80.9324
R1303 CSoutput.n390 CSoutput.n389 80.9324
R1304 CSoutput.n392 CSoutput.n391 80.9324
R1305 CSoutput.n394 CSoutput.n393 80.9324
R1306 CSoutput.n396 CSoutput.n395 80.9324
R1307 CSoutput.n398 CSoutput.n397 80.9324
R1308 CSoutput.n400 CSoutput.n399 80.9324
R1309 CSoutput.n402 CSoutput.n401 80.9324
R1310 CSoutput.n367 CSoutput.n366 80.9324
R1311 CSoutput.n369 CSoutput.n368 80.9324
R1312 CSoutput.n371 CSoutput.n370 80.9324
R1313 CSoutput.n373 CSoutput.n372 80.9324
R1314 CSoutput.n375 CSoutput.n374 80.9324
R1315 CSoutput.n377 CSoutput.n376 80.9324
R1316 CSoutput.n379 CSoutput.n378 80.9324
R1317 CSoutput.n381 CSoutput.n380 80.9324
R1318 CSoutput.n383 CSoutput.n382 80.9324
R1319 CSoutput.n25 CSoutput.n24 48.1486
R1320 CSoutput.n69 CSoutput.n3 48.1486
R1321 CSoutput.n38 CSoutput.n37 48.1486
R1322 CSoutput.n42 CSoutput.n41 48.1486
R1323 CSoutput.n51 CSoutput.n50 48.1486
R1324 CSoutput.n55 CSoutput.n54 48.1486
R1325 CSoutput.n22 CSoutput.n17 46.462
R1326 CSoutput.n72 CSoutput.n71 46.462
R1327 CSoutput.n20 CSoutput.n19 44.9055
R1328 CSoutput.n29 CSoutput.n28 43.7635
R1329 CSoutput.n65 CSoutput.n63 43.7635
R1330 CSoutput.n35 CSoutput.n13 41.7396
R1331 CSoutput.n57 CSoutput.n5 41.7396
R1332 CSoutput.n44 CSoutput.n9 37.0171
R1333 CSoutput.n48 CSoutput.n9 37.0171
R1334 CSoutput.n76 CSoutput.n75 34.9932
R1335 CSoutput.n31 CSoutput.n13 32.2947
R1336 CSoutput.n61 CSoutput.n5 32.2947
R1337 CSoutput.n30 CSoutput.n29 29.6014
R1338 CSoutput.n63 CSoutput.n62 29.6014
R1339 CSoutput.n19 CSoutput.n18 28.4085
R1340 CSoutput.n18 CSoutput.n17 25.1176
R1341 CSoutput.n72 CSoutput.n1 25.1176
R1342 CSoutput.n43 CSoutput.n42 22.0922
R1343 CSoutput.n50 CSoutput.n49 22.0922
R1344 CSoutput.n77 CSoutput.n76 21.8586
R1345 CSoutput.n37 CSoutput.n36 18.9681
R1346 CSoutput.n56 CSoutput.n55 18.9681
R1347 CSoutput.n25 CSoutput.n15 17.6292
R1348 CSoutput.n64 CSoutput.n3 17.6292
R1349 CSoutput.n24 CSoutput.n23 15.844
R1350 CSoutput.n70 CSoutput.n69 15.844
R1351 CSoutput.n38 CSoutput.n11 14.5051
R1352 CSoutput.n54 CSoutput.n7 14.5051
R1353 CSoutput.n405 CSoutput.n78 11.6139
R1354 CSoutput.n41 CSoutput.n11 11.3811
R1355 CSoutput.n51 CSoutput.n7 11.3811
R1356 CSoutput.n23 CSoutput.n22 10.0422
R1357 CSoutput.n71 CSoutput.n70 10.0422
R1358 CSoutput.n307 CSoutput.n291 9.25285
R1359 CSoutput.n109 CSoutput.n93 9.25285
R1360 CSoutput.n364 CSoutput.n324 9.05363
R1361 CSoutput.n363 CSoutput.n343 8.97993
R1362 CSoutput.n403 CSoutput.n383 8.97993
R1363 CSoutput.n28 CSoutput.n15 8.25698
R1364 CSoutput.n65 CSoutput.n64 8.25698
R1365 CSoutput.n364 CSoutput.n363 7.89345
R1366 CSoutput.n404 CSoutput.n403 7.89345
R1367 CSoutput.n324 CSoutput.n323 7.12641
R1368 CSoutput.n126 CSoutput.n125 7.12641
R1369 CSoutput.n36 CSoutput.n35 6.91809
R1370 CSoutput.n57 CSoutput.n56 6.91809
R1371 CSoutput.n405 CSoutput.n126 5.46119
R1372 CSoutput.n363 CSoutput.n362 5.25266
R1373 CSoutput.n403 CSoutput.n402 5.25266
R1374 CSoutput.n323 CSoutput.n322 5.1449
R1375 CSoutput.n307 CSoutput.n306 5.1449
R1376 CSoutput.n125 CSoutput.n124 5.1449
R1377 CSoutput.n109 CSoutput.n108 5.1449
R1378 CSoutput.n217 CSoutput.n170 4.5005
R1379 CSoutput.n186 CSoutput.n170 4.5005
R1380 CSoutput.n181 CSoutput.n165 4.5005
R1381 CSoutput.n181 CSoutput.n167 4.5005
R1382 CSoutput.n181 CSoutput.n164 4.5005
R1383 CSoutput.n181 CSoutput.n168 4.5005
R1384 CSoutput.n181 CSoutput.n163 4.5005
R1385 CSoutput.n181 CSoutput.t196 4.5005
R1386 CSoutput.n181 CSoutput.n162 4.5005
R1387 CSoutput.n181 CSoutput.n169 4.5005
R1388 CSoutput.n181 CSoutput.n170 4.5005
R1389 CSoutput.n179 CSoutput.n165 4.5005
R1390 CSoutput.n179 CSoutput.n167 4.5005
R1391 CSoutput.n179 CSoutput.n164 4.5005
R1392 CSoutput.n179 CSoutput.n168 4.5005
R1393 CSoutput.n179 CSoutput.n163 4.5005
R1394 CSoutput.n179 CSoutput.t196 4.5005
R1395 CSoutput.n179 CSoutput.n162 4.5005
R1396 CSoutput.n179 CSoutput.n169 4.5005
R1397 CSoutput.n179 CSoutput.n170 4.5005
R1398 CSoutput.n178 CSoutput.n165 4.5005
R1399 CSoutput.n178 CSoutput.n167 4.5005
R1400 CSoutput.n178 CSoutput.n164 4.5005
R1401 CSoutput.n178 CSoutput.n168 4.5005
R1402 CSoutput.n178 CSoutput.n163 4.5005
R1403 CSoutput.n178 CSoutput.t196 4.5005
R1404 CSoutput.n178 CSoutput.n162 4.5005
R1405 CSoutput.n178 CSoutput.n169 4.5005
R1406 CSoutput.n178 CSoutput.n170 4.5005
R1407 CSoutput.n263 CSoutput.n165 4.5005
R1408 CSoutput.n263 CSoutput.n167 4.5005
R1409 CSoutput.n263 CSoutput.n164 4.5005
R1410 CSoutput.n263 CSoutput.n168 4.5005
R1411 CSoutput.n263 CSoutput.n163 4.5005
R1412 CSoutput.n263 CSoutput.t196 4.5005
R1413 CSoutput.n263 CSoutput.n162 4.5005
R1414 CSoutput.n263 CSoutput.n169 4.5005
R1415 CSoutput.n263 CSoutput.n170 4.5005
R1416 CSoutput.n261 CSoutput.n165 4.5005
R1417 CSoutput.n261 CSoutput.n167 4.5005
R1418 CSoutput.n261 CSoutput.n164 4.5005
R1419 CSoutput.n261 CSoutput.n168 4.5005
R1420 CSoutput.n261 CSoutput.n163 4.5005
R1421 CSoutput.n261 CSoutput.t196 4.5005
R1422 CSoutput.n261 CSoutput.n162 4.5005
R1423 CSoutput.n261 CSoutput.n169 4.5005
R1424 CSoutput.n259 CSoutput.n165 4.5005
R1425 CSoutput.n259 CSoutput.n167 4.5005
R1426 CSoutput.n259 CSoutput.n164 4.5005
R1427 CSoutput.n259 CSoutput.n168 4.5005
R1428 CSoutput.n259 CSoutput.n163 4.5005
R1429 CSoutput.n259 CSoutput.t196 4.5005
R1430 CSoutput.n259 CSoutput.n162 4.5005
R1431 CSoutput.n259 CSoutput.n169 4.5005
R1432 CSoutput.n189 CSoutput.n165 4.5005
R1433 CSoutput.n189 CSoutput.n167 4.5005
R1434 CSoutput.n189 CSoutput.n164 4.5005
R1435 CSoutput.n189 CSoutput.n168 4.5005
R1436 CSoutput.n189 CSoutput.n163 4.5005
R1437 CSoutput.n189 CSoutput.t196 4.5005
R1438 CSoutput.n189 CSoutput.n162 4.5005
R1439 CSoutput.n189 CSoutput.n169 4.5005
R1440 CSoutput.n189 CSoutput.n170 4.5005
R1441 CSoutput.n188 CSoutput.n165 4.5005
R1442 CSoutput.n188 CSoutput.n167 4.5005
R1443 CSoutput.n188 CSoutput.n164 4.5005
R1444 CSoutput.n188 CSoutput.n168 4.5005
R1445 CSoutput.n188 CSoutput.n163 4.5005
R1446 CSoutput.n188 CSoutput.t196 4.5005
R1447 CSoutput.n188 CSoutput.n162 4.5005
R1448 CSoutput.n188 CSoutput.n169 4.5005
R1449 CSoutput.n188 CSoutput.n170 4.5005
R1450 CSoutput.n192 CSoutput.n165 4.5005
R1451 CSoutput.n192 CSoutput.n167 4.5005
R1452 CSoutput.n192 CSoutput.n164 4.5005
R1453 CSoutput.n192 CSoutput.n168 4.5005
R1454 CSoutput.n192 CSoutput.n163 4.5005
R1455 CSoutput.n192 CSoutput.t196 4.5005
R1456 CSoutput.n192 CSoutput.n162 4.5005
R1457 CSoutput.n192 CSoutput.n169 4.5005
R1458 CSoutput.n192 CSoutput.n170 4.5005
R1459 CSoutput.n191 CSoutput.n165 4.5005
R1460 CSoutput.n191 CSoutput.n167 4.5005
R1461 CSoutput.n191 CSoutput.n164 4.5005
R1462 CSoutput.n191 CSoutput.n168 4.5005
R1463 CSoutput.n191 CSoutput.n163 4.5005
R1464 CSoutput.n191 CSoutput.t196 4.5005
R1465 CSoutput.n191 CSoutput.n162 4.5005
R1466 CSoutput.n191 CSoutput.n169 4.5005
R1467 CSoutput.n191 CSoutput.n170 4.5005
R1468 CSoutput.n174 CSoutput.n165 4.5005
R1469 CSoutput.n174 CSoutput.n167 4.5005
R1470 CSoutput.n174 CSoutput.n164 4.5005
R1471 CSoutput.n174 CSoutput.n168 4.5005
R1472 CSoutput.n174 CSoutput.n163 4.5005
R1473 CSoutput.n174 CSoutput.t196 4.5005
R1474 CSoutput.n174 CSoutput.n162 4.5005
R1475 CSoutput.n174 CSoutput.n169 4.5005
R1476 CSoutput.n174 CSoutput.n170 4.5005
R1477 CSoutput.n266 CSoutput.n165 4.5005
R1478 CSoutput.n266 CSoutput.n167 4.5005
R1479 CSoutput.n266 CSoutput.n164 4.5005
R1480 CSoutput.n266 CSoutput.n168 4.5005
R1481 CSoutput.n266 CSoutput.n163 4.5005
R1482 CSoutput.n266 CSoutput.t196 4.5005
R1483 CSoutput.n266 CSoutput.n162 4.5005
R1484 CSoutput.n266 CSoutput.n169 4.5005
R1485 CSoutput.n266 CSoutput.n170 4.5005
R1486 CSoutput.n253 CSoutput.n224 4.5005
R1487 CSoutput.n253 CSoutput.n230 4.5005
R1488 CSoutput.n211 CSoutput.n200 4.5005
R1489 CSoutput.n211 CSoutput.n202 4.5005
R1490 CSoutput.n211 CSoutput.n199 4.5005
R1491 CSoutput.n211 CSoutput.n203 4.5005
R1492 CSoutput.n211 CSoutput.n198 4.5005
R1493 CSoutput.n211 CSoutput.t190 4.5005
R1494 CSoutput.n211 CSoutput.n197 4.5005
R1495 CSoutput.n211 CSoutput.n204 4.5005
R1496 CSoutput.n253 CSoutput.n211 4.5005
R1497 CSoutput.n232 CSoutput.n200 4.5005
R1498 CSoutput.n232 CSoutput.n202 4.5005
R1499 CSoutput.n232 CSoutput.n199 4.5005
R1500 CSoutput.n232 CSoutput.n203 4.5005
R1501 CSoutput.n232 CSoutput.n198 4.5005
R1502 CSoutput.n232 CSoutput.t190 4.5005
R1503 CSoutput.n232 CSoutput.n197 4.5005
R1504 CSoutput.n232 CSoutput.n204 4.5005
R1505 CSoutput.n253 CSoutput.n232 4.5005
R1506 CSoutput.n210 CSoutput.n200 4.5005
R1507 CSoutput.n210 CSoutput.n202 4.5005
R1508 CSoutput.n210 CSoutput.n199 4.5005
R1509 CSoutput.n210 CSoutput.n203 4.5005
R1510 CSoutput.n210 CSoutput.n198 4.5005
R1511 CSoutput.n210 CSoutput.t190 4.5005
R1512 CSoutput.n210 CSoutput.n197 4.5005
R1513 CSoutput.n210 CSoutput.n204 4.5005
R1514 CSoutput.n253 CSoutput.n210 4.5005
R1515 CSoutput.n234 CSoutput.n200 4.5005
R1516 CSoutput.n234 CSoutput.n202 4.5005
R1517 CSoutput.n234 CSoutput.n199 4.5005
R1518 CSoutput.n234 CSoutput.n203 4.5005
R1519 CSoutput.n234 CSoutput.n198 4.5005
R1520 CSoutput.n234 CSoutput.t190 4.5005
R1521 CSoutput.n234 CSoutput.n197 4.5005
R1522 CSoutput.n234 CSoutput.n204 4.5005
R1523 CSoutput.n253 CSoutput.n234 4.5005
R1524 CSoutput.n200 CSoutput.n195 4.5005
R1525 CSoutput.n202 CSoutput.n195 4.5005
R1526 CSoutput.n199 CSoutput.n195 4.5005
R1527 CSoutput.n203 CSoutput.n195 4.5005
R1528 CSoutput.n198 CSoutput.n195 4.5005
R1529 CSoutput.t190 CSoutput.n195 4.5005
R1530 CSoutput.n197 CSoutput.n195 4.5005
R1531 CSoutput.n204 CSoutput.n195 4.5005
R1532 CSoutput.n256 CSoutput.n200 4.5005
R1533 CSoutput.n256 CSoutput.n202 4.5005
R1534 CSoutput.n256 CSoutput.n199 4.5005
R1535 CSoutput.n256 CSoutput.n203 4.5005
R1536 CSoutput.n256 CSoutput.n198 4.5005
R1537 CSoutput.n256 CSoutput.t190 4.5005
R1538 CSoutput.n256 CSoutput.n197 4.5005
R1539 CSoutput.n256 CSoutput.n204 4.5005
R1540 CSoutput.n254 CSoutput.n200 4.5005
R1541 CSoutput.n254 CSoutput.n202 4.5005
R1542 CSoutput.n254 CSoutput.n199 4.5005
R1543 CSoutput.n254 CSoutput.n203 4.5005
R1544 CSoutput.n254 CSoutput.n198 4.5005
R1545 CSoutput.n254 CSoutput.t190 4.5005
R1546 CSoutput.n254 CSoutput.n197 4.5005
R1547 CSoutput.n254 CSoutput.n204 4.5005
R1548 CSoutput.n254 CSoutput.n253 4.5005
R1549 CSoutput.n236 CSoutput.n200 4.5005
R1550 CSoutput.n236 CSoutput.n202 4.5005
R1551 CSoutput.n236 CSoutput.n199 4.5005
R1552 CSoutput.n236 CSoutput.n203 4.5005
R1553 CSoutput.n236 CSoutput.n198 4.5005
R1554 CSoutput.n236 CSoutput.t190 4.5005
R1555 CSoutput.n236 CSoutput.n197 4.5005
R1556 CSoutput.n236 CSoutput.n204 4.5005
R1557 CSoutput.n253 CSoutput.n236 4.5005
R1558 CSoutput.n208 CSoutput.n200 4.5005
R1559 CSoutput.n208 CSoutput.n202 4.5005
R1560 CSoutput.n208 CSoutput.n199 4.5005
R1561 CSoutput.n208 CSoutput.n203 4.5005
R1562 CSoutput.n208 CSoutput.n198 4.5005
R1563 CSoutput.n208 CSoutput.t190 4.5005
R1564 CSoutput.n208 CSoutput.n197 4.5005
R1565 CSoutput.n208 CSoutput.n204 4.5005
R1566 CSoutput.n253 CSoutput.n208 4.5005
R1567 CSoutput.n238 CSoutput.n200 4.5005
R1568 CSoutput.n238 CSoutput.n202 4.5005
R1569 CSoutput.n238 CSoutput.n199 4.5005
R1570 CSoutput.n238 CSoutput.n203 4.5005
R1571 CSoutput.n238 CSoutput.n198 4.5005
R1572 CSoutput.n238 CSoutput.t190 4.5005
R1573 CSoutput.n238 CSoutput.n197 4.5005
R1574 CSoutput.n238 CSoutput.n204 4.5005
R1575 CSoutput.n253 CSoutput.n238 4.5005
R1576 CSoutput.n207 CSoutput.n200 4.5005
R1577 CSoutput.n207 CSoutput.n202 4.5005
R1578 CSoutput.n207 CSoutput.n199 4.5005
R1579 CSoutput.n207 CSoutput.n203 4.5005
R1580 CSoutput.n207 CSoutput.n198 4.5005
R1581 CSoutput.n207 CSoutput.t190 4.5005
R1582 CSoutput.n207 CSoutput.n197 4.5005
R1583 CSoutput.n207 CSoutput.n204 4.5005
R1584 CSoutput.n253 CSoutput.n207 4.5005
R1585 CSoutput.n252 CSoutput.n200 4.5005
R1586 CSoutput.n252 CSoutput.n202 4.5005
R1587 CSoutput.n252 CSoutput.n199 4.5005
R1588 CSoutput.n252 CSoutput.n203 4.5005
R1589 CSoutput.n252 CSoutput.n198 4.5005
R1590 CSoutput.n252 CSoutput.t190 4.5005
R1591 CSoutput.n252 CSoutput.n197 4.5005
R1592 CSoutput.n252 CSoutput.n204 4.5005
R1593 CSoutput.n253 CSoutput.n252 4.5005
R1594 CSoutput.n251 CSoutput.n136 4.5005
R1595 CSoutput.n152 CSoutput.n136 4.5005
R1596 CSoutput.n147 CSoutput.n131 4.5005
R1597 CSoutput.n147 CSoutput.n133 4.5005
R1598 CSoutput.n147 CSoutput.n130 4.5005
R1599 CSoutput.n147 CSoutput.n134 4.5005
R1600 CSoutput.n147 CSoutput.n129 4.5005
R1601 CSoutput.n147 CSoutput.t187 4.5005
R1602 CSoutput.n147 CSoutput.n128 4.5005
R1603 CSoutput.n147 CSoutput.n135 4.5005
R1604 CSoutput.n147 CSoutput.n136 4.5005
R1605 CSoutput.n145 CSoutput.n131 4.5005
R1606 CSoutput.n145 CSoutput.n133 4.5005
R1607 CSoutput.n145 CSoutput.n130 4.5005
R1608 CSoutput.n145 CSoutput.n134 4.5005
R1609 CSoutput.n145 CSoutput.n129 4.5005
R1610 CSoutput.n145 CSoutput.t187 4.5005
R1611 CSoutput.n145 CSoutput.n128 4.5005
R1612 CSoutput.n145 CSoutput.n135 4.5005
R1613 CSoutput.n145 CSoutput.n136 4.5005
R1614 CSoutput.n144 CSoutput.n131 4.5005
R1615 CSoutput.n144 CSoutput.n133 4.5005
R1616 CSoutput.n144 CSoutput.n130 4.5005
R1617 CSoutput.n144 CSoutput.n134 4.5005
R1618 CSoutput.n144 CSoutput.n129 4.5005
R1619 CSoutput.n144 CSoutput.t187 4.5005
R1620 CSoutput.n144 CSoutput.n128 4.5005
R1621 CSoutput.n144 CSoutput.n135 4.5005
R1622 CSoutput.n144 CSoutput.n136 4.5005
R1623 CSoutput.n273 CSoutput.n131 4.5005
R1624 CSoutput.n273 CSoutput.n133 4.5005
R1625 CSoutput.n273 CSoutput.n130 4.5005
R1626 CSoutput.n273 CSoutput.n134 4.5005
R1627 CSoutput.n273 CSoutput.n129 4.5005
R1628 CSoutput.n273 CSoutput.t187 4.5005
R1629 CSoutput.n273 CSoutput.n128 4.5005
R1630 CSoutput.n273 CSoutput.n135 4.5005
R1631 CSoutput.n273 CSoutput.n136 4.5005
R1632 CSoutput.n271 CSoutput.n131 4.5005
R1633 CSoutput.n271 CSoutput.n133 4.5005
R1634 CSoutput.n271 CSoutput.n130 4.5005
R1635 CSoutput.n271 CSoutput.n134 4.5005
R1636 CSoutput.n271 CSoutput.n129 4.5005
R1637 CSoutput.n271 CSoutput.t187 4.5005
R1638 CSoutput.n271 CSoutput.n128 4.5005
R1639 CSoutput.n271 CSoutput.n135 4.5005
R1640 CSoutput.n269 CSoutput.n131 4.5005
R1641 CSoutput.n269 CSoutput.n133 4.5005
R1642 CSoutput.n269 CSoutput.n130 4.5005
R1643 CSoutput.n269 CSoutput.n134 4.5005
R1644 CSoutput.n269 CSoutput.n129 4.5005
R1645 CSoutput.n269 CSoutput.t187 4.5005
R1646 CSoutput.n269 CSoutput.n128 4.5005
R1647 CSoutput.n269 CSoutput.n135 4.5005
R1648 CSoutput.n155 CSoutput.n131 4.5005
R1649 CSoutput.n155 CSoutput.n133 4.5005
R1650 CSoutput.n155 CSoutput.n130 4.5005
R1651 CSoutput.n155 CSoutput.n134 4.5005
R1652 CSoutput.n155 CSoutput.n129 4.5005
R1653 CSoutput.n155 CSoutput.t187 4.5005
R1654 CSoutput.n155 CSoutput.n128 4.5005
R1655 CSoutput.n155 CSoutput.n135 4.5005
R1656 CSoutput.n155 CSoutput.n136 4.5005
R1657 CSoutput.n154 CSoutput.n131 4.5005
R1658 CSoutput.n154 CSoutput.n133 4.5005
R1659 CSoutput.n154 CSoutput.n130 4.5005
R1660 CSoutput.n154 CSoutput.n134 4.5005
R1661 CSoutput.n154 CSoutput.n129 4.5005
R1662 CSoutput.n154 CSoutput.t187 4.5005
R1663 CSoutput.n154 CSoutput.n128 4.5005
R1664 CSoutput.n154 CSoutput.n135 4.5005
R1665 CSoutput.n154 CSoutput.n136 4.5005
R1666 CSoutput.n158 CSoutput.n131 4.5005
R1667 CSoutput.n158 CSoutput.n133 4.5005
R1668 CSoutput.n158 CSoutput.n130 4.5005
R1669 CSoutput.n158 CSoutput.n134 4.5005
R1670 CSoutput.n158 CSoutput.n129 4.5005
R1671 CSoutput.n158 CSoutput.t187 4.5005
R1672 CSoutput.n158 CSoutput.n128 4.5005
R1673 CSoutput.n158 CSoutput.n135 4.5005
R1674 CSoutput.n158 CSoutput.n136 4.5005
R1675 CSoutput.n157 CSoutput.n131 4.5005
R1676 CSoutput.n157 CSoutput.n133 4.5005
R1677 CSoutput.n157 CSoutput.n130 4.5005
R1678 CSoutput.n157 CSoutput.n134 4.5005
R1679 CSoutput.n157 CSoutput.n129 4.5005
R1680 CSoutput.n157 CSoutput.t187 4.5005
R1681 CSoutput.n157 CSoutput.n128 4.5005
R1682 CSoutput.n157 CSoutput.n135 4.5005
R1683 CSoutput.n157 CSoutput.n136 4.5005
R1684 CSoutput.n140 CSoutput.n131 4.5005
R1685 CSoutput.n140 CSoutput.n133 4.5005
R1686 CSoutput.n140 CSoutput.n130 4.5005
R1687 CSoutput.n140 CSoutput.n134 4.5005
R1688 CSoutput.n140 CSoutput.n129 4.5005
R1689 CSoutput.n140 CSoutput.t187 4.5005
R1690 CSoutput.n140 CSoutput.n128 4.5005
R1691 CSoutput.n140 CSoutput.n135 4.5005
R1692 CSoutput.n140 CSoutput.n136 4.5005
R1693 CSoutput.n276 CSoutput.n131 4.5005
R1694 CSoutput.n276 CSoutput.n133 4.5005
R1695 CSoutput.n276 CSoutput.n130 4.5005
R1696 CSoutput.n276 CSoutput.n134 4.5005
R1697 CSoutput.n276 CSoutput.n129 4.5005
R1698 CSoutput.n276 CSoutput.t187 4.5005
R1699 CSoutput.n276 CSoutput.n128 4.5005
R1700 CSoutput.n276 CSoutput.n135 4.5005
R1701 CSoutput.n276 CSoutput.n136 4.5005
R1702 CSoutput.n323 CSoutput.n307 4.10845
R1703 CSoutput.n125 CSoutput.n109 4.10845
R1704 CSoutput.n321 CSoutput.t158 4.06363
R1705 CSoutput.n321 CSoutput.t4 4.06363
R1706 CSoutput.n319 CSoutput.t39 4.06363
R1707 CSoutput.n319 CSoutput.t15 4.06363
R1708 CSoutput.n317 CSoutput.t53 4.06363
R1709 CSoutput.n317 CSoutput.t12 4.06363
R1710 CSoutput.n315 CSoutput.t169 4.06363
R1711 CSoutput.n315 CSoutput.t174 4.06363
R1712 CSoutput.n313 CSoutput.t26 4.06363
R1713 CSoutput.n313 CSoutput.t43 4.06363
R1714 CSoutput.n311 CSoutput.t70 4.06363
R1715 CSoutput.n311 CSoutput.t22 4.06363
R1716 CSoutput.n309 CSoutput.t64 4.06363
R1717 CSoutput.n309 CSoutput.t54 4.06363
R1718 CSoutput.n308 CSoutput.t19 4.06363
R1719 CSoutput.n308 CSoutput.t56 4.06363
R1720 CSoutput.n305 CSoutput.t59 4.06363
R1721 CSoutput.n305 CSoutput.t35 4.06363
R1722 CSoutput.n303 CSoutput.t76 4.06363
R1723 CSoutput.n303 CSoutput.t10 4.06363
R1724 CSoutput.n301 CSoutput.t52 4.06363
R1725 CSoutput.n301 CSoutput.t13 4.06363
R1726 CSoutput.n299 CSoutput.t75 4.06363
R1727 CSoutput.n299 CSoutput.t60 4.06363
R1728 CSoutput.n297 CSoutput.t5 4.06363
R1729 CSoutput.n297 CSoutput.t77 4.06363
R1730 CSoutput.n295 CSoutput.t170 4.06363
R1731 CSoutput.n295 CSoutput.t45 4.06363
R1732 CSoutput.n293 CSoutput.t57 4.06363
R1733 CSoutput.n293 CSoutput.t67 4.06363
R1734 CSoutput.n292 CSoutput.t162 4.06363
R1735 CSoutput.n292 CSoutput.t171 4.06363
R1736 CSoutput.n290 CSoutput.t165 4.06363
R1737 CSoutput.n290 CSoutput.t55 4.06363
R1738 CSoutput.n288 CSoutput.t42 4.06363
R1739 CSoutput.n288 CSoutput.t23 4.06363
R1740 CSoutput.n286 CSoutput.t37 4.06363
R1741 CSoutput.n286 CSoutput.t28 4.06363
R1742 CSoutput.n284 CSoutput.t41 4.06363
R1743 CSoutput.n284 CSoutput.t159 4.06363
R1744 CSoutput.n282 CSoutput.t36 4.06363
R1745 CSoutput.n282 CSoutput.t161 4.06363
R1746 CSoutput.n280 CSoutput.t44 4.06363
R1747 CSoutput.n280 CSoutput.t51 4.06363
R1748 CSoutput.n278 CSoutput.t7 4.06363
R1749 CSoutput.n278 CSoutput.t160 4.06363
R1750 CSoutput.n277 CSoutput.t173 4.06363
R1751 CSoutput.n277 CSoutput.t20 4.06363
R1752 CSoutput.n110 CSoutput.t32 4.06363
R1753 CSoutput.n110 CSoutput.t33 4.06363
R1754 CSoutput.n111 CSoutput.t31 4.06363
R1755 CSoutput.n111 CSoutput.t1 4.06363
R1756 CSoutput.n113 CSoutput.t16 4.06363
R1757 CSoutput.n113 CSoutput.t49 4.06363
R1758 CSoutput.n115 CSoutput.t40 4.06363
R1759 CSoutput.n115 CSoutput.t47 4.06363
R1760 CSoutput.n117 CSoutput.t172 4.06363
R1761 CSoutput.n117 CSoutput.t163 4.06363
R1762 CSoutput.n119 CSoutput.t17 4.06363
R1763 CSoutput.n119 CSoutput.t3 4.06363
R1764 CSoutput.n121 CSoutput.t168 4.06363
R1765 CSoutput.n121 CSoutput.t66 4.06363
R1766 CSoutput.n123 CSoutput.t166 4.06363
R1767 CSoutput.n123 CSoutput.t69 4.06363
R1768 CSoutput.n94 CSoutput.t62 4.06363
R1769 CSoutput.n94 CSoutput.t18 4.06363
R1770 CSoutput.n95 CSoutput.t29 4.06363
R1771 CSoutput.n95 CSoutput.t68 4.06363
R1772 CSoutput.n97 CSoutput.t34 4.06363
R1773 CSoutput.n97 CSoutput.t27 4.06363
R1774 CSoutput.n99 CSoutput.t8 4.06363
R1775 CSoutput.n99 CSoutput.t9 4.06363
R1776 CSoutput.n101 CSoutput.t11 4.06363
R1777 CSoutput.n101 CSoutput.t6 4.06363
R1778 CSoutput.n103 CSoutput.t65 4.06363
R1779 CSoutput.n103 CSoutput.t74 4.06363
R1780 CSoutput.n105 CSoutput.t46 4.06363
R1781 CSoutput.n105 CSoutput.t0 4.06363
R1782 CSoutput.n107 CSoutput.t164 4.06363
R1783 CSoutput.n107 CSoutput.t30 4.06363
R1784 CSoutput.n79 CSoutput.t167 4.06363
R1785 CSoutput.n79 CSoutput.t72 4.06363
R1786 CSoutput.n80 CSoutput.t63 4.06363
R1787 CSoutput.n80 CSoutput.t14 4.06363
R1788 CSoutput.n82 CSoutput.t38 4.06363
R1789 CSoutput.n82 CSoutput.t61 4.06363
R1790 CSoutput.n84 CSoutput.t24 4.06363
R1791 CSoutput.n84 CSoutput.t21 4.06363
R1792 CSoutput.n86 CSoutput.t25 4.06363
R1793 CSoutput.n86 CSoutput.t73 4.06363
R1794 CSoutput.n88 CSoutput.t50 4.06363
R1795 CSoutput.n88 CSoutput.t58 4.06363
R1796 CSoutput.n90 CSoutput.t175 4.06363
R1797 CSoutput.n90 CSoutput.t2 4.06363
R1798 CSoutput.n92 CSoutput.t48 4.06363
R1799 CSoutput.n92 CSoutput.t71 4.06363
R1800 CSoutput.n44 CSoutput.n43 3.79402
R1801 CSoutput.n49 CSoutput.n48 3.79402
R1802 CSoutput.n405 CSoutput.n404 3.57343
R1803 CSoutput.n404 CSoutput.n364 3.42304
R1804 CSoutput.n361 CSoutput.t139 2.82907
R1805 CSoutput.n361 CSoutput.t95 2.82907
R1806 CSoutput.n359 CSoutput.t118 2.82907
R1807 CSoutput.n359 CSoutput.t146 2.82907
R1808 CSoutput.n357 CSoutput.t79 2.82907
R1809 CSoutput.n357 CSoutput.t97 2.82907
R1810 CSoutput.n355 CSoutput.t109 2.82907
R1811 CSoutput.n355 CSoutput.t127 2.82907
R1812 CSoutput.n353 CSoutput.t87 2.82907
R1813 CSoutput.n353 CSoutput.t98 2.82907
R1814 CSoutput.n351 CSoutput.t102 2.82907
R1815 CSoutput.n351 CSoutput.t117 2.82907
R1816 CSoutput.n349 CSoutput.t140 2.82907
R1817 CSoutput.n349 CSoutput.t99 2.82907
R1818 CSoutput.n347 CSoutput.t105 2.82907
R1819 CSoutput.n347 CSoutput.t121 2.82907
R1820 CSoutput.n345 CSoutput.t83 2.82907
R1821 CSoutput.n345 CSoutput.t86 2.82907
R1822 CSoutput.n344 CSoutput.t96 2.82907
R1823 CSoutput.n344 CSoutput.t129 2.82907
R1824 CSoutput.n342 CSoutput.t80 2.82907
R1825 CSoutput.n342 CSoutput.t111 2.82907
R1826 CSoutput.n340 CSoutput.t138 2.82907
R1827 CSoutput.n340 CSoutput.t93 2.82907
R1828 CSoutput.n338 CSoutput.t103 2.82907
R1829 CSoutput.n338 CSoutput.t119 2.82907
R1830 CSoutput.n336 CSoutput.t128 2.82907
R1831 CSoutput.n336 CSoutput.t130 2.82907
R1832 CSoutput.n334 CSoutput.t107 2.82907
R1833 CSoutput.n334 CSoutput.t110 2.82907
R1834 CSoutput.n332 CSoutput.t104 2.82907
R1835 CSoutput.n332 CSoutput.t137 2.82907
R1836 CSoutput.n330 CSoutput.t81 2.82907
R1837 CSoutput.n330 CSoutput.t114 2.82907
R1838 CSoutput.n328 CSoutput.t123 2.82907
R1839 CSoutput.n328 CSoutput.t152 2.82907
R1840 CSoutput.n326 CSoutput.t89 2.82907
R1841 CSoutput.n326 CSoutput.t90 2.82907
R1842 CSoutput.n325 CSoutput.t113 2.82907
R1843 CSoutput.n325 CSoutput.t133 2.82907
R1844 CSoutput.n384 CSoutput.t155 2.82907
R1845 CSoutput.n384 CSoutput.t126 2.82907
R1846 CSoutput.n385 CSoutput.t88 2.82907
R1847 CSoutput.n385 CSoutput.t149 2.82907
R1848 CSoutput.n387 CSoutput.t144 2.82907
R1849 CSoutput.n387 CSoutput.t136 2.82907
R1850 CSoutput.n389 CSoutput.t85 2.82907
R1851 CSoutput.n389 CSoutput.t153 2.82907
R1852 CSoutput.n391 CSoutput.t131 2.82907
R1853 CSoutput.n391 CSoutput.t115 2.82907
R1854 CSoutput.n393 CSoutput.t108 2.82907
R1855 CSoutput.n393 CSoutput.t91 2.82907
R1856 CSoutput.n395 CSoutput.t154 2.82907
R1857 CSoutput.n395 CSoutput.t122 2.82907
R1858 CSoutput.n397 CSoutput.t112 2.82907
R1859 CSoutput.n397 CSoutput.t100 2.82907
R1860 CSoutput.n399 CSoutput.t142 2.82907
R1861 CSoutput.n399 CSoutput.t132 2.82907
R1862 CSoutput.n401 CSoutput.t106 2.82907
R1863 CSoutput.n401 CSoutput.t145 2.82907
R1864 CSoutput.n365 CSoutput.t150 2.82907
R1865 CSoutput.n365 CSoutput.t156 2.82907
R1866 CSoutput.n366 CSoutput.t120 2.82907
R1867 CSoutput.n366 CSoutput.t94 2.82907
R1868 CSoutput.n368 CSoutput.t84 2.82907
R1869 CSoutput.n368 CSoutput.t151 2.82907
R1870 CSoutput.n370 CSoutput.t157 2.82907
R1871 CSoutput.n370 CSoutput.t147 2.82907
R1872 CSoutput.n372 CSoutput.t143 2.82907
R1873 CSoutput.n372 CSoutput.t135 2.82907
R1874 CSoutput.n374 CSoutput.t125 2.82907
R1875 CSoutput.n374 CSoutput.t101 2.82907
R1876 CSoutput.n376 CSoutput.t148 2.82907
R1877 CSoutput.n376 CSoutput.t78 2.82907
R1878 CSoutput.n378 CSoutput.t134 2.82907
R1879 CSoutput.n378 CSoutput.t116 2.82907
R1880 CSoutput.n380 CSoutput.t82 2.82907
R1881 CSoutput.n380 CSoutput.t141 2.82907
R1882 CSoutput.n382 CSoutput.t124 2.82907
R1883 CSoutput.n382 CSoutput.t92 2.82907
R1884 CSoutput.n75 CSoutput.n1 2.45513
R1885 CSoutput.n324 CSoutput.n126 2.36742
R1886 CSoutput.n217 CSoutput.n215 2.251
R1887 CSoutput.n217 CSoutput.n214 2.251
R1888 CSoutput.n217 CSoutput.n213 2.251
R1889 CSoutput.n217 CSoutput.n212 2.251
R1890 CSoutput.n186 CSoutput.n185 2.251
R1891 CSoutput.n186 CSoutput.n184 2.251
R1892 CSoutput.n186 CSoutput.n183 2.251
R1893 CSoutput.n186 CSoutput.n182 2.251
R1894 CSoutput.n259 CSoutput.n258 2.251
R1895 CSoutput.n224 CSoutput.n222 2.251
R1896 CSoutput.n224 CSoutput.n221 2.251
R1897 CSoutput.n224 CSoutput.n220 2.251
R1898 CSoutput.n242 CSoutput.n224 2.251
R1899 CSoutput.n230 CSoutput.n229 2.251
R1900 CSoutput.n230 CSoutput.n228 2.251
R1901 CSoutput.n230 CSoutput.n227 2.251
R1902 CSoutput.n230 CSoutput.n226 2.251
R1903 CSoutput.n256 CSoutput.n196 2.251
R1904 CSoutput.n251 CSoutput.n249 2.251
R1905 CSoutput.n251 CSoutput.n248 2.251
R1906 CSoutput.n251 CSoutput.n247 2.251
R1907 CSoutput.n251 CSoutput.n246 2.251
R1908 CSoutput.n152 CSoutput.n151 2.251
R1909 CSoutput.n152 CSoutput.n150 2.251
R1910 CSoutput.n152 CSoutput.n149 2.251
R1911 CSoutput.n152 CSoutput.n148 2.251
R1912 CSoutput.n269 CSoutput.n268 2.251
R1913 CSoutput.n186 CSoutput.n166 2.2505
R1914 CSoutput.n181 CSoutput.n166 2.2505
R1915 CSoutput.n179 CSoutput.n166 2.2505
R1916 CSoutput.n178 CSoutput.n166 2.2505
R1917 CSoutput.n263 CSoutput.n166 2.2505
R1918 CSoutput.n261 CSoutput.n166 2.2505
R1919 CSoutput.n259 CSoutput.n166 2.2505
R1920 CSoutput.n189 CSoutput.n166 2.2505
R1921 CSoutput.n188 CSoutput.n166 2.2505
R1922 CSoutput.n192 CSoutput.n166 2.2505
R1923 CSoutput.n191 CSoutput.n166 2.2505
R1924 CSoutput.n174 CSoutput.n166 2.2505
R1925 CSoutput.n266 CSoutput.n166 2.2505
R1926 CSoutput.n266 CSoutput.n265 2.2505
R1927 CSoutput.n230 CSoutput.n201 2.2505
R1928 CSoutput.n211 CSoutput.n201 2.2505
R1929 CSoutput.n232 CSoutput.n201 2.2505
R1930 CSoutput.n210 CSoutput.n201 2.2505
R1931 CSoutput.n234 CSoutput.n201 2.2505
R1932 CSoutput.n201 CSoutput.n195 2.2505
R1933 CSoutput.n256 CSoutput.n201 2.2505
R1934 CSoutput.n254 CSoutput.n201 2.2505
R1935 CSoutput.n236 CSoutput.n201 2.2505
R1936 CSoutput.n208 CSoutput.n201 2.2505
R1937 CSoutput.n238 CSoutput.n201 2.2505
R1938 CSoutput.n207 CSoutput.n201 2.2505
R1939 CSoutput.n252 CSoutput.n201 2.2505
R1940 CSoutput.n252 CSoutput.n205 2.2505
R1941 CSoutput.n152 CSoutput.n132 2.2505
R1942 CSoutput.n147 CSoutput.n132 2.2505
R1943 CSoutput.n145 CSoutput.n132 2.2505
R1944 CSoutput.n144 CSoutput.n132 2.2505
R1945 CSoutput.n273 CSoutput.n132 2.2505
R1946 CSoutput.n271 CSoutput.n132 2.2505
R1947 CSoutput.n269 CSoutput.n132 2.2505
R1948 CSoutput.n155 CSoutput.n132 2.2505
R1949 CSoutput.n154 CSoutput.n132 2.2505
R1950 CSoutput.n158 CSoutput.n132 2.2505
R1951 CSoutput.n157 CSoutput.n132 2.2505
R1952 CSoutput.n140 CSoutput.n132 2.2505
R1953 CSoutput.n276 CSoutput.n132 2.2505
R1954 CSoutput.n276 CSoutput.n275 2.2505
R1955 CSoutput.n194 CSoutput.n187 2.25024
R1956 CSoutput.n194 CSoutput.n180 2.25024
R1957 CSoutput.n262 CSoutput.n194 2.25024
R1958 CSoutput.n194 CSoutput.n190 2.25024
R1959 CSoutput.n194 CSoutput.n193 2.25024
R1960 CSoutput.n194 CSoutput.n161 2.25024
R1961 CSoutput.n244 CSoutput.n241 2.25024
R1962 CSoutput.n244 CSoutput.n240 2.25024
R1963 CSoutput.n244 CSoutput.n239 2.25024
R1964 CSoutput.n244 CSoutput.n206 2.25024
R1965 CSoutput.n244 CSoutput.n243 2.25024
R1966 CSoutput.n245 CSoutput.n244 2.25024
R1967 CSoutput.n160 CSoutput.n153 2.25024
R1968 CSoutput.n160 CSoutput.n146 2.25024
R1969 CSoutput.n272 CSoutput.n160 2.25024
R1970 CSoutput.n160 CSoutput.n156 2.25024
R1971 CSoutput.n160 CSoutput.n159 2.25024
R1972 CSoutput.n160 CSoutput.n127 2.25024
R1973 CSoutput.n261 CSoutput.n171 1.50111
R1974 CSoutput.n209 CSoutput.n195 1.50111
R1975 CSoutput.n271 CSoutput.n137 1.50111
R1976 CSoutput.n217 CSoutput.n216 1.501
R1977 CSoutput.n224 CSoutput.n223 1.501
R1978 CSoutput.n251 CSoutput.n250 1.501
R1979 CSoutput.n265 CSoutput.n176 1.12536
R1980 CSoutput.n265 CSoutput.n177 1.12536
R1981 CSoutput.n265 CSoutput.n264 1.12536
R1982 CSoutput.n225 CSoutput.n205 1.12536
R1983 CSoutput.n231 CSoutput.n205 1.12536
R1984 CSoutput.n233 CSoutput.n205 1.12536
R1985 CSoutput.n275 CSoutput.n142 1.12536
R1986 CSoutput.n275 CSoutput.n143 1.12536
R1987 CSoutput.n275 CSoutput.n274 1.12536
R1988 CSoutput.n265 CSoutput.n172 1.12536
R1989 CSoutput.n265 CSoutput.n173 1.12536
R1990 CSoutput.n265 CSoutput.n175 1.12536
R1991 CSoutput.n255 CSoutput.n205 1.12536
R1992 CSoutput.n235 CSoutput.n205 1.12536
R1993 CSoutput.n237 CSoutput.n205 1.12536
R1994 CSoutput.n275 CSoutput.n138 1.12536
R1995 CSoutput.n275 CSoutput.n139 1.12536
R1996 CSoutput.n275 CSoutput.n141 1.12536
R1997 CSoutput.n31 CSoutput.n30 0.669944
R1998 CSoutput.n62 CSoutput.n61 0.669944
R1999 CSoutput.n348 CSoutput.n346 0.573776
R2000 CSoutput.n350 CSoutput.n348 0.573776
R2001 CSoutput.n352 CSoutput.n350 0.573776
R2002 CSoutput.n354 CSoutput.n352 0.573776
R2003 CSoutput.n356 CSoutput.n354 0.573776
R2004 CSoutput.n358 CSoutput.n356 0.573776
R2005 CSoutput.n360 CSoutput.n358 0.573776
R2006 CSoutput.n362 CSoutput.n360 0.573776
R2007 CSoutput.n329 CSoutput.n327 0.573776
R2008 CSoutput.n331 CSoutput.n329 0.573776
R2009 CSoutput.n333 CSoutput.n331 0.573776
R2010 CSoutput.n335 CSoutput.n333 0.573776
R2011 CSoutput.n337 CSoutput.n335 0.573776
R2012 CSoutput.n339 CSoutput.n337 0.573776
R2013 CSoutput.n341 CSoutput.n339 0.573776
R2014 CSoutput.n343 CSoutput.n341 0.573776
R2015 CSoutput.n402 CSoutput.n400 0.573776
R2016 CSoutput.n400 CSoutput.n398 0.573776
R2017 CSoutput.n398 CSoutput.n396 0.573776
R2018 CSoutput.n396 CSoutput.n394 0.573776
R2019 CSoutput.n394 CSoutput.n392 0.573776
R2020 CSoutput.n392 CSoutput.n390 0.573776
R2021 CSoutput.n390 CSoutput.n388 0.573776
R2022 CSoutput.n388 CSoutput.n386 0.573776
R2023 CSoutput.n383 CSoutput.n381 0.573776
R2024 CSoutput.n381 CSoutput.n379 0.573776
R2025 CSoutput.n379 CSoutput.n377 0.573776
R2026 CSoutput.n377 CSoutput.n375 0.573776
R2027 CSoutput.n375 CSoutput.n373 0.573776
R2028 CSoutput.n373 CSoutput.n371 0.573776
R2029 CSoutput.n371 CSoutput.n369 0.573776
R2030 CSoutput.n369 CSoutput.n367 0.573776
R2031 CSoutput.n405 CSoutput.n276 0.53442
R2032 CSoutput.n312 CSoutput.n310 0.358259
R2033 CSoutput.n314 CSoutput.n312 0.358259
R2034 CSoutput.n316 CSoutput.n314 0.358259
R2035 CSoutput.n318 CSoutput.n316 0.358259
R2036 CSoutput.n320 CSoutput.n318 0.358259
R2037 CSoutput.n322 CSoutput.n320 0.358259
R2038 CSoutput.n296 CSoutput.n294 0.358259
R2039 CSoutput.n298 CSoutput.n296 0.358259
R2040 CSoutput.n300 CSoutput.n298 0.358259
R2041 CSoutput.n302 CSoutput.n300 0.358259
R2042 CSoutput.n304 CSoutput.n302 0.358259
R2043 CSoutput.n306 CSoutput.n304 0.358259
R2044 CSoutput.n281 CSoutput.n279 0.358259
R2045 CSoutput.n283 CSoutput.n281 0.358259
R2046 CSoutput.n285 CSoutput.n283 0.358259
R2047 CSoutput.n287 CSoutput.n285 0.358259
R2048 CSoutput.n289 CSoutput.n287 0.358259
R2049 CSoutput.n291 CSoutput.n289 0.358259
R2050 CSoutput.n124 CSoutput.n122 0.358259
R2051 CSoutput.n122 CSoutput.n120 0.358259
R2052 CSoutput.n120 CSoutput.n118 0.358259
R2053 CSoutput.n118 CSoutput.n116 0.358259
R2054 CSoutput.n116 CSoutput.n114 0.358259
R2055 CSoutput.n114 CSoutput.n112 0.358259
R2056 CSoutput.n108 CSoutput.n106 0.358259
R2057 CSoutput.n106 CSoutput.n104 0.358259
R2058 CSoutput.n104 CSoutput.n102 0.358259
R2059 CSoutput.n102 CSoutput.n100 0.358259
R2060 CSoutput.n100 CSoutput.n98 0.358259
R2061 CSoutput.n98 CSoutput.n96 0.358259
R2062 CSoutput.n93 CSoutput.n91 0.358259
R2063 CSoutput.n91 CSoutput.n89 0.358259
R2064 CSoutput.n89 CSoutput.n87 0.358259
R2065 CSoutput.n87 CSoutput.n85 0.358259
R2066 CSoutput.n85 CSoutput.n83 0.358259
R2067 CSoutput.n83 CSoutput.n81 0.358259
R2068 CSoutput.n21 CSoutput.n20 0.169105
R2069 CSoutput.n21 CSoutput.n16 0.169105
R2070 CSoutput.n26 CSoutput.n16 0.169105
R2071 CSoutput.n27 CSoutput.n26 0.169105
R2072 CSoutput.n27 CSoutput.n14 0.169105
R2073 CSoutput.n32 CSoutput.n14 0.169105
R2074 CSoutput.n33 CSoutput.n32 0.169105
R2075 CSoutput.n34 CSoutput.n33 0.169105
R2076 CSoutput.n34 CSoutput.n12 0.169105
R2077 CSoutput.n39 CSoutput.n12 0.169105
R2078 CSoutput.n40 CSoutput.n39 0.169105
R2079 CSoutput.n40 CSoutput.n10 0.169105
R2080 CSoutput.n45 CSoutput.n10 0.169105
R2081 CSoutput.n46 CSoutput.n45 0.169105
R2082 CSoutput.n47 CSoutput.n46 0.169105
R2083 CSoutput.n47 CSoutput.n8 0.169105
R2084 CSoutput.n52 CSoutput.n8 0.169105
R2085 CSoutput.n53 CSoutput.n52 0.169105
R2086 CSoutput.n53 CSoutput.n6 0.169105
R2087 CSoutput.n58 CSoutput.n6 0.169105
R2088 CSoutput.n59 CSoutput.n58 0.169105
R2089 CSoutput.n60 CSoutput.n59 0.169105
R2090 CSoutput.n60 CSoutput.n4 0.169105
R2091 CSoutput.n66 CSoutput.n4 0.169105
R2092 CSoutput.n67 CSoutput.n66 0.169105
R2093 CSoutput.n68 CSoutput.n67 0.169105
R2094 CSoutput.n68 CSoutput.n2 0.169105
R2095 CSoutput.n73 CSoutput.n2 0.169105
R2096 CSoutput.n74 CSoutput.n73 0.169105
R2097 CSoutput.n74 CSoutput.n0 0.169105
R2098 CSoutput.n78 CSoutput.n0 0.169105
R2099 CSoutput.n219 CSoutput.n218 0.0910737
R2100 CSoutput.n270 CSoutput.n267 0.0723685
R2101 CSoutput.n224 CSoutput.n219 0.0522944
R2102 CSoutput.n267 CSoutput.n266 0.0499135
R2103 CSoutput.n218 CSoutput.n217 0.0499135
R2104 CSoutput.n252 CSoutput.n251 0.0464294
R2105 CSoutput.n260 CSoutput.n257 0.0391444
R2106 CSoutput.n219 CSoutput.t176 0.023435
R2107 CSoutput.n267 CSoutput.t180 0.02262
R2108 CSoutput.n218 CSoutput.t183 0.02262
R2109 CSoutput CSoutput.n405 0.0052
R2110 CSoutput.n189 CSoutput.n172 0.00365111
R2111 CSoutput.n192 CSoutput.n173 0.00365111
R2112 CSoutput.n175 CSoutput.n174 0.00365111
R2113 CSoutput.n217 CSoutput.n176 0.00365111
R2114 CSoutput.n181 CSoutput.n177 0.00365111
R2115 CSoutput.n264 CSoutput.n178 0.00365111
R2116 CSoutput.n255 CSoutput.n254 0.00365111
R2117 CSoutput.n235 CSoutput.n208 0.00365111
R2118 CSoutput.n237 CSoutput.n207 0.00365111
R2119 CSoutput.n225 CSoutput.n224 0.00365111
R2120 CSoutput.n231 CSoutput.n211 0.00365111
R2121 CSoutput.n233 CSoutput.n210 0.00365111
R2122 CSoutput.n155 CSoutput.n138 0.00365111
R2123 CSoutput.n158 CSoutput.n139 0.00365111
R2124 CSoutput.n141 CSoutput.n140 0.00365111
R2125 CSoutput.n251 CSoutput.n142 0.00365111
R2126 CSoutput.n147 CSoutput.n143 0.00365111
R2127 CSoutput.n274 CSoutput.n144 0.00365111
R2128 CSoutput.n186 CSoutput.n176 0.00340054
R2129 CSoutput.n179 CSoutput.n177 0.00340054
R2130 CSoutput.n264 CSoutput.n263 0.00340054
R2131 CSoutput.n259 CSoutput.n172 0.00340054
R2132 CSoutput.n188 CSoutput.n173 0.00340054
R2133 CSoutput.n191 CSoutput.n175 0.00340054
R2134 CSoutput.n230 CSoutput.n225 0.00340054
R2135 CSoutput.n232 CSoutput.n231 0.00340054
R2136 CSoutput.n234 CSoutput.n233 0.00340054
R2137 CSoutput.n256 CSoutput.n255 0.00340054
R2138 CSoutput.n236 CSoutput.n235 0.00340054
R2139 CSoutput.n238 CSoutput.n237 0.00340054
R2140 CSoutput.n152 CSoutput.n142 0.00340054
R2141 CSoutput.n145 CSoutput.n143 0.00340054
R2142 CSoutput.n274 CSoutput.n273 0.00340054
R2143 CSoutput.n269 CSoutput.n138 0.00340054
R2144 CSoutput.n154 CSoutput.n139 0.00340054
R2145 CSoutput.n157 CSoutput.n141 0.00340054
R2146 CSoutput.n187 CSoutput.n181 0.00252698
R2147 CSoutput.n180 CSoutput.n178 0.00252698
R2148 CSoutput.n262 CSoutput.n261 0.00252698
R2149 CSoutput.n190 CSoutput.n188 0.00252698
R2150 CSoutput.n193 CSoutput.n191 0.00252698
R2151 CSoutput.n266 CSoutput.n161 0.00252698
R2152 CSoutput.n187 CSoutput.n186 0.00252698
R2153 CSoutput.n180 CSoutput.n179 0.00252698
R2154 CSoutput.n263 CSoutput.n262 0.00252698
R2155 CSoutput.n190 CSoutput.n189 0.00252698
R2156 CSoutput.n193 CSoutput.n192 0.00252698
R2157 CSoutput.n174 CSoutput.n161 0.00252698
R2158 CSoutput.n241 CSoutput.n211 0.00252698
R2159 CSoutput.n240 CSoutput.n210 0.00252698
R2160 CSoutput.n239 CSoutput.n195 0.00252698
R2161 CSoutput.n236 CSoutput.n206 0.00252698
R2162 CSoutput.n243 CSoutput.n238 0.00252698
R2163 CSoutput.n252 CSoutput.n245 0.00252698
R2164 CSoutput.n241 CSoutput.n230 0.00252698
R2165 CSoutput.n240 CSoutput.n232 0.00252698
R2166 CSoutput.n239 CSoutput.n234 0.00252698
R2167 CSoutput.n254 CSoutput.n206 0.00252698
R2168 CSoutput.n243 CSoutput.n208 0.00252698
R2169 CSoutput.n245 CSoutput.n207 0.00252698
R2170 CSoutput.n153 CSoutput.n147 0.00252698
R2171 CSoutput.n146 CSoutput.n144 0.00252698
R2172 CSoutput.n272 CSoutput.n271 0.00252698
R2173 CSoutput.n156 CSoutput.n154 0.00252698
R2174 CSoutput.n159 CSoutput.n157 0.00252698
R2175 CSoutput.n276 CSoutput.n127 0.00252698
R2176 CSoutput.n153 CSoutput.n152 0.00252698
R2177 CSoutput.n146 CSoutput.n145 0.00252698
R2178 CSoutput.n273 CSoutput.n272 0.00252698
R2179 CSoutput.n156 CSoutput.n155 0.00252698
R2180 CSoutput.n159 CSoutput.n158 0.00252698
R2181 CSoutput.n140 CSoutput.n127 0.00252698
R2182 CSoutput.n261 CSoutput.n260 0.0020275
R2183 CSoutput.n260 CSoutput.n259 0.0020275
R2184 CSoutput.n257 CSoutput.n195 0.0020275
R2185 CSoutput.n257 CSoutput.n256 0.0020275
R2186 CSoutput.n271 CSoutput.n270 0.0020275
R2187 CSoutput.n270 CSoutput.n269 0.0020275
R2188 CSoutput.n171 CSoutput.n170 0.00166668
R2189 CSoutput.n253 CSoutput.n209 0.00166668
R2190 CSoutput.n137 CSoutput.n136 0.00166668
R2191 CSoutput.n275 CSoutput.n137 0.00133328
R2192 CSoutput.n209 CSoutput.n205 0.00133328
R2193 CSoutput.n265 CSoutput.n171 0.00133328
R2194 CSoutput.n268 CSoutput.n160 0.001
R2195 CSoutput.n246 CSoutput.n160 0.001
R2196 CSoutput.n148 CSoutput.n128 0.001
R2197 CSoutput.n247 CSoutput.n128 0.001
R2198 CSoutput.n149 CSoutput.n129 0.001
R2199 CSoutput.n248 CSoutput.n129 0.001
R2200 CSoutput.n150 CSoutput.n130 0.001
R2201 CSoutput.n249 CSoutput.n130 0.001
R2202 CSoutput.n151 CSoutput.n131 0.001
R2203 CSoutput.n250 CSoutput.n131 0.001
R2204 CSoutput.n244 CSoutput.n196 0.001
R2205 CSoutput.n244 CSoutput.n242 0.001
R2206 CSoutput.n226 CSoutput.n197 0.001
R2207 CSoutput.n220 CSoutput.n197 0.001
R2208 CSoutput.n227 CSoutput.n198 0.001
R2209 CSoutput.n221 CSoutput.n198 0.001
R2210 CSoutput.n228 CSoutput.n199 0.001
R2211 CSoutput.n222 CSoutput.n199 0.001
R2212 CSoutput.n229 CSoutput.n200 0.001
R2213 CSoutput.n223 CSoutput.n200 0.001
R2214 CSoutput.n258 CSoutput.n194 0.001
R2215 CSoutput.n212 CSoutput.n194 0.001
R2216 CSoutput.n182 CSoutput.n162 0.001
R2217 CSoutput.n213 CSoutput.n162 0.001
R2218 CSoutput.n183 CSoutput.n163 0.001
R2219 CSoutput.n214 CSoutput.n163 0.001
R2220 CSoutput.n184 CSoutput.n164 0.001
R2221 CSoutput.n215 CSoutput.n164 0.001
R2222 CSoutput.n185 CSoutput.n165 0.001
R2223 CSoutput.n216 CSoutput.n165 0.001
R2224 CSoutput.n216 CSoutput.n166 0.001
R2225 CSoutput.n215 CSoutput.n167 0.001
R2226 CSoutput.n214 CSoutput.n168 0.001
R2227 CSoutput.n213 CSoutput.t196 0.001
R2228 CSoutput.n212 CSoutput.n169 0.001
R2229 CSoutput.n185 CSoutput.n167 0.001
R2230 CSoutput.n184 CSoutput.n168 0.001
R2231 CSoutput.n183 CSoutput.t196 0.001
R2232 CSoutput.n182 CSoutput.n169 0.001
R2233 CSoutput.n258 CSoutput.n170 0.001
R2234 CSoutput.n223 CSoutput.n201 0.001
R2235 CSoutput.n222 CSoutput.n202 0.001
R2236 CSoutput.n221 CSoutput.n203 0.001
R2237 CSoutput.n220 CSoutput.t190 0.001
R2238 CSoutput.n242 CSoutput.n204 0.001
R2239 CSoutput.n229 CSoutput.n202 0.001
R2240 CSoutput.n228 CSoutput.n203 0.001
R2241 CSoutput.n227 CSoutput.t190 0.001
R2242 CSoutput.n226 CSoutput.n204 0.001
R2243 CSoutput.n253 CSoutput.n196 0.001
R2244 CSoutput.n250 CSoutput.n132 0.001
R2245 CSoutput.n249 CSoutput.n133 0.001
R2246 CSoutput.n248 CSoutput.n134 0.001
R2247 CSoutput.n247 CSoutput.t187 0.001
R2248 CSoutput.n246 CSoutput.n135 0.001
R2249 CSoutput.n151 CSoutput.n133 0.001
R2250 CSoutput.n150 CSoutput.n134 0.001
R2251 CSoutput.n149 CSoutput.t187 0.001
R2252 CSoutput.n148 CSoutput.n135 0.001
R2253 CSoutput.n268 CSoutput.n136 0.001
R2254 gnd.n2241 gnd.n2240 978.75
R2255 gnd.n4168 gnd.n4167 939.716
R2256 gnd.n5094 gnd.n5093 771.183
R2257 gnd.n6094 gnd.n6093 771.183
R2258 gnd.n6335 gnd.n935 771.183
R2259 gnd.n6675 gnd.n632 771.183
R2260 gnd.n4075 gnd.n1401 766.379
R2261 gnd.n4078 gnd.n4077 766.379
R2262 gnd.n3380 gnd.n3283 766.379
R2263 gnd.n3376 gnd.n3281 766.379
R2264 gnd.n4166 gnd.n1423 756.769
R2265 gnd.n2775 gnd.n2774 756.769
R2266 gnd.n3473 gnd.n3190 756.769
R2267 gnd.n3471 gnd.n3193 756.769
R2268 gnd.n7277 gnd.n125 751.963
R2269 gnd.n7435 gnd.n7434 751.963
R2270 gnd.n6833 gnd.n517 751.963
R2271 gnd.n5956 gnd.n479 751.963
R2272 gnd.n4998 gnd.n985 751.963
R2273 gnd.n6304 gnd.n6303 751.963
R2274 gnd.n4235 gnd.n4170 751.963
R2275 gnd.n4483 gnd.n1399 751.963
R2276 gnd.n7432 gnd.n127 732.745
R2277 gnd.n195 gnd.n123 732.745
R2278 gnd.n6836 gnd.n6835 732.745
R2279 gnd.n6908 gnd.n484 732.745
R2280 gnd.n6301 gnd.n987 732.745
R2281 gnd.n6232 gnd.n983 732.745
R2282 gnd.n4402 gnd.n4169 732.745
R2283 gnd.n4481 gnd.n4285 732.745
R2284 gnd.n2552 gnd.n1600 723.135
R2285 gnd.n2242 gnd.n1908 723.135
R2286 gnd.n7080 gnd.n343 723.135
R2287 gnd.n1476 gnd.n1210 723.135
R2288 gnd.n1600 gnd.n1599 585
R2289 gnd.n2554 gnd.n1600 585
R2290 gnd.n2557 gnd.n2556 585
R2291 gnd.n2556 gnd.n2555 585
R2292 gnd.n1597 gnd.n1596 585
R2293 gnd.n1596 gnd.n1595 585
R2294 gnd.n2562 gnd.n2561 585
R2295 gnd.n2563 gnd.n2562 585
R2296 gnd.n1594 gnd.n1593 585
R2297 gnd.n2564 gnd.n1594 585
R2298 gnd.n2567 gnd.n2566 585
R2299 gnd.n2566 gnd.n2565 585
R2300 gnd.n1591 gnd.n1590 585
R2301 gnd.n1590 gnd.n1589 585
R2302 gnd.n2572 gnd.n2571 585
R2303 gnd.n2573 gnd.n2572 585
R2304 gnd.n1588 gnd.n1587 585
R2305 gnd.n2574 gnd.n1588 585
R2306 gnd.n2577 gnd.n2576 585
R2307 gnd.n2576 gnd.n2575 585
R2308 gnd.n1585 gnd.n1584 585
R2309 gnd.n1584 gnd.n1583 585
R2310 gnd.n2582 gnd.n2581 585
R2311 gnd.n2583 gnd.n2582 585
R2312 gnd.n1582 gnd.n1581 585
R2313 gnd.n2584 gnd.n1582 585
R2314 gnd.n2587 gnd.n2586 585
R2315 gnd.n2586 gnd.n2585 585
R2316 gnd.n1579 gnd.n1578 585
R2317 gnd.n1578 gnd.n1577 585
R2318 gnd.n2592 gnd.n2591 585
R2319 gnd.n2593 gnd.n2592 585
R2320 gnd.n1576 gnd.n1575 585
R2321 gnd.n2594 gnd.n1576 585
R2322 gnd.n2597 gnd.n2596 585
R2323 gnd.n2596 gnd.n2595 585
R2324 gnd.n1573 gnd.n1572 585
R2325 gnd.n1572 gnd.n1571 585
R2326 gnd.n2602 gnd.n2601 585
R2327 gnd.n2603 gnd.n2602 585
R2328 gnd.n1570 gnd.n1569 585
R2329 gnd.n2604 gnd.n1570 585
R2330 gnd.n2607 gnd.n2606 585
R2331 gnd.n2606 gnd.n2605 585
R2332 gnd.n1567 gnd.n1566 585
R2333 gnd.n1566 gnd.n1565 585
R2334 gnd.n2612 gnd.n2611 585
R2335 gnd.n2613 gnd.n2612 585
R2336 gnd.n1564 gnd.n1563 585
R2337 gnd.n2614 gnd.n1564 585
R2338 gnd.n2617 gnd.n2616 585
R2339 gnd.n2616 gnd.n2615 585
R2340 gnd.n1561 gnd.n1560 585
R2341 gnd.n1560 gnd.n1559 585
R2342 gnd.n2622 gnd.n2621 585
R2343 gnd.n2623 gnd.n2622 585
R2344 gnd.n1558 gnd.n1557 585
R2345 gnd.n2624 gnd.n1558 585
R2346 gnd.n2627 gnd.n2626 585
R2347 gnd.n2626 gnd.n2625 585
R2348 gnd.n1555 gnd.n1554 585
R2349 gnd.n1554 gnd.n1553 585
R2350 gnd.n2632 gnd.n2631 585
R2351 gnd.n2633 gnd.n2632 585
R2352 gnd.n1552 gnd.n1551 585
R2353 gnd.n2634 gnd.n1552 585
R2354 gnd.n2637 gnd.n2636 585
R2355 gnd.n2636 gnd.n2635 585
R2356 gnd.n1549 gnd.n1548 585
R2357 gnd.n1548 gnd.n1547 585
R2358 gnd.n2642 gnd.n2641 585
R2359 gnd.n2643 gnd.n2642 585
R2360 gnd.n1546 gnd.n1545 585
R2361 gnd.n2644 gnd.n1546 585
R2362 gnd.n2647 gnd.n2646 585
R2363 gnd.n2646 gnd.n2645 585
R2364 gnd.n1543 gnd.n1542 585
R2365 gnd.n1542 gnd.n1541 585
R2366 gnd.n2652 gnd.n2651 585
R2367 gnd.n2653 gnd.n2652 585
R2368 gnd.n1540 gnd.n1539 585
R2369 gnd.n2654 gnd.n1540 585
R2370 gnd.n2657 gnd.n2656 585
R2371 gnd.n2656 gnd.n2655 585
R2372 gnd.n1537 gnd.n1536 585
R2373 gnd.n1536 gnd.n1535 585
R2374 gnd.n2662 gnd.n2661 585
R2375 gnd.n2663 gnd.n2662 585
R2376 gnd.n1534 gnd.n1533 585
R2377 gnd.n2664 gnd.n1534 585
R2378 gnd.n2667 gnd.n2666 585
R2379 gnd.n2666 gnd.n2665 585
R2380 gnd.n1531 gnd.n1530 585
R2381 gnd.n1530 gnd.n1529 585
R2382 gnd.n2672 gnd.n2671 585
R2383 gnd.n2673 gnd.n2672 585
R2384 gnd.n1528 gnd.n1527 585
R2385 gnd.n2674 gnd.n1528 585
R2386 gnd.n2677 gnd.n2676 585
R2387 gnd.n2676 gnd.n2675 585
R2388 gnd.n1525 gnd.n1524 585
R2389 gnd.n1524 gnd.n1523 585
R2390 gnd.n2682 gnd.n2681 585
R2391 gnd.n2683 gnd.n2682 585
R2392 gnd.n1522 gnd.n1521 585
R2393 gnd.n2684 gnd.n1522 585
R2394 gnd.n2687 gnd.n2686 585
R2395 gnd.n2686 gnd.n2685 585
R2396 gnd.n1519 gnd.n1518 585
R2397 gnd.n1518 gnd.n1517 585
R2398 gnd.n2692 gnd.n2691 585
R2399 gnd.n2693 gnd.n2692 585
R2400 gnd.n1516 gnd.n1515 585
R2401 gnd.n2694 gnd.n1516 585
R2402 gnd.n2697 gnd.n2696 585
R2403 gnd.n2696 gnd.n2695 585
R2404 gnd.n1513 gnd.n1512 585
R2405 gnd.n1512 gnd.n1511 585
R2406 gnd.n2702 gnd.n2701 585
R2407 gnd.n2703 gnd.n2702 585
R2408 gnd.n1510 gnd.n1509 585
R2409 gnd.n2704 gnd.n1510 585
R2410 gnd.n2707 gnd.n2706 585
R2411 gnd.n2706 gnd.n2705 585
R2412 gnd.n1507 gnd.n1506 585
R2413 gnd.n1506 gnd.n1505 585
R2414 gnd.n2712 gnd.n2711 585
R2415 gnd.n2713 gnd.n2712 585
R2416 gnd.n1504 gnd.n1503 585
R2417 gnd.n2714 gnd.n1504 585
R2418 gnd.n2717 gnd.n2716 585
R2419 gnd.n2716 gnd.n2715 585
R2420 gnd.n1501 gnd.n1500 585
R2421 gnd.n1500 gnd.n1499 585
R2422 gnd.n2722 gnd.n2721 585
R2423 gnd.n2723 gnd.n2722 585
R2424 gnd.n1498 gnd.n1497 585
R2425 gnd.n2724 gnd.n1498 585
R2426 gnd.n2727 gnd.n2726 585
R2427 gnd.n2726 gnd.n2725 585
R2428 gnd.n1495 gnd.n1494 585
R2429 gnd.n1494 gnd.n1493 585
R2430 gnd.n2732 gnd.n2731 585
R2431 gnd.n2733 gnd.n2732 585
R2432 gnd.n1492 gnd.n1491 585
R2433 gnd.n2734 gnd.n1492 585
R2434 gnd.n2737 gnd.n2736 585
R2435 gnd.n2736 gnd.n2735 585
R2436 gnd.n1489 gnd.n1488 585
R2437 gnd.n1488 gnd.n1487 585
R2438 gnd.n2742 gnd.n2741 585
R2439 gnd.n2743 gnd.n2742 585
R2440 gnd.n1486 gnd.n1485 585
R2441 gnd.n2744 gnd.n1486 585
R2442 gnd.n2747 gnd.n2746 585
R2443 gnd.n2746 gnd.n2745 585
R2444 gnd.n1483 gnd.n1482 585
R2445 gnd.n1482 gnd.n1481 585
R2446 gnd.n2752 gnd.n2751 585
R2447 gnd.n2753 gnd.n2752 585
R2448 gnd.n1480 gnd.n1479 585
R2449 gnd.n2754 gnd.n1480 585
R2450 gnd.n2757 gnd.n2756 585
R2451 gnd.n2756 gnd.n2755 585
R2452 gnd.n1477 gnd.n1475 585
R2453 gnd.n1475 gnd.n1474 585
R2454 gnd.n2765 gnd.n2764 585
R2455 gnd.n2766 gnd.n2765 585
R2456 gnd.n2552 gnd.n2551 585
R2457 gnd.n2553 gnd.n2552 585
R2458 gnd.n1603 gnd.n1602 585
R2459 gnd.n1602 gnd.n1601 585
R2460 gnd.n2547 gnd.n2546 585
R2461 gnd.n2546 gnd.n2545 585
R2462 gnd.n1606 gnd.n1605 585
R2463 gnd.n2544 gnd.n1606 585
R2464 gnd.n2542 gnd.n2541 585
R2465 gnd.n2543 gnd.n2542 585
R2466 gnd.n2540 gnd.n1608 585
R2467 gnd.n1608 gnd.n1607 585
R2468 gnd.n2539 gnd.n2538 585
R2469 gnd.n2538 gnd.n2537 585
R2470 gnd.n1613 gnd.n1612 585
R2471 gnd.n2536 gnd.n1613 585
R2472 gnd.n2534 gnd.n2533 585
R2473 gnd.n2535 gnd.n2534 585
R2474 gnd.n2532 gnd.n1615 585
R2475 gnd.n1615 gnd.n1614 585
R2476 gnd.n2531 gnd.n2530 585
R2477 gnd.n2530 gnd.n2529 585
R2478 gnd.n1621 gnd.n1620 585
R2479 gnd.n2528 gnd.n1621 585
R2480 gnd.n2526 gnd.n2525 585
R2481 gnd.n2527 gnd.n2526 585
R2482 gnd.n2524 gnd.n1623 585
R2483 gnd.n1623 gnd.n1622 585
R2484 gnd.n2523 gnd.n2522 585
R2485 gnd.n2522 gnd.n2521 585
R2486 gnd.n1629 gnd.n1628 585
R2487 gnd.n2520 gnd.n1629 585
R2488 gnd.n2518 gnd.n2517 585
R2489 gnd.n2519 gnd.n2518 585
R2490 gnd.n2516 gnd.n1631 585
R2491 gnd.n1631 gnd.n1630 585
R2492 gnd.n2515 gnd.n2514 585
R2493 gnd.n2514 gnd.n2513 585
R2494 gnd.n1637 gnd.n1636 585
R2495 gnd.n2512 gnd.n1637 585
R2496 gnd.n2510 gnd.n2509 585
R2497 gnd.n2511 gnd.n2510 585
R2498 gnd.n2508 gnd.n1639 585
R2499 gnd.n1639 gnd.n1638 585
R2500 gnd.n2507 gnd.n2506 585
R2501 gnd.n2506 gnd.n2505 585
R2502 gnd.n1645 gnd.n1644 585
R2503 gnd.n2504 gnd.n1645 585
R2504 gnd.n2502 gnd.n2501 585
R2505 gnd.n2503 gnd.n2502 585
R2506 gnd.n2500 gnd.n1647 585
R2507 gnd.n1647 gnd.n1646 585
R2508 gnd.n2499 gnd.n2498 585
R2509 gnd.n2498 gnd.n2497 585
R2510 gnd.n1653 gnd.n1652 585
R2511 gnd.n2496 gnd.n1653 585
R2512 gnd.n2494 gnd.n2493 585
R2513 gnd.n2495 gnd.n2494 585
R2514 gnd.n2492 gnd.n1655 585
R2515 gnd.n1655 gnd.n1654 585
R2516 gnd.n2491 gnd.n2490 585
R2517 gnd.n2490 gnd.n2489 585
R2518 gnd.n1661 gnd.n1660 585
R2519 gnd.n2488 gnd.n1661 585
R2520 gnd.n2486 gnd.n2485 585
R2521 gnd.n2487 gnd.n2486 585
R2522 gnd.n2484 gnd.n1663 585
R2523 gnd.n1663 gnd.n1662 585
R2524 gnd.n2483 gnd.n2482 585
R2525 gnd.n2482 gnd.n2481 585
R2526 gnd.n1669 gnd.n1668 585
R2527 gnd.n2480 gnd.n1669 585
R2528 gnd.n2478 gnd.n2477 585
R2529 gnd.n2479 gnd.n2478 585
R2530 gnd.n2476 gnd.n1671 585
R2531 gnd.n1671 gnd.n1670 585
R2532 gnd.n2475 gnd.n2474 585
R2533 gnd.n2474 gnd.n2473 585
R2534 gnd.n1677 gnd.n1676 585
R2535 gnd.n2472 gnd.n1677 585
R2536 gnd.n2470 gnd.n2469 585
R2537 gnd.n2471 gnd.n2470 585
R2538 gnd.n2468 gnd.n1679 585
R2539 gnd.n1679 gnd.n1678 585
R2540 gnd.n2467 gnd.n2466 585
R2541 gnd.n2466 gnd.n2465 585
R2542 gnd.n1685 gnd.n1684 585
R2543 gnd.n2464 gnd.n1685 585
R2544 gnd.n2462 gnd.n2461 585
R2545 gnd.n2463 gnd.n2462 585
R2546 gnd.n2460 gnd.n1687 585
R2547 gnd.n1687 gnd.n1686 585
R2548 gnd.n2459 gnd.n2458 585
R2549 gnd.n2458 gnd.n2457 585
R2550 gnd.n1693 gnd.n1692 585
R2551 gnd.n2456 gnd.n1693 585
R2552 gnd.n2454 gnd.n2453 585
R2553 gnd.n2455 gnd.n2454 585
R2554 gnd.n2452 gnd.n1695 585
R2555 gnd.n1695 gnd.n1694 585
R2556 gnd.n2451 gnd.n2450 585
R2557 gnd.n2450 gnd.n2449 585
R2558 gnd.n1701 gnd.n1700 585
R2559 gnd.n2448 gnd.n1701 585
R2560 gnd.n2446 gnd.n2445 585
R2561 gnd.n2447 gnd.n2446 585
R2562 gnd.n2444 gnd.n1703 585
R2563 gnd.n1703 gnd.n1702 585
R2564 gnd.n2443 gnd.n2442 585
R2565 gnd.n2442 gnd.n2441 585
R2566 gnd.n1709 gnd.n1708 585
R2567 gnd.n2440 gnd.n1709 585
R2568 gnd.n2438 gnd.n2437 585
R2569 gnd.n2439 gnd.n2438 585
R2570 gnd.n2436 gnd.n1711 585
R2571 gnd.n1711 gnd.n1710 585
R2572 gnd.n2435 gnd.n2434 585
R2573 gnd.n2434 gnd.n2433 585
R2574 gnd.n1717 gnd.n1716 585
R2575 gnd.n2432 gnd.n1717 585
R2576 gnd.n2430 gnd.n2429 585
R2577 gnd.n2431 gnd.n2430 585
R2578 gnd.n2428 gnd.n1719 585
R2579 gnd.n1719 gnd.n1718 585
R2580 gnd.n2427 gnd.n2426 585
R2581 gnd.n2426 gnd.n2425 585
R2582 gnd.n1725 gnd.n1724 585
R2583 gnd.n2424 gnd.n1725 585
R2584 gnd.n2422 gnd.n2421 585
R2585 gnd.n2423 gnd.n2422 585
R2586 gnd.n2420 gnd.n1727 585
R2587 gnd.n1727 gnd.n1726 585
R2588 gnd.n2419 gnd.n2418 585
R2589 gnd.n2418 gnd.n2417 585
R2590 gnd.n1733 gnd.n1732 585
R2591 gnd.n2416 gnd.n1733 585
R2592 gnd.n2414 gnd.n2413 585
R2593 gnd.n2415 gnd.n2414 585
R2594 gnd.n2412 gnd.n1735 585
R2595 gnd.n1735 gnd.n1734 585
R2596 gnd.n2411 gnd.n2410 585
R2597 gnd.n2410 gnd.n2409 585
R2598 gnd.n1741 gnd.n1740 585
R2599 gnd.n2408 gnd.n1741 585
R2600 gnd.n2406 gnd.n2405 585
R2601 gnd.n2407 gnd.n2406 585
R2602 gnd.n2404 gnd.n1743 585
R2603 gnd.n1743 gnd.n1742 585
R2604 gnd.n2403 gnd.n2402 585
R2605 gnd.n2402 gnd.n2401 585
R2606 gnd.n1749 gnd.n1748 585
R2607 gnd.n2400 gnd.n1749 585
R2608 gnd.n2398 gnd.n2397 585
R2609 gnd.n2399 gnd.n2398 585
R2610 gnd.n2396 gnd.n1751 585
R2611 gnd.n1751 gnd.n1750 585
R2612 gnd.n2395 gnd.n2394 585
R2613 gnd.n2394 gnd.n2393 585
R2614 gnd.n1757 gnd.n1756 585
R2615 gnd.n2392 gnd.n1757 585
R2616 gnd.n2390 gnd.n2389 585
R2617 gnd.n2391 gnd.n2390 585
R2618 gnd.n2388 gnd.n1759 585
R2619 gnd.n1759 gnd.n1758 585
R2620 gnd.n2387 gnd.n2386 585
R2621 gnd.n2386 gnd.n2385 585
R2622 gnd.n1765 gnd.n1764 585
R2623 gnd.n2384 gnd.n1765 585
R2624 gnd.n2382 gnd.n2381 585
R2625 gnd.n2383 gnd.n2382 585
R2626 gnd.n2380 gnd.n1767 585
R2627 gnd.n1767 gnd.n1766 585
R2628 gnd.n2379 gnd.n2378 585
R2629 gnd.n2378 gnd.n2377 585
R2630 gnd.n1773 gnd.n1772 585
R2631 gnd.n2376 gnd.n1773 585
R2632 gnd.n2374 gnd.n2373 585
R2633 gnd.n2375 gnd.n2374 585
R2634 gnd.n2372 gnd.n1775 585
R2635 gnd.n1775 gnd.n1774 585
R2636 gnd.n2371 gnd.n2370 585
R2637 gnd.n2370 gnd.n2369 585
R2638 gnd.n1781 gnd.n1780 585
R2639 gnd.n2368 gnd.n1781 585
R2640 gnd.n2366 gnd.n2365 585
R2641 gnd.n2367 gnd.n2366 585
R2642 gnd.n2364 gnd.n1783 585
R2643 gnd.n1783 gnd.n1782 585
R2644 gnd.n2363 gnd.n2362 585
R2645 gnd.n2362 gnd.n2361 585
R2646 gnd.n1789 gnd.n1788 585
R2647 gnd.n2360 gnd.n1789 585
R2648 gnd.n2358 gnd.n2357 585
R2649 gnd.n2359 gnd.n2358 585
R2650 gnd.n2356 gnd.n1791 585
R2651 gnd.n1791 gnd.n1790 585
R2652 gnd.n2355 gnd.n2354 585
R2653 gnd.n2354 gnd.n2353 585
R2654 gnd.n1797 gnd.n1796 585
R2655 gnd.n2352 gnd.n1797 585
R2656 gnd.n2350 gnd.n2349 585
R2657 gnd.n2351 gnd.n2350 585
R2658 gnd.n2348 gnd.n1799 585
R2659 gnd.n1799 gnd.n1798 585
R2660 gnd.n2347 gnd.n2346 585
R2661 gnd.n2346 gnd.n2345 585
R2662 gnd.n1805 gnd.n1804 585
R2663 gnd.n2344 gnd.n1805 585
R2664 gnd.n2342 gnd.n2341 585
R2665 gnd.n2343 gnd.n2342 585
R2666 gnd.n2340 gnd.n1807 585
R2667 gnd.n1807 gnd.n1806 585
R2668 gnd.n2339 gnd.n2338 585
R2669 gnd.n2338 gnd.n2337 585
R2670 gnd.n1813 gnd.n1812 585
R2671 gnd.n2336 gnd.n1813 585
R2672 gnd.n2334 gnd.n2333 585
R2673 gnd.n2335 gnd.n2334 585
R2674 gnd.n2332 gnd.n1815 585
R2675 gnd.n1815 gnd.n1814 585
R2676 gnd.n2331 gnd.n2330 585
R2677 gnd.n2330 gnd.n2329 585
R2678 gnd.n1821 gnd.n1820 585
R2679 gnd.n2328 gnd.n1821 585
R2680 gnd.n2326 gnd.n2325 585
R2681 gnd.n2327 gnd.n2326 585
R2682 gnd.n2324 gnd.n1823 585
R2683 gnd.n1823 gnd.n1822 585
R2684 gnd.n2323 gnd.n2322 585
R2685 gnd.n2322 gnd.n2321 585
R2686 gnd.n1829 gnd.n1828 585
R2687 gnd.n2320 gnd.n1829 585
R2688 gnd.n2318 gnd.n2317 585
R2689 gnd.n2319 gnd.n2318 585
R2690 gnd.n2316 gnd.n1831 585
R2691 gnd.n1831 gnd.n1830 585
R2692 gnd.n2315 gnd.n2314 585
R2693 gnd.n2314 gnd.n2313 585
R2694 gnd.n1837 gnd.n1836 585
R2695 gnd.n2312 gnd.n1837 585
R2696 gnd.n2310 gnd.n2309 585
R2697 gnd.n2311 gnd.n2310 585
R2698 gnd.n2308 gnd.n1839 585
R2699 gnd.n1839 gnd.n1838 585
R2700 gnd.n2307 gnd.n2306 585
R2701 gnd.n2306 gnd.n2305 585
R2702 gnd.n1845 gnd.n1844 585
R2703 gnd.n2304 gnd.n1845 585
R2704 gnd.n2302 gnd.n2301 585
R2705 gnd.n2303 gnd.n2302 585
R2706 gnd.n2300 gnd.n1847 585
R2707 gnd.n1847 gnd.n1846 585
R2708 gnd.n2299 gnd.n2298 585
R2709 gnd.n2298 gnd.n2297 585
R2710 gnd.n1853 gnd.n1852 585
R2711 gnd.n2296 gnd.n1853 585
R2712 gnd.n2294 gnd.n2293 585
R2713 gnd.n2295 gnd.n2294 585
R2714 gnd.n2292 gnd.n1855 585
R2715 gnd.n1855 gnd.n1854 585
R2716 gnd.n2291 gnd.n2290 585
R2717 gnd.n2290 gnd.n2289 585
R2718 gnd.n1861 gnd.n1860 585
R2719 gnd.n2288 gnd.n1861 585
R2720 gnd.n2286 gnd.n2285 585
R2721 gnd.n2287 gnd.n2286 585
R2722 gnd.n2284 gnd.n1863 585
R2723 gnd.n1863 gnd.n1862 585
R2724 gnd.n2283 gnd.n2282 585
R2725 gnd.n2282 gnd.n2281 585
R2726 gnd.n1869 gnd.n1868 585
R2727 gnd.n2280 gnd.n1869 585
R2728 gnd.n2278 gnd.n2277 585
R2729 gnd.n2279 gnd.n2278 585
R2730 gnd.n2276 gnd.n1871 585
R2731 gnd.n1871 gnd.n1870 585
R2732 gnd.n2275 gnd.n2274 585
R2733 gnd.n2274 gnd.n2273 585
R2734 gnd.n1877 gnd.n1876 585
R2735 gnd.n2272 gnd.n1877 585
R2736 gnd.n2270 gnd.n2269 585
R2737 gnd.n2271 gnd.n2270 585
R2738 gnd.n2268 gnd.n1879 585
R2739 gnd.n1879 gnd.n1878 585
R2740 gnd.n2267 gnd.n2266 585
R2741 gnd.n2266 gnd.n2265 585
R2742 gnd.n1885 gnd.n1884 585
R2743 gnd.n2264 gnd.n1885 585
R2744 gnd.n2262 gnd.n2261 585
R2745 gnd.n2263 gnd.n2262 585
R2746 gnd.n2260 gnd.n1887 585
R2747 gnd.n1887 gnd.n1886 585
R2748 gnd.n2259 gnd.n2258 585
R2749 gnd.n2258 gnd.n2257 585
R2750 gnd.n1893 gnd.n1892 585
R2751 gnd.n2256 gnd.n1893 585
R2752 gnd.n2254 gnd.n2253 585
R2753 gnd.n2255 gnd.n2254 585
R2754 gnd.n2252 gnd.n1895 585
R2755 gnd.n1895 gnd.n1894 585
R2756 gnd.n2251 gnd.n2250 585
R2757 gnd.n2250 gnd.n2249 585
R2758 gnd.n1901 gnd.n1900 585
R2759 gnd.n2248 gnd.n1901 585
R2760 gnd.n2246 gnd.n2245 585
R2761 gnd.n2247 gnd.n2246 585
R2762 gnd.n2244 gnd.n1903 585
R2763 gnd.n1903 gnd.n1902 585
R2764 gnd.n2243 gnd.n2242 585
R2765 gnd.n2242 gnd.n2241 585
R2766 gnd.n344 gnd.n342 585
R2767 gnd.n2068 gnd.n342 585
R2768 gnd.n2074 gnd.n2070 585
R2769 gnd.n2070 gnd.n2069 585
R2770 gnd.n2076 gnd.n2075 585
R2771 gnd.n2077 gnd.n2076 585
R2772 gnd.n2067 gnd.n2066 585
R2773 gnd.n2078 gnd.n2067 585
R2774 gnd.n2081 gnd.n2080 585
R2775 gnd.n2080 gnd.n2079 585
R2776 gnd.n2082 gnd.n2061 585
R2777 gnd.n2061 gnd.n2060 585
R2778 gnd.n2084 gnd.n2083 585
R2779 gnd.n2085 gnd.n2084 585
R2780 gnd.n2059 gnd.n2058 585
R2781 gnd.n2086 gnd.n2059 585
R2782 gnd.n2089 gnd.n2088 585
R2783 gnd.n2088 gnd.n2087 585
R2784 gnd.n2090 gnd.n2053 585
R2785 gnd.n2053 gnd.n2052 585
R2786 gnd.n2092 gnd.n2091 585
R2787 gnd.n2093 gnd.n2092 585
R2788 gnd.n2051 gnd.n2050 585
R2789 gnd.n2094 gnd.n2051 585
R2790 gnd.n2097 gnd.n2096 585
R2791 gnd.n2096 gnd.n2095 585
R2792 gnd.n2098 gnd.n2045 585
R2793 gnd.n2045 gnd.n2044 585
R2794 gnd.n2100 gnd.n2099 585
R2795 gnd.n2101 gnd.n2100 585
R2796 gnd.n2043 gnd.n2042 585
R2797 gnd.n2102 gnd.n2043 585
R2798 gnd.n2105 gnd.n2104 585
R2799 gnd.n2104 gnd.n2103 585
R2800 gnd.n2106 gnd.n2037 585
R2801 gnd.n2037 gnd.n2036 585
R2802 gnd.n2108 gnd.n2107 585
R2803 gnd.n2109 gnd.n2108 585
R2804 gnd.n2035 gnd.n2034 585
R2805 gnd.n2110 gnd.n2035 585
R2806 gnd.n2113 gnd.n2112 585
R2807 gnd.n2112 gnd.n2111 585
R2808 gnd.n2114 gnd.n2029 585
R2809 gnd.n2029 gnd.n2028 585
R2810 gnd.n2116 gnd.n2115 585
R2811 gnd.n2117 gnd.n2116 585
R2812 gnd.n2027 gnd.n2026 585
R2813 gnd.n2118 gnd.n2027 585
R2814 gnd.n2121 gnd.n2120 585
R2815 gnd.n2120 gnd.n2119 585
R2816 gnd.n2122 gnd.n2021 585
R2817 gnd.n2021 gnd.n2020 585
R2818 gnd.n2124 gnd.n2123 585
R2819 gnd.n2125 gnd.n2124 585
R2820 gnd.n2019 gnd.n2018 585
R2821 gnd.n2126 gnd.n2019 585
R2822 gnd.n2129 gnd.n2128 585
R2823 gnd.n2128 gnd.n2127 585
R2824 gnd.n2130 gnd.n2013 585
R2825 gnd.n2013 gnd.n2012 585
R2826 gnd.n2132 gnd.n2131 585
R2827 gnd.n2133 gnd.n2132 585
R2828 gnd.n2011 gnd.n2010 585
R2829 gnd.n2134 gnd.n2011 585
R2830 gnd.n2137 gnd.n2136 585
R2831 gnd.n2136 gnd.n2135 585
R2832 gnd.n2138 gnd.n2005 585
R2833 gnd.n2005 gnd.n2004 585
R2834 gnd.n2140 gnd.n2139 585
R2835 gnd.n2141 gnd.n2140 585
R2836 gnd.n2003 gnd.n2002 585
R2837 gnd.n2142 gnd.n2003 585
R2838 gnd.n2145 gnd.n2144 585
R2839 gnd.n2144 gnd.n2143 585
R2840 gnd.n2146 gnd.n1997 585
R2841 gnd.n1997 gnd.n1996 585
R2842 gnd.n2148 gnd.n2147 585
R2843 gnd.n2149 gnd.n2148 585
R2844 gnd.n1995 gnd.n1994 585
R2845 gnd.n2150 gnd.n1995 585
R2846 gnd.n2153 gnd.n2152 585
R2847 gnd.n2152 gnd.n2151 585
R2848 gnd.n2154 gnd.n1989 585
R2849 gnd.n1989 gnd.n1988 585
R2850 gnd.n2156 gnd.n2155 585
R2851 gnd.n2157 gnd.n2156 585
R2852 gnd.n1987 gnd.n1986 585
R2853 gnd.n2158 gnd.n1987 585
R2854 gnd.n2161 gnd.n2160 585
R2855 gnd.n2160 gnd.n2159 585
R2856 gnd.n2162 gnd.n1981 585
R2857 gnd.n1981 gnd.n1980 585
R2858 gnd.n2164 gnd.n2163 585
R2859 gnd.n2165 gnd.n2164 585
R2860 gnd.n1979 gnd.n1978 585
R2861 gnd.n2166 gnd.n1979 585
R2862 gnd.n2169 gnd.n2168 585
R2863 gnd.n2168 gnd.n2167 585
R2864 gnd.n2170 gnd.n1973 585
R2865 gnd.n1973 gnd.n1972 585
R2866 gnd.n2172 gnd.n2171 585
R2867 gnd.n2173 gnd.n2172 585
R2868 gnd.n1971 gnd.n1970 585
R2869 gnd.n2174 gnd.n1971 585
R2870 gnd.n2177 gnd.n2176 585
R2871 gnd.n2176 gnd.n2175 585
R2872 gnd.n2178 gnd.n1965 585
R2873 gnd.n1965 gnd.n1964 585
R2874 gnd.n2180 gnd.n2179 585
R2875 gnd.n2181 gnd.n2180 585
R2876 gnd.n1963 gnd.n1962 585
R2877 gnd.n2182 gnd.n1963 585
R2878 gnd.n2185 gnd.n2184 585
R2879 gnd.n2184 gnd.n2183 585
R2880 gnd.n2186 gnd.n1957 585
R2881 gnd.n1957 gnd.n1956 585
R2882 gnd.n2188 gnd.n2187 585
R2883 gnd.n2189 gnd.n2188 585
R2884 gnd.n1955 gnd.n1954 585
R2885 gnd.n2190 gnd.n1955 585
R2886 gnd.n2193 gnd.n2192 585
R2887 gnd.n2192 gnd.n2191 585
R2888 gnd.n2194 gnd.n1949 585
R2889 gnd.n1949 gnd.n1948 585
R2890 gnd.n2196 gnd.n2195 585
R2891 gnd.n2197 gnd.n2196 585
R2892 gnd.n1947 gnd.n1946 585
R2893 gnd.n2198 gnd.n1947 585
R2894 gnd.n2201 gnd.n2200 585
R2895 gnd.n2200 gnd.n2199 585
R2896 gnd.n2202 gnd.n1941 585
R2897 gnd.n1941 gnd.n1940 585
R2898 gnd.n2204 gnd.n2203 585
R2899 gnd.n2205 gnd.n2204 585
R2900 gnd.n1939 gnd.n1938 585
R2901 gnd.n2206 gnd.n1939 585
R2902 gnd.n2209 gnd.n2208 585
R2903 gnd.n2208 gnd.n2207 585
R2904 gnd.n2210 gnd.n1933 585
R2905 gnd.n1933 gnd.n1932 585
R2906 gnd.n2212 gnd.n2211 585
R2907 gnd.n2213 gnd.n2212 585
R2908 gnd.n1931 gnd.n1930 585
R2909 gnd.n2214 gnd.n1931 585
R2910 gnd.n2217 gnd.n2216 585
R2911 gnd.n2216 gnd.n2215 585
R2912 gnd.n2218 gnd.n1925 585
R2913 gnd.n1925 gnd.n1924 585
R2914 gnd.n2220 gnd.n2219 585
R2915 gnd.n2221 gnd.n2220 585
R2916 gnd.n1923 gnd.n1922 585
R2917 gnd.n2222 gnd.n1923 585
R2918 gnd.n2225 gnd.n2224 585
R2919 gnd.n2224 gnd.n2223 585
R2920 gnd.n2226 gnd.n1918 585
R2921 gnd.n1918 gnd.n1917 585
R2922 gnd.n2228 gnd.n2227 585
R2923 gnd.n2229 gnd.n2228 585
R2924 gnd.n1916 gnd.n1915 585
R2925 gnd.n2230 gnd.n1916 585
R2926 gnd.n2233 gnd.n2232 585
R2927 gnd.n2232 gnd.n2231 585
R2928 gnd.n1912 gnd.n1910 585
R2929 gnd.n1910 gnd.n1909 585
R2930 gnd.n2238 gnd.n2237 585
R2931 gnd.n2239 gnd.n2238 585
R2932 gnd.n1911 gnd.n1908 585
R2933 gnd.n2240 gnd.n1908 585
R2934 gnd.n6222 gnd.n985 585
R2935 gnd.n6302 gnd.n985 585
R2936 gnd.n6224 gnd.n6223 585
R2937 gnd.n6225 gnd.n6224 585
R2938 gnd.n1063 gnd.n1062 585
R2939 gnd.n4801 gnd.n1062 585
R2940 gnd.n4984 gnd.n4983 585
R2941 gnd.n4983 gnd.n4982 585
R2942 gnd.n1066 gnd.n1065 585
R2943 gnd.n4799 gnd.n1066 585
R2944 gnd.n4971 gnd.n4970 585
R2945 gnd.n4972 gnd.n4971 585
R2946 gnd.n1082 gnd.n1081 585
R2947 gnd.n4788 gnd.n1081 585
R2948 gnd.n4966 gnd.n4965 585
R2949 gnd.n4965 gnd.n4964 585
R2950 gnd.n1085 gnd.n1084 585
R2951 gnd.n4740 gnd.n1085 585
R2952 gnd.n4955 gnd.n4954 585
R2953 gnd.n4956 gnd.n4955 585
R2954 gnd.n1098 gnd.n1097 585
R2955 gnd.n4746 gnd.n1097 585
R2956 gnd.n4950 gnd.n4949 585
R2957 gnd.n4949 gnd.n4948 585
R2958 gnd.n1101 gnd.n1100 585
R2959 gnd.n4732 gnd.n1101 585
R2960 gnd.n4939 gnd.n4938 585
R2961 gnd.n4940 gnd.n4939 585
R2962 gnd.n1116 gnd.n1115 585
R2963 gnd.n4728 gnd.n1115 585
R2964 gnd.n4934 gnd.n4933 585
R2965 gnd.n4933 gnd.n4932 585
R2966 gnd.n1119 gnd.n1118 585
R2967 gnd.n4701 gnd.n1119 585
R2968 gnd.n4923 gnd.n4922 585
R2969 gnd.n4924 gnd.n4923 585
R2970 gnd.n1132 gnd.n1131 585
R2971 gnd.n4707 gnd.n1131 585
R2972 gnd.n4918 gnd.n4917 585
R2973 gnd.n4917 gnd.n4916 585
R2974 gnd.n1135 gnd.n1134 585
R2975 gnd.n4692 gnd.n1135 585
R2976 gnd.n4907 gnd.n4906 585
R2977 gnd.n4908 gnd.n4907 585
R2978 gnd.n1150 gnd.n1149 585
R2979 gnd.n4688 gnd.n1149 585
R2980 gnd.n4902 gnd.n4901 585
R2981 gnd.n4901 gnd.n4900 585
R2982 gnd.n1153 gnd.n1152 585
R2983 gnd.n4661 gnd.n1153 585
R2984 gnd.n4891 gnd.n4890 585
R2985 gnd.n4892 gnd.n4891 585
R2986 gnd.n1166 gnd.n1165 585
R2987 gnd.n4844 gnd.n1165 585
R2988 gnd.n4886 gnd.n4885 585
R2989 gnd.n4885 gnd.n4884 585
R2990 gnd.n1169 gnd.n1168 585
R2991 gnd.n4653 gnd.n1169 585
R2992 gnd.n4858 gnd.n4857 585
R2993 gnd.n4857 gnd.n4856 585
R2994 gnd.n4859 gnd.n1203 585
R2995 gnd.n4645 gnd.n1203 585
R2996 gnd.n4861 gnd.n4860 585
R2997 gnd.n4862 gnd.n4861 585
R2998 gnd.n1195 gnd.n1194 585
R2999 gnd.n1198 gnd.n1195 585
R3000 gnd.n4872 gnd.n4871 585
R3001 gnd.n4871 gnd.n4870 585
R3002 gnd.n4873 gnd.n1189 585
R3003 gnd.n1189 gnd.n1187 585
R3004 gnd.n4875 gnd.n4874 585
R3005 gnd.n4876 gnd.n4875 585
R3006 gnd.n1190 gnd.n1188 585
R3007 gnd.n4629 gnd.n1188 585
R3008 gnd.n1307 gnd.n1306 585
R3009 gnd.n1306 gnd.n1279 585
R3010 gnd.n1308 gnd.n1286 585
R3011 gnd.n4611 gnd.n1286 585
R3012 gnd.n4598 gnd.n4597 585
R3013 gnd.n4597 gnd.n4596 585
R3014 gnd.n4599 gnd.n1298 585
R3015 gnd.n1298 gnd.n1296 585
R3016 gnd.n4601 gnd.n4600 585
R3017 gnd.n4602 gnd.n4601 585
R3018 gnd.n1299 gnd.n1297 585
R3019 gnd.n4585 gnd.n1297 585
R3020 gnd.n4557 gnd.n4556 585
R3021 gnd.n4556 gnd.n1314 585
R3022 gnd.n4558 gnd.n1322 585
R3023 gnd.n4572 gnd.n1322 585
R3024 gnd.n4559 gnd.n1332 585
R3025 gnd.n1332 gnd.n1320 585
R3026 gnd.n4561 gnd.n4560 585
R3027 gnd.n4562 gnd.n4561 585
R3028 gnd.n1333 gnd.n1331 585
R3029 gnd.n1340 gnd.n1331 585
R3030 gnd.n4548 gnd.n4547 585
R3031 gnd.n4547 gnd.n4546 585
R3032 gnd.n1336 gnd.n1335 585
R3033 gnd.n1337 gnd.n1336 585
R3034 gnd.n4537 gnd.n4536 585
R3035 gnd.n4538 gnd.n4537 585
R3036 gnd.n1350 gnd.n1349 585
R3037 gnd.n1349 gnd.n1346 585
R3038 gnd.n4532 gnd.n4531 585
R3039 gnd.n4531 gnd.n4530 585
R3040 gnd.n1353 gnd.n1352 585
R3041 gnd.n1354 gnd.n1353 585
R3042 gnd.n4521 gnd.n4520 585
R3043 gnd.n4522 gnd.n4521 585
R3044 gnd.n1365 gnd.n1364 585
R3045 gnd.n1372 gnd.n1364 585
R3046 gnd.n4516 gnd.n4515 585
R3047 gnd.n4515 gnd.n4514 585
R3048 gnd.n1368 gnd.n1367 585
R3049 gnd.n1369 gnd.n1368 585
R3050 gnd.n4505 gnd.n4504 585
R3051 gnd.n4506 gnd.n4505 585
R3052 gnd.n1382 gnd.n1381 585
R3053 gnd.n1381 gnd.n1378 585
R3054 gnd.n4500 gnd.n4499 585
R3055 gnd.n4499 gnd.n4498 585
R3056 gnd.n1385 gnd.n1384 585
R3057 gnd.n1386 gnd.n1385 585
R3058 gnd.n4489 gnd.n4488 585
R3059 gnd.n4490 gnd.n4489 585
R3060 gnd.n1397 gnd.n1396 585
R3061 gnd.n4284 gnd.n1396 585
R3062 gnd.n4484 gnd.n4483 585
R3063 gnd.n4483 gnd.n4482 585
R3064 gnd.n4191 gnd.n1399 585
R3065 gnd.n4194 gnd.n4192 585
R3066 gnd.n4197 gnd.n4196 585
R3067 gnd.n4189 gnd.n4188 585
R3068 gnd.n4202 gnd.n4201 585
R3069 gnd.n4204 gnd.n4187 585
R3070 gnd.n4207 gnd.n4206 585
R3071 gnd.n4185 gnd.n4184 585
R3072 gnd.n4212 gnd.n4211 585
R3073 gnd.n4214 gnd.n4183 585
R3074 gnd.n4217 gnd.n4216 585
R3075 gnd.n4181 gnd.n4180 585
R3076 gnd.n4222 gnd.n4221 585
R3077 gnd.n4224 gnd.n4179 585
R3078 gnd.n4227 gnd.n4226 585
R3079 gnd.n4177 gnd.n4176 585
R3080 gnd.n4232 gnd.n4231 585
R3081 gnd.n4234 gnd.n4175 585
R3082 gnd.n4236 gnd.n4235 585
R3083 gnd.n4235 gnd.n4168 585
R3084 gnd.n6305 gnd.n6304 585
R3085 gnd.n5051 gnd.n978 585
R3086 gnd.n5055 gnd.n5052 585
R3087 gnd.n5056 gnd.n5049 585
R3088 gnd.n5048 gnd.n5039 585
R3089 gnd.n5063 gnd.n5038 585
R3090 gnd.n5064 gnd.n5037 585
R3091 gnd.n5035 gnd.n5029 585
R3092 gnd.n5071 gnd.n5028 585
R3093 gnd.n5072 gnd.n5026 585
R3094 gnd.n5025 gnd.n5016 585
R3095 gnd.n5079 gnd.n5015 585
R3096 gnd.n5080 gnd.n5014 585
R3097 gnd.n5012 gnd.n5006 585
R3098 gnd.n5087 gnd.n5005 585
R3099 gnd.n5088 gnd.n5003 585
R3100 gnd.n5002 gnd.n4997 585
R3101 gnd.n5000 gnd.n4999 585
R3102 gnd.n4998 gnd.n4988 585
R3103 gnd.n4998 gnd.n992 585
R3104 gnd.n6303 gnd.n981 585
R3105 gnd.n6303 gnd.n6302 585
R3106 gnd.n4803 gnd.n980 585
R3107 gnd.n6225 gnd.n980 585
R3108 gnd.n4806 gnd.n4802 585
R3109 gnd.n4802 gnd.n4801 585
R3110 gnd.n4807 gnd.n1069 585
R3111 gnd.n4982 gnd.n1069 585
R3112 gnd.n4808 gnd.n4800 585
R3113 gnd.n4800 gnd.n4799 585
R3114 gnd.n1241 gnd.n1079 585
R3115 gnd.n4972 gnd.n1079 585
R3116 gnd.n4812 gnd.n1240 585
R3117 gnd.n4788 gnd.n1240 585
R3118 gnd.n4813 gnd.n1088 585
R3119 gnd.n4964 gnd.n1088 585
R3120 gnd.n4814 gnd.n1239 585
R3121 gnd.n4740 gnd.n1239 585
R3122 gnd.n1237 gnd.n1095 585
R3123 gnd.n4956 gnd.n1095 585
R3124 gnd.n4818 gnd.n1236 585
R3125 gnd.n4746 gnd.n1236 585
R3126 gnd.n4819 gnd.n1104 585
R3127 gnd.n4948 gnd.n1104 585
R3128 gnd.n4820 gnd.n1235 585
R3129 gnd.n4732 gnd.n1235 585
R3130 gnd.n1233 gnd.n1113 585
R3131 gnd.n4940 gnd.n1113 585
R3132 gnd.n4824 gnd.n1232 585
R3133 gnd.n4728 gnd.n1232 585
R3134 gnd.n4825 gnd.n1122 585
R3135 gnd.n4932 gnd.n1122 585
R3136 gnd.n4826 gnd.n1231 585
R3137 gnd.n4701 gnd.n1231 585
R3138 gnd.n1229 gnd.n1129 585
R3139 gnd.n4924 gnd.n1129 585
R3140 gnd.n4830 gnd.n1228 585
R3141 gnd.n4707 gnd.n1228 585
R3142 gnd.n4831 gnd.n1138 585
R3143 gnd.n4916 gnd.n1138 585
R3144 gnd.n4832 gnd.n1227 585
R3145 gnd.n4692 gnd.n1227 585
R3146 gnd.n1225 gnd.n1147 585
R3147 gnd.n4908 gnd.n1147 585
R3148 gnd.n4836 gnd.n1224 585
R3149 gnd.n4688 gnd.n1224 585
R3150 gnd.n4837 gnd.n1156 585
R3151 gnd.n4900 gnd.n1156 585
R3152 gnd.n4838 gnd.n1223 585
R3153 gnd.n4661 gnd.n1223 585
R3154 gnd.n1220 gnd.n1163 585
R3155 gnd.n4892 gnd.n1163 585
R3156 gnd.n4843 gnd.n4842 585
R3157 gnd.n4844 gnd.n4843 585
R3158 gnd.n1219 gnd.n1172 585
R3159 gnd.n4884 gnd.n1172 585
R3160 gnd.n4652 gnd.n4651 585
R3161 gnd.n4653 gnd.n4652 585
R3162 gnd.n1269 gnd.n1209 585
R3163 gnd.n4856 gnd.n1209 585
R3164 gnd.n4647 gnd.n4646 585
R3165 gnd.n4646 gnd.n4645 585
R3166 gnd.n1271 gnd.n1202 585
R3167 gnd.n4862 gnd.n1202 585
R3168 gnd.n4622 gnd.n4620 585
R3169 gnd.n4620 gnd.n1198 585
R3170 gnd.n4623 gnd.n1197 585
R3171 gnd.n4870 gnd.n1197 585
R3172 gnd.n4625 gnd.n4624 585
R3173 gnd.n4624 gnd.n1187 585
R3174 gnd.n4626 gnd.n1186 585
R3175 gnd.n4876 gnd.n1186 585
R3176 gnd.n4628 gnd.n4627 585
R3177 gnd.n4629 gnd.n4628 585
R3178 gnd.n1281 gnd.n1280 585
R3179 gnd.n1280 gnd.n1279 585
R3180 gnd.n4613 gnd.n4612 585
R3181 gnd.n4612 gnd.n4611 585
R3182 gnd.n1284 gnd.n1283 585
R3183 gnd.n4596 gnd.n1284 585
R3184 gnd.n4581 gnd.n4580 585
R3185 gnd.n4580 gnd.n1296 585
R3186 gnd.n4582 gnd.n1295 585
R3187 gnd.n4602 gnd.n1295 585
R3188 gnd.n4584 gnd.n4583 585
R3189 gnd.n4585 gnd.n4584 585
R3190 gnd.n1316 gnd.n1315 585
R3191 gnd.n1315 gnd.n1314 585
R3192 gnd.n4574 gnd.n4573 585
R3193 gnd.n4573 gnd.n4572 585
R3194 gnd.n1319 gnd.n1318 585
R3195 gnd.n1320 gnd.n1319 585
R3196 gnd.n4257 gnd.n1330 585
R3197 gnd.n4562 gnd.n1330 585
R3198 gnd.n4259 gnd.n4258 585
R3199 gnd.n4258 gnd.n1340 585
R3200 gnd.n4260 gnd.n1339 585
R3201 gnd.n4546 gnd.n1339 585
R3202 gnd.n4262 gnd.n4261 585
R3203 gnd.n4261 gnd.n1337 585
R3204 gnd.n4263 gnd.n1348 585
R3205 gnd.n4538 gnd.n1348 585
R3206 gnd.n4265 gnd.n4264 585
R3207 gnd.n4264 gnd.n1346 585
R3208 gnd.n4266 gnd.n1356 585
R3209 gnd.n4530 gnd.n1356 585
R3210 gnd.n4268 gnd.n4267 585
R3211 gnd.n4267 gnd.n1354 585
R3212 gnd.n4269 gnd.n1363 585
R3213 gnd.n4522 gnd.n1363 585
R3214 gnd.n4271 gnd.n4270 585
R3215 gnd.n4270 gnd.n1372 585
R3216 gnd.n4272 gnd.n1371 585
R3217 gnd.n4514 gnd.n1371 585
R3218 gnd.n4274 gnd.n4273 585
R3219 gnd.n4273 gnd.n1369 585
R3220 gnd.n4275 gnd.n1380 585
R3221 gnd.n4506 gnd.n1380 585
R3222 gnd.n4277 gnd.n4276 585
R3223 gnd.n4276 gnd.n1378 585
R3224 gnd.n4278 gnd.n1388 585
R3225 gnd.n4498 gnd.n1388 585
R3226 gnd.n4280 gnd.n4279 585
R3227 gnd.n4279 gnd.n1386 585
R3228 gnd.n4281 gnd.n1395 585
R3229 gnd.n4490 gnd.n1395 585
R3230 gnd.n4283 gnd.n4282 585
R3231 gnd.n4284 gnd.n4283 585
R3232 gnd.n4171 gnd.n4170 585
R3233 gnd.n4482 gnd.n4170 585
R3234 gnd.n7337 gnd.n125 585
R3235 gnd.n7433 gnd.n125 585
R3236 gnd.n7338 gnd.n7275 585
R3237 gnd.n7275 gnd.n122 585
R3238 gnd.n7339 gnd.n203 585
R3239 gnd.n7353 gnd.n203 585
R3240 gnd.n215 gnd.n213 585
R3241 gnd.n213 gnd.n202 585
R3242 gnd.n7344 gnd.n7343 585
R3243 gnd.n7345 gnd.n7344 585
R3244 gnd.n214 gnd.n212 585
R3245 gnd.n212 gnd.n209 585
R3246 gnd.n7271 gnd.n7270 585
R3247 gnd.n7270 gnd.n7269 585
R3248 gnd.n218 gnd.n217 585
R3249 gnd.n228 gnd.n218 585
R3250 gnd.n7260 gnd.n7259 585
R3251 gnd.n7261 gnd.n7260 585
R3252 gnd.n230 gnd.n229 585
R3253 gnd.n229 gnd.n225 585
R3254 gnd.n7255 gnd.n7254 585
R3255 gnd.n7254 gnd.n7253 585
R3256 gnd.n233 gnd.n232 585
R3257 gnd.n234 gnd.n233 585
R3258 gnd.n7244 gnd.n7243 585
R3259 gnd.n7245 gnd.n7244 585
R3260 gnd.n245 gnd.n244 585
R3261 gnd.n250 gnd.n244 585
R3262 gnd.n7239 gnd.n7238 585
R3263 gnd.n7238 gnd.n7237 585
R3264 gnd.n248 gnd.n247 585
R3265 gnd.n259 gnd.n248 585
R3266 gnd.n7228 gnd.n7227 585
R3267 gnd.n7229 gnd.n7228 585
R3268 gnd.n261 gnd.n260 585
R3269 gnd.n260 gnd.n256 585
R3270 gnd.n7223 gnd.n7222 585
R3271 gnd.n7222 gnd.n7221 585
R3272 gnd.n264 gnd.n263 585
R3273 gnd.n265 gnd.n264 585
R3274 gnd.n7212 gnd.n7211 585
R3275 gnd.n7213 gnd.n7212 585
R3276 gnd.n275 gnd.n274 585
R3277 gnd.n280 gnd.n274 585
R3278 gnd.n7207 gnd.n7206 585
R3279 gnd.n7206 gnd.n7205 585
R3280 gnd.n278 gnd.n277 585
R3281 gnd.n289 gnd.n278 585
R3282 gnd.n7196 gnd.n7195 585
R3283 gnd.n7197 gnd.n7196 585
R3284 gnd.n291 gnd.n290 585
R3285 gnd.n290 gnd.n286 585
R3286 gnd.n7191 gnd.n7190 585
R3287 gnd.n7190 gnd.n7189 585
R3288 gnd.n294 gnd.n293 585
R3289 gnd.n295 gnd.n294 585
R3290 gnd.n7167 gnd.n7166 585
R3291 gnd.n7166 gnd.n7165 585
R3292 gnd.n7168 gnd.n323 585
R3293 gnd.n7161 gnd.n323 585
R3294 gnd.n329 gnd.n321 585
R3295 gnd.n330 gnd.n329 585
R3296 gnd.n7172 gnd.n320 585
R3297 gnd.n7088 gnd.n320 585
R3298 gnd.n7173 gnd.n319 585
R3299 gnd.n336 gnd.n319 585
R3300 gnd.n7174 gnd.n318 585
R3301 gnd.n7082 gnd.n318 585
R3302 gnd.n315 gnd.n313 585
R3303 gnd.n7062 gnd.n313 585
R3304 gnd.n7179 gnd.n7178 585
R3305 gnd.n7180 gnd.n7179 585
R3306 gnd.n314 gnd.n312 585
R3307 gnd.n7071 gnd.n312 585
R3308 gnd.n7033 gnd.n7031 585
R3309 gnd.n7031 gnd.n349 585
R3310 gnd.n7034 gnd.n362 585
R3311 gnd.n7050 gnd.n362 585
R3312 gnd.n7035 gnd.n7030 585
R3313 gnd.n7030 gnd.n7029 585
R3314 gnd.n376 gnd.n374 585
R3315 gnd.n6790 gnd.n374 585
R3316 gnd.n7040 gnd.n7039 585
R3317 gnd.n7041 gnd.n7040 585
R3318 gnd.n375 gnd.n373 585
R3319 gnd.n7019 gnd.n373 585
R3320 gnd.n6984 gnd.n395 585
R3321 gnd.n6998 gnd.n395 585
R3322 gnd.n408 gnd.n406 585
R3323 gnd.n6798 gnd.n406 585
R3324 gnd.n6989 gnd.n6988 585
R3325 gnd.n6990 gnd.n6989 585
R3326 gnd.n407 gnd.n405 585
R3327 gnd.n6777 gnd.n405 585
R3328 gnd.n6981 gnd.n6980 585
R3329 gnd.n6980 gnd.n6979 585
R3330 gnd.n411 gnd.n410 585
R3331 gnd.n6758 gnd.n411 585
R3332 gnd.n6970 gnd.n6969 585
R3333 gnd.n6971 gnd.n6970 585
R3334 gnd.n424 gnd.n423 585
R3335 gnd.n6764 gnd.n423 585
R3336 gnd.n6965 gnd.n6964 585
R3337 gnd.n6964 gnd.n6963 585
R3338 gnd.n427 gnd.n426 585
R3339 gnd.n6750 gnd.n427 585
R3340 gnd.n6954 gnd.n6953 585
R3341 gnd.n6955 gnd.n6954 585
R3342 gnd.n442 gnd.n441 585
R3343 gnd.n6746 gnd.n441 585
R3344 gnd.n6949 gnd.n6948 585
R3345 gnd.n6948 gnd.n6947 585
R3346 gnd.n445 gnd.n444 585
R3347 gnd.n6719 gnd.n445 585
R3348 gnd.n6938 gnd.n6937 585
R3349 gnd.n6939 gnd.n6938 585
R3350 gnd.n458 gnd.n457 585
R3351 gnd.n6725 gnd.n457 585
R3352 gnd.n6933 gnd.n6932 585
R3353 gnd.n6932 gnd.n6931 585
R3354 gnd.n461 gnd.n460 585
R3355 gnd.n6710 gnd.n461 585
R3356 gnd.n6922 gnd.n6921 585
R3357 gnd.n6923 gnd.n6922 585
R3358 gnd.n476 gnd.n475 585
R3359 gnd.n6706 gnd.n475 585
R3360 gnd.n6917 gnd.n6916 585
R3361 gnd.n6916 gnd.n6915 585
R3362 gnd.n479 gnd.n478 585
R3363 gnd.n6834 gnd.n479 585
R3364 gnd.n5957 gnd.n5956 585
R3365 gnd.n5959 gnd.n5958 585
R3366 gnd.n6089 gnd.n5960 585
R3367 gnd.n6088 gnd.n5961 585
R3368 gnd.n5963 gnd.n5962 585
R3369 gnd.n6081 gnd.n5971 585
R3370 gnd.n6080 gnd.n5972 585
R3371 gnd.n5979 gnd.n5973 585
R3372 gnd.n6073 gnd.n5980 585
R3373 gnd.n6072 gnd.n5981 585
R3374 gnd.n5983 gnd.n5982 585
R3375 gnd.n6065 gnd.n5991 585
R3376 gnd.n6064 gnd.n5992 585
R3377 gnd.n5999 gnd.n5993 585
R3378 gnd.n6057 gnd.n6000 585
R3379 gnd.n6056 gnd.n6001 585
R3380 gnd.n6003 gnd.n6002 585
R3381 gnd.n6049 gnd.n6046 585
R3382 gnd.n6045 gnd.n517 585
R3383 gnd.n6906 gnd.n517 585
R3384 gnd.n7436 gnd.n7435 585
R3385 gnd.n7308 gnd.n120 585
R3386 gnd.n7310 gnd.n7309 585
R3387 gnd.n7306 gnd.n7305 585
R3388 gnd.n7314 gnd.n7304 585
R3389 gnd.n7315 gnd.n7302 585
R3390 gnd.n7316 gnd.n7301 585
R3391 gnd.n7299 gnd.n7297 585
R3392 gnd.n7320 gnd.n7296 585
R3393 gnd.n7321 gnd.n7294 585
R3394 gnd.n7322 gnd.n7293 585
R3395 gnd.n7291 gnd.n7289 585
R3396 gnd.n7326 gnd.n7288 585
R3397 gnd.n7327 gnd.n7286 585
R3398 gnd.n7328 gnd.n7285 585
R3399 gnd.n7283 gnd.n7281 585
R3400 gnd.n7332 gnd.n7280 585
R3401 gnd.n7333 gnd.n7278 585
R3402 gnd.n7334 gnd.n7277 585
R3403 gnd.n7277 gnd.n124 585
R3404 gnd.n7434 gnd.n116 585
R3405 gnd.n7434 gnd.n7433 585
R3406 gnd.n7440 gnd.n115 585
R3407 gnd.n122 gnd.n115 585
R3408 gnd.n7441 gnd.n114 585
R3409 gnd.n7353 gnd.n114 585
R3410 gnd.n7442 gnd.n113 585
R3411 gnd.n202 gnd.n113 585
R3412 gnd.n211 gnd.n111 585
R3413 gnd.n7345 gnd.n211 585
R3414 gnd.n7446 gnd.n110 585
R3415 gnd.n209 gnd.n110 585
R3416 gnd.n7447 gnd.n109 585
R3417 gnd.n7269 gnd.n109 585
R3418 gnd.n7448 gnd.n108 585
R3419 gnd.n228 gnd.n108 585
R3420 gnd.n227 gnd.n106 585
R3421 gnd.n7261 gnd.n227 585
R3422 gnd.n7452 gnd.n105 585
R3423 gnd.n225 gnd.n105 585
R3424 gnd.n7453 gnd.n104 585
R3425 gnd.n7253 gnd.n104 585
R3426 gnd.n7454 gnd.n103 585
R3427 gnd.n234 gnd.n103 585
R3428 gnd.n243 gnd.n101 585
R3429 gnd.n7245 gnd.n243 585
R3430 gnd.n7458 gnd.n100 585
R3431 gnd.n250 gnd.n100 585
R3432 gnd.n7459 gnd.n99 585
R3433 gnd.n7237 gnd.n99 585
R3434 gnd.n7460 gnd.n98 585
R3435 gnd.n259 gnd.n98 585
R3436 gnd.n258 gnd.n96 585
R3437 gnd.n7229 gnd.n258 585
R3438 gnd.n7464 gnd.n95 585
R3439 gnd.n256 gnd.n95 585
R3440 gnd.n7465 gnd.n94 585
R3441 gnd.n7221 gnd.n94 585
R3442 gnd.n7466 gnd.n93 585
R3443 gnd.n265 gnd.n93 585
R3444 gnd.n273 gnd.n91 585
R3445 gnd.n7213 gnd.n273 585
R3446 gnd.n7470 gnd.n90 585
R3447 gnd.n280 gnd.n90 585
R3448 gnd.n7471 gnd.n89 585
R3449 gnd.n7205 gnd.n89 585
R3450 gnd.n7472 gnd.n88 585
R3451 gnd.n289 gnd.n88 585
R3452 gnd.n288 gnd.n86 585
R3453 gnd.n7197 gnd.n288 585
R3454 gnd.n7476 gnd.n85 585
R3455 gnd.n286 gnd.n85 585
R3456 gnd.n7477 gnd.n84 585
R3457 gnd.n7189 gnd.n84 585
R3458 gnd.n7478 gnd.n83 585
R3459 gnd.n295 gnd.n83 585
R3460 gnd.n325 gnd.n81 585
R3461 gnd.n7165 gnd.n325 585
R3462 gnd.n7482 gnd.n80 585
R3463 gnd.n7161 gnd.n80 585
R3464 gnd.n7483 gnd.n79 585
R3465 gnd.n330 gnd.n79 585
R3466 gnd.n7484 gnd.n78 585
R3467 gnd.n7088 gnd.n78 585
R3468 gnd.n340 gnd.n76 585
R3469 gnd.n340 gnd.n336 585
R3470 gnd.n7064 gnd.n341 585
R3471 gnd.n7082 gnd.n341 585
R3472 gnd.n7065 gnd.n7063 585
R3473 gnd.n7063 gnd.n7062 585
R3474 gnd.n353 gnd.n310 585
R3475 gnd.n7180 gnd.n310 585
R3476 gnd.n7070 gnd.n7069 585
R3477 gnd.n7071 gnd.n7070 585
R3478 gnd.n352 gnd.n351 585
R3479 gnd.n351 gnd.n349 585
R3480 gnd.n382 gnd.n360 585
R3481 gnd.n7050 gnd.n360 585
R3482 gnd.n7028 gnd.n7027 585
R3483 gnd.n7029 gnd.n7028 585
R3484 gnd.n381 gnd.n380 585
R3485 gnd.n6790 gnd.n380 585
R3486 gnd.n7022 gnd.n371 585
R3487 gnd.n7041 gnd.n371 585
R3488 gnd.n7021 gnd.n7020 585
R3489 gnd.n7020 gnd.n7019 585
R3490 gnd.n385 gnd.n384 585
R3491 gnd.n6998 gnd.n385 585
R3492 gnd.n6802 gnd.n6799 585
R3493 gnd.n6799 gnd.n6798 585
R3494 gnd.n6803 gnd.n403 585
R3495 gnd.n6990 gnd.n403 585
R3496 gnd.n6804 gnd.n584 585
R3497 gnd.n6777 gnd.n584 585
R3498 gnd.n582 gnd.n414 585
R3499 gnd.n6979 gnd.n414 585
R3500 gnd.n6808 gnd.n581 585
R3501 gnd.n6758 gnd.n581 585
R3502 gnd.n6809 gnd.n421 585
R3503 gnd.n6971 gnd.n421 585
R3504 gnd.n6810 gnd.n580 585
R3505 gnd.n6764 gnd.n580 585
R3506 gnd.n578 gnd.n430 585
R3507 gnd.n6963 gnd.n430 585
R3508 gnd.n6814 gnd.n577 585
R3509 gnd.n6750 gnd.n577 585
R3510 gnd.n6815 gnd.n439 585
R3511 gnd.n6955 gnd.n439 585
R3512 gnd.n6816 gnd.n576 585
R3513 gnd.n6746 gnd.n576 585
R3514 gnd.n574 gnd.n448 585
R3515 gnd.n6947 gnd.n448 585
R3516 gnd.n6820 gnd.n573 585
R3517 gnd.n6719 gnd.n573 585
R3518 gnd.n6821 gnd.n455 585
R3519 gnd.n6939 gnd.n455 585
R3520 gnd.n6822 gnd.n572 585
R3521 gnd.n6725 gnd.n572 585
R3522 gnd.n570 gnd.n464 585
R3523 gnd.n6931 gnd.n464 585
R3524 gnd.n6826 gnd.n569 585
R3525 gnd.n6710 gnd.n569 585
R3526 gnd.n6827 gnd.n473 585
R3527 gnd.n6923 gnd.n473 585
R3528 gnd.n6828 gnd.n568 585
R3529 gnd.n6706 gnd.n568 585
R3530 gnd.n565 gnd.n482 585
R3531 gnd.n6915 gnd.n482 585
R3532 gnd.n6833 gnd.n6832 585
R3533 gnd.n6834 gnd.n6833 585
R3534 gnd.n4075 gnd.n4074 585
R3535 gnd.n4076 gnd.n4075 585
R3536 gnd.n2769 gnd.n2768 585
R3537 gnd.n2776 gnd.n2768 585
R3538 gnd.n4057 gnd.n4056 585
R3539 gnd.n4058 gnd.n4057 585
R3540 gnd.n2787 gnd.n2786 585
R3541 gnd.n2786 gnd.n2782 585
R3542 gnd.n4047 gnd.n4046 585
R3543 gnd.n4048 gnd.n4047 585
R3544 gnd.n2795 gnd.n2794 585
R3545 gnd.n2800 gnd.n2794 585
R3546 gnd.n3769 gnd.n2812 585
R3547 gnd.n2812 gnd.n2799 585
R3548 gnd.n3771 gnd.n3770 585
R3549 gnd.n3772 gnd.n3771 585
R3550 gnd.n2813 gnd.n2811 585
R3551 gnd.n2811 gnd.n2807 585
R3552 gnd.n3760 gnd.n3759 585
R3553 gnd.n3761 gnd.n3760 585
R3554 gnd.n2820 gnd.n2819 585
R3555 gnd.n2825 gnd.n2819 585
R3556 gnd.n3738 gnd.n2838 585
R3557 gnd.n2838 gnd.n2824 585
R3558 gnd.n3740 gnd.n3739 585
R3559 gnd.n3741 gnd.n3740 585
R3560 gnd.n2839 gnd.n2837 585
R3561 gnd.n2837 gnd.n2833 585
R3562 gnd.n3729 gnd.n3728 585
R3563 gnd.n3730 gnd.n3729 585
R3564 gnd.n2846 gnd.n2845 585
R3565 gnd.n2850 gnd.n2845 585
R3566 gnd.n3707 gnd.n2862 585
R3567 gnd.n3000 gnd.n2862 585
R3568 gnd.n3709 gnd.n3708 585
R3569 gnd.n3710 gnd.n3709 585
R3570 gnd.n2863 gnd.n2861 585
R3571 gnd.n2861 gnd.n2858 585
R3572 gnd.n3698 gnd.n3697 585
R3573 gnd.n3699 gnd.n3698 585
R3574 gnd.n2870 gnd.n2869 585
R3575 gnd.n2875 gnd.n2869 585
R3576 gnd.n3676 gnd.n2888 585
R3577 gnd.n2888 gnd.n2874 585
R3578 gnd.n3678 gnd.n3677 585
R3579 gnd.n3679 gnd.n3678 585
R3580 gnd.n2889 gnd.n2887 585
R3581 gnd.n2887 gnd.n2883 585
R3582 gnd.n3667 gnd.n3666 585
R3583 gnd.n3668 gnd.n3667 585
R3584 gnd.n2897 gnd.n2896 585
R3585 gnd.n2902 gnd.n2896 585
R3586 gnd.n3645 gnd.n2914 585
R3587 gnd.n2914 gnd.n2901 585
R3588 gnd.n3647 gnd.n3646 585
R3589 gnd.n3648 gnd.n3647 585
R3590 gnd.n2915 gnd.n2913 585
R3591 gnd.n2913 gnd.n2909 585
R3592 gnd.n3636 gnd.n3635 585
R3593 gnd.n3637 gnd.n3636 585
R3594 gnd.n2922 gnd.n2921 585
R3595 gnd.n3025 gnd.n2921 585
R3596 gnd.n3614 gnd.n2937 585
R3597 gnd.n2937 gnd.n2926 585
R3598 gnd.n3616 gnd.n3615 585
R3599 gnd.n3617 gnd.n3616 585
R3600 gnd.n2938 gnd.n2936 585
R3601 gnd.n3606 gnd.n2936 585
R3602 gnd.n3106 gnd.n3105 585
R3603 gnd.n3106 gnd.n2943 585
R3604 gnd.n3593 gnd.n3592 585
R3605 gnd.n3592 gnd.n3591 585
R3606 gnd.n3594 gnd.n3098 585
R3607 gnd.n3571 gnd.n3098 585
R3608 gnd.n3596 gnd.n3595 585
R3609 gnd.n3597 gnd.n3596 585
R3610 gnd.n3099 gnd.n3097 585
R3611 gnd.n3579 gnd.n3097 585
R3612 gnd.n3563 gnd.n3562 585
R3613 gnd.n3562 gnd.n3116 585
R3614 gnd.n3561 gnd.n3121 585
R3615 gnd.n3561 gnd.n3560 585
R3616 gnd.n3546 gnd.n3122 585
R3617 gnd.n3130 gnd.n3122 585
R3618 gnd.n3548 gnd.n3547 585
R3619 gnd.n3549 gnd.n3548 585
R3620 gnd.n3133 gnd.n3132 585
R3621 gnd.n3140 gnd.n3132 585
R3622 gnd.n3521 gnd.n3520 585
R3623 gnd.n3522 gnd.n3521 585
R3624 gnd.n3152 gnd.n3151 585
R3625 gnd.n3151 gnd.n3147 585
R3626 gnd.n3511 gnd.n3510 585
R3627 gnd.n3512 gnd.n3511 585
R3628 gnd.n3162 gnd.n3161 585
R3629 gnd.n3167 gnd.n3161 585
R3630 gnd.n3489 gnd.n3180 585
R3631 gnd.n3180 gnd.n3166 585
R3632 gnd.n3491 gnd.n3490 585
R3633 gnd.n3492 gnd.n3491 585
R3634 gnd.n3181 gnd.n3179 585
R3635 gnd.n3179 gnd.n3175 585
R3636 gnd.n3480 gnd.n3479 585
R3637 gnd.n3481 gnd.n3480 585
R3638 gnd.n3188 gnd.n3187 585
R3639 gnd.n3192 gnd.n3187 585
R3640 gnd.n3457 gnd.n3209 585
R3641 gnd.n3209 gnd.n3191 585
R3642 gnd.n3459 gnd.n3458 585
R3643 gnd.n3460 gnd.n3459 585
R3644 gnd.n3210 gnd.n3208 585
R3645 gnd.n3208 gnd.n3199 585
R3646 gnd.n3452 gnd.n3451 585
R3647 gnd.n3451 gnd.n3450 585
R3648 gnd.n3257 gnd.n3256 585
R3649 gnd.n3258 gnd.n3257 585
R3650 gnd.n3411 gnd.n3410 585
R3651 gnd.n3412 gnd.n3411 585
R3652 gnd.n3267 gnd.n3266 585
R3653 gnd.n3266 gnd.n3265 585
R3654 gnd.n3406 gnd.n3405 585
R3655 gnd.n3405 gnd.n3404 585
R3656 gnd.n3270 gnd.n3269 585
R3657 gnd.n3271 gnd.n3270 585
R3658 gnd.n3395 gnd.n3394 585
R3659 gnd.n3396 gnd.n3395 585
R3660 gnd.n3278 gnd.n3277 585
R3661 gnd.n3387 gnd.n3277 585
R3662 gnd.n3390 gnd.n3389 585
R3663 gnd.n3389 gnd.n3388 585
R3664 gnd.n3281 gnd.n3280 585
R3665 gnd.n3282 gnd.n3281 585
R3666 gnd.n3376 gnd.n3375 585
R3667 gnd.n3374 gnd.n3300 585
R3668 gnd.n3373 gnd.n3299 585
R3669 gnd.n3378 gnd.n3299 585
R3670 gnd.n3372 gnd.n3371 585
R3671 gnd.n3370 gnd.n3369 585
R3672 gnd.n3368 gnd.n3367 585
R3673 gnd.n3366 gnd.n3365 585
R3674 gnd.n3364 gnd.n3363 585
R3675 gnd.n3362 gnd.n3361 585
R3676 gnd.n3360 gnd.n3359 585
R3677 gnd.n3358 gnd.n3357 585
R3678 gnd.n3356 gnd.n3355 585
R3679 gnd.n3354 gnd.n3353 585
R3680 gnd.n3352 gnd.n3351 585
R3681 gnd.n3350 gnd.n3349 585
R3682 gnd.n3348 gnd.n3347 585
R3683 gnd.n3346 gnd.n3345 585
R3684 gnd.n3344 gnd.n3343 585
R3685 gnd.n3342 gnd.n3341 585
R3686 gnd.n3340 gnd.n3339 585
R3687 gnd.n3338 gnd.n3337 585
R3688 gnd.n3336 gnd.n3335 585
R3689 gnd.n3334 gnd.n3333 585
R3690 gnd.n3332 gnd.n3331 585
R3691 gnd.n3330 gnd.n3329 585
R3692 gnd.n3287 gnd.n3286 585
R3693 gnd.n3381 gnd.n3380 585
R3694 gnd.n4079 gnd.n4078 585
R3695 gnd.n4081 gnd.n4080 585
R3696 gnd.n4083 gnd.n4082 585
R3697 gnd.n4085 gnd.n4084 585
R3698 gnd.n4087 gnd.n4086 585
R3699 gnd.n4089 gnd.n4088 585
R3700 gnd.n4091 gnd.n4090 585
R3701 gnd.n4093 gnd.n4092 585
R3702 gnd.n4095 gnd.n4094 585
R3703 gnd.n4097 gnd.n4096 585
R3704 gnd.n4099 gnd.n4098 585
R3705 gnd.n4101 gnd.n4100 585
R3706 gnd.n4103 gnd.n4102 585
R3707 gnd.n4105 gnd.n4104 585
R3708 gnd.n4107 gnd.n4106 585
R3709 gnd.n4109 gnd.n4108 585
R3710 gnd.n4111 gnd.n4110 585
R3711 gnd.n4113 gnd.n4112 585
R3712 gnd.n4115 gnd.n4114 585
R3713 gnd.n4117 gnd.n4116 585
R3714 gnd.n4119 gnd.n4118 585
R3715 gnd.n4121 gnd.n4120 585
R3716 gnd.n4123 gnd.n4122 585
R3717 gnd.n4125 gnd.n4124 585
R3718 gnd.n4127 gnd.n4126 585
R3719 gnd.n4128 gnd.n1443 585
R3720 gnd.n4129 gnd.n1401 585
R3721 gnd.n4167 gnd.n1401 585
R3722 gnd.n4077 gnd.n1473 585
R3723 gnd.n4077 gnd.n4076 585
R3724 gnd.n2976 gnd.n1472 585
R3725 gnd.n2776 gnd.n1472 585
R3726 gnd.n2977 gnd.n2784 585
R3727 gnd.n4058 gnd.n2784 585
R3728 gnd.n2979 gnd.n2978 585
R3729 gnd.n2978 gnd.n2782 585
R3730 gnd.n2980 gnd.n2793 585
R3731 gnd.n4048 gnd.n2793 585
R3732 gnd.n2982 gnd.n2981 585
R3733 gnd.n2982 gnd.n2800 585
R3734 gnd.n2984 gnd.n2983 585
R3735 gnd.n2983 gnd.n2799 585
R3736 gnd.n2985 gnd.n2809 585
R3737 gnd.n3772 gnd.n2809 585
R3738 gnd.n2987 gnd.n2986 585
R3739 gnd.n2986 gnd.n2807 585
R3740 gnd.n2988 gnd.n2818 585
R3741 gnd.n3761 gnd.n2818 585
R3742 gnd.n2990 gnd.n2989 585
R3743 gnd.n2990 gnd.n2825 585
R3744 gnd.n2992 gnd.n2991 585
R3745 gnd.n2991 gnd.n2824 585
R3746 gnd.n2993 gnd.n2835 585
R3747 gnd.n3741 gnd.n2835 585
R3748 gnd.n2995 gnd.n2994 585
R3749 gnd.n2994 gnd.n2833 585
R3750 gnd.n2996 gnd.n2844 585
R3751 gnd.n3730 gnd.n2844 585
R3752 gnd.n2998 gnd.n2997 585
R3753 gnd.n2998 gnd.n2850 585
R3754 gnd.n3002 gnd.n3001 585
R3755 gnd.n3001 gnd.n3000 585
R3756 gnd.n3003 gnd.n2860 585
R3757 gnd.n3710 gnd.n2860 585
R3758 gnd.n3005 gnd.n3004 585
R3759 gnd.n3004 gnd.n2858 585
R3760 gnd.n3006 gnd.n2868 585
R3761 gnd.n3699 gnd.n2868 585
R3762 gnd.n3008 gnd.n3007 585
R3763 gnd.n3008 gnd.n2875 585
R3764 gnd.n3010 gnd.n3009 585
R3765 gnd.n3009 gnd.n2874 585
R3766 gnd.n3011 gnd.n2885 585
R3767 gnd.n3679 gnd.n2885 585
R3768 gnd.n3013 gnd.n3012 585
R3769 gnd.n3012 gnd.n2883 585
R3770 gnd.n3014 gnd.n2895 585
R3771 gnd.n3668 gnd.n2895 585
R3772 gnd.n3016 gnd.n3015 585
R3773 gnd.n3016 gnd.n2902 585
R3774 gnd.n3018 gnd.n3017 585
R3775 gnd.n3017 gnd.n2901 585
R3776 gnd.n3019 gnd.n2911 585
R3777 gnd.n3648 gnd.n2911 585
R3778 gnd.n3021 gnd.n3020 585
R3779 gnd.n3020 gnd.n2909 585
R3780 gnd.n3022 gnd.n2920 585
R3781 gnd.n3637 gnd.n2920 585
R3782 gnd.n3027 gnd.n3026 585
R3783 gnd.n3026 gnd.n3025 585
R3784 gnd.n3023 gnd.n2946 585
R3785 gnd.n3023 gnd.n2926 585
R3786 gnd.n3603 gnd.n2934 585
R3787 gnd.n3617 gnd.n2934 585
R3788 gnd.n3605 gnd.n3604 585
R3789 gnd.n3606 gnd.n3605 585
R3790 gnd.n3107 gnd.n2944 585
R3791 gnd.n2944 gnd.n2943 585
R3792 gnd.n3109 gnd.n3108 585
R3793 gnd.n3591 gnd.n3109 585
R3794 gnd.n3094 gnd.n3092 585
R3795 gnd.n3571 gnd.n3094 585
R3796 gnd.n3599 gnd.n3598 585
R3797 gnd.n3598 gnd.n3597 585
R3798 gnd.n3093 gnd.n3091 585
R3799 gnd.n3579 gnd.n3093 585
R3800 gnd.n3556 gnd.n3125 585
R3801 gnd.n3125 gnd.n3116 585
R3802 gnd.n3558 gnd.n3557 585
R3803 gnd.n3560 gnd.n3558 585
R3804 gnd.n3126 gnd.n3124 585
R3805 gnd.n3130 gnd.n3124 585
R3806 gnd.n3551 gnd.n3550 585
R3807 gnd.n3550 gnd.n3549 585
R3808 gnd.n3129 gnd.n3128 585
R3809 gnd.n3140 gnd.n3129 585
R3810 gnd.n3430 gnd.n3149 585
R3811 gnd.n3522 gnd.n3149 585
R3812 gnd.n3432 gnd.n3431 585
R3813 gnd.n3431 gnd.n3147 585
R3814 gnd.n3433 gnd.n3160 585
R3815 gnd.n3512 gnd.n3160 585
R3816 gnd.n3435 gnd.n3434 585
R3817 gnd.n3435 gnd.n3167 585
R3818 gnd.n3437 gnd.n3436 585
R3819 gnd.n3436 gnd.n3166 585
R3820 gnd.n3438 gnd.n3177 585
R3821 gnd.n3492 gnd.n3177 585
R3822 gnd.n3440 gnd.n3439 585
R3823 gnd.n3439 gnd.n3175 585
R3824 gnd.n3441 gnd.n3186 585
R3825 gnd.n3481 gnd.n3186 585
R3826 gnd.n3443 gnd.n3442 585
R3827 gnd.n3443 gnd.n3192 585
R3828 gnd.n3445 gnd.n3444 585
R3829 gnd.n3444 gnd.n3191 585
R3830 gnd.n3446 gnd.n3207 585
R3831 gnd.n3460 gnd.n3207 585
R3832 gnd.n3447 gnd.n3260 585
R3833 gnd.n3260 gnd.n3199 585
R3834 gnd.n3449 gnd.n3448 585
R3835 gnd.n3450 gnd.n3449 585
R3836 gnd.n3261 gnd.n3259 585
R3837 gnd.n3259 gnd.n3258 585
R3838 gnd.n3414 gnd.n3413 585
R3839 gnd.n3413 gnd.n3412 585
R3840 gnd.n3264 gnd.n3263 585
R3841 gnd.n3265 gnd.n3264 585
R3842 gnd.n3403 gnd.n3402 585
R3843 gnd.n3404 gnd.n3403 585
R3844 gnd.n3273 gnd.n3272 585
R3845 gnd.n3272 gnd.n3271 585
R3846 gnd.n3398 gnd.n3397 585
R3847 gnd.n3397 gnd.n3396 585
R3848 gnd.n3276 gnd.n3275 585
R3849 gnd.n3387 gnd.n3276 585
R3850 gnd.n3386 gnd.n3385 585
R3851 gnd.n3388 gnd.n3386 585
R3852 gnd.n3284 gnd.n3283 585
R3853 gnd.n3283 gnd.n3282 585
R3854 gnd.n4066 gnd.n1423 585
R3855 gnd.n1423 gnd.n1400 585
R3856 gnd.n4068 gnd.n4067 585
R3857 gnd.n4069 gnd.n4068 585
R3858 gnd.n2778 gnd.n2777 585
R3859 gnd.n2785 gnd.n2777 585
R3860 gnd.n4061 gnd.n4060 585
R3861 gnd.n4060 gnd.n4059 585
R3862 gnd.n2781 gnd.n2780 585
R3863 gnd.n4049 gnd.n2781 585
R3864 gnd.n3780 gnd.n2802 585
R3865 gnd.n2802 gnd.n2792 585
R3866 gnd.n3782 gnd.n3781 585
R3867 gnd.n3783 gnd.n3782 585
R3868 gnd.n2803 gnd.n2801 585
R3869 gnd.n2810 gnd.n2801 585
R3870 gnd.n3775 gnd.n3774 585
R3871 gnd.n3774 gnd.n3773 585
R3872 gnd.n2806 gnd.n2805 585
R3873 gnd.n3762 gnd.n2806 585
R3874 gnd.n3749 gnd.n2828 585
R3875 gnd.n2828 gnd.n2827 585
R3876 gnd.n3751 gnd.n3750 585
R3877 gnd.n3752 gnd.n3751 585
R3878 gnd.n2829 gnd.n2826 585
R3879 gnd.n2836 gnd.n2826 585
R3880 gnd.n3744 gnd.n3743 585
R3881 gnd.n3743 gnd.n3742 585
R3882 gnd.n2832 gnd.n2831 585
R3883 gnd.n3731 gnd.n2832 585
R3884 gnd.n3718 gnd.n2853 585
R3885 gnd.n2853 gnd.n2852 585
R3886 gnd.n3720 gnd.n3719 585
R3887 gnd.n3721 gnd.n3720 585
R3888 gnd.n2854 gnd.n2851 585
R3889 gnd.n2999 gnd.n2851 585
R3890 gnd.n3713 gnd.n3712 585
R3891 gnd.n3712 gnd.n3711 585
R3892 gnd.n2857 gnd.n2856 585
R3893 gnd.n3700 gnd.n2857 585
R3894 gnd.n3687 gnd.n2878 585
R3895 gnd.n2878 gnd.n2877 585
R3896 gnd.n3689 gnd.n3688 585
R3897 gnd.n3690 gnd.n3689 585
R3898 gnd.n2879 gnd.n2876 585
R3899 gnd.n2886 gnd.n2876 585
R3900 gnd.n3682 gnd.n3681 585
R3901 gnd.n3681 gnd.n3680 585
R3902 gnd.n2882 gnd.n2881 585
R3903 gnd.n3669 gnd.n2882 585
R3904 gnd.n3656 gnd.n2904 585
R3905 gnd.n2904 gnd.n2894 585
R3906 gnd.n3658 gnd.n3657 585
R3907 gnd.n3659 gnd.n3658 585
R3908 gnd.n2905 gnd.n2903 585
R3909 gnd.n2912 gnd.n2903 585
R3910 gnd.n3651 gnd.n3650 585
R3911 gnd.n3650 gnd.n3649 585
R3912 gnd.n2908 gnd.n2907 585
R3913 gnd.n3638 gnd.n2908 585
R3914 gnd.n3625 gnd.n2928 585
R3915 gnd.n3024 gnd.n2928 585
R3916 gnd.n3627 gnd.n3626 585
R3917 gnd.n3628 gnd.n3627 585
R3918 gnd.n2929 gnd.n2927 585
R3919 gnd.n2935 gnd.n2927 585
R3920 gnd.n3620 gnd.n3619 585
R3921 gnd.n3619 gnd.n3618 585
R3922 gnd.n2932 gnd.n2931 585
R3923 gnd.n3607 gnd.n2932 585
R3924 gnd.n3589 gnd.n3588 585
R3925 gnd.n3590 gnd.n3589 585
R3926 gnd.n3111 gnd.n3110 585
R3927 gnd.n3572 gnd.n3110 585
R3928 gnd.n3584 gnd.n3583 585
R3929 gnd.n3583 gnd.n3096 585
R3930 gnd.n3582 gnd.n3113 585
R3931 gnd.n3582 gnd.n3095 585
R3932 gnd.n3581 gnd.n3115 585
R3933 gnd.n3581 gnd.n3580 585
R3934 gnd.n3533 gnd.n3114 585
R3935 gnd.n3559 gnd.n3114 585
R3936 gnd.n3535 gnd.n3534 585
R3937 gnd.n3534 gnd.n3123 585
R3938 gnd.n3536 gnd.n3142 585
R3939 gnd.n3142 gnd.n3131 585
R3940 gnd.n3538 gnd.n3537 585
R3941 gnd.n3539 gnd.n3538 585
R3942 gnd.n3143 gnd.n3141 585
R3943 gnd.n3150 gnd.n3141 585
R3944 gnd.n3525 gnd.n3524 585
R3945 gnd.n3524 gnd.n3523 585
R3946 gnd.n3146 gnd.n3145 585
R3947 gnd.n3513 gnd.n3146 585
R3948 gnd.n3500 gnd.n3170 585
R3949 gnd.n3170 gnd.n3169 585
R3950 gnd.n3502 gnd.n3501 585
R3951 gnd.n3503 gnd.n3502 585
R3952 gnd.n3171 gnd.n3168 585
R3953 gnd.n3178 gnd.n3168 585
R3954 gnd.n3495 gnd.n3494 585
R3955 gnd.n3494 gnd.n3493 585
R3956 gnd.n3174 gnd.n3173 585
R3957 gnd.n3482 gnd.n3174 585
R3958 gnd.n3469 gnd.n3195 585
R3959 gnd.n3195 gnd.n3194 585
R3960 gnd.n3471 gnd.n3470 585
R3961 gnd.n3472 gnd.n3471 585
R3962 gnd.n3465 gnd.n3193 585
R3963 gnd.n3464 gnd.n3463 585
R3964 gnd.n3198 gnd.n3197 585
R3965 gnd.n3461 gnd.n3198 585
R3966 gnd.n3220 gnd.n3219 585
R3967 gnd.n3223 gnd.n3222 585
R3968 gnd.n3221 gnd.n3216 585
R3969 gnd.n3228 gnd.n3227 585
R3970 gnd.n3230 gnd.n3229 585
R3971 gnd.n3233 gnd.n3232 585
R3972 gnd.n3231 gnd.n3214 585
R3973 gnd.n3238 gnd.n3237 585
R3974 gnd.n3240 gnd.n3239 585
R3975 gnd.n3243 gnd.n3242 585
R3976 gnd.n3241 gnd.n3212 585
R3977 gnd.n3248 gnd.n3247 585
R3978 gnd.n3252 gnd.n3249 585
R3979 gnd.n3253 gnd.n3190 585
R3980 gnd.n2774 gnd.n1438 585
R3981 gnd.n4135 gnd.n4134 585
R3982 gnd.n4137 gnd.n4136 585
R3983 gnd.n4139 gnd.n4138 585
R3984 gnd.n4141 gnd.n4140 585
R3985 gnd.n4143 gnd.n4142 585
R3986 gnd.n4145 gnd.n4144 585
R3987 gnd.n4147 gnd.n4146 585
R3988 gnd.n4149 gnd.n4148 585
R3989 gnd.n4151 gnd.n4150 585
R3990 gnd.n4153 gnd.n4152 585
R3991 gnd.n4155 gnd.n4154 585
R3992 gnd.n4157 gnd.n4156 585
R3993 gnd.n4160 gnd.n4159 585
R3994 gnd.n4158 gnd.n1426 585
R3995 gnd.n4164 gnd.n1424 585
R3996 gnd.n4166 gnd.n4165 585
R3997 gnd.n4167 gnd.n4166 585
R3998 gnd.n2775 gnd.n2772 585
R3999 gnd.n2775 gnd.n1400 585
R4000 gnd.n4071 gnd.n4070 585
R4001 gnd.n4070 gnd.n4069 585
R4002 gnd.n2773 gnd.n2771 585
R4003 gnd.n2785 gnd.n2773 585
R4004 gnd.n4052 gnd.n2783 585
R4005 gnd.n4059 gnd.n2783 585
R4006 gnd.n4051 gnd.n4050 585
R4007 gnd.n4050 gnd.n4049 585
R4008 gnd.n2791 gnd.n2789 585
R4009 gnd.n2792 gnd.n2791 585
R4010 gnd.n3785 gnd.n3784 585
R4011 gnd.n3784 gnd.n3783 585
R4012 gnd.n2798 gnd.n2797 585
R4013 gnd.n2810 gnd.n2798 585
R4014 gnd.n3765 gnd.n2808 585
R4015 gnd.n3773 gnd.n2808 585
R4016 gnd.n3764 gnd.n3763 585
R4017 gnd.n3763 gnd.n3762 585
R4018 gnd.n2817 gnd.n2815 585
R4019 gnd.n2827 gnd.n2817 585
R4020 gnd.n3754 gnd.n3753 585
R4021 gnd.n3753 gnd.n3752 585
R4022 gnd.n2823 gnd.n2822 585
R4023 gnd.n2836 gnd.n2823 585
R4024 gnd.n3734 gnd.n2834 585
R4025 gnd.n3742 gnd.n2834 585
R4026 gnd.n3733 gnd.n3732 585
R4027 gnd.n3732 gnd.n3731 585
R4028 gnd.n2843 gnd.n2841 585
R4029 gnd.n2852 gnd.n2843 585
R4030 gnd.n3723 gnd.n3722 585
R4031 gnd.n3722 gnd.n3721 585
R4032 gnd.n2849 gnd.n2848 585
R4033 gnd.n2999 gnd.n2849 585
R4034 gnd.n3703 gnd.n2859 585
R4035 gnd.n3711 gnd.n2859 585
R4036 gnd.n3702 gnd.n3701 585
R4037 gnd.n3701 gnd.n3700 585
R4038 gnd.n2867 gnd.n2865 585
R4039 gnd.n2877 gnd.n2867 585
R4040 gnd.n3692 gnd.n3691 585
R4041 gnd.n3691 gnd.n3690 585
R4042 gnd.n2873 gnd.n2872 585
R4043 gnd.n2886 gnd.n2873 585
R4044 gnd.n3672 gnd.n2884 585
R4045 gnd.n3680 gnd.n2884 585
R4046 gnd.n3671 gnd.n3670 585
R4047 gnd.n3670 gnd.n3669 585
R4048 gnd.n2893 gnd.n2891 585
R4049 gnd.n2894 gnd.n2893 585
R4050 gnd.n3661 gnd.n3660 585
R4051 gnd.n3660 gnd.n3659 585
R4052 gnd.n2900 gnd.n2899 585
R4053 gnd.n2912 gnd.n2900 585
R4054 gnd.n3641 gnd.n2910 585
R4055 gnd.n3649 gnd.n2910 585
R4056 gnd.n3640 gnd.n3639 585
R4057 gnd.n3639 gnd.n3638 585
R4058 gnd.n2919 gnd.n2917 585
R4059 gnd.n3024 gnd.n2919 585
R4060 gnd.n3630 gnd.n3629 585
R4061 gnd.n3629 gnd.n3628 585
R4062 gnd.n2925 gnd.n2924 585
R4063 gnd.n2935 gnd.n2925 585
R4064 gnd.n3610 gnd.n2933 585
R4065 gnd.n3618 gnd.n2933 585
R4066 gnd.n3609 gnd.n3608 585
R4067 gnd.n3608 gnd.n3607 585
R4068 gnd.n2942 gnd.n2940 585
R4069 gnd.n3590 gnd.n2942 585
R4070 gnd.n3573 gnd.n3570 585
R4071 gnd.n3573 gnd.n3572 585
R4072 gnd.n3575 gnd.n3574 585
R4073 gnd.n3574 gnd.n3096 585
R4074 gnd.n3576 gnd.n3118 585
R4075 gnd.n3118 gnd.n3095 585
R4076 gnd.n3578 gnd.n3577 585
R4077 gnd.n3580 gnd.n3578 585
R4078 gnd.n3119 gnd.n3117 585
R4079 gnd.n3559 gnd.n3117 585
R4080 gnd.n3543 gnd.n3542 585
R4081 gnd.n3542 gnd.n3123 585
R4082 gnd.n3541 gnd.n3137 585
R4083 gnd.n3541 gnd.n3131 585
R4084 gnd.n3540 gnd.n3139 585
R4085 gnd.n3540 gnd.n3539 585
R4086 gnd.n3517 gnd.n3138 585
R4087 gnd.n3150 gnd.n3138 585
R4088 gnd.n3516 gnd.n3148 585
R4089 gnd.n3523 gnd.n3148 585
R4090 gnd.n3515 gnd.n3514 585
R4091 gnd.n3514 gnd.n3513 585
R4092 gnd.n3159 gnd.n3156 585
R4093 gnd.n3169 gnd.n3159 585
R4094 gnd.n3505 gnd.n3504 585
R4095 gnd.n3504 gnd.n3503 585
R4096 gnd.n3165 gnd.n3164 585
R4097 gnd.n3178 gnd.n3165 585
R4098 gnd.n3485 gnd.n3176 585
R4099 gnd.n3493 gnd.n3176 585
R4100 gnd.n3484 gnd.n3483 585
R4101 gnd.n3483 gnd.n3482 585
R4102 gnd.n3185 gnd.n3183 585
R4103 gnd.n3194 gnd.n3185 585
R4104 gnd.n3474 gnd.n3473 585
R4105 gnd.n3473 gnd.n3472 585
R4106 gnd.n6301 gnd.n6300 585
R4107 gnd.n6302 gnd.n6301 585
R4108 gnd.n988 gnd.n986 585
R4109 gnd.n6225 gnd.n986 585
R4110 gnd.n4979 gnd.n1072 585
R4111 gnd.n4801 gnd.n1072 585
R4112 gnd.n4981 gnd.n4980 585
R4113 gnd.n4982 gnd.n4981 585
R4114 gnd.n1073 gnd.n1071 585
R4115 gnd.n4799 gnd.n1071 585
R4116 gnd.n4974 gnd.n4973 585
R4117 gnd.n4973 gnd.n4972 585
R4118 gnd.n1076 gnd.n1075 585
R4119 gnd.n4788 gnd.n1076 585
R4120 gnd.n4963 gnd.n4962 585
R4121 gnd.n4964 gnd.n4963 585
R4122 gnd.n1090 gnd.n1089 585
R4123 gnd.n4740 gnd.n1089 585
R4124 gnd.n4958 gnd.n4957 585
R4125 gnd.n4957 gnd.n4956 585
R4126 gnd.n1093 gnd.n1092 585
R4127 gnd.n4746 gnd.n1093 585
R4128 gnd.n4947 gnd.n4946 585
R4129 gnd.n4948 gnd.n4947 585
R4130 gnd.n1107 gnd.n1106 585
R4131 gnd.n4732 gnd.n1106 585
R4132 gnd.n4942 gnd.n4941 585
R4133 gnd.n4941 gnd.n4940 585
R4134 gnd.n1110 gnd.n1109 585
R4135 gnd.n4728 gnd.n1110 585
R4136 gnd.n4931 gnd.n4930 585
R4137 gnd.n4932 gnd.n4931 585
R4138 gnd.n1124 gnd.n1123 585
R4139 gnd.n4701 gnd.n1123 585
R4140 gnd.n4926 gnd.n4925 585
R4141 gnd.n4925 gnd.n4924 585
R4142 gnd.n1127 gnd.n1126 585
R4143 gnd.n4707 gnd.n1127 585
R4144 gnd.n4915 gnd.n4914 585
R4145 gnd.n4916 gnd.n4915 585
R4146 gnd.n1141 gnd.n1140 585
R4147 gnd.n4692 gnd.n1140 585
R4148 gnd.n4910 gnd.n4909 585
R4149 gnd.n4909 gnd.n4908 585
R4150 gnd.n1144 gnd.n1143 585
R4151 gnd.n4688 gnd.n1144 585
R4152 gnd.n4899 gnd.n4898 585
R4153 gnd.n4900 gnd.n4899 585
R4154 gnd.n1158 gnd.n1157 585
R4155 gnd.n4661 gnd.n1157 585
R4156 gnd.n4894 gnd.n4893 585
R4157 gnd.n4893 gnd.n4892 585
R4158 gnd.n1161 gnd.n1160 585
R4159 gnd.n4844 gnd.n1161 585
R4160 gnd.n4883 gnd.n4882 585
R4161 gnd.n4884 gnd.n4883 585
R4162 gnd.n1175 gnd.n1174 585
R4163 gnd.n4653 gnd.n1174 585
R4164 gnd.n4855 gnd.n4854 585
R4165 gnd.n4856 gnd.n4855 585
R4166 gnd.n4853 gnd.n1199 585
R4167 gnd.n4645 gnd.n1199 585
R4168 gnd.n4864 gnd.n4863 585
R4169 gnd.n4863 gnd.n4862 585
R4170 gnd.n4866 gnd.n4865 585
R4171 gnd.n4866 gnd.n1198 585
R4172 gnd.n4869 gnd.n4868 585
R4173 gnd.n4870 gnd.n4869 585
R4174 gnd.n4867 gnd.n1184 585
R4175 gnd.n1187 gnd.n1184 585
R4176 gnd.n4878 gnd.n4877 585
R4177 gnd.n4877 gnd.n4876 585
R4178 gnd.n4879 gnd.n1183 585
R4179 gnd.n4629 gnd.n1183 585
R4180 gnd.n1288 gnd.n1182 585
R4181 gnd.n1288 gnd.n1279 585
R4182 gnd.n4610 gnd.n4609 585
R4183 gnd.n4611 gnd.n4610 585
R4184 gnd.n4608 gnd.n1287 585
R4185 gnd.n4596 gnd.n1287 585
R4186 gnd.n1293 gnd.n1289 585
R4187 gnd.n1296 gnd.n1293 585
R4188 gnd.n4604 gnd.n4603 585
R4189 gnd.n4603 gnd.n4602 585
R4190 gnd.n1292 gnd.n1291 585
R4191 gnd.n4585 gnd.n1292 585
R4192 gnd.n4569 gnd.n1324 585
R4193 gnd.n1324 gnd.n1314 585
R4194 gnd.n4571 gnd.n4570 585
R4195 gnd.n4572 gnd.n4571 585
R4196 gnd.n1325 gnd.n1323 585
R4197 gnd.n1323 gnd.n1320 585
R4198 gnd.n4564 gnd.n4563 585
R4199 gnd.n4563 gnd.n4562 585
R4200 gnd.n1328 gnd.n1327 585
R4201 gnd.n1340 gnd.n1328 585
R4202 gnd.n4545 gnd.n4544 585
R4203 gnd.n4546 gnd.n4545 585
R4204 gnd.n1342 gnd.n1341 585
R4205 gnd.n1341 gnd.n1337 585
R4206 gnd.n4540 gnd.n4539 585
R4207 gnd.n4539 gnd.n4538 585
R4208 gnd.n1345 gnd.n1344 585
R4209 gnd.n1346 gnd.n1345 585
R4210 gnd.n4529 gnd.n4528 585
R4211 gnd.n4530 gnd.n4529 585
R4212 gnd.n1358 gnd.n1357 585
R4213 gnd.n1357 gnd.n1354 585
R4214 gnd.n4524 gnd.n4523 585
R4215 gnd.n4523 gnd.n4522 585
R4216 gnd.n1361 gnd.n1360 585
R4217 gnd.n1372 gnd.n1361 585
R4218 gnd.n4513 gnd.n4512 585
R4219 gnd.n4514 gnd.n4513 585
R4220 gnd.n1374 gnd.n1373 585
R4221 gnd.n1373 gnd.n1369 585
R4222 gnd.n4508 gnd.n4507 585
R4223 gnd.n4507 gnd.n4506 585
R4224 gnd.n1377 gnd.n1376 585
R4225 gnd.n1378 gnd.n1377 585
R4226 gnd.n4497 gnd.n4496 585
R4227 gnd.n4498 gnd.n4497 585
R4228 gnd.n1390 gnd.n1389 585
R4229 gnd.n1389 gnd.n1386 585
R4230 gnd.n4492 gnd.n4491 585
R4231 gnd.n4491 gnd.n4490 585
R4232 gnd.n1393 gnd.n1392 585
R4233 gnd.n4284 gnd.n1393 585
R4234 gnd.n4481 gnd.n4480 585
R4235 gnd.n4482 gnd.n4481 585
R4236 gnd.n4477 gnd.n4285 585
R4237 gnd.n4476 gnd.n4475 585
R4238 gnd.n4473 gnd.n4287 585
R4239 gnd.n4473 gnd.n4168 585
R4240 gnd.n4472 gnd.n4471 585
R4241 gnd.n4470 gnd.n4469 585
R4242 gnd.n4468 gnd.n4292 585
R4243 gnd.n4466 gnd.n4465 585
R4244 gnd.n4464 gnd.n4293 585
R4245 gnd.n4463 gnd.n4462 585
R4246 gnd.n4460 gnd.n4298 585
R4247 gnd.n4458 gnd.n4457 585
R4248 gnd.n4456 gnd.n4299 585
R4249 gnd.n4455 gnd.n4454 585
R4250 gnd.n4452 gnd.n4304 585
R4251 gnd.n4450 gnd.n4449 585
R4252 gnd.n4448 gnd.n4305 585
R4253 gnd.n4447 gnd.n4446 585
R4254 gnd.n4444 gnd.n4310 585
R4255 gnd.n4442 gnd.n4441 585
R4256 gnd.n4440 gnd.n4311 585
R4257 gnd.n4439 gnd.n4438 585
R4258 gnd.n4436 gnd.n4319 585
R4259 gnd.n4434 gnd.n4433 585
R4260 gnd.n4432 gnd.n4320 585
R4261 gnd.n4431 gnd.n4430 585
R4262 gnd.n4428 gnd.n4325 585
R4263 gnd.n4426 gnd.n4425 585
R4264 gnd.n4424 gnd.n4326 585
R4265 gnd.n4423 gnd.n4422 585
R4266 gnd.n4420 gnd.n4331 585
R4267 gnd.n4418 gnd.n4417 585
R4268 gnd.n4416 gnd.n4332 585
R4269 gnd.n4415 gnd.n4414 585
R4270 gnd.n4412 gnd.n4337 585
R4271 gnd.n4410 gnd.n4409 585
R4272 gnd.n4408 gnd.n4338 585
R4273 gnd.n4407 gnd.n4343 585
R4274 gnd.n4400 gnd.n4346 585
R4275 gnd.n4403 gnd.n4402 585
R4276 gnd.n6232 gnd.n6231 585
R4277 gnd.n6234 gnd.n1055 585
R4278 gnd.n6236 gnd.n6235 585
R4279 gnd.n6237 gnd.n1048 585
R4280 gnd.n6239 gnd.n6238 585
R4281 gnd.n6241 gnd.n1046 585
R4282 gnd.n6243 gnd.n6242 585
R4283 gnd.n6244 gnd.n1041 585
R4284 gnd.n6246 gnd.n6245 585
R4285 gnd.n6248 gnd.n1039 585
R4286 gnd.n6250 gnd.n6249 585
R4287 gnd.n6251 gnd.n1034 585
R4288 gnd.n6253 gnd.n6252 585
R4289 gnd.n6255 gnd.n1032 585
R4290 gnd.n6257 gnd.n6256 585
R4291 gnd.n6258 gnd.n1027 585
R4292 gnd.n6260 gnd.n6259 585
R4293 gnd.n6262 gnd.n1025 585
R4294 gnd.n6264 gnd.n6263 585
R4295 gnd.n6265 gnd.n1019 585
R4296 gnd.n6267 gnd.n6266 585
R4297 gnd.n6271 gnd.n1014 585
R4298 gnd.n6273 gnd.n6272 585
R4299 gnd.n6274 gnd.n1009 585
R4300 gnd.n6276 gnd.n6275 585
R4301 gnd.n6278 gnd.n1007 585
R4302 gnd.n6280 gnd.n6279 585
R4303 gnd.n6281 gnd.n1002 585
R4304 gnd.n6283 gnd.n6282 585
R4305 gnd.n6285 gnd.n1000 585
R4306 gnd.n6287 gnd.n6286 585
R4307 gnd.n6288 gnd.n994 585
R4308 gnd.n6290 gnd.n6289 585
R4309 gnd.n6292 gnd.n993 585
R4310 gnd.n6293 gnd.n991 585
R4311 gnd.n6296 gnd.n6295 585
R4312 gnd.n6297 gnd.n987 585
R4313 gnd.n992 gnd.n987 585
R4314 gnd.n6228 gnd.n983 585
R4315 gnd.n6302 gnd.n983 585
R4316 gnd.n6227 gnd.n6226 585
R4317 gnd.n6226 gnd.n6225 585
R4318 gnd.n1060 gnd.n1059 585
R4319 gnd.n4801 gnd.n1060 585
R4320 gnd.n4796 gnd.n1068 585
R4321 gnd.n4982 gnd.n1068 585
R4322 gnd.n4798 gnd.n4797 585
R4323 gnd.n4799 gnd.n4798 585
R4324 gnd.n1243 gnd.n1078 585
R4325 gnd.n4972 gnd.n1078 585
R4326 gnd.n4790 gnd.n4789 585
R4327 gnd.n4789 gnd.n4788 585
R4328 gnd.n1245 gnd.n1087 585
R4329 gnd.n4964 gnd.n1087 585
R4330 gnd.n4742 gnd.n4741 585
R4331 gnd.n4741 gnd.n4740 585
R4332 gnd.n4743 gnd.n1094 585
R4333 gnd.n4956 gnd.n1094 585
R4334 gnd.n4745 gnd.n4744 585
R4335 gnd.n4746 gnd.n4745 585
R4336 gnd.n1252 gnd.n1103 585
R4337 gnd.n4948 gnd.n1103 585
R4338 gnd.n4734 gnd.n4733 585
R4339 gnd.n4733 gnd.n4732 585
R4340 gnd.n4731 gnd.n1112 585
R4341 gnd.n4940 gnd.n1112 585
R4342 gnd.n4730 gnd.n4729 585
R4343 gnd.n4729 gnd.n4728 585
R4344 gnd.n1254 gnd.n1121 585
R4345 gnd.n4932 gnd.n1121 585
R4346 gnd.n4703 gnd.n4702 585
R4347 gnd.n4702 gnd.n4701 585
R4348 gnd.n4704 gnd.n1128 585
R4349 gnd.n4924 gnd.n1128 585
R4350 gnd.n4706 gnd.n4705 585
R4351 gnd.n4707 gnd.n4706 585
R4352 gnd.n1262 gnd.n1137 585
R4353 gnd.n4916 gnd.n1137 585
R4354 gnd.n4694 gnd.n4693 585
R4355 gnd.n4693 gnd.n4692 585
R4356 gnd.n4691 gnd.n1146 585
R4357 gnd.n4908 gnd.n1146 585
R4358 gnd.n4690 gnd.n4689 585
R4359 gnd.n4689 gnd.n4688 585
R4360 gnd.n1264 gnd.n1155 585
R4361 gnd.n4900 gnd.n1155 585
R4362 gnd.n4663 gnd.n4662 585
R4363 gnd.n4662 gnd.n4661 585
R4364 gnd.n4660 gnd.n1162 585
R4365 gnd.n4892 gnd.n1162 585
R4366 gnd.n4659 gnd.n1218 585
R4367 gnd.n4844 gnd.n1218 585
R4368 gnd.n1266 gnd.n1171 585
R4369 gnd.n4884 gnd.n1171 585
R4370 gnd.n4655 gnd.n4654 585
R4371 gnd.n4654 gnd.n4653 585
R4372 gnd.n1268 gnd.n1208 585
R4373 gnd.n4856 gnd.n1208 585
R4374 gnd.n4644 gnd.n4643 585
R4375 gnd.n4645 gnd.n4644 585
R4376 gnd.n1272 gnd.n1201 585
R4377 gnd.n4862 gnd.n1201 585
R4378 gnd.n4639 gnd.n4638 585
R4379 gnd.n4638 gnd.n1198 585
R4380 gnd.n4637 gnd.n1196 585
R4381 gnd.n4870 gnd.n1196 585
R4382 gnd.n4636 gnd.n4635 585
R4383 gnd.n4635 gnd.n1187 585
R4384 gnd.n1275 gnd.n1185 585
R4385 gnd.n4876 gnd.n1185 585
R4386 gnd.n4631 gnd.n4630 585
R4387 gnd.n4630 gnd.n4629 585
R4388 gnd.n1278 gnd.n1277 585
R4389 gnd.n1279 gnd.n1278 585
R4390 gnd.n4593 gnd.n1285 585
R4391 gnd.n4611 gnd.n1285 585
R4392 gnd.n4595 gnd.n4594 585
R4393 gnd.n4596 gnd.n4595 585
R4394 gnd.n1310 gnd.n1309 585
R4395 gnd.n1309 gnd.n1296 585
R4396 gnd.n4588 gnd.n1294 585
R4397 gnd.n4602 gnd.n1294 585
R4398 gnd.n4587 gnd.n4586 585
R4399 gnd.n4586 gnd.n4585 585
R4400 gnd.n1313 gnd.n1312 585
R4401 gnd.n1314 gnd.n1313 585
R4402 gnd.n4369 gnd.n1321 585
R4403 gnd.n4572 gnd.n1321 585
R4404 gnd.n4371 gnd.n4370 585
R4405 gnd.n4370 gnd.n1320 585
R4406 gnd.n4372 gnd.n1329 585
R4407 gnd.n4562 gnd.n1329 585
R4408 gnd.n4374 gnd.n4373 585
R4409 gnd.n4373 gnd.n1340 585
R4410 gnd.n4375 gnd.n1338 585
R4411 gnd.n4546 gnd.n1338 585
R4412 gnd.n4377 gnd.n4376 585
R4413 gnd.n4376 gnd.n1337 585
R4414 gnd.n4378 gnd.n1347 585
R4415 gnd.n4538 gnd.n1347 585
R4416 gnd.n4380 gnd.n4379 585
R4417 gnd.n4379 gnd.n1346 585
R4418 gnd.n4381 gnd.n1355 585
R4419 gnd.n4530 gnd.n1355 585
R4420 gnd.n4383 gnd.n4382 585
R4421 gnd.n4382 gnd.n1354 585
R4422 gnd.n4384 gnd.n1362 585
R4423 gnd.n4522 gnd.n1362 585
R4424 gnd.n4386 gnd.n4385 585
R4425 gnd.n4385 gnd.n1372 585
R4426 gnd.n4387 gnd.n1370 585
R4427 gnd.n4514 gnd.n1370 585
R4428 gnd.n4389 gnd.n4388 585
R4429 gnd.n4388 gnd.n1369 585
R4430 gnd.n4390 gnd.n1379 585
R4431 gnd.n4506 gnd.n1379 585
R4432 gnd.n4392 gnd.n4391 585
R4433 gnd.n4391 gnd.n1378 585
R4434 gnd.n4393 gnd.n1387 585
R4435 gnd.n4498 gnd.n1387 585
R4436 gnd.n4395 gnd.n4394 585
R4437 gnd.n4394 gnd.n1386 585
R4438 gnd.n4396 gnd.n1394 585
R4439 gnd.n4490 gnd.n1394 585
R4440 gnd.n4397 gnd.n4348 585
R4441 gnd.n4348 gnd.n4284 585
R4442 gnd.n4398 gnd.n4169 585
R4443 gnd.n4482 gnd.n4169 585
R4444 gnd.n7432 gnd.n7431 585
R4445 gnd.n7433 gnd.n7432 585
R4446 gnd.n128 gnd.n126 585
R4447 gnd.n126 gnd.n122 585
R4448 gnd.n7352 gnd.n7351 585
R4449 gnd.n7353 gnd.n7352 585
R4450 gnd.n205 gnd.n204 585
R4451 gnd.n204 gnd.n202 585
R4452 gnd.n7347 gnd.n7346 585
R4453 gnd.n7346 gnd.n7345 585
R4454 gnd.n208 gnd.n207 585
R4455 gnd.n209 gnd.n208 585
R4456 gnd.n7268 gnd.n7267 585
R4457 gnd.n7269 gnd.n7268 585
R4458 gnd.n221 gnd.n220 585
R4459 gnd.n228 gnd.n220 585
R4460 gnd.n7263 gnd.n7262 585
R4461 gnd.n7262 gnd.n7261 585
R4462 gnd.n224 gnd.n223 585
R4463 gnd.n225 gnd.n224 585
R4464 gnd.n7252 gnd.n7251 585
R4465 gnd.n7253 gnd.n7252 585
R4466 gnd.n238 gnd.n237 585
R4467 gnd.n237 gnd.n234 585
R4468 gnd.n7247 gnd.n7246 585
R4469 gnd.n7246 gnd.n7245 585
R4470 gnd.n241 gnd.n240 585
R4471 gnd.n250 gnd.n241 585
R4472 gnd.n7236 gnd.n7235 585
R4473 gnd.n7237 gnd.n7236 585
R4474 gnd.n252 gnd.n251 585
R4475 gnd.n259 gnd.n251 585
R4476 gnd.n7231 gnd.n7230 585
R4477 gnd.n7230 gnd.n7229 585
R4478 gnd.n255 gnd.n254 585
R4479 gnd.n256 gnd.n255 585
R4480 gnd.n7220 gnd.n7219 585
R4481 gnd.n7221 gnd.n7220 585
R4482 gnd.n268 gnd.n267 585
R4483 gnd.n267 gnd.n265 585
R4484 gnd.n7215 gnd.n7214 585
R4485 gnd.n7214 gnd.n7213 585
R4486 gnd.n271 gnd.n270 585
R4487 gnd.n280 gnd.n271 585
R4488 gnd.n7204 gnd.n7203 585
R4489 gnd.n7205 gnd.n7204 585
R4490 gnd.n282 gnd.n281 585
R4491 gnd.n289 gnd.n281 585
R4492 gnd.n7199 gnd.n7198 585
R4493 gnd.n7198 gnd.n7197 585
R4494 gnd.n285 gnd.n284 585
R4495 gnd.n286 gnd.n285 585
R4496 gnd.n7188 gnd.n7187 585
R4497 gnd.n7189 gnd.n7188 585
R4498 gnd.n298 gnd.n297 585
R4499 gnd.n297 gnd.n295 585
R4500 gnd.n7164 gnd.n7163 585
R4501 gnd.n7165 gnd.n7164 585
R4502 gnd.n7162 gnd.n328 585
R4503 gnd.n7162 gnd.n7161 585
R4504 gnd.n327 gnd.n326 585
R4505 gnd.n330 gnd.n326 585
R4506 gnd.n7087 gnd.n7086 585
R4507 gnd.n7088 gnd.n7087 585
R4508 gnd.n7085 gnd.n7084 585
R4509 gnd.n7084 gnd.n336 585
R4510 gnd.n7083 gnd.n338 585
R4511 gnd.n7083 gnd.n7082 585
R4512 gnd.n337 gnd.n307 585
R4513 gnd.n7062 gnd.n307 585
R4514 gnd.n7182 gnd.n7181 585
R4515 gnd.n7181 gnd.n7180 585
R4516 gnd.n7183 gnd.n306 585
R4517 gnd.n7071 gnd.n306 585
R4518 gnd.n364 gnd.n305 585
R4519 gnd.n364 gnd.n349 585
R4520 gnd.n7049 gnd.n7048 585
R4521 gnd.n7050 gnd.n7049 585
R4522 gnd.n7047 gnd.n363 585
R4523 gnd.n7029 gnd.n363 585
R4524 gnd.n369 gnd.n365 585
R4525 gnd.n6790 gnd.n369 585
R4526 gnd.n7043 gnd.n7042 585
R4527 gnd.n7042 gnd.n7041 585
R4528 gnd.n368 gnd.n367 585
R4529 gnd.n7019 gnd.n368 585
R4530 gnd.n6997 gnd.n6996 585
R4531 gnd.n6998 gnd.n6997 585
R4532 gnd.n397 gnd.n396 585
R4533 gnd.n6798 gnd.n396 585
R4534 gnd.n6992 gnd.n6991 585
R4535 gnd.n6991 gnd.n6990 585
R4536 gnd.n400 gnd.n399 585
R4537 gnd.n6777 gnd.n400 585
R4538 gnd.n6978 gnd.n6977 585
R4539 gnd.n6979 gnd.n6978 585
R4540 gnd.n416 gnd.n415 585
R4541 gnd.n6758 gnd.n415 585
R4542 gnd.n6973 gnd.n6972 585
R4543 gnd.n6972 gnd.n6971 585
R4544 gnd.n419 gnd.n418 585
R4545 gnd.n6764 gnd.n419 585
R4546 gnd.n6962 gnd.n6961 585
R4547 gnd.n6963 gnd.n6962 585
R4548 gnd.n433 gnd.n432 585
R4549 gnd.n6750 gnd.n432 585
R4550 gnd.n6957 gnd.n6956 585
R4551 gnd.n6956 gnd.n6955 585
R4552 gnd.n436 gnd.n435 585
R4553 gnd.n6746 gnd.n436 585
R4554 gnd.n6946 gnd.n6945 585
R4555 gnd.n6947 gnd.n6946 585
R4556 gnd.n450 gnd.n449 585
R4557 gnd.n6719 gnd.n449 585
R4558 gnd.n6941 gnd.n6940 585
R4559 gnd.n6940 gnd.n6939 585
R4560 gnd.n453 gnd.n452 585
R4561 gnd.n6725 gnd.n453 585
R4562 gnd.n6930 gnd.n6929 585
R4563 gnd.n6931 gnd.n6930 585
R4564 gnd.n467 gnd.n466 585
R4565 gnd.n6710 gnd.n466 585
R4566 gnd.n6925 gnd.n6924 585
R4567 gnd.n6924 gnd.n6923 585
R4568 gnd.n470 gnd.n469 585
R4569 gnd.n6706 gnd.n470 585
R4570 gnd.n6914 gnd.n6913 585
R4571 gnd.n6915 gnd.n6914 585
R4572 gnd.n485 gnd.n484 585
R4573 gnd.n6834 gnd.n484 585
R4574 gnd.n6909 gnd.n6908 585
R4575 gnd.n488 gnd.n487 585
R4576 gnd.n6905 gnd.n6904 585
R4577 gnd.n6906 gnd.n6905 585
R4578 gnd.n6903 gnd.n519 585
R4579 gnd.n6902 gnd.n6901 585
R4580 gnd.n6900 gnd.n6899 585
R4581 gnd.n6898 gnd.n6897 585
R4582 gnd.n6896 gnd.n6895 585
R4583 gnd.n6894 gnd.n6893 585
R4584 gnd.n6892 gnd.n6891 585
R4585 gnd.n6890 gnd.n6889 585
R4586 gnd.n6888 gnd.n6887 585
R4587 gnd.n6886 gnd.n6885 585
R4588 gnd.n6884 gnd.n6883 585
R4589 gnd.n6882 gnd.n6881 585
R4590 gnd.n6880 gnd.n6879 585
R4591 gnd.n6877 gnd.n6876 585
R4592 gnd.n6875 gnd.n6874 585
R4593 gnd.n6873 gnd.n6872 585
R4594 gnd.n6871 gnd.n6870 585
R4595 gnd.n6869 gnd.n6868 585
R4596 gnd.n6867 gnd.n6866 585
R4597 gnd.n6865 gnd.n6864 585
R4598 gnd.n6863 gnd.n6862 585
R4599 gnd.n6861 gnd.n6860 585
R4600 gnd.n6859 gnd.n6858 585
R4601 gnd.n6857 gnd.n6856 585
R4602 gnd.n6855 gnd.n6854 585
R4603 gnd.n6853 gnd.n6852 585
R4604 gnd.n6851 gnd.n6850 585
R4605 gnd.n6849 gnd.n6848 585
R4606 gnd.n6847 gnd.n6846 585
R4607 gnd.n6845 gnd.n6844 585
R4608 gnd.n6843 gnd.n6842 585
R4609 gnd.n6841 gnd.n557 585
R4610 gnd.n561 gnd.n558 585
R4611 gnd.n6837 gnd.n6836 585
R4612 gnd.n196 gnd.n195 585
R4613 gnd.n7361 gnd.n191 585
R4614 gnd.n7363 gnd.n7362 585
R4615 gnd.n7365 gnd.n189 585
R4616 gnd.n7367 gnd.n7366 585
R4617 gnd.n7368 gnd.n184 585
R4618 gnd.n7370 gnd.n7369 585
R4619 gnd.n7372 gnd.n182 585
R4620 gnd.n7374 gnd.n7373 585
R4621 gnd.n7375 gnd.n177 585
R4622 gnd.n7377 gnd.n7376 585
R4623 gnd.n7379 gnd.n175 585
R4624 gnd.n7381 gnd.n7380 585
R4625 gnd.n7382 gnd.n170 585
R4626 gnd.n7384 gnd.n7383 585
R4627 gnd.n7386 gnd.n168 585
R4628 gnd.n7388 gnd.n7387 585
R4629 gnd.n7389 gnd.n163 585
R4630 gnd.n7391 gnd.n7390 585
R4631 gnd.n7393 gnd.n161 585
R4632 gnd.n7395 gnd.n7394 585
R4633 gnd.n7399 gnd.n156 585
R4634 gnd.n7401 gnd.n7400 585
R4635 gnd.n7403 gnd.n154 585
R4636 gnd.n7405 gnd.n7404 585
R4637 gnd.n7406 gnd.n149 585
R4638 gnd.n7408 gnd.n7407 585
R4639 gnd.n7410 gnd.n147 585
R4640 gnd.n7412 gnd.n7411 585
R4641 gnd.n7413 gnd.n142 585
R4642 gnd.n7415 gnd.n7414 585
R4643 gnd.n7417 gnd.n140 585
R4644 gnd.n7419 gnd.n7418 585
R4645 gnd.n7420 gnd.n135 585
R4646 gnd.n7422 gnd.n7421 585
R4647 gnd.n7424 gnd.n133 585
R4648 gnd.n7426 gnd.n7425 585
R4649 gnd.n7427 gnd.n131 585
R4650 gnd.n7428 gnd.n127 585
R4651 gnd.n127 gnd.n124 585
R4652 gnd.n7357 gnd.n123 585
R4653 gnd.n7433 gnd.n123 585
R4654 gnd.n7356 gnd.n7355 585
R4655 gnd.n7355 gnd.n122 585
R4656 gnd.n7354 gnd.n200 585
R4657 gnd.n7354 gnd.n7353 585
R4658 gnd.n7121 gnd.n201 585
R4659 gnd.n202 gnd.n201 585
R4660 gnd.n7122 gnd.n210 585
R4661 gnd.n7345 gnd.n210 585
R4662 gnd.n7124 gnd.n7123 585
R4663 gnd.n7123 gnd.n209 585
R4664 gnd.n7125 gnd.n219 585
R4665 gnd.n7269 gnd.n219 585
R4666 gnd.n7127 gnd.n7126 585
R4667 gnd.n7126 gnd.n228 585
R4668 gnd.n7128 gnd.n226 585
R4669 gnd.n7261 gnd.n226 585
R4670 gnd.n7130 gnd.n7129 585
R4671 gnd.n7129 gnd.n225 585
R4672 gnd.n7131 gnd.n235 585
R4673 gnd.n7253 gnd.n235 585
R4674 gnd.n7133 gnd.n7132 585
R4675 gnd.n7132 gnd.n234 585
R4676 gnd.n7134 gnd.n242 585
R4677 gnd.n7245 gnd.n242 585
R4678 gnd.n7136 gnd.n7135 585
R4679 gnd.n7135 gnd.n250 585
R4680 gnd.n7137 gnd.n249 585
R4681 gnd.n7237 gnd.n249 585
R4682 gnd.n7139 gnd.n7138 585
R4683 gnd.n7138 gnd.n259 585
R4684 gnd.n7140 gnd.n257 585
R4685 gnd.n7229 gnd.n257 585
R4686 gnd.n7142 gnd.n7141 585
R4687 gnd.n7141 gnd.n256 585
R4688 gnd.n7143 gnd.n266 585
R4689 gnd.n7221 gnd.n266 585
R4690 gnd.n7145 gnd.n7144 585
R4691 gnd.n7144 gnd.n265 585
R4692 gnd.n7146 gnd.n272 585
R4693 gnd.n7213 gnd.n272 585
R4694 gnd.n7148 gnd.n7147 585
R4695 gnd.n7147 gnd.n280 585
R4696 gnd.n7149 gnd.n279 585
R4697 gnd.n7205 gnd.n279 585
R4698 gnd.n7151 gnd.n7150 585
R4699 gnd.n7150 gnd.n289 585
R4700 gnd.n7152 gnd.n287 585
R4701 gnd.n7197 gnd.n287 585
R4702 gnd.n7154 gnd.n7153 585
R4703 gnd.n7153 gnd.n286 585
R4704 gnd.n7155 gnd.n296 585
R4705 gnd.n7189 gnd.n296 585
R4706 gnd.n7157 gnd.n7156 585
R4707 gnd.n7156 gnd.n295 585
R4708 gnd.n7158 gnd.n324 585
R4709 gnd.n7165 gnd.n324 585
R4710 gnd.n7160 gnd.n7159 585
R4711 gnd.n7161 gnd.n7160 585
R4712 gnd.n332 gnd.n331 585
R4713 gnd.n331 gnd.n330 585
R4714 gnd.n7090 gnd.n7089 585
R4715 gnd.n7089 gnd.n7088 585
R4716 gnd.n335 gnd.n334 585
R4717 gnd.n336 gnd.n335 585
R4718 gnd.n7059 gnd.n339 585
R4719 gnd.n7082 gnd.n339 585
R4720 gnd.n7061 gnd.n7060 585
R4721 gnd.n7062 gnd.n7061 585
R4722 gnd.n355 gnd.n309 585
R4723 gnd.n7180 gnd.n309 585
R4724 gnd.n7054 gnd.n350 585
R4725 gnd.n7071 gnd.n350 585
R4726 gnd.n7053 gnd.n7052 585
R4727 gnd.n7052 gnd.n349 585
R4728 gnd.n7051 gnd.n357 585
R4729 gnd.n7051 gnd.n7050 585
R4730 gnd.n6789 gnd.n358 585
R4731 gnd.n7029 gnd.n358 585
R4732 gnd.n6792 gnd.n6791 585
R4733 gnd.n6791 gnd.n6790 585
R4734 gnd.n6793 gnd.n370 585
R4735 gnd.n7041 gnd.n370 585
R4736 gnd.n6794 gnd.n387 585
R4737 gnd.n7019 gnd.n387 585
R4738 gnd.n6795 gnd.n394 585
R4739 gnd.n6998 gnd.n394 585
R4740 gnd.n6797 gnd.n6796 585
R4741 gnd.n6798 gnd.n6797 585
R4742 gnd.n585 gnd.n402 585
R4743 gnd.n6990 gnd.n402 585
R4744 gnd.n6779 gnd.n6778 585
R4745 gnd.n6778 gnd.n6777 585
R4746 gnd.n587 gnd.n413 585
R4747 gnd.n6979 gnd.n413 585
R4748 gnd.n6760 gnd.n6759 585
R4749 gnd.n6759 gnd.n6758 585
R4750 gnd.n6761 gnd.n420 585
R4751 gnd.n6971 gnd.n420 585
R4752 gnd.n6763 gnd.n6762 585
R4753 gnd.n6764 gnd.n6763 585
R4754 gnd.n594 gnd.n429 585
R4755 gnd.n6963 gnd.n429 585
R4756 gnd.n6752 gnd.n6751 585
R4757 gnd.n6751 gnd.n6750 585
R4758 gnd.n6749 gnd.n438 585
R4759 gnd.n6955 gnd.n438 585
R4760 gnd.n6748 gnd.n6747 585
R4761 gnd.n6747 gnd.n6746 585
R4762 gnd.n596 gnd.n447 585
R4763 gnd.n6947 gnd.n447 585
R4764 gnd.n6721 gnd.n6720 585
R4765 gnd.n6720 gnd.n6719 585
R4766 gnd.n6722 gnd.n454 585
R4767 gnd.n6939 gnd.n454 585
R4768 gnd.n6724 gnd.n6723 585
R4769 gnd.n6725 gnd.n6724 585
R4770 gnd.n6701 gnd.n463 585
R4771 gnd.n6931 gnd.n463 585
R4772 gnd.n6712 gnd.n6711 585
R4773 gnd.n6711 gnd.n6710 585
R4774 gnd.n6709 gnd.n472 585
R4775 gnd.n6923 gnd.n472 585
R4776 gnd.n6708 gnd.n6707 585
R4777 gnd.n6707 gnd.n6706 585
R4778 gnd.n6703 gnd.n481 585
R4779 gnd.n6915 gnd.n481 585
R4780 gnd.n6835 gnd.n563 585
R4781 gnd.n6835 gnd.n6834 585
R4782 gnd.n5931 gnd.n5164 585
R4783 gnd.n5164 gnd.n681 585
R4784 gnd.n5933 gnd.n5932 585
R4785 gnd.n5934 gnd.n5933 585
R4786 gnd.n5165 gnd.n5163 585
R4787 gnd.n5163 gnd.n690 585
R4788 gnd.n5802 gnd.n5801 585
R4789 gnd.n5803 gnd.n5802 585
R4790 gnd.n5800 gnd.n5237 585
R4791 gnd.n5796 gnd.n5237 585
R4792 gnd.n5799 gnd.n5798 585
R4793 gnd.n5798 gnd.n5797 585
R4794 gnd.n5239 gnd.n5238 585
R4795 gnd.n5239 gnd.n696 585
R4796 gnd.n5787 gnd.n5786 585
R4797 gnd.n5788 gnd.n5787 585
R4798 gnd.n5785 gnd.n5244 585
R4799 gnd.n5244 gnd.n705 585
R4800 gnd.n5784 gnd.n5783 585
R4801 gnd.n5783 gnd.n703 585
R4802 gnd.n5782 gnd.n5245 585
R4803 gnd.n5782 gnd.n5781 585
R4804 gnd.n5770 gnd.n5246 585
R4805 gnd.n5246 gnd.n712 585
R4806 gnd.n5772 gnd.n5771 585
R4807 gnd.n5773 gnd.n5772 585
R4808 gnd.n5769 gnd.n5253 585
R4809 gnd.n5253 gnd.n5252 585
R4810 gnd.n5768 gnd.n5767 585
R4811 gnd.n5767 gnd.n720 585
R4812 gnd.n5766 gnd.n5254 585
R4813 gnd.n5766 gnd.n718 585
R4814 gnd.n5765 gnd.n5256 585
R4815 gnd.n5765 gnd.n5764 585
R4816 gnd.n5751 gnd.n5255 585
R4817 gnd.n5255 gnd.n726 585
R4818 gnd.n5753 gnd.n5752 585
R4819 gnd.n5754 gnd.n5753 585
R4820 gnd.n5750 gnd.n5262 585
R4821 gnd.n5262 gnd.t151 585
R4822 gnd.n5749 gnd.n5748 585
R4823 gnd.n5748 gnd.n733 585
R4824 gnd.n5747 gnd.n5263 585
R4825 gnd.n5747 gnd.n5746 585
R4826 gnd.n5734 gnd.n5264 585
R4827 gnd.n5266 gnd.n5264 585
R4828 gnd.n5735 gnd.n5273 585
R4829 gnd.n5273 gnd.n740 585
R4830 gnd.n5737 gnd.n5736 585
R4831 gnd.n5738 gnd.n5737 585
R4832 gnd.n5733 gnd.n5272 585
R4833 gnd.n5272 gnd.n749 585
R4834 gnd.n5732 gnd.n5731 585
R4835 gnd.n5731 gnd.n747 585
R4836 gnd.n5730 gnd.n5274 585
R4837 gnd.n5730 gnd.n5729 585
R4838 gnd.n5716 gnd.n5275 585
R4839 gnd.n5275 gnd.n757 585
R4840 gnd.n5717 gnd.n5283 585
R4841 gnd.n5283 gnd.n755 585
R4842 gnd.n5719 gnd.n5718 585
R4843 gnd.n5720 gnd.n5719 585
R4844 gnd.n5715 gnd.n5282 585
R4845 gnd.n5282 gnd.n765 585
R4846 gnd.n5714 gnd.n5713 585
R4847 gnd.n5713 gnd.n763 585
R4848 gnd.n5712 gnd.n5284 585
R4849 gnd.n5712 gnd.n5711 585
R4850 gnd.n5698 gnd.n5285 585
R4851 gnd.n5285 gnd.n773 585
R4852 gnd.n5699 gnd.n5294 585
R4853 gnd.n5294 gnd.n771 585
R4854 gnd.n5701 gnd.n5700 585
R4855 gnd.n5702 gnd.n5701 585
R4856 gnd.n5697 gnd.n5293 585
R4857 gnd.n5293 gnd.n5292 585
R4858 gnd.n5696 gnd.n5695 585
R4859 gnd.n5695 gnd.n779 585
R4860 gnd.n5694 gnd.n5295 585
R4861 gnd.n5694 gnd.n5693 585
R4862 gnd.n5680 gnd.n5296 585
R4863 gnd.n5296 gnd.n788 585
R4864 gnd.n5681 gnd.n5304 585
R4865 gnd.n5304 gnd.n786 585
R4866 gnd.n5683 gnd.n5682 585
R4867 gnd.n5684 gnd.n5683 585
R4868 gnd.n5679 gnd.n5303 585
R4869 gnd.n5303 gnd.n795 585
R4870 gnd.n5678 gnd.n5677 585
R4871 gnd.n5677 gnd.n5676 585
R4872 gnd.n5306 gnd.n5305 585
R4873 gnd.n5308 gnd.n5306 585
R4874 gnd.n5663 gnd.n5662 585
R4875 gnd.n5662 gnd.n803 585
R4876 gnd.n5664 gnd.n5315 585
R4877 gnd.n5315 gnd.n801 585
R4878 gnd.n5666 gnd.n5665 585
R4879 gnd.n5667 gnd.n5666 585
R4880 gnd.n5661 gnd.n5314 585
R4881 gnd.n5314 gnd.n811 585
R4882 gnd.n5660 gnd.n5659 585
R4883 gnd.n5659 gnd.n809 585
R4884 gnd.n5658 gnd.n5316 585
R4885 gnd.n5658 gnd.n5657 585
R4886 gnd.n5643 gnd.n5317 585
R4887 gnd.n5317 gnd.n819 585
R4888 gnd.n5644 gnd.n5324 585
R4889 gnd.n5324 gnd.n817 585
R4890 gnd.n5646 gnd.n5645 585
R4891 gnd.n5647 gnd.n5646 585
R4892 gnd.n5642 gnd.n5323 585
R4893 gnd.n5323 gnd.n827 585
R4894 gnd.n5641 gnd.n5640 585
R4895 gnd.n5640 gnd.n825 585
R4896 gnd.n5639 gnd.n5325 585
R4897 gnd.n5639 gnd.n5638 585
R4898 gnd.n5626 gnd.n5326 585
R4899 gnd.n5326 gnd.n834 585
R4900 gnd.n5628 gnd.n5627 585
R4901 gnd.n5629 gnd.n5628 585
R4902 gnd.n5625 gnd.n5333 585
R4903 gnd.n5333 gnd.n5332 585
R4904 gnd.n5624 gnd.n5623 585
R4905 gnd.n5623 gnd.n841 585
R4906 gnd.n5622 gnd.n5334 585
R4907 gnd.n5622 gnd.t26 585
R4908 gnd.n5621 gnd.n5336 585
R4909 gnd.n5621 gnd.n5620 585
R4910 gnd.n5607 gnd.n5335 585
R4911 gnd.n5335 gnd.n848 585
R4912 gnd.n5609 gnd.n5608 585
R4913 gnd.n5610 gnd.n5609 585
R4914 gnd.n5606 gnd.n5342 585
R4915 gnd.n5342 gnd.n856 585
R4916 gnd.n5605 gnd.n5604 585
R4917 gnd.n5604 gnd.n854 585
R4918 gnd.n5603 gnd.n5343 585
R4919 gnd.n5603 gnd.n5602 585
R4920 gnd.n5590 gnd.n5344 585
R4921 gnd.n5346 gnd.n5344 585
R4922 gnd.n5591 gnd.n5353 585
R4923 gnd.n5353 gnd.n862 585
R4924 gnd.n5593 gnd.n5592 585
R4925 gnd.n5594 gnd.n5593 585
R4926 gnd.n5589 gnd.n5352 585
R4927 gnd.n5352 gnd.n871 585
R4928 gnd.n5588 gnd.n5587 585
R4929 gnd.n5587 gnd.n869 585
R4930 gnd.n5586 gnd.n5354 585
R4931 gnd.n5586 gnd.n5585 585
R4932 gnd.n5572 gnd.n5355 585
R4933 gnd.n5355 gnd.n879 585
R4934 gnd.n5573 gnd.n5363 585
R4935 gnd.n5363 gnd.n877 585
R4936 gnd.n5575 gnd.n5574 585
R4937 gnd.n5576 gnd.n5575 585
R4938 gnd.n5571 gnd.n5362 585
R4939 gnd.n5362 gnd.n887 585
R4940 gnd.n5570 gnd.n5569 585
R4941 gnd.n5569 gnd.n885 585
R4942 gnd.n5568 gnd.n5364 585
R4943 gnd.n5568 gnd.n5567 585
R4944 gnd.n5429 gnd.n5365 585
R4945 gnd.n5367 gnd.n5365 585
R4946 gnd.n5432 gnd.n5431 585
R4947 gnd.n5434 gnd.n5408 585
R4948 gnd.n5435 gnd.n5407 585
R4949 gnd.n5435 gnd.n893 585
R4950 gnd.n5438 gnd.n5437 585
R4951 gnd.n5439 gnd.n5406 585
R4952 gnd.n5441 gnd.n5440 585
R4953 gnd.n5443 gnd.n5405 585
R4954 gnd.n5446 gnd.n5445 585
R4955 gnd.n5447 gnd.n5404 585
R4956 gnd.n5449 gnd.n5448 585
R4957 gnd.n5451 gnd.n5403 585
R4958 gnd.n5454 gnd.n5453 585
R4959 gnd.n5455 gnd.n5402 585
R4960 gnd.n5457 gnd.n5456 585
R4961 gnd.n5459 gnd.n5401 585
R4962 gnd.n5462 gnd.n5461 585
R4963 gnd.n5463 gnd.n5400 585
R4964 gnd.n5465 gnd.n5464 585
R4965 gnd.n5467 gnd.n5399 585
R4966 gnd.n5470 gnd.n5469 585
R4967 gnd.n5471 gnd.n5398 585
R4968 gnd.n5473 gnd.n5472 585
R4969 gnd.n5475 gnd.n5397 585
R4970 gnd.n5478 gnd.n5477 585
R4971 gnd.n5479 gnd.n5396 585
R4972 gnd.n5481 gnd.n5480 585
R4973 gnd.n5483 gnd.n5395 585
R4974 gnd.n5486 gnd.n5485 585
R4975 gnd.n5487 gnd.n5392 585
R4976 gnd.n5490 gnd.n5489 585
R4977 gnd.n5492 gnd.n5391 585
R4978 gnd.n5493 gnd.n5389 585
R4979 gnd.n5496 gnd.n5388 585
R4980 gnd.n5498 gnd.n5497 585
R4981 gnd.n5500 gnd.n5387 585
R4982 gnd.n5503 gnd.n5502 585
R4983 gnd.n5505 gnd.n5384 585
R4984 gnd.n5507 gnd.n5506 585
R4985 gnd.n5509 gnd.n5383 585
R4986 gnd.n5512 gnd.n5511 585
R4987 gnd.n5513 gnd.n5382 585
R4988 gnd.n5515 gnd.n5514 585
R4989 gnd.n5517 gnd.n5381 585
R4990 gnd.n5520 gnd.n5519 585
R4991 gnd.n5521 gnd.n5380 585
R4992 gnd.n5523 gnd.n5522 585
R4993 gnd.n5525 gnd.n5379 585
R4994 gnd.n5528 gnd.n5527 585
R4995 gnd.n5529 gnd.n5378 585
R4996 gnd.n5531 gnd.n5530 585
R4997 gnd.n5533 gnd.n5377 585
R4998 gnd.n5536 gnd.n5535 585
R4999 gnd.n5537 gnd.n5376 585
R5000 gnd.n5539 gnd.n5538 585
R5001 gnd.n5541 gnd.n5375 585
R5002 gnd.n5544 gnd.n5543 585
R5003 gnd.n5545 gnd.n5374 585
R5004 gnd.n5547 gnd.n5546 585
R5005 gnd.n5549 gnd.n5373 585
R5006 gnd.n5552 gnd.n5551 585
R5007 gnd.n5553 gnd.n5372 585
R5008 gnd.n5555 gnd.n5554 585
R5009 gnd.n5557 gnd.n5371 585
R5010 gnd.n5558 gnd.n5370 585
R5011 gnd.n5561 gnd.n5560 585
R5012 gnd.n5812 gnd.n5811 585
R5013 gnd.n5813 gnd.n5234 585
R5014 gnd.n5815 gnd.n5814 585
R5015 gnd.n5817 gnd.n5232 585
R5016 gnd.n5819 gnd.n5818 585
R5017 gnd.n5820 gnd.n5231 585
R5018 gnd.n5822 gnd.n5821 585
R5019 gnd.n5824 gnd.n5229 585
R5020 gnd.n5826 gnd.n5825 585
R5021 gnd.n5827 gnd.n5228 585
R5022 gnd.n5829 gnd.n5828 585
R5023 gnd.n5831 gnd.n5226 585
R5024 gnd.n5833 gnd.n5832 585
R5025 gnd.n5834 gnd.n5225 585
R5026 gnd.n5836 gnd.n5835 585
R5027 gnd.n5838 gnd.n5223 585
R5028 gnd.n5840 gnd.n5839 585
R5029 gnd.n5841 gnd.n5222 585
R5030 gnd.n5843 gnd.n5842 585
R5031 gnd.n5845 gnd.n5220 585
R5032 gnd.n5847 gnd.n5846 585
R5033 gnd.n5848 gnd.n5219 585
R5034 gnd.n5850 gnd.n5849 585
R5035 gnd.n5852 gnd.n5217 585
R5036 gnd.n5854 gnd.n5853 585
R5037 gnd.n5855 gnd.n5216 585
R5038 gnd.n5857 gnd.n5856 585
R5039 gnd.n5859 gnd.n5214 585
R5040 gnd.n5861 gnd.n5860 585
R5041 gnd.n5863 gnd.n5211 585
R5042 gnd.n5865 gnd.n5864 585
R5043 gnd.n5867 gnd.n5210 585
R5044 gnd.n5868 gnd.n683 585
R5045 gnd.n5871 gnd.n534 585
R5046 gnd.n5873 gnd.n5872 585
R5047 gnd.n5875 gnd.n5208 585
R5048 gnd.n5877 gnd.n5876 585
R5049 gnd.n5879 gnd.n5205 585
R5050 gnd.n5881 gnd.n5880 585
R5051 gnd.n5883 gnd.n5203 585
R5052 gnd.n5885 gnd.n5884 585
R5053 gnd.n5886 gnd.n5202 585
R5054 gnd.n5888 gnd.n5887 585
R5055 gnd.n5890 gnd.n5200 585
R5056 gnd.n5892 gnd.n5891 585
R5057 gnd.n5893 gnd.n5199 585
R5058 gnd.n5895 gnd.n5894 585
R5059 gnd.n5897 gnd.n5197 585
R5060 gnd.n5899 gnd.n5898 585
R5061 gnd.n5900 gnd.n5196 585
R5062 gnd.n5902 gnd.n5901 585
R5063 gnd.n5904 gnd.n5194 585
R5064 gnd.n5906 gnd.n5905 585
R5065 gnd.n5907 gnd.n5193 585
R5066 gnd.n5909 gnd.n5908 585
R5067 gnd.n5911 gnd.n5191 585
R5068 gnd.n5913 gnd.n5912 585
R5069 gnd.n5914 gnd.n5190 585
R5070 gnd.n5916 gnd.n5915 585
R5071 gnd.n5918 gnd.n5188 585
R5072 gnd.n5920 gnd.n5919 585
R5073 gnd.n5921 gnd.n5187 585
R5074 gnd.n5923 gnd.n5922 585
R5075 gnd.n5925 gnd.n5186 585
R5076 gnd.n5926 gnd.n5185 585
R5077 gnd.n5929 gnd.n5928 585
R5078 gnd.n5810 gnd.n5808 585
R5079 gnd.n5810 gnd.n681 585
R5080 gnd.n5807 gnd.n5162 585
R5081 gnd.n5934 gnd.n5162 585
R5082 gnd.n5806 gnd.n5805 585
R5083 gnd.n5805 gnd.n690 585
R5084 gnd.n5804 gnd.n5235 585
R5085 gnd.n5804 gnd.n5803 585
R5086 gnd.n5792 gnd.n5236 585
R5087 gnd.n5796 gnd.n5236 585
R5088 gnd.n5794 gnd.n5793 585
R5089 gnd.n5797 gnd.n5794 585
R5090 gnd.n5791 gnd.n5240 585
R5091 gnd.n5240 gnd.n696 585
R5092 gnd.n5790 gnd.n5789 585
R5093 gnd.n5789 gnd.n5788 585
R5094 gnd.n5242 gnd.n5241 585
R5095 gnd.n5242 gnd.n705 585
R5096 gnd.n5777 gnd.n5248 585
R5097 gnd.n5248 gnd.n703 585
R5098 gnd.n5779 gnd.n5778 585
R5099 gnd.n5781 gnd.n5779 585
R5100 gnd.n5776 gnd.n5247 585
R5101 gnd.n5247 gnd.n712 585
R5102 gnd.n5775 gnd.n5774 585
R5103 gnd.n5774 gnd.n5773 585
R5104 gnd.n5250 gnd.n5249 585
R5105 gnd.n5252 gnd.n5250 585
R5106 gnd.n5759 gnd.n5758 585
R5107 gnd.n5758 gnd.n720 585
R5108 gnd.n5760 gnd.n5258 585
R5109 gnd.n5258 gnd.n718 585
R5110 gnd.n5762 gnd.n5761 585
R5111 gnd.n5764 gnd.n5762 585
R5112 gnd.n5757 gnd.n5257 585
R5113 gnd.n5257 gnd.n726 585
R5114 gnd.n5756 gnd.n5755 585
R5115 gnd.n5755 gnd.n5754 585
R5116 gnd.n5260 gnd.n5259 585
R5117 gnd.n5260 gnd.t151 585
R5118 gnd.n5743 gnd.n5268 585
R5119 gnd.n5268 gnd.n733 585
R5120 gnd.n5745 gnd.n5744 585
R5121 gnd.n5746 gnd.n5745 585
R5122 gnd.n5742 gnd.n5267 585
R5123 gnd.n5267 gnd.n5266 585
R5124 gnd.n5741 gnd.n5740 585
R5125 gnd.n5740 gnd.n740 585
R5126 gnd.n5739 gnd.n5269 585
R5127 gnd.n5739 gnd.n5738 585
R5128 gnd.n5725 gnd.n5270 585
R5129 gnd.n5270 gnd.n749 585
R5130 gnd.n5726 gnd.n5278 585
R5131 gnd.n5278 gnd.n747 585
R5132 gnd.n5728 gnd.n5727 585
R5133 gnd.n5729 gnd.n5728 585
R5134 gnd.n5724 gnd.n5277 585
R5135 gnd.n5277 gnd.n757 585
R5136 gnd.n5723 gnd.n5722 585
R5137 gnd.n5722 gnd.n755 585
R5138 gnd.n5721 gnd.n5279 585
R5139 gnd.n5721 gnd.n5720 585
R5140 gnd.n5707 gnd.n5280 585
R5141 gnd.n5280 gnd.n765 585
R5142 gnd.n5708 gnd.n5288 585
R5143 gnd.n5288 gnd.n763 585
R5144 gnd.n5710 gnd.n5709 585
R5145 gnd.n5711 gnd.n5710 585
R5146 gnd.n5706 gnd.n5287 585
R5147 gnd.n5287 gnd.n773 585
R5148 gnd.n5705 gnd.n5704 585
R5149 gnd.n5704 gnd.n771 585
R5150 gnd.n5703 gnd.n5289 585
R5151 gnd.n5703 gnd.n5702 585
R5152 gnd.n5689 gnd.n5290 585
R5153 gnd.n5292 gnd.n5290 585
R5154 gnd.n5690 gnd.n5299 585
R5155 gnd.n5299 gnd.n779 585
R5156 gnd.n5692 gnd.n5691 585
R5157 gnd.n5693 gnd.n5692 585
R5158 gnd.n5688 gnd.n5298 585
R5159 gnd.n5298 gnd.n788 585
R5160 gnd.n5687 gnd.n5686 585
R5161 gnd.n5686 gnd.n786 585
R5162 gnd.n5685 gnd.n5300 585
R5163 gnd.n5685 gnd.n5684 585
R5164 gnd.n5673 gnd.n5301 585
R5165 gnd.n5301 gnd.n795 585
R5166 gnd.n5675 gnd.n5674 585
R5167 gnd.n5676 gnd.n5675 585
R5168 gnd.n5672 gnd.n5309 585
R5169 gnd.n5309 gnd.n5308 585
R5170 gnd.n5671 gnd.n5670 585
R5171 gnd.n5670 gnd.n803 585
R5172 gnd.n5669 gnd.n5310 585
R5173 gnd.n5669 gnd.n801 585
R5174 gnd.n5668 gnd.n5312 585
R5175 gnd.n5668 gnd.n5667 585
R5176 gnd.n5652 gnd.n5311 585
R5177 gnd.n5311 gnd.n811 585
R5178 gnd.n5653 gnd.n5319 585
R5179 gnd.n5319 gnd.n809 585
R5180 gnd.n5655 gnd.n5654 585
R5181 gnd.n5657 gnd.n5655 585
R5182 gnd.n5651 gnd.n5318 585
R5183 gnd.n5318 gnd.n819 585
R5184 gnd.n5650 gnd.n5649 585
R5185 gnd.n5649 gnd.n817 585
R5186 gnd.n5648 gnd.n5320 585
R5187 gnd.n5648 gnd.n5647 585
R5188 gnd.n5633 gnd.n5321 585
R5189 gnd.n5321 gnd.n827 585
R5190 gnd.n5634 gnd.n5328 585
R5191 gnd.n5328 gnd.n825 585
R5192 gnd.n5636 gnd.n5635 585
R5193 gnd.n5638 gnd.n5636 585
R5194 gnd.n5632 gnd.n5327 585
R5195 gnd.n5327 gnd.n834 585
R5196 gnd.n5631 gnd.n5630 585
R5197 gnd.n5630 gnd.n5629 585
R5198 gnd.n5330 gnd.n5329 585
R5199 gnd.n5332 gnd.n5330 585
R5200 gnd.n5615 gnd.n5614 585
R5201 gnd.n5614 gnd.n841 585
R5202 gnd.n5616 gnd.n5338 585
R5203 gnd.n5338 gnd.t26 585
R5204 gnd.n5618 gnd.n5617 585
R5205 gnd.n5620 gnd.n5618 585
R5206 gnd.n5613 gnd.n5337 585
R5207 gnd.n5337 gnd.n848 585
R5208 gnd.n5612 gnd.n5611 585
R5209 gnd.n5611 gnd.n5610 585
R5210 gnd.n5340 gnd.n5339 585
R5211 gnd.n5340 gnd.n856 585
R5212 gnd.n5599 gnd.n5348 585
R5213 gnd.n5348 gnd.n854 585
R5214 gnd.n5601 gnd.n5600 585
R5215 gnd.n5602 gnd.n5601 585
R5216 gnd.n5598 gnd.n5347 585
R5217 gnd.n5347 gnd.n5346 585
R5218 gnd.n5597 gnd.n5596 585
R5219 gnd.n5596 gnd.n862 585
R5220 gnd.n5595 gnd.n5349 585
R5221 gnd.n5595 gnd.n5594 585
R5222 gnd.n5581 gnd.n5350 585
R5223 gnd.n5350 gnd.n871 585
R5224 gnd.n5582 gnd.n5358 585
R5225 gnd.n5358 gnd.n869 585
R5226 gnd.n5584 gnd.n5583 585
R5227 gnd.n5585 gnd.n5584 585
R5228 gnd.n5580 gnd.n5357 585
R5229 gnd.n5357 gnd.n879 585
R5230 gnd.n5579 gnd.n5578 585
R5231 gnd.n5578 gnd.n877 585
R5232 gnd.n5577 gnd.n5359 585
R5233 gnd.n5577 gnd.n5576 585
R5234 gnd.n5563 gnd.n5360 585
R5235 gnd.n5360 gnd.n887 585
R5236 gnd.n5564 gnd.n5369 585
R5237 gnd.n5369 gnd.n885 585
R5238 gnd.n5566 gnd.n5565 585
R5239 gnd.n5567 gnd.n5566 585
R5240 gnd.n5562 gnd.n5368 585
R5241 gnd.n5368 gnd.n5367 585
R5242 gnd.n2763 gnd.n1476 585
R5243 gnd.n1476 gnd.n1200 585
R5244 gnd.n7080 gnd.n7079 585
R5245 gnd.n7081 gnd.n7080 585
R5246 gnd.n7076 gnd.n343 585
R5247 gnd.n343 gnd.n311 585
R5248 gnd.n7075 gnd.n7074 585
R5249 gnd.n7074 gnd.n308 585
R5250 gnd.n7073 gnd.n346 585
R5251 gnd.n7073 gnd.n7072 585
R5252 gnd.n7010 gnd.n348 585
R5253 gnd.n361 gnd.n348 585
R5254 gnd.n7012 gnd.n7011 585
R5255 gnd.n7012 gnd.n359 585
R5256 gnd.n7014 gnd.n7013 585
R5257 gnd.n7013 gnd.n379 585
R5258 gnd.n7015 gnd.n389 585
R5259 gnd.n389 gnd.n372 585
R5260 gnd.n7017 gnd.n7016 585
R5261 gnd.n7018 gnd.n7017 585
R5262 gnd.n390 gnd.n388 585
R5263 gnd.n388 gnd.n386 585
R5264 gnd.n7001 gnd.n7000 585
R5265 gnd.n7000 gnd.n6999 585
R5266 gnd.n393 gnd.n392 585
R5267 gnd.n404 gnd.n393 585
R5268 gnd.n6773 gnd.n589 585
R5269 gnd.n589 gnd.n401 585
R5270 gnd.n6775 gnd.n6774 585
R5271 gnd.n6776 gnd.n6775 585
R5272 gnd.n590 gnd.n588 585
R5273 gnd.n588 gnd.n412 585
R5274 gnd.n6768 gnd.n6767 585
R5275 gnd.n6767 gnd.n422 585
R5276 gnd.n6766 gnd.n592 585
R5277 gnd.n6766 gnd.n6765 585
R5278 gnd.n6737 gnd.n593 585
R5279 gnd.n593 gnd.n431 585
R5280 gnd.n6739 gnd.n6738 585
R5281 gnd.n6739 gnd.n428 585
R5282 gnd.n6741 gnd.n6740 585
R5283 gnd.n6740 gnd.n440 585
R5284 gnd.n6742 gnd.n599 585
R5285 gnd.n599 gnd.n437 585
R5286 gnd.n6744 gnd.n6743 585
R5287 gnd.n6745 gnd.n6744 585
R5288 gnd.n600 gnd.n598 585
R5289 gnd.n598 gnd.n446 585
R5290 gnd.n6729 gnd.n6728 585
R5291 gnd.n6728 gnd.n456 585
R5292 gnd.n6727 gnd.n602 585
R5293 gnd.n6727 gnd.n6726 585
R5294 gnd.n6700 gnd.n6699 585
R5295 gnd.n6700 gnd.n465 585
R5296 gnd.n604 gnd.n603 585
R5297 gnd.n603 gnd.n462 585
R5298 gnd.n6695 gnd.n6694 585
R5299 gnd.n6694 gnd.n474 585
R5300 gnd.n6693 gnd.n606 585
R5301 gnd.n6693 gnd.n471 585
R5302 gnd.n6692 gnd.n6691 585
R5303 gnd.n6692 gnd.n483 585
R5304 gnd.n608 gnd.n607 585
R5305 gnd.n607 gnd.n480 585
R5306 gnd.n6687 gnd.n6686 585
R5307 gnd.n6686 gnd.n564 585
R5308 gnd.n6685 gnd.n610 585
R5309 gnd.n6685 gnd.n518 585
R5310 gnd.n6684 gnd.n6683 585
R5311 gnd.n6684 gnd.n489 585
R5312 gnd.n612 gnd.n611 585
R5313 gnd.n6676 gnd.n611 585
R5314 gnd.n6679 gnd.n6678 585
R5315 gnd.n6678 gnd.n6677 585
R5316 gnd.n615 gnd.n614 585
R5317 gnd.n616 gnd.n615 585
R5318 gnd.n6665 gnd.n641 585
R5319 gnd.n641 gnd.n639 585
R5320 gnd.n6667 gnd.n6666 585
R5321 gnd.n6668 gnd.n6667 585
R5322 gnd.n642 gnd.n640 585
R5323 gnd.n648 gnd.n640 585
R5324 gnd.n6660 gnd.n6659 585
R5325 gnd.n6659 gnd.n6658 585
R5326 gnd.n645 gnd.n644 585
R5327 gnd.n646 gnd.n645 585
R5328 gnd.n6648 gnd.n6647 585
R5329 gnd.n6649 gnd.n6648 585
R5330 gnd.n657 gnd.n656 585
R5331 gnd.n656 gnd.n654 585
R5332 gnd.n6643 gnd.n6642 585
R5333 gnd.n6642 gnd.n6641 585
R5334 gnd.n660 gnd.n659 585
R5335 gnd.n661 gnd.n660 585
R5336 gnd.n6632 gnd.n6631 585
R5337 gnd.n6633 gnd.n6632 585
R5338 gnd.n671 gnd.n670 585
R5339 gnd.n670 gnd.n668 585
R5340 gnd.n6627 gnd.n6626 585
R5341 gnd.n6626 gnd.n6625 585
R5342 gnd.n674 gnd.n673 585
R5343 gnd.n5937 gnd.n674 585
R5344 gnd.n6616 gnd.n6615 585
R5345 gnd.n6617 gnd.n6616 585
R5346 gnd.n685 gnd.n684 585
R5347 gnd.n5935 gnd.n684 585
R5348 gnd.n6611 gnd.n6610 585
R5349 gnd.n6610 gnd.n6609 585
R5350 gnd.n688 gnd.n687 585
R5351 gnd.n5795 gnd.n688 585
R5352 gnd.n6600 gnd.n6599 585
R5353 gnd.n6601 gnd.n6600 585
R5354 gnd.n699 gnd.n698 585
R5355 gnd.n5243 gnd.n698 585
R5356 gnd.n6595 gnd.n6594 585
R5357 gnd.n6594 gnd.n6593 585
R5358 gnd.n702 gnd.n701 585
R5359 gnd.n5780 gnd.n702 585
R5360 gnd.n6584 gnd.n6583 585
R5361 gnd.n6585 gnd.n6584 585
R5362 gnd.n714 gnd.n713 585
R5363 gnd.n5251 gnd.n713 585
R5364 gnd.n6579 gnd.n6578 585
R5365 gnd.n6578 gnd.n6577 585
R5366 gnd.n717 gnd.n716 585
R5367 gnd.n5763 gnd.n717 585
R5368 gnd.n6568 gnd.n6567 585
R5369 gnd.n6569 gnd.n6568 585
R5370 gnd.n729 gnd.n728 585
R5371 gnd.n5261 gnd.n728 585
R5372 gnd.n6563 gnd.n6562 585
R5373 gnd.n6562 gnd.n6561 585
R5374 gnd.n732 gnd.n731 585
R5375 gnd.n5265 gnd.n732 585
R5376 gnd.n6552 gnd.n6551 585
R5377 gnd.n6553 gnd.n6552 585
R5378 gnd.n743 gnd.n742 585
R5379 gnd.n5271 gnd.n742 585
R5380 gnd.n6547 gnd.n6546 585
R5381 gnd.n6546 gnd.n6545 585
R5382 gnd.n746 gnd.n745 585
R5383 gnd.n5276 gnd.n746 585
R5384 gnd.n6536 gnd.n6535 585
R5385 gnd.n6537 gnd.n6536 585
R5386 gnd.n759 gnd.n758 585
R5387 gnd.n5281 gnd.n758 585
R5388 gnd.n6531 gnd.n6530 585
R5389 gnd.n6530 gnd.n6529 585
R5390 gnd.n762 gnd.n761 585
R5391 gnd.n5286 gnd.n762 585
R5392 gnd.n6520 gnd.n6519 585
R5393 gnd.n6521 gnd.n6520 585
R5394 gnd.n775 gnd.n774 585
R5395 gnd.n5291 gnd.n774 585
R5396 gnd.n6515 gnd.n6514 585
R5397 gnd.n6514 gnd.n6513 585
R5398 gnd.n778 gnd.n777 585
R5399 gnd.n5297 gnd.n778 585
R5400 gnd.n6504 gnd.n6503 585
R5401 gnd.n6505 gnd.n6504 585
R5402 gnd.n790 gnd.n789 585
R5403 gnd.n5302 gnd.n789 585
R5404 gnd.n6499 gnd.n6498 585
R5405 gnd.n6498 gnd.n6497 585
R5406 gnd.n793 gnd.n792 585
R5407 gnd.n5307 gnd.n793 585
R5408 gnd.n6488 gnd.n6487 585
R5409 gnd.n6489 gnd.n6488 585
R5410 gnd.n805 gnd.n804 585
R5411 gnd.n5313 gnd.n804 585
R5412 gnd.n6483 gnd.n6482 585
R5413 gnd.n6482 gnd.n6481 585
R5414 gnd.n808 gnd.n807 585
R5415 gnd.n5656 gnd.n808 585
R5416 gnd.n6472 gnd.n6471 585
R5417 gnd.n6473 gnd.n6472 585
R5418 gnd.n821 gnd.n820 585
R5419 gnd.n5322 gnd.n820 585
R5420 gnd.n6467 gnd.n6466 585
R5421 gnd.n6466 gnd.n6465 585
R5422 gnd.n824 gnd.n823 585
R5423 gnd.n5637 gnd.n824 585
R5424 gnd.n6456 gnd.n6455 585
R5425 gnd.n6457 gnd.n6456 585
R5426 gnd.n836 gnd.n835 585
R5427 gnd.n5331 gnd.n835 585
R5428 gnd.n6451 gnd.n6450 585
R5429 gnd.n6450 gnd.n6449 585
R5430 gnd.n839 gnd.n838 585
R5431 gnd.n5619 gnd.n839 585
R5432 gnd.n6440 gnd.n6439 585
R5433 gnd.n6441 gnd.n6440 585
R5434 gnd.n850 gnd.n849 585
R5435 gnd.n5341 gnd.n849 585
R5436 gnd.n6435 gnd.n6434 585
R5437 gnd.n6434 gnd.n6433 585
R5438 gnd.n853 gnd.n852 585
R5439 gnd.n5345 gnd.n853 585
R5440 gnd.n6424 gnd.n6423 585
R5441 gnd.n6425 gnd.n6424 585
R5442 gnd.n865 gnd.n864 585
R5443 gnd.n5351 gnd.n864 585
R5444 gnd.n6419 gnd.n6418 585
R5445 gnd.n6418 gnd.n6417 585
R5446 gnd.n868 gnd.n867 585
R5447 gnd.n5356 gnd.n868 585
R5448 gnd.n6408 gnd.n6407 585
R5449 gnd.n6409 gnd.n6408 585
R5450 gnd.n881 gnd.n880 585
R5451 gnd.n5361 gnd.n880 585
R5452 gnd.n6403 gnd.n6402 585
R5453 gnd.n6402 gnd.n6401 585
R5454 gnd.n884 gnd.n883 585
R5455 gnd.n5366 gnd.n884 585
R5456 gnd.n6392 gnd.n6391 585
R5457 gnd.n6393 gnd.n6392 585
R5458 gnd.n896 gnd.n895 585
R5459 gnd.n901 gnd.n895 585
R5460 gnd.n6387 gnd.n6386 585
R5461 gnd.n6386 gnd.n6385 585
R5462 gnd.n899 gnd.n898 585
R5463 gnd.n909 gnd.n899 585
R5464 gnd.n6376 gnd.n6375 585
R5465 gnd.n6377 gnd.n6376 585
R5466 gnd.n911 gnd.n910 585
R5467 gnd.n910 gnd.n907 585
R5468 gnd.n6371 gnd.n6370 585
R5469 gnd.n6370 gnd.n6369 585
R5470 gnd.n914 gnd.n913 585
R5471 gnd.n923 gnd.n914 585
R5472 gnd.n6360 gnd.n6359 585
R5473 gnd.n6361 gnd.n6360 585
R5474 gnd.n925 gnd.n924 585
R5475 gnd.n924 gnd.n921 585
R5476 gnd.n6355 gnd.n6354 585
R5477 gnd.n6354 gnd.n6353 585
R5478 gnd.n928 gnd.n927 585
R5479 gnd.n929 gnd.n928 585
R5480 gnd.n6344 gnd.n6343 585
R5481 gnd.n6345 gnd.n6344 585
R5482 gnd.n939 gnd.n938 585
R5483 gnd.n938 gnd.n936 585
R5484 gnd.n6339 gnd.n6338 585
R5485 gnd.n6338 gnd.n6337 585
R5486 gnd.n942 gnd.n941 585
R5487 gnd.n6336 gnd.n942 585
R5488 gnd.n4770 gnd.n4769 585
R5489 gnd.n4769 gnd.n943 585
R5490 gnd.n4771 gnd.n4764 585
R5491 gnd.n4764 gnd.n4763 585
R5492 gnd.n4774 gnd.n4772 585
R5493 gnd.n4774 gnd.n4773 585
R5494 gnd.n4775 gnd.n4762 585
R5495 gnd.n4775 gnd.n984 585
R5496 gnd.n4777 gnd.n4776 585
R5497 gnd.n4776 gnd.n982 585
R5498 gnd.n4778 gnd.n4757 585
R5499 gnd.n4757 gnd.n1061 585
R5500 gnd.n4780 gnd.n4779 585
R5501 gnd.n4780 gnd.n1070 585
R5502 gnd.n4781 gnd.n4756 585
R5503 gnd.n4781 gnd.n1067 585
R5504 gnd.n4783 gnd.n4782 585
R5505 gnd.n4782 gnd.n1080 585
R5506 gnd.n4784 gnd.n1247 585
R5507 gnd.n1247 gnd.n1077 585
R5508 gnd.n4786 gnd.n4785 585
R5509 gnd.n4787 gnd.n4786 585
R5510 gnd.n1248 gnd.n1246 585
R5511 gnd.n1246 gnd.n1086 585
R5512 gnd.n4750 gnd.n4749 585
R5513 gnd.n4749 gnd.n1096 585
R5514 gnd.n4748 gnd.n1250 585
R5515 gnd.n4748 gnd.n4747 585
R5516 gnd.n4719 gnd.n1251 585
R5517 gnd.n1251 gnd.n1105 585
R5518 gnd.n4721 gnd.n4720 585
R5519 gnd.n4721 gnd.n1102 585
R5520 gnd.n4723 gnd.n4722 585
R5521 gnd.n4722 gnd.n1114 585
R5522 gnd.n4724 gnd.n1257 585
R5523 gnd.n1257 gnd.n1111 585
R5524 gnd.n4726 gnd.n4725 585
R5525 gnd.n4727 gnd.n4726 585
R5526 gnd.n1258 gnd.n1256 585
R5527 gnd.n1256 gnd.n1120 585
R5528 gnd.n4711 gnd.n4710 585
R5529 gnd.n4710 gnd.n1130 585
R5530 gnd.n4709 gnd.n1260 585
R5531 gnd.n4709 gnd.n4708 585
R5532 gnd.n4679 gnd.n1261 585
R5533 gnd.n1261 gnd.n1139 585
R5534 gnd.n4681 gnd.n4680 585
R5535 gnd.n4681 gnd.n1136 585
R5536 gnd.n4683 gnd.n4682 585
R5537 gnd.n4682 gnd.n1148 585
R5538 gnd.n4684 gnd.n4668 585
R5539 gnd.n4668 gnd.n1145 585
R5540 gnd.n4686 gnd.n4685 585
R5541 gnd.n4687 gnd.n4686 585
R5542 gnd.n4669 gnd.n4667 585
R5543 gnd.n4667 gnd.n1154 585
R5544 gnd.n4671 gnd.n1217 585
R5545 gnd.n1217 gnd.n1164 585
R5546 gnd.n4846 gnd.n1216 585
R5547 gnd.n4846 gnd.n4845 585
R5548 gnd.n4848 gnd.n4847 585
R5549 gnd.n4847 gnd.n1173 585
R5550 gnd.n4849 gnd.n1211 585
R5551 gnd.n1211 gnd.n1170 585
R5552 gnd.n4851 gnd.n4850 585
R5553 gnd.n4852 gnd.n4851 585
R5554 gnd.n1212 gnd.n1210 585
R5555 gnd.n1210 gnd.n1207 585
R5556 gnd.n6095 gnd.n6094 585
R5557 gnd.n6094 gnd.n639 585
R5558 gnd.n6096 gnd.n638 585
R5559 gnd.n6668 gnd.n638 585
R5560 gnd.n6097 gnd.n5949 585
R5561 gnd.n5949 gnd.n648 585
R5562 gnd.n5947 gnd.n647 585
R5563 gnd.n6658 gnd.n647 585
R5564 gnd.n6101 gnd.n5946 585
R5565 gnd.n5946 gnd.n646 585
R5566 gnd.n6102 gnd.n655 585
R5567 gnd.n6649 gnd.n655 585
R5568 gnd.n6103 gnd.n5945 585
R5569 gnd.n5945 gnd.n654 585
R5570 gnd.n5943 gnd.n662 585
R5571 gnd.n6641 gnd.n662 585
R5572 gnd.n6107 gnd.n5942 585
R5573 gnd.n5942 gnd.n661 585
R5574 gnd.n6108 gnd.n669 585
R5575 gnd.n6633 gnd.n669 585
R5576 gnd.n6109 gnd.n5941 585
R5577 gnd.n5941 gnd.n668 585
R5578 gnd.n5939 gnd.n675 585
R5579 gnd.n6625 gnd.n675 585
R5580 gnd.n6113 gnd.n5938 585
R5581 gnd.n5938 gnd.n5937 585
R5582 gnd.n6114 gnd.n682 585
R5583 gnd.n6617 gnd.n682 585
R5584 gnd.n6115 gnd.n5936 585
R5585 gnd.n5936 gnd.n5935 585
R5586 gnd.n5160 gnd.n689 585
R5587 gnd.n6609 gnd.n689 585
R5588 gnd.n6119 gnd.n5159 585
R5589 gnd.n5795 gnd.n5159 585
R5590 gnd.n6120 gnd.n697 585
R5591 gnd.n6601 gnd.n697 585
R5592 gnd.n6121 gnd.n5158 585
R5593 gnd.n5243 gnd.n5158 585
R5594 gnd.n5156 gnd.n704 585
R5595 gnd.n6593 gnd.n704 585
R5596 gnd.n6125 gnd.n5155 585
R5597 gnd.n5780 gnd.n5155 585
R5598 gnd.n6126 gnd.n711 585
R5599 gnd.n6585 gnd.n711 585
R5600 gnd.n6127 gnd.n5154 585
R5601 gnd.n5251 gnd.n5154 585
R5602 gnd.n5152 gnd.n719 585
R5603 gnd.n6577 gnd.n719 585
R5604 gnd.n6131 gnd.n5151 585
R5605 gnd.n5763 gnd.n5151 585
R5606 gnd.n6132 gnd.n727 585
R5607 gnd.n6569 gnd.n727 585
R5608 gnd.n6133 gnd.n5150 585
R5609 gnd.n5261 gnd.n5150 585
R5610 gnd.n5148 gnd.n734 585
R5611 gnd.n6561 gnd.n734 585
R5612 gnd.n6137 gnd.n5147 585
R5613 gnd.n5265 gnd.n5147 585
R5614 gnd.n6138 gnd.n741 585
R5615 gnd.n6553 gnd.n741 585
R5616 gnd.n6139 gnd.n5146 585
R5617 gnd.n5271 gnd.n5146 585
R5618 gnd.n5144 gnd.n748 585
R5619 gnd.n6545 gnd.n748 585
R5620 gnd.n6143 gnd.n5143 585
R5621 gnd.n5276 gnd.n5143 585
R5622 gnd.n6144 gnd.n756 585
R5623 gnd.n6537 gnd.n756 585
R5624 gnd.n6145 gnd.n5142 585
R5625 gnd.n5281 gnd.n5142 585
R5626 gnd.n5140 gnd.n764 585
R5627 gnd.n6529 gnd.n764 585
R5628 gnd.n6149 gnd.n5139 585
R5629 gnd.n5286 gnd.n5139 585
R5630 gnd.n6150 gnd.n772 585
R5631 gnd.n6521 gnd.n772 585
R5632 gnd.n6151 gnd.n5138 585
R5633 gnd.n5291 gnd.n5138 585
R5634 gnd.n5136 gnd.n780 585
R5635 gnd.n6513 gnd.n780 585
R5636 gnd.n6155 gnd.n5135 585
R5637 gnd.n5297 gnd.n5135 585
R5638 gnd.n6156 gnd.n787 585
R5639 gnd.n6505 gnd.n787 585
R5640 gnd.n6157 gnd.n5134 585
R5641 gnd.n5302 gnd.n5134 585
R5642 gnd.n5132 gnd.n794 585
R5643 gnd.n6497 gnd.n794 585
R5644 gnd.n6161 gnd.n5131 585
R5645 gnd.n5307 gnd.n5131 585
R5646 gnd.n6162 gnd.n802 585
R5647 gnd.n6489 gnd.n802 585
R5648 gnd.n6163 gnd.n5130 585
R5649 gnd.n5313 gnd.n5130 585
R5650 gnd.n5128 gnd.n810 585
R5651 gnd.n6481 gnd.n810 585
R5652 gnd.n6167 gnd.n5127 585
R5653 gnd.n5656 gnd.n5127 585
R5654 gnd.n6168 gnd.n818 585
R5655 gnd.n6473 gnd.n818 585
R5656 gnd.n6169 gnd.n5126 585
R5657 gnd.n5322 gnd.n5126 585
R5658 gnd.n5124 gnd.n826 585
R5659 gnd.n6465 gnd.n826 585
R5660 gnd.n6173 gnd.n5123 585
R5661 gnd.n5637 gnd.n5123 585
R5662 gnd.n6174 gnd.n833 585
R5663 gnd.n6457 gnd.n833 585
R5664 gnd.n6175 gnd.n5122 585
R5665 gnd.n5331 gnd.n5122 585
R5666 gnd.n5120 gnd.n840 585
R5667 gnd.n6449 gnd.n840 585
R5668 gnd.n6179 gnd.n5119 585
R5669 gnd.n5619 gnd.n5119 585
R5670 gnd.n6180 gnd.n847 585
R5671 gnd.n6441 gnd.n847 585
R5672 gnd.n6181 gnd.n5118 585
R5673 gnd.n5341 gnd.n5118 585
R5674 gnd.n5116 gnd.n855 585
R5675 gnd.n6433 gnd.n855 585
R5676 gnd.n6185 gnd.n5115 585
R5677 gnd.n5345 gnd.n5115 585
R5678 gnd.n6186 gnd.n863 585
R5679 gnd.n6425 gnd.n863 585
R5680 gnd.n6187 gnd.n5114 585
R5681 gnd.n5351 gnd.n5114 585
R5682 gnd.n5112 gnd.n870 585
R5683 gnd.n6417 gnd.n870 585
R5684 gnd.n6191 gnd.n5111 585
R5685 gnd.n5356 gnd.n5111 585
R5686 gnd.n6192 gnd.n878 585
R5687 gnd.n6409 gnd.n878 585
R5688 gnd.n6193 gnd.n5110 585
R5689 gnd.n5361 gnd.n5110 585
R5690 gnd.n5108 gnd.n886 585
R5691 gnd.n6401 gnd.n886 585
R5692 gnd.n6197 gnd.n5107 585
R5693 gnd.n5366 gnd.n5107 585
R5694 gnd.n6198 gnd.n894 585
R5695 gnd.n6393 gnd.n894 585
R5696 gnd.n6199 gnd.n5106 585
R5697 gnd.n5106 gnd.n901 585
R5698 gnd.n5104 gnd.n900 585
R5699 gnd.n6385 gnd.n900 585
R5700 gnd.n6203 gnd.n5103 585
R5701 gnd.n5103 gnd.n909 585
R5702 gnd.n6204 gnd.n908 585
R5703 gnd.n6377 gnd.n908 585
R5704 gnd.n6205 gnd.n5102 585
R5705 gnd.n5102 gnd.n907 585
R5706 gnd.n5100 gnd.n915 585
R5707 gnd.n6369 gnd.n915 585
R5708 gnd.n6209 gnd.n5099 585
R5709 gnd.n5099 gnd.n923 585
R5710 gnd.n6210 gnd.n922 585
R5711 gnd.n6361 gnd.n922 585
R5712 gnd.n6211 gnd.n5098 585
R5713 gnd.n5098 gnd.n921 585
R5714 gnd.n5096 gnd.n930 585
R5715 gnd.n6353 gnd.n930 585
R5716 gnd.n6215 gnd.n5095 585
R5717 gnd.n5095 gnd.n929 585
R5718 gnd.n6216 gnd.n937 585
R5719 gnd.n6345 gnd.n937 585
R5720 gnd.n6217 gnd.n5094 585
R5721 gnd.n5094 gnd.n936 585
R5722 gnd.n5093 gnd.n5092 585
R5723 gnd.n5091 gnd.n4992 585
R5724 gnd.n4994 gnd.n4993 585
R5725 gnd.n5084 gnd.n5008 585
R5726 gnd.n5083 gnd.n5009 585
R5727 gnd.n5018 gnd.n5010 585
R5728 gnd.n5076 gnd.n5019 585
R5729 gnd.n5075 gnd.n5020 585
R5730 gnd.n5022 gnd.n5021 585
R5731 gnd.n5068 gnd.n5031 585
R5732 gnd.n5067 gnd.n5032 585
R5733 gnd.n5041 gnd.n5033 585
R5734 gnd.n5060 gnd.n5042 585
R5735 gnd.n5059 gnd.n5043 585
R5736 gnd.n5045 gnd.n5044 585
R5737 gnd.n973 gnd.n972 585
R5738 gnd.n6308 gnd.n974 585
R5739 gnd.n6310 gnd.n6309 585
R5740 gnd.n6312 gnd.n6311 585
R5741 gnd.n968 gnd.n967 585
R5742 gnd.n6317 gnd.n969 585
R5743 gnd.n6319 gnd.n6318 585
R5744 gnd.n6321 gnd.n6320 585
R5745 gnd.n964 gnd.n963 585
R5746 gnd.n6325 gnd.n965 585
R5747 gnd.n6328 gnd.n6327 585
R5748 gnd.n6330 gnd.n6329 585
R5749 gnd.n959 gnd.n958 585
R5750 gnd.n6335 gnd.n6334 585
R5751 gnd.n6336 gnd.n6335 585
R5752 gnd.n6671 gnd.n632 585
R5753 gnd.n639 gnd.n632 585
R5754 gnd.n6670 gnd.n6669 585
R5755 gnd.n6669 gnd.n6668 585
R5756 gnd.n637 gnd.n636 585
R5757 gnd.n648 gnd.n637 585
R5758 gnd.n6657 gnd.n6656 585
R5759 gnd.n6658 gnd.n6657 585
R5760 gnd.n650 gnd.n649 585
R5761 gnd.n649 gnd.n646 585
R5762 gnd.n6651 gnd.n6650 585
R5763 gnd.n6650 gnd.n6649 585
R5764 gnd.n653 gnd.n652 585
R5765 gnd.n654 gnd.n653 585
R5766 gnd.n6640 gnd.n6639 585
R5767 gnd.n6641 gnd.n6640 585
R5768 gnd.n664 gnd.n663 585
R5769 gnd.n663 gnd.n661 585
R5770 gnd.n6635 gnd.n6634 585
R5771 gnd.n6634 gnd.n6633 585
R5772 gnd.n667 gnd.n666 585
R5773 gnd.n668 gnd.n667 585
R5774 gnd.n6624 gnd.n6623 585
R5775 gnd.n6625 gnd.n6624 585
R5776 gnd.n677 gnd.n676 585
R5777 gnd.n5937 gnd.n676 585
R5778 gnd.n6619 gnd.n6618 585
R5779 gnd.n6618 gnd.n6617 585
R5780 gnd.n680 gnd.n679 585
R5781 gnd.n5935 gnd.n680 585
R5782 gnd.n6608 gnd.n6607 585
R5783 gnd.n6609 gnd.n6608 585
R5784 gnd.n692 gnd.n691 585
R5785 gnd.n5795 gnd.n691 585
R5786 gnd.n6603 gnd.n6602 585
R5787 gnd.n6602 gnd.n6601 585
R5788 gnd.n695 gnd.n694 585
R5789 gnd.n5243 gnd.n695 585
R5790 gnd.n6592 gnd.n6591 585
R5791 gnd.n6593 gnd.n6592 585
R5792 gnd.n707 gnd.n706 585
R5793 gnd.n5780 gnd.n706 585
R5794 gnd.n6587 gnd.n6586 585
R5795 gnd.n6586 gnd.n6585 585
R5796 gnd.n710 gnd.n709 585
R5797 gnd.n5251 gnd.n710 585
R5798 gnd.n6576 gnd.n6575 585
R5799 gnd.n6577 gnd.n6576 585
R5800 gnd.n722 gnd.n721 585
R5801 gnd.n5763 gnd.n721 585
R5802 gnd.n6571 gnd.n6570 585
R5803 gnd.n6570 gnd.n6569 585
R5804 gnd.n725 gnd.n724 585
R5805 gnd.n5261 gnd.n725 585
R5806 gnd.n6560 gnd.n6559 585
R5807 gnd.n6561 gnd.n6560 585
R5808 gnd.n736 gnd.n735 585
R5809 gnd.n5265 gnd.n735 585
R5810 gnd.n6555 gnd.n6554 585
R5811 gnd.n6554 gnd.n6553 585
R5812 gnd.n739 gnd.n738 585
R5813 gnd.n5271 gnd.n739 585
R5814 gnd.n6544 gnd.n6543 585
R5815 gnd.n6545 gnd.n6544 585
R5816 gnd.n751 gnd.n750 585
R5817 gnd.n5276 gnd.n750 585
R5818 gnd.n6539 gnd.n6538 585
R5819 gnd.n6538 gnd.n6537 585
R5820 gnd.n754 gnd.n753 585
R5821 gnd.n5281 gnd.n754 585
R5822 gnd.n6528 gnd.n6527 585
R5823 gnd.n6529 gnd.n6528 585
R5824 gnd.n767 gnd.n766 585
R5825 gnd.n5286 gnd.n766 585
R5826 gnd.n6523 gnd.n6522 585
R5827 gnd.n6522 gnd.n6521 585
R5828 gnd.n770 gnd.n769 585
R5829 gnd.n5291 gnd.n770 585
R5830 gnd.n6512 gnd.n6511 585
R5831 gnd.n6513 gnd.n6512 585
R5832 gnd.n782 gnd.n781 585
R5833 gnd.n5297 gnd.n781 585
R5834 gnd.n6507 gnd.n6506 585
R5835 gnd.n6506 gnd.n6505 585
R5836 gnd.n785 gnd.n784 585
R5837 gnd.n5302 gnd.n785 585
R5838 gnd.n6496 gnd.n6495 585
R5839 gnd.n6497 gnd.n6496 585
R5840 gnd.n797 gnd.n796 585
R5841 gnd.n5307 gnd.n796 585
R5842 gnd.n6491 gnd.n6490 585
R5843 gnd.n6490 gnd.n6489 585
R5844 gnd.n800 gnd.n799 585
R5845 gnd.n5313 gnd.n800 585
R5846 gnd.n6480 gnd.n6479 585
R5847 gnd.n6481 gnd.n6480 585
R5848 gnd.n813 gnd.n812 585
R5849 gnd.n5656 gnd.n812 585
R5850 gnd.n6475 gnd.n6474 585
R5851 gnd.n6474 gnd.n6473 585
R5852 gnd.n816 gnd.n815 585
R5853 gnd.n5322 gnd.n816 585
R5854 gnd.n6464 gnd.n6463 585
R5855 gnd.n6465 gnd.n6464 585
R5856 gnd.n829 gnd.n828 585
R5857 gnd.n5637 gnd.n828 585
R5858 gnd.n6459 gnd.n6458 585
R5859 gnd.n6458 gnd.n6457 585
R5860 gnd.n832 gnd.n831 585
R5861 gnd.n5331 gnd.n832 585
R5862 gnd.n6448 gnd.n6447 585
R5863 gnd.n6449 gnd.n6448 585
R5864 gnd.n843 gnd.n842 585
R5865 gnd.n5619 gnd.n842 585
R5866 gnd.n6443 gnd.n6442 585
R5867 gnd.n6442 gnd.n6441 585
R5868 gnd.n846 gnd.n845 585
R5869 gnd.n5341 gnd.n846 585
R5870 gnd.n6432 gnd.n6431 585
R5871 gnd.n6433 gnd.n6432 585
R5872 gnd.n858 gnd.n857 585
R5873 gnd.n5345 gnd.n857 585
R5874 gnd.n6427 gnd.n6426 585
R5875 gnd.n6426 gnd.n6425 585
R5876 gnd.n861 gnd.n860 585
R5877 gnd.n5351 gnd.n861 585
R5878 gnd.n6416 gnd.n6415 585
R5879 gnd.n6417 gnd.n6416 585
R5880 gnd.n873 gnd.n872 585
R5881 gnd.n5356 gnd.n872 585
R5882 gnd.n6411 gnd.n6410 585
R5883 gnd.n6410 gnd.n6409 585
R5884 gnd.n876 gnd.n875 585
R5885 gnd.n5361 gnd.n876 585
R5886 gnd.n6400 gnd.n6399 585
R5887 gnd.n6401 gnd.n6400 585
R5888 gnd.n889 gnd.n888 585
R5889 gnd.n5366 gnd.n888 585
R5890 gnd.n6395 gnd.n6394 585
R5891 gnd.n6394 gnd.n6393 585
R5892 gnd.n892 gnd.n891 585
R5893 gnd.n901 gnd.n892 585
R5894 gnd.n6384 gnd.n6383 585
R5895 gnd.n6385 gnd.n6384 585
R5896 gnd.n903 gnd.n902 585
R5897 gnd.n909 gnd.n902 585
R5898 gnd.n6379 gnd.n6378 585
R5899 gnd.n6378 gnd.n6377 585
R5900 gnd.n906 gnd.n905 585
R5901 gnd.n907 gnd.n906 585
R5902 gnd.n6368 gnd.n6367 585
R5903 gnd.n6369 gnd.n6368 585
R5904 gnd.n917 gnd.n916 585
R5905 gnd.n923 gnd.n916 585
R5906 gnd.n6363 gnd.n6362 585
R5907 gnd.n6362 gnd.n6361 585
R5908 gnd.n920 gnd.n919 585
R5909 gnd.n921 gnd.n920 585
R5910 gnd.n6352 gnd.n6351 585
R5911 gnd.n6353 gnd.n6352 585
R5912 gnd.n932 gnd.n931 585
R5913 gnd.n931 gnd.n929 585
R5914 gnd.n6347 gnd.n6346 585
R5915 gnd.n6346 gnd.n6345 585
R5916 gnd.n935 gnd.n934 585
R5917 gnd.n936 gnd.n935 585
R5918 gnd.n6675 gnd.n6674 585
R5919 gnd.n6677 gnd.n6675 585
R5920 gnd.n633 gnd.n631 585
R5921 gnd.n6029 gnd.n6028 585
R5922 gnd.n6030 gnd.n6027 585
R5923 gnd.n6022 gnd.n6021 585
R5924 gnd.n6034 gnd.n6020 585
R5925 gnd.n6035 gnd.n6019 585
R5926 gnd.n6036 gnd.n6018 585
R5927 gnd.n6016 gnd.n6015 585
R5928 gnd.n6040 gnd.n6014 585
R5929 gnd.n6041 gnd.n6013 585
R5930 gnd.n6042 gnd.n6012 585
R5931 gnd.n6009 gnd.n6008 585
R5932 gnd.n6052 gnd.n6007 585
R5933 gnd.n6053 gnd.n6006 585
R5934 gnd.n6005 gnd.n5997 585
R5935 gnd.n6060 gnd.n5996 585
R5936 gnd.n6061 gnd.n5995 585
R5937 gnd.n5989 gnd.n5988 585
R5938 gnd.n6068 gnd.n5987 585
R5939 gnd.n6069 gnd.n5986 585
R5940 gnd.n5985 gnd.n5977 585
R5941 gnd.n6076 gnd.n5976 585
R5942 gnd.n6077 gnd.n5975 585
R5943 gnd.n5969 gnd.n5968 585
R5944 gnd.n6084 gnd.n5967 585
R5945 gnd.n6085 gnd.n5966 585
R5946 gnd.n5965 gnd.n5951 585
R5947 gnd.n6093 gnd.n6092 585
R5948 gnd.n5928 gnd.n5164 511.721
R5949 gnd.n5811 gnd.n5810 511.721
R5950 gnd.n5560 gnd.n5368 511.721
R5951 gnd.n5432 gnd.n5365 511.721
R5952 gnd.n2554 gnd.n2553 414.56
R5953 gnd.n5385 gnd.t121 389.64
R5954 gnd.n5212 gnd.t67 389.64
R5955 gnd.n5393 gnd.t34 389.64
R5956 gnd.n5206 gnd.t124 389.64
R5957 gnd.n961 gnd.t111 371.625
R5958 gnd.n118 gnd.t52 371.625
R5959 gnd.n6047 gnd.t85 371.625
R5960 gnd.n976 gnd.t101 371.625
R5961 gnd.n537 gnd.t78 371.625
R5962 gnd.n559 gnd.t56 371.625
R5963 gnd.n197 gnd.t130 371.625
R5964 gnd.n7396 gnd.t139 371.625
R5965 gnd.n4312 gnd.t75 371.625
R5966 gnd.n4344 gnd.t42 371.625
R5967 gnd.n4173 gnd.t108 371.625
R5968 gnd.n1053 gnd.t71 371.625
R5969 gnd.n1016 gnd.t98 371.625
R5970 gnd.n6024 gnd.t88 371.625
R5971 gnd.n3250 gnd.t38 323.425
R5972 gnd.n1439 gnd.t81 323.425
R5973 gnd.n4037 gnd.n4011 289.615
R5974 gnd.n4005 gnd.n3979 289.615
R5975 gnd.n3973 gnd.n3947 289.615
R5976 gnd.n3942 gnd.n3916 289.615
R5977 gnd.n3910 gnd.n3884 289.615
R5978 gnd.n3878 gnd.n3852 289.615
R5979 gnd.n3846 gnd.n3820 289.615
R5980 gnd.n3815 gnd.n3789 289.615
R5981 gnd.n3324 gnd.t104 279.217
R5982 gnd.n1465 gnd.t60 279.217
R5983 gnd.n5415 gnd.t51 260.649
R5984 gnd.n5177 gnd.t94 260.649
R5985 gnd.n5433 gnd.n893 256.663
R5986 gnd.n5436 gnd.n893 256.663
R5987 gnd.n5442 gnd.n893 256.663
R5988 gnd.n5444 gnd.n893 256.663
R5989 gnd.n5450 gnd.n893 256.663
R5990 gnd.n5452 gnd.n893 256.663
R5991 gnd.n5458 gnd.n893 256.663
R5992 gnd.n5460 gnd.n893 256.663
R5993 gnd.n5466 gnd.n893 256.663
R5994 gnd.n5468 gnd.n893 256.663
R5995 gnd.n5474 gnd.n893 256.663
R5996 gnd.n5476 gnd.n893 256.663
R5997 gnd.n5482 gnd.n893 256.663
R5998 gnd.n5484 gnd.n893 256.663
R5999 gnd.n5491 gnd.n893 256.663
R6000 gnd.n5494 gnd.n893 256.663
R6001 gnd.n5496 gnd.n5495 256.663
R6002 gnd.n5390 gnd.n893 256.663
R6003 gnd.n5499 gnd.n893 256.663
R6004 gnd.n5501 gnd.n893 256.663
R6005 gnd.n5508 gnd.n893 256.663
R6006 gnd.n5510 gnd.n893 256.663
R6007 gnd.n5516 gnd.n893 256.663
R6008 gnd.n5518 gnd.n893 256.663
R6009 gnd.n5524 gnd.n893 256.663
R6010 gnd.n5526 gnd.n893 256.663
R6011 gnd.n5532 gnd.n893 256.663
R6012 gnd.n5534 gnd.n893 256.663
R6013 gnd.n5540 gnd.n893 256.663
R6014 gnd.n5542 gnd.n893 256.663
R6015 gnd.n5548 gnd.n893 256.663
R6016 gnd.n5550 gnd.n893 256.663
R6017 gnd.n5556 gnd.n893 256.663
R6018 gnd.n5559 gnd.n893 256.663
R6019 gnd.n5809 gnd.n683 256.663
R6020 gnd.n5816 gnd.n683 256.663
R6021 gnd.n5233 gnd.n683 256.663
R6022 gnd.n5823 gnd.n683 256.663
R6023 gnd.n5230 gnd.n683 256.663
R6024 gnd.n5830 gnd.n683 256.663
R6025 gnd.n5227 gnd.n683 256.663
R6026 gnd.n5837 gnd.n683 256.663
R6027 gnd.n5224 gnd.n683 256.663
R6028 gnd.n5844 gnd.n683 256.663
R6029 gnd.n5221 gnd.n683 256.663
R6030 gnd.n5851 gnd.n683 256.663
R6031 gnd.n5218 gnd.n683 256.663
R6032 gnd.n5858 gnd.n683 256.663
R6033 gnd.n5215 gnd.n683 256.663
R6034 gnd.n5866 gnd.n683 256.663
R6035 gnd.n5869 gnd.n534 256.663
R6036 gnd.n5870 gnd.n683 256.663
R6037 gnd.n5874 gnd.n683 256.663
R6038 gnd.n5209 gnd.n683 256.663
R6039 gnd.n5882 gnd.n683 256.663
R6040 gnd.n5204 gnd.n683 256.663
R6041 gnd.n5889 gnd.n683 256.663
R6042 gnd.n5201 gnd.n683 256.663
R6043 gnd.n5896 gnd.n683 256.663
R6044 gnd.n5198 gnd.n683 256.663
R6045 gnd.n5903 gnd.n683 256.663
R6046 gnd.n5195 gnd.n683 256.663
R6047 gnd.n5910 gnd.n683 256.663
R6048 gnd.n5192 gnd.n683 256.663
R6049 gnd.n5917 gnd.n683 256.663
R6050 gnd.n5189 gnd.n683 256.663
R6051 gnd.n5924 gnd.n683 256.663
R6052 gnd.n5927 gnd.n683 256.663
R6053 gnd.n4193 gnd.n4168 242.672
R6054 gnd.n4195 gnd.n4168 242.672
R6055 gnd.n4203 gnd.n4168 242.672
R6056 gnd.n4205 gnd.n4168 242.672
R6057 gnd.n4213 gnd.n4168 242.672
R6058 gnd.n4215 gnd.n4168 242.672
R6059 gnd.n4223 gnd.n4168 242.672
R6060 gnd.n4225 gnd.n4168 242.672
R6061 gnd.n4233 gnd.n4168 242.672
R6062 gnd.n992 gnd.n979 242.672
R6063 gnd.n5050 gnd.n992 242.672
R6064 gnd.n5047 gnd.n992 242.672
R6065 gnd.n5036 gnd.n992 242.672
R6066 gnd.n5027 gnd.n992 242.672
R6067 gnd.n5024 gnd.n992 242.672
R6068 gnd.n5013 gnd.n992 242.672
R6069 gnd.n5004 gnd.n992 242.672
R6070 gnd.n5001 gnd.n992 242.672
R6071 gnd.n6906 gnd.n508 242.672
R6072 gnd.n6906 gnd.n509 242.672
R6073 gnd.n6906 gnd.n510 242.672
R6074 gnd.n6906 gnd.n511 242.672
R6075 gnd.n6906 gnd.n512 242.672
R6076 gnd.n6906 gnd.n513 242.672
R6077 gnd.n6906 gnd.n514 242.672
R6078 gnd.n6906 gnd.n515 242.672
R6079 gnd.n6906 gnd.n516 242.672
R6080 gnd.n124 gnd.n121 242.672
R6081 gnd.n7307 gnd.n124 242.672
R6082 gnd.n7303 gnd.n124 242.672
R6083 gnd.n7300 gnd.n124 242.672
R6084 gnd.n7295 gnd.n124 242.672
R6085 gnd.n7292 gnd.n124 242.672
R6086 gnd.n7287 gnd.n124 242.672
R6087 gnd.n7284 gnd.n124 242.672
R6088 gnd.n7279 gnd.n124 242.672
R6089 gnd.n3378 gnd.n3377 242.672
R6090 gnd.n3378 gnd.n3288 242.672
R6091 gnd.n3378 gnd.n3289 242.672
R6092 gnd.n3378 gnd.n3290 242.672
R6093 gnd.n3378 gnd.n3291 242.672
R6094 gnd.n3378 gnd.n3292 242.672
R6095 gnd.n3378 gnd.n3293 242.672
R6096 gnd.n3378 gnd.n3294 242.672
R6097 gnd.n3378 gnd.n3295 242.672
R6098 gnd.n3378 gnd.n3296 242.672
R6099 gnd.n3378 gnd.n3297 242.672
R6100 gnd.n3378 gnd.n3298 242.672
R6101 gnd.n3379 gnd.n3378 242.672
R6102 gnd.n4167 gnd.n1414 242.672
R6103 gnd.n4167 gnd.n1413 242.672
R6104 gnd.n4167 gnd.n1412 242.672
R6105 gnd.n4167 gnd.n1411 242.672
R6106 gnd.n4167 gnd.n1410 242.672
R6107 gnd.n4167 gnd.n1409 242.672
R6108 gnd.n4167 gnd.n1408 242.672
R6109 gnd.n4167 gnd.n1407 242.672
R6110 gnd.n4167 gnd.n1406 242.672
R6111 gnd.n4167 gnd.n1405 242.672
R6112 gnd.n4167 gnd.n1404 242.672
R6113 gnd.n4167 gnd.n1403 242.672
R6114 gnd.n4167 gnd.n1402 242.672
R6115 gnd.n3462 gnd.n3461 242.672
R6116 gnd.n3461 gnd.n3200 242.672
R6117 gnd.n3461 gnd.n3201 242.672
R6118 gnd.n3461 gnd.n3202 242.672
R6119 gnd.n3461 gnd.n3203 242.672
R6120 gnd.n3461 gnd.n3204 242.672
R6121 gnd.n3461 gnd.n3205 242.672
R6122 gnd.n3461 gnd.n3206 242.672
R6123 gnd.n4167 gnd.n1415 242.672
R6124 gnd.n4167 gnd.n1416 242.672
R6125 gnd.n4167 gnd.n1417 242.672
R6126 gnd.n4167 gnd.n1418 242.672
R6127 gnd.n4167 gnd.n1419 242.672
R6128 gnd.n4167 gnd.n1420 242.672
R6129 gnd.n4167 gnd.n1421 242.672
R6130 gnd.n4167 gnd.n1422 242.672
R6131 gnd.n4474 gnd.n4168 242.672
R6132 gnd.n4288 gnd.n4168 242.672
R6133 gnd.n4467 gnd.n4168 242.672
R6134 gnd.n4461 gnd.n4168 242.672
R6135 gnd.n4459 gnd.n4168 242.672
R6136 gnd.n4453 gnd.n4168 242.672
R6137 gnd.n4451 gnd.n4168 242.672
R6138 gnd.n4445 gnd.n4168 242.672
R6139 gnd.n4443 gnd.n4168 242.672
R6140 gnd.n4437 gnd.n4168 242.672
R6141 gnd.n4435 gnd.n4168 242.672
R6142 gnd.n4429 gnd.n4168 242.672
R6143 gnd.n4427 gnd.n4168 242.672
R6144 gnd.n4421 gnd.n4168 242.672
R6145 gnd.n4419 gnd.n4168 242.672
R6146 gnd.n4413 gnd.n4168 242.672
R6147 gnd.n4411 gnd.n4168 242.672
R6148 gnd.n4342 gnd.n4168 242.672
R6149 gnd.n4401 gnd.n4168 242.672
R6150 gnd.n6233 gnd.n992 242.672
R6151 gnd.n1056 gnd.n992 242.672
R6152 gnd.n6240 gnd.n992 242.672
R6153 gnd.n1047 gnd.n992 242.672
R6154 gnd.n6247 gnd.n992 242.672
R6155 gnd.n1040 gnd.n992 242.672
R6156 gnd.n6254 gnd.n992 242.672
R6157 gnd.n1033 gnd.n992 242.672
R6158 gnd.n6261 gnd.n992 242.672
R6159 gnd.n1026 gnd.n992 242.672
R6160 gnd.n6268 gnd.n992 242.672
R6161 gnd.n6269 gnd.n1018 242.672
R6162 gnd.n6270 gnd.n992 242.672
R6163 gnd.n1015 gnd.n992 242.672
R6164 gnd.n6277 gnd.n992 242.672
R6165 gnd.n1008 gnd.n992 242.672
R6166 gnd.n6284 gnd.n992 242.672
R6167 gnd.n1001 gnd.n992 242.672
R6168 gnd.n6291 gnd.n992 242.672
R6169 gnd.n6294 gnd.n992 242.672
R6170 gnd.n6907 gnd.n6906 242.672
R6171 gnd.n6906 gnd.n490 242.672
R6172 gnd.n6906 gnd.n491 242.672
R6173 gnd.n6906 gnd.n492 242.672
R6174 gnd.n6906 gnd.n493 242.672
R6175 gnd.n6906 gnd.n494 242.672
R6176 gnd.n6906 gnd.n495 242.672
R6177 gnd.n6906 gnd.n496 242.672
R6178 gnd.n6878 gnd.n535 242.672
R6179 gnd.n6906 gnd.n497 242.672
R6180 gnd.n6906 gnd.n498 242.672
R6181 gnd.n6906 gnd.n499 242.672
R6182 gnd.n6906 gnd.n500 242.672
R6183 gnd.n6906 gnd.n501 242.672
R6184 gnd.n6906 gnd.n502 242.672
R6185 gnd.n6906 gnd.n503 242.672
R6186 gnd.n6906 gnd.n504 242.672
R6187 gnd.n6906 gnd.n505 242.672
R6188 gnd.n6906 gnd.n506 242.672
R6189 gnd.n6906 gnd.n507 242.672
R6190 gnd.n194 gnd.n124 242.672
R6191 gnd.n7364 gnd.n124 242.672
R6192 gnd.n190 gnd.n124 242.672
R6193 gnd.n7371 gnd.n124 242.672
R6194 gnd.n183 gnd.n124 242.672
R6195 gnd.n7378 gnd.n124 242.672
R6196 gnd.n176 gnd.n124 242.672
R6197 gnd.n7385 gnd.n124 242.672
R6198 gnd.n169 gnd.n124 242.672
R6199 gnd.n7392 gnd.n124 242.672
R6200 gnd.n162 gnd.n124 242.672
R6201 gnd.n7402 gnd.n124 242.672
R6202 gnd.n155 gnd.n124 242.672
R6203 gnd.n7409 gnd.n124 242.672
R6204 gnd.n148 gnd.n124 242.672
R6205 gnd.n7416 gnd.n124 242.672
R6206 gnd.n141 gnd.n124 242.672
R6207 gnd.n7423 gnd.n124 242.672
R6208 gnd.n134 gnd.n124 242.672
R6209 gnd.n6336 gnd.n944 242.672
R6210 gnd.n6336 gnd.n945 242.672
R6211 gnd.n6336 gnd.n946 242.672
R6212 gnd.n6336 gnd.n947 242.672
R6213 gnd.n6336 gnd.n948 242.672
R6214 gnd.n6336 gnd.n949 242.672
R6215 gnd.n6336 gnd.n950 242.672
R6216 gnd.n6336 gnd.n951 242.672
R6217 gnd.n6336 gnd.n952 242.672
R6218 gnd.n6336 gnd.n953 242.672
R6219 gnd.n6336 gnd.n954 242.672
R6220 gnd.n6336 gnd.n955 242.672
R6221 gnd.n6336 gnd.n956 242.672
R6222 gnd.n6336 gnd.n957 242.672
R6223 gnd.n6677 gnd.n630 242.672
R6224 gnd.n6677 gnd.n629 242.672
R6225 gnd.n6677 gnd.n628 242.672
R6226 gnd.n6677 gnd.n627 242.672
R6227 gnd.n6677 gnd.n626 242.672
R6228 gnd.n6677 gnd.n625 242.672
R6229 gnd.n6677 gnd.n624 242.672
R6230 gnd.n6677 gnd.n623 242.672
R6231 gnd.n6677 gnd.n622 242.672
R6232 gnd.n6677 gnd.n621 242.672
R6233 gnd.n6677 gnd.n620 242.672
R6234 gnd.n6677 gnd.n619 242.672
R6235 gnd.n6677 gnd.n618 242.672
R6236 gnd.n6677 gnd.n617 242.672
R6237 gnd.n131 gnd.n127 240.244
R6238 gnd.n7425 gnd.n7424 240.244
R6239 gnd.n7422 gnd.n135 240.244
R6240 gnd.n7418 gnd.n7417 240.244
R6241 gnd.n7415 gnd.n142 240.244
R6242 gnd.n7411 gnd.n7410 240.244
R6243 gnd.n7408 gnd.n149 240.244
R6244 gnd.n7404 gnd.n7403 240.244
R6245 gnd.n7401 gnd.n156 240.244
R6246 gnd.n7394 gnd.n7393 240.244
R6247 gnd.n7391 gnd.n163 240.244
R6248 gnd.n7387 gnd.n7386 240.244
R6249 gnd.n7384 gnd.n170 240.244
R6250 gnd.n7380 gnd.n7379 240.244
R6251 gnd.n7377 gnd.n177 240.244
R6252 gnd.n7373 gnd.n7372 240.244
R6253 gnd.n7370 gnd.n184 240.244
R6254 gnd.n7366 gnd.n7365 240.244
R6255 gnd.n7363 gnd.n191 240.244
R6256 gnd.n6835 gnd.n481 240.244
R6257 gnd.n6707 gnd.n481 240.244
R6258 gnd.n6707 gnd.n472 240.244
R6259 gnd.n6711 gnd.n472 240.244
R6260 gnd.n6711 gnd.n463 240.244
R6261 gnd.n6724 gnd.n463 240.244
R6262 gnd.n6724 gnd.n454 240.244
R6263 gnd.n6720 gnd.n454 240.244
R6264 gnd.n6720 gnd.n447 240.244
R6265 gnd.n6747 gnd.n447 240.244
R6266 gnd.n6747 gnd.n438 240.244
R6267 gnd.n6751 gnd.n438 240.244
R6268 gnd.n6751 gnd.n429 240.244
R6269 gnd.n6763 gnd.n429 240.244
R6270 gnd.n6763 gnd.n420 240.244
R6271 gnd.n6759 gnd.n420 240.244
R6272 gnd.n6759 gnd.n413 240.244
R6273 gnd.n6778 gnd.n413 240.244
R6274 gnd.n6778 gnd.n402 240.244
R6275 gnd.n6797 gnd.n402 240.244
R6276 gnd.n6797 gnd.n394 240.244
R6277 gnd.n394 gnd.n387 240.244
R6278 gnd.n387 gnd.n370 240.244
R6279 gnd.n6791 gnd.n370 240.244
R6280 gnd.n6791 gnd.n358 240.244
R6281 gnd.n7051 gnd.n358 240.244
R6282 gnd.n7052 gnd.n7051 240.244
R6283 gnd.n7052 gnd.n350 240.244
R6284 gnd.n350 gnd.n309 240.244
R6285 gnd.n7061 gnd.n309 240.244
R6286 gnd.n7061 gnd.n339 240.244
R6287 gnd.n339 gnd.n335 240.244
R6288 gnd.n7089 gnd.n335 240.244
R6289 gnd.n7089 gnd.n331 240.244
R6290 gnd.n7160 gnd.n331 240.244
R6291 gnd.n7160 gnd.n324 240.244
R6292 gnd.n7156 gnd.n324 240.244
R6293 gnd.n7156 gnd.n296 240.244
R6294 gnd.n7153 gnd.n296 240.244
R6295 gnd.n7153 gnd.n287 240.244
R6296 gnd.n7150 gnd.n287 240.244
R6297 gnd.n7150 gnd.n279 240.244
R6298 gnd.n7147 gnd.n279 240.244
R6299 gnd.n7147 gnd.n272 240.244
R6300 gnd.n7144 gnd.n272 240.244
R6301 gnd.n7144 gnd.n266 240.244
R6302 gnd.n7141 gnd.n266 240.244
R6303 gnd.n7141 gnd.n257 240.244
R6304 gnd.n7138 gnd.n257 240.244
R6305 gnd.n7138 gnd.n249 240.244
R6306 gnd.n7135 gnd.n249 240.244
R6307 gnd.n7135 gnd.n242 240.244
R6308 gnd.n7132 gnd.n242 240.244
R6309 gnd.n7132 gnd.n235 240.244
R6310 gnd.n7129 gnd.n235 240.244
R6311 gnd.n7129 gnd.n226 240.244
R6312 gnd.n7126 gnd.n226 240.244
R6313 gnd.n7126 gnd.n219 240.244
R6314 gnd.n7123 gnd.n219 240.244
R6315 gnd.n7123 gnd.n210 240.244
R6316 gnd.n210 gnd.n201 240.244
R6317 gnd.n7354 gnd.n201 240.244
R6318 gnd.n7355 gnd.n7354 240.244
R6319 gnd.n7355 gnd.n123 240.244
R6320 gnd.n6905 gnd.n488 240.244
R6321 gnd.n6905 gnd.n519 240.244
R6322 gnd.n6901 gnd.n6900 240.244
R6323 gnd.n6897 gnd.n6896 240.244
R6324 gnd.n6893 gnd.n6892 240.244
R6325 gnd.n6889 gnd.n6888 240.244
R6326 gnd.n6885 gnd.n6884 240.244
R6327 gnd.n6881 gnd.n6880 240.244
R6328 gnd.n6876 gnd.n6875 240.244
R6329 gnd.n6872 gnd.n6871 240.244
R6330 gnd.n6868 gnd.n6867 240.244
R6331 gnd.n6864 gnd.n6863 240.244
R6332 gnd.n6860 gnd.n6859 240.244
R6333 gnd.n6856 gnd.n6855 240.244
R6334 gnd.n6852 gnd.n6851 240.244
R6335 gnd.n6848 gnd.n6847 240.244
R6336 gnd.n6844 gnd.n6843 240.244
R6337 gnd.n558 gnd.n557 240.244
R6338 gnd.n6914 gnd.n484 240.244
R6339 gnd.n6914 gnd.n470 240.244
R6340 gnd.n6924 gnd.n470 240.244
R6341 gnd.n6924 gnd.n466 240.244
R6342 gnd.n6930 gnd.n466 240.244
R6343 gnd.n6930 gnd.n453 240.244
R6344 gnd.n6940 gnd.n453 240.244
R6345 gnd.n6940 gnd.n449 240.244
R6346 gnd.n6946 gnd.n449 240.244
R6347 gnd.n6946 gnd.n436 240.244
R6348 gnd.n6956 gnd.n436 240.244
R6349 gnd.n6956 gnd.n432 240.244
R6350 gnd.n6962 gnd.n432 240.244
R6351 gnd.n6962 gnd.n419 240.244
R6352 gnd.n6972 gnd.n419 240.244
R6353 gnd.n6972 gnd.n415 240.244
R6354 gnd.n6978 gnd.n415 240.244
R6355 gnd.n6978 gnd.n400 240.244
R6356 gnd.n6991 gnd.n400 240.244
R6357 gnd.n6991 gnd.n396 240.244
R6358 gnd.n6997 gnd.n396 240.244
R6359 gnd.n6997 gnd.n368 240.244
R6360 gnd.n7042 gnd.n368 240.244
R6361 gnd.n7042 gnd.n369 240.244
R6362 gnd.n369 gnd.n363 240.244
R6363 gnd.n7049 gnd.n363 240.244
R6364 gnd.n7049 gnd.n364 240.244
R6365 gnd.n364 gnd.n306 240.244
R6366 gnd.n7181 gnd.n306 240.244
R6367 gnd.n7181 gnd.n307 240.244
R6368 gnd.n7083 gnd.n307 240.244
R6369 gnd.n7084 gnd.n7083 240.244
R6370 gnd.n7087 gnd.n7084 240.244
R6371 gnd.n7087 gnd.n326 240.244
R6372 gnd.n7162 gnd.n326 240.244
R6373 gnd.n7164 gnd.n7162 240.244
R6374 gnd.n7164 gnd.n297 240.244
R6375 gnd.n7188 gnd.n297 240.244
R6376 gnd.n7188 gnd.n285 240.244
R6377 gnd.n7198 gnd.n285 240.244
R6378 gnd.n7198 gnd.n281 240.244
R6379 gnd.n7204 gnd.n281 240.244
R6380 gnd.n7204 gnd.n271 240.244
R6381 gnd.n7214 gnd.n271 240.244
R6382 gnd.n7214 gnd.n267 240.244
R6383 gnd.n7220 gnd.n267 240.244
R6384 gnd.n7220 gnd.n255 240.244
R6385 gnd.n7230 gnd.n255 240.244
R6386 gnd.n7230 gnd.n251 240.244
R6387 gnd.n7236 gnd.n251 240.244
R6388 gnd.n7236 gnd.n241 240.244
R6389 gnd.n7246 gnd.n241 240.244
R6390 gnd.n7246 gnd.n237 240.244
R6391 gnd.n7252 gnd.n237 240.244
R6392 gnd.n7252 gnd.n224 240.244
R6393 gnd.n7262 gnd.n224 240.244
R6394 gnd.n7262 gnd.n220 240.244
R6395 gnd.n7268 gnd.n220 240.244
R6396 gnd.n7268 gnd.n208 240.244
R6397 gnd.n7346 gnd.n208 240.244
R6398 gnd.n7346 gnd.n204 240.244
R6399 gnd.n7352 gnd.n204 240.244
R6400 gnd.n7352 gnd.n126 240.244
R6401 gnd.n7432 gnd.n126 240.244
R6402 gnd.n6295 gnd.n987 240.244
R6403 gnd.n6293 gnd.n6292 240.244
R6404 gnd.n6290 gnd.n994 240.244
R6405 gnd.n6286 gnd.n6285 240.244
R6406 gnd.n6283 gnd.n1002 240.244
R6407 gnd.n6279 gnd.n6278 240.244
R6408 gnd.n6276 gnd.n1009 240.244
R6409 gnd.n6272 gnd.n6271 240.244
R6410 gnd.n6267 gnd.n1019 240.244
R6411 gnd.n6263 gnd.n6262 240.244
R6412 gnd.n6260 gnd.n1027 240.244
R6413 gnd.n6256 gnd.n6255 240.244
R6414 gnd.n6253 gnd.n1034 240.244
R6415 gnd.n6249 gnd.n6248 240.244
R6416 gnd.n6246 gnd.n1041 240.244
R6417 gnd.n6242 gnd.n6241 240.244
R6418 gnd.n6239 gnd.n1048 240.244
R6419 gnd.n6235 gnd.n6234 240.244
R6420 gnd.n4348 gnd.n4169 240.244
R6421 gnd.n4348 gnd.n1394 240.244
R6422 gnd.n4394 gnd.n1394 240.244
R6423 gnd.n4394 gnd.n1387 240.244
R6424 gnd.n4391 gnd.n1387 240.244
R6425 gnd.n4391 gnd.n1379 240.244
R6426 gnd.n4388 gnd.n1379 240.244
R6427 gnd.n4388 gnd.n1370 240.244
R6428 gnd.n4385 gnd.n1370 240.244
R6429 gnd.n4385 gnd.n1362 240.244
R6430 gnd.n4382 gnd.n1362 240.244
R6431 gnd.n4382 gnd.n1355 240.244
R6432 gnd.n4379 gnd.n1355 240.244
R6433 gnd.n4379 gnd.n1347 240.244
R6434 gnd.n4376 gnd.n1347 240.244
R6435 gnd.n4376 gnd.n1338 240.244
R6436 gnd.n4373 gnd.n1338 240.244
R6437 gnd.n4373 gnd.n1329 240.244
R6438 gnd.n4370 gnd.n1329 240.244
R6439 gnd.n4370 gnd.n1321 240.244
R6440 gnd.n1321 gnd.n1313 240.244
R6441 gnd.n4586 gnd.n1313 240.244
R6442 gnd.n4586 gnd.n1294 240.244
R6443 gnd.n1309 gnd.n1294 240.244
R6444 gnd.n4595 gnd.n1309 240.244
R6445 gnd.n4595 gnd.n1285 240.244
R6446 gnd.n1285 gnd.n1278 240.244
R6447 gnd.n4630 gnd.n1278 240.244
R6448 gnd.n4630 gnd.n1185 240.244
R6449 gnd.n4635 gnd.n1185 240.244
R6450 gnd.n4635 gnd.n1196 240.244
R6451 gnd.n4638 gnd.n1196 240.244
R6452 gnd.n4638 gnd.n1201 240.244
R6453 gnd.n4644 gnd.n1201 240.244
R6454 gnd.n4644 gnd.n1208 240.244
R6455 gnd.n4654 gnd.n1208 240.244
R6456 gnd.n4654 gnd.n1171 240.244
R6457 gnd.n1218 gnd.n1171 240.244
R6458 gnd.n1218 gnd.n1162 240.244
R6459 gnd.n4662 gnd.n1162 240.244
R6460 gnd.n4662 gnd.n1155 240.244
R6461 gnd.n4689 gnd.n1155 240.244
R6462 gnd.n4689 gnd.n1146 240.244
R6463 gnd.n4693 gnd.n1146 240.244
R6464 gnd.n4693 gnd.n1137 240.244
R6465 gnd.n4706 gnd.n1137 240.244
R6466 gnd.n4706 gnd.n1128 240.244
R6467 gnd.n4702 gnd.n1128 240.244
R6468 gnd.n4702 gnd.n1121 240.244
R6469 gnd.n4729 gnd.n1121 240.244
R6470 gnd.n4729 gnd.n1112 240.244
R6471 gnd.n4733 gnd.n1112 240.244
R6472 gnd.n4733 gnd.n1103 240.244
R6473 gnd.n4745 gnd.n1103 240.244
R6474 gnd.n4745 gnd.n1094 240.244
R6475 gnd.n4741 gnd.n1094 240.244
R6476 gnd.n4741 gnd.n1087 240.244
R6477 gnd.n4789 gnd.n1087 240.244
R6478 gnd.n4789 gnd.n1078 240.244
R6479 gnd.n4798 gnd.n1078 240.244
R6480 gnd.n4798 gnd.n1068 240.244
R6481 gnd.n1068 gnd.n1060 240.244
R6482 gnd.n6226 gnd.n1060 240.244
R6483 gnd.n6226 gnd.n983 240.244
R6484 gnd.n4475 gnd.n4473 240.244
R6485 gnd.n4473 gnd.n4472 240.244
R6486 gnd.n4469 gnd.n4468 240.244
R6487 gnd.n4466 gnd.n4293 240.244
R6488 gnd.n4462 gnd.n4460 240.244
R6489 gnd.n4458 gnd.n4299 240.244
R6490 gnd.n4454 gnd.n4452 240.244
R6491 gnd.n4450 gnd.n4305 240.244
R6492 gnd.n4446 gnd.n4444 240.244
R6493 gnd.n4442 gnd.n4311 240.244
R6494 gnd.n4438 gnd.n4436 240.244
R6495 gnd.n4434 gnd.n4320 240.244
R6496 gnd.n4430 gnd.n4428 240.244
R6497 gnd.n4426 gnd.n4326 240.244
R6498 gnd.n4422 gnd.n4420 240.244
R6499 gnd.n4418 gnd.n4332 240.244
R6500 gnd.n4414 gnd.n4412 240.244
R6501 gnd.n4410 gnd.n4338 240.244
R6502 gnd.n4400 gnd.n4343 240.244
R6503 gnd.n4481 gnd.n1393 240.244
R6504 gnd.n4491 gnd.n1393 240.244
R6505 gnd.n4491 gnd.n1389 240.244
R6506 gnd.n4497 gnd.n1389 240.244
R6507 gnd.n4497 gnd.n1377 240.244
R6508 gnd.n4507 gnd.n1377 240.244
R6509 gnd.n4507 gnd.n1373 240.244
R6510 gnd.n4513 gnd.n1373 240.244
R6511 gnd.n4513 gnd.n1361 240.244
R6512 gnd.n4523 gnd.n1361 240.244
R6513 gnd.n4523 gnd.n1357 240.244
R6514 gnd.n4529 gnd.n1357 240.244
R6515 gnd.n4529 gnd.n1345 240.244
R6516 gnd.n4539 gnd.n1345 240.244
R6517 gnd.n4539 gnd.n1341 240.244
R6518 gnd.n4545 gnd.n1341 240.244
R6519 gnd.n4545 gnd.n1328 240.244
R6520 gnd.n4563 gnd.n1328 240.244
R6521 gnd.n4563 gnd.n1323 240.244
R6522 gnd.n4571 gnd.n1323 240.244
R6523 gnd.n4571 gnd.n1324 240.244
R6524 gnd.n1324 gnd.n1292 240.244
R6525 gnd.n4603 gnd.n1292 240.244
R6526 gnd.n4603 gnd.n1293 240.244
R6527 gnd.n1293 gnd.n1287 240.244
R6528 gnd.n4610 gnd.n1287 240.244
R6529 gnd.n4610 gnd.n1288 240.244
R6530 gnd.n1288 gnd.n1183 240.244
R6531 gnd.n4877 gnd.n1183 240.244
R6532 gnd.n4877 gnd.n1184 240.244
R6533 gnd.n4869 gnd.n1184 240.244
R6534 gnd.n4869 gnd.n4866 240.244
R6535 gnd.n4866 gnd.n4863 240.244
R6536 gnd.n4863 gnd.n1199 240.244
R6537 gnd.n4855 gnd.n1199 240.244
R6538 gnd.n4855 gnd.n1174 240.244
R6539 gnd.n4883 gnd.n1174 240.244
R6540 gnd.n4883 gnd.n1161 240.244
R6541 gnd.n4893 gnd.n1161 240.244
R6542 gnd.n4893 gnd.n1157 240.244
R6543 gnd.n4899 gnd.n1157 240.244
R6544 gnd.n4899 gnd.n1144 240.244
R6545 gnd.n4909 gnd.n1144 240.244
R6546 gnd.n4909 gnd.n1140 240.244
R6547 gnd.n4915 gnd.n1140 240.244
R6548 gnd.n4915 gnd.n1127 240.244
R6549 gnd.n4925 gnd.n1127 240.244
R6550 gnd.n4925 gnd.n1123 240.244
R6551 gnd.n4931 gnd.n1123 240.244
R6552 gnd.n4931 gnd.n1110 240.244
R6553 gnd.n4941 gnd.n1110 240.244
R6554 gnd.n4941 gnd.n1106 240.244
R6555 gnd.n4947 gnd.n1106 240.244
R6556 gnd.n4947 gnd.n1093 240.244
R6557 gnd.n4957 gnd.n1093 240.244
R6558 gnd.n4957 gnd.n1089 240.244
R6559 gnd.n4963 gnd.n1089 240.244
R6560 gnd.n4963 gnd.n1076 240.244
R6561 gnd.n4973 gnd.n1076 240.244
R6562 gnd.n4973 gnd.n1071 240.244
R6563 gnd.n4981 gnd.n1071 240.244
R6564 gnd.n4981 gnd.n1072 240.244
R6565 gnd.n1072 gnd.n986 240.244
R6566 gnd.n6301 gnd.n986 240.244
R6567 gnd.n4166 gnd.n1424 240.244
R6568 gnd.n4159 gnd.n4158 240.244
R6569 gnd.n4156 gnd.n4155 240.244
R6570 gnd.n4152 gnd.n4151 240.244
R6571 gnd.n4148 gnd.n4147 240.244
R6572 gnd.n4144 gnd.n4143 240.244
R6573 gnd.n4140 gnd.n4139 240.244
R6574 gnd.n4136 gnd.n4135 240.244
R6575 gnd.n3473 gnd.n3185 240.244
R6576 gnd.n3483 gnd.n3185 240.244
R6577 gnd.n3483 gnd.n3176 240.244
R6578 gnd.n3176 gnd.n3165 240.244
R6579 gnd.n3504 gnd.n3165 240.244
R6580 gnd.n3504 gnd.n3159 240.244
R6581 gnd.n3514 gnd.n3159 240.244
R6582 gnd.n3514 gnd.n3148 240.244
R6583 gnd.n3148 gnd.n3138 240.244
R6584 gnd.n3540 gnd.n3138 240.244
R6585 gnd.n3541 gnd.n3540 240.244
R6586 gnd.n3542 gnd.n3541 240.244
R6587 gnd.n3542 gnd.n3117 240.244
R6588 gnd.n3578 gnd.n3117 240.244
R6589 gnd.n3578 gnd.n3118 240.244
R6590 gnd.n3574 gnd.n3118 240.244
R6591 gnd.n3574 gnd.n3573 240.244
R6592 gnd.n3573 gnd.n2942 240.244
R6593 gnd.n3608 gnd.n2942 240.244
R6594 gnd.n3608 gnd.n2933 240.244
R6595 gnd.n2933 gnd.n2925 240.244
R6596 gnd.n3629 gnd.n2925 240.244
R6597 gnd.n3629 gnd.n2919 240.244
R6598 gnd.n3639 gnd.n2919 240.244
R6599 gnd.n3639 gnd.n2910 240.244
R6600 gnd.n2910 gnd.n2900 240.244
R6601 gnd.n3660 gnd.n2900 240.244
R6602 gnd.n3660 gnd.n2893 240.244
R6603 gnd.n3670 gnd.n2893 240.244
R6604 gnd.n3670 gnd.n2884 240.244
R6605 gnd.n2884 gnd.n2873 240.244
R6606 gnd.n3691 gnd.n2873 240.244
R6607 gnd.n3691 gnd.n2867 240.244
R6608 gnd.n3701 gnd.n2867 240.244
R6609 gnd.n3701 gnd.n2859 240.244
R6610 gnd.n2859 gnd.n2849 240.244
R6611 gnd.n3722 gnd.n2849 240.244
R6612 gnd.n3722 gnd.n2843 240.244
R6613 gnd.n3732 gnd.n2843 240.244
R6614 gnd.n3732 gnd.n2834 240.244
R6615 gnd.n2834 gnd.n2823 240.244
R6616 gnd.n3753 gnd.n2823 240.244
R6617 gnd.n3753 gnd.n2817 240.244
R6618 gnd.n3763 gnd.n2817 240.244
R6619 gnd.n3763 gnd.n2808 240.244
R6620 gnd.n2808 gnd.n2798 240.244
R6621 gnd.n3784 gnd.n2798 240.244
R6622 gnd.n3784 gnd.n2791 240.244
R6623 gnd.n4050 gnd.n2791 240.244
R6624 gnd.n4050 gnd.n2783 240.244
R6625 gnd.n2783 gnd.n2773 240.244
R6626 gnd.n4070 gnd.n2773 240.244
R6627 gnd.n4070 gnd.n2775 240.244
R6628 gnd.n3463 gnd.n3198 240.244
R6629 gnd.n3219 gnd.n3198 240.244
R6630 gnd.n3222 gnd.n3221 240.244
R6631 gnd.n3229 gnd.n3228 240.244
R6632 gnd.n3232 gnd.n3231 240.244
R6633 gnd.n3239 gnd.n3238 240.244
R6634 gnd.n3242 gnd.n3241 240.244
R6635 gnd.n3249 gnd.n3248 240.244
R6636 gnd.n3471 gnd.n3195 240.244
R6637 gnd.n3195 gnd.n3174 240.244
R6638 gnd.n3494 gnd.n3174 240.244
R6639 gnd.n3494 gnd.n3168 240.244
R6640 gnd.n3502 gnd.n3168 240.244
R6641 gnd.n3502 gnd.n3170 240.244
R6642 gnd.n3170 gnd.n3146 240.244
R6643 gnd.n3524 gnd.n3146 240.244
R6644 gnd.n3524 gnd.n3141 240.244
R6645 gnd.n3538 gnd.n3141 240.244
R6646 gnd.n3538 gnd.n3142 240.244
R6647 gnd.n3534 gnd.n3142 240.244
R6648 gnd.n3534 gnd.n3114 240.244
R6649 gnd.n3581 gnd.n3114 240.244
R6650 gnd.n3582 gnd.n3581 240.244
R6651 gnd.n3583 gnd.n3582 240.244
R6652 gnd.n3583 gnd.n3110 240.244
R6653 gnd.n3589 gnd.n3110 240.244
R6654 gnd.n3589 gnd.n2932 240.244
R6655 gnd.n3619 gnd.n2932 240.244
R6656 gnd.n3619 gnd.n2927 240.244
R6657 gnd.n3627 gnd.n2927 240.244
R6658 gnd.n3627 gnd.n2928 240.244
R6659 gnd.n2928 gnd.n2908 240.244
R6660 gnd.n3650 gnd.n2908 240.244
R6661 gnd.n3650 gnd.n2903 240.244
R6662 gnd.n3658 gnd.n2903 240.244
R6663 gnd.n3658 gnd.n2904 240.244
R6664 gnd.n2904 gnd.n2882 240.244
R6665 gnd.n3681 gnd.n2882 240.244
R6666 gnd.n3681 gnd.n2876 240.244
R6667 gnd.n3689 gnd.n2876 240.244
R6668 gnd.n3689 gnd.n2878 240.244
R6669 gnd.n2878 gnd.n2857 240.244
R6670 gnd.n3712 gnd.n2857 240.244
R6671 gnd.n3712 gnd.n2851 240.244
R6672 gnd.n3720 gnd.n2851 240.244
R6673 gnd.n3720 gnd.n2853 240.244
R6674 gnd.n2853 gnd.n2832 240.244
R6675 gnd.n3743 gnd.n2832 240.244
R6676 gnd.n3743 gnd.n2826 240.244
R6677 gnd.n3751 gnd.n2826 240.244
R6678 gnd.n3751 gnd.n2828 240.244
R6679 gnd.n2828 gnd.n2806 240.244
R6680 gnd.n3774 gnd.n2806 240.244
R6681 gnd.n3774 gnd.n2801 240.244
R6682 gnd.n3782 gnd.n2801 240.244
R6683 gnd.n3782 gnd.n2802 240.244
R6684 gnd.n2802 gnd.n2781 240.244
R6685 gnd.n4060 gnd.n2781 240.244
R6686 gnd.n4060 gnd.n2777 240.244
R6687 gnd.n4068 gnd.n2777 240.244
R6688 gnd.n4068 gnd.n1423 240.244
R6689 gnd.n1443 gnd.n1401 240.244
R6690 gnd.n4126 gnd.n4125 240.244
R6691 gnd.n4122 gnd.n4121 240.244
R6692 gnd.n4118 gnd.n4117 240.244
R6693 gnd.n4114 gnd.n4113 240.244
R6694 gnd.n4110 gnd.n4109 240.244
R6695 gnd.n4106 gnd.n4105 240.244
R6696 gnd.n4102 gnd.n4101 240.244
R6697 gnd.n4098 gnd.n4097 240.244
R6698 gnd.n4094 gnd.n4093 240.244
R6699 gnd.n4090 gnd.n4089 240.244
R6700 gnd.n4086 gnd.n4085 240.244
R6701 gnd.n4082 gnd.n4081 240.244
R6702 gnd.n3386 gnd.n3283 240.244
R6703 gnd.n3386 gnd.n3276 240.244
R6704 gnd.n3397 gnd.n3276 240.244
R6705 gnd.n3397 gnd.n3272 240.244
R6706 gnd.n3403 gnd.n3272 240.244
R6707 gnd.n3403 gnd.n3264 240.244
R6708 gnd.n3413 gnd.n3264 240.244
R6709 gnd.n3413 gnd.n3259 240.244
R6710 gnd.n3449 gnd.n3259 240.244
R6711 gnd.n3449 gnd.n3260 240.244
R6712 gnd.n3260 gnd.n3207 240.244
R6713 gnd.n3444 gnd.n3207 240.244
R6714 gnd.n3444 gnd.n3443 240.244
R6715 gnd.n3443 gnd.n3186 240.244
R6716 gnd.n3439 gnd.n3186 240.244
R6717 gnd.n3439 gnd.n3177 240.244
R6718 gnd.n3436 gnd.n3177 240.244
R6719 gnd.n3436 gnd.n3435 240.244
R6720 gnd.n3435 gnd.n3160 240.244
R6721 gnd.n3431 gnd.n3160 240.244
R6722 gnd.n3431 gnd.n3149 240.244
R6723 gnd.n3149 gnd.n3129 240.244
R6724 gnd.n3550 gnd.n3129 240.244
R6725 gnd.n3550 gnd.n3124 240.244
R6726 gnd.n3558 gnd.n3124 240.244
R6727 gnd.n3558 gnd.n3125 240.244
R6728 gnd.n3125 gnd.n3093 240.244
R6729 gnd.n3598 gnd.n3093 240.244
R6730 gnd.n3598 gnd.n3094 240.244
R6731 gnd.n3109 gnd.n3094 240.244
R6732 gnd.n3109 gnd.n2944 240.244
R6733 gnd.n3605 gnd.n2944 240.244
R6734 gnd.n3605 gnd.n2934 240.244
R6735 gnd.n3023 gnd.n2934 240.244
R6736 gnd.n3026 gnd.n3023 240.244
R6737 gnd.n3026 gnd.n2920 240.244
R6738 gnd.n3020 gnd.n2920 240.244
R6739 gnd.n3020 gnd.n2911 240.244
R6740 gnd.n3017 gnd.n2911 240.244
R6741 gnd.n3017 gnd.n3016 240.244
R6742 gnd.n3016 gnd.n2895 240.244
R6743 gnd.n3012 gnd.n2895 240.244
R6744 gnd.n3012 gnd.n2885 240.244
R6745 gnd.n3009 gnd.n2885 240.244
R6746 gnd.n3009 gnd.n3008 240.244
R6747 gnd.n3008 gnd.n2868 240.244
R6748 gnd.n3004 gnd.n2868 240.244
R6749 gnd.n3004 gnd.n2860 240.244
R6750 gnd.n3001 gnd.n2860 240.244
R6751 gnd.n3001 gnd.n2998 240.244
R6752 gnd.n2998 gnd.n2844 240.244
R6753 gnd.n2994 gnd.n2844 240.244
R6754 gnd.n2994 gnd.n2835 240.244
R6755 gnd.n2991 gnd.n2835 240.244
R6756 gnd.n2991 gnd.n2990 240.244
R6757 gnd.n2990 gnd.n2818 240.244
R6758 gnd.n2986 gnd.n2818 240.244
R6759 gnd.n2986 gnd.n2809 240.244
R6760 gnd.n2983 gnd.n2809 240.244
R6761 gnd.n2983 gnd.n2982 240.244
R6762 gnd.n2982 gnd.n2793 240.244
R6763 gnd.n2978 gnd.n2793 240.244
R6764 gnd.n2978 gnd.n2784 240.244
R6765 gnd.n2784 gnd.n1472 240.244
R6766 gnd.n4077 gnd.n1472 240.244
R6767 gnd.n3300 gnd.n3299 240.244
R6768 gnd.n3371 gnd.n3299 240.244
R6769 gnd.n3369 gnd.n3368 240.244
R6770 gnd.n3365 gnd.n3364 240.244
R6771 gnd.n3361 gnd.n3360 240.244
R6772 gnd.n3357 gnd.n3356 240.244
R6773 gnd.n3353 gnd.n3352 240.244
R6774 gnd.n3349 gnd.n3348 240.244
R6775 gnd.n3345 gnd.n3344 240.244
R6776 gnd.n3341 gnd.n3340 240.244
R6777 gnd.n3337 gnd.n3336 240.244
R6778 gnd.n3333 gnd.n3332 240.244
R6779 gnd.n3329 gnd.n3287 240.244
R6780 gnd.n3389 gnd.n3281 240.244
R6781 gnd.n3389 gnd.n3277 240.244
R6782 gnd.n3395 gnd.n3277 240.244
R6783 gnd.n3395 gnd.n3270 240.244
R6784 gnd.n3405 gnd.n3270 240.244
R6785 gnd.n3405 gnd.n3266 240.244
R6786 gnd.n3411 gnd.n3266 240.244
R6787 gnd.n3411 gnd.n3257 240.244
R6788 gnd.n3451 gnd.n3257 240.244
R6789 gnd.n3451 gnd.n3208 240.244
R6790 gnd.n3459 gnd.n3208 240.244
R6791 gnd.n3459 gnd.n3209 240.244
R6792 gnd.n3209 gnd.n3187 240.244
R6793 gnd.n3480 gnd.n3187 240.244
R6794 gnd.n3480 gnd.n3179 240.244
R6795 gnd.n3491 gnd.n3179 240.244
R6796 gnd.n3491 gnd.n3180 240.244
R6797 gnd.n3180 gnd.n3161 240.244
R6798 gnd.n3511 gnd.n3161 240.244
R6799 gnd.n3511 gnd.n3151 240.244
R6800 gnd.n3521 gnd.n3151 240.244
R6801 gnd.n3521 gnd.n3132 240.244
R6802 gnd.n3548 gnd.n3132 240.244
R6803 gnd.n3548 gnd.n3122 240.244
R6804 gnd.n3561 gnd.n3122 240.244
R6805 gnd.n3562 gnd.n3561 240.244
R6806 gnd.n3562 gnd.n3097 240.244
R6807 gnd.n3596 gnd.n3097 240.244
R6808 gnd.n3596 gnd.n3098 240.244
R6809 gnd.n3592 gnd.n3098 240.244
R6810 gnd.n3592 gnd.n3106 240.244
R6811 gnd.n3106 gnd.n2936 240.244
R6812 gnd.n3616 gnd.n2936 240.244
R6813 gnd.n3616 gnd.n2937 240.244
R6814 gnd.n2937 gnd.n2921 240.244
R6815 gnd.n3636 gnd.n2921 240.244
R6816 gnd.n3636 gnd.n2913 240.244
R6817 gnd.n3647 gnd.n2913 240.244
R6818 gnd.n3647 gnd.n2914 240.244
R6819 gnd.n2914 gnd.n2896 240.244
R6820 gnd.n3667 gnd.n2896 240.244
R6821 gnd.n3667 gnd.n2887 240.244
R6822 gnd.n3678 gnd.n2887 240.244
R6823 gnd.n3678 gnd.n2888 240.244
R6824 gnd.n2888 gnd.n2869 240.244
R6825 gnd.n3698 gnd.n2869 240.244
R6826 gnd.n3698 gnd.n2861 240.244
R6827 gnd.n3709 gnd.n2861 240.244
R6828 gnd.n3709 gnd.n2862 240.244
R6829 gnd.n2862 gnd.n2845 240.244
R6830 gnd.n3729 gnd.n2845 240.244
R6831 gnd.n3729 gnd.n2837 240.244
R6832 gnd.n3740 gnd.n2837 240.244
R6833 gnd.n3740 gnd.n2838 240.244
R6834 gnd.n2838 gnd.n2819 240.244
R6835 gnd.n3760 gnd.n2819 240.244
R6836 gnd.n3760 gnd.n2811 240.244
R6837 gnd.n3771 gnd.n2811 240.244
R6838 gnd.n3771 gnd.n2812 240.244
R6839 gnd.n2812 gnd.n2794 240.244
R6840 gnd.n4047 gnd.n2794 240.244
R6841 gnd.n4047 gnd.n2786 240.244
R6842 gnd.n4057 gnd.n2786 240.244
R6843 gnd.n4057 gnd.n2768 240.244
R6844 gnd.n4075 gnd.n2768 240.244
R6845 gnd.n7278 gnd.n7277 240.244
R6846 gnd.n7283 gnd.n7280 240.244
R6847 gnd.n7286 gnd.n7285 240.244
R6848 gnd.n7291 gnd.n7288 240.244
R6849 gnd.n7294 gnd.n7293 240.244
R6850 gnd.n7299 gnd.n7296 240.244
R6851 gnd.n7302 gnd.n7301 240.244
R6852 gnd.n7306 gnd.n7304 240.244
R6853 gnd.n7309 gnd.n7308 240.244
R6854 gnd.n6833 gnd.n482 240.244
R6855 gnd.n568 gnd.n482 240.244
R6856 gnd.n568 gnd.n473 240.244
R6857 gnd.n569 gnd.n473 240.244
R6858 gnd.n569 gnd.n464 240.244
R6859 gnd.n572 gnd.n464 240.244
R6860 gnd.n572 gnd.n455 240.244
R6861 gnd.n573 gnd.n455 240.244
R6862 gnd.n573 gnd.n448 240.244
R6863 gnd.n576 gnd.n448 240.244
R6864 gnd.n576 gnd.n439 240.244
R6865 gnd.n577 gnd.n439 240.244
R6866 gnd.n577 gnd.n430 240.244
R6867 gnd.n580 gnd.n430 240.244
R6868 gnd.n580 gnd.n421 240.244
R6869 gnd.n581 gnd.n421 240.244
R6870 gnd.n581 gnd.n414 240.244
R6871 gnd.n584 gnd.n414 240.244
R6872 gnd.n584 gnd.n403 240.244
R6873 gnd.n6799 gnd.n403 240.244
R6874 gnd.n6799 gnd.n385 240.244
R6875 gnd.n7020 gnd.n385 240.244
R6876 gnd.n7020 gnd.n371 240.244
R6877 gnd.n380 gnd.n371 240.244
R6878 gnd.n7028 gnd.n380 240.244
R6879 gnd.n7028 gnd.n360 240.244
R6880 gnd.n360 gnd.n351 240.244
R6881 gnd.n7070 gnd.n351 240.244
R6882 gnd.n7070 gnd.n310 240.244
R6883 gnd.n7063 gnd.n310 240.244
R6884 gnd.n7063 gnd.n341 240.244
R6885 gnd.n341 gnd.n340 240.244
R6886 gnd.n340 gnd.n78 240.244
R6887 gnd.n79 gnd.n78 240.244
R6888 gnd.n80 gnd.n79 240.244
R6889 gnd.n325 gnd.n80 240.244
R6890 gnd.n325 gnd.n83 240.244
R6891 gnd.n84 gnd.n83 240.244
R6892 gnd.n85 gnd.n84 240.244
R6893 gnd.n288 gnd.n85 240.244
R6894 gnd.n288 gnd.n88 240.244
R6895 gnd.n89 gnd.n88 240.244
R6896 gnd.n90 gnd.n89 240.244
R6897 gnd.n273 gnd.n90 240.244
R6898 gnd.n273 gnd.n93 240.244
R6899 gnd.n94 gnd.n93 240.244
R6900 gnd.n95 gnd.n94 240.244
R6901 gnd.n258 gnd.n95 240.244
R6902 gnd.n258 gnd.n98 240.244
R6903 gnd.n99 gnd.n98 240.244
R6904 gnd.n100 gnd.n99 240.244
R6905 gnd.n243 gnd.n100 240.244
R6906 gnd.n243 gnd.n103 240.244
R6907 gnd.n104 gnd.n103 240.244
R6908 gnd.n105 gnd.n104 240.244
R6909 gnd.n227 gnd.n105 240.244
R6910 gnd.n227 gnd.n108 240.244
R6911 gnd.n109 gnd.n108 240.244
R6912 gnd.n110 gnd.n109 240.244
R6913 gnd.n211 gnd.n110 240.244
R6914 gnd.n211 gnd.n113 240.244
R6915 gnd.n114 gnd.n113 240.244
R6916 gnd.n115 gnd.n114 240.244
R6917 gnd.n7434 gnd.n115 240.244
R6918 gnd.n5960 gnd.n5959 240.244
R6919 gnd.n5962 gnd.n5961 240.244
R6920 gnd.n5972 gnd.n5971 240.244
R6921 gnd.n5980 gnd.n5979 240.244
R6922 gnd.n5982 gnd.n5981 240.244
R6923 gnd.n5992 gnd.n5991 240.244
R6924 gnd.n6000 gnd.n5999 240.244
R6925 gnd.n6002 gnd.n6001 240.244
R6926 gnd.n6046 gnd.n517 240.244
R6927 gnd.n6916 gnd.n479 240.244
R6928 gnd.n6916 gnd.n475 240.244
R6929 gnd.n6922 gnd.n475 240.244
R6930 gnd.n6922 gnd.n461 240.244
R6931 gnd.n6932 gnd.n461 240.244
R6932 gnd.n6932 gnd.n457 240.244
R6933 gnd.n6938 gnd.n457 240.244
R6934 gnd.n6938 gnd.n445 240.244
R6935 gnd.n6948 gnd.n445 240.244
R6936 gnd.n6948 gnd.n441 240.244
R6937 gnd.n6954 gnd.n441 240.244
R6938 gnd.n6954 gnd.n427 240.244
R6939 gnd.n6964 gnd.n427 240.244
R6940 gnd.n6964 gnd.n423 240.244
R6941 gnd.n6970 gnd.n423 240.244
R6942 gnd.n6970 gnd.n411 240.244
R6943 gnd.n6980 gnd.n411 240.244
R6944 gnd.n6980 gnd.n405 240.244
R6945 gnd.n6989 gnd.n405 240.244
R6946 gnd.n6989 gnd.n406 240.244
R6947 gnd.n406 gnd.n395 240.244
R6948 gnd.n395 gnd.n373 240.244
R6949 gnd.n7040 gnd.n373 240.244
R6950 gnd.n7040 gnd.n374 240.244
R6951 gnd.n7030 gnd.n374 240.244
R6952 gnd.n7030 gnd.n362 240.244
R6953 gnd.n7031 gnd.n362 240.244
R6954 gnd.n7031 gnd.n312 240.244
R6955 gnd.n7179 gnd.n312 240.244
R6956 gnd.n7179 gnd.n313 240.244
R6957 gnd.n318 gnd.n313 240.244
R6958 gnd.n319 gnd.n318 240.244
R6959 gnd.n320 gnd.n319 240.244
R6960 gnd.n329 gnd.n320 240.244
R6961 gnd.n329 gnd.n323 240.244
R6962 gnd.n7166 gnd.n323 240.244
R6963 gnd.n7166 gnd.n294 240.244
R6964 gnd.n7190 gnd.n294 240.244
R6965 gnd.n7190 gnd.n290 240.244
R6966 gnd.n7196 gnd.n290 240.244
R6967 gnd.n7196 gnd.n278 240.244
R6968 gnd.n7206 gnd.n278 240.244
R6969 gnd.n7206 gnd.n274 240.244
R6970 gnd.n7212 gnd.n274 240.244
R6971 gnd.n7212 gnd.n264 240.244
R6972 gnd.n7222 gnd.n264 240.244
R6973 gnd.n7222 gnd.n260 240.244
R6974 gnd.n7228 gnd.n260 240.244
R6975 gnd.n7228 gnd.n248 240.244
R6976 gnd.n7238 gnd.n248 240.244
R6977 gnd.n7238 gnd.n244 240.244
R6978 gnd.n7244 gnd.n244 240.244
R6979 gnd.n7244 gnd.n233 240.244
R6980 gnd.n7254 gnd.n233 240.244
R6981 gnd.n7254 gnd.n229 240.244
R6982 gnd.n7260 gnd.n229 240.244
R6983 gnd.n7260 gnd.n218 240.244
R6984 gnd.n7270 gnd.n218 240.244
R6985 gnd.n7270 gnd.n212 240.244
R6986 gnd.n7344 gnd.n212 240.244
R6987 gnd.n7344 gnd.n213 240.244
R6988 gnd.n213 gnd.n203 240.244
R6989 gnd.n7275 gnd.n203 240.244
R6990 gnd.n7275 gnd.n125 240.244
R6991 gnd.n5000 gnd.n4998 240.244
R6992 gnd.n5003 gnd.n5002 240.244
R6993 gnd.n5012 gnd.n5005 240.244
R6994 gnd.n5015 gnd.n5014 240.244
R6995 gnd.n5026 gnd.n5025 240.244
R6996 gnd.n5035 gnd.n5028 240.244
R6997 gnd.n5038 gnd.n5037 240.244
R6998 gnd.n5049 gnd.n5048 240.244
R6999 gnd.n5052 gnd.n5051 240.244
R7000 gnd.n4283 gnd.n4170 240.244
R7001 gnd.n4283 gnd.n1395 240.244
R7002 gnd.n4279 gnd.n1395 240.244
R7003 gnd.n4279 gnd.n1388 240.244
R7004 gnd.n4276 gnd.n1388 240.244
R7005 gnd.n4276 gnd.n1380 240.244
R7006 gnd.n4273 gnd.n1380 240.244
R7007 gnd.n4273 gnd.n1371 240.244
R7008 gnd.n4270 gnd.n1371 240.244
R7009 gnd.n4270 gnd.n1363 240.244
R7010 gnd.n4267 gnd.n1363 240.244
R7011 gnd.n4267 gnd.n1356 240.244
R7012 gnd.n4264 gnd.n1356 240.244
R7013 gnd.n4264 gnd.n1348 240.244
R7014 gnd.n4261 gnd.n1348 240.244
R7015 gnd.n4261 gnd.n1339 240.244
R7016 gnd.n4258 gnd.n1339 240.244
R7017 gnd.n4258 gnd.n1330 240.244
R7018 gnd.n1330 gnd.n1319 240.244
R7019 gnd.n4573 gnd.n1319 240.244
R7020 gnd.n4573 gnd.n1315 240.244
R7021 gnd.n4584 gnd.n1315 240.244
R7022 gnd.n4584 gnd.n1295 240.244
R7023 gnd.n4580 gnd.n1295 240.244
R7024 gnd.n4580 gnd.n1284 240.244
R7025 gnd.n4612 gnd.n1284 240.244
R7026 gnd.n4612 gnd.n1280 240.244
R7027 gnd.n4628 gnd.n1280 240.244
R7028 gnd.n4628 gnd.n1186 240.244
R7029 gnd.n4624 gnd.n1186 240.244
R7030 gnd.n4624 gnd.n1197 240.244
R7031 gnd.n4620 gnd.n1197 240.244
R7032 gnd.n4620 gnd.n1202 240.244
R7033 gnd.n4646 gnd.n1202 240.244
R7034 gnd.n4646 gnd.n1209 240.244
R7035 gnd.n4652 gnd.n1209 240.244
R7036 gnd.n4652 gnd.n1172 240.244
R7037 gnd.n4843 gnd.n1172 240.244
R7038 gnd.n4843 gnd.n1163 240.244
R7039 gnd.n1223 gnd.n1163 240.244
R7040 gnd.n1223 gnd.n1156 240.244
R7041 gnd.n1224 gnd.n1156 240.244
R7042 gnd.n1224 gnd.n1147 240.244
R7043 gnd.n1227 gnd.n1147 240.244
R7044 gnd.n1227 gnd.n1138 240.244
R7045 gnd.n1228 gnd.n1138 240.244
R7046 gnd.n1228 gnd.n1129 240.244
R7047 gnd.n1231 gnd.n1129 240.244
R7048 gnd.n1231 gnd.n1122 240.244
R7049 gnd.n1232 gnd.n1122 240.244
R7050 gnd.n1232 gnd.n1113 240.244
R7051 gnd.n1235 gnd.n1113 240.244
R7052 gnd.n1235 gnd.n1104 240.244
R7053 gnd.n1236 gnd.n1104 240.244
R7054 gnd.n1236 gnd.n1095 240.244
R7055 gnd.n1239 gnd.n1095 240.244
R7056 gnd.n1239 gnd.n1088 240.244
R7057 gnd.n1240 gnd.n1088 240.244
R7058 gnd.n1240 gnd.n1079 240.244
R7059 gnd.n4800 gnd.n1079 240.244
R7060 gnd.n4800 gnd.n1069 240.244
R7061 gnd.n4802 gnd.n1069 240.244
R7062 gnd.n4802 gnd.n980 240.244
R7063 gnd.n6303 gnd.n980 240.244
R7064 gnd.n4196 gnd.n4194 240.244
R7065 gnd.n4202 gnd.n4188 240.244
R7066 gnd.n4206 gnd.n4204 240.244
R7067 gnd.n4212 gnd.n4184 240.244
R7068 gnd.n4216 gnd.n4214 240.244
R7069 gnd.n4222 gnd.n4180 240.244
R7070 gnd.n4226 gnd.n4224 240.244
R7071 gnd.n4232 gnd.n4176 240.244
R7072 gnd.n4235 gnd.n4234 240.244
R7073 gnd.n4483 gnd.n1396 240.244
R7074 gnd.n4489 gnd.n1396 240.244
R7075 gnd.n4489 gnd.n1385 240.244
R7076 gnd.n4499 gnd.n1385 240.244
R7077 gnd.n4499 gnd.n1381 240.244
R7078 gnd.n4505 gnd.n1381 240.244
R7079 gnd.n4505 gnd.n1368 240.244
R7080 gnd.n4515 gnd.n1368 240.244
R7081 gnd.n4515 gnd.n1364 240.244
R7082 gnd.n4521 gnd.n1364 240.244
R7083 gnd.n4521 gnd.n1353 240.244
R7084 gnd.n4531 gnd.n1353 240.244
R7085 gnd.n4531 gnd.n1349 240.244
R7086 gnd.n4537 gnd.n1349 240.244
R7087 gnd.n4537 gnd.n1336 240.244
R7088 gnd.n4547 gnd.n1336 240.244
R7089 gnd.n4547 gnd.n1331 240.244
R7090 gnd.n4561 gnd.n1331 240.244
R7091 gnd.n4561 gnd.n1332 240.244
R7092 gnd.n1332 gnd.n1322 240.244
R7093 gnd.n4556 gnd.n1322 240.244
R7094 gnd.n4556 gnd.n1297 240.244
R7095 gnd.n4601 gnd.n1297 240.244
R7096 gnd.n4601 gnd.n1298 240.244
R7097 gnd.n4597 gnd.n1298 240.244
R7098 gnd.n4597 gnd.n1286 240.244
R7099 gnd.n1306 gnd.n1286 240.244
R7100 gnd.n1306 gnd.n1188 240.244
R7101 gnd.n4875 gnd.n1188 240.244
R7102 gnd.n4875 gnd.n1189 240.244
R7103 gnd.n4871 gnd.n1189 240.244
R7104 gnd.n4871 gnd.n1195 240.244
R7105 gnd.n4861 gnd.n1195 240.244
R7106 gnd.n4861 gnd.n1203 240.244
R7107 gnd.n4857 gnd.n1203 240.244
R7108 gnd.n4857 gnd.n1169 240.244
R7109 gnd.n4885 gnd.n1169 240.244
R7110 gnd.n4885 gnd.n1165 240.244
R7111 gnd.n4891 gnd.n1165 240.244
R7112 gnd.n4891 gnd.n1153 240.244
R7113 gnd.n4901 gnd.n1153 240.244
R7114 gnd.n4901 gnd.n1149 240.244
R7115 gnd.n4907 gnd.n1149 240.244
R7116 gnd.n4907 gnd.n1135 240.244
R7117 gnd.n4917 gnd.n1135 240.244
R7118 gnd.n4917 gnd.n1131 240.244
R7119 gnd.n4923 gnd.n1131 240.244
R7120 gnd.n4923 gnd.n1119 240.244
R7121 gnd.n4933 gnd.n1119 240.244
R7122 gnd.n4933 gnd.n1115 240.244
R7123 gnd.n4939 gnd.n1115 240.244
R7124 gnd.n4939 gnd.n1101 240.244
R7125 gnd.n4949 gnd.n1101 240.244
R7126 gnd.n4949 gnd.n1097 240.244
R7127 gnd.n4955 gnd.n1097 240.244
R7128 gnd.n4955 gnd.n1085 240.244
R7129 gnd.n4965 gnd.n1085 240.244
R7130 gnd.n4965 gnd.n1081 240.244
R7131 gnd.n4971 gnd.n1081 240.244
R7132 gnd.n4971 gnd.n1066 240.244
R7133 gnd.n4983 gnd.n1066 240.244
R7134 gnd.n4983 gnd.n1062 240.244
R7135 gnd.n6224 gnd.n1062 240.244
R7136 gnd.n6224 gnd.n985 240.244
R7137 gnd.n2552 gnd.n1602 240.244
R7138 gnd.n2546 gnd.n1602 240.244
R7139 gnd.n2546 gnd.n1606 240.244
R7140 gnd.n2542 gnd.n1606 240.244
R7141 gnd.n2542 gnd.n1608 240.244
R7142 gnd.n2538 gnd.n1608 240.244
R7143 gnd.n2538 gnd.n1613 240.244
R7144 gnd.n2534 gnd.n1613 240.244
R7145 gnd.n2534 gnd.n1615 240.244
R7146 gnd.n2530 gnd.n1615 240.244
R7147 gnd.n2530 gnd.n1621 240.244
R7148 gnd.n2526 gnd.n1621 240.244
R7149 gnd.n2526 gnd.n1623 240.244
R7150 gnd.n2522 gnd.n1623 240.244
R7151 gnd.n2522 gnd.n1629 240.244
R7152 gnd.n2518 gnd.n1629 240.244
R7153 gnd.n2518 gnd.n1631 240.244
R7154 gnd.n2514 gnd.n1631 240.244
R7155 gnd.n2514 gnd.n1637 240.244
R7156 gnd.n2510 gnd.n1637 240.244
R7157 gnd.n2510 gnd.n1639 240.244
R7158 gnd.n2506 gnd.n1639 240.244
R7159 gnd.n2506 gnd.n1645 240.244
R7160 gnd.n2502 gnd.n1645 240.244
R7161 gnd.n2502 gnd.n1647 240.244
R7162 gnd.n2498 gnd.n1647 240.244
R7163 gnd.n2498 gnd.n1653 240.244
R7164 gnd.n2494 gnd.n1653 240.244
R7165 gnd.n2494 gnd.n1655 240.244
R7166 gnd.n2490 gnd.n1655 240.244
R7167 gnd.n2490 gnd.n1661 240.244
R7168 gnd.n2486 gnd.n1661 240.244
R7169 gnd.n2486 gnd.n1663 240.244
R7170 gnd.n2482 gnd.n1663 240.244
R7171 gnd.n2482 gnd.n1669 240.244
R7172 gnd.n2478 gnd.n1669 240.244
R7173 gnd.n2478 gnd.n1671 240.244
R7174 gnd.n2474 gnd.n1671 240.244
R7175 gnd.n2474 gnd.n1677 240.244
R7176 gnd.n2470 gnd.n1677 240.244
R7177 gnd.n2470 gnd.n1679 240.244
R7178 gnd.n2466 gnd.n1679 240.244
R7179 gnd.n2466 gnd.n1685 240.244
R7180 gnd.n2462 gnd.n1685 240.244
R7181 gnd.n2462 gnd.n1687 240.244
R7182 gnd.n2458 gnd.n1687 240.244
R7183 gnd.n2458 gnd.n1693 240.244
R7184 gnd.n2454 gnd.n1693 240.244
R7185 gnd.n2454 gnd.n1695 240.244
R7186 gnd.n2450 gnd.n1695 240.244
R7187 gnd.n2450 gnd.n1701 240.244
R7188 gnd.n2446 gnd.n1701 240.244
R7189 gnd.n2446 gnd.n1703 240.244
R7190 gnd.n2442 gnd.n1703 240.244
R7191 gnd.n2442 gnd.n1709 240.244
R7192 gnd.n2438 gnd.n1709 240.244
R7193 gnd.n2438 gnd.n1711 240.244
R7194 gnd.n2434 gnd.n1711 240.244
R7195 gnd.n2434 gnd.n1717 240.244
R7196 gnd.n2430 gnd.n1717 240.244
R7197 gnd.n2430 gnd.n1719 240.244
R7198 gnd.n2426 gnd.n1719 240.244
R7199 gnd.n2426 gnd.n1725 240.244
R7200 gnd.n2422 gnd.n1725 240.244
R7201 gnd.n2422 gnd.n1727 240.244
R7202 gnd.n2418 gnd.n1727 240.244
R7203 gnd.n2418 gnd.n1733 240.244
R7204 gnd.n2414 gnd.n1733 240.244
R7205 gnd.n2414 gnd.n1735 240.244
R7206 gnd.n2410 gnd.n1735 240.244
R7207 gnd.n2410 gnd.n1741 240.244
R7208 gnd.n2406 gnd.n1741 240.244
R7209 gnd.n2406 gnd.n1743 240.244
R7210 gnd.n2402 gnd.n1743 240.244
R7211 gnd.n2402 gnd.n1749 240.244
R7212 gnd.n2398 gnd.n1749 240.244
R7213 gnd.n2398 gnd.n1751 240.244
R7214 gnd.n2394 gnd.n1751 240.244
R7215 gnd.n2394 gnd.n1757 240.244
R7216 gnd.n2390 gnd.n1757 240.244
R7217 gnd.n2390 gnd.n1759 240.244
R7218 gnd.n2386 gnd.n1759 240.244
R7219 gnd.n2386 gnd.n1765 240.244
R7220 gnd.n2382 gnd.n1765 240.244
R7221 gnd.n2382 gnd.n1767 240.244
R7222 gnd.n2378 gnd.n1767 240.244
R7223 gnd.n2378 gnd.n1773 240.244
R7224 gnd.n2374 gnd.n1773 240.244
R7225 gnd.n2374 gnd.n1775 240.244
R7226 gnd.n2370 gnd.n1775 240.244
R7227 gnd.n2370 gnd.n1781 240.244
R7228 gnd.n2366 gnd.n1781 240.244
R7229 gnd.n2366 gnd.n1783 240.244
R7230 gnd.n2362 gnd.n1783 240.244
R7231 gnd.n2362 gnd.n1789 240.244
R7232 gnd.n2358 gnd.n1789 240.244
R7233 gnd.n2358 gnd.n1791 240.244
R7234 gnd.n2354 gnd.n1791 240.244
R7235 gnd.n2354 gnd.n1797 240.244
R7236 gnd.n2350 gnd.n1797 240.244
R7237 gnd.n2350 gnd.n1799 240.244
R7238 gnd.n2346 gnd.n1799 240.244
R7239 gnd.n2346 gnd.n1805 240.244
R7240 gnd.n2342 gnd.n1805 240.244
R7241 gnd.n2342 gnd.n1807 240.244
R7242 gnd.n2338 gnd.n1807 240.244
R7243 gnd.n2338 gnd.n1813 240.244
R7244 gnd.n2334 gnd.n1813 240.244
R7245 gnd.n2334 gnd.n1815 240.244
R7246 gnd.n2330 gnd.n1815 240.244
R7247 gnd.n2330 gnd.n1821 240.244
R7248 gnd.n2326 gnd.n1821 240.244
R7249 gnd.n2326 gnd.n1823 240.244
R7250 gnd.n2322 gnd.n1823 240.244
R7251 gnd.n2322 gnd.n1829 240.244
R7252 gnd.n2318 gnd.n1829 240.244
R7253 gnd.n2318 gnd.n1831 240.244
R7254 gnd.n2314 gnd.n1831 240.244
R7255 gnd.n2314 gnd.n1837 240.244
R7256 gnd.n2310 gnd.n1837 240.244
R7257 gnd.n2310 gnd.n1839 240.244
R7258 gnd.n2306 gnd.n1839 240.244
R7259 gnd.n2306 gnd.n1845 240.244
R7260 gnd.n2302 gnd.n1845 240.244
R7261 gnd.n2302 gnd.n1847 240.244
R7262 gnd.n2298 gnd.n1847 240.244
R7263 gnd.n2298 gnd.n1853 240.244
R7264 gnd.n2294 gnd.n1853 240.244
R7265 gnd.n2294 gnd.n1855 240.244
R7266 gnd.n2290 gnd.n1855 240.244
R7267 gnd.n2290 gnd.n1861 240.244
R7268 gnd.n2286 gnd.n1861 240.244
R7269 gnd.n2286 gnd.n1863 240.244
R7270 gnd.n2282 gnd.n1863 240.244
R7271 gnd.n2282 gnd.n1869 240.244
R7272 gnd.n2278 gnd.n1869 240.244
R7273 gnd.n2278 gnd.n1871 240.244
R7274 gnd.n2274 gnd.n1871 240.244
R7275 gnd.n2274 gnd.n1877 240.244
R7276 gnd.n2270 gnd.n1877 240.244
R7277 gnd.n2270 gnd.n1879 240.244
R7278 gnd.n2266 gnd.n1879 240.244
R7279 gnd.n2266 gnd.n1885 240.244
R7280 gnd.n2262 gnd.n1885 240.244
R7281 gnd.n2262 gnd.n1887 240.244
R7282 gnd.n2258 gnd.n1887 240.244
R7283 gnd.n2258 gnd.n1893 240.244
R7284 gnd.n2254 gnd.n1893 240.244
R7285 gnd.n2254 gnd.n1895 240.244
R7286 gnd.n2250 gnd.n1895 240.244
R7287 gnd.n2250 gnd.n1901 240.244
R7288 gnd.n2246 gnd.n1901 240.244
R7289 gnd.n2246 gnd.n1903 240.244
R7290 gnd.n2242 gnd.n1903 240.244
R7291 gnd.n2238 gnd.n1908 240.244
R7292 gnd.n2238 gnd.n1910 240.244
R7293 gnd.n2232 gnd.n1910 240.244
R7294 gnd.n2232 gnd.n1916 240.244
R7295 gnd.n2228 gnd.n1916 240.244
R7296 gnd.n2228 gnd.n1918 240.244
R7297 gnd.n2224 gnd.n1918 240.244
R7298 gnd.n2224 gnd.n1923 240.244
R7299 gnd.n2220 gnd.n1923 240.244
R7300 gnd.n2220 gnd.n1925 240.244
R7301 gnd.n2216 gnd.n1925 240.244
R7302 gnd.n2216 gnd.n1931 240.244
R7303 gnd.n2212 gnd.n1931 240.244
R7304 gnd.n2212 gnd.n1933 240.244
R7305 gnd.n2208 gnd.n1933 240.244
R7306 gnd.n2208 gnd.n1939 240.244
R7307 gnd.n2204 gnd.n1939 240.244
R7308 gnd.n2204 gnd.n1941 240.244
R7309 gnd.n2200 gnd.n1941 240.244
R7310 gnd.n2200 gnd.n1947 240.244
R7311 gnd.n2196 gnd.n1947 240.244
R7312 gnd.n2196 gnd.n1949 240.244
R7313 gnd.n2192 gnd.n1949 240.244
R7314 gnd.n2192 gnd.n1955 240.244
R7315 gnd.n2188 gnd.n1955 240.244
R7316 gnd.n2188 gnd.n1957 240.244
R7317 gnd.n2184 gnd.n1957 240.244
R7318 gnd.n2184 gnd.n1963 240.244
R7319 gnd.n2180 gnd.n1963 240.244
R7320 gnd.n2180 gnd.n1965 240.244
R7321 gnd.n2176 gnd.n1965 240.244
R7322 gnd.n2176 gnd.n1971 240.244
R7323 gnd.n2172 gnd.n1971 240.244
R7324 gnd.n2172 gnd.n1973 240.244
R7325 gnd.n2168 gnd.n1973 240.244
R7326 gnd.n2168 gnd.n1979 240.244
R7327 gnd.n2164 gnd.n1979 240.244
R7328 gnd.n2164 gnd.n1981 240.244
R7329 gnd.n2160 gnd.n1981 240.244
R7330 gnd.n2160 gnd.n1987 240.244
R7331 gnd.n2156 gnd.n1987 240.244
R7332 gnd.n2156 gnd.n1989 240.244
R7333 gnd.n2152 gnd.n1989 240.244
R7334 gnd.n2152 gnd.n1995 240.244
R7335 gnd.n2148 gnd.n1995 240.244
R7336 gnd.n2148 gnd.n1997 240.244
R7337 gnd.n2144 gnd.n1997 240.244
R7338 gnd.n2144 gnd.n2003 240.244
R7339 gnd.n2140 gnd.n2003 240.244
R7340 gnd.n2140 gnd.n2005 240.244
R7341 gnd.n2136 gnd.n2005 240.244
R7342 gnd.n2136 gnd.n2011 240.244
R7343 gnd.n2132 gnd.n2011 240.244
R7344 gnd.n2132 gnd.n2013 240.244
R7345 gnd.n2128 gnd.n2013 240.244
R7346 gnd.n2128 gnd.n2019 240.244
R7347 gnd.n2124 gnd.n2019 240.244
R7348 gnd.n2124 gnd.n2021 240.244
R7349 gnd.n2120 gnd.n2021 240.244
R7350 gnd.n2120 gnd.n2027 240.244
R7351 gnd.n2116 gnd.n2027 240.244
R7352 gnd.n2116 gnd.n2029 240.244
R7353 gnd.n2112 gnd.n2029 240.244
R7354 gnd.n2112 gnd.n2035 240.244
R7355 gnd.n2108 gnd.n2035 240.244
R7356 gnd.n2108 gnd.n2037 240.244
R7357 gnd.n2104 gnd.n2037 240.244
R7358 gnd.n2104 gnd.n2043 240.244
R7359 gnd.n2100 gnd.n2043 240.244
R7360 gnd.n2100 gnd.n2045 240.244
R7361 gnd.n2096 gnd.n2045 240.244
R7362 gnd.n2096 gnd.n2051 240.244
R7363 gnd.n2092 gnd.n2051 240.244
R7364 gnd.n2092 gnd.n2053 240.244
R7365 gnd.n2088 gnd.n2053 240.244
R7366 gnd.n2088 gnd.n2059 240.244
R7367 gnd.n2084 gnd.n2059 240.244
R7368 gnd.n2084 gnd.n2061 240.244
R7369 gnd.n2080 gnd.n2061 240.244
R7370 gnd.n2080 gnd.n2067 240.244
R7371 gnd.n2076 gnd.n2067 240.244
R7372 gnd.n2076 gnd.n2070 240.244
R7373 gnd.n2070 gnd.n342 240.244
R7374 gnd.n7080 gnd.n342 240.244
R7375 gnd.n4851 gnd.n1210 240.244
R7376 gnd.n4851 gnd.n1211 240.244
R7377 gnd.n4847 gnd.n1211 240.244
R7378 gnd.n4847 gnd.n4846 240.244
R7379 gnd.n4846 gnd.n1217 240.244
R7380 gnd.n4667 gnd.n1217 240.244
R7381 gnd.n4686 gnd.n4667 240.244
R7382 gnd.n4686 gnd.n4668 240.244
R7383 gnd.n4682 gnd.n4668 240.244
R7384 gnd.n4682 gnd.n4681 240.244
R7385 gnd.n4681 gnd.n1261 240.244
R7386 gnd.n4709 gnd.n1261 240.244
R7387 gnd.n4710 gnd.n4709 240.244
R7388 gnd.n4710 gnd.n1256 240.244
R7389 gnd.n4726 gnd.n1256 240.244
R7390 gnd.n4726 gnd.n1257 240.244
R7391 gnd.n4722 gnd.n1257 240.244
R7392 gnd.n4722 gnd.n4721 240.244
R7393 gnd.n4721 gnd.n1251 240.244
R7394 gnd.n4748 gnd.n1251 240.244
R7395 gnd.n4749 gnd.n4748 240.244
R7396 gnd.n4749 gnd.n1246 240.244
R7397 gnd.n4786 gnd.n1246 240.244
R7398 gnd.n4786 gnd.n1247 240.244
R7399 gnd.n4782 gnd.n1247 240.244
R7400 gnd.n4782 gnd.n4781 240.244
R7401 gnd.n4781 gnd.n4780 240.244
R7402 gnd.n4780 gnd.n4757 240.244
R7403 gnd.n4776 gnd.n4757 240.244
R7404 gnd.n4776 gnd.n4775 240.244
R7405 gnd.n4775 gnd.n4774 240.244
R7406 gnd.n4774 gnd.n4764 240.244
R7407 gnd.n4769 gnd.n4764 240.244
R7408 gnd.n4769 gnd.n942 240.244
R7409 gnd.n6338 gnd.n942 240.244
R7410 gnd.n6338 gnd.n938 240.244
R7411 gnd.n6344 gnd.n938 240.244
R7412 gnd.n6344 gnd.n928 240.244
R7413 gnd.n6354 gnd.n928 240.244
R7414 gnd.n6354 gnd.n924 240.244
R7415 gnd.n6360 gnd.n924 240.244
R7416 gnd.n6360 gnd.n914 240.244
R7417 gnd.n6370 gnd.n914 240.244
R7418 gnd.n6370 gnd.n910 240.244
R7419 gnd.n6376 gnd.n910 240.244
R7420 gnd.n6376 gnd.n899 240.244
R7421 gnd.n6386 gnd.n899 240.244
R7422 gnd.n6386 gnd.n895 240.244
R7423 gnd.n6392 gnd.n895 240.244
R7424 gnd.n6392 gnd.n884 240.244
R7425 gnd.n6402 gnd.n884 240.244
R7426 gnd.n6402 gnd.n880 240.244
R7427 gnd.n6408 gnd.n880 240.244
R7428 gnd.n6408 gnd.n868 240.244
R7429 gnd.n6418 gnd.n868 240.244
R7430 gnd.n6418 gnd.n864 240.244
R7431 gnd.n6424 gnd.n864 240.244
R7432 gnd.n6424 gnd.n853 240.244
R7433 gnd.n6434 gnd.n853 240.244
R7434 gnd.n6434 gnd.n849 240.244
R7435 gnd.n6440 gnd.n849 240.244
R7436 gnd.n6440 gnd.n839 240.244
R7437 gnd.n6450 gnd.n839 240.244
R7438 gnd.n6450 gnd.n835 240.244
R7439 gnd.n6456 gnd.n835 240.244
R7440 gnd.n6456 gnd.n824 240.244
R7441 gnd.n6466 gnd.n824 240.244
R7442 gnd.n6466 gnd.n820 240.244
R7443 gnd.n6472 gnd.n820 240.244
R7444 gnd.n6472 gnd.n808 240.244
R7445 gnd.n6482 gnd.n808 240.244
R7446 gnd.n6482 gnd.n804 240.244
R7447 gnd.n6488 gnd.n804 240.244
R7448 gnd.n6488 gnd.n793 240.244
R7449 gnd.n6498 gnd.n793 240.244
R7450 gnd.n6498 gnd.n789 240.244
R7451 gnd.n6504 gnd.n789 240.244
R7452 gnd.n6504 gnd.n778 240.244
R7453 gnd.n6514 gnd.n778 240.244
R7454 gnd.n6514 gnd.n774 240.244
R7455 gnd.n6520 gnd.n774 240.244
R7456 gnd.n6520 gnd.n762 240.244
R7457 gnd.n6530 gnd.n762 240.244
R7458 gnd.n6530 gnd.n758 240.244
R7459 gnd.n6536 gnd.n758 240.244
R7460 gnd.n6536 gnd.n746 240.244
R7461 gnd.n6546 gnd.n746 240.244
R7462 gnd.n6546 gnd.n742 240.244
R7463 gnd.n6552 gnd.n742 240.244
R7464 gnd.n6552 gnd.n732 240.244
R7465 gnd.n6562 gnd.n732 240.244
R7466 gnd.n6562 gnd.n728 240.244
R7467 gnd.n6568 gnd.n728 240.244
R7468 gnd.n6568 gnd.n717 240.244
R7469 gnd.n6578 gnd.n717 240.244
R7470 gnd.n6578 gnd.n713 240.244
R7471 gnd.n6584 gnd.n713 240.244
R7472 gnd.n6584 gnd.n702 240.244
R7473 gnd.n6594 gnd.n702 240.244
R7474 gnd.n6594 gnd.n698 240.244
R7475 gnd.n6600 gnd.n698 240.244
R7476 gnd.n6600 gnd.n688 240.244
R7477 gnd.n6610 gnd.n688 240.244
R7478 gnd.n6610 gnd.n684 240.244
R7479 gnd.n6616 gnd.n684 240.244
R7480 gnd.n6616 gnd.n674 240.244
R7481 gnd.n6626 gnd.n674 240.244
R7482 gnd.n6626 gnd.n670 240.244
R7483 gnd.n6632 gnd.n670 240.244
R7484 gnd.n6632 gnd.n660 240.244
R7485 gnd.n6642 gnd.n660 240.244
R7486 gnd.n6642 gnd.n656 240.244
R7487 gnd.n6648 gnd.n656 240.244
R7488 gnd.n6648 gnd.n645 240.244
R7489 gnd.n6659 gnd.n645 240.244
R7490 gnd.n6659 gnd.n640 240.244
R7491 gnd.n6667 gnd.n640 240.244
R7492 gnd.n6667 gnd.n641 240.244
R7493 gnd.n641 gnd.n615 240.244
R7494 gnd.n6678 gnd.n615 240.244
R7495 gnd.n6678 gnd.n611 240.244
R7496 gnd.n6684 gnd.n611 240.244
R7497 gnd.n6685 gnd.n6684 240.244
R7498 gnd.n6686 gnd.n6685 240.244
R7499 gnd.n6686 gnd.n607 240.244
R7500 gnd.n6692 gnd.n607 240.244
R7501 gnd.n6693 gnd.n6692 240.244
R7502 gnd.n6694 gnd.n6693 240.244
R7503 gnd.n6694 gnd.n603 240.244
R7504 gnd.n6700 gnd.n603 240.244
R7505 gnd.n6727 gnd.n6700 240.244
R7506 gnd.n6728 gnd.n6727 240.244
R7507 gnd.n6728 gnd.n598 240.244
R7508 gnd.n6744 gnd.n598 240.244
R7509 gnd.n6744 gnd.n599 240.244
R7510 gnd.n6740 gnd.n599 240.244
R7511 gnd.n6740 gnd.n6739 240.244
R7512 gnd.n6739 gnd.n593 240.244
R7513 gnd.n6766 gnd.n593 240.244
R7514 gnd.n6767 gnd.n6766 240.244
R7515 gnd.n6767 gnd.n588 240.244
R7516 gnd.n6775 gnd.n588 240.244
R7517 gnd.n6775 gnd.n589 240.244
R7518 gnd.n589 gnd.n393 240.244
R7519 gnd.n7000 gnd.n393 240.244
R7520 gnd.n7000 gnd.n388 240.244
R7521 gnd.n7017 gnd.n388 240.244
R7522 gnd.n7017 gnd.n389 240.244
R7523 gnd.n7013 gnd.n389 240.244
R7524 gnd.n7013 gnd.n7012 240.244
R7525 gnd.n7012 gnd.n348 240.244
R7526 gnd.n7073 gnd.n348 240.244
R7527 gnd.n7074 gnd.n7073 240.244
R7528 gnd.n7074 gnd.n343 240.244
R7529 gnd.n2556 gnd.n1600 240.244
R7530 gnd.n2556 gnd.n1596 240.244
R7531 gnd.n2562 gnd.n1596 240.244
R7532 gnd.n2562 gnd.n1594 240.244
R7533 gnd.n2566 gnd.n1594 240.244
R7534 gnd.n2566 gnd.n1590 240.244
R7535 gnd.n2572 gnd.n1590 240.244
R7536 gnd.n2572 gnd.n1588 240.244
R7537 gnd.n2576 gnd.n1588 240.244
R7538 gnd.n2576 gnd.n1584 240.244
R7539 gnd.n2582 gnd.n1584 240.244
R7540 gnd.n2582 gnd.n1582 240.244
R7541 gnd.n2586 gnd.n1582 240.244
R7542 gnd.n2586 gnd.n1578 240.244
R7543 gnd.n2592 gnd.n1578 240.244
R7544 gnd.n2592 gnd.n1576 240.244
R7545 gnd.n2596 gnd.n1576 240.244
R7546 gnd.n2596 gnd.n1572 240.244
R7547 gnd.n2602 gnd.n1572 240.244
R7548 gnd.n2602 gnd.n1570 240.244
R7549 gnd.n2606 gnd.n1570 240.244
R7550 gnd.n2606 gnd.n1566 240.244
R7551 gnd.n2612 gnd.n1566 240.244
R7552 gnd.n2612 gnd.n1564 240.244
R7553 gnd.n2616 gnd.n1564 240.244
R7554 gnd.n2616 gnd.n1560 240.244
R7555 gnd.n2622 gnd.n1560 240.244
R7556 gnd.n2622 gnd.n1558 240.244
R7557 gnd.n2626 gnd.n1558 240.244
R7558 gnd.n2626 gnd.n1554 240.244
R7559 gnd.n2632 gnd.n1554 240.244
R7560 gnd.n2632 gnd.n1552 240.244
R7561 gnd.n2636 gnd.n1552 240.244
R7562 gnd.n2636 gnd.n1548 240.244
R7563 gnd.n2642 gnd.n1548 240.244
R7564 gnd.n2642 gnd.n1546 240.244
R7565 gnd.n2646 gnd.n1546 240.244
R7566 gnd.n2646 gnd.n1542 240.244
R7567 gnd.n2652 gnd.n1542 240.244
R7568 gnd.n2652 gnd.n1540 240.244
R7569 gnd.n2656 gnd.n1540 240.244
R7570 gnd.n2656 gnd.n1536 240.244
R7571 gnd.n2662 gnd.n1536 240.244
R7572 gnd.n2662 gnd.n1534 240.244
R7573 gnd.n2666 gnd.n1534 240.244
R7574 gnd.n2666 gnd.n1530 240.244
R7575 gnd.n2672 gnd.n1530 240.244
R7576 gnd.n2672 gnd.n1528 240.244
R7577 gnd.n2676 gnd.n1528 240.244
R7578 gnd.n2676 gnd.n1524 240.244
R7579 gnd.n2682 gnd.n1524 240.244
R7580 gnd.n2682 gnd.n1522 240.244
R7581 gnd.n2686 gnd.n1522 240.244
R7582 gnd.n2686 gnd.n1518 240.244
R7583 gnd.n2692 gnd.n1518 240.244
R7584 gnd.n2692 gnd.n1516 240.244
R7585 gnd.n2696 gnd.n1516 240.244
R7586 gnd.n2696 gnd.n1512 240.244
R7587 gnd.n2702 gnd.n1512 240.244
R7588 gnd.n2702 gnd.n1510 240.244
R7589 gnd.n2706 gnd.n1510 240.244
R7590 gnd.n2706 gnd.n1506 240.244
R7591 gnd.n2712 gnd.n1506 240.244
R7592 gnd.n2712 gnd.n1504 240.244
R7593 gnd.n2716 gnd.n1504 240.244
R7594 gnd.n2716 gnd.n1500 240.244
R7595 gnd.n2722 gnd.n1500 240.244
R7596 gnd.n2722 gnd.n1498 240.244
R7597 gnd.n2726 gnd.n1498 240.244
R7598 gnd.n2726 gnd.n1494 240.244
R7599 gnd.n2732 gnd.n1494 240.244
R7600 gnd.n2732 gnd.n1492 240.244
R7601 gnd.n2736 gnd.n1492 240.244
R7602 gnd.n2736 gnd.n1488 240.244
R7603 gnd.n2742 gnd.n1488 240.244
R7604 gnd.n2742 gnd.n1486 240.244
R7605 gnd.n2746 gnd.n1486 240.244
R7606 gnd.n2746 gnd.n1482 240.244
R7607 gnd.n2752 gnd.n1482 240.244
R7608 gnd.n2752 gnd.n1480 240.244
R7609 gnd.n2756 gnd.n1480 240.244
R7610 gnd.n2756 gnd.n1475 240.244
R7611 gnd.n2765 gnd.n1475 240.244
R7612 gnd.n2765 gnd.n1476 240.244
R7613 gnd.n5094 gnd.n937 240.244
R7614 gnd.n5095 gnd.n937 240.244
R7615 gnd.n5095 gnd.n930 240.244
R7616 gnd.n5098 gnd.n930 240.244
R7617 gnd.n5098 gnd.n922 240.244
R7618 gnd.n5099 gnd.n922 240.244
R7619 gnd.n5099 gnd.n915 240.244
R7620 gnd.n5102 gnd.n915 240.244
R7621 gnd.n5102 gnd.n908 240.244
R7622 gnd.n5103 gnd.n908 240.244
R7623 gnd.n5103 gnd.n900 240.244
R7624 gnd.n5106 gnd.n900 240.244
R7625 gnd.n5106 gnd.n894 240.244
R7626 gnd.n5107 gnd.n894 240.244
R7627 gnd.n5107 gnd.n886 240.244
R7628 gnd.n5110 gnd.n886 240.244
R7629 gnd.n5110 gnd.n878 240.244
R7630 gnd.n5111 gnd.n878 240.244
R7631 gnd.n5111 gnd.n870 240.244
R7632 gnd.n5114 gnd.n870 240.244
R7633 gnd.n5114 gnd.n863 240.244
R7634 gnd.n5115 gnd.n863 240.244
R7635 gnd.n5115 gnd.n855 240.244
R7636 gnd.n5118 gnd.n855 240.244
R7637 gnd.n5118 gnd.n847 240.244
R7638 gnd.n5119 gnd.n847 240.244
R7639 gnd.n5119 gnd.n840 240.244
R7640 gnd.n5122 gnd.n840 240.244
R7641 gnd.n5122 gnd.n833 240.244
R7642 gnd.n5123 gnd.n833 240.244
R7643 gnd.n5123 gnd.n826 240.244
R7644 gnd.n5126 gnd.n826 240.244
R7645 gnd.n5126 gnd.n818 240.244
R7646 gnd.n5127 gnd.n818 240.244
R7647 gnd.n5127 gnd.n810 240.244
R7648 gnd.n5130 gnd.n810 240.244
R7649 gnd.n5130 gnd.n802 240.244
R7650 gnd.n5131 gnd.n802 240.244
R7651 gnd.n5131 gnd.n794 240.244
R7652 gnd.n5134 gnd.n794 240.244
R7653 gnd.n5134 gnd.n787 240.244
R7654 gnd.n5135 gnd.n787 240.244
R7655 gnd.n5135 gnd.n780 240.244
R7656 gnd.n5138 gnd.n780 240.244
R7657 gnd.n5138 gnd.n772 240.244
R7658 gnd.n5139 gnd.n772 240.244
R7659 gnd.n5139 gnd.n764 240.244
R7660 gnd.n5142 gnd.n764 240.244
R7661 gnd.n5142 gnd.n756 240.244
R7662 gnd.n5143 gnd.n756 240.244
R7663 gnd.n5143 gnd.n748 240.244
R7664 gnd.n5146 gnd.n748 240.244
R7665 gnd.n5146 gnd.n741 240.244
R7666 gnd.n5147 gnd.n741 240.244
R7667 gnd.n5147 gnd.n734 240.244
R7668 gnd.n5150 gnd.n734 240.244
R7669 gnd.n5150 gnd.n727 240.244
R7670 gnd.n5151 gnd.n727 240.244
R7671 gnd.n5151 gnd.n719 240.244
R7672 gnd.n5154 gnd.n719 240.244
R7673 gnd.n5154 gnd.n711 240.244
R7674 gnd.n5155 gnd.n711 240.244
R7675 gnd.n5155 gnd.n704 240.244
R7676 gnd.n5158 gnd.n704 240.244
R7677 gnd.n5158 gnd.n697 240.244
R7678 gnd.n5159 gnd.n697 240.244
R7679 gnd.n5159 gnd.n689 240.244
R7680 gnd.n5936 gnd.n689 240.244
R7681 gnd.n5936 gnd.n682 240.244
R7682 gnd.n5938 gnd.n682 240.244
R7683 gnd.n5938 gnd.n675 240.244
R7684 gnd.n5941 gnd.n675 240.244
R7685 gnd.n5941 gnd.n669 240.244
R7686 gnd.n5942 gnd.n669 240.244
R7687 gnd.n5942 gnd.n662 240.244
R7688 gnd.n5945 gnd.n662 240.244
R7689 gnd.n5945 gnd.n655 240.244
R7690 gnd.n5946 gnd.n655 240.244
R7691 gnd.n5946 gnd.n647 240.244
R7692 gnd.n5949 gnd.n647 240.244
R7693 gnd.n5949 gnd.n638 240.244
R7694 gnd.n6094 gnd.n638 240.244
R7695 gnd.n4993 gnd.n4992 240.244
R7696 gnd.n5009 gnd.n5008 240.244
R7697 gnd.n5019 gnd.n5018 240.244
R7698 gnd.n5021 gnd.n5020 240.244
R7699 gnd.n5032 gnd.n5031 240.244
R7700 gnd.n5042 gnd.n5041 240.244
R7701 gnd.n5044 gnd.n5043 240.244
R7702 gnd.n974 gnd.n973 240.244
R7703 gnd.n6311 gnd.n6310 240.244
R7704 gnd.n969 gnd.n968 240.244
R7705 gnd.n6320 gnd.n6319 240.244
R7706 gnd.n965 gnd.n964 240.244
R7707 gnd.n6329 gnd.n6328 240.244
R7708 gnd.n6335 gnd.n958 240.244
R7709 gnd.n6346 gnd.n935 240.244
R7710 gnd.n6346 gnd.n931 240.244
R7711 gnd.n6352 gnd.n931 240.244
R7712 gnd.n6352 gnd.n920 240.244
R7713 gnd.n6362 gnd.n920 240.244
R7714 gnd.n6362 gnd.n916 240.244
R7715 gnd.n6368 gnd.n916 240.244
R7716 gnd.n6368 gnd.n906 240.244
R7717 gnd.n6378 gnd.n906 240.244
R7718 gnd.n6378 gnd.n902 240.244
R7719 gnd.n6384 gnd.n902 240.244
R7720 gnd.n6384 gnd.n892 240.244
R7721 gnd.n6394 gnd.n892 240.244
R7722 gnd.n6394 gnd.n888 240.244
R7723 gnd.n6400 gnd.n888 240.244
R7724 gnd.n6400 gnd.n876 240.244
R7725 gnd.n6410 gnd.n876 240.244
R7726 gnd.n6410 gnd.n872 240.244
R7727 gnd.n6416 gnd.n872 240.244
R7728 gnd.n6416 gnd.n861 240.244
R7729 gnd.n6426 gnd.n861 240.244
R7730 gnd.n6426 gnd.n857 240.244
R7731 gnd.n6432 gnd.n857 240.244
R7732 gnd.n6432 gnd.n846 240.244
R7733 gnd.n6442 gnd.n846 240.244
R7734 gnd.n6442 gnd.n842 240.244
R7735 gnd.n6448 gnd.n842 240.244
R7736 gnd.n6448 gnd.n832 240.244
R7737 gnd.n6458 gnd.n832 240.244
R7738 gnd.n6458 gnd.n828 240.244
R7739 gnd.n6464 gnd.n828 240.244
R7740 gnd.n6464 gnd.n816 240.244
R7741 gnd.n6474 gnd.n816 240.244
R7742 gnd.n6474 gnd.n812 240.244
R7743 gnd.n6480 gnd.n812 240.244
R7744 gnd.n6480 gnd.n800 240.244
R7745 gnd.n6490 gnd.n800 240.244
R7746 gnd.n6490 gnd.n796 240.244
R7747 gnd.n6496 gnd.n796 240.244
R7748 gnd.n6496 gnd.n785 240.244
R7749 gnd.n6506 gnd.n785 240.244
R7750 gnd.n6506 gnd.n781 240.244
R7751 gnd.n6512 gnd.n781 240.244
R7752 gnd.n6512 gnd.n770 240.244
R7753 gnd.n6522 gnd.n770 240.244
R7754 gnd.n6522 gnd.n766 240.244
R7755 gnd.n6528 gnd.n766 240.244
R7756 gnd.n6528 gnd.n754 240.244
R7757 gnd.n6538 gnd.n754 240.244
R7758 gnd.n6538 gnd.n750 240.244
R7759 gnd.n6544 gnd.n750 240.244
R7760 gnd.n6544 gnd.n739 240.244
R7761 gnd.n6554 gnd.n739 240.244
R7762 gnd.n6554 gnd.n735 240.244
R7763 gnd.n6560 gnd.n735 240.244
R7764 gnd.n6560 gnd.n725 240.244
R7765 gnd.n6570 gnd.n725 240.244
R7766 gnd.n6570 gnd.n721 240.244
R7767 gnd.n6576 gnd.n721 240.244
R7768 gnd.n6576 gnd.n710 240.244
R7769 gnd.n6586 gnd.n710 240.244
R7770 gnd.n6586 gnd.n706 240.244
R7771 gnd.n6592 gnd.n706 240.244
R7772 gnd.n6592 gnd.n695 240.244
R7773 gnd.n6602 gnd.n695 240.244
R7774 gnd.n6602 gnd.n691 240.244
R7775 gnd.n6608 gnd.n691 240.244
R7776 gnd.n6608 gnd.n680 240.244
R7777 gnd.n6618 gnd.n680 240.244
R7778 gnd.n6618 gnd.n676 240.244
R7779 gnd.n6624 gnd.n676 240.244
R7780 gnd.n6624 gnd.n667 240.244
R7781 gnd.n6634 gnd.n667 240.244
R7782 gnd.n6634 gnd.n663 240.244
R7783 gnd.n6640 gnd.n663 240.244
R7784 gnd.n6640 gnd.n653 240.244
R7785 gnd.n6650 gnd.n653 240.244
R7786 gnd.n6650 gnd.n649 240.244
R7787 gnd.n6657 gnd.n649 240.244
R7788 gnd.n6657 gnd.n637 240.244
R7789 gnd.n6669 gnd.n637 240.244
R7790 gnd.n6669 gnd.n632 240.244
R7791 gnd.n5966 gnd.n5965 240.244
R7792 gnd.n5968 gnd.n5967 240.244
R7793 gnd.n5976 gnd.n5975 240.244
R7794 gnd.n5986 gnd.n5985 240.244
R7795 gnd.n5988 gnd.n5987 240.244
R7796 gnd.n5996 gnd.n5995 240.244
R7797 gnd.n6006 gnd.n6005 240.244
R7798 gnd.n6008 gnd.n6007 240.244
R7799 gnd.n6013 gnd.n6012 240.244
R7800 gnd.n6015 gnd.n6014 240.244
R7801 gnd.n6019 gnd.n6018 240.244
R7802 gnd.n6021 gnd.n6020 240.244
R7803 gnd.n6028 gnd.n6027 240.244
R7804 gnd.n6675 gnd.n631 240.244
R7805 gnd.n5415 gnd.n5414 240.132
R7806 gnd.n5177 gnd.n5176 240.132
R7807 gnd.n2553 gnd.n1601 225.874
R7808 gnd.n2545 gnd.n1601 225.874
R7809 gnd.n2545 gnd.n2544 225.874
R7810 gnd.n2544 gnd.n2543 225.874
R7811 gnd.n2543 gnd.n1607 225.874
R7812 gnd.n2537 gnd.n1607 225.874
R7813 gnd.n2537 gnd.n2536 225.874
R7814 gnd.n2536 gnd.n2535 225.874
R7815 gnd.n2535 gnd.n1614 225.874
R7816 gnd.n2529 gnd.n1614 225.874
R7817 gnd.n2529 gnd.n2528 225.874
R7818 gnd.n2528 gnd.n2527 225.874
R7819 gnd.n2527 gnd.n1622 225.874
R7820 gnd.n2521 gnd.n1622 225.874
R7821 gnd.n2521 gnd.n2520 225.874
R7822 gnd.n2520 gnd.n2519 225.874
R7823 gnd.n2519 gnd.n1630 225.874
R7824 gnd.n2513 gnd.n1630 225.874
R7825 gnd.n2513 gnd.n2512 225.874
R7826 gnd.n2512 gnd.n2511 225.874
R7827 gnd.n2511 gnd.n1638 225.874
R7828 gnd.n2505 gnd.n1638 225.874
R7829 gnd.n2505 gnd.n2504 225.874
R7830 gnd.n2504 gnd.n2503 225.874
R7831 gnd.n2503 gnd.n1646 225.874
R7832 gnd.n2497 gnd.n1646 225.874
R7833 gnd.n2497 gnd.n2496 225.874
R7834 gnd.n2496 gnd.n2495 225.874
R7835 gnd.n2495 gnd.n1654 225.874
R7836 gnd.n2489 gnd.n1654 225.874
R7837 gnd.n2489 gnd.n2488 225.874
R7838 gnd.n2488 gnd.n2487 225.874
R7839 gnd.n2487 gnd.n1662 225.874
R7840 gnd.n2481 gnd.n1662 225.874
R7841 gnd.n2481 gnd.n2480 225.874
R7842 gnd.n2480 gnd.n2479 225.874
R7843 gnd.n2479 gnd.n1670 225.874
R7844 gnd.n2473 gnd.n1670 225.874
R7845 gnd.n2473 gnd.n2472 225.874
R7846 gnd.n2472 gnd.n2471 225.874
R7847 gnd.n2471 gnd.n1678 225.874
R7848 gnd.n2465 gnd.n1678 225.874
R7849 gnd.n2465 gnd.n2464 225.874
R7850 gnd.n2464 gnd.n2463 225.874
R7851 gnd.n2463 gnd.n1686 225.874
R7852 gnd.n2457 gnd.n1686 225.874
R7853 gnd.n2457 gnd.n2456 225.874
R7854 gnd.n2456 gnd.n2455 225.874
R7855 gnd.n2455 gnd.n1694 225.874
R7856 gnd.n2449 gnd.n1694 225.874
R7857 gnd.n2449 gnd.n2448 225.874
R7858 gnd.n2448 gnd.n2447 225.874
R7859 gnd.n2447 gnd.n1702 225.874
R7860 gnd.n2441 gnd.n1702 225.874
R7861 gnd.n2441 gnd.n2440 225.874
R7862 gnd.n2440 gnd.n2439 225.874
R7863 gnd.n2439 gnd.n1710 225.874
R7864 gnd.n2433 gnd.n1710 225.874
R7865 gnd.n2433 gnd.n2432 225.874
R7866 gnd.n2432 gnd.n2431 225.874
R7867 gnd.n2431 gnd.n1718 225.874
R7868 gnd.n2425 gnd.n1718 225.874
R7869 gnd.n2425 gnd.n2424 225.874
R7870 gnd.n2424 gnd.n2423 225.874
R7871 gnd.n2423 gnd.n1726 225.874
R7872 gnd.n2417 gnd.n1726 225.874
R7873 gnd.n2417 gnd.n2416 225.874
R7874 gnd.n2416 gnd.n2415 225.874
R7875 gnd.n2415 gnd.n1734 225.874
R7876 gnd.n2409 gnd.n1734 225.874
R7877 gnd.n2409 gnd.n2408 225.874
R7878 gnd.n2408 gnd.n2407 225.874
R7879 gnd.n2407 gnd.n1742 225.874
R7880 gnd.n2401 gnd.n1742 225.874
R7881 gnd.n2401 gnd.n2400 225.874
R7882 gnd.n2400 gnd.n2399 225.874
R7883 gnd.n2399 gnd.n1750 225.874
R7884 gnd.n2393 gnd.n1750 225.874
R7885 gnd.n2393 gnd.n2392 225.874
R7886 gnd.n2392 gnd.n2391 225.874
R7887 gnd.n2391 gnd.n1758 225.874
R7888 gnd.n2385 gnd.n1758 225.874
R7889 gnd.n2385 gnd.n2384 225.874
R7890 gnd.n2384 gnd.n2383 225.874
R7891 gnd.n2383 gnd.n1766 225.874
R7892 gnd.n2377 gnd.n1766 225.874
R7893 gnd.n2377 gnd.n2376 225.874
R7894 gnd.n2376 gnd.n2375 225.874
R7895 gnd.n2375 gnd.n1774 225.874
R7896 gnd.n2369 gnd.n1774 225.874
R7897 gnd.n2369 gnd.n2368 225.874
R7898 gnd.n2368 gnd.n2367 225.874
R7899 gnd.n2367 gnd.n1782 225.874
R7900 gnd.n2361 gnd.n1782 225.874
R7901 gnd.n2361 gnd.n2360 225.874
R7902 gnd.n2360 gnd.n2359 225.874
R7903 gnd.n2359 gnd.n1790 225.874
R7904 gnd.n2353 gnd.n1790 225.874
R7905 gnd.n2353 gnd.n2352 225.874
R7906 gnd.n2352 gnd.n2351 225.874
R7907 gnd.n2351 gnd.n1798 225.874
R7908 gnd.n2345 gnd.n1798 225.874
R7909 gnd.n2345 gnd.n2344 225.874
R7910 gnd.n2344 gnd.n2343 225.874
R7911 gnd.n2343 gnd.n1806 225.874
R7912 gnd.n2337 gnd.n1806 225.874
R7913 gnd.n2337 gnd.n2336 225.874
R7914 gnd.n2336 gnd.n2335 225.874
R7915 gnd.n2335 gnd.n1814 225.874
R7916 gnd.n2329 gnd.n1814 225.874
R7917 gnd.n2329 gnd.n2328 225.874
R7918 gnd.n2328 gnd.n2327 225.874
R7919 gnd.n2327 gnd.n1822 225.874
R7920 gnd.n2321 gnd.n1822 225.874
R7921 gnd.n2321 gnd.n2320 225.874
R7922 gnd.n2320 gnd.n2319 225.874
R7923 gnd.n2319 gnd.n1830 225.874
R7924 gnd.n2313 gnd.n1830 225.874
R7925 gnd.n2313 gnd.n2312 225.874
R7926 gnd.n2312 gnd.n2311 225.874
R7927 gnd.n2311 gnd.n1838 225.874
R7928 gnd.n2305 gnd.n1838 225.874
R7929 gnd.n2305 gnd.n2304 225.874
R7930 gnd.n2304 gnd.n2303 225.874
R7931 gnd.n2303 gnd.n1846 225.874
R7932 gnd.n2297 gnd.n1846 225.874
R7933 gnd.n2297 gnd.n2296 225.874
R7934 gnd.n2296 gnd.n2295 225.874
R7935 gnd.n2295 gnd.n1854 225.874
R7936 gnd.n2289 gnd.n1854 225.874
R7937 gnd.n2289 gnd.n2288 225.874
R7938 gnd.n2288 gnd.n2287 225.874
R7939 gnd.n2287 gnd.n1862 225.874
R7940 gnd.n2281 gnd.n1862 225.874
R7941 gnd.n2281 gnd.n2280 225.874
R7942 gnd.n2280 gnd.n2279 225.874
R7943 gnd.n2279 gnd.n1870 225.874
R7944 gnd.n2273 gnd.n1870 225.874
R7945 gnd.n2273 gnd.n2272 225.874
R7946 gnd.n2272 gnd.n2271 225.874
R7947 gnd.n2271 gnd.n1878 225.874
R7948 gnd.n2265 gnd.n1878 225.874
R7949 gnd.n2265 gnd.n2264 225.874
R7950 gnd.n2264 gnd.n2263 225.874
R7951 gnd.n2263 gnd.n1886 225.874
R7952 gnd.n2257 gnd.n1886 225.874
R7953 gnd.n2257 gnd.n2256 225.874
R7954 gnd.n2256 gnd.n2255 225.874
R7955 gnd.n2255 gnd.n1894 225.874
R7956 gnd.n2249 gnd.n1894 225.874
R7957 gnd.n2249 gnd.n2248 225.874
R7958 gnd.n2248 gnd.n2247 225.874
R7959 gnd.n2247 gnd.n1902 225.874
R7960 gnd.n2241 gnd.n1902 225.874
R7961 gnd.n3324 gnd.t107 224.174
R7962 gnd.n1465 gnd.t62 224.174
R7963 gnd.n535 gnd.n496 199.319
R7964 gnd.n535 gnd.n497 199.319
R7965 gnd.n6270 gnd.n6269 199.319
R7966 gnd.n6269 gnd.n6268 199.319
R7967 gnd.n5416 gnd.n5413 186.49
R7968 gnd.n5178 gnd.n5175 186.49
R7969 gnd.n4038 gnd.n4037 185
R7970 gnd.n4036 gnd.n4035 185
R7971 gnd.n4015 gnd.n4014 185
R7972 gnd.n4030 gnd.n4029 185
R7973 gnd.n4028 gnd.n4027 185
R7974 gnd.n4019 gnd.n4018 185
R7975 gnd.n4022 gnd.n4021 185
R7976 gnd.n4006 gnd.n4005 185
R7977 gnd.n4004 gnd.n4003 185
R7978 gnd.n3983 gnd.n3982 185
R7979 gnd.n3998 gnd.n3997 185
R7980 gnd.n3996 gnd.n3995 185
R7981 gnd.n3987 gnd.n3986 185
R7982 gnd.n3990 gnd.n3989 185
R7983 gnd.n3974 gnd.n3973 185
R7984 gnd.n3972 gnd.n3971 185
R7985 gnd.n3951 gnd.n3950 185
R7986 gnd.n3966 gnd.n3965 185
R7987 gnd.n3964 gnd.n3963 185
R7988 gnd.n3955 gnd.n3954 185
R7989 gnd.n3958 gnd.n3957 185
R7990 gnd.n3943 gnd.n3942 185
R7991 gnd.n3941 gnd.n3940 185
R7992 gnd.n3920 gnd.n3919 185
R7993 gnd.n3935 gnd.n3934 185
R7994 gnd.n3933 gnd.n3932 185
R7995 gnd.n3924 gnd.n3923 185
R7996 gnd.n3927 gnd.n3926 185
R7997 gnd.n3911 gnd.n3910 185
R7998 gnd.n3909 gnd.n3908 185
R7999 gnd.n3888 gnd.n3887 185
R8000 gnd.n3903 gnd.n3902 185
R8001 gnd.n3901 gnd.n3900 185
R8002 gnd.n3892 gnd.n3891 185
R8003 gnd.n3895 gnd.n3894 185
R8004 gnd.n3879 gnd.n3878 185
R8005 gnd.n3877 gnd.n3876 185
R8006 gnd.n3856 gnd.n3855 185
R8007 gnd.n3871 gnd.n3870 185
R8008 gnd.n3869 gnd.n3868 185
R8009 gnd.n3860 gnd.n3859 185
R8010 gnd.n3863 gnd.n3862 185
R8011 gnd.n3847 gnd.n3846 185
R8012 gnd.n3845 gnd.n3844 185
R8013 gnd.n3824 gnd.n3823 185
R8014 gnd.n3839 gnd.n3838 185
R8015 gnd.n3837 gnd.n3836 185
R8016 gnd.n3828 gnd.n3827 185
R8017 gnd.n3831 gnd.n3830 185
R8018 gnd.n3816 gnd.n3815 185
R8019 gnd.n3814 gnd.n3813 185
R8020 gnd.n3793 gnd.n3792 185
R8021 gnd.n3808 gnd.n3807 185
R8022 gnd.n3806 gnd.n3805 185
R8023 gnd.n3797 gnd.n3796 185
R8024 gnd.n3800 gnd.n3799 185
R8025 gnd.n3325 gnd.t106 178.987
R8026 gnd.n1466 gnd.t63 178.987
R8027 gnd.n1 gnd.t343 170.774
R8028 gnd.n7 gnd.t166 170.103
R8029 gnd.n6 gnd.t345 170.103
R8030 gnd.n5 gnd.t339 170.103
R8031 gnd.n4 gnd.t153 170.103
R8032 gnd.n3 gnd.t347 170.103
R8033 gnd.n2 gnd.t146 170.103
R8034 gnd.n1 gnd.t168 170.103
R8035 gnd.n5926 gnd.n5925 163.367
R8036 gnd.n5923 gnd.n5187 163.367
R8037 gnd.n5919 gnd.n5918 163.367
R8038 gnd.n5916 gnd.n5190 163.367
R8039 gnd.n5912 gnd.n5911 163.367
R8040 gnd.n5909 gnd.n5193 163.367
R8041 gnd.n5905 gnd.n5904 163.367
R8042 gnd.n5902 gnd.n5196 163.367
R8043 gnd.n5898 gnd.n5897 163.367
R8044 gnd.n5895 gnd.n5199 163.367
R8045 gnd.n5891 gnd.n5890 163.367
R8046 gnd.n5888 gnd.n5202 163.367
R8047 gnd.n5884 gnd.n5883 163.367
R8048 gnd.n5881 gnd.n5205 163.367
R8049 gnd.n5876 gnd.n5875 163.367
R8050 gnd.n5873 gnd.n5871 163.367
R8051 gnd.n5868 gnd.n5867 163.367
R8052 gnd.n5865 gnd.n5211 163.367
R8053 gnd.n5860 gnd.n5859 163.367
R8054 gnd.n5857 gnd.n5216 163.367
R8055 gnd.n5853 gnd.n5852 163.367
R8056 gnd.n5850 gnd.n5219 163.367
R8057 gnd.n5846 gnd.n5845 163.367
R8058 gnd.n5843 gnd.n5222 163.367
R8059 gnd.n5839 gnd.n5838 163.367
R8060 gnd.n5836 gnd.n5225 163.367
R8061 gnd.n5832 gnd.n5831 163.367
R8062 gnd.n5829 gnd.n5228 163.367
R8063 gnd.n5825 gnd.n5824 163.367
R8064 gnd.n5822 gnd.n5231 163.367
R8065 gnd.n5818 gnd.n5817 163.367
R8066 gnd.n5815 gnd.n5234 163.367
R8067 gnd.n5566 gnd.n5368 163.367
R8068 gnd.n5566 gnd.n5369 163.367
R8069 gnd.n5369 gnd.n5360 163.367
R8070 gnd.n5577 gnd.n5360 163.367
R8071 gnd.n5578 gnd.n5577 163.367
R8072 gnd.n5578 gnd.n5357 163.367
R8073 gnd.n5584 gnd.n5357 163.367
R8074 gnd.n5584 gnd.n5358 163.367
R8075 gnd.n5358 gnd.n5350 163.367
R8076 gnd.n5595 gnd.n5350 163.367
R8077 gnd.n5596 gnd.n5595 163.367
R8078 gnd.n5596 gnd.n5347 163.367
R8079 gnd.n5601 gnd.n5347 163.367
R8080 gnd.n5601 gnd.n5348 163.367
R8081 gnd.n5348 gnd.n5340 163.367
R8082 gnd.n5611 gnd.n5340 163.367
R8083 gnd.n5611 gnd.n5337 163.367
R8084 gnd.n5618 gnd.n5337 163.367
R8085 gnd.n5618 gnd.n5338 163.367
R8086 gnd.n5614 gnd.n5338 163.367
R8087 gnd.n5614 gnd.n5330 163.367
R8088 gnd.n5630 gnd.n5330 163.367
R8089 gnd.n5630 gnd.n5327 163.367
R8090 gnd.n5636 gnd.n5327 163.367
R8091 gnd.n5636 gnd.n5328 163.367
R8092 gnd.n5328 gnd.n5321 163.367
R8093 gnd.n5648 gnd.n5321 163.367
R8094 gnd.n5649 gnd.n5648 163.367
R8095 gnd.n5649 gnd.n5318 163.367
R8096 gnd.n5655 gnd.n5318 163.367
R8097 gnd.n5655 gnd.n5319 163.367
R8098 gnd.n5319 gnd.n5311 163.367
R8099 gnd.n5668 gnd.n5311 163.367
R8100 gnd.n5669 gnd.n5668 163.367
R8101 gnd.n5670 gnd.n5669 163.367
R8102 gnd.n5670 gnd.n5309 163.367
R8103 gnd.n5675 gnd.n5309 163.367
R8104 gnd.n5675 gnd.n5301 163.367
R8105 gnd.n5685 gnd.n5301 163.367
R8106 gnd.n5686 gnd.n5685 163.367
R8107 gnd.n5686 gnd.n5298 163.367
R8108 gnd.n5692 gnd.n5298 163.367
R8109 gnd.n5692 gnd.n5299 163.367
R8110 gnd.n5299 gnd.n5290 163.367
R8111 gnd.n5703 gnd.n5290 163.367
R8112 gnd.n5704 gnd.n5703 163.367
R8113 gnd.n5704 gnd.n5287 163.367
R8114 gnd.n5710 gnd.n5287 163.367
R8115 gnd.n5710 gnd.n5288 163.367
R8116 gnd.n5288 gnd.n5280 163.367
R8117 gnd.n5721 gnd.n5280 163.367
R8118 gnd.n5722 gnd.n5721 163.367
R8119 gnd.n5722 gnd.n5277 163.367
R8120 gnd.n5728 gnd.n5277 163.367
R8121 gnd.n5728 gnd.n5278 163.367
R8122 gnd.n5278 gnd.n5270 163.367
R8123 gnd.n5739 gnd.n5270 163.367
R8124 gnd.n5740 gnd.n5739 163.367
R8125 gnd.n5740 gnd.n5267 163.367
R8126 gnd.n5745 gnd.n5267 163.367
R8127 gnd.n5745 gnd.n5268 163.367
R8128 gnd.n5268 gnd.n5260 163.367
R8129 gnd.n5755 gnd.n5260 163.367
R8130 gnd.n5755 gnd.n5257 163.367
R8131 gnd.n5762 gnd.n5257 163.367
R8132 gnd.n5762 gnd.n5258 163.367
R8133 gnd.n5758 gnd.n5258 163.367
R8134 gnd.n5758 gnd.n5250 163.367
R8135 gnd.n5774 gnd.n5250 163.367
R8136 gnd.n5774 gnd.n5247 163.367
R8137 gnd.n5779 gnd.n5247 163.367
R8138 gnd.n5779 gnd.n5248 163.367
R8139 gnd.n5248 gnd.n5242 163.367
R8140 gnd.n5789 gnd.n5242 163.367
R8141 gnd.n5789 gnd.n5240 163.367
R8142 gnd.n5794 gnd.n5240 163.367
R8143 gnd.n5794 gnd.n5236 163.367
R8144 gnd.n5804 gnd.n5236 163.367
R8145 gnd.n5805 gnd.n5804 163.367
R8146 gnd.n5805 gnd.n5162 163.367
R8147 gnd.n5810 gnd.n5162 163.367
R8148 gnd.n5435 gnd.n5434 163.367
R8149 gnd.n5437 gnd.n5435 163.367
R8150 gnd.n5441 gnd.n5406 163.367
R8151 gnd.n5445 gnd.n5443 163.367
R8152 gnd.n5449 gnd.n5404 163.367
R8153 gnd.n5453 gnd.n5451 163.367
R8154 gnd.n5457 gnd.n5402 163.367
R8155 gnd.n5461 gnd.n5459 163.367
R8156 gnd.n5465 gnd.n5400 163.367
R8157 gnd.n5469 gnd.n5467 163.367
R8158 gnd.n5473 gnd.n5398 163.367
R8159 gnd.n5477 gnd.n5475 163.367
R8160 gnd.n5481 gnd.n5396 163.367
R8161 gnd.n5485 gnd.n5483 163.367
R8162 gnd.n5490 gnd.n5392 163.367
R8163 gnd.n5493 gnd.n5492 163.367
R8164 gnd.n5498 gnd.n5388 163.367
R8165 gnd.n5502 gnd.n5500 163.367
R8166 gnd.n5507 gnd.n5384 163.367
R8167 gnd.n5511 gnd.n5509 163.367
R8168 gnd.n5515 gnd.n5382 163.367
R8169 gnd.n5519 gnd.n5517 163.367
R8170 gnd.n5523 gnd.n5380 163.367
R8171 gnd.n5527 gnd.n5525 163.367
R8172 gnd.n5531 gnd.n5378 163.367
R8173 gnd.n5535 gnd.n5533 163.367
R8174 gnd.n5539 gnd.n5376 163.367
R8175 gnd.n5543 gnd.n5541 163.367
R8176 gnd.n5547 gnd.n5374 163.367
R8177 gnd.n5551 gnd.n5549 163.367
R8178 gnd.n5555 gnd.n5372 163.367
R8179 gnd.n5558 gnd.n5557 163.367
R8180 gnd.n5568 gnd.n5365 163.367
R8181 gnd.n5569 gnd.n5568 163.367
R8182 gnd.n5569 gnd.n5362 163.367
R8183 gnd.n5575 gnd.n5362 163.367
R8184 gnd.n5575 gnd.n5363 163.367
R8185 gnd.n5363 gnd.n5355 163.367
R8186 gnd.n5586 gnd.n5355 163.367
R8187 gnd.n5587 gnd.n5586 163.367
R8188 gnd.n5587 gnd.n5352 163.367
R8189 gnd.n5593 gnd.n5352 163.367
R8190 gnd.n5593 gnd.n5353 163.367
R8191 gnd.n5353 gnd.n5344 163.367
R8192 gnd.n5603 gnd.n5344 163.367
R8193 gnd.n5604 gnd.n5603 163.367
R8194 gnd.n5604 gnd.n5342 163.367
R8195 gnd.n5609 gnd.n5342 163.367
R8196 gnd.n5609 gnd.n5335 163.367
R8197 gnd.n5621 gnd.n5335 163.367
R8198 gnd.n5622 gnd.n5621 163.367
R8199 gnd.n5623 gnd.n5622 163.367
R8200 gnd.n5623 gnd.n5333 163.367
R8201 gnd.n5628 gnd.n5333 163.367
R8202 gnd.n5628 gnd.n5326 163.367
R8203 gnd.n5639 gnd.n5326 163.367
R8204 gnd.n5640 gnd.n5639 163.367
R8205 gnd.n5640 gnd.n5323 163.367
R8206 gnd.n5646 gnd.n5323 163.367
R8207 gnd.n5646 gnd.n5324 163.367
R8208 gnd.n5324 gnd.n5317 163.367
R8209 gnd.n5658 gnd.n5317 163.367
R8210 gnd.n5659 gnd.n5658 163.367
R8211 gnd.n5659 gnd.n5314 163.367
R8212 gnd.n5666 gnd.n5314 163.367
R8213 gnd.n5666 gnd.n5315 163.367
R8214 gnd.n5662 gnd.n5315 163.367
R8215 gnd.n5662 gnd.n5306 163.367
R8216 gnd.n5677 gnd.n5306 163.367
R8217 gnd.n5677 gnd.n5303 163.367
R8218 gnd.n5683 gnd.n5303 163.367
R8219 gnd.n5683 gnd.n5304 163.367
R8220 gnd.n5304 gnd.n5296 163.367
R8221 gnd.n5694 gnd.n5296 163.367
R8222 gnd.n5695 gnd.n5694 163.367
R8223 gnd.n5695 gnd.n5293 163.367
R8224 gnd.n5701 gnd.n5293 163.367
R8225 gnd.n5701 gnd.n5294 163.367
R8226 gnd.n5294 gnd.n5285 163.367
R8227 gnd.n5712 gnd.n5285 163.367
R8228 gnd.n5713 gnd.n5712 163.367
R8229 gnd.n5713 gnd.n5282 163.367
R8230 gnd.n5719 gnd.n5282 163.367
R8231 gnd.n5719 gnd.n5283 163.367
R8232 gnd.n5283 gnd.n5275 163.367
R8233 gnd.n5730 gnd.n5275 163.367
R8234 gnd.n5731 gnd.n5730 163.367
R8235 gnd.n5731 gnd.n5272 163.367
R8236 gnd.n5737 gnd.n5272 163.367
R8237 gnd.n5737 gnd.n5273 163.367
R8238 gnd.n5273 gnd.n5264 163.367
R8239 gnd.n5747 gnd.n5264 163.367
R8240 gnd.n5748 gnd.n5747 163.367
R8241 gnd.n5748 gnd.n5262 163.367
R8242 gnd.n5753 gnd.n5262 163.367
R8243 gnd.n5753 gnd.n5255 163.367
R8244 gnd.n5765 gnd.n5255 163.367
R8245 gnd.n5766 gnd.n5765 163.367
R8246 gnd.n5767 gnd.n5766 163.367
R8247 gnd.n5767 gnd.n5253 163.367
R8248 gnd.n5772 gnd.n5253 163.367
R8249 gnd.n5772 gnd.n5246 163.367
R8250 gnd.n5782 gnd.n5246 163.367
R8251 gnd.n5783 gnd.n5782 163.367
R8252 gnd.n5783 gnd.n5244 163.367
R8253 gnd.n5787 gnd.n5244 163.367
R8254 gnd.n5787 gnd.n5239 163.367
R8255 gnd.n5798 gnd.n5239 163.367
R8256 gnd.n5798 gnd.n5237 163.367
R8257 gnd.n5802 gnd.n5237 163.367
R8258 gnd.n5802 gnd.n5163 163.367
R8259 gnd.n5933 gnd.n5163 163.367
R8260 gnd.n5933 gnd.n5164 163.367
R8261 gnd.n5184 gnd.n5183 156.462
R8262 gnd.n3978 gnd.n3946 153.042
R8263 gnd.n4042 gnd.n4041 152.079
R8264 gnd.n4010 gnd.n4009 152.079
R8265 gnd.n3978 gnd.n3977 152.079
R8266 gnd.n5421 gnd.n5420 152
R8267 gnd.n5422 gnd.n5411 152
R8268 gnd.n5424 gnd.n5423 152
R8269 gnd.n5426 gnd.n5409 152
R8270 gnd.n5428 gnd.n5427 152
R8271 gnd.n5182 gnd.n5166 152
R8272 gnd.n5174 gnd.n5167 152
R8273 gnd.n5173 gnd.n5172 152
R8274 gnd.n5171 gnd.n5168 152
R8275 gnd.n5169 gnd.t92 150.546
R8276 gnd.t157 gnd.n4020 147.661
R8277 gnd.t31 gnd.n3988 147.661
R8278 gnd.t155 gnd.n3956 147.661
R8279 gnd.t170 gnd.n3925 147.661
R8280 gnd.t143 gnd.n3893 147.661
R8281 gnd.t175 gnd.n3861 147.661
R8282 gnd.t173 gnd.n3829 147.661
R8283 gnd.t1 gnd.n3798 147.661
R8284 gnd.n5870 gnd.n5869 143.351
R8285 gnd.n5495 gnd.n5494 143.351
R8286 gnd.n5495 gnd.n5390 143.351
R8287 gnd.n5418 gnd.t133 130.484
R8288 gnd.n5427 gnd.t49 126.766
R8289 gnd.n5425 gnd.t118 126.766
R8290 gnd.n5411 gnd.t64 126.766
R8291 gnd.n5419 gnd.t95 126.766
R8292 gnd.n5170 gnd.t136 126.766
R8293 gnd.n5172 gnd.t115 126.766
R8294 gnd.n5181 gnd.t46 126.766
R8295 gnd.n5183 gnd.t127 126.766
R8296 gnd.n6878 gnd.n534 108.609
R8297 gnd.n5496 gnd.n1018 108.609
R8298 gnd.n4037 gnd.n4036 104.615
R8299 gnd.n4036 gnd.n4014 104.615
R8300 gnd.n4029 gnd.n4014 104.615
R8301 gnd.n4029 gnd.n4028 104.615
R8302 gnd.n4028 gnd.n4018 104.615
R8303 gnd.n4021 gnd.n4018 104.615
R8304 gnd.n4005 gnd.n4004 104.615
R8305 gnd.n4004 gnd.n3982 104.615
R8306 gnd.n3997 gnd.n3982 104.615
R8307 gnd.n3997 gnd.n3996 104.615
R8308 gnd.n3996 gnd.n3986 104.615
R8309 gnd.n3989 gnd.n3986 104.615
R8310 gnd.n3973 gnd.n3972 104.615
R8311 gnd.n3972 gnd.n3950 104.615
R8312 gnd.n3965 gnd.n3950 104.615
R8313 gnd.n3965 gnd.n3964 104.615
R8314 gnd.n3964 gnd.n3954 104.615
R8315 gnd.n3957 gnd.n3954 104.615
R8316 gnd.n3942 gnd.n3941 104.615
R8317 gnd.n3941 gnd.n3919 104.615
R8318 gnd.n3934 gnd.n3919 104.615
R8319 gnd.n3934 gnd.n3933 104.615
R8320 gnd.n3933 gnd.n3923 104.615
R8321 gnd.n3926 gnd.n3923 104.615
R8322 gnd.n3910 gnd.n3909 104.615
R8323 gnd.n3909 gnd.n3887 104.615
R8324 gnd.n3902 gnd.n3887 104.615
R8325 gnd.n3902 gnd.n3901 104.615
R8326 gnd.n3901 gnd.n3891 104.615
R8327 gnd.n3894 gnd.n3891 104.615
R8328 gnd.n3878 gnd.n3877 104.615
R8329 gnd.n3877 gnd.n3855 104.615
R8330 gnd.n3870 gnd.n3855 104.615
R8331 gnd.n3870 gnd.n3869 104.615
R8332 gnd.n3869 gnd.n3859 104.615
R8333 gnd.n3862 gnd.n3859 104.615
R8334 gnd.n3846 gnd.n3845 104.615
R8335 gnd.n3845 gnd.n3823 104.615
R8336 gnd.n3838 gnd.n3823 104.615
R8337 gnd.n3838 gnd.n3837 104.615
R8338 gnd.n3837 gnd.n3827 104.615
R8339 gnd.n3830 gnd.n3827 104.615
R8340 gnd.n3815 gnd.n3814 104.615
R8341 gnd.n3814 gnd.n3792 104.615
R8342 gnd.n3807 gnd.n3792 104.615
R8343 gnd.n3807 gnd.n3806 104.615
R8344 gnd.n3806 gnd.n3796 104.615
R8345 gnd.n3799 gnd.n3796 104.615
R8346 gnd.n3250 gnd.t41 100.632
R8347 gnd.n1439 gnd.t83 100.632
R8348 gnd.n7425 gnd.n134 99.6594
R8349 gnd.n7423 gnd.n7422 99.6594
R8350 gnd.n7418 gnd.n141 99.6594
R8351 gnd.n7416 gnd.n7415 99.6594
R8352 gnd.n7411 gnd.n148 99.6594
R8353 gnd.n7409 gnd.n7408 99.6594
R8354 gnd.n7404 gnd.n155 99.6594
R8355 gnd.n7402 gnd.n7401 99.6594
R8356 gnd.n7394 gnd.n162 99.6594
R8357 gnd.n7392 gnd.n7391 99.6594
R8358 gnd.n7387 gnd.n169 99.6594
R8359 gnd.n7385 gnd.n7384 99.6594
R8360 gnd.n7380 gnd.n176 99.6594
R8361 gnd.n7378 gnd.n7377 99.6594
R8362 gnd.n7373 gnd.n183 99.6594
R8363 gnd.n7371 gnd.n7370 99.6594
R8364 gnd.n7366 gnd.n190 99.6594
R8365 gnd.n7364 gnd.n7363 99.6594
R8366 gnd.n195 gnd.n194 99.6594
R8367 gnd.n6908 gnd.n6907 99.6594
R8368 gnd.n519 gnd.n490 99.6594
R8369 gnd.n6900 gnd.n491 99.6594
R8370 gnd.n6896 gnd.n492 99.6594
R8371 gnd.n6892 gnd.n493 99.6594
R8372 gnd.n6888 gnd.n494 99.6594
R8373 gnd.n6884 gnd.n495 99.6594
R8374 gnd.n6880 gnd.n496 99.6594
R8375 gnd.n6875 gnd.n498 99.6594
R8376 gnd.n6871 gnd.n499 99.6594
R8377 gnd.n6867 gnd.n500 99.6594
R8378 gnd.n6863 gnd.n501 99.6594
R8379 gnd.n6859 gnd.n502 99.6594
R8380 gnd.n6855 gnd.n503 99.6594
R8381 gnd.n6851 gnd.n504 99.6594
R8382 gnd.n6847 gnd.n505 99.6594
R8383 gnd.n6843 gnd.n506 99.6594
R8384 gnd.n558 gnd.n507 99.6594
R8385 gnd.n6294 gnd.n6293 99.6594
R8386 gnd.n6291 gnd.n6290 99.6594
R8387 gnd.n6286 gnd.n1001 99.6594
R8388 gnd.n6284 gnd.n6283 99.6594
R8389 gnd.n6279 gnd.n1008 99.6594
R8390 gnd.n6277 gnd.n6276 99.6594
R8391 gnd.n6272 gnd.n1015 99.6594
R8392 gnd.n6268 gnd.n6267 99.6594
R8393 gnd.n6263 gnd.n1026 99.6594
R8394 gnd.n6261 gnd.n6260 99.6594
R8395 gnd.n6256 gnd.n1033 99.6594
R8396 gnd.n6254 gnd.n6253 99.6594
R8397 gnd.n6249 gnd.n1040 99.6594
R8398 gnd.n6247 gnd.n6246 99.6594
R8399 gnd.n6242 gnd.n1047 99.6594
R8400 gnd.n6240 gnd.n6239 99.6594
R8401 gnd.n6235 gnd.n1056 99.6594
R8402 gnd.n6233 gnd.n6232 99.6594
R8403 gnd.n4474 gnd.n4285 99.6594
R8404 gnd.n4472 gnd.n4288 99.6594
R8405 gnd.n4468 gnd.n4467 99.6594
R8406 gnd.n4461 gnd.n4293 99.6594
R8407 gnd.n4460 gnd.n4459 99.6594
R8408 gnd.n4453 gnd.n4299 99.6594
R8409 gnd.n4452 gnd.n4451 99.6594
R8410 gnd.n4445 gnd.n4305 99.6594
R8411 gnd.n4444 gnd.n4443 99.6594
R8412 gnd.n4437 gnd.n4311 99.6594
R8413 gnd.n4436 gnd.n4435 99.6594
R8414 gnd.n4429 gnd.n4320 99.6594
R8415 gnd.n4428 gnd.n4427 99.6594
R8416 gnd.n4421 gnd.n4326 99.6594
R8417 gnd.n4420 gnd.n4419 99.6594
R8418 gnd.n4413 gnd.n4332 99.6594
R8419 gnd.n4412 gnd.n4411 99.6594
R8420 gnd.n4342 gnd.n4338 99.6594
R8421 gnd.n4401 gnd.n4400 99.6594
R8422 gnd.n4158 gnd.n1422 99.6594
R8423 gnd.n4156 gnd.n1421 99.6594
R8424 gnd.n4152 gnd.n1420 99.6594
R8425 gnd.n4148 gnd.n1419 99.6594
R8426 gnd.n4144 gnd.n1418 99.6594
R8427 gnd.n4140 gnd.n1417 99.6594
R8428 gnd.n4136 gnd.n1416 99.6594
R8429 gnd.n2774 gnd.n1415 99.6594
R8430 gnd.n3462 gnd.n3193 99.6594
R8431 gnd.n3219 gnd.n3200 99.6594
R8432 gnd.n3221 gnd.n3201 99.6594
R8433 gnd.n3229 gnd.n3202 99.6594
R8434 gnd.n3231 gnd.n3203 99.6594
R8435 gnd.n3239 gnd.n3204 99.6594
R8436 gnd.n3241 gnd.n3205 99.6594
R8437 gnd.n3249 gnd.n3206 99.6594
R8438 gnd.n4126 gnd.n1402 99.6594
R8439 gnd.n4122 gnd.n1403 99.6594
R8440 gnd.n4118 gnd.n1404 99.6594
R8441 gnd.n4114 gnd.n1405 99.6594
R8442 gnd.n4110 gnd.n1406 99.6594
R8443 gnd.n4106 gnd.n1407 99.6594
R8444 gnd.n4102 gnd.n1408 99.6594
R8445 gnd.n4098 gnd.n1409 99.6594
R8446 gnd.n4094 gnd.n1410 99.6594
R8447 gnd.n4090 gnd.n1411 99.6594
R8448 gnd.n4086 gnd.n1412 99.6594
R8449 gnd.n4082 gnd.n1413 99.6594
R8450 gnd.n4078 gnd.n1414 99.6594
R8451 gnd.n3377 gnd.n3376 99.6594
R8452 gnd.n3371 gnd.n3288 99.6594
R8453 gnd.n3368 gnd.n3289 99.6594
R8454 gnd.n3364 gnd.n3290 99.6594
R8455 gnd.n3360 gnd.n3291 99.6594
R8456 gnd.n3356 gnd.n3292 99.6594
R8457 gnd.n3352 gnd.n3293 99.6594
R8458 gnd.n3348 gnd.n3294 99.6594
R8459 gnd.n3344 gnd.n3295 99.6594
R8460 gnd.n3340 gnd.n3296 99.6594
R8461 gnd.n3336 gnd.n3297 99.6594
R8462 gnd.n3332 gnd.n3298 99.6594
R8463 gnd.n3379 gnd.n3287 99.6594
R8464 gnd.n7280 gnd.n7279 99.6594
R8465 gnd.n7285 gnd.n7284 99.6594
R8466 gnd.n7288 gnd.n7287 99.6594
R8467 gnd.n7293 gnd.n7292 99.6594
R8468 gnd.n7296 gnd.n7295 99.6594
R8469 gnd.n7301 gnd.n7300 99.6594
R8470 gnd.n7304 gnd.n7303 99.6594
R8471 gnd.n7309 gnd.n7307 99.6594
R8472 gnd.n7435 gnd.n121 99.6594
R8473 gnd.n5956 gnd.n508 99.6594
R8474 gnd.n5960 gnd.n509 99.6594
R8475 gnd.n5962 gnd.n510 99.6594
R8476 gnd.n5972 gnd.n511 99.6594
R8477 gnd.n5980 gnd.n512 99.6594
R8478 gnd.n5982 gnd.n513 99.6594
R8479 gnd.n5992 gnd.n514 99.6594
R8480 gnd.n6000 gnd.n515 99.6594
R8481 gnd.n6002 gnd.n516 99.6594
R8482 gnd.n5002 gnd.n5001 99.6594
R8483 gnd.n5005 gnd.n5004 99.6594
R8484 gnd.n5014 gnd.n5013 99.6594
R8485 gnd.n5025 gnd.n5024 99.6594
R8486 gnd.n5028 gnd.n5027 99.6594
R8487 gnd.n5037 gnd.n5036 99.6594
R8488 gnd.n5048 gnd.n5047 99.6594
R8489 gnd.n5052 gnd.n5050 99.6594
R8490 gnd.n6304 gnd.n979 99.6594
R8491 gnd.n4193 gnd.n1399 99.6594
R8492 gnd.n4196 gnd.n4195 99.6594
R8493 gnd.n4203 gnd.n4202 99.6594
R8494 gnd.n4206 gnd.n4205 99.6594
R8495 gnd.n4213 gnd.n4212 99.6594
R8496 gnd.n4216 gnd.n4215 99.6594
R8497 gnd.n4223 gnd.n4222 99.6594
R8498 gnd.n4226 gnd.n4225 99.6594
R8499 gnd.n4233 gnd.n4232 99.6594
R8500 gnd.n4194 gnd.n4193 99.6594
R8501 gnd.n4195 gnd.n4188 99.6594
R8502 gnd.n4204 gnd.n4203 99.6594
R8503 gnd.n4205 gnd.n4184 99.6594
R8504 gnd.n4214 gnd.n4213 99.6594
R8505 gnd.n4215 gnd.n4180 99.6594
R8506 gnd.n4224 gnd.n4223 99.6594
R8507 gnd.n4225 gnd.n4176 99.6594
R8508 gnd.n4234 gnd.n4233 99.6594
R8509 gnd.n5051 gnd.n979 99.6594
R8510 gnd.n5050 gnd.n5049 99.6594
R8511 gnd.n5047 gnd.n5038 99.6594
R8512 gnd.n5036 gnd.n5035 99.6594
R8513 gnd.n5027 gnd.n5026 99.6594
R8514 gnd.n5024 gnd.n5015 99.6594
R8515 gnd.n5013 gnd.n5012 99.6594
R8516 gnd.n5004 gnd.n5003 99.6594
R8517 gnd.n5001 gnd.n5000 99.6594
R8518 gnd.n5959 gnd.n508 99.6594
R8519 gnd.n5961 gnd.n509 99.6594
R8520 gnd.n5971 gnd.n510 99.6594
R8521 gnd.n5979 gnd.n511 99.6594
R8522 gnd.n5981 gnd.n512 99.6594
R8523 gnd.n5991 gnd.n513 99.6594
R8524 gnd.n5999 gnd.n514 99.6594
R8525 gnd.n6001 gnd.n515 99.6594
R8526 gnd.n6046 gnd.n516 99.6594
R8527 gnd.n7308 gnd.n121 99.6594
R8528 gnd.n7307 gnd.n7306 99.6594
R8529 gnd.n7303 gnd.n7302 99.6594
R8530 gnd.n7300 gnd.n7299 99.6594
R8531 gnd.n7295 gnd.n7294 99.6594
R8532 gnd.n7292 gnd.n7291 99.6594
R8533 gnd.n7287 gnd.n7286 99.6594
R8534 gnd.n7284 gnd.n7283 99.6594
R8535 gnd.n7279 gnd.n7278 99.6594
R8536 gnd.n3377 gnd.n3300 99.6594
R8537 gnd.n3369 gnd.n3288 99.6594
R8538 gnd.n3365 gnd.n3289 99.6594
R8539 gnd.n3361 gnd.n3290 99.6594
R8540 gnd.n3357 gnd.n3291 99.6594
R8541 gnd.n3353 gnd.n3292 99.6594
R8542 gnd.n3349 gnd.n3293 99.6594
R8543 gnd.n3345 gnd.n3294 99.6594
R8544 gnd.n3341 gnd.n3295 99.6594
R8545 gnd.n3337 gnd.n3296 99.6594
R8546 gnd.n3333 gnd.n3297 99.6594
R8547 gnd.n3329 gnd.n3298 99.6594
R8548 gnd.n3380 gnd.n3379 99.6594
R8549 gnd.n4081 gnd.n1414 99.6594
R8550 gnd.n4085 gnd.n1413 99.6594
R8551 gnd.n4089 gnd.n1412 99.6594
R8552 gnd.n4093 gnd.n1411 99.6594
R8553 gnd.n4097 gnd.n1410 99.6594
R8554 gnd.n4101 gnd.n1409 99.6594
R8555 gnd.n4105 gnd.n1408 99.6594
R8556 gnd.n4109 gnd.n1407 99.6594
R8557 gnd.n4113 gnd.n1406 99.6594
R8558 gnd.n4117 gnd.n1405 99.6594
R8559 gnd.n4121 gnd.n1404 99.6594
R8560 gnd.n4125 gnd.n1403 99.6594
R8561 gnd.n1443 gnd.n1402 99.6594
R8562 gnd.n3463 gnd.n3462 99.6594
R8563 gnd.n3222 gnd.n3200 99.6594
R8564 gnd.n3228 gnd.n3201 99.6594
R8565 gnd.n3232 gnd.n3202 99.6594
R8566 gnd.n3238 gnd.n3203 99.6594
R8567 gnd.n3242 gnd.n3204 99.6594
R8568 gnd.n3248 gnd.n3205 99.6594
R8569 gnd.n3206 gnd.n3190 99.6594
R8570 gnd.n4135 gnd.n1415 99.6594
R8571 gnd.n4139 gnd.n1416 99.6594
R8572 gnd.n4143 gnd.n1417 99.6594
R8573 gnd.n4147 gnd.n1418 99.6594
R8574 gnd.n4151 gnd.n1419 99.6594
R8575 gnd.n4155 gnd.n1420 99.6594
R8576 gnd.n4159 gnd.n1421 99.6594
R8577 gnd.n1424 gnd.n1422 99.6594
R8578 gnd.n4475 gnd.n4474 99.6594
R8579 gnd.n4469 gnd.n4288 99.6594
R8580 gnd.n4467 gnd.n4466 99.6594
R8581 gnd.n4462 gnd.n4461 99.6594
R8582 gnd.n4459 gnd.n4458 99.6594
R8583 gnd.n4454 gnd.n4453 99.6594
R8584 gnd.n4451 gnd.n4450 99.6594
R8585 gnd.n4446 gnd.n4445 99.6594
R8586 gnd.n4443 gnd.n4442 99.6594
R8587 gnd.n4438 gnd.n4437 99.6594
R8588 gnd.n4435 gnd.n4434 99.6594
R8589 gnd.n4430 gnd.n4429 99.6594
R8590 gnd.n4427 gnd.n4426 99.6594
R8591 gnd.n4422 gnd.n4421 99.6594
R8592 gnd.n4419 gnd.n4418 99.6594
R8593 gnd.n4414 gnd.n4413 99.6594
R8594 gnd.n4411 gnd.n4410 99.6594
R8595 gnd.n4343 gnd.n4342 99.6594
R8596 gnd.n4402 gnd.n4401 99.6594
R8597 gnd.n6234 gnd.n6233 99.6594
R8598 gnd.n1056 gnd.n1048 99.6594
R8599 gnd.n6241 gnd.n6240 99.6594
R8600 gnd.n1047 gnd.n1041 99.6594
R8601 gnd.n6248 gnd.n6247 99.6594
R8602 gnd.n1040 gnd.n1034 99.6594
R8603 gnd.n6255 gnd.n6254 99.6594
R8604 gnd.n1033 gnd.n1027 99.6594
R8605 gnd.n6262 gnd.n6261 99.6594
R8606 gnd.n1026 gnd.n1019 99.6594
R8607 gnd.n6271 gnd.n6270 99.6594
R8608 gnd.n1015 gnd.n1009 99.6594
R8609 gnd.n6278 gnd.n6277 99.6594
R8610 gnd.n1008 gnd.n1002 99.6594
R8611 gnd.n6285 gnd.n6284 99.6594
R8612 gnd.n1001 gnd.n994 99.6594
R8613 gnd.n6292 gnd.n6291 99.6594
R8614 gnd.n6295 gnd.n6294 99.6594
R8615 gnd.n6907 gnd.n488 99.6594
R8616 gnd.n6901 gnd.n490 99.6594
R8617 gnd.n6897 gnd.n491 99.6594
R8618 gnd.n6893 gnd.n492 99.6594
R8619 gnd.n6889 gnd.n493 99.6594
R8620 gnd.n6885 gnd.n494 99.6594
R8621 gnd.n6881 gnd.n495 99.6594
R8622 gnd.n6876 gnd.n497 99.6594
R8623 gnd.n6872 gnd.n498 99.6594
R8624 gnd.n6868 gnd.n499 99.6594
R8625 gnd.n6864 gnd.n500 99.6594
R8626 gnd.n6860 gnd.n501 99.6594
R8627 gnd.n6856 gnd.n502 99.6594
R8628 gnd.n6852 gnd.n503 99.6594
R8629 gnd.n6848 gnd.n504 99.6594
R8630 gnd.n6844 gnd.n505 99.6594
R8631 gnd.n557 gnd.n506 99.6594
R8632 gnd.n6836 gnd.n507 99.6594
R8633 gnd.n194 gnd.n191 99.6594
R8634 gnd.n7365 gnd.n7364 99.6594
R8635 gnd.n190 gnd.n184 99.6594
R8636 gnd.n7372 gnd.n7371 99.6594
R8637 gnd.n183 gnd.n177 99.6594
R8638 gnd.n7379 gnd.n7378 99.6594
R8639 gnd.n176 gnd.n170 99.6594
R8640 gnd.n7386 gnd.n7385 99.6594
R8641 gnd.n169 gnd.n163 99.6594
R8642 gnd.n7393 gnd.n7392 99.6594
R8643 gnd.n162 gnd.n156 99.6594
R8644 gnd.n7403 gnd.n7402 99.6594
R8645 gnd.n155 gnd.n149 99.6594
R8646 gnd.n7410 gnd.n7409 99.6594
R8647 gnd.n148 gnd.n142 99.6594
R8648 gnd.n7417 gnd.n7416 99.6594
R8649 gnd.n141 gnd.n135 99.6594
R8650 gnd.n7424 gnd.n7423 99.6594
R8651 gnd.n134 gnd.n131 99.6594
R8652 gnd.n5093 gnd.n944 99.6594
R8653 gnd.n4993 gnd.n945 99.6594
R8654 gnd.n5009 gnd.n946 99.6594
R8655 gnd.n5019 gnd.n947 99.6594
R8656 gnd.n5021 gnd.n948 99.6594
R8657 gnd.n5032 gnd.n949 99.6594
R8658 gnd.n5042 gnd.n950 99.6594
R8659 gnd.n5044 gnd.n951 99.6594
R8660 gnd.n974 gnd.n952 99.6594
R8661 gnd.n6311 gnd.n953 99.6594
R8662 gnd.n969 gnd.n954 99.6594
R8663 gnd.n6320 gnd.n955 99.6594
R8664 gnd.n965 gnd.n956 99.6594
R8665 gnd.n6329 gnd.n957 99.6594
R8666 gnd.n4992 gnd.n944 99.6594
R8667 gnd.n5008 gnd.n945 99.6594
R8668 gnd.n5018 gnd.n946 99.6594
R8669 gnd.n5020 gnd.n947 99.6594
R8670 gnd.n5031 gnd.n948 99.6594
R8671 gnd.n5041 gnd.n949 99.6594
R8672 gnd.n5043 gnd.n950 99.6594
R8673 gnd.n973 gnd.n951 99.6594
R8674 gnd.n6310 gnd.n952 99.6594
R8675 gnd.n968 gnd.n953 99.6594
R8676 gnd.n6319 gnd.n954 99.6594
R8677 gnd.n964 gnd.n955 99.6594
R8678 gnd.n6328 gnd.n956 99.6594
R8679 gnd.n958 gnd.n957 99.6594
R8680 gnd.n6093 gnd.n617 99.6594
R8681 gnd.n5966 gnd.n618 99.6594
R8682 gnd.n5968 gnd.n619 99.6594
R8683 gnd.n5976 gnd.n620 99.6594
R8684 gnd.n5986 gnd.n621 99.6594
R8685 gnd.n5988 gnd.n622 99.6594
R8686 gnd.n5996 gnd.n623 99.6594
R8687 gnd.n6006 gnd.n624 99.6594
R8688 gnd.n6008 gnd.n625 99.6594
R8689 gnd.n6013 gnd.n626 99.6594
R8690 gnd.n6015 gnd.n627 99.6594
R8691 gnd.n6019 gnd.n628 99.6594
R8692 gnd.n6021 gnd.n629 99.6594
R8693 gnd.n6028 gnd.n630 99.6594
R8694 gnd.n631 gnd.n630 99.6594
R8695 gnd.n6027 gnd.n629 99.6594
R8696 gnd.n6020 gnd.n628 99.6594
R8697 gnd.n6018 gnd.n627 99.6594
R8698 gnd.n6014 gnd.n626 99.6594
R8699 gnd.n6012 gnd.n625 99.6594
R8700 gnd.n6007 gnd.n624 99.6594
R8701 gnd.n6005 gnd.n623 99.6594
R8702 gnd.n5995 gnd.n622 99.6594
R8703 gnd.n5987 gnd.n621 99.6594
R8704 gnd.n5985 gnd.n620 99.6594
R8705 gnd.n5975 gnd.n619 99.6594
R8706 gnd.n5967 gnd.n618 99.6594
R8707 gnd.n5965 gnd.n617 99.6594
R8708 gnd.n961 gnd.t114 98.63
R8709 gnd.n118 gnd.t54 98.63
R8710 gnd.n6047 gnd.t87 98.63
R8711 gnd.n976 gnd.t102 98.63
R8712 gnd.n537 gnd.t80 98.63
R8713 gnd.n559 gnd.t59 98.63
R8714 gnd.n197 gnd.t131 98.63
R8715 gnd.n7396 gnd.t140 98.63
R8716 gnd.n4312 gnd.t77 98.63
R8717 gnd.n4344 gnd.t45 98.63
R8718 gnd.n4173 gnd.t110 98.63
R8719 gnd.n1053 gnd.t73 98.63
R8720 gnd.n1016 gnd.t99 98.63
R8721 gnd.n6024 gnd.t90 98.63
R8722 gnd.n5385 gnd.t123 96.6984
R8723 gnd.n5212 gnd.t69 96.6984
R8724 gnd.n5393 gnd.t37 96.6906
R8725 gnd.n5206 gnd.t125 96.6906
R8726 gnd.n2240 gnd.n2239 89.3769
R8727 gnd.n2239 gnd.n1909 89.3769
R8728 gnd.n2231 gnd.n1909 89.3769
R8729 gnd.n2231 gnd.n2230 89.3769
R8730 gnd.n2230 gnd.n2229 89.3769
R8731 gnd.n2229 gnd.n1917 89.3769
R8732 gnd.n2223 gnd.n1917 89.3769
R8733 gnd.n2223 gnd.n2222 89.3769
R8734 gnd.n2222 gnd.n2221 89.3769
R8735 gnd.n2221 gnd.n1924 89.3769
R8736 gnd.n2215 gnd.n1924 89.3769
R8737 gnd.n2215 gnd.n2214 89.3769
R8738 gnd.n2214 gnd.n2213 89.3769
R8739 gnd.n2213 gnd.n1932 89.3769
R8740 gnd.n2207 gnd.n1932 89.3769
R8741 gnd.n2207 gnd.n2206 89.3769
R8742 gnd.n2206 gnd.n2205 89.3769
R8743 gnd.n2205 gnd.n1940 89.3769
R8744 gnd.n2199 gnd.n1940 89.3769
R8745 gnd.n2199 gnd.n2198 89.3769
R8746 gnd.n2198 gnd.n2197 89.3769
R8747 gnd.n2197 gnd.n1948 89.3769
R8748 gnd.n2191 gnd.n1948 89.3769
R8749 gnd.n2191 gnd.n2190 89.3769
R8750 gnd.n2190 gnd.n2189 89.3769
R8751 gnd.n2189 gnd.n1956 89.3769
R8752 gnd.n2183 gnd.n1956 89.3769
R8753 gnd.n2183 gnd.n2182 89.3769
R8754 gnd.n2182 gnd.n2181 89.3769
R8755 gnd.n2181 gnd.n1964 89.3769
R8756 gnd.n2175 gnd.n1964 89.3769
R8757 gnd.n2175 gnd.n2174 89.3769
R8758 gnd.n2174 gnd.n2173 89.3769
R8759 gnd.n2173 gnd.n1972 89.3769
R8760 gnd.n2167 gnd.n1972 89.3769
R8761 gnd.n2167 gnd.n2166 89.3769
R8762 gnd.n2166 gnd.n2165 89.3769
R8763 gnd.n2165 gnd.n1980 89.3769
R8764 gnd.n2159 gnd.n1980 89.3769
R8765 gnd.n2159 gnd.n2158 89.3769
R8766 gnd.n2158 gnd.n2157 89.3769
R8767 gnd.n2157 gnd.n1988 89.3769
R8768 gnd.n2151 gnd.n1988 89.3769
R8769 gnd.n2151 gnd.n2150 89.3769
R8770 gnd.n2150 gnd.n2149 89.3769
R8771 gnd.n2149 gnd.n1996 89.3769
R8772 gnd.n2143 gnd.n1996 89.3769
R8773 gnd.n2143 gnd.n2142 89.3769
R8774 gnd.n2142 gnd.n2141 89.3769
R8775 gnd.n2141 gnd.n2004 89.3769
R8776 gnd.n2135 gnd.n2004 89.3769
R8777 gnd.n2135 gnd.n2134 89.3769
R8778 gnd.n2134 gnd.n2133 89.3769
R8779 gnd.n2133 gnd.n2012 89.3769
R8780 gnd.n2127 gnd.n2012 89.3769
R8781 gnd.n2127 gnd.n2126 89.3769
R8782 gnd.n2126 gnd.n2125 89.3769
R8783 gnd.n2125 gnd.n2020 89.3769
R8784 gnd.n2119 gnd.n2020 89.3769
R8785 gnd.n2119 gnd.n2118 89.3769
R8786 gnd.n2118 gnd.n2117 89.3769
R8787 gnd.n2117 gnd.n2028 89.3769
R8788 gnd.n2111 gnd.n2028 89.3769
R8789 gnd.n2111 gnd.n2110 89.3769
R8790 gnd.n2110 gnd.n2109 89.3769
R8791 gnd.n2109 gnd.n2036 89.3769
R8792 gnd.n2103 gnd.n2036 89.3769
R8793 gnd.n2103 gnd.n2102 89.3769
R8794 gnd.n2102 gnd.n2101 89.3769
R8795 gnd.n2101 gnd.n2044 89.3769
R8796 gnd.n2095 gnd.n2044 89.3769
R8797 gnd.n2095 gnd.n2094 89.3769
R8798 gnd.n2094 gnd.n2093 89.3769
R8799 gnd.n2093 gnd.n2052 89.3769
R8800 gnd.n2087 gnd.n2052 89.3769
R8801 gnd.n2087 gnd.n2086 89.3769
R8802 gnd.n2086 gnd.n2085 89.3769
R8803 gnd.n2085 gnd.n2060 89.3769
R8804 gnd.n2079 gnd.n2060 89.3769
R8805 gnd.n2079 gnd.n2078 89.3769
R8806 gnd.n2078 gnd.n2077 89.3769
R8807 gnd.n2077 gnd.n2069 89.3769
R8808 gnd.n2069 gnd.n2068 89.3769
R8809 gnd.n5418 gnd.n5417 81.8399
R8810 gnd.n3251 gnd.t40 74.8376
R8811 gnd.n1440 gnd.t84 74.8376
R8812 gnd.n5386 gnd.t122 72.8438
R8813 gnd.n5213 gnd.t70 72.8438
R8814 gnd.n5419 gnd.n5412 72.8411
R8815 gnd.n5425 gnd.n5410 72.8411
R8816 gnd.n5181 gnd.n5180 72.8411
R8817 gnd.n962 gnd.t113 72.836
R8818 gnd.n5394 gnd.t36 72.836
R8819 gnd.n5207 gnd.t126 72.836
R8820 gnd.n119 gnd.t55 72.836
R8821 gnd.n6048 gnd.t86 72.836
R8822 gnd.n977 gnd.t103 72.836
R8823 gnd.n538 gnd.t79 72.836
R8824 gnd.n560 gnd.t58 72.836
R8825 gnd.n198 gnd.t132 72.836
R8826 gnd.n7397 gnd.t141 72.836
R8827 gnd.n4313 gnd.t76 72.836
R8828 gnd.n4345 gnd.t44 72.836
R8829 gnd.n4174 gnd.t109 72.836
R8830 gnd.n1054 gnd.t74 72.836
R8831 gnd.n1017 gnd.t100 72.836
R8832 gnd.n6025 gnd.t91 72.836
R8833 gnd.n5927 gnd.n5926 71.676
R8834 gnd.n5924 gnd.n5923 71.676
R8835 gnd.n5919 gnd.n5189 71.676
R8836 gnd.n5917 gnd.n5916 71.676
R8837 gnd.n5912 gnd.n5192 71.676
R8838 gnd.n5910 gnd.n5909 71.676
R8839 gnd.n5905 gnd.n5195 71.676
R8840 gnd.n5903 gnd.n5902 71.676
R8841 gnd.n5898 gnd.n5198 71.676
R8842 gnd.n5896 gnd.n5895 71.676
R8843 gnd.n5891 gnd.n5201 71.676
R8844 gnd.n5889 gnd.n5888 71.676
R8845 gnd.n5884 gnd.n5204 71.676
R8846 gnd.n5882 gnd.n5881 71.676
R8847 gnd.n5876 gnd.n5209 71.676
R8848 gnd.n5874 gnd.n5873 71.676
R8849 gnd.n5869 gnd.n5868 71.676
R8850 gnd.n5866 gnd.n5865 71.676
R8851 gnd.n5860 gnd.n5215 71.676
R8852 gnd.n5858 gnd.n5857 71.676
R8853 gnd.n5853 gnd.n5218 71.676
R8854 gnd.n5851 gnd.n5850 71.676
R8855 gnd.n5846 gnd.n5221 71.676
R8856 gnd.n5844 gnd.n5843 71.676
R8857 gnd.n5839 gnd.n5224 71.676
R8858 gnd.n5837 gnd.n5836 71.676
R8859 gnd.n5832 gnd.n5227 71.676
R8860 gnd.n5830 gnd.n5829 71.676
R8861 gnd.n5825 gnd.n5230 71.676
R8862 gnd.n5823 gnd.n5822 71.676
R8863 gnd.n5818 gnd.n5233 71.676
R8864 gnd.n5816 gnd.n5815 71.676
R8865 gnd.n5811 gnd.n5809 71.676
R8866 gnd.n5433 gnd.n5432 71.676
R8867 gnd.n5437 gnd.n5436 71.676
R8868 gnd.n5442 gnd.n5441 71.676
R8869 gnd.n5445 gnd.n5444 71.676
R8870 gnd.n5450 gnd.n5449 71.676
R8871 gnd.n5453 gnd.n5452 71.676
R8872 gnd.n5458 gnd.n5457 71.676
R8873 gnd.n5461 gnd.n5460 71.676
R8874 gnd.n5466 gnd.n5465 71.676
R8875 gnd.n5469 gnd.n5468 71.676
R8876 gnd.n5474 gnd.n5473 71.676
R8877 gnd.n5477 gnd.n5476 71.676
R8878 gnd.n5482 gnd.n5481 71.676
R8879 gnd.n5485 gnd.n5484 71.676
R8880 gnd.n5491 gnd.n5490 71.676
R8881 gnd.n5494 gnd.n5493 71.676
R8882 gnd.n5499 gnd.n5498 71.676
R8883 gnd.n5502 gnd.n5501 71.676
R8884 gnd.n5508 gnd.n5507 71.676
R8885 gnd.n5511 gnd.n5510 71.676
R8886 gnd.n5516 gnd.n5515 71.676
R8887 gnd.n5519 gnd.n5518 71.676
R8888 gnd.n5524 gnd.n5523 71.676
R8889 gnd.n5527 gnd.n5526 71.676
R8890 gnd.n5532 gnd.n5531 71.676
R8891 gnd.n5535 gnd.n5534 71.676
R8892 gnd.n5540 gnd.n5539 71.676
R8893 gnd.n5543 gnd.n5542 71.676
R8894 gnd.n5548 gnd.n5547 71.676
R8895 gnd.n5551 gnd.n5550 71.676
R8896 gnd.n5556 gnd.n5555 71.676
R8897 gnd.n5559 gnd.n5558 71.676
R8898 gnd.n5434 gnd.n5433 71.676
R8899 gnd.n5436 gnd.n5406 71.676
R8900 gnd.n5443 gnd.n5442 71.676
R8901 gnd.n5444 gnd.n5404 71.676
R8902 gnd.n5451 gnd.n5450 71.676
R8903 gnd.n5452 gnd.n5402 71.676
R8904 gnd.n5459 gnd.n5458 71.676
R8905 gnd.n5460 gnd.n5400 71.676
R8906 gnd.n5467 gnd.n5466 71.676
R8907 gnd.n5468 gnd.n5398 71.676
R8908 gnd.n5475 gnd.n5474 71.676
R8909 gnd.n5476 gnd.n5396 71.676
R8910 gnd.n5483 gnd.n5482 71.676
R8911 gnd.n5484 gnd.n5392 71.676
R8912 gnd.n5492 gnd.n5491 71.676
R8913 gnd.n5390 gnd.n5388 71.676
R8914 gnd.n5500 gnd.n5499 71.676
R8915 gnd.n5501 gnd.n5384 71.676
R8916 gnd.n5509 gnd.n5508 71.676
R8917 gnd.n5510 gnd.n5382 71.676
R8918 gnd.n5517 gnd.n5516 71.676
R8919 gnd.n5518 gnd.n5380 71.676
R8920 gnd.n5525 gnd.n5524 71.676
R8921 gnd.n5526 gnd.n5378 71.676
R8922 gnd.n5533 gnd.n5532 71.676
R8923 gnd.n5534 gnd.n5376 71.676
R8924 gnd.n5541 gnd.n5540 71.676
R8925 gnd.n5542 gnd.n5374 71.676
R8926 gnd.n5549 gnd.n5548 71.676
R8927 gnd.n5550 gnd.n5372 71.676
R8928 gnd.n5557 gnd.n5556 71.676
R8929 gnd.n5560 gnd.n5559 71.676
R8930 gnd.n5809 gnd.n5234 71.676
R8931 gnd.n5817 gnd.n5816 71.676
R8932 gnd.n5233 gnd.n5231 71.676
R8933 gnd.n5824 gnd.n5823 71.676
R8934 gnd.n5230 gnd.n5228 71.676
R8935 gnd.n5831 gnd.n5830 71.676
R8936 gnd.n5227 gnd.n5225 71.676
R8937 gnd.n5838 gnd.n5837 71.676
R8938 gnd.n5224 gnd.n5222 71.676
R8939 gnd.n5845 gnd.n5844 71.676
R8940 gnd.n5221 gnd.n5219 71.676
R8941 gnd.n5852 gnd.n5851 71.676
R8942 gnd.n5218 gnd.n5216 71.676
R8943 gnd.n5859 gnd.n5858 71.676
R8944 gnd.n5215 gnd.n5211 71.676
R8945 gnd.n5867 gnd.n5866 71.676
R8946 gnd.n5871 gnd.n5870 71.676
R8947 gnd.n5875 gnd.n5874 71.676
R8948 gnd.n5209 gnd.n5205 71.676
R8949 gnd.n5883 gnd.n5882 71.676
R8950 gnd.n5204 gnd.n5202 71.676
R8951 gnd.n5890 gnd.n5889 71.676
R8952 gnd.n5201 gnd.n5199 71.676
R8953 gnd.n5897 gnd.n5896 71.676
R8954 gnd.n5198 gnd.n5196 71.676
R8955 gnd.n5904 gnd.n5903 71.676
R8956 gnd.n5195 gnd.n5193 71.676
R8957 gnd.n5911 gnd.n5910 71.676
R8958 gnd.n5192 gnd.n5190 71.676
R8959 gnd.n5918 gnd.n5917 71.676
R8960 gnd.n5189 gnd.n5187 71.676
R8961 gnd.n5925 gnd.n5924 71.676
R8962 gnd.n5928 gnd.n5927 71.676
R8963 gnd.n8 gnd.t33 69.1507
R8964 gnd.n14 gnd.t341 68.4792
R8965 gnd.n13 gnd.t5 68.4792
R8966 gnd.n12 gnd.t149 68.4792
R8967 gnd.n11 gnd.t161 68.4792
R8968 gnd.n10 gnd.t164 68.4792
R8969 gnd.n9 gnd.t159 68.4792
R8970 gnd.n8 gnd.t3 68.4792
R8971 gnd.n3378 gnd.n3282 64.369
R8972 gnd.n5504 gnd.n5386 59.5399
R8973 gnd.n5862 gnd.n5213 59.5399
R8974 gnd.n5488 gnd.n5394 59.5399
R8975 gnd.n5878 gnd.n5207 59.5399
R8976 gnd.n5430 gnd.n5428 59.1804
R8977 gnd.n4167 gnd.n1400 57.3586
R8978 gnd.n3069 gnd.t185 56.607
R8979 gnd.n56 gnd.t311 56.607
R8980 gnd.n3030 gnd.t265 56.407
R8981 gnd.n3049 gnd.t238 56.407
R8982 gnd.n17 gnd.t304 56.407
R8983 gnd.n36 gnd.t275 56.407
R8984 gnd.n3086 gnd.t247 55.8337
R8985 gnd.n3047 gnd.t289 55.8337
R8986 gnd.n3066 gnd.t262 55.8337
R8987 gnd.n73 gnd.t321 55.8337
R8988 gnd.n34 gnd.t302 55.8337
R8989 gnd.n53 gnd.t272 55.8337
R8990 gnd.n5416 gnd.n5415 54.358
R8991 gnd.n5178 gnd.n5177 54.358
R8992 gnd.n2068 gnd.n236 53.6263
R8993 gnd.n3069 gnd.n3068 53.0052
R8994 gnd.n3071 gnd.n3070 53.0052
R8995 gnd.n3073 gnd.n3072 53.0052
R8996 gnd.n3075 gnd.n3074 53.0052
R8997 gnd.n3077 gnd.n3076 53.0052
R8998 gnd.n3079 gnd.n3078 53.0052
R8999 gnd.n3081 gnd.n3080 53.0052
R9000 gnd.n3083 gnd.n3082 53.0052
R9001 gnd.n3085 gnd.n3084 53.0052
R9002 gnd.n3030 gnd.n3029 53.0052
R9003 gnd.n3032 gnd.n3031 53.0052
R9004 gnd.n3034 gnd.n3033 53.0052
R9005 gnd.n3036 gnd.n3035 53.0052
R9006 gnd.n3038 gnd.n3037 53.0052
R9007 gnd.n3040 gnd.n3039 53.0052
R9008 gnd.n3042 gnd.n3041 53.0052
R9009 gnd.n3044 gnd.n3043 53.0052
R9010 gnd.n3046 gnd.n3045 53.0052
R9011 gnd.n3049 gnd.n3048 53.0052
R9012 gnd.n3051 gnd.n3050 53.0052
R9013 gnd.n3053 gnd.n3052 53.0052
R9014 gnd.n3055 gnd.n3054 53.0052
R9015 gnd.n3057 gnd.n3056 53.0052
R9016 gnd.n3059 gnd.n3058 53.0052
R9017 gnd.n3061 gnd.n3060 53.0052
R9018 gnd.n3063 gnd.n3062 53.0052
R9019 gnd.n3065 gnd.n3064 53.0052
R9020 gnd.n72 gnd.n71 53.0052
R9021 gnd.n70 gnd.n69 53.0052
R9022 gnd.n68 gnd.n67 53.0052
R9023 gnd.n66 gnd.n65 53.0052
R9024 gnd.n64 gnd.n63 53.0052
R9025 gnd.n62 gnd.n61 53.0052
R9026 gnd.n60 gnd.n59 53.0052
R9027 gnd.n58 gnd.n57 53.0052
R9028 gnd.n56 gnd.n55 53.0052
R9029 gnd.n33 gnd.n32 53.0052
R9030 gnd.n31 gnd.n30 53.0052
R9031 gnd.n29 gnd.n28 53.0052
R9032 gnd.n27 gnd.n26 53.0052
R9033 gnd.n25 gnd.n24 53.0052
R9034 gnd.n23 gnd.n22 53.0052
R9035 gnd.n21 gnd.n20 53.0052
R9036 gnd.n19 gnd.n18 53.0052
R9037 gnd.n17 gnd.n16 53.0052
R9038 gnd.n52 gnd.n51 53.0052
R9039 gnd.n50 gnd.n49 53.0052
R9040 gnd.n48 gnd.n47 53.0052
R9041 gnd.n46 gnd.n45 53.0052
R9042 gnd.n44 gnd.n43 53.0052
R9043 gnd.n42 gnd.n41 53.0052
R9044 gnd.n40 gnd.n39 53.0052
R9045 gnd.n38 gnd.n37 53.0052
R9046 gnd.n36 gnd.n35 53.0052
R9047 gnd.n5169 gnd.n5168 52.4801
R9048 gnd.n4021 gnd.t157 52.3082
R9049 gnd.n3989 gnd.t31 52.3082
R9050 gnd.n3957 gnd.t155 52.3082
R9051 gnd.n3926 gnd.t170 52.3082
R9052 gnd.n3894 gnd.t143 52.3082
R9053 gnd.n3862 gnd.t175 52.3082
R9054 gnd.n3830 gnd.t173 52.3082
R9055 gnd.n3799 gnd.t1 52.3082
R9056 gnd.n4482 gnd.n4168 51.6227
R9057 gnd.n7433 gnd.n124 51.6227
R9058 gnd.n3851 gnd.n3819 51.4173
R9059 gnd.n3915 gnd.n3914 50.455
R9060 gnd.n3883 gnd.n3882 50.455
R9061 gnd.n3851 gnd.n3850 50.455
R9062 gnd.n3325 gnd.n3324 45.1884
R9063 gnd.n1466 gnd.n1465 45.1884
R9064 gnd.n5930 gnd.n5184 44.3322
R9065 gnd.n5419 gnd.n5418 44.3189
R9066 gnd.n6326 gnd.n962 42.2793
R9067 gnd.n3326 gnd.n3325 42.2793
R9068 gnd.n1467 gnd.n1466 42.2793
R9069 gnd.n3252 gnd.n3251 42.2793
R9070 gnd.n4134 gnd.n1440 42.2793
R9071 gnd.n120 gnd.n119 42.2793
R9072 gnd.n6049 gnd.n6048 42.2793
R9073 gnd.n978 gnd.n977 42.2793
R9074 gnd.n561 gnd.n560 42.2793
R9075 gnd.n7361 gnd.n198 42.2793
R9076 gnd.n7398 gnd.n7397 42.2793
R9077 gnd.n4314 gnd.n4313 42.2793
R9078 gnd.n4346 gnd.n4345 42.2793
R9079 gnd.n4175 gnd.n4174 42.2793
R9080 gnd.n1055 gnd.n1054 42.2793
R9081 gnd.n6026 gnd.n6025 42.2793
R9082 gnd.n5417 gnd.n5416 41.6274
R9083 gnd.n5179 gnd.n5178 41.6274
R9084 gnd.n5426 gnd.n5425 40.8975
R9085 gnd.n5182 gnd.n5181 40.8975
R9086 gnd.n6878 gnd.n538 36.9518
R9087 gnd.n1018 gnd.n1017 36.9518
R9088 gnd.n5425 gnd.n5424 35.055
R9089 gnd.n5420 gnd.n5419 35.055
R9090 gnd.n5171 gnd.n5170 35.055
R9091 gnd.n5181 gnd.n5167 35.055
R9092 gnd.n5812 gnd.n5808 33.2493
R9093 gnd.n5562 gnd.n5561 33.2493
R9094 gnd.n2555 gnd.n2554 32.6173
R9095 gnd.n2555 gnd.n1595 32.6173
R9096 gnd.n2563 gnd.n1595 32.6173
R9097 gnd.n2564 gnd.n2563 32.6173
R9098 gnd.n2565 gnd.n2564 32.6173
R9099 gnd.n2565 gnd.n1589 32.6173
R9100 gnd.n2573 gnd.n1589 32.6173
R9101 gnd.n2574 gnd.n2573 32.6173
R9102 gnd.n2575 gnd.n2574 32.6173
R9103 gnd.n2575 gnd.n1583 32.6173
R9104 gnd.n2583 gnd.n1583 32.6173
R9105 gnd.n2584 gnd.n2583 32.6173
R9106 gnd.n2585 gnd.n2584 32.6173
R9107 gnd.n2585 gnd.n1577 32.6173
R9108 gnd.n2593 gnd.n1577 32.6173
R9109 gnd.n2594 gnd.n2593 32.6173
R9110 gnd.n2595 gnd.n2594 32.6173
R9111 gnd.n2595 gnd.n1571 32.6173
R9112 gnd.n2603 gnd.n1571 32.6173
R9113 gnd.n2604 gnd.n2603 32.6173
R9114 gnd.n2605 gnd.n2604 32.6173
R9115 gnd.n2605 gnd.n1565 32.6173
R9116 gnd.n2613 gnd.n1565 32.6173
R9117 gnd.n2614 gnd.n2613 32.6173
R9118 gnd.n2615 gnd.n2614 32.6173
R9119 gnd.n2615 gnd.n1559 32.6173
R9120 gnd.n2623 gnd.n1559 32.6173
R9121 gnd.n2624 gnd.n2623 32.6173
R9122 gnd.n2625 gnd.n2624 32.6173
R9123 gnd.n2625 gnd.n1553 32.6173
R9124 gnd.n2633 gnd.n1553 32.6173
R9125 gnd.n2634 gnd.n2633 32.6173
R9126 gnd.n2635 gnd.n2634 32.6173
R9127 gnd.n2635 gnd.n1547 32.6173
R9128 gnd.n2643 gnd.n1547 32.6173
R9129 gnd.n2644 gnd.n2643 32.6173
R9130 gnd.n2645 gnd.n2644 32.6173
R9131 gnd.n2645 gnd.n1541 32.6173
R9132 gnd.n2653 gnd.n1541 32.6173
R9133 gnd.n2654 gnd.n2653 32.6173
R9134 gnd.n2655 gnd.n2654 32.6173
R9135 gnd.n2655 gnd.n1535 32.6173
R9136 gnd.n2663 gnd.n1535 32.6173
R9137 gnd.n2664 gnd.n2663 32.6173
R9138 gnd.n2665 gnd.n2664 32.6173
R9139 gnd.n2665 gnd.n1529 32.6173
R9140 gnd.n2673 gnd.n1529 32.6173
R9141 gnd.n2674 gnd.n2673 32.6173
R9142 gnd.n2675 gnd.n2674 32.6173
R9143 gnd.n2675 gnd.n1523 32.6173
R9144 gnd.n2683 gnd.n1523 32.6173
R9145 gnd.n2684 gnd.n2683 32.6173
R9146 gnd.n2685 gnd.n2684 32.6173
R9147 gnd.n2685 gnd.n1517 32.6173
R9148 gnd.n2693 gnd.n1517 32.6173
R9149 gnd.n2694 gnd.n2693 32.6173
R9150 gnd.n2695 gnd.n2694 32.6173
R9151 gnd.n2695 gnd.n1511 32.6173
R9152 gnd.n2703 gnd.n1511 32.6173
R9153 gnd.n2704 gnd.n2703 32.6173
R9154 gnd.n2705 gnd.n2704 32.6173
R9155 gnd.n2705 gnd.n1505 32.6173
R9156 gnd.n2713 gnd.n1505 32.6173
R9157 gnd.n2714 gnd.n2713 32.6173
R9158 gnd.n2715 gnd.n2714 32.6173
R9159 gnd.n2715 gnd.n1499 32.6173
R9160 gnd.n2723 gnd.n1499 32.6173
R9161 gnd.n2724 gnd.n2723 32.6173
R9162 gnd.n2725 gnd.n2724 32.6173
R9163 gnd.n2725 gnd.n1493 32.6173
R9164 gnd.n2733 gnd.n1493 32.6173
R9165 gnd.n2734 gnd.n2733 32.6173
R9166 gnd.n2735 gnd.n2734 32.6173
R9167 gnd.n2735 gnd.n1487 32.6173
R9168 gnd.n2743 gnd.n1487 32.6173
R9169 gnd.n2744 gnd.n2743 32.6173
R9170 gnd.n2745 gnd.n2744 32.6173
R9171 gnd.n2745 gnd.n1481 32.6173
R9172 gnd.n2753 gnd.n1481 32.6173
R9173 gnd.n2754 gnd.n2753 32.6173
R9174 gnd.n2755 gnd.n2754 32.6173
R9175 gnd.n2755 gnd.n1474 32.6173
R9176 gnd.n2766 gnd.n1474 32.6173
R9177 gnd.n3388 gnd.n3282 31.8661
R9178 gnd.n3388 gnd.n3387 31.8661
R9179 gnd.n3396 gnd.n3271 31.8661
R9180 gnd.n3404 gnd.n3271 31.8661
R9181 gnd.n3404 gnd.n3265 31.8661
R9182 gnd.n3412 gnd.n3265 31.8661
R9183 gnd.n3412 gnd.n3258 31.8661
R9184 gnd.n3450 gnd.n3258 31.8661
R9185 gnd.n3460 gnd.n3191 31.8661
R9186 gnd.n4482 gnd.n4284 31.8661
R9187 gnd.n4490 gnd.n1386 31.8661
R9188 gnd.n4498 gnd.n1386 31.8661
R9189 gnd.n4498 gnd.n1378 31.8661
R9190 gnd.n4506 gnd.n1378 31.8661
R9191 gnd.n4514 gnd.n1369 31.8661
R9192 gnd.n4514 gnd.n1372 31.8661
R9193 gnd.n4522 gnd.n1354 31.8661
R9194 gnd.n4530 gnd.n1354 31.8661
R9195 gnd.n4538 gnd.n1346 31.8661
R9196 gnd.n4546 gnd.n1337 31.8661
R9197 gnd.n4546 gnd.n1340 31.8661
R9198 gnd.n4562 gnd.n1320 31.8661
R9199 gnd.n4572 gnd.n1320 31.8661
R9200 gnd.n4585 gnd.n1314 31.8661
R9201 gnd.n4602 gnd.n1296 31.8661
R9202 gnd.n4596 gnd.n1296 31.8661
R9203 gnd.n4611 gnd.n1279 31.8661
R9204 gnd.n4629 gnd.n1279 31.8661
R9205 gnd.n4876 gnd.n1187 31.8661
R9206 gnd.n4870 gnd.n1198 31.8661
R9207 gnd.n4773 gnd.n984 31.8661
R9208 gnd.n4763 gnd.n943 31.8661
R9209 gnd.n6336 gnd.n943 31.8661
R9210 gnd.n6337 gnd.n6336 31.8661
R9211 gnd.n6337 gnd.n936 31.8661
R9212 gnd.n6345 gnd.n936 31.8661
R9213 gnd.n6353 gnd.n929 31.8661
R9214 gnd.n6353 gnd.n921 31.8661
R9215 gnd.n6361 gnd.n921 31.8661
R9216 gnd.n6361 gnd.n923 31.8661
R9217 gnd.n6369 gnd.n907 31.8661
R9218 gnd.n6377 gnd.n907 31.8661
R9219 gnd.n6377 gnd.n909 31.8661
R9220 gnd.n6385 gnd.n901 31.8661
R9221 gnd.n6633 gnd.n668 31.8661
R9222 gnd.n6633 gnd.n661 31.8661
R9223 gnd.n6641 gnd.n661 31.8661
R9224 gnd.n6649 gnd.n654 31.8661
R9225 gnd.n6649 gnd.n646 31.8661
R9226 gnd.n6658 gnd.n646 31.8661
R9227 gnd.n6658 gnd.n648 31.8661
R9228 gnd.n6668 gnd.n639 31.8661
R9229 gnd.n639 gnd.n616 31.8661
R9230 gnd.n6677 gnd.n616 31.8661
R9231 gnd.n6677 gnd.n6676 31.8661
R9232 gnd.n6676 gnd.n489 31.8661
R9233 gnd.n564 gnd.n518 31.8661
R9234 gnd.n7088 gnd.n336 31.8661
R9235 gnd.n7161 gnd.n330 31.8661
R9236 gnd.n7165 gnd.n295 31.8661
R9237 gnd.n7189 gnd.n295 31.8661
R9238 gnd.n7197 gnd.n286 31.8661
R9239 gnd.n7197 gnd.n289 31.8661
R9240 gnd.n7205 gnd.n280 31.8661
R9241 gnd.n7213 gnd.n265 31.8661
R9242 gnd.n7221 gnd.n265 31.8661
R9243 gnd.n7229 gnd.n256 31.8661
R9244 gnd.n7229 gnd.n259 31.8661
R9245 gnd.n7237 gnd.n250 31.8661
R9246 gnd.n7245 gnd.n234 31.8661
R9247 gnd.n7253 gnd.n234 31.8661
R9248 gnd.n7261 gnd.n225 31.8661
R9249 gnd.n7261 gnd.n228 31.8661
R9250 gnd.n7269 gnd.n209 31.8661
R9251 gnd.n7345 gnd.n209 31.8661
R9252 gnd.n7345 gnd.n202 31.8661
R9253 gnd.n7353 gnd.n202 31.8661
R9254 gnd.n7433 gnd.n122 31.8661
R9255 gnd.n4876 gnd.t236 31.5474
R9256 gnd.n7161 gnd.t300 31.5474
R9257 gnd.t269 gnd.n1314 30.9101
R9258 gnd.n909 gnd.t32 30.9101
R9259 gnd.t165 gnd.n668 30.9101
R9260 gnd.n280 gnd.t229 30.9101
R9261 gnd.n6625 gnd.t128 30.5915
R9262 gnd.t219 gnd.n1346 30.2728
R9263 gnd.n250 gnd.t200 30.2728
R9264 gnd.n4284 gnd.t43 28.3609
R9265 gnd.n6393 gnd.n893 28.3609
R9266 gnd.n6617 gnd.n683 28.3609
R9267 gnd.t53 gnd.n122 28.3609
R9268 gnd.n4763 gnd.n992 27.4049
R9269 gnd.n6906 gnd.n489 27.4049
R9270 gnd.n962 gnd.n961 25.7944
R9271 gnd.n3251 gnd.n3250 25.7944
R9272 gnd.n1440 gnd.n1439 25.7944
R9273 gnd.n119 gnd.n118 25.7944
R9274 gnd.n6048 gnd.n6047 25.7944
R9275 gnd.n977 gnd.n976 25.7944
R9276 gnd.n538 gnd.n537 25.7944
R9277 gnd.n560 gnd.n559 25.7944
R9278 gnd.n198 gnd.n197 25.7944
R9279 gnd.n7397 gnd.n7396 25.7944
R9280 gnd.n4313 gnd.n4312 25.7944
R9281 gnd.n4345 gnd.n4344 25.7944
R9282 gnd.n4174 gnd.n4173 25.7944
R9283 gnd.n1054 gnd.n1053 25.7944
R9284 gnd.n1017 gnd.n1016 25.7944
R9285 gnd.n6025 gnd.n6024 25.7944
R9286 gnd.n3472 gnd.n3192 24.8557
R9287 gnd.n3482 gnd.n3175 24.8557
R9288 gnd.n3178 gnd.n3166 24.8557
R9289 gnd.n3503 gnd.n3167 24.8557
R9290 gnd.n3513 gnd.n3147 24.8557
R9291 gnd.n3523 gnd.n3522 24.8557
R9292 gnd.n3131 gnd.n3130 24.8557
R9293 gnd.n3560 gnd.n3123 24.8557
R9294 gnd.n3559 gnd.n3116 24.8557
R9295 gnd.n3597 gnd.n3095 24.8557
R9296 gnd.n3571 gnd.n3096 24.8557
R9297 gnd.n3590 gnd.n2943 24.8557
R9298 gnd.n3607 gnd.n3606 24.8557
R9299 gnd.n3618 gnd.n3617 24.8557
R9300 gnd.n2935 gnd.n2926 24.8557
R9301 gnd.n3638 gnd.n2909 24.8557
R9302 gnd.n2912 gnd.n2901 24.8557
R9303 gnd.n3659 gnd.n2902 24.8557
R9304 gnd.n3668 gnd.n2894 24.8557
R9305 gnd.n3669 gnd.n2883 24.8557
R9306 gnd.n2886 gnd.n2874 24.8557
R9307 gnd.n3690 gnd.n2875 24.8557
R9308 gnd.n3700 gnd.n2858 24.8557
R9309 gnd.n3711 gnd.n3710 24.8557
R9310 gnd.n3000 gnd.n2999 24.8557
R9311 gnd.n3721 gnd.n2850 24.8557
R9312 gnd.n3731 gnd.n2833 24.8557
R9313 gnd.n3742 gnd.n3741 24.8557
R9314 gnd.n3752 gnd.n2825 24.8557
R9315 gnd.n3762 gnd.n2807 24.8557
R9316 gnd.n3773 gnd.n3772 24.8557
R9317 gnd.n3783 gnd.n2800 24.8557
R9318 gnd.n4048 gnd.n2792 24.8557
R9319 gnd.n4049 gnd.n2782 24.8557
R9320 gnd.n5386 gnd.n5385 23.855
R9321 gnd.n5213 gnd.n5212 23.855
R9322 gnd.n5394 gnd.n5393 23.855
R9323 gnd.n5207 gnd.n5206 23.855
R9324 gnd.n3493 gnd.t0 23.2624
R9325 gnd.n4506 gnd.t246 23.2624
R9326 gnd.n7269 gnd.t271 23.2624
R9327 gnd.n3194 gnd.t39 22.6251
R9328 gnd.n4538 gnd.t217 22.6251
R9329 gnd.n7237 gnd.t186 22.6251
R9330 gnd.n4585 gnd.t194 21.9878
R9331 gnd.n7205 gnd.t241 21.9878
R9332 gnd.n5585 gnd.n869 21.6691
R9333 gnd.n5594 gnd.n862 21.6691
R9334 gnd.n5602 gnd.n854 21.6691
R9335 gnd.n5620 gnd.n848 21.6691
R9336 gnd.n5332 gnd.n841 21.6691
R9337 gnd.n5667 gnd.n811 21.6691
R9338 gnd.n5308 gnd.n803 21.6691
R9339 gnd.n5684 gnd.n795 21.6691
R9340 gnd.n5693 gnd.n779 21.6691
R9341 gnd.n5702 gnd.n771 21.6691
R9342 gnd.n5711 gnd.n763 21.6691
R9343 gnd.n5746 gnd.n733 21.6691
R9344 gnd.n5754 gnd.n726 21.6691
R9345 gnd.n5252 gnd.n720 21.6691
R9346 gnd.n5781 gnd.n712 21.6691
R9347 gnd.n5934 gnd.n690 21.6691
R9348 gnd.t169 gnd.n3199 21.3504
R9349 gnd.t198 gnd.n1187 21.3504
R9350 gnd.n1200 gnd.n1198 21.3504
R9351 gnd.n4645 gnd.t221 21.3504
R9352 gnd.n7062 gnd.t210 21.3504
R9353 gnd.n7081 gnd.n336 21.3504
R9354 gnd.t290 gnd.n330 21.3504
R9355 gnd.n5430 gnd.n5429 21.0737
R9356 gnd.n5931 gnd.n5930 21.0737
R9357 gnd.n6433 gnd.n856 21.0318
R9358 gnd.n5302 gnd.n786 21.0318
R9359 gnd.n5297 gnd.n788 21.0318
R9360 gnd.n6577 gnd.n718 21.0318
R9361 gnd.t14 gnd.n2824 20.7131
R9362 gnd.n4611 gnd.t180 20.7131
R9363 gnd.n6369 gnd.t342 20.7131
R9364 gnd.n6641 gnd.t340 20.7131
R9365 gnd.n7189 gnd.t248 20.7131
R9366 gnd.t68 gnd.n5796 20.3945
R9367 gnd.n3699 gnd.t16 20.0758
R9368 gnd.n4562 gnd.t250 20.0758
R9369 gnd.n7221 gnd.t282 20.0758
R9370 gnd.n5413 gnd.t97 19.8005
R9371 gnd.n5413 gnd.t135 19.8005
R9372 gnd.n5414 gnd.t120 19.8005
R9373 gnd.n5414 gnd.t66 19.8005
R9374 gnd.n5175 gnd.t48 19.8005
R9375 gnd.n5175 gnd.t129 19.8005
R9376 gnd.n5176 gnd.t138 19.8005
R9377 gnd.n5176 gnd.t117 19.8005
R9378 gnd.n5567 gnd.t119 19.7572
R9379 gnd.n6449 gnd.t26 19.7572
R9380 gnd.n5676 gnd.n5307 19.7572
R9381 gnd.n5292 gnd.n5291 19.7572
R9382 gnd.n6561 gnd.t151 19.7572
R9383 gnd.n2767 gnd.n2766 19.5706
R9384 gnd.n5410 gnd.n5409 19.5087
R9385 gnd.n5423 gnd.n5410 19.5087
R9386 gnd.n5421 gnd.n5412 19.5087
R9387 gnd.n5180 gnd.n5174 19.5087
R9388 gnd.t18 gnd.n3648 19.4385
R9389 gnd.n4522 gnd.t196 19.4385
R9390 gnd.n6347 gnd.n934 19.3944
R9391 gnd.n6347 gnd.n932 19.3944
R9392 gnd.n6351 gnd.n932 19.3944
R9393 gnd.n6351 gnd.n919 19.3944
R9394 gnd.n6363 gnd.n919 19.3944
R9395 gnd.n6363 gnd.n917 19.3944
R9396 gnd.n6367 gnd.n917 19.3944
R9397 gnd.n6367 gnd.n905 19.3944
R9398 gnd.n6379 gnd.n905 19.3944
R9399 gnd.n6379 gnd.n903 19.3944
R9400 gnd.n6383 gnd.n903 19.3944
R9401 gnd.n6383 gnd.n891 19.3944
R9402 gnd.n6395 gnd.n891 19.3944
R9403 gnd.n6395 gnd.n889 19.3944
R9404 gnd.n6399 gnd.n889 19.3944
R9405 gnd.n6399 gnd.n875 19.3944
R9406 gnd.n6411 gnd.n875 19.3944
R9407 gnd.n6411 gnd.n873 19.3944
R9408 gnd.n6415 gnd.n873 19.3944
R9409 gnd.n6415 gnd.n860 19.3944
R9410 gnd.n6427 gnd.n860 19.3944
R9411 gnd.n6427 gnd.n858 19.3944
R9412 gnd.n6431 gnd.n858 19.3944
R9413 gnd.n6431 gnd.n845 19.3944
R9414 gnd.n6443 gnd.n845 19.3944
R9415 gnd.n6443 gnd.n843 19.3944
R9416 gnd.n6447 gnd.n843 19.3944
R9417 gnd.n6447 gnd.n831 19.3944
R9418 gnd.n6459 gnd.n831 19.3944
R9419 gnd.n6459 gnd.n829 19.3944
R9420 gnd.n6463 gnd.n829 19.3944
R9421 gnd.n6463 gnd.n815 19.3944
R9422 gnd.n6475 gnd.n815 19.3944
R9423 gnd.n6475 gnd.n813 19.3944
R9424 gnd.n6479 gnd.n813 19.3944
R9425 gnd.n6479 gnd.n799 19.3944
R9426 gnd.n6491 gnd.n799 19.3944
R9427 gnd.n6491 gnd.n797 19.3944
R9428 gnd.n6495 gnd.n797 19.3944
R9429 gnd.n6495 gnd.n784 19.3944
R9430 gnd.n6507 gnd.n784 19.3944
R9431 gnd.n6507 gnd.n782 19.3944
R9432 gnd.n6511 gnd.n782 19.3944
R9433 gnd.n6511 gnd.n769 19.3944
R9434 gnd.n6523 gnd.n769 19.3944
R9435 gnd.n6523 gnd.n767 19.3944
R9436 gnd.n6527 gnd.n767 19.3944
R9437 gnd.n6527 gnd.n753 19.3944
R9438 gnd.n6539 gnd.n753 19.3944
R9439 gnd.n6539 gnd.n751 19.3944
R9440 gnd.n6543 gnd.n751 19.3944
R9441 gnd.n6543 gnd.n738 19.3944
R9442 gnd.n6555 gnd.n738 19.3944
R9443 gnd.n6555 gnd.n736 19.3944
R9444 gnd.n6559 gnd.n736 19.3944
R9445 gnd.n6559 gnd.n724 19.3944
R9446 gnd.n6571 gnd.n724 19.3944
R9447 gnd.n6571 gnd.n722 19.3944
R9448 gnd.n6575 gnd.n722 19.3944
R9449 gnd.n6575 gnd.n709 19.3944
R9450 gnd.n6587 gnd.n709 19.3944
R9451 gnd.n6587 gnd.n707 19.3944
R9452 gnd.n6591 gnd.n707 19.3944
R9453 gnd.n6591 gnd.n694 19.3944
R9454 gnd.n6603 gnd.n694 19.3944
R9455 gnd.n6603 gnd.n692 19.3944
R9456 gnd.n6607 gnd.n692 19.3944
R9457 gnd.n6607 gnd.n679 19.3944
R9458 gnd.n6619 gnd.n679 19.3944
R9459 gnd.n6619 gnd.n677 19.3944
R9460 gnd.n6623 gnd.n677 19.3944
R9461 gnd.n6623 gnd.n666 19.3944
R9462 gnd.n6635 gnd.n666 19.3944
R9463 gnd.n6635 gnd.n664 19.3944
R9464 gnd.n6639 gnd.n664 19.3944
R9465 gnd.n6639 gnd.n652 19.3944
R9466 gnd.n6651 gnd.n652 19.3944
R9467 gnd.n6651 gnd.n650 19.3944
R9468 gnd.n6656 gnd.n650 19.3944
R9469 gnd.n6656 gnd.n636 19.3944
R9470 gnd.n6670 gnd.n636 19.3944
R9471 gnd.n6671 gnd.n6670 19.3944
R9472 gnd.n6330 gnd.n6327 19.3944
R9473 gnd.n6330 gnd.n959 19.3944
R9474 gnd.n6334 gnd.n959 19.3944
R9475 gnd.n5092 gnd.n5091 19.3944
R9476 gnd.n5091 gnd.n4994 19.3944
R9477 gnd.n5084 gnd.n4994 19.3944
R9478 gnd.n5084 gnd.n5083 19.3944
R9479 gnd.n5083 gnd.n5010 19.3944
R9480 gnd.n5076 gnd.n5010 19.3944
R9481 gnd.n5076 gnd.n5075 19.3944
R9482 gnd.n5075 gnd.n5022 19.3944
R9483 gnd.n5068 gnd.n5022 19.3944
R9484 gnd.n5068 gnd.n5067 19.3944
R9485 gnd.n5067 gnd.n5033 19.3944
R9486 gnd.n5060 gnd.n5033 19.3944
R9487 gnd.n5060 gnd.n5059 19.3944
R9488 gnd.n5059 gnd.n5045 19.3944
R9489 gnd.n5045 gnd.n972 19.3944
R9490 gnd.n6308 gnd.n972 19.3944
R9491 gnd.n6309 gnd.n6308 19.3944
R9492 gnd.n6312 gnd.n6309 19.3944
R9493 gnd.n6312 gnd.n967 19.3944
R9494 gnd.n6317 gnd.n967 19.3944
R9495 gnd.n6318 gnd.n6317 19.3944
R9496 gnd.n6321 gnd.n6318 19.3944
R9497 gnd.n6321 gnd.n963 19.3944
R9498 gnd.n6325 gnd.n963 19.3944
R9499 gnd.n3375 gnd.n3374 19.3944
R9500 gnd.n3374 gnd.n3373 19.3944
R9501 gnd.n3373 gnd.n3372 19.3944
R9502 gnd.n3372 gnd.n3370 19.3944
R9503 gnd.n3370 gnd.n3367 19.3944
R9504 gnd.n3367 gnd.n3366 19.3944
R9505 gnd.n3366 gnd.n3363 19.3944
R9506 gnd.n3363 gnd.n3362 19.3944
R9507 gnd.n3362 gnd.n3359 19.3944
R9508 gnd.n3359 gnd.n3358 19.3944
R9509 gnd.n3358 gnd.n3355 19.3944
R9510 gnd.n3355 gnd.n3354 19.3944
R9511 gnd.n3354 gnd.n3351 19.3944
R9512 gnd.n3351 gnd.n3350 19.3944
R9513 gnd.n3350 gnd.n3347 19.3944
R9514 gnd.n3347 gnd.n3346 19.3944
R9515 gnd.n3346 gnd.n3343 19.3944
R9516 gnd.n3343 gnd.n3342 19.3944
R9517 gnd.n3342 gnd.n3339 19.3944
R9518 gnd.n3339 gnd.n3338 19.3944
R9519 gnd.n3338 gnd.n3335 19.3944
R9520 gnd.n3335 gnd.n3334 19.3944
R9521 gnd.n3331 gnd.n3330 19.3944
R9522 gnd.n3330 gnd.n3286 19.3944
R9523 gnd.n3381 gnd.n3286 19.3944
R9524 gnd.n4084 gnd.n4083 19.3944
R9525 gnd.n4083 gnd.n4080 19.3944
R9526 gnd.n4080 gnd.n4079 19.3944
R9527 gnd.n4129 gnd.n4128 19.3944
R9528 gnd.n4128 gnd.n4127 19.3944
R9529 gnd.n4127 gnd.n4124 19.3944
R9530 gnd.n4124 gnd.n4123 19.3944
R9531 gnd.n4123 gnd.n4120 19.3944
R9532 gnd.n4120 gnd.n4119 19.3944
R9533 gnd.n4119 gnd.n4116 19.3944
R9534 gnd.n4116 gnd.n4115 19.3944
R9535 gnd.n4115 gnd.n4112 19.3944
R9536 gnd.n4112 gnd.n4111 19.3944
R9537 gnd.n4111 gnd.n4108 19.3944
R9538 gnd.n4108 gnd.n4107 19.3944
R9539 gnd.n4107 gnd.n4104 19.3944
R9540 gnd.n4104 gnd.n4103 19.3944
R9541 gnd.n4103 gnd.n4100 19.3944
R9542 gnd.n4100 gnd.n4099 19.3944
R9543 gnd.n4099 gnd.n4096 19.3944
R9544 gnd.n4096 gnd.n4095 19.3944
R9545 gnd.n4095 gnd.n4092 19.3944
R9546 gnd.n4092 gnd.n4091 19.3944
R9547 gnd.n4091 gnd.n4088 19.3944
R9548 gnd.n4088 gnd.n4087 19.3944
R9549 gnd.n3474 gnd.n3183 19.3944
R9550 gnd.n3484 gnd.n3183 19.3944
R9551 gnd.n3485 gnd.n3484 19.3944
R9552 gnd.n3485 gnd.n3164 19.3944
R9553 gnd.n3505 gnd.n3164 19.3944
R9554 gnd.n3505 gnd.n3156 19.3944
R9555 gnd.n3515 gnd.n3156 19.3944
R9556 gnd.n3516 gnd.n3515 19.3944
R9557 gnd.n3517 gnd.n3516 19.3944
R9558 gnd.n3517 gnd.n3139 19.3944
R9559 gnd.n3139 gnd.n3137 19.3944
R9560 gnd.n3543 gnd.n3137 19.3944
R9561 gnd.n3543 gnd.n3119 19.3944
R9562 gnd.n3577 gnd.n3119 19.3944
R9563 gnd.n3577 gnd.n3576 19.3944
R9564 gnd.n3576 gnd.n3575 19.3944
R9565 gnd.n3575 gnd.n3570 19.3944
R9566 gnd.n3570 gnd.n2940 19.3944
R9567 gnd.n3609 gnd.n2940 19.3944
R9568 gnd.n3610 gnd.n3609 19.3944
R9569 gnd.n3610 gnd.n2924 19.3944
R9570 gnd.n3630 gnd.n2924 19.3944
R9571 gnd.n3630 gnd.n2917 19.3944
R9572 gnd.n3640 gnd.n2917 19.3944
R9573 gnd.n3641 gnd.n3640 19.3944
R9574 gnd.n3641 gnd.n2899 19.3944
R9575 gnd.n3661 gnd.n2899 19.3944
R9576 gnd.n3661 gnd.n2891 19.3944
R9577 gnd.n3671 gnd.n2891 19.3944
R9578 gnd.n3672 gnd.n3671 19.3944
R9579 gnd.n3672 gnd.n2872 19.3944
R9580 gnd.n3692 gnd.n2872 19.3944
R9581 gnd.n3692 gnd.n2865 19.3944
R9582 gnd.n3702 gnd.n2865 19.3944
R9583 gnd.n3703 gnd.n3702 19.3944
R9584 gnd.n3703 gnd.n2848 19.3944
R9585 gnd.n3723 gnd.n2848 19.3944
R9586 gnd.n3723 gnd.n2841 19.3944
R9587 gnd.n3733 gnd.n2841 19.3944
R9588 gnd.n3734 gnd.n3733 19.3944
R9589 gnd.n3734 gnd.n2822 19.3944
R9590 gnd.n3754 gnd.n2822 19.3944
R9591 gnd.n3754 gnd.n2815 19.3944
R9592 gnd.n3764 gnd.n2815 19.3944
R9593 gnd.n3765 gnd.n3764 19.3944
R9594 gnd.n3765 gnd.n2797 19.3944
R9595 gnd.n3785 gnd.n2797 19.3944
R9596 gnd.n3785 gnd.n2789 19.3944
R9597 gnd.n4051 gnd.n2789 19.3944
R9598 gnd.n4052 gnd.n4051 19.3944
R9599 gnd.n4052 gnd.n2771 19.3944
R9600 gnd.n4071 gnd.n2771 19.3944
R9601 gnd.n4071 gnd.n2772 19.3944
R9602 gnd.n3465 gnd.n3464 19.3944
R9603 gnd.n3464 gnd.n3197 19.3944
R9604 gnd.n3220 gnd.n3197 19.3944
R9605 gnd.n3223 gnd.n3220 19.3944
R9606 gnd.n3223 gnd.n3216 19.3944
R9607 gnd.n3227 gnd.n3216 19.3944
R9608 gnd.n3230 gnd.n3227 19.3944
R9609 gnd.n3233 gnd.n3230 19.3944
R9610 gnd.n3233 gnd.n3214 19.3944
R9611 gnd.n3237 gnd.n3214 19.3944
R9612 gnd.n3240 gnd.n3237 19.3944
R9613 gnd.n3243 gnd.n3240 19.3944
R9614 gnd.n3243 gnd.n3212 19.3944
R9615 gnd.n3247 gnd.n3212 19.3944
R9616 gnd.n3470 gnd.n3469 19.3944
R9617 gnd.n3469 gnd.n3173 19.3944
R9618 gnd.n3495 gnd.n3173 19.3944
R9619 gnd.n3495 gnd.n3171 19.3944
R9620 gnd.n3501 gnd.n3171 19.3944
R9621 gnd.n3501 gnd.n3500 19.3944
R9622 gnd.n3500 gnd.n3145 19.3944
R9623 gnd.n3525 gnd.n3145 19.3944
R9624 gnd.n3525 gnd.n3143 19.3944
R9625 gnd.n3537 gnd.n3143 19.3944
R9626 gnd.n3537 gnd.n3536 19.3944
R9627 gnd.n3536 gnd.n3535 19.3944
R9628 gnd.n3535 gnd.n3533 19.3944
R9629 gnd.n3533 gnd.n3115 19.3944
R9630 gnd.n3115 gnd.n3113 19.3944
R9631 gnd.n3584 gnd.n3113 19.3944
R9632 gnd.n3584 gnd.n3111 19.3944
R9633 gnd.n3588 gnd.n3111 19.3944
R9634 gnd.n3588 gnd.n2931 19.3944
R9635 gnd.n3620 gnd.n2931 19.3944
R9636 gnd.n3620 gnd.n2929 19.3944
R9637 gnd.n3626 gnd.n2929 19.3944
R9638 gnd.n3626 gnd.n3625 19.3944
R9639 gnd.n3625 gnd.n2907 19.3944
R9640 gnd.n3651 gnd.n2907 19.3944
R9641 gnd.n3651 gnd.n2905 19.3944
R9642 gnd.n3657 gnd.n2905 19.3944
R9643 gnd.n3657 gnd.n3656 19.3944
R9644 gnd.n3656 gnd.n2881 19.3944
R9645 gnd.n3682 gnd.n2881 19.3944
R9646 gnd.n3682 gnd.n2879 19.3944
R9647 gnd.n3688 gnd.n2879 19.3944
R9648 gnd.n3688 gnd.n3687 19.3944
R9649 gnd.n3687 gnd.n2856 19.3944
R9650 gnd.n3713 gnd.n2856 19.3944
R9651 gnd.n3713 gnd.n2854 19.3944
R9652 gnd.n3719 gnd.n2854 19.3944
R9653 gnd.n3719 gnd.n3718 19.3944
R9654 gnd.n3718 gnd.n2831 19.3944
R9655 gnd.n3744 gnd.n2831 19.3944
R9656 gnd.n3744 gnd.n2829 19.3944
R9657 gnd.n3750 gnd.n2829 19.3944
R9658 gnd.n3750 gnd.n3749 19.3944
R9659 gnd.n3749 gnd.n2805 19.3944
R9660 gnd.n3775 gnd.n2805 19.3944
R9661 gnd.n3775 gnd.n2803 19.3944
R9662 gnd.n3781 gnd.n2803 19.3944
R9663 gnd.n3781 gnd.n3780 19.3944
R9664 gnd.n3780 gnd.n2780 19.3944
R9665 gnd.n4061 gnd.n2780 19.3944
R9666 gnd.n4061 gnd.n2778 19.3944
R9667 gnd.n4067 gnd.n2778 19.3944
R9668 gnd.n4067 gnd.n4066 19.3944
R9669 gnd.n4165 gnd.n4164 19.3944
R9670 gnd.n4164 gnd.n1426 19.3944
R9671 gnd.n4160 gnd.n1426 19.3944
R9672 gnd.n4160 gnd.n4157 19.3944
R9673 gnd.n4157 gnd.n4154 19.3944
R9674 gnd.n4154 gnd.n4153 19.3944
R9675 gnd.n4153 gnd.n4150 19.3944
R9676 gnd.n4150 gnd.n4149 19.3944
R9677 gnd.n4149 gnd.n4146 19.3944
R9678 gnd.n4146 gnd.n4145 19.3944
R9679 gnd.n4145 gnd.n4142 19.3944
R9680 gnd.n4142 gnd.n4141 19.3944
R9681 gnd.n4141 gnd.n4138 19.3944
R9682 gnd.n4138 gnd.n4137 19.3944
R9683 gnd.n3385 gnd.n3284 19.3944
R9684 gnd.n3385 gnd.n3275 19.3944
R9685 gnd.n3398 gnd.n3275 19.3944
R9686 gnd.n3398 gnd.n3273 19.3944
R9687 gnd.n3402 gnd.n3273 19.3944
R9688 gnd.n3402 gnd.n3263 19.3944
R9689 gnd.n3414 gnd.n3263 19.3944
R9690 gnd.n3414 gnd.n3261 19.3944
R9691 gnd.n3448 gnd.n3261 19.3944
R9692 gnd.n3448 gnd.n3447 19.3944
R9693 gnd.n3447 gnd.n3446 19.3944
R9694 gnd.n3446 gnd.n3445 19.3944
R9695 gnd.n3445 gnd.n3442 19.3944
R9696 gnd.n3442 gnd.n3441 19.3944
R9697 gnd.n3441 gnd.n3440 19.3944
R9698 gnd.n3440 gnd.n3438 19.3944
R9699 gnd.n3438 gnd.n3437 19.3944
R9700 gnd.n3437 gnd.n3434 19.3944
R9701 gnd.n3434 gnd.n3433 19.3944
R9702 gnd.n3433 gnd.n3432 19.3944
R9703 gnd.n3432 gnd.n3430 19.3944
R9704 gnd.n3430 gnd.n3128 19.3944
R9705 gnd.n3551 gnd.n3128 19.3944
R9706 gnd.n3551 gnd.n3126 19.3944
R9707 gnd.n3557 gnd.n3126 19.3944
R9708 gnd.n3557 gnd.n3556 19.3944
R9709 gnd.n3556 gnd.n3091 19.3944
R9710 gnd.n3599 gnd.n3091 19.3944
R9711 gnd.n3599 gnd.n3092 19.3944
R9712 gnd.n3108 gnd.n3107 19.3944
R9713 gnd.n3604 gnd.n3603 19.3944
R9714 gnd.n3027 gnd.n2946 19.3944
R9715 gnd.n3022 gnd.n3021 19.3944
R9716 gnd.n3021 gnd.n3019 19.3944
R9717 gnd.n3019 gnd.n3018 19.3944
R9718 gnd.n3018 gnd.n3015 19.3944
R9719 gnd.n3015 gnd.n3014 19.3944
R9720 gnd.n3014 gnd.n3013 19.3944
R9721 gnd.n3013 gnd.n3011 19.3944
R9722 gnd.n3011 gnd.n3010 19.3944
R9723 gnd.n3010 gnd.n3007 19.3944
R9724 gnd.n3007 gnd.n3006 19.3944
R9725 gnd.n3006 gnd.n3005 19.3944
R9726 gnd.n3005 gnd.n3003 19.3944
R9727 gnd.n3003 gnd.n3002 19.3944
R9728 gnd.n3002 gnd.n2997 19.3944
R9729 gnd.n2997 gnd.n2996 19.3944
R9730 gnd.n2996 gnd.n2995 19.3944
R9731 gnd.n2995 gnd.n2993 19.3944
R9732 gnd.n2993 gnd.n2992 19.3944
R9733 gnd.n2992 gnd.n2989 19.3944
R9734 gnd.n2989 gnd.n2988 19.3944
R9735 gnd.n2988 gnd.n2987 19.3944
R9736 gnd.n2987 gnd.n2985 19.3944
R9737 gnd.n2985 gnd.n2984 19.3944
R9738 gnd.n2984 gnd.n2981 19.3944
R9739 gnd.n2981 gnd.n2980 19.3944
R9740 gnd.n2980 gnd.n2979 19.3944
R9741 gnd.n2979 gnd.n2977 19.3944
R9742 gnd.n2977 gnd.n2976 19.3944
R9743 gnd.n2976 gnd.n1473 19.3944
R9744 gnd.n3390 gnd.n3280 19.3944
R9745 gnd.n3390 gnd.n3278 19.3944
R9746 gnd.n3394 gnd.n3278 19.3944
R9747 gnd.n3394 gnd.n3269 19.3944
R9748 gnd.n3406 gnd.n3269 19.3944
R9749 gnd.n3406 gnd.n3267 19.3944
R9750 gnd.n3410 gnd.n3267 19.3944
R9751 gnd.n3410 gnd.n3256 19.3944
R9752 gnd.n3452 gnd.n3256 19.3944
R9753 gnd.n3452 gnd.n3210 19.3944
R9754 gnd.n3458 gnd.n3210 19.3944
R9755 gnd.n3458 gnd.n3457 19.3944
R9756 gnd.n3457 gnd.n3188 19.3944
R9757 gnd.n3479 gnd.n3188 19.3944
R9758 gnd.n3479 gnd.n3181 19.3944
R9759 gnd.n3490 gnd.n3181 19.3944
R9760 gnd.n3490 gnd.n3489 19.3944
R9761 gnd.n3489 gnd.n3162 19.3944
R9762 gnd.n3510 gnd.n3162 19.3944
R9763 gnd.n3510 gnd.n3152 19.3944
R9764 gnd.n3520 gnd.n3152 19.3944
R9765 gnd.n3520 gnd.n3133 19.3944
R9766 gnd.n3547 gnd.n3133 19.3944
R9767 gnd.n3547 gnd.n3546 19.3944
R9768 gnd.n3546 gnd.n3121 19.3944
R9769 gnd.n3563 gnd.n3121 19.3944
R9770 gnd.n3563 gnd.n3099 19.3944
R9771 gnd.n3595 gnd.n3099 19.3944
R9772 gnd.n3595 gnd.n3594 19.3944
R9773 gnd.n3594 gnd.n3593 19.3944
R9774 gnd.n3593 gnd.n3105 19.3944
R9775 gnd.n3105 gnd.n2938 19.3944
R9776 gnd.n3615 gnd.n2938 19.3944
R9777 gnd.n3615 gnd.n3614 19.3944
R9778 gnd.n3614 gnd.n2922 19.3944
R9779 gnd.n3635 gnd.n2922 19.3944
R9780 gnd.n3635 gnd.n2915 19.3944
R9781 gnd.n3646 gnd.n2915 19.3944
R9782 gnd.n3646 gnd.n3645 19.3944
R9783 gnd.n3645 gnd.n2897 19.3944
R9784 gnd.n3666 gnd.n2897 19.3944
R9785 gnd.n3666 gnd.n2889 19.3944
R9786 gnd.n3677 gnd.n2889 19.3944
R9787 gnd.n3677 gnd.n3676 19.3944
R9788 gnd.n3676 gnd.n2870 19.3944
R9789 gnd.n3697 gnd.n2870 19.3944
R9790 gnd.n3697 gnd.n2863 19.3944
R9791 gnd.n3708 gnd.n2863 19.3944
R9792 gnd.n3708 gnd.n3707 19.3944
R9793 gnd.n3707 gnd.n2846 19.3944
R9794 gnd.n3728 gnd.n2846 19.3944
R9795 gnd.n3728 gnd.n2839 19.3944
R9796 gnd.n3739 gnd.n2839 19.3944
R9797 gnd.n3739 gnd.n3738 19.3944
R9798 gnd.n3738 gnd.n2820 19.3944
R9799 gnd.n3759 gnd.n2820 19.3944
R9800 gnd.n3759 gnd.n2813 19.3944
R9801 gnd.n3770 gnd.n2813 19.3944
R9802 gnd.n3770 gnd.n3769 19.3944
R9803 gnd.n3769 gnd.n2795 19.3944
R9804 gnd.n4046 gnd.n2795 19.3944
R9805 gnd.n4046 gnd.n2787 19.3944
R9806 gnd.n4056 gnd.n2787 19.3944
R9807 gnd.n4056 gnd.n2769 19.3944
R9808 gnd.n4074 gnd.n2769 19.3944
R9809 gnd.n6832 gnd.n565 19.3944
R9810 gnd.n6828 gnd.n565 19.3944
R9811 gnd.n6828 gnd.n6827 19.3944
R9812 gnd.n6827 gnd.n6826 19.3944
R9813 gnd.n6826 gnd.n570 19.3944
R9814 gnd.n6822 gnd.n570 19.3944
R9815 gnd.n6822 gnd.n6821 19.3944
R9816 gnd.n6821 gnd.n6820 19.3944
R9817 gnd.n6820 gnd.n574 19.3944
R9818 gnd.n6816 gnd.n574 19.3944
R9819 gnd.n6816 gnd.n6815 19.3944
R9820 gnd.n6815 gnd.n6814 19.3944
R9821 gnd.n6814 gnd.n578 19.3944
R9822 gnd.n6810 gnd.n578 19.3944
R9823 gnd.n6810 gnd.n6809 19.3944
R9824 gnd.n6809 gnd.n6808 19.3944
R9825 gnd.n6808 gnd.n582 19.3944
R9826 gnd.n6804 gnd.n582 19.3944
R9827 gnd.n6804 gnd.n6803 19.3944
R9828 gnd.n6803 gnd.n6802 19.3944
R9829 gnd.n6802 gnd.n384 19.3944
R9830 gnd.n7021 gnd.n384 19.3944
R9831 gnd.n7022 gnd.n7021 19.3944
R9832 gnd.n7022 gnd.n381 19.3944
R9833 gnd.n7027 gnd.n381 19.3944
R9834 gnd.n7027 gnd.n382 19.3944
R9835 gnd.n382 gnd.n352 19.3944
R9836 gnd.n7069 gnd.n352 19.3944
R9837 gnd.n7069 gnd.n353 19.3944
R9838 gnd.n7065 gnd.n353 19.3944
R9839 gnd.n7065 gnd.n7064 19.3944
R9840 gnd.n7064 gnd.n76 19.3944
R9841 gnd.n7484 gnd.n76 19.3944
R9842 gnd.n7484 gnd.n7483 19.3944
R9843 gnd.n7483 gnd.n7482 19.3944
R9844 gnd.n7482 gnd.n81 19.3944
R9845 gnd.n7478 gnd.n81 19.3944
R9846 gnd.n7478 gnd.n7477 19.3944
R9847 gnd.n7477 gnd.n7476 19.3944
R9848 gnd.n7476 gnd.n86 19.3944
R9849 gnd.n7472 gnd.n86 19.3944
R9850 gnd.n7472 gnd.n7471 19.3944
R9851 gnd.n7471 gnd.n7470 19.3944
R9852 gnd.n7470 gnd.n91 19.3944
R9853 gnd.n7466 gnd.n91 19.3944
R9854 gnd.n7466 gnd.n7465 19.3944
R9855 gnd.n7465 gnd.n7464 19.3944
R9856 gnd.n7464 gnd.n96 19.3944
R9857 gnd.n7460 gnd.n96 19.3944
R9858 gnd.n7460 gnd.n7459 19.3944
R9859 gnd.n7459 gnd.n7458 19.3944
R9860 gnd.n7458 gnd.n101 19.3944
R9861 gnd.n7454 gnd.n101 19.3944
R9862 gnd.n7454 gnd.n7453 19.3944
R9863 gnd.n7453 gnd.n7452 19.3944
R9864 gnd.n7452 gnd.n106 19.3944
R9865 gnd.n7448 gnd.n106 19.3944
R9866 gnd.n7448 gnd.n7447 19.3944
R9867 gnd.n7447 gnd.n7446 19.3944
R9868 gnd.n7446 gnd.n111 19.3944
R9869 gnd.n7442 gnd.n111 19.3944
R9870 gnd.n7442 gnd.n7441 19.3944
R9871 gnd.n7441 gnd.n7440 19.3944
R9872 gnd.n7440 gnd.n116 19.3944
R9873 gnd.n7334 gnd.n7333 19.3944
R9874 gnd.n7333 gnd.n7332 19.3944
R9875 gnd.n7332 gnd.n7281 19.3944
R9876 gnd.n7328 gnd.n7281 19.3944
R9877 gnd.n7328 gnd.n7327 19.3944
R9878 gnd.n7327 gnd.n7326 19.3944
R9879 gnd.n7326 gnd.n7289 19.3944
R9880 gnd.n7322 gnd.n7289 19.3944
R9881 gnd.n7322 gnd.n7321 19.3944
R9882 gnd.n7321 gnd.n7320 19.3944
R9883 gnd.n7320 gnd.n7297 19.3944
R9884 gnd.n7316 gnd.n7297 19.3944
R9885 gnd.n7316 gnd.n7315 19.3944
R9886 gnd.n7315 gnd.n7314 19.3944
R9887 gnd.n7314 gnd.n7305 19.3944
R9888 gnd.n7310 gnd.n7305 19.3944
R9889 gnd.n5958 gnd.n5957 19.3944
R9890 gnd.n6089 gnd.n5958 19.3944
R9891 gnd.n6089 gnd.n6088 19.3944
R9892 gnd.n6088 gnd.n5963 19.3944
R9893 gnd.n6081 gnd.n5963 19.3944
R9894 gnd.n6081 gnd.n6080 19.3944
R9895 gnd.n6080 gnd.n5973 19.3944
R9896 gnd.n6073 gnd.n5973 19.3944
R9897 gnd.n6073 gnd.n6072 19.3944
R9898 gnd.n6072 gnd.n5983 19.3944
R9899 gnd.n6065 gnd.n5983 19.3944
R9900 gnd.n6065 gnd.n6064 19.3944
R9901 gnd.n6064 gnd.n5993 19.3944
R9902 gnd.n6057 gnd.n5993 19.3944
R9903 gnd.n6057 gnd.n6056 19.3944
R9904 gnd.n6056 gnd.n6003 19.3944
R9905 gnd.n6917 gnd.n478 19.3944
R9906 gnd.n6917 gnd.n476 19.3944
R9907 gnd.n6921 gnd.n476 19.3944
R9908 gnd.n6921 gnd.n460 19.3944
R9909 gnd.n6933 gnd.n460 19.3944
R9910 gnd.n6933 gnd.n458 19.3944
R9911 gnd.n6937 gnd.n458 19.3944
R9912 gnd.n6937 gnd.n444 19.3944
R9913 gnd.n6949 gnd.n444 19.3944
R9914 gnd.n6949 gnd.n442 19.3944
R9915 gnd.n6953 gnd.n442 19.3944
R9916 gnd.n6953 gnd.n426 19.3944
R9917 gnd.n6965 gnd.n426 19.3944
R9918 gnd.n6965 gnd.n424 19.3944
R9919 gnd.n6969 gnd.n424 19.3944
R9920 gnd.n6969 gnd.n410 19.3944
R9921 gnd.n6981 gnd.n410 19.3944
R9922 gnd.n6981 gnd.n407 19.3944
R9923 gnd.n6988 gnd.n407 19.3944
R9924 gnd.n6988 gnd.n408 19.3944
R9925 gnd.n6984 gnd.n408 19.3944
R9926 gnd.n6984 gnd.n375 19.3944
R9927 gnd.n7039 gnd.n375 19.3944
R9928 gnd.n7039 gnd.n376 19.3944
R9929 gnd.n7035 gnd.n376 19.3944
R9930 gnd.n7035 gnd.n7034 19.3944
R9931 gnd.n7034 gnd.n7033 19.3944
R9932 gnd.n7033 gnd.n314 19.3944
R9933 gnd.n7178 gnd.n314 19.3944
R9934 gnd.n7178 gnd.n315 19.3944
R9935 gnd.n7174 gnd.n315 19.3944
R9936 gnd.n7174 gnd.n7173 19.3944
R9937 gnd.n7173 gnd.n7172 19.3944
R9938 gnd.n7172 gnd.n321 19.3944
R9939 gnd.n7168 gnd.n321 19.3944
R9940 gnd.n7168 gnd.n7167 19.3944
R9941 gnd.n7167 gnd.n293 19.3944
R9942 gnd.n7191 gnd.n293 19.3944
R9943 gnd.n7191 gnd.n291 19.3944
R9944 gnd.n7195 gnd.n291 19.3944
R9945 gnd.n7195 gnd.n277 19.3944
R9946 gnd.n7207 gnd.n277 19.3944
R9947 gnd.n7207 gnd.n275 19.3944
R9948 gnd.n7211 gnd.n275 19.3944
R9949 gnd.n7211 gnd.n263 19.3944
R9950 gnd.n7223 gnd.n263 19.3944
R9951 gnd.n7223 gnd.n261 19.3944
R9952 gnd.n7227 gnd.n261 19.3944
R9953 gnd.n7227 gnd.n247 19.3944
R9954 gnd.n7239 gnd.n247 19.3944
R9955 gnd.n7239 gnd.n245 19.3944
R9956 gnd.n7243 gnd.n245 19.3944
R9957 gnd.n7243 gnd.n232 19.3944
R9958 gnd.n7255 gnd.n232 19.3944
R9959 gnd.n7255 gnd.n230 19.3944
R9960 gnd.n7259 gnd.n230 19.3944
R9961 gnd.n7259 gnd.n217 19.3944
R9962 gnd.n7271 gnd.n217 19.3944
R9963 gnd.n7271 gnd.n214 19.3944
R9964 gnd.n7343 gnd.n214 19.3944
R9965 gnd.n7343 gnd.n215 19.3944
R9966 gnd.n7339 gnd.n215 19.3944
R9967 gnd.n7339 gnd.n7338 19.3944
R9968 gnd.n7338 gnd.n7337 19.3944
R9969 gnd.n4999 gnd.n4988 19.3944
R9970 gnd.n4999 gnd.n4997 19.3944
R9971 gnd.n5088 gnd.n4997 19.3944
R9972 gnd.n5088 gnd.n5087 19.3944
R9973 gnd.n5087 gnd.n5006 19.3944
R9974 gnd.n5080 gnd.n5006 19.3944
R9975 gnd.n5080 gnd.n5079 19.3944
R9976 gnd.n5079 gnd.n5016 19.3944
R9977 gnd.n5072 gnd.n5016 19.3944
R9978 gnd.n5072 gnd.n5071 19.3944
R9979 gnd.n5071 gnd.n5029 19.3944
R9980 gnd.n5064 gnd.n5029 19.3944
R9981 gnd.n5064 gnd.n5063 19.3944
R9982 gnd.n5063 gnd.n5039 19.3944
R9983 gnd.n5056 gnd.n5039 19.3944
R9984 gnd.n5056 gnd.n5055 19.3944
R9985 gnd.n4850 gnd.n1212 19.3944
R9986 gnd.n4850 gnd.n4849 19.3944
R9987 gnd.n4849 gnd.n4848 19.3944
R9988 gnd.n4848 gnd.n1216 19.3944
R9989 gnd.n4671 gnd.n1216 19.3944
R9990 gnd.n4671 gnd.n4669 19.3944
R9991 gnd.n4685 gnd.n4669 19.3944
R9992 gnd.n4685 gnd.n4684 19.3944
R9993 gnd.n4684 gnd.n4683 19.3944
R9994 gnd.n4683 gnd.n4680 19.3944
R9995 gnd.n4680 gnd.n4679 19.3944
R9996 gnd.n4679 gnd.n1260 19.3944
R9997 gnd.n4711 gnd.n1260 19.3944
R9998 gnd.n4711 gnd.n1258 19.3944
R9999 gnd.n4725 gnd.n1258 19.3944
R10000 gnd.n4725 gnd.n4724 19.3944
R10001 gnd.n4724 gnd.n4723 19.3944
R10002 gnd.n4723 gnd.n4720 19.3944
R10003 gnd.n4720 gnd.n4719 19.3944
R10004 gnd.n4719 gnd.n1250 19.3944
R10005 gnd.n4750 gnd.n1250 19.3944
R10006 gnd.n4750 gnd.n1248 19.3944
R10007 gnd.n4785 gnd.n1248 19.3944
R10008 gnd.n4785 gnd.n4784 19.3944
R10009 gnd.n4784 gnd.n4783 19.3944
R10010 gnd.n4783 gnd.n4756 19.3944
R10011 gnd.n4779 gnd.n4756 19.3944
R10012 gnd.n4779 gnd.n4778 19.3944
R10013 gnd.n4778 gnd.n4777 19.3944
R10014 gnd.n4777 gnd.n4762 19.3944
R10015 gnd.n4772 gnd.n4762 19.3944
R10016 gnd.n4772 gnd.n4771 19.3944
R10017 gnd.n4771 gnd.n4770 19.3944
R10018 gnd.n4770 gnd.n941 19.3944
R10019 gnd.n6339 gnd.n941 19.3944
R10020 gnd.n6339 gnd.n939 19.3944
R10021 gnd.n6343 gnd.n939 19.3944
R10022 gnd.n6343 gnd.n927 19.3944
R10023 gnd.n6355 gnd.n927 19.3944
R10024 gnd.n6355 gnd.n925 19.3944
R10025 gnd.n6359 gnd.n925 19.3944
R10026 gnd.n6359 gnd.n913 19.3944
R10027 gnd.n6371 gnd.n913 19.3944
R10028 gnd.n6371 gnd.n911 19.3944
R10029 gnd.n6375 gnd.n911 19.3944
R10030 gnd.n6375 gnd.n898 19.3944
R10031 gnd.n6387 gnd.n898 19.3944
R10032 gnd.n6387 gnd.n896 19.3944
R10033 gnd.n6391 gnd.n896 19.3944
R10034 gnd.n6391 gnd.n883 19.3944
R10035 gnd.n6403 gnd.n883 19.3944
R10036 gnd.n6403 gnd.n881 19.3944
R10037 gnd.n6407 gnd.n881 19.3944
R10038 gnd.n6407 gnd.n867 19.3944
R10039 gnd.n6419 gnd.n867 19.3944
R10040 gnd.n6419 gnd.n865 19.3944
R10041 gnd.n6423 gnd.n865 19.3944
R10042 gnd.n6423 gnd.n852 19.3944
R10043 gnd.n6435 gnd.n852 19.3944
R10044 gnd.n6435 gnd.n850 19.3944
R10045 gnd.n6439 gnd.n850 19.3944
R10046 gnd.n6439 gnd.n838 19.3944
R10047 gnd.n6451 gnd.n838 19.3944
R10048 gnd.n6451 gnd.n836 19.3944
R10049 gnd.n6455 gnd.n836 19.3944
R10050 gnd.n6455 gnd.n823 19.3944
R10051 gnd.n6467 gnd.n823 19.3944
R10052 gnd.n6467 gnd.n821 19.3944
R10053 gnd.n6471 gnd.n821 19.3944
R10054 gnd.n6471 gnd.n807 19.3944
R10055 gnd.n6483 gnd.n807 19.3944
R10056 gnd.n6483 gnd.n805 19.3944
R10057 gnd.n6487 gnd.n805 19.3944
R10058 gnd.n6487 gnd.n792 19.3944
R10059 gnd.n6499 gnd.n792 19.3944
R10060 gnd.n6499 gnd.n790 19.3944
R10061 gnd.n6503 gnd.n790 19.3944
R10062 gnd.n6503 gnd.n777 19.3944
R10063 gnd.n6515 gnd.n777 19.3944
R10064 gnd.n6515 gnd.n775 19.3944
R10065 gnd.n6519 gnd.n775 19.3944
R10066 gnd.n6519 gnd.n761 19.3944
R10067 gnd.n6531 gnd.n761 19.3944
R10068 gnd.n6531 gnd.n759 19.3944
R10069 gnd.n6535 gnd.n759 19.3944
R10070 gnd.n6535 gnd.n745 19.3944
R10071 gnd.n6547 gnd.n745 19.3944
R10072 gnd.n6547 gnd.n743 19.3944
R10073 gnd.n6551 gnd.n743 19.3944
R10074 gnd.n6551 gnd.n731 19.3944
R10075 gnd.n6563 gnd.n731 19.3944
R10076 gnd.n6563 gnd.n729 19.3944
R10077 gnd.n6567 gnd.n729 19.3944
R10078 gnd.n6567 gnd.n716 19.3944
R10079 gnd.n6579 gnd.n716 19.3944
R10080 gnd.n6579 gnd.n714 19.3944
R10081 gnd.n6583 gnd.n714 19.3944
R10082 gnd.n6583 gnd.n701 19.3944
R10083 gnd.n6595 gnd.n701 19.3944
R10084 gnd.n6595 gnd.n699 19.3944
R10085 gnd.n6599 gnd.n699 19.3944
R10086 gnd.n6599 gnd.n687 19.3944
R10087 gnd.n6611 gnd.n687 19.3944
R10088 gnd.n6611 gnd.n685 19.3944
R10089 gnd.n6615 gnd.n685 19.3944
R10090 gnd.n6615 gnd.n673 19.3944
R10091 gnd.n6627 gnd.n673 19.3944
R10092 gnd.n6627 gnd.n671 19.3944
R10093 gnd.n6631 gnd.n671 19.3944
R10094 gnd.n6631 gnd.n659 19.3944
R10095 gnd.n6643 gnd.n659 19.3944
R10096 gnd.n6643 gnd.n657 19.3944
R10097 gnd.n6647 gnd.n657 19.3944
R10098 gnd.n6647 gnd.n644 19.3944
R10099 gnd.n6660 gnd.n644 19.3944
R10100 gnd.n6660 gnd.n642 19.3944
R10101 gnd.n6666 gnd.n642 19.3944
R10102 gnd.n6666 gnd.n6665 19.3944
R10103 gnd.n6665 gnd.n614 19.3944
R10104 gnd.n6679 gnd.n614 19.3944
R10105 gnd.n6679 gnd.n612 19.3944
R10106 gnd.n6683 gnd.n612 19.3944
R10107 gnd.n6683 gnd.n610 19.3944
R10108 gnd.n6687 gnd.n610 19.3944
R10109 gnd.n6687 gnd.n608 19.3944
R10110 gnd.n6691 gnd.n608 19.3944
R10111 gnd.n6691 gnd.n606 19.3944
R10112 gnd.n6695 gnd.n606 19.3944
R10113 gnd.n6695 gnd.n604 19.3944
R10114 gnd.n6699 gnd.n604 19.3944
R10115 gnd.n6699 gnd.n602 19.3944
R10116 gnd.n6729 gnd.n602 19.3944
R10117 gnd.n6729 gnd.n600 19.3944
R10118 gnd.n6743 gnd.n600 19.3944
R10119 gnd.n6743 gnd.n6742 19.3944
R10120 gnd.n6742 gnd.n6741 19.3944
R10121 gnd.n6741 gnd.n6738 19.3944
R10122 gnd.n6738 gnd.n6737 19.3944
R10123 gnd.n6737 gnd.n592 19.3944
R10124 gnd.n6768 gnd.n592 19.3944
R10125 gnd.n6768 gnd.n590 19.3944
R10126 gnd.n6774 gnd.n590 19.3944
R10127 gnd.n6774 gnd.n6773 19.3944
R10128 gnd.n6773 gnd.n392 19.3944
R10129 gnd.n7001 gnd.n392 19.3944
R10130 gnd.n7001 gnd.n390 19.3944
R10131 gnd.n7016 gnd.n390 19.3944
R10132 gnd.n7016 gnd.n7015 19.3944
R10133 gnd.n7015 gnd.n7014 19.3944
R10134 gnd.n7014 gnd.n7011 19.3944
R10135 gnd.n7011 gnd.n7010 19.3944
R10136 gnd.n7010 gnd.n346 19.3944
R10137 gnd.n7075 gnd.n346 19.3944
R10138 gnd.n7076 gnd.n7075 19.3944
R10139 gnd.n2237 gnd.n1911 19.3944
R10140 gnd.n2237 gnd.n1912 19.3944
R10141 gnd.n2233 gnd.n1912 19.3944
R10142 gnd.n2233 gnd.n1915 19.3944
R10143 gnd.n2227 gnd.n1915 19.3944
R10144 gnd.n2227 gnd.n2226 19.3944
R10145 gnd.n2226 gnd.n2225 19.3944
R10146 gnd.n2225 gnd.n1922 19.3944
R10147 gnd.n2219 gnd.n1922 19.3944
R10148 gnd.n2219 gnd.n2218 19.3944
R10149 gnd.n2218 gnd.n2217 19.3944
R10150 gnd.n2217 gnd.n1930 19.3944
R10151 gnd.n2211 gnd.n1930 19.3944
R10152 gnd.n2211 gnd.n2210 19.3944
R10153 gnd.n2210 gnd.n2209 19.3944
R10154 gnd.n2209 gnd.n1938 19.3944
R10155 gnd.n2203 gnd.n1938 19.3944
R10156 gnd.n2203 gnd.n2202 19.3944
R10157 gnd.n2202 gnd.n2201 19.3944
R10158 gnd.n2201 gnd.n1946 19.3944
R10159 gnd.n2195 gnd.n1946 19.3944
R10160 gnd.n2195 gnd.n2194 19.3944
R10161 gnd.n2194 gnd.n2193 19.3944
R10162 gnd.n2193 gnd.n1954 19.3944
R10163 gnd.n2187 gnd.n1954 19.3944
R10164 gnd.n2187 gnd.n2186 19.3944
R10165 gnd.n2186 gnd.n2185 19.3944
R10166 gnd.n2185 gnd.n1962 19.3944
R10167 gnd.n2179 gnd.n1962 19.3944
R10168 gnd.n2179 gnd.n2178 19.3944
R10169 gnd.n2178 gnd.n2177 19.3944
R10170 gnd.n2177 gnd.n1970 19.3944
R10171 gnd.n2171 gnd.n1970 19.3944
R10172 gnd.n2171 gnd.n2170 19.3944
R10173 gnd.n2170 gnd.n2169 19.3944
R10174 gnd.n2169 gnd.n1978 19.3944
R10175 gnd.n2163 gnd.n1978 19.3944
R10176 gnd.n2163 gnd.n2162 19.3944
R10177 gnd.n2162 gnd.n2161 19.3944
R10178 gnd.n2161 gnd.n1986 19.3944
R10179 gnd.n2155 gnd.n1986 19.3944
R10180 gnd.n2155 gnd.n2154 19.3944
R10181 gnd.n2154 gnd.n2153 19.3944
R10182 gnd.n2153 gnd.n1994 19.3944
R10183 gnd.n2147 gnd.n1994 19.3944
R10184 gnd.n2147 gnd.n2146 19.3944
R10185 gnd.n2146 gnd.n2145 19.3944
R10186 gnd.n2145 gnd.n2002 19.3944
R10187 gnd.n2139 gnd.n2002 19.3944
R10188 gnd.n2139 gnd.n2138 19.3944
R10189 gnd.n2138 gnd.n2137 19.3944
R10190 gnd.n2137 gnd.n2010 19.3944
R10191 gnd.n2131 gnd.n2010 19.3944
R10192 gnd.n2131 gnd.n2130 19.3944
R10193 gnd.n2130 gnd.n2129 19.3944
R10194 gnd.n2129 gnd.n2018 19.3944
R10195 gnd.n2123 gnd.n2018 19.3944
R10196 gnd.n2123 gnd.n2122 19.3944
R10197 gnd.n2122 gnd.n2121 19.3944
R10198 gnd.n2121 gnd.n2026 19.3944
R10199 gnd.n2115 gnd.n2026 19.3944
R10200 gnd.n2115 gnd.n2114 19.3944
R10201 gnd.n2114 gnd.n2113 19.3944
R10202 gnd.n2113 gnd.n2034 19.3944
R10203 gnd.n2107 gnd.n2034 19.3944
R10204 gnd.n2107 gnd.n2106 19.3944
R10205 gnd.n2106 gnd.n2105 19.3944
R10206 gnd.n2105 gnd.n2042 19.3944
R10207 gnd.n2099 gnd.n2042 19.3944
R10208 gnd.n2099 gnd.n2098 19.3944
R10209 gnd.n2098 gnd.n2097 19.3944
R10210 gnd.n2097 gnd.n2050 19.3944
R10211 gnd.n2091 gnd.n2050 19.3944
R10212 gnd.n2091 gnd.n2090 19.3944
R10213 gnd.n2090 gnd.n2089 19.3944
R10214 gnd.n2089 gnd.n2058 19.3944
R10215 gnd.n2083 gnd.n2058 19.3944
R10216 gnd.n2083 gnd.n2082 19.3944
R10217 gnd.n2082 gnd.n2081 19.3944
R10218 gnd.n2081 gnd.n2066 19.3944
R10219 gnd.n2075 gnd.n2066 19.3944
R10220 gnd.n2075 gnd.n2074 19.3944
R10221 gnd.n2074 gnd.n344 19.3944
R10222 gnd.n7079 gnd.n344 19.3944
R10223 gnd.n2551 gnd.n1603 19.3944
R10224 gnd.n2547 gnd.n1603 19.3944
R10225 gnd.n2547 gnd.n1605 19.3944
R10226 gnd.n2541 gnd.n1605 19.3944
R10227 gnd.n2541 gnd.n2540 19.3944
R10228 gnd.n2540 gnd.n2539 19.3944
R10229 gnd.n2539 gnd.n1612 19.3944
R10230 gnd.n2533 gnd.n1612 19.3944
R10231 gnd.n2533 gnd.n2532 19.3944
R10232 gnd.n2532 gnd.n2531 19.3944
R10233 gnd.n2531 gnd.n1620 19.3944
R10234 gnd.n2525 gnd.n1620 19.3944
R10235 gnd.n2525 gnd.n2524 19.3944
R10236 gnd.n2524 gnd.n2523 19.3944
R10237 gnd.n2523 gnd.n1628 19.3944
R10238 gnd.n2517 gnd.n1628 19.3944
R10239 gnd.n2517 gnd.n2516 19.3944
R10240 gnd.n2516 gnd.n2515 19.3944
R10241 gnd.n2515 gnd.n1636 19.3944
R10242 gnd.n2509 gnd.n1636 19.3944
R10243 gnd.n2509 gnd.n2508 19.3944
R10244 gnd.n2508 gnd.n2507 19.3944
R10245 gnd.n2507 gnd.n1644 19.3944
R10246 gnd.n2501 gnd.n1644 19.3944
R10247 gnd.n2501 gnd.n2500 19.3944
R10248 gnd.n2500 gnd.n2499 19.3944
R10249 gnd.n2499 gnd.n1652 19.3944
R10250 gnd.n2493 gnd.n1652 19.3944
R10251 gnd.n2493 gnd.n2492 19.3944
R10252 gnd.n2492 gnd.n2491 19.3944
R10253 gnd.n2491 gnd.n1660 19.3944
R10254 gnd.n2485 gnd.n1660 19.3944
R10255 gnd.n2485 gnd.n2484 19.3944
R10256 gnd.n2484 gnd.n2483 19.3944
R10257 gnd.n2483 gnd.n1668 19.3944
R10258 gnd.n2477 gnd.n1668 19.3944
R10259 gnd.n2477 gnd.n2476 19.3944
R10260 gnd.n2476 gnd.n2475 19.3944
R10261 gnd.n2475 gnd.n1676 19.3944
R10262 gnd.n2469 gnd.n1676 19.3944
R10263 gnd.n2469 gnd.n2468 19.3944
R10264 gnd.n2468 gnd.n2467 19.3944
R10265 gnd.n2467 gnd.n1684 19.3944
R10266 gnd.n2461 gnd.n1684 19.3944
R10267 gnd.n2461 gnd.n2460 19.3944
R10268 gnd.n2460 gnd.n2459 19.3944
R10269 gnd.n2459 gnd.n1692 19.3944
R10270 gnd.n2453 gnd.n1692 19.3944
R10271 gnd.n2453 gnd.n2452 19.3944
R10272 gnd.n2452 gnd.n2451 19.3944
R10273 gnd.n2451 gnd.n1700 19.3944
R10274 gnd.n2445 gnd.n1700 19.3944
R10275 gnd.n2445 gnd.n2444 19.3944
R10276 gnd.n2444 gnd.n2443 19.3944
R10277 gnd.n2443 gnd.n1708 19.3944
R10278 gnd.n2437 gnd.n1708 19.3944
R10279 gnd.n2437 gnd.n2436 19.3944
R10280 gnd.n2436 gnd.n2435 19.3944
R10281 gnd.n2435 gnd.n1716 19.3944
R10282 gnd.n2429 gnd.n1716 19.3944
R10283 gnd.n2429 gnd.n2428 19.3944
R10284 gnd.n2428 gnd.n2427 19.3944
R10285 gnd.n2427 gnd.n1724 19.3944
R10286 gnd.n2421 gnd.n1724 19.3944
R10287 gnd.n2421 gnd.n2420 19.3944
R10288 gnd.n2420 gnd.n2419 19.3944
R10289 gnd.n2419 gnd.n1732 19.3944
R10290 gnd.n2413 gnd.n1732 19.3944
R10291 gnd.n2413 gnd.n2412 19.3944
R10292 gnd.n2412 gnd.n2411 19.3944
R10293 gnd.n2411 gnd.n1740 19.3944
R10294 gnd.n2405 gnd.n1740 19.3944
R10295 gnd.n2405 gnd.n2404 19.3944
R10296 gnd.n2404 gnd.n2403 19.3944
R10297 gnd.n2403 gnd.n1748 19.3944
R10298 gnd.n2397 gnd.n1748 19.3944
R10299 gnd.n2397 gnd.n2396 19.3944
R10300 gnd.n2396 gnd.n2395 19.3944
R10301 gnd.n2395 gnd.n1756 19.3944
R10302 gnd.n2389 gnd.n1756 19.3944
R10303 gnd.n2389 gnd.n2388 19.3944
R10304 gnd.n2388 gnd.n2387 19.3944
R10305 gnd.n2387 gnd.n1764 19.3944
R10306 gnd.n2381 gnd.n1764 19.3944
R10307 gnd.n2381 gnd.n2380 19.3944
R10308 gnd.n2380 gnd.n2379 19.3944
R10309 gnd.n2379 gnd.n1772 19.3944
R10310 gnd.n2373 gnd.n1772 19.3944
R10311 gnd.n2373 gnd.n2372 19.3944
R10312 gnd.n2372 gnd.n2371 19.3944
R10313 gnd.n2371 gnd.n1780 19.3944
R10314 gnd.n2365 gnd.n1780 19.3944
R10315 gnd.n2365 gnd.n2364 19.3944
R10316 gnd.n2364 gnd.n2363 19.3944
R10317 gnd.n2363 gnd.n1788 19.3944
R10318 gnd.n2357 gnd.n1788 19.3944
R10319 gnd.n2357 gnd.n2356 19.3944
R10320 gnd.n2356 gnd.n2355 19.3944
R10321 gnd.n2355 gnd.n1796 19.3944
R10322 gnd.n2349 gnd.n1796 19.3944
R10323 gnd.n2349 gnd.n2348 19.3944
R10324 gnd.n2348 gnd.n2347 19.3944
R10325 gnd.n2347 gnd.n1804 19.3944
R10326 gnd.n2341 gnd.n1804 19.3944
R10327 gnd.n2341 gnd.n2340 19.3944
R10328 gnd.n2340 gnd.n2339 19.3944
R10329 gnd.n2339 gnd.n1812 19.3944
R10330 gnd.n2333 gnd.n1812 19.3944
R10331 gnd.n2333 gnd.n2332 19.3944
R10332 gnd.n2332 gnd.n2331 19.3944
R10333 gnd.n2331 gnd.n1820 19.3944
R10334 gnd.n2325 gnd.n1820 19.3944
R10335 gnd.n2325 gnd.n2324 19.3944
R10336 gnd.n2324 gnd.n2323 19.3944
R10337 gnd.n2323 gnd.n1828 19.3944
R10338 gnd.n2317 gnd.n1828 19.3944
R10339 gnd.n2317 gnd.n2316 19.3944
R10340 gnd.n2316 gnd.n2315 19.3944
R10341 gnd.n2315 gnd.n1836 19.3944
R10342 gnd.n2309 gnd.n1836 19.3944
R10343 gnd.n2309 gnd.n2308 19.3944
R10344 gnd.n2308 gnd.n2307 19.3944
R10345 gnd.n2307 gnd.n1844 19.3944
R10346 gnd.n2301 gnd.n1844 19.3944
R10347 gnd.n2301 gnd.n2300 19.3944
R10348 gnd.n2300 gnd.n2299 19.3944
R10349 gnd.n2299 gnd.n1852 19.3944
R10350 gnd.n2293 gnd.n1852 19.3944
R10351 gnd.n2293 gnd.n2292 19.3944
R10352 gnd.n2292 gnd.n2291 19.3944
R10353 gnd.n2291 gnd.n1860 19.3944
R10354 gnd.n2285 gnd.n1860 19.3944
R10355 gnd.n2285 gnd.n2284 19.3944
R10356 gnd.n2284 gnd.n2283 19.3944
R10357 gnd.n2283 gnd.n1868 19.3944
R10358 gnd.n2277 gnd.n1868 19.3944
R10359 gnd.n2277 gnd.n2276 19.3944
R10360 gnd.n2276 gnd.n2275 19.3944
R10361 gnd.n2275 gnd.n1876 19.3944
R10362 gnd.n2269 gnd.n1876 19.3944
R10363 gnd.n2269 gnd.n2268 19.3944
R10364 gnd.n2268 gnd.n2267 19.3944
R10365 gnd.n2267 gnd.n1884 19.3944
R10366 gnd.n2261 gnd.n1884 19.3944
R10367 gnd.n2261 gnd.n2260 19.3944
R10368 gnd.n2260 gnd.n2259 19.3944
R10369 gnd.n2259 gnd.n1892 19.3944
R10370 gnd.n2253 gnd.n1892 19.3944
R10371 gnd.n2253 gnd.n2252 19.3944
R10372 gnd.n2252 gnd.n2251 19.3944
R10373 gnd.n2251 gnd.n1900 19.3944
R10374 gnd.n2245 gnd.n1900 19.3944
R10375 gnd.n2245 gnd.n2244 19.3944
R10376 gnd.n2244 gnd.n2243 19.3944
R10377 gnd.n6909 gnd.n487 19.3944
R10378 gnd.n6904 gnd.n487 19.3944
R10379 gnd.n6904 gnd.n6903 19.3944
R10380 gnd.n6903 gnd.n6902 19.3944
R10381 gnd.n6902 gnd.n6899 19.3944
R10382 gnd.n6899 gnd.n6898 19.3944
R10383 gnd.n6898 gnd.n6895 19.3944
R10384 gnd.n6895 gnd.n6894 19.3944
R10385 gnd.n6894 gnd.n6891 19.3944
R10386 gnd.n6891 gnd.n6890 19.3944
R10387 gnd.n6890 gnd.n6887 19.3944
R10388 gnd.n6887 gnd.n6886 19.3944
R10389 gnd.n6886 gnd.n6883 19.3944
R10390 gnd.n6883 gnd.n6882 19.3944
R10391 gnd.n6882 gnd.n6879 19.3944
R10392 gnd.n6877 gnd.n6874 19.3944
R10393 gnd.n6874 gnd.n6873 19.3944
R10394 gnd.n6873 gnd.n6870 19.3944
R10395 gnd.n6870 gnd.n6869 19.3944
R10396 gnd.n6869 gnd.n6866 19.3944
R10397 gnd.n6866 gnd.n6865 19.3944
R10398 gnd.n6865 gnd.n6862 19.3944
R10399 gnd.n6862 gnd.n6861 19.3944
R10400 gnd.n6861 gnd.n6858 19.3944
R10401 gnd.n6858 gnd.n6857 19.3944
R10402 gnd.n6857 gnd.n6854 19.3944
R10403 gnd.n6854 gnd.n6853 19.3944
R10404 gnd.n6853 gnd.n6850 19.3944
R10405 gnd.n6850 gnd.n6849 19.3944
R10406 gnd.n6849 gnd.n6846 19.3944
R10407 gnd.n6846 gnd.n6845 19.3944
R10408 gnd.n6845 gnd.n6842 19.3944
R10409 gnd.n6842 gnd.n6841 19.3944
R10410 gnd.n6703 gnd.n563 19.3944
R10411 gnd.n6708 gnd.n6703 19.3944
R10412 gnd.n6709 gnd.n6708 19.3944
R10413 gnd.n6712 gnd.n6709 19.3944
R10414 gnd.n6712 gnd.n6701 19.3944
R10415 gnd.n6723 gnd.n6701 19.3944
R10416 gnd.n6723 gnd.n6722 19.3944
R10417 gnd.n6722 gnd.n6721 19.3944
R10418 gnd.n6721 gnd.n596 19.3944
R10419 gnd.n6748 gnd.n596 19.3944
R10420 gnd.n6749 gnd.n6748 19.3944
R10421 gnd.n6752 gnd.n6749 19.3944
R10422 gnd.n6752 gnd.n594 19.3944
R10423 gnd.n6762 gnd.n594 19.3944
R10424 gnd.n6762 gnd.n6761 19.3944
R10425 gnd.n6761 gnd.n6760 19.3944
R10426 gnd.n6760 gnd.n587 19.3944
R10427 gnd.n6779 gnd.n587 19.3944
R10428 gnd.n6779 gnd.n585 19.3944
R10429 gnd.n6796 gnd.n585 19.3944
R10430 gnd.n6796 gnd.n6795 19.3944
R10431 gnd.n6795 gnd.n6794 19.3944
R10432 gnd.n6794 gnd.n6793 19.3944
R10433 gnd.n6793 gnd.n6792 19.3944
R10434 gnd.n6792 gnd.n6789 19.3944
R10435 gnd.n6789 gnd.n357 19.3944
R10436 gnd.n7053 gnd.n357 19.3944
R10437 gnd.n7054 gnd.n7053 19.3944
R10438 gnd.n7054 gnd.n355 19.3944
R10439 gnd.n7060 gnd.n355 19.3944
R10440 gnd.n7060 gnd.n7059 19.3944
R10441 gnd.n7059 gnd.n334 19.3944
R10442 gnd.n7090 gnd.n334 19.3944
R10443 gnd.n7090 gnd.n332 19.3944
R10444 gnd.n7159 gnd.n332 19.3944
R10445 gnd.n7159 gnd.n7158 19.3944
R10446 gnd.n7158 gnd.n7157 19.3944
R10447 gnd.n7157 gnd.n7155 19.3944
R10448 gnd.n7155 gnd.n7154 19.3944
R10449 gnd.n7154 gnd.n7152 19.3944
R10450 gnd.n7152 gnd.n7151 19.3944
R10451 gnd.n7151 gnd.n7149 19.3944
R10452 gnd.n7149 gnd.n7148 19.3944
R10453 gnd.n7148 gnd.n7146 19.3944
R10454 gnd.n7146 gnd.n7145 19.3944
R10455 gnd.n7145 gnd.n7143 19.3944
R10456 gnd.n7143 gnd.n7142 19.3944
R10457 gnd.n7142 gnd.n7140 19.3944
R10458 gnd.n7140 gnd.n7139 19.3944
R10459 gnd.n7139 gnd.n7137 19.3944
R10460 gnd.n7137 gnd.n7136 19.3944
R10461 gnd.n7136 gnd.n7134 19.3944
R10462 gnd.n7134 gnd.n7133 19.3944
R10463 gnd.n7133 gnd.n7131 19.3944
R10464 gnd.n7131 gnd.n7130 19.3944
R10465 gnd.n7130 gnd.n7128 19.3944
R10466 gnd.n7128 gnd.n7127 19.3944
R10467 gnd.n7127 gnd.n7125 19.3944
R10468 gnd.n7125 gnd.n7124 19.3944
R10469 gnd.n7124 gnd.n7122 19.3944
R10470 gnd.n7122 gnd.n7121 19.3944
R10471 gnd.n7121 gnd.n200 19.3944
R10472 gnd.n7356 gnd.n200 19.3944
R10473 gnd.n7357 gnd.n7356 19.3944
R10474 gnd.n7395 gnd.n161 19.3944
R10475 gnd.n7390 gnd.n161 19.3944
R10476 gnd.n7390 gnd.n7389 19.3944
R10477 gnd.n7389 gnd.n7388 19.3944
R10478 gnd.n7388 gnd.n168 19.3944
R10479 gnd.n7383 gnd.n168 19.3944
R10480 gnd.n7383 gnd.n7382 19.3944
R10481 gnd.n7382 gnd.n7381 19.3944
R10482 gnd.n7381 gnd.n175 19.3944
R10483 gnd.n7376 gnd.n175 19.3944
R10484 gnd.n7376 gnd.n7375 19.3944
R10485 gnd.n7375 gnd.n7374 19.3944
R10486 gnd.n7374 gnd.n182 19.3944
R10487 gnd.n7369 gnd.n182 19.3944
R10488 gnd.n7369 gnd.n7368 19.3944
R10489 gnd.n7368 gnd.n7367 19.3944
R10490 gnd.n7367 gnd.n189 19.3944
R10491 gnd.n7362 gnd.n189 19.3944
R10492 gnd.n7428 gnd.n7427 19.3944
R10493 gnd.n7427 gnd.n7426 19.3944
R10494 gnd.n7426 gnd.n133 19.3944
R10495 gnd.n7421 gnd.n133 19.3944
R10496 gnd.n7421 gnd.n7420 19.3944
R10497 gnd.n7420 gnd.n7419 19.3944
R10498 gnd.n7419 gnd.n140 19.3944
R10499 gnd.n7414 gnd.n140 19.3944
R10500 gnd.n7414 gnd.n7413 19.3944
R10501 gnd.n7413 gnd.n7412 19.3944
R10502 gnd.n7412 gnd.n147 19.3944
R10503 gnd.n7407 gnd.n147 19.3944
R10504 gnd.n7407 gnd.n7406 19.3944
R10505 gnd.n7406 gnd.n7405 19.3944
R10506 gnd.n7405 gnd.n154 19.3944
R10507 gnd.n7400 gnd.n154 19.3944
R10508 gnd.n7400 gnd.n7399 19.3944
R10509 gnd.n6913 gnd.n485 19.3944
R10510 gnd.n6913 gnd.n469 19.3944
R10511 gnd.n6925 gnd.n469 19.3944
R10512 gnd.n6925 gnd.n467 19.3944
R10513 gnd.n6929 gnd.n467 19.3944
R10514 gnd.n6929 gnd.n452 19.3944
R10515 gnd.n6941 gnd.n452 19.3944
R10516 gnd.n6941 gnd.n450 19.3944
R10517 gnd.n6945 gnd.n450 19.3944
R10518 gnd.n6945 gnd.n435 19.3944
R10519 gnd.n6957 gnd.n435 19.3944
R10520 gnd.n6957 gnd.n433 19.3944
R10521 gnd.n6961 gnd.n433 19.3944
R10522 gnd.n6961 gnd.n418 19.3944
R10523 gnd.n6973 gnd.n418 19.3944
R10524 gnd.n6973 gnd.n416 19.3944
R10525 gnd.n6977 gnd.n416 19.3944
R10526 gnd.n6977 gnd.n399 19.3944
R10527 gnd.n6992 gnd.n399 19.3944
R10528 gnd.n6992 gnd.n397 19.3944
R10529 gnd.n6996 gnd.n397 19.3944
R10530 gnd.n6996 gnd.n367 19.3944
R10531 gnd.n7043 gnd.n367 19.3944
R10532 gnd.n7043 gnd.n365 19.3944
R10533 gnd.n7047 gnd.n365 19.3944
R10534 gnd.n7048 gnd.n7047 19.3944
R10535 gnd.n7048 gnd.n305 19.3944
R10536 gnd.n7183 gnd.n7182 19.3944
R10537 gnd.n338 gnd.n337 19.3944
R10538 gnd.n7086 gnd.n7085 19.3944
R10539 gnd.n328 gnd.n327 19.3944
R10540 gnd.n7163 gnd.n298 19.3944
R10541 gnd.n7187 gnd.n298 19.3944
R10542 gnd.n7187 gnd.n284 19.3944
R10543 gnd.n7199 gnd.n284 19.3944
R10544 gnd.n7199 gnd.n282 19.3944
R10545 gnd.n7203 gnd.n282 19.3944
R10546 gnd.n7203 gnd.n270 19.3944
R10547 gnd.n7215 gnd.n270 19.3944
R10548 gnd.n7215 gnd.n268 19.3944
R10549 gnd.n7219 gnd.n268 19.3944
R10550 gnd.n7219 gnd.n254 19.3944
R10551 gnd.n7231 gnd.n254 19.3944
R10552 gnd.n7231 gnd.n252 19.3944
R10553 gnd.n7235 gnd.n252 19.3944
R10554 gnd.n7235 gnd.n240 19.3944
R10555 gnd.n7247 gnd.n240 19.3944
R10556 gnd.n7247 gnd.n238 19.3944
R10557 gnd.n7251 gnd.n238 19.3944
R10558 gnd.n7251 gnd.n223 19.3944
R10559 gnd.n7263 gnd.n223 19.3944
R10560 gnd.n7263 gnd.n221 19.3944
R10561 gnd.n7267 gnd.n221 19.3944
R10562 gnd.n7267 gnd.n207 19.3944
R10563 gnd.n7347 gnd.n207 19.3944
R10564 gnd.n7347 gnd.n205 19.3944
R10565 gnd.n7351 gnd.n205 19.3944
R10566 gnd.n7351 gnd.n128 19.3944
R10567 gnd.n7431 gnd.n128 19.3944
R10568 gnd.n4477 gnd.n4476 19.3944
R10569 gnd.n4476 gnd.n4287 19.3944
R10570 gnd.n4471 gnd.n4287 19.3944
R10571 gnd.n4471 gnd.n4470 19.3944
R10572 gnd.n4470 gnd.n4292 19.3944
R10573 gnd.n4465 gnd.n4292 19.3944
R10574 gnd.n4465 gnd.n4464 19.3944
R10575 gnd.n4464 gnd.n4463 19.3944
R10576 gnd.n4463 gnd.n4298 19.3944
R10577 gnd.n4457 gnd.n4298 19.3944
R10578 gnd.n4457 gnd.n4456 19.3944
R10579 gnd.n4456 gnd.n4455 19.3944
R10580 gnd.n4455 gnd.n4304 19.3944
R10581 gnd.n4449 gnd.n4304 19.3944
R10582 gnd.n4449 gnd.n4448 19.3944
R10583 gnd.n4448 gnd.n4447 19.3944
R10584 gnd.n4447 gnd.n4310 19.3944
R10585 gnd.n4441 gnd.n4440 19.3944
R10586 gnd.n4440 gnd.n4439 19.3944
R10587 gnd.n4439 gnd.n4319 19.3944
R10588 gnd.n4433 gnd.n4319 19.3944
R10589 gnd.n4433 gnd.n4432 19.3944
R10590 gnd.n4432 gnd.n4431 19.3944
R10591 gnd.n4431 gnd.n4325 19.3944
R10592 gnd.n4425 gnd.n4325 19.3944
R10593 gnd.n4425 gnd.n4424 19.3944
R10594 gnd.n4424 gnd.n4423 19.3944
R10595 gnd.n4423 gnd.n4331 19.3944
R10596 gnd.n4417 gnd.n4331 19.3944
R10597 gnd.n4417 gnd.n4416 19.3944
R10598 gnd.n4416 gnd.n4415 19.3944
R10599 gnd.n4415 gnd.n4337 19.3944
R10600 gnd.n4409 gnd.n4337 19.3944
R10601 gnd.n4409 gnd.n4408 19.3944
R10602 gnd.n4408 gnd.n4407 19.3944
R10603 gnd.n4484 gnd.n1397 19.3944
R10604 gnd.n4488 gnd.n1397 19.3944
R10605 gnd.n4488 gnd.n1384 19.3944
R10606 gnd.n4500 gnd.n1384 19.3944
R10607 gnd.n4500 gnd.n1382 19.3944
R10608 gnd.n4504 gnd.n1382 19.3944
R10609 gnd.n4504 gnd.n1367 19.3944
R10610 gnd.n4516 gnd.n1367 19.3944
R10611 gnd.n4516 gnd.n1365 19.3944
R10612 gnd.n4520 gnd.n1365 19.3944
R10613 gnd.n4520 gnd.n1352 19.3944
R10614 gnd.n4532 gnd.n1352 19.3944
R10615 gnd.n4532 gnd.n1350 19.3944
R10616 gnd.n4536 gnd.n1350 19.3944
R10617 gnd.n4536 gnd.n1335 19.3944
R10618 gnd.n4548 gnd.n1335 19.3944
R10619 gnd.n4548 gnd.n1333 19.3944
R10620 gnd.n4560 gnd.n1333 19.3944
R10621 gnd.n4560 gnd.n4559 19.3944
R10622 gnd.n4559 gnd.n4558 19.3944
R10623 gnd.n4558 gnd.n4557 19.3944
R10624 gnd.n4557 gnd.n1299 19.3944
R10625 gnd.n4600 gnd.n1299 19.3944
R10626 gnd.n4600 gnd.n4599 19.3944
R10627 gnd.n4599 gnd.n4598 19.3944
R10628 gnd.n4598 gnd.n1308 19.3944
R10629 gnd.n1308 gnd.n1307 19.3944
R10630 gnd.n1307 gnd.n1190 19.3944
R10631 gnd.n4874 gnd.n1190 19.3944
R10632 gnd.n4874 gnd.n4873 19.3944
R10633 gnd.n4873 gnd.n4872 19.3944
R10634 gnd.n4872 gnd.n1194 19.3944
R10635 gnd.n4860 gnd.n1194 19.3944
R10636 gnd.n4860 gnd.n4859 19.3944
R10637 gnd.n4859 gnd.n4858 19.3944
R10638 gnd.n4858 gnd.n1168 19.3944
R10639 gnd.n4886 gnd.n1168 19.3944
R10640 gnd.n4886 gnd.n1166 19.3944
R10641 gnd.n4890 gnd.n1166 19.3944
R10642 gnd.n4890 gnd.n1152 19.3944
R10643 gnd.n4902 gnd.n1152 19.3944
R10644 gnd.n4902 gnd.n1150 19.3944
R10645 gnd.n4906 gnd.n1150 19.3944
R10646 gnd.n4906 gnd.n1134 19.3944
R10647 gnd.n4918 gnd.n1134 19.3944
R10648 gnd.n4918 gnd.n1132 19.3944
R10649 gnd.n4922 gnd.n1132 19.3944
R10650 gnd.n4922 gnd.n1118 19.3944
R10651 gnd.n4934 gnd.n1118 19.3944
R10652 gnd.n4934 gnd.n1116 19.3944
R10653 gnd.n4938 gnd.n1116 19.3944
R10654 gnd.n4938 gnd.n1100 19.3944
R10655 gnd.n4950 gnd.n1100 19.3944
R10656 gnd.n4950 gnd.n1098 19.3944
R10657 gnd.n4954 gnd.n1098 19.3944
R10658 gnd.n4954 gnd.n1084 19.3944
R10659 gnd.n4966 gnd.n1084 19.3944
R10660 gnd.n4966 gnd.n1082 19.3944
R10661 gnd.n4970 gnd.n1082 19.3944
R10662 gnd.n4970 gnd.n1065 19.3944
R10663 gnd.n4984 gnd.n1065 19.3944
R10664 gnd.n4984 gnd.n1063 19.3944
R10665 gnd.n6223 gnd.n1063 19.3944
R10666 gnd.n6223 gnd.n6222 19.3944
R10667 gnd.n4192 gnd.n4191 19.3944
R10668 gnd.n4197 gnd.n4192 19.3944
R10669 gnd.n4197 gnd.n4189 19.3944
R10670 gnd.n4201 gnd.n4189 19.3944
R10671 gnd.n4201 gnd.n4187 19.3944
R10672 gnd.n4207 gnd.n4187 19.3944
R10673 gnd.n4207 gnd.n4185 19.3944
R10674 gnd.n4211 gnd.n4185 19.3944
R10675 gnd.n4211 gnd.n4183 19.3944
R10676 gnd.n4217 gnd.n4183 19.3944
R10677 gnd.n4217 gnd.n4181 19.3944
R10678 gnd.n4221 gnd.n4181 19.3944
R10679 gnd.n4221 gnd.n4179 19.3944
R10680 gnd.n4227 gnd.n4179 19.3944
R10681 gnd.n4227 gnd.n4177 19.3944
R10682 gnd.n4231 gnd.n4177 19.3944
R10683 gnd.n4282 gnd.n4171 19.3944
R10684 gnd.n4282 gnd.n4281 19.3944
R10685 gnd.n4281 gnd.n4280 19.3944
R10686 gnd.n4280 gnd.n4278 19.3944
R10687 gnd.n4278 gnd.n4277 19.3944
R10688 gnd.n4277 gnd.n4275 19.3944
R10689 gnd.n4275 gnd.n4274 19.3944
R10690 gnd.n4274 gnd.n4272 19.3944
R10691 gnd.n4272 gnd.n4271 19.3944
R10692 gnd.n4271 gnd.n4269 19.3944
R10693 gnd.n4269 gnd.n4268 19.3944
R10694 gnd.n4268 gnd.n4266 19.3944
R10695 gnd.n4266 gnd.n4265 19.3944
R10696 gnd.n4265 gnd.n4263 19.3944
R10697 gnd.n4263 gnd.n4262 19.3944
R10698 gnd.n4262 gnd.n4260 19.3944
R10699 gnd.n4260 gnd.n4259 19.3944
R10700 gnd.n4259 gnd.n4257 19.3944
R10701 gnd.n4257 gnd.n1318 19.3944
R10702 gnd.n4574 gnd.n1318 19.3944
R10703 gnd.n4574 gnd.n1316 19.3944
R10704 gnd.n4583 gnd.n1316 19.3944
R10705 gnd.n4583 gnd.n4582 19.3944
R10706 gnd.n4582 gnd.n4581 19.3944
R10707 gnd.n4581 gnd.n1283 19.3944
R10708 gnd.n4613 gnd.n1283 19.3944
R10709 gnd.n4613 gnd.n1281 19.3944
R10710 gnd.n4627 gnd.n1281 19.3944
R10711 gnd.n4627 gnd.n4626 19.3944
R10712 gnd.n4626 gnd.n4625 19.3944
R10713 gnd.n4625 gnd.n4623 19.3944
R10714 gnd.n4623 gnd.n4622 19.3944
R10715 gnd.n4622 gnd.n1271 19.3944
R10716 gnd.n4647 gnd.n1271 19.3944
R10717 gnd.n4647 gnd.n1269 19.3944
R10718 gnd.n4651 gnd.n1269 19.3944
R10719 gnd.n4651 gnd.n1219 19.3944
R10720 gnd.n4842 gnd.n1219 19.3944
R10721 gnd.n4842 gnd.n1220 19.3944
R10722 gnd.n4838 gnd.n1220 19.3944
R10723 gnd.n4838 gnd.n4837 19.3944
R10724 gnd.n4837 gnd.n4836 19.3944
R10725 gnd.n4836 gnd.n1225 19.3944
R10726 gnd.n4832 gnd.n1225 19.3944
R10727 gnd.n4832 gnd.n4831 19.3944
R10728 gnd.n4831 gnd.n4830 19.3944
R10729 gnd.n4830 gnd.n1229 19.3944
R10730 gnd.n4826 gnd.n1229 19.3944
R10731 gnd.n4826 gnd.n4825 19.3944
R10732 gnd.n4825 gnd.n4824 19.3944
R10733 gnd.n4824 gnd.n1233 19.3944
R10734 gnd.n4820 gnd.n1233 19.3944
R10735 gnd.n4820 gnd.n4819 19.3944
R10736 gnd.n4819 gnd.n4818 19.3944
R10737 gnd.n4818 gnd.n1237 19.3944
R10738 gnd.n4814 gnd.n1237 19.3944
R10739 gnd.n4814 gnd.n4813 19.3944
R10740 gnd.n4813 gnd.n4812 19.3944
R10741 gnd.n4812 gnd.n1241 19.3944
R10742 gnd.n4808 gnd.n1241 19.3944
R10743 gnd.n4808 gnd.n4807 19.3944
R10744 gnd.n4807 gnd.n4806 19.3944
R10745 gnd.n4806 gnd.n4803 19.3944
R10746 gnd.n4803 gnd.n981 19.3944
R10747 gnd.n4398 gnd.n4397 19.3944
R10748 gnd.n4397 gnd.n4396 19.3944
R10749 gnd.n4396 gnd.n4395 19.3944
R10750 gnd.n4395 gnd.n4393 19.3944
R10751 gnd.n4393 gnd.n4392 19.3944
R10752 gnd.n4392 gnd.n4390 19.3944
R10753 gnd.n4390 gnd.n4389 19.3944
R10754 gnd.n4389 gnd.n4387 19.3944
R10755 gnd.n4387 gnd.n4386 19.3944
R10756 gnd.n4386 gnd.n4384 19.3944
R10757 gnd.n4384 gnd.n4383 19.3944
R10758 gnd.n4383 gnd.n4381 19.3944
R10759 gnd.n4381 gnd.n4380 19.3944
R10760 gnd.n4380 gnd.n4378 19.3944
R10761 gnd.n4378 gnd.n4377 19.3944
R10762 gnd.n4377 gnd.n4375 19.3944
R10763 gnd.n4375 gnd.n4374 19.3944
R10764 gnd.n4374 gnd.n4372 19.3944
R10765 gnd.n4372 gnd.n4371 19.3944
R10766 gnd.n4371 gnd.n4369 19.3944
R10767 gnd.n4369 gnd.n1312 19.3944
R10768 gnd.n4587 gnd.n1312 19.3944
R10769 gnd.n4588 gnd.n4587 19.3944
R10770 gnd.n4588 gnd.n1310 19.3944
R10771 gnd.n4594 gnd.n1310 19.3944
R10772 gnd.n4594 gnd.n4593 19.3944
R10773 gnd.n4593 gnd.n1277 19.3944
R10774 gnd.n4631 gnd.n1277 19.3944
R10775 gnd.n4631 gnd.n1275 19.3944
R10776 gnd.n4636 gnd.n1275 19.3944
R10777 gnd.n4637 gnd.n4636 19.3944
R10778 gnd.n4639 gnd.n4637 19.3944
R10779 gnd.n4639 gnd.n1272 19.3944
R10780 gnd.n4643 gnd.n1272 19.3944
R10781 gnd.n4643 gnd.n1268 19.3944
R10782 gnd.n4655 gnd.n1268 19.3944
R10783 gnd.n4655 gnd.n1266 19.3944
R10784 gnd.n4659 gnd.n1266 19.3944
R10785 gnd.n4660 gnd.n4659 19.3944
R10786 gnd.n4663 gnd.n4660 19.3944
R10787 gnd.n4663 gnd.n1264 19.3944
R10788 gnd.n4690 gnd.n1264 19.3944
R10789 gnd.n4691 gnd.n4690 19.3944
R10790 gnd.n4694 gnd.n4691 19.3944
R10791 gnd.n4694 gnd.n1262 19.3944
R10792 gnd.n4705 gnd.n1262 19.3944
R10793 gnd.n4705 gnd.n4704 19.3944
R10794 gnd.n4704 gnd.n4703 19.3944
R10795 gnd.n4703 gnd.n1254 19.3944
R10796 gnd.n4730 gnd.n1254 19.3944
R10797 gnd.n4731 gnd.n4730 19.3944
R10798 gnd.n4734 gnd.n4731 19.3944
R10799 gnd.n4734 gnd.n1252 19.3944
R10800 gnd.n4744 gnd.n1252 19.3944
R10801 gnd.n4744 gnd.n4743 19.3944
R10802 gnd.n4743 gnd.n4742 19.3944
R10803 gnd.n4742 gnd.n1245 19.3944
R10804 gnd.n4790 gnd.n1245 19.3944
R10805 gnd.n4790 gnd.n1243 19.3944
R10806 gnd.n4797 gnd.n1243 19.3944
R10807 gnd.n4797 gnd.n4796 19.3944
R10808 gnd.n4796 gnd.n1059 19.3944
R10809 gnd.n6227 gnd.n1059 19.3944
R10810 gnd.n6228 gnd.n6227 19.3944
R10811 gnd.n6266 gnd.n6265 19.3944
R10812 gnd.n6265 gnd.n6264 19.3944
R10813 gnd.n6264 gnd.n1025 19.3944
R10814 gnd.n6259 gnd.n1025 19.3944
R10815 gnd.n6259 gnd.n6258 19.3944
R10816 gnd.n6258 gnd.n6257 19.3944
R10817 gnd.n6257 gnd.n1032 19.3944
R10818 gnd.n6252 gnd.n1032 19.3944
R10819 gnd.n6252 gnd.n6251 19.3944
R10820 gnd.n6251 gnd.n6250 19.3944
R10821 gnd.n6250 gnd.n1039 19.3944
R10822 gnd.n6245 gnd.n1039 19.3944
R10823 gnd.n6245 gnd.n6244 19.3944
R10824 gnd.n6244 gnd.n6243 19.3944
R10825 gnd.n6243 gnd.n1046 19.3944
R10826 gnd.n6238 gnd.n1046 19.3944
R10827 gnd.n6238 gnd.n6237 19.3944
R10828 gnd.n6237 gnd.n6236 19.3944
R10829 gnd.n6297 gnd.n6296 19.3944
R10830 gnd.n6296 gnd.n991 19.3944
R10831 gnd.n993 gnd.n991 19.3944
R10832 gnd.n6289 gnd.n993 19.3944
R10833 gnd.n6289 gnd.n6288 19.3944
R10834 gnd.n6288 gnd.n6287 19.3944
R10835 gnd.n6287 gnd.n1000 19.3944
R10836 gnd.n6282 gnd.n1000 19.3944
R10837 gnd.n6282 gnd.n6281 19.3944
R10838 gnd.n6281 gnd.n6280 19.3944
R10839 gnd.n6280 gnd.n1007 19.3944
R10840 gnd.n6275 gnd.n1007 19.3944
R10841 gnd.n6275 gnd.n6274 19.3944
R10842 gnd.n6274 gnd.n6273 19.3944
R10843 gnd.n6273 gnd.n1014 19.3944
R10844 gnd.n4480 gnd.n1392 19.3944
R10845 gnd.n4492 gnd.n1392 19.3944
R10846 gnd.n4492 gnd.n1390 19.3944
R10847 gnd.n4496 gnd.n1390 19.3944
R10848 gnd.n4496 gnd.n1376 19.3944
R10849 gnd.n4508 gnd.n1376 19.3944
R10850 gnd.n4508 gnd.n1374 19.3944
R10851 gnd.n4512 gnd.n1374 19.3944
R10852 gnd.n4512 gnd.n1360 19.3944
R10853 gnd.n4524 gnd.n1360 19.3944
R10854 gnd.n4524 gnd.n1358 19.3944
R10855 gnd.n4528 gnd.n1358 19.3944
R10856 gnd.n4528 gnd.n1344 19.3944
R10857 gnd.n4540 gnd.n1344 19.3944
R10858 gnd.n4540 gnd.n1342 19.3944
R10859 gnd.n4544 gnd.n1342 19.3944
R10860 gnd.n4544 gnd.n1327 19.3944
R10861 gnd.n4564 gnd.n1327 19.3944
R10862 gnd.n4564 gnd.n1325 19.3944
R10863 gnd.n4570 gnd.n1325 19.3944
R10864 gnd.n4570 gnd.n4569 19.3944
R10865 gnd.n4569 gnd.n1291 19.3944
R10866 gnd.n4604 gnd.n1291 19.3944
R10867 gnd.n4604 gnd.n1289 19.3944
R10868 gnd.n4608 gnd.n1289 19.3944
R10869 gnd.n4609 gnd.n4608 19.3944
R10870 gnd.n4609 gnd.n1182 19.3944
R10871 gnd.n4879 gnd.n4878 19.3944
R10872 gnd.n4868 gnd.n4867 19.3944
R10873 gnd.n4865 gnd.n4864 19.3944
R10874 gnd.n4854 gnd.n4853 19.3944
R10875 gnd.n4882 gnd.n1175 19.3944
R10876 gnd.n4882 gnd.n1160 19.3944
R10877 gnd.n4894 gnd.n1160 19.3944
R10878 gnd.n4894 gnd.n1158 19.3944
R10879 gnd.n4898 gnd.n1158 19.3944
R10880 gnd.n4898 gnd.n1143 19.3944
R10881 gnd.n4910 gnd.n1143 19.3944
R10882 gnd.n4910 gnd.n1141 19.3944
R10883 gnd.n4914 gnd.n1141 19.3944
R10884 gnd.n4914 gnd.n1126 19.3944
R10885 gnd.n4926 gnd.n1126 19.3944
R10886 gnd.n4926 gnd.n1124 19.3944
R10887 gnd.n4930 gnd.n1124 19.3944
R10888 gnd.n4930 gnd.n1109 19.3944
R10889 gnd.n4942 gnd.n1109 19.3944
R10890 gnd.n4942 gnd.n1107 19.3944
R10891 gnd.n4946 gnd.n1107 19.3944
R10892 gnd.n4946 gnd.n1092 19.3944
R10893 gnd.n4958 gnd.n1092 19.3944
R10894 gnd.n4958 gnd.n1090 19.3944
R10895 gnd.n4962 gnd.n1090 19.3944
R10896 gnd.n4962 gnd.n1075 19.3944
R10897 gnd.n4974 gnd.n1075 19.3944
R10898 gnd.n4974 gnd.n1073 19.3944
R10899 gnd.n4980 gnd.n1073 19.3944
R10900 gnd.n4980 gnd.n4979 19.3944
R10901 gnd.n4979 gnd.n988 19.3944
R10902 gnd.n6300 gnd.n988 19.3944
R10903 gnd.n2557 gnd.n1599 19.3944
R10904 gnd.n2557 gnd.n1597 19.3944
R10905 gnd.n2561 gnd.n1597 19.3944
R10906 gnd.n2561 gnd.n1593 19.3944
R10907 gnd.n2567 gnd.n1593 19.3944
R10908 gnd.n2567 gnd.n1591 19.3944
R10909 gnd.n2571 gnd.n1591 19.3944
R10910 gnd.n2571 gnd.n1587 19.3944
R10911 gnd.n2577 gnd.n1587 19.3944
R10912 gnd.n2577 gnd.n1585 19.3944
R10913 gnd.n2581 gnd.n1585 19.3944
R10914 gnd.n2581 gnd.n1581 19.3944
R10915 gnd.n2587 gnd.n1581 19.3944
R10916 gnd.n2587 gnd.n1579 19.3944
R10917 gnd.n2591 gnd.n1579 19.3944
R10918 gnd.n2591 gnd.n1575 19.3944
R10919 gnd.n2597 gnd.n1575 19.3944
R10920 gnd.n2597 gnd.n1573 19.3944
R10921 gnd.n2601 gnd.n1573 19.3944
R10922 gnd.n2601 gnd.n1569 19.3944
R10923 gnd.n2607 gnd.n1569 19.3944
R10924 gnd.n2607 gnd.n1567 19.3944
R10925 gnd.n2611 gnd.n1567 19.3944
R10926 gnd.n2611 gnd.n1563 19.3944
R10927 gnd.n2617 gnd.n1563 19.3944
R10928 gnd.n2617 gnd.n1561 19.3944
R10929 gnd.n2621 gnd.n1561 19.3944
R10930 gnd.n2621 gnd.n1557 19.3944
R10931 gnd.n2627 gnd.n1557 19.3944
R10932 gnd.n2627 gnd.n1555 19.3944
R10933 gnd.n2631 gnd.n1555 19.3944
R10934 gnd.n2631 gnd.n1551 19.3944
R10935 gnd.n2637 gnd.n1551 19.3944
R10936 gnd.n2637 gnd.n1549 19.3944
R10937 gnd.n2641 gnd.n1549 19.3944
R10938 gnd.n2641 gnd.n1545 19.3944
R10939 gnd.n2647 gnd.n1545 19.3944
R10940 gnd.n2647 gnd.n1543 19.3944
R10941 gnd.n2651 gnd.n1543 19.3944
R10942 gnd.n2651 gnd.n1539 19.3944
R10943 gnd.n2657 gnd.n1539 19.3944
R10944 gnd.n2657 gnd.n1537 19.3944
R10945 gnd.n2661 gnd.n1537 19.3944
R10946 gnd.n2661 gnd.n1533 19.3944
R10947 gnd.n2667 gnd.n1533 19.3944
R10948 gnd.n2667 gnd.n1531 19.3944
R10949 gnd.n2671 gnd.n1531 19.3944
R10950 gnd.n2671 gnd.n1527 19.3944
R10951 gnd.n2677 gnd.n1527 19.3944
R10952 gnd.n2677 gnd.n1525 19.3944
R10953 gnd.n2681 gnd.n1525 19.3944
R10954 gnd.n2681 gnd.n1521 19.3944
R10955 gnd.n2687 gnd.n1521 19.3944
R10956 gnd.n2687 gnd.n1519 19.3944
R10957 gnd.n2691 gnd.n1519 19.3944
R10958 gnd.n2691 gnd.n1515 19.3944
R10959 gnd.n2697 gnd.n1515 19.3944
R10960 gnd.n2697 gnd.n1513 19.3944
R10961 gnd.n2701 gnd.n1513 19.3944
R10962 gnd.n2701 gnd.n1509 19.3944
R10963 gnd.n2707 gnd.n1509 19.3944
R10964 gnd.n2707 gnd.n1507 19.3944
R10965 gnd.n2711 gnd.n1507 19.3944
R10966 gnd.n2711 gnd.n1503 19.3944
R10967 gnd.n2717 gnd.n1503 19.3944
R10968 gnd.n2717 gnd.n1501 19.3944
R10969 gnd.n2721 gnd.n1501 19.3944
R10970 gnd.n2721 gnd.n1497 19.3944
R10971 gnd.n2727 gnd.n1497 19.3944
R10972 gnd.n2727 gnd.n1495 19.3944
R10973 gnd.n2731 gnd.n1495 19.3944
R10974 gnd.n2731 gnd.n1491 19.3944
R10975 gnd.n2737 gnd.n1491 19.3944
R10976 gnd.n2737 gnd.n1489 19.3944
R10977 gnd.n2741 gnd.n1489 19.3944
R10978 gnd.n2741 gnd.n1485 19.3944
R10979 gnd.n2747 gnd.n1485 19.3944
R10980 gnd.n2747 gnd.n1483 19.3944
R10981 gnd.n2751 gnd.n1483 19.3944
R10982 gnd.n2751 gnd.n1479 19.3944
R10983 gnd.n2757 gnd.n1479 19.3944
R10984 gnd.n2757 gnd.n1477 19.3944
R10985 gnd.n2764 gnd.n1477 19.3944
R10986 gnd.n2764 gnd.n2763 19.3944
R10987 gnd.n6217 gnd.n6216 19.3944
R10988 gnd.n6216 gnd.n6215 19.3944
R10989 gnd.n6215 gnd.n5096 19.3944
R10990 gnd.n6211 gnd.n5096 19.3944
R10991 gnd.n6211 gnd.n6210 19.3944
R10992 gnd.n6210 gnd.n6209 19.3944
R10993 gnd.n6209 gnd.n5100 19.3944
R10994 gnd.n6205 gnd.n5100 19.3944
R10995 gnd.n6205 gnd.n6204 19.3944
R10996 gnd.n6204 gnd.n6203 19.3944
R10997 gnd.n6203 gnd.n5104 19.3944
R10998 gnd.n6199 gnd.n5104 19.3944
R10999 gnd.n6199 gnd.n6198 19.3944
R11000 gnd.n6198 gnd.n6197 19.3944
R11001 gnd.n6197 gnd.n5108 19.3944
R11002 gnd.n6193 gnd.n5108 19.3944
R11003 gnd.n6193 gnd.n6192 19.3944
R11004 gnd.n6192 gnd.n6191 19.3944
R11005 gnd.n6191 gnd.n5112 19.3944
R11006 gnd.n6187 gnd.n5112 19.3944
R11007 gnd.n6187 gnd.n6186 19.3944
R11008 gnd.n6186 gnd.n6185 19.3944
R11009 gnd.n6185 gnd.n5116 19.3944
R11010 gnd.n6181 gnd.n5116 19.3944
R11011 gnd.n6181 gnd.n6180 19.3944
R11012 gnd.n6180 gnd.n6179 19.3944
R11013 gnd.n6179 gnd.n5120 19.3944
R11014 gnd.n6175 gnd.n5120 19.3944
R11015 gnd.n6175 gnd.n6174 19.3944
R11016 gnd.n6174 gnd.n6173 19.3944
R11017 gnd.n6173 gnd.n5124 19.3944
R11018 gnd.n6169 gnd.n5124 19.3944
R11019 gnd.n6169 gnd.n6168 19.3944
R11020 gnd.n6168 gnd.n6167 19.3944
R11021 gnd.n6167 gnd.n5128 19.3944
R11022 gnd.n6163 gnd.n5128 19.3944
R11023 gnd.n6163 gnd.n6162 19.3944
R11024 gnd.n6162 gnd.n6161 19.3944
R11025 gnd.n6161 gnd.n5132 19.3944
R11026 gnd.n6157 gnd.n5132 19.3944
R11027 gnd.n6157 gnd.n6156 19.3944
R11028 gnd.n6156 gnd.n6155 19.3944
R11029 gnd.n6155 gnd.n5136 19.3944
R11030 gnd.n6151 gnd.n5136 19.3944
R11031 gnd.n6151 gnd.n6150 19.3944
R11032 gnd.n6150 gnd.n6149 19.3944
R11033 gnd.n6149 gnd.n5140 19.3944
R11034 gnd.n6145 gnd.n5140 19.3944
R11035 gnd.n6145 gnd.n6144 19.3944
R11036 gnd.n6144 gnd.n6143 19.3944
R11037 gnd.n6143 gnd.n5144 19.3944
R11038 gnd.n6139 gnd.n5144 19.3944
R11039 gnd.n6139 gnd.n6138 19.3944
R11040 gnd.n6138 gnd.n6137 19.3944
R11041 gnd.n6137 gnd.n5148 19.3944
R11042 gnd.n6133 gnd.n5148 19.3944
R11043 gnd.n6133 gnd.n6132 19.3944
R11044 gnd.n6132 gnd.n6131 19.3944
R11045 gnd.n6131 gnd.n5152 19.3944
R11046 gnd.n6127 gnd.n5152 19.3944
R11047 gnd.n6127 gnd.n6126 19.3944
R11048 gnd.n6126 gnd.n6125 19.3944
R11049 gnd.n6125 gnd.n5156 19.3944
R11050 gnd.n6121 gnd.n5156 19.3944
R11051 gnd.n6121 gnd.n6120 19.3944
R11052 gnd.n6120 gnd.n6119 19.3944
R11053 gnd.n6119 gnd.n5160 19.3944
R11054 gnd.n6115 gnd.n5160 19.3944
R11055 gnd.n6115 gnd.n6114 19.3944
R11056 gnd.n6114 gnd.n6113 19.3944
R11057 gnd.n6113 gnd.n5939 19.3944
R11058 gnd.n6109 gnd.n5939 19.3944
R11059 gnd.n6109 gnd.n6108 19.3944
R11060 gnd.n6108 gnd.n6107 19.3944
R11061 gnd.n6107 gnd.n5943 19.3944
R11062 gnd.n6103 gnd.n5943 19.3944
R11063 gnd.n6103 gnd.n6102 19.3944
R11064 gnd.n6102 gnd.n6101 19.3944
R11065 gnd.n6101 gnd.n5947 19.3944
R11066 gnd.n6097 gnd.n5947 19.3944
R11067 gnd.n6097 gnd.n6096 19.3944
R11068 gnd.n6096 gnd.n6095 19.3944
R11069 gnd.n6030 gnd.n6029 19.3944
R11070 gnd.n6029 gnd.n633 19.3944
R11071 gnd.n6674 gnd.n633 19.3944
R11072 gnd.n6092 gnd.n5951 19.3944
R11073 gnd.n6085 gnd.n5951 19.3944
R11074 gnd.n6085 gnd.n6084 19.3944
R11075 gnd.n6084 gnd.n5969 19.3944
R11076 gnd.n6077 gnd.n5969 19.3944
R11077 gnd.n6077 gnd.n6076 19.3944
R11078 gnd.n6076 gnd.n5977 19.3944
R11079 gnd.n6069 gnd.n5977 19.3944
R11080 gnd.n6069 gnd.n6068 19.3944
R11081 gnd.n6068 gnd.n5989 19.3944
R11082 gnd.n6061 gnd.n5989 19.3944
R11083 gnd.n6061 gnd.n6060 19.3944
R11084 gnd.n6060 gnd.n5997 19.3944
R11085 gnd.n6053 gnd.n5997 19.3944
R11086 gnd.n6053 gnd.n6052 19.3944
R11087 gnd.n6052 gnd.n6009 19.3944
R11088 gnd.n6042 gnd.n6009 19.3944
R11089 gnd.n6042 gnd.n6041 19.3944
R11090 gnd.n6041 gnd.n6040 19.3944
R11091 gnd.n6040 gnd.n6016 19.3944
R11092 gnd.n6036 gnd.n6016 19.3944
R11093 gnd.n6036 gnd.n6035 19.3944
R11094 gnd.n6035 gnd.n6034 19.3944
R11095 gnd.n6034 gnd.n6022 19.3944
R11096 gnd.n3591 gnd.t23 18.8012
R11097 gnd.n3024 gnd.t30 18.8012
R11098 gnd.n3461 gnd.n3460 18.4825
R11099 gnd.n6417 gnd.n871 18.4825
R11100 gnd.t6 gnd.n819 18.4825
R11101 gnd.t8 gnd.n755 18.4825
R11102 gnd.n6593 gnd.n703 18.4825
R11103 gnd.n6879 gnd.n6878 18.4247
R11104 gnd.n1018 gnd.n1014 18.4247
R11105 gnd.n7310 gnd.n120 18.2308
R11106 gnd.n6049 gnd.n6003 18.2308
R11107 gnd.n5055 gnd.n978 18.2308
R11108 gnd.n4231 gnd.n4175 18.2308
R11109 gnd.t13 gnd.n3140 18.1639
R11110 gnd.n3169 gnd.t21 17.5266
R11111 gnd.n4069 gnd.n2767 17.2079
R11112 gnd.n5367 gnd.n5366 17.2079
R11113 gnd.n6409 gnd.n879 17.2079
R11114 gnd.n6465 gnd.n825 17.2079
R11115 gnd.n6545 gnd.n749 17.2079
R11116 gnd.n6601 gnd.n696 17.2079
R11117 gnd.n7253 gnd.n236 17.2079
R11118 gnd.n3580 gnd.t17 16.8893
R11119 gnd.n4856 gnd.n1207 16.5706
R11120 gnd.n4884 gnd.n1170 16.5706
R11121 gnd.n4844 gnd.n1173 16.5706
R11122 gnd.n4661 gnd.n1164 16.5706
R11123 gnd.n4900 gnd.n1154 16.5706
R11124 gnd.n4688 gnd.n4687 16.5706
R11125 gnd.n4908 gnd.n1145 16.5706
R11126 gnd.n4916 gnd.n1136 16.5706
R11127 gnd.n4707 gnd.n1139 16.5706
R11128 gnd.n4701 gnd.n1130 16.5706
R11129 gnd.n4932 gnd.n1120 16.5706
R11130 gnd.n4728 gnd.n4727 16.5706
R11131 gnd.n4940 gnd.n1111 16.5706
R11132 gnd.n4948 gnd.n1102 16.5706
R11133 gnd.n4746 gnd.n1105 16.5706
R11134 gnd.n4740 gnd.n1096 16.5706
R11135 gnd.n4964 gnd.n1086 16.5706
R11136 gnd.n4788 gnd.n4787 16.5706
R11137 gnd.n4972 gnd.n1077 16.5706
R11138 gnd.n4799 gnd.n1080 16.5706
R11139 gnd.n4982 gnd.n1067 16.5706
R11140 gnd.n4801 gnd.n1070 16.5706
R11141 gnd.n6225 gnd.n1061 16.5706
R11142 gnd.n6302 gnd.n982 16.5706
R11143 gnd.n5647 gnd.t171 16.5706
R11144 gnd.n5729 gnd.t147 16.5706
R11145 gnd.n6834 gnd.n480 16.5706
R11146 gnd.n6915 gnd.n483 16.5706
R11147 gnd.n6706 gnd.n471 16.5706
R11148 gnd.n6923 gnd.n474 16.5706
R11149 gnd.n6710 gnd.n462 16.5706
R11150 gnd.n6931 gnd.n465 16.5706
R11151 gnd.n6726 gnd.n6725 16.5706
R11152 gnd.n6939 gnd.n456 16.5706
R11153 gnd.n6719 gnd.n446 16.5706
R11154 gnd.n6746 gnd.n437 16.5706
R11155 gnd.n6955 gnd.n440 16.5706
R11156 gnd.n6963 gnd.n431 16.5706
R11157 gnd.n6765 gnd.n6764 16.5706
R11158 gnd.n6971 gnd.n422 16.5706
R11159 gnd.n6758 gnd.n412 16.5706
R11160 gnd.n6777 gnd.n401 16.5706
R11161 gnd.n6990 gnd.n404 16.5706
R11162 gnd.n6998 gnd.n386 16.5706
R11163 gnd.n7019 gnd.n7018 16.5706
R11164 gnd.n7041 gnd.n372 16.5706
R11165 gnd.n6790 gnd.n379 16.5706
R11166 gnd.n7050 gnd.n361 16.5706
R11167 gnd.n7072 gnd.n349 16.5706
R11168 gnd.n7180 gnd.n311 16.5706
R11169 gnd.n3396 gnd.t105 16.2519
R11170 gnd.n3628 gnd.t15 16.2519
R11171 gnd.n4852 gnd.t188 16.2519
R11172 gnd.n6345 gnd.t112 16.2519
R11173 gnd.n6668 gnd.t89 16.2519
R11174 gnd.t286 gnd.n308 16.2519
R11175 gnd.n6401 gnd.n887 15.9333
R11176 gnd.n5322 gnd.n817 15.9333
R11177 gnd.n6473 gnd.n817 15.9333
R11178 gnd.n6537 gnd.n757 15.9333
R11179 gnd.n5276 gnd.n757 15.9333
R11180 gnd.n4022 gnd.n4020 15.6674
R11181 gnd.n3990 gnd.n3988 15.6674
R11182 gnd.n3958 gnd.n3956 15.6674
R11183 gnd.n3927 gnd.n3925 15.6674
R11184 gnd.n3895 gnd.n3893 15.6674
R11185 gnd.n3863 gnd.n3861 15.6674
R11186 gnd.n3831 gnd.n3829 15.6674
R11187 gnd.n3800 gnd.n3798 15.6674
R11188 gnd.n3387 gnd.t105 15.6146
R11189 gnd.t61 gnd.n4058 15.6146
R11190 gnd.t82 gnd.n2776 15.6146
R11191 gnd.t190 gnd.n1148 15.6146
R11192 gnd.t112 gnd.n929 15.6146
R11193 gnd.n5610 gnd.t145 15.6146
R11194 gnd.n5764 gnd.t148 15.6146
R11195 gnd.n648 gnd.t89 15.6146
R11196 gnd.n6999 gnd.t231 15.6146
R11197 gnd.n4645 gnd.n1207 15.296
R11198 gnd.n4856 gnd.n4852 15.296
R11199 gnd.n4653 gnd.n1170 15.296
R11200 gnd.n4884 gnd.n1173 15.296
R11201 gnd.n4845 gnd.n4844 15.296
R11202 gnd.n4892 gnd.n1164 15.296
R11203 gnd.n4661 gnd.n1154 15.296
R11204 gnd.n4688 gnd.n1145 15.296
R11205 gnd.n4908 gnd.n1148 15.296
R11206 gnd.n4692 gnd.n1136 15.296
R11207 gnd.n4916 gnd.n1139 15.296
R11208 gnd.n4708 gnd.n4707 15.296
R11209 gnd.n4924 gnd.n1130 15.296
R11210 gnd.n4701 gnd.n1120 15.296
R11211 gnd.n4728 gnd.n1111 15.296
R11212 gnd.n4940 gnd.n1114 15.296
R11213 gnd.n4732 gnd.n1102 15.296
R11214 gnd.n4948 gnd.n1105 15.296
R11215 gnd.n4747 gnd.n4746 15.296
R11216 gnd.n4956 gnd.n1096 15.296
R11217 gnd.n4740 gnd.n1086 15.296
R11218 gnd.n4788 gnd.n1077 15.296
R11219 gnd.n4972 gnd.n1080 15.296
R11220 gnd.n4799 gnd.n1067 15.296
R11221 gnd.n4982 gnd.n1070 15.296
R11222 gnd.n6225 gnd.n982 15.296
R11223 gnd.n6302 gnd.n984 15.296
R11224 gnd.n6834 gnd.n564 15.296
R11225 gnd.n6915 gnd.n480 15.296
R11226 gnd.n6923 gnd.n471 15.296
R11227 gnd.n6710 gnd.n474 15.296
R11228 gnd.n6931 gnd.n462 15.296
R11229 gnd.n6725 gnd.n465 15.296
R11230 gnd.n6719 gnd.n456 15.296
R11231 gnd.n6947 gnd.n446 15.296
R11232 gnd.n6746 gnd.n6745 15.296
R11233 gnd.n6955 gnd.n437 15.296
R11234 gnd.n6750 gnd.n440 15.296
R11235 gnd.n6963 gnd.n428 15.296
R11236 gnd.n6764 gnd.n431 15.296
R11237 gnd.n6758 gnd.n422 15.296
R11238 gnd.n6979 gnd.n412 15.296
R11239 gnd.n6777 gnd.n6776 15.296
R11240 gnd.n6990 gnd.n401 15.296
R11241 gnd.n6798 gnd.n404 15.296
R11242 gnd.n6999 gnd.n6998 15.296
R11243 gnd.n7019 gnd.n386 15.296
R11244 gnd.n6790 gnd.n372 15.296
R11245 gnd.n7029 gnd.n379 15.296
R11246 gnd.n7050 gnd.n359 15.296
R11247 gnd.n361 gnd.n349 15.296
R11248 gnd.n7072 gnd.n7071 15.296
R11249 gnd.n7180 gnd.n308 15.296
R11250 gnd.n7062 gnd.n311 15.296
R11251 gnd.n5170 gnd.n5169 15.0827
R11252 gnd.n5417 gnd.n5412 15.0481
R11253 gnd.n5180 gnd.n5179 15.0481
R11254 gnd.n2852 gnd.t22 14.9773
R11255 gnd.t206 gnd.n1114 14.9773
R11256 gnd.t346 gnd.n809 14.9773
R11257 gnd.t160 gnd.n765 14.9773
R11258 gnd.t294 gnd.n428 14.9773
R11259 gnd.n5356 gnd.n879 14.6587
R11260 gnd.n6425 gnd.t28 14.6587
R11261 gnd.n5637 gnd.n825 14.6587
R11262 gnd.n6481 gnd.n809 14.6587
R11263 gnd.n6529 gnd.n765 14.6587
R11264 gnd.n5271 gnd.n749 14.6587
R11265 gnd.n6585 gnd.t150 14.6587
R11266 gnd.n5243 gnd.n696 14.6587
R11267 gnd.n6617 gnd.n681 14.6587
R11268 gnd.n2827 gnd.t142 14.34
R11269 gnd.n2810 gnd.t20 14.34
R11270 gnd.n3549 gnd.t154 13.7027
R11271 gnd.n3253 gnd.n3252 13.5763
R11272 gnd.n4134 gnd.n1438 13.5763
R11273 gnd.n6841 gnd.n561 13.5763
R11274 gnd.n7362 gnd.n7361 13.5763
R11275 gnd.n4407 gnd.n4346 13.5763
R11276 gnd.n6236 gnd.n1055 13.5763
R11277 gnd.n3461 gnd.n3199 13.384
R11278 gnd.n5629 gnd.n5331 13.384
R11279 gnd.n5629 gnd.t9 13.384
R11280 gnd.n6489 gnd.n801 13.384
R11281 gnd.n6521 gnd.n773 13.384
R11282 gnd.n5266 gnd.t27 13.384
R11283 gnd.n5266 gnd.n5265 13.384
R11284 gnd.n5780 gnd.n703 13.384
R11285 gnd.n5428 gnd.n5409 13.1884
R11286 gnd.n5423 gnd.n5422 13.1884
R11287 gnd.n5422 gnd.n5421 13.1884
R11288 gnd.n5173 gnd.n5168 13.1884
R11289 gnd.n5174 gnd.n5173 13.1884
R11290 gnd.n5424 gnd.n5411 13.146
R11291 gnd.n5420 gnd.n5411 13.146
R11292 gnd.n5172 gnd.n5171 13.146
R11293 gnd.n5172 gnd.n5167 13.146
R11294 gnd.n5361 gnd.t167 13.0654
R11295 gnd.n5795 gnd.t4 13.0654
R11296 gnd.n4023 gnd.n4019 12.8005
R11297 gnd.n3991 gnd.n3987 12.8005
R11298 gnd.n3959 gnd.n3955 12.8005
R11299 gnd.n3928 gnd.n3924 12.8005
R11300 gnd.n3896 gnd.n3892 12.8005
R11301 gnd.n3864 gnd.n3860 12.8005
R11302 gnd.n3832 gnd.n3828 12.8005
R11303 gnd.n3801 gnd.n3797 12.8005
R11304 gnd.t65 gnd.t35 12.7467
R11305 gnd.n1372 gnd.t196 12.4281
R11306 gnd.n4956 gnd.t208 12.4281
R11307 gnd.n6947 gnd.t225 12.4281
R11308 gnd.t212 gnd.n225 12.4281
R11309 gnd.n3252 gnd.n3247 12.4126
R11310 gnd.n4137 gnd.n4134 12.4126
R11311 gnd.n6837 gnd.n561 12.4126
R11312 gnd.n7361 gnd.n196 12.4126
R11313 gnd.n4403 gnd.n4346 12.4126
R11314 gnd.n6231 gnd.n1055 12.4126
R11315 gnd.n5431 gnd.n5430 12.1761
R11316 gnd.n5930 gnd.n5929 12.1761
R11317 gnd.n5346 gnd.n5345 12.1094
R11318 gnd.n5619 gnd.t26 12.1094
R11319 gnd.n5261 gnd.t151 12.1094
R11320 gnd.n5773 gnd.n5251 12.1094
R11321 gnd.n5788 gnd.t93 12.1094
R11322 gnd.n5935 gnd.t47 12.1094
R11323 gnd.n4027 gnd.n4026 12.0247
R11324 gnd.n3995 gnd.n3994 12.0247
R11325 gnd.n3963 gnd.n3962 12.0247
R11326 gnd.n3932 gnd.n3931 12.0247
R11327 gnd.n3900 gnd.n3899 12.0247
R11328 gnd.n3868 gnd.n3867 12.0247
R11329 gnd.n3836 gnd.n3835 12.0247
R11330 gnd.n3805 gnd.n3804 12.0247
R11331 gnd.n1340 gnd.t250 11.7908
R11332 gnd.n4924 gnd.t227 11.7908
R11333 gnd.t72 gnd.n1061 11.7908
R11334 gnd.t57 gnd.n483 11.7908
R11335 gnd.n6979 gnd.t258 11.7908
R11336 gnd.t282 gnd.n256 11.7908
R11337 gnd.n5367 gnd.t50 11.4721
R11338 gnd.t7 gnd.n801 11.4721
R11339 gnd.t144 gnd.n773 11.4721
R11340 gnd.n4030 gnd.n4017 11.249
R11341 gnd.n3998 gnd.n3985 11.249
R11342 gnd.n3966 gnd.n3953 11.249
R11343 gnd.n3935 gnd.n3922 11.249
R11344 gnd.n3903 gnd.n3890 11.249
R11345 gnd.n3871 gnd.n3858 11.249
R11346 gnd.n3839 gnd.n3826 11.249
R11347 gnd.n3808 gnd.n3795 11.249
R11348 gnd.n3539 gnd.t154 11.1535
R11349 gnd.n4596 gnd.t180 11.1535
R11350 gnd.n4892 gnd.t182 11.1535
R11351 gnd.n923 gnd.t342 11.1535
R11352 gnd.t158 gnd.n834 11.1535
R11353 gnd.t338 gnd.n740 11.1535
R11354 gnd.t340 gnd.n654 11.1535
R11355 gnd.n7029 gnd.t276 11.1535
R11356 gnd.t248 gnd.n286 11.1535
R11357 gnd.n5610 gnd.n5341 10.8348
R11358 gnd.n6505 gnd.n786 10.8348
R11359 gnd.n6505 gnd.n788 10.8348
R11360 gnd.n5764 gnd.n5763 10.8348
R11361 gnd.n5864 gnd.n5210 10.6151
R11362 gnd.n5864 gnd.n5863 10.6151
R11363 gnd.n5861 gnd.n5214 10.6151
R11364 gnd.n5856 gnd.n5214 10.6151
R11365 gnd.n5856 gnd.n5855 10.6151
R11366 gnd.n5855 gnd.n5854 10.6151
R11367 gnd.n5854 gnd.n5217 10.6151
R11368 gnd.n5849 gnd.n5217 10.6151
R11369 gnd.n5849 gnd.n5848 10.6151
R11370 gnd.n5848 gnd.n5847 10.6151
R11371 gnd.n5847 gnd.n5220 10.6151
R11372 gnd.n5842 gnd.n5220 10.6151
R11373 gnd.n5842 gnd.n5841 10.6151
R11374 gnd.n5841 gnd.n5840 10.6151
R11375 gnd.n5840 gnd.n5223 10.6151
R11376 gnd.n5835 gnd.n5223 10.6151
R11377 gnd.n5835 gnd.n5834 10.6151
R11378 gnd.n5834 gnd.n5833 10.6151
R11379 gnd.n5833 gnd.n5226 10.6151
R11380 gnd.n5828 gnd.n5226 10.6151
R11381 gnd.n5828 gnd.n5827 10.6151
R11382 gnd.n5827 gnd.n5826 10.6151
R11383 gnd.n5826 gnd.n5229 10.6151
R11384 gnd.n5821 gnd.n5229 10.6151
R11385 gnd.n5821 gnd.n5820 10.6151
R11386 gnd.n5820 gnd.n5819 10.6151
R11387 gnd.n5819 gnd.n5232 10.6151
R11388 gnd.n5814 gnd.n5232 10.6151
R11389 gnd.n5814 gnd.n5813 10.6151
R11390 gnd.n5813 gnd.n5812 10.6151
R11391 gnd.n5565 gnd.n5562 10.6151
R11392 gnd.n5565 gnd.n5564 10.6151
R11393 gnd.n5564 gnd.n5563 10.6151
R11394 gnd.n5563 gnd.n5359 10.6151
R11395 gnd.n5579 gnd.n5359 10.6151
R11396 gnd.n5580 gnd.n5579 10.6151
R11397 gnd.n5583 gnd.n5580 10.6151
R11398 gnd.n5583 gnd.n5582 10.6151
R11399 gnd.n5582 gnd.n5581 10.6151
R11400 gnd.n5581 gnd.n5349 10.6151
R11401 gnd.n5597 gnd.n5349 10.6151
R11402 gnd.n5598 gnd.n5597 10.6151
R11403 gnd.n5600 gnd.n5598 10.6151
R11404 gnd.n5600 gnd.n5599 10.6151
R11405 gnd.n5599 gnd.n5339 10.6151
R11406 gnd.n5612 gnd.n5339 10.6151
R11407 gnd.n5613 gnd.n5612 10.6151
R11408 gnd.n5617 gnd.n5613 10.6151
R11409 gnd.n5617 gnd.n5616 10.6151
R11410 gnd.n5616 gnd.n5615 10.6151
R11411 gnd.n5615 gnd.n5329 10.6151
R11412 gnd.n5631 gnd.n5329 10.6151
R11413 gnd.n5632 gnd.n5631 10.6151
R11414 gnd.n5635 gnd.n5632 10.6151
R11415 gnd.n5635 gnd.n5634 10.6151
R11416 gnd.n5634 gnd.n5633 10.6151
R11417 gnd.n5633 gnd.n5320 10.6151
R11418 gnd.n5650 gnd.n5320 10.6151
R11419 gnd.n5651 gnd.n5650 10.6151
R11420 gnd.n5654 gnd.n5651 10.6151
R11421 gnd.n5654 gnd.n5653 10.6151
R11422 gnd.n5653 gnd.n5652 10.6151
R11423 gnd.n5652 gnd.n5312 10.6151
R11424 gnd.n5312 gnd.n5310 10.6151
R11425 gnd.n5671 gnd.n5310 10.6151
R11426 gnd.n5672 gnd.n5671 10.6151
R11427 gnd.n5674 gnd.n5672 10.6151
R11428 gnd.n5674 gnd.n5673 10.6151
R11429 gnd.n5673 gnd.n5300 10.6151
R11430 gnd.n5687 gnd.n5300 10.6151
R11431 gnd.n5688 gnd.n5687 10.6151
R11432 gnd.n5691 gnd.n5688 10.6151
R11433 gnd.n5691 gnd.n5690 10.6151
R11434 gnd.n5690 gnd.n5689 10.6151
R11435 gnd.n5689 gnd.n5289 10.6151
R11436 gnd.n5705 gnd.n5289 10.6151
R11437 gnd.n5706 gnd.n5705 10.6151
R11438 gnd.n5709 gnd.n5706 10.6151
R11439 gnd.n5709 gnd.n5708 10.6151
R11440 gnd.n5708 gnd.n5707 10.6151
R11441 gnd.n5707 gnd.n5279 10.6151
R11442 gnd.n5723 gnd.n5279 10.6151
R11443 gnd.n5724 gnd.n5723 10.6151
R11444 gnd.n5727 gnd.n5724 10.6151
R11445 gnd.n5727 gnd.n5726 10.6151
R11446 gnd.n5726 gnd.n5725 10.6151
R11447 gnd.n5725 gnd.n5269 10.6151
R11448 gnd.n5741 gnd.n5269 10.6151
R11449 gnd.n5742 gnd.n5741 10.6151
R11450 gnd.n5744 gnd.n5742 10.6151
R11451 gnd.n5744 gnd.n5743 10.6151
R11452 gnd.n5743 gnd.n5259 10.6151
R11453 gnd.n5756 gnd.n5259 10.6151
R11454 gnd.n5757 gnd.n5756 10.6151
R11455 gnd.n5761 gnd.n5757 10.6151
R11456 gnd.n5761 gnd.n5760 10.6151
R11457 gnd.n5760 gnd.n5759 10.6151
R11458 gnd.n5759 gnd.n5249 10.6151
R11459 gnd.n5775 gnd.n5249 10.6151
R11460 gnd.n5776 gnd.n5775 10.6151
R11461 gnd.n5778 gnd.n5776 10.6151
R11462 gnd.n5778 gnd.n5777 10.6151
R11463 gnd.n5777 gnd.n5241 10.6151
R11464 gnd.n5790 gnd.n5241 10.6151
R11465 gnd.n5791 gnd.n5790 10.6151
R11466 gnd.n5793 gnd.n5791 10.6151
R11467 gnd.n5793 gnd.n5792 10.6151
R11468 gnd.n5792 gnd.n5235 10.6151
R11469 gnd.n5806 gnd.n5235 10.6151
R11470 gnd.n5807 gnd.n5806 10.6151
R11471 gnd.n5808 gnd.n5807 10.6151
R11472 gnd.n5497 gnd.n5387 10.6151
R11473 gnd.n5503 gnd.n5387 10.6151
R11474 gnd.n5506 gnd.n5505 10.6151
R11475 gnd.n5506 gnd.n5383 10.6151
R11476 gnd.n5512 gnd.n5383 10.6151
R11477 gnd.n5513 gnd.n5512 10.6151
R11478 gnd.n5514 gnd.n5513 10.6151
R11479 gnd.n5514 gnd.n5381 10.6151
R11480 gnd.n5520 gnd.n5381 10.6151
R11481 gnd.n5521 gnd.n5520 10.6151
R11482 gnd.n5522 gnd.n5521 10.6151
R11483 gnd.n5522 gnd.n5379 10.6151
R11484 gnd.n5528 gnd.n5379 10.6151
R11485 gnd.n5529 gnd.n5528 10.6151
R11486 gnd.n5530 gnd.n5529 10.6151
R11487 gnd.n5530 gnd.n5377 10.6151
R11488 gnd.n5536 gnd.n5377 10.6151
R11489 gnd.n5537 gnd.n5536 10.6151
R11490 gnd.n5538 gnd.n5537 10.6151
R11491 gnd.n5538 gnd.n5375 10.6151
R11492 gnd.n5544 gnd.n5375 10.6151
R11493 gnd.n5545 gnd.n5544 10.6151
R11494 gnd.n5546 gnd.n5545 10.6151
R11495 gnd.n5546 gnd.n5373 10.6151
R11496 gnd.n5552 gnd.n5373 10.6151
R11497 gnd.n5553 gnd.n5552 10.6151
R11498 gnd.n5554 gnd.n5553 10.6151
R11499 gnd.n5554 gnd.n5371 10.6151
R11500 gnd.n5371 gnd.n5370 10.6151
R11501 gnd.n5561 gnd.n5370 10.6151
R11502 gnd.n5431 gnd.n5408 10.6151
R11503 gnd.n5408 gnd.n5407 10.6151
R11504 gnd.n5438 gnd.n5407 10.6151
R11505 gnd.n5439 gnd.n5438 10.6151
R11506 gnd.n5440 gnd.n5439 10.6151
R11507 gnd.n5440 gnd.n5405 10.6151
R11508 gnd.n5446 gnd.n5405 10.6151
R11509 gnd.n5447 gnd.n5446 10.6151
R11510 gnd.n5448 gnd.n5447 10.6151
R11511 gnd.n5448 gnd.n5403 10.6151
R11512 gnd.n5454 gnd.n5403 10.6151
R11513 gnd.n5455 gnd.n5454 10.6151
R11514 gnd.n5456 gnd.n5455 10.6151
R11515 gnd.n5456 gnd.n5401 10.6151
R11516 gnd.n5462 gnd.n5401 10.6151
R11517 gnd.n5463 gnd.n5462 10.6151
R11518 gnd.n5464 gnd.n5463 10.6151
R11519 gnd.n5464 gnd.n5399 10.6151
R11520 gnd.n5470 gnd.n5399 10.6151
R11521 gnd.n5471 gnd.n5470 10.6151
R11522 gnd.n5472 gnd.n5471 10.6151
R11523 gnd.n5472 gnd.n5397 10.6151
R11524 gnd.n5478 gnd.n5397 10.6151
R11525 gnd.n5479 gnd.n5478 10.6151
R11526 gnd.n5480 gnd.n5479 10.6151
R11527 gnd.n5480 gnd.n5395 10.6151
R11528 gnd.n5486 gnd.n5395 10.6151
R11529 gnd.n5487 gnd.n5486 10.6151
R11530 gnd.n5489 gnd.n5391 10.6151
R11531 gnd.n5391 gnd.n5389 10.6151
R11532 gnd.n5929 gnd.n5185 10.6151
R11533 gnd.n5186 gnd.n5185 10.6151
R11534 gnd.n5922 gnd.n5186 10.6151
R11535 gnd.n5922 gnd.n5921 10.6151
R11536 gnd.n5921 gnd.n5920 10.6151
R11537 gnd.n5920 gnd.n5188 10.6151
R11538 gnd.n5915 gnd.n5188 10.6151
R11539 gnd.n5915 gnd.n5914 10.6151
R11540 gnd.n5914 gnd.n5913 10.6151
R11541 gnd.n5913 gnd.n5191 10.6151
R11542 gnd.n5908 gnd.n5191 10.6151
R11543 gnd.n5908 gnd.n5907 10.6151
R11544 gnd.n5907 gnd.n5906 10.6151
R11545 gnd.n5906 gnd.n5194 10.6151
R11546 gnd.n5901 gnd.n5194 10.6151
R11547 gnd.n5901 gnd.n5900 10.6151
R11548 gnd.n5900 gnd.n5899 10.6151
R11549 gnd.n5899 gnd.n5197 10.6151
R11550 gnd.n5894 gnd.n5197 10.6151
R11551 gnd.n5894 gnd.n5893 10.6151
R11552 gnd.n5893 gnd.n5892 10.6151
R11553 gnd.n5892 gnd.n5200 10.6151
R11554 gnd.n5887 gnd.n5200 10.6151
R11555 gnd.n5887 gnd.n5886 10.6151
R11556 gnd.n5886 gnd.n5885 10.6151
R11557 gnd.n5885 gnd.n5203 10.6151
R11558 gnd.n5880 gnd.n5203 10.6151
R11559 gnd.n5880 gnd.n5879 10.6151
R11560 gnd.n5877 gnd.n5208 10.6151
R11561 gnd.n5872 gnd.n5208 10.6151
R11562 gnd.n5429 gnd.n5364 10.6151
R11563 gnd.n5570 gnd.n5364 10.6151
R11564 gnd.n5571 gnd.n5570 10.6151
R11565 gnd.n5574 gnd.n5571 10.6151
R11566 gnd.n5574 gnd.n5573 10.6151
R11567 gnd.n5573 gnd.n5572 10.6151
R11568 gnd.n5572 gnd.n5354 10.6151
R11569 gnd.n5588 gnd.n5354 10.6151
R11570 gnd.n5589 gnd.n5588 10.6151
R11571 gnd.n5592 gnd.n5589 10.6151
R11572 gnd.n5592 gnd.n5591 10.6151
R11573 gnd.n5591 gnd.n5590 10.6151
R11574 gnd.n5590 gnd.n5343 10.6151
R11575 gnd.n5605 gnd.n5343 10.6151
R11576 gnd.n5606 gnd.n5605 10.6151
R11577 gnd.n5608 gnd.n5606 10.6151
R11578 gnd.n5608 gnd.n5607 10.6151
R11579 gnd.n5607 gnd.n5336 10.6151
R11580 gnd.n5336 gnd.n5334 10.6151
R11581 gnd.n5624 gnd.n5334 10.6151
R11582 gnd.n5625 gnd.n5624 10.6151
R11583 gnd.n5627 gnd.n5625 10.6151
R11584 gnd.n5627 gnd.n5626 10.6151
R11585 gnd.n5626 gnd.n5325 10.6151
R11586 gnd.n5641 gnd.n5325 10.6151
R11587 gnd.n5642 gnd.n5641 10.6151
R11588 gnd.n5645 gnd.n5642 10.6151
R11589 gnd.n5645 gnd.n5644 10.6151
R11590 gnd.n5644 gnd.n5643 10.6151
R11591 gnd.n5643 gnd.n5316 10.6151
R11592 gnd.n5660 gnd.n5316 10.6151
R11593 gnd.n5661 gnd.n5660 10.6151
R11594 gnd.n5665 gnd.n5661 10.6151
R11595 gnd.n5665 gnd.n5664 10.6151
R11596 gnd.n5664 gnd.n5663 10.6151
R11597 gnd.n5663 gnd.n5305 10.6151
R11598 gnd.n5678 gnd.n5305 10.6151
R11599 gnd.n5679 gnd.n5678 10.6151
R11600 gnd.n5682 gnd.n5679 10.6151
R11601 gnd.n5682 gnd.n5681 10.6151
R11602 gnd.n5681 gnd.n5680 10.6151
R11603 gnd.n5680 gnd.n5295 10.6151
R11604 gnd.n5696 gnd.n5295 10.6151
R11605 gnd.n5697 gnd.n5696 10.6151
R11606 gnd.n5700 gnd.n5697 10.6151
R11607 gnd.n5700 gnd.n5699 10.6151
R11608 gnd.n5699 gnd.n5698 10.6151
R11609 gnd.n5698 gnd.n5284 10.6151
R11610 gnd.n5714 gnd.n5284 10.6151
R11611 gnd.n5715 gnd.n5714 10.6151
R11612 gnd.n5718 gnd.n5715 10.6151
R11613 gnd.n5718 gnd.n5717 10.6151
R11614 gnd.n5717 gnd.n5716 10.6151
R11615 gnd.n5716 gnd.n5274 10.6151
R11616 gnd.n5732 gnd.n5274 10.6151
R11617 gnd.n5733 gnd.n5732 10.6151
R11618 gnd.n5736 gnd.n5733 10.6151
R11619 gnd.n5736 gnd.n5735 10.6151
R11620 gnd.n5735 gnd.n5734 10.6151
R11621 gnd.n5734 gnd.n5263 10.6151
R11622 gnd.n5749 gnd.n5263 10.6151
R11623 gnd.n5750 gnd.n5749 10.6151
R11624 gnd.n5752 gnd.n5750 10.6151
R11625 gnd.n5752 gnd.n5751 10.6151
R11626 gnd.n5751 gnd.n5256 10.6151
R11627 gnd.n5256 gnd.n5254 10.6151
R11628 gnd.n5768 gnd.n5254 10.6151
R11629 gnd.n5769 gnd.n5768 10.6151
R11630 gnd.n5771 gnd.n5769 10.6151
R11631 gnd.n5771 gnd.n5770 10.6151
R11632 gnd.n5770 gnd.n5245 10.6151
R11633 gnd.n5784 gnd.n5245 10.6151
R11634 gnd.n5785 gnd.n5784 10.6151
R11635 gnd.n5786 gnd.n5785 10.6151
R11636 gnd.n5786 gnd.n5238 10.6151
R11637 gnd.n5799 gnd.n5238 10.6151
R11638 gnd.n5800 gnd.n5799 10.6151
R11639 gnd.n5801 gnd.n5800 10.6151
R11640 gnd.n5801 gnd.n5165 10.6151
R11641 gnd.n5932 gnd.n5165 10.6151
R11642 gnd.n5932 gnd.n5931 10.6151
R11643 gnd.n3450 gnd.t169 10.5161
R11644 gnd.n3761 gnd.t142 10.5161
R11645 gnd.t20 gnd.n2799 10.5161
R11646 gnd.n4870 gnd.t198 10.5161
R11647 gnd.n4862 gnd.n1200 10.5161
R11648 gnd.n4862 gnd.t221 10.5161
R11649 gnd.n5638 gnd.t158 10.5161
R11650 gnd.n5738 gnd.t338 10.5161
R11651 gnd.n7082 gnd.t210 10.5161
R11652 gnd.n7082 gnd.n7081 10.5161
R11653 gnd.n7088 gnd.t290 10.5161
R11654 gnd.n4031 gnd.n4015 10.4732
R11655 gnd.n3999 gnd.n3983 10.4732
R11656 gnd.n3967 gnd.n3951 10.4732
R11657 gnd.n3936 gnd.n3920 10.4732
R11658 gnd.n3904 gnd.n3888 10.4732
R11659 gnd.n3872 gnd.n3856 10.4732
R11660 gnd.n3840 gnd.n3824 10.4732
R11661 gnd.n3809 gnd.n3793 10.4732
R11662 gnd.n3730 gnd.t22 9.87883
R11663 gnd.n4602 gnd.t194 9.87883
R11664 gnd.n4900 gnd.t202 9.87883
R11665 gnd.n6497 gnd.t163 9.87883
R11666 gnd.n6513 gnd.t152 9.87883
R11667 gnd.n7041 gnd.t215 9.87883
R11668 gnd.n289 gnd.t241 9.87883
R11669 gnd.n7487 gnd.n74 9.81789
R11670 gnd.n4035 gnd.n4034 9.69747
R11671 gnd.n4003 gnd.n4002 9.69747
R11672 gnd.n3971 gnd.n3970 9.69747
R11673 gnd.n3940 gnd.n3939 9.69747
R11674 gnd.n3908 gnd.n3907 9.69747
R11675 gnd.n3876 gnd.n3875 9.69747
R11676 gnd.n3844 gnd.n3843 9.69747
R11677 gnd.n3813 gnd.n3812 9.69747
R11678 gnd.n5602 gnd.n5345 9.56018
R11679 gnd.n5620 gnd.n5619 9.56018
R11680 gnd.n6497 gnd.n795 9.56018
R11681 gnd.n6513 gnd.n779 9.56018
R11682 gnd.n5754 gnd.n5261 9.56018
R11683 gnd.n5252 gnd.n5251 9.56018
R11684 gnd.t93 gnd.n705 9.56018
R11685 gnd.n6220 gnd.n4988 9.45599
R11686 gnd.n5957 gnd.n5955 9.45599
R11687 gnd.n4041 gnd.n4040 9.45567
R11688 gnd.n4009 gnd.n4008 9.45567
R11689 gnd.n3977 gnd.n3976 9.45567
R11690 gnd.n3946 gnd.n3945 9.45567
R11691 gnd.n3914 gnd.n3913 9.45567
R11692 gnd.n3882 gnd.n3881 9.45567
R11693 gnd.n3850 gnd.n3849 9.45567
R11694 gnd.n3819 gnd.n3818 9.45567
R11695 gnd.n3088 gnd.n3087 9.39724
R11696 gnd.n4040 gnd.n4039 9.3005
R11697 gnd.n4013 gnd.n4012 9.3005
R11698 gnd.n4034 gnd.n4033 9.3005
R11699 gnd.n4032 gnd.n4031 9.3005
R11700 gnd.n4017 gnd.n4016 9.3005
R11701 gnd.n4026 gnd.n4025 9.3005
R11702 gnd.n4024 gnd.n4023 9.3005
R11703 gnd.n4008 gnd.n4007 9.3005
R11704 gnd.n3981 gnd.n3980 9.3005
R11705 gnd.n4002 gnd.n4001 9.3005
R11706 gnd.n4000 gnd.n3999 9.3005
R11707 gnd.n3985 gnd.n3984 9.3005
R11708 gnd.n3994 gnd.n3993 9.3005
R11709 gnd.n3992 gnd.n3991 9.3005
R11710 gnd.n3976 gnd.n3975 9.3005
R11711 gnd.n3949 gnd.n3948 9.3005
R11712 gnd.n3970 gnd.n3969 9.3005
R11713 gnd.n3968 gnd.n3967 9.3005
R11714 gnd.n3953 gnd.n3952 9.3005
R11715 gnd.n3962 gnd.n3961 9.3005
R11716 gnd.n3960 gnd.n3959 9.3005
R11717 gnd.n3945 gnd.n3944 9.3005
R11718 gnd.n3918 gnd.n3917 9.3005
R11719 gnd.n3939 gnd.n3938 9.3005
R11720 gnd.n3937 gnd.n3936 9.3005
R11721 gnd.n3922 gnd.n3921 9.3005
R11722 gnd.n3931 gnd.n3930 9.3005
R11723 gnd.n3929 gnd.n3928 9.3005
R11724 gnd.n3913 gnd.n3912 9.3005
R11725 gnd.n3886 gnd.n3885 9.3005
R11726 gnd.n3907 gnd.n3906 9.3005
R11727 gnd.n3905 gnd.n3904 9.3005
R11728 gnd.n3890 gnd.n3889 9.3005
R11729 gnd.n3899 gnd.n3898 9.3005
R11730 gnd.n3897 gnd.n3896 9.3005
R11731 gnd.n3881 gnd.n3880 9.3005
R11732 gnd.n3854 gnd.n3853 9.3005
R11733 gnd.n3875 gnd.n3874 9.3005
R11734 gnd.n3873 gnd.n3872 9.3005
R11735 gnd.n3858 gnd.n3857 9.3005
R11736 gnd.n3867 gnd.n3866 9.3005
R11737 gnd.n3865 gnd.n3864 9.3005
R11738 gnd.n3849 gnd.n3848 9.3005
R11739 gnd.n3822 gnd.n3821 9.3005
R11740 gnd.n3843 gnd.n3842 9.3005
R11741 gnd.n3841 gnd.n3840 9.3005
R11742 gnd.n3826 gnd.n3825 9.3005
R11743 gnd.n3835 gnd.n3834 9.3005
R11744 gnd.n3833 gnd.n3832 9.3005
R11745 gnd.n3818 gnd.n3817 9.3005
R11746 gnd.n3791 gnd.n3790 9.3005
R11747 gnd.n3812 gnd.n3811 9.3005
R11748 gnd.n3810 gnd.n3809 9.3005
R11749 gnd.n3795 gnd.n3794 9.3005
R11750 gnd.n3804 gnd.n3803 9.3005
R11751 gnd.n3802 gnd.n3801 9.3005
R11752 gnd.n4164 gnd.n4163 9.3005
R11753 gnd.n4162 gnd.n1426 9.3005
R11754 gnd.n4161 gnd.n4160 9.3005
R11755 gnd.n4157 gnd.n1427 9.3005
R11756 gnd.n4154 gnd.n1428 9.3005
R11757 gnd.n4153 gnd.n1429 9.3005
R11758 gnd.n4150 gnd.n1430 9.3005
R11759 gnd.n4149 gnd.n1431 9.3005
R11760 gnd.n4146 gnd.n1432 9.3005
R11761 gnd.n4145 gnd.n1433 9.3005
R11762 gnd.n4142 gnd.n1434 9.3005
R11763 gnd.n4141 gnd.n1435 9.3005
R11764 gnd.n4138 gnd.n1436 9.3005
R11765 gnd.n4137 gnd.n1437 9.3005
R11766 gnd.n4134 gnd.n4133 9.3005
R11767 gnd.n4132 gnd.n1438 9.3005
R11768 gnd.n4165 gnd.n1425 9.3005
R11769 gnd.n3469 gnd.n3468 9.3005
R11770 gnd.n3173 gnd.n3172 9.3005
R11771 gnd.n3496 gnd.n3495 9.3005
R11772 gnd.n3497 gnd.n3171 9.3005
R11773 gnd.n3501 gnd.n3498 9.3005
R11774 gnd.n3500 gnd.n3499 9.3005
R11775 gnd.n3145 gnd.n3144 9.3005
R11776 gnd.n3526 gnd.n3525 9.3005
R11777 gnd.n3527 gnd.n3143 9.3005
R11778 gnd.n3537 gnd.n3528 9.3005
R11779 gnd.n3536 gnd.n3529 9.3005
R11780 gnd.n3535 gnd.n3530 9.3005
R11781 gnd.n3533 gnd.n3532 9.3005
R11782 gnd.n3531 gnd.n3115 9.3005
R11783 gnd.n3113 gnd.n3112 9.3005
R11784 gnd.n3585 gnd.n3584 9.3005
R11785 gnd.n3586 gnd.n3111 9.3005
R11786 gnd.n3588 gnd.n3587 9.3005
R11787 gnd.n2931 gnd.n2930 9.3005
R11788 gnd.n3621 gnd.n3620 9.3005
R11789 gnd.n3622 gnd.n2929 9.3005
R11790 gnd.n3626 gnd.n3623 9.3005
R11791 gnd.n3625 gnd.n3624 9.3005
R11792 gnd.n2907 gnd.n2906 9.3005
R11793 gnd.n3652 gnd.n3651 9.3005
R11794 gnd.n3653 gnd.n2905 9.3005
R11795 gnd.n3657 gnd.n3654 9.3005
R11796 gnd.n3656 gnd.n3655 9.3005
R11797 gnd.n2881 gnd.n2880 9.3005
R11798 gnd.n3683 gnd.n3682 9.3005
R11799 gnd.n3684 gnd.n2879 9.3005
R11800 gnd.n3688 gnd.n3685 9.3005
R11801 gnd.n3687 gnd.n3686 9.3005
R11802 gnd.n2856 gnd.n2855 9.3005
R11803 gnd.n3714 gnd.n3713 9.3005
R11804 gnd.n3715 gnd.n2854 9.3005
R11805 gnd.n3719 gnd.n3716 9.3005
R11806 gnd.n3718 gnd.n3717 9.3005
R11807 gnd.n2831 gnd.n2830 9.3005
R11808 gnd.n3745 gnd.n3744 9.3005
R11809 gnd.n3746 gnd.n2829 9.3005
R11810 gnd.n3750 gnd.n3747 9.3005
R11811 gnd.n3749 gnd.n3748 9.3005
R11812 gnd.n2805 gnd.n2804 9.3005
R11813 gnd.n3776 gnd.n3775 9.3005
R11814 gnd.n3777 gnd.n2803 9.3005
R11815 gnd.n3781 gnd.n3778 9.3005
R11816 gnd.n3780 gnd.n3779 9.3005
R11817 gnd.n2780 gnd.n2779 9.3005
R11818 gnd.n4062 gnd.n4061 9.3005
R11819 gnd.n4063 gnd.n2778 9.3005
R11820 gnd.n4067 gnd.n4064 9.3005
R11821 gnd.n4066 gnd.n4065 9.3005
R11822 gnd.n3470 gnd.n3467 9.3005
R11823 gnd.n3252 gnd.n3211 9.3005
R11824 gnd.n3247 gnd.n3246 9.3005
R11825 gnd.n3245 gnd.n3212 9.3005
R11826 gnd.n3244 gnd.n3243 9.3005
R11827 gnd.n3240 gnd.n3213 9.3005
R11828 gnd.n3237 gnd.n3236 9.3005
R11829 gnd.n3235 gnd.n3214 9.3005
R11830 gnd.n3234 gnd.n3233 9.3005
R11831 gnd.n3230 gnd.n3215 9.3005
R11832 gnd.n3227 gnd.n3226 9.3005
R11833 gnd.n3225 gnd.n3216 9.3005
R11834 gnd.n3224 gnd.n3223 9.3005
R11835 gnd.n3220 gnd.n3218 9.3005
R11836 gnd.n3217 gnd.n3197 9.3005
R11837 gnd.n3464 gnd.n3196 9.3005
R11838 gnd.n3466 gnd.n3465 9.3005
R11839 gnd.n3254 gnd.n3253 9.3005
R11840 gnd.n3477 gnd.n3183 9.3005
R11841 gnd.n3484 gnd.n3184 9.3005
R11842 gnd.n3486 gnd.n3485 9.3005
R11843 gnd.n3487 gnd.n3164 9.3005
R11844 gnd.n3506 gnd.n3505 9.3005
R11845 gnd.n3508 gnd.n3156 9.3005
R11846 gnd.n3515 gnd.n3158 9.3005
R11847 gnd.n3516 gnd.n3153 9.3005
R11848 gnd.n3518 gnd.n3517 9.3005
R11849 gnd.n3154 gnd.n3139 9.3005
R11850 gnd.n3137 gnd.n3135 9.3005
R11851 gnd.n3544 gnd.n3543 9.3005
R11852 gnd.n3120 gnd.n3119 9.3005
R11853 gnd.n3577 gnd.n3565 9.3005
R11854 gnd.n3576 gnd.n3567 9.3005
R11855 gnd.n3575 gnd.n3568 9.3005
R11856 gnd.n3570 gnd.n3569 9.3005
R11857 gnd.n3103 gnd.n2940 9.3005
R11858 gnd.n3609 gnd.n2941 9.3005
R11859 gnd.n3611 gnd.n3610 9.3005
R11860 gnd.n3612 gnd.n2924 9.3005
R11861 gnd.n3631 gnd.n3630 9.3005
R11862 gnd.n3633 gnd.n2917 9.3005
R11863 gnd.n3640 gnd.n2918 9.3005
R11864 gnd.n3642 gnd.n3641 9.3005
R11865 gnd.n3643 gnd.n2899 9.3005
R11866 gnd.n3662 gnd.n3661 9.3005
R11867 gnd.n3664 gnd.n2891 9.3005
R11868 gnd.n3671 gnd.n2892 9.3005
R11869 gnd.n3673 gnd.n3672 9.3005
R11870 gnd.n3674 gnd.n2872 9.3005
R11871 gnd.n3693 gnd.n3692 9.3005
R11872 gnd.n3695 gnd.n2865 9.3005
R11873 gnd.n3702 gnd.n2866 9.3005
R11874 gnd.n3704 gnd.n3703 9.3005
R11875 gnd.n3705 gnd.n2848 9.3005
R11876 gnd.n3724 gnd.n3723 9.3005
R11877 gnd.n3726 gnd.n2841 9.3005
R11878 gnd.n3733 gnd.n2842 9.3005
R11879 gnd.n3735 gnd.n3734 9.3005
R11880 gnd.n3736 gnd.n2822 9.3005
R11881 gnd.n3755 gnd.n3754 9.3005
R11882 gnd.n3757 gnd.n2815 9.3005
R11883 gnd.n3764 gnd.n2816 9.3005
R11884 gnd.n3766 gnd.n3765 9.3005
R11885 gnd.n3767 gnd.n2797 9.3005
R11886 gnd.n3786 gnd.n3785 9.3005
R11887 gnd.n3788 gnd.n2789 9.3005
R11888 gnd.n4051 gnd.n2790 9.3005
R11889 gnd.n4053 gnd.n4052 9.3005
R11890 gnd.n4054 gnd.n2771 9.3005
R11891 gnd.n4072 gnd.n4071 9.3005
R11892 gnd.n2772 gnd.n1441 9.3005
R11893 gnd.n3475 gnd.n3474 9.3005
R11894 gnd.n4128 gnd.n1442 9.3005
R11895 gnd.n4127 gnd.n1444 9.3005
R11896 gnd.n4124 gnd.n1445 9.3005
R11897 gnd.n4123 gnd.n1446 9.3005
R11898 gnd.n4120 gnd.n1447 9.3005
R11899 gnd.n4119 gnd.n1448 9.3005
R11900 gnd.n4116 gnd.n1449 9.3005
R11901 gnd.n4115 gnd.n1450 9.3005
R11902 gnd.n4112 gnd.n1451 9.3005
R11903 gnd.n4111 gnd.n1452 9.3005
R11904 gnd.n4108 gnd.n1453 9.3005
R11905 gnd.n4107 gnd.n1454 9.3005
R11906 gnd.n4104 gnd.n1455 9.3005
R11907 gnd.n4103 gnd.n1456 9.3005
R11908 gnd.n4100 gnd.n1457 9.3005
R11909 gnd.n4099 gnd.n1458 9.3005
R11910 gnd.n4096 gnd.n1459 9.3005
R11911 gnd.n4095 gnd.n1460 9.3005
R11912 gnd.n4092 gnd.n1461 9.3005
R11913 gnd.n4091 gnd.n1462 9.3005
R11914 gnd.n4088 gnd.n1463 9.3005
R11915 gnd.n4087 gnd.n1464 9.3005
R11916 gnd.n4084 gnd.n1468 9.3005
R11917 gnd.n4083 gnd.n1469 9.3005
R11918 gnd.n4080 gnd.n1470 9.3005
R11919 gnd.n4079 gnd.n1471 9.3005
R11920 gnd.n4130 gnd.n4129 9.3005
R11921 gnd.n3021 gnd.n2947 9.3005
R11922 gnd.n3019 gnd.n2948 9.3005
R11923 gnd.n3018 gnd.n2949 9.3005
R11924 gnd.n3015 gnd.n2950 9.3005
R11925 gnd.n3014 gnd.n2951 9.3005
R11926 gnd.n3013 gnd.n2952 9.3005
R11927 gnd.n3011 gnd.n2953 9.3005
R11928 gnd.n3010 gnd.n2954 9.3005
R11929 gnd.n3007 gnd.n2955 9.3005
R11930 gnd.n3006 gnd.n2956 9.3005
R11931 gnd.n3005 gnd.n2957 9.3005
R11932 gnd.n3003 gnd.n2958 9.3005
R11933 gnd.n3002 gnd.n2959 9.3005
R11934 gnd.n2997 gnd.n2960 9.3005
R11935 gnd.n2996 gnd.n2961 9.3005
R11936 gnd.n2995 gnd.n2962 9.3005
R11937 gnd.n2993 gnd.n2963 9.3005
R11938 gnd.n2992 gnd.n2964 9.3005
R11939 gnd.n2989 gnd.n2965 9.3005
R11940 gnd.n2988 gnd.n2966 9.3005
R11941 gnd.n2987 gnd.n2967 9.3005
R11942 gnd.n2985 gnd.n2968 9.3005
R11943 gnd.n2984 gnd.n2969 9.3005
R11944 gnd.n2981 gnd.n2970 9.3005
R11945 gnd.n2980 gnd.n2971 9.3005
R11946 gnd.n2979 gnd.n2972 9.3005
R11947 gnd.n2977 gnd.n2973 9.3005
R11948 gnd.n2976 gnd.n2975 9.3005
R11949 gnd.n2974 gnd.n1473 9.3005
R11950 gnd.n3385 gnd.n3384 9.3005
R11951 gnd.n3275 gnd.n3274 9.3005
R11952 gnd.n3399 gnd.n3398 9.3005
R11953 gnd.n3400 gnd.n3273 9.3005
R11954 gnd.n3402 gnd.n3401 9.3005
R11955 gnd.n3263 gnd.n3262 9.3005
R11956 gnd.n3415 gnd.n3414 9.3005
R11957 gnd.n3416 gnd.n3261 9.3005
R11958 gnd.n3448 gnd.n3417 9.3005
R11959 gnd.n3447 gnd.n3418 9.3005
R11960 gnd.n3446 gnd.n3419 9.3005
R11961 gnd.n3445 gnd.n3420 9.3005
R11962 gnd.n3442 gnd.n3421 9.3005
R11963 gnd.n3441 gnd.n3422 9.3005
R11964 gnd.n3440 gnd.n3423 9.3005
R11965 gnd.n3438 gnd.n3424 9.3005
R11966 gnd.n3437 gnd.n3425 9.3005
R11967 gnd.n3434 gnd.n3426 9.3005
R11968 gnd.n3433 gnd.n3427 9.3005
R11969 gnd.n3432 gnd.n3428 9.3005
R11970 gnd.n3430 gnd.n3429 9.3005
R11971 gnd.n3128 gnd.n3127 9.3005
R11972 gnd.n3552 gnd.n3551 9.3005
R11973 gnd.n3553 gnd.n3126 9.3005
R11974 gnd.n3557 gnd.n3554 9.3005
R11975 gnd.n3556 gnd.n3555 9.3005
R11976 gnd.n3091 gnd.n3090 9.3005
R11977 gnd.n3600 gnd.n3599 9.3005
R11978 gnd.n3383 gnd.n3284 9.3005
R11979 gnd.n3286 gnd.n3285 9.3005
R11980 gnd.n3330 gnd.n3328 9.3005
R11981 gnd.n3331 gnd.n3327 9.3005
R11982 gnd.n3334 gnd.n3323 9.3005
R11983 gnd.n3335 gnd.n3322 9.3005
R11984 gnd.n3338 gnd.n3321 9.3005
R11985 gnd.n3339 gnd.n3320 9.3005
R11986 gnd.n3342 gnd.n3319 9.3005
R11987 gnd.n3343 gnd.n3318 9.3005
R11988 gnd.n3346 gnd.n3317 9.3005
R11989 gnd.n3347 gnd.n3316 9.3005
R11990 gnd.n3350 gnd.n3315 9.3005
R11991 gnd.n3351 gnd.n3314 9.3005
R11992 gnd.n3354 gnd.n3313 9.3005
R11993 gnd.n3355 gnd.n3312 9.3005
R11994 gnd.n3358 gnd.n3311 9.3005
R11995 gnd.n3359 gnd.n3310 9.3005
R11996 gnd.n3362 gnd.n3309 9.3005
R11997 gnd.n3363 gnd.n3308 9.3005
R11998 gnd.n3366 gnd.n3307 9.3005
R11999 gnd.n3367 gnd.n3306 9.3005
R12000 gnd.n3370 gnd.n3305 9.3005
R12001 gnd.n3372 gnd.n3304 9.3005
R12002 gnd.n3373 gnd.n3303 9.3005
R12003 gnd.n3374 gnd.n3302 9.3005
R12004 gnd.n3375 gnd.n3301 9.3005
R12005 gnd.n3382 gnd.n3381 9.3005
R12006 gnd.n3391 gnd.n3390 9.3005
R12007 gnd.n3392 gnd.n3278 9.3005
R12008 gnd.n3394 gnd.n3393 9.3005
R12009 gnd.n3269 gnd.n3268 9.3005
R12010 gnd.n3407 gnd.n3406 9.3005
R12011 gnd.n3408 gnd.n3267 9.3005
R12012 gnd.n3410 gnd.n3409 9.3005
R12013 gnd.n3256 gnd.n3255 9.3005
R12014 gnd.n3453 gnd.n3452 9.3005
R12015 gnd.n3454 gnd.n3210 9.3005
R12016 gnd.n3458 gnd.n3456 9.3005
R12017 gnd.n3457 gnd.n3189 9.3005
R12018 gnd.n3476 gnd.n3188 9.3005
R12019 gnd.n3479 gnd.n3478 9.3005
R12020 gnd.n3182 gnd.n3181 9.3005
R12021 gnd.n3490 gnd.n3488 9.3005
R12022 gnd.n3489 gnd.n3163 9.3005
R12023 gnd.n3507 gnd.n3162 9.3005
R12024 gnd.n3510 gnd.n3509 9.3005
R12025 gnd.n3157 gnd.n3152 9.3005
R12026 gnd.n3520 gnd.n3519 9.3005
R12027 gnd.n3155 gnd.n3133 9.3005
R12028 gnd.n3547 gnd.n3134 9.3005
R12029 gnd.n3546 gnd.n3545 9.3005
R12030 gnd.n3136 gnd.n3121 9.3005
R12031 gnd.n3564 gnd.n3563 9.3005
R12032 gnd.n3566 gnd.n3099 9.3005
R12033 gnd.n3595 gnd.n3100 9.3005
R12034 gnd.n3594 gnd.n3101 9.3005
R12035 gnd.n3593 gnd.n3102 9.3005
R12036 gnd.n3105 gnd.n3104 9.3005
R12037 gnd.n2939 gnd.n2938 9.3005
R12038 gnd.n3615 gnd.n3613 9.3005
R12039 gnd.n3614 gnd.n2923 9.3005
R12040 gnd.n3632 gnd.n2922 9.3005
R12041 gnd.n3635 gnd.n3634 9.3005
R12042 gnd.n2916 gnd.n2915 9.3005
R12043 gnd.n3646 gnd.n3644 9.3005
R12044 gnd.n3645 gnd.n2898 9.3005
R12045 gnd.n3663 gnd.n2897 9.3005
R12046 gnd.n3666 gnd.n3665 9.3005
R12047 gnd.n2890 gnd.n2889 9.3005
R12048 gnd.n3677 gnd.n3675 9.3005
R12049 gnd.n3676 gnd.n2871 9.3005
R12050 gnd.n3694 gnd.n2870 9.3005
R12051 gnd.n3697 gnd.n3696 9.3005
R12052 gnd.n2864 gnd.n2863 9.3005
R12053 gnd.n3708 gnd.n3706 9.3005
R12054 gnd.n3707 gnd.n2847 9.3005
R12055 gnd.n3725 gnd.n2846 9.3005
R12056 gnd.n3728 gnd.n3727 9.3005
R12057 gnd.n2840 gnd.n2839 9.3005
R12058 gnd.n3739 gnd.n3737 9.3005
R12059 gnd.n3738 gnd.n2821 9.3005
R12060 gnd.n3756 gnd.n2820 9.3005
R12061 gnd.n3759 gnd.n3758 9.3005
R12062 gnd.n2814 gnd.n2813 9.3005
R12063 gnd.n3770 gnd.n3768 9.3005
R12064 gnd.n3769 gnd.n2796 9.3005
R12065 gnd.n3787 gnd.n2795 9.3005
R12066 gnd.n4046 gnd.n4045 9.3005
R12067 gnd.n2788 gnd.n2787 9.3005
R12068 gnd.n4056 gnd.n4055 9.3005
R12069 gnd.n2770 gnd.n2769 9.3005
R12070 gnd.n4074 gnd.n4073 9.3005
R12071 gnd.n3280 gnd.n3279 9.3005
R12072 gnd.n2551 gnd.n2550 9.3005
R12073 gnd.n2549 gnd.n1603 9.3005
R12074 gnd.n2548 gnd.n2547 9.3005
R12075 gnd.n1605 gnd.n1604 9.3005
R12076 gnd.n2541 gnd.n1609 9.3005
R12077 gnd.n2540 gnd.n1610 9.3005
R12078 gnd.n2539 gnd.n1611 9.3005
R12079 gnd.n1616 gnd.n1612 9.3005
R12080 gnd.n2533 gnd.n1617 9.3005
R12081 gnd.n2532 gnd.n1618 9.3005
R12082 gnd.n2531 gnd.n1619 9.3005
R12083 gnd.n1624 gnd.n1620 9.3005
R12084 gnd.n2525 gnd.n1625 9.3005
R12085 gnd.n2524 gnd.n1626 9.3005
R12086 gnd.n2523 gnd.n1627 9.3005
R12087 gnd.n1632 gnd.n1628 9.3005
R12088 gnd.n2517 gnd.n1633 9.3005
R12089 gnd.n2516 gnd.n1634 9.3005
R12090 gnd.n2515 gnd.n1635 9.3005
R12091 gnd.n1640 gnd.n1636 9.3005
R12092 gnd.n2509 gnd.n1641 9.3005
R12093 gnd.n2508 gnd.n1642 9.3005
R12094 gnd.n2507 gnd.n1643 9.3005
R12095 gnd.n1648 gnd.n1644 9.3005
R12096 gnd.n2501 gnd.n1649 9.3005
R12097 gnd.n2500 gnd.n1650 9.3005
R12098 gnd.n2499 gnd.n1651 9.3005
R12099 gnd.n1656 gnd.n1652 9.3005
R12100 gnd.n2493 gnd.n1657 9.3005
R12101 gnd.n2492 gnd.n1658 9.3005
R12102 gnd.n2491 gnd.n1659 9.3005
R12103 gnd.n1664 gnd.n1660 9.3005
R12104 gnd.n2485 gnd.n1665 9.3005
R12105 gnd.n2484 gnd.n1666 9.3005
R12106 gnd.n2483 gnd.n1667 9.3005
R12107 gnd.n1672 gnd.n1668 9.3005
R12108 gnd.n2477 gnd.n1673 9.3005
R12109 gnd.n2476 gnd.n1674 9.3005
R12110 gnd.n2475 gnd.n1675 9.3005
R12111 gnd.n1680 gnd.n1676 9.3005
R12112 gnd.n2469 gnd.n1681 9.3005
R12113 gnd.n2468 gnd.n1682 9.3005
R12114 gnd.n2467 gnd.n1683 9.3005
R12115 gnd.n1688 gnd.n1684 9.3005
R12116 gnd.n2461 gnd.n1689 9.3005
R12117 gnd.n2460 gnd.n1690 9.3005
R12118 gnd.n2459 gnd.n1691 9.3005
R12119 gnd.n1696 gnd.n1692 9.3005
R12120 gnd.n2453 gnd.n1697 9.3005
R12121 gnd.n2452 gnd.n1698 9.3005
R12122 gnd.n2451 gnd.n1699 9.3005
R12123 gnd.n1704 gnd.n1700 9.3005
R12124 gnd.n2445 gnd.n1705 9.3005
R12125 gnd.n2444 gnd.n1706 9.3005
R12126 gnd.n2443 gnd.n1707 9.3005
R12127 gnd.n1712 gnd.n1708 9.3005
R12128 gnd.n2437 gnd.n1713 9.3005
R12129 gnd.n2436 gnd.n1714 9.3005
R12130 gnd.n2435 gnd.n1715 9.3005
R12131 gnd.n1720 gnd.n1716 9.3005
R12132 gnd.n2429 gnd.n1721 9.3005
R12133 gnd.n2428 gnd.n1722 9.3005
R12134 gnd.n2427 gnd.n1723 9.3005
R12135 gnd.n1728 gnd.n1724 9.3005
R12136 gnd.n2421 gnd.n1729 9.3005
R12137 gnd.n2420 gnd.n1730 9.3005
R12138 gnd.n2419 gnd.n1731 9.3005
R12139 gnd.n1736 gnd.n1732 9.3005
R12140 gnd.n2413 gnd.n1737 9.3005
R12141 gnd.n2412 gnd.n1738 9.3005
R12142 gnd.n2411 gnd.n1739 9.3005
R12143 gnd.n1744 gnd.n1740 9.3005
R12144 gnd.n2405 gnd.n1745 9.3005
R12145 gnd.n2404 gnd.n1746 9.3005
R12146 gnd.n2403 gnd.n1747 9.3005
R12147 gnd.n1752 gnd.n1748 9.3005
R12148 gnd.n2397 gnd.n1753 9.3005
R12149 gnd.n2396 gnd.n1754 9.3005
R12150 gnd.n2395 gnd.n1755 9.3005
R12151 gnd.n1760 gnd.n1756 9.3005
R12152 gnd.n2389 gnd.n1761 9.3005
R12153 gnd.n2388 gnd.n1762 9.3005
R12154 gnd.n2387 gnd.n1763 9.3005
R12155 gnd.n1768 gnd.n1764 9.3005
R12156 gnd.n2381 gnd.n1769 9.3005
R12157 gnd.n2380 gnd.n1770 9.3005
R12158 gnd.n2379 gnd.n1771 9.3005
R12159 gnd.n1776 gnd.n1772 9.3005
R12160 gnd.n2373 gnd.n1777 9.3005
R12161 gnd.n2372 gnd.n1778 9.3005
R12162 gnd.n2371 gnd.n1779 9.3005
R12163 gnd.n1784 gnd.n1780 9.3005
R12164 gnd.n2365 gnd.n1785 9.3005
R12165 gnd.n2364 gnd.n1786 9.3005
R12166 gnd.n2363 gnd.n1787 9.3005
R12167 gnd.n1792 gnd.n1788 9.3005
R12168 gnd.n2357 gnd.n1793 9.3005
R12169 gnd.n2356 gnd.n1794 9.3005
R12170 gnd.n2355 gnd.n1795 9.3005
R12171 gnd.n1800 gnd.n1796 9.3005
R12172 gnd.n2349 gnd.n1801 9.3005
R12173 gnd.n2348 gnd.n1802 9.3005
R12174 gnd.n2347 gnd.n1803 9.3005
R12175 gnd.n1808 gnd.n1804 9.3005
R12176 gnd.n2341 gnd.n1809 9.3005
R12177 gnd.n2340 gnd.n1810 9.3005
R12178 gnd.n2339 gnd.n1811 9.3005
R12179 gnd.n1816 gnd.n1812 9.3005
R12180 gnd.n2333 gnd.n1817 9.3005
R12181 gnd.n2332 gnd.n1818 9.3005
R12182 gnd.n2331 gnd.n1819 9.3005
R12183 gnd.n1824 gnd.n1820 9.3005
R12184 gnd.n2325 gnd.n1825 9.3005
R12185 gnd.n2324 gnd.n1826 9.3005
R12186 gnd.n2323 gnd.n1827 9.3005
R12187 gnd.n1832 gnd.n1828 9.3005
R12188 gnd.n2317 gnd.n1833 9.3005
R12189 gnd.n2316 gnd.n1834 9.3005
R12190 gnd.n2315 gnd.n1835 9.3005
R12191 gnd.n1840 gnd.n1836 9.3005
R12192 gnd.n2309 gnd.n1841 9.3005
R12193 gnd.n2308 gnd.n1842 9.3005
R12194 gnd.n2307 gnd.n1843 9.3005
R12195 gnd.n1848 gnd.n1844 9.3005
R12196 gnd.n2301 gnd.n1849 9.3005
R12197 gnd.n2300 gnd.n1850 9.3005
R12198 gnd.n2299 gnd.n1851 9.3005
R12199 gnd.n1856 gnd.n1852 9.3005
R12200 gnd.n2293 gnd.n1857 9.3005
R12201 gnd.n2292 gnd.n1858 9.3005
R12202 gnd.n2291 gnd.n1859 9.3005
R12203 gnd.n1864 gnd.n1860 9.3005
R12204 gnd.n2285 gnd.n1865 9.3005
R12205 gnd.n2284 gnd.n1866 9.3005
R12206 gnd.n2283 gnd.n1867 9.3005
R12207 gnd.n1872 gnd.n1868 9.3005
R12208 gnd.n2277 gnd.n1873 9.3005
R12209 gnd.n2276 gnd.n1874 9.3005
R12210 gnd.n2275 gnd.n1875 9.3005
R12211 gnd.n1880 gnd.n1876 9.3005
R12212 gnd.n2269 gnd.n1881 9.3005
R12213 gnd.n2268 gnd.n1882 9.3005
R12214 gnd.n2267 gnd.n1883 9.3005
R12215 gnd.n1888 gnd.n1884 9.3005
R12216 gnd.n2261 gnd.n1889 9.3005
R12217 gnd.n2260 gnd.n1890 9.3005
R12218 gnd.n2259 gnd.n1891 9.3005
R12219 gnd.n1896 gnd.n1892 9.3005
R12220 gnd.n2253 gnd.n1897 9.3005
R12221 gnd.n2252 gnd.n1898 9.3005
R12222 gnd.n2251 gnd.n1899 9.3005
R12223 gnd.n1904 gnd.n1900 9.3005
R12224 gnd.n2245 gnd.n1905 9.3005
R12225 gnd.n2244 gnd.n1906 9.3005
R12226 gnd.n2243 gnd.n1907 9.3005
R12227 gnd.n2237 gnd.n2236 9.3005
R12228 gnd.n2235 gnd.n1912 9.3005
R12229 gnd.n2234 gnd.n2233 9.3005
R12230 gnd.n1915 gnd.n1914 9.3005
R12231 gnd.n2227 gnd.n1919 9.3005
R12232 gnd.n2226 gnd.n1920 9.3005
R12233 gnd.n2225 gnd.n1921 9.3005
R12234 gnd.n1926 gnd.n1922 9.3005
R12235 gnd.n2219 gnd.n1927 9.3005
R12236 gnd.n2218 gnd.n1928 9.3005
R12237 gnd.n2217 gnd.n1929 9.3005
R12238 gnd.n1934 gnd.n1930 9.3005
R12239 gnd.n2211 gnd.n1935 9.3005
R12240 gnd.n2210 gnd.n1936 9.3005
R12241 gnd.n2209 gnd.n1937 9.3005
R12242 gnd.n1942 gnd.n1938 9.3005
R12243 gnd.n2203 gnd.n1943 9.3005
R12244 gnd.n2202 gnd.n1944 9.3005
R12245 gnd.n2201 gnd.n1945 9.3005
R12246 gnd.n1950 gnd.n1946 9.3005
R12247 gnd.n2195 gnd.n1951 9.3005
R12248 gnd.n2194 gnd.n1952 9.3005
R12249 gnd.n2193 gnd.n1953 9.3005
R12250 gnd.n1958 gnd.n1954 9.3005
R12251 gnd.n2187 gnd.n1959 9.3005
R12252 gnd.n2186 gnd.n1960 9.3005
R12253 gnd.n2185 gnd.n1961 9.3005
R12254 gnd.n1966 gnd.n1962 9.3005
R12255 gnd.n2179 gnd.n1967 9.3005
R12256 gnd.n2178 gnd.n1968 9.3005
R12257 gnd.n2177 gnd.n1969 9.3005
R12258 gnd.n1974 gnd.n1970 9.3005
R12259 gnd.n2171 gnd.n1975 9.3005
R12260 gnd.n2170 gnd.n1976 9.3005
R12261 gnd.n2169 gnd.n1977 9.3005
R12262 gnd.n1982 gnd.n1978 9.3005
R12263 gnd.n2163 gnd.n1983 9.3005
R12264 gnd.n2162 gnd.n1984 9.3005
R12265 gnd.n2161 gnd.n1985 9.3005
R12266 gnd.n1990 gnd.n1986 9.3005
R12267 gnd.n2155 gnd.n1991 9.3005
R12268 gnd.n2154 gnd.n1992 9.3005
R12269 gnd.n2153 gnd.n1993 9.3005
R12270 gnd.n1998 gnd.n1994 9.3005
R12271 gnd.n2147 gnd.n1999 9.3005
R12272 gnd.n2146 gnd.n2000 9.3005
R12273 gnd.n2145 gnd.n2001 9.3005
R12274 gnd.n2006 gnd.n2002 9.3005
R12275 gnd.n2139 gnd.n2007 9.3005
R12276 gnd.n2138 gnd.n2008 9.3005
R12277 gnd.n2137 gnd.n2009 9.3005
R12278 gnd.n2014 gnd.n2010 9.3005
R12279 gnd.n2131 gnd.n2015 9.3005
R12280 gnd.n2130 gnd.n2016 9.3005
R12281 gnd.n2129 gnd.n2017 9.3005
R12282 gnd.n2022 gnd.n2018 9.3005
R12283 gnd.n2123 gnd.n2023 9.3005
R12284 gnd.n2122 gnd.n2024 9.3005
R12285 gnd.n2121 gnd.n2025 9.3005
R12286 gnd.n2030 gnd.n2026 9.3005
R12287 gnd.n2115 gnd.n2031 9.3005
R12288 gnd.n2114 gnd.n2032 9.3005
R12289 gnd.n2113 gnd.n2033 9.3005
R12290 gnd.n2038 gnd.n2034 9.3005
R12291 gnd.n2107 gnd.n2039 9.3005
R12292 gnd.n2106 gnd.n2040 9.3005
R12293 gnd.n2105 gnd.n2041 9.3005
R12294 gnd.n2046 gnd.n2042 9.3005
R12295 gnd.n2099 gnd.n2047 9.3005
R12296 gnd.n2098 gnd.n2048 9.3005
R12297 gnd.n2097 gnd.n2049 9.3005
R12298 gnd.n2054 gnd.n2050 9.3005
R12299 gnd.n2091 gnd.n2055 9.3005
R12300 gnd.n2090 gnd.n2056 9.3005
R12301 gnd.n2089 gnd.n2057 9.3005
R12302 gnd.n2062 gnd.n2058 9.3005
R12303 gnd.n2083 gnd.n2063 9.3005
R12304 gnd.n2082 gnd.n2064 9.3005
R12305 gnd.n2081 gnd.n2065 9.3005
R12306 gnd.n2071 gnd.n2066 9.3005
R12307 gnd.n2075 gnd.n2072 9.3005
R12308 gnd.n2074 gnd.n2073 9.3005
R12309 gnd.n345 gnd.n344 9.3005
R12310 gnd.n7079 gnd.n7078 9.3005
R12311 gnd.n1913 gnd.n1911 9.3005
R12312 gnd.n7427 gnd.n130 9.3005
R12313 gnd.n7426 gnd.n132 9.3005
R12314 gnd.n136 gnd.n133 9.3005
R12315 gnd.n7421 gnd.n137 9.3005
R12316 gnd.n7420 gnd.n138 9.3005
R12317 gnd.n7419 gnd.n139 9.3005
R12318 gnd.n143 gnd.n140 9.3005
R12319 gnd.n7414 gnd.n144 9.3005
R12320 gnd.n7413 gnd.n145 9.3005
R12321 gnd.n7412 gnd.n146 9.3005
R12322 gnd.n150 gnd.n147 9.3005
R12323 gnd.n7407 gnd.n151 9.3005
R12324 gnd.n7406 gnd.n152 9.3005
R12325 gnd.n7405 gnd.n153 9.3005
R12326 gnd.n157 gnd.n154 9.3005
R12327 gnd.n7400 gnd.n158 9.3005
R12328 gnd.n7399 gnd.n159 9.3005
R12329 gnd.n7395 gnd.n160 9.3005
R12330 gnd.n164 gnd.n161 9.3005
R12331 gnd.n7390 gnd.n165 9.3005
R12332 gnd.n7389 gnd.n166 9.3005
R12333 gnd.n7388 gnd.n167 9.3005
R12334 gnd.n171 gnd.n168 9.3005
R12335 gnd.n7383 gnd.n172 9.3005
R12336 gnd.n7382 gnd.n173 9.3005
R12337 gnd.n7381 gnd.n174 9.3005
R12338 gnd.n178 gnd.n175 9.3005
R12339 gnd.n7376 gnd.n179 9.3005
R12340 gnd.n7375 gnd.n180 9.3005
R12341 gnd.n7374 gnd.n181 9.3005
R12342 gnd.n185 gnd.n182 9.3005
R12343 gnd.n7369 gnd.n186 9.3005
R12344 gnd.n7368 gnd.n187 9.3005
R12345 gnd.n7367 gnd.n188 9.3005
R12346 gnd.n192 gnd.n189 9.3005
R12347 gnd.n7362 gnd.n193 9.3005
R12348 gnd.n7361 gnd.n7360 9.3005
R12349 gnd.n7359 gnd.n196 9.3005
R12350 gnd.n7429 gnd.n7428 9.3005
R12351 gnd.n6704 gnd.n6703 9.3005
R12352 gnd.n6708 gnd.n6705 9.3005
R12353 gnd.n6709 gnd.n6702 9.3005
R12354 gnd.n6713 gnd.n6712 9.3005
R12355 gnd.n6714 gnd.n6701 9.3005
R12356 gnd.n6723 gnd.n6715 9.3005
R12357 gnd.n6722 gnd.n6716 9.3005
R12358 gnd.n6721 gnd.n6718 9.3005
R12359 gnd.n6717 gnd.n596 9.3005
R12360 gnd.n6748 gnd.n597 9.3005
R12361 gnd.n6749 gnd.n595 9.3005
R12362 gnd.n6753 gnd.n6752 9.3005
R12363 gnd.n6754 gnd.n594 9.3005
R12364 gnd.n6762 gnd.n6755 9.3005
R12365 gnd.n6761 gnd.n6756 9.3005
R12366 gnd.n6760 gnd.n6757 9.3005
R12367 gnd.n587 gnd.n586 9.3005
R12368 gnd.n6780 gnd.n6779 9.3005
R12369 gnd.n6781 gnd.n585 9.3005
R12370 gnd.n6796 gnd.n6782 9.3005
R12371 gnd.n6795 gnd.n6783 9.3005
R12372 gnd.n6794 gnd.n6784 9.3005
R12373 gnd.n6793 gnd.n6785 9.3005
R12374 gnd.n6792 gnd.n6786 9.3005
R12375 gnd.n6789 gnd.n6788 9.3005
R12376 gnd.n6787 gnd.n357 9.3005
R12377 gnd.n7053 gnd.n356 9.3005
R12378 gnd.n7055 gnd.n7054 9.3005
R12379 gnd.n7056 gnd.n355 9.3005
R12380 gnd.n7060 gnd.n7057 9.3005
R12381 gnd.n7059 gnd.n7058 9.3005
R12382 gnd.n334 gnd.n333 9.3005
R12383 gnd.n7091 gnd.n7090 9.3005
R12384 gnd.n7092 gnd.n332 9.3005
R12385 gnd.n7159 gnd.n7093 9.3005
R12386 gnd.n7158 gnd.n7094 9.3005
R12387 gnd.n7157 gnd.n7095 9.3005
R12388 gnd.n7155 gnd.n7096 9.3005
R12389 gnd.n7154 gnd.n7097 9.3005
R12390 gnd.n7152 gnd.n7098 9.3005
R12391 gnd.n7151 gnd.n7099 9.3005
R12392 gnd.n7149 gnd.n7100 9.3005
R12393 gnd.n7148 gnd.n7101 9.3005
R12394 gnd.n7146 gnd.n7102 9.3005
R12395 gnd.n7145 gnd.n7103 9.3005
R12396 gnd.n7143 gnd.n7104 9.3005
R12397 gnd.n7142 gnd.n7105 9.3005
R12398 gnd.n7140 gnd.n7106 9.3005
R12399 gnd.n7139 gnd.n7107 9.3005
R12400 gnd.n7137 gnd.n7108 9.3005
R12401 gnd.n7136 gnd.n7109 9.3005
R12402 gnd.n7134 gnd.n7110 9.3005
R12403 gnd.n7133 gnd.n7111 9.3005
R12404 gnd.n7131 gnd.n7112 9.3005
R12405 gnd.n7130 gnd.n7113 9.3005
R12406 gnd.n7128 gnd.n7114 9.3005
R12407 gnd.n7127 gnd.n7115 9.3005
R12408 gnd.n7125 gnd.n7116 9.3005
R12409 gnd.n7124 gnd.n7117 9.3005
R12410 gnd.n7122 gnd.n7118 9.3005
R12411 gnd.n7121 gnd.n7120 9.3005
R12412 gnd.n7119 gnd.n200 9.3005
R12413 gnd.n7356 gnd.n199 9.3005
R12414 gnd.n7358 gnd.n7357 9.3005
R12415 gnd.n563 gnd.n562 9.3005
R12416 gnd.n6841 gnd.n6840 9.3005
R12417 gnd.n6842 gnd.n556 9.3005
R12418 gnd.n6845 gnd.n555 9.3005
R12419 gnd.n6846 gnd.n554 9.3005
R12420 gnd.n6849 gnd.n553 9.3005
R12421 gnd.n6850 gnd.n552 9.3005
R12422 gnd.n6853 gnd.n551 9.3005
R12423 gnd.n6854 gnd.n550 9.3005
R12424 gnd.n6857 gnd.n549 9.3005
R12425 gnd.n6858 gnd.n548 9.3005
R12426 gnd.n6861 gnd.n547 9.3005
R12427 gnd.n6862 gnd.n546 9.3005
R12428 gnd.n6865 gnd.n545 9.3005
R12429 gnd.n6866 gnd.n544 9.3005
R12430 gnd.n6869 gnd.n543 9.3005
R12431 gnd.n6870 gnd.n542 9.3005
R12432 gnd.n6873 gnd.n541 9.3005
R12433 gnd.n6874 gnd.n540 9.3005
R12434 gnd.n6877 gnd.n539 9.3005
R12435 gnd.n6879 gnd.n533 9.3005
R12436 gnd.n6882 gnd.n532 9.3005
R12437 gnd.n6883 gnd.n531 9.3005
R12438 gnd.n6886 gnd.n530 9.3005
R12439 gnd.n6887 gnd.n529 9.3005
R12440 gnd.n6890 gnd.n528 9.3005
R12441 gnd.n6891 gnd.n527 9.3005
R12442 gnd.n6894 gnd.n526 9.3005
R12443 gnd.n6895 gnd.n525 9.3005
R12444 gnd.n6898 gnd.n524 9.3005
R12445 gnd.n6899 gnd.n523 9.3005
R12446 gnd.n6902 gnd.n522 9.3005
R12447 gnd.n6903 gnd.n521 9.3005
R12448 gnd.n6904 gnd.n520 9.3005
R12449 gnd.n487 gnd.n486 9.3005
R12450 gnd.n6910 gnd.n6909 9.3005
R12451 gnd.n6839 gnd.n561 9.3005
R12452 gnd.n6838 gnd.n6837 9.3005
R12453 gnd.n6913 gnd.n6912 9.3005
R12454 gnd.n469 gnd.n468 9.3005
R12455 gnd.n6926 gnd.n6925 9.3005
R12456 gnd.n6927 gnd.n467 9.3005
R12457 gnd.n6929 gnd.n6928 9.3005
R12458 gnd.n452 gnd.n451 9.3005
R12459 gnd.n6942 gnd.n6941 9.3005
R12460 gnd.n6943 gnd.n450 9.3005
R12461 gnd.n6945 gnd.n6944 9.3005
R12462 gnd.n435 gnd.n434 9.3005
R12463 gnd.n6958 gnd.n6957 9.3005
R12464 gnd.n6959 gnd.n433 9.3005
R12465 gnd.n6961 gnd.n6960 9.3005
R12466 gnd.n418 gnd.n417 9.3005
R12467 gnd.n6974 gnd.n6973 9.3005
R12468 gnd.n6975 gnd.n416 9.3005
R12469 gnd.n6977 gnd.n6976 9.3005
R12470 gnd.n399 gnd.n398 9.3005
R12471 gnd.n6993 gnd.n6992 9.3005
R12472 gnd.n6994 gnd.n397 9.3005
R12473 gnd.n6996 gnd.n6995 9.3005
R12474 gnd.n367 gnd.n366 9.3005
R12475 gnd.n7044 gnd.n7043 9.3005
R12476 gnd.n7045 gnd.n365 9.3005
R12477 gnd.n7047 gnd.n7046 9.3005
R12478 gnd.n7048 gnd.n299 9.3005
R12479 gnd.n7187 gnd.n7186 9.3005
R12480 gnd.n284 gnd.n283 9.3005
R12481 gnd.n7200 gnd.n7199 9.3005
R12482 gnd.n7201 gnd.n282 9.3005
R12483 gnd.n7203 gnd.n7202 9.3005
R12484 gnd.n270 gnd.n269 9.3005
R12485 gnd.n7216 gnd.n7215 9.3005
R12486 gnd.n7217 gnd.n268 9.3005
R12487 gnd.n7219 gnd.n7218 9.3005
R12488 gnd.n254 gnd.n253 9.3005
R12489 gnd.n7232 gnd.n7231 9.3005
R12490 gnd.n7233 gnd.n252 9.3005
R12491 gnd.n7235 gnd.n7234 9.3005
R12492 gnd.n240 gnd.n239 9.3005
R12493 gnd.n7248 gnd.n7247 9.3005
R12494 gnd.n7249 gnd.n238 9.3005
R12495 gnd.n7251 gnd.n7250 9.3005
R12496 gnd.n223 gnd.n222 9.3005
R12497 gnd.n7264 gnd.n7263 9.3005
R12498 gnd.n7265 gnd.n221 9.3005
R12499 gnd.n7267 gnd.n7266 9.3005
R12500 gnd.n207 gnd.n206 9.3005
R12501 gnd.n7348 gnd.n7347 9.3005
R12502 gnd.n7349 gnd.n205 9.3005
R12503 gnd.n7351 gnd.n7350 9.3005
R12504 gnd.n129 gnd.n128 9.3005
R12505 gnd.n7431 gnd.n7430 9.3005
R12506 gnd.n6911 gnd.n485 9.3005
R12507 gnd.n7185 gnd.n298 9.3005
R12508 gnd.n7008 gnd.n346 9.3005
R12509 gnd.n7075 gnd.n347 9.3005
R12510 gnd.n7077 gnd.n7076 9.3005
R12511 gnd.n4848 gnd.n1215 9.3005
R12512 gnd.n4670 gnd.n1216 9.3005
R12513 gnd.n4672 gnd.n4671 9.3005
R12514 gnd.n4673 gnd.n4669 9.3005
R12515 gnd.n4685 gnd.n4674 9.3005
R12516 gnd.n4684 gnd.n4675 9.3005
R12517 gnd.n4683 gnd.n4676 9.3005
R12518 gnd.n4680 gnd.n4677 9.3005
R12519 gnd.n4679 gnd.n4678 9.3005
R12520 gnd.n1260 gnd.n1259 9.3005
R12521 gnd.n4712 gnd.n4711 9.3005
R12522 gnd.n4713 gnd.n1258 9.3005
R12523 gnd.n4725 gnd.n4714 9.3005
R12524 gnd.n4724 gnd.n4715 9.3005
R12525 gnd.n4723 gnd.n4716 9.3005
R12526 gnd.n4720 gnd.n4717 9.3005
R12527 gnd.n4719 gnd.n4718 9.3005
R12528 gnd.n1250 gnd.n1249 9.3005
R12529 gnd.n4751 gnd.n4750 9.3005
R12530 gnd.n4752 gnd.n1248 9.3005
R12531 gnd.n4785 gnd.n4753 9.3005
R12532 gnd.n4784 gnd.n4754 9.3005
R12533 gnd.n4783 gnd.n4755 9.3005
R12534 gnd.n4758 gnd.n4756 9.3005
R12535 gnd.n4779 gnd.n4759 9.3005
R12536 gnd.n4778 gnd.n4760 9.3005
R12537 gnd.n4777 gnd.n4761 9.3005
R12538 gnd.n4765 gnd.n4762 9.3005
R12539 gnd.n4772 gnd.n4766 9.3005
R12540 gnd.n4771 gnd.n4767 9.3005
R12541 gnd.n4770 gnd.n4768 9.3005
R12542 gnd.n941 gnd.n940 9.3005
R12543 gnd.n6340 gnd.n6339 9.3005
R12544 gnd.n6341 gnd.n939 9.3005
R12545 gnd.n6343 gnd.n6342 9.3005
R12546 gnd.n927 gnd.n926 9.3005
R12547 gnd.n6356 gnd.n6355 9.3005
R12548 gnd.n6357 gnd.n925 9.3005
R12549 gnd.n6359 gnd.n6358 9.3005
R12550 gnd.n913 gnd.n912 9.3005
R12551 gnd.n6372 gnd.n6371 9.3005
R12552 gnd.n6373 gnd.n911 9.3005
R12553 gnd.n6375 gnd.n6374 9.3005
R12554 gnd.n898 gnd.n897 9.3005
R12555 gnd.n6388 gnd.n6387 9.3005
R12556 gnd.n6389 gnd.n896 9.3005
R12557 gnd.n6391 gnd.n6390 9.3005
R12558 gnd.n883 gnd.n882 9.3005
R12559 gnd.n6404 gnd.n6403 9.3005
R12560 gnd.n6405 gnd.n881 9.3005
R12561 gnd.n6407 gnd.n6406 9.3005
R12562 gnd.n867 gnd.n866 9.3005
R12563 gnd.n6420 gnd.n6419 9.3005
R12564 gnd.n6421 gnd.n865 9.3005
R12565 gnd.n6423 gnd.n6422 9.3005
R12566 gnd.n852 gnd.n851 9.3005
R12567 gnd.n6436 gnd.n6435 9.3005
R12568 gnd.n6437 gnd.n850 9.3005
R12569 gnd.n6439 gnd.n6438 9.3005
R12570 gnd.n838 gnd.n837 9.3005
R12571 gnd.n6452 gnd.n6451 9.3005
R12572 gnd.n6453 gnd.n836 9.3005
R12573 gnd.n6455 gnd.n6454 9.3005
R12574 gnd.n823 gnd.n822 9.3005
R12575 gnd.n6468 gnd.n6467 9.3005
R12576 gnd.n6469 gnd.n821 9.3005
R12577 gnd.n6471 gnd.n6470 9.3005
R12578 gnd.n807 gnd.n806 9.3005
R12579 gnd.n6484 gnd.n6483 9.3005
R12580 gnd.n6485 gnd.n805 9.3005
R12581 gnd.n6487 gnd.n6486 9.3005
R12582 gnd.n792 gnd.n791 9.3005
R12583 gnd.n6500 gnd.n6499 9.3005
R12584 gnd.n6501 gnd.n790 9.3005
R12585 gnd.n6503 gnd.n6502 9.3005
R12586 gnd.n777 gnd.n776 9.3005
R12587 gnd.n6516 gnd.n6515 9.3005
R12588 gnd.n6517 gnd.n775 9.3005
R12589 gnd.n6519 gnd.n6518 9.3005
R12590 gnd.n761 gnd.n760 9.3005
R12591 gnd.n6532 gnd.n6531 9.3005
R12592 gnd.n6533 gnd.n759 9.3005
R12593 gnd.n6535 gnd.n6534 9.3005
R12594 gnd.n745 gnd.n744 9.3005
R12595 gnd.n6548 gnd.n6547 9.3005
R12596 gnd.n6549 gnd.n743 9.3005
R12597 gnd.n6551 gnd.n6550 9.3005
R12598 gnd.n731 gnd.n730 9.3005
R12599 gnd.n6564 gnd.n6563 9.3005
R12600 gnd.n6565 gnd.n729 9.3005
R12601 gnd.n6567 gnd.n6566 9.3005
R12602 gnd.n716 gnd.n715 9.3005
R12603 gnd.n6580 gnd.n6579 9.3005
R12604 gnd.n6581 gnd.n714 9.3005
R12605 gnd.n6583 gnd.n6582 9.3005
R12606 gnd.n701 gnd.n700 9.3005
R12607 gnd.n6596 gnd.n6595 9.3005
R12608 gnd.n6597 gnd.n699 9.3005
R12609 gnd.n6599 gnd.n6598 9.3005
R12610 gnd.n687 gnd.n686 9.3005
R12611 gnd.n6612 gnd.n6611 9.3005
R12612 gnd.n6613 gnd.n685 9.3005
R12613 gnd.n6615 gnd.n6614 9.3005
R12614 gnd.n673 gnd.n672 9.3005
R12615 gnd.n6628 gnd.n6627 9.3005
R12616 gnd.n6629 gnd.n671 9.3005
R12617 gnd.n6631 gnd.n6630 9.3005
R12618 gnd.n659 gnd.n658 9.3005
R12619 gnd.n6644 gnd.n6643 9.3005
R12620 gnd.n6645 gnd.n657 9.3005
R12621 gnd.n6647 gnd.n6646 9.3005
R12622 gnd.n644 gnd.n643 9.3005
R12623 gnd.n6661 gnd.n6660 9.3005
R12624 gnd.n6662 gnd.n642 9.3005
R12625 gnd.n6666 gnd.n6663 9.3005
R12626 gnd.n6665 gnd.n6664 9.3005
R12627 gnd.n614 gnd.n613 9.3005
R12628 gnd.n6680 gnd.n6679 9.3005
R12629 gnd.n6681 gnd.n612 9.3005
R12630 gnd.n6683 gnd.n6682 9.3005
R12631 gnd.n610 gnd.n609 9.3005
R12632 gnd.n6688 gnd.n6687 9.3005
R12633 gnd.n6689 gnd.n608 9.3005
R12634 gnd.n6691 gnd.n6690 9.3005
R12635 gnd.n606 gnd.n605 9.3005
R12636 gnd.n6696 gnd.n6695 9.3005
R12637 gnd.n6697 gnd.n604 9.3005
R12638 gnd.n6699 gnd.n6698 9.3005
R12639 gnd.n602 gnd.n601 9.3005
R12640 gnd.n6730 gnd.n6729 9.3005
R12641 gnd.n6731 gnd.n600 9.3005
R12642 gnd.n6743 gnd.n6732 9.3005
R12643 gnd.n6742 gnd.n6733 9.3005
R12644 gnd.n6741 gnd.n6734 9.3005
R12645 gnd.n6738 gnd.n6735 9.3005
R12646 gnd.n6737 gnd.n6736 9.3005
R12647 gnd.n592 gnd.n591 9.3005
R12648 gnd.n6769 gnd.n6768 9.3005
R12649 gnd.n6770 gnd.n590 9.3005
R12650 gnd.n6774 gnd.n6771 9.3005
R12651 gnd.n6773 gnd.n6772 9.3005
R12652 gnd.n392 gnd.n391 9.3005
R12653 gnd.n7002 gnd.n7001 9.3005
R12654 gnd.n7003 gnd.n390 9.3005
R12655 gnd.n7016 gnd.n7004 9.3005
R12656 gnd.n7015 gnd.n7005 9.3005
R12657 gnd.n7014 gnd.n7006 9.3005
R12658 gnd.n7011 gnd.n7007 9.3005
R12659 gnd.n7010 gnd.n7009 9.3005
R12660 gnd.n4622 gnd.n4621 9.3005
R12661 gnd.n4282 gnd.n4239 9.3005
R12662 gnd.n4281 gnd.n4240 9.3005
R12663 gnd.n4280 gnd.n4241 9.3005
R12664 gnd.n4278 gnd.n4242 9.3005
R12665 gnd.n4277 gnd.n4243 9.3005
R12666 gnd.n4275 gnd.n4244 9.3005
R12667 gnd.n4274 gnd.n4245 9.3005
R12668 gnd.n4272 gnd.n4246 9.3005
R12669 gnd.n4271 gnd.n4247 9.3005
R12670 gnd.n4269 gnd.n4248 9.3005
R12671 gnd.n4268 gnd.n4249 9.3005
R12672 gnd.n4266 gnd.n4250 9.3005
R12673 gnd.n4265 gnd.n4251 9.3005
R12674 gnd.n4263 gnd.n4252 9.3005
R12675 gnd.n4262 gnd.n4253 9.3005
R12676 gnd.n4260 gnd.n4254 9.3005
R12677 gnd.n4259 gnd.n4255 9.3005
R12678 gnd.n4257 gnd.n4256 9.3005
R12679 gnd.n1318 gnd.n1317 9.3005
R12680 gnd.n4575 gnd.n4574 9.3005
R12681 gnd.n4576 gnd.n1316 9.3005
R12682 gnd.n4583 gnd.n4577 9.3005
R12683 gnd.n4582 gnd.n4578 9.3005
R12684 gnd.n4581 gnd.n4579 9.3005
R12685 gnd.n1283 gnd.n1282 9.3005
R12686 gnd.n4614 gnd.n4613 9.3005
R12687 gnd.n4615 gnd.n1281 9.3005
R12688 gnd.n4627 gnd.n4616 9.3005
R12689 gnd.n4626 gnd.n4617 9.3005
R12690 gnd.n4625 gnd.n4618 9.3005
R12691 gnd.n4623 gnd.n4619 9.3005
R12692 gnd.n4238 gnd.n4171 9.3005
R12693 gnd.n4231 gnd.n4230 9.3005
R12694 gnd.n4229 gnd.n4177 9.3005
R12695 gnd.n4228 gnd.n4227 9.3005
R12696 gnd.n4179 gnd.n4178 9.3005
R12697 gnd.n4221 gnd.n4220 9.3005
R12698 gnd.n4219 gnd.n4181 9.3005
R12699 gnd.n4218 gnd.n4217 9.3005
R12700 gnd.n4183 gnd.n4182 9.3005
R12701 gnd.n4211 gnd.n4210 9.3005
R12702 gnd.n4209 gnd.n4185 9.3005
R12703 gnd.n4208 gnd.n4207 9.3005
R12704 gnd.n4187 gnd.n4186 9.3005
R12705 gnd.n4201 gnd.n4200 9.3005
R12706 gnd.n4199 gnd.n4189 9.3005
R12707 gnd.n4198 gnd.n4197 9.3005
R12708 gnd.n4192 gnd.n4190 9.3005
R12709 gnd.n4191 gnd.n1398 9.3005
R12710 gnd.n4175 gnd.n4172 9.3005
R12711 gnd.n4237 gnd.n4236 9.3005
R12712 gnd.n4486 gnd.n1397 9.3005
R12713 gnd.n4488 gnd.n4487 9.3005
R12714 gnd.n1384 gnd.n1383 9.3005
R12715 gnd.n4501 gnd.n4500 9.3005
R12716 gnd.n4502 gnd.n1382 9.3005
R12717 gnd.n4504 gnd.n4503 9.3005
R12718 gnd.n1367 gnd.n1366 9.3005
R12719 gnd.n4517 gnd.n4516 9.3005
R12720 gnd.n4518 gnd.n1365 9.3005
R12721 gnd.n4520 gnd.n4519 9.3005
R12722 gnd.n1352 gnd.n1351 9.3005
R12723 gnd.n4533 gnd.n4532 9.3005
R12724 gnd.n4534 gnd.n1350 9.3005
R12725 gnd.n4536 gnd.n4535 9.3005
R12726 gnd.n1335 gnd.n1334 9.3005
R12727 gnd.n4549 gnd.n4548 9.3005
R12728 gnd.n4550 gnd.n1333 9.3005
R12729 gnd.n4560 gnd.n4551 9.3005
R12730 gnd.n4559 gnd.n4552 9.3005
R12731 gnd.n4558 gnd.n4553 9.3005
R12732 gnd.n4557 gnd.n4555 9.3005
R12733 gnd.n4554 gnd.n1299 9.3005
R12734 gnd.n4600 gnd.n1300 9.3005
R12735 gnd.n4599 gnd.n1301 9.3005
R12736 gnd.n4598 gnd.n1302 9.3005
R12737 gnd.n1308 gnd.n1303 9.3005
R12738 gnd.n1307 gnd.n1305 9.3005
R12739 gnd.n1304 gnd.n1190 9.3005
R12740 gnd.n4874 gnd.n1191 9.3005
R12741 gnd.n4873 gnd.n1192 9.3005
R12742 gnd.n4872 gnd.n1193 9.3005
R12743 gnd.n1273 gnd.n1194 9.3005
R12744 gnd.n4860 gnd.n1204 9.3005
R12745 gnd.n4859 gnd.n1205 9.3005
R12746 gnd.n4858 gnd.n1206 9.3005
R12747 gnd.n1168 gnd.n1167 9.3005
R12748 gnd.n4887 gnd.n4886 9.3005
R12749 gnd.n4888 gnd.n1166 9.3005
R12750 gnd.n4890 gnd.n4889 9.3005
R12751 gnd.n1152 gnd.n1151 9.3005
R12752 gnd.n4903 gnd.n4902 9.3005
R12753 gnd.n4904 gnd.n1150 9.3005
R12754 gnd.n4906 gnd.n4905 9.3005
R12755 gnd.n1134 gnd.n1133 9.3005
R12756 gnd.n4919 gnd.n4918 9.3005
R12757 gnd.n4920 gnd.n1132 9.3005
R12758 gnd.n4922 gnd.n4921 9.3005
R12759 gnd.n1118 gnd.n1117 9.3005
R12760 gnd.n4935 gnd.n4934 9.3005
R12761 gnd.n4936 gnd.n1116 9.3005
R12762 gnd.n4938 gnd.n4937 9.3005
R12763 gnd.n1100 gnd.n1099 9.3005
R12764 gnd.n4951 gnd.n4950 9.3005
R12765 gnd.n4952 gnd.n1098 9.3005
R12766 gnd.n4954 gnd.n4953 9.3005
R12767 gnd.n1084 gnd.n1083 9.3005
R12768 gnd.n4967 gnd.n4966 9.3005
R12769 gnd.n4968 gnd.n1082 9.3005
R12770 gnd.n4970 gnd.n4969 9.3005
R12771 gnd.n1065 gnd.n1064 9.3005
R12772 gnd.n4985 gnd.n4984 9.3005
R12773 gnd.n4986 gnd.n1063 9.3005
R12774 gnd.n6223 gnd.n4987 9.3005
R12775 gnd.n6222 gnd.n6221 9.3005
R12776 gnd.n4485 gnd.n4484 9.3005
R12777 gnd.n1020 gnd.n1014 9.3005
R12778 gnd.n6273 gnd.n1013 9.3005
R12779 gnd.n6274 gnd.n1012 9.3005
R12780 gnd.n6275 gnd.n1011 9.3005
R12781 gnd.n1010 gnd.n1007 9.3005
R12782 gnd.n6280 gnd.n1006 9.3005
R12783 gnd.n6281 gnd.n1005 9.3005
R12784 gnd.n6282 gnd.n1004 9.3005
R12785 gnd.n1003 gnd.n1000 9.3005
R12786 gnd.n6287 gnd.n999 9.3005
R12787 gnd.n6288 gnd.n998 9.3005
R12788 gnd.n6289 gnd.n997 9.3005
R12789 gnd.n996 gnd.n993 9.3005
R12790 gnd.n995 gnd.n991 9.3005
R12791 gnd.n6296 gnd.n990 9.3005
R12792 gnd.n6298 gnd.n6297 9.3005
R12793 gnd.n6265 gnd.n1023 9.3005
R12794 gnd.n6264 gnd.n1024 9.3005
R12795 gnd.n1028 gnd.n1025 9.3005
R12796 gnd.n6259 gnd.n1029 9.3005
R12797 gnd.n6258 gnd.n1030 9.3005
R12798 gnd.n6257 gnd.n1031 9.3005
R12799 gnd.n1035 gnd.n1032 9.3005
R12800 gnd.n6252 gnd.n1036 9.3005
R12801 gnd.n6251 gnd.n1037 9.3005
R12802 gnd.n6250 gnd.n1038 9.3005
R12803 gnd.n1042 gnd.n1039 9.3005
R12804 gnd.n6245 gnd.n1043 9.3005
R12805 gnd.n6244 gnd.n1044 9.3005
R12806 gnd.n6243 gnd.n1045 9.3005
R12807 gnd.n1049 gnd.n1046 9.3005
R12808 gnd.n6238 gnd.n1050 9.3005
R12809 gnd.n6237 gnd.n1051 9.3005
R12810 gnd.n6236 gnd.n1052 9.3005
R12811 gnd.n1057 gnd.n1055 9.3005
R12812 gnd.n6231 gnd.n6230 9.3005
R12813 gnd.n6266 gnd.n1022 9.3005
R12814 gnd.n4397 gnd.n4347 9.3005
R12815 gnd.n4396 gnd.n4349 9.3005
R12816 gnd.n4395 gnd.n4350 9.3005
R12817 gnd.n4393 gnd.n4351 9.3005
R12818 gnd.n4392 gnd.n4352 9.3005
R12819 gnd.n4390 gnd.n4353 9.3005
R12820 gnd.n4389 gnd.n4354 9.3005
R12821 gnd.n4387 gnd.n4355 9.3005
R12822 gnd.n4386 gnd.n4356 9.3005
R12823 gnd.n4384 gnd.n4357 9.3005
R12824 gnd.n4383 gnd.n4358 9.3005
R12825 gnd.n4381 gnd.n4359 9.3005
R12826 gnd.n4380 gnd.n4360 9.3005
R12827 gnd.n4378 gnd.n4361 9.3005
R12828 gnd.n4377 gnd.n4362 9.3005
R12829 gnd.n4375 gnd.n4363 9.3005
R12830 gnd.n4374 gnd.n4364 9.3005
R12831 gnd.n4372 gnd.n4365 9.3005
R12832 gnd.n4371 gnd.n4366 9.3005
R12833 gnd.n4369 gnd.n4368 9.3005
R12834 gnd.n4367 gnd.n1312 9.3005
R12835 gnd.n4587 gnd.n1311 9.3005
R12836 gnd.n4589 gnd.n4588 9.3005
R12837 gnd.n4590 gnd.n1310 9.3005
R12838 gnd.n4594 gnd.n4591 9.3005
R12839 gnd.n4593 gnd.n4592 9.3005
R12840 gnd.n1277 gnd.n1276 9.3005
R12841 gnd.n4632 gnd.n4631 9.3005
R12842 gnd.n4633 gnd.n1275 9.3005
R12843 gnd.n4636 gnd.n4634 9.3005
R12844 gnd.n4637 gnd.n1274 9.3005
R12845 gnd.n4640 gnd.n4639 9.3005
R12846 gnd.n4641 gnd.n1272 9.3005
R12847 gnd.n4643 gnd.n4642 9.3005
R12848 gnd.n1268 gnd.n1267 9.3005
R12849 gnd.n4656 gnd.n4655 9.3005
R12850 gnd.n4657 gnd.n1266 9.3005
R12851 gnd.n4659 gnd.n4658 9.3005
R12852 gnd.n4660 gnd.n1265 9.3005
R12853 gnd.n4664 gnd.n4663 9.3005
R12854 gnd.n4665 gnd.n1264 9.3005
R12855 gnd.n4690 gnd.n4666 9.3005
R12856 gnd.n4691 gnd.n1263 9.3005
R12857 gnd.n4695 gnd.n4694 9.3005
R12858 gnd.n4696 gnd.n1262 9.3005
R12859 gnd.n4705 gnd.n4697 9.3005
R12860 gnd.n4704 gnd.n4698 9.3005
R12861 gnd.n4703 gnd.n4700 9.3005
R12862 gnd.n4699 gnd.n1254 9.3005
R12863 gnd.n4730 gnd.n1255 9.3005
R12864 gnd.n4731 gnd.n1253 9.3005
R12865 gnd.n4735 gnd.n4734 9.3005
R12866 gnd.n4736 gnd.n1252 9.3005
R12867 gnd.n4744 gnd.n4737 9.3005
R12868 gnd.n4743 gnd.n4738 9.3005
R12869 gnd.n4742 gnd.n4739 9.3005
R12870 gnd.n1245 gnd.n1244 9.3005
R12871 gnd.n4791 gnd.n4790 9.3005
R12872 gnd.n4792 gnd.n1243 9.3005
R12873 gnd.n4797 gnd.n4793 9.3005
R12874 gnd.n4796 gnd.n4795 9.3005
R12875 gnd.n4794 gnd.n1059 9.3005
R12876 gnd.n6227 gnd.n1058 9.3005
R12877 gnd.n6229 gnd.n6228 9.3005
R12878 gnd.n4399 gnd.n4398 9.3005
R12879 gnd.n4407 gnd.n4406 9.3005
R12880 gnd.n4408 gnd.n4341 9.3005
R12881 gnd.n4409 gnd.n4340 9.3005
R12882 gnd.n4339 gnd.n4337 9.3005
R12883 gnd.n4415 gnd.n4336 9.3005
R12884 gnd.n4416 gnd.n4335 9.3005
R12885 gnd.n4417 gnd.n4334 9.3005
R12886 gnd.n4333 gnd.n4331 9.3005
R12887 gnd.n4423 gnd.n4330 9.3005
R12888 gnd.n4424 gnd.n4329 9.3005
R12889 gnd.n4425 gnd.n4328 9.3005
R12890 gnd.n4327 gnd.n4325 9.3005
R12891 gnd.n4431 gnd.n4324 9.3005
R12892 gnd.n4432 gnd.n4323 9.3005
R12893 gnd.n4433 gnd.n4322 9.3005
R12894 gnd.n4321 gnd.n4319 9.3005
R12895 gnd.n4439 gnd.n4318 9.3005
R12896 gnd.n4440 gnd.n4317 9.3005
R12897 gnd.n4441 gnd.n4316 9.3005
R12898 gnd.n4315 gnd.n4310 9.3005
R12899 gnd.n4447 gnd.n4309 9.3005
R12900 gnd.n4448 gnd.n4308 9.3005
R12901 gnd.n4449 gnd.n4307 9.3005
R12902 gnd.n4306 gnd.n4304 9.3005
R12903 gnd.n4455 gnd.n4303 9.3005
R12904 gnd.n4456 gnd.n4302 9.3005
R12905 gnd.n4457 gnd.n4301 9.3005
R12906 gnd.n4300 gnd.n4298 9.3005
R12907 gnd.n4463 gnd.n4297 9.3005
R12908 gnd.n4464 gnd.n4296 9.3005
R12909 gnd.n4465 gnd.n4295 9.3005
R12910 gnd.n4294 gnd.n4292 9.3005
R12911 gnd.n4470 gnd.n4291 9.3005
R12912 gnd.n4471 gnd.n4290 9.3005
R12913 gnd.n4289 gnd.n4287 9.3005
R12914 gnd.n4476 gnd.n4286 9.3005
R12915 gnd.n4478 gnd.n4477 9.3005
R12916 gnd.n4405 gnd.n4346 9.3005
R12917 gnd.n4404 gnd.n4403 9.3005
R12918 gnd.n1392 gnd.n1391 9.3005
R12919 gnd.n4493 gnd.n4492 9.3005
R12920 gnd.n4494 gnd.n1390 9.3005
R12921 gnd.n4496 gnd.n4495 9.3005
R12922 gnd.n1376 gnd.n1375 9.3005
R12923 gnd.n4509 gnd.n4508 9.3005
R12924 gnd.n4510 gnd.n1374 9.3005
R12925 gnd.n4512 gnd.n4511 9.3005
R12926 gnd.n1360 gnd.n1359 9.3005
R12927 gnd.n4525 gnd.n4524 9.3005
R12928 gnd.n4526 gnd.n1358 9.3005
R12929 gnd.n4528 gnd.n4527 9.3005
R12930 gnd.n1344 gnd.n1343 9.3005
R12931 gnd.n4541 gnd.n4540 9.3005
R12932 gnd.n4542 gnd.n1342 9.3005
R12933 gnd.n4544 gnd.n4543 9.3005
R12934 gnd.n1327 gnd.n1326 9.3005
R12935 gnd.n4565 gnd.n4564 9.3005
R12936 gnd.n4566 gnd.n1325 9.3005
R12937 gnd.n4570 gnd.n4567 9.3005
R12938 gnd.n4569 gnd.n4568 9.3005
R12939 gnd.n1291 gnd.n1290 9.3005
R12940 gnd.n4605 gnd.n4604 9.3005
R12941 gnd.n4606 gnd.n1289 9.3005
R12942 gnd.n4608 gnd.n4607 9.3005
R12943 gnd.n4609 gnd.n1176 9.3005
R12944 gnd.n1160 gnd.n1159 9.3005
R12945 gnd.n4895 gnd.n4894 9.3005
R12946 gnd.n4896 gnd.n1158 9.3005
R12947 gnd.n4898 gnd.n4897 9.3005
R12948 gnd.n1143 gnd.n1142 9.3005
R12949 gnd.n4911 gnd.n4910 9.3005
R12950 gnd.n4912 gnd.n1141 9.3005
R12951 gnd.n4914 gnd.n4913 9.3005
R12952 gnd.n1126 gnd.n1125 9.3005
R12953 gnd.n4927 gnd.n4926 9.3005
R12954 gnd.n4928 gnd.n1124 9.3005
R12955 gnd.n4930 gnd.n4929 9.3005
R12956 gnd.n1109 gnd.n1108 9.3005
R12957 gnd.n4943 gnd.n4942 9.3005
R12958 gnd.n4944 gnd.n1107 9.3005
R12959 gnd.n4946 gnd.n4945 9.3005
R12960 gnd.n1092 gnd.n1091 9.3005
R12961 gnd.n4959 gnd.n4958 9.3005
R12962 gnd.n4960 gnd.n1090 9.3005
R12963 gnd.n4962 gnd.n4961 9.3005
R12964 gnd.n1075 gnd.n1074 9.3005
R12965 gnd.n4975 gnd.n4974 9.3005
R12966 gnd.n4976 gnd.n1073 9.3005
R12967 gnd.n4980 gnd.n4977 9.3005
R12968 gnd.n4979 gnd.n4978 9.3005
R12969 gnd.n989 gnd.n988 9.3005
R12970 gnd.n6300 gnd.n6299 9.3005
R12971 gnd.n4480 gnd.n4479 9.3005
R12972 gnd.n4882 gnd.n4881 9.3005
R12973 gnd.n4850 gnd.n1213 9.3005
R12974 gnd.n4849 gnd.n1214 9.3005
R12975 gnd.n2761 gnd.n1212 9.3005
R12976 gnd.n2764 gnd.n2760 9.3005
R12977 gnd.n2759 gnd.n1477 9.3005
R12978 gnd.n2758 gnd.n2757 9.3005
R12979 gnd.n1479 gnd.n1478 9.3005
R12980 gnd.n2751 gnd.n2750 9.3005
R12981 gnd.n2749 gnd.n1483 9.3005
R12982 gnd.n2748 gnd.n2747 9.3005
R12983 gnd.n1485 gnd.n1484 9.3005
R12984 gnd.n2741 gnd.n2740 9.3005
R12985 gnd.n2739 gnd.n1489 9.3005
R12986 gnd.n2738 gnd.n2737 9.3005
R12987 gnd.n1491 gnd.n1490 9.3005
R12988 gnd.n2731 gnd.n2730 9.3005
R12989 gnd.n2729 gnd.n1495 9.3005
R12990 gnd.n2728 gnd.n2727 9.3005
R12991 gnd.n1497 gnd.n1496 9.3005
R12992 gnd.n2721 gnd.n2720 9.3005
R12993 gnd.n2719 gnd.n1501 9.3005
R12994 gnd.n2718 gnd.n2717 9.3005
R12995 gnd.n1503 gnd.n1502 9.3005
R12996 gnd.n2711 gnd.n2710 9.3005
R12997 gnd.n2709 gnd.n1507 9.3005
R12998 gnd.n2708 gnd.n2707 9.3005
R12999 gnd.n1509 gnd.n1508 9.3005
R13000 gnd.n2701 gnd.n2700 9.3005
R13001 gnd.n2699 gnd.n1513 9.3005
R13002 gnd.n2698 gnd.n2697 9.3005
R13003 gnd.n1515 gnd.n1514 9.3005
R13004 gnd.n2691 gnd.n2690 9.3005
R13005 gnd.n2689 gnd.n1519 9.3005
R13006 gnd.n2688 gnd.n2687 9.3005
R13007 gnd.n1521 gnd.n1520 9.3005
R13008 gnd.n2681 gnd.n2680 9.3005
R13009 gnd.n2679 gnd.n1525 9.3005
R13010 gnd.n2678 gnd.n2677 9.3005
R13011 gnd.n1527 gnd.n1526 9.3005
R13012 gnd.n2671 gnd.n2670 9.3005
R13013 gnd.n2669 gnd.n1531 9.3005
R13014 gnd.n2668 gnd.n2667 9.3005
R13015 gnd.n1533 gnd.n1532 9.3005
R13016 gnd.n2661 gnd.n2660 9.3005
R13017 gnd.n2659 gnd.n1537 9.3005
R13018 gnd.n2658 gnd.n2657 9.3005
R13019 gnd.n1539 gnd.n1538 9.3005
R13020 gnd.n2651 gnd.n2650 9.3005
R13021 gnd.n2649 gnd.n1543 9.3005
R13022 gnd.n2648 gnd.n2647 9.3005
R13023 gnd.n1545 gnd.n1544 9.3005
R13024 gnd.n2641 gnd.n2640 9.3005
R13025 gnd.n2639 gnd.n1549 9.3005
R13026 gnd.n2638 gnd.n2637 9.3005
R13027 gnd.n1551 gnd.n1550 9.3005
R13028 gnd.n2631 gnd.n2630 9.3005
R13029 gnd.n2629 gnd.n1555 9.3005
R13030 gnd.n2628 gnd.n2627 9.3005
R13031 gnd.n1557 gnd.n1556 9.3005
R13032 gnd.n2621 gnd.n2620 9.3005
R13033 gnd.n2619 gnd.n1561 9.3005
R13034 gnd.n2618 gnd.n2617 9.3005
R13035 gnd.n1563 gnd.n1562 9.3005
R13036 gnd.n2611 gnd.n2610 9.3005
R13037 gnd.n2609 gnd.n1567 9.3005
R13038 gnd.n2608 gnd.n2607 9.3005
R13039 gnd.n1569 gnd.n1568 9.3005
R13040 gnd.n2601 gnd.n2600 9.3005
R13041 gnd.n2599 gnd.n1573 9.3005
R13042 gnd.n2598 gnd.n2597 9.3005
R13043 gnd.n1575 gnd.n1574 9.3005
R13044 gnd.n2591 gnd.n2590 9.3005
R13045 gnd.n2589 gnd.n1579 9.3005
R13046 gnd.n2588 gnd.n2587 9.3005
R13047 gnd.n1581 gnd.n1580 9.3005
R13048 gnd.n2581 gnd.n2580 9.3005
R13049 gnd.n2579 gnd.n1585 9.3005
R13050 gnd.n2578 gnd.n2577 9.3005
R13051 gnd.n1587 gnd.n1586 9.3005
R13052 gnd.n2571 gnd.n2570 9.3005
R13053 gnd.n2569 gnd.n1591 9.3005
R13054 gnd.n2568 gnd.n2567 9.3005
R13055 gnd.n1593 gnd.n1592 9.3005
R13056 gnd.n2561 gnd.n2560 9.3005
R13057 gnd.n2559 gnd.n1597 9.3005
R13058 gnd.n2558 gnd.n2557 9.3005
R13059 gnd.n1599 gnd.n1598 9.3005
R13060 gnd.n2763 gnd.n2762 9.3005
R13061 gnd.n5953 gnd.n5951 9.3005
R13062 gnd.n6086 gnd.n6085 9.3005
R13063 gnd.n6084 gnd.n6083 9.3005
R13064 gnd.n5970 gnd.n5969 9.3005
R13065 gnd.n6078 gnd.n6077 9.3005
R13066 gnd.n6076 gnd.n6075 9.3005
R13067 gnd.n5978 gnd.n5977 9.3005
R13068 gnd.n6070 gnd.n6069 9.3005
R13069 gnd.n6068 gnd.n6067 9.3005
R13070 gnd.n5990 gnd.n5989 9.3005
R13071 gnd.n6062 gnd.n6061 9.3005
R13072 gnd.n6060 gnd.n6059 9.3005
R13073 gnd.n5998 gnd.n5997 9.3005
R13074 gnd.n6054 gnd.n6053 9.3005
R13075 gnd.n6052 gnd.n6051 9.3005
R13076 gnd.n6010 gnd.n6009 9.3005
R13077 gnd.n6043 gnd.n6042 9.3005
R13078 gnd.n6041 gnd.n6011 9.3005
R13079 gnd.n6092 gnd.n6091 9.3005
R13080 gnd.n6004 gnd.n6003 9.3005
R13081 gnd.n6056 gnd.n6055 9.3005
R13082 gnd.n6058 gnd.n6057 9.3005
R13083 gnd.n5994 gnd.n5993 9.3005
R13084 gnd.n6064 gnd.n6063 9.3005
R13085 gnd.n6066 gnd.n6065 9.3005
R13086 gnd.n5984 gnd.n5983 9.3005
R13087 gnd.n6072 gnd.n6071 9.3005
R13088 gnd.n6074 gnd.n6073 9.3005
R13089 gnd.n5974 gnd.n5973 9.3005
R13090 gnd.n6080 gnd.n6079 9.3005
R13091 gnd.n6082 gnd.n6081 9.3005
R13092 gnd.n5964 gnd.n5963 9.3005
R13093 gnd.n6088 gnd.n6087 9.3005
R13094 gnd.n6090 gnd.n6089 9.3005
R13095 gnd.n5958 gnd.n5952 9.3005
R13096 gnd.n6050 gnd.n6049 9.3005
R13097 gnd.n6045 gnd.n6044 9.3005
R13098 gnd.n6040 gnd.n6039 9.3005
R13099 gnd.n6038 gnd.n6016 9.3005
R13100 gnd.n6037 gnd.n6036 9.3005
R13101 gnd.n6035 gnd.n6017 9.3005
R13102 gnd.n6034 gnd.n6033 9.3005
R13103 gnd.n6032 gnd.n6022 9.3005
R13104 gnd.n6031 gnd.n6030 9.3005
R13105 gnd.n6029 gnd.n6023 9.3005
R13106 gnd.n634 gnd.n633 9.3005
R13107 gnd.n6674 gnd.n6673 9.3005
R13108 gnd.n6348 gnd.n6347 9.3005
R13109 gnd.n6349 gnd.n932 9.3005
R13110 gnd.n6351 gnd.n6350 9.3005
R13111 gnd.n919 gnd.n918 9.3005
R13112 gnd.n6364 gnd.n6363 9.3005
R13113 gnd.n6365 gnd.n917 9.3005
R13114 gnd.n6367 gnd.n6366 9.3005
R13115 gnd.n905 gnd.n904 9.3005
R13116 gnd.n6380 gnd.n6379 9.3005
R13117 gnd.n6381 gnd.n903 9.3005
R13118 gnd.n6383 gnd.n6382 9.3005
R13119 gnd.n891 gnd.n890 9.3005
R13120 gnd.n6396 gnd.n6395 9.3005
R13121 gnd.n6397 gnd.n889 9.3005
R13122 gnd.n6399 gnd.n6398 9.3005
R13123 gnd.n875 gnd.n874 9.3005
R13124 gnd.n6412 gnd.n6411 9.3005
R13125 gnd.n6413 gnd.n873 9.3005
R13126 gnd.n6415 gnd.n6414 9.3005
R13127 gnd.n860 gnd.n859 9.3005
R13128 gnd.n6428 gnd.n6427 9.3005
R13129 gnd.n6429 gnd.n858 9.3005
R13130 gnd.n6431 gnd.n6430 9.3005
R13131 gnd.n845 gnd.n844 9.3005
R13132 gnd.n6444 gnd.n6443 9.3005
R13133 gnd.n6445 gnd.n843 9.3005
R13134 gnd.n6447 gnd.n6446 9.3005
R13135 gnd.n831 gnd.n830 9.3005
R13136 gnd.n6460 gnd.n6459 9.3005
R13137 gnd.n6461 gnd.n829 9.3005
R13138 gnd.n6463 gnd.n6462 9.3005
R13139 gnd.n815 gnd.n814 9.3005
R13140 gnd.n6476 gnd.n6475 9.3005
R13141 gnd.n6477 gnd.n813 9.3005
R13142 gnd.n6479 gnd.n6478 9.3005
R13143 gnd.n799 gnd.n798 9.3005
R13144 gnd.n6492 gnd.n6491 9.3005
R13145 gnd.n6493 gnd.n797 9.3005
R13146 gnd.n6495 gnd.n6494 9.3005
R13147 gnd.n784 gnd.n783 9.3005
R13148 gnd.n6508 gnd.n6507 9.3005
R13149 gnd.n6509 gnd.n782 9.3005
R13150 gnd.n6511 gnd.n6510 9.3005
R13151 gnd.n769 gnd.n768 9.3005
R13152 gnd.n6524 gnd.n6523 9.3005
R13153 gnd.n6525 gnd.n767 9.3005
R13154 gnd.n6527 gnd.n6526 9.3005
R13155 gnd.n753 gnd.n752 9.3005
R13156 gnd.n6540 gnd.n6539 9.3005
R13157 gnd.n6541 gnd.n751 9.3005
R13158 gnd.n6543 gnd.n6542 9.3005
R13159 gnd.n738 gnd.n737 9.3005
R13160 gnd.n6556 gnd.n6555 9.3005
R13161 gnd.n6557 gnd.n736 9.3005
R13162 gnd.n6559 gnd.n6558 9.3005
R13163 gnd.n724 gnd.n723 9.3005
R13164 gnd.n6572 gnd.n6571 9.3005
R13165 gnd.n6573 gnd.n722 9.3005
R13166 gnd.n6575 gnd.n6574 9.3005
R13167 gnd.n709 gnd.n708 9.3005
R13168 gnd.n6588 gnd.n6587 9.3005
R13169 gnd.n6589 gnd.n707 9.3005
R13170 gnd.n6591 gnd.n6590 9.3005
R13171 gnd.n694 gnd.n693 9.3005
R13172 gnd.n6604 gnd.n6603 9.3005
R13173 gnd.n6605 gnd.n692 9.3005
R13174 gnd.n6607 gnd.n6606 9.3005
R13175 gnd.n679 gnd.n678 9.3005
R13176 gnd.n6620 gnd.n6619 9.3005
R13177 gnd.n6621 gnd.n677 9.3005
R13178 gnd.n6623 gnd.n6622 9.3005
R13179 gnd.n666 gnd.n665 9.3005
R13180 gnd.n6636 gnd.n6635 9.3005
R13181 gnd.n6637 gnd.n664 9.3005
R13182 gnd.n6639 gnd.n6638 9.3005
R13183 gnd.n652 gnd.n651 9.3005
R13184 gnd.n6652 gnd.n6651 9.3005
R13185 gnd.n6653 gnd.n650 9.3005
R13186 gnd.n6656 gnd.n6655 9.3005
R13187 gnd.n6654 gnd.n636 9.3005
R13188 gnd.n6670 gnd.n635 9.3005
R13189 gnd.n6672 gnd.n6671 9.3005
R13190 gnd.n934 gnd.n933 9.3005
R13191 gnd.n6332 gnd.n959 9.3005
R13192 gnd.n6331 gnd.n6330 9.3005
R13193 gnd.n6327 gnd.n960 9.3005
R13194 gnd.n6325 gnd.n6324 9.3005
R13195 gnd.n6323 gnd.n963 9.3005
R13196 gnd.n6322 gnd.n6321 9.3005
R13197 gnd.n6318 gnd.n966 9.3005
R13198 gnd.n6317 gnd.n6316 9.3005
R13199 gnd.n6315 gnd.n967 9.3005
R13200 gnd.n6334 gnd.n6333 9.3005
R13201 gnd.n1271 gnd.n1270 9.3005
R13202 gnd.n4648 gnd.n4647 9.3005
R13203 gnd.n4649 gnd.n1269 9.3005
R13204 gnd.n4651 gnd.n4650 9.3005
R13205 gnd.n1221 gnd.n1219 9.3005
R13206 gnd.n4842 gnd.n4841 9.3005
R13207 gnd.n4840 gnd.n1220 9.3005
R13208 gnd.n4839 gnd.n4838 9.3005
R13209 gnd.n4837 gnd.n1222 9.3005
R13210 gnd.n4836 gnd.n4835 9.3005
R13211 gnd.n4834 gnd.n1225 9.3005
R13212 gnd.n4833 gnd.n4832 9.3005
R13213 gnd.n4831 gnd.n1226 9.3005
R13214 gnd.n4830 gnd.n4829 9.3005
R13215 gnd.n4828 gnd.n1229 9.3005
R13216 gnd.n4827 gnd.n4826 9.3005
R13217 gnd.n4825 gnd.n1230 9.3005
R13218 gnd.n4824 gnd.n4823 9.3005
R13219 gnd.n4822 gnd.n1233 9.3005
R13220 gnd.n4821 gnd.n4820 9.3005
R13221 gnd.n4819 gnd.n1234 9.3005
R13222 gnd.n4818 gnd.n4817 9.3005
R13223 gnd.n4816 gnd.n1237 9.3005
R13224 gnd.n4815 gnd.n4814 9.3005
R13225 gnd.n4813 gnd.n1238 9.3005
R13226 gnd.n4812 gnd.n4811 9.3005
R13227 gnd.n4810 gnd.n1241 9.3005
R13228 gnd.n4809 gnd.n4808 9.3005
R13229 gnd.n4807 gnd.n1242 9.3005
R13230 gnd.n4806 gnd.n4805 9.3005
R13231 gnd.n4804 gnd.n4803 9.3005
R13232 gnd.n981 gnd.n970 9.3005
R13233 gnd.n6313 gnd.n6312 9.3005
R13234 gnd.n6309 gnd.n971 9.3005
R13235 gnd.n6308 gnd.n6307 9.3005
R13236 gnd.n5053 gnd.n972 9.3005
R13237 gnd.n5046 gnd.n5045 9.3005
R13238 gnd.n5059 gnd.n5058 9.3005
R13239 gnd.n5061 gnd.n5060 9.3005
R13240 gnd.n5034 gnd.n5033 9.3005
R13241 gnd.n5067 gnd.n5066 9.3005
R13242 gnd.n5069 gnd.n5068 9.3005
R13243 gnd.n5023 gnd.n5022 9.3005
R13244 gnd.n5075 gnd.n5074 9.3005
R13245 gnd.n5077 gnd.n5076 9.3005
R13246 gnd.n5011 gnd.n5010 9.3005
R13247 gnd.n5083 gnd.n5082 9.3005
R13248 gnd.n5085 gnd.n5084 9.3005
R13249 gnd.n4996 gnd.n4994 9.3005
R13250 gnd.n5091 gnd.n5090 9.3005
R13251 gnd.n5092 gnd.n4991 9.3005
R13252 gnd.n4999 gnd.n4989 9.3005
R13253 gnd.n4997 gnd.n4995 9.3005
R13254 gnd.n5089 gnd.n5088 9.3005
R13255 gnd.n5087 gnd.n5086 9.3005
R13256 gnd.n5007 gnd.n5006 9.3005
R13257 gnd.n5081 gnd.n5080 9.3005
R13258 gnd.n5079 gnd.n5078 9.3005
R13259 gnd.n5017 gnd.n5016 9.3005
R13260 gnd.n5073 gnd.n5072 9.3005
R13261 gnd.n5071 gnd.n5070 9.3005
R13262 gnd.n5030 gnd.n5029 9.3005
R13263 gnd.n5065 gnd.n5064 9.3005
R13264 gnd.n5063 gnd.n5062 9.3005
R13265 gnd.n5040 gnd.n5039 9.3005
R13266 gnd.n5057 gnd.n5056 9.3005
R13267 gnd.n5055 gnd.n5054 9.3005
R13268 gnd.n978 gnd.n975 9.3005
R13269 gnd.n6306 gnd.n6305 9.3005
R13270 gnd.n6216 gnd.n4990 9.3005
R13271 gnd.n6215 gnd.n6214 9.3005
R13272 gnd.n6213 gnd.n5096 9.3005
R13273 gnd.n6212 gnd.n6211 9.3005
R13274 gnd.n6210 gnd.n5097 9.3005
R13275 gnd.n6209 gnd.n6208 9.3005
R13276 gnd.n6207 gnd.n5100 9.3005
R13277 gnd.n6206 gnd.n6205 9.3005
R13278 gnd.n6204 gnd.n5101 9.3005
R13279 gnd.n6203 gnd.n6202 9.3005
R13280 gnd.n6201 gnd.n5104 9.3005
R13281 gnd.n6200 gnd.n6199 9.3005
R13282 gnd.n6198 gnd.n5105 9.3005
R13283 gnd.n6197 gnd.n6196 9.3005
R13284 gnd.n6195 gnd.n5108 9.3005
R13285 gnd.n6194 gnd.n6193 9.3005
R13286 gnd.n6192 gnd.n5109 9.3005
R13287 gnd.n6191 gnd.n6190 9.3005
R13288 gnd.n6189 gnd.n5112 9.3005
R13289 gnd.n6188 gnd.n6187 9.3005
R13290 gnd.n6186 gnd.n5113 9.3005
R13291 gnd.n6185 gnd.n6184 9.3005
R13292 gnd.n6183 gnd.n5116 9.3005
R13293 gnd.n6182 gnd.n6181 9.3005
R13294 gnd.n6180 gnd.n5117 9.3005
R13295 gnd.n6179 gnd.n6178 9.3005
R13296 gnd.n6177 gnd.n5120 9.3005
R13297 gnd.n6176 gnd.n6175 9.3005
R13298 gnd.n6174 gnd.n5121 9.3005
R13299 gnd.n6173 gnd.n6172 9.3005
R13300 gnd.n6171 gnd.n5124 9.3005
R13301 gnd.n6170 gnd.n6169 9.3005
R13302 gnd.n6168 gnd.n5125 9.3005
R13303 gnd.n6167 gnd.n6166 9.3005
R13304 gnd.n6165 gnd.n5128 9.3005
R13305 gnd.n6164 gnd.n6163 9.3005
R13306 gnd.n6162 gnd.n5129 9.3005
R13307 gnd.n6161 gnd.n6160 9.3005
R13308 gnd.n6159 gnd.n5132 9.3005
R13309 gnd.n6158 gnd.n6157 9.3005
R13310 gnd.n6156 gnd.n5133 9.3005
R13311 gnd.n6155 gnd.n6154 9.3005
R13312 gnd.n6153 gnd.n5136 9.3005
R13313 gnd.n6152 gnd.n6151 9.3005
R13314 gnd.n6150 gnd.n5137 9.3005
R13315 gnd.n6149 gnd.n6148 9.3005
R13316 gnd.n6147 gnd.n5140 9.3005
R13317 gnd.n6146 gnd.n6145 9.3005
R13318 gnd.n6144 gnd.n5141 9.3005
R13319 gnd.n6143 gnd.n6142 9.3005
R13320 gnd.n6141 gnd.n5144 9.3005
R13321 gnd.n6140 gnd.n6139 9.3005
R13322 gnd.n6138 gnd.n5145 9.3005
R13323 gnd.n6137 gnd.n6136 9.3005
R13324 gnd.n6135 gnd.n5148 9.3005
R13325 gnd.n6134 gnd.n6133 9.3005
R13326 gnd.n6132 gnd.n5149 9.3005
R13327 gnd.n6131 gnd.n6130 9.3005
R13328 gnd.n6129 gnd.n5152 9.3005
R13329 gnd.n6128 gnd.n6127 9.3005
R13330 gnd.n6126 gnd.n5153 9.3005
R13331 gnd.n6125 gnd.n6124 9.3005
R13332 gnd.n6123 gnd.n5156 9.3005
R13333 gnd.n6122 gnd.n6121 9.3005
R13334 gnd.n6120 gnd.n5157 9.3005
R13335 gnd.n6119 gnd.n6118 9.3005
R13336 gnd.n6117 gnd.n5160 9.3005
R13337 gnd.n6116 gnd.n6115 9.3005
R13338 gnd.n6114 gnd.n5161 9.3005
R13339 gnd.n6113 gnd.n6112 9.3005
R13340 gnd.n6111 gnd.n5939 9.3005
R13341 gnd.n6110 gnd.n6109 9.3005
R13342 gnd.n6108 gnd.n5940 9.3005
R13343 gnd.n6107 gnd.n6106 9.3005
R13344 gnd.n6105 gnd.n5943 9.3005
R13345 gnd.n6104 gnd.n6103 9.3005
R13346 gnd.n6102 gnd.n5944 9.3005
R13347 gnd.n6101 gnd.n6100 9.3005
R13348 gnd.n6099 gnd.n5947 9.3005
R13349 gnd.n6098 gnd.n6097 9.3005
R13350 gnd.n6096 gnd.n5948 9.3005
R13351 gnd.n6095 gnd.n5950 9.3005
R13352 gnd.n6218 gnd.n6217 9.3005
R13353 gnd.n6918 gnd.n6917 9.3005
R13354 gnd.n6919 gnd.n476 9.3005
R13355 gnd.n6921 gnd.n6920 9.3005
R13356 gnd.n460 gnd.n459 9.3005
R13357 gnd.n6934 gnd.n6933 9.3005
R13358 gnd.n6935 gnd.n458 9.3005
R13359 gnd.n6937 gnd.n6936 9.3005
R13360 gnd.n444 gnd.n443 9.3005
R13361 gnd.n6950 gnd.n6949 9.3005
R13362 gnd.n6951 gnd.n442 9.3005
R13363 gnd.n6953 gnd.n6952 9.3005
R13364 gnd.n426 gnd.n425 9.3005
R13365 gnd.n6966 gnd.n6965 9.3005
R13366 gnd.n6967 gnd.n424 9.3005
R13367 gnd.n6969 gnd.n6968 9.3005
R13368 gnd.n410 gnd.n409 9.3005
R13369 gnd.n6982 gnd.n6981 9.3005
R13370 gnd.n6983 gnd.n407 9.3005
R13371 gnd.n6988 gnd.n6987 9.3005
R13372 gnd.n6986 gnd.n408 9.3005
R13373 gnd.n6985 gnd.n6984 9.3005
R13374 gnd.n377 gnd.n375 9.3005
R13375 gnd.n7039 gnd.n7038 9.3005
R13376 gnd.n7037 gnd.n376 9.3005
R13377 gnd.n7036 gnd.n7035 9.3005
R13378 gnd.n7034 gnd.n378 9.3005
R13379 gnd.n7033 gnd.n7032 9.3005
R13380 gnd.n316 gnd.n314 9.3005
R13381 gnd.n7178 gnd.n7177 9.3005
R13382 gnd.n7176 gnd.n315 9.3005
R13383 gnd.n7175 gnd.n7174 9.3005
R13384 gnd.n7173 gnd.n317 9.3005
R13385 gnd.n7172 gnd.n7171 9.3005
R13386 gnd.n7170 gnd.n321 9.3005
R13387 gnd.n7169 gnd.n7168 9.3005
R13388 gnd.n7167 gnd.n322 9.3005
R13389 gnd.n293 gnd.n292 9.3005
R13390 gnd.n7192 gnd.n7191 9.3005
R13391 gnd.n7193 gnd.n291 9.3005
R13392 gnd.n7195 gnd.n7194 9.3005
R13393 gnd.n277 gnd.n276 9.3005
R13394 gnd.n7208 gnd.n7207 9.3005
R13395 gnd.n7209 gnd.n275 9.3005
R13396 gnd.n7211 gnd.n7210 9.3005
R13397 gnd.n263 gnd.n262 9.3005
R13398 gnd.n7224 gnd.n7223 9.3005
R13399 gnd.n7225 gnd.n261 9.3005
R13400 gnd.n7227 gnd.n7226 9.3005
R13401 gnd.n247 gnd.n246 9.3005
R13402 gnd.n7240 gnd.n7239 9.3005
R13403 gnd.n7241 gnd.n245 9.3005
R13404 gnd.n7243 gnd.n7242 9.3005
R13405 gnd.n232 gnd.n231 9.3005
R13406 gnd.n7256 gnd.n7255 9.3005
R13407 gnd.n7257 gnd.n230 9.3005
R13408 gnd.n7259 gnd.n7258 9.3005
R13409 gnd.n217 gnd.n216 9.3005
R13410 gnd.n7272 gnd.n7271 9.3005
R13411 gnd.n7273 gnd.n214 9.3005
R13412 gnd.n7343 gnd.n7342 9.3005
R13413 gnd.n7341 gnd.n215 9.3005
R13414 gnd.n7340 gnd.n7339 9.3005
R13415 gnd.n7338 gnd.n7274 9.3005
R13416 gnd.n7337 gnd.n7336 9.3005
R13417 gnd.n478 gnd.n477 9.3005
R13418 gnd.n7333 gnd.n7276 9.3005
R13419 gnd.n7332 gnd.n7331 9.3005
R13420 gnd.n7330 gnd.n7281 9.3005
R13421 gnd.n7329 gnd.n7328 9.3005
R13422 gnd.n7327 gnd.n7282 9.3005
R13423 gnd.n7326 gnd.n7325 9.3005
R13424 gnd.n7324 gnd.n7289 9.3005
R13425 gnd.n7323 gnd.n7322 9.3005
R13426 gnd.n7321 gnd.n7290 9.3005
R13427 gnd.n7320 gnd.n7319 9.3005
R13428 gnd.n7318 gnd.n7297 9.3005
R13429 gnd.n7317 gnd.n7316 9.3005
R13430 gnd.n7315 gnd.n7298 9.3005
R13431 gnd.n7314 gnd.n7313 9.3005
R13432 gnd.n7312 gnd.n7305 9.3005
R13433 gnd.n7311 gnd.n7310 9.3005
R13434 gnd.n120 gnd.n117 9.3005
R13435 gnd.n7437 gnd.n7436 9.3005
R13436 gnd.n7335 gnd.n7334 9.3005
R13437 gnd.n6830 gnd.n565 9.3005
R13438 gnd.n6829 gnd.n6828 9.3005
R13439 gnd.n6827 gnd.n567 9.3005
R13440 gnd.n6826 gnd.n6825 9.3005
R13441 gnd.n6824 gnd.n570 9.3005
R13442 gnd.n6823 gnd.n6822 9.3005
R13443 gnd.n6821 gnd.n571 9.3005
R13444 gnd.n6820 gnd.n6819 9.3005
R13445 gnd.n6818 gnd.n574 9.3005
R13446 gnd.n6817 gnd.n6816 9.3005
R13447 gnd.n6815 gnd.n575 9.3005
R13448 gnd.n6814 gnd.n6813 9.3005
R13449 gnd.n6812 gnd.n578 9.3005
R13450 gnd.n6811 gnd.n6810 9.3005
R13451 gnd.n6809 gnd.n579 9.3005
R13452 gnd.n6808 gnd.n6807 9.3005
R13453 gnd.n6806 gnd.n582 9.3005
R13454 gnd.n6805 gnd.n6804 9.3005
R13455 gnd.n6803 gnd.n583 9.3005
R13456 gnd.n6802 gnd.n6801 9.3005
R13457 gnd.n6800 gnd.n384 9.3005
R13458 gnd.n7021 gnd.n383 9.3005
R13459 gnd.n7023 gnd.n7022 9.3005
R13460 gnd.n7024 gnd.n381 9.3005
R13461 gnd.n7027 gnd.n7026 9.3005
R13462 gnd.n7025 gnd.n382 9.3005
R13463 gnd.n354 gnd.n352 9.3005
R13464 gnd.n7069 gnd.n7068 9.3005
R13465 gnd.n7067 gnd.n353 9.3005
R13466 gnd.n7066 gnd.n7065 9.3005
R13467 gnd.n7064 gnd.n75 9.3005
R13468 gnd.n7486 gnd.n76 9.3005
R13469 gnd.n7485 gnd.n7484 9.3005
R13470 gnd.n7483 gnd.n77 9.3005
R13471 gnd.n7482 gnd.n7481 9.3005
R13472 gnd.n7480 gnd.n81 9.3005
R13473 gnd.n7479 gnd.n7478 9.3005
R13474 gnd.n7477 gnd.n82 9.3005
R13475 gnd.n7476 gnd.n7475 9.3005
R13476 gnd.n7474 gnd.n86 9.3005
R13477 gnd.n7473 gnd.n7472 9.3005
R13478 gnd.n7471 gnd.n87 9.3005
R13479 gnd.n7470 gnd.n7469 9.3005
R13480 gnd.n7468 gnd.n91 9.3005
R13481 gnd.n7467 gnd.n7466 9.3005
R13482 gnd.n7465 gnd.n92 9.3005
R13483 gnd.n7464 gnd.n7463 9.3005
R13484 gnd.n7462 gnd.n96 9.3005
R13485 gnd.n7461 gnd.n7460 9.3005
R13486 gnd.n7459 gnd.n97 9.3005
R13487 gnd.n7458 gnd.n7457 9.3005
R13488 gnd.n7456 gnd.n101 9.3005
R13489 gnd.n7455 gnd.n7454 9.3005
R13490 gnd.n7453 gnd.n102 9.3005
R13491 gnd.n7452 gnd.n7451 9.3005
R13492 gnd.n7450 gnd.n106 9.3005
R13493 gnd.n7449 gnd.n7448 9.3005
R13494 gnd.n7447 gnd.n107 9.3005
R13495 gnd.n7446 gnd.n7445 9.3005
R13496 gnd.n7444 gnd.n111 9.3005
R13497 gnd.n7443 gnd.n7442 9.3005
R13498 gnd.n7441 gnd.n112 9.3005
R13499 gnd.n7440 gnd.n7439 9.3005
R13500 gnd.n7438 gnd.n116 9.3005
R13501 gnd.n6832 gnd.n6831 9.3005
R13502 gnd.t24 gnd.n3679 9.24152
R13503 gnd.n4059 gnd.t61 9.24152
R13504 gnd.n2785 gnd.t82 9.24152
R13505 gnd.t217 gnd.n1337 9.24152
R13506 gnd.n4932 gnd.t178 9.24152
R13507 gnd.n6971 gnd.t192 9.24152
R13508 gnd.n259 gnd.t186 9.24152
R13509 gnd.t174 gnd.t24 8.92286
R13510 gnd.n6609 gnd.t116 8.92286
R13511 gnd.n4038 gnd.n4013 8.92171
R13512 gnd.n4006 gnd.n3981 8.92171
R13513 gnd.n3974 gnd.n3949 8.92171
R13514 gnd.n3943 gnd.n3918 8.92171
R13515 gnd.n3911 gnd.n3886 8.92171
R13516 gnd.n3879 gnd.n3854 8.92171
R13517 gnd.n3847 gnd.n3822 8.92171
R13518 gnd.n3816 gnd.n3791 8.92171
R13519 gnd.n5184 gnd.n5166 8.72777
R13520 gnd.n3025 gnd.t15 8.60421
R13521 gnd.t246 gnd.n1369 8.60421
R13522 gnd.n4964 gnd.t184 8.60421
R13523 gnd.n6939 gnd.t274 8.60421
R13524 gnd.n228 gnd.t271 8.60421
R13525 gnd.n3067 gnd.n3047 8.43467
R13526 gnd.n54 gnd.n34 8.43467
R13527 gnd.n4621 gnd.n0 8.41456
R13528 gnd.n7487 gnd.n7486 8.41456
R13529 gnd.n5351 gnd.t134 8.28555
R13530 gnd.t29 gnd.n856 8.28555
R13531 gnd.n5332 gnd.n5331 8.28555
R13532 gnd.n6489 gnd.n803 8.28555
R13533 gnd.n6521 gnd.n771 8.28555
R13534 gnd.n5746 gnd.n5265 8.28555
R13535 gnd.t162 gnd.n718 8.28555
R13536 gnd.n4039 gnd.n4011 8.14595
R13537 gnd.n4007 gnd.n3979 8.14595
R13538 gnd.n3975 gnd.n3947 8.14595
R13539 gnd.n3944 gnd.n3916 8.14595
R13540 gnd.n3912 gnd.n3884 8.14595
R13541 gnd.n3880 gnd.n3852 8.14595
R13542 gnd.n3848 gnd.n3820 8.14595
R13543 gnd.n3817 gnd.n3789 8.14595
R13544 gnd.n4044 gnd.n4043 7.97301
R13545 gnd.t17 gnd.n3579 7.9669
R13546 gnd.n7436 gnd.n120 7.75808
R13547 gnd.n6049 gnd.n6045 7.75808
R13548 gnd.n6305 gnd.n978 7.75808
R13549 gnd.n4236 gnd.n4175 7.75808
R13550 gnd.n4076 gnd.n2767 7.64824
R13551 gnd.n5576 gnd.t65 7.64824
R13552 gnd.n3512 gnd.t21 7.32958
R13553 gnd.n5427 gnd.n5426 7.30353
R13554 gnd.n5183 gnd.n5182 7.30353
R13555 gnd.n3472 gnd.n3191 7.01093
R13556 gnd.n3194 gnd.n3192 7.01093
R13557 gnd.n3482 gnd.n3481 7.01093
R13558 gnd.n3493 gnd.n3175 7.01093
R13559 gnd.n3492 gnd.n3178 7.01093
R13560 gnd.n3503 gnd.n3166 7.01093
R13561 gnd.n3169 gnd.n3167 7.01093
R13562 gnd.n3513 gnd.n3512 7.01093
R13563 gnd.n3523 gnd.n3147 7.01093
R13564 gnd.n3522 gnd.n3150 7.01093
R13565 gnd.n3539 gnd.n3140 7.01093
R13566 gnd.n3549 gnd.n3131 7.01093
R13567 gnd.n3560 gnd.n3559 7.01093
R13568 gnd.n3580 gnd.n3116 7.01093
R13569 gnd.n3579 gnd.n3095 7.01093
R13570 gnd.n3597 gnd.n3096 7.01093
R13571 gnd.n3591 gnd.n3590 7.01093
R13572 gnd.n3607 gnd.n2943 7.01093
R13573 gnd.n3617 gnd.n2935 7.01093
R13574 gnd.n3628 gnd.n2926 7.01093
R13575 gnd.n3025 gnd.n3024 7.01093
R13576 gnd.n3638 gnd.n3637 7.01093
R13577 gnd.n3649 gnd.n2909 7.01093
R13578 gnd.n3648 gnd.n2912 7.01093
R13579 gnd.n3659 gnd.n2901 7.01093
R13580 gnd.n3669 gnd.n3668 7.01093
R13581 gnd.n3680 gnd.n2883 7.01093
R13582 gnd.n3679 gnd.n2886 7.01093
R13583 gnd.n3690 gnd.n2874 7.01093
R13584 gnd.n2877 gnd.n2875 7.01093
R13585 gnd.n3700 gnd.n3699 7.01093
R13586 gnd.n3711 gnd.n2858 7.01093
R13587 gnd.n2852 gnd.n2850 7.01093
R13588 gnd.n3731 gnd.n3730 7.01093
R13589 gnd.n3742 gnd.n2833 7.01093
R13590 gnd.n3741 gnd.n2836 7.01093
R13591 gnd.n3752 gnd.n2824 7.01093
R13592 gnd.n2827 gnd.n2825 7.01093
R13593 gnd.n3773 gnd.n2807 7.01093
R13594 gnd.n3772 gnd.n2810 7.01093
R13595 gnd.n3783 gnd.n2799 7.01093
R13596 gnd.n2800 gnd.n2792 7.01093
R13597 gnd.n4049 gnd.n4048 7.01093
R13598 gnd.n4059 gnd.n2782 7.01093
R13599 gnd.n4058 gnd.n2785 7.01093
R13600 gnd.n4069 gnd.n2776 7.01093
R13601 gnd.n4076 gnd.n1400 7.01093
R13602 gnd.n5638 gnd.n5637 7.01093
R13603 gnd.n6481 gnd.n811 7.01093
R13604 gnd.n5313 gnd.t7 7.01093
R13605 gnd.n5286 gnd.t144 7.01093
R13606 gnd.n6529 gnd.n763 7.01093
R13607 gnd.n5738 gnd.n5271 7.01093
R13608 gnd.n5788 gnd.n5243 7.01093
R13609 gnd.n5803 gnd.t116 7.01093
R13610 gnd.n3150 gnd.t13 6.69227
R13611 gnd.n3680 gnd.t174 6.69227
R13612 gnd.n3762 gnd.t12 6.69227
R13613 gnd.n4787 gnd.t184 6.69227
R13614 gnd.t2 gnd.n5351 6.69227
R13615 gnd.t344 gnd.n5780 6.69227
R13616 gnd.n6726 gnd.t274 6.69227
R13617 gnd.n5863 gnd.n5862 6.5566
R13618 gnd.n5504 gnd.n5503 6.5566
R13619 gnd.n5489 gnd.n5488 6.5566
R13620 gnd.n5878 gnd.n5877 6.5566
R13621 gnd.n6327 gnd.n6326 6.20656
R13622 gnd.n7398 gnd.n7395 6.20656
R13623 gnd.n4441 gnd.n4314 6.20656
R13624 gnd.n6030 gnd.n6026 6.20656
R13625 gnd.t172 gnd.n3571 6.05496
R13626 gnd.n3572 gnd.t23 6.05496
R13627 gnd.n3637 gnd.t30 6.05496
R13628 gnd.n2999 gnd.t19 6.05496
R13629 gnd.n4727 gnd.t178 6.05496
R13630 gnd.n6765 gnd.t192 6.05496
R13631 gnd.n4041 gnd.n4011 5.81868
R13632 gnd.n4009 gnd.n3979 5.81868
R13633 gnd.n3977 gnd.n3947 5.81868
R13634 gnd.n3946 gnd.n3916 5.81868
R13635 gnd.n3914 gnd.n3884 5.81868
R13636 gnd.n3882 gnd.n3852 5.81868
R13637 gnd.n3850 gnd.n3820 5.81868
R13638 gnd.n3819 gnd.n3789 5.81868
R13639 gnd.n6401 gnd.n885 5.73631
R13640 gnd.n5576 gnd.n5361 5.73631
R13641 gnd.n5647 gnd.n5322 5.73631
R13642 gnd.n6473 gnd.n819 5.73631
R13643 gnd.n6537 gnd.n755 5.73631
R13644 gnd.n5729 gnd.n5276 5.73631
R13645 gnd.n5796 gnd.n5795 5.73631
R13646 gnd.n6609 gnd.n690 5.73631
R13647 gnd.n5210 gnd.n534 5.62001
R13648 gnd.n5497 gnd.n5496 5.62001
R13649 gnd.n5496 gnd.n5389 5.62001
R13650 gnd.n5872 gnd.n534 5.62001
R13651 gnd.n3331 gnd.n3326 5.4308
R13652 gnd.n4084 gnd.n1467 5.4308
R13653 gnd.n3649 gnd.t18 5.41765
R13654 gnd.t25 gnd.n2894 5.41765
R13655 gnd.n3721 gnd.t156 5.41765
R13656 gnd.n4845 gnd.t182 5.41765
R13657 gnd.n4687 gnd.t202 5.41765
R13658 gnd.n6441 gnd.t145 5.41765
R13659 gnd.n6569 gnd.t148 5.41765
R13660 gnd.n7018 gnd.t215 5.41765
R13661 gnd.t276 gnd.n359 5.41765
R13662 gnd.t134 gnd.n871 5.09899
R13663 gnd.n5346 gnd.t28 5.09899
R13664 gnd.n6457 gnd.t9 5.09899
R13665 gnd.t171 gnd.n827 5.09899
R13666 gnd.t147 gnd.n747 5.09899
R13667 gnd.n6553 gnd.t27 5.09899
R13668 gnd.n5773 gnd.t150 5.09899
R13669 gnd.t47 gnd.n681 5.09899
R13670 gnd.n4039 gnd.n4038 5.04292
R13671 gnd.n4007 gnd.n4006 5.04292
R13672 gnd.n3975 gnd.n3974 5.04292
R13673 gnd.n3944 gnd.n3943 5.04292
R13674 gnd.n3912 gnd.n3911 5.04292
R13675 gnd.n3880 gnd.n3879 5.04292
R13676 gnd.n3848 gnd.n3847 5.04292
R13677 gnd.n3817 gnd.n3816 5.04292
R13678 gnd.n3087 gnd.n3086 4.82753
R13679 gnd.n74 gnd.n73 4.82753
R13680 gnd.n3618 gnd.t10 4.78034
R13681 gnd.n2877 gnd.t16 4.78034
R13682 gnd.n4708 gnd.t227 4.78034
R13683 gnd.n6776 gnd.t258 4.78034
R13684 gnd.n3092 gnd.n3089 4.74817
R13685 gnd.n3604 gnd.n2945 4.74817
R13686 gnd.n3602 gnd.n2946 4.74817
R13687 gnd.n3028 gnd.n3022 4.74817
R13688 gnd.n3108 gnd.n3089 4.74817
R13689 gnd.n3107 gnd.n2945 4.74817
R13690 gnd.n3603 gnd.n3602 4.74817
R13691 gnd.n3028 gnd.n3027 4.74817
R13692 gnd.n7184 gnd.n7183 4.74817
R13693 gnd.n337 gnd.n304 4.74817
R13694 gnd.n7085 gnd.n303 4.74817
R13695 gnd.n327 gnd.n302 4.74817
R13696 gnd.n7163 gnd.n301 4.74817
R13697 gnd.n7184 gnd.n305 4.74817
R13698 gnd.n7182 gnd.n304 4.74817
R13699 gnd.n338 gnd.n303 4.74817
R13700 gnd.n7086 gnd.n302 4.74817
R13701 gnd.n328 gnd.n301 4.74817
R13702 gnd.n4880 gnd.n4879 4.74817
R13703 gnd.n4867 gnd.n1181 4.74817
R13704 gnd.n4865 gnd.n1180 4.74817
R13705 gnd.n4853 gnd.n1179 4.74817
R13706 gnd.n1178 gnd.n1175 4.74817
R13707 gnd.n4880 gnd.n1182 4.74817
R13708 gnd.n4878 gnd.n1181 4.74817
R13709 gnd.n4868 gnd.n1180 4.74817
R13710 gnd.n4864 gnd.n1179 4.74817
R13711 gnd.n4854 gnd.n1178 4.74817
R13712 gnd.n3067 gnd.n3066 4.7074
R13713 gnd.n54 gnd.n53 4.7074
R13714 gnd.n3087 gnd.n3067 4.65959
R13715 gnd.n74 gnd.n54 4.65959
R13716 gnd.n6878 gnd.n536 4.6132
R13717 gnd.n1021 gnd.n1018 4.6132
R13718 gnd.n4773 gnd.n992 4.46168
R13719 gnd.n5567 gnd.n5366 4.46168
R13720 gnd.n6409 gnd.n877 4.46168
R13721 gnd.n5585 gnd.t96 4.46168
R13722 gnd.n6465 gnd.n827 4.46168
R13723 gnd.n5657 gnd.n5656 4.46168
R13724 gnd.n5720 gnd.n5281 4.46168
R13725 gnd.n6545 gnd.n747 4.46168
R13726 gnd.n5935 gnd.n5934 4.46168
R13727 gnd.n6906 gnd.n518 4.46168
R13728 gnd.n5179 gnd.n5166 4.46111
R13729 gnd.n4024 gnd.n4020 4.38594
R13730 gnd.n3992 gnd.n3988 4.38594
R13731 gnd.n3960 gnd.n3956 4.38594
R13732 gnd.n3929 gnd.n3925 4.38594
R13733 gnd.n3897 gnd.n3893 4.38594
R13734 gnd.n3865 gnd.n3861 4.38594
R13735 gnd.n3833 gnd.n3829 4.38594
R13736 gnd.n3802 gnd.n3798 4.38594
R13737 gnd.n4035 gnd.n4013 4.26717
R13738 gnd.n4003 gnd.n3981 4.26717
R13739 gnd.n3971 gnd.n3949 4.26717
R13740 gnd.n3940 gnd.n3918 4.26717
R13741 gnd.n3908 gnd.n3886 4.26717
R13742 gnd.n3876 gnd.n3854 4.26717
R13743 gnd.n3844 gnd.n3822 4.26717
R13744 gnd.n3813 gnd.n3791 4.26717
R13745 gnd.t11 gnd.n3123 4.14303
R13746 gnd.n2836 gnd.t14 4.14303
R13747 gnd.n4747 gnd.t208 4.14303
R13748 gnd.n6745 gnd.t225 4.14303
R13749 gnd.n4043 gnd.n4042 4.08274
R13750 gnd.n5862 gnd.n5861 4.05904
R13751 gnd.n5505 gnd.n5504 4.05904
R13752 gnd.n5488 gnd.n5487 4.05904
R13753 gnd.n5879 gnd.n5878 4.05904
R13754 gnd.n15 gnd.n7 3.99943
R13755 gnd.n4043 gnd.n3915 3.70378
R13756 gnd.n3601 gnd.n3088 3.65935
R13757 gnd.n15 gnd.n14 3.60163
R13758 gnd.n4490 gnd.t43 3.50571
R13759 gnd.n4801 gnd.t72 3.50571
R13760 gnd.n901 gnd.n893 3.50571
R13761 gnd.n5937 gnd.n683 3.50571
R13762 gnd.n6706 gnd.t57 3.50571
R13763 gnd.n7353 gnd.t53 3.50571
R13764 gnd.n4034 gnd.n4015 3.49141
R13765 gnd.n4002 gnd.n3983 3.49141
R13766 gnd.n3970 gnd.n3951 3.49141
R13767 gnd.n3939 gnd.n3920 3.49141
R13768 gnd.n3907 gnd.n3888 3.49141
R13769 gnd.n3875 gnd.n3856 3.49141
R13770 gnd.n3843 gnd.n3824 3.49141
R13771 gnd.n3812 gnd.n3793 3.49141
R13772 gnd.n6393 gnd.t50 3.18706
R13773 gnd.n6417 gnd.n869 3.18706
R13774 gnd.n6457 gnd.n834 3.18706
R13775 gnd.n5657 gnd.t6 3.18706
R13776 gnd.n5667 gnd.n5313 3.18706
R13777 gnd.n5711 gnd.n5286 3.18706
R13778 gnd.n5720 gnd.t8 3.18706
R13779 gnd.n6553 gnd.n740 3.18706
R13780 gnd.n6593 gnd.n705 3.18706
R13781 gnd.n3130 gnd.t11 2.8684
R13782 gnd.t167 gnd.n887 2.8684
R13783 gnd.n5803 gnd.t4 2.8684
R13784 gnd.n3068 gnd.t318 2.82907
R13785 gnd.n3068 gnd.t264 2.82907
R13786 gnd.n3070 gnd.t303 2.82907
R13787 gnd.n3070 gnd.t179 2.82907
R13788 gnd.n3072 gnd.t214 2.82907
R13789 gnd.n3072 gnd.t191 2.82907
R13790 gnd.n3074 gnd.t189 2.82907
R13791 gnd.n3074 gnd.t329 2.82907
R13792 gnd.n3076 gnd.t199 2.82907
R13793 gnd.n3076 gnd.t254 2.82907
R13794 gnd.n3078 gnd.t293 2.82907
R13795 gnd.n3078 gnd.t237 2.82907
R13796 gnd.n3080 gnd.t270 2.82907
R13797 gnd.n3080 gnd.t195 2.82907
R13798 gnd.n3082 gnd.t240 2.82907
R13799 gnd.n3082 gnd.t322 2.82907
R13800 gnd.n3084 gnd.t297 2.82907
R13801 gnd.n3084 gnd.t296 2.82907
R13802 gnd.n3029 gnd.t207 2.82907
R13803 gnd.n3029 gnd.t235 2.82907
R13804 gnd.n3031 gnd.t253 2.82907
R13805 gnd.n3031 gnd.t319 2.82907
R13806 gnd.n3033 gnd.t233 2.82907
R13807 gnd.n3033 gnd.t224 2.82907
R13808 gnd.n3035 gnd.t278 2.82907
R13809 gnd.n3035 gnd.t183 2.82907
R13810 gnd.n3037 gnd.t324 2.82907
R13811 gnd.n3037 gnd.t243 2.82907
R13812 gnd.n3039 gnd.t260 2.82907
R13813 gnd.n3039 gnd.t292 2.82907
R13814 gnd.n3041 gnd.t308 2.82907
R13815 gnd.n3041 gnd.t234 2.82907
R13816 gnd.n3043 gnd.t244 2.82907
R13817 gnd.n3043 gnd.t273 2.82907
R13818 gnd.n3045 gnd.t197 2.82907
R13819 gnd.n3045 gnd.t220 2.82907
R13820 gnd.n3048 gnd.t328 2.82907
R13821 gnd.n3048 gnd.t209 2.82907
R13822 gnd.n3050 gnd.t228 2.82907
R13823 gnd.n3050 gnd.t285 2.82907
R13824 gnd.n3052 gnd.t203 2.82907
R13825 gnd.n3052 gnd.t337 2.82907
R13826 gnd.n3054 gnd.t252 2.82907
R13827 gnd.n3054 gnd.t239 2.82907
R13828 gnd.n3056 gnd.t309 2.82907
R13829 gnd.n3056 gnd.t222 2.82907
R13830 gnd.n3058 gnd.t181 2.82907
R13831 gnd.n3058 gnd.t263 2.82907
R13832 gnd.n3060 gnd.t279 2.82907
R13833 gnd.n3060 gnd.t204 2.82907
R13834 gnd.n3062 gnd.t218 2.82907
R13835 gnd.n3062 gnd.t251 2.82907
R13836 gnd.n3064 gnd.t325 2.82907
R13837 gnd.n3064 gnd.t334 2.82907
R13838 gnd.n71 gnd.t205 2.82907
R13839 gnd.n71 gnd.t223 2.82907
R13840 gnd.n69 gnd.t283 2.82907
R13841 gnd.n69 gnd.t187 2.82907
R13842 gnd.n67 gnd.t316 2.82907
R13843 gnd.n67 gnd.t230 2.82907
R13844 gnd.n65 gnd.t336 2.82907
R13845 gnd.n65 gnd.t249 2.82907
R13846 gnd.n63 gnd.t211 2.82907
R13847 gnd.n63 gnd.t327 2.82907
R13848 gnd.n61 gnd.t298 2.82907
R13849 gnd.n61 gnd.t312 2.82907
R13850 gnd.n59 gnd.t314 2.82907
R13851 gnd.n59 gnd.t333 2.82907
R13852 gnd.n57 gnd.t310 2.82907
R13853 gnd.n57 gnd.t259 2.82907
R13854 gnd.n55 gnd.t226 2.82907
R13855 gnd.n55 gnd.t295 2.82907
R13856 gnd.n32 gnd.t201 2.82907
R13857 gnd.n32 gnd.t213 2.82907
R13858 gnd.n30 gnd.t305 2.82907
R13859 gnd.n30 gnd.t281 2.82907
R13860 gnd.n28 gnd.t266 2.82907
R13861 gnd.n28 gnd.t330 2.82907
R13862 gnd.n26 gnd.t306 2.82907
R13863 gnd.n26 gnd.t299 2.82907
R13864 gnd.n24 gnd.t280 2.82907
R13865 gnd.n24 gnd.t317 2.82907
R13866 gnd.n22 gnd.t307 2.82907
R13867 gnd.n22 gnd.t313 2.82907
R13868 gnd.n20 gnd.t257 2.82907
R13869 gnd.n20 gnd.t216 2.82907
R13870 gnd.n18 gnd.t193 2.82907
R13871 gnd.n18 gnd.t288 2.82907
R13872 gnd.n16 gnd.t268 2.82907
R13873 gnd.n16 gnd.t335 2.82907
R13874 gnd.n51 gnd.t326 2.82907
R13875 gnd.n51 gnd.t331 2.82907
R13876 gnd.n49 gnd.t284 2.82907
R13877 gnd.n49 gnd.t256 2.82907
R13878 gnd.n47 gnd.t242 2.82907
R13879 gnd.n47 gnd.t315 2.82907
R13880 gnd.n45 gnd.t301 2.82907
R13881 gnd.n45 gnd.t267 2.82907
R13882 gnd.n43 gnd.t255 2.82907
R13883 gnd.n43 gnd.t291 2.82907
R13884 gnd.n41 gnd.t277 2.82907
R13885 gnd.n41 gnd.t287 2.82907
R13886 gnd.n39 gnd.t232 2.82907
R13887 gnd.n39 gnd.t332 2.82907
R13888 gnd.n37 gnd.t323 2.82907
R13889 gnd.n37 gnd.t261 2.82907
R13890 gnd.n35 gnd.t245 2.82907
R13891 gnd.n35 gnd.t320 2.82907
R13892 gnd.n4031 gnd.n4030 2.71565
R13893 gnd.n3999 gnd.n3998 2.71565
R13894 gnd.n3967 gnd.n3966 2.71565
R13895 gnd.n3936 gnd.n3935 2.71565
R13896 gnd.n3904 gnd.n3903 2.71565
R13897 gnd.n3872 gnd.n3871 2.71565
R13898 gnd.n3840 gnd.n3839 2.71565
R13899 gnd.n3809 gnd.n3808 2.71565
R13900 gnd.t96 gnd.n5356 2.54975
R13901 gnd.n5341 gnd.t29 2.54975
R13902 gnd.n5763 gnd.t162 2.54975
R13903 gnd.n5797 gnd.t137 2.54975
R13904 gnd.n3601 gnd.n3089 2.27742
R13905 gnd.n3601 gnd.n2945 2.27742
R13906 gnd.n3602 gnd.n3601 2.27742
R13907 gnd.n3601 gnd.n3028 2.27742
R13908 gnd.n7185 gnd.n7184 2.27742
R13909 gnd.n7185 gnd.n304 2.27742
R13910 gnd.n7185 gnd.n303 2.27742
R13911 gnd.n7185 gnd.n302 2.27742
R13912 gnd.n7185 gnd.n301 2.27742
R13913 gnd.n4881 gnd.n4880 2.27742
R13914 gnd.n4881 gnd.n1181 2.27742
R13915 gnd.n4881 gnd.n1180 2.27742
R13916 gnd.n4881 gnd.n1179 2.27742
R13917 gnd.n4881 gnd.n1178 2.27742
R13918 gnd.n3481 gnd.t39 2.23109
R13919 gnd.n3606 gnd.t10 2.23109
R13920 gnd.n5656 gnd.t346 2.23109
R13921 gnd.n5281 gnd.t160 2.23109
R13922 gnd.n236 gnd.t212 2.23109
R13923 gnd.n4027 gnd.n4017 1.93989
R13924 gnd.n3995 gnd.n3985 1.93989
R13925 gnd.n3963 gnd.n3953 1.93989
R13926 gnd.n3932 gnd.n3922 1.93989
R13927 gnd.n3900 gnd.n3890 1.93989
R13928 gnd.n3868 gnd.n3858 1.93989
R13929 gnd.n3836 gnd.n3826 1.93989
R13930 gnd.n3805 gnd.n3795 1.93989
R13931 gnd.t119 gnd.n885 1.91244
R13932 gnd.n6425 gnd.n862 1.91244
R13933 gnd.n6449 gnd.n841 1.91244
R13934 gnd.n5308 gnd.n5307 1.91244
R13935 gnd.n5676 gnd.t177 1.91244
R13936 gnd.n5292 gnd.t176 1.91244
R13937 gnd.n5702 gnd.n5291 1.91244
R13938 gnd.n6561 gnd.n733 1.91244
R13939 gnd.n6585 gnd.n712 1.91244
R13940 gnd.n6601 gnd.t137 1.91244
R13941 gnd.t0 gnd.n3492 1.59378
R13942 gnd.n2902 gnd.t25 1.59378
R13943 gnd.n3000 gnd.t156 1.59378
R13944 gnd.n4530 gnd.t219 1.59378
R13945 gnd.n4732 gnd.t206 1.59378
R13946 gnd.n5594 gnd.t2 1.59378
R13947 gnd.n5781 gnd.t344 1.59378
R13948 gnd.n6750 gnd.t294 1.59378
R13949 gnd.n7245 gnd.t200 1.59378
R13950 gnd.t35 gnd.n877 1.27512
R13951 gnd.n5797 gnd.t68 1.27512
R13952 gnd.n5937 gnd.t128 1.27512
R13953 gnd.n3334 gnd.n3326 1.16414
R13954 gnd.n4087 gnd.n1467 1.16414
R13955 gnd.n4026 gnd.n4019 1.16414
R13956 gnd.n3994 gnd.n3987 1.16414
R13957 gnd.n3962 gnd.n3955 1.16414
R13958 gnd.n3931 gnd.n3924 1.16414
R13959 gnd.n3899 gnd.n3892 1.16414
R13960 gnd.n3867 gnd.n3860 1.16414
R13961 gnd.n3835 gnd.n3828 1.16414
R13962 gnd.n3804 gnd.n3797 1.16414
R13963 gnd.n6878 gnd.n6877 0.970197
R13964 gnd.n6266 gnd.n1018 0.970197
R13965 gnd.n4010 gnd.n3978 0.962709
R13966 gnd.n4042 gnd.n4010 0.962709
R13967 gnd.n3883 gnd.n3851 0.962709
R13968 gnd.n3915 gnd.n3883 0.962709
R13969 gnd.n3572 gnd.t172 0.956468
R13970 gnd.n3710 gnd.t19 0.956468
R13971 gnd.n4572 gnd.t269 0.956468
R13972 gnd.n4692 gnd.t190 0.956468
R13973 gnd.n6385 gnd.t32 0.956468
R13974 gnd.n6625 gnd.t165 0.956468
R13975 gnd.n6798 gnd.t231 0.956468
R13976 gnd.n7213 gnd.t229 0.956468
R13977 gnd.n3079 gnd.n3077 0.773756
R13978 gnd.n66 gnd.n64 0.773756
R13979 gnd.n3086 gnd.n3085 0.773756
R13980 gnd.n3085 gnd.n3083 0.773756
R13981 gnd.n3083 gnd.n3081 0.773756
R13982 gnd.n3081 gnd.n3079 0.773756
R13983 gnd.n3077 gnd.n3075 0.773756
R13984 gnd.n3075 gnd.n3073 0.773756
R13985 gnd.n3073 gnd.n3071 0.773756
R13986 gnd.n3071 gnd.n3069 0.773756
R13987 gnd.n58 gnd.n56 0.773756
R13988 gnd.n60 gnd.n58 0.773756
R13989 gnd.n62 gnd.n60 0.773756
R13990 gnd.n64 gnd.n62 0.773756
R13991 gnd.n68 gnd.n66 0.773756
R13992 gnd.n70 gnd.n68 0.773756
R13993 gnd.n72 gnd.n70 0.773756
R13994 gnd.n73 gnd.n72 0.773756
R13995 gnd.n2 gnd.n1 0.672012
R13996 gnd.n3 gnd.n2 0.672012
R13997 gnd.n4 gnd.n3 0.672012
R13998 gnd.n5 gnd.n4 0.672012
R13999 gnd.n6 gnd.n5 0.672012
R14000 gnd.n7 gnd.n6 0.672012
R14001 gnd.n9 gnd.n8 0.672012
R14002 gnd.n10 gnd.n9 0.672012
R14003 gnd.n11 gnd.n10 0.672012
R14004 gnd.n12 gnd.n11 0.672012
R14005 gnd.n13 gnd.n12 0.672012
R14006 gnd.n14 gnd.n13 0.672012
R14007 gnd.n6433 gnd.n854 0.637812
R14008 gnd.n6441 gnd.n848 0.637812
R14009 gnd.n5684 gnd.n5302 0.637812
R14010 gnd.n5693 gnd.n5297 0.637812
R14011 gnd.n6569 gnd.n726 0.637812
R14012 gnd.n6577 gnd.n720 0.637812
R14013 gnd.n7488 gnd.n7487 0.63688
R14014 gnd gnd.n0 0.634843
R14015 gnd.n3047 gnd.n3046 0.573776
R14016 gnd.n3046 gnd.n3044 0.573776
R14017 gnd.n3044 gnd.n3042 0.573776
R14018 gnd.n3042 gnd.n3040 0.573776
R14019 gnd.n3040 gnd.n3038 0.573776
R14020 gnd.n3038 gnd.n3036 0.573776
R14021 gnd.n3036 gnd.n3034 0.573776
R14022 gnd.n3034 gnd.n3032 0.573776
R14023 gnd.n3032 gnd.n3030 0.573776
R14024 gnd.n3066 gnd.n3065 0.573776
R14025 gnd.n3065 gnd.n3063 0.573776
R14026 gnd.n3063 gnd.n3061 0.573776
R14027 gnd.n3061 gnd.n3059 0.573776
R14028 gnd.n3059 gnd.n3057 0.573776
R14029 gnd.n3057 gnd.n3055 0.573776
R14030 gnd.n3055 gnd.n3053 0.573776
R14031 gnd.n3053 gnd.n3051 0.573776
R14032 gnd.n3051 gnd.n3049 0.573776
R14033 gnd.n19 gnd.n17 0.573776
R14034 gnd.n21 gnd.n19 0.573776
R14035 gnd.n23 gnd.n21 0.573776
R14036 gnd.n25 gnd.n23 0.573776
R14037 gnd.n27 gnd.n25 0.573776
R14038 gnd.n29 gnd.n27 0.573776
R14039 gnd.n31 gnd.n29 0.573776
R14040 gnd.n33 gnd.n31 0.573776
R14041 gnd.n34 gnd.n33 0.573776
R14042 gnd.n38 gnd.n36 0.573776
R14043 gnd.n40 gnd.n38 0.573776
R14044 gnd.n42 gnd.n40 0.573776
R14045 gnd.n44 gnd.n42 0.573776
R14046 gnd.n46 gnd.n44 0.573776
R14047 gnd.n48 gnd.n46 0.573776
R14048 gnd.n50 gnd.n48 0.573776
R14049 gnd.n52 gnd.n50 0.573776
R14050 gnd.n53 gnd.n52 0.573776
R14051 gnd.n7185 gnd.n300 0.5435
R14052 gnd.n4881 gnd.n1177 0.5435
R14053 gnd.n6219 gnd.n6218 0.523366
R14054 gnd.n5954 gnd.n5950 0.523366
R14055 gnd.n6673 gnd.n6672 0.489829
R14056 gnd.n6333 gnd.n933 0.489829
R14057 gnd.n2974 gnd.n1471 0.486781
R14058 gnd.n3383 gnd.n3382 0.48678
R14059 gnd.n4065 gnd.n1425 0.480683
R14060 gnd.n3467 gnd.n3466 0.480683
R14061 gnd.n4238 gnd.n4237 0.477634
R14062 gnd.n4485 gnd.n1398 0.477634
R14063 gnd.n7336 gnd.n7335 0.477634
R14064 gnd.n7438 gnd.n7437 0.477634
R14065 gnd.n7430 gnd.n7429 0.465439
R14066 gnd.n7359 gnd.n7358 0.465439
R14067 gnd.n6838 gnd.n562 0.465439
R14068 gnd.n6911 gnd.n6910 0.465439
R14069 gnd.n6299 gnd.n6298 0.465439
R14070 gnd.n6230 gnd.n6229 0.465439
R14071 gnd.n4404 gnd.n4399 0.465439
R14072 gnd.n4479 gnd.n4478 0.465439
R14073 gnd.n2550 gnd.n1598 0.459342
R14074 gnd.n1913 gnd.n1907 0.459342
R14075 gnd.n7078 gnd.n7077 0.459342
R14076 gnd.n2762 gnd.n2761 0.459342
R14077 gnd.n6326 gnd.n6325 0.388379
R14078 gnd.n4023 gnd.n4022 0.388379
R14079 gnd.n3991 gnd.n3990 0.388379
R14080 gnd.n3959 gnd.n3958 0.388379
R14081 gnd.n3928 gnd.n3927 0.388379
R14082 gnd.n3896 gnd.n3895 0.388379
R14083 gnd.n3864 gnd.n3863 0.388379
R14084 gnd.n3832 gnd.n3831 0.388379
R14085 gnd.n3801 gnd.n3800 0.388379
R14086 gnd.n7399 gnd.n7398 0.388379
R14087 gnd.n4314 gnd.n4310 0.388379
R14088 gnd.n6026 gnd.n6022 0.388379
R14089 gnd.n6221 gnd.n6220 0.377553
R14090 gnd.n5955 gnd.n477 0.377553
R14091 gnd.n7488 gnd.n15 0.374463
R14092 gnd.t12 gnd.n3761 0.319156
R14093 gnd.n4629 gnd.t236 0.319156
R14094 gnd.n4653 gnd.t188 0.319156
R14095 gnd.t177 gnd.t163 0.319156
R14096 gnd.t176 gnd.t152 0.319156
R14097 gnd.n7071 gnd.t286 0.319156
R14098 gnd.n7165 gnd.t300 0.319156
R14099 gnd.n3301 gnd.n3279 0.311721
R14100 gnd gnd.n7488 0.295112
R14101 gnd.n4132 gnd.n4131 0.268793
R14102 gnd.n6314 gnd.n970 0.247451
R14103 gnd.n6831 gnd.n566 0.247451
R14104 gnd.n4131 gnd.n4130 0.241354
R14105 gnd.n536 gnd.n533 0.229039
R14106 gnd.n539 gnd.n536 0.229039
R14107 gnd.n1021 gnd.n1020 0.229039
R14108 gnd.n1022 gnd.n1021 0.229039
R14109 gnd.n3088 gnd.n0 0.210825
R14110 gnd.n3455 gnd.n3254 0.206293
R14111 gnd.n4040 gnd.n4012 0.155672
R14112 gnd.n4033 gnd.n4012 0.155672
R14113 gnd.n4033 gnd.n4032 0.155672
R14114 gnd.n4032 gnd.n4016 0.155672
R14115 gnd.n4025 gnd.n4016 0.155672
R14116 gnd.n4025 gnd.n4024 0.155672
R14117 gnd.n4008 gnd.n3980 0.155672
R14118 gnd.n4001 gnd.n3980 0.155672
R14119 gnd.n4001 gnd.n4000 0.155672
R14120 gnd.n4000 gnd.n3984 0.155672
R14121 gnd.n3993 gnd.n3984 0.155672
R14122 gnd.n3993 gnd.n3992 0.155672
R14123 gnd.n3976 gnd.n3948 0.155672
R14124 gnd.n3969 gnd.n3948 0.155672
R14125 gnd.n3969 gnd.n3968 0.155672
R14126 gnd.n3968 gnd.n3952 0.155672
R14127 gnd.n3961 gnd.n3952 0.155672
R14128 gnd.n3961 gnd.n3960 0.155672
R14129 gnd.n3945 gnd.n3917 0.155672
R14130 gnd.n3938 gnd.n3917 0.155672
R14131 gnd.n3938 gnd.n3937 0.155672
R14132 gnd.n3937 gnd.n3921 0.155672
R14133 gnd.n3930 gnd.n3921 0.155672
R14134 gnd.n3930 gnd.n3929 0.155672
R14135 gnd.n3913 gnd.n3885 0.155672
R14136 gnd.n3906 gnd.n3885 0.155672
R14137 gnd.n3906 gnd.n3905 0.155672
R14138 gnd.n3905 gnd.n3889 0.155672
R14139 gnd.n3898 gnd.n3889 0.155672
R14140 gnd.n3898 gnd.n3897 0.155672
R14141 gnd.n3881 gnd.n3853 0.155672
R14142 gnd.n3874 gnd.n3853 0.155672
R14143 gnd.n3874 gnd.n3873 0.155672
R14144 gnd.n3873 gnd.n3857 0.155672
R14145 gnd.n3866 gnd.n3857 0.155672
R14146 gnd.n3866 gnd.n3865 0.155672
R14147 gnd.n3849 gnd.n3821 0.155672
R14148 gnd.n3842 gnd.n3821 0.155672
R14149 gnd.n3842 gnd.n3841 0.155672
R14150 gnd.n3841 gnd.n3825 0.155672
R14151 gnd.n3834 gnd.n3825 0.155672
R14152 gnd.n3834 gnd.n3833 0.155672
R14153 gnd.n3818 gnd.n3790 0.155672
R14154 gnd.n3811 gnd.n3790 0.155672
R14155 gnd.n3811 gnd.n3810 0.155672
R14156 gnd.n3810 gnd.n3794 0.155672
R14157 gnd.n3803 gnd.n3794 0.155672
R14158 gnd.n3803 gnd.n3802 0.155672
R14159 gnd.n4163 gnd.n1425 0.152939
R14160 gnd.n4163 gnd.n4162 0.152939
R14161 gnd.n4162 gnd.n4161 0.152939
R14162 gnd.n4161 gnd.n1427 0.152939
R14163 gnd.n1428 gnd.n1427 0.152939
R14164 gnd.n1429 gnd.n1428 0.152939
R14165 gnd.n1430 gnd.n1429 0.152939
R14166 gnd.n1431 gnd.n1430 0.152939
R14167 gnd.n1432 gnd.n1431 0.152939
R14168 gnd.n1433 gnd.n1432 0.152939
R14169 gnd.n1434 gnd.n1433 0.152939
R14170 gnd.n1435 gnd.n1434 0.152939
R14171 gnd.n1436 gnd.n1435 0.152939
R14172 gnd.n1437 gnd.n1436 0.152939
R14173 gnd.n4133 gnd.n1437 0.152939
R14174 gnd.n4133 gnd.n4132 0.152939
R14175 gnd.n3468 gnd.n3467 0.152939
R14176 gnd.n3468 gnd.n3172 0.152939
R14177 gnd.n3496 gnd.n3172 0.152939
R14178 gnd.n3497 gnd.n3496 0.152939
R14179 gnd.n3498 gnd.n3497 0.152939
R14180 gnd.n3499 gnd.n3498 0.152939
R14181 gnd.n3499 gnd.n3144 0.152939
R14182 gnd.n3526 gnd.n3144 0.152939
R14183 gnd.n3527 gnd.n3526 0.152939
R14184 gnd.n3528 gnd.n3527 0.152939
R14185 gnd.n3529 gnd.n3528 0.152939
R14186 gnd.n3530 gnd.n3529 0.152939
R14187 gnd.n3532 gnd.n3530 0.152939
R14188 gnd.n3532 gnd.n3531 0.152939
R14189 gnd.n3531 gnd.n3112 0.152939
R14190 gnd.n3585 gnd.n3112 0.152939
R14191 gnd.n3586 gnd.n3585 0.152939
R14192 gnd.n3587 gnd.n3586 0.152939
R14193 gnd.n3587 gnd.n2930 0.152939
R14194 gnd.n3621 gnd.n2930 0.152939
R14195 gnd.n3622 gnd.n3621 0.152939
R14196 gnd.n3623 gnd.n3622 0.152939
R14197 gnd.n3624 gnd.n3623 0.152939
R14198 gnd.n3624 gnd.n2906 0.152939
R14199 gnd.n3652 gnd.n2906 0.152939
R14200 gnd.n3653 gnd.n3652 0.152939
R14201 gnd.n3654 gnd.n3653 0.152939
R14202 gnd.n3655 gnd.n3654 0.152939
R14203 gnd.n3655 gnd.n2880 0.152939
R14204 gnd.n3683 gnd.n2880 0.152939
R14205 gnd.n3684 gnd.n3683 0.152939
R14206 gnd.n3685 gnd.n3684 0.152939
R14207 gnd.n3686 gnd.n3685 0.152939
R14208 gnd.n3686 gnd.n2855 0.152939
R14209 gnd.n3714 gnd.n2855 0.152939
R14210 gnd.n3715 gnd.n3714 0.152939
R14211 gnd.n3716 gnd.n3715 0.152939
R14212 gnd.n3717 gnd.n3716 0.152939
R14213 gnd.n3717 gnd.n2830 0.152939
R14214 gnd.n3745 gnd.n2830 0.152939
R14215 gnd.n3746 gnd.n3745 0.152939
R14216 gnd.n3747 gnd.n3746 0.152939
R14217 gnd.n3748 gnd.n3747 0.152939
R14218 gnd.n3748 gnd.n2804 0.152939
R14219 gnd.n3776 gnd.n2804 0.152939
R14220 gnd.n3777 gnd.n3776 0.152939
R14221 gnd.n3778 gnd.n3777 0.152939
R14222 gnd.n3779 gnd.n3778 0.152939
R14223 gnd.n3779 gnd.n2779 0.152939
R14224 gnd.n4062 gnd.n2779 0.152939
R14225 gnd.n4063 gnd.n4062 0.152939
R14226 gnd.n4064 gnd.n4063 0.152939
R14227 gnd.n4065 gnd.n4064 0.152939
R14228 gnd.n3466 gnd.n3196 0.152939
R14229 gnd.n3217 gnd.n3196 0.152939
R14230 gnd.n3218 gnd.n3217 0.152939
R14231 gnd.n3224 gnd.n3218 0.152939
R14232 gnd.n3225 gnd.n3224 0.152939
R14233 gnd.n3226 gnd.n3225 0.152939
R14234 gnd.n3226 gnd.n3215 0.152939
R14235 gnd.n3234 gnd.n3215 0.152939
R14236 gnd.n3235 gnd.n3234 0.152939
R14237 gnd.n3236 gnd.n3235 0.152939
R14238 gnd.n3236 gnd.n3213 0.152939
R14239 gnd.n3244 gnd.n3213 0.152939
R14240 gnd.n3245 gnd.n3244 0.152939
R14241 gnd.n3246 gnd.n3245 0.152939
R14242 gnd.n3246 gnd.n3211 0.152939
R14243 gnd.n3254 gnd.n3211 0.152939
R14244 gnd.n4130 gnd.n1442 0.152939
R14245 gnd.n1444 gnd.n1442 0.152939
R14246 gnd.n1445 gnd.n1444 0.152939
R14247 gnd.n1446 gnd.n1445 0.152939
R14248 gnd.n1447 gnd.n1446 0.152939
R14249 gnd.n1448 gnd.n1447 0.152939
R14250 gnd.n1449 gnd.n1448 0.152939
R14251 gnd.n1450 gnd.n1449 0.152939
R14252 gnd.n1451 gnd.n1450 0.152939
R14253 gnd.n1452 gnd.n1451 0.152939
R14254 gnd.n1453 gnd.n1452 0.152939
R14255 gnd.n1454 gnd.n1453 0.152939
R14256 gnd.n1455 gnd.n1454 0.152939
R14257 gnd.n1456 gnd.n1455 0.152939
R14258 gnd.n1457 gnd.n1456 0.152939
R14259 gnd.n1458 gnd.n1457 0.152939
R14260 gnd.n1459 gnd.n1458 0.152939
R14261 gnd.n1460 gnd.n1459 0.152939
R14262 gnd.n1461 gnd.n1460 0.152939
R14263 gnd.n1462 gnd.n1461 0.152939
R14264 gnd.n1463 gnd.n1462 0.152939
R14265 gnd.n1464 gnd.n1463 0.152939
R14266 gnd.n1468 gnd.n1464 0.152939
R14267 gnd.n1469 gnd.n1468 0.152939
R14268 gnd.n1470 gnd.n1469 0.152939
R14269 gnd.n1471 gnd.n1470 0.152939
R14270 gnd.n2948 gnd.n2947 0.152939
R14271 gnd.n2949 gnd.n2948 0.152939
R14272 gnd.n2950 gnd.n2949 0.152939
R14273 gnd.n2951 gnd.n2950 0.152939
R14274 gnd.n2952 gnd.n2951 0.152939
R14275 gnd.n2953 gnd.n2952 0.152939
R14276 gnd.n2954 gnd.n2953 0.152939
R14277 gnd.n2955 gnd.n2954 0.152939
R14278 gnd.n2956 gnd.n2955 0.152939
R14279 gnd.n2957 gnd.n2956 0.152939
R14280 gnd.n2958 gnd.n2957 0.152939
R14281 gnd.n2959 gnd.n2958 0.152939
R14282 gnd.n2960 gnd.n2959 0.152939
R14283 gnd.n2961 gnd.n2960 0.152939
R14284 gnd.n2962 gnd.n2961 0.152939
R14285 gnd.n2963 gnd.n2962 0.152939
R14286 gnd.n2964 gnd.n2963 0.152939
R14287 gnd.n2965 gnd.n2964 0.152939
R14288 gnd.n2966 gnd.n2965 0.152939
R14289 gnd.n2967 gnd.n2966 0.152939
R14290 gnd.n2968 gnd.n2967 0.152939
R14291 gnd.n2969 gnd.n2968 0.152939
R14292 gnd.n2970 gnd.n2969 0.152939
R14293 gnd.n2971 gnd.n2970 0.152939
R14294 gnd.n2972 gnd.n2971 0.152939
R14295 gnd.n2973 gnd.n2972 0.152939
R14296 gnd.n2975 gnd.n2973 0.152939
R14297 gnd.n2975 gnd.n2974 0.152939
R14298 gnd.n3384 gnd.n3383 0.152939
R14299 gnd.n3384 gnd.n3274 0.152939
R14300 gnd.n3399 gnd.n3274 0.152939
R14301 gnd.n3400 gnd.n3399 0.152939
R14302 gnd.n3401 gnd.n3400 0.152939
R14303 gnd.n3401 gnd.n3262 0.152939
R14304 gnd.n3415 gnd.n3262 0.152939
R14305 gnd.n3416 gnd.n3415 0.152939
R14306 gnd.n3417 gnd.n3416 0.152939
R14307 gnd.n3418 gnd.n3417 0.152939
R14308 gnd.n3419 gnd.n3418 0.152939
R14309 gnd.n3420 gnd.n3419 0.152939
R14310 gnd.n3421 gnd.n3420 0.152939
R14311 gnd.n3422 gnd.n3421 0.152939
R14312 gnd.n3423 gnd.n3422 0.152939
R14313 gnd.n3424 gnd.n3423 0.152939
R14314 gnd.n3425 gnd.n3424 0.152939
R14315 gnd.n3426 gnd.n3425 0.152939
R14316 gnd.n3427 gnd.n3426 0.152939
R14317 gnd.n3428 gnd.n3427 0.152939
R14318 gnd.n3429 gnd.n3428 0.152939
R14319 gnd.n3429 gnd.n3127 0.152939
R14320 gnd.n3552 gnd.n3127 0.152939
R14321 gnd.n3553 gnd.n3552 0.152939
R14322 gnd.n3554 gnd.n3553 0.152939
R14323 gnd.n3555 gnd.n3554 0.152939
R14324 gnd.n3555 gnd.n3090 0.152939
R14325 gnd.n3600 gnd.n3090 0.152939
R14326 gnd.n3302 gnd.n3301 0.152939
R14327 gnd.n3303 gnd.n3302 0.152939
R14328 gnd.n3304 gnd.n3303 0.152939
R14329 gnd.n3305 gnd.n3304 0.152939
R14330 gnd.n3306 gnd.n3305 0.152939
R14331 gnd.n3307 gnd.n3306 0.152939
R14332 gnd.n3308 gnd.n3307 0.152939
R14333 gnd.n3309 gnd.n3308 0.152939
R14334 gnd.n3310 gnd.n3309 0.152939
R14335 gnd.n3311 gnd.n3310 0.152939
R14336 gnd.n3312 gnd.n3311 0.152939
R14337 gnd.n3313 gnd.n3312 0.152939
R14338 gnd.n3314 gnd.n3313 0.152939
R14339 gnd.n3315 gnd.n3314 0.152939
R14340 gnd.n3316 gnd.n3315 0.152939
R14341 gnd.n3317 gnd.n3316 0.152939
R14342 gnd.n3318 gnd.n3317 0.152939
R14343 gnd.n3319 gnd.n3318 0.152939
R14344 gnd.n3320 gnd.n3319 0.152939
R14345 gnd.n3321 gnd.n3320 0.152939
R14346 gnd.n3322 gnd.n3321 0.152939
R14347 gnd.n3323 gnd.n3322 0.152939
R14348 gnd.n3327 gnd.n3323 0.152939
R14349 gnd.n3328 gnd.n3327 0.152939
R14350 gnd.n3328 gnd.n3285 0.152939
R14351 gnd.n3382 gnd.n3285 0.152939
R14352 gnd.n2550 gnd.n2549 0.152939
R14353 gnd.n2549 gnd.n2548 0.152939
R14354 gnd.n2548 gnd.n1604 0.152939
R14355 gnd.n1609 gnd.n1604 0.152939
R14356 gnd.n1610 gnd.n1609 0.152939
R14357 gnd.n1611 gnd.n1610 0.152939
R14358 gnd.n1616 gnd.n1611 0.152939
R14359 gnd.n1617 gnd.n1616 0.152939
R14360 gnd.n1618 gnd.n1617 0.152939
R14361 gnd.n1619 gnd.n1618 0.152939
R14362 gnd.n1624 gnd.n1619 0.152939
R14363 gnd.n1625 gnd.n1624 0.152939
R14364 gnd.n1626 gnd.n1625 0.152939
R14365 gnd.n1627 gnd.n1626 0.152939
R14366 gnd.n1632 gnd.n1627 0.152939
R14367 gnd.n1633 gnd.n1632 0.152939
R14368 gnd.n1634 gnd.n1633 0.152939
R14369 gnd.n1635 gnd.n1634 0.152939
R14370 gnd.n1640 gnd.n1635 0.152939
R14371 gnd.n1641 gnd.n1640 0.152939
R14372 gnd.n1642 gnd.n1641 0.152939
R14373 gnd.n1643 gnd.n1642 0.152939
R14374 gnd.n1648 gnd.n1643 0.152939
R14375 gnd.n1649 gnd.n1648 0.152939
R14376 gnd.n1650 gnd.n1649 0.152939
R14377 gnd.n1651 gnd.n1650 0.152939
R14378 gnd.n1656 gnd.n1651 0.152939
R14379 gnd.n1657 gnd.n1656 0.152939
R14380 gnd.n1658 gnd.n1657 0.152939
R14381 gnd.n1659 gnd.n1658 0.152939
R14382 gnd.n1664 gnd.n1659 0.152939
R14383 gnd.n1665 gnd.n1664 0.152939
R14384 gnd.n1666 gnd.n1665 0.152939
R14385 gnd.n1667 gnd.n1666 0.152939
R14386 gnd.n1672 gnd.n1667 0.152939
R14387 gnd.n1673 gnd.n1672 0.152939
R14388 gnd.n1674 gnd.n1673 0.152939
R14389 gnd.n1675 gnd.n1674 0.152939
R14390 gnd.n1680 gnd.n1675 0.152939
R14391 gnd.n1681 gnd.n1680 0.152939
R14392 gnd.n1682 gnd.n1681 0.152939
R14393 gnd.n1683 gnd.n1682 0.152939
R14394 gnd.n1688 gnd.n1683 0.152939
R14395 gnd.n1689 gnd.n1688 0.152939
R14396 gnd.n1690 gnd.n1689 0.152939
R14397 gnd.n1691 gnd.n1690 0.152939
R14398 gnd.n1696 gnd.n1691 0.152939
R14399 gnd.n1697 gnd.n1696 0.152939
R14400 gnd.n1698 gnd.n1697 0.152939
R14401 gnd.n1699 gnd.n1698 0.152939
R14402 gnd.n1704 gnd.n1699 0.152939
R14403 gnd.n1705 gnd.n1704 0.152939
R14404 gnd.n1706 gnd.n1705 0.152939
R14405 gnd.n1707 gnd.n1706 0.152939
R14406 gnd.n1712 gnd.n1707 0.152939
R14407 gnd.n1713 gnd.n1712 0.152939
R14408 gnd.n1714 gnd.n1713 0.152939
R14409 gnd.n1715 gnd.n1714 0.152939
R14410 gnd.n1720 gnd.n1715 0.152939
R14411 gnd.n1721 gnd.n1720 0.152939
R14412 gnd.n1722 gnd.n1721 0.152939
R14413 gnd.n1723 gnd.n1722 0.152939
R14414 gnd.n1728 gnd.n1723 0.152939
R14415 gnd.n1729 gnd.n1728 0.152939
R14416 gnd.n1730 gnd.n1729 0.152939
R14417 gnd.n1731 gnd.n1730 0.152939
R14418 gnd.n1736 gnd.n1731 0.152939
R14419 gnd.n1737 gnd.n1736 0.152939
R14420 gnd.n1738 gnd.n1737 0.152939
R14421 gnd.n1739 gnd.n1738 0.152939
R14422 gnd.n1744 gnd.n1739 0.152939
R14423 gnd.n1745 gnd.n1744 0.152939
R14424 gnd.n1746 gnd.n1745 0.152939
R14425 gnd.n1747 gnd.n1746 0.152939
R14426 gnd.n1752 gnd.n1747 0.152939
R14427 gnd.n1753 gnd.n1752 0.152939
R14428 gnd.n1754 gnd.n1753 0.152939
R14429 gnd.n1755 gnd.n1754 0.152939
R14430 gnd.n1760 gnd.n1755 0.152939
R14431 gnd.n1761 gnd.n1760 0.152939
R14432 gnd.n1762 gnd.n1761 0.152939
R14433 gnd.n1763 gnd.n1762 0.152939
R14434 gnd.n1768 gnd.n1763 0.152939
R14435 gnd.n1769 gnd.n1768 0.152939
R14436 gnd.n1770 gnd.n1769 0.152939
R14437 gnd.n1771 gnd.n1770 0.152939
R14438 gnd.n1776 gnd.n1771 0.152939
R14439 gnd.n1777 gnd.n1776 0.152939
R14440 gnd.n1778 gnd.n1777 0.152939
R14441 gnd.n1779 gnd.n1778 0.152939
R14442 gnd.n1784 gnd.n1779 0.152939
R14443 gnd.n1785 gnd.n1784 0.152939
R14444 gnd.n1786 gnd.n1785 0.152939
R14445 gnd.n1787 gnd.n1786 0.152939
R14446 gnd.n1792 gnd.n1787 0.152939
R14447 gnd.n1793 gnd.n1792 0.152939
R14448 gnd.n1794 gnd.n1793 0.152939
R14449 gnd.n1795 gnd.n1794 0.152939
R14450 gnd.n1800 gnd.n1795 0.152939
R14451 gnd.n1801 gnd.n1800 0.152939
R14452 gnd.n1802 gnd.n1801 0.152939
R14453 gnd.n1803 gnd.n1802 0.152939
R14454 gnd.n1808 gnd.n1803 0.152939
R14455 gnd.n1809 gnd.n1808 0.152939
R14456 gnd.n1810 gnd.n1809 0.152939
R14457 gnd.n1811 gnd.n1810 0.152939
R14458 gnd.n1816 gnd.n1811 0.152939
R14459 gnd.n1817 gnd.n1816 0.152939
R14460 gnd.n1818 gnd.n1817 0.152939
R14461 gnd.n1819 gnd.n1818 0.152939
R14462 gnd.n1824 gnd.n1819 0.152939
R14463 gnd.n1825 gnd.n1824 0.152939
R14464 gnd.n1826 gnd.n1825 0.152939
R14465 gnd.n1827 gnd.n1826 0.152939
R14466 gnd.n1832 gnd.n1827 0.152939
R14467 gnd.n1833 gnd.n1832 0.152939
R14468 gnd.n1834 gnd.n1833 0.152939
R14469 gnd.n1835 gnd.n1834 0.152939
R14470 gnd.n1840 gnd.n1835 0.152939
R14471 gnd.n1841 gnd.n1840 0.152939
R14472 gnd.n1842 gnd.n1841 0.152939
R14473 gnd.n1843 gnd.n1842 0.152939
R14474 gnd.n1848 gnd.n1843 0.152939
R14475 gnd.n1849 gnd.n1848 0.152939
R14476 gnd.n1850 gnd.n1849 0.152939
R14477 gnd.n1851 gnd.n1850 0.152939
R14478 gnd.n1856 gnd.n1851 0.152939
R14479 gnd.n1857 gnd.n1856 0.152939
R14480 gnd.n1858 gnd.n1857 0.152939
R14481 gnd.n1859 gnd.n1858 0.152939
R14482 gnd.n1864 gnd.n1859 0.152939
R14483 gnd.n1865 gnd.n1864 0.152939
R14484 gnd.n1866 gnd.n1865 0.152939
R14485 gnd.n1867 gnd.n1866 0.152939
R14486 gnd.n1872 gnd.n1867 0.152939
R14487 gnd.n1873 gnd.n1872 0.152939
R14488 gnd.n1874 gnd.n1873 0.152939
R14489 gnd.n1875 gnd.n1874 0.152939
R14490 gnd.n1880 gnd.n1875 0.152939
R14491 gnd.n1881 gnd.n1880 0.152939
R14492 gnd.n1882 gnd.n1881 0.152939
R14493 gnd.n1883 gnd.n1882 0.152939
R14494 gnd.n1888 gnd.n1883 0.152939
R14495 gnd.n1889 gnd.n1888 0.152939
R14496 gnd.n1890 gnd.n1889 0.152939
R14497 gnd.n1891 gnd.n1890 0.152939
R14498 gnd.n1896 gnd.n1891 0.152939
R14499 gnd.n1897 gnd.n1896 0.152939
R14500 gnd.n1898 gnd.n1897 0.152939
R14501 gnd.n1899 gnd.n1898 0.152939
R14502 gnd.n1904 gnd.n1899 0.152939
R14503 gnd.n1905 gnd.n1904 0.152939
R14504 gnd.n1906 gnd.n1905 0.152939
R14505 gnd.n1907 gnd.n1906 0.152939
R14506 gnd.n2236 gnd.n1913 0.152939
R14507 gnd.n2236 gnd.n2235 0.152939
R14508 gnd.n2235 gnd.n2234 0.152939
R14509 gnd.n2234 gnd.n1914 0.152939
R14510 gnd.n1919 gnd.n1914 0.152939
R14511 gnd.n1920 gnd.n1919 0.152939
R14512 gnd.n1921 gnd.n1920 0.152939
R14513 gnd.n1926 gnd.n1921 0.152939
R14514 gnd.n1927 gnd.n1926 0.152939
R14515 gnd.n1928 gnd.n1927 0.152939
R14516 gnd.n1929 gnd.n1928 0.152939
R14517 gnd.n1934 gnd.n1929 0.152939
R14518 gnd.n1935 gnd.n1934 0.152939
R14519 gnd.n1936 gnd.n1935 0.152939
R14520 gnd.n1937 gnd.n1936 0.152939
R14521 gnd.n1942 gnd.n1937 0.152939
R14522 gnd.n1943 gnd.n1942 0.152939
R14523 gnd.n1944 gnd.n1943 0.152939
R14524 gnd.n1945 gnd.n1944 0.152939
R14525 gnd.n1950 gnd.n1945 0.152939
R14526 gnd.n1951 gnd.n1950 0.152939
R14527 gnd.n1952 gnd.n1951 0.152939
R14528 gnd.n1953 gnd.n1952 0.152939
R14529 gnd.n1958 gnd.n1953 0.152939
R14530 gnd.n1959 gnd.n1958 0.152939
R14531 gnd.n1960 gnd.n1959 0.152939
R14532 gnd.n1961 gnd.n1960 0.152939
R14533 gnd.n1966 gnd.n1961 0.152939
R14534 gnd.n1967 gnd.n1966 0.152939
R14535 gnd.n1968 gnd.n1967 0.152939
R14536 gnd.n1969 gnd.n1968 0.152939
R14537 gnd.n1974 gnd.n1969 0.152939
R14538 gnd.n1975 gnd.n1974 0.152939
R14539 gnd.n1976 gnd.n1975 0.152939
R14540 gnd.n1977 gnd.n1976 0.152939
R14541 gnd.n1982 gnd.n1977 0.152939
R14542 gnd.n1983 gnd.n1982 0.152939
R14543 gnd.n1984 gnd.n1983 0.152939
R14544 gnd.n1985 gnd.n1984 0.152939
R14545 gnd.n1990 gnd.n1985 0.152939
R14546 gnd.n1991 gnd.n1990 0.152939
R14547 gnd.n1992 gnd.n1991 0.152939
R14548 gnd.n1993 gnd.n1992 0.152939
R14549 gnd.n1998 gnd.n1993 0.152939
R14550 gnd.n1999 gnd.n1998 0.152939
R14551 gnd.n2000 gnd.n1999 0.152939
R14552 gnd.n2001 gnd.n2000 0.152939
R14553 gnd.n2006 gnd.n2001 0.152939
R14554 gnd.n2007 gnd.n2006 0.152939
R14555 gnd.n2008 gnd.n2007 0.152939
R14556 gnd.n2009 gnd.n2008 0.152939
R14557 gnd.n2014 gnd.n2009 0.152939
R14558 gnd.n2015 gnd.n2014 0.152939
R14559 gnd.n2016 gnd.n2015 0.152939
R14560 gnd.n2017 gnd.n2016 0.152939
R14561 gnd.n2022 gnd.n2017 0.152939
R14562 gnd.n2023 gnd.n2022 0.152939
R14563 gnd.n2024 gnd.n2023 0.152939
R14564 gnd.n2025 gnd.n2024 0.152939
R14565 gnd.n2030 gnd.n2025 0.152939
R14566 gnd.n2031 gnd.n2030 0.152939
R14567 gnd.n2032 gnd.n2031 0.152939
R14568 gnd.n2033 gnd.n2032 0.152939
R14569 gnd.n2038 gnd.n2033 0.152939
R14570 gnd.n2039 gnd.n2038 0.152939
R14571 gnd.n2040 gnd.n2039 0.152939
R14572 gnd.n2041 gnd.n2040 0.152939
R14573 gnd.n2046 gnd.n2041 0.152939
R14574 gnd.n2047 gnd.n2046 0.152939
R14575 gnd.n2048 gnd.n2047 0.152939
R14576 gnd.n2049 gnd.n2048 0.152939
R14577 gnd.n2054 gnd.n2049 0.152939
R14578 gnd.n2055 gnd.n2054 0.152939
R14579 gnd.n2056 gnd.n2055 0.152939
R14580 gnd.n2057 gnd.n2056 0.152939
R14581 gnd.n2062 gnd.n2057 0.152939
R14582 gnd.n2063 gnd.n2062 0.152939
R14583 gnd.n2064 gnd.n2063 0.152939
R14584 gnd.n2065 gnd.n2064 0.152939
R14585 gnd.n2071 gnd.n2065 0.152939
R14586 gnd.n2072 gnd.n2071 0.152939
R14587 gnd.n2073 gnd.n2072 0.152939
R14588 gnd.n2073 gnd.n345 0.152939
R14589 gnd.n7078 gnd.n345 0.152939
R14590 gnd.n7186 gnd.n7185 0.152939
R14591 gnd.n7186 gnd.n283 0.152939
R14592 gnd.n7200 gnd.n283 0.152939
R14593 gnd.n7201 gnd.n7200 0.152939
R14594 gnd.n7202 gnd.n7201 0.152939
R14595 gnd.n7202 gnd.n269 0.152939
R14596 gnd.n7216 gnd.n269 0.152939
R14597 gnd.n7217 gnd.n7216 0.152939
R14598 gnd.n7218 gnd.n7217 0.152939
R14599 gnd.n7218 gnd.n253 0.152939
R14600 gnd.n7232 gnd.n253 0.152939
R14601 gnd.n7233 gnd.n7232 0.152939
R14602 gnd.n7234 gnd.n7233 0.152939
R14603 gnd.n7234 gnd.n239 0.152939
R14604 gnd.n7248 gnd.n239 0.152939
R14605 gnd.n7249 gnd.n7248 0.152939
R14606 gnd.n7250 gnd.n7249 0.152939
R14607 gnd.n7250 gnd.n222 0.152939
R14608 gnd.n7264 gnd.n222 0.152939
R14609 gnd.n7265 gnd.n7264 0.152939
R14610 gnd.n7266 gnd.n7265 0.152939
R14611 gnd.n7266 gnd.n206 0.152939
R14612 gnd.n7348 gnd.n206 0.152939
R14613 gnd.n7349 gnd.n7348 0.152939
R14614 gnd.n7350 gnd.n7349 0.152939
R14615 gnd.n7350 gnd.n129 0.152939
R14616 gnd.n7430 gnd.n129 0.152939
R14617 gnd.n7429 gnd.n130 0.152939
R14618 gnd.n132 gnd.n130 0.152939
R14619 gnd.n136 gnd.n132 0.152939
R14620 gnd.n137 gnd.n136 0.152939
R14621 gnd.n138 gnd.n137 0.152939
R14622 gnd.n139 gnd.n138 0.152939
R14623 gnd.n143 gnd.n139 0.152939
R14624 gnd.n144 gnd.n143 0.152939
R14625 gnd.n145 gnd.n144 0.152939
R14626 gnd.n146 gnd.n145 0.152939
R14627 gnd.n150 gnd.n146 0.152939
R14628 gnd.n151 gnd.n150 0.152939
R14629 gnd.n152 gnd.n151 0.152939
R14630 gnd.n153 gnd.n152 0.152939
R14631 gnd.n157 gnd.n153 0.152939
R14632 gnd.n158 gnd.n157 0.152939
R14633 gnd.n159 gnd.n158 0.152939
R14634 gnd.n160 gnd.n159 0.152939
R14635 gnd.n164 gnd.n160 0.152939
R14636 gnd.n165 gnd.n164 0.152939
R14637 gnd.n166 gnd.n165 0.152939
R14638 gnd.n167 gnd.n166 0.152939
R14639 gnd.n171 gnd.n167 0.152939
R14640 gnd.n172 gnd.n171 0.152939
R14641 gnd.n173 gnd.n172 0.152939
R14642 gnd.n174 gnd.n173 0.152939
R14643 gnd.n178 gnd.n174 0.152939
R14644 gnd.n179 gnd.n178 0.152939
R14645 gnd.n180 gnd.n179 0.152939
R14646 gnd.n181 gnd.n180 0.152939
R14647 gnd.n185 gnd.n181 0.152939
R14648 gnd.n186 gnd.n185 0.152939
R14649 gnd.n187 gnd.n186 0.152939
R14650 gnd.n188 gnd.n187 0.152939
R14651 gnd.n192 gnd.n188 0.152939
R14652 gnd.n193 gnd.n192 0.152939
R14653 gnd.n7360 gnd.n193 0.152939
R14654 gnd.n7360 gnd.n7359 0.152939
R14655 gnd.n6704 gnd.n562 0.152939
R14656 gnd.n6705 gnd.n6704 0.152939
R14657 gnd.n6705 gnd.n6702 0.152939
R14658 gnd.n6713 gnd.n6702 0.152939
R14659 gnd.n6714 gnd.n6713 0.152939
R14660 gnd.n6715 gnd.n6714 0.152939
R14661 gnd.n6716 gnd.n6715 0.152939
R14662 gnd.n6718 gnd.n6716 0.152939
R14663 gnd.n6718 gnd.n6717 0.152939
R14664 gnd.n6717 gnd.n597 0.152939
R14665 gnd.n597 gnd.n595 0.152939
R14666 gnd.n6753 gnd.n595 0.152939
R14667 gnd.n6754 gnd.n6753 0.152939
R14668 gnd.n6755 gnd.n6754 0.152939
R14669 gnd.n6756 gnd.n6755 0.152939
R14670 gnd.n6757 gnd.n6756 0.152939
R14671 gnd.n6757 gnd.n586 0.152939
R14672 gnd.n6780 gnd.n586 0.152939
R14673 gnd.n6781 gnd.n6780 0.152939
R14674 gnd.n6782 gnd.n6781 0.152939
R14675 gnd.n6783 gnd.n6782 0.152939
R14676 gnd.n6784 gnd.n6783 0.152939
R14677 gnd.n6785 gnd.n6784 0.152939
R14678 gnd.n6786 gnd.n6785 0.152939
R14679 gnd.n6788 gnd.n6786 0.152939
R14680 gnd.n6788 gnd.n6787 0.152939
R14681 gnd.n6787 gnd.n356 0.152939
R14682 gnd.n7055 gnd.n356 0.152939
R14683 gnd.n7056 gnd.n7055 0.152939
R14684 gnd.n7057 gnd.n7056 0.152939
R14685 gnd.n7058 gnd.n7057 0.152939
R14686 gnd.n7058 gnd.n333 0.152939
R14687 gnd.n7091 gnd.n333 0.152939
R14688 gnd.n7092 gnd.n7091 0.152939
R14689 gnd.n7093 gnd.n7092 0.152939
R14690 gnd.n7094 gnd.n7093 0.152939
R14691 gnd.n7095 gnd.n7094 0.152939
R14692 gnd.n7096 gnd.n7095 0.152939
R14693 gnd.n7097 gnd.n7096 0.152939
R14694 gnd.n7098 gnd.n7097 0.152939
R14695 gnd.n7099 gnd.n7098 0.152939
R14696 gnd.n7100 gnd.n7099 0.152939
R14697 gnd.n7101 gnd.n7100 0.152939
R14698 gnd.n7102 gnd.n7101 0.152939
R14699 gnd.n7103 gnd.n7102 0.152939
R14700 gnd.n7104 gnd.n7103 0.152939
R14701 gnd.n7105 gnd.n7104 0.152939
R14702 gnd.n7106 gnd.n7105 0.152939
R14703 gnd.n7107 gnd.n7106 0.152939
R14704 gnd.n7108 gnd.n7107 0.152939
R14705 gnd.n7109 gnd.n7108 0.152939
R14706 gnd.n7110 gnd.n7109 0.152939
R14707 gnd.n7111 gnd.n7110 0.152939
R14708 gnd.n7112 gnd.n7111 0.152939
R14709 gnd.n7113 gnd.n7112 0.152939
R14710 gnd.n7114 gnd.n7113 0.152939
R14711 gnd.n7115 gnd.n7114 0.152939
R14712 gnd.n7116 gnd.n7115 0.152939
R14713 gnd.n7117 gnd.n7116 0.152939
R14714 gnd.n7118 gnd.n7117 0.152939
R14715 gnd.n7120 gnd.n7118 0.152939
R14716 gnd.n7120 gnd.n7119 0.152939
R14717 gnd.n7119 gnd.n199 0.152939
R14718 gnd.n7358 gnd.n199 0.152939
R14719 gnd.n6910 gnd.n486 0.152939
R14720 gnd.n520 gnd.n486 0.152939
R14721 gnd.n521 gnd.n520 0.152939
R14722 gnd.n522 gnd.n521 0.152939
R14723 gnd.n523 gnd.n522 0.152939
R14724 gnd.n524 gnd.n523 0.152939
R14725 gnd.n525 gnd.n524 0.152939
R14726 gnd.n526 gnd.n525 0.152939
R14727 gnd.n527 gnd.n526 0.152939
R14728 gnd.n528 gnd.n527 0.152939
R14729 gnd.n529 gnd.n528 0.152939
R14730 gnd.n530 gnd.n529 0.152939
R14731 gnd.n531 gnd.n530 0.152939
R14732 gnd.n532 gnd.n531 0.152939
R14733 gnd.n533 gnd.n532 0.152939
R14734 gnd.n540 gnd.n539 0.152939
R14735 gnd.n541 gnd.n540 0.152939
R14736 gnd.n542 gnd.n541 0.152939
R14737 gnd.n543 gnd.n542 0.152939
R14738 gnd.n544 gnd.n543 0.152939
R14739 gnd.n545 gnd.n544 0.152939
R14740 gnd.n546 gnd.n545 0.152939
R14741 gnd.n547 gnd.n546 0.152939
R14742 gnd.n548 gnd.n547 0.152939
R14743 gnd.n549 gnd.n548 0.152939
R14744 gnd.n550 gnd.n549 0.152939
R14745 gnd.n551 gnd.n550 0.152939
R14746 gnd.n552 gnd.n551 0.152939
R14747 gnd.n553 gnd.n552 0.152939
R14748 gnd.n554 gnd.n553 0.152939
R14749 gnd.n555 gnd.n554 0.152939
R14750 gnd.n556 gnd.n555 0.152939
R14751 gnd.n6840 gnd.n556 0.152939
R14752 gnd.n6840 gnd.n6839 0.152939
R14753 gnd.n6839 gnd.n6838 0.152939
R14754 gnd.n6912 gnd.n6911 0.152939
R14755 gnd.n6912 gnd.n468 0.152939
R14756 gnd.n6926 gnd.n468 0.152939
R14757 gnd.n6927 gnd.n6926 0.152939
R14758 gnd.n6928 gnd.n6927 0.152939
R14759 gnd.n6928 gnd.n451 0.152939
R14760 gnd.n6942 gnd.n451 0.152939
R14761 gnd.n6943 gnd.n6942 0.152939
R14762 gnd.n6944 gnd.n6943 0.152939
R14763 gnd.n6944 gnd.n434 0.152939
R14764 gnd.n6958 gnd.n434 0.152939
R14765 gnd.n6959 gnd.n6958 0.152939
R14766 gnd.n6960 gnd.n6959 0.152939
R14767 gnd.n6960 gnd.n417 0.152939
R14768 gnd.n6974 gnd.n417 0.152939
R14769 gnd.n6975 gnd.n6974 0.152939
R14770 gnd.n6976 gnd.n6975 0.152939
R14771 gnd.n6976 gnd.n398 0.152939
R14772 gnd.n6993 gnd.n398 0.152939
R14773 gnd.n6994 gnd.n6993 0.152939
R14774 gnd.n6995 gnd.n6994 0.152939
R14775 gnd.n6995 gnd.n366 0.152939
R14776 gnd.n7044 gnd.n366 0.152939
R14777 gnd.n7045 gnd.n7044 0.152939
R14778 gnd.n7046 gnd.n7045 0.152939
R14779 gnd.n7046 gnd.n299 0.152939
R14780 gnd.n7185 gnd.n299 0.152939
R14781 gnd.n7009 gnd.n7008 0.152939
R14782 gnd.n7008 gnd.n347 0.152939
R14783 gnd.n1215 gnd.n1214 0.152939
R14784 gnd.n4670 gnd.n1215 0.152939
R14785 gnd.n4672 gnd.n4670 0.152939
R14786 gnd.n4673 gnd.n4672 0.152939
R14787 gnd.n4674 gnd.n4673 0.152939
R14788 gnd.n4675 gnd.n4674 0.152939
R14789 gnd.n4676 gnd.n4675 0.152939
R14790 gnd.n4677 gnd.n4676 0.152939
R14791 gnd.n4678 gnd.n4677 0.152939
R14792 gnd.n4678 gnd.n1259 0.152939
R14793 gnd.n4712 gnd.n1259 0.152939
R14794 gnd.n4713 gnd.n4712 0.152939
R14795 gnd.n4714 gnd.n4713 0.152939
R14796 gnd.n4715 gnd.n4714 0.152939
R14797 gnd.n4716 gnd.n4715 0.152939
R14798 gnd.n4717 gnd.n4716 0.152939
R14799 gnd.n4718 gnd.n4717 0.152939
R14800 gnd.n4718 gnd.n1249 0.152939
R14801 gnd.n4751 gnd.n1249 0.152939
R14802 gnd.n4752 gnd.n4751 0.152939
R14803 gnd.n4753 gnd.n4752 0.152939
R14804 gnd.n4754 gnd.n4753 0.152939
R14805 gnd.n4755 gnd.n4754 0.152939
R14806 gnd.n4758 gnd.n4755 0.152939
R14807 gnd.n4759 gnd.n4758 0.152939
R14808 gnd.n4760 gnd.n4759 0.152939
R14809 gnd.n4761 gnd.n4760 0.152939
R14810 gnd.n4765 gnd.n4761 0.152939
R14811 gnd.n4766 gnd.n4765 0.152939
R14812 gnd.n4767 gnd.n4766 0.152939
R14813 gnd.n4768 gnd.n4767 0.152939
R14814 gnd.n4768 gnd.n940 0.152939
R14815 gnd.n6340 gnd.n940 0.152939
R14816 gnd.n6341 gnd.n6340 0.152939
R14817 gnd.n6342 gnd.n6341 0.152939
R14818 gnd.n6342 gnd.n926 0.152939
R14819 gnd.n6356 gnd.n926 0.152939
R14820 gnd.n6357 gnd.n6356 0.152939
R14821 gnd.n6358 gnd.n6357 0.152939
R14822 gnd.n6358 gnd.n912 0.152939
R14823 gnd.n6372 gnd.n912 0.152939
R14824 gnd.n6373 gnd.n6372 0.152939
R14825 gnd.n6374 gnd.n6373 0.152939
R14826 gnd.n6374 gnd.n897 0.152939
R14827 gnd.n6388 gnd.n897 0.152939
R14828 gnd.n6389 gnd.n6388 0.152939
R14829 gnd.n6390 gnd.n6389 0.152939
R14830 gnd.n6390 gnd.n882 0.152939
R14831 gnd.n6404 gnd.n882 0.152939
R14832 gnd.n6405 gnd.n6404 0.152939
R14833 gnd.n6406 gnd.n6405 0.152939
R14834 gnd.n6406 gnd.n866 0.152939
R14835 gnd.n6420 gnd.n866 0.152939
R14836 gnd.n6421 gnd.n6420 0.152939
R14837 gnd.n6422 gnd.n6421 0.152939
R14838 gnd.n6422 gnd.n851 0.152939
R14839 gnd.n6436 gnd.n851 0.152939
R14840 gnd.n6437 gnd.n6436 0.152939
R14841 gnd.n6438 gnd.n6437 0.152939
R14842 gnd.n6438 gnd.n837 0.152939
R14843 gnd.n6452 gnd.n837 0.152939
R14844 gnd.n6453 gnd.n6452 0.152939
R14845 gnd.n6454 gnd.n6453 0.152939
R14846 gnd.n6454 gnd.n822 0.152939
R14847 gnd.n6468 gnd.n822 0.152939
R14848 gnd.n6469 gnd.n6468 0.152939
R14849 gnd.n6470 gnd.n6469 0.152939
R14850 gnd.n6470 gnd.n806 0.152939
R14851 gnd.n6484 gnd.n806 0.152939
R14852 gnd.n6485 gnd.n6484 0.152939
R14853 gnd.n6486 gnd.n6485 0.152939
R14854 gnd.n6486 gnd.n791 0.152939
R14855 gnd.n6500 gnd.n791 0.152939
R14856 gnd.n6501 gnd.n6500 0.152939
R14857 gnd.n6502 gnd.n6501 0.152939
R14858 gnd.n6502 gnd.n776 0.152939
R14859 gnd.n6516 gnd.n776 0.152939
R14860 gnd.n6517 gnd.n6516 0.152939
R14861 gnd.n6518 gnd.n6517 0.152939
R14862 gnd.n6518 gnd.n760 0.152939
R14863 gnd.n6532 gnd.n760 0.152939
R14864 gnd.n6533 gnd.n6532 0.152939
R14865 gnd.n6534 gnd.n6533 0.152939
R14866 gnd.n6534 gnd.n744 0.152939
R14867 gnd.n6548 gnd.n744 0.152939
R14868 gnd.n6549 gnd.n6548 0.152939
R14869 gnd.n6550 gnd.n6549 0.152939
R14870 gnd.n6550 gnd.n730 0.152939
R14871 gnd.n6564 gnd.n730 0.152939
R14872 gnd.n6565 gnd.n6564 0.152939
R14873 gnd.n6566 gnd.n6565 0.152939
R14874 gnd.n6566 gnd.n715 0.152939
R14875 gnd.n6580 gnd.n715 0.152939
R14876 gnd.n6581 gnd.n6580 0.152939
R14877 gnd.n6582 gnd.n6581 0.152939
R14878 gnd.n6582 gnd.n700 0.152939
R14879 gnd.n6596 gnd.n700 0.152939
R14880 gnd.n6597 gnd.n6596 0.152939
R14881 gnd.n6598 gnd.n6597 0.152939
R14882 gnd.n6598 gnd.n686 0.152939
R14883 gnd.n6612 gnd.n686 0.152939
R14884 gnd.n6613 gnd.n6612 0.152939
R14885 gnd.n6614 gnd.n6613 0.152939
R14886 gnd.n6614 gnd.n672 0.152939
R14887 gnd.n6628 gnd.n672 0.152939
R14888 gnd.n6629 gnd.n6628 0.152939
R14889 gnd.n6630 gnd.n6629 0.152939
R14890 gnd.n6630 gnd.n658 0.152939
R14891 gnd.n6644 gnd.n658 0.152939
R14892 gnd.n6645 gnd.n6644 0.152939
R14893 gnd.n6646 gnd.n6645 0.152939
R14894 gnd.n6646 gnd.n643 0.152939
R14895 gnd.n6661 gnd.n643 0.152939
R14896 gnd.n6662 gnd.n6661 0.152939
R14897 gnd.n6663 gnd.n6662 0.152939
R14898 gnd.n6664 gnd.n6663 0.152939
R14899 gnd.n6664 gnd.n613 0.152939
R14900 gnd.n6680 gnd.n613 0.152939
R14901 gnd.n6681 gnd.n6680 0.152939
R14902 gnd.n6682 gnd.n6681 0.152939
R14903 gnd.n6682 gnd.n609 0.152939
R14904 gnd.n6688 gnd.n609 0.152939
R14905 gnd.n6689 gnd.n6688 0.152939
R14906 gnd.n6690 gnd.n6689 0.152939
R14907 gnd.n6690 gnd.n605 0.152939
R14908 gnd.n6696 gnd.n605 0.152939
R14909 gnd.n6697 gnd.n6696 0.152939
R14910 gnd.n6698 gnd.n6697 0.152939
R14911 gnd.n6698 gnd.n601 0.152939
R14912 gnd.n6730 gnd.n601 0.152939
R14913 gnd.n6731 gnd.n6730 0.152939
R14914 gnd.n6732 gnd.n6731 0.152939
R14915 gnd.n6733 gnd.n6732 0.152939
R14916 gnd.n6734 gnd.n6733 0.152939
R14917 gnd.n6735 gnd.n6734 0.152939
R14918 gnd.n6736 gnd.n6735 0.152939
R14919 gnd.n6736 gnd.n591 0.152939
R14920 gnd.n6769 gnd.n591 0.152939
R14921 gnd.n6770 gnd.n6769 0.152939
R14922 gnd.n6771 gnd.n6770 0.152939
R14923 gnd.n6772 gnd.n6771 0.152939
R14924 gnd.n6772 gnd.n391 0.152939
R14925 gnd.n7002 gnd.n391 0.152939
R14926 gnd.n7003 gnd.n7002 0.152939
R14927 gnd.n7004 gnd.n7003 0.152939
R14928 gnd.n7005 gnd.n7004 0.152939
R14929 gnd.n7006 gnd.n7005 0.152939
R14930 gnd.n7007 gnd.n7006 0.152939
R14931 gnd.n7009 gnd.n7007 0.152939
R14932 gnd.n4239 gnd.n4238 0.152939
R14933 gnd.n4240 gnd.n4239 0.152939
R14934 gnd.n4241 gnd.n4240 0.152939
R14935 gnd.n4242 gnd.n4241 0.152939
R14936 gnd.n4243 gnd.n4242 0.152939
R14937 gnd.n4244 gnd.n4243 0.152939
R14938 gnd.n4245 gnd.n4244 0.152939
R14939 gnd.n4246 gnd.n4245 0.152939
R14940 gnd.n4247 gnd.n4246 0.152939
R14941 gnd.n4248 gnd.n4247 0.152939
R14942 gnd.n4249 gnd.n4248 0.152939
R14943 gnd.n4250 gnd.n4249 0.152939
R14944 gnd.n4251 gnd.n4250 0.152939
R14945 gnd.n4252 gnd.n4251 0.152939
R14946 gnd.n4253 gnd.n4252 0.152939
R14947 gnd.n4254 gnd.n4253 0.152939
R14948 gnd.n4255 gnd.n4254 0.152939
R14949 gnd.n4256 gnd.n4255 0.152939
R14950 gnd.n4256 gnd.n1317 0.152939
R14951 gnd.n4575 gnd.n1317 0.152939
R14952 gnd.n4576 gnd.n4575 0.152939
R14953 gnd.n4577 gnd.n4576 0.152939
R14954 gnd.n4578 gnd.n4577 0.152939
R14955 gnd.n4579 gnd.n4578 0.152939
R14956 gnd.n4579 gnd.n1282 0.152939
R14957 gnd.n4614 gnd.n1282 0.152939
R14958 gnd.n4615 gnd.n4614 0.152939
R14959 gnd.n4616 gnd.n4615 0.152939
R14960 gnd.n4617 gnd.n4616 0.152939
R14961 gnd.n4618 gnd.n4617 0.152939
R14962 gnd.n4619 gnd.n4618 0.152939
R14963 gnd.n4190 gnd.n1398 0.152939
R14964 gnd.n4198 gnd.n4190 0.152939
R14965 gnd.n4199 gnd.n4198 0.152939
R14966 gnd.n4200 gnd.n4199 0.152939
R14967 gnd.n4200 gnd.n4186 0.152939
R14968 gnd.n4208 gnd.n4186 0.152939
R14969 gnd.n4209 gnd.n4208 0.152939
R14970 gnd.n4210 gnd.n4209 0.152939
R14971 gnd.n4210 gnd.n4182 0.152939
R14972 gnd.n4218 gnd.n4182 0.152939
R14973 gnd.n4219 gnd.n4218 0.152939
R14974 gnd.n4220 gnd.n4219 0.152939
R14975 gnd.n4220 gnd.n4178 0.152939
R14976 gnd.n4228 gnd.n4178 0.152939
R14977 gnd.n4229 gnd.n4228 0.152939
R14978 gnd.n4230 gnd.n4229 0.152939
R14979 gnd.n4230 gnd.n4172 0.152939
R14980 gnd.n4237 gnd.n4172 0.152939
R14981 gnd.n4486 gnd.n4485 0.152939
R14982 gnd.n4487 gnd.n4486 0.152939
R14983 gnd.n4487 gnd.n1383 0.152939
R14984 gnd.n4501 gnd.n1383 0.152939
R14985 gnd.n4502 gnd.n4501 0.152939
R14986 gnd.n4503 gnd.n4502 0.152939
R14987 gnd.n4503 gnd.n1366 0.152939
R14988 gnd.n4517 gnd.n1366 0.152939
R14989 gnd.n4518 gnd.n4517 0.152939
R14990 gnd.n4519 gnd.n4518 0.152939
R14991 gnd.n4519 gnd.n1351 0.152939
R14992 gnd.n4533 gnd.n1351 0.152939
R14993 gnd.n4534 gnd.n4533 0.152939
R14994 gnd.n4535 gnd.n4534 0.152939
R14995 gnd.n4535 gnd.n1334 0.152939
R14996 gnd.n4549 gnd.n1334 0.152939
R14997 gnd.n4550 gnd.n4549 0.152939
R14998 gnd.n4551 gnd.n4550 0.152939
R14999 gnd.n4552 gnd.n4551 0.152939
R15000 gnd.n4553 gnd.n4552 0.152939
R15001 gnd.n4555 gnd.n4553 0.152939
R15002 gnd.n4555 gnd.n4554 0.152939
R15003 gnd.n4554 gnd.n1300 0.152939
R15004 gnd.n1301 gnd.n1300 0.152939
R15005 gnd.n1302 gnd.n1301 0.152939
R15006 gnd.n1303 gnd.n1302 0.152939
R15007 gnd.n1305 gnd.n1303 0.152939
R15008 gnd.n1305 gnd.n1304 0.152939
R15009 gnd.n1304 gnd.n1191 0.152939
R15010 gnd.n1192 gnd.n1191 0.152939
R15011 gnd.n1193 gnd.n1192 0.152939
R15012 gnd.n1273 gnd.n1193 0.152939
R15013 gnd.n1273 gnd.n1204 0.152939
R15014 gnd.n1205 gnd.n1204 0.152939
R15015 gnd.n1206 gnd.n1205 0.152939
R15016 gnd.n1206 gnd.n1167 0.152939
R15017 gnd.n4887 gnd.n1167 0.152939
R15018 gnd.n4888 gnd.n4887 0.152939
R15019 gnd.n4889 gnd.n4888 0.152939
R15020 gnd.n4889 gnd.n1151 0.152939
R15021 gnd.n4903 gnd.n1151 0.152939
R15022 gnd.n4904 gnd.n4903 0.152939
R15023 gnd.n4905 gnd.n4904 0.152939
R15024 gnd.n4905 gnd.n1133 0.152939
R15025 gnd.n4919 gnd.n1133 0.152939
R15026 gnd.n4920 gnd.n4919 0.152939
R15027 gnd.n4921 gnd.n4920 0.152939
R15028 gnd.n4921 gnd.n1117 0.152939
R15029 gnd.n4935 gnd.n1117 0.152939
R15030 gnd.n4936 gnd.n4935 0.152939
R15031 gnd.n4937 gnd.n4936 0.152939
R15032 gnd.n4937 gnd.n1099 0.152939
R15033 gnd.n4951 gnd.n1099 0.152939
R15034 gnd.n4952 gnd.n4951 0.152939
R15035 gnd.n4953 gnd.n4952 0.152939
R15036 gnd.n4953 gnd.n1083 0.152939
R15037 gnd.n4967 gnd.n1083 0.152939
R15038 gnd.n4968 gnd.n4967 0.152939
R15039 gnd.n4969 gnd.n4968 0.152939
R15040 gnd.n4969 gnd.n1064 0.152939
R15041 gnd.n4985 gnd.n1064 0.152939
R15042 gnd.n4986 gnd.n4985 0.152939
R15043 gnd.n4987 gnd.n4986 0.152939
R15044 gnd.n6221 gnd.n4987 0.152939
R15045 gnd.n4881 gnd.n1159 0.152939
R15046 gnd.n4895 gnd.n1159 0.152939
R15047 gnd.n4896 gnd.n4895 0.152939
R15048 gnd.n4897 gnd.n4896 0.152939
R15049 gnd.n4897 gnd.n1142 0.152939
R15050 gnd.n4911 gnd.n1142 0.152939
R15051 gnd.n4912 gnd.n4911 0.152939
R15052 gnd.n4913 gnd.n4912 0.152939
R15053 gnd.n4913 gnd.n1125 0.152939
R15054 gnd.n4927 gnd.n1125 0.152939
R15055 gnd.n4928 gnd.n4927 0.152939
R15056 gnd.n4929 gnd.n4928 0.152939
R15057 gnd.n4929 gnd.n1108 0.152939
R15058 gnd.n4943 gnd.n1108 0.152939
R15059 gnd.n4944 gnd.n4943 0.152939
R15060 gnd.n4945 gnd.n4944 0.152939
R15061 gnd.n4945 gnd.n1091 0.152939
R15062 gnd.n4959 gnd.n1091 0.152939
R15063 gnd.n4960 gnd.n4959 0.152939
R15064 gnd.n4961 gnd.n4960 0.152939
R15065 gnd.n4961 gnd.n1074 0.152939
R15066 gnd.n4975 gnd.n1074 0.152939
R15067 gnd.n4976 gnd.n4975 0.152939
R15068 gnd.n4977 gnd.n4976 0.152939
R15069 gnd.n4978 gnd.n4977 0.152939
R15070 gnd.n4978 gnd.n989 0.152939
R15071 gnd.n6299 gnd.n989 0.152939
R15072 gnd.n6298 gnd.n990 0.152939
R15073 gnd.n995 gnd.n990 0.152939
R15074 gnd.n996 gnd.n995 0.152939
R15075 gnd.n997 gnd.n996 0.152939
R15076 gnd.n998 gnd.n997 0.152939
R15077 gnd.n999 gnd.n998 0.152939
R15078 gnd.n1003 gnd.n999 0.152939
R15079 gnd.n1004 gnd.n1003 0.152939
R15080 gnd.n1005 gnd.n1004 0.152939
R15081 gnd.n1006 gnd.n1005 0.152939
R15082 gnd.n1010 gnd.n1006 0.152939
R15083 gnd.n1011 gnd.n1010 0.152939
R15084 gnd.n1012 gnd.n1011 0.152939
R15085 gnd.n1013 gnd.n1012 0.152939
R15086 gnd.n1020 gnd.n1013 0.152939
R15087 gnd.n1023 gnd.n1022 0.152939
R15088 gnd.n1024 gnd.n1023 0.152939
R15089 gnd.n1028 gnd.n1024 0.152939
R15090 gnd.n1029 gnd.n1028 0.152939
R15091 gnd.n1030 gnd.n1029 0.152939
R15092 gnd.n1031 gnd.n1030 0.152939
R15093 gnd.n1035 gnd.n1031 0.152939
R15094 gnd.n1036 gnd.n1035 0.152939
R15095 gnd.n1037 gnd.n1036 0.152939
R15096 gnd.n1038 gnd.n1037 0.152939
R15097 gnd.n1042 gnd.n1038 0.152939
R15098 gnd.n1043 gnd.n1042 0.152939
R15099 gnd.n1044 gnd.n1043 0.152939
R15100 gnd.n1045 gnd.n1044 0.152939
R15101 gnd.n1049 gnd.n1045 0.152939
R15102 gnd.n1050 gnd.n1049 0.152939
R15103 gnd.n1051 gnd.n1050 0.152939
R15104 gnd.n1052 gnd.n1051 0.152939
R15105 gnd.n1057 gnd.n1052 0.152939
R15106 gnd.n6230 gnd.n1057 0.152939
R15107 gnd.n4399 gnd.n4347 0.152939
R15108 gnd.n4349 gnd.n4347 0.152939
R15109 gnd.n4350 gnd.n4349 0.152939
R15110 gnd.n4351 gnd.n4350 0.152939
R15111 gnd.n4352 gnd.n4351 0.152939
R15112 gnd.n4353 gnd.n4352 0.152939
R15113 gnd.n4354 gnd.n4353 0.152939
R15114 gnd.n4355 gnd.n4354 0.152939
R15115 gnd.n4356 gnd.n4355 0.152939
R15116 gnd.n4357 gnd.n4356 0.152939
R15117 gnd.n4358 gnd.n4357 0.152939
R15118 gnd.n4359 gnd.n4358 0.152939
R15119 gnd.n4360 gnd.n4359 0.152939
R15120 gnd.n4361 gnd.n4360 0.152939
R15121 gnd.n4362 gnd.n4361 0.152939
R15122 gnd.n4363 gnd.n4362 0.152939
R15123 gnd.n4364 gnd.n4363 0.152939
R15124 gnd.n4365 gnd.n4364 0.152939
R15125 gnd.n4366 gnd.n4365 0.152939
R15126 gnd.n4368 gnd.n4366 0.152939
R15127 gnd.n4368 gnd.n4367 0.152939
R15128 gnd.n4367 gnd.n1311 0.152939
R15129 gnd.n4589 gnd.n1311 0.152939
R15130 gnd.n4590 gnd.n4589 0.152939
R15131 gnd.n4591 gnd.n4590 0.152939
R15132 gnd.n4592 gnd.n4591 0.152939
R15133 gnd.n4592 gnd.n1276 0.152939
R15134 gnd.n4632 gnd.n1276 0.152939
R15135 gnd.n4633 gnd.n4632 0.152939
R15136 gnd.n4634 gnd.n4633 0.152939
R15137 gnd.n4634 gnd.n1274 0.152939
R15138 gnd.n4640 gnd.n1274 0.152939
R15139 gnd.n4641 gnd.n4640 0.152939
R15140 gnd.n4642 gnd.n4641 0.152939
R15141 gnd.n4642 gnd.n1267 0.152939
R15142 gnd.n4656 gnd.n1267 0.152939
R15143 gnd.n4657 gnd.n4656 0.152939
R15144 gnd.n4658 gnd.n4657 0.152939
R15145 gnd.n4658 gnd.n1265 0.152939
R15146 gnd.n4664 gnd.n1265 0.152939
R15147 gnd.n4665 gnd.n4664 0.152939
R15148 gnd.n4666 gnd.n4665 0.152939
R15149 gnd.n4666 gnd.n1263 0.152939
R15150 gnd.n4695 gnd.n1263 0.152939
R15151 gnd.n4696 gnd.n4695 0.152939
R15152 gnd.n4697 gnd.n4696 0.152939
R15153 gnd.n4698 gnd.n4697 0.152939
R15154 gnd.n4700 gnd.n4698 0.152939
R15155 gnd.n4700 gnd.n4699 0.152939
R15156 gnd.n4699 gnd.n1255 0.152939
R15157 gnd.n1255 gnd.n1253 0.152939
R15158 gnd.n4735 gnd.n1253 0.152939
R15159 gnd.n4736 gnd.n4735 0.152939
R15160 gnd.n4737 gnd.n4736 0.152939
R15161 gnd.n4738 gnd.n4737 0.152939
R15162 gnd.n4739 gnd.n4738 0.152939
R15163 gnd.n4739 gnd.n1244 0.152939
R15164 gnd.n4791 gnd.n1244 0.152939
R15165 gnd.n4792 gnd.n4791 0.152939
R15166 gnd.n4793 gnd.n4792 0.152939
R15167 gnd.n4795 gnd.n4793 0.152939
R15168 gnd.n4795 gnd.n4794 0.152939
R15169 gnd.n4794 gnd.n1058 0.152939
R15170 gnd.n6229 gnd.n1058 0.152939
R15171 gnd.n4478 gnd.n4286 0.152939
R15172 gnd.n4289 gnd.n4286 0.152939
R15173 gnd.n4290 gnd.n4289 0.152939
R15174 gnd.n4291 gnd.n4290 0.152939
R15175 gnd.n4294 gnd.n4291 0.152939
R15176 gnd.n4295 gnd.n4294 0.152939
R15177 gnd.n4296 gnd.n4295 0.152939
R15178 gnd.n4297 gnd.n4296 0.152939
R15179 gnd.n4300 gnd.n4297 0.152939
R15180 gnd.n4301 gnd.n4300 0.152939
R15181 gnd.n4302 gnd.n4301 0.152939
R15182 gnd.n4303 gnd.n4302 0.152939
R15183 gnd.n4306 gnd.n4303 0.152939
R15184 gnd.n4307 gnd.n4306 0.152939
R15185 gnd.n4308 gnd.n4307 0.152939
R15186 gnd.n4309 gnd.n4308 0.152939
R15187 gnd.n4315 gnd.n4309 0.152939
R15188 gnd.n4316 gnd.n4315 0.152939
R15189 gnd.n4317 gnd.n4316 0.152939
R15190 gnd.n4318 gnd.n4317 0.152939
R15191 gnd.n4321 gnd.n4318 0.152939
R15192 gnd.n4322 gnd.n4321 0.152939
R15193 gnd.n4323 gnd.n4322 0.152939
R15194 gnd.n4324 gnd.n4323 0.152939
R15195 gnd.n4327 gnd.n4324 0.152939
R15196 gnd.n4328 gnd.n4327 0.152939
R15197 gnd.n4329 gnd.n4328 0.152939
R15198 gnd.n4330 gnd.n4329 0.152939
R15199 gnd.n4333 gnd.n4330 0.152939
R15200 gnd.n4334 gnd.n4333 0.152939
R15201 gnd.n4335 gnd.n4334 0.152939
R15202 gnd.n4336 gnd.n4335 0.152939
R15203 gnd.n4339 gnd.n4336 0.152939
R15204 gnd.n4340 gnd.n4339 0.152939
R15205 gnd.n4341 gnd.n4340 0.152939
R15206 gnd.n4406 gnd.n4341 0.152939
R15207 gnd.n4406 gnd.n4405 0.152939
R15208 gnd.n4405 gnd.n4404 0.152939
R15209 gnd.n4479 gnd.n1391 0.152939
R15210 gnd.n4493 gnd.n1391 0.152939
R15211 gnd.n4494 gnd.n4493 0.152939
R15212 gnd.n4495 gnd.n4494 0.152939
R15213 gnd.n4495 gnd.n1375 0.152939
R15214 gnd.n4509 gnd.n1375 0.152939
R15215 gnd.n4510 gnd.n4509 0.152939
R15216 gnd.n4511 gnd.n4510 0.152939
R15217 gnd.n4511 gnd.n1359 0.152939
R15218 gnd.n4525 gnd.n1359 0.152939
R15219 gnd.n4526 gnd.n4525 0.152939
R15220 gnd.n4527 gnd.n4526 0.152939
R15221 gnd.n4527 gnd.n1343 0.152939
R15222 gnd.n4541 gnd.n1343 0.152939
R15223 gnd.n4542 gnd.n4541 0.152939
R15224 gnd.n4543 gnd.n4542 0.152939
R15225 gnd.n4543 gnd.n1326 0.152939
R15226 gnd.n4565 gnd.n1326 0.152939
R15227 gnd.n4566 gnd.n4565 0.152939
R15228 gnd.n4567 gnd.n4566 0.152939
R15229 gnd.n4568 gnd.n4567 0.152939
R15230 gnd.n4568 gnd.n1290 0.152939
R15231 gnd.n4605 gnd.n1290 0.152939
R15232 gnd.n4606 gnd.n4605 0.152939
R15233 gnd.n4607 gnd.n4606 0.152939
R15234 gnd.n4607 gnd.n1176 0.152939
R15235 gnd.n4881 gnd.n1176 0.152939
R15236 gnd.n1214 gnd.n1213 0.152939
R15237 gnd.n2558 gnd.n1598 0.152939
R15238 gnd.n2559 gnd.n2558 0.152939
R15239 gnd.n2560 gnd.n2559 0.152939
R15240 gnd.n2560 gnd.n1592 0.152939
R15241 gnd.n2568 gnd.n1592 0.152939
R15242 gnd.n2569 gnd.n2568 0.152939
R15243 gnd.n2570 gnd.n2569 0.152939
R15244 gnd.n2570 gnd.n1586 0.152939
R15245 gnd.n2578 gnd.n1586 0.152939
R15246 gnd.n2579 gnd.n2578 0.152939
R15247 gnd.n2580 gnd.n2579 0.152939
R15248 gnd.n2580 gnd.n1580 0.152939
R15249 gnd.n2588 gnd.n1580 0.152939
R15250 gnd.n2589 gnd.n2588 0.152939
R15251 gnd.n2590 gnd.n2589 0.152939
R15252 gnd.n2590 gnd.n1574 0.152939
R15253 gnd.n2598 gnd.n1574 0.152939
R15254 gnd.n2599 gnd.n2598 0.152939
R15255 gnd.n2600 gnd.n2599 0.152939
R15256 gnd.n2600 gnd.n1568 0.152939
R15257 gnd.n2608 gnd.n1568 0.152939
R15258 gnd.n2609 gnd.n2608 0.152939
R15259 gnd.n2610 gnd.n2609 0.152939
R15260 gnd.n2610 gnd.n1562 0.152939
R15261 gnd.n2618 gnd.n1562 0.152939
R15262 gnd.n2619 gnd.n2618 0.152939
R15263 gnd.n2620 gnd.n2619 0.152939
R15264 gnd.n2620 gnd.n1556 0.152939
R15265 gnd.n2628 gnd.n1556 0.152939
R15266 gnd.n2629 gnd.n2628 0.152939
R15267 gnd.n2630 gnd.n2629 0.152939
R15268 gnd.n2630 gnd.n1550 0.152939
R15269 gnd.n2638 gnd.n1550 0.152939
R15270 gnd.n2639 gnd.n2638 0.152939
R15271 gnd.n2640 gnd.n2639 0.152939
R15272 gnd.n2640 gnd.n1544 0.152939
R15273 gnd.n2648 gnd.n1544 0.152939
R15274 gnd.n2649 gnd.n2648 0.152939
R15275 gnd.n2650 gnd.n2649 0.152939
R15276 gnd.n2650 gnd.n1538 0.152939
R15277 gnd.n2658 gnd.n1538 0.152939
R15278 gnd.n2659 gnd.n2658 0.152939
R15279 gnd.n2660 gnd.n2659 0.152939
R15280 gnd.n2660 gnd.n1532 0.152939
R15281 gnd.n2668 gnd.n1532 0.152939
R15282 gnd.n2669 gnd.n2668 0.152939
R15283 gnd.n2670 gnd.n2669 0.152939
R15284 gnd.n2670 gnd.n1526 0.152939
R15285 gnd.n2678 gnd.n1526 0.152939
R15286 gnd.n2679 gnd.n2678 0.152939
R15287 gnd.n2680 gnd.n2679 0.152939
R15288 gnd.n2680 gnd.n1520 0.152939
R15289 gnd.n2688 gnd.n1520 0.152939
R15290 gnd.n2689 gnd.n2688 0.152939
R15291 gnd.n2690 gnd.n2689 0.152939
R15292 gnd.n2690 gnd.n1514 0.152939
R15293 gnd.n2698 gnd.n1514 0.152939
R15294 gnd.n2699 gnd.n2698 0.152939
R15295 gnd.n2700 gnd.n2699 0.152939
R15296 gnd.n2700 gnd.n1508 0.152939
R15297 gnd.n2708 gnd.n1508 0.152939
R15298 gnd.n2709 gnd.n2708 0.152939
R15299 gnd.n2710 gnd.n2709 0.152939
R15300 gnd.n2710 gnd.n1502 0.152939
R15301 gnd.n2718 gnd.n1502 0.152939
R15302 gnd.n2719 gnd.n2718 0.152939
R15303 gnd.n2720 gnd.n2719 0.152939
R15304 gnd.n2720 gnd.n1496 0.152939
R15305 gnd.n2728 gnd.n1496 0.152939
R15306 gnd.n2729 gnd.n2728 0.152939
R15307 gnd.n2730 gnd.n2729 0.152939
R15308 gnd.n2730 gnd.n1490 0.152939
R15309 gnd.n2738 gnd.n1490 0.152939
R15310 gnd.n2739 gnd.n2738 0.152939
R15311 gnd.n2740 gnd.n2739 0.152939
R15312 gnd.n2740 gnd.n1484 0.152939
R15313 gnd.n2748 gnd.n1484 0.152939
R15314 gnd.n2749 gnd.n2748 0.152939
R15315 gnd.n2750 gnd.n2749 0.152939
R15316 gnd.n2750 gnd.n1478 0.152939
R15317 gnd.n2758 gnd.n1478 0.152939
R15318 gnd.n2759 gnd.n2758 0.152939
R15319 gnd.n2760 gnd.n2759 0.152939
R15320 gnd.n2762 gnd.n2760 0.152939
R15321 gnd.n6039 gnd.n6038 0.152939
R15322 gnd.n6038 gnd.n6037 0.152939
R15323 gnd.n6037 gnd.n6017 0.152939
R15324 gnd.n6033 gnd.n6017 0.152939
R15325 gnd.n6033 gnd.n6032 0.152939
R15326 gnd.n6032 gnd.n6031 0.152939
R15327 gnd.n6031 gnd.n6023 0.152939
R15328 gnd.n6023 gnd.n634 0.152939
R15329 gnd.n6673 gnd.n634 0.152939
R15330 gnd.n6348 gnd.n933 0.152939
R15331 gnd.n6349 gnd.n6348 0.152939
R15332 gnd.n6350 gnd.n6349 0.152939
R15333 gnd.n6350 gnd.n918 0.152939
R15334 gnd.n6364 gnd.n918 0.152939
R15335 gnd.n6365 gnd.n6364 0.152939
R15336 gnd.n6366 gnd.n6365 0.152939
R15337 gnd.n6366 gnd.n904 0.152939
R15338 gnd.n6380 gnd.n904 0.152939
R15339 gnd.n6381 gnd.n6380 0.152939
R15340 gnd.n6382 gnd.n6381 0.152939
R15341 gnd.n6382 gnd.n890 0.152939
R15342 gnd.n6396 gnd.n890 0.152939
R15343 gnd.n6397 gnd.n6396 0.152939
R15344 gnd.n6398 gnd.n6397 0.152939
R15345 gnd.n6398 gnd.n874 0.152939
R15346 gnd.n6412 gnd.n874 0.152939
R15347 gnd.n6413 gnd.n6412 0.152939
R15348 gnd.n6414 gnd.n6413 0.152939
R15349 gnd.n6414 gnd.n859 0.152939
R15350 gnd.n6428 gnd.n859 0.152939
R15351 gnd.n6429 gnd.n6428 0.152939
R15352 gnd.n6430 gnd.n6429 0.152939
R15353 gnd.n6430 gnd.n844 0.152939
R15354 gnd.n6444 gnd.n844 0.152939
R15355 gnd.n6445 gnd.n6444 0.152939
R15356 gnd.n6446 gnd.n6445 0.152939
R15357 gnd.n6446 gnd.n830 0.152939
R15358 gnd.n6460 gnd.n830 0.152939
R15359 gnd.n6461 gnd.n6460 0.152939
R15360 gnd.n6462 gnd.n6461 0.152939
R15361 gnd.n6462 gnd.n814 0.152939
R15362 gnd.n6476 gnd.n814 0.152939
R15363 gnd.n6477 gnd.n6476 0.152939
R15364 gnd.n6478 gnd.n6477 0.152939
R15365 gnd.n6478 gnd.n798 0.152939
R15366 gnd.n6492 gnd.n798 0.152939
R15367 gnd.n6493 gnd.n6492 0.152939
R15368 gnd.n6494 gnd.n6493 0.152939
R15369 gnd.n6494 gnd.n783 0.152939
R15370 gnd.n6508 gnd.n783 0.152939
R15371 gnd.n6509 gnd.n6508 0.152939
R15372 gnd.n6510 gnd.n6509 0.152939
R15373 gnd.n6510 gnd.n768 0.152939
R15374 gnd.n6524 gnd.n768 0.152939
R15375 gnd.n6525 gnd.n6524 0.152939
R15376 gnd.n6526 gnd.n6525 0.152939
R15377 gnd.n6526 gnd.n752 0.152939
R15378 gnd.n6540 gnd.n752 0.152939
R15379 gnd.n6541 gnd.n6540 0.152939
R15380 gnd.n6542 gnd.n6541 0.152939
R15381 gnd.n6542 gnd.n737 0.152939
R15382 gnd.n6556 gnd.n737 0.152939
R15383 gnd.n6557 gnd.n6556 0.152939
R15384 gnd.n6558 gnd.n6557 0.152939
R15385 gnd.n6558 gnd.n723 0.152939
R15386 gnd.n6572 gnd.n723 0.152939
R15387 gnd.n6573 gnd.n6572 0.152939
R15388 gnd.n6574 gnd.n6573 0.152939
R15389 gnd.n6574 gnd.n708 0.152939
R15390 gnd.n6588 gnd.n708 0.152939
R15391 gnd.n6589 gnd.n6588 0.152939
R15392 gnd.n6590 gnd.n6589 0.152939
R15393 gnd.n6590 gnd.n693 0.152939
R15394 gnd.n6604 gnd.n693 0.152939
R15395 gnd.n6605 gnd.n6604 0.152939
R15396 gnd.n6606 gnd.n6605 0.152939
R15397 gnd.n6606 gnd.n678 0.152939
R15398 gnd.n6620 gnd.n678 0.152939
R15399 gnd.n6621 gnd.n6620 0.152939
R15400 gnd.n6622 gnd.n6621 0.152939
R15401 gnd.n6622 gnd.n665 0.152939
R15402 gnd.n6636 gnd.n665 0.152939
R15403 gnd.n6637 gnd.n6636 0.152939
R15404 gnd.n6638 gnd.n6637 0.152939
R15405 gnd.n6638 gnd.n651 0.152939
R15406 gnd.n6652 gnd.n651 0.152939
R15407 gnd.n6653 gnd.n6652 0.152939
R15408 gnd.n6655 gnd.n6653 0.152939
R15409 gnd.n6655 gnd.n6654 0.152939
R15410 gnd.n6654 gnd.n635 0.152939
R15411 gnd.n6672 gnd.n635 0.152939
R15412 gnd.n6316 gnd.n6315 0.152939
R15413 gnd.n6316 gnd.n966 0.152939
R15414 gnd.n6322 gnd.n966 0.152939
R15415 gnd.n6323 gnd.n6322 0.152939
R15416 gnd.n6324 gnd.n6323 0.152939
R15417 gnd.n6324 gnd.n960 0.152939
R15418 gnd.n6331 gnd.n960 0.152939
R15419 gnd.n6332 gnd.n6331 0.152939
R15420 gnd.n6333 gnd.n6332 0.152939
R15421 gnd.n4648 gnd.n1270 0.152939
R15422 gnd.n4649 gnd.n4648 0.152939
R15423 gnd.n4650 gnd.n4649 0.152939
R15424 gnd.n4650 gnd.n1221 0.152939
R15425 gnd.n4841 gnd.n1221 0.152939
R15426 gnd.n4841 gnd.n4840 0.152939
R15427 gnd.n4840 gnd.n4839 0.152939
R15428 gnd.n4839 gnd.n1222 0.152939
R15429 gnd.n4835 gnd.n1222 0.152939
R15430 gnd.n4835 gnd.n4834 0.152939
R15431 gnd.n4834 gnd.n4833 0.152939
R15432 gnd.n4833 gnd.n1226 0.152939
R15433 gnd.n4829 gnd.n1226 0.152939
R15434 gnd.n4829 gnd.n4828 0.152939
R15435 gnd.n4828 gnd.n4827 0.152939
R15436 gnd.n4827 gnd.n1230 0.152939
R15437 gnd.n4823 gnd.n1230 0.152939
R15438 gnd.n4823 gnd.n4822 0.152939
R15439 gnd.n4822 gnd.n4821 0.152939
R15440 gnd.n4821 gnd.n1234 0.152939
R15441 gnd.n4817 gnd.n1234 0.152939
R15442 gnd.n4817 gnd.n4816 0.152939
R15443 gnd.n4816 gnd.n4815 0.152939
R15444 gnd.n4815 gnd.n1238 0.152939
R15445 gnd.n4811 gnd.n1238 0.152939
R15446 gnd.n4811 gnd.n4810 0.152939
R15447 gnd.n4810 gnd.n4809 0.152939
R15448 gnd.n4809 gnd.n1242 0.152939
R15449 gnd.n4805 gnd.n1242 0.152939
R15450 gnd.n4805 gnd.n4804 0.152939
R15451 gnd.n4804 gnd.n970 0.152939
R15452 gnd.n6218 gnd.n4990 0.152939
R15453 gnd.n6214 gnd.n4990 0.152939
R15454 gnd.n6214 gnd.n6213 0.152939
R15455 gnd.n6213 gnd.n6212 0.152939
R15456 gnd.n6212 gnd.n5097 0.152939
R15457 gnd.n6208 gnd.n5097 0.152939
R15458 gnd.n6208 gnd.n6207 0.152939
R15459 gnd.n6207 gnd.n6206 0.152939
R15460 gnd.n6206 gnd.n5101 0.152939
R15461 gnd.n6202 gnd.n5101 0.152939
R15462 gnd.n6202 gnd.n6201 0.152939
R15463 gnd.n6201 gnd.n6200 0.152939
R15464 gnd.n6200 gnd.n5105 0.152939
R15465 gnd.n6196 gnd.n5105 0.152939
R15466 gnd.n6196 gnd.n6195 0.152939
R15467 gnd.n6195 gnd.n6194 0.152939
R15468 gnd.n6194 gnd.n5109 0.152939
R15469 gnd.n6190 gnd.n5109 0.152939
R15470 gnd.n6190 gnd.n6189 0.152939
R15471 gnd.n6189 gnd.n6188 0.152939
R15472 gnd.n6188 gnd.n5113 0.152939
R15473 gnd.n6184 gnd.n5113 0.152939
R15474 gnd.n6184 gnd.n6183 0.152939
R15475 gnd.n6183 gnd.n6182 0.152939
R15476 gnd.n6182 gnd.n5117 0.152939
R15477 gnd.n6178 gnd.n5117 0.152939
R15478 gnd.n6178 gnd.n6177 0.152939
R15479 gnd.n6177 gnd.n6176 0.152939
R15480 gnd.n6176 gnd.n5121 0.152939
R15481 gnd.n6172 gnd.n5121 0.152939
R15482 gnd.n6172 gnd.n6171 0.152939
R15483 gnd.n6171 gnd.n6170 0.152939
R15484 gnd.n6170 gnd.n5125 0.152939
R15485 gnd.n6166 gnd.n5125 0.152939
R15486 gnd.n6166 gnd.n6165 0.152939
R15487 gnd.n6165 gnd.n6164 0.152939
R15488 gnd.n6164 gnd.n5129 0.152939
R15489 gnd.n6160 gnd.n5129 0.152939
R15490 gnd.n6160 gnd.n6159 0.152939
R15491 gnd.n6159 gnd.n6158 0.152939
R15492 gnd.n6158 gnd.n5133 0.152939
R15493 gnd.n6154 gnd.n5133 0.152939
R15494 gnd.n6154 gnd.n6153 0.152939
R15495 gnd.n6153 gnd.n6152 0.152939
R15496 gnd.n6152 gnd.n5137 0.152939
R15497 gnd.n6148 gnd.n5137 0.152939
R15498 gnd.n6148 gnd.n6147 0.152939
R15499 gnd.n6147 gnd.n6146 0.152939
R15500 gnd.n6146 gnd.n5141 0.152939
R15501 gnd.n6142 gnd.n5141 0.152939
R15502 gnd.n6142 gnd.n6141 0.152939
R15503 gnd.n6141 gnd.n6140 0.152939
R15504 gnd.n6140 gnd.n5145 0.152939
R15505 gnd.n6136 gnd.n5145 0.152939
R15506 gnd.n6136 gnd.n6135 0.152939
R15507 gnd.n6135 gnd.n6134 0.152939
R15508 gnd.n6134 gnd.n5149 0.152939
R15509 gnd.n6130 gnd.n5149 0.152939
R15510 gnd.n6130 gnd.n6129 0.152939
R15511 gnd.n6129 gnd.n6128 0.152939
R15512 gnd.n6128 gnd.n5153 0.152939
R15513 gnd.n6124 gnd.n5153 0.152939
R15514 gnd.n6124 gnd.n6123 0.152939
R15515 gnd.n6123 gnd.n6122 0.152939
R15516 gnd.n6122 gnd.n5157 0.152939
R15517 gnd.n6118 gnd.n5157 0.152939
R15518 gnd.n6118 gnd.n6117 0.152939
R15519 gnd.n6117 gnd.n6116 0.152939
R15520 gnd.n6116 gnd.n5161 0.152939
R15521 gnd.n6112 gnd.n5161 0.152939
R15522 gnd.n6112 gnd.n6111 0.152939
R15523 gnd.n6111 gnd.n6110 0.152939
R15524 gnd.n6110 gnd.n5940 0.152939
R15525 gnd.n6106 gnd.n5940 0.152939
R15526 gnd.n6106 gnd.n6105 0.152939
R15527 gnd.n6105 gnd.n6104 0.152939
R15528 gnd.n6104 gnd.n5944 0.152939
R15529 gnd.n6100 gnd.n5944 0.152939
R15530 gnd.n6100 gnd.n6099 0.152939
R15531 gnd.n6099 gnd.n6098 0.152939
R15532 gnd.n6098 gnd.n5948 0.152939
R15533 gnd.n5950 gnd.n5948 0.152939
R15534 gnd.n6918 gnd.n477 0.152939
R15535 gnd.n6919 gnd.n6918 0.152939
R15536 gnd.n6920 gnd.n6919 0.152939
R15537 gnd.n6920 gnd.n459 0.152939
R15538 gnd.n6934 gnd.n459 0.152939
R15539 gnd.n6935 gnd.n6934 0.152939
R15540 gnd.n6936 gnd.n6935 0.152939
R15541 gnd.n6936 gnd.n443 0.152939
R15542 gnd.n6950 gnd.n443 0.152939
R15543 gnd.n6951 gnd.n6950 0.152939
R15544 gnd.n6952 gnd.n6951 0.152939
R15545 gnd.n6952 gnd.n425 0.152939
R15546 gnd.n6966 gnd.n425 0.152939
R15547 gnd.n6967 gnd.n6966 0.152939
R15548 gnd.n6968 gnd.n6967 0.152939
R15549 gnd.n6968 gnd.n409 0.152939
R15550 gnd.n6982 gnd.n409 0.152939
R15551 gnd.n6983 gnd.n6982 0.152939
R15552 gnd.n6987 gnd.n6983 0.152939
R15553 gnd.n6987 gnd.n6986 0.152939
R15554 gnd.n6986 gnd.n6985 0.152939
R15555 gnd.n6985 gnd.n377 0.152939
R15556 gnd.n7038 gnd.n377 0.152939
R15557 gnd.n7038 gnd.n7037 0.152939
R15558 gnd.n7037 gnd.n7036 0.152939
R15559 gnd.n7036 gnd.n378 0.152939
R15560 gnd.n7032 gnd.n378 0.152939
R15561 gnd.n7032 gnd.n316 0.152939
R15562 gnd.n7177 gnd.n316 0.152939
R15563 gnd.n7177 gnd.n7176 0.152939
R15564 gnd.n7176 gnd.n7175 0.152939
R15565 gnd.n7175 gnd.n317 0.152939
R15566 gnd.n7171 gnd.n317 0.152939
R15567 gnd.n7171 gnd.n7170 0.152939
R15568 gnd.n7170 gnd.n7169 0.152939
R15569 gnd.n7169 gnd.n322 0.152939
R15570 gnd.n322 gnd.n292 0.152939
R15571 gnd.n7192 gnd.n292 0.152939
R15572 gnd.n7193 gnd.n7192 0.152939
R15573 gnd.n7194 gnd.n7193 0.152939
R15574 gnd.n7194 gnd.n276 0.152939
R15575 gnd.n7208 gnd.n276 0.152939
R15576 gnd.n7209 gnd.n7208 0.152939
R15577 gnd.n7210 gnd.n7209 0.152939
R15578 gnd.n7210 gnd.n262 0.152939
R15579 gnd.n7224 gnd.n262 0.152939
R15580 gnd.n7225 gnd.n7224 0.152939
R15581 gnd.n7226 gnd.n7225 0.152939
R15582 gnd.n7226 gnd.n246 0.152939
R15583 gnd.n7240 gnd.n246 0.152939
R15584 gnd.n7241 gnd.n7240 0.152939
R15585 gnd.n7242 gnd.n7241 0.152939
R15586 gnd.n7242 gnd.n231 0.152939
R15587 gnd.n7256 gnd.n231 0.152939
R15588 gnd.n7257 gnd.n7256 0.152939
R15589 gnd.n7258 gnd.n7257 0.152939
R15590 gnd.n7258 gnd.n216 0.152939
R15591 gnd.n7272 gnd.n216 0.152939
R15592 gnd.n7273 gnd.n7272 0.152939
R15593 gnd.n7342 gnd.n7273 0.152939
R15594 gnd.n7342 gnd.n7341 0.152939
R15595 gnd.n7341 gnd.n7340 0.152939
R15596 gnd.n7340 gnd.n7274 0.152939
R15597 gnd.n7336 gnd.n7274 0.152939
R15598 gnd.n7335 gnd.n7276 0.152939
R15599 gnd.n7331 gnd.n7276 0.152939
R15600 gnd.n7331 gnd.n7330 0.152939
R15601 gnd.n7330 gnd.n7329 0.152939
R15602 gnd.n7329 gnd.n7282 0.152939
R15603 gnd.n7325 gnd.n7282 0.152939
R15604 gnd.n7325 gnd.n7324 0.152939
R15605 gnd.n7324 gnd.n7323 0.152939
R15606 gnd.n7323 gnd.n7290 0.152939
R15607 gnd.n7319 gnd.n7290 0.152939
R15608 gnd.n7319 gnd.n7318 0.152939
R15609 gnd.n7318 gnd.n7317 0.152939
R15610 gnd.n7317 gnd.n7298 0.152939
R15611 gnd.n7313 gnd.n7298 0.152939
R15612 gnd.n7313 gnd.n7312 0.152939
R15613 gnd.n7312 gnd.n7311 0.152939
R15614 gnd.n7311 gnd.n117 0.152939
R15615 gnd.n7437 gnd.n117 0.152939
R15616 gnd.n6831 gnd.n6830 0.152939
R15617 gnd.n6830 gnd.n6829 0.152939
R15618 gnd.n6829 gnd.n567 0.152939
R15619 gnd.n6825 gnd.n567 0.152939
R15620 gnd.n6825 gnd.n6824 0.152939
R15621 gnd.n6824 gnd.n6823 0.152939
R15622 gnd.n6823 gnd.n571 0.152939
R15623 gnd.n6819 gnd.n571 0.152939
R15624 gnd.n6819 gnd.n6818 0.152939
R15625 gnd.n6818 gnd.n6817 0.152939
R15626 gnd.n6817 gnd.n575 0.152939
R15627 gnd.n6813 gnd.n575 0.152939
R15628 gnd.n6813 gnd.n6812 0.152939
R15629 gnd.n6812 gnd.n6811 0.152939
R15630 gnd.n6811 gnd.n579 0.152939
R15631 gnd.n6807 gnd.n579 0.152939
R15632 gnd.n6807 gnd.n6806 0.152939
R15633 gnd.n6806 gnd.n6805 0.152939
R15634 gnd.n6805 gnd.n583 0.152939
R15635 gnd.n6801 gnd.n583 0.152939
R15636 gnd.n6801 gnd.n6800 0.152939
R15637 gnd.n6800 gnd.n383 0.152939
R15638 gnd.n7023 gnd.n383 0.152939
R15639 gnd.n7024 gnd.n7023 0.152939
R15640 gnd.n7026 gnd.n7024 0.152939
R15641 gnd.n7026 gnd.n7025 0.152939
R15642 gnd.n7025 gnd.n354 0.152939
R15643 gnd.n7068 gnd.n354 0.152939
R15644 gnd.n7068 gnd.n7067 0.152939
R15645 gnd.n7067 gnd.n7066 0.152939
R15646 gnd.n7066 gnd.n75 0.152939
R15647 gnd.n7486 gnd.n75 0.152939
R15648 gnd.n7486 gnd.n7485 0.152939
R15649 gnd.n7485 gnd.n77 0.152939
R15650 gnd.n7481 gnd.n77 0.152939
R15651 gnd.n7481 gnd.n7480 0.152939
R15652 gnd.n7480 gnd.n7479 0.152939
R15653 gnd.n7479 gnd.n82 0.152939
R15654 gnd.n7475 gnd.n82 0.152939
R15655 gnd.n7475 gnd.n7474 0.152939
R15656 gnd.n7474 gnd.n7473 0.152939
R15657 gnd.n7473 gnd.n87 0.152939
R15658 gnd.n7469 gnd.n87 0.152939
R15659 gnd.n7469 gnd.n7468 0.152939
R15660 gnd.n7468 gnd.n7467 0.152939
R15661 gnd.n7467 gnd.n92 0.152939
R15662 gnd.n7463 gnd.n92 0.152939
R15663 gnd.n7463 gnd.n7462 0.152939
R15664 gnd.n7462 gnd.n7461 0.152939
R15665 gnd.n7461 gnd.n97 0.152939
R15666 gnd.n7457 gnd.n97 0.152939
R15667 gnd.n7457 gnd.n7456 0.152939
R15668 gnd.n7456 gnd.n7455 0.152939
R15669 gnd.n7455 gnd.n102 0.152939
R15670 gnd.n7451 gnd.n102 0.152939
R15671 gnd.n7451 gnd.n7450 0.152939
R15672 gnd.n7450 gnd.n7449 0.152939
R15673 gnd.n7449 gnd.n107 0.152939
R15674 gnd.n7445 gnd.n107 0.152939
R15675 gnd.n7445 gnd.n7444 0.152939
R15676 gnd.n7444 gnd.n7443 0.152939
R15677 gnd.n7443 gnd.n112 0.152939
R15678 gnd.n7439 gnd.n112 0.152939
R15679 gnd.n7439 gnd.n7438 0.152939
R15680 gnd.n6039 gnd.n566 0.151415
R15681 gnd.n6315 gnd.n6314 0.151415
R15682 gnd.n4621 gnd.n4619 0.145814
R15683 gnd.n4621 gnd.n1270 0.145814
R15684 gnd.n347 gnd.n300 0.130073
R15685 gnd.n1213 gnd.n1177 0.130073
R15686 gnd.n3601 gnd.n2947 0.0767195
R15687 gnd.n3601 gnd.n3600 0.0767195
R15688 gnd.n6220 gnd.n6219 0.063
R15689 gnd.n5955 gnd.n5954 0.063
R15690 gnd.n4131 gnd.n1441 0.0477147
R15691 gnd.n3391 gnd.n3279 0.0442063
R15692 gnd.n3392 gnd.n3391 0.0442063
R15693 gnd.n3393 gnd.n3392 0.0442063
R15694 gnd.n3393 gnd.n3268 0.0442063
R15695 gnd.n3407 gnd.n3268 0.0442063
R15696 gnd.n3408 gnd.n3407 0.0442063
R15697 gnd.n3409 gnd.n3408 0.0442063
R15698 gnd.n3409 gnd.n3255 0.0442063
R15699 gnd.n3453 gnd.n3255 0.0442063
R15700 gnd.n3454 gnd.n3453 0.0442063
R15701 gnd.n3456 gnd.n3189 0.0344674
R15702 gnd.n6043 gnd.n6011 0.0344674
R15703 gnd.n6313 gnd.n971 0.0344674
R15704 gnd.n3476 gnd.n3475 0.0269946
R15705 gnd.n3478 gnd.n3477 0.0269946
R15706 gnd.n3184 gnd.n3182 0.0269946
R15707 gnd.n3488 gnd.n3486 0.0269946
R15708 gnd.n3487 gnd.n3163 0.0269946
R15709 gnd.n3507 gnd.n3506 0.0269946
R15710 gnd.n3509 gnd.n3508 0.0269946
R15711 gnd.n3158 gnd.n3157 0.0269946
R15712 gnd.n3519 gnd.n3153 0.0269946
R15713 gnd.n3518 gnd.n3155 0.0269946
R15714 gnd.n3154 gnd.n3134 0.0269946
R15715 gnd.n3545 gnd.n3135 0.0269946
R15716 gnd.n3544 gnd.n3136 0.0269946
R15717 gnd.n3564 gnd.n3120 0.0269946
R15718 gnd.n3566 gnd.n3565 0.0269946
R15719 gnd.n3567 gnd.n3100 0.0269946
R15720 gnd.n3568 gnd.n3101 0.0269946
R15721 gnd.n3569 gnd.n3102 0.0269946
R15722 gnd.n3104 gnd.n3103 0.0269946
R15723 gnd.n2941 gnd.n2939 0.0269946
R15724 gnd.n3613 gnd.n3611 0.0269946
R15725 gnd.n3612 gnd.n2923 0.0269946
R15726 gnd.n3632 gnd.n3631 0.0269946
R15727 gnd.n3634 gnd.n3633 0.0269946
R15728 gnd.n2918 gnd.n2916 0.0269946
R15729 gnd.n3644 gnd.n3642 0.0269946
R15730 gnd.n3643 gnd.n2898 0.0269946
R15731 gnd.n3663 gnd.n3662 0.0269946
R15732 gnd.n3665 gnd.n3664 0.0269946
R15733 gnd.n2892 gnd.n2890 0.0269946
R15734 gnd.n3675 gnd.n3673 0.0269946
R15735 gnd.n3674 gnd.n2871 0.0269946
R15736 gnd.n3694 gnd.n3693 0.0269946
R15737 gnd.n3696 gnd.n3695 0.0269946
R15738 gnd.n2866 gnd.n2864 0.0269946
R15739 gnd.n3706 gnd.n3704 0.0269946
R15740 gnd.n3705 gnd.n2847 0.0269946
R15741 gnd.n3725 gnd.n3724 0.0269946
R15742 gnd.n3727 gnd.n3726 0.0269946
R15743 gnd.n2842 gnd.n2840 0.0269946
R15744 gnd.n3737 gnd.n3735 0.0269946
R15745 gnd.n3736 gnd.n2821 0.0269946
R15746 gnd.n3756 gnd.n3755 0.0269946
R15747 gnd.n3758 gnd.n3757 0.0269946
R15748 gnd.n2816 gnd.n2814 0.0269946
R15749 gnd.n3768 gnd.n3766 0.0269946
R15750 gnd.n3767 gnd.n2796 0.0269946
R15751 gnd.n3787 gnd.n3786 0.0269946
R15752 gnd.n2790 gnd.n2788 0.0269946
R15753 gnd.n4055 gnd.n4053 0.0269946
R15754 gnd.n4054 gnd.n2770 0.0269946
R15755 gnd.n4073 gnd.n4072 0.0269946
R15756 gnd.n5954 gnd.n5952 0.0246168
R15757 gnd.n6219 gnd.n4989 0.0246168
R15758 gnd.n7077 gnd.n300 0.0233659
R15759 gnd.n2761 gnd.n1177 0.0233659
R15760 gnd.n3456 gnd.n3455 0.0202011
R15761 gnd.n6091 gnd.n5952 0.0174837
R15762 gnd.n6091 gnd.n6090 0.0174837
R15763 gnd.n6090 gnd.n5953 0.0174837
R15764 gnd.n6087 gnd.n5953 0.0174837
R15765 gnd.n6087 gnd.n6086 0.0174837
R15766 gnd.n6086 gnd.n5964 0.0174837
R15767 gnd.n6083 gnd.n5964 0.0174837
R15768 gnd.n6083 gnd.n6082 0.0174837
R15769 gnd.n6082 gnd.n5970 0.0174837
R15770 gnd.n6079 gnd.n5970 0.0174837
R15771 gnd.n6079 gnd.n6078 0.0174837
R15772 gnd.n6078 gnd.n5974 0.0174837
R15773 gnd.n6075 gnd.n5974 0.0174837
R15774 gnd.n6075 gnd.n6074 0.0174837
R15775 gnd.n6074 gnd.n5978 0.0174837
R15776 gnd.n6071 gnd.n5978 0.0174837
R15777 gnd.n6071 gnd.n6070 0.0174837
R15778 gnd.n6070 gnd.n5984 0.0174837
R15779 gnd.n6067 gnd.n5984 0.0174837
R15780 gnd.n6067 gnd.n6066 0.0174837
R15781 gnd.n6066 gnd.n5990 0.0174837
R15782 gnd.n6063 gnd.n5990 0.0174837
R15783 gnd.n6063 gnd.n6062 0.0174837
R15784 gnd.n6062 gnd.n5994 0.0174837
R15785 gnd.n6059 gnd.n5994 0.0174837
R15786 gnd.n6059 gnd.n6058 0.0174837
R15787 gnd.n6058 gnd.n5998 0.0174837
R15788 gnd.n6055 gnd.n5998 0.0174837
R15789 gnd.n6055 gnd.n6054 0.0174837
R15790 gnd.n6054 gnd.n6004 0.0174837
R15791 gnd.n6051 gnd.n6004 0.0174837
R15792 gnd.n6051 gnd.n6050 0.0174837
R15793 gnd.n6050 gnd.n6010 0.0174837
R15794 gnd.n6044 gnd.n6010 0.0174837
R15795 gnd.n6044 gnd.n6043 0.0174837
R15796 gnd.n4991 gnd.n4989 0.0174837
R15797 gnd.n4995 gnd.n4991 0.0174837
R15798 gnd.n5090 gnd.n4995 0.0174837
R15799 gnd.n5090 gnd.n5089 0.0174837
R15800 gnd.n5089 gnd.n4996 0.0174837
R15801 gnd.n5086 gnd.n4996 0.0174837
R15802 gnd.n5086 gnd.n5085 0.0174837
R15803 gnd.n5085 gnd.n5007 0.0174837
R15804 gnd.n5082 gnd.n5007 0.0174837
R15805 gnd.n5082 gnd.n5081 0.0174837
R15806 gnd.n5081 gnd.n5011 0.0174837
R15807 gnd.n5078 gnd.n5011 0.0174837
R15808 gnd.n5078 gnd.n5077 0.0174837
R15809 gnd.n5077 gnd.n5017 0.0174837
R15810 gnd.n5074 gnd.n5017 0.0174837
R15811 gnd.n5074 gnd.n5073 0.0174837
R15812 gnd.n5073 gnd.n5023 0.0174837
R15813 gnd.n5070 gnd.n5023 0.0174837
R15814 gnd.n5070 gnd.n5069 0.0174837
R15815 gnd.n5069 gnd.n5030 0.0174837
R15816 gnd.n5066 gnd.n5030 0.0174837
R15817 gnd.n5066 gnd.n5065 0.0174837
R15818 gnd.n5065 gnd.n5034 0.0174837
R15819 gnd.n5062 gnd.n5034 0.0174837
R15820 gnd.n5062 gnd.n5061 0.0174837
R15821 gnd.n5061 gnd.n5040 0.0174837
R15822 gnd.n5058 gnd.n5040 0.0174837
R15823 gnd.n5058 gnd.n5057 0.0174837
R15824 gnd.n5057 gnd.n5046 0.0174837
R15825 gnd.n5054 gnd.n5046 0.0174837
R15826 gnd.n5054 gnd.n5053 0.0174837
R15827 gnd.n5053 gnd.n975 0.0174837
R15828 gnd.n6307 gnd.n975 0.0174837
R15829 gnd.n6307 gnd.n6306 0.0174837
R15830 gnd.n6306 gnd.n971 0.0174837
R15831 gnd.n3455 gnd.n3454 0.0148637
R15832 gnd.n4044 gnd.n3788 0.0144266
R15833 gnd.n4045 gnd.n4044 0.0130679
R15834 gnd.n3475 gnd.n3189 0.00797283
R15835 gnd.n3477 gnd.n3476 0.00797283
R15836 gnd.n3478 gnd.n3184 0.00797283
R15837 gnd.n3486 gnd.n3182 0.00797283
R15838 gnd.n3488 gnd.n3487 0.00797283
R15839 gnd.n3506 gnd.n3163 0.00797283
R15840 gnd.n3508 gnd.n3507 0.00797283
R15841 gnd.n3509 gnd.n3158 0.00797283
R15842 gnd.n3157 gnd.n3153 0.00797283
R15843 gnd.n3519 gnd.n3518 0.00797283
R15844 gnd.n3155 gnd.n3154 0.00797283
R15845 gnd.n3135 gnd.n3134 0.00797283
R15846 gnd.n3545 gnd.n3544 0.00797283
R15847 gnd.n3136 gnd.n3120 0.00797283
R15848 gnd.n3565 gnd.n3564 0.00797283
R15849 gnd.n3567 gnd.n3566 0.00797283
R15850 gnd.n3568 gnd.n3100 0.00797283
R15851 gnd.n3569 gnd.n3101 0.00797283
R15852 gnd.n3103 gnd.n3102 0.00797283
R15853 gnd.n3104 gnd.n2941 0.00797283
R15854 gnd.n3611 gnd.n2939 0.00797283
R15855 gnd.n3613 gnd.n3612 0.00797283
R15856 gnd.n3631 gnd.n2923 0.00797283
R15857 gnd.n3633 gnd.n3632 0.00797283
R15858 gnd.n3634 gnd.n2918 0.00797283
R15859 gnd.n3642 gnd.n2916 0.00797283
R15860 gnd.n3644 gnd.n3643 0.00797283
R15861 gnd.n3662 gnd.n2898 0.00797283
R15862 gnd.n3664 gnd.n3663 0.00797283
R15863 gnd.n3665 gnd.n2892 0.00797283
R15864 gnd.n3673 gnd.n2890 0.00797283
R15865 gnd.n3675 gnd.n3674 0.00797283
R15866 gnd.n3693 gnd.n2871 0.00797283
R15867 gnd.n3695 gnd.n3694 0.00797283
R15868 gnd.n3696 gnd.n2866 0.00797283
R15869 gnd.n3704 gnd.n2864 0.00797283
R15870 gnd.n3706 gnd.n3705 0.00797283
R15871 gnd.n3724 gnd.n2847 0.00797283
R15872 gnd.n3726 gnd.n3725 0.00797283
R15873 gnd.n3727 gnd.n2842 0.00797283
R15874 gnd.n3735 gnd.n2840 0.00797283
R15875 gnd.n3737 gnd.n3736 0.00797283
R15876 gnd.n3755 gnd.n2821 0.00797283
R15877 gnd.n3757 gnd.n3756 0.00797283
R15878 gnd.n3758 gnd.n2816 0.00797283
R15879 gnd.n3766 gnd.n2814 0.00797283
R15880 gnd.n3768 gnd.n3767 0.00797283
R15881 gnd.n3786 gnd.n2796 0.00797283
R15882 gnd.n3788 gnd.n3787 0.00797283
R15883 gnd.n4045 gnd.n2790 0.00797283
R15884 gnd.n4053 gnd.n2788 0.00797283
R15885 gnd.n4055 gnd.n4054 0.00797283
R15886 gnd.n4072 gnd.n2770 0.00797283
R15887 gnd.n4073 gnd.n1441 0.00797283
R15888 gnd.n333 gnd.n317 0.00433921
R15889 gnd.n4640 gnd.n1273 0.00433921
R15890 gnd.n6011 gnd.n566 0.000839674
R15891 gnd.n6314 gnd.n6313 0.000839674
R15892 a_n6972_8799.n173 a_n6972_8799.t50 485.149
R15893 a_n6972_8799.n189 a_n6972_8799.t62 485.149
R15894 a_n6972_8799.n206 a_n6972_8799.t110 485.149
R15895 a_n6972_8799.n122 a_n6972_8799.t106 485.149
R15896 a_n6972_8799.n138 a_n6972_8799.t117 485.149
R15897 a_n6972_8799.n155 a_n6972_8799.t109 485.149
R15898 a_n6972_8799.n183 a_n6972_8799.t71 464.166
R15899 a_n6972_8799.n182 a_n6972_8799.t70 464.166
R15900 a_n6972_8799.n168 a_n6972_8799.t48 464.166
R15901 a_n6972_8799.n181 a_n6972_8799.t107 464.166
R15902 a_n6972_8799.n180 a_n6972_8799.t72 464.166
R15903 a_n6972_8799.n169 a_n6972_8799.t54 464.166
R15904 a_n6972_8799.n179 a_n6972_8799.t111 464.166
R15905 a_n6972_8799.n178 a_n6972_8799.t86 464.166
R15906 a_n6972_8799.n170 a_n6972_8799.t84 464.166
R15907 a_n6972_8799.n177 a_n6972_8799.t31 464.166
R15908 a_n6972_8799.n176 a_n6972_8799.t90 464.166
R15909 a_n6972_8799.n171 a_n6972_8799.t89 464.166
R15910 a_n6972_8799.n175 a_n6972_8799.t33 464.166
R15911 a_n6972_8799.n174 a_n6972_8799.t32 464.166
R15912 a_n6972_8799.n172 a_n6972_8799.t103 464.166
R15913 a_n6972_8799.n199 a_n6972_8799.t78 464.166
R15914 a_n6972_8799.n198 a_n6972_8799.t77 464.166
R15915 a_n6972_8799.n184 a_n6972_8799.t61 464.166
R15916 a_n6972_8799.n197 a_n6972_8799.t119 464.166
R15917 a_n6972_8799.n196 a_n6972_8799.t83 464.166
R15918 a_n6972_8799.n185 a_n6972_8799.t63 464.166
R15919 a_n6972_8799.n195 a_n6972_8799.t123 464.166
R15920 a_n6972_8799.n194 a_n6972_8799.t96 464.166
R15921 a_n6972_8799.n186 a_n6972_8799.t95 464.166
R15922 a_n6972_8799.n193 a_n6972_8799.t40 464.166
R15923 a_n6972_8799.n192 a_n6972_8799.t99 464.166
R15924 a_n6972_8799.n187 a_n6972_8799.t98 464.166
R15925 a_n6972_8799.n191 a_n6972_8799.t44 464.166
R15926 a_n6972_8799.n190 a_n6972_8799.t43 464.166
R15927 a_n6972_8799.n188 a_n6972_8799.t114 464.166
R15928 a_n6972_8799.n216 a_n6972_8799.t122 464.166
R15929 a_n6972_8799.n215 a_n6972_8799.t42 464.166
R15930 a_n6972_8799.n201 a_n6972_8799.t82 464.166
R15931 a_n6972_8799.n214 a_n6972_8799.t30 464.166
R15932 a_n6972_8799.n213 a_n6972_8799.t102 464.166
R15933 a_n6972_8799.n202 a_n6972_8799.t52 464.166
R15934 a_n6972_8799.n212 a_n6972_8799.t88 464.166
R15935 a_n6972_8799.n211 a_n6972_8799.t35 464.166
R15936 a_n6972_8799.n203 a_n6972_8799.t56 464.166
R15937 a_n6972_8799.n210 a_n6972_8799.t118 464.166
R15938 a_n6972_8799.n209 a_n6972_8799.t94 464.166
R15939 a_n6972_8799.n204 a_n6972_8799.t113 464.166
R15940 a_n6972_8799.n208 a_n6972_8799.t80 464.166
R15941 a_n6972_8799.n207 a_n6972_8799.t97 464.166
R15942 a_n6972_8799.n205 a_n6972_8799.t46 464.166
R15943 a_n6972_8799.n121 a_n6972_8799.t68 464.166
R15944 a_n6972_8799.n124 a_n6972_8799.t69 464.166
R15945 a_n6972_8799.n120 a_n6972_8799.t92 464.166
R15946 a_n6972_8799.n125 a_n6972_8799.t59 464.166
R15947 a_n6972_8799.n126 a_n6972_8799.t60 464.166
R15948 a_n6972_8799.n127 a_n6972_8799.t91 464.166
R15949 a_n6972_8799.n128 a_n6972_8799.t28 464.166
R15950 a_n6972_8799.n119 a_n6972_8799.t57 464.166
R15951 a_n6972_8799.n129 a_n6972_8799.t74 464.166
R15952 a_n6972_8799.n130 a_n6972_8799.t108 464.166
R15953 a_n6972_8799.n131 a_n6972_8799.t39 464.166
R15954 a_n6972_8799.n132 a_n6972_8799.t55 464.166
R15955 a_n6972_8799.n118 a_n6972_8799.t105 464.166
R15956 a_n6972_8799.n133 a_n6972_8799.t36 464.166
R15957 a_n6972_8799.n137 a_n6972_8799.t75 464.166
R15958 a_n6972_8799.n140 a_n6972_8799.t76 464.166
R15959 a_n6972_8799.n136 a_n6972_8799.t104 464.166
R15960 a_n6972_8799.n141 a_n6972_8799.t66 464.166
R15961 a_n6972_8799.n142 a_n6972_8799.t67 464.166
R15962 a_n6972_8799.n143 a_n6972_8799.t100 464.166
R15963 a_n6972_8799.n144 a_n6972_8799.t38 464.166
R15964 a_n6972_8799.n135 a_n6972_8799.t65 464.166
R15965 a_n6972_8799.n145 a_n6972_8799.t85 464.166
R15966 a_n6972_8799.n146 a_n6972_8799.t120 464.166
R15967 a_n6972_8799.n147 a_n6972_8799.t53 464.166
R15968 a_n6972_8799.n148 a_n6972_8799.t64 464.166
R15969 a_n6972_8799.n134 a_n6972_8799.t115 464.166
R15970 a_n6972_8799.n149 a_n6972_8799.t47 464.166
R15971 a_n6972_8799.n154 a_n6972_8799.t45 464.166
R15972 a_n6972_8799.n157 a_n6972_8799.t29 464.166
R15973 a_n6972_8799.n153 a_n6972_8799.t79 464.166
R15974 a_n6972_8799.n158 a_n6972_8799.t112 464.166
R15975 a_n6972_8799.n159 a_n6972_8799.t93 464.166
R15976 a_n6972_8799.n160 a_n6972_8799.t116 464.166
R15977 a_n6972_8799.n161 a_n6972_8799.t73 464.166
R15978 a_n6972_8799.n152 a_n6972_8799.t34 464.166
R15979 a_n6972_8799.n162 a_n6972_8799.t87 464.166
R15980 a_n6972_8799.n163 a_n6972_8799.t51 464.166
R15981 a_n6972_8799.n164 a_n6972_8799.t101 464.166
R15982 a_n6972_8799.n165 a_n6972_8799.t58 464.166
R15983 a_n6972_8799.n151 a_n6972_8799.t81 464.166
R15984 a_n6972_8799.n166 a_n6972_8799.t41 464.166
R15985 a_n6972_8799.n51 a_n6972_8799.n33 74.4178
R15986 a_n6972_8799.n174 a_n6972_8799.n51 12.4674
R15987 a_n6972_8799.n50 a_n6972_8799.n33 80.107
R15988 a_n6972_8799.n50 a_n6972_8799.n175 1.08907
R15989 a_n6972_8799.n34 a_n6972_8799.n49 75.3623
R15990 a_n6972_8799.n48 a_n6972_8799.n34 70.3058
R15991 a_n6972_8799.n36 a_n6972_8799.n47 70.1674
R15992 a_n6972_8799.n47 a_n6972_8799.n170 20.9683
R15993 a_n6972_8799.n46 a_n6972_8799.n36 75.0448
R15994 a_n6972_8799.n178 a_n6972_8799.n46 11.2134
R15995 a_n6972_8799.n45 a_n6972_8799.n35 80.4688
R15996 a_n6972_8799.n35 a_n6972_8799.n44 74.73
R15997 a_n6972_8799.n43 a_n6972_8799.n37 70.1674
R15998 a_n6972_8799.n181 a_n6972_8799.n43 20.9683
R15999 a_n6972_8799.n37 a_n6972_8799.n42 70.5844
R16000 a_n6972_8799.n42 a_n6972_8799.n168 20.1342
R16001 a_n6972_8799.n41 a_n6972_8799.n38 75.6825
R16002 a_n6972_8799.n182 a_n6972_8799.n41 9.93802
R16003 a_n6972_8799.n38 a_n6972_8799.n183 161.3
R16004 a_n6972_8799.n62 a_n6972_8799.n27 74.4178
R16005 a_n6972_8799.n190 a_n6972_8799.n62 12.4674
R16006 a_n6972_8799.n61 a_n6972_8799.n27 80.107
R16007 a_n6972_8799.n61 a_n6972_8799.n191 1.08907
R16008 a_n6972_8799.n28 a_n6972_8799.n60 75.3623
R16009 a_n6972_8799.n59 a_n6972_8799.n28 70.3058
R16010 a_n6972_8799.n30 a_n6972_8799.n58 70.1674
R16011 a_n6972_8799.n58 a_n6972_8799.n186 20.9683
R16012 a_n6972_8799.n57 a_n6972_8799.n30 75.0448
R16013 a_n6972_8799.n194 a_n6972_8799.n57 11.2134
R16014 a_n6972_8799.n56 a_n6972_8799.n29 80.4688
R16015 a_n6972_8799.n29 a_n6972_8799.n55 74.73
R16016 a_n6972_8799.n54 a_n6972_8799.n31 70.1674
R16017 a_n6972_8799.n197 a_n6972_8799.n54 20.9683
R16018 a_n6972_8799.n31 a_n6972_8799.n53 70.5844
R16019 a_n6972_8799.n53 a_n6972_8799.n184 20.1342
R16020 a_n6972_8799.n52 a_n6972_8799.n32 75.6825
R16021 a_n6972_8799.n198 a_n6972_8799.n52 9.93802
R16022 a_n6972_8799.n32 a_n6972_8799.n199 161.3
R16023 a_n6972_8799.n73 a_n6972_8799.n21 74.4178
R16024 a_n6972_8799.n207 a_n6972_8799.n73 12.4674
R16025 a_n6972_8799.n72 a_n6972_8799.n21 80.107
R16026 a_n6972_8799.n72 a_n6972_8799.n208 1.08907
R16027 a_n6972_8799.n22 a_n6972_8799.n71 75.3623
R16028 a_n6972_8799.n70 a_n6972_8799.n22 70.3058
R16029 a_n6972_8799.n24 a_n6972_8799.n69 70.1674
R16030 a_n6972_8799.n69 a_n6972_8799.n203 20.9683
R16031 a_n6972_8799.n68 a_n6972_8799.n24 75.0448
R16032 a_n6972_8799.n211 a_n6972_8799.n68 11.2134
R16033 a_n6972_8799.n67 a_n6972_8799.n23 80.4688
R16034 a_n6972_8799.n23 a_n6972_8799.n66 74.73
R16035 a_n6972_8799.n65 a_n6972_8799.n25 70.1674
R16036 a_n6972_8799.n214 a_n6972_8799.n65 20.9683
R16037 a_n6972_8799.n25 a_n6972_8799.n64 70.5844
R16038 a_n6972_8799.n64 a_n6972_8799.n201 20.1342
R16039 a_n6972_8799.n63 a_n6972_8799.n26 75.6825
R16040 a_n6972_8799.n215 a_n6972_8799.n63 9.93802
R16041 a_n6972_8799.n26 a_n6972_8799.n216 161.3
R16042 a_n6972_8799.n16 a_n6972_8799.n84 70.1674
R16043 a_n6972_8799.n133 a_n6972_8799.n84 20.9683
R16044 a_n6972_8799.n83 a_n6972_8799.n16 74.4178
R16045 a_n6972_8799.n83 a_n6972_8799.n118 12.4674
R16046 a_n6972_8799.n15 a_n6972_8799.n82 80.107
R16047 a_n6972_8799.n132 a_n6972_8799.n82 1.08907
R16048 a_n6972_8799.n81 a_n6972_8799.n15 75.3623
R16049 a_n6972_8799.n17 a_n6972_8799.n80 70.3058
R16050 a_n6972_8799.n79 a_n6972_8799.n17 70.1674
R16051 a_n6972_8799.n79 a_n6972_8799.n119 20.9683
R16052 a_n6972_8799.n18 a_n6972_8799.n78 75.0448
R16053 a_n6972_8799.n128 a_n6972_8799.n78 11.2134
R16054 a_n6972_8799.n77 a_n6972_8799.n18 80.4688
R16055 a_n6972_8799.n19 a_n6972_8799.n76 74.73
R16056 a_n6972_8799.n75 a_n6972_8799.n19 70.1674
R16057 a_n6972_8799.n75 a_n6972_8799.n120 20.9683
R16058 a_n6972_8799.n20 a_n6972_8799.n74 70.5844
R16059 a_n6972_8799.n124 a_n6972_8799.n74 20.1342
R16060 a_n6972_8799.n123 a_n6972_8799.n20 161.3
R16061 a_n6972_8799.n10 a_n6972_8799.n95 70.1674
R16062 a_n6972_8799.n149 a_n6972_8799.n95 20.9683
R16063 a_n6972_8799.n94 a_n6972_8799.n10 74.4178
R16064 a_n6972_8799.n94 a_n6972_8799.n134 12.4674
R16065 a_n6972_8799.n9 a_n6972_8799.n93 80.107
R16066 a_n6972_8799.n148 a_n6972_8799.n93 1.08907
R16067 a_n6972_8799.n92 a_n6972_8799.n9 75.3623
R16068 a_n6972_8799.n11 a_n6972_8799.n91 70.3058
R16069 a_n6972_8799.n90 a_n6972_8799.n11 70.1674
R16070 a_n6972_8799.n90 a_n6972_8799.n135 20.9683
R16071 a_n6972_8799.n12 a_n6972_8799.n89 75.0448
R16072 a_n6972_8799.n144 a_n6972_8799.n89 11.2134
R16073 a_n6972_8799.n88 a_n6972_8799.n12 80.4688
R16074 a_n6972_8799.n13 a_n6972_8799.n87 74.73
R16075 a_n6972_8799.n86 a_n6972_8799.n13 70.1674
R16076 a_n6972_8799.n86 a_n6972_8799.n136 20.9683
R16077 a_n6972_8799.n14 a_n6972_8799.n85 70.5844
R16078 a_n6972_8799.n140 a_n6972_8799.n85 20.1342
R16079 a_n6972_8799.n139 a_n6972_8799.n14 161.3
R16080 a_n6972_8799.n4 a_n6972_8799.n106 70.1674
R16081 a_n6972_8799.n166 a_n6972_8799.n106 20.9683
R16082 a_n6972_8799.n105 a_n6972_8799.n4 74.4178
R16083 a_n6972_8799.n105 a_n6972_8799.n151 12.4674
R16084 a_n6972_8799.n3 a_n6972_8799.n104 80.107
R16085 a_n6972_8799.n165 a_n6972_8799.n104 1.08907
R16086 a_n6972_8799.n103 a_n6972_8799.n3 75.3623
R16087 a_n6972_8799.n5 a_n6972_8799.n102 70.3058
R16088 a_n6972_8799.n101 a_n6972_8799.n5 70.1674
R16089 a_n6972_8799.n101 a_n6972_8799.n152 20.9683
R16090 a_n6972_8799.n6 a_n6972_8799.n100 75.0448
R16091 a_n6972_8799.n161 a_n6972_8799.n100 11.2134
R16092 a_n6972_8799.n99 a_n6972_8799.n6 80.4688
R16093 a_n6972_8799.n7 a_n6972_8799.n98 74.73
R16094 a_n6972_8799.n97 a_n6972_8799.n7 70.1674
R16095 a_n6972_8799.n97 a_n6972_8799.n153 20.9683
R16096 a_n6972_8799.n8 a_n6972_8799.n96 70.5844
R16097 a_n6972_8799.n157 a_n6972_8799.n96 20.1342
R16098 a_n6972_8799.n156 a_n6972_8799.n8 161.3
R16099 a_n6972_8799.n39 a_n6972_8799.n107 98.9633
R16100 a_n6972_8799.n40 a_n6972_8799.n222 98.9631
R16101 a_n6972_8799.n40 a_n6972_8799.n221 98.6055
R16102 a_n6972_8799.n39 a_n6972_8799.n109 98.6055
R16103 a_n6972_8799.n39 a_n6972_8799.n108 98.6055
R16104 a_n6972_8799.n223 a_n6972_8799.n40 98.6054
R16105 a_n6972_8799.n1 a_n6972_8799.n110 81.4626
R16106 a_n6972_8799.n2 a_n6972_8799.n114 81.4626
R16107 a_n6972_8799.n2 a_n6972_8799.n112 81.4626
R16108 a_n6972_8799.n0 a_n6972_8799.n116 80.9324
R16109 a_n6972_8799.n1 a_n6972_8799.n117 80.9324
R16110 a_n6972_8799.n1 a_n6972_8799.n111 80.9324
R16111 a_n6972_8799.n2 a_n6972_8799.n115 80.9324
R16112 a_n6972_8799.n2 a_n6972_8799.n113 80.9324
R16113 a_n6972_8799.n33 a_n6972_8799.n173 70.4033
R16114 a_n6972_8799.n27 a_n6972_8799.n189 70.4033
R16115 a_n6972_8799.n21 a_n6972_8799.n206 70.4033
R16116 a_n6972_8799.n20 a_n6972_8799.n122 70.4033
R16117 a_n6972_8799.n14 a_n6972_8799.n138 70.4033
R16118 a_n6972_8799.n8 a_n6972_8799.n155 70.4033
R16119 a_n6972_8799.n183 a_n6972_8799.n182 48.2005
R16120 a_n6972_8799.n43 a_n6972_8799.n180 20.9683
R16121 a_n6972_8799.n179 a_n6972_8799.n178 48.2005
R16122 a_n6972_8799.n177 a_n6972_8799.n47 20.9683
R16123 a_n6972_8799.n175 a_n6972_8799.n171 48.2005
R16124 a_n6972_8799.n199 a_n6972_8799.n198 48.2005
R16125 a_n6972_8799.n54 a_n6972_8799.n196 20.9683
R16126 a_n6972_8799.n195 a_n6972_8799.n194 48.2005
R16127 a_n6972_8799.n193 a_n6972_8799.n58 20.9683
R16128 a_n6972_8799.n191 a_n6972_8799.n187 48.2005
R16129 a_n6972_8799.n216 a_n6972_8799.n215 48.2005
R16130 a_n6972_8799.n65 a_n6972_8799.n213 20.9683
R16131 a_n6972_8799.n212 a_n6972_8799.n211 48.2005
R16132 a_n6972_8799.n210 a_n6972_8799.n69 20.9683
R16133 a_n6972_8799.n208 a_n6972_8799.n204 48.2005
R16134 a_n6972_8799.n125 a_n6972_8799.n75 20.9683
R16135 a_n6972_8799.n128 a_n6972_8799.n127 48.2005
R16136 a_n6972_8799.n129 a_n6972_8799.n79 20.9683
R16137 a_n6972_8799.n132 a_n6972_8799.n131 48.2005
R16138 a_n6972_8799.t37 a_n6972_8799.n84 485.135
R16139 a_n6972_8799.n141 a_n6972_8799.n86 20.9683
R16140 a_n6972_8799.n144 a_n6972_8799.n143 48.2005
R16141 a_n6972_8799.n145 a_n6972_8799.n90 20.9683
R16142 a_n6972_8799.n148 a_n6972_8799.n147 48.2005
R16143 a_n6972_8799.t49 a_n6972_8799.n95 485.135
R16144 a_n6972_8799.n158 a_n6972_8799.n97 20.9683
R16145 a_n6972_8799.n161 a_n6972_8799.n160 48.2005
R16146 a_n6972_8799.n162 a_n6972_8799.n101 20.9683
R16147 a_n6972_8799.n165 a_n6972_8799.n164 48.2005
R16148 a_n6972_8799.t121 a_n6972_8799.n106 485.135
R16149 a_n6972_8799.n45 a_n6972_8799.n169 47.835
R16150 a_n6972_8799.n48 a_n6972_8799.n176 20.6913
R16151 a_n6972_8799.n56 a_n6972_8799.n185 47.835
R16152 a_n6972_8799.n59 a_n6972_8799.n192 20.6913
R16153 a_n6972_8799.n67 a_n6972_8799.n202 47.835
R16154 a_n6972_8799.n70 a_n6972_8799.n209 20.6913
R16155 a_n6972_8799.n126 a_n6972_8799.n77 47.835
R16156 a_n6972_8799.n130 a_n6972_8799.n80 20.6913
R16157 a_n6972_8799.n142 a_n6972_8799.n88 47.835
R16158 a_n6972_8799.n146 a_n6972_8799.n91 20.6913
R16159 a_n6972_8799.n159 a_n6972_8799.n99 47.835
R16160 a_n6972_8799.n163 a_n6972_8799.n102 20.6913
R16161 a_n6972_8799.n181 a_n6972_8799.n42 22.3251
R16162 a_n6972_8799.n197 a_n6972_8799.n53 22.3251
R16163 a_n6972_8799.n214 a_n6972_8799.n64 22.3251
R16164 a_n6972_8799.n120 a_n6972_8799.n74 22.3251
R16165 a_n6972_8799.n136 a_n6972_8799.n85 22.3251
R16166 a_n6972_8799.n153 a_n6972_8799.n96 22.3251
R16167 a_n6972_8799.n51 a_n6972_8799.n172 33.6462
R16168 a_n6972_8799.n62 a_n6972_8799.n188 33.6462
R16169 a_n6972_8799.n73 a_n6972_8799.n205 33.6462
R16170 a_n6972_8799.n124 a_n6972_8799.n123 27.0217
R16171 a_n6972_8799.n133 a_n6972_8799.n83 33.6462
R16172 a_n6972_8799.n140 a_n6972_8799.n139 27.0217
R16173 a_n6972_8799.n149 a_n6972_8799.n94 33.6462
R16174 a_n6972_8799.n157 a_n6972_8799.n156 27.0217
R16175 a_n6972_8799.n166 a_n6972_8799.n105 33.6462
R16176 a_n6972_8799.n44 a_n6972_8799.n169 11.843
R16177 a_n6972_8799.n176 a_n6972_8799.n49 36.139
R16178 a_n6972_8799.n55 a_n6972_8799.n185 11.843
R16179 a_n6972_8799.n192 a_n6972_8799.n60 36.139
R16180 a_n6972_8799.n66 a_n6972_8799.n202 11.843
R16181 a_n6972_8799.n209 a_n6972_8799.n71 36.139
R16182 a_n6972_8799.n126 a_n6972_8799.n76 11.843
R16183 a_n6972_8799.n130 a_n6972_8799.n81 36.139
R16184 a_n6972_8799.n142 a_n6972_8799.n87 11.843
R16185 a_n6972_8799.n146 a_n6972_8799.n92 36.139
R16186 a_n6972_8799.n159 a_n6972_8799.n98 11.843
R16187 a_n6972_8799.n163 a_n6972_8799.n103 36.139
R16188 a_n6972_8799.n46 a_n6972_8799.n170 35.3134
R16189 a_n6972_8799.n57 a_n6972_8799.n186 35.3134
R16190 a_n6972_8799.n68 a_n6972_8799.n203 35.3134
R16191 a_n6972_8799.n119 a_n6972_8799.n78 35.3134
R16192 a_n6972_8799.n135 a_n6972_8799.n89 35.3134
R16193 a_n6972_8799.n152 a_n6972_8799.n100 35.3134
R16194 a_n6972_8799.n180 a_n6972_8799.n44 34.4824
R16195 a_n6972_8799.n49 a_n6972_8799.n171 10.5784
R16196 a_n6972_8799.n196 a_n6972_8799.n55 34.4824
R16197 a_n6972_8799.n60 a_n6972_8799.n187 10.5784
R16198 a_n6972_8799.n213 a_n6972_8799.n66 34.4824
R16199 a_n6972_8799.n71 a_n6972_8799.n204 10.5784
R16200 a_n6972_8799.n76 a_n6972_8799.n125 34.4824
R16201 a_n6972_8799.n131 a_n6972_8799.n81 10.5784
R16202 a_n6972_8799.n87 a_n6972_8799.n141 34.4824
R16203 a_n6972_8799.n147 a_n6972_8799.n92 10.5784
R16204 a_n6972_8799.n98 a_n6972_8799.n158 34.4824
R16205 a_n6972_8799.n164 a_n6972_8799.n103 10.5784
R16206 a_n6972_8799.n41 a_n6972_8799.n168 36.9592
R16207 a_n6972_8799.n52 a_n6972_8799.n184 36.9592
R16208 a_n6972_8799.n63 a_n6972_8799.n201 36.9592
R16209 a_n6972_8799.n123 a_n6972_8799.n121 21.1793
R16210 a_n6972_8799.n139 a_n6972_8799.n137 21.1793
R16211 a_n6972_8799.n156 a_n6972_8799.n154 21.1793
R16212 a_n6972_8799.n173 a_n6972_8799.n172 20.9576
R16213 a_n6972_8799.n189 a_n6972_8799.n188 20.9576
R16214 a_n6972_8799.n206 a_n6972_8799.n205 20.9576
R16215 a_n6972_8799.n122 a_n6972_8799.n121 20.9576
R16216 a_n6972_8799.n138 a_n6972_8799.n137 20.9576
R16217 a_n6972_8799.n155 a_n6972_8799.n154 20.9576
R16218 a_n6972_8799.n219 a_n6972_8799.n1 12.3339
R16219 a_n6972_8799.n220 a_n6972_8799.n219 11.4887
R16220 a_n6972_8799.n200 a_n6972_8799.n38 9.07815
R16221 a_n6972_8799.n150 a_n6972_8799.n16 9.07815
R16222 a_n6972_8799.n218 a_n6972_8799.n167 6.86264
R16223 a_n6972_8799.n218 a_n6972_8799.n217 6.52017
R16224 a_n6972_8799.n200 a_n6972_8799.n32 4.9702
R16225 a_n6972_8799.n217 a_n6972_8799.n26 4.9702
R16226 a_n6972_8799.n150 a_n6972_8799.n10 4.9702
R16227 a_n6972_8799.n167 a_n6972_8799.n4 4.9702
R16228 a_n6972_8799.n217 a_n6972_8799.n200 4.10845
R16229 a_n6972_8799.n167 a_n6972_8799.n150 4.10845
R16230 a_n6972_8799.n222 a_n6972_8799.t23 3.61217
R16231 a_n6972_8799.n222 a_n6972_8799.t3 3.61217
R16232 a_n6972_8799.n221 a_n6972_8799.t20 3.61217
R16233 a_n6972_8799.n221 a_n6972_8799.t21 3.61217
R16234 a_n6972_8799.n109 a_n6972_8799.t24 3.61217
R16235 a_n6972_8799.n109 a_n6972_8799.t16 3.61217
R16236 a_n6972_8799.n108 a_n6972_8799.t22 3.61217
R16237 a_n6972_8799.n108 a_n6972_8799.t27 3.61217
R16238 a_n6972_8799.n107 a_n6972_8799.t5 3.61217
R16239 a_n6972_8799.n107 a_n6972_8799.t25 3.61217
R16240 a_n6972_8799.t2 a_n6972_8799.n223 3.61217
R16241 a_n6972_8799.n223 a_n6972_8799.t26 3.61217
R16242 a_n6972_8799.n219 a_n6972_8799.n218 3.4105
R16243 a_n6972_8799.n116 a_n6972_8799.t4 2.82907
R16244 a_n6972_8799.n116 a_n6972_8799.t7 2.82907
R16245 a_n6972_8799.n117 a_n6972_8799.t12 2.82907
R16246 a_n6972_8799.n117 a_n6972_8799.t1 2.82907
R16247 a_n6972_8799.n111 a_n6972_8799.t8 2.82907
R16248 a_n6972_8799.n111 a_n6972_8799.t10 2.82907
R16249 a_n6972_8799.n110 a_n6972_8799.t15 2.82907
R16250 a_n6972_8799.n110 a_n6972_8799.t6 2.82907
R16251 a_n6972_8799.n114 a_n6972_8799.t9 2.82907
R16252 a_n6972_8799.n114 a_n6972_8799.t17 2.82907
R16253 a_n6972_8799.n115 a_n6972_8799.t18 2.82907
R16254 a_n6972_8799.n115 a_n6972_8799.t11 2.82907
R16255 a_n6972_8799.n113 a_n6972_8799.t19 2.82907
R16256 a_n6972_8799.n113 a_n6972_8799.t14 2.82907
R16257 a_n6972_8799.n112 a_n6972_8799.t13 2.82907
R16258 a_n6972_8799.n112 a_n6972_8799.t0 2.82907
R16259 a_n6972_8799.n50 a_n6972_8799.n174 47.0982
R16260 a_n6972_8799.n61 a_n6972_8799.n190 47.0982
R16261 a_n6972_8799.n72 a_n6972_8799.n207 47.0982
R16262 a_n6972_8799.n118 a_n6972_8799.n82 47.0982
R16263 a_n6972_8799.n134 a_n6972_8799.n93 47.0982
R16264 a_n6972_8799.n151 a_n6972_8799.n104 47.0982
R16265 a_n6972_8799.n0 a_n6972_8799.n2 33.2634
R16266 a_n6972_8799.n40 a_n6972_8799.n220 31.0217
R16267 a_n6972_8799.n45 a_n6972_8799.n179 0.365327
R16268 a_n6972_8799.n177 a_n6972_8799.n48 21.4216
R16269 a_n6972_8799.n56 a_n6972_8799.n195 0.365327
R16270 a_n6972_8799.n193 a_n6972_8799.n59 21.4216
R16271 a_n6972_8799.n67 a_n6972_8799.n212 0.365327
R16272 a_n6972_8799.n210 a_n6972_8799.n70 21.4216
R16273 a_n6972_8799.n127 a_n6972_8799.n77 0.365327
R16274 a_n6972_8799.n80 a_n6972_8799.n129 21.4216
R16275 a_n6972_8799.n143 a_n6972_8799.n88 0.365327
R16276 a_n6972_8799.n91 a_n6972_8799.n145 21.4216
R16277 a_n6972_8799.n160 a_n6972_8799.n99 0.365327
R16278 a_n6972_8799.n102 a_n6972_8799.n162 21.4216
R16279 a_n6972_8799.n220 a_n6972_8799.n39 18.1434
R16280 a_n6972_8799.n34 a_n6972_8799.n33 1.13686
R16281 a_n6972_8799.n28 a_n6972_8799.n27 1.13686
R16282 a_n6972_8799.n22 a_n6972_8799.n21 1.13686
R16283 a_n6972_8799.n16 a_n6972_8799.n15 1.13686
R16284 a_n6972_8799.n10 a_n6972_8799.n9 1.13686
R16285 a_n6972_8799.n4 a_n6972_8799.n3 1.13686
R16286 a_n6972_8799.n1 a_n6972_8799.n0 1.06084
R16287 a_n6972_8799.n38 a_n6972_8799.n37 0.758076
R16288 a_n6972_8799.n35 a_n6972_8799.n37 0.758076
R16289 a_n6972_8799.n36 a_n6972_8799.n35 0.758076
R16290 a_n6972_8799.n36 a_n6972_8799.n34 0.758076
R16291 a_n6972_8799.n32 a_n6972_8799.n31 0.758076
R16292 a_n6972_8799.n29 a_n6972_8799.n31 0.758076
R16293 a_n6972_8799.n30 a_n6972_8799.n29 0.758076
R16294 a_n6972_8799.n30 a_n6972_8799.n28 0.758076
R16295 a_n6972_8799.n26 a_n6972_8799.n25 0.758076
R16296 a_n6972_8799.n23 a_n6972_8799.n25 0.758076
R16297 a_n6972_8799.n24 a_n6972_8799.n23 0.758076
R16298 a_n6972_8799.n24 a_n6972_8799.n22 0.758076
R16299 a_n6972_8799.n19 a_n6972_8799.n20 0.758076
R16300 a_n6972_8799.n18 a_n6972_8799.n19 0.758076
R16301 a_n6972_8799.n17 a_n6972_8799.n18 0.758076
R16302 a_n6972_8799.n15 a_n6972_8799.n17 0.758076
R16303 a_n6972_8799.n13 a_n6972_8799.n14 0.758076
R16304 a_n6972_8799.n12 a_n6972_8799.n13 0.758076
R16305 a_n6972_8799.n11 a_n6972_8799.n12 0.758076
R16306 a_n6972_8799.n9 a_n6972_8799.n11 0.758076
R16307 a_n6972_8799.n7 a_n6972_8799.n8 0.758076
R16308 a_n6972_8799.n6 a_n6972_8799.n7 0.758076
R16309 a_n6972_8799.n5 a_n6972_8799.n6 0.758076
R16310 a_n6972_8799.n3 a_n6972_8799.n5 0.758076
R16311 vdd.n315 vdd.n279 756.745
R16312 vdd.n260 vdd.n224 756.745
R16313 vdd.n217 vdd.n181 756.745
R16314 vdd.n162 vdd.n126 756.745
R16315 vdd.n120 vdd.n84 756.745
R16316 vdd.n65 vdd.n29 756.745
R16317 vdd.n1684 vdd.n1648 756.745
R16318 vdd.n1739 vdd.n1703 756.745
R16319 vdd.n1586 vdd.n1550 756.745
R16320 vdd.n1641 vdd.n1605 756.745
R16321 vdd.n1489 vdd.n1453 756.745
R16322 vdd.n1544 vdd.n1508 756.745
R16323 vdd.n2094 vdd.t54 640.208
R16324 vdd.n936 vdd.t39 640.208
R16325 vdd.n2068 vdd.t0 640.208
R16326 vdd.n928 vdd.t64 640.208
R16327 vdd.n2839 vdd.t26 640.208
R16328 vdd.n2559 vdd.t61 640.208
R16329 vdd.n804 vdd.t43 640.208
R16330 vdd.n2556 vdd.t47 640.208
R16331 vdd.n768 vdd.t51 640.208
R16332 vdd.n998 vdd.t57 640.208
R16333 vdd.n1148 vdd.t12 592.009
R16334 vdd.n1304 vdd.t23 592.009
R16335 vdd.n1340 vdd.t30 592.009
R16336 vdd.n2250 vdd.t19 592.009
R16337 vdd.n1887 vdd.t33 592.009
R16338 vdd.n1847 vdd.t36 592.009
R16339 vdd.n405 vdd.t8 592.009
R16340 vdd.n419 vdd.t67 592.009
R16341 vdd.n431 vdd.t73 592.009
R16342 vdd.n723 vdd.t4 592.009
R16343 vdd.n686 vdd.t16 592.009
R16344 vdd.n3013 vdd.t70 592.009
R16345 vdd.n316 vdd.n315 585
R16346 vdd.n314 vdd.n281 585
R16347 vdd.n313 vdd.n312 585
R16348 vdd.n284 vdd.n282 585
R16349 vdd.n307 vdd.n306 585
R16350 vdd.n305 vdd.n304 585
R16351 vdd.n288 vdd.n287 585
R16352 vdd.n299 vdd.n298 585
R16353 vdd.n297 vdd.n296 585
R16354 vdd.n292 vdd.n291 585
R16355 vdd.n261 vdd.n260 585
R16356 vdd.n259 vdd.n226 585
R16357 vdd.n258 vdd.n257 585
R16358 vdd.n229 vdd.n227 585
R16359 vdd.n252 vdd.n251 585
R16360 vdd.n250 vdd.n249 585
R16361 vdd.n233 vdd.n232 585
R16362 vdd.n244 vdd.n243 585
R16363 vdd.n242 vdd.n241 585
R16364 vdd.n237 vdd.n236 585
R16365 vdd.n218 vdd.n217 585
R16366 vdd.n216 vdd.n183 585
R16367 vdd.n215 vdd.n214 585
R16368 vdd.n186 vdd.n184 585
R16369 vdd.n209 vdd.n208 585
R16370 vdd.n207 vdd.n206 585
R16371 vdd.n190 vdd.n189 585
R16372 vdd.n201 vdd.n200 585
R16373 vdd.n199 vdd.n198 585
R16374 vdd.n194 vdd.n193 585
R16375 vdd.n163 vdd.n162 585
R16376 vdd.n161 vdd.n128 585
R16377 vdd.n160 vdd.n159 585
R16378 vdd.n131 vdd.n129 585
R16379 vdd.n154 vdd.n153 585
R16380 vdd.n152 vdd.n151 585
R16381 vdd.n135 vdd.n134 585
R16382 vdd.n146 vdd.n145 585
R16383 vdd.n144 vdd.n143 585
R16384 vdd.n139 vdd.n138 585
R16385 vdd.n121 vdd.n120 585
R16386 vdd.n119 vdd.n86 585
R16387 vdd.n118 vdd.n117 585
R16388 vdd.n89 vdd.n87 585
R16389 vdd.n112 vdd.n111 585
R16390 vdd.n110 vdd.n109 585
R16391 vdd.n93 vdd.n92 585
R16392 vdd.n104 vdd.n103 585
R16393 vdd.n102 vdd.n101 585
R16394 vdd.n97 vdd.n96 585
R16395 vdd.n66 vdd.n65 585
R16396 vdd.n64 vdd.n31 585
R16397 vdd.n63 vdd.n62 585
R16398 vdd.n34 vdd.n32 585
R16399 vdd.n57 vdd.n56 585
R16400 vdd.n55 vdd.n54 585
R16401 vdd.n38 vdd.n37 585
R16402 vdd.n49 vdd.n48 585
R16403 vdd.n47 vdd.n46 585
R16404 vdd.n42 vdd.n41 585
R16405 vdd.n1685 vdd.n1684 585
R16406 vdd.n1683 vdd.n1650 585
R16407 vdd.n1682 vdd.n1681 585
R16408 vdd.n1653 vdd.n1651 585
R16409 vdd.n1676 vdd.n1675 585
R16410 vdd.n1674 vdd.n1673 585
R16411 vdd.n1657 vdd.n1656 585
R16412 vdd.n1668 vdd.n1667 585
R16413 vdd.n1666 vdd.n1665 585
R16414 vdd.n1661 vdd.n1660 585
R16415 vdd.n1740 vdd.n1739 585
R16416 vdd.n1738 vdd.n1705 585
R16417 vdd.n1737 vdd.n1736 585
R16418 vdd.n1708 vdd.n1706 585
R16419 vdd.n1731 vdd.n1730 585
R16420 vdd.n1729 vdd.n1728 585
R16421 vdd.n1712 vdd.n1711 585
R16422 vdd.n1723 vdd.n1722 585
R16423 vdd.n1721 vdd.n1720 585
R16424 vdd.n1716 vdd.n1715 585
R16425 vdd.n1587 vdd.n1586 585
R16426 vdd.n1585 vdd.n1552 585
R16427 vdd.n1584 vdd.n1583 585
R16428 vdd.n1555 vdd.n1553 585
R16429 vdd.n1578 vdd.n1577 585
R16430 vdd.n1576 vdd.n1575 585
R16431 vdd.n1559 vdd.n1558 585
R16432 vdd.n1570 vdd.n1569 585
R16433 vdd.n1568 vdd.n1567 585
R16434 vdd.n1563 vdd.n1562 585
R16435 vdd.n1642 vdd.n1641 585
R16436 vdd.n1640 vdd.n1607 585
R16437 vdd.n1639 vdd.n1638 585
R16438 vdd.n1610 vdd.n1608 585
R16439 vdd.n1633 vdd.n1632 585
R16440 vdd.n1631 vdd.n1630 585
R16441 vdd.n1614 vdd.n1613 585
R16442 vdd.n1625 vdd.n1624 585
R16443 vdd.n1623 vdd.n1622 585
R16444 vdd.n1618 vdd.n1617 585
R16445 vdd.n1490 vdd.n1489 585
R16446 vdd.n1488 vdd.n1455 585
R16447 vdd.n1487 vdd.n1486 585
R16448 vdd.n1458 vdd.n1456 585
R16449 vdd.n1481 vdd.n1480 585
R16450 vdd.n1479 vdd.n1478 585
R16451 vdd.n1462 vdd.n1461 585
R16452 vdd.n1473 vdd.n1472 585
R16453 vdd.n1471 vdd.n1470 585
R16454 vdd.n1466 vdd.n1465 585
R16455 vdd.n1545 vdd.n1544 585
R16456 vdd.n1543 vdd.n1510 585
R16457 vdd.n1542 vdd.n1541 585
R16458 vdd.n1513 vdd.n1511 585
R16459 vdd.n1536 vdd.n1535 585
R16460 vdd.n1534 vdd.n1533 585
R16461 vdd.n1517 vdd.n1516 585
R16462 vdd.n1528 vdd.n1527 585
R16463 vdd.n1526 vdd.n1525 585
R16464 vdd.n1521 vdd.n1520 585
R16465 vdd.n445 vdd.n370 462.44
R16466 vdd.n3251 vdd.n372 462.44
R16467 vdd.n3146 vdd.n657 462.44
R16468 vdd.n3144 vdd.n660 462.44
R16469 vdd.n2245 vdd.n1047 462.44
R16470 vdd.n2248 vdd.n2247 462.44
R16471 vdd.n1375 vdd.n1145 462.44
R16472 vdd.n1372 vdd.n1143 462.44
R16473 vdd.n293 vdd.t214 329.043
R16474 vdd.n238 vdd.t190 329.043
R16475 vdd.n195 vdd.t202 329.043
R16476 vdd.n140 vdd.t179 329.043
R16477 vdd.n98 vdd.t136 329.043
R16478 vdd.n43 vdd.t113 329.043
R16479 vdd.n1662 vdd.t228 329.043
R16480 vdd.n1717 vdd.t140 329.043
R16481 vdd.n1564 vdd.t215 329.043
R16482 vdd.n1619 vdd.t123 329.043
R16483 vdd.n1467 vdd.t115 329.043
R16484 vdd.n1522 vdd.t137 329.043
R16485 vdd.n1148 vdd.t15 319.788
R16486 vdd.n1304 vdd.t25 319.788
R16487 vdd.n1340 vdd.t32 319.788
R16488 vdd.n2250 vdd.t21 319.788
R16489 vdd.n1887 vdd.t34 319.788
R16490 vdd.n1847 vdd.t37 319.788
R16491 vdd.n405 vdd.t10 319.788
R16492 vdd.n419 vdd.t68 319.788
R16493 vdd.n431 vdd.t74 319.788
R16494 vdd.n723 vdd.t7 319.788
R16495 vdd.n686 vdd.t18 319.788
R16496 vdd.n3013 vdd.t72 319.788
R16497 vdd.n1149 vdd.t14 303.69
R16498 vdd.n1305 vdd.t24 303.69
R16499 vdd.n1341 vdd.t31 303.69
R16500 vdd.n2251 vdd.t22 303.69
R16501 vdd.n1888 vdd.t35 303.69
R16502 vdd.n1848 vdd.t38 303.69
R16503 vdd.n406 vdd.t11 303.69
R16504 vdd.n420 vdd.t69 303.69
R16505 vdd.n432 vdd.t75 303.69
R16506 vdd.n724 vdd.t6 303.69
R16507 vdd.n687 vdd.t17 303.69
R16508 vdd.n3014 vdd.t71 303.69
R16509 vdd.n2782 vdd.n884 297.074
R16510 vdd.n2975 vdd.n778 297.074
R16511 vdd.n2912 vdd.n775 297.074
R16512 vdd.n2705 vdd.n885 297.074
R16513 vdd.n2520 vdd.n925 297.074
R16514 vdd.n2451 vdd.n2450 297.074
R16515 vdd.n2197 vdd.n1021 297.074
R16516 vdd.n2293 vdd.n1019 297.074
R16517 vdd.n2891 vdd.n776 297.074
R16518 vdd.n2978 vdd.n2977 297.074
R16519 vdd.n2554 vdd.n886 297.074
R16520 vdd.n2780 vdd.n887 297.074
R16521 vdd.n2448 vdd.n934 297.074
R16522 vdd.n932 vdd.n907 297.074
R16523 vdd.n2134 vdd.n1022 297.074
R16524 vdd.n2291 vdd.n1023 297.074
R16525 vdd.n2893 vdd.n776 185
R16526 vdd.n2976 vdd.n776 185
R16527 vdd.n2895 vdd.n2894 185
R16528 vdd.n2894 vdd.n774 185
R16529 vdd.n2896 vdd.n810 185
R16530 vdd.n2906 vdd.n810 185
R16531 vdd.n2897 vdd.n819 185
R16532 vdd.n819 vdd.n817 185
R16533 vdd.n2899 vdd.n2898 185
R16534 vdd.n2900 vdd.n2899 185
R16535 vdd.n2852 vdd.n818 185
R16536 vdd.n818 vdd.n814 185
R16537 vdd.n2851 vdd.n2850 185
R16538 vdd.n2850 vdd.n2849 185
R16539 vdd.n821 vdd.n820 185
R16540 vdd.n822 vdd.n821 185
R16541 vdd.n2842 vdd.n2841 185
R16542 vdd.n2843 vdd.n2842 185
R16543 vdd.n2838 vdd.n831 185
R16544 vdd.n831 vdd.n828 185
R16545 vdd.n2837 vdd.n2836 185
R16546 vdd.n2836 vdd.n2835 185
R16547 vdd.n833 vdd.n832 185
R16548 vdd.n841 vdd.n833 185
R16549 vdd.n2828 vdd.n2827 185
R16550 vdd.n2829 vdd.n2828 185
R16551 vdd.n2826 vdd.n842 185
R16552 vdd.n2677 vdd.n842 185
R16553 vdd.n2825 vdd.n2824 185
R16554 vdd.n2824 vdd.n2823 185
R16555 vdd.n844 vdd.n843 185
R16556 vdd.n845 vdd.n844 185
R16557 vdd.n2816 vdd.n2815 185
R16558 vdd.n2817 vdd.n2816 185
R16559 vdd.n2814 vdd.n854 185
R16560 vdd.n854 vdd.n851 185
R16561 vdd.n2813 vdd.n2812 185
R16562 vdd.n2812 vdd.n2811 185
R16563 vdd.n856 vdd.n855 185
R16564 vdd.n864 vdd.n856 185
R16565 vdd.n2804 vdd.n2803 185
R16566 vdd.n2805 vdd.n2804 185
R16567 vdd.n2802 vdd.n865 185
R16568 vdd.n871 vdd.n865 185
R16569 vdd.n2801 vdd.n2800 185
R16570 vdd.n2800 vdd.n2799 185
R16571 vdd.n867 vdd.n866 185
R16572 vdd.n868 vdd.n867 185
R16573 vdd.n2792 vdd.n2791 185
R16574 vdd.n2793 vdd.n2792 185
R16575 vdd.n2790 vdd.n877 185
R16576 vdd.n2698 vdd.n877 185
R16577 vdd.n2789 vdd.n2788 185
R16578 vdd.n2788 vdd.n2787 185
R16579 vdd.n879 vdd.n878 185
R16580 vdd.t248 vdd.n879 185
R16581 vdd.n2780 vdd.n2779 185
R16582 vdd.n2781 vdd.n2780 185
R16583 vdd.n2778 vdd.n887 185
R16584 vdd.n2777 vdd.n2776 185
R16585 vdd.n889 vdd.n888 185
R16586 vdd.n2563 vdd.n2562 185
R16587 vdd.n2565 vdd.n2564 185
R16588 vdd.n2567 vdd.n2566 185
R16589 vdd.n2569 vdd.n2568 185
R16590 vdd.n2571 vdd.n2570 185
R16591 vdd.n2573 vdd.n2572 185
R16592 vdd.n2575 vdd.n2574 185
R16593 vdd.n2577 vdd.n2576 185
R16594 vdd.n2579 vdd.n2578 185
R16595 vdd.n2581 vdd.n2580 185
R16596 vdd.n2583 vdd.n2582 185
R16597 vdd.n2585 vdd.n2584 185
R16598 vdd.n2587 vdd.n2586 185
R16599 vdd.n2589 vdd.n2588 185
R16600 vdd.n2591 vdd.n2590 185
R16601 vdd.n2593 vdd.n2592 185
R16602 vdd.n2595 vdd.n2594 185
R16603 vdd.n2597 vdd.n2596 185
R16604 vdd.n2599 vdd.n2598 185
R16605 vdd.n2601 vdd.n2600 185
R16606 vdd.n2603 vdd.n2602 185
R16607 vdd.n2605 vdd.n2604 185
R16608 vdd.n2607 vdd.n2606 185
R16609 vdd.n2609 vdd.n2608 185
R16610 vdd.n2611 vdd.n2610 185
R16611 vdd.n2613 vdd.n2612 185
R16612 vdd.n2615 vdd.n2614 185
R16613 vdd.n2617 vdd.n2616 185
R16614 vdd.n2619 vdd.n2618 185
R16615 vdd.n2621 vdd.n2620 185
R16616 vdd.n2623 vdd.n2622 185
R16617 vdd.n2624 vdd.n2554 185
R16618 vdd.n2774 vdd.n2554 185
R16619 vdd.n2979 vdd.n2978 185
R16620 vdd.n2980 vdd.n767 185
R16621 vdd.n2982 vdd.n2981 185
R16622 vdd.n2984 vdd.n765 185
R16623 vdd.n2986 vdd.n2985 185
R16624 vdd.n2987 vdd.n764 185
R16625 vdd.n2989 vdd.n2988 185
R16626 vdd.n2991 vdd.n762 185
R16627 vdd.n2993 vdd.n2992 185
R16628 vdd.n2994 vdd.n761 185
R16629 vdd.n2996 vdd.n2995 185
R16630 vdd.n2998 vdd.n759 185
R16631 vdd.n3000 vdd.n2999 185
R16632 vdd.n3001 vdd.n758 185
R16633 vdd.n3003 vdd.n3002 185
R16634 vdd.n3005 vdd.n757 185
R16635 vdd.n3006 vdd.n754 185
R16636 vdd.n3009 vdd.n3008 185
R16637 vdd.n755 vdd.n753 185
R16638 vdd.n2865 vdd.n2864 185
R16639 vdd.n2867 vdd.n2866 185
R16640 vdd.n2869 vdd.n2861 185
R16641 vdd.n2871 vdd.n2870 185
R16642 vdd.n2872 vdd.n2860 185
R16643 vdd.n2874 vdd.n2873 185
R16644 vdd.n2876 vdd.n2858 185
R16645 vdd.n2878 vdd.n2877 185
R16646 vdd.n2879 vdd.n2857 185
R16647 vdd.n2881 vdd.n2880 185
R16648 vdd.n2883 vdd.n2855 185
R16649 vdd.n2885 vdd.n2884 185
R16650 vdd.n2886 vdd.n2854 185
R16651 vdd.n2888 vdd.n2887 185
R16652 vdd.n2890 vdd.n2853 185
R16653 vdd.n2892 vdd.n2891 185
R16654 vdd.n2891 vdd.n756 185
R16655 vdd.n2977 vdd.n771 185
R16656 vdd.n2977 vdd.n2976 185
R16657 vdd.n2629 vdd.n773 185
R16658 vdd.n774 vdd.n773 185
R16659 vdd.n2630 vdd.n809 185
R16660 vdd.n2906 vdd.n809 185
R16661 vdd.n2632 vdd.n2631 185
R16662 vdd.n2631 vdd.n817 185
R16663 vdd.n2633 vdd.n816 185
R16664 vdd.n2900 vdd.n816 185
R16665 vdd.n2635 vdd.n2634 185
R16666 vdd.n2634 vdd.n814 185
R16667 vdd.n2636 vdd.n824 185
R16668 vdd.n2849 vdd.n824 185
R16669 vdd.n2638 vdd.n2637 185
R16670 vdd.n2637 vdd.n822 185
R16671 vdd.n2639 vdd.n830 185
R16672 vdd.n2843 vdd.n830 185
R16673 vdd.n2641 vdd.n2640 185
R16674 vdd.n2640 vdd.n828 185
R16675 vdd.n2642 vdd.n835 185
R16676 vdd.n2835 vdd.n835 185
R16677 vdd.n2644 vdd.n2643 185
R16678 vdd.n2643 vdd.n841 185
R16679 vdd.n2645 vdd.n840 185
R16680 vdd.n2829 vdd.n840 185
R16681 vdd.n2679 vdd.n2678 185
R16682 vdd.n2678 vdd.n2677 185
R16683 vdd.n2680 vdd.n847 185
R16684 vdd.n2823 vdd.n847 185
R16685 vdd.n2682 vdd.n2681 185
R16686 vdd.n2681 vdd.n845 185
R16687 vdd.n2683 vdd.n853 185
R16688 vdd.n2817 vdd.n853 185
R16689 vdd.n2685 vdd.n2684 185
R16690 vdd.n2684 vdd.n851 185
R16691 vdd.n2686 vdd.n858 185
R16692 vdd.n2811 vdd.n858 185
R16693 vdd.n2688 vdd.n2687 185
R16694 vdd.n2687 vdd.n864 185
R16695 vdd.n2689 vdd.n863 185
R16696 vdd.n2805 vdd.n863 185
R16697 vdd.n2691 vdd.n2690 185
R16698 vdd.n2690 vdd.n871 185
R16699 vdd.n2692 vdd.n870 185
R16700 vdd.n2799 vdd.n870 185
R16701 vdd.n2694 vdd.n2693 185
R16702 vdd.n2693 vdd.n868 185
R16703 vdd.n2695 vdd.n876 185
R16704 vdd.n2793 vdd.n876 185
R16705 vdd.n2697 vdd.n2696 185
R16706 vdd.n2698 vdd.n2697 185
R16707 vdd.n2628 vdd.n881 185
R16708 vdd.n2787 vdd.n881 185
R16709 vdd.n2627 vdd.n2626 185
R16710 vdd.n2626 vdd.t248 185
R16711 vdd.n2625 vdd.n886 185
R16712 vdd.n2781 vdd.n886 185
R16713 vdd.n2245 vdd.n2244 185
R16714 vdd.n2246 vdd.n2245 185
R16715 vdd.n1048 vdd.n1046 185
R16716 vdd.n1046 vdd.n1044 185
R16717 vdd.n1814 vdd.n1813 185
R16718 vdd.n1813 vdd.n1812 185
R16719 vdd.n1051 vdd.n1050 185
R16720 vdd.n1052 vdd.n1051 185
R16721 vdd.n1801 vdd.n1800 185
R16722 vdd.n1802 vdd.n1801 185
R16723 vdd.n1060 vdd.n1059 185
R16724 vdd.n1793 vdd.n1059 185
R16725 vdd.n1796 vdd.n1795 185
R16726 vdd.n1795 vdd.n1794 185
R16727 vdd.n1063 vdd.n1062 185
R16728 vdd.n1069 vdd.n1063 185
R16729 vdd.n1784 vdd.n1783 185
R16730 vdd.n1785 vdd.n1784 185
R16731 vdd.n1071 vdd.n1070 185
R16732 vdd.n1776 vdd.n1070 185
R16733 vdd.n1779 vdd.n1778 185
R16734 vdd.n1778 vdd.n1777 185
R16735 vdd.n1074 vdd.n1073 185
R16736 vdd.n1075 vdd.n1074 185
R16737 vdd.n1767 vdd.n1766 185
R16738 vdd.n1768 vdd.n1767 185
R16739 vdd.n1083 vdd.n1082 185
R16740 vdd.n1082 vdd.n1081 185
R16741 vdd.n1762 vdd.n1761 185
R16742 vdd.n1761 vdd.n1760 185
R16743 vdd.n1086 vdd.n1085 185
R16744 vdd.n1092 vdd.n1086 185
R16745 vdd.n1751 vdd.n1750 185
R16746 vdd.n1752 vdd.n1751 185
R16747 vdd.n1094 vdd.n1093 185
R16748 vdd.n1448 vdd.n1093 185
R16749 vdd.n1451 vdd.n1450 185
R16750 vdd.n1450 vdd.n1449 185
R16751 vdd.n1097 vdd.n1096 185
R16752 vdd.n1104 vdd.n1097 185
R16753 vdd.n1439 vdd.n1438 185
R16754 vdd.n1440 vdd.n1439 185
R16755 vdd.n1106 vdd.n1105 185
R16756 vdd.n1105 vdd.n1103 185
R16757 vdd.n1434 vdd.n1433 185
R16758 vdd.n1433 vdd.n1432 185
R16759 vdd.n1109 vdd.n1108 185
R16760 vdd.n1110 vdd.n1109 185
R16761 vdd.n1423 vdd.n1422 185
R16762 vdd.n1424 vdd.n1423 185
R16763 vdd.n1117 vdd.n1116 185
R16764 vdd.n1415 vdd.n1116 185
R16765 vdd.n1418 vdd.n1417 185
R16766 vdd.n1417 vdd.n1416 185
R16767 vdd.n1120 vdd.n1119 185
R16768 vdd.n1126 vdd.n1120 185
R16769 vdd.n1406 vdd.n1405 185
R16770 vdd.n1407 vdd.n1406 185
R16771 vdd.n1128 vdd.n1127 185
R16772 vdd.n1398 vdd.n1127 185
R16773 vdd.n1401 vdd.n1400 185
R16774 vdd.n1400 vdd.n1399 185
R16775 vdd.n1131 vdd.n1130 185
R16776 vdd.n1132 vdd.n1131 185
R16777 vdd.n1389 vdd.n1388 185
R16778 vdd.n1390 vdd.n1389 185
R16779 vdd.n1140 vdd.n1139 185
R16780 vdd.n1139 vdd.n1138 185
R16781 vdd.n1384 vdd.n1383 185
R16782 vdd.n1383 vdd.n1382 185
R16783 vdd.n1143 vdd.n1142 185
R16784 vdd.n1144 vdd.n1143 185
R16785 vdd.n1372 vdd.n1371 185
R16786 vdd.n1370 vdd.n1183 185
R16787 vdd.n1185 vdd.n1182 185
R16788 vdd.n1374 vdd.n1182 185
R16789 vdd.n1366 vdd.n1187 185
R16790 vdd.n1365 vdd.n1188 185
R16791 vdd.n1364 vdd.n1189 185
R16792 vdd.n1192 vdd.n1190 185
R16793 vdd.n1360 vdd.n1193 185
R16794 vdd.n1359 vdd.n1194 185
R16795 vdd.n1358 vdd.n1195 185
R16796 vdd.n1198 vdd.n1196 185
R16797 vdd.n1354 vdd.n1199 185
R16798 vdd.n1353 vdd.n1200 185
R16799 vdd.n1352 vdd.n1201 185
R16800 vdd.n1204 vdd.n1202 185
R16801 vdd.n1348 vdd.n1205 185
R16802 vdd.n1347 vdd.n1206 185
R16803 vdd.n1346 vdd.n1207 185
R16804 vdd.n1338 vdd.n1208 185
R16805 vdd.n1342 vdd.n1339 185
R16806 vdd.n1337 vdd.n1210 185
R16807 vdd.n1336 vdd.n1211 185
R16808 vdd.n1214 vdd.n1212 185
R16809 vdd.n1332 vdd.n1215 185
R16810 vdd.n1331 vdd.n1216 185
R16811 vdd.n1330 vdd.n1217 185
R16812 vdd.n1220 vdd.n1218 185
R16813 vdd.n1326 vdd.n1221 185
R16814 vdd.n1325 vdd.n1222 185
R16815 vdd.n1324 vdd.n1223 185
R16816 vdd.n1226 vdd.n1224 185
R16817 vdd.n1320 vdd.n1227 185
R16818 vdd.n1319 vdd.n1228 185
R16819 vdd.n1318 vdd.n1229 185
R16820 vdd.n1232 vdd.n1230 185
R16821 vdd.n1314 vdd.n1233 185
R16822 vdd.n1313 vdd.n1234 185
R16823 vdd.n1312 vdd.n1235 185
R16824 vdd.n1238 vdd.n1236 185
R16825 vdd.n1308 vdd.n1239 185
R16826 vdd.n1307 vdd.n1240 185
R16827 vdd.n1306 vdd.n1303 185
R16828 vdd.n1243 vdd.n1241 185
R16829 vdd.n1299 vdd.n1244 185
R16830 vdd.n1298 vdd.n1245 185
R16831 vdd.n1297 vdd.n1246 185
R16832 vdd.n1249 vdd.n1247 185
R16833 vdd.n1293 vdd.n1250 185
R16834 vdd.n1292 vdd.n1251 185
R16835 vdd.n1291 vdd.n1252 185
R16836 vdd.n1255 vdd.n1253 185
R16837 vdd.n1287 vdd.n1256 185
R16838 vdd.n1286 vdd.n1257 185
R16839 vdd.n1285 vdd.n1258 185
R16840 vdd.n1261 vdd.n1259 185
R16841 vdd.n1281 vdd.n1262 185
R16842 vdd.n1280 vdd.n1263 185
R16843 vdd.n1279 vdd.n1264 185
R16844 vdd.n1267 vdd.n1265 185
R16845 vdd.n1275 vdd.n1268 185
R16846 vdd.n1274 vdd.n1269 185
R16847 vdd.n1273 vdd.n1270 185
R16848 vdd.n1271 vdd.n1151 185
R16849 vdd.n1376 vdd.n1375 185
R16850 vdd.n1375 vdd.n1374 185
R16851 vdd.n2249 vdd.n2248 185
R16852 vdd.n2253 vdd.n1040 185
R16853 vdd.n1916 vdd.n1039 185
R16854 vdd.n1919 vdd.n1918 185
R16855 vdd.n1921 vdd.n1920 185
R16856 vdd.n1924 vdd.n1923 185
R16857 vdd.n1926 vdd.n1925 185
R16858 vdd.n1928 vdd.n1914 185
R16859 vdd.n1930 vdd.n1929 185
R16860 vdd.n1931 vdd.n1908 185
R16861 vdd.n1933 vdd.n1932 185
R16862 vdd.n1935 vdd.n1906 185
R16863 vdd.n1937 vdd.n1936 185
R16864 vdd.n1938 vdd.n1901 185
R16865 vdd.n1940 vdd.n1939 185
R16866 vdd.n1942 vdd.n1899 185
R16867 vdd.n1944 vdd.n1943 185
R16868 vdd.n1945 vdd.n1895 185
R16869 vdd.n1947 vdd.n1946 185
R16870 vdd.n1949 vdd.n1892 185
R16871 vdd.n1951 vdd.n1950 185
R16872 vdd.n1893 vdd.n1886 185
R16873 vdd.n1955 vdd.n1890 185
R16874 vdd.n1956 vdd.n1882 185
R16875 vdd.n1958 vdd.n1957 185
R16876 vdd.n1960 vdd.n1880 185
R16877 vdd.n1962 vdd.n1961 185
R16878 vdd.n1963 vdd.n1875 185
R16879 vdd.n1965 vdd.n1964 185
R16880 vdd.n1967 vdd.n1873 185
R16881 vdd.n1969 vdd.n1968 185
R16882 vdd.n1970 vdd.n1868 185
R16883 vdd.n1972 vdd.n1971 185
R16884 vdd.n1974 vdd.n1866 185
R16885 vdd.n1976 vdd.n1975 185
R16886 vdd.n1977 vdd.n1861 185
R16887 vdd.n1979 vdd.n1978 185
R16888 vdd.n1981 vdd.n1859 185
R16889 vdd.n1983 vdd.n1982 185
R16890 vdd.n1984 vdd.n1855 185
R16891 vdd.n1986 vdd.n1985 185
R16892 vdd.n1988 vdd.n1852 185
R16893 vdd.n1990 vdd.n1989 185
R16894 vdd.n1853 vdd.n1846 185
R16895 vdd.n1994 vdd.n1850 185
R16896 vdd.n1995 vdd.n1842 185
R16897 vdd.n1997 vdd.n1996 185
R16898 vdd.n1999 vdd.n1840 185
R16899 vdd.n2001 vdd.n2000 185
R16900 vdd.n2002 vdd.n1835 185
R16901 vdd.n2004 vdd.n2003 185
R16902 vdd.n2006 vdd.n1833 185
R16903 vdd.n2008 vdd.n2007 185
R16904 vdd.n2009 vdd.n1828 185
R16905 vdd.n2011 vdd.n2010 185
R16906 vdd.n2013 vdd.n1827 185
R16907 vdd.n2014 vdd.n1824 185
R16908 vdd.n2017 vdd.n2016 185
R16909 vdd.n1826 vdd.n1822 185
R16910 vdd.n2234 vdd.n1820 185
R16911 vdd.n2236 vdd.n2235 185
R16912 vdd.n2238 vdd.n1818 185
R16913 vdd.n2240 vdd.n2239 185
R16914 vdd.n2241 vdd.n1047 185
R16915 vdd.n2247 vdd.n1043 185
R16916 vdd.n2247 vdd.n2246 185
R16917 vdd.n1055 vdd.n1042 185
R16918 vdd.n1044 vdd.n1042 185
R16919 vdd.n1811 vdd.n1810 185
R16920 vdd.n1812 vdd.n1811 185
R16921 vdd.n1054 vdd.n1053 185
R16922 vdd.n1053 vdd.n1052 185
R16923 vdd.n1804 vdd.n1803 185
R16924 vdd.n1803 vdd.n1802 185
R16925 vdd.n1058 vdd.n1057 185
R16926 vdd.n1793 vdd.n1058 185
R16927 vdd.n1792 vdd.n1791 185
R16928 vdd.n1794 vdd.n1792 185
R16929 vdd.n1065 vdd.n1064 185
R16930 vdd.n1069 vdd.n1064 185
R16931 vdd.n1787 vdd.n1786 185
R16932 vdd.n1786 vdd.n1785 185
R16933 vdd.n1068 vdd.n1067 185
R16934 vdd.n1776 vdd.n1068 185
R16935 vdd.n1775 vdd.n1774 185
R16936 vdd.n1777 vdd.n1775 185
R16937 vdd.n1077 vdd.n1076 185
R16938 vdd.n1076 vdd.n1075 185
R16939 vdd.n1770 vdd.n1769 185
R16940 vdd.n1769 vdd.n1768 185
R16941 vdd.n1080 vdd.n1079 185
R16942 vdd.n1081 vdd.n1080 185
R16943 vdd.n1759 vdd.n1758 185
R16944 vdd.n1760 vdd.n1759 185
R16945 vdd.n1088 vdd.n1087 185
R16946 vdd.n1092 vdd.n1087 185
R16947 vdd.n1754 vdd.n1753 185
R16948 vdd.n1753 vdd.n1752 185
R16949 vdd.n1091 vdd.n1090 185
R16950 vdd.n1448 vdd.n1091 185
R16951 vdd.n1447 vdd.n1446 185
R16952 vdd.n1449 vdd.n1447 185
R16953 vdd.n1099 vdd.n1098 185
R16954 vdd.n1104 vdd.n1098 185
R16955 vdd.n1442 vdd.n1441 185
R16956 vdd.n1441 vdd.n1440 185
R16957 vdd.n1102 vdd.n1101 185
R16958 vdd.n1103 vdd.n1102 185
R16959 vdd.n1431 vdd.n1430 185
R16960 vdd.n1432 vdd.n1431 185
R16961 vdd.n1112 vdd.n1111 185
R16962 vdd.n1111 vdd.n1110 185
R16963 vdd.n1426 vdd.n1425 185
R16964 vdd.n1425 vdd.n1424 185
R16965 vdd.n1115 vdd.n1114 185
R16966 vdd.n1415 vdd.n1115 185
R16967 vdd.n1414 vdd.n1413 185
R16968 vdd.n1416 vdd.n1414 185
R16969 vdd.n1122 vdd.n1121 185
R16970 vdd.n1126 vdd.n1121 185
R16971 vdd.n1409 vdd.n1408 185
R16972 vdd.n1408 vdd.n1407 185
R16973 vdd.n1125 vdd.n1124 185
R16974 vdd.n1398 vdd.n1125 185
R16975 vdd.n1397 vdd.n1396 185
R16976 vdd.n1399 vdd.n1397 185
R16977 vdd.n1134 vdd.n1133 185
R16978 vdd.n1133 vdd.n1132 185
R16979 vdd.n1392 vdd.n1391 185
R16980 vdd.n1391 vdd.n1390 185
R16981 vdd.n1137 vdd.n1136 185
R16982 vdd.n1138 vdd.n1137 185
R16983 vdd.n1381 vdd.n1380 185
R16984 vdd.n1382 vdd.n1381 185
R16985 vdd.n1146 vdd.n1145 185
R16986 vdd.n1145 vdd.n1144 185
R16987 vdd.n927 vdd.n925 185
R16988 vdd.n2449 vdd.n925 185
R16989 vdd.n2371 vdd.n944 185
R16990 vdd.n944 vdd.t262 185
R16991 vdd.n2373 vdd.n2372 185
R16992 vdd.n2374 vdd.n2373 185
R16993 vdd.n2370 vdd.n943 185
R16994 vdd.n2073 vdd.n943 185
R16995 vdd.n2369 vdd.n2368 185
R16996 vdd.n2368 vdd.n2367 185
R16997 vdd.n946 vdd.n945 185
R16998 vdd.n947 vdd.n946 185
R16999 vdd.n2358 vdd.n2357 185
R17000 vdd.n2359 vdd.n2358 185
R17001 vdd.n2356 vdd.n957 185
R17002 vdd.n957 vdd.n954 185
R17003 vdd.n2355 vdd.n2354 185
R17004 vdd.n2354 vdd.n2353 185
R17005 vdd.n959 vdd.n958 185
R17006 vdd.n960 vdd.n959 185
R17007 vdd.n2346 vdd.n2345 185
R17008 vdd.n2347 vdd.n2346 185
R17009 vdd.n2344 vdd.n968 185
R17010 vdd.n973 vdd.n968 185
R17011 vdd.n2343 vdd.n2342 185
R17012 vdd.n2342 vdd.n2341 185
R17013 vdd.n970 vdd.n969 185
R17014 vdd.n979 vdd.n970 185
R17015 vdd.n2334 vdd.n2333 185
R17016 vdd.n2335 vdd.n2334 185
R17017 vdd.n2332 vdd.n980 185
R17018 vdd.n2174 vdd.n980 185
R17019 vdd.n2331 vdd.n2330 185
R17020 vdd.n2330 vdd.n2329 185
R17021 vdd.n982 vdd.n981 185
R17022 vdd.n983 vdd.n982 185
R17023 vdd.n2322 vdd.n2321 185
R17024 vdd.n2323 vdd.n2322 185
R17025 vdd.n2320 vdd.n992 185
R17026 vdd.n992 vdd.n989 185
R17027 vdd.n2319 vdd.n2318 185
R17028 vdd.n2318 vdd.n2317 185
R17029 vdd.n994 vdd.n993 185
R17030 vdd.n1004 vdd.n994 185
R17031 vdd.n2309 vdd.n2308 185
R17032 vdd.n2310 vdd.n2309 185
R17033 vdd.n2307 vdd.n1005 185
R17034 vdd.n1005 vdd.n1001 185
R17035 vdd.n2306 vdd.n2305 185
R17036 vdd.n2305 vdd.n2304 185
R17037 vdd.n1007 vdd.n1006 185
R17038 vdd.n1008 vdd.n1007 185
R17039 vdd.n2297 vdd.n2296 185
R17040 vdd.n2298 vdd.n2297 185
R17041 vdd.n2295 vdd.n1017 185
R17042 vdd.n1017 vdd.n1014 185
R17043 vdd.n2294 vdd.n2293 185
R17044 vdd.n2293 vdd.n2292 185
R17045 vdd.n1019 vdd.n1018 185
R17046 vdd.n2029 vdd.n2028 185
R17047 vdd.n2030 vdd.n2026 185
R17048 vdd.n2026 vdd.n1020 185
R17049 vdd.n2032 vdd.n2031 185
R17050 vdd.n2034 vdd.n2025 185
R17051 vdd.n2037 vdd.n2036 185
R17052 vdd.n2038 vdd.n2024 185
R17053 vdd.n2040 vdd.n2039 185
R17054 vdd.n2042 vdd.n2023 185
R17055 vdd.n2045 vdd.n2044 185
R17056 vdd.n2046 vdd.n2022 185
R17057 vdd.n2048 vdd.n2047 185
R17058 vdd.n2050 vdd.n2021 185
R17059 vdd.n2053 vdd.n2052 185
R17060 vdd.n2054 vdd.n2020 185
R17061 vdd.n2056 vdd.n2055 185
R17062 vdd.n2058 vdd.n2019 185
R17063 vdd.n2231 vdd.n2059 185
R17064 vdd.n2230 vdd.n2229 185
R17065 vdd.n2227 vdd.n2060 185
R17066 vdd.n2225 vdd.n2224 185
R17067 vdd.n2223 vdd.n2061 185
R17068 vdd.n2222 vdd.n2221 185
R17069 vdd.n2219 vdd.n2062 185
R17070 vdd.n2217 vdd.n2216 185
R17071 vdd.n2215 vdd.n2063 185
R17072 vdd.n2214 vdd.n2213 185
R17073 vdd.n2211 vdd.n2064 185
R17074 vdd.n2209 vdd.n2208 185
R17075 vdd.n2207 vdd.n2065 185
R17076 vdd.n2206 vdd.n2205 185
R17077 vdd.n2203 vdd.n2066 185
R17078 vdd.n2201 vdd.n2200 185
R17079 vdd.n2199 vdd.n2067 185
R17080 vdd.n2198 vdd.n2197 185
R17081 vdd.n2452 vdd.n2451 185
R17082 vdd.n2454 vdd.n2453 185
R17083 vdd.n2456 vdd.n2455 185
R17084 vdd.n2459 vdd.n2458 185
R17085 vdd.n2461 vdd.n2460 185
R17086 vdd.n2463 vdd.n2462 185
R17087 vdd.n2465 vdd.n2464 185
R17088 vdd.n2467 vdd.n2466 185
R17089 vdd.n2469 vdd.n2468 185
R17090 vdd.n2471 vdd.n2470 185
R17091 vdd.n2473 vdd.n2472 185
R17092 vdd.n2475 vdd.n2474 185
R17093 vdd.n2477 vdd.n2476 185
R17094 vdd.n2479 vdd.n2478 185
R17095 vdd.n2481 vdd.n2480 185
R17096 vdd.n2483 vdd.n2482 185
R17097 vdd.n2485 vdd.n2484 185
R17098 vdd.n2487 vdd.n2486 185
R17099 vdd.n2489 vdd.n2488 185
R17100 vdd.n2491 vdd.n2490 185
R17101 vdd.n2493 vdd.n2492 185
R17102 vdd.n2495 vdd.n2494 185
R17103 vdd.n2497 vdd.n2496 185
R17104 vdd.n2499 vdd.n2498 185
R17105 vdd.n2501 vdd.n2500 185
R17106 vdd.n2503 vdd.n2502 185
R17107 vdd.n2505 vdd.n2504 185
R17108 vdd.n2507 vdd.n2506 185
R17109 vdd.n2509 vdd.n2508 185
R17110 vdd.n2511 vdd.n2510 185
R17111 vdd.n2513 vdd.n2512 185
R17112 vdd.n2515 vdd.n2514 185
R17113 vdd.n2517 vdd.n2516 185
R17114 vdd.n2518 vdd.n926 185
R17115 vdd.n2520 vdd.n2519 185
R17116 vdd.n2521 vdd.n2520 185
R17117 vdd.n2450 vdd.n930 185
R17118 vdd.n2450 vdd.n2449 185
R17119 vdd.n2071 vdd.n931 185
R17120 vdd.t262 vdd.n931 185
R17121 vdd.n2072 vdd.n941 185
R17122 vdd.n2374 vdd.n941 185
R17123 vdd.n2075 vdd.n2074 185
R17124 vdd.n2074 vdd.n2073 185
R17125 vdd.n2076 vdd.n948 185
R17126 vdd.n2367 vdd.n948 185
R17127 vdd.n2078 vdd.n2077 185
R17128 vdd.n2077 vdd.n947 185
R17129 vdd.n2079 vdd.n955 185
R17130 vdd.n2359 vdd.n955 185
R17131 vdd.n2081 vdd.n2080 185
R17132 vdd.n2080 vdd.n954 185
R17133 vdd.n2082 vdd.n961 185
R17134 vdd.n2353 vdd.n961 185
R17135 vdd.n2084 vdd.n2083 185
R17136 vdd.n2083 vdd.n960 185
R17137 vdd.n2085 vdd.n966 185
R17138 vdd.n2347 vdd.n966 185
R17139 vdd.n2087 vdd.n2086 185
R17140 vdd.n2086 vdd.n973 185
R17141 vdd.n2088 vdd.n971 185
R17142 vdd.n2341 vdd.n971 185
R17143 vdd.n2090 vdd.n2089 185
R17144 vdd.n2089 vdd.n979 185
R17145 vdd.n2091 vdd.n977 185
R17146 vdd.n2335 vdd.n977 185
R17147 vdd.n2176 vdd.n2175 185
R17148 vdd.n2175 vdd.n2174 185
R17149 vdd.n2177 vdd.n984 185
R17150 vdd.n2329 vdd.n984 185
R17151 vdd.n2179 vdd.n2178 185
R17152 vdd.n2178 vdd.n983 185
R17153 vdd.n2180 vdd.n990 185
R17154 vdd.n2323 vdd.n990 185
R17155 vdd.n2182 vdd.n2181 185
R17156 vdd.n2181 vdd.n989 185
R17157 vdd.n2183 vdd.n995 185
R17158 vdd.n2317 vdd.n995 185
R17159 vdd.n2185 vdd.n2184 185
R17160 vdd.n2184 vdd.n1004 185
R17161 vdd.n2186 vdd.n1002 185
R17162 vdd.n2310 vdd.n1002 185
R17163 vdd.n2188 vdd.n2187 185
R17164 vdd.n2187 vdd.n1001 185
R17165 vdd.n2189 vdd.n1009 185
R17166 vdd.n2304 vdd.n1009 185
R17167 vdd.n2191 vdd.n2190 185
R17168 vdd.n2190 vdd.n1008 185
R17169 vdd.n2192 vdd.n1015 185
R17170 vdd.n2298 vdd.n1015 185
R17171 vdd.n2194 vdd.n2193 185
R17172 vdd.n2193 vdd.n1014 185
R17173 vdd.n2195 vdd.n1021 185
R17174 vdd.n2292 vdd.n1021 185
R17175 vdd.n370 vdd.n369 185
R17176 vdd.n3254 vdd.n370 185
R17177 vdd.n3257 vdd.n3256 185
R17178 vdd.n3256 vdd.n3255 185
R17179 vdd.n3258 vdd.n364 185
R17180 vdd.n364 vdd.n363 185
R17181 vdd.n3260 vdd.n3259 185
R17182 vdd.n3261 vdd.n3260 185
R17183 vdd.n359 vdd.n358 185
R17184 vdd.n3262 vdd.n359 185
R17185 vdd.n3265 vdd.n3264 185
R17186 vdd.n3264 vdd.n3263 185
R17187 vdd.n3266 vdd.n353 185
R17188 vdd.n3236 vdd.n353 185
R17189 vdd.n3268 vdd.n3267 185
R17190 vdd.n3269 vdd.n3268 185
R17191 vdd.n348 vdd.n347 185
R17192 vdd.n3270 vdd.n348 185
R17193 vdd.n3273 vdd.n3272 185
R17194 vdd.n3272 vdd.n3271 185
R17195 vdd.n3274 vdd.n342 185
R17196 vdd.n349 vdd.n342 185
R17197 vdd.n3276 vdd.n3275 185
R17198 vdd.n3277 vdd.n3276 185
R17199 vdd.n338 vdd.n337 185
R17200 vdd.n3278 vdd.n338 185
R17201 vdd.n3281 vdd.n3280 185
R17202 vdd.n3280 vdd.n3279 185
R17203 vdd.n3282 vdd.n333 185
R17204 vdd.n333 vdd.n332 185
R17205 vdd.n3284 vdd.n3283 185
R17206 vdd.n3285 vdd.n3284 185
R17207 vdd.n327 vdd.n325 185
R17208 vdd.n3286 vdd.n327 185
R17209 vdd.n3289 vdd.n3288 185
R17210 vdd.n3288 vdd.n3287 185
R17211 vdd.n326 vdd.n324 185
R17212 vdd.n328 vdd.n326 185
R17213 vdd.n3212 vdd.n3211 185
R17214 vdd.n3213 vdd.n3212 185
R17215 vdd.n615 vdd.n614 185
R17216 vdd.n614 vdd.n613 185
R17217 vdd.n3207 vdd.n3206 185
R17218 vdd.n3206 vdd.n3205 185
R17219 vdd.n618 vdd.n617 185
R17220 vdd.n624 vdd.n618 185
R17221 vdd.n3193 vdd.n3192 185
R17222 vdd.n3194 vdd.n3193 185
R17223 vdd.n626 vdd.n625 185
R17224 vdd.n3185 vdd.n625 185
R17225 vdd.n3188 vdd.n3187 185
R17226 vdd.n3187 vdd.n3186 185
R17227 vdd.n629 vdd.n628 185
R17228 vdd.n636 vdd.n629 185
R17229 vdd.n3176 vdd.n3175 185
R17230 vdd.n3177 vdd.n3176 185
R17231 vdd.n638 vdd.n637 185
R17232 vdd.n637 vdd.n635 185
R17233 vdd.n3171 vdd.n3170 185
R17234 vdd.n3170 vdd.n3169 185
R17235 vdd.n641 vdd.n640 185
R17236 vdd.n642 vdd.n641 185
R17237 vdd.n3160 vdd.n3159 185
R17238 vdd.n3161 vdd.n3160 185
R17239 vdd.n650 vdd.n649 185
R17240 vdd.n649 vdd.n648 185
R17241 vdd.n3155 vdd.n3154 185
R17242 vdd.n3154 vdd.n3153 185
R17243 vdd.n653 vdd.n652 185
R17244 vdd.n659 vdd.n653 185
R17245 vdd.n3144 vdd.n3143 185
R17246 vdd.n3145 vdd.n3144 185
R17247 vdd.n3140 vdd.n660 185
R17248 vdd.n3139 vdd.n3138 185
R17249 vdd.n3136 vdd.n662 185
R17250 vdd.n3136 vdd.n658 185
R17251 vdd.n3135 vdd.n3134 185
R17252 vdd.n3133 vdd.n3132 185
R17253 vdd.n3131 vdd.n3130 185
R17254 vdd.n3129 vdd.n3128 185
R17255 vdd.n3127 vdd.n668 185
R17256 vdd.n3125 vdd.n3124 185
R17257 vdd.n3123 vdd.n669 185
R17258 vdd.n3122 vdd.n3121 185
R17259 vdd.n3119 vdd.n674 185
R17260 vdd.n3117 vdd.n3116 185
R17261 vdd.n3115 vdd.n675 185
R17262 vdd.n3114 vdd.n3113 185
R17263 vdd.n3111 vdd.n680 185
R17264 vdd.n3109 vdd.n3108 185
R17265 vdd.n3107 vdd.n681 185
R17266 vdd.n3106 vdd.n3105 185
R17267 vdd.n3103 vdd.n688 185
R17268 vdd.n3101 vdd.n3100 185
R17269 vdd.n3099 vdd.n689 185
R17270 vdd.n3098 vdd.n3097 185
R17271 vdd.n3095 vdd.n694 185
R17272 vdd.n3093 vdd.n3092 185
R17273 vdd.n3091 vdd.n695 185
R17274 vdd.n3090 vdd.n3089 185
R17275 vdd.n3087 vdd.n700 185
R17276 vdd.n3085 vdd.n3084 185
R17277 vdd.n3083 vdd.n701 185
R17278 vdd.n3082 vdd.n3081 185
R17279 vdd.n3079 vdd.n706 185
R17280 vdd.n3077 vdd.n3076 185
R17281 vdd.n3075 vdd.n707 185
R17282 vdd.n3074 vdd.n3073 185
R17283 vdd.n3071 vdd.n712 185
R17284 vdd.n3069 vdd.n3068 185
R17285 vdd.n3067 vdd.n713 185
R17286 vdd.n3066 vdd.n3065 185
R17287 vdd.n3063 vdd.n718 185
R17288 vdd.n3061 vdd.n3060 185
R17289 vdd.n3059 vdd.n719 185
R17290 vdd.n728 vdd.n722 185
R17291 vdd.n3055 vdd.n3054 185
R17292 vdd.n3052 vdd.n726 185
R17293 vdd.n3051 vdd.n3050 185
R17294 vdd.n3049 vdd.n3048 185
R17295 vdd.n3047 vdd.n732 185
R17296 vdd.n3045 vdd.n3044 185
R17297 vdd.n3043 vdd.n733 185
R17298 vdd.n3042 vdd.n3041 185
R17299 vdd.n3039 vdd.n738 185
R17300 vdd.n3037 vdd.n3036 185
R17301 vdd.n3035 vdd.n739 185
R17302 vdd.n3034 vdd.n3033 185
R17303 vdd.n3031 vdd.n744 185
R17304 vdd.n3029 vdd.n3028 185
R17305 vdd.n3027 vdd.n745 185
R17306 vdd.n3026 vdd.n3025 185
R17307 vdd.n3023 vdd.n3022 185
R17308 vdd.n3021 vdd.n3020 185
R17309 vdd.n3019 vdd.n3018 185
R17310 vdd.n3017 vdd.n3016 185
R17311 vdd.n3012 vdd.n657 185
R17312 vdd.n658 vdd.n657 185
R17313 vdd.n3251 vdd.n3250 185
R17314 vdd.n599 vdd.n404 185
R17315 vdd.n598 vdd.n597 185
R17316 vdd.n596 vdd.n595 185
R17317 vdd.n594 vdd.n409 185
R17318 vdd.n590 vdd.n589 185
R17319 vdd.n588 vdd.n587 185
R17320 vdd.n586 vdd.n585 185
R17321 vdd.n584 vdd.n411 185
R17322 vdd.n580 vdd.n579 185
R17323 vdd.n578 vdd.n577 185
R17324 vdd.n576 vdd.n575 185
R17325 vdd.n574 vdd.n413 185
R17326 vdd.n570 vdd.n569 185
R17327 vdd.n568 vdd.n567 185
R17328 vdd.n566 vdd.n565 185
R17329 vdd.n564 vdd.n415 185
R17330 vdd.n560 vdd.n559 185
R17331 vdd.n558 vdd.n557 185
R17332 vdd.n556 vdd.n555 185
R17333 vdd.n554 vdd.n417 185
R17334 vdd.n550 vdd.n549 185
R17335 vdd.n548 vdd.n547 185
R17336 vdd.n546 vdd.n545 185
R17337 vdd.n544 vdd.n421 185
R17338 vdd.n540 vdd.n539 185
R17339 vdd.n538 vdd.n537 185
R17340 vdd.n536 vdd.n535 185
R17341 vdd.n534 vdd.n423 185
R17342 vdd.n530 vdd.n529 185
R17343 vdd.n528 vdd.n527 185
R17344 vdd.n526 vdd.n525 185
R17345 vdd.n524 vdd.n425 185
R17346 vdd.n520 vdd.n519 185
R17347 vdd.n518 vdd.n517 185
R17348 vdd.n516 vdd.n515 185
R17349 vdd.n514 vdd.n427 185
R17350 vdd.n510 vdd.n509 185
R17351 vdd.n508 vdd.n507 185
R17352 vdd.n506 vdd.n505 185
R17353 vdd.n504 vdd.n429 185
R17354 vdd.n500 vdd.n499 185
R17355 vdd.n498 vdd.n497 185
R17356 vdd.n496 vdd.n495 185
R17357 vdd.n494 vdd.n433 185
R17358 vdd.n490 vdd.n489 185
R17359 vdd.n488 vdd.n487 185
R17360 vdd.n486 vdd.n485 185
R17361 vdd.n484 vdd.n435 185
R17362 vdd.n480 vdd.n479 185
R17363 vdd.n478 vdd.n477 185
R17364 vdd.n476 vdd.n475 185
R17365 vdd.n474 vdd.n437 185
R17366 vdd.n470 vdd.n469 185
R17367 vdd.n468 vdd.n467 185
R17368 vdd.n466 vdd.n465 185
R17369 vdd.n464 vdd.n439 185
R17370 vdd.n460 vdd.n459 185
R17371 vdd.n458 vdd.n457 185
R17372 vdd.n456 vdd.n455 185
R17373 vdd.n454 vdd.n441 185
R17374 vdd.n450 vdd.n449 185
R17375 vdd.n448 vdd.n447 185
R17376 vdd.n446 vdd.n445 185
R17377 vdd.n3247 vdd.n372 185
R17378 vdd.n3254 vdd.n372 185
R17379 vdd.n3246 vdd.n371 185
R17380 vdd.n3255 vdd.n371 185
R17381 vdd.n3245 vdd.n3244 185
R17382 vdd.n3244 vdd.n363 185
R17383 vdd.n602 vdd.n362 185
R17384 vdd.n3261 vdd.n362 185
R17385 vdd.n3240 vdd.n361 185
R17386 vdd.n3262 vdd.n361 185
R17387 vdd.n3239 vdd.n360 185
R17388 vdd.n3263 vdd.n360 185
R17389 vdd.n3238 vdd.n3237 185
R17390 vdd.n3237 vdd.n3236 185
R17391 vdd.n604 vdd.n352 185
R17392 vdd.n3269 vdd.n352 185
R17393 vdd.n3232 vdd.n351 185
R17394 vdd.n3270 vdd.n351 185
R17395 vdd.n3231 vdd.n350 185
R17396 vdd.n3271 vdd.n350 185
R17397 vdd.n3230 vdd.n3229 185
R17398 vdd.n3229 vdd.n349 185
R17399 vdd.n606 vdd.n341 185
R17400 vdd.n3277 vdd.n341 185
R17401 vdd.n3225 vdd.n340 185
R17402 vdd.n3278 vdd.n340 185
R17403 vdd.n3224 vdd.n339 185
R17404 vdd.n3279 vdd.n339 185
R17405 vdd.n3223 vdd.n3222 185
R17406 vdd.n3222 vdd.n332 185
R17407 vdd.n608 vdd.n331 185
R17408 vdd.n3285 vdd.n331 185
R17409 vdd.n3218 vdd.n330 185
R17410 vdd.n3286 vdd.n330 185
R17411 vdd.n3217 vdd.n329 185
R17412 vdd.n3287 vdd.n329 185
R17413 vdd.n3216 vdd.n3215 185
R17414 vdd.n3215 vdd.n328 185
R17415 vdd.n3214 vdd.n610 185
R17416 vdd.n3214 vdd.n3213 185
R17417 vdd.n3202 vdd.n612 185
R17418 vdd.n613 vdd.n612 185
R17419 vdd.n3204 vdd.n3203 185
R17420 vdd.n3205 vdd.n3204 185
R17421 vdd.n620 vdd.n619 185
R17422 vdd.n624 vdd.n619 185
R17423 vdd.n3196 vdd.n3195 185
R17424 vdd.n3195 vdd.n3194 185
R17425 vdd.n623 vdd.n622 185
R17426 vdd.n3185 vdd.n623 185
R17427 vdd.n3184 vdd.n3183 185
R17428 vdd.n3186 vdd.n3184 185
R17429 vdd.n631 vdd.n630 185
R17430 vdd.n636 vdd.n630 185
R17431 vdd.n3179 vdd.n3178 185
R17432 vdd.n3178 vdd.n3177 185
R17433 vdd.n634 vdd.n633 185
R17434 vdd.n635 vdd.n634 185
R17435 vdd.n3168 vdd.n3167 185
R17436 vdd.n3169 vdd.n3168 185
R17437 vdd.n644 vdd.n643 185
R17438 vdd.n643 vdd.n642 185
R17439 vdd.n3163 vdd.n3162 185
R17440 vdd.n3162 vdd.n3161 185
R17441 vdd.n647 vdd.n646 185
R17442 vdd.n648 vdd.n647 185
R17443 vdd.n3152 vdd.n3151 185
R17444 vdd.n3153 vdd.n3152 185
R17445 vdd.n655 vdd.n654 185
R17446 vdd.n659 vdd.n654 185
R17447 vdd.n3147 vdd.n3146 185
R17448 vdd.n3146 vdd.n3145 185
R17449 vdd.n884 vdd.n883 185
R17450 vdd.n2772 vdd.n2771 185
R17451 vdd.n2770 vdd.n2555 185
R17452 vdd.n2774 vdd.n2555 185
R17453 vdd.n2769 vdd.n2768 185
R17454 vdd.n2767 vdd.n2766 185
R17455 vdd.n2765 vdd.n2764 185
R17456 vdd.n2763 vdd.n2762 185
R17457 vdd.n2761 vdd.n2760 185
R17458 vdd.n2759 vdd.n2758 185
R17459 vdd.n2757 vdd.n2756 185
R17460 vdd.n2755 vdd.n2754 185
R17461 vdd.n2753 vdd.n2752 185
R17462 vdd.n2751 vdd.n2750 185
R17463 vdd.n2749 vdd.n2748 185
R17464 vdd.n2747 vdd.n2746 185
R17465 vdd.n2745 vdd.n2744 185
R17466 vdd.n2743 vdd.n2742 185
R17467 vdd.n2741 vdd.n2740 185
R17468 vdd.n2739 vdd.n2738 185
R17469 vdd.n2737 vdd.n2736 185
R17470 vdd.n2735 vdd.n2734 185
R17471 vdd.n2733 vdd.n2732 185
R17472 vdd.n2731 vdd.n2730 185
R17473 vdd.n2729 vdd.n2728 185
R17474 vdd.n2727 vdd.n2726 185
R17475 vdd.n2725 vdd.n2724 185
R17476 vdd.n2723 vdd.n2722 185
R17477 vdd.n2721 vdd.n2720 185
R17478 vdd.n2719 vdd.n2718 185
R17479 vdd.n2717 vdd.n2716 185
R17480 vdd.n2715 vdd.n2714 185
R17481 vdd.n2713 vdd.n2712 185
R17482 vdd.n2710 vdd.n2709 185
R17483 vdd.n2708 vdd.n2707 185
R17484 vdd.n2706 vdd.n2705 185
R17485 vdd.n2913 vdd.n2912 185
R17486 vdd.n2914 vdd.n803 185
R17487 vdd.n2916 vdd.n2915 185
R17488 vdd.n2918 vdd.n801 185
R17489 vdd.n2920 vdd.n2919 185
R17490 vdd.n2921 vdd.n800 185
R17491 vdd.n2923 vdd.n2922 185
R17492 vdd.n2925 vdd.n798 185
R17493 vdd.n2927 vdd.n2926 185
R17494 vdd.n2928 vdd.n797 185
R17495 vdd.n2930 vdd.n2929 185
R17496 vdd.n2932 vdd.n795 185
R17497 vdd.n2934 vdd.n2933 185
R17498 vdd.n2935 vdd.n794 185
R17499 vdd.n2937 vdd.n2936 185
R17500 vdd.n2939 vdd.n792 185
R17501 vdd.n2941 vdd.n2940 185
R17502 vdd.n2943 vdd.n791 185
R17503 vdd.n2945 vdd.n2944 185
R17504 vdd.n2947 vdd.n789 185
R17505 vdd.n2949 vdd.n2948 185
R17506 vdd.n2950 vdd.n788 185
R17507 vdd.n2952 vdd.n2951 185
R17508 vdd.n2954 vdd.n786 185
R17509 vdd.n2956 vdd.n2955 185
R17510 vdd.n2957 vdd.n785 185
R17511 vdd.n2959 vdd.n2958 185
R17512 vdd.n2961 vdd.n783 185
R17513 vdd.n2963 vdd.n2962 185
R17514 vdd.n2964 vdd.n782 185
R17515 vdd.n2966 vdd.n2965 185
R17516 vdd.n2968 vdd.n781 185
R17517 vdd.n2969 vdd.n780 185
R17518 vdd.n2972 vdd.n2971 185
R17519 vdd.n2973 vdd.n778 185
R17520 vdd.n778 vdd.n756 185
R17521 vdd.n2910 vdd.n775 185
R17522 vdd.n2976 vdd.n775 185
R17523 vdd.n2909 vdd.n2908 185
R17524 vdd.n2908 vdd.n774 185
R17525 vdd.n2907 vdd.n807 185
R17526 vdd.n2907 vdd.n2906 185
R17527 vdd.n2661 vdd.n808 185
R17528 vdd.n817 vdd.n808 185
R17529 vdd.n2662 vdd.n815 185
R17530 vdd.n2900 vdd.n815 185
R17531 vdd.n2664 vdd.n2663 185
R17532 vdd.n2663 vdd.n814 185
R17533 vdd.n2665 vdd.n823 185
R17534 vdd.n2849 vdd.n823 185
R17535 vdd.n2667 vdd.n2666 185
R17536 vdd.n2666 vdd.n822 185
R17537 vdd.n2668 vdd.n829 185
R17538 vdd.n2843 vdd.n829 185
R17539 vdd.n2670 vdd.n2669 185
R17540 vdd.n2669 vdd.n828 185
R17541 vdd.n2671 vdd.n834 185
R17542 vdd.n2835 vdd.n834 185
R17543 vdd.n2673 vdd.n2672 185
R17544 vdd.n2672 vdd.n841 185
R17545 vdd.n2674 vdd.n839 185
R17546 vdd.n2829 vdd.n839 185
R17547 vdd.n2676 vdd.n2675 185
R17548 vdd.n2677 vdd.n2676 185
R17549 vdd.n2660 vdd.n846 185
R17550 vdd.n2823 vdd.n846 185
R17551 vdd.n2659 vdd.n2658 185
R17552 vdd.n2658 vdd.n845 185
R17553 vdd.n2657 vdd.n852 185
R17554 vdd.n2817 vdd.n852 185
R17555 vdd.n2656 vdd.n2655 185
R17556 vdd.n2655 vdd.n851 185
R17557 vdd.n2654 vdd.n857 185
R17558 vdd.n2811 vdd.n857 185
R17559 vdd.n2653 vdd.n2652 185
R17560 vdd.n2652 vdd.n864 185
R17561 vdd.n2651 vdd.n862 185
R17562 vdd.n2805 vdd.n862 185
R17563 vdd.n2650 vdd.n2649 185
R17564 vdd.n2649 vdd.n871 185
R17565 vdd.n2648 vdd.n869 185
R17566 vdd.n2799 vdd.n869 185
R17567 vdd.n2647 vdd.n2646 185
R17568 vdd.n2646 vdd.n868 185
R17569 vdd.n2558 vdd.n875 185
R17570 vdd.n2793 vdd.n875 185
R17571 vdd.n2700 vdd.n2699 185
R17572 vdd.n2699 vdd.n2698 185
R17573 vdd.n2701 vdd.n880 185
R17574 vdd.n2787 vdd.n880 185
R17575 vdd.n2703 vdd.n2702 185
R17576 vdd.n2702 vdd.t248 185
R17577 vdd.n2704 vdd.n885 185
R17578 vdd.n2781 vdd.n885 185
R17579 vdd.n2783 vdd.n2782 185
R17580 vdd.n2782 vdd.n2781 185
R17581 vdd.n2784 vdd.n882 185
R17582 vdd.n882 vdd.t248 185
R17583 vdd.n2786 vdd.n2785 185
R17584 vdd.n2787 vdd.n2786 185
R17585 vdd.n874 vdd.n873 185
R17586 vdd.n2698 vdd.n874 185
R17587 vdd.n2795 vdd.n2794 185
R17588 vdd.n2794 vdd.n2793 185
R17589 vdd.n2796 vdd.n872 185
R17590 vdd.n872 vdd.n868 185
R17591 vdd.n2798 vdd.n2797 185
R17592 vdd.n2799 vdd.n2798 185
R17593 vdd.n861 vdd.n860 185
R17594 vdd.n871 vdd.n861 185
R17595 vdd.n2807 vdd.n2806 185
R17596 vdd.n2806 vdd.n2805 185
R17597 vdd.n2808 vdd.n859 185
R17598 vdd.n864 vdd.n859 185
R17599 vdd.n2810 vdd.n2809 185
R17600 vdd.n2811 vdd.n2810 185
R17601 vdd.n850 vdd.n849 185
R17602 vdd.n851 vdd.n850 185
R17603 vdd.n2819 vdd.n2818 185
R17604 vdd.n2818 vdd.n2817 185
R17605 vdd.n2820 vdd.n848 185
R17606 vdd.n848 vdd.n845 185
R17607 vdd.n2822 vdd.n2821 185
R17608 vdd.n2823 vdd.n2822 185
R17609 vdd.n838 vdd.n837 185
R17610 vdd.n2677 vdd.n838 185
R17611 vdd.n2831 vdd.n2830 185
R17612 vdd.n2830 vdd.n2829 185
R17613 vdd.n2832 vdd.n836 185
R17614 vdd.n841 vdd.n836 185
R17615 vdd.n2834 vdd.n2833 185
R17616 vdd.n2835 vdd.n2834 185
R17617 vdd.n827 vdd.n826 185
R17618 vdd.n828 vdd.n827 185
R17619 vdd.n2845 vdd.n2844 185
R17620 vdd.n2844 vdd.n2843 185
R17621 vdd.n2846 vdd.n825 185
R17622 vdd.n825 vdd.n822 185
R17623 vdd.n2848 vdd.n2847 185
R17624 vdd.n2849 vdd.n2848 185
R17625 vdd.n813 vdd.n812 185
R17626 vdd.n814 vdd.n813 185
R17627 vdd.n2902 vdd.n2901 185
R17628 vdd.n2901 vdd.n2900 185
R17629 vdd.n2903 vdd.n811 185
R17630 vdd.n817 vdd.n811 185
R17631 vdd.n2905 vdd.n2904 185
R17632 vdd.n2906 vdd.n2905 185
R17633 vdd.n779 vdd.n777 185
R17634 vdd.n777 vdd.n774 185
R17635 vdd.n2975 vdd.n2974 185
R17636 vdd.n2976 vdd.n2975 185
R17637 vdd.n2448 vdd.n2447 185
R17638 vdd.n2449 vdd.n2448 185
R17639 vdd.n935 vdd.n933 185
R17640 vdd.n933 vdd.t262 185
R17641 vdd.n2363 vdd.n942 185
R17642 vdd.n2374 vdd.n942 185
R17643 vdd.n2364 vdd.n951 185
R17644 vdd.n2073 vdd.n951 185
R17645 vdd.n2366 vdd.n2365 185
R17646 vdd.n2367 vdd.n2366 185
R17647 vdd.n2362 vdd.n950 185
R17648 vdd.n950 vdd.n947 185
R17649 vdd.n2361 vdd.n2360 185
R17650 vdd.n2360 vdd.n2359 185
R17651 vdd.n953 vdd.n952 185
R17652 vdd.n954 vdd.n953 185
R17653 vdd.n2352 vdd.n2351 185
R17654 vdd.n2353 vdd.n2352 185
R17655 vdd.n2350 vdd.n963 185
R17656 vdd.n963 vdd.n960 185
R17657 vdd.n2349 vdd.n2348 185
R17658 vdd.n2348 vdd.n2347 185
R17659 vdd.n965 vdd.n964 185
R17660 vdd.n973 vdd.n965 185
R17661 vdd.n2340 vdd.n2339 185
R17662 vdd.n2341 vdd.n2340 185
R17663 vdd.n2338 vdd.n974 185
R17664 vdd.n979 vdd.n974 185
R17665 vdd.n2337 vdd.n2336 185
R17666 vdd.n2336 vdd.n2335 185
R17667 vdd.n976 vdd.n975 185
R17668 vdd.n2174 vdd.n976 185
R17669 vdd.n2328 vdd.n2327 185
R17670 vdd.n2329 vdd.n2328 185
R17671 vdd.n2326 vdd.n986 185
R17672 vdd.n986 vdd.n983 185
R17673 vdd.n2325 vdd.n2324 185
R17674 vdd.n2324 vdd.n2323 185
R17675 vdd.n988 vdd.n987 185
R17676 vdd.n989 vdd.n988 185
R17677 vdd.n2316 vdd.n2315 185
R17678 vdd.n2317 vdd.n2316 185
R17679 vdd.n2313 vdd.n997 185
R17680 vdd.n1004 vdd.n997 185
R17681 vdd.n2312 vdd.n2311 185
R17682 vdd.n2311 vdd.n2310 185
R17683 vdd.n1000 vdd.n999 185
R17684 vdd.n1001 vdd.n1000 185
R17685 vdd.n2303 vdd.n2302 185
R17686 vdd.n2304 vdd.n2303 185
R17687 vdd.n2301 vdd.n1011 185
R17688 vdd.n1011 vdd.n1008 185
R17689 vdd.n2300 vdd.n2299 185
R17690 vdd.n2299 vdd.n2298 185
R17691 vdd.n1013 vdd.n1012 185
R17692 vdd.n1014 vdd.n1013 185
R17693 vdd.n2291 vdd.n2290 185
R17694 vdd.n2292 vdd.n2291 185
R17695 vdd.n2379 vdd.n907 185
R17696 vdd.n2521 vdd.n907 185
R17697 vdd.n2381 vdd.n2380 185
R17698 vdd.n2383 vdd.n2382 185
R17699 vdd.n2385 vdd.n2384 185
R17700 vdd.n2387 vdd.n2386 185
R17701 vdd.n2389 vdd.n2388 185
R17702 vdd.n2391 vdd.n2390 185
R17703 vdd.n2393 vdd.n2392 185
R17704 vdd.n2395 vdd.n2394 185
R17705 vdd.n2397 vdd.n2396 185
R17706 vdd.n2399 vdd.n2398 185
R17707 vdd.n2401 vdd.n2400 185
R17708 vdd.n2403 vdd.n2402 185
R17709 vdd.n2405 vdd.n2404 185
R17710 vdd.n2407 vdd.n2406 185
R17711 vdd.n2409 vdd.n2408 185
R17712 vdd.n2411 vdd.n2410 185
R17713 vdd.n2413 vdd.n2412 185
R17714 vdd.n2415 vdd.n2414 185
R17715 vdd.n2417 vdd.n2416 185
R17716 vdd.n2419 vdd.n2418 185
R17717 vdd.n2421 vdd.n2420 185
R17718 vdd.n2423 vdd.n2422 185
R17719 vdd.n2425 vdd.n2424 185
R17720 vdd.n2427 vdd.n2426 185
R17721 vdd.n2429 vdd.n2428 185
R17722 vdd.n2431 vdd.n2430 185
R17723 vdd.n2433 vdd.n2432 185
R17724 vdd.n2435 vdd.n2434 185
R17725 vdd.n2437 vdd.n2436 185
R17726 vdd.n2439 vdd.n2438 185
R17727 vdd.n2441 vdd.n2440 185
R17728 vdd.n2443 vdd.n2442 185
R17729 vdd.n2445 vdd.n2444 185
R17730 vdd.n2446 vdd.n934 185
R17731 vdd.n2378 vdd.n932 185
R17732 vdd.n2449 vdd.n932 185
R17733 vdd.n2377 vdd.n2376 185
R17734 vdd.n2376 vdd.t262 185
R17735 vdd.n2375 vdd.n939 185
R17736 vdd.n2375 vdd.n2374 185
R17737 vdd.n2155 vdd.n940 185
R17738 vdd.n2073 vdd.n940 185
R17739 vdd.n2156 vdd.n949 185
R17740 vdd.n2367 vdd.n949 185
R17741 vdd.n2158 vdd.n2157 185
R17742 vdd.n2157 vdd.n947 185
R17743 vdd.n2159 vdd.n956 185
R17744 vdd.n2359 vdd.n956 185
R17745 vdd.n2161 vdd.n2160 185
R17746 vdd.n2160 vdd.n954 185
R17747 vdd.n2162 vdd.n962 185
R17748 vdd.n2353 vdd.n962 185
R17749 vdd.n2164 vdd.n2163 185
R17750 vdd.n2163 vdd.n960 185
R17751 vdd.n2165 vdd.n967 185
R17752 vdd.n2347 vdd.n967 185
R17753 vdd.n2167 vdd.n2166 185
R17754 vdd.n2166 vdd.n973 185
R17755 vdd.n2168 vdd.n972 185
R17756 vdd.n2341 vdd.n972 185
R17757 vdd.n2170 vdd.n2169 185
R17758 vdd.n2169 vdd.n979 185
R17759 vdd.n2171 vdd.n978 185
R17760 vdd.n2335 vdd.n978 185
R17761 vdd.n2173 vdd.n2172 185
R17762 vdd.n2174 vdd.n2173 185
R17763 vdd.n2154 vdd.n985 185
R17764 vdd.n2329 vdd.n985 185
R17765 vdd.n2153 vdd.n2152 185
R17766 vdd.n2152 vdd.n983 185
R17767 vdd.n2151 vdd.n991 185
R17768 vdd.n2323 vdd.n991 185
R17769 vdd.n2150 vdd.n2149 185
R17770 vdd.n2149 vdd.n989 185
R17771 vdd.n2148 vdd.n996 185
R17772 vdd.n2317 vdd.n996 185
R17773 vdd.n2147 vdd.n2146 185
R17774 vdd.n2146 vdd.n1004 185
R17775 vdd.n2145 vdd.n1003 185
R17776 vdd.n2310 vdd.n1003 185
R17777 vdd.n2144 vdd.n2143 185
R17778 vdd.n2143 vdd.n1001 185
R17779 vdd.n2142 vdd.n1010 185
R17780 vdd.n2304 vdd.n1010 185
R17781 vdd.n2141 vdd.n2140 185
R17782 vdd.n2140 vdd.n1008 185
R17783 vdd.n2139 vdd.n1016 185
R17784 vdd.n2298 vdd.n1016 185
R17785 vdd.n2138 vdd.n2137 185
R17786 vdd.n2137 vdd.n1014 185
R17787 vdd.n2136 vdd.n1022 185
R17788 vdd.n2292 vdd.n1022 185
R17789 vdd.n2289 vdd.n1023 185
R17790 vdd.n2288 vdd.n2287 185
R17791 vdd.n2285 vdd.n1024 185
R17792 vdd.n2283 vdd.n2282 185
R17793 vdd.n2281 vdd.n1025 185
R17794 vdd.n2280 vdd.n2279 185
R17795 vdd.n2277 vdd.n1026 185
R17796 vdd.n2275 vdd.n2274 185
R17797 vdd.n2273 vdd.n1027 185
R17798 vdd.n2272 vdd.n2271 185
R17799 vdd.n2269 vdd.n1028 185
R17800 vdd.n2267 vdd.n2266 185
R17801 vdd.n2265 vdd.n1029 185
R17802 vdd.n2264 vdd.n2263 185
R17803 vdd.n2261 vdd.n1030 185
R17804 vdd.n2259 vdd.n2258 185
R17805 vdd.n2257 vdd.n1031 185
R17806 vdd.n2256 vdd.n1033 185
R17807 vdd.n2101 vdd.n1034 185
R17808 vdd.n2104 vdd.n2103 185
R17809 vdd.n2106 vdd.n2105 185
R17810 vdd.n2108 vdd.n2100 185
R17811 vdd.n2111 vdd.n2110 185
R17812 vdd.n2112 vdd.n2099 185
R17813 vdd.n2114 vdd.n2113 185
R17814 vdd.n2116 vdd.n2098 185
R17815 vdd.n2119 vdd.n2118 185
R17816 vdd.n2120 vdd.n2097 185
R17817 vdd.n2122 vdd.n2121 185
R17818 vdd.n2124 vdd.n2096 185
R17819 vdd.n2127 vdd.n2126 185
R17820 vdd.n2128 vdd.n2093 185
R17821 vdd.n2131 vdd.n2130 185
R17822 vdd.n2133 vdd.n2092 185
R17823 vdd.n2135 vdd.n2134 185
R17824 vdd.n2134 vdd.n1020 185
R17825 vdd.n315 vdd.n314 171.744
R17826 vdd.n314 vdd.n313 171.744
R17827 vdd.n313 vdd.n282 171.744
R17828 vdd.n306 vdd.n282 171.744
R17829 vdd.n306 vdd.n305 171.744
R17830 vdd.n305 vdd.n287 171.744
R17831 vdd.n298 vdd.n287 171.744
R17832 vdd.n298 vdd.n297 171.744
R17833 vdd.n297 vdd.n291 171.744
R17834 vdd.n260 vdd.n259 171.744
R17835 vdd.n259 vdd.n258 171.744
R17836 vdd.n258 vdd.n227 171.744
R17837 vdd.n251 vdd.n227 171.744
R17838 vdd.n251 vdd.n250 171.744
R17839 vdd.n250 vdd.n232 171.744
R17840 vdd.n243 vdd.n232 171.744
R17841 vdd.n243 vdd.n242 171.744
R17842 vdd.n242 vdd.n236 171.744
R17843 vdd.n217 vdd.n216 171.744
R17844 vdd.n216 vdd.n215 171.744
R17845 vdd.n215 vdd.n184 171.744
R17846 vdd.n208 vdd.n184 171.744
R17847 vdd.n208 vdd.n207 171.744
R17848 vdd.n207 vdd.n189 171.744
R17849 vdd.n200 vdd.n189 171.744
R17850 vdd.n200 vdd.n199 171.744
R17851 vdd.n199 vdd.n193 171.744
R17852 vdd.n162 vdd.n161 171.744
R17853 vdd.n161 vdd.n160 171.744
R17854 vdd.n160 vdd.n129 171.744
R17855 vdd.n153 vdd.n129 171.744
R17856 vdd.n153 vdd.n152 171.744
R17857 vdd.n152 vdd.n134 171.744
R17858 vdd.n145 vdd.n134 171.744
R17859 vdd.n145 vdd.n144 171.744
R17860 vdd.n144 vdd.n138 171.744
R17861 vdd.n120 vdd.n119 171.744
R17862 vdd.n119 vdd.n118 171.744
R17863 vdd.n118 vdd.n87 171.744
R17864 vdd.n111 vdd.n87 171.744
R17865 vdd.n111 vdd.n110 171.744
R17866 vdd.n110 vdd.n92 171.744
R17867 vdd.n103 vdd.n92 171.744
R17868 vdd.n103 vdd.n102 171.744
R17869 vdd.n102 vdd.n96 171.744
R17870 vdd.n65 vdd.n64 171.744
R17871 vdd.n64 vdd.n63 171.744
R17872 vdd.n63 vdd.n32 171.744
R17873 vdd.n56 vdd.n32 171.744
R17874 vdd.n56 vdd.n55 171.744
R17875 vdd.n55 vdd.n37 171.744
R17876 vdd.n48 vdd.n37 171.744
R17877 vdd.n48 vdd.n47 171.744
R17878 vdd.n47 vdd.n41 171.744
R17879 vdd.n1684 vdd.n1683 171.744
R17880 vdd.n1683 vdd.n1682 171.744
R17881 vdd.n1682 vdd.n1651 171.744
R17882 vdd.n1675 vdd.n1651 171.744
R17883 vdd.n1675 vdd.n1674 171.744
R17884 vdd.n1674 vdd.n1656 171.744
R17885 vdd.n1667 vdd.n1656 171.744
R17886 vdd.n1667 vdd.n1666 171.744
R17887 vdd.n1666 vdd.n1660 171.744
R17888 vdd.n1739 vdd.n1738 171.744
R17889 vdd.n1738 vdd.n1737 171.744
R17890 vdd.n1737 vdd.n1706 171.744
R17891 vdd.n1730 vdd.n1706 171.744
R17892 vdd.n1730 vdd.n1729 171.744
R17893 vdd.n1729 vdd.n1711 171.744
R17894 vdd.n1722 vdd.n1711 171.744
R17895 vdd.n1722 vdd.n1721 171.744
R17896 vdd.n1721 vdd.n1715 171.744
R17897 vdd.n1586 vdd.n1585 171.744
R17898 vdd.n1585 vdd.n1584 171.744
R17899 vdd.n1584 vdd.n1553 171.744
R17900 vdd.n1577 vdd.n1553 171.744
R17901 vdd.n1577 vdd.n1576 171.744
R17902 vdd.n1576 vdd.n1558 171.744
R17903 vdd.n1569 vdd.n1558 171.744
R17904 vdd.n1569 vdd.n1568 171.744
R17905 vdd.n1568 vdd.n1562 171.744
R17906 vdd.n1641 vdd.n1640 171.744
R17907 vdd.n1640 vdd.n1639 171.744
R17908 vdd.n1639 vdd.n1608 171.744
R17909 vdd.n1632 vdd.n1608 171.744
R17910 vdd.n1632 vdd.n1631 171.744
R17911 vdd.n1631 vdd.n1613 171.744
R17912 vdd.n1624 vdd.n1613 171.744
R17913 vdd.n1624 vdd.n1623 171.744
R17914 vdd.n1623 vdd.n1617 171.744
R17915 vdd.n1489 vdd.n1488 171.744
R17916 vdd.n1488 vdd.n1487 171.744
R17917 vdd.n1487 vdd.n1456 171.744
R17918 vdd.n1480 vdd.n1456 171.744
R17919 vdd.n1480 vdd.n1479 171.744
R17920 vdd.n1479 vdd.n1461 171.744
R17921 vdd.n1472 vdd.n1461 171.744
R17922 vdd.n1472 vdd.n1471 171.744
R17923 vdd.n1471 vdd.n1465 171.744
R17924 vdd.n1544 vdd.n1543 171.744
R17925 vdd.n1543 vdd.n1542 171.744
R17926 vdd.n1542 vdd.n1511 171.744
R17927 vdd.n1535 vdd.n1511 171.744
R17928 vdd.n1535 vdd.n1534 171.744
R17929 vdd.n1534 vdd.n1516 171.744
R17930 vdd.n1527 vdd.n1516 171.744
R17931 vdd.n1527 vdd.n1526 171.744
R17932 vdd.n1526 vdd.n1520 171.744
R17933 vdd.n449 vdd.n448 146.341
R17934 vdd.n455 vdd.n454 146.341
R17935 vdd.n459 vdd.n458 146.341
R17936 vdd.n465 vdd.n464 146.341
R17937 vdd.n469 vdd.n468 146.341
R17938 vdd.n475 vdd.n474 146.341
R17939 vdd.n479 vdd.n478 146.341
R17940 vdd.n485 vdd.n484 146.341
R17941 vdd.n489 vdd.n488 146.341
R17942 vdd.n495 vdd.n494 146.341
R17943 vdd.n499 vdd.n498 146.341
R17944 vdd.n505 vdd.n504 146.341
R17945 vdd.n509 vdd.n508 146.341
R17946 vdd.n515 vdd.n514 146.341
R17947 vdd.n519 vdd.n518 146.341
R17948 vdd.n525 vdd.n524 146.341
R17949 vdd.n529 vdd.n528 146.341
R17950 vdd.n535 vdd.n534 146.341
R17951 vdd.n539 vdd.n538 146.341
R17952 vdd.n545 vdd.n544 146.341
R17953 vdd.n549 vdd.n548 146.341
R17954 vdd.n555 vdd.n554 146.341
R17955 vdd.n559 vdd.n558 146.341
R17956 vdd.n565 vdd.n564 146.341
R17957 vdd.n569 vdd.n568 146.341
R17958 vdd.n575 vdd.n574 146.341
R17959 vdd.n579 vdd.n578 146.341
R17960 vdd.n585 vdd.n584 146.341
R17961 vdd.n589 vdd.n588 146.341
R17962 vdd.n595 vdd.n594 146.341
R17963 vdd.n597 vdd.n404 146.341
R17964 vdd.n3146 vdd.n654 146.341
R17965 vdd.n3152 vdd.n654 146.341
R17966 vdd.n3152 vdd.n647 146.341
R17967 vdd.n3162 vdd.n647 146.341
R17968 vdd.n3162 vdd.n643 146.341
R17969 vdd.n3168 vdd.n643 146.341
R17970 vdd.n3168 vdd.n634 146.341
R17971 vdd.n3178 vdd.n634 146.341
R17972 vdd.n3178 vdd.n630 146.341
R17973 vdd.n3184 vdd.n630 146.341
R17974 vdd.n3184 vdd.n623 146.341
R17975 vdd.n3195 vdd.n623 146.341
R17976 vdd.n3195 vdd.n619 146.341
R17977 vdd.n3204 vdd.n619 146.341
R17978 vdd.n3204 vdd.n612 146.341
R17979 vdd.n3214 vdd.n612 146.341
R17980 vdd.n3215 vdd.n3214 146.341
R17981 vdd.n3215 vdd.n329 146.341
R17982 vdd.n330 vdd.n329 146.341
R17983 vdd.n331 vdd.n330 146.341
R17984 vdd.n3222 vdd.n331 146.341
R17985 vdd.n3222 vdd.n339 146.341
R17986 vdd.n340 vdd.n339 146.341
R17987 vdd.n341 vdd.n340 146.341
R17988 vdd.n3229 vdd.n341 146.341
R17989 vdd.n3229 vdd.n350 146.341
R17990 vdd.n351 vdd.n350 146.341
R17991 vdd.n352 vdd.n351 146.341
R17992 vdd.n3237 vdd.n352 146.341
R17993 vdd.n3237 vdd.n360 146.341
R17994 vdd.n361 vdd.n360 146.341
R17995 vdd.n362 vdd.n361 146.341
R17996 vdd.n3244 vdd.n362 146.341
R17997 vdd.n3244 vdd.n371 146.341
R17998 vdd.n372 vdd.n371 146.341
R17999 vdd.n3138 vdd.n3136 146.341
R18000 vdd.n3136 vdd.n3135 146.341
R18001 vdd.n3132 vdd.n3131 146.341
R18002 vdd.n3128 vdd.n3127 146.341
R18003 vdd.n3125 vdd.n669 146.341
R18004 vdd.n3121 vdd.n3119 146.341
R18005 vdd.n3117 vdd.n675 146.341
R18006 vdd.n3113 vdd.n3111 146.341
R18007 vdd.n3109 vdd.n681 146.341
R18008 vdd.n3105 vdd.n3103 146.341
R18009 vdd.n3101 vdd.n689 146.341
R18010 vdd.n3097 vdd.n3095 146.341
R18011 vdd.n3093 vdd.n695 146.341
R18012 vdd.n3089 vdd.n3087 146.341
R18013 vdd.n3085 vdd.n701 146.341
R18014 vdd.n3081 vdd.n3079 146.341
R18015 vdd.n3077 vdd.n707 146.341
R18016 vdd.n3073 vdd.n3071 146.341
R18017 vdd.n3069 vdd.n713 146.341
R18018 vdd.n3065 vdd.n3063 146.341
R18019 vdd.n3061 vdd.n719 146.341
R18020 vdd.n3054 vdd.n728 146.341
R18021 vdd.n3052 vdd.n3051 146.341
R18022 vdd.n3048 vdd.n3047 146.341
R18023 vdd.n3045 vdd.n733 146.341
R18024 vdd.n3041 vdd.n3039 146.341
R18025 vdd.n3037 vdd.n739 146.341
R18026 vdd.n3033 vdd.n3031 146.341
R18027 vdd.n3029 vdd.n745 146.341
R18028 vdd.n3025 vdd.n3023 146.341
R18029 vdd.n3020 vdd.n3019 146.341
R18030 vdd.n3016 vdd.n657 146.341
R18031 vdd.n3144 vdd.n653 146.341
R18032 vdd.n3154 vdd.n653 146.341
R18033 vdd.n3154 vdd.n649 146.341
R18034 vdd.n3160 vdd.n649 146.341
R18035 vdd.n3160 vdd.n641 146.341
R18036 vdd.n3170 vdd.n641 146.341
R18037 vdd.n3170 vdd.n637 146.341
R18038 vdd.n3176 vdd.n637 146.341
R18039 vdd.n3176 vdd.n629 146.341
R18040 vdd.n3187 vdd.n629 146.341
R18041 vdd.n3187 vdd.n625 146.341
R18042 vdd.n3193 vdd.n625 146.341
R18043 vdd.n3193 vdd.n618 146.341
R18044 vdd.n3206 vdd.n618 146.341
R18045 vdd.n3206 vdd.n614 146.341
R18046 vdd.n3212 vdd.n614 146.341
R18047 vdd.n3212 vdd.n326 146.341
R18048 vdd.n3288 vdd.n326 146.341
R18049 vdd.n3288 vdd.n327 146.341
R18050 vdd.n3284 vdd.n327 146.341
R18051 vdd.n3284 vdd.n333 146.341
R18052 vdd.n3280 vdd.n333 146.341
R18053 vdd.n3280 vdd.n338 146.341
R18054 vdd.n3276 vdd.n338 146.341
R18055 vdd.n3276 vdd.n342 146.341
R18056 vdd.n3272 vdd.n342 146.341
R18057 vdd.n3272 vdd.n348 146.341
R18058 vdd.n3268 vdd.n348 146.341
R18059 vdd.n3268 vdd.n353 146.341
R18060 vdd.n3264 vdd.n353 146.341
R18061 vdd.n3264 vdd.n359 146.341
R18062 vdd.n3260 vdd.n359 146.341
R18063 vdd.n3260 vdd.n364 146.341
R18064 vdd.n3256 vdd.n364 146.341
R18065 vdd.n3256 vdd.n370 146.341
R18066 vdd.n2239 vdd.n2238 146.341
R18067 vdd.n2236 vdd.n1820 146.341
R18068 vdd.n2016 vdd.n1826 146.341
R18069 vdd.n2014 vdd.n2013 146.341
R18070 vdd.n2011 vdd.n1828 146.341
R18071 vdd.n2007 vdd.n2006 146.341
R18072 vdd.n2004 vdd.n1835 146.341
R18073 vdd.n2000 vdd.n1999 146.341
R18074 vdd.n1997 vdd.n1842 146.341
R18075 vdd.n1853 vdd.n1850 146.341
R18076 vdd.n1989 vdd.n1988 146.341
R18077 vdd.n1986 vdd.n1855 146.341
R18078 vdd.n1982 vdd.n1981 146.341
R18079 vdd.n1979 vdd.n1861 146.341
R18080 vdd.n1975 vdd.n1974 146.341
R18081 vdd.n1972 vdd.n1868 146.341
R18082 vdd.n1968 vdd.n1967 146.341
R18083 vdd.n1965 vdd.n1875 146.341
R18084 vdd.n1961 vdd.n1960 146.341
R18085 vdd.n1958 vdd.n1882 146.341
R18086 vdd.n1893 vdd.n1890 146.341
R18087 vdd.n1950 vdd.n1949 146.341
R18088 vdd.n1947 vdd.n1895 146.341
R18089 vdd.n1943 vdd.n1942 146.341
R18090 vdd.n1940 vdd.n1901 146.341
R18091 vdd.n1936 vdd.n1935 146.341
R18092 vdd.n1933 vdd.n1908 146.341
R18093 vdd.n1929 vdd.n1928 146.341
R18094 vdd.n1926 vdd.n1923 146.341
R18095 vdd.n1921 vdd.n1918 146.341
R18096 vdd.n1916 vdd.n1040 146.341
R18097 vdd.n1381 vdd.n1145 146.341
R18098 vdd.n1381 vdd.n1137 146.341
R18099 vdd.n1391 vdd.n1137 146.341
R18100 vdd.n1391 vdd.n1133 146.341
R18101 vdd.n1397 vdd.n1133 146.341
R18102 vdd.n1397 vdd.n1125 146.341
R18103 vdd.n1408 vdd.n1125 146.341
R18104 vdd.n1408 vdd.n1121 146.341
R18105 vdd.n1414 vdd.n1121 146.341
R18106 vdd.n1414 vdd.n1115 146.341
R18107 vdd.n1425 vdd.n1115 146.341
R18108 vdd.n1425 vdd.n1111 146.341
R18109 vdd.n1431 vdd.n1111 146.341
R18110 vdd.n1431 vdd.n1102 146.341
R18111 vdd.n1441 vdd.n1102 146.341
R18112 vdd.n1441 vdd.n1098 146.341
R18113 vdd.n1447 vdd.n1098 146.341
R18114 vdd.n1447 vdd.n1091 146.341
R18115 vdd.n1753 vdd.n1091 146.341
R18116 vdd.n1753 vdd.n1087 146.341
R18117 vdd.n1759 vdd.n1087 146.341
R18118 vdd.n1759 vdd.n1080 146.341
R18119 vdd.n1769 vdd.n1080 146.341
R18120 vdd.n1769 vdd.n1076 146.341
R18121 vdd.n1775 vdd.n1076 146.341
R18122 vdd.n1775 vdd.n1068 146.341
R18123 vdd.n1786 vdd.n1068 146.341
R18124 vdd.n1786 vdd.n1064 146.341
R18125 vdd.n1792 vdd.n1064 146.341
R18126 vdd.n1792 vdd.n1058 146.341
R18127 vdd.n1803 vdd.n1058 146.341
R18128 vdd.n1803 vdd.n1053 146.341
R18129 vdd.n1811 vdd.n1053 146.341
R18130 vdd.n1811 vdd.n1042 146.341
R18131 vdd.n2247 vdd.n1042 146.341
R18132 vdd.n1183 vdd.n1182 146.341
R18133 vdd.n1187 vdd.n1182 146.341
R18134 vdd.n1189 vdd.n1188 146.341
R18135 vdd.n1193 vdd.n1192 146.341
R18136 vdd.n1195 vdd.n1194 146.341
R18137 vdd.n1199 vdd.n1198 146.341
R18138 vdd.n1201 vdd.n1200 146.341
R18139 vdd.n1205 vdd.n1204 146.341
R18140 vdd.n1207 vdd.n1206 146.341
R18141 vdd.n1339 vdd.n1338 146.341
R18142 vdd.n1211 vdd.n1210 146.341
R18143 vdd.n1215 vdd.n1214 146.341
R18144 vdd.n1217 vdd.n1216 146.341
R18145 vdd.n1221 vdd.n1220 146.341
R18146 vdd.n1223 vdd.n1222 146.341
R18147 vdd.n1227 vdd.n1226 146.341
R18148 vdd.n1229 vdd.n1228 146.341
R18149 vdd.n1233 vdd.n1232 146.341
R18150 vdd.n1235 vdd.n1234 146.341
R18151 vdd.n1239 vdd.n1238 146.341
R18152 vdd.n1303 vdd.n1240 146.341
R18153 vdd.n1244 vdd.n1243 146.341
R18154 vdd.n1246 vdd.n1245 146.341
R18155 vdd.n1250 vdd.n1249 146.341
R18156 vdd.n1252 vdd.n1251 146.341
R18157 vdd.n1256 vdd.n1255 146.341
R18158 vdd.n1258 vdd.n1257 146.341
R18159 vdd.n1262 vdd.n1261 146.341
R18160 vdd.n1264 vdd.n1263 146.341
R18161 vdd.n1268 vdd.n1267 146.341
R18162 vdd.n1270 vdd.n1269 146.341
R18163 vdd.n1375 vdd.n1151 146.341
R18164 vdd.n1383 vdd.n1143 146.341
R18165 vdd.n1383 vdd.n1139 146.341
R18166 vdd.n1389 vdd.n1139 146.341
R18167 vdd.n1389 vdd.n1131 146.341
R18168 vdd.n1400 vdd.n1131 146.341
R18169 vdd.n1400 vdd.n1127 146.341
R18170 vdd.n1406 vdd.n1127 146.341
R18171 vdd.n1406 vdd.n1120 146.341
R18172 vdd.n1417 vdd.n1120 146.341
R18173 vdd.n1417 vdd.n1116 146.341
R18174 vdd.n1423 vdd.n1116 146.341
R18175 vdd.n1423 vdd.n1109 146.341
R18176 vdd.n1433 vdd.n1109 146.341
R18177 vdd.n1433 vdd.n1105 146.341
R18178 vdd.n1439 vdd.n1105 146.341
R18179 vdd.n1439 vdd.n1097 146.341
R18180 vdd.n1450 vdd.n1097 146.341
R18181 vdd.n1450 vdd.n1093 146.341
R18182 vdd.n1751 vdd.n1093 146.341
R18183 vdd.n1751 vdd.n1086 146.341
R18184 vdd.n1761 vdd.n1086 146.341
R18185 vdd.n1761 vdd.n1082 146.341
R18186 vdd.n1767 vdd.n1082 146.341
R18187 vdd.n1767 vdd.n1074 146.341
R18188 vdd.n1778 vdd.n1074 146.341
R18189 vdd.n1778 vdd.n1070 146.341
R18190 vdd.n1784 vdd.n1070 146.341
R18191 vdd.n1784 vdd.n1063 146.341
R18192 vdd.n1795 vdd.n1063 146.341
R18193 vdd.n1795 vdd.n1059 146.341
R18194 vdd.n1801 vdd.n1059 146.341
R18195 vdd.n1801 vdd.n1051 146.341
R18196 vdd.n1813 vdd.n1051 146.341
R18197 vdd.n1813 vdd.n1046 146.341
R18198 vdd.n2245 vdd.n1046 146.341
R18199 vdd.n1045 vdd.n1020 141.707
R18200 vdd.n756 vdd.n658 141.707
R18201 vdd.n2094 vdd.t56 127.284
R18202 vdd.n936 vdd.t41 127.284
R18203 vdd.n2068 vdd.t3 127.284
R18204 vdd.n928 vdd.t65 127.284
R18205 vdd.n2839 vdd.t28 127.284
R18206 vdd.n2839 vdd.t29 127.284
R18207 vdd.n2559 vdd.t63 127.284
R18208 vdd.n804 vdd.t45 127.284
R18209 vdd.n2556 vdd.t50 127.284
R18210 vdd.n768 vdd.t52 127.284
R18211 vdd.n998 vdd.t59 127.284
R18212 vdd.n998 vdd.t60 127.284
R18213 vdd.n22 vdd.n20 117.314
R18214 vdd.n17 vdd.n15 117.314
R18215 vdd.n27 vdd.n26 116.927
R18216 vdd.n24 vdd.n23 116.927
R18217 vdd.n22 vdd.n21 116.927
R18218 vdd.n17 vdd.n16 116.927
R18219 vdd.n19 vdd.n18 116.927
R18220 vdd.n27 vdd.n25 116.927
R18221 vdd.n2095 vdd.t55 111.188
R18222 vdd.n937 vdd.t42 111.188
R18223 vdd.n2069 vdd.t2 111.188
R18224 vdd.n929 vdd.t66 111.188
R18225 vdd.n2560 vdd.t62 111.188
R18226 vdd.n805 vdd.t46 111.188
R18227 vdd.n2557 vdd.t49 111.188
R18228 vdd.n769 vdd.t53 111.188
R18229 vdd.n2782 vdd.n882 99.5127
R18230 vdd.n2786 vdd.n882 99.5127
R18231 vdd.n2786 vdd.n874 99.5127
R18232 vdd.n2794 vdd.n874 99.5127
R18233 vdd.n2794 vdd.n872 99.5127
R18234 vdd.n2798 vdd.n872 99.5127
R18235 vdd.n2798 vdd.n861 99.5127
R18236 vdd.n2806 vdd.n861 99.5127
R18237 vdd.n2806 vdd.n859 99.5127
R18238 vdd.n2810 vdd.n859 99.5127
R18239 vdd.n2810 vdd.n850 99.5127
R18240 vdd.n2818 vdd.n850 99.5127
R18241 vdd.n2818 vdd.n848 99.5127
R18242 vdd.n2822 vdd.n848 99.5127
R18243 vdd.n2822 vdd.n838 99.5127
R18244 vdd.n2830 vdd.n838 99.5127
R18245 vdd.n2830 vdd.n836 99.5127
R18246 vdd.n2834 vdd.n836 99.5127
R18247 vdd.n2834 vdd.n827 99.5127
R18248 vdd.n2844 vdd.n827 99.5127
R18249 vdd.n2844 vdd.n825 99.5127
R18250 vdd.n2848 vdd.n825 99.5127
R18251 vdd.n2848 vdd.n813 99.5127
R18252 vdd.n2901 vdd.n813 99.5127
R18253 vdd.n2901 vdd.n811 99.5127
R18254 vdd.n2905 vdd.n811 99.5127
R18255 vdd.n2905 vdd.n777 99.5127
R18256 vdd.n2975 vdd.n777 99.5127
R18257 vdd.n2971 vdd.n778 99.5127
R18258 vdd.n2969 vdd.n2968 99.5127
R18259 vdd.n2966 vdd.n782 99.5127
R18260 vdd.n2962 vdd.n2961 99.5127
R18261 vdd.n2959 vdd.n785 99.5127
R18262 vdd.n2955 vdd.n2954 99.5127
R18263 vdd.n2952 vdd.n788 99.5127
R18264 vdd.n2948 vdd.n2947 99.5127
R18265 vdd.n2945 vdd.n791 99.5127
R18266 vdd.n2940 vdd.n2939 99.5127
R18267 vdd.n2937 vdd.n794 99.5127
R18268 vdd.n2933 vdd.n2932 99.5127
R18269 vdd.n2930 vdd.n797 99.5127
R18270 vdd.n2926 vdd.n2925 99.5127
R18271 vdd.n2923 vdd.n800 99.5127
R18272 vdd.n2919 vdd.n2918 99.5127
R18273 vdd.n2916 vdd.n803 99.5127
R18274 vdd.n2702 vdd.n885 99.5127
R18275 vdd.n2702 vdd.n880 99.5127
R18276 vdd.n2699 vdd.n880 99.5127
R18277 vdd.n2699 vdd.n875 99.5127
R18278 vdd.n2646 vdd.n875 99.5127
R18279 vdd.n2646 vdd.n869 99.5127
R18280 vdd.n2649 vdd.n869 99.5127
R18281 vdd.n2649 vdd.n862 99.5127
R18282 vdd.n2652 vdd.n862 99.5127
R18283 vdd.n2652 vdd.n857 99.5127
R18284 vdd.n2655 vdd.n857 99.5127
R18285 vdd.n2655 vdd.n852 99.5127
R18286 vdd.n2658 vdd.n852 99.5127
R18287 vdd.n2658 vdd.n846 99.5127
R18288 vdd.n2676 vdd.n846 99.5127
R18289 vdd.n2676 vdd.n839 99.5127
R18290 vdd.n2672 vdd.n839 99.5127
R18291 vdd.n2672 vdd.n834 99.5127
R18292 vdd.n2669 vdd.n834 99.5127
R18293 vdd.n2669 vdd.n829 99.5127
R18294 vdd.n2666 vdd.n829 99.5127
R18295 vdd.n2666 vdd.n823 99.5127
R18296 vdd.n2663 vdd.n823 99.5127
R18297 vdd.n2663 vdd.n815 99.5127
R18298 vdd.n815 vdd.n808 99.5127
R18299 vdd.n2907 vdd.n808 99.5127
R18300 vdd.n2908 vdd.n2907 99.5127
R18301 vdd.n2908 vdd.n775 99.5127
R18302 vdd.n2772 vdd.n2555 99.5127
R18303 vdd.n2768 vdd.n2555 99.5127
R18304 vdd.n2766 vdd.n2765 99.5127
R18305 vdd.n2762 vdd.n2761 99.5127
R18306 vdd.n2758 vdd.n2757 99.5127
R18307 vdd.n2754 vdd.n2753 99.5127
R18308 vdd.n2750 vdd.n2749 99.5127
R18309 vdd.n2746 vdd.n2745 99.5127
R18310 vdd.n2742 vdd.n2741 99.5127
R18311 vdd.n2738 vdd.n2737 99.5127
R18312 vdd.n2734 vdd.n2733 99.5127
R18313 vdd.n2730 vdd.n2729 99.5127
R18314 vdd.n2726 vdd.n2725 99.5127
R18315 vdd.n2722 vdd.n2721 99.5127
R18316 vdd.n2718 vdd.n2717 99.5127
R18317 vdd.n2714 vdd.n2713 99.5127
R18318 vdd.n2709 vdd.n2708 99.5127
R18319 vdd.n2520 vdd.n926 99.5127
R18320 vdd.n2516 vdd.n2515 99.5127
R18321 vdd.n2512 vdd.n2511 99.5127
R18322 vdd.n2508 vdd.n2507 99.5127
R18323 vdd.n2504 vdd.n2503 99.5127
R18324 vdd.n2500 vdd.n2499 99.5127
R18325 vdd.n2496 vdd.n2495 99.5127
R18326 vdd.n2492 vdd.n2491 99.5127
R18327 vdd.n2488 vdd.n2487 99.5127
R18328 vdd.n2484 vdd.n2483 99.5127
R18329 vdd.n2480 vdd.n2479 99.5127
R18330 vdd.n2476 vdd.n2475 99.5127
R18331 vdd.n2472 vdd.n2471 99.5127
R18332 vdd.n2468 vdd.n2467 99.5127
R18333 vdd.n2464 vdd.n2463 99.5127
R18334 vdd.n2460 vdd.n2459 99.5127
R18335 vdd.n2455 vdd.n2454 99.5127
R18336 vdd.n2193 vdd.n1021 99.5127
R18337 vdd.n2193 vdd.n1015 99.5127
R18338 vdd.n2190 vdd.n1015 99.5127
R18339 vdd.n2190 vdd.n1009 99.5127
R18340 vdd.n2187 vdd.n1009 99.5127
R18341 vdd.n2187 vdd.n1002 99.5127
R18342 vdd.n2184 vdd.n1002 99.5127
R18343 vdd.n2184 vdd.n995 99.5127
R18344 vdd.n2181 vdd.n995 99.5127
R18345 vdd.n2181 vdd.n990 99.5127
R18346 vdd.n2178 vdd.n990 99.5127
R18347 vdd.n2178 vdd.n984 99.5127
R18348 vdd.n2175 vdd.n984 99.5127
R18349 vdd.n2175 vdd.n977 99.5127
R18350 vdd.n2089 vdd.n977 99.5127
R18351 vdd.n2089 vdd.n971 99.5127
R18352 vdd.n2086 vdd.n971 99.5127
R18353 vdd.n2086 vdd.n966 99.5127
R18354 vdd.n2083 vdd.n966 99.5127
R18355 vdd.n2083 vdd.n961 99.5127
R18356 vdd.n2080 vdd.n961 99.5127
R18357 vdd.n2080 vdd.n955 99.5127
R18358 vdd.n2077 vdd.n955 99.5127
R18359 vdd.n2077 vdd.n948 99.5127
R18360 vdd.n2074 vdd.n948 99.5127
R18361 vdd.n2074 vdd.n941 99.5127
R18362 vdd.n941 vdd.n931 99.5127
R18363 vdd.n2450 vdd.n931 99.5127
R18364 vdd.n2028 vdd.n2026 99.5127
R18365 vdd.n2032 vdd.n2026 99.5127
R18366 vdd.n2036 vdd.n2034 99.5127
R18367 vdd.n2040 vdd.n2024 99.5127
R18368 vdd.n2044 vdd.n2042 99.5127
R18369 vdd.n2048 vdd.n2022 99.5127
R18370 vdd.n2052 vdd.n2050 99.5127
R18371 vdd.n2056 vdd.n2020 99.5127
R18372 vdd.n2059 vdd.n2058 99.5127
R18373 vdd.n2229 vdd.n2227 99.5127
R18374 vdd.n2225 vdd.n2061 99.5127
R18375 vdd.n2221 vdd.n2219 99.5127
R18376 vdd.n2217 vdd.n2063 99.5127
R18377 vdd.n2213 vdd.n2211 99.5127
R18378 vdd.n2209 vdd.n2065 99.5127
R18379 vdd.n2205 vdd.n2203 99.5127
R18380 vdd.n2201 vdd.n2067 99.5127
R18381 vdd.n2293 vdd.n1017 99.5127
R18382 vdd.n2297 vdd.n1017 99.5127
R18383 vdd.n2297 vdd.n1007 99.5127
R18384 vdd.n2305 vdd.n1007 99.5127
R18385 vdd.n2305 vdd.n1005 99.5127
R18386 vdd.n2309 vdd.n1005 99.5127
R18387 vdd.n2309 vdd.n994 99.5127
R18388 vdd.n2318 vdd.n994 99.5127
R18389 vdd.n2318 vdd.n992 99.5127
R18390 vdd.n2322 vdd.n992 99.5127
R18391 vdd.n2322 vdd.n982 99.5127
R18392 vdd.n2330 vdd.n982 99.5127
R18393 vdd.n2330 vdd.n980 99.5127
R18394 vdd.n2334 vdd.n980 99.5127
R18395 vdd.n2334 vdd.n970 99.5127
R18396 vdd.n2342 vdd.n970 99.5127
R18397 vdd.n2342 vdd.n968 99.5127
R18398 vdd.n2346 vdd.n968 99.5127
R18399 vdd.n2346 vdd.n959 99.5127
R18400 vdd.n2354 vdd.n959 99.5127
R18401 vdd.n2354 vdd.n957 99.5127
R18402 vdd.n2358 vdd.n957 99.5127
R18403 vdd.n2358 vdd.n946 99.5127
R18404 vdd.n2368 vdd.n946 99.5127
R18405 vdd.n2368 vdd.n943 99.5127
R18406 vdd.n2373 vdd.n943 99.5127
R18407 vdd.n2373 vdd.n944 99.5127
R18408 vdd.n944 vdd.n925 99.5127
R18409 vdd.n2891 vdd.n2890 99.5127
R18410 vdd.n2888 vdd.n2854 99.5127
R18411 vdd.n2884 vdd.n2883 99.5127
R18412 vdd.n2881 vdd.n2857 99.5127
R18413 vdd.n2877 vdd.n2876 99.5127
R18414 vdd.n2874 vdd.n2860 99.5127
R18415 vdd.n2870 vdd.n2869 99.5127
R18416 vdd.n2867 vdd.n2864 99.5127
R18417 vdd.n3008 vdd.n755 99.5127
R18418 vdd.n3006 vdd.n3005 99.5127
R18419 vdd.n3003 vdd.n758 99.5127
R18420 vdd.n2999 vdd.n2998 99.5127
R18421 vdd.n2996 vdd.n761 99.5127
R18422 vdd.n2992 vdd.n2991 99.5127
R18423 vdd.n2989 vdd.n764 99.5127
R18424 vdd.n2985 vdd.n2984 99.5127
R18425 vdd.n2982 vdd.n767 99.5127
R18426 vdd.n2626 vdd.n886 99.5127
R18427 vdd.n2626 vdd.n881 99.5127
R18428 vdd.n2697 vdd.n881 99.5127
R18429 vdd.n2697 vdd.n876 99.5127
R18430 vdd.n2693 vdd.n876 99.5127
R18431 vdd.n2693 vdd.n870 99.5127
R18432 vdd.n2690 vdd.n870 99.5127
R18433 vdd.n2690 vdd.n863 99.5127
R18434 vdd.n2687 vdd.n863 99.5127
R18435 vdd.n2687 vdd.n858 99.5127
R18436 vdd.n2684 vdd.n858 99.5127
R18437 vdd.n2684 vdd.n853 99.5127
R18438 vdd.n2681 vdd.n853 99.5127
R18439 vdd.n2681 vdd.n847 99.5127
R18440 vdd.n2678 vdd.n847 99.5127
R18441 vdd.n2678 vdd.n840 99.5127
R18442 vdd.n2643 vdd.n840 99.5127
R18443 vdd.n2643 vdd.n835 99.5127
R18444 vdd.n2640 vdd.n835 99.5127
R18445 vdd.n2640 vdd.n830 99.5127
R18446 vdd.n2637 vdd.n830 99.5127
R18447 vdd.n2637 vdd.n824 99.5127
R18448 vdd.n2634 vdd.n824 99.5127
R18449 vdd.n2634 vdd.n816 99.5127
R18450 vdd.n2631 vdd.n816 99.5127
R18451 vdd.n2631 vdd.n809 99.5127
R18452 vdd.n809 vdd.n773 99.5127
R18453 vdd.n2977 vdd.n773 99.5127
R18454 vdd.n2776 vdd.n889 99.5127
R18455 vdd.n2564 vdd.n2563 99.5127
R18456 vdd.n2568 vdd.n2567 99.5127
R18457 vdd.n2572 vdd.n2571 99.5127
R18458 vdd.n2576 vdd.n2575 99.5127
R18459 vdd.n2580 vdd.n2579 99.5127
R18460 vdd.n2584 vdd.n2583 99.5127
R18461 vdd.n2588 vdd.n2587 99.5127
R18462 vdd.n2592 vdd.n2591 99.5127
R18463 vdd.n2596 vdd.n2595 99.5127
R18464 vdd.n2600 vdd.n2599 99.5127
R18465 vdd.n2604 vdd.n2603 99.5127
R18466 vdd.n2608 vdd.n2607 99.5127
R18467 vdd.n2612 vdd.n2611 99.5127
R18468 vdd.n2616 vdd.n2615 99.5127
R18469 vdd.n2620 vdd.n2619 99.5127
R18470 vdd.n2622 vdd.n2554 99.5127
R18471 vdd.n2780 vdd.n879 99.5127
R18472 vdd.n2788 vdd.n879 99.5127
R18473 vdd.n2788 vdd.n877 99.5127
R18474 vdd.n2792 vdd.n877 99.5127
R18475 vdd.n2792 vdd.n867 99.5127
R18476 vdd.n2800 vdd.n867 99.5127
R18477 vdd.n2800 vdd.n865 99.5127
R18478 vdd.n2804 vdd.n865 99.5127
R18479 vdd.n2804 vdd.n856 99.5127
R18480 vdd.n2812 vdd.n856 99.5127
R18481 vdd.n2812 vdd.n854 99.5127
R18482 vdd.n2816 vdd.n854 99.5127
R18483 vdd.n2816 vdd.n844 99.5127
R18484 vdd.n2824 vdd.n844 99.5127
R18485 vdd.n2824 vdd.n842 99.5127
R18486 vdd.n2828 vdd.n842 99.5127
R18487 vdd.n2828 vdd.n833 99.5127
R18488 vdd.n2836 vdd.n833 99.5127
R18489 vdd.n2836 vdd.n831 99.5127
R18490 vdd.n2842 vdd.n831 99.5127
R18491 vdd.n2842 vdd.n821 99.5127
R18492 vdd.n2850 vdd.n821 99.5127
R18493 vdd.n2850 vdd.n818 99.5127
R18494 vdd.n2899 vdd.n818 99.5127
R18495 vdd.n2899 vdd.n819 99.5127
R18496 vdd.n819 vdd.n810 99.5127
R18497 vdd.n2894 vdd.n810 99.5127
R18498 vdd.n2894 vdd.n776 99.5127
R18499 vdd.n2444 vdd.n2443 99.5127
R18500 vdd.n2440 vdd.n2439 99.5127
R18501 vdd.n2436 vdd.n2435 99.5127
R18502 vdd.n2432 vdd.n2431 99.5127
R18503 vdd.n2428 vdd.n2427 99.5127
R18504 vdd.n2424 vdd.n2423 99.5127
R18505 vdd.n2420 vdd.n2419 99.5127
R18506 vdd.n2416 vdd.n2415 99.5127
R18507 vdd.n2412 vdd.n2411 99.5127
R18508 vdd.n2408 vdd.n2407 99.5127
R18509 vdd.n2404 vdd.n2403 99.5127
R18510 vdd.n2400 vdd.n2399 99.5127
R18511 vdd.n2396 vdd.n2395 99.5127
R18512 vdd.n2392 vdd.n2391 99.5127
R18513 vdd.n2388 vdd.n2387 99.5127
R18514 vdd.n2384 vdd.n2383 99.5127
R18515 vdd.n2380 vdd.n907 99.5127
R18516 vdd.n2137 vdd.n1022 99.5127
R18517 vdd.n2137 vdd.n1016 99.5127
R18518 vdd.n2140 vdd.n1016 99.5127
R18519 vdd.n2140 vdd.n1010 99.5127
R18520 vdd.n2143 vdd.n1010 99.5127
R18521 vdd.n2143 vdd.n1003 99.5127
R18522 vdd.n2146 vdd.n1003 99.5127
R18523 vdd.n2146 vdd.n996 99.5127
R18524 vdd.n2149 vdd.n996 99.5127
R18525 vdd.n2149 vdd.n991 99.5127
R18526 vdd.n2152 vdd.n991 99.5127
R18527 vdd.n2152 vdd.n985 99.5127
R18528 vdd.n2173 vdd.n985 99.5127
R18529 vdd.n2173 vdd.n978 99.5127
R18530 vdd.n2169 vdd.n978 99.5127
R18531 vdd.n2169 vdd.n972 99.5127
R18532 vdd.n2166 vdd.n972 99.5127
R18533 vdd.n2166 vdd.n967 99.5127
R18534 vdd.n2163 vdd.n967 99.5127
R18535 vdd.n2163 vdd.n962 99.5127
R18536 vdd.n2160 vdd.n962 99.5127
R18537 vdd.n2160 vdd.n956 99.5127
R18538 vdd.n2157 vdd.n956 99.5127
R18539 vdd.n2157 vdd.n949 99.5127
R18540 vdd.n949 vdd.n940 99.5127
R18541 vdd.n2375 vdd.n940 99.5127
R18542 vdd.n2376 vdd.n2375 99.5127
R18543 vdd.n2376 vdd.n932 99.5127
R18544 vdd.n2287 vdd.n2285 99.5127
R18545 vdd.n2283 vdd.n1025 99.5127
R18546 vdd.n2279 vdd.n2277 99.5127
R18547 vdd.n2275 vdd.n1027 99.5127
R18548 vdd.n2271 vdd.n2269 99.5127
R18549 vdd.n2267 vdd.n1029 99.5127
R18550 vdd.n2263 vdd.n2261 99.5127
R18551 vdd.n2259 vdd.n1031 99.5127
R18552 vdd.n2101 vdd.n1033 99.5127
R18553 vdd.n2106 vdd.n2103 99.5127
R18554 vdd.n2110 vdd.n2108 99.5127
R18555 vdd.n2114 vdd.n2099 99.5127
R18556 vdd.n2118 vdd.n2116 99.5127
R18557 vdd.n2122 vdd.n2097 99.5127
R18558 vdd.n2126 vdd.n2124 99.5127
R18559 vdd.n2131 vdd.n2093 99.5127
R18560 vdd.n2134 vdd.n2133 99.5127
R18561 vdd.n2291 vdd.n1013 99.5127
R18562 vdd.n2299 vdd.n1013 99.5127
R18563 vdd.n2299 vdd.n1011 99.5127
R18564 vdd.n2303 vdd.n1011 99.5127
R18565 vdd.n2303 vdd.n1000 99.5127
R18566 vdd.n2311 vdd.n1000 99.5127
R18567 vdd.n2311 vdd.n997 99.5127
R18568 vdd.n2316 vdd.n997 99.5127
R18569 vdd.n2316 vdd.n988 99.5127
R18570 vdd.n2324 vdd.n988 99.5127
R18571 vdd.n2324 vdd.n986 99.5127
R18572 vdd.n2328 vdd.n986 99.5127
R18573 vdd.n2328 vdd.n976 99.5127
R18574 vdd.n2336 vdd.n976 99.5127
R18575 vdd.n2336 vdd.n974 99.5127
R18576 vdd.n2340 vdd.n974 99.5127
R18577 vdd.n2340 vdd.n965 99.5127
R18578 vdd.n2348 vdd.n965 99.5127
R18579 vdd.n2348 vdd.n963 99.5127
R18580 vdd.n2352 vdd.n963 99.5127
R18581 vdd.n2352 vdd.n953 99.5127
R18582 vdd.n2360 vdd.n953 99.5127
R18583 vdd.n2360 vdd.n950 99.5127
R18584 vdd.n2366 vdd.n950 99.5127
R18585 vdd.n2366 vdd.n951 99.5127
R18586 vdd.n951 vdd.n942 99.5127
R18587 vdd.n942 vdd.n933 99.5127
R18588 vdd.n2448 vdd.n933 99.5127
R18589 vdd.n9 vdd.n7 98.9633
R18590 vdd.n2 vdd.n0 98.9633
R18591 vdd.n9 vdd.n8 98.6055
R18592 vdd.n11 vdd.n10 98.6055
R18593 vdd.n13 vdd.n12 98.6055
R18594 vdd.n6 vdd.n5 98.6055
R18595 vdd.n4 vdd.n3 98.6055
R18596 vdd.n2 vdd.n1 98.6055
R18597 vdd.t214 vdd.n291 85.8723
R18598 vdd.t190 vdd.n236 85.8723
R18599 vdd.t202 vdd.n193 85.8723
R18600 vdd.t179 vdd.n138 85.8723
R18601 vdd.t136 vdd.n96 85.8723
R18602 vdd.t113 vdd.n41 85.8723
R18603 vdd.t228 vdd.n1660 85.8723
R18604 vdd.t140 vdd.n1715 85.8723
R18605 vdd.t215 vdd.n1562 85.8723
R18606 vdd.t123 vdd.n1617 85.8723
R18607 vdd.t115 vdd.n1465 85.8723
R18608 vdd.t137 vdd.n1520 85.8723
R18609 vdd.n2840 vdd.n2839 78.546
R18610 vdd.n2314 vdd.n998 78.546
R18611 vdd.n278 vdd.n277 75.1835
R18612 vdd.n276 vdd.n275 75.1835
R18613 vdd.n274 vdd.n273 75.1835
R18614 vdd.n272 vdd.n271 75.1835
R18615 vdd.n270 vdd.n269 75.1835
R18616 vdd.n268 vdd.n267 75.1835
R18617 vdd.n266 vdd.n265 75.1835
R18618 vdd.n180 vdd.n179 75.1835
R18619 vdd.n178 vdd.n177 75.1835
R18620 vdd.n176 vdd.n175 75.1835
R18621 vdd.n174 vdd.n173 75.1835
R18622 vdd.n172 vdd.n171 75.1835
R18623 vdd.n170 vdd.n169 75.1835
R18624 vdd.n168 vdd.n167 75.1835
R18625 vdd.n83 vdd.n82 75.1835
R18626 vdd.n81 vdd.n80 75.1835
R18627 vdd.n79 vdd.n78 75.1835
R18628 vdd.n77 vdd.n76 75.1835
R18629 vdd.n75 vdd.n74 75.1835
R18630 vdd.n73 vdd.n72 75.1835
R18631 vdd.n71 vdd.n70 75.1835
R18632 vdd.n1690 vdd.n1689 75.1835
R18633 vdd.n1692 vdd.n1691 75.1835
R18634 vdd.n1694 vdd.n1693 75.1835
R18635 vdd.n1696 vdd.n1695 75.1835
R18636 vdd.n1698 vdd.n1697 75.1835
R18637 vdd.n1700 vdd.n1699 75.1835
R18638 vdd.n1702 vdd.n1701 75.1835
R18639 vdd.n1592 vdd.n1591 75.1835
R18640 vdd.n1594 vdd.n1593 75.1835
R18641 vdd.n1596 vdd.n1595 75.1835
R18642 vdd.n1598 vdd.n1597 75.1835
R18643 vdd.n1600 vdd.n1599 75.1835
R18644 vdd.n1602 vdd.n1601 75.1835
R18645 vdd.n1604 vdd.n1603 75.1835
R18646 vdd.n1495 vdd.n1494 75.1835
R18647 vdd.n1497 vdd.n1496 75.1835
R18648 vdd.n1499 vdd.n1498 75.1835
R18649 vdd.n1501 vdd.n1500 75.1835
R18650 vdd.n1503 vdd.n1502 75.1835
R18651 vdd.n1505 vdd.n1504 75.1835
R18652 vdd.n1507 vdd.n1506 75.1835
R18653 vdd.n2775 vdd.n2774 72.8958
R18654 vdd.n2774 vdd.n2538 72.8958
R18655 vdd.n2774 vdd.n2539 72.8958
R18656 vdd.n2774 vdd.n2540 72.8958
R18657 vdd.n2774 vdd.n2541 72.8958
R18658 vdd.n2774 vdd.n2542 72.8958
R18659 vdd.n2774 vdd.n2543 72.8958
R18660 vdd.n2774 vdd.n2544 72.8958
R18661 vdd.n2774 vdd.n2545 72.8958
R18662 vdd.n2774 vdd.n2546 72.8958
R18663 vdd.n2774 vdd.n2547 72.8958
R18664 vdd.n2774 vdd.n2548 72.8958
R18665 vdd.n2774 vdd.n2549 72.8958
R18666 vdd.n2774 vdd.n2550 72.8958
R18667 vdd.n2774 vdd.n2551 72.8958
R18668 vdd.n2774 vdd.n2552 72.8958
R18669 vdd.n2774 vdd.n2553 72.8958
R18670 vdd.n772 vdd.n756 72.8958
R18671 vdd.n2983 vdd.n756 72.8958
R18672 vdd.n766 vdd.n756 72.8958
R18673 vdd.n2990 vdd.n756 72.8958
R18674 vdd.n763 vdd.n756 72.8958
R18675 vdd.n2997 vdd.n756 72.8958
R18676 vdd.n760 vdd.n756 72.8958
R18677 vdd.n3004 vdd.n756 72.8958
R18678 vdd.n3007 vdd.n756 72.8958
R18679 vdd.n2863 vdd.n756 72.8958
R18680 vdd.n2868 vdd.n756 72.8958
R18681 vdd.n2862 vdd.n756 72.8958
R18682 vdd.n2875 vdd.n756 72.8958
R18683 vdd.n2859 vdd.n756 72.8958
R18684 vdd.n2882 vdd.n756 72.8958
R18685 vdd.n2856 vdd.n756 72.8958
R18686 vdd.n2889 vdd.n756 72.8958
R18687 vdd.n2027 vdd.n1020 72.8958
R18688 vdd.n2033 vdd.n1020 72.8958
R18689 vdd.n2035 vdd.n1020 72.8958
R18690 vdd.n2041 vdd.n1020 72.8958
R18691 vdd.n2043 vdd.n1020 72.8958
R18692 vdd.n2049 vdd.n1020 72.8958
R18693 vdd.n2051 vdd.n1020 72.8958
R18694 vdd.n2057 vdd.n1020 72.8958
R18695 vdd.n2228 vdd.n1020 72.8958
R18696 vdd.n2226 vdd.n1020 72.8958
R18697 vdd.n2220 vdd.n1020 72.8958
R18698 vdd.n2218 vdd.n1020 72.8958
R18699 vdd.n2212 vdd.n1020 72.8958
R18700 vdd.n2210 vdd.n1020 72.8958
R18701 vdd.n2204 vdd.n1020 72.8958
R18702 vdd.n2202 vdd.n1020 72.8958
R18703 vdd.n2196 vdd.n1020 72.8958
R18704 vdd.n2521 vdd.n908 72.8958
R18705 vdd.n2521 vdd.n909 72.8958
R18706 vdd.n2521 vdd.n910 72.8958
R18707 vdd.n2521 vdd.n911 72.8958
R18708 vdd.n2521 vdd.n912 72.8958
R18709 vdd.n2521 vdd.n913 72.8958
R18710 vdd.n2521 vdd.n914 72.8958
R18711 vdd.n2521 vdd.n915 72.8958
R18712 vdd.n2521 vdd.n916 72.8958
R18713 vdd.n2521 vdd.n917 72.8958
R18714 vdd.n2521 vdd.n918 72.8958
R18715 vdd.n2521 vdd.n919 72.8958
R18716 vdd.n2521 vdd.n920 72.8958
R18717 vdd.n2521 vdd.n921 72.8958
R18718 vdd.n2521 vdd.n922 72.8958
R18719 vdd.n2521 vdd.n923 72.8958
R18720 vdd.n2521 vdd.n924 72.8958
R18721 vdd.n2774 vdd.n2773 72.8958
R18722 vdd.n2774 vdd.n2522 72.8958
R18723 vdd.n2774 vdd.n2523 72.8958
R18724 vdd.n2774 vdd.n2524 72.8958
R18725 vdd.n2774 vdd.n2525 72.8958
R18726 vdd.n2774 vdd.n2526 72.8958
R18727 vdd.n2774 vdd.n2527 72.8958
R18728 vdd.n2774 vdd.n2528 72.8958
R18729 vdd.n2774 vdd.n2529 72.8958
R18730 vdd.n2774 vdd.n2530 72.8958
R18731 vdd.n2774 vdd.n2531 72.8958
R18732 vdd.n2774 vdd.n2532 72.8958
R18733 vdd.n2774 vdd.n2533 72.8958
R18734 vdd.n2774 vdd.n2534 72.8958
R18735 vdd.n2774 vdd.n2535 72.8958
R18736 vdd.n2774 vdd.n2536 72.8958
R18737 vdd.n2774 vdd.n2537 72.8958
R18738 vdd.n2911 vdd.n756 72.8958
R18739 vdd.n2917 vdd.n756 72.8958
R18740 vdd.n802 vdd.n756 72.8958
R18741 vdd.n2924 vdd.n756 72.8958
R18742 vdd.n799 vdd.n756 72.8958
R18743 vdd.n2931 vdd.n756 72.8958
R18744 vdd.n796 vdd.n756 72.8958
R18745 vdd.n2938 vdd.n756 72.8958
R18746 vdd.n793 vdd.n756 72.8958
R18747 vdd.n2946 vdd.n756 72.8958
R18748 vdd.n790 vdd.n756 72.8958
R18749 vdd.n2953 vdd.n756 72.8958
R18750 vdd.n787 vdd.n756 72.8958
R18751 vdd.n2960 vdd.n756 72.8958
R18752 vdd.n784 vdd.n756 72.8958
R18753 vdd.n2967 vdd.n756 72.8958
R18754 vdd.n2970 vdd.n756 72.8958
R18755 vdd.n2521 vdd.n906 72.8958
R18756 vdd.n2521 vdd.n905 72.8958
R18757 vdd.n2521 vdd.n904 72.8958
R18758 vdd.n2521 vdd.n903 72.8958
R18759 vdd.n2521 vdd.n902 72.8958
R18760 vdd.n2521 vdd.n901 72.8958
R18761 vdd.n2521 vdd.n900 72.8958
R18762 vdd.n2521 vdd.n899 72.8958
R18763 vdd.n2521 vdd.n898 72.8958
R18764 vdd.n2521 vdd.n897 72.8958
R18765 vdd.n2521 vdd.n896 72.8958
R18766 vdd.n2521 vdd.n895 72.8958
R18767 vdd.n2521 vdd.n894 72.8958
R18768 vdd.n2521 vdd.n893 72.8958
R18769 vdd.n2521 vdd.n892 72.8958
R18770 vdd.n2521 vdd.n891 72.8958
R18771 vdd.n2521 vdd.n890 72.8958
R18772 vdd.n2286 vdd.n1020 72.8958
R18773 vdd.n2284 vdd.n1020 72.8958
R18774 vdd.n2278 vdd.n1020 72.8958
R18775 vdd.n2276 vdd.n1020 72.8958
R18776 vdd.n2270 vdd.n1020 72.8958
R18777 vdd.n2268 vdd.n1020 72.8958
R18778 vdd.n2262 vdd.n1020 72.8958
R18779 vdd.n2260 vdd.n1020 72.8958
R18780 vdd.n1032 vdd.n1020 72.8958
R18781 vdd.n2102 vdd.n1020 72.8958
R18782 vdd.n2107 vdd.n1020 72.8958
R18783 vdd.n2109 vdd.n1020 72.8958
R18784 vdd.n2115 vdd.n1020 72.8958
R18785 vdd.n2117 vdd.n1020 72.8958
R18786 vdd.n2123 vdd.n1020 72.8958
R18787 vdd.n2125 vdd.n1020 72.8958
R18788 vdd.n2132 vdd.n1020 72.8958
R18789 vdd.n1374 vdd.n1373 66.2847
R18790 vdd.n1374 vdd.n1152 66.2847
R18791 vdd.n1374 vdd.n1153 66.2847
R18792 vdd.n1374 vdd.n1154 66.2847
R18793 vdd.n1374 vdd.n1155 66.2847
R18794 vdd.n1374 vdd.n1156 66.2847
R18795 vdd.n1374 vdd.n1157 66.2847
R18796 vdd.n1374 vdd.n1158 66.2847
R18797 vdd.n1374 vdd.n1159 66.2847
R18798 vdd.n1374 vdd.n1160 66.2847
R18799 vdd.n1374 vdd.n1161 66.2847
R18800 vdd.n1374 vdd.n1162 66.2847
R18801 vdd.n1374 vdd.n1163 66.2847
R18802 vdd.n1374 vdd.n1164 66.2847
R18803 vdd.n1374 vdd.n1165 66.2847
R18804 vdd.n1374 vdd.n1166 66.2847
R18805 vdd.n1374 vdd.n1167 66.2847
R18806 vdd.n1374 vdd.n1168 66.2847
R18807 vdd.n1374 vdd.n1169 66.2847
R18808 vdd.n1374 vdd.n1170 66.2847
R18809 vdd.n1374 vdd.n1171 66.2847
R18810 vdd.n1374 vdd.n1172 66.2847
R18811 vdd.n1374 vdd.n1173 66.2847
R18812 vdd.n1374 vdd.n1174 66.2847
R18813 vdd.n1374 vdd.n1175 66.2847
R18814 vdd.n1374 vdd.n1176 66.2847
R18815 vdd.n1374 vdd.n1177 66.2847
R18816 vdd.n1374 vdd.n1178 66.2847
R18817 vdd.n1374 vdd.n1179 66.2847
R18818 vdd.n1374 vdd.n1180 66.2847
R18819 vdd.n1374 vdd.n1181 66.2847
R18820 vdd.n1045 vdd.n1041 66.2847
R18821 vdd.n1917 vdd.n1045 66.2847
R18822 vdd.n1922 vdd.n1045 66.2847
R18823 vdd.n1927 vdd.n1045 66.2847
R18824 vdd.n1915 vdd.n1045 66.2847
R18825 vdd.n1934 vdd.n1045 66.2847
R18826 vdd.n1907 vdd.n1045 66.2847
R18827 vdd.n1941 vdd.n1045 66.2847
R18828 vdd.n1900 vdd.n1045 66.2847
R18829 vdd.n1948 vdd.n1045 66.2847
R18830 vdd.n1894 vdd.n1045 66.2847
R18831 vdd.n1889 vdd.n1045 66.2847
R18832 vdd.n1959 vdd.n1045 66.2847
R18833 vdd.n1881 vdd.n1045 66.2847
R18834 vdd.n1966 vdd.n1045 66.2847
R18835 vdd.n1874 vdd.n1045 66.2847
R18836 vdd.n1973 vdd.n1045 66.2847
R18837 vdd.n1867 vdd.n1045 66.2847
R18838 vdd.n1980 vdd.n1045 66.2847
R18839 vdd.n1860 vdd.n1045 66.2847
R18840 vdd.n1987 vdd.n1045 66.2847
R18841 vdd.n1854 vdd.n1045 66.2847
R18842 vdd.n1849 vdd.n1045 66.2847
R18843 vdd.n1998 vdd.n1045 66.2847
R18844 vdd.n1841 vdd.n1045 66.2847
R18845 vdd.n2005 vdd.n1045 66.2847
R18846 vdd.n1834 vdd.n1045 66.2847
R18847 vdd.n2012 vdd.n1045 66.2847
R18848 vdd.n2015 vdd.n1045 66.2847
R18849 vdd.n1825 vdd.n1045 66.2847
R18850 vdd.n2237 vdd.n1045 66.2847
R18851 vdd.n1819 vdd.n1045 66.2847
R18852 vdd.n3137 vdd.n658 66.2847
R18853 vdd.n663 vdd.n658 66.2847
R18854 vdd.n666 vdd.n658 66.2847
R18855 vdd.n3126 vdd.n658 66.2847
R18856 vdd.n3120 vdd.n658 66.2847
R18857 vdd.n3118 vdd.n658 66.2847
R18858 vdd.n3112 vdd.n658 66.2847
R18859 vdd.n3110 vdd.n658 66.2847
R18860 vdd.n3104 vdd.n658 66.2847
R18861 vdd.n3102 vdd.n658 66.2847
R18862 vdd.n3096 vdd.n658 66.2847
R18863 vdd.n3094 vdd.n658 66.2847
R18864 vdd.n3088 vdd.n658 66.2847
R18865 vdd.n3086 vdd.n658 66.2847
R18866 vdd.n3080 vdd.n658 66.2847
R18867 vdd.n3078 vdd.n658 66.2847
R18868 vdd.n3072 vdd.n658 66.2847
R18869 vdd.n3070 vdd.n658 66.2847
R18870 vdd.n3064 vdd.n658 66.2847
R18871 vdd.n3062 vdd.n658 66.2847
R18872 vdd.n727 vdd.n658 66.2847
R18873 vdd.n3053 vdd.n658 66.2847
R18874 vdd.n729 vdd.n658 66.2847
R18875 vdd.n3046 vdd.n658 66.2847
R18876 vdd.n3040 vdd.n658 66.2847
R18877 vdd.n3038 vdd.n658 66.2847
R18878 vdd.n3032 vdd.n658 66.2847
R18879 vdd.n3030 vdd.n658 66.2847
R18880 vdd.n3024 vdd.n658 66.2847
R18881 vdd.n750 vdd.n658 66.2847
R18882 vdd.n752 vdd.n658 66.2847
R18883 vdd.n3253 vdd.n3252 66.2847
R18884 vdd.n3253 vdd.n403 66.2847
R18885 vdd.n3253 vdd.n402 66.2847
R18886 vdd.n3253 vdd.n401 66.2847
R18887 vdd.n3253 vdd.n400 66.2847
R18888 vdd.n3253 vdd.n399 66.2847
R18889 vdd.n3253 vdd.n398 66.2847
R18890 vdd.n3253 vdd.n397 66.2847
R18891 vdd.n3253 vdd.n396 66.2847
R18892 vdd.n3253 vdd.n395 66.2847
R18893 vdd.n3253 vdd.n394 66.2847
R18894 vdd.n3253 vdd.n393 66.2847
R18895 vdd.n3253 vdd.n392 66.2847
R18896 vdd.n3253 vdd.n391 66.2847
R18897 vdd.n3253 vdd.n390 66.2847
R18898 vdd.n3253 vdd.n389 66.2847
R18899 vdd.n3253 vdd.n388 66.2847
R18900 vdd.n3253 vdd.n387 66.2847
R18901 vdd.n3253 vdd.n386 66.2847
R18902 vdd.n3253 vdd.n385 66.2847
R18903 vdd.n3253 vdd.n384 66.2847
R18904 vdd.n3253 vdd.n383 66.2847
R18905 vdd.n3253 vdd.n382 66.2847
R18906 vdd.n3253 vdd.n381 66.2847
R18907 vdd.n3253 vdd.n380 66.2847
R18908 vdd.n3253 vdd.n379 66.2847
R18909 vdd.n3253 vdd.n378 66.2847
R18910 vdd.n3253 vdd.n377 66.2847
R18911 vdd.n3253 vdd.n376 66.2847
R18912 vdd.n3253 vdd.n375 66.2847
R18913 vdd.n3253 vdd.n374 66.2847
R18914 vdd.n3253 vdd.n373 66.2847
R18915 vdd.n448 vdd.n373 52.4337
R18916 vdd.n454 vdd.n374 52.4337
R18917 vdd.n458 vdd.n375 52.4337
R18918 vdd.n464 vdd.n376 52.4337
R18919 vdd.n468 vdd.n377 52.4337
R18920 vdd.n474 vdd.n378 52.4337
R18921 vdd.n478 vdd.n379 52.4337
R18922 vdd.n484 vdd.n380 52.4337
R18923 vdd.n488 vdd.n381 52.4337
R18924 vdd.n494 vdd.n382 52.4337
R18925 vdd.n498 vdd.n383 52.4337
R18926 vdd.n504 vdd.n384 52.4337
R18927 vdd.n508 vdd.n385 52.4337
R18928 vdd.n514 vdd.n386 52.4337
R18929 vdd.n518 vdd.n387 52.4337
R18930 vdd.n524 vdd.n388 52.4337
R18931 vdd.n528 vdd.n389 52.4337
R18932 vdd.n534 vdd.n390 52.4337
R18933 vdd.n538 vdd.n391 52.4337
R18934 vdd.n544 vdd.n392 52.4337
R18935 vdd.n548 vdd.n393 52.4337
R18936 vdd.n554 vdd.n394 52.4337
R18937 vdd.n558 vdd.n395 52.4337
R18938 vdd.n564 vdd.n396 52.4337
R18939 vdd.n568 vdd.n397 52.4337
R18940 vdd.n574 vdd.n398 52.4337
R18941 vdd.n578 vdd.n399 52.4337
R18942 vdd.n584 vdd.n400 52.4337
R18943 vdd.n588 vdd.n401 52.4337
R18944 vdd.n594 vdd.n402 52.4337
R18945 vdd.n597 vdd.n403 52.4337
R18946 vdd.n3252 vdd.n3251 52.4337
R18947 vdd.n3137 vdd.n660 52.4337
R18948 vdd.n3135 vdd.n663 52.4337
R18949 vdd.n3131 vdd.n666 52.4337
R18950 vdd.n3127 vdd.n3126 52.4337
R18951 vdd.n3120 vdd.n669 52.4337
R18952 vdd.n3119 vdd.n3118 52.4337
R18953 vdd.n3112 vdd.n675 52.4337
R18954 vdd.n3111 vdd.n3110 52.4337
R18955 vdd.n3104 vdd.n681 52.4337
R18956 vdd.n3103 vdd.n3102 52.4337
R18957 vdd.n3096 vdd.n689 52.4337
R18958 vdd.n3095 vdd.n3094 52.4337
R18959 vdd.n3088 vdd.n695 52.4337
R18960 vdd.n3087 vdd.n3086 52.4337
R18961 vdd.n3080 vdd.n701 52.4337
R18962 vdd.n3079 vdd.n3078 52.4337
R18963 vdd.n3072 vdd.n707 52.4337
R18964 vdd.n3071 vdd.n3070 52.4337
R18965 vdd.n3064 vdd.n713 52.4337
R18966 vdd.n3063 vdd.n3062 52.4337
R18967 vdd.n727 vdd.n719 52.4337
R18968 vdd.n3054 vdd.n3053 52.4337
R18969 vdd.n3051 vdd.n729 52.4337
R18970 vdd.n3047 vdd.n3046 52.4337
R18971 vdd.n3040 vdd.n733 52.4337
R18972 vdd.n3039 vdd.n3038 52.4337
R18973 vdd.n3032 vdd.n739 52.4337
R18974 vdd.n3031 vdd.n3030 52.4337
R18975 vdd.n3024 vdd.n745 52.4337
R18976 vdd.n3023 vdd.n750 52.4337
R18977 vdd.n3019 vdd.n752 52.4337
R18978 vdd.n2239 vdd.n1819 52.4337
R18979 vdd.n2237 vdd.n2236 52.4337
R18980 vdd.n1826 vdd.n1825 52.4337
R18981 vdd.n2015 vdd.n2014 52.4337
R18982 vdd.n2012 vdd.n2011 52.4337
R18983 vdd.n2007 vdd.n1834 52.4337
R18984 vdd.n2005 vdd.n2004 52.4337
R18985 vdd.n2000 vdd.n1841 52.4337
R18986 vdd.n1998 vdd.n1997 52.4337
R18987 vdd.n1850 vdd.n1849 52.4337
R18988 vdd.n1989 vdd.n1854 52.4337
R18989 vdd.n1987 vdd.n1986 52.4337
R18990 vdd.n1982 vdd.n1860 52.4337
R18991 vdd.n1980 vdd.n1979 52.4337
R18992 vdd.n1975 vdd.n1867 52.4337
R18993 vdd.n1973 vdd.n1972 52.4337
R18994 vdd.n1968 vdd.n1874 52.4337
R18995 vdd.n1966 vdd.n1965 52.4337
R18996 vdd.n1961 vdd.n1881 52.4337
R18997 vdd.n1959 vdd.n1958 52.4337
R18998 vdd.n1890 vdd.n1889 52.4337
R18999 vdd.n1950 vdd.n1894 52.4337
R19000 vdd.n1948 vdd.n1947 52.4337
R19001 vdd.n1943 vdd.n1900 52.4337
R19002 vdd.n1941 vdd.n1940 52.4337
R19003 vdd.n1936 vdd.n1907 52.4337
R19004 vdd.n1934 vdd.n1933 52.4337
R19005 vdd.n1929 vdd.n1915 52.4337
R19006 vdd.n1927 vdd.n1926 52.4337
R19007 vdd.n1922 vdd.n1921 52.4337
R19008 vdd.n1917 vdd.n1916 52.4337
R19009 vdd.n2248 vdd.n1041 52.4337
R19010 vdd.n1373 vdd.n1372 52.4337
R19011 vdd.n1187 vdd.n1152 52.4337
R19012 vdd.n1189 vdd.n1153 52.4337
R19013 vdd.n1193 vdd.n1154 52.4337
R19014 vdd.n1195 vdd.n1155 52.4337
R19015 vdd.n1199 vdd.n1156 52.4337
R19016 vdd.n1201 vdd.n1157 52.4337
R19017 vdd.n1205 vdd.n1158 52.4337
R19018 vdd.n1207 vdd.n1159 52.4337
R19019 vdd.n1339 vdd.n1160 52.4337
R19020 vdd.n1211 vdd.n1161 52.4337
R19021 vdd.n1215 vdd.n1162 52.4337
R19022 vdd.n1217 vdd.n1163 52.4337
R19023 vdd.n1221 vdd.n1164 52.4337
R19024 vdd.n1223 vdd.n1165 52.4337
R19025 vdd.n1227 vdd.n1166 52.4337
R19026 vdd.n1229 vdd.n1167 52.4337
R19027 vdd.n1233 vdd.n1168 52.4337
R19028 vdd.n1235 vdd.n1169 52.4337
R19029 vdd.n1239 vdd.n1170 52.4337
R19030 vdd.n1303 vdd.n1171 52.4337
R19031 vdd.n1244 vdd.n1172 52.4337
R19032 vdd.n1246 vdd.n1173 52.4337
R19033 vdd.n1250 vdd.n1174 52.4337
R19034 vdd.n1252 vdd.n1175 52.4337
R19035 vdd.n1256 vdd.n1176 52.4337
R19036 vdd.n1258 vdd.n1177 52.4337
R19037 vdd.n1262 vdd.n1178 52.4337
R19038 vdd.n1264 vdd.n1179 52.4337
R19039 vdd.n1268 vdd.n1180 52.4337
R19040 vdd.n1270 vdd.n1181 52.4337
R19041 vdd.n1373 vdd.n1183 52.4337
R19042 vdd.n1188 vdd.n1152 52.4337
R19043 vdd.n1192 vdd.n1153 52.4337
R19044 vdd.n1194 vdd.n1154 52.4337
R19045 vdd.n1198 vdd.n1155 52.4337
R19046 vdd.n1200 vdd.n1156 52.4337
R19047 vdd.n1204 vdd.n1157 52.4337
R19048 vdd.n1206 vdd.n1158 52.4337
R19049 vdd.n1338 vdd.n1159 52.4337
R19050 vdd.n1210 vdd.n1160 52.4337
R19051 vdd.n1214 vdd.n1161 52.4337
R19052 vdd.n1216 vdd.n1162 52.4337
R19053 vdd.n1220 vdd.n1163 52.4337
R19054 vdd.n1222 vdd.n1164 52.4337
R19055 vdd.n1226 vdd.n1165 52.4337
R19056 vdd.n1228 vdd.n1166 52.4337
R19057 vdd.n1232 vdd.n1167 52.4337
R19058 vdd.n1234 vdd.n1168 52.4337
R19059 vdd.n1238 vdd.n1169 52.4337
R19060 vdd.n1240 vdd.n1170 52.4337
R19061 vdd.n1243 vdd.n1171 52.4337
R19062 vdd.n1245 vdd.n1172 52.4337
R19063 vdd.n1249 vdd.n1173 52.4337
R19064 vdd.n1251 vdd.n1174 52.4337
R19065 vdd.n1255 vdd.n1175 52.4337
R19066 vdd.n1257 vdd.n1176 52.4337
R19067 vdd.n1261 vdd.n1177 52.4337
R19068 vdd.n1263 vdd.n1178 52.4337
R19069 vdd.n1267 vdd.n1179 52.4337
R19070 vdd.n1269 vdd.n1180 52.4337
R19071 vdd.n1181 vdd.n1151 52.4337
R19072 vdd.n1041 vdd.n1040 52.4337
R19073 vdd.n1918 vdd.n1917 52.4337
R19074 vdd.n1923 vdd.n1922 52.4337
R19075 vdd.n1928 vdd.n1927 52.4337
R19076 vdd.n1915 vdd.n1908 52.4337
R19077 vdd.n1935 vdd.n1934 52.4337
R19078 vdd.n1907 vdd.n1901 52.4337
R19079 vdd.n1942 vdd.n1941 52.4337
R19080 vdd.n1900 vdd.n1895 52.4337
R19081 vdd.n1949 vdd.n1948 52.4337
R19082 vdd.n1894 vdd.n1893 52.4337
R19083 vdd.n1889 vdd.n1882 52.4337
R19084 vdd.n1960 vdd.n1959 52.4337
R19085 vdd.n1881 vdd.n1875 52.4337
R19086 vdd.n1967 vdd.n1966 52.4337
R19087 vdd.n1874 vdd.n1868 52.4337
R19088 vdd.n1974 vdd.n1973 52.4337
R19089 vdd.n1867 vdd.n1861 52.4337
R19090 vdd.n1981 vdd.n1980 52.4337
R19091 vdd.n1860 vdd.n1855 52.4337
R19092 vdd.n1988 vdd.n1987 52.4337
R19093 vdd.n1854 vdd.n1853 52.4337
R19094 vdd.n1849 vdd.n1842 52.4337
R19095 vdd.n1999 vdd.n1998 52.4337
R19096 vdd.n1841 vdd.n1835 52.4337
R19097 vdd.n2006 vdd.n2005 52.4337
R19098 vdd.n1834 vdd.n1828 52.4337
R19099 vdd.n2013 vdd.n2012 52.4337
R19100 vdd.n2016 vdd.n2015 52.4337
R19101 vdd.n1825 vdd.n1820 52.4337
R19102 vdd.n2238 vdd.n2237 52.4337
R19103 vdd.n1819 vdd.n1047 52.4337
R19104 vdd.n3138 vdd.n3137 52.4337
R19105 vdd.n3132 vdd.n663 52.4337
R19106 vdd.n3128 vdd.n666 52.4337
R19107 vdd.n3126 vdd.n3125 52.4337
R19108 vdd.n3121 vdd.n3120 52.4337
R19109 vdd.n3118 vdd.n3117 52.4337
R19110 vdd.n3113 vdd.n3112 52.4337
R19111 vdd.n3110 vdd.n3109 52.4337
R19112 vdd.n3105 vdd.n3104 52.4337
R19113 vdd.n3102 vdd.n3101 52.4337
R19114 vdd.n3097 vdd.n3096 52.4337
R19115 vdd.n3094 vdd.n3093 52.4337
R19116 vdd.n3089 vdd.n3088 52.4337
R19117 vdd.n3086 vdd.n3085 52.4337
R19118 vdd.n3081 vdd.n3080 52.4337
R19119 vdd.n3078 vdd.n3077 52.4337
R19120 vdd.n3073 vdd.n3072 52.4337
R19121 vdd.n3070 vdd.n3069 52.4337
R19122 vdd.n3065 vdd.n3064 52.4337
R19123 vdd.n3062 vdd.n3061 52.4337
R19124 vdd.n728 vdd.n727 52.4337
R19125 vdd.n3053 vdd.n3052 52.4337
R19126 vdd.n3048 vdd.n729 52.4337
R19127 vdd.n3046 vdd.n3045 52.4337
R19128 vdd.n3041 vdd.n3040 52.4337
R19129 vdd.n3038 vdd.n3037 52.4337
R19130 vdd.n3033 vdd.n3032 52.4337
R19131 vdd.n3030 vdd.n3029 52.4337
R19132 vdd.n3025 vdd.n3024 52.4337
R19133 vdd.n3020 vdd.n750 52.4337
R19134 vdd.n3016 vdd.n752 52.4337
R19135 vdd.n3252 vdd.n404 52.4337
R19136 vdd.n595 vdd.n403 52.4337
R19137 vdd.n589 vdd.n402 52.4337
R19138 vdd.n585 vdd.n401 52.4337
R19139 vdd.n579 vdd.n400 52.4337
R19140 vdd.n575 vdd.n399 52.4337
R19141 vdd.n569 vdd.n398 52.4337
R19142 vdd.n565 vdd.n397 52.4337
R19143 vdd.n559 vdd.n396 52.4337
R19144 vdd.n555 vdd.n395 52.4337
R19145 vdd.n549 vdd.n394 52.4337
R19146 vdd.n545 vdd.n393 52.4337
R19147 vdd.n539 vdd.n392 52.4337
R19148 vdd.n535 vdd.n391 52.4337
R19149 vdd.n529 vdd.n390 52.4337
R19150 vdd.n525 vdd.n389 52.4337
R19151 vdd.n519 vdd.n388 52.4337
R19152 vdd.n515 vdd.n387 52.4337
R19153 vdd.n509 vdd.n386 52.4337
R19154 vdd.n505 vdd.n385 52.4337
R19155 vdd.n499 vdd.n384 52.4337
R19156 vdd.n495 vdd.n383 52.4337
R19157 vdd.n489 vdd.n382 52.4337
R19158 vdd.n485 vdd.n381 52.4337
R19159 vdd.n479 vdd.n380 52.4337
R19160 vdd.n475 vdd.n379 52.4337
R19161 vdd.n469 vdd.n378 52.4337
R19162 vdd.n465 vdd.n377 52.4337
R19163 vdd.n459 vdd.n376 52.4337
R19164 vdd.n455 vdd.n375 52.4337
R19165 vdd.n449 vdd.n374 52.4337
R19166 vdd.n445 vdd.n373 52.4337
R19167 vdd.t238 vdd.t252 51.4683
R19168 vdd.n266 vdd.n264 42.0461
R19169 vdd.n168 vdd.n166 42.0461
R19170 vdd.n71 vdd.n69 42.0461
R19171 vdd.n1690 vdd.n1688 42.0461
R19172 vdd.n1592 vdd.n1590 42.0461
R19173 vdd.n1495 vdd.n1493 42.0461
R19174 vdd.n320 vdd.n319 41.6884
R19175 vdd.n222 vdd.n221 41.6884
R19176 vdd.n125 vdd.n124 41.6884
R19177 vdd.n1744 vdd.n1743 41.6884
R19178 vdd.n1646 vdd.n1645 41.6884
R19179 vdd.n1549 vdd.n1548 41.6884
R19180 vdd.n1150 vdd.n1149 41.1157
R19181 vdd.n1306 vdd.n1305 41.1157
R19182 vdd.n1342 vdd.n1341 41.1157
R19183 vdd.n407 vdd.n406 41.1157
R19184 vdd.n547 vdd.n420 41.1157
R19185 vdd.n433 vdd.n432 41.1157
R19186 vdd.n2970 vdd.n2969 39.2114
R19187 vdd.n2967 vdd.n2966 39.2114
R19188 vdd.n2962 vdd.n784 39.2114
R19189 vdd.n2960 vdd.n2959 39.2114
R19190 vdd.n2955 vdd.n787 39.2114
R19191 vdd.n2953 vdd.n2952 39.2114
R19192 vdd.n2948 vdd.n790 39.2114
R19193 vdd.n2946 vdd.n2945 39.2114
R19194 vdd.n2940 vdd.n793 39.2114
R19195 vdd.n2938 vdd.n2937 39.2114
R19196 vdd.n2933 vdd.n796 39.2114
R19197 vdd.n2931 vdd.n2930 39.2114
R19198 vdd.n2926 vdd.n799 39.2114
R19199 vdd.n2924 vdd.n2923 39.2114
R19200 vdd.n2919 vdd.n802 39.2114
R19201 vdd.n2917 vdd.n2916 39.2114
R19202 vdd.n2912 vdd.n2911 39.2114
R19203 vdd.n2773 vdd.n884 39.2114
R19204 vdd.n2768 vdd.n2522 39.2114
R19205 vdd.n2765 vdd.n2523 39.2114
R19206 vdd.n2761 vdd.n2524 39.2114
R19207 vdd.n2757 vdd.n2525 39.2114
R19208 vdd.n2753 vdd.n2526 39.2114
R19209 vdd.n2749 vdd.n2527 39.2114
R19210 vdd.n2745 vdd.n2528 39.2114
R19211 vdd.n2741 vdd.n2529 39.2114
R19212 vdd.n2737 vdd.n2530 39.2114
R19213 vdd.n2733 vdd.n2531 39.2114
R19214 vdd.n2729 vdd.n2532 39.2114
R19215 vdd.n2725 vdd.n2533 39.2114
R19216 vdd.n2721 vdd.n2534 39.2114
R19217 vdd.n2717 vdd.n2535 39.2114
R19218 vdd.n2713 vdd.n2536 39.2114
R19219 vdd.n2708 vdd.n2537 39.2114
R19220 vdd.n2516 vdd.n924 39.2114
R19221 vdd.n2512 vdd.n923 39.2114
R19222 vdd.n2508 vdd.n922 39.2114
R19223 vdd.n2504 vdd.n921 39.2114
R19224 vdd.n2500 vdd.n920 39.2114
R19225 vdd.n2496 vdd.n919 39.2114
R19226 vdd.n2492 vdd.n918 39.2114
R19227 vdd.n2488 vdd.n917 39.2114
R19228 vdd.n2484 vdd.n916 39.2114
R19229 vdd.n2480 vdd.n915 39.2114
R19230 vdd.n2476 vdd.n914 39.2114
R19231 vdd.n2472 vdd.n913 39.2114
R19232 vdd.n2468 vdd.n912 39.2114
R19233 vdd.n2464 vdd.n911 39.2114
R19234 vdd.n2460 vdd.n910 39.2114
R19235 vdd.n2455 vdd.n909 39.2114
R19236 vdd.n2451 vdd.n908 39.2114
R19237 vdd.n2027 vdd.n1019 39.2114
R19238 vdd.n2033 vdd.n2032 39.2114
R19239 vdd.n2036 vdd.n2035 39.2114
R19240 vdd.n2041 vdd.n2040 39.2114
R19241 vdd.n2044 vdd.n2043 39.2114
R19242 vdd.n2049 vdd.n2048 39.2114
R19243 vdd.n2052 vdd.n2051 39.2114
R19244 vdd.n2057 vdd.n2056 39.2114
R19245 vdd.n2228 vdd.n2059 39.2114
R19246 vdd.n2227 vdd.n2226 39.2114
R19247 vdd.n2220 vdd.n2061 39.2114
R19248 vdd.n2219 vdd.n2218 39.2114
R19249 vdd.n2212 vdd.n2063 39.2114
R19250 vdd.n2211 vdd.n2210 39.2114
R19251 vdd.n2204 vdd.n2065 39.2114
R19252 vdd.n2203 vdd.n2202 39.2114
R19253 vdd.n2196 vdd.n2067 39.2114
R19254 vdd.n2889 vdd.n2888 39.2114
R19255 vdd.n2884 vdd.n2856 39.2114
R19256 vdd.n2882 vdd.n2881 39.2114
R19257 vdd.n2877 vdd.n2859 39.2114
R19258 vdd.n2875 vdd.n2874 39.2114
R19259 vdd.n2870 vdd.n2862 39.2114
R19260 vdd.n2868 vdd.n2867 39.2114
R19261 vdd.n2863 vdd.n755 39.2114
R19262 vdd.n3007 vdd.n3006 39.2114
R19263 vdd.n3004 vdd.n3003 39.2114
R19264 vdd.n2999 vdd.n760 39.2114
R19265 vdd.n2997 vdd.n2996 39.2114
R19266 vdd.n2992 vdd.n763 39.2114
R19267 vdd.n2990 vdd.n2989 39.2114
R19268 vdd.n2985 vdd.n766 39.2114
R19269 vdd.n2983 vdd.n2982 39.2114
R19270 vdd.n2978 vdd.n772 39.2114
R19271 vdd.n2775 vdd.n887 39.2114
R19272 vdd.n2538 vdd.n889 39.2114
R19273 vdd.n2564 vdd.n2539 39.2114
R19274 vdd.n2568 vdd.n2540 39.2114
R19275 vdd.n2572 vdd.n2541 39.2114
R19276 vdd.n2576 vdd.n2542 39.2114
R19277 vdd.n2580 vdd.n2543 39.2114
R19278 vdd.n2584 vdd.n2544 39.2114
R19279 vdd.n2588 vdd.n2545 39.2114
R19280 vdd.n2592 vdd.n2546 39.2114
R19281 vdd.n2596 vdd.n2547 39.2114
R19282 vdd.n2600 vdd.n2548 39.2114
R19283 vdd.n2604 vdd.n2549 39.2114
R19284 vdd.n2608 vdd.n2550 39.2114
R19285 vdd.n2612 vdd.n2551 39.2114
R19286 vdd.n2616 vdd.n2552 39.2114
R19287 vdd.n2620 vdd.n2553 39.2114
R19288 vdd.n2776 vdd.n2775 39.2114
R19289 vdd.n2563 vdd.n2538 39.2114
R19290 vdd.n2567 vdd.n2539 39.2114
R19291 vdd.n2571 vdd.n2540 39.2114
R19292 vdd.n2575 vdd.n2541 39.2114
R19293 vdd.n2579 vdd.n2542 39.2114
R19294 vdd.n2583 vdd.n2543 39.2114
R19295 vdd.n2587 vdd.n2544 39.2114
R19296 vdd.n2591 vdd.n2545 39.2114
R19297 vdd.n2595 vdd.n2546 39.2114
R19298 vdd.n2599 vdd.n2547 39.2114
R19299 vdd.n2603 vdd.n2548 39.2114
R19300 vdd.n2607 vdd.n2549 39.2114
R19301 vdd.n2611 vdd.n2550 39.2114
R19302 vdd.n2615 vdd.n2551 39.2114
R19303 vdd.n2619 vdd.n2552 39.2114
R19304 vdd.n2622 vdd.n2553 39.2114
R19305 vdd.n772 vdd.n767 39.2114
R19306 vdd.n2984 vdd.n2983 39.2114
R19307 vdd.n766 vdd.n764 39.2114
R19308 vdd.n2991 vdd.n2990 39.2114
R19309 vdd.n763 vdd.n761 39.2114
R19310 vdd.n2998 vdd.n2997 39.2114
R19311 vdd.n760 vdd.n758 39.2114
R19312 vdd.n3005 vdd.n3004 39.2114
R19313 vdd.n3008 vdd.n3007 39.2114
R19314 vdd.n2864 vdd.n2863 39.2114
R19315 vdd.n2869 vdd.n2868 39.2114
R19316 vdd.n2862 vdd.n2860 39.2114
R19317 vdd.n2876 vdd.n2875 39.2114
R19318 vdd.n2859 vdd.n2857 39.2114
R19319 vdd.n2883 vdd.n2882 39.2114
R19320 vdd.n2856 vdd.n2854 39.2114
R19321 vdd.n2890 vdd.n2889 39.2114
R19322 vdd.n2028 vdd.n2027 39.2114
R19323 vdd.n2034 vdd.n2033 39.2114
R19324 vdd.n2035 vdd.n2024 39.2114
R19325 vdd.n2042 vdd.n2041 39.2114
R19326 vdd.n2043 vdd.n2022 39.2114
R19327 vdd.n2050 vdd.n2049 39.2114
R19328 vdd.n2051 vdd.n2020 39.2114
R19329 vdd.n2058 vdd.n2057 39.2114
R19330 vdd.n2229 vdd.n2228 39.2114
R19331 vdd.n2226 vdd.n2225 39.2114
R19332 vdd.n2221 vdd.n2220 39.2114
R19333 vdd.n2218 vdd.n2217 39.2114
R19334 vdd.n2213 vdd.n2212 39.2114
R19335 vdd.n2210 vdd.n2209 39.2114
R19336 vdd.n2205 vdd.n2204 39.2114
R19337 vdd.n2202 vdd.n2201 39.2114
R19338 vdd.n2197 vdd.n2196 39.2114
R19339 vdd.n2454 vdd.n908 39.2114
R19340 vdd.n2459 vdd.n909 39.2114
R19341 vdd.n2463 vdd.n910 39.2114
R19342 vdd.n2467 vdd.n911 39.2114
R19343 vdd.n2471 vdd.n912 39.2114
R19344 vdd.n2475 vdd.n913 39.2114
R19345 vdd.n2479 vdd.n914 39.2114
R19346 vdd.n2483 vdd.n915 39.2114
R19347 vdd.n2487 vdd.n916 39.2114
R19348 vdd.n2491 vdd.n917 39.2114
R19349 vdd.n2495 vdd.n918 39.2114
R19350 vdd.n2499 vdd.n919 39.2114
R19351 vdd.n2503 vdd.n920 39.2114
R19352 vdd.n2507 vdd.n921 39.2114
R19353 vdd.n2511 vdd.n922 39.2114
R19354 vdd.n2515 vdd.n923 39.2114
R19355 vdd.n926 vdd.n924 39.2114
R19356 vdd.n2773 vdd.n2772 39.2114
R19357 vdd.n2766 vdd.n2522 39.2114
R19358 vdd.n2762 vdd.n2523 39.2114
R19359 vdd.n2758 vdd.n2524 39.2114
R19360 vdd.n2754 vdd.n2525 39.2114
R19361 vdd.n2750 vdd.n2526 39.2114
R19362 vdd.n2746 vdd.n2527 39.2114
R19363 vdd.n2742 vdd.n2528 39.2114
R19364 vdd.n2738 vdd.n2529 39.2114
R19365 vdd.n2734 vdd.n2530 39.2114
R19366 vdd.n2730 vdd.n2531 39.2114
R19367 vdd.n2726 vdd.n2532 39.2114
R19368 vdd.n2722 vdd.n2533 39.2114
R19369 vdd.n2718 vdd.n2534 39.2114
R19370 vdd.n2714 vdd.n2535 39.2114
R19371 vdd.n2709 vdd.n2536 39.2114
R19372 vdd.n2705 vdd.n2537 39.2114
R19373 vdd.n2911 vdd.n803 39.2114
R19374 vdd.n2918 vdd.n2917 39.2114
R19375 vdd.n802 vdd.n800 39.2114
R19376 vdd.n2925 vdd.n2924 39.2114
R19377 vdd.n799 vdd.n797 39.2114
R19378 vdd.n2932 vdd.n2931 39.2114
R19379 vdd.n796 vdd.n794 39.2114
R19380 vdd.n2939 vdd.n2938 39.2114
R19381 vdd.n793 vdd.n791 39.2114
R19382 vdd.n2947 vdd.n2946 39.2114
R19383 vdd.n790 vdd.n788 39.2114
R19384 vdd.n2954 vdd.n2953 39.2114
R19385 vdd.n787 vdd.n785 39.2114
R19386 vdd.n2961 vdd.n2960 39.2114
R19387 vdd.n784 vdd.n782 39.2114
R19388 vdd.n2968 vdd.n2967 39.2114
R19389 vdd.n2971 vdd.n2970 39.2114
R19390 vdd.n934 vdd.n890 39.2114
R19391 vdd.n2443 vdd.n891 39.2114
R19392 vdd.n2439 vdd.n892 39.2114
R19393 vdd.n2435 vdd.n893 39.2114
R19394 vdd.n2431 vdd.n894 39.2114
R19395 vdd.n2427 vdd.n895 39.2114
R19396 vdd.n2423 vdd.n896 39.2114
R19397 vdd.n2419 vdd.n897 39.2114
R19398 vdd.n2415 vdd.n898 39.2114
R19399 vdd.n2411 vdd.n899 39.2114
R19400 vdd.n2407 vdd.n900 39.2114
R19401 vdd.n2403 vdd.n901 39.2114
R19402 vdd.n2399 vdd.n902 39.2114
R19403 vdd.n2395 vdd.n903 39.2114
R19404 vdd.n2391 vdd.n904 39.2114
R19405 vdd.n2387 vdd.n905 39.2114
R19406 vdd.n2383 vdd.n906 39.2114
R19407 vdd.n2286 vdd.n1023 39.2114
R19408 vdd.n2285 vdd.n2284 39.2114
R19409 vdd.n2278 vdd.n1025 39.2114
R19410 vdd.n2277 vdd.n2276 39.2114
R19411 vdd.n2270 vdd.n1027 39.2114
R19412 vdd.n2269 vdd.n2268 39.2114
R19413 vdd.n2262 vdd.n1029 39.2114
R19414 vdd.n2261 vdd.n2260 39.2114
R19415 vdd.n1032 vdd.n1031 39.2114
R19416 vdd.n2102 vdd.n2101 39.2114
R19417 vdd.n2107 vdd.n2106 39.2114
R19418 vdd.n2110 vdd.n2109 39.2114
R19419 vdd.n2115 vdd.n2114 39.2114
R19420 vdd.n2118 vdd.n2117 39.2114
R19421 vdd.n2123 vdd.n2122 39.2114
R19422 vdd.n2126 vdd.n2125 39.2114
R19423 vdd.n2132 vdd.n2131 39.2114
R19424 vdd.n2380 vdd.n906 39.2114
R19425 vdd.n2384 vdd.n905 39.2114
R19426 vdd.n2388 vdd.n904 39.2114
R19427 vdd.n2392 vdd.n903 39.2114
R19428 vdd.n2396 vdd.n902 39.2114
R19429 vdd.n2400 vdd.n901 39.2114
R19430 vdd.n2404 vdd.n900 39.2114
R19431 vdd.n2408 vdd.n899 39.2114
R19432 vdd.n2412 vdd.n898 39.2114
R19433 vdd.n2416 vdd.n897 39.2114
R19434 vdd.n2420 vdd.n896 39.2114
R19435 vdd.n2424 vdd.n895 39.2114
R19436 vdd.n2428 vdd.n894 39.2114
R19437 vdd.n2432 vdd.n893 39.2114
R19438 vdd.n2436 vdd.n892 39.2114
R19439 vdd.n2440 vdd.n891 39.2114
R19440 vdd.n2444 vdd.n890 39.2114
R19441 vdd.n2287 vdd.n2286 39.2114
R19442 vdd.n2284 vdd.n2283 39.2114
R19443 vdd.n2279 vdd.n2278 39.2114
R19444 vdd.n2276 vdd.n2275 39.2114
R19445 vdd.n2271 vdd.n2270 39.2114
R19446 vdd.n2268 vdd.n2267 39.2114
R19447 vdd.n2263 vdd.n2262 39.2114
R19448 vdd.n2260 vdd.n2259 39.2114
R19449 vdd.n1033 vdd.n1032 39.2114
R19450 vdd.n2103 vdd.n2102 39.2114
R19451 vdd.n2108 vdd.n2107 39.2114
R19452 vdd.n2109 vdd.n2099 39.2114
R19453 vdd.n2116 vdd.n2115 39.2114
R19454 vdd.n2117 vdd.n2097 39.2114
R19455 vdd.n2124 vdd.n2123 39.2114
R19456 vdd.n2125 vdd.n2093 39.2114
R19457 vdd.n2133 vdd.n2132 39.2114
R19458 vdd.n2252 vdd.n2251 37.2369
R19459 vdd.n1955 vdd.n1888 37.2369
R19460 vdd.n1994 vdd.n1848 37.2369
R19461 vdd.n3059 vdd.n724 37.2369
R19462 vdd.n688 vdd.n687 37.2369
R19463 vdd.n3015 vdd.n3014 37.2369
R19464 vdd.n2294 vdd.n1018 31.6883
R19465 vdd.n2519 vdd.n927 31.6883
R19466 vdd.n2452 vdd.n930 31.6883
R19467 vdd.n2198 vdd.n2195 31.6883
R19468 vdd.n2706 vdd.n2704 31.6883
R19469 vdd.n2913 vdd.n2910 31.6883
R19470 vdd.n2783 vdd.n883 31.6883
R19471 vdd.n2974 vdd.n2973 31.6883
R19472 vdd.n2893 vdd.n2892 31.6883
R19473 vdd.n2979 vdd.n771 31.6883
R19474 vdd.n2625 vdd.n2624 31.6883
R19475 vdd.n2779 vdd.n2778 31.6883
R19476 vdd.n2290 vdd.n2289 31.6883
R19477 vdd.n2447 vdd.n2446 31.6883
R19478 vdd.n2379 vdd.n2378 31.6883
R19479 vdd.n2136 vdd.n2135 31.6883
R19480 vdd.n2129 vdd.n2095 30.449
R19481 vdd.n938 vdd.n937 30.449
R19482 vdd.n2070 vdd.n2069 30.449
R19483 vdd.n2457 vdd.n929 30.449
R19484 vdd.n2561 vdd.n2560 30.449
R19485 vdd.n806 vdd.n805 30.449
R19486 vdd.n2711 vdd.n2557 30.449
R19487 vdd.n770 vdd.n769 30.449
R19488 vdd.n1380 vdd.n1146 19.3944
R19489 vdd.n1380 vdd.n1136 19.3944
R19490 vdd.n1392 vdd.n1136 19.3944
R19491 vdd.n1392 vdd.n1134 19.3944
R19492 vdd.n1396 vdd.n1134 19.3944
R19493 vdd.n1396 vdd.n1124 19.3944
R19494 vdd.n1409 vdd.n1124 19.3944
R19495 vdd.n1409 vdd.n1122 19.3944
R19496 vdd.n1413 vdd.n1122 19.3944
R19497 vdd.n1413 vdd.n1114 19.3944
R19498 vdd.n1426 vdd.n1114 19.3944
R19499 vdd.n1426 vdd.n1112 19.3944
R19500 vdd.n1430 vdd.n1112 19.3944
R19501 vdd.n1430 vdd.n1101 19.3944
R19502 vdd.n1442 vdd.n1101 19.3944
R19503 vdd.n1442 vdd.n1099 19.3944
R19504 vdd.n1446 vdd.n1099 19.3944
R19505 vdd.n1446 vdd.n1090 19.3944
R19506 vdd.n1754 vdd.n1090 19.3944
R19507 vdd.n1754 vdd.n1088 19.3944
R19508 vdd.n1758 vdd.n1088 19.3944
R19509 vdd.n1758 vdd.n1079 19.3944
R19510 vdd.n1770 vdd.n1079 19.3944
R19511 vdd.n1770 vdd.n1077 19.3944
R19512 vdd.n1774 vdd.n1077 19.3944
R19513 vdd.n1774 vdd.n1067 19.3944
R19514 vdd.n1787 vdd.n1067 19.3944
R19515 vdd.n1787 vdd.n1065 19.3944
R19516 vdd.n1791 vdd.n1065 19.3944
R19517 vdd.n1791 vdd.n1057 19.3944
R19518 vdd.n1804 vdd.n1057 19.3944
R19519 vdd.n1804 vdd.n1054 19.3944
R19520 vdd.n1810 vdd.n1054 19.3944
R19521 vdd.n1810 vdd.n1055 19.3944
R19522 vdd.n1055 vdd.n1043 19.3944
R19523 vdd.n1299 vdd.n1241 19.3944
R19524 vdd.n1299 vdd.n1298 19.3944
R19525 vdd.n1298 vdd.n1297 19.3944
R19526 vdd.n1297 vdd.n1247 19.3944
R19527 vdd.n1293 vdd.n1247 19.3944
R19528 vdd.n1293 vdd.n1292 19.3944
R19529 vdd.n1292 vdd.n1291 19.3944
R19530 vdd.n1291 vdd.n1253 19.3944
R19531 vdd.n1287 vdd.n1253 19.3944
R19532 vdd.n1287 vdd.n1286 19.3944
R19533 vdd.n1286 vdd.n1285 19.3944
R19534 vdd.n1285 vdd.n1259 19.3944
R19535 vdd.n1281 vdd.n1259 19.3944
R19536 vdd.n1281 vdd.n1280 19.3944
R19537 vdd.n1280 vdd.n1279 19.3944
R19538 vdd.n1279 vdd.n1265 19.3944
R19539 vdd.n1275 vdd.n1265 19.3944
R19540 vdd.n1275 vdd.n1274 19.3944
R19541 vdd.n1274 vdd.n1273 19.3944
R19542 vdd.n1273 vdd.n1271 19.3944
R19543 vdd.n1337 vdd.n1336 19.3944
R19544 vdd.n1336 vdd.n1212 19.3944
R19545 vdd.n1332 vdd.n1212 19.3944
R19546 vdd.n1332 vdd.n1331 19.3944
R19547 vdd.n1331 vdd.n1330 19.3944
R19548 vdd.n1330 vdd.n1218 19.3944
R19549 vdd.n1326 vdd.n1218 19.3944
R19550 vdd.n1326 vdd.n1325 19.3944
R19551 vdd.n1325 vdd.n1324 19.3944
R19552 vdd.n1324 vdd.n1224 19.3944
R19553 vdd.n1320 vdd.n1224 19.3944
R19554 vdd.n1320 vdd.n1319 19.3944
R19555 vdd.n1319 vdd.n1318 19.3944
R19556 vdd.n1318 vdd.n1230 19.3944
R19557 vdd.n1314 vdd.n1230 19.3944
R19558 vdd.n1314 vdd.n1313 19.3944
R19559 vdd.n1313 vdd.n1312 19.3944
R19560 vdd.n1312 vdd.n1236 19.3944
R19561 vdd.n1308 vdd.n1236 19.3944
R19562 vdd.n1308 vdd.n1307 19.3944
R19563 vdd.n1371 vdd.n1370 19.3944
R19564 vdd.n1370 vdd.n1185 19.3944
R19565 vdd.n1366 vdd.n1185 19.3944
R19566 vdd.n1366 vdd.n1365 19.3944
R19567 vdd.n1365 vdd.n1364 19.3944
R19568 vdd.n1364 vdd.n1190 19.3944
R19569 vdd.n1360 vdd.n1190 19.3944
R19570 vdd.n1360 vdd.n1359 19.3944
R19571 vdd.n1359 vdd.n1358 19.3944
R19572 vdd.n1358 vdd.n1196 19.3944
R19573 vdd.n1354 vdd.n1196 19.3944
R19574 vdd.n1354 vdd.n1353 19.3944
R19575 vdd.n1353 vdd.n1352 19.3944
R19576 vdd.n1352 vdd.n1202 19.3944
R19577 vdd.n1348 vdd.n1202 19.3944
R19578 vdd.n1348 vdd.n1347 19.3944
R19579 vdd.n1347 vdd.n1346 19.3944
R19580 vdd.n1346 vdd.n1208 19.3944
R19581 vdd.n1951 vdd.n1886 19.3944
R19582 vdd.n1951 vdd.n1892 19.3944
R19583 vdd.n1946 vdd.n1892 19.3944
R19584 vdd.n1946 vdd.n1945 19.3944
R19585 vdd.n1945 vdd.n1944 19.3944
R19586 vdd.n1944 vdd.n1899 19.3944
R19587 vdd.n1939 vdd.n1899 19.3944
R19588 vdd.n1939 vdd.n1938 19.3944
R19589 vdd.n1938 vdd.n1937 19.3944
R19590 vdd.n1937 vdd.n1906 19.3944
R19591 vdd.n1932 vdd.n1906 19.3944
R19592 vdd.n1932 vdd.n1931 19.3944
R19593 vdd.n1931 vdd.n1930 19.3944
R19594 vdd.n1930 vdd.n1914 19.3944
R19595 vdd.n1925 vdd.n1914 19.3944
R19596 vdd.n1925 vdd.n1924 19.3944
R19597 vdd.n1920 vdd.n1919 19.3944
R19598 vdd.n2253 vdd.n1039 19.3944
R19599 vdd.n1990 vdd.n1846 19.3944
R19600 vdd.n1990 vdd.n1852 19.3944
R19601 vdd.n1985 vdd.n1852 19.3944
R19602 vdd.n1985 vdd.n1984 19.3944
R19603 vdd.n1984 vdd.n1983 19.3944
R19604 vdd.n1983 vdd.n1859 19.3944
R19605 vdd.n1978 vdd.n1859 19.3944
R19606 vdd.n1978 vdd.n1977 19.3944
R19607 vdd.n1977 vdd.n1976 19.3944
R19608 vdd.n1976 vdd.n1866 19.3944
R19609 vdd.n1971 vdd.n1866 19.3944
R19610 vdd.n1971 vdd.n1970 19.3944
R19611 vdd.n1970 vdd.n1969 19.3944
R19612 vdd.n1969 vdd.n1873 19.3944
R19613 vdd.n1964 vdd.n1873 19.3944
R19614 vdd.n1964 vdd.n1963 19.3944
R19615 vdd.n1963 vdd.n1962 19.3944
R19616 vdd.n1962 vdd.n1880 19.3944
R19617 vdd.n1957 vdd.n1880 19.3944
R19618 vdd.n1957 vdd.n1956 19.3944
R19619 vdd.n2241 vdd.n2240 19.3944
R19620 vdd.n2240 vdd.n1818 19.3944
R19621 vdd.n2235 vdd.n2234 19.3944
R19622 vdd.n2017 vdd.n1822 19.3944
R19623 vdd.n2017 vdd.n1824 19.3944
R19624 vdd.n1827 vdd.n1824 19.3944
R19625 vdd.n2010 vdd.n1827 19.3944
R19626 vdd.n2010 vdd.n2009 19.3944
R19627 vdd.n2009 vdd.n2008 19.3944
R19628 vdd.n2008 vdd.n1833 19.3944
R19629 vdd.n2003 vdd.n1833 19.3944
R19630 vdd.n2003 vdd.n2002 19.3944
R19631 vdd.n2002 vdd.n2001 19.3944
R19632 vdd.n2001 vdd.n1840 19.3944
R19633 vdd.n1996 vdd.n1840 19.3944
R19634 vdd.n1996 vdd.n1995 19.3944
R19635 vdd.n1384 vdd.n1142 19.3944
R19636 vdd.n1384 vdd.n1140 19.3944
R19637 vdd.n1388 vdd.n1140 19.3944
R19638 vdd.n1388 vdd.n1130 19.3944
R19639 vdd.n1401 vdd.n1130 19.3944
R19640 vdd.n1401 vdd.n1128 19.3944
R19641 vdd.n1405 vdd.n1128 19.3944
R19642 vdd.n1405 vdd.n1119 19.3944
R19643 vdd.n1418 vdd.n1119 19.3944
R19644 vdd.n1418 vdd.n1117 19.3944
R19645 vdd.n1422 vdd.n1117 19.3944
R19646 vdd.n1422 vdd.n1108 19.3944
R19647 vdd.n1434 vdd.n1108 19.3944
R19648 vdd.n1434 vdd.n1106 19.3944
R19649 vdd.n1438 vdd.n1106 19.3944
R19650 vdd.n1438 vdd.n1096 19.3944
R19651 vdd.n1451 vdd.n1096 19.3944
R19652 vdd.n1451 vdd.n1094 19.3944
R19653 vdd.n1750 vdd.n1094 19.3944
R19654 vdd.n1750 vdd.n1085 19.3944
R19655 vdd.n1762 vdd.n1085 19.3944
R19656 vdd.n1762 vdd.n1083 19.3944
R19657 vdd.n1766 vdd.n1083 19.3944
R19658 vdd.n1766 vdd.n1073 19.3944
R19659 vdd.n1779 vdd.n1073 19.3944
R19660 vdd.n1779 vdd.n1071 19.3944
R19661 vdd.n1783 vdd.n1071 19.3944
R19662 vdd.n1783 vdd.n1062 19.3944
R19663 vdd.n1796 vdd.n1062 19.3944
R19664 vdd.n1796 vdd.n1060 19.3944
R19665 vdd.n1800 vdd.n1060 19.3944
R19666 vdd.n1800 vdd.n1050 19.3944
R19667 vdd.n1814 vdd.n1050 19.3944
R19668 vdd.n1814 vdd.n1048 19.3944
R19669 vdd.n2244 vdd.n1048 19.3944
R19670 vdd.n3147 vdd.n655 19.3944
R19671 vdd.n3151 vdd.n655 19.3944
R19672 vdd.n3151 vdd.n646 19.3944
R19673 vdd.n3163 vdd.n646 19.3944
R19674 vdd.n3163 vdd.n644 19.3944
R19675 vdd.n3167 vdd.n644 19.3944
R19676 vdd.n3167 vdd.n633 19.3944
R19677 vdd.n3179 vdd.n633 19.3944
R19678 vdd.n3179 vdd.n631 19.3944
R19679 vdd.n3183 vdd.n631 19.3944
R19680 vdd.n3183 vdd.n622 19.3944
R19681 vdd.n3196 vdd.n622 19.3944
R19682 vdd.n3196 vdd.n620 19.3944
R19683 vdd.n3203 vdd.n620 19.3944
R19684 vdd.n3203 vdd.n3202 19.3944
R19685 vdd.n3202 vdd.n610 19.3944
R19686 vdd.n3216 vdd.n610 19.3944
R19687 vdd.n3217 vdd.n3216 19.3944
R19688 vdd.n3218 vdd.n3217 19.3944
R19689 vdd.n3218 vdd.n608 19.3944
R19690 vdd.n3223 vdd.n608 19.3944
R19691 vdd.n3224 vdd.n3223 19.3944
R19692 vdd.n3225 vdd.n3224 19.3944
R19693 vdd.n3225 vdd.n606 19.3944
R19694 vdd.n3230 vdd.n606 19.3944
R19695 vdd.n3231 vdd.n3230 19.3944
R19696 vdd.n3232 vdd.n3231 19.3944
R19697 vdd.n3232 vdd.n604 19.3944
R19698 vdd.n3238 vdd.n604 19.3944
R19699 vdd.n3239 vdd.n3238 19.3944
R19700 vdd.n3240 vdd.n3239 19.3944
R19701 vdd.n3240 vdd.n602 19.3944
R19702 vdd.n3245 vdd.n602 19.3944
R19703 vdd.n3246 vdd.n3245 19.3944
R19704 vdd.n3247 vdd.n3246 19.3944
R19705 vdd.n550 vdd.n417 19.3944
R19706 vdd.n556 vdd.n417 19.3944
R19707 vdd.n557 vdd.n556 19.3944
R19708 vdd.n560 vdd.n557 19.3944
R19709 vdd.n560 vdd.n415 19.3944
R19710 vdd.n566 vdd.n415 19.3944
R19711 vdd.n567 vdd.n566 19.3944
R19712 vdd.n570 vdd.n567 19.3944
R19713 vdd.n570 vdd.n413 19.3944
R19714 vdd.n576 vdd.n413 19.3944
R19715 vdd.n577 vdd.n576 19.3944
R19716 vdd.n580 vdd.n577 19.3944
R19717 vdd.n580 vdd.n411 19.3944
R19718 vdd.n586 vdd.n411 19.3944
R19719 vdd.n587 vdd.n586 19.3944
R19720 vdd.n590 vdd.n587 19.3944
R19721 vdd.n590 vdd.n409 19.3944
R19722 vdd.n596 vdd.n409 19.3944
R19723 vdd.n598 vdd.n596 19.3944
R19724 vdd.n599 vdd.n598 19.3944
R19725 vdd.n497 vdd.n496 19.3944
R19726 vdd.n500 vdd.n497 19.3944
R19727 vdd.n500 vdd.n429 19.3944
R19728 vdd.n506 vdd.n429 19.3944
R19729 vdd.n507 vdd.n506 19.3944
R19730 vdd.n510 vdd.n507 19.3944
R19731 vdd.n510 vdd.n427 19.3944
R19732 vdd.n516 vdd.n427 19.3944
R19733 vdd.n517 vdd.n516 19.3944
R19734 vdd.n520 vdd.n517 19.3944
R19735 vdd.n520 vdd.n425 19.3944
R19736 vdd.n526 vdd.n425 19.3944
R19737 vdd.n527 vdd.n526 19.3944
R19738 vdd.n530 vdd.n527 19.3944
R19739 vdd.n530 vdd.n423 19.3944
R19740 vdd.n536 vdd.n423 19.3944
R19741 vdd.n537 vdd.n536 19.3944
R19742 vdd.n540 vdd.n537 19.3944
R19743 vdd.n540 vdd.n421 19.3944
R19744 vdd.n546 vdd.n421 19.3944
R19745 vdd.n447 vdd.n446 19.3944
R19746 vdd.n450 vdd.n447 19.3944
R19747 vdd.n450 vdd.n441 19.3944
R19748 vdd.n456 vdd.n441 19.3944
R19749 vdd.n457 vdd.n456 19.3944
R19750 vdd.n460 vdd.n457 19.3944
R19751 vdd.n460 vdd.n439 19.3944
R19752 vdd.n466 vdd.n439 19.3944
R19753 vdd.n467 vdd.n466 19.3944
R19754 vdd.n470 vdd.n467 19.3944
R19755 vdd.n470 vdd.n437 19.3944
R19756 vdd.n476 vdd.n437 19.3944
R19757 vdd.n477 vdd.n476 19.3944
R19758 vdd.n480 vdd.n477 19.3944
R19759 vdd.n480 vdd.n435 19.3944
R19760 vdd.n486 vdd.n435 19.3944
R19761 vdd.n487 vdd.n486 19.3944
R19762 vdd.n490 vdd.n487 19.3944
R19763 vdd.n3143 vdd.n652 19.3944
R19764 vdd.n3155 vdd.n652 19.3944
R19765 vdd.n3155 vdd.n650 19.3944
R19766 vdd.n3159 vdd.n650 19.3944
R19767 vdd.n3159 vdd.n640 19.3944
R19768 vdd.n3171 vdd.n640 19.3944
R19769 vdd.n3171 vdd.n638 19.3944
R19770 vdd.n3175 vdd.n638 19.3944
R19771 vdd.n3175 vdd.n628 19.3944
R19772 vdd.n3188 vdd.n628 19.3944
R19773 vdd.n3188 vdd.n626 19.3944
R19774 vdd.n3192 vdd.n626 19.3944
R19775 vdd.n3192 vdd.n617 19.3944
R19776 vdd.n3207 vdd.n617 19.3944
R19777 vdd.n3207 vdd.n615 19.3944
R19778 vdd.n3211 vdd.n615 19.3944
R19779 vdd.n3211 vdd.n324 19.3944
R19780 vdd.n3289 vdd.n324 19.3944
R19781 vdd.n3289 vdd.n325 19.3944
R19782 vdd.n3283 vdd.n325 19.3944
R19783 vdd.n3283 vdd.n3282 19.3944
R19784 vdd.n3282 vdd.n3281 19.3944
R19785 vdd.n3281 vdd.n337 19.3944
R19786 vdd.n3275 vdd.n337 19.3944
R19787 vdd.n3275 vdd.n3274 19.3944
R19788 vdd.n3274 vdd.n3273 19.3944
R19789 vdd.n3273 vdd.n347 19.3944
R19790 vdd.n3267 vdd.n347 19.3944
R19791 vdd.n3267 vdd.n3266 19.3944
R19792 vdd.n3266 vdd.n3265 19.3944
R19793 vdd.n3265 vdd.n358 19.3944
R19794 vdd.n3259 vdd.n358 19.3944
R19795 vdd.n3259 vdd.n3258 19.3944
R19796 vdd.n3258 vdd.n3257 19.3944
R19797 vdd.n3257 vdd.n369 19.3944
R19798 vdd.n3100 vdd.n3099 19.3944
R19799 vdd.n3099 vdd.n3098 19.3944
R19800 vdd.n3098 vdd.n694 19.3944
R19801 vdd.n3092 vdd.n694 19.3944
R19802 vdd.n3092 vdd.n3091 19.3944
R19803 vdd.n3091 vdd.n3090 19.3944
R19804 vdd.n3090 vdd.n700 19.3944
R19805 vdd.n3084 vdd.n700 19.3944
R19806 vdd.n3084 vdd.n3083 19.3944
R19807 vdd.n3083 vdd.n3082 19.3944
R19808 vdd.n3082 vdd.n706 19.3944
R19809 vdd.n3076 vdd.n706 19.3944
R19810 vdd.n3076 vdd.n3075 19.3944
R19811 vdd.n3075 vdd.n3074 19.3944
R19812 vdd.n3074 vdd.n712 19.3944
R19813 vdd.n3068 vdd.n712 19.3944
R19814 vdd.n3068 vdd.n3067 19.3944
R19815 vdd.n3067 vdd.n3066 19.3944
R19816 vdd.n3066 vdd.n718 19.3944
R19817 vdd.n3060 vdd.n718 19.3944
R19818 vdd.n3140 vdd.n3139 19.3944
R19819 vdd.n3139 vdd.n662 19.3944
R19820 vdd.n3134 vdd.n3133 19.3944
R19821 vdd.n3130 vdd.n3129 19.3944
R19822 vdd.n3129 vdd.n668 19.3944
R19823 vdd.n3124 vdd.n668 19.3944
R19824 vdd.n3124 vdd.n3123 19.3944
R19825 vdd.n3123 vdd.n3122 19.3944
R19826 vdd.n3122 vdd.n674 19.3944
R19827 vdd.n3116 vdd.n674 19.3944
R19828 vdd.n3116 vdd.n3115 19.3944
R19829 vdd.n3115 vdd.n3114 19.3944
R19830 vdd.n3114 vdd.n680 19.3944
R19831 vdd.n3108 vdd.n680 19.3944
R19832 vdd.n3108 vdd.n3107 19.3944
R19833 vdd.n3107 vdd.n3106 19.3944
R19834 vdd.n3055 vdd.n722 19.3944
R19835 vdd.n3055 vdd.n726 19.3944
R19836 vdd.n3050 vdd.n726 19.3944
R19837 vdd.n3050 vdd.n3049 19.3944
R19838 vdd.n3049 vdd.n732 19.3944
R19839 vdd.n3044 vdd.n732 19.3944
R19840 vdd.n3044 vdd.n3043 19.3944
R19841 vdd.n3043 vdd.n3042 19.3944
R19842 vdd.n3042 vdd.n738 19.3944
R19843 vdd.n3036 vdd.n738 19.3944
R19844 vdd.n3036 vdd.n3035 19.3944
R19845 vdd.n3035 vdd.n3034 19.3944
R19846 vdd.n3034 vdd.n744 19.3944
R19847 vdd.n3028 vdd.n744 19.3944
R19848 vdd.n3028 vdd.n3027 19.3944
R19849 vdd.n3027 vdd.n3026 19.3944
R19850 vdd.n3022 vdd.n3021 19.3944
R19851 vdd.n3018 vdd.n3017 19.3944
R19852 vdd.n1306 vdd.n1241 19.0066
R19853 vdd.n1955 vdd.n1886 19.0066
R19854 vdd.n550 vdd.n547 19.0066
R19855 vdd.n3059 vdd.n722 19.0066
R19856 vdd.n1374 vdd.n1144 18.5924
R19857 vdd.n2246 vdd.n1045 18.5924
R19858 vdd.n3145 vdd.n658 18.5924
R19859 vdd.n3254 vdd.n3253 18.5924
R19860 vdd.n2095 vdd.n2094 16.0975
R19861 vdd.n937 vdd.n936 16.0975
R19862 vdd.n1149 vdd.n1148 16.0975
R19863 vdd.n1305 vdd.n1304 16.0975
R19864 vdd.n1341 vdd.n1340 16.0975
R19865 vdd.n2251 vdd.n2250 16.0975
R19866 vdd.n1888 vdd.n1887 16.0975
R19867 vdd.n1848 vdd.n1847 16.0975
R19868 vdd.n2069 vdd.n2068 16.0975
R19869 vdd.n929 vdd.n928 16.0975
R19870 vdd.n2560 vdd.n2559 16.0975
R19871 vdd.n406 vdd.n405 16.0975
R19872 vdd.n420 vdd.n419 16.0975
R19873 vdd.n432 vdd.n431 16.0975
R19874 vdd.n724 vdd.n723 16.0975
R19875 vdd.n687 vdd.n686 16.0975
R19876 vdd.n805 vdd.n804 16.0975
R19877 vdd.n2557 vdd.n2556 16.0975
R19878 vdd.n3014 vdd.n3013 16.0975
R19879 vdd.n769 vdd.n768 16.0975
R19880 vdd.t252 vdd.n2521 15.4182
R19881 vdd.n2774 vdd.t238 15.4182
R19882 vdd.n28 vdd.n27 14.8572
R19883 vdd.n2292 vdd.n1020 14.5112
R19884 vdd.n2976 vdd.n756 14.5112
R19885 vdd.n316 vdd.n281 13.1884
R19886 vdd.n261 vdd.n226 13.1884
R19887 vdd.n218 vdd.n183 13.1884
R19888 vdd.n163 vdd.n128 13.1884
R19889 vdd.n121 vdd.n86 13.1884
R19890 vdd.n66 vdd.n31 13.1884
R19891 vdd.n1685 vdd.n1650 13.1884
R19892 vdd.n1740 vdd.n1705 13.1884
R19893 vdd.n1587 vdd.n1552 13.1884
R19894 vdd.n1642 vdd.n1607 13.1884
R19895 vdd.n1490 vdd.n1455 13.1884
R19896 vdd.n1545 vdd.n1510 13.1884
R19897 vdd.n1342 vdd.n1337 12.9944
R19898 vdd.n1342 vdd.n1208 12.9944
R19899 vdd.n1994 vdd.n1846 12.9944
R19900 vdd.n1995 vdd.n1994 12.9944
R19901 vdd.n496 vdd.n433 12.9944
R19902 vdd.n490 vdd.n433 12.9944
R19903 vdd.n3100 vdd.n688 12.9944
R19904 vdd.n3106 vdd.n688 12.9944
R19905 vdd.n317 vdd.n279 12.8005
R19906 vdd.n312 vdd.n283 12.8005
R19907 vdd.n262 vdd.n224 12.8005
R19908 vdd.n257 vdd.n228 12.8005
R19909 vdd.n219 vdd.n181 12.8005
R19910 vdd.n214 vdd.n185 12.8005
R19911 vdd.n164 vdd.n126 12.8005
R19912 vdd.n159 vdd.n130 12.8005
R19913 vdd.n122 vdd.n84 12.8005
R19914 vdd.n117 vdd.n88 12.8005
R19915 vdd.n67 vdd.n29 12.8005
R19916 vdd.n62 vdd.n33 12.8005
R19917 vdd.n1686 vdd.n1648 12.8005
R19918 vdd.n1681 vdd.n1652 12.8005
R19919 vdd.n1741 vdd.n1703 12.8005
R19920 vdd.n1736 vdd.n1707 12.8005
R19921 vdd.n1588 vdd.n1550 12.8005
R19922 vdd.n1583 vdd.n1554 12.8005
R19923 vdd.n1643 vdd.n1605 12.8005
R19924 vdd.n1638 vdd.n1609 12.8005
R19925 vdd.n1491 vdd.n1453 12.8005
R19926 vdd.n1486 vdd.n1457 12.8005
R19927 vdd.n1546 vdd.n1508 12.8005
R19928 vdd.n1541 vdd.n1512 12.8005
R19929 vdd.n311 vdd.n284 12.0247
R19930 vdd.n256 vdd.n229 12.0247
R19931 vdd.n213 vdd.n186 12.0247
R19932 vdd.n158 vdd.n131 12.0247
R19933 vdd.n116 vdd.n89 12.0247
R19934 vdd.n61 vdd.n34 12.0247
R19935 vdd.n1680 vdd.n1653 12.0247
R19936 vdd.n1735 vdd.n1708 12.0247
R19937 vdd.n1582 vdd.n1555 12.0247
R19938 vdd.n1637 vdd.n1610 12.0247
R19939 vdd.n1485 vdd.n1458 12.0247
R19940 vdd.n1540 vdd.n1513 12.0247
R19941 vdd.n1382 vdd.n1144 11.337
R19942 vdd.n1390 vdd.n1138 11.337
R19943 vdd.n1390 vdd.n1132 11.337
R19944 vdd.n1399 vdd.n1132 11.337
R19945 vdd.n1407 vdd.n1126 11.337
R19946 vdd.n1416 vdd.n1415 11.337
R19947 vdd.n1432 vdd.n1110 11.337
R19948 vdd.n1440 vdd.n1103 11.337
R19949 vdd.n1449 vdd.n1448 11.337
R19950 vdd.n1752 vdd.n1092 11.337
R19951 vdd.n1768 vdd.n1081 11.337
R19952 vdd.n1777 vdd.n1075 11.337
R19953 vdd.n1785 vdd.n1069 11.337
R19954 vdd.n1794 vdd.n1793 11.337
R19955 vdd.n1802 vdd.n1052 11.337
R19956 vdd.n1812 vdd.n1052 11.337
R19957 vdd.n2246 vdd.n1044 11.337
R19958 vdd.n3145 vdd.n659 11.337
R19959 vdd.n3153 vdd.n648 11.337
R19960 vdd.n3161 vdd.n648 11.337
R19961 vdd.n3169 vdd.n642 11.337
R19962 vdd.n3177 vdd.n635 11.337
R19963 vdd.n3186 vdd.n3185 11.337
R19964 vdd.n3194 vdd.n624 11.337
R19965 vdd.n3213 vdd.n613 11.337
R19966 vdd.n3287 vdd.n328 11.337
R19967 vdd.n3285 vdd.n332 11.337
R19968 vdd.n3279 vdd.n3278 11.337
R19969 vdd.n3271 vdd.n349 11.337
R19970 vdd.n3270 vdd.n3269 11.337
R19971 vdd.n3263 vdd.n3262 11.337
R19972 vdd.n3262 vdd.n3261 11.337
R19973 vdd.n3261 vdd.n363 11.337
R19974 vdd.n3255 vdd.n3254 11.337
R19975 vdd.n308 vdd.n307 11.249
R19976 vdd.n253 vdd.n252 11.249
R19977 vdd.n210 vdd.n209 11.249
R19978 vdd.n155 vdd.n154 11.249
R19979 vdd.n113 vdd.n112 11.249
R19980 vdd.n58 vdd.n57 11.249
R19981 vdd.n1677 vdd.n1676 11.249
R19982 vdd.n1732 vdd.n1731 11.249
R19983 vdd.n1579 vdd.n1578 11.249
R19984 vdd.n1634 vdd.n1633 11.249
R19985 vdd.n1482 vdd.n1481 11.249
R19986 vdd.n1537 vdd.n1536 11.249
R19987 vdd.n2449 vdd.t258 11.1103
R19988 vdd.n2781 vdd.t250 11.1103
R19989 vdd.n1802 vdd.t114 10.7702
R19990 vdd.n3161 vdd.t112 10.7702
R19991 vdd.n293 vdd.n292 10.7238
R19992 vdd.n238 vdd.n237 10.7238
R19993 vdd.n195 vdd.n194 10.7238
R19994 vdd.n140 vdd.n139 10.7238
R19995 vdd.n98 vdd.n97 10.7238
R19996 vdd.n43 vdd.n42 10.7238
R19997 vdd.n1662 vdd.n1661 10.7238
R19998 vdd.n1717 vdd.n1716 10.7238
R19999 vdd.n1564 vdd.n1563 10.7238
R20000 vdd.n1619 vdd.n1618 10.7238
R20001 vdd.n1467 vdd.n1466 10.7238
R20002 vdd.n1522 vdd.n1521 10.7238
R20003 vdd.n2295 vdd.n2294 10.6151
R20004 vdd.n2296 vdd.n2295 10.6151
R20005 vdd.n2296 vdd.n1006 10.6151
R20006 vdd.n2306 vdd.n1006 10.6151
R20007 vdd.n2307 vdd.n2306 10.6151
R20008 vdd.n2308 vdd.n2307 10.6151
R20009 vdd.n2308 vdd.n993 10.6151
R20010 vdd.n2319 vdd.n993 10.6151
R20011 vdd.n2320 vdd.n2319 10.6151
R20012 vdd.n2321 vdd.n2320 10.6151
R20013 vdd.n2321 vdd.n981 10.6151
R20014 vdd.n2331 vdd.n981 10.6151
R20015 vdd.n2332 vdd.n2331 10.6151
R20016 vdd.n2333 vdd.n2332 10.6151
R20017 vdd.n2333 vdd.n969 10.6151
R20018 vdd.n2343 vdd.n969 10.6151
R20019 vdd.n2344 vdd.n2343 10.6151
R20020 vdd.n2345 vdd.n2344 10.6151
R20021 vdd.n2345 vdd.n958 10.6151
R20022 vdd.n2355 vdd.n958 10.6151
R20023 vdd.n2356 vdd.n2355 10.6151
R20024 vdd.n2357 vdd.n2356 10.6151
R20025 vdd.n2357 vdd.n945 10.6151
R20026 vdd.n2369 vdd.n945 10.6151
R20027 vdd.n2370 vdd.n2369 10.6151
R20028 vdd.n2372 vdd.n2370 10.6151
R20029 vdd.n2372 vdd.n2371 10.6151
R20030 vdd.n2371 vdd.n927 10.6151
R20031 vdd.n2519 vdd.n2518 10.6151
R20032 vdd.n2518 vdd.n2517 10.6151
R20033 vdd.n2517 vdd.n2514 10.6151
R20034 vdd.n2514 vdd.n2513 10.6151
R20035 vdd.n2513 vdd.n2510 10.6151
R20036 vdd.n2510 vdd.n2509 10.6151
R20037 vdd.n2509 vdd.n2506 10.6151
R20038 vdd.n2506 vdd.n2505 10.6151
R20039 vdd.n2505 vdd.n2502 10.6151
R20040 vdd.n2502 vdd.n2501 10.6151
R20041 vdd.n2501 vdd.n2498 10.6151
R20042 vdd.n2498 vdd.n2497 10.6151
R20043 vdd.n2497 vdd.n2494 10.6151
R20044 vdd.n2494 vdd.n2493 10.6151
R20045 vdd.n2493 vdd.n2490 10.6151
R20046 vdd.n2490 vdd.n2489 10.6151
R20047 vdd.n2489 vdd.n2486 10.6151
R20048 vdd.n2486 vdd.n2485 10.6151
R20049 vdd.n2485 vdd.n2482 10.6151
R20050 vdd.n2482 vdd.n2481 10.6151
R20051 vdd.n2481 vdd.n2478 10.6151
R20052 vdd.n2478 vdd.n2477 10.6151
R20053 vdd.n2477 vdd.n2474 10.6151
R20054 vdd.n2474 vdd.n2473 10.6151
R20055 vdd.n2473 vdd.n2470 10.6151
R20056 vdd.n2470 vdd.n2469 10.6151
R20057 vdd.n2469 vdd.n2466 10.6151
R20058 vdd.n2466 vdd.n2465 10.6151
R20059 vdd.n2465 vdd.n2462 10.6151
R20060 vdd.n2462 vdd.n2461 10.6151
R20061 vdd.n2461 vdd.n2458 10.6151
R20062 vdd.n2456 vdd.n2453 10.6151
R20063 vdd.n2453 vdd.n2452 10.6151
R20064 vdd.n2195 vdd.n2194 10.6151
R20065 vdd.n2194 vdd.n2192 10.6151
R20066 vdd.n2192 vdd.n2191 10.6151
R20067 vdd.n2191 vdd.n2189 10.6151
R20068 vdd.n2189 vdd.n2188 10.6151
R20069 vdd.n2188 vdd.n2186 10.6151
R20070 vdd.n2186 vdd.n2185 10.6151
R20071 vdd.n2185 vdd.n2183 10.6151
R20072 vdd.n2183 vdd.n2182 10.6151
R20073 vdd.n2182 vdd.n2180 10.6151
R20074 vdd.n2180 vdd.n2179 10.6151
R20075 vdd.n2179 vdd.n2177 10.6151
R20076 vdd.n2177 vdd.n2176 10.6151
R20077 vdd.n2176 vdd.n2091 10.6151
R20078 vdd.n2091 vdd.n2090 10.6151
R20079 vdd.n2090 vdd.n2088 10.6151
R20080 vdd.n2088 vdd.n2087 10.6151
R20081 vdd.n2087 vdd.n2085 10.6151
R20082 vdd.n2085 vdd.n2084 10.6151
R20083 vdd.n2084 vdd.n2082 10.6151
R20084 vdd.n2082 vdd.n2081 10.6151
R20085 vdd.n2081 vdd.n2079 10.6151
R20086 vdd.n2079 vdd.n2078 10.6151
R20087 vdd.n2078 vdd.n2076 10.6151
R20088 vdd.n2076 vdd.n2075 10.6151
R20089 vdd.n2075 vdd.n2072 10.6151
R20090 vdd.n2072 vdd.n2071 10.6151
R20091 vdd.n2071 vdd.n930 10.6151
R20092 vdd.n2029 vdd.n1018 10.6151
R20093 vdd.n2030 vdd.n2029 10.6151
R20094 vdd.n2031 vdd.n2030 10.6151
R20095 vdd.n2031 vdd.n2025 10.6151
R20096 vdd.n2037 vdd.n2025 10.6151
R20097 vdd.n2038 vdd.n2037 10.6151
R20098 vdd.n2039 vdd.n2038 10.6151
R20099 vdd.n2039 vdd.n2023 10.6151
R20100 vdd.n2045 vdd.n2023 10.6151
R20101 vdd.n2046 vdd.n2045 10.6151
R20102 vdd.n2047 vdd.n2046 10.6151
R20103 vdd.n2047 vdd.n2021 10.6151
R20104 vdd.n2053 vdd.n2021 10.6151
R20105 vdd.n2054 vdd.n2053 10.6151
R20106 vdd.n2055 vdd.n2054 10.6151
R20107 vdd.n2055 vdd.n2019 10.6151
R20108 vdd.n2231 vdd.n2019 10.6151
R20109 vdd.n2231 vdd.n2230 10.6151
R20110 vdd.n2230 vdd.n2060 10.6151
R20111 vdd.n2224 vdd.n2060 10.6151
R20112 vdd.n2224 vdd.n2223 10.6151
R20113 vdd.n2223 vdd.n2222 10.6151
R20114 vdd.n2222 vdd.n2062 10.6151
R20115 vdd.n2216 vdd.n2062 10.6151
R20116 vdd.n2216 vdd.n2215 10.6151
R20117 vdd.n2215 vdd.n2214 10.6151
R20118 vdd.n2214 vdd.n2064 10.6151
R20119 vdd.n2208 vdd.n2064 10.6151
R20120 vdd.n2208 vdd.n2207 10.6151
R20121 vdd.n2207 vdd.n2206 10.6151
R20122 vdd.n2206 vdd.n2066 10.6151
R20123 vdd.n2200 vdd.n2199 10.6151
R20124 vdd.n2199 vdd.n2198 10.6151
R20125 vdd.n2704 vdd.n2703 10.6151
R20126 vdd.n2703 vdd.n2701 10.6151
R20127 vdd.n2701 vdd.n2700 10.6151
R20128 vdd.n2700 vdd.n2558 10.6151
R20129 vdd.n2647 vdd.n2558 10.6151
R20130 vdd.n2648 vdd.n2647 10.6151
R20131 vdd.n2650 vdd.n2648 10.6151
R20132 vdd.n2651 vdd.n2650 10.6151
R20133 vdd.n2653 vdd.n2651 10.6151
R20134 vdd.n2654 vdd.n2653 10.6151
R20135 vdd.n2656 vdd.n2654 10.6151
R20136 vdd.n2657 vdd.n2656 10.6151
R20137 vdd.n2659 vdd.n2657 10.6151
R20138 vdd.n2660 vdd.n2659 10.6151
R20139 vdd.n2675 vdd.n2660 10.6151
R20140 vdd.n2675 vdd.n2674 10.6151
R20141 vdd.n2674 vdd.n2673 10.6151
R20142 vdd.n2673 vdd.n2671 10.6151
R20143 vdd.n2671 vdd.n2670 10.6151
R20144 vdd.n2670 vdd.n2668 10.6151
R20145 vdd.n2668 vdd.n2667 10.6151
R20146 vdd.n2667 vdd.n2665 10.6151
R20147 vdd.n2665 vdd.n2664 10.6151
R20148 vdd.n2664 vdd.n2662 10.6151
R20149 vdd.n2662 vdd.n2661 10.6151
R20150 vdd.n2661 vdd.n807 10.6151
R20151 vdd.n2909 vdd.n807 10.6151
R20152 vdd.n2910 vdd.n2909 10.6151
R20153 vdd.n2771 vdd.n883 10.6151
R20154 vdd.n2771 vdd.n2770 10.6151
R20155 vdd.n2770 vdd.n2769 10.6151
R20156 vdd.n2769 vdd.n2767 10.6151
R20157 vdd.n2767 vdd.n2764 10.6151
R20158 vdd.n2764 vdd.n2763 10.6151
R20159 vdd.n2763 vdd.n2760 10.6151
R20160 vdd.n2760 vdd.n2759 10.6151
R20161 vdd.n2759 vdd.n2756 10.6151
R20162 vdd.n2756 vdd.n2755 10.6151
R20163 vdd.n2755 vdd.n2752 10.6151
R20164 vdd.n2752 vdd.n2751 10.6151
R20165 vdd.n2751 vdd.n2748 10.6151
R20166 vdd.n2748 vdd.n2747 10.6151
R20167 vdd.n2747 vdd.n2744 10.6151
R20168 vdd.n2744 vdd.n2743 10.6151
R20169 vdd.n2743 vdd.n2740 10.6151
R20170 vdd.n2740 vdd.n2739 10.6151
R20171 vdd.n2739 vdd.n2736 10.6151
R20172 vdd.n2736 vdd.n2735 10.6151
R20173 vdd.n2735 vdd.n2732 10.6151
R20174 vdd.n2732 vdd.n2731 10.6151
R20175 vdd.n2731 vdd.n2728 10.6151
R20176 vdd.n2728 vdd.n2727 10.6151
R20177 vdd.n2727 vdd.n2724 10.6151
R20178 vdd.n2724 vdd.n2723 10.6151
R20179 vdd.n2723 vdd.n2720 10.6151
R20180 vdd.n2720 vdd.n2719 10.6151
R20181 vdd.n2719 vdd.n2716 10.6151
R20182 vdd.n2716 vdd.n2715 10.6151
R20183 vdd.n2715 vdd.n2712 10.6151
R20184 vdd.n2710 vdd.n2707 10.6151
R20185 vdd.n2707 vdd.n2706 10.6151
R20186 vdd.n2784 vdd.n2783 10.6151
R20187 vdd.n2785 vdd.n2784 10.6151
R20188 vdd.n2785 vdd.n873 10.6151
R20189 vdd.n2795 vdd.n873 10.6151
R20190 vdd.n2796 vdd.n2795 10.6151
R20191 vdd.n2797 vdd.n2796 10.6151
R20192 vdd.n2797 vdd.n860 10.6151
R20193 vdd.n2807 vdd.n860 10.6151
R20194 vdd.n2808 vdd.n2807 10.6151
R20195 vdd.n2809 vdd.n2808 10.6151
R20196 vdd.n2809 vdd.n849 10.6151
R20197 vdd.n2819 vdd.n849 10.6151
R20198 vdd.n2820 vdd.n2819 10.6151
R20199 vdd.n2821 vdd.n2820 10.6151
R20200 vdd.n2821 vdd.n837 10.6151
R20201 vdd.n2831 vdd.n837 10.6151
R20202 vdd.n2832 vdd.n2831 10.6151
R20203 vdd.n2833 vdd.n2832 10.6151
R20204 vdd.n2833 vdd.n826 10.6151
R20205 vdd.n2845 vdd.n826 10.6151
R20206 vdd.n2846 vdd.n2845 10.6151
R20207 vdd.n2847 vdd.n2846 10.6151
R20208 vdd.n2847 vdd.n812 10.6151
R20209 vdd.n2902 vdd.n812 10.6151
R20210 vdd.n2903 vdd.n2902 10.6151
R20211 vdd.n2904 vdd.n2903 10.6151
R20212 vdd.n2904 vdd.n779 10.6151
R20213 vdd.n2974 vdd.n779 10.6151
R20214 vdd.n2973 vdd.n2972 10.6151
R20215 vdd.n2972 vdd.n780 10.6151
R20216 vdd.n781 vdd.n780 10.6151
R20217 vdd.n2965 vdd.n781 10.6151
R20218 vdd.n2965 vdd.n2964 10.6151
R20219 vdd.n2964 vdd.n2963 10.6151
R20220 vdd.n2963 vdd.n783 10.6151
R20221 vdd.n2958 vdd.n783 10.6151
R20222 vdd.n2958 vdd.n2957 10.6151
R20223 vdd.n2957 vdd.n2956 10.6151
R20224 vdd.n2956 vdd.n786 10.6151
R20225 vdd.n2951 vdd.n786 10.6151
R20226 vdd.n2951 vdd.n2950 10.6151
R20227 vdd.n2950 vdd.n2949 10.6151
R20228 vdd.n2949 vdd.n789 10.6151
R20229 vdd.n2944 vdd.n789 10.6151
R20230 vdd.n2944 vdd.n2943 10.6151
R20231 vdd.n2943 vdd.n2941 10.6151
R20232 vdd.n2941 vdd.n792 10.6151
R20233 vdd.n2936 vdd.n792 10.6151
R20234 vdd.n2936 vdd.n2935 10.6151
R20235 vdd.n2935 vdd.n2934 10.6151
R20236 vdd.n2934 vdd.n795 10.6151
R20237 vdd.n2929 vdd.n795 10.6151
R20238 vdd.n2929 vdd.n2928 10.6151
R20239 vdd.n2928 vdd.n2927 10.6151
R20240 vdd.n2927 vdd.n798 10.6151
R20241 vdd.n2922 vdd.n798 10.6151
R20242 vdd.n2922 vdd.n2921 10.6151
R20243 vdd.n2921 vdd.n2920 10.6151
R20244 vdd.n2920 vdd.n801 10.6151
R20245 vdd.n2915 vdd.n2914 10.6151
R20246 vdd.n2914 vdd.n2913 10.6151
R20247 vdd.n2892 vdd.n2853 10.6151
R20248 vdd.n2887 vdd.n2853 10.6151
R20249 vdd.n2887 vdd.n2886 10.6151
R20250 vdd.n2886 vdd.n2885 10.6151
R20251 vdd.n2885 vdd.n2855 10.6151
R20252 vdd.n2880 vdd.n2855 10.6151
R20253 vdd.n2880 vdd.n2879 10.6151
R20254 vdd.n2879 vdd.n2878 10.6151
R20255 vdd.n2878 vdd.n2858 10.6151
R20256 vdd.n2873 vdd.n2858 10.6151
R20257 vdd.n2873 vdd.n2872 10.6151
R20258 vdd.n2872 vdd.n2871 10.6151
R20259 vdd.n2871 vdd.n2861 10.6151
R20260 vdd.n2866 vdd.n2861 10.6151
R20261 vdd.n2866 vdd.n2865 10.6151
R20262 vdd.n2865 vdd.n753 10.6151
R20263 vdd.n3009 vdd.n753 10.6151
R20264 vdd.n3009 vdd.n754 10.6151
R20265 vdd.n757 vdd.n754 10.6151
R20266 vdd.n3002 vdd.n757 10.6151
R20267 vdd.n3002 vdd.n3001 10.6151
R20268 vdd.n3001 vdd.n3000 10.6151
R20269 vdd.n3000 vdd.n759 10.6151
R20270 vdd.n2995 vdd.n759 10.6151
R20271 vdd.n2995 vdd.n2994 10.6151
R20272 vdd.n2994 vdd.n2993 10.6151
R20273 vdd.n2993 vdd.n762 10.6151
R20274 vdd.n2988 vdd.n762 10.6151
R20275 vdd.n2988 vdd.n2987 10.6151
R20276 vdd.n2987 vdd.n2986 10.6151
R20277 vdd.n2986 vdd.n765 10.6151
R20278 vdd.n2981 vdd.n2980 10.6151
R20279 vdd.n2980 vdd.n2979 10.6151
R20280 vdd.n2627 vdd.n2625 10.6151
R20281 vdd.n2628 vdd.n2627 10.6151
R20282 vdd.n2696 vdd.n2628 10.6151
R20283 vdd.n2696 vdd.n2695 10.6151
R20284 vdd.n2695 vdd.n2694 10.6151
R20285 vdd.n2694 vdd.n2692 10.6151
R20286 vdd.n2692 vdd.n2691 10.6151
R20287 vdd.n2691 vdd.n2689 10.6151
R20288 vdd.n2689 vdd.n2688 10.6151
R20289 vdd.n2688 vdd.n2686 10.6151
R20290 vdd.n2686 vdd.n2685 10.6151
R20291 vdd.n2685 vdd.n2683 10.6151
R20292 vdd.n2683 vdd.n2682 10.6151
R20293 vdd.n2682 vdd.n2680 10.6151
R20294 vdd.n2680 vdd.n2679 10.6151
R20295 vdd.n2679 vdd.n2645 10.6151
R20296 vdd.n2645 vdd.n2644 10.6151
R20297 vdd.n2644 vdd.n2642 10.6151
R20298 vdd.n2642 vdd.n2641 10.6151
R20299 vdd.n2641 vdd.n2639 10.6151
R20300 vdd.n2639 vdd.n2638 10.6151
R20301 vdd.n2638 vdd.n2636 10.6151
R20302 vdd.n2636 vdd.n2635 10.6151
R20303 vdd.n2635 vdd.n2633 10.6151
R20304 vdd.n2633 vdd.n2632 10.6151
R20305 vdd.n2632 vdd.n2630 10.6151
R20306 vdd.n2630 vdd.n2629 10.6151
R20307 vdd.n2629 vdd.n771 10.6151
R20308 vdd.n2778 vdd.n2777 10.6151
R20309 vdd.n2777 vdd.n888 10.6151
R20310 vdd.n2562 vdd.n888 10.6151
R20311 vdd.n2565 vdd.n2562 10.6151
R20312 vdd.n2566 vdd.n2565 10.6151
R20313 vdd.n2569 vdd.n2566 10.6151
R20314 vdd.n2570 vdd.n2569 10.6151
R20315 vdd.n2573 vdd.n2570 10.6151
R20316 vdd.n2574 vdd.n2573 10.6151
R20317 vdd.n2577 vdd.n2574 10.6151
R20318 vdd.n2578 vdd.n2577 10.6151
R20319 vdd.n2581 vdd.n2578 10.6151
R20320 vdd.n2582 vdd.n2581 10.6151
R20321 vdd.n2585 vdd.n2582 10.6151
R20322 vdd.n2586 vdd.n2585 10.6151
R20323 vdd.n2589 vdd.n2586 10.6151
R20324 vdd.n2590 vdd.n2589 10.6151
R20325 vdd.n2593 vdd.n2590 10.6151
R20326 vdd.n2594 vdd.n2593 10.6151
R20327 vdd.n2597 vdd.n2594 10.6151
R20328 vdd.n2598 vdd.n2597 10.6151
R20329 vdd.n2601 vdd.n2598 10.6151
R20330 vdd.n2602 vdd.n2601 10.6151
R20331 vdd.n2605 vdd.n2602 10.6151
R20332 vdd.n2606 vdd.n2605 10.6151
R20333 vdd.n2609 vdd.n2606 10.6151
R20334 vdd.n2610 vdd.n2609 10.6151
R20335 vdd.n2613 vdd.n2610 10.6151
R20336 vdd.n2614 vdd.n2613 10.6151
R20337 vdd.n2617 vdd.n2614 10.6151
R20338 vdd.n2618 vdd.n2617 10.6151
R20339 vdd.n2623 vdd.n2621 10.6151
R20340 vdd.n2624 vdd.n2623 10.6151
R20341 vdd.n2779 vdd.n878 10.6151
R20342 vdd.n2789 vdd.n878 10.6151
R20343 vdd.n2790 vdd.n2789 10.6151
R20344 vdd.n2791 vdd.n2790 10.6151
R20345 vdd.n2791 vdd.n866 10.6151
R20346 vdd.n2801 vdd.n866 10.6151
R20347 vdd.n2802 vdd.n2801 10.6151
R20348 vdd.n2803 vdd.n2802 10.6151
R20349 vdd.n2803 vdd.n855 10.6151
R20350 vdd.n2813 vdd.n855 10.6151
R20351 vdd.n2814 vdd.n2813 10.6151
R20352 vdd.n2815 vdd.n2814 10.6151
R20353 vdd.n2815 vdd.n843 10.6151
R20354 vdd.n2825 vdd.n843 10.6151
R20355 vdd.n2826 vdd.n2825 10.6151
R20356 vdd.n2827 vdd.n2826 10.6151
R20357 vdd.n2827 vdd.n832 10.6151
R20358 vdd.n2837 vdd.n832 10.6151
R20359 vdd.n2838 vdd.n2837 10.6151
R20360 vdd.n2841 vdd.n2838 10.6151
R20361 vdd.n2851 vdd.n820 10.6151
R20362 vdd.n2852 vdd.n2851 10.6151
R20363 vdd.n2898 vdd.n2852 10.6151
R20364 vdd.n2898 vdd.n2897 10.6151
R20365 vdd.n2897 vdd.n2896 10.6151
R20366 vdd.n2896 vdd.n2895 10.6151
R20367 vdd.n2895 vdd.n2893 10.6151
R20368 vdd.n2290 vdd.n1012 10.6151
R20369 vdd.n2300 vdd.n1012 10.6151
R20370 vdd.n2301 vdd.n2300 10.6151
R20371 vdd.n2302 vdd.n2301 10.6151
R20372 vdd.n2302 vdd.n999 10.6151
R20373 vdd.n2312 vdd.n999 10.6151
R20374 vdd.n2313 vdd.n2312 10.6151
R20375 vdd.n2315 vdd.n987 10.6151
R20376 vdd.n2325 vdd.n987 10.6151
R20377 vdd.n2326 vdd.n2325 10.6151
R20378 vdd.n2327 vdd.n2326 10.6151
R20379 vdd.n2327 vdd.n975 10.6151
R20380 vdd.n2337 vdd.n975 10.6151
R20381 vdd.n2338 vdd.n2337 10.6151
R20382 vdd.n2339 vdd.n2338 10.6151
R20383 vdd.n2339 vdd.n964 10.6151
R20384 vdd.n2349 vdd.n964 10.6151
R20385 vdd.n2350 vdd.n2349 10.6151
R20386 vdd.n2351 vdd.n2350 10.6151
R20387 vdd.n2351 vdd.n952 10.6151
R20388 vdd.n2361 vdd.n952 10.6151
R20389 vdd.n2362 vdd.n2361 10.6151
R20390 vdd.n2365 vdd.n2362 10.6151
R20391 vdd.n2365 vdd.n2364 10.6151
R20392 vdd.n2364 vdd.n2363 10.6151
R20393 vdd.n2363 vdd.n935 10.6151
R20394 vdd.n2447 vdd.n935 10.6151
R20395 vdd.n2446 vdd.n2445 10.6151
R20396 vdd.n2445 vdd.n2442 10.6151
R20397 vdd.n2442 vdd.n2441 10.6151
R20398 vdd.n2441 vdd.n2438 10.6151
R20399 vdd.n2438 vdd.n2437 10.6151
R20400 vdd.n2437 vdd.n2434 10.6151
R20401 vdd.n2434 vdd.n2433 10.6151
R20402 vdd.n2433 vdd.n2430 10.6151
R20403 vdd.n2430 vdd.n2429 10.6151
R20404 vdd.n2429 vdd.n2426 10.6151
R20405 vdd.n2426 vdd.n2425 10.6151
R20406 vdd.n2425 vdd.n2422 10.6151
R20407 vdd.n2422 vdd.n2421 10.6151
R20408 vdd.n2421 vdd.n2418 10.6151
R20409 vdd.n2418 vdd.n2417 10.6151
R20410 vdd.n2417 vdd.n2414 10.6151
R20411 vdd.n2414 vdd.n2413 10.6151
R20412 vdd.n2413 vdd.n2410 10.6151
R20413 vdd.n2410 vdd.n2409 10.6151
R20414 vdd.n2409 vdd.n2406 10.6151
R20415 vdd.n2406 vdd.n2405 10.6151
R20416 vdd.n2405 vdd.n2402 10.6151
R20417 vdd.n2402 vdd.n2401 10.6151
R20418 vdd.n2401 vdd.n2398 10.6151
R20419 vdd.n2398 vdd.n2397 10.6151
R20420 vdd.n2397 vdd.n2394 10.6151
R20421 vdd.n2394 vdd.n2393 10.6151
R20422 vdd.n2393 vdd.n2390 10.6151
R20423 vdd.n2390 vdd.n2389 10.6151
R20424 vdd.n2389 vdd.n2386 10.6151
R20425 vdd.n2386 vdd.n2385 10.6151
R20426 vdd.n2382 vdd.n2381 10.6151
R20427 vdd.n2381 vdd.n2379 10.6151
R20428 vdd.n2138 vdd.n2136 10.6151
R20429 vdd.n2139 vdd.n2138 10.6151
R20430 vdd.n2141 vdd.n2139 10.6151
R20431 vdd.n2142 vdd.n2141 10.6151
R20432 vdd.n2144 vdd.n2142 10.6151
R20433 vdd.n2145 vdd.n2144 10.6151
R20434 vdd.n2147 vdd.n2145 10.6151
R20435 vdd.n2148 vdd.n2147 10.6151
R20436 vdd.n2150 vdd.n2148 10.6151
R20437 vdd.n2151 vdd.n2150 10.6151
R20438 vdd.n2153 vdd.n2151 10.6151
R20439 vdd.n2154 vdd.n2153 10.6151
R20440 vdd.n2172 vdd.n2154 10.6151
R20441 vdd.n2172 vdd.n2171 10.6151
R20442 vdd.n2171 vdd.n2170 10.6151
R20443 vdd.n2170 vdd.n2168 10.6151
R20444 vdd.n2168 vdd.n2167 10.6151
R20445 vdd.n2167 vdd.n2165 10.6151
R20446 vdd.n2165 vdd.n2164 10.6151
R20447 vdd.n2164 vdd.n2162 10.6151
R20448 vdd.n2162 vdd.n2161 10.6151
R20449 vdd.n2161 vdd.n2159 10.6151
R20450 vdd.n2159 vdd.n2158 10.6151
R20451 vdd.n2158 vdd.n2156 10.6151
R20452 vdd.n2156 vdd.n2155 10.6151
R20453 vdd.n2155 vdd.n939 10.6151
R20454 vdd.n2377 vdd.n939 10.6151
R20455 vdd.n2378 vdd.n2377 10.6151
R20456 vdd.n2289 vdd.n2288 10.6151
R20457 vdd.n2288 vdd.n1024 10.6151
R20458 vdd.n2282 vdd.n1024 10.6151
R20459 vdd.n2282 vdd.n2281 10.6151
R20460 vdd.n2281 vdd.n2280 10.6151
R20461 vdd.n2280 vdd.n1026 10.6151
R20462 vdd.n2274 vdd.n1026 10.6151
R20463 vdd.n2274 vdd.n2273 10.6151
R20464 vdd.n2273 vdd.n2272 10.6151
R20465 vdd.n2272 vdd.n1028 10.6151
R20466 vdd.n2266 vdd.n1028 10.6151
R20467 vdd.n2266 vdd.n2265 10.6151
R20468 vdd.n2265 vdd.n2264 10.6151
R20469 vdd.n2264 vdd.n1030 10.6151
R20470 vdd.n2258 vdd.n1030 10.6151
R20471 vdd.n2258 vdd.n2257 10.6151
R20472 vdd.n2257 vdd.n2256 10.6151
R20473 vdd.n2256 vdd.n1034 10.6151
R20474 vdd.n2104 vdd.n1034 10.6151
R20475 vdd.n2105 vdd.n2104 10.6151
R20476 vdd.n2105 vdd.n2100 10.6151
R20477 vdd.n2111 vdd.n2100 10.6151
R20478 vdd.n2112 vdd.n2111 10.6151
R20479 vdd.n2113 vdd.n2112 10.6151
R20480 vdd.n2113 vdd.n2098 10.6151
R20481 vdd.n2119 vdd.n2098 10.6151
R20482 vdd.n2120 vdd.n2119 10.6151
R20483 vdd.n2121 vdd.n2120 10.6151
R20484 vdd.n2121 vdd.n2096 10.6151
R20485 vdd.n2127 vdd.n2096 10.6151
R20486 vdd.n2128 vdd.n2127 10.6151
R20487 vdd.n2130 vdd.n2092 10.6151
R20488 vdd.n2135 vdd.n2092 10.6151
R20489 vdd.t198 vdd.n1776 10.5435
R20490 vdd.n636 vdd.t118 10.5435
R20491 vdd.n304 vdd.n286 10.4732
R20492 vdd.n249 vdd.n231 10.4732
R20493 vdd.n206 vdd.n188 10.4732
R20494 vdd.n151 vdd.n133 10.4732
R20495 vdd.n109 vdd.n91 10.4732
R20496 vdd.n54 vdd.n36 10.4732
R20497 vdd.n1673 vdd.n1655 10.4732
R20498 vdd.n1728 vdd.n1710 10.4732
R20499 vdd.n1575 vdd.n1557 10.4732
R20500 vdd.n1630 vdd.n1612 10.4732
R20501 vdd.n1478 vdd.n1460 10.4732
R20502 vdd.n1533 vdd.n1515 10.4732
R20503 vdd.n1760 vdd.t167 10.3167
R20504 vdd.n3205 vdd.t110 10.3167
R20505 vdd.t124 vdd.n1104 10.09
R20506 vdd.n1812 vdd.t20 10.09
R20507 vdd.n3153 vdd.t5 10.09
R20508 vdd.n3286 vdd.t120 10.09
R20509 vdd.n1424 vdd.t142 9.86327
R20510 vdd.n3277 vdd.t176 9.86327
R20511 vdd.n303 vdd.n288 9.69747
R20512 vdd.n248 vdd.n233 9.69747
R20513 vdd.n205 vdd.n190 9.69747
R20514 vdd.n150 vdd.n135 9.69747
R20515 vdd.n108 vdd.n93 9.69747
R20516 vdd.n53 vdd.n38 9.69747
R20517 vdd.n1672 vdd.n1657 9.69747
R20518 vdd.n1727 vdd.n1712 9.69747
R20519 vdd.n1574 vdd.n1559 9.69747
R20520 vdd.n1629 vdd.n1614 9.69747
R20521 vdd.n1477 vdd.n1462 9.69747
R20522 vdd.n1532 vdd.n1517 9.69747
R20523 vdd.n2232 vdd.n2231 9.67831
R20524 vdd.n2943 vdd.n2942 9.67831
R20525 vdd.n3010 vdd.n3009 9.67831
R20526 vdd.n2256 vdd.n2255 9.67831
R20527 vdd.t122 vdd.n1398 9.63654
R20528 vdd.n3236 vdd.t135 9.63654
R20529 vdd.n319 vdd.n318 9.45567
R20530 vdd.n264 vdd.n263 9.45567
R20531 vdd.n221 vdd.n220 9.45567
R20532 vdd.n166 vdd.n165 9.45567
R20533 vdd.n124 vdd.n123 9.45567
R20534 vdd.n69 vdd.n68 9.45567
R20535 vdd.n1688 vdd.n1687 9.45567
R20536 vdd.n1743 vdd.n1742 9.45567
R20537 vdd.n1590 vdd.n1589 9.45567
R20538 vdd.n1645 vdd.n1644 9.45567
R20539 vdd.n1493 vdd.n1492 9.45567
R20540 vdd.n1548 vdd.n1547 9.45567
R20541 vdd.n1992 vdd.n1846 9.3005
R20542 vdd.n1991 vdd.n1990 9.3005
R20543 vdd.n1852 vdd.n1851 9.3005
R20544 vdd.n1985 vdd.n1856 9.3005
R20545 vdd.n1984 vdd.n1857 9.3005
R20546 vdd.n1983 vdd.n1858 9.3005
R20547 vdd.n1862 vdd.n1859 9.3005
R20548 vdd.n1978 vdd.n1863 9.3005
R20549 vdd.n1977 vdd.n1864 9.3005
R20550 vdd.n1976 vdd.n1865 9.3005
R20551 vdd.n1869 vdd.n1866 9.3005
R20552 vdd.n1971 vdd.n1870 9.3005
R20553 vdd.n1970 vdd.n1871 9.3005
R20554 vdd.n1969 vdd.n1872 9.3005
R20555 vdd.n1876 vdd.n1873 9.3005
R20556 vdd.n1964 vdd.n1877 9.3005
R20557 vdd.n1963 vdd.n1878 9.3005
R20558 vdd.n1962 vdd.n1879 9.3005
R20559 vdd.n1883 vdd.n1880 9.3005
R20560 vdd.n1957 vdd.n1884 9.3005
R20561 vdd.n1956 vdd.n1885 9.3005
R20562 vdd.n1955 vdd.n1954 9.3005
R20563 vdd.n1953 vdd.n1886 9.3005
R20564 vdd.n1952 vdd.n1951 9.3005
R20565 vdd.n1892 vdd.n1891 9.3005
R20566 vdd.n1946 vdd.n1896 9.3005
R20567 vdd.n1945 vdd.n1897 9.3005
R20568 vdd.n1944 vdd.n1898 9.3005
R20569 vdd.n1902 vdd.n1899 9.3005
R20570 vdd.n1939 vdd.n1903 9.3005
R20571 vdd.n1938 vdd.n1904 9.3005
R20572 vdd.n1937 vdd.n1905 9.3005
R20573 vdd.n1909 vdd.n1906 9.3005
R20574 vdd.n1932 vdd.n1910 9.3005
R20575 vdd.n1931 vdd.n1911 9.3005
R20576 vdd.n1930 vdd.n1912 9.3005
R20577 vdd.n1914 vdd.n1913 9.3005
R20578 vdd.n1925 vdd.n1035 9.3005
R20579 vdd.n1994 vdd.n1993 9.3005
R20580 vdd.n2018 vdd.n2017 9.3005
R20581 vdd.n1824 vdd.n1823 9.3005
R20582 vdd.n1829 vdd.n1827 9.3005
R20583 vdd.n2010 vdd.n1830 9.3005
R20584 vdd.n2009 vdd.n1831 9.3005
R20585 vdd.n2008 vdd.n1832 9.3005
R20586 vdd.n1836 vdd.n1833 9.3005
R20587 vdd.n2003 vdd.n1837 9.3005
R20588 vdd.n2002 vdd.n1838 9.3005
R20589 vdd.n2001 vdd.n1839 9.3005
R20590 vdd.n1843 vdd.n1840 9.3005
R20591 vdd.n1996 vdd.n1844 9.3005
R20592 vdd.n1995 vdd.n1845 9.3005
R20593 vdd.n2240 vdd.n1817 9.3005
R20594 vdd.n2242 vdd.n2241 9.3005
R20595 vdd.n1748 vdd.n1094 9.3005
R20596 vdd.n1750 vdd.n1749 9.3005
R20597 vdd.n1085 vdd.n1084 9.3005
R20598 vdd.n1763 vdd.n1762 9.3005
R20599 vdd.n1764 vdd.n1083 9.3005
R20600 vdd.n1766 vdd.n1765 9.3005
R20601 vdd.n1073 vdd.n1072 9.3005
R20602 vdd.n1780 vdd.n1779 9.3005
R20603 vdd.n1781 vdd.n1071 9.3005
R20604 vdd.n1783 vdd.n1782 9.3005
R20605 vdd.n1062 vdd.n1061 9.3005
R20606 vdd.n1797 vdd.n1796 9.3005
R20607 vdd.n1798 vdd.n1060 9.3005
R20608 vdd.n1800 vdd.n1799 9.3005
R20609 vdd.n1050 vdd.n1049 9.3005
R20610 vdd.n1815 vdd.n1814 9.3005
R20611 vdd.n1816 vdd.n1048 9.3005
R20612 vdd.n2244 vdd.n2243 9.3005
R20613 vdd.n295 vdd.n294 9.3005
R20614 vdd.n290 vdd.n289 9.3005
R20615 vdd.n301 vdd.n300 9.3005
R20616 vdd.n303 vdd.n302 9.3005
R20617 vdd.n286 vdd.n285 9.3005
R20618 vdd.n309 vdd.n308 9.3005
R20619 vdd.n311 vdd.n310 9.3005
R20620 vdd.n283 vdd.n280 9.3005
R20621 vdd.n318 vdd.n317 9.3005
R20622 vdd.n240 vdd.n239 9.3005
R20623 vdd.n235 vdd.n234 9.3005
R20624 vdd.n246 vdd.n245 9.3005
R20625 vdd.n248 vdd.n247 9.3005
R20626 vdd.n231 vdd.n230 9.3005
R20627 vdd.n254 vdd.n253 9.3005
R20628 vdd.n256 vdd.n255 9.3005
R20629 vdd.n228 vdd.n225 9.3005
R20630 vdd.n263 vdd.n262 9.3005
R20631 vdd.n197 vdd.n196 9.3005
R20632 vdd.n192 vdd.n191 9.3005
R20633 vdd.n203 vdd.n202 9.3005
R20634 vdd.n205 vdd.n204 9.3005
R20635 vdd.n188 vdd.n187 9.3005
R20636 vdd.n211 vdd.n210 9.3005
R20637 vdd.n213 vdd.n212 9.3005
R20638 vdd.n185 vdd.n182 9.3005
R20639 vdd.n220 vdd.n219 9.3005
R20640 vdd.n142 vdd.n141 9.3005
R20641 vdd.n137 vdd.n136 9.3005
R20642 vdd.n148 vdd.n147 9.3005
R20643 vdd.n150 vdd.n149 9.3005
R20644 vdd.n133 vdd.n132 9.3005
R20645 vdd.n156 vdd.n155 9.3005
R20646 vdd.n158 vdd.n157 9.3005
R20647 vdd.n130 vdd.n127 9.3005
R20648 vdd.n165 vdd.n164 9.3005
R20649 vdd.n100 vdd.n99 9.3005
R20650 vdd.n95 vdd.n94 9.3005
R20651 vdd.n106 vdd.n105 9.3005
R20652 vdd.n108 vdd.n107 9.3005
R20653 vdd.n91 vdd.n90 9.3005
R20654 vdd.n114 vdd.n113 9.3005
R20655 vdd.n116 vdd.n115 9.3005
R20656 vdd.n88 vdd.n85 9.3005
R20657 vdd.n123 vdd.n122 9.3005
R20658 vdd.n45 vdd.n44 9.3005
R20659 vdd.n40 vdd.n39 9.3005
R20660 vdd.n51 vdd.n50 9.3005
R20661 vdd.n53 vdd.n52 9.3005
R20662 vdd.n36 vdd.n35 9.3005
R20663 vdd.n59 vdd.n58 9.3005
R20664 vdd.n61 vdd.n60 9.3005
R20665 vdd.n33 vdd.n30 9.3005
R20666 vdd.n68 vdd.n67 9.3005
R20667 vdd.n3059 vdd.n3058 9.3005
R20668 vdd.n3060 vdd.n721 9.3005
R20669 vdd.n720 vdd.n718 9.3005
R20670 vdd.n3066 vdd.n717 9.3005
R20671 vdd.n3067 vdd.n716 9.3005
R20672 vdd.n3068 vdd.n715 9.3005
R20673 vdd.n714 vdd.n712 9.3005
R20674 vdd.n3074 vdd.n711 9.3005
R20675 vdd.n3075 vdd.n710 9.3005
R20676 vdd.n3076 vdd.n709 9.3005
R20677 vdd.n708 vdd.n706 9.3005
R20678 vdd.n3082 vdd.n705 9.3005
R20679 vdd.n3083 vdd.n704 9.3005
R20680 vdd.n3084 vdd.n703 9.3005
R20681 vdd.n702 vdd.n700 9.3005
R20682 vdd.n3090 vdd.n699 9.3005
R20683 vdd.n3091 vdd.n698 9.3005
R20684 vdd.n3092 vdd.n697 9.3005
R20685 vdd.n696 vdd.n694 9.3005
R20686 vdd.n3098 vdd.n693 9.3005
R20687 vdd.n3099 vdd.n692 9.3005
R20688 vdd.n3100 vdd.n691 9.3005
R20689 vdd.n690 vdd.n688 9.3005
R20690 vdd.n3106 vdd.n685 9.3005
R20691 vdd.n3107 vdd.n684 9.3005
R20692 vdd.n3108 vdd.n683 9.3005
R20693 vdd.n682 vdd.n680 9.3005
R20694 vdd.n3114 vdd.n679 9.3005
R20695 vdd.n3115 vdd.n678 9.3005
R20696 vdd.n3116 vdd.n677 9.3005
R20697 vdd.n676 vdd.n674 9.3005
R20698 vdd.n3122 vdd.n673 9.3005
R20699 vdd.n3123 vdd.n672 9.3005
R20700 vdd.n3124 vdd.n671 9.3005
R20701 vdd.n670 vdd.n668 9.3005
R20702 vdd.n3129 vdd.n667 9.3005
R20703 vdd.n3139 vdd.n661 9.3005
R20704 vdd.n3141 vdd.n3140 9.3005
R20705 vdd.n652 vdd.n651 9.3005
R20706 vdd.n3156 vdd.n3155 9.3005
R20707 vdd.n3157 vdd.n650 9.3005
R20708 vdd.n3159 vdd.n3158 9.3005
R20709 vdd.n640 vdd.n639 9.3005
R20710 vdd.n3172 vdd.n3171 9.3005
R20711 vdd.n3173 vdd.n638 9.3005
R20712 vdd.n3175 vdd.n3174 9.3005
R20713 vdd.n628 vdd.n627 9.3005
R20714 vdd.n3189 vdd.n3188 9.3005
R20715 vdd.n3190 vdd.n626 9.3005
R20716 vdd.n3192 vdd.n3191 9.3005
R20717 vdd.n617 vdd.n616 9.3005
R20718 vdd.n3208 vdd.n3207 9.3005
R20719 vdd.n3209 vdd.n615 9.3005
R20720 vdd.n3211 vdd.n3210 9.3005
R20721 vdd.n324 vdd.n322 9.3005
R20722 vdd.n3143 vdd.n3142 9.3005
R20723 vdd.n3290 vdd.n3289 9.3005
R20724 vdd.n325 vdd.n323 9.3005
R20725 vdd.n3283 vdd.n334 9.3005
R20726 vdd.n3282 vdd.n335 9.3005
R20727 vdd.n3281 vdd.n336 9.3005
R20728 vdd.n343 vdd.n337 9.3005
R20729 vdd.n3275 vdd.n344 9.3005
R20730 vdd.n3274 vdd.n345 9.3005
R20731 vdd.n3273 vdd.n346 9.3005
R20732 vdd.n354 vdd.n347 9.3005
R20733 vdd.n3267 vdd.n355 9.3005
R20734 vdd.n3266 vdd.n356 9.3005
R20735 vdd.n3265 vdd.n357 9.3005
R20736 vdd.n365 vdd.n358 9.3005
R20737 vdd.n3259 vdd.n366 9.3005
R20738 vdd.n3258 vdd.n367 9.3005
R20739 vdd.n3257 vdd.n368 9.3005
R20740 vdd.n443 vdd.n369 9.3005
R20741 vdd.n447 vdd.n442 9.3005
R20742 vdd.n451 vdd.n450 9.3005
R20743 vdd.n452 vdd.n441 9.3005
R20744 vdd.n456 vdd.n453 9.3005
R20745 vdd.n457 vdd.n440 9.3005
R20746 vdd.n461 vdd.n460 9.3005
R20747 vdd.n462 vdd.n439 9.3005
R20748 vdd.n466 vdd.n463 9.3005
R20749 vdd.n467 vdd.n438 9.3005
R20750 vdd.n471 vdd.n470 9.3005
R20751 vdd.n472 vdd.n437 9.3005
R20752 vdd.n476 vdd.n473 9.3005
R20753 vdd.n477 vdd.n436 9.3005
R20754 vdd.n481 vdd.n480 9.3005
R20755 vdd.n482 vdd.n435 9.3005
R20756 vdd.n486 vdd.n483 9.3005
R20757 vdd.n487 vdd.n434 9.3005
R20758 vdd.n491 vdd.n490 9.3005
R20759 vdd.n492 vdd.n433 9.3005
R20760 vdd.n496 vdd.n493 9.3005
R20761 vdd.n497 vdd.n430 9.3005
R20762 vdd.n501 vdd.n500 9.3005
R20763 vdd.n502 vdd.n429 9.3005
R20764 vdd.n506 vdd.n503 9.3005
R20765 vdd.n507 vdd.n428 9.3005
R20766 vdd.n511 vdd.n510 9.3005
R20767 vdd.n512 vdd.n427 9.3005
R20768 vdd.n516 vdd.n513 9.3005
R20769 vdd.n517 vdd.n426 9.3005
R20770 vdd.n521 vdd.n520 9.3005
R20771 vdd.n522 vdd.n425 9.3005
R20772 vdd.n526 vdd.n523 9.3005
R20773 vdd.n527 vdd.n424 9.3005
R20774 vdd.n531 vdd.n530 9.3005
R20775 vdd.n532 vdd.n423 9.3005
R20776 vdd.n536 vdd.n533 9.3005
R20777 vdd.n537 vdd.n422 9.3005
R20778 vdd.n541 vdd.n540 9.3005
R20779 vdd.n542 vdd.n421 9.3005
R20780 vdd.n546 vdd.n543 9.3005
R20781 vdd.n547 vdd.n418 9.3005
R20782 vdd.n551 vdd.n550 9.3005
R20783 vdd.n552 vdd.n417 9.3005
R20784 vdd.n556 vdd.n553 9.3005
R20785 vdd.n557 vdd.n416 9.3005
R20786 vdd.n561 vdd.n560 9.3005
R20787 vdd.n562 vdd.n415 9.3005
R20788 vdd.n566 vdd.n563 9.3005
R20789 vdd.n567 vdd.n414 9.3005
R20790 vdd.n571 vdd.n570 9.3005
R20791 vdd.n572 vdd.n413 9.3005
R20792 vdd.n576 vdd.n573 9.3005
R20793 vdd.n577 vdd.n412 9.3005
R20794 vdd.n581 vdd.n580 9.3005
R20795 vdd.n582 vdd.n411 9.3005
R20796 vdd.n586 vdd.n583 9.3005
R20797 vdd.n587 vdd.n410 9.3005
R20798 vdd.n591 vdd.n590 9.3005
R20799 vdd.n592 vdd.n409 9.3005
R20800 vdd.n596 vdd.n593 9.3005
R20801 vdd.n598 vdd.n408 9.3005
R20802 vdd.n600 vdd.n599 9.3005
R20803 vdd.n3250 vdd.n3249 9.3005
R20804 vdd.n446 vdd.n444 9.3005
R20805 vdd.n3149 vdd.n655 9.3005
R20806 vdd.n3151 vdd.n3150 9.3005
R20807 vdd.n646 vdd.n645 9.3005
R20808 vdd.n3164 vdd.n3163 9.3005
R20809 vdd.n3165 vdd.n644 9.3005
R20810 vdd.n3167 vdd.n3166 9.3005
R20811 vdd.n633 vdd.n632 9.3005
R20812 vdd.n3180 vdd.n3179 9.3005
R20813 vdd.n3181 vdd.n631 9.3005
R20814 vdd.n3183 vdd.n3182 9.3005
R20815 vdd.n622 vdd.n621 9.3005
R20816 vdd.n3197 vdd.n3196 9.3005
R20817 vdd.n3198 vdd.n620 9.3005
R20818 vdd.n3203 vdd.n3199 9.3005
R20819 vdd.n3202 vdd.n3201 9.3005
R20820 vdd.n3200 vdd.n610 9.3005
R20821 vdd.n3216 vdd.n611 9.3005
R20822 vdd.n3217 vdd.n609 9.3005
R20823 vdd.n3219 vdd.n3218 9.3005
R20824 vdd.n3220 vdd.n608 9.3005
R20825 vdd.n3223 vdd.n3221 9.3005
R20826 vdd.n3224 vdd.n607 9.3005
R20827 vdd.n3226 vdd.n3225 9.3005
R20828 vdd.n3227 vdd.n606 9.3005
R20829 vdd.n3230 vdd.n3228 9.3005
R20830 vdd.n3231 vdd.n605 9.3005
R20831 vdd.n3233 vdd.n3232 9.3005
R20832 vdd.n3234 vdd.n604 9.3005
R20833 vdd.n3238 vdd.n3235 9.3005
R20834 vdd.n3239 vdd.n603 9.3005
R20835 vdd.n3241 vdd.n3240 9.3005
R20836 vdd.n3242 vdd.n602 9.3005
R20837 vdd.n3245 vdd.n3243 9.3005
R20838 vdd.n3246 vdd.n601 9.3005
R20839 vdd.n3248 vdd.n3247 9.3005
R20840 vdd.n3148 vdd.n3147 9.3005
R20841 vdd.n3012 vdd.n656 9.3005
R20842 vdd.n3017 vdd.n3011 9.3005
R20843 vdd.n3027 vdd.n748 9.3005
R20844 vdd.n3028 vdd.n747 9.3005
R20845 vdd.n746 vdd.n744 9.3005
R20846 vdd.n3034 vdd.n743 9.3005
R20847 vdd.n3035 vdd.n742 9.3005
R20848 vdd.n3036 vdd.n741 9.3005
R20849 vdd.n740 vdd.n738 9.3005
R20850 vdd.n3042 vdd.n737 9.3005
R20851 vdd.n3043 vdd.n736 9.3005
R20852 vdd.n3044 vdd.n735 9.3005
R20853 vdd.n734 vdd.n732 9.3005
R20854 vdd.n3049 vdd.n731 9.3005
R20855 vdd.n3050 vdd.n730 9.3005
R20856 vdd.n726 vdd.n725 9.3005
R20857 vdd.n3056 vdd.n3055 9.3005
R20858 vdd.n3057 vdd.n722 9.3005
R20859 vdd.n2254 vdd.n2253 9.3005
R20860 vdd.n2249 vdd.n1038 9.3005
R20861 vdd.n1380 vdd.n1379 9.3005
R20862 vdd.n1136 vdd.n1135 9.3005
R20863 vdd.n1393 vdd.n1392 9.3005
R20864 vdd.n1394 vdd.n1134 9.3005
R20865 vdd.n1396 vdd.n1395 9.3005
R20866 vdd.n1124 vdd.n1123 9.3005
R20867 vdd.n1410 vdd.n1409 9.3005
R20868 vdd.n1411 vdd.n1122 9.3005
R20869 vdd.n1413 vdd.n1412 9.3005
R20870 vdd.n1114 vdd.n1113 9.3005
R20871 vdd.n1427 vdd.n1426 9.3005
R20872 vdd.n1428 vdd.n1112 9.3005
R20873 vdd.n1430 vdd.n1429 9.3005
R20874 vdd.n1101 vdd.n1100 9.3005
R20875 vdd.n1443 vdd.n1442 9.3005
R20876 vdd.n1444 vdd.n1099 9.3005
R20877 vdd.n1446 vdd.n1445 9.3005
R20878 vdd.n1090 vdd.n1089 9.3005
R20879 vdd.n1755 vdd.n1754 9.3005
R20880 vdd.n1756 vdd.n1088 9.3005
R20881 vdd.n1758 vdd.n1757 9.3005
R20882 vdd.n1079 vdd.n1078 9.3005
R20883 vdd.n1771 vdd.n1770 9.3005
R20884 vdd.n1772 vdd.n1077 9.3005
R20885 vdd.n1774 vdd.n1773 9.3005
R20886 vdd.n1067 vdd.n1066 9.3005
R20887 vdd.n1788 vdd.n1787 9.3005
R20888 vdd.n1789 vdd.n1065 9.3005
R20889 vdd.n1791 vdd.n1790 9.3005
R20890 vdd.n1057 vdd.n1056 9.3005
R20891 vdd.n1805 vdd.n1804 9.3005
R20892 vdd.n1806 vdd.n1054 9.3005
R20893 vdd.n1810 vdd.n1809 9.3005
R20894 vdd.n1808 vdd.n1055 9.3005
R20895 vdd.n1807 vdd.n1043 9.3005
R20896 vdd.n1378 vdd.n1146 9.3005
R20897 vdd.n1271 vdd.n1147 9.3005
R20898 vdd.n1273 vdd.n1272 9.3005
R20899 vdd.n1274 vdd.n1266 9.3005
R20900 vdd.n1276 vdd.n1275 9.3005
R20901 vdd.n1277 vdd.n1265 9.3005
R20902 vdd.n1279 vdd.n1278 9.3005
R20903 vdd.n1280 vdd.n1260 9.3005
R20904 vdd.n1282 vdd.n1281 9.3005
R20905 vdd.n1283 vdd.n1259 9.3005
R20906 vdd.n1285 vdd.n1284 9.3005
R20907 vdd.n1286 vdd.n1254 9.3005
R20908 vdd.n1288 vdd.n1287 9.3005
R20909 vdd.n1289 vdd.n1253 9.3005
R20910 vdd.n1291 vdd.n1290 9.3005
R20911 vdd.n1292 vdd.n1248 9.3005
R20912 vdd.n1294 vdd.n1293 9.3005
R20913 vdd.n1295 vdd.n1247 9.3005
R20914 vdd.n1297 vdd.n1296 9.3005
R20915 vdd.n1298 vdd.n1242 9.3005
R20916 vdd.n1300 vdd.n1299 9.3005
R20917 vdd.n1301 vdd.n1241 9.3005
R20918 vdd.n1306 vdd.n1302 9.3005
R20919 vdd.n1307 vdd.n1237 9.3005
R20920 vdd.n1309 vdd.n1308 9.3005
R20921 vdd.n1310 vdd.n1236 9.3005
R20922 vdd.n1312 vdd.n1311 9.3005
R20923 vdd.n1313 vdd.n1231 9.3005
R20924 vdd.n1315 vdd.n1314 9.3005
R20925 vdd.n1316 vdd.n1230 9.3005
R20926 vdd.n1318 vdd.n1317 9.3005
R20927 vdd.n1319 vdd.n1225 9.3005
R20928 vdd.n1321 vdd.n1320 9.3005
R20929 vdd.n1322 vdd.n1224 9.3005
R20930 vdd.n1324 vdd.n1323 9.3005
R20931 vdd.n1325 vdd.n1219 9.3005
R20932 vdd.n1327 vdd.n1326 9.3005
R20933 vdd.n1328 vdd.n1218 9.3005
R20934 vdd.n1330 vdd.n1329 9.3005
R20935 vdd.n1331 vdd.n1213 9.3005
R20936 vdd.n1333 vdd.n1332 9.3005
R20937 vdd.n1334 vdd.n1212 9.3005
R20938 vdd.n1336 vdd.n1335 9.3005
R20939 vdd.n1337 vdd.n1209 9.3005
R20940 vdd.n1343 vdd.n1342 9.3005
R20941 vdd.n1344 vdd.n1208 9.3005
R20942 vdd.n1346 vdd.n1345 9.3005
R20943 vdd.n1347 vdd.n1203 9.3005
R20944 vdd.n1349 vdd.n1348 9.3005
R20945 vdd.n1350 vdd.n1202 9.3005
R20946 vdd.n1352 vdd.n1351 9.3005
R20947 vdd.n1353 vdd.n1197 9.3005
R20948 vdd.n1355 vdd.n1354 9.3005
R20949 vdd.n1356 vdd.n1196 9.3005
R20950 vdd.n1358 vdd.n1357 9.3005
R20951 vdd.n1359 vdd.n1191 9.3005
R20952 vdd.n1361 vdd.n1360 9.3005
R20953 vdd.n1362 vdd.n1190 9.3005
R20954 vdd.n1364 vdd.n1363 9.3005
R20955 vdd.n1365 vdd.n1186 9.3005
R20956 vdd.n1367 vdd.n1366 9.3005
R20957 vdd.n1368 vdd.n1185 9.3005
R20958 vdd.n1370 vdd.n1369 9.3005
R20959 vdd.n1371 vdd.n1184 9.3005
R20960 vdd.n1377 vdd.n1376 9.3005
R20961 vdd.n1385 vdd.n1384 9.3005
R20962 vdd.n1386 vdd.n1140 9.3005
R20963 vdd.n1388 vdd.n1387 9.3005
R20964 vdd.n1130 vdd.n1129 9.3005
R20965 vdd.n1402 vdd.n1401 9.3005
R20966 vdd.n1403 vdd.n1128 9.3005
R20967 vdd.n1405 vdd.n1404 9.3005
R20968 vdd.n1119 vdd.n1118 9.3005
R20969 vdd.n1419 vdd.n1418 9.3005
R20970 vdd.n1420 vdd.n1117 9.3005
R20971 vdd.n1422 vdd.n1421 9.3005
R20972 vdd.n1108 vdd.n1107 9.3005
R20973 vdd.n1435 vdd.n1434 9.3005
R20974 vdd.n1436 vdd.n1106 9.3005
R20975 vdd.n1438 vdd.n1437 9.3005
R20976 vdd.n1096 vdd.n1095 9.3005
R20977 vdd.n1452 vdd.n1451 9.3005
R20978 vdd.n1142 vdd.n1141 9.3005
R20979 vdd.n1664 vdd.n1663 9.3005
R20980 vdd.n1659 vdd.n1658 9.3005
R20981 vdd.n1670 vdd.n1669 9.3005
R20982 vdd.n1672 vdd.n1671 9.3005
R20983 vdd.n1655 vdd.n1654 9.3005
R20984 vdd.n1678 vdd.n1677 9.3005
R20985 vdd.n1680 vdd.n1679 9.3005
R20986 vdd.n1652 vdd.n1649 9.3005
R20987 vdd.n1687 vdd.n1686 9.3005
R20988 vdd.n1719 vdd.n1718 9.3005
R20989 vdd.n1714 vdd.n1713 9.3005
R20990 vdd.n1725 vdd.n1724 9.3005
R20991 vdd.n1727 vdd.n1726 9.3005
R20992 vdd.n1710 vdd.n1709 9.3005
R20993 vdd.n1733 vdd.n1732 9.3005
R20994 vdd.n1735 vdd.n1734 9.3005
R20995 vdd.n1707 vdd.n1704 9.3005
R20996 vdd.n1742 vdd.n1741 9.3005
R20997 vdd.n1566 vdd.n1565 9.3005
R20998 vdd.n1561 vdd.n1560 9.3005
R20999 vdd.n1572 vdd.n1571 9.3005
R21000 vdd.n1574 vdd.n1573 9.3005
R21001 vdd.n1557 vdd.n1556 9.3005
R21002 vdd.n1580 vdd.n1579 9.3005
R21003 vdd.n1582 vdd.n1581 9.3005
R21004 vdd.n1554 vdd.n1551 9.3005
R21005 vdd.n1589 vdd.n1588 9.3005
R21006 vdd.n1621 vdd.n1620 9.3005
R21007 vdd.n1616 vdd.n1615 9.3005
R21008 vdd.n1627 vdd.n1626 9.3005
R21009 vdd.n1629 vdd.n1628 9.3005
R21010 vdd.n1612 vdd.n1611 9.3005
R21011 vdd.n1635 vdd.n1634 9.3005
R21012 vdd.n1637 vdd.n1636 9.3005
R21013 vdd.n1609 vdd.n1606 9.3005
R21014 vdd.n1644 vdd.n1643 9.3005
R21015 vdd.n1469 vdd.n1468 9.3005
R21016 vdd.n1464 vdd.n1463 9.3005
R21017 vdd.n1475 vdd.n1474 9.3005
R21018 vdd.n1477 vdd.n1476 9.3005
R21019 vdd.n1460 vdd.n1459 9.3005
R21020 vdd.n1483 vdd.n1482 9.3005
R21021 vdd.n1485 vdd.n1484 9.3005
R21022 vdd.n1457 vdd.n1454 9.3005
R21023 vdd.n1492 vdd.n1491 9.3005
R21024 vdd.n1524 vdd.n1523 9.3005
R21025 vdd.n1519 vdd.n1518 9.3005
R21026 vdd.n1530 vdd.n1529 9.3005
R21027 vdd.n1532 vdd.n1531 9.3005
R21028 vdd.n1515 vdd.n1514 9.3005
R21029 vdd.n1538 vdd.n1537 9.3005
R21030 vdd.n1540 vdd.n1539 9.3005
R21031 vdd.n1512 vdd.n1509 9.3005
R21032 vdd.n1547 vdd.n1546 9.3005
R21033 vdd.n1398 vdd.t184 9.18308
R21034 vdd.n3236 vdd.t128 9.18308
R21035 vdd.n1424 vdd.t132 8.95635
R21036 vdd.t130 vdd.n3277 8.95635
R21037 vdd.n300 vdd.n299 8.92171
R21038 vdd.n245 vdd.n244 8.92171
R21039 vdd.n202 vdd.n201 8.92171
R21040 vdd.n147 vdd.n146 8.92171
R21041 vdd.n105 vdd.n104 8.92171
R21042 vdd.n50 vdd.n49 8.92171
R21043 vdd.n1669 vdd.n1668 8.92171
R21044 vdd.n1724 vdd.n1723 8.92171
R21045 vdd.n1571 vdd.n1570 8.92171
R21046 vdd.n1626 vdd.n1625 8.92171
R21047 vdd.n1474 vdd.n1473 8.92171
R21048 vdd.n1529 vdd.n1528 8.92171
R21049 vdd.n223 vdd.n125 8.81535
R21050 vdd.n1647 vdd.n1549 8.81535
R21051 vdd.n1104 vdd.t187 8.72962
R21052 vdd.t157 vdd.n3286 8.72962
R21053 vdd.n1760 vdd.t116 8.50289
R21054 vdd.n3205 vdd.t200 8.50289
R21055 vdd.n28 vdd.n14 8.42249
R21056 vdd.n1776 vdd.t126 8.27616
R21057 vdd.t173 vdd.n636 8.27616
R21058 vdd.n3292 vdd.n3291 8.16225
R21059 vdd.n1747 vdd.n1746 8.16225
R21060 vdd.n296 vdd.n290 8.14595
R21061 vdd.n241 vdd.n235 8.14595
R21062 vdd.n198 vdd.n192 8.14595
R21063 vdd.n143 vdd.n137 8.14595
R21064 vdd.n101 vdd.n95 8.14595
R21065 vdd.n46 vdd.n40 8.14595
R21066 vdd.n1665 vdd.n1659 8.14595
R21067 vdd.n1720 vdd.n1714 8.14595
R21068 vdd.n1567 vdd.n1561 8.14595
R21069 vdd.n1622 vdd.n1616 8.14595
R21070 vdd.n1470 vdd.n1464 8.14595
R21071 vdd.n1525 vdd.n1519 8.14595
R21072 vdd.n2840 vdd.n820 8.11757
R21073 vdd.n2314 vdd.n2313 8.11757
R21074 vdd.t13 vdd.n1138 7.8227
R21075 vdd.t9 vdd.n363 7.8227
R21076 vdd.n2292 vdd.n1014 7.70933
R21077 vdd.n2298 vdd.n1014 7.70933
R21078 vdd.n2304 vdd.n1008 7.70933
R21079 vdd.n2304 vdd.n1001 7.70933
R21080 vdd.n2310 vdd.n1001 7.70933
R21081 vdd.n2310 vdd.n1004 7.70933
R21082 vdd.n2317 vdd.n989 7.70933
R21083 vdd.n2323 vdd.n989 7.70933
R21084 vdd.n2329 vdd.n983 7.70933
R21085 vdd.n2335 vdd.n979 7.70933
R21086 vdd.n2341 vdd.n973 7.70933
R21087 vdd.n2353 vdd.n960 7.70933
R21088 vdd.n2359 vdd.n954 7.70933
R21089 vdd.n2359 vdd.n947 7.70933
R21090 vdd.n2367 vdd.n947 7.70933
R21091 vdd.n2374 vdd.t262 7.70933
R21092 vdd.n2449 vdd.t262 7.70933
R21093 vdd.n2781 vdd.t248 7.70933
R21094 vdd.n2787 vdd.t248 7.70933
R21095 vdd.n2793 vdd.n868 7.70933
R21096 vdd.n2799 vdd.n868 7.70933
R21097 vdd.n2799 vdd.n871 7.70933
R21098 vdd.n2805 vdd.n864 7.70933
R21099 vdd.n2817 vdd.n851 7.70933
R21100 vdd.n2823 vdd.n845 7.70933
R21101 vdd.n2829 vdd.n841 7.70933
R21102 vdd.n2835 vdd.n828 7.70933
R21103 vdd.n2843 vdd.n828 7.70933
R21104 vdd.n2849 vdd.n822 7.70933
R21105 vdd.n2849 vdd.n814 7.70933
R21106 vdd.n2900 vdd.n814 7.70933
R21107 vdd.n2900 vdd.n817 7.70933
R21108 vdd.n2906 vdd.n774 7.70933
R21109 vdd.n2976 vdd.n774 7.70933
R21110 vdd.n295 vdd.n292 7.3702
R21111 vdd.n240 vdd.n237 7.3702
R21112 vdd.n197 vdd.n194 7.3702
R21113 vdd.n142 vdd.n139 7.3702
R21114 vdd.n100 vdd.n97 7.3702
R21115 vdd.n45 vdd.n42 7.3702
R21116 vdd.n1664 vdd.n1661 7.3702
R21117 vdd.n1719 vdd.n1716 7.3702
R21118 vdd.n1566 vdd.n1563 7.3702
R21119 vdd.n1621 vdd.n1618 7.3702
R21120 vdd.n1469 vdd.n1466 7.3702
R21121 vdd.n1524 vdd.n1521 7.3702
R21122 vdd.n1307 vdd.n1306 6.98232
R21123 vdd.n1956 vdd.n1955 6.98232
R21124 vdd.n547 vdd.n546 6.98232
R21125 vdd.n3060 vdd.n3059 6.98232
R21126 vdd.n1794 vdd.t217 6.91577
R21127 vdd.n3169 vdd.t180 6.91577
R21128 vdd.t147 vdd.n1075 6.68904
R21129 vdd.n3185 vdd.t145 6.68904
R21130 vdd.n1752 vdd.t196 6.46231
R21131 vdd.n3213 vdd.t155 6.46231
R21132 vdd.n3292 vdd.n321 6.32949
R21133 vdd.n1746 vdd.n1745 6.32949
R21134 vdd.t160 vdd.n1103 6.23558
R21135 vdd.t150 vdd.n332 6.23558
R21136 vdd.n1416 vdd.t182 6.00885
R21137 vdd.n2329 vdd.t99 6.00885
R21138 vdd.n2829 vdd.t93 6.00885
R21139 vdd.n3271 vdd.t153 6.00885
R21140 vdd.n1004 vdd.t58 5.89549
R21141 vdd.t27 vdd.n822 5.89549
R21142 vdd.n296 vdd.n295 5.81868
R21143 vdd.n241 vdd.n240 5.81868
R21144 vdd.n198 vdd.n197 5.81868
R21145 vdd.n143 vdd.n142 5.81868
R21146 vdd.n101 vdd.n100 5.81868
R21147 vdd.n46 vdd.n45 5.81868
R21148 vdd.n1665 vdd.n1664 5.81868
R21149 vdd.n1720 vdd.n1719 5.81868
R21150 vdd.n1567 vdd.n1566 5.81868
R21151 vdd.n1622 vdd.n1621 5.81868
R21152 vdd.n1470 vdd.n1469 5.81868
R21153 vdd.n1525 vdd.n1524 5.81868
R21154 vdd.t1 vdd.n1008 5.78212
R21155 vdd.n2073 vdd.t40 5.78212
R21156 vdd.n2698 vdd.t48 5.78212
R21157 vdd.n817 vdd.t44 5.78212
R21158 vdd.n2457 vdd.n2456 5.77611
R21159 vdd.n2200 vdd.n2070 5.77611
R21160 vdd.n2711 vdd.n2710 5.77611
R21161 vdd.n2915 vdd.n806 5.77611
R21162 vdd.n2981 vdd.n770 5.77611
R21163 vdd.n2621 vdd.n2561 5.77611
R21164 vdd.n2382 vdd.n938 5.77611
R21165 vdd.n2130 vdd.n2129 5.77611
R21166 vdd.n1376 vdd.n1150 5.62474
R21167 vdd.n2252 vdd.n2249 5.62474
R21168 vdd.n3250 vdd.n407 5.62474
R21169 vdd.n3015 vdd.n3012 5.62474
R21170 vdd.t100 vdd.n960 5.44203
R21171 vdd.n864 vdd.t260 5.44203
R21172 vdd.n1126 vdd.t182 5.32866
R21173 vdd.t153 vdd.n3270 5.32866
R21174 vdd.n1432 vdd.t160 5.10193
R21175 vdd.t106 vdd.n983 5.10193
R21176 vdd.n973 vdd.t108 5.10193
R21177 vdd.t109 vdd.n851 5.10193
R21178 vdd.n841 vdd.t92 5.10193
R21179 vdd.n3279 vdd.t150 5.10193
R21180 vdd.n299 vdd.n290 5.04292
R21181 vdd.n244 vdd.n235 5.04292
R21182 vdd.n201 vdd.n192 5.04292
R21183 vdd.n146 vdd.n137 5.04292
R21184 vdd.n104 vdd.n95 5.04292
R21185 vdd.n49 vdd.n40 5.04292
R21186 vdd.n1668 vdd.n1659 5.04292
R21187 vdd.n1723 vdd.n1714 5.04292
R21188 vdd.n1570 vdd.n1561 5.04292
R21189 vdd.n1625 vdd.n1616 5.04292
R21190 vdd.n1473 vdd.n1464 5.04292
R21191 vdd.n1528 vdd.n1519 5.04292
R21192 vdd.n1448 vdd.t196 4.8752
R21193 vdd.t107 vdd.t242 4.8752
R21194 vdd.t98 vdd.t254 4.8752
R21195 vdd.t240 vdd.t104 4.8752
R21196 vdd.t94 vdd.t97 4.8752
R21197 vdd.t155 vdd.n328 4.8752
R21198 vdd.n2458 vdd.n2457 4.83952
R21199 vdd.n2070 vdd.n2066 4.83952
R21200 vdd.n2712 vdd.n2711 4.83952
R21201 vdd.n806 vdd.n801 4.83952
R21202 vdd.n770 vdd.n765 4.83952
R21203 vdd.n2618 vdd.n2561 4.83952
R21204 vdd.n2385 vdd.n938 4.83952
R21205 vdd.n2129 vdd.n2128 4.83952
R21206 vdd.n1924 vdd.n1036 4.74817
R21207 vdd.n1919 vdd.n1037 4.74817
R21208 vdd.n1821 vdd.n1818 4.74817
R21209 vdd.n2233 vdd.n1822 4.74817
R21210 vdd.n2235 vdd.n1821 4.74817
R21211 vdd.n2234 vdd.n2233 4.74817
R21212 vdd.n664 vdd.n662 4.74817
R21213 vdd.n3130 vdd.n665 4.74817
R21214 vdd.n3133 vdd.n665 4.74817
R21215 vdd.n3134 vdd.n664 4.74817
R21216 vdd.n3022 vdd.n749 4.74817
R21217 vdd.n3018 vdd.n751 4.74817
R21218 vdd.n3021 vdd.n751 4.74817
R21219 vdd.n3026 vdd.n749 4.74817
R21220 vdd.n1920 vdd.n1036 4.74817
R21221 vdd.n1039 vdd.n1037 4.74817
R21222 vdd.n321 vdd.n320 4.7074
R21223 vdd.n223 vdd.n222 4.7074
R21224 vdd.n1745 vdd.n1744 4.7074
R21225 vdd.n1647 vdd.n1646 4.7074
R21226 vdd.n1768 vdd.t147 4.64847
R21227 vdd.n3194 vdd.t145 4.64847
R21228 vdd.n2335 vdd.t256 4.53511
R21229 vdd.n2823 vdd.t246 4.53511
R21230 vdd.n1069 vdd.t217 4.42174
R21231 vdd.t180 vdd.n635 4.42174
R21232 vdd.n2367 vdd.t244 4.30838
R21233 vdd.n2793 vdd.t102 4.30838
R21234 vdd.n300 vdd.n288 4.26717
R21235 vdd.n245 vdd.n233 4.26717
R21236 vdd.n202 vdd.n190 4.26717
R21237 vdd.n147 vdd.n135 4.26717
R21238 vdd.n105 vdd.n93 4.26717
R21239 vdd.n50 vdd.n38 4.26717
R21240 vdd.n1669 vdd.n1657 4.26717
R21241 vdd.n1724 vdd.n1712 4.26717
R21242 vdd.n1571 vdd.n1559 4.26717
R21243 vdd.n1626 vdd.n1614 4.26717
R21244 vdd.n1474 vdd.n1462 4.26717
R21245 vdd.n1529 vdd.n1517 4.26717
R21246 vdd.n321 vdd.n223 4.10845
R21247 vdd.n1745 vdd.n1647 4.10845
R21248 vdd.n277 vdd.t233 4.06363
R21249 vdd.n277 vdd.t144 4.06363
R21250 vdd.n275 vdd.t165 4.06363
R21251 vdd.n275 vdd.t232 4.06363
R21252 vdd.n273 vdd.t234 4.06363
R21253 vdd.n273 vdd.t164 4.06363
R21254 vdd.n271 vdd.t169 4.06363
R21255 vdd.n271 vdd.t171 4.06363
R21256 vdd.n269 vdd.t210 4.06363
R21257 vdd.n269 vdd.t134 4.06363
R21258 vdd.n267 vdd.t139 4.06363
R21259 vdd.n267 vdd.t189 4.06363
R21260 vdd.n265 vdd.t191 4.06363
R21261 vdd.n265 vdd.t216 4.06363
R21262 vdd.n179 vdd.t222 4.06363
R21263 vdd.n179 vdd.t129 4.06363
R21264 vdd.n177 vdd.t152 4.06363
R21265 vdd.n177 vdd.t221 4.06363
R21266 vdd.n175 vdd.t225 4.06363
R21267 vdd.n175 vdd.t151 4.06363
R21268 vdd.n173 vdd.t156 4.06363
R21269 vdd.n173 vdd.t158 4.06363
R21270 vdd.n171 vdd.t201 4.06363
R21271 vdd.n171 vdd.t111 4.06363
R21272 vdd.n169 vdd.t119 4.06363
R21273 vdd.n169 vdd.t172 4.06363
R21274 vdd.n167 vdd.t181 4.06363
R21275 vdd.n167 vdd.t203 4.06363
R21276 vdd.n82 vdd.t154 4.06363
R21277 vdd.n82 vdd.t219 4.06363
R21278 vdd.n80 vdd.t131 4.06363
R21279 vdd.n80 vdd.t177 4.06363
R21280 vdd.n78 vdd.t121 4.06363
R21281 vdd.n78 vdd.t159 4.06363
R21282 vdd.n76 vdd.t230 4.06363
R21283 vdd.n76 vdd.t208 4.06363
R21284 vdd.n74 vdd.t212 4.06363
R21285 vdd.n74 vdd.t166 4.06363
R21286 vdd.n72 vdd.t235 4.06363
R21287 vdd.n72 vdd.t146 4.06363
R21288 vdd.n70 vdd.t223 4.06363
R21289 vdd.n70 vdd.t174 4.06363
R21290 vdd.n1689 vdd.t141 4.06363
R21291 vdd.n1689 vdd.t229 4.06363
R21292 vdd.n1691 vdd.t226 4.06363
R21293 vdd.n1691 vdd.t209 4.06363
R21294 vdd.n1693 vdd.t186 4.06363
R21295 vdd.n1693 vdd.t138 4.06363
R21296 vdd.n1695 vdd.t237 4.06363
R21297 vdd.n1695 vdd.t207 4.06363
R21298 vdd.n1697 vdd.t204 4.06363
R21299 vdd.n1697 vdd.t163 4.06363
R21300 vdd.n1699 vdd.t162 4.06363
R21301 vdd.n1699 vdd.t205 4.06363
R21302 vdd.n1701 vdd.t193 4.06363
R21303 vdd.n1701 vdd.t192 4.06363
R21304 vdd.n1591 vdd.t127 4.06363
R21305 vdd.n1591 vdd.t218 4.06363
R21306 vdd.n1593 vdd.t211 4.06363
R21307 vdd.n1593 vdd.t199 4.06363
R21308 vdd.n1595 vdd.t170 4.06363
R21309 vdd.n1595 vdd.t117 4.06363
R21310 vdd.n1597 vdd.t227 4.06363
R21311 vdd.n1597 vdd.t197 4.06363
R21312 vdd.n1599 vdd.t194 4.06363
R21313 vdd.n1599 vdd.t149 4.06363
R21314 vdd.n1601 vdd.t143 4.06363
R21315 vdd.n1601 vdd.t195 4.06363
R21316 vdd.n1603 vdd.t185 4.06363
R21317 vdd.n1603 vdd.t183 4.06363
R21318 vdd.n1494 vdd.t175 4.06363
R21319 vdd.n1494 vdd.t224 4.06363
R21320 vdd.n1496 vdd.t148 4.06363
R21321 vdd.n1496 vdd.t206 4.06363
R21322 vdd.n1498 vdd.t168 4.06363
R21323 vdd.n1498 vdd.t213 4.06363
R21324 vdd.n1500 vdd.t188 4.06363
R21325 vdd.n1500 vdd.t231 4.06363
R21326 vdd.n1502 vdd.t161 4.06363
R21327 vdd.n1502 vdd.t125 4.06363
R21328 vdd.n1504 vdd.t178 4.06363
R21329 vdd.n1504 vdd.t133 4.06363
R21330 vdd.n1506 vdd.t220 4.06363
R21331 vdd.n1506 vdd.t236 4.06363
R21332 vdd.n26 vdd.t80 3.9605
R21333 vdd.n26 vdd.t77 3.9605
R21334 vdd.n23 vdd.t76 3.9605
R21335 vdd.n23 vdd.t79 3.9605
R21336 vdd.n21 vdd.t87 3.9605
R21337 vdd.n21 vdd.t78 3.9605
R21338 vdd.n20 vdd.t82 3.9605
R21339 vdd.n20 vdd.t85 3.9605
R21340 vdd.n15 vdd.t91 3.9605
R21341 vdd.n15 vdd.t90 3.9605
R21342 vdd.n16 vdd.t83 3.9605
R21343 vdd.n16 vdd.t89 3.9605
R21344 vdd.n18 vdd.t84 3.9605
R21345 vdd.n18 vdd.t81 3.9605
R21346 vdd.n25 vdd.t88 3.9605
R21347 vdd.n25 vdd.t86 3.9605
R21348 vdd.n7 vdd.t95 3.61217
R21349 vdd.n7 vdd.t247 3.61217
R21350 vdd.n8 vdd.t241 3.61217
R21351 vdd.n8 vdd.t261 3.61217
R21352 vdd.n10 vdd.t249 3.61217
R21353 vdd.n10 vdd.t103 3.61217
R21354 vdd.n12 vdd.t239 3.61217
R21355 vdd.n12 vdd.t251 3.61217
R21356 vdd.n5 vdd.t259 3.61217
R21357 vdd.n5 vdd.t253 3.61217
R21358 vdd.n3 vdd.t245 3.61217
R21359 vdd.n3 vdd.t263 3.61217
R21360 vdd.n1 vdd.t101 3.61217
R21361 vdd.n1 vdd.t255 3.61217
R21362 vdd.n0 vdd.t257 3.61217
R21363 vdd.n0 vdd.t243 3.61217
R21364 vdd.n1382 vdd.t13 3.51482
R21365 vdd.n3255 vdd.t9 3.51482
R21366 vdd.n304 vdd.n303 3.49141
R21367 vdd.n249 vdd.n248 3.49141
R21368 vdd.n206 vdd.n205 3.49141
R21369 vdd.n151 vdd.n150 3.49141
R21370 vdd.n109 vdd.n108 3.49141
R21371 vdd.n54 vdd.n53 3.49141
R21372 vdd.n1673 vdd.n1672 3.49141
R21373 vdd.n1728 vdd.n1727 3.49141
R21374 vdd.n1575 vdd.n1574 3.49141
R21375 vdd.n1630 vdd.n1629 3.49141
R21376 vdd.n1478 vdd.n1477 3.49141
R21377 vdd.n1533 vdd.n1532 3.49141
R21378 vdd.n2073 vdd.t244 3.40145
R21379 vdd.n2521 vdd.t258 3.40145
R21380 vdd.n2774 vdd.t250 3.40145
R21381 vdd.n2698 vdd.t102 3.40145
R21382 vdd.n2174 vdd.t256 3.17472
R21383 vdd.n2677 vdd.t246 3.17472
R21384 vdd.n1785 vdd.t126 3.06136
R21385 vdd.n3177 vdd.t173 3.06136
R21386 vdd.t116 vdd.n1081 2.83463
R21387 vdd.n624 vdd.t200 2.83463
R21388 vdd.n307 vdd.n286 2.71565
R21389 vdd.n252 vdd.n231 2.71565
R21390 vdd.n209 vdd.n188 2.71565
R21391 vdd.n154 vdd.n133 2.71565
R21392 vdd.n112 vdd.n91 2.71565
R21393 vdd.n57 vdd.n36 2.71565
R21394 vdd.n1676 vdd.n1655 2.71565
R21395 vdd.n1731 vdd.n1710 2.71565
R21396 vdd.n1578 vdd.n1557 2.71565
R21397 vdd.n1633 vdd.n1612 2.71565
R21398 vdd.n1481 vdd.n1460 2.71565
R21399 vdd.n1536 vdd.n1515 2.71565
R21400 vdd.n1449 vdd.t187 2.6079
R21401 vdd.n2323 vdd.t106 2.6079
R21402 vdd.n2347 vdd.t108 2.6079
R21403 vdd.n2811 vdd.t109 2.6079
R21404 vdd.n2835 vdd.t92 2.6079
R21405 vdd.n3287 vdd.t157 2.6079
R21406 vdd.n2841 vdd.n2840 2.49806
R21407 vdd.n2315 vdd.n2314 2.49806
R21408 vdd.n294 vdd.n293 2.4129
R21409 vdd.n239 vdd.n238 2.4129
R21410 vdd.n196 vdd.n195 2.4129
R21411 vdd.n141 vdd.n140 2.4129
R21412 vdd.n99 vdd.n98 2.4129
R21413 vdd.n44 vdd.n43 2.4129
R21414 vdd.n1663 vdd.n1662 2.4129
R21415 vdd.n1718 vdd.n1717 2.4129
R21416 vdd.n1565 vdd.n1564 2.4129
R21417 vdd.n1620 vdd.n1619 2.4129
R21418 vdd.n1468 vdd.n1467 2.4129
R21419 vdd.n1523 vdd.n1522 2.4129
R21420 vdd.t132 vdd.n1110 2.38117
R21421 vdd.n3278 vdd.t130 2.38117
R21422 vdd.n2232 vdd.n1821 2.27742
R21423 vdd.n2233 vdd.n2232 2.27742
R21424 vdd.n2942 vdd.n665 2.27742
R21425 vdd.n2942 vdd.n664 2.27742
R21426 vdd.n3010 vdd.n751 2.27742
R21427 vdd.n3010 vdd.n749 2.27742
R21428 vdd.n2255 vdd.n1036 2.27742
R21429 vdd.n2255 vdd.n1037 2.27742
R21430 vdd.n2347 vdd.t100 2.2678
R21431 vdd.n2811 vdd.t260 2.2678
R21432 vdd.n1407 vdd.t184 2.15444
R21433 vdd.n3269 vdd.t128 2.15444
R21434 vdd.t254 vdd.n954 2.04107
R21435 vdd.n871 vdd.t240 2.04107
R21436 vdd.n308 vdd.n284 1.93989
R21437 vdd.n253 vdd.n229 1.93989
R21438 vdd.n210 vdd.n186 1.93989
R21439 vdd.n155 vdd.n131 1.93989
R21440 vdd.n113 vdd.n89 1.93989
R21441 vdd.n58 vdd.n34 1.93989
R21442 vdd.n1677 vdd.n1653 1.93989
R21443 vdd.n1732 vdd.n1708 1.93989
R21444 vdd.n1579 vdd.n1555 1.93989
R21445 vdd.n1634 vdd.n1610 1.93989
R21446 vdd.n1482 vdd.n1458 1.93989
R21447 vdd.n1537 vdd.n1513 1.93989
R21448 vdd.n2298 vdd.t1 1.92771
R21449 vdd.n2374 vdd.t40 1.92771
R21450 vdd.n2787 vdd.t48 1.92771
R21451 vdd.n2906 vdd.t44 1.92771
R21452 vdd.n1399 vdd.t122 1.70098
R21453 vdd.n2174 vdd.t99 1.70098
R21454 vdd.n979 vdd.t107 1.70098
R21455 vdd.t97 vdd.n845 1.70098
R21456 vdd.n2677 vdd.t93 1.70098
R21457 vdd.n3263 vdd.t135 1.70098
R21458 vdd.n1415 vdd.t142 1.47425
R21459 vdd.n349 vdd.t176 1.47425
R21460 vdd.n1440 vdd.t124 1.24752
R21461 vdd.t20 vdd.n1044 1.24752
R21462 vdd.n659 vdd.t5 1.24752
R21463 vdd.t120 vdd.n3285 1.24752
R21464 vdd.n319 vdd.n279 1.16414
R21465 vdd.n312 vdd.n311 1.16414
R21466 vdd.n264 vdd.n224 1.16414
R21467 vdd.n257 vdd.n256 1.16414
R21468 vdd.n221 vdd.n181 1.16414
R21469 vdd.n214 vdd.n213 1.16414
R21470 vdd.n166 vdd.n126 1.16414
R21471 vdd.n159 vdd.n158 1.16414
R21472 vdd.n124 vdd.n84 1.16414
R21473 vdd.n117 vdd.n116 1.16414
R21474 vdd.n69 vdd.n29 1.16414
R21475 vdd.n62 vdd.n61 1.16414
R21476 vdd.n1688 vdd.n1648 1.16414
R21477 vdd.n1681 vdd.n1680 1.16414
R21478 vdd.n1743 vdd.n1703 1.16414
R21479 vdd.n1736 vdd.n1735 1.16414
R21480 vdd.n1590 vdd.n1550 1.16414
R21481 vdd.n1583 vdd.n1582 1.16414
R21482 vdd.n1645 vdd.n1605 1.16414
R21483 vdd.n1638 vdd.n1637 1.16414
R21484 vdd.n1493 vdd.n1453 1.16414
R21485 vdd.n1486 vdd.n1485 1.16414
R21486 vdd.n1548 vdd.n1508 1.16414
R21487 vdd.n1541 vdd.n1540 1.16414
R21488 vdd.n2341 vdd.t242 1.13415
R21489 vdd.n2817 vdd.t94 1.13415
R21490 vdd.n1092 vdd.t167 1.02079
R21491 vdd.t58 vdd.t105 1.02079
R21492 vdd.t96 vdd.t27 1.02079
R21493 vdd.t110 vdd.n613 1.02079
R21494 vdd.n1271 vdd.n1150 0.970197
R21495 vdd.n2253 vdd.n2252 0.970197
R21496 vdd.n599 vdd.n407 0.970197
R21497 vdd.n3017 vdd.n3015 0.970197
R21498 vdd.n1746 vdd.n28 0.852297
R21499 vdd vdd.n3292 0.844463
R21500 vdd.n1777 vdd.t198 0.794056
R21501 vdd.n2317 vdd.t105 0.794056
R21502 vdd.n2353 vdd.t98 0.794056
R21503 vdd.n2805 vdd.t104 0.794056
R21504 vdd.n2843 vdd.t96 0.794056
R21505 vdd.n3186 vdd.t118 0.794056
R21506 vdd.n1793 vdd.t114 0.567326
R21507 vdd.t112 vdd.n642 0.567326
R21508 vdd.n2243 vdd.n2242 0.482207
R21509 vdd.n3142 vdd.n3141 0.482207
R21510 vdd.n444 vdd.n443 0.482207
R21511 vdd.n3249 vdd.n3248 0.482207
R21512 vdd.n3148 vdd.n656 0.482207
R21513 vdd.n1807 vdd.n1038 0.482207
R21514 vdd.n1378 vdd.n1377 0.482207
R21515 vdd.n1184 vdd.n1141 0.482207
R21516 vdd.n4 vdd.n2 0.459552
R21517 vdd.n11 vdd.n9 0.459552
R21518 vdd.n317 vdd.n316 0.388379
R21519 vdd.n283 vdd.n281 0.388379
R21520 vdd.n262 vdd.n261 0.388379
R21521 vdd.n228 vdd.n226 0.388379
R21522 vdd.n219 vdd.n218 0.388379
R21523 vdd.n185 vdd.n183 0.388379
R21524 vdd.n164 vdd.n163 0.388379
R21525 vdd.n130 vdd.n128 0.388379
R21526 vdd.n122 vdd.n121 0.388379
R21527 vdd.n88 vdd.n86 0.388379
R21528 vdd.n67 vdd.n66 0.388379
R21529 vdd.n33 vdd.n31 0.388379
R21530 vdd.n1686 vdd.n1685 0.388379
R21531 vdd.n1652 vdd.n1650 0.388379
R21532 vdd.n1741 vdd.n1740 0.388379
R21533 vdd.n1707 vdd.n1705 0.388379
R21534 vdd.n1588 vdd.n1587 0.388379
R21535 vdd.n1554 vdd.n1552 0.388379
R21536 vdd.n1643 vdd.n1642 0.388379
R21537 vdd.n1609 vdd.n1607 0.388379
R21538 vdd.n1491 vdd.n1490 0.388379
R21539 vdd.n1457 vdd.n1455 0.388379
R21540 vdd.n1546 vdd.n1545 0.388379
R21541 vdd.n1512 vdd.n1510 0.388379
R21542 vdd.n19 vdd.n17 0.387128
R21543 vdd.n24 vdd.n22 0.387128
R21544 vdd.n6 vdd.n4 0.358259
R21545 vdd.n13 vdd.n11 0.358259
R21546 vdd.n268 vdd.n266 0.358259
R21547 vdd.n270 vdd.n268 0.358259
R21548 vdd.n272 vdd.n270 0.358259
R21549 vdd.n274 vdd.n272 0.358259
R21550 vdd.n276 vdd.n274 0.358259
R21551 vdd.n278 vdd.n276 0.358259
R21552 vdd.n320 vdd.n278 0.358259
R21553 vdd.n170 vdd.n168 0.358259
R21554 vdd.n172 vdd.n170 0.358259
R21555 vdd.n174 vdd.n172 0.358259
R21556 vdd.n176 vdd.n174 0.358259
R21557 vdd.n178 vdd.n176 0.358259
R21558 vdd.n180 vdd.n178 0.358259
R21559 vdd.n222 vdd.n180 0.358259
R21560 vdd.n73 vdd.n71 0.358259
R21561 vdd.n75 vdd.n73 0.358259
R21562 vdd.n77 vdd.n75 0.358259
R21563 vdd.n79 vdd.n77 0.358259
R21564 vdd.n81 vdd.n79 0.358259
R21565 vdd.n83 vdd.n81 0.358259
R21566 vdd.n125 vdd.n83 0.358259
R21567 vdd.n1744 vdd.n1702 0.358259
R21568 vdd.n1702 vdd.n1700 0.358259
R21569 vdd.n1700 vdd.n1698 0.358259
R21570 vdd.n1698 vdd.n1696 0.358259
R21571 vdd.n1696 vdd.n1694 0.358259
R21572 vdd.n1694 vdd.n1692 0.358259
R21573 vdd.n1692 vdd.n1690 0.358259
R21574 vdd.n1646 vdd.n1604 0.358259
R21575 vdd.n1604 vdd.n1602 0.358259
R21576 vdd.n1602 vdd.n1600 0.358259
R21577 vdd.n1600 vdd.n1598 0.358259
R21578 vdd.n1598 vdd.n1596 0.358259
R21579 vdd.n1596 vdd.n1594 0.358259
R21580 vdd.n1594 vdd.n1592 0.358259
R21581 vdd.n1549 vdd.n1507 0.358259
R21582 vdd.n1507 vdd.n1505 0.358259
R21583 vdd.n1505 vdd.n1503 0.358259
R21584 vdd.n1503 vdd.n1501 0.358259
R21585 vdd.n1501 vdd.n1499 0.358259
R21586 vdd.n1499 vdd.n1497 0.358259
R21587 vdd.n1497 vdd.n1495 0.358259
R21588 vdd.n14 vdd.n6 0.334552
R21589 vdd.n14 vdd.n13 0.334552
R21590 vdd.n27 vdd.n19 0.21707
R21591 vdd.n27 vdd.n24 0.21707
R21592 vdd.n318 vdd.n280 0.155672
R21593 vdd.n310 vdd.n280 0.155672
R21594 vdd.n310 vdd.n309 0.155672
R21595 vdd.n309 vdd.n285 0.155672
R21596 vdd.n302 vdd.n285 0.155672
R21597 vdd.n302 vdd.n301 0.155672
R21598 vdd.n301 vdd.n289 0.155672
R21599 vdd.n294 vdd.n289 0.155672
R21600 vdd.n263 vdd.n225 0.155672
R21601 vdd.n255 vdd.n225 0.155672
R21602 vdd.n255 vdd.n254 0.155672
R21603 vdd.n254 vdd.n230 0.155672
R21604 vdd.n247 vdd.n230 0.155672
R21605 vdd.n247 vdd.n246 0.155672
R21606 vdd.n246 vdd.n234 0.155672
R21607 vdd.n239 vdd.n234 0.155672
R21608 vdd.n220 vdd.n182 0.155672
R21609 vdd.n212 vdd.n182 0.155672
R21610 vdd.n212 vdd.n211 0.155672
R21611 vdd.n211 vdd.n187 0.155672
R21612 vdd.n204 vdd.n187 0.155672
R21613 vdd.n204 vdd.n203 0.155672
R21614 vdd.n203 vdd.n191 0.155672
R21615 vdd.n196 vdd.n191 0.155672
R21616 vdd.n165 vdd.n127 0.155672
R21617 vdd.n157 vdd.n127 0.155672
R21618 vdd.n157 vdd.n156 0.155672
R21619 vdd.n156 vdd.n132 0.155672
R21620 vdd.n149 vdd.n132 0.155672
R21621 vdd.n149 vdd.n148 0.155672
R21622 vdd.n148 vdd.n136 0.155672
R21623 vdd.n141 vdd.n136 0.155672
R21624 vdd.n123 vdd.n85 0.155672
R21625 vdd.n115 vdd.n85 0.155672
R21626 vdd.n115 vdd.n114 0.155672
R21627 vdd.n114 vdd.n90 0.155672
R21628 vdd.n107 vdd.n90 0.155672
R21629 vdd.n107 vdd.n106 0.155672
R21630 vdd.n106 vdd.n94 0.155672
R21631 vdd.n99 vdd.n94 0.155672
R21632 vdd.n68 vdd.n30 0.155672
R21633 vdd.n60 vdd.n30 0.155672
R21634 vdd.n60 vdd.n59 0.155672
R21635 vdd.n59 vdd.n35 0.155672
R21636 vdd.n52 vdd.n35 0.155672
R21637 vdd.n52 vdd.n51 0.155672
R21638 vdd.n51 vdd.n39 0.155672
R21639 vdd.n44 vdd.n39 0.155672
R21640 vdd.n1687 vdd.n1649 0.155672
R21641 vdd.n1679 vdd.n1649 0.155672
R21642 vdd.n1679 vdd.n1678 0.155672
R21643 vdd.n1678 vdd.n1654 0.155672
R21644 vdd.n1671 vdd.n1654 0.155672
R21645 vdd.n1671 vdd.n1670 0.155672
R21646 vdd.n1670 vdd.n1658 0.155672
R21647 vdd.n1663 vdd.n1658 0.155672
R21648 vdd.n1742 vdd.n1704 0.155672
R21649 vdd.n1734 vdd.n1704 0.155672
R21650 vdd.n1734 vdd.n1733 0.155672
R21651 vdd.n1733 vdd.n1709 0.155672
R21652 vdd.n1726 vdd.n1709 0.155672
R21653 vdd.n1726 vdd.n1725 0.155672
R21654 vdd.n1725 vdd.n1713 0.155672
R21655 vdd.n1718 vdd.n1713 0.155672
R21656 vdd.n1589 vdd.n1551 0.155672
R21657 vdd.n1581 vdd.n1551 0.155672
R21658 vdd.n1581 vdd.n1580 0.155672
R21659 vdd.n1580 vdd.n1556 0.155672
R21660 vdd.n1573 vdd.n1556 0.155672
R21661 vdd.n1573 vdd.n1572 0.155672
R21662 vdd.n1572 vdd.n1560 0.155672
R21663 vdd.n1565 vdd.n1560 0.155672
R21664 vdd.n1644 vdd.n1606 0.155672
R21665 vdd.n1636 vdd.n1606 0.155672
R21666 vdd.n1636 vdd.n1635 0.155672
R21667 vdd.n1635 vdd.n1611 0.155672
R21668 vdd.n1628 vdd.n1611 0.155672
R21669 vdd.n1628 vdd.n1627 0.155672
R21670 vdd.n1627 vdd.n1615 0.155672
R21671 vdd.n1620 vdd.n1615 0.155672
R21672 vdd.n1492 vdd.n1454 0.155672
R21673 vdd.n1484 vdd.n1454 0.155672
R21674 vdd.n1484 vdd.n1483 0.155672
R21675 vdd.n1483 vdd.n1459 0.155672
R21676 vdd.n1476 vdd.n1459 0.155672
R21677 vdd.n1476 vdd.n1475 0.155672
R21678 vdd.n1475 vdd.n1463 0.155672
R21679 vdd.n1468 vdd.n1463 0.155672
R21680 vdd.n1547 vdd.n1509 0.155672
R21681 vdd.n1539 vdd.n1509 0.155672
R21682 vdd.n1539 vdd.n1538 0.155672
R21683 vdd.n1538 vdd.n1514 0.155672
R21684 vdd.n1531 vdd.n1514 0.155672
R21685 vdd.n1531 vdd.n1530 0.155672
R21686 vdd.n1530 vdd.n1518 0.155672
R21687 vdd.n1523 vdd.n1518 0.155672
R21688 vdd.n2018 vdd.n1823 0.152939
R21689 vdd.n1829 vdd.n1823 0.152939
R21690 vdd.n1830 vdd.n1829 0.152939
R21691 vdd.n1831 vdd.n1830 0.152939
R21692 vdd.n1832 vdd.n1831 0.152939
R21693 vdd.n1836 vdd.n1832 0.152939
R21694 vdd.n1837 vdd.n1836 0.152939
R21695 vdd.n1838 vdd.n1837 0.152939
R21696 vdd.n1839 vdd.n1838 0.152939
R21697 vdd.n1843 vdd.n1839 0.152939
R21698 vdd.n1844 vdd.n1843 0.152939
R21699 vdd.n1845 vdd.n1844 0.152939
R21700 vdd.n1993 vdd.n1845 0.152939
R21701 vdd.n1993 vdd.n1992 0.152939
R21702 vdd.n1992 vdd.n1991 0.152939
R21703 vdd.n1991 vdd.n1851 0.152939
R21704 vdd.n1856 vdd.n1851 0.152939
R21705 vdd.n1857 vdd.n1856 0.152939
R21706 vdd.n1858 vdd.n1857 0.152939
R21707 vdd.n1862 vdd.n1858 0.152939
R21708 vdd.n1863 vdd.n1862 0.152939
R21709 vdd.n1864 vdd.n1863 0.152939
R21710 vdd.n1865 vdd.n1864 0.152939
R21711 vdd.n1869 vdd.n1865 0.152939
R21712 vdd.n1870 vdd.n1869 0.152939
R21713 vdd.n1871 vdd.n1870 0.152939
R21714 vdd.n1872 vdd.n1871 0.152939
R21715 vdd.n1876 vdd.n1872 0.152939
R21716 vdd.n1877 vdd.n1876 0.152939
R21717 vdd.n1878 vdd.n1877 0.152939
R21718 vdd.n1879 vdd.n1878 0.152939
R21719 vdd.n1883 vdd.n1879 0.152939
R21720 vdd.n1884 vdd.n1883 0.152939
R21721 vdd.n1885 vdd.n1884 0.152939
R21722 vdd.n1954 vdd.n1885 0.152939
R21723 vdd.n1954 vdd.n1953 0.152939
R21724 vdd.n1953 vdd.n1952 0.152939
R21725 vdd.n1952 vdd.n1891 0.152939
R21726 vdd.n1896 vdd.n1891 0.152939
R21727 vdd.n1897 vdd.n1896 0.152939
R21728 vdd.n1898 vdd.n1897 0.152939
R21729 vdd.n1902 vdd.n1898 0.152939
R21730 vdd.n1903 vdd.n1902 0.152939
R21731 vdd.n1904 vdd.n1903 0.152939
R21732 vdd.n1905 vdd.n1904 0.152939
R21733 vdd.n1909 vdd.n1905 0.152939
R21734 vdd.n1910 vdd.n1909 0.152939
R21735 vdd.n1911 vdd.n1910 0.152939
R21736 vdd.n1912 vdd.n1911 0.152939
R21737 vdd.n1913 vdd.n1912 0.152939
R21738 vdd.n1913 vdd.n1035 0.152939
R21739 vdd.n2242 vdd.n1817 0.152939
R21740 vdd.n1749 vdd.n1748 0.152939
R21741 vdd.n1749 vdd.n1084 0.152939
R21742 vdd.n1763 vdd.n1084 0.152939
R21743 vdd.n1764 vdd.n1763 0.152939
R21744 vdd.n1765 vdd.n1764 0.152939
R21745 vdd.n1765 vdd.n1072 0.152939
R21746 vdd.n1780 vdd.n1072 0.152939
R21747 vdd.n1781 vdd.n1780 0.152939
R21748 vdd.n1782 vdd.n1781 0.152939
R21749 vdd.n1782 vdd.n1061 0.152939
R21750 vdd.n1797 vdd.n1061 0.152939
R21751 vdd.n1798 vdd.n1797 0.152939
R21752 vdd.n1799 vdd.n1798 0.152939
R21753 vdd.n1799 vdd.n1049 0.152939
R21754 vdd.n1815 vdd.n1049 0.152939
R21755 vdd.n1816 vdd.n1815 0.152939
R21756 vdd.n2243 vdd.n1816 0.152939
R21757 vdd.n670 vdd.n667 0.152939
R21758 vdd.n671 vdd.n670 0.152939
R21759 vdd.n672 vdd.n671 0.152939
R21760 vdd.n673 vdd.n672 0.152939
R21761 vdd.n676 vdd.n673 0.152939
R21762 vdd.n677 vdd.n676 0.152939
R21763 vdd.n678 vdd.n677 0.152939
R21764 vdd.n679 vdd.n678 0.152939
R21765 vdd.n682 vdd.n679 0.152939
R21766 vdd.n683 vdd.n682 0.152939
R21767 vdd.n684 vdd.n683 0.152939
R21768 vdd.n685 vdd.n684 0.152939
R21769 vdd.n690 vdd.n685 0.152939
R21770 vdd.n691 vdd.n690 0.152939
R21771 vdd.n692 vdd.n691 0.152939
R21772 vdd.n693 vdd.n692 0.152939
R21773 vdd.n696 vdd.n693 0.152939
R21774 vdd.n697 vdd.n696 0.152939
R21775 vdd.n698 vdd.n697 0.152939
R21776 vdd.n699 vdd.n698 0.152939
R21777 vdd.n702 vdd.n699 0.152939
R21778 vdd.n703 vdd.n702 0.152939
R21779 vdd.n704 vdd.n703 0.152939
R21780 vdd.n705 vdd.n704 0.152939
R21781 vdd.n708 vdd.n705 0.152939
R21782 vdd.n709 vdd.n708 0.152939
R21783 vdd.n710 vdd.n709 0.152939
R21784 vdd.n711 vdd.n710 0.152939
R21785 vdd.n714 vdd.n711 0.152939
R21786 vdd.n715 vdd.n714 0.152939
R21787 vdd.n716 vdd.n715 0.152939
R21788 vdd.n717 vdd.n716 0.152939
R21789 vdd.n720 vdd.n717 0.152939
R21790 vdd.n721 vdd.n720 0.152939
R21791 vdd.n3058 vdd.n721 0.152939
R21792 vdd.n3058 vdd.n3057 0.152939
R21793 vdd.n3057 vdd.n3056 0.152939
R21794 vdd.n3056 vdd.n725 0.152939
R21795 vdd.n730 vdd.n725 0.152939
R21796 vdd.n731 vdd.n730 0.152939
R21797 vdd.n734 vdd.n731 0.152939
R21798 vdd.n735 vdd.n734 0.152939
R21799 vdd.n736 vdd.n735 0.152939
R21800 vdd.n737 vdd.n736 0.152939
R21801 vdd.n740 vdd.n737 0.152939
R21802 vdd.n741 vdd.n740 0.152939
R21803 vdd.n742 vdd.n741 0.152939
R21804 vdd.n743 vdd.n742 0.152939
R21805 vdd.n746 vdd.n743 0.152939
R21806 vdd.n747 vdd.n746 0.152939
R21807 vdd.n748 vdd.n747 0.152939
R21808 vdd.n3141 vdd.n661 0.152939
R21809 vdd.n3142 vdd.n651 0.152939
R21810 vdd.n3156 vdd.n651 0.152939
R21811 vdd.n3157 vdd.n3156 0.152939
R21812 vdd.n3158 vdd.n3157 0.152939
R21813 vdd.n3158 vdd.n639 0.152939
R21814 vdd.n3172 vdd.n639 0.152939
R21815 vdd.n3173 vdd.n3172 0.152939
R21816 vdd.n3174 vdd.n3173 0.152939
R21817 vdd.n3174 vdd.n627 0.152939
R21818 vdd.n3189 vdd.n627 0.152939
R21819 vdd.n3190 vdd.n3189 0.152939
R21820 vdd.n3191 vdd.n3190 0.152939
R21821 vdd.n3191 vdd.n616 0.152939
R21822 vdd.n3208 vdd.n616 0.152939
R21823 vdd.n3209 vdd.n3208 0.152939
R21824 vdd.n3210 vdd.n3209 0.152939
R21825 vdd.n3210 vdd.n322 0.152939
R21826 vdd.n3290 vdd.n323 0.152939
R21827 vdd.n334 vdd.n323 0.152939
R21828 vdd.n335 vdd.n334 0.152939
R21829 vdd.n336 vdd.n335 0.152939
R21830 vdd.n343 vdd.n336 0.152939
R21831 vdd.n344 vdd.n343 0.152939
R21832 vdd.n345 vdd.n344 0.152939
R21833 vdd.n346 vdd.n345 0.152939
R21834 vdd.n354 vdd.n346 0.152939
R21835 vdd.n355 vdd.n354 0.152939
R21836 vdd.n356 vdd.n355 0.152939
R21837 vdd.n357 vdd.n356 0.152939
R21838 vdd.n365 vdd.n357 0.152939
R21839 vdd.n366 vdd.n365 0.152939
R21840 vdd.n367 vdd.n366 0.152939
R21841 vdd.n368 vdd.n367 0.152939
R21842 vdd.n443 vdd.n368 0.152939
R21843 vdd.n444 vdd.n442 0.152939
R21844 vdd.n451 vdd.n442 0.152939
R21845 vdd.n452 vdd.n451 0.152939
R21846 vdd.n453 vdd.n452 0.152939
R21847 vdd.n453 vdd.n440 0.152939
R21848 vdd.n461 vdd.n440 0.152939
R21849 vdd.n462 vdd.n461 0.152939
R21850 vdd.n463 vdd.n462 0.152939
R21851 vdd.n463 vdd.n438 0.152939
R21852 vdd.n471 vdd.n438 0.152939
R21853 vdd.n472 vdd.n471 0.152939
R21854 vdd.n473 vdd.n472 0.152939
R21855 vdd.n473 vdd.n436 0.152939
R21856 vdd.n481 vdd.n436 0.152939
R21857 vdd.n482 vdd.n481 0.152939
R21858 vdd.n483 vdd.n482 0.152939
R21859 vdd.n483 vdd.n434 0.152939
R21860 vdd.n491 vdd.n434 0.152939
R21861 vdd.n492 vdd.n491 0.152939
R21862 vdd.n493 vdd.n492 0.152939
R21863 vdd.n493 vdd.n430 0.152939
R21864 vdd.n501 vdd.n430 0.152939
R21865 vdd.n502 vdd.n501 0.152939
R21866 vdd.n503 vdd.n502 0.152939
R21867 vdd.n503 vdd.n428 0.152939
R21868 vdd.n511 vdd.n428 0.152939
R21869 vdd.n512 vdd.n511 0.152939
R21870 vdd.n513 vdd.n512 0.152939
R21871 vdd.n513 vdd.n426 0.152939
R21872 vdd.n521 vdd.n426 0.152939
R21873 vdd.n522 vdd.n521 0.152939
R21874 vdd.n523 vdd.n522 0.152939
R21875 vdd.n523 vdd.n424 0.152939
R21876 vdd.n531 vdd.n424 0.152939
R21877 vdd.n532 vdd.n531 0.152939
R21878 vdd.n533 vdd.n532 0.152939
R21879 vdd.n533 vdd.n422 0.152939
R21880 vdd.n541 vdd.n422 0.152939
R21881 vdd.n542 vdd.n541 0.152939
R21882 vdd.n543 vdd.n542 0.152939
R21883 vdd.n543 vdd.n418 0.152939
R21884 vdd.n551 vdd.n418 0.152939
R21885 vdd.n552 vdd.n551 0.152939
R21886 vdd.n553 vdd.n552 0.152939
R21887 vdd.n553 vdd.n416 0.152939
R21888 vdd.n561 vdd.n416 0.152939
R21889 vdd.n562 vdd.n561 0.152939
R21890 vdd.n563 vdd.n562 0.152939
R21891 vdd.n563 vdd.n414 0.152939
R21892 vdd.n571 vdd.n414 0.152939
R21893 vdd.n572 vdd.n571 0.152939
R21894 vdd.n573 vdd.n572 0.152939
R21895 vdd.n573 vdd.n412 0.152939
R21896 vdd.n581 vdd.n412 0.152939
R21897 vdd.n582 vdd.n581 0.152939
R21898 vdd.n583 vdd.n582 0.152939
R21899 vdd.n583 vdd.n410 0.152939
R21900 vdd.n591 vdd.n410 0.152939
R21901 vdd.n592 vdd.n591 0.152939
R21902 vdd.n593 vdd.n592 0.152939
R21903 vdd.n593 vdd.n408 0.152939
R21904 vdd.n600 vdd.n408 0.152939
R21905 vdd.n3249 vdd.n600 0.152939
R21906 vdd.n3149 vdd.n3148 0.152939
R21907 vdd.n3150 vdd.n3149 0.152939
R21908 vdd.n3150 vdd.n645 0.152939
R21909 vdd.n3164 vdd.n645 0.152939
R21910 vdd.n3165 vdd.n3164 0.152939
R21911 vdd.n3166 vdd.n3165 0.152939
R21912 vdd.n3166 vdd.n632 0.152939
R21913 vdd.n3180 vdd.n632 0.152939
R21914 vdd.n3181 vdd.n3180 0.152939
R21915 vdd.n3182 vdd.n3181 0.152939
R21916 vdd.n3182 vdd.n621 0.152939
R21917 vdd.n3197 vdd.n621 0.152939
R21918 vdd.n3198 vdd.n3197 0.152939
R21919 vdd.n3199 vdd.n3198 0.152939
R21920 vdd.n3201 vdd.n3199 0.152939
R21921 vdd.n3201 vdd.n3200 0.152939
R21922 vdd.n3200 vdd.n611 0.152939
R21923 vdd.n611 vdd.n609 0.152939
R21924 vdd.n3219 vdd.n609 0.152939
R21925 vdd.n3220 vdd.n3219 0.152939
R21926 vdd.n3221 vdd.n3220 0.152939
R21927 vdd.n3221 vdd.n607 0.152939
R21928 vdd.n3226 vdd.n607 0.152939
R21929 vdd.n3227 vdd.n3226 0.152939
R21930 vdd.n3228 vdd.n3227 0.152939
R21931 vdd.n3228 vdd.n605 0.152939
R21932 vdd.n3233 vdd.n605 0.152939
R21933 vdd.n3234 vdd.n3233 0.152939
R21934 vdd.n3235 vdd.n3234 0.152939
R21935 vdd.n3235 vdd.n603 0.152939
R21936 vdd.n3241 vdd.n603 0.152939
R21937 vdd.n3242 vdd.n3241 0.152939
R21938 vdd.n3243 vdd.n3242 0.152939
R21939 vdd.n3243 vdd.n601 0.152939
R21940 vdd.n3248 vdd.n601 0.152939
R21941 vdd.n3011 vdd.n656 0.152939
R21942 vdd.n2254 vdd.n1038 0.152939
R21943 vdd.n1379 vdd.n1378 0.152939
R21944 vdd.n1379 vdd.n1135 0.152939
R21945 vdd.n1393 vdd.n1135 0.152939
R21946 vdd.n1394 vdd.n1393 0.152939
R21947 vdd.n1395 vdd.n1394 0.152939
R21948 vdd.n1395 vdd.n1123 0.152939
R21949 vdd.n1410 vdd.n1123 0.152939
R21950 vdd.n1411 vdd.n1410 0.152939
R21951 vdd.n1412 vdd.n1411 0.152939
R21952 vdd.n1412 vdd.n1113 0.152939
R21953 vdd.n1427 vdd.n1113 0.152939
R21954 vdd.n1428 vdd.n1427 0.152939
R21955 vdd.n1429 vdd.n1428 0.152939
R21956 vdd.n1429 vdd.n1100 0.152939
R21957 vdd.n1443 vdd.n1100 0.152939
R21958 vdd.n1444 vdd.n1443 0.152939
R21959 vdd.n1445 vdd.n1444 0.152939
R21960 vdd.n1445 vdd.n1089 0.152939
R21961 vdd.n1755 vdd.n1089 0.152939
R21962 vdd.n1756 vdd.n1755 0.152939
R21963 vdd.n1757 vdd.n1756 0.152939
R21964 vdd.n1757 vdd.n1078 0.152939
R21965 vdd.n1771 vdd.n1078 0.152939
R21966 vdd.n1772 vdd.n1771 0.152939
R21967 vdd.n1773 vdd.n1772 0.152939
R21968 vdd.n1773 vdd.n1066 0.152939
R21969 vdd.n1788 vdd.n1066 0.152939
R21970 vdd.n1789 vdd.n1788 0.152939
R21971 vdd.n1790 vdd.n1789 0.152939
R21972 vdd.n1790 vdd.n1056 0.152939
R21973 vdd.n1805 vdd.n1056 0.152939
R21974 vdd.n1806 vdd.n1805 0.152939
R21975 vdd.n1809 vdd.n1806 0.152939
R21976 vdd.n1809 vdd.n1808 0.152939
R21977 vdd.n1808 vdd.n1807 0.152939
R21978 vdd.n1369 vdd.n1184 0.152939
R21979 vdd.n1369 vdd.n1368 0.152939
R21980 vdd.n1368 vdd.n1367 0.152939
R21981 vdd.n1367 vdd.n1186 0.152939
R21982 vdd.n1363 vdd.n1186 0.152939
R21983 vdd.n1363 vdd.n1362 0.152939
R21984 vdd.n1362 vdd.n1361 0.152939
R21985 vdd.n1361 vdd.n1191 0.152939
R21986 vdd.n1357 vdd.n1191 0.152939
R21987 vdd.n1357 vdd.n1356 0.152939
R21988 vdd.n1356 vdd.n1355 0.152939
R21989 vdd.n1355 vdd.n1197 0.152939
R21990 vdd.n1351 vdd.n1197 0.152939
R21991 vdd.n1351 vdd.n1350 0.152939
R21992 vdd.n1350 vdd.n1349 0.152939
R21993 vdd.n1349 vdd.n1203 0.152939
R21994 vdd.n1345 vdd.n1203 0.152939
R21995 vdd.n1345 vdd.n1344 0.152939
R21996 vdd.n1344 vdd.n1343 0.152939
R21997 vdd.n1343 vdd.n1209 0.152939
R21998 vdd.n1335 vdd.n1209 0.152939
R21999 vdd.n1335 vdd.n1334 0.152939
R22000 vdd.n1334 vdd.n1333 0.152939
R22001 vdd.n1333 vdd.n1213 0.152939
R22002 vdd.n1329 vdd.n1213 0.152939
R22003 vdd.n1329 vdd.n1328 0.152939
R22004 vdd.n1328 vdd.n1327 0.152939
R22005 vdd.n1327 vdd.n1219 0.152939
R22006 vdd.n1323 vdd.n1219 0.152939
R22007 vdd.n1323 vdd.n1322 0.152939
R22008 vdd.n1322 vdd.n1321 0.152939
R22009 vdd.n1321 vdd.n1225 0.152939
R22010 vdd.n1317 vdd.n1225 0.152939
R22011 vdd.n1317 vdd.n1316 0.152939
R22012 vdd.n1316 vdd.n1315 0.152939
R22013 vdd.n1315 vdd.n1231 0.152939
R22014 vdd.n1311 vdd.n1231 0.152939
R22015 vdd.n1311 vdd.n1310 0.152939
R22016 vdd.n1310 vdd.n1309 0.152939
R22017 vdd.n1309 vdd.n1237 0.152939
R22018 vdd.n1302 vdd.n1237 0.152939
R22019 vdd.n1302 vdd.n1301 0.152939
R22020 vdd.n1301 vdd.n1300 0.152939
R22021 vdd.n1300 vdd.n1242 0.152939
R22022 vdd.n1296 vdd.n1242 0.152939
R22023 vdd.n1296 vdd.n1295 0.152939
R22024 vdd.n1295 vdd.n1294 0.152939
R22025 vdd.n1294 vdd.n1248 0.152939
R22026 vdd.n1290 vdd.n1248 0.152939
R22027 vdd.n1290 vdd.n1289 0.152939
R22028 vdd.n1289 vdd.n1288 0.152939
R22029 vdd.n1288 vdd.n1254 0.152939
R22030 vdd.n1284 vdd.n1254 0.152939
R22031 vdd.n1284 vdd.n1283 0.152939
R22032 vdd.n1283 vdd.n1282 0.152939
R22033 vdd.n1282 vdd.n1260 0.152939
R22034 vdd.n1278 vdd.n1260 0.152939
R22035 vdd.n1278 vdd.n1277 0.152939
R22036 vdd.n1277 vdd.n1276 0.152939
R22037 vdd.n1276 vdd.n1266 0.152939
R22038 vdd.n1272 vdd.n1266 0.152939
R22039 vdd.n1272 vdd.n1147 0.152939
R22040 vdd.n1377 vdd.n1147 0.152939
R22041 vdd.n1385 vdd.n1141 0.152939
R22042 vdd.n1386 vdd.n1385 0.152939
R22043 vdd.n1387 vdd.n1386 0.152939
R22044 vdd.n1387 vdd.n1129 0.152939
R22045 vdd.n1402 vdd.n1129 0.152939
R22046 vdd.n1403 vdd.n1402 0.152939
R22047 vdd.n1404 vdd.n1403 0.152939
R22048 vdd.n1404 vdd.n1118 0.152939
R22049 vdd.n1419 vdd.n1118 0.152939
R22050 vdd.n1420 vdd.n1419 0.152939
R22051 vdd.n1421 vdd.n1420 0.152939
R22052 vdd.n1421 vdd.n1107 0.152939
R22053 vdd.n1435 vdd.n1107 0.152939
R22054 vdd.n1436 vdd.n1435 0.152939
R22055 vdd.n1437 vdd.n1436 0.152939
R22056 vdd.n1437 vdd.n1095 0.152939
R22057 vdd.n1452 vdd.n1095 0.152939
R22058 vdd.n2232 vdd.n1817 0.110256
R22059 vdd.n2942 vdd.n661 0.110256
R22060 vdd.n3011 vdd.n3010 0.110256
R22061 vdd.n2255 vdd.n2254 0.110256
R22062 vdd.n1748 vdd.n1747 0.0695946
R22063 vdd.n3291 vdd.n322 0.0695946
R22064 vdd.n3291 vdd.n3290 0.0695946
R22065 vdd.n1747 vdd.n1452 0.0695946
R22066 vdd.n2232 vdd.n2018 0.0431829
R22067 vdd.n2255 vdd.n1035 0.0431829
R22068 vdd.n2942 vdd.n667 0.0431829
R22069 vdd.n3010 vdd.n748 0.0431829
R22070 vdd vdd.n28 0.00833333
R22071 a_n1986_13878.n6 a_n1986_13878.t66 539.01
R22072 a_n1986_13878.n66 a_n1986_13878.t49 512.366
R22073 a_n1986_13878.n65 a_n1986_13878.t53 512.366
R22074 a_n1986_13878.n63 a_n1986_13878.t43 512.366
R22075 a_n1986_13878.n64 a_n1986_13878.t58 512.366
R22076 a_n1986_13878.n50 a_n1986_13878.t19 533.058
R22077 a_n1986_13878.n8 a_n1986_13878.t11 539.01
R22078 a_n1986_13878.n69 a_n1986_13878.t17 512.366
R22079 a_n1986_13878.n68 a_n1986_13878.t13 512.366
R22080 a_n1986_13878.n54 a_n1986_13878.t29 512.366
R22081 a_n1986_13878.n67 a_n1986_13878.t27 512.366
R22082 a_n1986_13878.n20 a_n1986_13878.t9 539.01
R22083 a_n1986_13878.n90 a_n1986_13878.t25 512.366
R22084 a_n1986_13878.n91 a_n1986_13878.t21 512.366
R22085 a_n1986_13878.n52 a_n1986_13878.t15 512.366
R22086 a_n1986_13878.n92 a_n1986_13878.t7 512.366
R22087 a_n1986_13878.n24 a_n1986_13878.t61 539.01
R22088 a_n1986_13878.n87 a_n1986_13878.t62 512.366
R22089 a_n1986_13878.n88 a_n1986_13878.t41 512.366
R22090 a_n1986_13878.n53 a_n1986_13878.t48 512.366
R22091 a_n1986_13878.n89 a_n1986_13878.t57 512.366
R22092 a_n1986_13878.n79 a_n1986_13878.t55 512.366
R22093 a_n1986_13878.n78 a_n1986_13878.t46 512.366
R22094 a_n1986_13878.n77 a_n1986_13878.t40 512.366
R22095 a_n1986_13878.n81 a_n1986_13878.t63 512.366
R22096 a_n1986_13878.n80 a_n1986_13878.t52 512.366
R22097 a_n1986_13878.n76 a_n1986_13878.t51 512.366
R22098 a_n1986_13878.n83 a_n1986_13878.t59 512.366
R22099 a_n1986_13878.n82 a_n1986_13878.t44 512.366
R22100 a_n1986_13878.n75 a_n1986_13878.t45 512.366
R22101 a_n1986_13878.n85 a_n1986_13878.t47 512.366
R22102 a_n1986_13878.n84 a_n1986_13878.t56 512.366
R22103 a_n1986_13878.n74 a_n1986_13878.t67 512.366
R22104 a_n1986_13878.n49 a_n1986_13878.n4 70.3058
R22105 a_n1986_13878.n17 a_n1986_13878.n34 70.3058
R22106 a_n1986_13878.n21 a_n1986_13878.n31 70.3058
R22107 a_n1986_13878.n30 a_n1986_13878.n22 70.1674
R22108 a_n1986_13878.n30 a_n1986_13878.n53 20.9683
R22109 a_n1986_13878.n22 a_n1986_13878.n29 75.0448
R22110 a_n1986_13878.n88 a_n1986_13878.n29 11.2134
R22111 a_n1986_13878.n23 a_n1986_13878.n24 44.8194
R22112 a_n1986_13878.n33 a_n1986_13878.n18 70.1674
R22113 a_n1986_13878.n33 a_n1986_13878.n52 20.9683
R22114 a_n1986_13878.n18 a_n1986_13878.n32 75.0448
R22115 a_n1986_13878.n91 a_n1986_13878.n32 11.2134
R22116 a_n1986_13878.n19 a_n1986_13878.n20 44.8194
R22117 a_n1986_13878.n9 a_n1986_13878.n43 70.1674
R22118 a_n1986_13878.n11 a_n1986_13878.n40 70.1674
R22119 a_n1986_13878.n13 a_n1986_13878.n38 70.1674
R22120 a_n1986_13878.n15 a_n1986_13878.n36 70.1674
R22121 a_n1986_13878.n36 a_n1986_13878.n74 20.9683
R22122 a_n1986_13878.n35 a_n1986_13878.n16 75.0448
R22123 a_n1986_13878.n84 a_n1986_13878.n35 11.2134
R22124 a_n1986_13878.n16 a_n1986_13878.n85 161.3
R22125 a_n1986_13878.n38 a_n1986_13878.n75 20.9683
R22126 a_n1986_13878.n37 a_n1986_13878.n14 75.0448
R22127 a_n1986_13878.n82 a_n1986_13878.n37 11.2134
R22128 a_n1986_13878.n14 a_n1986_13878.n83 161.3
R22129 a_n1986_13878.n40 a_n1986_13878.n76 20.9683
R22130 a_n1986_13878.n39 a_n1986_13878.n12 75.0448
R22131 a_n1986_13878.n80 a_n1986_13878.n39 11.2134
R22132 a_n1986_13878.n12 a_n1986_13878.n81 161.3
R22133 a_n1986_13878.n43 a_n1986_13878.n77 20.9683
R22134 a_n1986_13878.n41 a_n1986_13878.n10 75.0448
R22135 a_n1986_13878.n78 a_n1986_13878.n41 11.2134
R22136 a_n1986_13878.n10 a_n1986_13878.n79 161.3
R22137 a_n1986_13878.n28 a_n1986_13878.n46 70.1674
R22138 a_n1986_13878.n46 a_n1986_13878.n54 20.9683
R22139 a_n1986_13878.n45 a_n1986_13878.n44 75.0448
R22140 a_n1986_13878.n68 a_n1986_13878.n45 11.2134
R22141 a_n1986_13878.n7 a_n1986_13878.n8 44.8194
R22142 a_n1986_13878.n50 a_n1986_13878.n28 70.3058
R22143 a_n1986_13878.n5 a_n1986_13878.n48 70.1674
R22144 a_n1986_13878.n48 a_n1986_13878.n63 20.9683
R22145 a_n1986_13878.n47 a_n1986_13878.n5 75.0448
R22146 a_n1986_13878.n65 a_n1986_13878.n47 11.2134
R22147 a_n1986_13878.n3 a_n1986_13878.n6 44.8194
R22148 a_n1986_13878.n1 a_n1986_13878.n61 81.4626
R22149 a_n1986_13878.n2 a_n1986_13878.n57 81.4626
R22150 a_n1986_13878.n2 a_n1986_13878.n55 81.4626
R22151 a_n1986_13878.n1 a_n1986_13878.n62 80.9324
R22152 a_n1986_13878.n1 a_n1986_13878.n60 80.9324
R22153 a_n1986_13878.n0 a_n1986_13878.n59 80.9324
R22154 a_n1986_13878.n2 a_n1986_13878.n58 80.9324
R22155 a_n1986_13878.n2 a_n1986_13878.n56 80.9324
R22156 a_n1986_13878.n26 a_n1986_13878.t10 74.6477
R22157 a_n1986_13878.n25 a_n1986_13878.t20 74.6477
R22158 a_n1986_13878.n72 a_n1986_13878.t12 74.2899
R22159 a_n1986_13878.n27 a_n1986_13878.t24 74.2897
R22160 a_n1986_13878.n26 a_n1986_13878.n51 70.6783
R22161 a_n1986_13878.n25 a_n1986_13878.n70 70.6783
R22162 a_n1986_13878.n25 a_n1986_13878.n71 70.6783
R22163 a_n1986_13878.n94 a_n1986_13878.n27 70.6782
R22164 a_n1986_13878.n66 a_n1986_13878.n65 48.2005
R22165 a_n1986_13878.n64 a_n1986_13878.n48 20.9683
R22166 a_n1986_13878.n69 a_n1986_13878.n68 48.2005
R22167 a_n1986_13878.n67 a_n1986_13878.n46 20.9683
R22168 a_n1986_13878.n91 a_n1986_13878.n90 48.2005
R22169 a_n1986_13878.n92 a_n1986_13878.n33 20.9683
R22170 a_n1986_13878.n88 a_n1986_13878.n87 48.2005
R22171 a_n1986_13878.n89 a_n1986_13878.n30 20.9683
R22172 a_n1986_13878.n79 a_n1986_13878.n78 48.2005
R22173 a_n1986_13878.t60 a_n1986_13878.n43 533.335
R22174 a_n1986_13878.n81 a_n1986_13878.n80 48.2005
R22175 a_n1986_13878.t65 a_n1986_13878.n40 533.335
R22176 a_n1986_13878.n83 a_n1986_13878.n82 48.2005
R22177 a_n1986_13878.t54 a_n1986_13878.n38 533.335
R22178 a_n1986_13878.n85 a_n1986_13878.n84 48.2005
R22179 a_n1986_13878.t50 a_n1986_13878.n36 533.335
R22180 a_n1986_13878.n49 a_n1986_13878.t64 533.058
R22181 a_n1986_13878.t23 a_n1986_13878.n34 533.058
R22182 a_n1986_13878.t42 a_n1986_13878.n31 533.058
R22183 a_n1986_13878.n47 a_n1986_13878.n63 35.3134
R22184 a_n1986_13878.n45 a_n1986_13878.n54 35.3134
R22185 a_n1986_13878.n52 a_n1986_13878.n32 35.3134
R22186 a_n1986_13878.n53 a_n1986_13878.n29 35.3134
R22187 a_n1986_13878.n41 a_n1986_13878.n77 35.3134
R22188 a_n1986_13878.n39 a_n1986_13878.n76 35.3134
R22189 a_n1986_13878.n37 a_n1986_13878.n75 35.3134
R22190 a_n1986_13878.n35 a_n1986_13878.n74 35.3134
R22191 a_n1986_13878.n0 a_n1986_13878.n2 32.5247
R22192 a_n1986_13878.n28 a_n1986_13878.n1 23.891
R22193 a_n1986_13878.n23 a_n1986_13878.n86 12.046
R22194 a_n1986_13878.n4 a_n1986_13878.n42 11.8414
R22195 a_n1986_13878.n73 a_n1986_13878.n7 10.5365
R22196 a_n1986_13878.n27 a_n1986_13878.n93 9.50122
R22197 a_n1986_13878.n9 a_n1986_13878.n42 7.47588
R22198 a_n1986_13878.n86 a_n1986_13878.n16 7.47588
R22199 a_n1986_13878.n93 a_n1986_13878.n17 6.70126
R22200 a_n1986_13878.n73 a_n1986_13878.n72 5.65783
R22201 a_n1986_13878.n93 a_n1986_13878.n42 5.3452
R22202 a_n1986_13878.n19 a_n1986_13878.n21 3.95126
R22203 a_n1986_13878.n28 a_n1986_13878.n3 3.95126
R22204 a_n1986_13878.n51 a_n1986_13878.t26 3.61217
R22205 a_n1986_13878.n51 a_n1986_13878.t22 3.61217
R22206 a_n1986_13878.n70 a_n1986_13878.t30 3.61217
R22207 a_n1986_13878.n70 a_n1986_13878.t28 3.61217
R22208 a_n1986_13878.n71 a_n1986_13878.t18 3.61217
R22209 a_n1986_13878.n71 a_n1986_13878.t14 3.61217
R22210 a_n1986_13878.n94 a_n1986_13878.t16 3.61217
R22211 a_n1986_13878.t8 a_n1986_13878.n94 3.61217
R22212 a_n1986_13878.n61 a_n1986_13878.t1 2.82907
R22213 a_n1986_13878.n61 a_n1986_13878.t39 2.82907
R22214 a_n1986_13878.n62 a_n1986_13878.t35 2.82907
R22215 a_n1986_13878.n62 a_n1986_13878.t0 2.82907
R22216 a_n1986_13878.n60 a_n1986_13878.t4 2.82907
R22217 a_n1986_13878.n60 a_n1986_13878.t3 2.82907
R22218 a_n1986_13878.n59 a_n1986_13878.t6 2.82907
R22219 a_n1986_13878.n59 a_n1986_13878.t36 2.82907
R22220 a_n1986_13878.n57 a_n1986_13878.t38 2.82907
R22221 a_n1986_13878.n57 a_n1986_13878.t33 2.82907
R22222 a_n1986_13878.n58 a_n1986_13878.t5 2.82907
R22223 a_n1986_13878.n58 a_n1986_13878.t34 2.82907
R22224 a_n1986_13878.n56 a_n1986_13878.t2 2.82907
R22225 a_n1986_13878.n56 a_n1986_13878.t32 2.82907
R22226 a_n1986_13878.n55 a_n1986_13878.t37 2.82907
R22227 a_n1986_13878.n55 a_n1986_13878.t31 2.82907
R22228 a_n1986_13878.n86 a_n1986_13878.n73 1.30542
R22229 a_n1986_13878.n13 a_n1986_13878.n12 1.04595
R22230 a_n1986_13878.n6 a_n1986_13878.n66 13.657
R22231 a_n1986_13878.n64 a_n1986_13878.n49 21.4216
R22232 a_n1986_13878.n8 a_n1986_13878.n69 13.657
R22233 a_n1986_13878.n67 a_n1986_13878.n50 21.4216
R22234 a_n1986_13878.n90 a_n1986_13878.n20 13.657
R22235 a_n1986_13878.n34 a_n1986_13878.n92 21.4216
R22236 a_n1986_13878.n87 a_n1986_13878.n24 13.657
R22237 a_n1986_13878.n31 a_n1986_13878.n89 21.4216
R22238 a_n1986_13878.n1 a_n1986_13878.n0 1.06084
R22239 a_n1986_13878.n23 a_n1986_13878.n22 0.758076
R22240 a_n1986_13878.n22 a_n1986_13878.n21 0.758076
R22241 a_n1986_13878.n19 a_n1986_13878.n18 0.758076
R22242 a_n1986_13878.n18 a_n1986_13878.n17 0.758076
R22243 a_n1986_13878.n16 a_n1986_13878.n15 0.758076
R22244 a_n1986_13878.n14 a_n1986_13878.n13 0.758076
R22245 a_n1986_13878.n12 a_n1986_13878.n11 0.758076
R22246 a_n1986_13878.n10 a_n1986_13878.n9 0.758076
R22247 a_n1986_13878.n44 a_n1986_13878.n7 0.758076
R22248 a_n1986_13878.n5 a_n1986_13878.n3 0.758076
R22249 a_n1986_13878.n5 a_n1986_13878.n4 0.758076
R22250 a_n1986_13878.n44 a_n1986_13878.n28 0.720197
R22251 a_n1986_13878.n27 a_n1986_13878.n26 0.716017
R22252 a_n1986_13878.n72 a_n1986_13878.n25 0.716017
R22253 a_n1986_13878.n15 a_n1986_13878.n14 0.67853
R22254 a_n1986_13878.n11 a_n1986_13878.n10 0.67853
R22255 a_n1808_13878.n2 a_n1808_13878.n0 98.9633
R22256 a_n1808_13878.n5 a_n1808_13878.n3 98.7517
R22257 a_n1808_13878.n2 a_n1808_13878.n1 98.6055
R22258 a_n1808_13878.n7 a_n1808_13878.n6 98.6055
R22259 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R22260 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R22261 a_n1808_13878.n9 a_n1808_13878.t1 74.6477
R22262 a_n1808_13878.n14 a_n1808_13878.t2 74.2899
R22263 a_n1808_13878.n11 a_n1808_13878.t3 74.2899
R22264 a_n1808_13878.n10 a_n1808_13878.t0 74.2899
R22265 a_n1808_13878.n13 a_n1808_13878.n12 70.6783
R22266 a_n1808_13878.n9 a_n1808_13878.n8 70.6783
R22267 a_n1808_13878.n15 a_n1808_13878.n7 13.5694
R22268 a_n1808_13878.n16 a_n1808_13878.n15 11.5762
R22269 a_n1808_13878.n15 a_n1808_13878.n14 6.2408
R22270 a_n1808_13878.n1 a_n1808_13878.t8 3.61217
R22271 a_n1808_13878.n1 a_n1808_13878.t13 3.61217
R22272 a_n1808_13878.n0 a_n1808_13878.t15 3.61217
R22273 a_n1808_13878.n0 a_n1808_13878.t19 3.61217
R22274 a_n1808_13878.n12 a_n1808_13878.t6 3.61217
R22275 a_n1808_13878.n12 a_n1808_13878.t7 3.61217
R22276 a_n1808_13878.n8 a_n1808_13878.t4 3.61217
R22277 a_n1808_13878.n8 a_n1808_13878.t5 3.61217
R22278 a_n1808_13878.n6 a_n1808_13878.t14 3.61217
R22279 a_n1808_13878.n6 a_n1808_13878.t9 3.61217
R22280 a_n1808_13878.n4 a_n1808_13878.t16 3.61217
R22281 a_n1808_13878.n4 a_n1808_13878.t11 3.61217
R22282 a_n1808_13878.n3 a_n1808_13878.t10 3.61217
R22283 a_n1808_13878.n3 a_n1808_13878.t12 3.61217
R22284 a_n1808_13878.n17 a_n1808_13878.t17 3.61217
R22285 a_n1808_13878.t18 a_n1808_13878.n17 3.61217
R22286 a_n1808_13878.n10 a_n1808_13878.n9 0.358259
R22287 a_n1808_13878.n13 a_n1808_13878.n11 0.358259
R22288 a_n1808_13878.n14 a_n1808_13878.n13 0.358259
R22289 a_n1808_13878.n16 a_n1808_13878.n2 0.358259
R22290 a_n1808_13878.n7 a_n1808_13878.n5 0.146627
R22291 a_n1808_13878.n11 a_n1808_13878.n10 0.101793
R22292 outputibias.n27 outputibias.n1 289.615
R22293 outputibias.n58 outputibias.n32 289.615
R22294 outputibias.n90 outputibias.n64 289.615
R22295 outputibias.n122 outputibias.n96 289.615
R22296 outputibias.n28 outputibias.n27 185
R22297 outputibias.n26 outputibias.n25 185
R22298 outputibias.n5 outputibias.n4 185
R22299 outputibias.n20 outputibias.n19 185
R22300 outputibias.n18 outputibias.n17 185
R22301 outputibias.n9 outputibias.n8 185
R22302 outputibias.n12 outputibias.n11 185
R22303 outputibias.n59 outputibias.n58 185
R22304 outputibias.n57 outputibias.n56 185
R22305 outputibias.n36 outputibias.n35 185
R22306 outputibias.n51 outputibias.n50 185
R22307 outputibias.n49 outputibias.n48 185
R22308 outputibias.n40 outputibias.n39 185
R22309 outputibias.n43 outputibias.n42 185
R22310 outputibias.n91 outputibias.n90 185
R22311 outputibias.n89 outputibias.n88 185
R22312 outputibias.n68 outputibias.n67 185
R22313 outputibias.n83 outputibias.n82 185
R22314 outputibias.n81 outputibias.n80 185
R22315 outputibias.n72 outputibias.n71 185
R22316 outputibias.n75 outputibias.n74 185
R22317 outputibias.n123 outputibias.n122 185
R22318 outputibias.n121 outputibias.n120 185
R22319 outputibias.n100 outputibias.n99 185
R22320 outputibias.n115 outputibias.n114 185
R22321 outputibias.n113 outputibias.n112 185
R22322 outputibias.n104 outputibias.n103 185
R22323 outputibias.n107 outputibias.n106 185
R22324 outputibias.n0 outputibias.t9 178.945
R22325 outputibias.n133 outputibias.t10 177.018
R22326 outputibias.n132 outputibias.t11 177.018
R22327 outputibias.n0 outputibias.t8 177.018
R22328 outputibias.t7 outputibias.n10 147.661
R22329 outputibias.t1 outputibias.n41 147.661
R22330 outputibias.t3 outputibias.n73 147.661
R22331 outputibias.t5 outputibias.n105 147.661
R22332 outputibias.n128 outputibias.t6 132.363
R22333 outputibias.n128 outputibias.t0 130.436
R22334 outputibias.n129 outputibias.t2 130.436
R22335 outputibias.n130 outputibias.t4 130.436
R22336 outputibias.n27 outputibias.n26 104.615
R22337 outputibias.n26 outputibias.n4 104.615
R22338 outputibias.n19 outputibias.n4 104.615
R22339 outputibias.n19 outputibias.n18 104.615
R22340 outputibias.n18 outputibias.n8 104.615
R22341 outputibias.n11 outputibias.n8 104.615
R22342 outputibias.n58 outputibias.n57 104.615
R22343 outputibias.n57 outputibias.n35 104.615
R22344 outputibias.n50 outputibias.n35 104.615
R22345 outputibias.n50 outputibias.n49 104.615
R22346 outputibias.n49 outputibias.n39 104.615
R22347 outputibias.n42 outputibias.n39 104.615
R22348 outputibias.n90 outputibias.n89 104.615
R22349 outputibias.n89 outputibias.n67 104.615
R22350 outputibias.n82 outputibias.n67 104.615
R22351 outputibias.n82 outputibias.n81 104.615
R22352 outputibias.n81 outputibias.n71 104.615
R22353 outputibias.n74 outputibias.n71 104.615
R22354 outputibias.n122 outputibias.n121 104.615
R22355 outputibias.n121 outputibias.n99 104.615
R22356 outputibias.n114 outputibias.n99 104.615
R22357 outputibias.n114 outputibias.n113 104.615
R22358 outputibias.n113 outputibias.n103 104.615
R22359 outputibias.n106 outputibias.n103 104.615
R22360 outputibias.n63 outputibias.n31 95.6354
R22361 outputibias.n63 outputibias.n62 94.6732
R22362 outputibias.n95 outputibias.n94 94.6732
R22363 outputibias.n127 outputibias.n126 94.6732
R22364 outputibias.n11 outputibias.t7 52.3082
R22365 outputibias.n42 outputibias.t1 52.3082
R22366 outputibias.n74 outputibias.t3 52.3082
R22367 outputibias.n106 outputibias.t5 52.3082
R22368 outputibias.n12 outputibias.n10 15.6674
R22369 outputibias.n43 outputibias.n41 15.6674
R22370 outputibias.n75 outputibias.n73 15.6674
R22371 outputibias.n107 outputibias.n105 15.6674
R22372 outputibias.n13 outputibias.n9 12.8005
R22373 outputibias.n44 outputibias.n40 12.8005
R22374 outputibias.n76 outputibias.n72 12.8005
R22375 outputibias.n108 outputibias.n104 12.8005
R22376 outputibias.n17 outputibias.n16 12.0247
R22377 outputibias.n48 outputibias.n47 12.0247
R22378 outputibias.n80 outputibias.n79 12.0247
R22379 outputibias.n112 outputibias.n111 12.0247
R22380 outputibias.n20 outputibias.n7 11.249
R22381 outputibias.n51 outputibias.n38 11.249
R22382 outputibias.n83 outputibias.n70 11.249
R22383 outputibias.n115 outputibias.n102 11.249
R22384 outputibias.n21 outputibias.n5 10.4732
R22385 outputibias.n52 outputibias.n36 10.4732
R22386 outputibias.n84 outputibias.n68 10.4732
R22387 outputibias.n116 outputibias.n100 10.4732
R22388 outputibias.n25 outputibias.n24 9.69747
R22389 outputibias.n56 outputibias.n55 9.69747
R22390 outputibias.n88 outputibias.n87 9.69747
R22391 outputibias.n120 outputibias.n119 9.69747
R22392 outputibias.n31 outputibias.n30 9.45567
R22393 outputibias.n62 outputibias.n61 9.45567
R22394 outputibias.n94 outputibias.n93 9.45567
R22395 outputibias.n126 outputibias.n125 9.45567
R22396 outputibias.n30 outputibias.n29 9.3005
R22397 outputibias.n3 outputibias.n2 9.3005
R22398 outputibias.n24 outputibias.n23 9.3005
R22399 outputibias.n22 outputibias.n21 9.3005
R22400 outputibias.n7 outputibias.n6 9.3005
R22401 outputibias.n16 outputibias.n15 9.3005
R22402 outputibias.n14 outputibias.n13 9.3005
R22403 outputibias.n61 outputibias.n60 9.3005
R22404 outputibias.n34 outputibias.n33 9.3005
R22405 outputibias.n55 outputibias.n54 9.3005
R22406 outputibias.n53 outputibias.n52 9.3005
R22407 outputibias.n38 outputibias.n37 9.3005
R22408 outputibias.n47 outputibias.n46 9.3005
R22409 outputibias.n45 outputibias.n44 9.3005
R22410 outputibias.n93 outputibias.n92 9.3005
R22411 outputibias.n66 outputibias.n65 9.3005
R22412 outputibias.n87 outputibias.n86 9.3005
R22413 outputibias.n85 outputibias.n84 9.3005
R22414 outputibias.n70 outputibias.n69 9.3005
R22415 outputibias.n79 outputibias.n78 9.3005
R22416 outputibias.n77 outputibias.n76 9.3005
R22417 outputibias.n125 outputibias.n124 9.3005
R22418 outputibias.n98 outputibias.n97 9.3005
R22419 outputibias.n119 outputibias.n118 9.3005
R22420 outputibias.n117 outputibias.n116 9.3005
R22421 outputibias.n102 outputibias.n101 9.3005
R22422 outputibias.n111 outputibias.n110 9.3005
R22423 outputibias.n109 outputibias.n108 9.3005
R22424 outputibias.n28 outputibias.n3 8.92171
R22425 outputibias.n59 outputibias.n34 8.92171
R22426 outputibias.n91 outputibias.n66 8.92171
R22427 outputibias.n123 outputibias.n98 8.92171
R22428 outputibias.n29 outputibias.n1 8.14595
R22429 outputibias.n60 outputibias.n32 8.14595
R22430 outputibias.n92 outputibias.n64 8.14595
R22431 outputibias.n124 outputibias.n96 8.14595
R22432 outputibias.n31 outputibias.n1 5.81868
R22433 outputibias.n62 outputibias.n32 5.81868
R22434 outputibias.n94 outputibias.n64 5.81868
R22435 outputibias.n126 outputibias.n96 5.81868
R22436 outputibias.n131 outputibias.n130 5.20947
R22437 outputibias.n29 outputibias.n28 5.04292
R22438 outputibias.n60 outputibias.n59 5.04292
R22439 outputibias.n92 outputibias.n91 5.04292
R22440 outputibias.n124 outputibias.n123 5.04292
R22441 outputibias.n131 outputibias.n127 4.42209
R22442 outputibias.n14 outputibias.n10 4.38594
R22443 outputibias.n45 outputibias.n41 4.38594
R22444 outputibias.n77 outputibias.n73 4.38594
R22445 outputibias.n109 outputibias.n105 4.38594
R22446 outputibias.n132 outputibias.n131 4.28454
R22447 outputibias.n25 outputibias.n3 4.26717
R22448 outputibias.n56 outputibias.n34 4.26717
R22449 outputibias.n88 outputibias.n66 4.26717
R22450 outputibias.n120 outputibias.n98 4.26717
R22451 outputibias.n24 outputibias.n5 3.49141
R22452 outputibias.n55 outputibias.n36 3.49141
R22453 outputibias.n87 outputibias.n68 3.49141
R22454 outputibias.n119 outputibias.n100 3.49141
R22455 outputibias.n21 outputibias.n20 2.71565
R22456 outputibias.n52 outputibias.n51 2.71565
R22457 outputibias.n84 outputibias.n83 2.71565
R22458 outputibias.n116 outputibias.n115 2.71565
R22459 outputibias.n17 outputibias.n7 1.93989
R22460 outputibias.n48 outputibias.n38 1.93989
R22461 outputibias.n80 outputibias.n70 1.93989
R22462 outputibias.n112 outputibias.n102 1.93989
R22463 outputibias.n130 outputibias.n129 1.9266
R22464 outputibias.n129 outputibias.n128 1.9266
R22465 outputibias.n133 outputibias.n132 1.92658
R22466 outputibias.n134 outputibias.n133 1.29913
R22467 outputibias.n16 outputibias.n9 1.16414
R22468 outputibias.n47 outputibias.n40 1.16414
R22469 outputibias.n79 outputibias.n72 1.16414
R22470 outputibias.n111 outputibias.n104 1.16414
R22471 outputibias.n127 outputibias.n95 0.962709
R22472 outputibias.n95 outputibias.n63 0.962709
R22473 outputibias.n13 outputibias.n12 0.388379
R22474 outputibias.n44 outputibias.n43 0.388379
R22475 outputibias.n76 outputibias.n75 0.388379
R22476 outputibias.n108 outputibias.n107 0.388379
R22477 outputibias.n134 outputibias.n0 0.337251
R22478 outputibias outputibias.n134 0.302375
R22479 outputibias.n30 outputibias.n2 0.155672
R22480 outputibias.n23 outputibias.n2 0.155672
R22481 outputibias.n23 outputibias.n22 0.155672
R22482 outputibias.n22 outputibias.n6 0.155672
R22483 outputibias.n15 outputibias.n6 0.155672
R22484 outputibias.n15 outputibias.n14 0.155672
R22485 outputibias.n61 outputibias.n33 0.155672
R22486 outputibias.n54 outputibias.n33 0.155672
R22487 outputibias.n54 outputibias.n53 0.155672
R22488 outputibias.n53 outputibias.n37 0.155672
R22489 outputibias.n46 outputibias.n37 0.155672
R22490 outputibias.n46 outputibias.n45 0.155672
R22491 outputibias.n93 outputibias.n65 0.155672
R22492 outputibias.n86 outputibias.n65 0.155672
R22493 outputibias.n86 outputibias.n85 0.155672
R22494 outputibias.n85 outputibias.n69 0.155672
R22495 outputibias.n78 outputibias.n69 0.155672
R22496 outputibias.n78 outputibias.n77 0.155672
R22497 outputibias.n125 outputibias.n97 0.155672
R22498 outputibias.n118 outputibias.n97 0.155672
R22499 outputibias.n118 outputibias.n117 0.155672
R22500 outputibias.n117 outputibias.n101 0.155672
R22501 outputibias.n110 outputibias.n101 0.155672
R22502 outputibias.n110 outputibias.n109 0.155672
R22503 plus.n46 plus.t9 252.611
R22504 plus.n9 plus.t11 252.611
R22505 plus.n76 plus.t4 243.97
R22506 plus.n72 plus.t12 231.093
R22507 plus.n35 plus.t7 231.093
R22508 plus.n76 plus.n75 223.454
R22509 plus.n78 plus.n77 223.454
R22510 plus.n47 plus.t5 187.445
R22511 plus.n44 plus.t18 187.445
R22512 plus.n42 plus.t17 187.445
R22513 plus.n59 plus.t13 187.445
R22514 plus.n65 plus.t14 187.445
R22515 plus.n38 plus.t10 187.445
R22516 plus.n1 plus.t6 187.445
R22517 plus.n28 plus.t16 187.445
R22518 plus.n22 plus.t15 187.445
R22519 plus.n5 plus.t20 187.445
R22520 plus.n7 plus.t19 187.445
R22521 plus.n10 plus.t8 187.445
R22522 plus.n73 plus.n72 161.3
R22523 plus.n71 plus.n37 161.3
R22524 plus.n70 plus.n69 161.3
R22525 plus.n68 plus.n67 161.3
R22526 plus.n66 plus.n39 161.3
R22527 plus.n64 plus.n63 161.3
R22528 plus.n62 plus.n40 161.3
R22529 plus.n61 plus.n60 161.3
R22530 plus.n58 plus.n41 161.3
R22531 plus.n57 plus.n56 161.3
R22532 plus.n55 plus.n54 161.3
R22533 plus.n53 plus.n43 161.3
R22534 plus.n52 plus.n51 161.3
R22535 plus.n50 plus.n49 161.3
R22536 plus.n48 plus.n45 161.3
R22537 plus.n11 plus.n8 161.3
R22538 plus.n13 plus.n12 161.3
R22539 plus.n15 plus.n14 161.3
R22540 plus.n16 plus.n6 161.3
R22541 plus.n18 plus.n17 161.3
R22542 plus.n20 plus.n19 161.3
R22543 plus.n21 plus.n4 161.3
R22544 plus.n24 plus.n23 161.3
R22545 plus.n25 plus.n3 161.3
R22546 plus.n27 plus.n26 161.3
R22547 plus.n29 plus.n2 161.3
R22548 plus.n31 plus.n30 161.3
R22549 plus.n33 plus.n32 161.3
R22550 plus.n34 plus.n0 161.3
R22551 plus.n36 plus.n35 161.3
R22552 plus.n49 plus.n48 56.5617
R22553 plus.n58 plus.n57 56.5617
R22554 plus.n67 plus.n66 56.5617
R22555 plus.n30 plus.n29 56.5617
R22556 plus.n21 plus.n20 56.5617
R22557 plus.n12 plus.n11 56.5617
R22558 plus.n71 plus.n70 46.3896
R22559 plus.n34 plus.n33 46.3896
R22560 plus.n46 plus.n45 42.8164
R22561 plus.n9 plus.n8 42.8164
R22562 plus.n54 plus.n53 42.5146
R22563 plus.n60 plus.n40 42.5146
R22564 plus.n23 plus.n3 42.5146
R22565 plus.n17 plus.n16 42.5146
R22566 plus.n53 plus.n52 38.6395
R22567 plus.n64 plus.n40 38.6395
R22568 plus.n27 plus.n3 38.6395
R22569 plus.n16 plus.n15 38.6395
R22570 plus.n47 plus.n46 38.2514
R22571 plus.n10 plus.n9 38.2514
R22572 plus.n74 plus.n73 31.491
R22573 plus.n49 plus.n44 19.9199
R22574 plus.n66 plus.n65 19.9199
R22575 plus.n29 plus.n28 19.9199
R22576 plus.n12 plus.n7 19.9199
R22577 plus.n75 plus.t1 19.8005
R22578 plus.n75 plus.t2 19.8005
R22579 plus.n77 plus.t0 19.8005
R22580 plus.n77 plus.t3 19.8005
R22581 plus.n57 plus.n42 17.9525
R22582 plus.n59 plus.n58 17.9525
R22583 plus.n22 plus.n21 17.9525
R22584 plus.n20 plus.n5 17.9525
R22585 plus.n48 plus.n47 15.9852
R22586 plus.n67 plus.n38 15.9852
R22587 plus.n30 plus.n1 15.9852
R22588 plus.n11 plus.n10 15.9852
R22589 plus.n72 plus.n71 15.3369
R22590 plus.n35 plus.n34 15.3369
R22591 plus plus.n79 14.7609
R22592 plus.n74 plus.n36 11.9494
R22593 plus.n70 plus.n38 8.60764
R22594 plus.n33 plus.n1 8.60764
R22595 plus.n54 plus.n42 6.6403
R22596 plus.n60 plus.n59 6.6403
R22597 plus.n23 plus.n22 6.6403
R22598 plus.n17 plus.n5 6.6403
R22599 plus.n79 plus.n78 5.40567
R22600 plus.n52 plus.n44 4.67295
R22601 plus.n65 plus.n64 4.67295
R22602 plus.n28 plus.n27 4.67295
R22603 plus.n15 plus.n7 4.67295
R22604 plus.n79 plus.n74 1.188
R22605 plus.n78 plus.n76 0.716017
R22606 plus.n50 plus.n45 0.189894
R22607 plus.n51 plus.n50 0.189894
R22608 plus.n51 plus.n43 0.189894
R22609 plus.n55 plus.n43 0.189894
R22610 plus.n56 plus.n55 0.189894
R22611 plus.n56 plus.n41 0.189894
R22612 plus.n61 plus.n41 0.189894
R22613 plus.n62 plus.n61 0.189894
R22614 plus.n63 plus.n62 0.189894
R22615 plus.n63 plus.n39 0.189894
R22616 plus.n68 plus.n39 0.189894
R22617 plus.n69 plus.n68 0.189894
R22618 plus.n69 plus.n37 0.189894
R22619 plus.n73 plus.n37 0.189894
R22620 plus.n36 plus.n0 0.189894
R22621 plus.n32 plus.n0 0.189894
R22622 plus.n32 plus.n31 0.189894
R22623 plus.n31 plus.n2 0.189894
R22624 plus.n26 plus.n2 0.189894
R22625 plus.n26 plus.n25 0.189894
R22626 plus.n25 plus.n24 0.189894
R22627 plus.n24 plus.n4 0.189894
R22628 plus.n19 plus.n4 0.189894
R22629 plus.n19 plus.n18 0.189894
R22630 plus.n18 plus.n6 0.189894
R22631 plus.n14 plus.n6 0.189894
R22632 plus.n14 plus.n13 0.189894
R22633 plus.n13 plus.n8 0.189894
R22634 a_n2903_n3924.n0 a_n2903_n3924.t36 214.981
R22635 a_n2903_n3924.n2 a_n2903_n3924.t12 214.452
R22636 a_n2903_n3924.n11 a_n2903_n3924.t37 214.321
R22637 a_n2903_n3924.n12 a_n2903_n3924.t35 214.321
R22638 a_n2903_n3924.n13 a_n2903_n3924.t11 214.321
R22639 a_n2903_n3924.n14 a_n2903_n3924.t38 214.321
R22640 a_n2903_n3924.n15 a_n2903_n3924.t8 214.321
R22641 a_n2903_n3924.n0 a_n2903_n3924.t13 214.321
R22642 a_n2903_n3924.n1 a_n2903_n3924.t26 55.8337
R22643 a_n2903_n3924.n3 a_n2903_n3924.t39 55.8337
R22644 a_n2903_n3924.n10 a_n2903_n3924.t6 55.8337
R22645 a_n2903_n3924.n34 a_n2903_n3924.t23 55.8335
R22646 a_n2903_n3924.n32 a_n2903_n3924.t10 55.8335
R22647 a_n2903_n3924.n25 a_n2903_n3924.t33 55.8335
R22648 a_n2903_n3924.n24 a_n2903_n3924.t24 55.8335
R22649 a_n2903_n3924.n17 a_n2903_n3924.t28 55.8335
R22650 a_n2903_n3924.n36 a_n2903_n3924.n35 53.0052
R22651 a_n2903_n3924.n38 a_n2903_n3924.n37 53.0052
R22652 a_n2903_n3924.n5 a_n2903_n3924.n4 53.0052
R22653 a_n2903_n3924.n7 a_n2903_n3924.n6 53.0052
R22654 a_n2903_n3924.n9 a_n2903_n3924.n8 53.0052
R22655 a_n2903_n3924.n31 a_n2903_n3924.n30 53.0051
R22656 a_n2903_n3924.n29 a_n2903_n3924.n28 53.0051
R22657 a_n2903_n3924.n27 a_n2903_n3924.n26 53.0051
R22658 a_n2903_n3924.n23 a_n2903_n3924.n22 53.0051
R22659 a_n2903_n3924.n21 a_n2903_n3924.n20 53.0051
R22660 a_n2903_n3924.n19 a_n2903_n3924.n18 53.0051
R22661 a_n2903_n3924.n40 a_n2903_n3924.n39 53.0051
R22662 a_n2903_n3924.n16 a_n2903_n3924.n10 12.2417
R22663 a_n2903_n3924.n34 a_n2903_n3924.n33 12.2417
R22664 a_n2903_n3924.n17 a_n2903_n3924.n16 5.16214
R22665 a_n2903_n3924.n33 a_n2903_n3924.n32 5.16214
R22666 a_n2903_n3924.n35 a_n2903_n3924.t21 2.82907
R22667 a_n2903_n3924.n35 a_n2903_n3924.t25 2.82907
R22668 a_n2903_n3924.n37 a_n2903_n3924.t18 2.82907
R22669 a_n2903_n3924.n37 a_n2903_n3924.t22 2.82907
R22670 a_n2903_n3924.n4 a_n2903_n3924.t0 2.82907
R22671 a_n2903_n3924.n4 a_n2903_n3924.t1 2.82907
R22672 a_n2903_n3924.n6 a_n2903_n3924.t3 2.82907
R22673 a_n2903_n3924.n6 a_n2903_n3924.t31 2.82907
R22674 a_n2903_n3924.n8 a_n2903_n3924.t32 2.82907
R22675 a_n2903_n3924.n8 a_n2903_n3924.t4 2.82907
R22676 a_n2903_n3924.n30 a_n2903_n3924.t14 2.82907
R22677 a_n2903_n3924.n30 a_n2903_n3924.t34 2.82907
R22678 a_n2903_n3924.n28 a_n2903_n3924.t9 2.82907
R22679 a_n2903_n3924.n28 a_n2903_n3924.t5 2.82907
R22680 a_n2903_n3924.n26 a_n2903_n3924.t7 2.82907
R22681 a_n2903_n3924.n26 a_n2903_n3924.t2 2.82907
R22682 a_n2903_n3924.n22 a_n2903_n3924.t16 2.82907
R22683 a_n2903_n3924.n22 a_n2903_n3924.t27 2.82907
R22684 a_n2903_n3924.n20 a_n2903_n3924.t20 2.82907
R22685 a_n2903_n3924.n20 a_n2903_n3924.t15 2.82907
R22686 a_n2903_n3924.n18 a_n2903_n3924.t29 2.82907
R22687 a_n2903_n3924.n18 a_n2903_n3924.t19 2.82907
R22688 a_n2903_n3924.t30 a_n2903_n3924.n40 2.82907
R22689 a_n2903_n3924.n40 a_n2903_n3924.t17 2.82907
R22690 a_n2903_n3924.n33 a_n2903_n3924.n2 1.95694
R22691 a_n2903_n3924.n16 a_n2903_n3924.n0 1.95694
R22692 a_n2903_n3924.n0 a_n2903_n3924.n15 0.684366
R22693 a_n2903_n3924.n15 a_n2903_n3924.n14 0.672012
R22694 a_n2903_n3924.n14 a_n2903_n3924.n13 0.672012
R22695 a_n2903_n3924.n13 a_n2903_n3924.n12 0.672012
R22696 a_n2903_n3924.n12 a_n2903_n3924.n11 0.672012
R22697 a_n2903_n3924.n11 a_n2903_n3924.n2 0.541924
R22698 a_n2903_n3924.n19 a_n2903_n3924.n17 0.530672
R22699 a_n2903_n3924.n21 a_n2903_n3924.n19 0.530672
R22700 a_n2903_n3924.n23 a_n2903_n3924.n21 0.530672
R22701 a_n2903_n3924.n24 a_n2903_n3924.n23 0.530672
R22702 a_n2903_n3924.n27 a_n2903_n3924.n25 0.530672
R22703 a_n2903_n3924.n29 a_n2903_n3924.n27 0.530672
R22704 a_n2903_n3924.n31 a_n2903_n3924.n29 0.530672
R22705 a_n2903_n3924.n32 a_n2903_n3924.n31 0.530672
R22706 a_n2903_n3924.n10 a_n2903_n3924.n9 0.530672
R22707 a_n2903_n3924.n9 a_n2903_n3924.n7 0.530672
R22708 a_n2903_n3924.n7 a_n2903_n3924.n5 0.530672
R22709 a_n2903_n3924.n5 a_n2903_n3924.n3 0.530672
R22710 a_n2903_n3924.n39 a_n2903_n3924.n1 0.530672
R22711 a_n2903_n3924.n39 a_n2903_n3924.n38 0.530672
R22712 a_n2903_n3924.n38 a_n2903_n3924.n36 0.530672
R22713 a_n2903_n3924.n36 a_n2903_n3924.n34 0.530672
R22714 a_n2903_n3924.n25 a_n2903_n3924.n24 0.235414
R22715 a_n2903_n3924.n3 a_n2903_n3924.n1 0.235414
R22716 a_n1986_8322.n6 a_n1986_8322.t5 74.6477
R22717 a_n1986_8322.n1 a_n1986_8322.t11 74.6477
R22718 a_n1986_8322.t20 a_n1986_8322.n18 74.6476
R22719 a_n1986_8322.n14 a_n1986_8322.t13 74.2899
R22720 a_n1986_8322.n7 a_n1986_8322.t3 74.2899
R22721 a_n1986_8322.n8 a_n1986_8322.t6 74.2899
R22722 a_n1986_8322.n11 a_n1986_8322.t7 74.2899
R22723 a_n1986_8322.n4 a_n1986_8322.t10 74.2899
R22724 a_n1986_8322.n18 a_n1986_8322.n17 70.6783
R22725 a_n1986_8322.n16 a_n1986_8322.n15 70.6783
R22726 a_n1986_8322.n6 a_n1986_8322.n5 70.6783
R22727 a_n1986_8322.n10 a_n1986_8322.n9 70.6783
R22728 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R22729 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R22730 a_n1986_8322.n12 a_n1986_8322.n4 22.7556
R22731 a_n1986_8322.n13 a_n1986_8322.t1 10.1306
R22732 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R22733 a_n1986_8322.n14 a_n1986_8322.n13 5.83671
R22734 a_n1986_8322.n13 a_n1986_8322.n12 5.3452
R22735 a_n1986_8322.n17 a_n1986_8322.t18 3.61217
R22736 a_n1986_8322.n17 a_n1986_8322.t15 3.61217
R22737 a_n1986_8322.n15 a_n1986_8322.t12 3.61217
R22738 a_n1986_8322.n15 a_n1986_8322.t21 3.61217
R22739 a_n1986_8322.n5 a_n1986_8322.t9 3.61217
R22740 a_n1986_8322.n5 a_n1986_8322.t8 3.61217
R22741 a_n1986_8322.n9 a_n1986_8322.t4 3.61217
R22742 a_n1986_8322.n9 a_n1986_8322.t2 3.61217
R22743 a_n1986_8322.n0 a_n1986_8322.t19 3.61217
R22744 a_n1986_8322.n0 a_n1986_8322.t14 3.61217
R22745 a_n1986_8322.n2 a_n1986_8322.t17 3.61217
R22746 a_n1986_8322.n2 a_n1986_8322.t16 3.61217
R22747 a_n1986_8322.n11 a_n1986_8322.n10 0.358259
R22748 a_n1986_8322.n10 a_n1986_8322.n8 0.358259
R22749 a_n1986_8322.n7 a_n1986_8322.n6 0.358259
R22750 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R22751 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R22752 a_n1986_8322.n16 a_n1986_8322.n14 0.358259
R22753 a_n1986_8322.n18 a_n1986_8322.n16 0.358259
R22754 a_n1986_8322.n8 a_n1986_8322.n7 0.101793
R22755 a_n1986_8322.t1 a_n1986_8322.t0 0.057021
R22756 minus.n46 minus.t20 252.611
R22757 minus.n9 minus.t13 252.611
R22758 minus.n78 minus.t3 243.255
R22759 minus.n72 minus.t15 231.093
R22760 minus.n35 minus.t17 231.093
R22761 minus.n77 minus.n75 224.169
R22762 minus.n77 minus.n76 223.454
R22763 minus.n38 minus.t12 187.445
R22764 minus.n65 minus.t7 187.445
R22765 minus.n59 minus.t6 187.445
R22766 minus.n42 minus.t11 187.445
R22767 minus.n44 minus.t10 187.445
R22768 minus.n47 minus.t16 187.445
R22769 minus.n10 minus.t9 187.445
R22770 minus.n7 minus.t8 187.445
R22771 minus.n5 minus.t5 187.445
R22772 minus.n22 minus.t18 187.445
R22773 minus.n28 minus.t19 187.445
R22774 minus.n1 minus.t14 187.445
R22775 minus.n48 minus.n45 161.3
R22776 minus.n50 minus.n49 161.3
R22777 minus.n52 minus.n51 161.3
R22778 minus.n53 minus.n43 161.3
R22779 minus.n55 minus.n54 161.3
R22780 minus.n57 minus.n56 161.3
R22781 minus.n58 minus.n41 161.3
R22782 minus.n61 minus.n60 161.3
R22783 minus.n62 minus.n40 161.3
R22784 minus.n64 minus.n63 161.3
R22785 minus.n66 minus.n39 161.3
R22786 minus.n68 minus.n67 161.3
R22787 minus.n70 minus.n69 161.3
R22788 minus.n71 minus.n37 161.3
R22789 minus.n73 minus.n72 161.3
R22790 minus.n36 minus.n35 161.3
R22791 minus.n34 minus.n0 161.3
R22792 minus.n33 minus.n32 161.3
R22793 minus.n31 minus.n30 161.3
R22794 minus.n29 minus.n2 161.3
R22795 minus.n27 minus.n26 161.3
R22796 minus.n25 minus.n3 161.3
R22797 minus.n24 minus.n23 161.3
R22798 minus.n21 minus.n4 161.3
R22799 minus.n20 minus.n19 161.3
R22800 minus.n18 minus.n17 161.3
R22801 minus.n16 minus.n6 161.3
R22802 minus.n15 minus.n14 161.3
R22803 minus.n13 minus.n12 161.3
R22804 minus.n11 minus.n8 161.3
R22805 minus.n67 minus.n66 56.5617
R22806 minus.n58 minus.n57 56.5617
R22807 minus.n49 minus.n48 56.5617
R22808 minus.n12 minus.n11 56.5617
R22809 minus.n21 minus.n20 56.5617
R22810 minus.n30 minus.n29 56.5617
R22811 minus.n71 minus.n70 46.3896
R22812 minus.n34 minus.n33 46.3896
R22813 minus.n46 minus.n45 42.8164
R22814 minus.n9 minus.n8 42.8164
R22815 minus.n60 minus.n40 42.5146
R22816 minus.n54 minus.n53 42.5146
R22817 minus.n17 minus.n16 42.5146
R22818 minus.n23 minus.n3 42.5146
R22819 minus.n64 minus.n40 38.6395
R22820 minus.n53 minus.n52 38.6395
R22821 minus.n16 minus.n15 38.6395
R22822 minus.n27 minus.n3 38.6395
R22823 minus.n47 minus.n46 38.2514
R22824 minus.n10 minus.n9 38.2514
R22825 minus.n74 minus.n73 31.7069
R22826 minus.n66 minus.n65 19.9199
R22827 minus.n49 minus.n44 19.9199
R22828 minus.n12 minus.n7 19.9199
R22829 minus.n29 minus.n28 19.9199
R22830 minus.n76 minus.t2 19.8005
R22831 minus.n76 minus.t0 19.8005
R22832 minus.n75 minus.t1 19.8005
R22833 minus.n75 minus.t4 19.8005
R22834 minus.n59 minus.n58 17.9525
R22835 minus.n57 minus.n42 17.9525
R22836 minus.n20 minus.n5 17.9525
R22837 minus.n22 minus.n21 17.9525
R22838 minus.n67 minus.n38 15.9852
R22839 minus.n48 minus.n47 15.9852
R22840 minus.n11 minus.n10 15.9852
R22841 minus.n30 minus.n1 15.9852
R22842 minus.n72 minus.n71 15.3369
R22843 minus.n35 minus.n34 15.3369
R22844 minus.n74 minus.n36 12.1653
R22845 minus minus.n79 11.8887
R22846 minus.n70 minus.n38 8.60764
R22847 minus.n33 minus.n1 8.60764
R22848 minus.n60 minus.n59 6.6403
R22849 minus.n54 minus.n42 6.6403
R22850 minus.n17 minus.n5 6.6403
R22851 minus.n23 minus.n22 6.6403
R22852 minus.n79 minus.n78 4.80222
R22853 minus.n65 minus.n64 4.67295
R22854 minus.n52 minus.n44 4.67295
R22855 minus.n15 minus.n7 4.67295
R22856 minus.n28 minus.n27 4.67295
R22857 minus.n79 minus.n74 0.972091
R22858 minus.n78 minus.n77 0.716017
R22859 minus.n73 minus.n37 0.189894
R22860 minus.n69 minus.n37 0.189894
R22861 minus.n69 minus.n68 0.189894
R22862 minus.n68 minus.n39 0.189894
R22863 minus.n63 minus.n39 0.189894
R22864 minus.n63 minus.n62 0.189894
R22865 minus.n62 minus.n61 0.189894
R22866 minus.n61 minus.n41 0.189894
R22867 minus.n56 minus.n41 0.189894
R22868 minus.n56 minus.n55 0.189894
R22869 minus.n55 minus.n43 0.189894
R22870 minus.n51 minus.n43 0.189894
R22871 minus.n51 minus.n50 0.189894
R22872 minus.n50 minus.n45 0.189894
R22873 minus.n13 minus.n8 0.189894
R22874 minus.n14 minus.n13 0.189894
R22875 minus.n14 minus.n6 0.189894
R22876 minus.n18 minus.n6 0.189894
R22877 minus.n19 minus.n18 0.189894
R22878 minus.n19 minus.n4 0.189894
R22879 minus.n24 minus.n4 0.189894
R22880 minus.n25 minus.n24 0.189894
R22881 minus.n26 minus.n25 0.189894
R22882 minus.n26 minus.n2 0.189894
R22883 minus.n31 minus.n2 0.189894
R22884 minus.n32 minus.n31 0.189894
R22885 minus.n32 minus.n0 0.189894
R22886 minus.n36 minus.n0 0.189894
R22887 output.n41 output.n15 289.615
R22888 output.n72 output.n46 289.615
R22889 output.n104 output.n78 289.615
R22890 output.n136 output.n110 289.615
R22891 output.n77 output.n45 197.26
R22892 output.n77 output.n76 196.298
R22893 output.n109 output.n108 196.298
R22894 output.n141 output.n140 196.298
R22895 output.n42 output.n41 185
R22896 output.n40 output.n39 185
R22897 output.n19 output.n18 185
R22898 output.n34 output.n33 185
R22899 output.n32 output.n31 185
R22900 output.n23 output.n22 185
R22901 output.n26 output.n25 185
R22902 output.n73 output.n72 185
R22903 output.n71 output.n70 185
R22904 output.n50 output.n49 185
R22905 output.n65 output.n64 185
R22906 output.n63 output.n62 185
R22907 output.n54 output.n53 185
R22908 output.n57 output.n56 185
R22909 output.n105 output.n104 185
R22910 output.n103 output.n102 185
R22911 output.n82 output.n81 185
R22912 output.n97 output.n96 185
R22913 output.n95 output.n94 185
R22914 output.n86 output.n85 185
R22915 output.n89 output.n88 185
R22916 output.n137 output.n136 185
R22917 output.n135 output.n134 185
R22918 output.n114 output.n113 185
R22919 output.n129 output.n128 185
R22920 output.n127 output.n126 185
R22921 output.n118 output.n117 185
R22922 output.n121 output.n120 185
R22923 output.t18 output.n24 147.661
R22924 output.t19 output.n55 147.661
R22925 output.t17 output.n87 147.661
R22926 output.t16 output.n119 147.661
R22927 output.n41 output.n40 104.615
R22928 output.n40 output.n18 104.615
R22929 output.n33 output.n18 104.615
R22930 output.n33 output.n32 104.615
R22931 output.n32 output.n22 104.615
R22932 output.n25 output.n22 104.615
R22933 output.n72 output.n71 104.615
R22934 output.n71 output.n49 104.615
R22935 output.n64 output.n49 104.615
R22936 output.n64 output.n63 104.615
R22937 output.n63 output.n53 104.615
R22938 output.n56 output.n53 104.615
R22939 output.n104 output.n103 104.615
R22940 output.n103 output.n81 104.615
R22941 output.n96 output.n81 104.615
R22942 output.n96 output.n95 104.615
R22943 output.n95 output.n85 104.615
R22944 output.n88 output.n85 104.615
R22945 output.n136 output.n135 104.615
R22946 output.n135 output.n113 104.615
R22947 output.n128 output.n113 104.615
R22948 output.n128 output.n127 104.615
R22949 output.n127 output.n117 104.615
R22950 output.n120 output.n117 104.615
R22951 output.n1 output.t10 77.056
R22952 output.n14 output.t11 76.6694
R22953 output.n1 output.n0 72.7095
R22954 output.n3 output.n2 72.7095
R22955 output.n5 output.n4 72.7095
R22956 output.n7 output.n6 72.7095
R22957 output.n9 output.n8 72.7095
R22958 output.n11 output.n10 72.7095
R22959 output.n13 output.n12 72.7095
R22960 output.n25 output.t18 52.3082
R22961 output.n56 output.t19 52.3082
R22962 output.n88 output.t17 52.3082
R22963 output.n120 output.t16 52.3082
R22964 output.n26 output.n24 15.6674
R22965 output.n57 output.n55 15.6674
R22966 output.n89 output.n87 15.6674
R22967 output.n121 output.n119 15.6674
R22968 output.n27 output.n23 12.8005
R22969 output.n58 output.n54 12.8005
R22970 output.n90 output.n86 12.8005
R22971 output.n122 output.n118 12.8005
R22972 output.n31 output.n30 12.0247
R22973 output.n62 output.n61 12.0247
R22974 output.n94 output.n93 12.0247
R22975 output.n126 output.n125 12.0247
R22976 output.n34 output.n21 11.249
R22977 output.n65 output.n52 11.249
R22978 output.n97 output.n84 11.249
R22979 output.n129 output.n116 11.249
R22980 output.n35 output.n19 10.4732
R22981 output.n66 output.n50 10.4732
R22982 output.n98 output.n82 10.4732
R22983 output.n130 output.n114 10.4732
R22984 output.n39 output.n38 9.69747
R22985 output.n70 output.n69 9.69747
R22986 output.n102 output.n101 9.69747
R22987 output.n134 output.n133 9.69747
R22988 output.n45 output.n44 9.45567
R22989 output.n76 output.n75 9.45567
R22990 output.n108 output.n107 9.45567
R22991 output.n140 output.n139 9.45567
R22992 output.n44 output.n43 9.3005
R22993 output.n17 output.n16 9.3005
R22994 output.n38 output.n37 9.3005
R22995 output.n36 output.n35 9.3005
R22996 output.n21 output.n20 9.3005
R22997 output.n30 output.n29 9.3005
R22998 output.n28 output.n27 9.3005
R22999 output.n75 output.n74 9.3005
R23000 output.n48 output.n47 9.3005
R23001 output.n69 output.n68 9.3005
R23002 output.n67 output.n66 9.3005
R23003 output.n52 output.n51 9.3005
R23004 output.n61 output.n60 9.3005
R23005 output.n59 output.n58 9.3005
R23006 output.n107 output.n106 9.3005
R23007 output.n80 output.n79 9.3005
R23008 output.n101 output.n100 9.3005
R23009 output.n99 output.n98 9.3005
R23010 output.n84 output.n83 9.3005
R23011 output.n93 output.n92 9.3005
R23012 output.n91 output.n90 9.3005
R23013 output.n139 output.n138 9.3005
R23014 output.n112 output.n111 9.3005
R23015 output.n133 output.n132 9.3005
R23016 output.n131 output.n130 9.3005
R23017 output.n116 output.n115 9.3005
R23018 output.n125 output.n124 9.3005
R23019 output.n123 output.n122 9.3005
R23020 output.n42 output.n17 8.92171
R23021 output.n73 output.n48 8.92171
R23022 output.n105 output.n80 8.92171
R23023 output.n137 output.n112 8.92171
R23024 output output.n141 8.15037
R23025 output.n43 output.n15 8.14595
R23026 output.n74 output.n46 8.14595
R23027 output.n106 output.n78 8.14595
R23028 output.n138 output.n110 8.14595
R23029 output.n45 output.n15 5.81868
R23030 output.n76 output.n46 5.81868
R23031 output.n108 output.n78 5.81868
R23032 output.n140 output.n110 5.81868
R23033 output.n43 output.n42 5.04292
R23034 output.n74 output.n73 5.04292
R23035 output.n106 output.n105 5.04292
R23036 output.n138 output.n137 5.04292
R23037 output.n28 output.n24 4.38594
R23038 output.n59 output.n55 4.38594
R23039 output.n91 output.n87 4.38594
R23040 output.n123 output.n119 4.38594
R23041 output.n39 output.n17 4.26717
R23042 output.n70 output.n48 4.26717
R23043 output.n102 output.n80 4.26717
R23044 output.n134 output.n112 4.26717
R23045 output.n0 output.t4 3.9605
R23046 output.n0 output.t2 3.9605
R23047 output.n2 output.t9 3.9605
R23048 output.n2 output.t12 3.9605
R23049 output.n4 output.t14 3.9605
R23050 output.n4 output.t6 3.9605
R23051 output.n6 output.t8 3.9605
R23052 output.n6 output.t15 3.9605
R23053 output.n8 output.t0 3.9605
R23054 output.n8 output.t5 3.9605
R23055 output.n10 output.t7 3.9605
R23056 output.n10 output.t13 3.9605
R23057 output.n12 output.t3 3.9605
R23058 output.n12 output.t1 3.9605
R23059 output.n38 output.n19 3.49141
R23060 output.n69 output.n50 3.49141
R23061 output.n101 output.n82 3.49141
R23062 output.n133 output.n114 3.49141
R23063 output.n35 output.n34 2.71565
R23064 output.n66 output.n65 2.71565
R23065 output.n98 output.n97 2.71565
R23066 output.n130 output.n129 2.71565
R23067 output.n31 output.n21 1.93989
R23068 output.n62 output.n52 1.93989
R23069 output.n94 output.n84 1.93989
R23070 output.n126 output.n116 1.93989
R23071 output.n30 output.n23 1.16414
R23072 output.n61 output.n54 1.16414
R23073 output.n93 output.n86 1.16414
R23074 output.n125 output.n118 1.16414
R23075 output.n141 output.n109 0.962709
R23076 output.n109 output.n77 0.962709
R23077 output.n27 output.n26 0.388379
R23078 output.n58 output.n57 0.388379
R23079 output.n90 output.n89 0.388379
R23080 output.n122 output.n121 0.388379
R23081 output.n14 output.n13 0.387128
R23082 output.n13 output.n11 0.387128
R23083 output.n11 output.n9 0.387128
R23084 output.n9 output.n7 0.387128
R23085 output.n7 output.n5 0.387128
R23086 output.n5 output.n3 0.387128
R23087 output.n3 output.n1 0.387128
R23088 output.n44 output.n16 0.155672
R23089 output.n37 output.n16 0.155672
R23090 output.n37 output.n36 0.155672
R23091 output.n36 output.n20 0.155672
R23092 output.n29 output.n20 0.155672
R23093 output.n29 output.n28 0.155672
R23094 output.n75 output.n47 0.155672
R23095 output.n68 output.n47 0.155672
R23096 output.n68 output.n67 0.155672
R23097 output.n67 output.n51 0.155672
R23098 output.n60 output.n51 0.155672
R23099 output.n60 output.n59 0.155672
R23100 output.n107 output.n79 0.155672
R23101 output.n100 output.n79 0.155672
R23102 output.n100 output.n99 0.155672
R23103 output.n99 output.n83 0.155672
R23104 output.n92 output.n83 0.155672
R23105 output.n92 output.n91 0.155672
R23106 output.n139 output.n111 0.155672
R23107 output.n132 output.n111 0.155672
R23108 output.n132 output.n131 0.155672
R23109 output.n131 output.n115 0.155672
R23110 output.n124 output.n115 0.155672
R23111 output.n124 output.n123 0.155672
R23112 output output.n14 0.126227
R23113 diffpairibias.n0 diffpairibias.t18 436.822
R23114 diffpairibias.n21 diffpairibias.t19 435.479
R23115 diffpairibias.n20 diffpairibias.t16 435.479
R23116 diffpairibias.n19 diffpairibias.t17 435.479
R23117 diffpairibias.n18 diffpairibias.t21 435.479
R23118 diffpairibias.n0 diffpairibias.t22 435.479
R23119 diffpairibias.n1 diffpairibias.t20 435.479
R23120 diffpairibias.n2 diffpairibias.t23 435.479
R23121 diffpairibias.n10 diffpairibias.t0 377.536
R23122 diffpairibias.n10 diffpairibias.t8 376.193
R23123 diffpairibias.n11 diffpairibias.t10 376.193
R23124 diffpairibias.n12 diffpairibias.t6 376.193
R23125 diffpairibias.n13 diffpairibias.t2 376.193
R23126 diffpairibias.n14 diffpairibias.t12 376.193
R23127 diffpairibias.n15 diffpairibias.t4 376.193
R23128 diffpairibias.n16 diffpairibias.t14 376.193
R23129 diffpairibias.n3 diffpairibias.t1 113.368
R23130 diffpairibias.n3 diffpairibias.t9 112.698
R23131 diffpairibias.n4 diffpairibias.t11 112.698
R23132 diffpairibias.n5 diffpairibias.t7 112.698
R23133 diffpairibias.n6 diffpairibias.t3 112.698
R23134 diffpairibias.n7 diffpairibias.t13 112.698
R23135 diffpairibias.n8 diffpairibias.t5 112.698
R23136 diffpairibias.n9 diffpairibias.t15 112.698
R23137 diffpairibias.n17 diffpairibias.n16 4.77242
R23138 diffpairibias.n17 diffpairibias.n9 4.30807
R23139 diffpairibias.n18 diffpairibias.n17 4.13945
R23140 diffpairibias.n16 diffpairibias.n15 1.34352
R23141 diffpairibias.n15 diffpairibias.n14 1.34352
R23142 diffpairibias.n14 diffpairibias.n13 1.34352
R23143 diffpairibias.n13 diffpairibias.n12 1.34352
R23144 diffpairibias.n12 diffpairibias.n11 1.34352
R23145 diffpairibias.n11 diffpairibias.n10 1.34352
R23146 diffpairibias.n2 diffpairibias.n1 1.34352
R23147 diffpairibias.n1 diffpairibias.n0 1.34352
R23148 diffpairibias.n19 diffpairibias.n18 1.34352
R23149 diffpairibias.n20 diffpairibias.n19 1.34352
R23150 diffpairibias.n21 diffpairibias.n20 1.34352
R23151 diffpairibias.n22 diffpairibias.n21 0.862419
R23152 diffpairibias diffpairibias.n22 0.684875
R23153 diffpairibias.n9 diffpairibias.n8 0.672012
R23154 diffpairibias.n8 diffpairibias.n7 0.672012
R23155 diffpairibias.n7 diffpairibias.n6 0.672012
R23156 diffpairibias.n6 diffpairibias.n5 0.672012
R23157 diffpairibias.n5 diffpairibias.n4 0.672012
R23158 diffpairibias.n4 diffpairibias.n3 0.672012
R23159 diffpairibias.n22 diffpairibias.n2 0.190907
C0 CSoutput outputibias 0.032386f
C1 vdd CSoutput 0.116309p
C2 minus diffpairibias 3.46e-19
C3 commonsourceibias output 0.006808f
C4 CSoutput minus 3.04887f
C5 vdd plus 0.081525f
C6 commonsourceibias outputibias 0.003832f
C7 plus diffpairibias 2.47e-19
C8 vdd commonsourceibias 0.004218f
C9 CSoutput plus 0.876783f
C10 commonsourceibias diffpairibias 0.052851f
C11 CSoutput commonsourceibias 44.9728f
C12 minus plus 9.55164f
C13 minus commonsourceibias 0.323289f
C14 plus commonsourceibias 0.277692f
C15 output outputibias 2.34152f
C16 vdd output 7.23429f
C17 CSoutput output 6.13571f
C18 diffpairibias gnd 48.96854f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.181391p
C22 plus gnd 33.576103f
C23 minus gnd 28.21859f
C24 CSoutput gnd 0.114582p
C25 vdd gnd 0.408747p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 output.t10 gnd 0.464308f
C74 output.t4 gnd 0.044422f
C75 output.t2 gnd 0.044422f
C76 output.n0 gnd 0.364624f
C77 output.n1 gnd 0.614102f
C78 output.t9 gnd 0.044422f
C79 output.t12 gnd 0.044422f
C80 output.n2 gnd 0.364624f
C81 output.n3 gnd 0.350265f
C82 output.t14 gnd 0.044422f
C83 output.t6 gnd 0.044422f
C84 output.n4 gnd 0.364624f
C85 output.n5 gnd 0.350265f
C86 output.t8 gnd 0.044422f
C87 output.t15 gnd 0.044422f
C88 output.n6 gnd 0.364624f
C89 output.n7 gnd 0.350265f
C90 output.t0 gnd 0.044422f
C91 output.t5 gnd 0.044422f
C92 output.n8 gnd 0.364624f
C93 output.n9 gnd 0.350265f
C94 output.t7 gnd 0.044422f
C95 output.t13 gnd 0.044422f
C96 output.n10 gnd 0.364624f
C97 output.n11 gnd 0.350265f
C98 output.t3 gnd 0.044422f
C99 output.t1 gnd 0.044422f
C100 output.n12 gnd 0.364624f
C101 output.n13 gnd 0.350265f
C102 output.t11 gnd 0.462979f
C103 output.n14 gnd 0.28994f
C104 output.n15 gnd 0.015803f
C105 output.n16 gnd 0.011243f
C106 output.n17 gnd 0.006041f
C107 output.n18 gnd 0.01428f
C108 output.n19 gnd 0.006397f
C109 output.n20 gnd 0.011243f
C110 output.n21 gnd 0.006041f
C111 output.n22 gnd 0.01428f
C112 output.n23 gnd 0.006397f
C113 output.n24 gnd 0.048111f
C114 output.t18 gnd 0.023274f
C115 output.n25 gnd 0.01071f
C116 output.n26 gnd 0.008435f
C117 output.n27 gnd 0.006041f
C118 output.n28 gnd 0.267512f
C119 output.n29 gnd 0.011243f
C120 output.n30 gnd 0.006041f
C121 output.n31 gnd 0.006397f
C122 output.n32 gnd 0.01428f
C123 output.n33 gnd 0.01428f
C124 output.n34 gnd 0.006397f
C125 output.n35 gnd 0.006041f
C126 output.n36 gnd 0.011243f
C127 output.n37 gnd 0.011243f
C128 output.n38 gnd 0.006041f
C129 output.n39 gnd 0.006397f
C130 output.n40 gnd 0.01428f
C131 output.n41 gnd 0.030913f
C132 output.n42 gnd 0.006397f
C133 output.n43 gnd 0.006041f
C134 output.n44 gnd 0.025987f
C135 output.n45 gnd 0.097665f
C136 output.n46 gnd 0.015803f
C137 output.n47 gnd 0.011243f
C138 output.n48 gnd 0.006041f
C139 output.n49 gnd 0.01428f
C140 output.n50 gnd 0.006397f
C141 output.n51 gnd 0.011243f
C142 output.n52 gnd 0.006041f
C143 output.n53 gnd 0.01428f
C144 output.n54 gnd 0.006397f
C145 output.n55 gnd 0.048111f
C146 output.t19 gnd 0.023274f
C147 output.n56 gnd 0.01071f
C148 output.n57 gnd 0.008435f
C149 output.n58 gnd 0.006041f
C150 output.n59 gnd 0.267512f
C151 output.n60 gnd 0.011243f
C152 output.n61 gnd 0.006041f
C153 output.n62 gnd 0.006397f
C154 output.n63 gnd 0.01428f
C155 output.n64 gnd 0.01428f
C156 output.n65 gnd 0.006397f
C157 output.n66 gnd 0.006041f
C158 output.n67 gnd 0.011243f
C159 output.n68 gnd 0.011243f
C160 output.n69 gnd 0.006041f
C161 output.n70 gnd 0.006397f
C162 output.n71 gnd 0.01428f
C163 output.n72 gnd 0.030913f
C164 output.n73 gnd 0.006397f
C165 output.n74 gnd 0.006041f
C166 output.n75 gnd 0.025987f
C167 output.n76 gnd 0.09306f
C168 output.n77 gnd 1.65264f
C169 output.n78 gnd 0.015803f
C170 output.n79 gnd 0.011243f
C171 output.n80 gnd 0.006041f
C172 output.n81 gnd 0.01428f
C173 output.n82 gnd 0.006397f
C174 output.n83 gnd 0.011243f
C175 output.n84 gnd 0.006041f
C176 output.n85 gnd 0.01428f
C177 output.n86 gnd 0.006397f
C178 output.n87 gnd 0.048111f
C179 output.t17 gnd 0.023274f
C180 output.n88 gnd 0.01071f
C181 output.n89 gnd 0.008435f
C182 output.n90 gnd 0.006041f
C183 output.n91 gnd 0.267512f
C184 output.n92 gnd 0.011243f
C185 output.n93 gnd 0.006041f
C186 output.n94 gnd 0.006397f
C187 output.n95 gnd 0.01428f
C188 output.n96 gnd 0.01428f
C189 output.n97 gnd 0.006397f
C190 output.n98 gnd 0.006041f
C191 output.n99 gnd 0.011243f
C192 output.n100 gnd 0.011243f
C193 output.n101 gnd 0.006041f
C194 output.n102 gnd 0.006397f
C195 output.n103 gnd 0.01428f
C196 output.n104 gnd 0.030913f
C197 output.n105 gnd 0.006397f
C198 output.n106 gnd 0.006041f
C199 output.n107 gnd 0.025987f
C200 output.n108 gnd 0.09306f
C201 output.n109 gnd 0.713089f
C202 output.n110 gnd 0.015803f
C203 output.n111 gnd 0.011243f
C204 output.n112 gnd 0.006041f
C205 output.n113 gnd 0.01428f
C206 output.n114 gnd 0.006397f
C207 output.n115 gnd 0.011243f
C208 output.n116 gnd 0.006041f
C209 output.n117 gnd 0.01428f
C210 output.n118 gnd 0.006397f
C211 output.n119 gnd 0.048111f
C212 output.t16 gnd 0.023274f
C213 output.n120 gnd 0.01071f
C214 output.n121 gnd 0.008435f
C215 output.n122 gnd 0.006041f
C216 output.n123 gnd 0.267512f
C217 output.n124 gnd 0.011243f
C218 output.n125 gnd 0.006041f
C219 output.n126 gnd 0.006397f
C220 output.n127 gnd 0.01428f
C221 output.n128 gnd 0.01428f
C222 output.n129 gnd 0.006397f
C223 output.n130 gnd 0.006041f
C224 output.n131 gnd 0.011243f
C225 output.n132 gnd 0.011243f
C226 output.n133 gnd 0.006041f
C227 output.n134 gnd 0.006397f
C228 output.n135 gnd 0.01428f
C229 output.n136 gnd 0.030913f
C230 output.n137 gnd 0.006397f
C231 output.n138 gnd 0.006041f
C232 output.n139 gnd 0.025987f
C233 output.n140 gnd 0.09306f
C234 output.n141 gnd 1.67353f
C235 minus.n0 gnd 0.02942f
C236 minus.t14 gnd 0.494688f
C237 minus.n1 gnd 0.200074f
C238 minus.n2 gnd 0.02942f
C239 minus.t19 gnd 0.494688f
C240 minus.n3 gnd 0.023912f
C241 minus.n4 gnd 0.02942f
C242 minus.t18 gnd 0.494688f
C243 minus.t5 gnd 0.494688f
C244 minus.n5 gnd 0.200074f
C245 minus.n6 gnd 0.02942f
C246 minus.t8 gnd 0.494688f
C247 minus.n7 gnd 0.200074f
C248 minus.n8 gnd 0.126287f
C249 minus.t9 gnd 0.494688f
C250 minus.t13 gnd 0.555405f
C251 minus.n9 gnd 0.232141f
C252 minus.n10 gnd 0.231054f
C253 minus.n11 gnd 0.036596f
C254 minus.n12 gnd 0.034393f
C255 minus.n13 gnd 0.02942f
C256 minus.n14 gnd 0.02942f
C257 minus.n15 gnd 0.036853f
C258 minus.n16 gnd 0.023912f
C259 minus.n17 gnd 0.037847f
C260 minus.n18 gnd 0.02942f
C261 minus.n19 gnd 0.02942f
C262 minus.n20 gnd 0.035494f
C263 minus.n21 gnd 0.035494f
C264 minus.n22 gnd 0.200074f
C265 minus.n23 gnd 0.037847f
C266 minus.n24 gnd 0.02942f
C267 minus.n25 gnd 0.02942f
C268 minus.n26 gnd 0.02942f
C269 minus.n27 gnd 0.036853f
C270 minus.n28 gnd 0.200074f
C271 minus.n29 gnd 0.034393f
C272 minus.n30 gnd 0.036596f
C273 minus.n31 gnd 0.02942f
C274 minus.n32 gnd 0.02942f
C275 minus.n33 gnd 0.038315f
C276 minus.n34 gnd 0.012185f
C277 minus.t17 gnd 0.535005f
C278 minus.n35 gnd 0.232377f
C279 minus.n36 gnd 0.345687f
C280 minus.n37 gnd 0.02942f
C281 minus.t15 gnd 0.535005f
C282 minus.t12 gnd 0.494688f
C283 minus.n38 gnd 0.200074f
C284 minus.n39 gnd 0.02942f
C285 minus.t7 gnd 0.494688f
C286 minus.n40 gnd 0.023912f
C287 minus.n41 gnd 0.02942f
C288 minus.t6 gnd 0.494688f
C289 minus.t11 gnd 0.494688f
C290 minus.n42 gnd 0.200074f
C291 minus.n43 gnd 0.02942f
C292 minus.t10 gnd 0.494688f
C293 minus.n44 gnd 0.200074f
C294 minus.n45 gnd 0.126287f
C295 minus.t16 gnd 0.494688f
C296 minus.t20 gnd 0.555405f
C297 minus.n46 gnd 0.232141f
C298 minus.n47 gnd 0.231054f
C299 minus.n48 gnd 0.036596f
C300 minus.n49 gnd 0.034393f
C301 minus.n50 gnd 0.02942f
C302 minus.n51 gnd 0.02942f
C303 minus.n52 gnd 0.036853f
C304 minus.n53 gnd 0.023912f
C305 minus.n54 gnd 0.037847f
C306 minus.n55 gnd 0.02942f
C307 minus.n56 gnd 0.02942f
C308 minus.n57 gnd 0.035494f
C309 minus.n58 gnd 0.035494f
C310 minus.n59 gnd 0.200074f
C311 minus.n60 gnd 0.037847f
C312 minus.n61 gnd 0.02942f
C313 minus.n62 gnd 0.02942f
C314 minus.n63 gnd 0.02942f
C315 minus.n64 gnd 0.036853f
C316 minus.n65 gnd 0.200074f
C317 minus.n66 gnd 0.034393f
C318 minus.n67 gnd 0.036596f
C319 minus.n68 gnd 0.02942f
C320 minus.n69 gnd 0.02942f
C321 minus.n70 gnd 0.038315f
C322 minus.n71 gnd 0.012185f
C323 minus.n72 gnd 0.232377f
C324 minus.n73 gnd 0.916705f
C325 minus.n74 gnd 1.37788f
C326 minus.t1 gnd 0.009069f
C327 minus.t4 gnd 0.009069f
C328 minus.n75 gnd 0.029822f
C329 minus.t2 gnd 0.009069f
C330 minus.t0 gnd 0.009069f
C331 minus.n76 gnd 0.029413f
C332 minus.n77 gnd 0.251028f
C333 minus.t3 gnd 0.050478f
C334 minus.n78 gnd 0.136984f
C335 minus.n79 gnd 2.0791f
C336 a_n1986_8322.t0 gnd 49.3545f
C337 a_n1986_8322.t1 gnd 76.194405f
C338 a_n1986_8322.t11 gnd 0.875731f
C339 a_n1986_8322.t19 gnd 0.093526f
C340 a_n1986_8322.t14 gnd 0.093526f
C341 a_n1986_8322.n0 gnd 0.658798f
C342 a_n1986_8322.n1 gnd 0.736109f
C343 a_n1986_8322.t17 gnd 0.093526f
C344 a_n1986_8322.t16 gnd 0.093526f
C345 a_n1986_8322.n2 gnd 0.658798f
C346 a_n1986_8322.n3 gnd 0.374008f
C347 a_n1986_8322.t10 gnd 0.873987f
C348 a_n1986_8322.n4 gnd 1.39886f
C349 a_n1986_8322.t5 gnd 0.875731f
C350 a_n1986_8322.t9 gnd 0.093526f
C351 a_n1986_8322.t8 gnd 0.093526f
C352 a_n1986_8322.n5 gnd 0.658798f
C353 a_n1986_8322.n6 gnd 0.736109f
C354 a_n1986_8322.t3 gnd 0.873987f
C355 a_n1986_8322.n7 gnd 0.37042f
C356 a_n1986_8322.t6 gnd 0.873987f
C357 a_n1986_8322.n8 gnd 0.37042f
C358 a_n1986_8322.t4 gnd 0.093526f
C359 a_n1986_8322.t2 gnd 0.093526f
C360 a_n1986_8322.n9 gnd 0.658798f
C361 a_n1986_8322.n10 gnd 0.374008f
C362 a_n1986_8322.t7 gnd 0.873987f
C363 a_n1986_8322.n11 gnd 0.872256f
C364 a_n1986_8322.n12 gnd 1.5906f
C365 a_n1986_8322.n13 gnd 3.77945f
C366 a_n1986_8322.t13 gnd 0.873987f
C367 a_n1986_8322.n14 gnd 0.766467f
C368 a_n1986_8322.t12 gnd 0.093526f
C369 a_n1986_8322.t21 gnd 0.093526f
C370 a_n1986_8322.n15 gnd 0.658798f
C371 a_n1986_8322.n16 gnd 0.374008f
C372 a_n1986_8322.t18 gnd 0.093526f
C373 a_n1986_8322.t15 gnd 0.093526f
C374 a_n1986_8322.n17 gnd 0.658798f
C375 a_n1986_8322.n18 gnd 0.736108f
C376 a_n1986_8322.t20 gnd 0.875732f
C377 a_n2903_n3924.n0 gnd 1.45586f
C378 a_n2903_n3924.t17 gnd 0.088483f
C379 a_n2903_n3924.t26 gnd 0.919619f
C380 a_n2903_n3924.n1 gnd 0.347657f
C381 a_n2903_n3924.t12 gnd 1.14306f
C382 a_n2903_n3924.n2 gnd 1.19083f
C383 a_n2903_n3924.t39 gnd 0.919619f
C384 a_n2903_n3924.n3 gnd 0.347657f
C385 a_n2903_n3924.t0 gnd 0.088483f
C386 a_n2903_n3924.t1 gnd 0.088483f
C387 a_n2903_n3924.n4 gnd 0.722655f
C388 a_n2903_n3924.n5 gnd 0.364177f
C389 a_n2903_n3924.t3 gnd 0.088483f
C390 a_n2903_n3924.t31 gnd 0.088483f
C391 a_n2903_n3924.n6 gnd 0.722655f
C392 a_n2903_n3924.n7 gnd 0.364177f
C393 a_n2903_n3924.t32 gnd 0.088483f
C394 a_n2903_n3924.t4 gnd 0.088483f
C395 a_n2903_n3924.n8 gnd 0.722655f
C396 a_n2903_n3924.n9 gnd 0.364177f
C397 a_n2903_n3924.t6 gnd 0.919619f
C398 a_n2903_n3924.n10 gnd 0.860834f
C399 a_n2903_n3924.t36 gnd 1.14419f
C400 a_n2903_n3924.t37 gnd 1.14261f
C401 a_n2903_n3924.n11 gnd 0.745791f
C402 a_n2903_n3924.t35 gnd 1.14261f
C403 a_n2903_n3924.n12 gnd 0.804756f
C404 a_n2903_n3924.t11 gnd 1.14261f
C405 a_n2903_n3924.n13 gnd 0.804756f
C406 a_n2903_n3924.t38 gnd 1.14261f
C407 a_n2903_n3924.n14 gnd 0.804756f
C408 a_n2903_n3924.t8 gnd 1.14261f
C409 a_n2903_n3924.n15 gnd 0.804756f
C410 a_n2903_n3924.t13 gnd 1.14261f
C411 a_n2903_n3924.n16 gnd 0.834168f
C412 a_n2903_n3924.t28 gnd 0.919616f
C413 a_n2903_n3924.n17 gnd 0.571219f
C414 a_n2903_n3924.t29 gnd 0.088483f
C415 a_n2903_n3924.t19 gnd 0.088483f
C416 a_n2903_n3924.n18 gnd 0.722654f
C417 a_n2903_n3924.n19 gnd 0.364178f
C418 a_n2903_n3924.t20 gnd 0.088483f
C419 a_n2903_n3924.t15 gnd 0.088483f
C420 a_n2903_n3924.n20 gnd 0.722654f
C421 a_n2903_n3924.n21 gnd 0.364178f
C422 a_n2903_n3924.t16 gnd 0.088483f
C423 a_n2903_n3924.t27 gnd 0.088483f
C424 a_n2903_n3924.n22 gnd 0.722654f
C425 a_n2903_n3924.n23 gnd 0.364178f
C426 a_n2903_n3924.t24 gnd 0.919616f
C427 a_n2903_n3924.n24 gnd 0.347661f
C428 a_n2903_n3924.t33 gnd 0.919616f
C429 a_n2903_n3924.n25 gnd 0.347661f
C430 a_n2903_n3924.t7 gnd 0.088483f
C431 a_n2903_n3924.t2 gnd 0.088483f
C432 a_n2903_n3924.n26 gnd 0.722654f
C433 a_n2903_n3924.n27 gnd 0.364178f
C434 a_n2903_n3924.t9 gnd 0.088483f
C435 a_n2903_n3924.t5 gnd 0.088483f
C436 a_n2903_n3924.n28 gnd 0.722654f
C437 a_n2903_n3924.n29 gnd 0.364178f
C438 a_n2903_n3924.t14 gnd 0.088483f
C439 a_n2903_n3924.t34 gnd 0.088483f
C440 a_n2903_n3924.n30 gnd 0.722654f
C441 a_n2903_n3924.n31 gnd 0.364178f
C442 a_n2903_n3924.t10 gnd 0.919616f
C443 a_n2903_n3924.n32 gnd 0.571219f
C444 a_n2903_n3924.n33 gnd 0.834168f
C445 a_n2903_n3924.t23 gnd 0.919616f
C446 a_n2903_n3924.n34 gnd 0.860837f
C447 a_n2903_n3924.t21 gnd 0.088483f
C448 a_n2903_n3924.t25 gnd 0.088483f
C449 a_n2903_n3924.n35 gnd 0.722655f
C450 a_n2903_n3924.n36 gnd 0.364177f
C451 a_n2903_n3924.t18 gnd 0.088483f
C452 a_n2903_n3924.t22 gnd 0.088483f
C453 a_n2903_n3924.n37 gnd 0.722655f
C454 a_n2903_n3924.n38 gnd 0.364177f
C455 a_n2903_n3924.n39 gnd 0.364176f
C456 a_n2903_n3924.n40 gnd 0.722656f
C457 a_n2903_n3924.t30 gnd 0.088483f
C458 plus.n0 gnd 0.021643f
C459 plus.t7 gnd 0.393587f
C460 plus.t6 gnd 0.363927f
C461 plus.n1 gnd 0.147188f
C462 plus.n2 gnd 0.021643f
C463 plus.t16 gnd 0.363927f
C464 plus.n3 gnd 0.017591f
C465 plus.n4 gnd 0.021643f
C466 plus.t15 gnd 0.363927f
C467 plus.t20 gnd 0.363927f
C468 plus.n5 gnd 0.147188f
C469 plus.n6 gnd 0.021643f
C470 plus.t19 gnd 0.363927f
C471 plus.n7 gnd 0.147188f
C472 plus.n8 gnd 0.092906f
C473 plus.t8 gnd 0.363927f
C474 plus.t11 gnd 0.408595f
C475 plus.n9 gnd 0.170779f
C476 plus.n10 gnd 0.16998f
C477 plus.n11 gnd 0.026922f
C478 plus.n12 gnd 0.025302f
C479 plus.n13 gnd 0.021643f
C480 plus.n14 gnd 0.021643f
C481 plus.n15 gnd 0.027112f
C482 plus.n16 gnd 0.017591f
C483 plus.n17 gnd 0.027843f
C484 plus.n18 gnd 0.021643f
C485 plus.n19 gnd 0.021643f
C486 plus.n20 gnd 0.026112f
C487 plus.n21 gnd 0.026112f
C488 plus.n22 gnd 0.147188f
C489 plus.n23 gnd 0.027843f
C490 plus.n24 gnd 0.021643f
C491 plus.n25 gnd 0.021643f
C492 plus.n26 gnd 0.021643f
C493 plus.n27 gnd 0.027112f
C494 plus.n28 gnd 0.147188f
C495 plus.n29 gnd 0.025302f
C496 plus.n30 gnd 0.026922f
C497 plus.n31 gnd 0.021643f
C498 plus.n32 gnd 0.021643f
C499 plus.n33 gnd 0.028188f
C500 plus.n34 gnd 0.008964f
C501 plus.n35 gnd 0.170953f
C502 plus.n36 gnd 0.248746f
C503 plus.n37 gnd 0.021643f
C504 plus.t10 gnd 0.363927f
C505 plus.n38 gnd 0.147188f
C506 plus.n39 gnd 0.021643f
C507 plus.t14 gnd 0.363927f
C508 plus.n40 gnd 0.017591f
C509 plus.n41 gnd 0.021643f
C510 plus.t13 gnd 0.363927f
C511 plus.t17 gnd 0.363927f
C512 plus.n42 gnd 0.147188f
C513 plus.n43 gnd 0.021643f
C514 plus.t18 gnd 0.363927f
C515 plus.n44 gnd 0.147188f
C516 plus.n45 gnd 0.092906f
C517 plus.t5 gnd 0.363927f
C518 plus.t9 gnd 0.408595f
C519 plus.n46 gnd 0.170779f
C520 plus.n47 gnd 0.16998f
C521 plus.n48 gnd 0.026922f
C522 plus.n49 gnd 0.025302f
C523 plus.n50 gnd 0.021643f
C524 plus.n51 gnd 0.021643f
C525 plus.n52 gnd 0.027112f
C526 plus.n53 gnd 0.017591f
C527 plus.n54 gnd 0.027843f
C528 plus.n55 gnd 0.021643f
C529 plus.n56 gnd 0.021643f
C530 plus.n57 gnd 0.026112f
C531 plus.n58 gnd 0.026112f
C532 plus.n59 gnd 0.147188f
C533 plus.n60 gnd 0.027843f
C534 plus.n61 gnd 0.021643f
C535 plus.n62 gnd 0.021643f
C536 plus.n63 gnd 0.021643f
C537 plus.n64 gnd 0.027112f
C538 plus.n65 gnd 0.147188f
C539 plus.n66 gnd 0.025302f
C540 plus.n67 gnd 0.026922f
C541 plus.n68 gnd 0.021643f
C542 plus.n69 gnd 0.021643f
C543 plus.n70 gnd 0.028188f
C544 plus.n71 gnd 0.008964f
C545 plus.t12 gnd 0.393587f
C546 plus.n72 gnd 0.170953f
C547 plus.n73 gnd 0.665721f
C548 plus.n74 gnd 1.00509f
C549 plus.t4 gnd 0.037363f
C550 plus.t1 gnd 0.006672f
C551 plus.t2 gnd 0.006672f
C552 plus.n75 gnd 0.021638f
C553 plus.n76 gnd 0.167981f
C554 plus.t0 gnd 0.006672f
C555 plus.t3 gnd 0.006672f
C556 plus.n77 gnd 0.021638f
C557 plus.n78 gnd 0.12609f
C558 plus.n79 gnd 2.65796f
C559 outputibias.t8 gnd 0.11477f
C560 outputibias.t9 gnd 0.115567f
C561 outputibias.n0 gnd 0.130108f
C562 outputibias.n1 gnd 0.001372f
C563 outputibias.n2 gnd 9.76e-19
C564 outputibias.n3 gnd 5.24e-19
C565 outputibias.n4 gnd 0.001239f
C566 outputibias.n5 gnd 5.55e-19
C567 outputibias.n6 gnd 9.76e-19
C568 outputibias.n7 gnd 5.24e-19
C569 outputibias.n8 gnd 0.001239f
C570 outputibias.n9 gnd 5.55e-19
C571 outputibias.n10 gnd 0.004176f
C572 outputibias.t7 gnd 0.00202f
C573 outputibias.n11 gnd 9.3e-19
C574 outputibias.n12 gnd 7.32e-19
C575 outputibias.n13 gnd 5.24e-19
C576 outputibias.n14 gnd 0.02322f
C577 outputibias.n15 gnd 9.76e-19
C578 outputibias.n16 gnd 5.24e-19
C579 outputibias.n17 gnd 5.55e-19
C580 outputibias.n18 gnd 0.001239f
C581 outputibias.n19 gnd 0.001239f
C582 outputibias.n20 gnd 5.55e-19
C583 outputibias.n21 gnd 5.24e-19
C584 outputibias.n22 gnd 9.76e-19
C585 outputibias.n23 gnd 9.76e-19
C586 outputibias.n24 gnd 5.24e-19
C587 outputibias.n25 gnd 5.55e-19
C588 outputibias.n26 gnd 0.001239f
C589 outputibias.n27 gnd 0.002683f
C590 outputibias.n28 gnd 5.55e-19
C591 outputibias.n29 gnd 5.24e-19
C592 outputibias.n30 gnd 0.002256f
C593 outputibias.n31 gnd 0.005781f
C594 outputibias.n32 gnd 0.001372f
C595 outputibias.n33 gnd 9.76e-19
C596 outputibias.n34 gnd 5.24e-19
C597 outputibias.n35 gnd 0.001239f
C598 outputibias.n36 gnd 5.55e-19
C599 outputibias.n37 gnd 9.76e-19
C600 outputibias.n38 gnd 5.24e-19
C601 outputibias.n39 gnd 0.001239f
C602 outputibias.n40 gnd 5.55e-19
C603 outputibias.n41 gnd 0.004176f
C604 outputibias.t1 gnd 0.00202f
C605 outputibias.n42 gnd 9.3e-19
C606 outputibias.n43 gnd 7.32e-19
C607 outputibias.n44 gnd 5.24e-19
C608 outputibias.n45 gnd 0.02322f
C609 outputibias.n46 gnd 9.76e-19
C610 outputibias.n47 gnd 5.24e-19
C611 outputibias.n48 gnd 5.55e-19
C612 outputibias.n49 gnd 0.001239f
C613 outputibias.n50 gnd 0.001239f
C614 outputibias.n51 gnd 5.55e-19
C615 outputibias.n52 gnd 5.24e-19
C616 outputibias.n53 gnd 9.76e-19
C617 outputibias.n54 gnd 9.76e-19
C618 outputibias.n55 gnd 5.24e-19
C619 outputibias.n56 gnd 5.55e-19
C620 outputibias.n57 gnd 0.001239f
C621 outputibias.n58 gnd 0.002683f
C622 outputibias.n59 gnd 5.55e-19
C623 outputibias.n60 gnd 5.24e-19
C624 outputibias.n61 gnd 0.002256f
C625 outputibias.n62 gnd 0.005197f
C626 outputibias.n63 gnd 0.121892f
C627 outputibias.n64 gnd 0.001372f
C628 outputibias.n65 gnd 9.76e-19
C629 outputibias.n66 gnd 5.24e-19
C630 outputibias.n67 gnd 0.001239f
C631 outputibias.n68 gnd 5.55e-19
C632 outputibias.n69 gnd 9.76e-19
C633 outputibias.n70 gnd 5.24e-19
C634 outputibias.n71 gnd 0.001239f
C635 outputibias.n72 gnd 5.55e-19
C636 outputibias.n73 gnd 0.004176f
C637 outputibias.t3 gnd 0.00202f
C638 outputibias.n74 gnd 9.3e-19
C639 outputibias.n75 gnd 7.32e-19
C640 outputibias.n76 gnd 5.24e-19
C641 outputibias.n77 gnd 0.02322f
C642 outputibias.n78 gnd 9.76e-19
C643 outputibias.n79 gnd 5.24e-19
C644 outputibias.n80 gnd 5.55e-19
C645 outputibias.n81 gnd 0.001239f
C646 outputibias.n82 gnd 0.001239f
C647 outputibias.n83 gnd 5.55e-19
C648 outputibias.n84 gnd 5.24e-19
C649 outputibias.n85 gnd 9.76e-19
C650 outputibias.n86 gnd 9.76e-19
C651 outputibias.n87 gnd 5.24e-19
C652 outputibias.n88 gnd 5.55e-19
C653 outputibias.n89 gnd 0.001239f
C654 outputibias.n90 gnd 0.002683f
C655 outputibias.n91 gnd 5.55e-19
C656 outputibias.n92 gnd 5.24e-19
C657 outputibias.n93 gnd 0.002256f
C658 outputibias.n94 gnd 0.005197f
C659 outputibias.n95 gnd 0.064513f
C660 outputibias.n96 gnd 0.001372f
C661 outputibias.n97 gnd 9.76e-19
C662 outputibias.n98 gnd 5.24e-19
C663 outputibias.n99 gnd 0.001239f
C664 outputibias.n100 gnd 5.55e-19
C665 outputibias.n101 gnd 9.76e-19
C666 outputibias.n102 gnd 5.24e-19
C667 outputibias.n103 gnd 0.001239f
C668 outputibias.n104 gnd 5.55e-19
C669 outputibias.n105 gnd 0.004176f
C670 outputibias.t5 gnd 0.00202f
C671 outputibias.n106 gnd 9.3e-19
C672 outputibias.n107 gnd 7.32e-19
C673 outputibias.n108 gnd 5.24e-19
C674 outputibias.n109 gnd 0.02322f
C675 outputibias.n110 gnd 9.76e-19
C676 outputibias.n111 gnd 5.24e-19
C677 outputibias.n112 gnd 5.55e-19
C678 outputibias.n113 gnd 0.001239f
C679 outputibias.n114 gnd 0.001239f
C680 outputibias.n115 gnd 5.55e-19
C681 outputibias.n116 gnd 5.24e-19
C682 outputibias.n117 gnd 9.76e-19
C683 outputibias.n118 gnd 9.76e-19
C684 outputibias.n119 gnd 5.24e-19
C685 outputibias.n120 gnd 5.55e-19
C686 outputibias.n121 gnd 0.001239f
C687 outputibias.n122 gnd 0.002683f
C688 outputibias.n123 gnd 5.55e-19
C689 outputibias.n124 gnd 5.24e-19
C690 outputibias.n125 gnd 0.002256f
C691 outputibias.n126 gnd 0.005197f
C692 outputibias.n127 gnd 0.084814f
C693 outputibias.t4 gnd 0.108319f
C694 outputibias.t2 gnd 0.108319f
C695 outputibias.t0 gnd 0.108319f
C696 outputibias.t6 gnd 0.109238f
C697 outputibias.n128 gnd 0.134674f
C698 outputibias.n129 gnd 0.07244f
C699 outputibias.n130 gnd 0.079818f
C700 outputibias.n131 gnd 0.164901f
C701 outputibias.t11 gnd 0.11477f
C702 outputibias.n132 gnd 0.067481f
C703 outputibias.t10 gnd 0.11477f
C704 outputibias.n133 gnd 0.065115f
C705 outputibias.n134 gnd 0.029159f
C706 a_n1808_13878.t17 gnd 0.185195f
C707 a_n1808_13878.t15 gnd 0.185195f
C708 a_n1808_13878.t19 gnd 0.185195f
C709 a_n1808_13878.n0 gnd 1.46067f
C710 a_n1808_13878.t8 gnd 0.185195f
C711 a_n1808_13878.t13 gnd 0.185195f
C712 a_n1808_13878.n1 gnd 1.45825f
C713 a_n1808_13878.n2 gnd 1.31079f
C714 a_n1808_13878.t10 gnd 0.185195f
C715 a_n1808_13878.t12 gnd 0.185195f
C716 a_n1808_13878.n3 gnd 1.4598f
C717 a_n1808_13878.t16 gnd 0.185195f
C718 a_n1808_13878.t11 gnd 0.185195f
C719 a_n1808_13878.n4 gnd 1.45825f
C720 a_n1808_13878.n5 gnd 2.03762f
C721 a_n1808_13878.t14 gnd 0.185195f
C722 a_n1808_13878.t9 gnd 0.185195f
C723 a_n1808_13878.n6 gnd 1.45825f
C724 a_n1808_13878.n7 gnd 3.69301f
C725 a_n1808_13878.t1 gnd 1.73408f
C726 a_n1808_13878.t4 gnd 0.185195f
C727 a_n1808_13878.t5 gnd 0.185195f
C728 a_n1808_13878.n8 gnd 1.30452f
C729 a_n1808_13878.n9 gnd 1.4576f
C730 a_n1808_13878.t0 gnd 1.73062f
C731 a_n1808_13878.n10 gnd 0.733487f
C732 a_n1808_13878.t3 gnd 1.73062f
C733 a_n1808_13878.n11 gnd 0.733487f
C734 a_n1808_13878.t6 gnd 0.185195f
C735 a_n1808_13878.t7 gnd 0.185195f
C736 a_n1808_13878.n12 gnd 1.30452f
C737 a_n1808_13878.n13 gnd 0.74059f
C738 a_n1808_13878.t2 gnd 1.73062f
C739 a_n1808_13878.n14 gnd 1.7272f
C740 a_n1808_13878.n15 gnd 2.51438f
C741 a_n1808_13878.n16 gnd 1.80025f
C742 a_n1808_13878.n17 gnd 1.45826f
C743 a_n1808_13878.t18 gnd 0.185195f
C744 a_n1986_13878.n0 gnd 2.75605f
C745 a_n1986_13878.n1 gnd 3.98159f
C746 a_n1986_13878.n2 gnd 3.8498f
C747 a_n1986_13878.n3 gnd 0.485058f
C748 a_n1986_13878.n4 gnd 0.654433f
C749 a_n1986_13878.n5 gnd 0.212692f
C750 a_n1986_13878.n6 gnd 0.278259f
C751 a_n1986_13878.n7 gnd 0.629578f
C752 a_n1986_13878.n8 gnd 0.278259f
C753 a_n1986_13878.n9 gnd 0.518119f
C754 a_n1986_13878.n10 gnd 0.20181f
C755 a_n1986_13878.n11 gnd 0.148637f
C756 a_n1986_13878.n12 gnd 0.233609f
C757 a_n1986_13878.n13 gnd 0.180436f
C758 a_n1986_13878.n14 gnd 0.20181f
C759 a_n1986_13878.n15 gnd 0.148637f
C760 a_n1986_13878.n16 gnd 0.571292f
C761 a_n1986_13878.n17 gnd 0.425782f
C762 a_n1986_13878.n18 gnd 0.212692f
C763 a_n1986_13878.n19 gnd 0.485058f
C764 a_n1986_13878.n20 gnd 0.278259f
C765 a_n1986_13878.n21 gnd 0.431885f
C766 a_n1986_13878.n22 gnd 0.212692f
C767 a_n1986_13878.n23 gnd 0.720523f
C768 a_n1986_13878.n24 gnd 0.278259f
C769 a_n1986_13878.n25 gnd 1.75107f
C770 a_n1986_13878.n26 gnd 1.16112f
C771 a_n1986_13878.n27 gnd 1.88684f
C772 a_n1986_13878.n28 gnd 3.1659f
C773 a_n1986_13878.n29 gnd 0.008235f
C774 a_n1986_13878.n31 gnd 0.281365f
C775 a_n1986_13878.n32 gnd 0.008235f
C776 a_n1986_13878.n34 gnd 0.281365f
C777 a_n1986_13878.n35 gnd 0.008235f
C778 a_n1986_13878.n36 gnd 0.280966f
C779 a_n1986_13878.n37 gnd 0.008235f
C780 a_n1986_13878.n38 gnd 0.280966f
C781 a_n1986_13878.n39 gnd 0.008235f
C782 a_n1986_13878.n40 gnd 0.280966f
C783 a_n1986_13878.n41 gnd 0.008235f
C784 a_n1986_13878.n42 gnd 1.3183f
C785 a_n1986_13878.n43 gnd 0.280966f
C786 a_n1986_13878.n44 gnd 0.106346f
C787 a_n1986_13878.n45 gnd 0.008235f
C788 a_n1986_13878.n47 gnd 0.008235f
C789 a_n1986_13878.n49 gnd 0.281365f
C790 a_n1986_13878.n50 gnd 0.281365f
C791 a_n1986_13878.t16 gnd 0.147525f
C792 a_n1986_13878.t10 gnd 1.38135f
C793 a_n1986_13878.t26 gnd 0.147525f
C794 a_n1986_13878.t22 gnd 0.147525f
C795 a_n1986_13878.n51 gnd 1.03917f
C796 a_n1986_13878.t15 gnd 0.686217f
C797 a_n1986_13878.n52 gnd 0.301704f
C798 a_n1986_13878.t7 gnd 0.686217f
C799 a_n1986_13878.t25 gnd 0.686217f
C800 a_n1986_13878.t48 gnd 0.686217f
C801 a_n1986_13878.n53 gnd 0.301704f
C802 a_n1986_13878.t57 gnd 0.686217f
C803 a_n1986_13878.t62 gnd 0.686217f
C804 a_n1986_13878.t11 gnd 0.700669f
C805 a_n1986_13878.t17 gnd 0.686217f
C806 a_n1986_13878.t13 gnd 0.686217f
C807 a_n1986_13878.t29 gnd 0.686217f
C808 a_n1986_13878.n54 gnd 0.301704f
C809 a_n1986_13878.t27 gnd 0.686217f
C810 a_n1986_13878.t19 gnd 0.697562f
C811 a_n1986_13878.t37 gnd 0.114742f
C812 a_n1986_13878.t31 gnd 0.114742f
C813 a_n1986_13878.n55 gnd 1.01689f
C814 a_n1986_13878.t2 gnd 0.114742f
C815 a_n1986_13878.t32 gnd 0.114742f
C816 a_n1986_13878.n56 gnd 1.0139f
C817 a_n1986_13878.t38 gnd 0.114742f
C818 a_n1986_13878.t33 gnd 0.114742f
C819 a_n1986_13878.n57 gnd 1.01689f
C820 a_n1986_13878.t5 gnd 0.114742f
C821 a_n1986_13878.t34 gnd 0.114742f
C822 a_n1986_13878.n58 gnd 1.0139f
C823 a_n1986_13878.t6 gnd 0.114742f
C824 a_n1986_13878.t36 gnd 0.114742f
C825 a_n1986_13878.n59 gnd 1.0139f
C826 a_n1986_13878.t4 gnd 0.114742f
C827 a_n1986_13878.t3 gnd 0.114742f
C828 a_n1986_13878.n60 gnd 1.0139f
C829 a_n1986_13878.t1 gnd 0.114742f
C830 a_n1986_13878.t39 gnd 0.114742f
C831 a_n1986_13878.n61 gnd 1.01689f
C832 a_n1986_13878.t35 gnd 0.114742f
C833 a_n1986_13878.t0 gnd 0.114742f
C834 a_n1986_13878.n62 gnd 1.0139f
C835 a_n1986_13878.t66 gnd 0.700669f
C836 a_n1986_13878.t49 gnd 0.686217f
C837 a_n1986_13878.t53 gnd 0.686217f
C838 a_n1986_13878.t43 gnd 0.686217f
C839 a_n1986_13878.n63 gnd 0.301704f
C840 a_n1986_13878.t58 gnd 0.686217f
C841 a_n1986_13878.t64 gnd 0.697562f
C842 a_n1986_13878.n64 gnd 0.304282f
C843 a_n1986_13878.n65 gnd 0.297873f
C844 a_n1986_13878.n66 gnd 0.304282f
C845 a_n1986_13878.n67 gnd 0.304282f
C846 a_n1986_13878.n68 gnd 0.297873f
C847 a_n1986_13878.n69 gnd 0.304282f
C848 a_n1986_13878.t20 gnd 1.38135f
C849 a_n1986_13878.t30 gnd 0.147525f
C850 a_n1986_13878.t28 gnd 0.147525f
C851 a_n1986_13878.n70 gnd 1.03917f
C852 a_n1986_13878.t18 gnd 0.147525f
C853 a_n1986_13878.t14 gnd 0.147525f
C854 a_n1986_13878.n71 gnd 1.03917f
C855 a_n1986_13878.t12 gnd 1.3786f
C856 a_n1986_13878.n72 gnd 1.12735f
C857 a_n1986_13878.n73 gnd 0.775089f
C858 a_n1986_13878.t47 gnd 0.686217f
C859 a_n1986_13878.t56 gnd 0.686217f
C860 a_n1986_13878.t67 gnd 0.686217f
C861 a_n1986_13878.n74 gnd 0.301704f
C862 a_n1986_13878.t59 gnd 0.686217f
C863 a_n1986_13878.t44 gnd 0.686217f
C864 a_n1986_13878.t45 gnd 0.686217f
C865 a_n1986_13878.n75 gnd 0.301704f
C866 a_n1986_13878.t63 gnd 0.686217f
C867 a_n1986_13878.t52 gnd 0.686217f
C868 a_n1986_13878.t51 gnd 0.686217f
C869 a_n1986_13878.n76 gnd 0.301704f
C870 a_n1986_13878.t55 gnd 0.686217f
C871 a_n1986_13878.t46 gnd 0.686217f
C872 a_n1986_13878.t40 gnd 0.686217f
C873 a_n1986_13878.n77 gnd 0.301704f
C874 a_n1986_13878.t60 gnd 0.697715f
C875 a_n1986_13878.n78 gnd 0.297873f
C876 a_n1986_13878.n79 gnd 0.292464f
C877 a_n1986_13878.t65 gnd 0.697715f
C878 a_n1986_13878.n80 gnd 0.297873f
C879 a_n1986_13878.n81 gnd 0.292464f
C880 a_n1986_13878.t54 gnd 0.697715f
C881 a_n1986_13878.n82 gnd 0.297873f
C882 a_n1986_13878.n83 gnd 0.292464f
C883 a_n1986_13878.t50 gnd 0.697715f
C884 a_n1986_13878.n84 gnd 0.297873f
C885 a_n1986_13878.n85 gnd 0.292464f
C886 a_n1986_13878.n86 gnd 0.991154f
C887 a_n1986_13878.t61 gnd 0.700669f
C888 a_n1986_13878.n87 gnd 0.304282f
C889 a_n1986_13878.t41 gnd 0.686217f
C890 a_n1986_13878.n88 gnd 0.297873f
C891 a_n1986_13878.n89 gnd 0.304282f
C892 a_n1986_13878.t42 gnd 0.697562f
C893 a_n1986_13878.t9 gnd 0.700669f
C894 a_n1986_13878.n90 gnd 0.304282f
C895 a_n1986_13878.t21 gnd 0.686217f
C896 a_n1986_13878.n91 gnd 0.297873f
C897 a_n1986_13878.n92 gnd 0.304282f
C898 a_n1986_13878.t23 gnd 0.697562f
C899 a_n1986_13878.n93 gnd 1.115f
C900 a_n1986_13878.t24 gnd 1.3786f
C901 a_n1986_13878.n94 gnd 1.03917f
C902 a_n1986_13878.t8 gnd 0.147525f
C903 vdd.t257 gnd 0.038364f
C904 vdd.t243 gnd 0.038364f
C905 vdd.n0 gnd 0.30258f
C906 vdd.t101 gnd 0.038364f
C907 vdd.t255 gnd 0.038364f
C908 vdd.n1 gnd 0.302081f
C909 vdd.n2 gnd 0.278576f
C910 vdd.t245 gnd 0.038364f
C911 vdd.t263 gnd 0.038364f
C912 vdd.n3 gnd 0.302081f
C913 vdd.n4 gnd 0.140886f
C914 vdd.t259 gnd 0.038364f
C915 vdd.t253 gnd 0.038364f
C916 vdd.n5 gnd 0.302081f
C917 vdd.n6 gnd 0.132196f
C918 vdd.t95 gnd 0.038364f
C919 vdd.t247 gnd 0.038364f
C920 vdd.n7 gnd 0.30258f
C921 vdd.t241 gnd 0.038364f
C922 vdd.t261 gnd 0.038364f
C923 vdd.n8 gnd 0.302081f
C924 vdd.n9 gnd 0.278576f
C925 vdd.t249 gnd 0.038364f
C926 vdd.t103 gnd 0.038364f
C927 vdd.n10 gnd 0.302081f
C928 vdd.n11 gnd 0.140886f
C929 vdd.t239 gnd 0.038364f
C930 vdd.t251 gnd 0.038364f
C931 vdd.n12 gnd 0.302081f
C932 vdd.n13 gnd 0.132196f
C933 vdd.n14 gnd 0.09346f
C934 vdd.t91 gnd 0.021313f
C935 vdd.t90 gnd 0.021313f
C936 vdd.n15 gnd 0.196178f
C937 vdd.t83 gnd 0.021313f
C938 vdd.t89 gnd 0.021313f
C939 vdd.n16 gnd 0.195604f
C940 vdd.n17 gnd 0.340413f
C941 vdd.t84 gnd 0.021313f
C942 vdd.t81 gnd 0.021313f
C943 vdd.n18 gnd 0.195604f
C944 vdd.n19 gnd 0.140833f
C945 vdd.t82 gnd 0.021313f
C946 vdd.t85 gnd 0.021313f
C947 vdd.n20 gnd 0.196178f
C948 vdd.t87 gnd 0.021313f
C949 vdd.t78 gnd 0.021313f
C950 vdd.n21 gnd 0.195604f
C951 vdd.n22 gnd 0.340413f
C952 vdd.t76 gnd 0.021313f
C953 vdd.t79 gnd 0.021313f
C954 vdd.n23 gnd 0.195604f
C955 vdd.n24 gnd 0.140833f
C956 vdd.t88 gnd 0.021313f
C957 vdd.t86 gnd 0.021313f
C958 vdd.n25 gnd 0.195604f
C959 vdd.t80 gnd 0.021313f
C960 vdd.t77 gnd 0.021313f
C961 vdd.n26 gnd 0.195604f
C962 vdd.n27 gnd 22.769402f
C963 vdd.n28 gnd 8.49977f
C964 vdd.n29 gnd 0.005813f
C965 vdd.n30 gnd 0.005394f
C966 vdd.n31 gnd 0.002984f
C967 vdd.n32 gnd 0.006851f
C968 vdd.n33 gnd 0.002899f
C969 vdd.n34 gnd 0.003069f
C970 vdd.n35 gnd 0.005394f
C971 vdd.n36 gnd 0.002899f
C972 vdd.n37 gnd 0.006851f
C973 vdd.n38 gnd 0.003069f
C974 vdd.n39 gnd 0.005394f
C975 vdd.n40 gnd 0.002899f
C976 vdd.n41 gnd 0.005138f
C977 vdd.n42 gnd 0.005154f
C978 vdd.t113 gnd 0.014719f
C979 vdd.n43 gnd 0.03275f
C980 vdd.n44 gnd 0.170439f
C981 vdd.n45 gnd 0.002899f
C982 vdd.n46 gnd 0.003069f
C983 vdd.n47 gnd 0.006851f
C984 vdd.n48 gnd 0.006851f
C985 vdd.n49 gnd 0.003069f
C986 vdd.n50 gnd 0.002899f
C987 vdd.n51 gnd 0.005394f
C988 vdd.n52 gnd 0.005394f
C989 vdd.n53 gnd 0.002899f
C990 vdd.n54 gnd 0.003069f
C991 vdd.n55 gnd 0.006851f
C992 vdd.n56 gnd 0.006851f
C993 vdd.n57 gnd 0.003069f
C994 vdd.n58 gnd 0.002899f
C995 vdd.n59 gnd 0.005394f
C996 vdd.n60 gnd 0.005394f
C997 vdd.n61 gnd 0.002899f
C998 vdd.n62 gnd 0.003069f
C999 vdd.n63 gnd 0.006851f
C1000 vdd.n64 gnd 0.006851f
C1001 vdd.n65 gnd 0.016198f
C1002 vdd.n66 gnd 0.002984f
C1003 vdd.n67 gnd 0.002899f
C1004 vdd.n68 gnd 0.013942f
C1005 vdd.n69 gnd 0.009734f
C1006 vdd.t223 gnd 0.034101f
C1007 vdd.t174 gnd 0.034101f
C1008 vdd.n70 gnd 0.234366f
C1009 vdd.n71 gnd 0.184293f
C1010 vdd.t235 gnd 0.034101f
C1011 vdd.t146 gnd 0.034101f
C1012 vdd.n72 gnd 0.234366f
C1013 vdd.n73 gnd 0.148723f
C1014 vdd.t212 gnd 0.034101f
C1015 vdd.t166 gnd 0.034101f
C1016 vdd.n74 gnd 0.234366f
C1017 vdd.n75 gnd 0.148723f
C1018 vdd.t230 gnd 0.034101f
C1019 vdd.t208 gnd 0.034101f
C1020 vdd.n76 gnd 0.234366f
C1021 vdd.n77 gnd 0.148723f
C1022 vdd.t121 gnd 0.034101f
C1023 vdd.t159 gnd 0.034101f
C1024 vdd.n78 gnd 0.234366f
C1025 vdd.n79 gnd 0.148723f
C1026 vdd.t131 gnd 0.034101f
C1027 vdd.t177 gnd 0.034101f
C1028 vdd.n80 gnd 0.234366f
C1029 vdd.n81 gnd 0.148723f
C1030 vdd.t154 gnd 0.034101f
C1031 vdd.t219 gnd 0.034101f
C1032 vdd.n82 gnd 0.234366f
C1033 vdd.n83 gnd 0.148723f
C1034 vdd.n84 gnd 0.005813f
C1035 vdd.n85 gnd 0.005394f
C1036 vdd.n86 gnd 0.002984f
C1037 vdd.n87 gnd 0.006851f
C1038 vdd.n88 gnd 0.002899f
C1039 vdd.n89 gnd 0.003069f
C1040 vdd.n90 gnd 0.005394f
C1041 vdd.n91 gnd 0.002899f
C1042 vdd.n92 gnd 0.006851f
C1043 vdd.n93 gnd 0.003069f
C1044 vdd.n94 gnd 0.005394f
C1045 vdd.n95 gnd 0.002899f
C1046 vdd.n96 gnd 0.005138f
C1047 vdd.n97 gnd 0.005154f
C1048 vdd.t136 gnd 0.014719f
C1049 vdd.n98 gnd 0.03275f
C1050 vdd.n99 gnd 0.170439f
C1051 vdd.n100 gnd 0.002899f
C1052 vdd.n101 gnd 0.003069f
C1053 vdd.n102 gnd 0.006851f
C1054 vdd.n103 gnd 0.006851f
C1055 vdd.n104 gnd 0.003069f
C1056 vdd.n105 gnd 0.002899f
C1057 vdd.n106 gnd 0.005394f
C1058 vdd.n107 gnd 0.005394f
C1059 vdd.n108 gnd 0.002899f
C1060 vdd.n109 gnd 0.003069f
C1061 vdd.n110 gnd 0.006851f
C1062 vdd.n111 gnd 0.006851f
C1063 vdd.n112 gnd 0.003069f
C1064 vdd.n113 gnd 0.002899f
C1065 vdd.n114 gnd 0.005394f
C1066 vdd.n115 gnd 0.005394f
C1067 vdd.n116 gnd 0.002899f
C1068 vdd.n117 gnd 0.003069f
C1069 vdd.n118 gnd 0.006851f
C1070 vdd.n119 gnd 0.006851f
C1071 vdd.n120 gnd 0.016198f
C1072 vdd.n121 gnd 0.002984f
C1073 vdd.n122 gnd 0.002899f
C1074 vdd.n123 gnd 0.013942f
C1075 vdd.n124 gnd 0.009428f
C1076 vdd.n125 gnd 0.110651f
C1077 vdd.n126 gnd 0.005813f
C1078 vdd.n127 gnd 0.005394f
C1079 vdd.n128 gnd 0.002984f
C1080 vdd.n129 gnd 0.006851f
C1081 vdd.n130 gnd 0.002899f
C1082 vdd.n131 gnd 0.003069f
C1083 vdd.n132 gnd 0.005394f
C1084 vdd.n133 gnd 0.002899f
C1085 vdd.n134 gnd 0.006851f
C1086 vdd.n135 gnd 0.003069f
C1087 vdd.n136 gnd 0.005394f
C1088 vdd.n137 gnd 0.002899f
C1089 vdd.n138 gnd 0.005138f
C1090 vdd.n139 gnd 0.005154f
C1091 vdd.t179 gnd 0.014719f
C1092 vdd.n140 gnd 0.03275f
C1093 vdd.n141 gnd 0.170439f
C1094 vdd.n142 gnd 0.002899f
C1095 vdd.n143 gnd 0.003069f
C1096 vdd.n144 gnd 0.006851f
C1097 vdd.n145 gnd 0.006851f
C1098 vdd.n146 gnd 0.003069f
C1099 vdd.n147 gnd 0.002899f
C1100 vdd.n148 gnd 0.005394f
C1101 vdd.n149 gnd 0.005394f
C1102 vdd.n150 gnd 0.002899f
C1103 vdd.n151 gnd 0.003069f
C1104 vdd.n152 gnd 0.006851f
C1105 vdd.n153 gnd 0.006851f
C1106 vdd.n154 gnd 0.003069f
C1107 vdd.n155 gnd 0.002899f
C1108 vdd.n156 gnd 0.005394f
C1109 vdd.n157 gnd 0.005394f
C1110 vdd.n158 gnd 0.002899f
C1111 vdd.n159 gnd 0.003069f
C1112 vdd.n160 gnd 0.006851f
C1113 vdd.n161 gnd 0.006851f
C1114 vdd.n162 gnd 0.016198f
C1115 vdd.n163 gnd 0.002984f
C1116 vdd.n164 gnd 0.002899f
C1117 vdd.n165 gnd 0.013942f
C1118 vdd.n166 gnd 0.009734f
C1119 vdd.t181 gnd 0.034101f
C1120 vdd.t203 gnd 0.034101f
C1121 vdd.n167 gnd 0.234366f
C1122 vdd.n168 gnd 0.184293f
C1123 vdd.t119 gnd 0.034101f
C1124 vdd.t172 gnd 0.034101f
C1125 vdd.n169 gnd 0.234366f
C1126 vdd.n170 gnd 0.148723f
C1127 vdd.t201 gnd 0.034101f
C1128 vdd.t111 gnd 0.034101f
C1129 vdd.n171 gnd 0.234366f
C1130 vdd.n172 gnd 0.148723f
C1131 vdd.t156 gnd 0.034101f
C1132 vdd.t158 gnd 0.034101f
C1133 vdd.n173 gnd 0.234366f
C1134 vdd.n174 gnd 0.148723f
C1135 vdd.t225 gnd 0.034101f
C1136 vdd.t151 gnd 0.034101f
C1137 vdd.n175 gnd 0.234366f
C1138 vdd.n176 gnd 0.148723f
C1139 vdd.t152 gnd 0.034101f
C1140 vdd.t221 gnd 0.034101f
C1141 vdd.n177 gnd 0.234366f
C1142 vdd.n178 gnd 0.148723f
C1143 vdd.t222 gnd 0.034101f
C1144 vdd.t129 gnd 0.034101f
C1145 vdd.n179 gnd 0.234366f
C1146 vdd.n180 gnd 0.148723f
C1147 vdd.n181 gnd 0.005813f
C1148 vdd.n182 gnd 0.005394f
C1149 vdd.n183 gnd 0.002984f
C1150 vdd.n184 gnd 0.006851f
C1151 vdd.n185 gnd 0.002899f
C1152 vdd.n186 gnd 0.003069f
C1153 vdd.n187 gnd 0.005394f
C1154 vdd.n188 gnd 0.002899f
C1155 vdd.n189 gnd 0.006851f
C1156 vdd.n190 gnd 0.003069f
C1157 vdd.n191 gnd 0.005394f
C1158 vdd.n192 gnd 0.002899f
C1159 vdd.n193 gnd 0.005138f
C1160 vdd.n194 gnd 0.005154f
C1161 vdd.t202 gnd 0.014719f
C1162 vdd.n195 gnd 0.03275f
C1163 vdd.n196 gnd 0.170439f
C1164 vdd.n197 gnd 0.002899f
C1165 vdd.n198 gnd 0.003069f
C1166 vdd.n199 gnd 0.006851f
C1167 vdd.n200 gnd 0.006851f
C1168 vdd.n201 gnd 0.003069f
C1169 vdd.n202 gnd 0.002899f
C1170 vdd.n203 gnd 0.005394f
C1171 vdd.n204 gnd 0.005394f
C1172 vdd.n205 gnd 0.002899f
C1173 vdd.n206 gnd 0.003069f
C1174 vdd.n207 gnd 0.006851f
C1175 vdd.n208 gnd 0.006851f
C1176 vdd.n209 gnd 0.003069f
C1177 vdd.n210 gnd 0.002899f
C1178 vdd.n211 gnd 0.005394f
C1179 vdd.n212 gnd 0.005394f
C1180 vdd.n213 gnd 0.002899f
C1181 vdd.n214 gnd 0.003069f
C1182 vdd.n215 gnd 0.006851f
C1183 vdd.n216 gnd 0.006851f
C1184 vdd.n217 gnd 0.016198f
C1185 vdd.n218 gnd 0.002984f
C1186 vdd.n219 gnd 0.002899f
C1187 vdd.n220 gnd 0.013942f
C1188 vdd.n221 gnd 0.009428f
C1189 vdd.n222 gnd 0.065826f
C1190 vdd.n223 gnd 0.237189f
C1191 vdd.n224 gnd 0.005813f
C1192 vdd.n225 gnd 0.005394f
C1193 vdd.n226 gnd 0.002984f
C1194 vdd.n227 gnd 0.006851f
C1195 vdd.n228 gnd 0.002899f
C1196 vdd.n229 gnd 0.003069f
C1197 vdd.n230 gnd 0.005394f
C1198 vdd.n231 gnd 0.002899f
C1199 vdd.n232 gnd 0.006851f
C1200 vdd.n233 gnd 0.003069f
C1201 vdd.n234 gnd 0.005394f
C1202 vdd.n235 gnd 0.002899f
C1203 vdd.n236 gnd 0.005138f
C1204 vdd.n237 gnd 0.005154f
C1205 vdd.t190 gnd 0.014719f
C1206 vdd.n238 gnd 0.03275f
C1207 vdd.n239 gnd 0.170439f
C1208 vdd.n240 gnd 0.002899f
C1209 vdd.n241 gnd 0.003069f
C1210 vdd.n242 gnd 0.006851f
C1211 vdd.n243 gnd 0.006851f
C1212 vdd.n244 gnd 0.003069f
C1213 vdd.n245 gnd 0.002899f
C1214 vdd.n246 gnd 0.005394f
C1215 vdd.n247 gnd 0.005394f
C1216 vdd.n248 gnd 0.002899f
C1217 vdd.n249 gnd 0.003069f
C1218 vdd.n250 gnd 0.006851f
C1219 vdd.n251 gnd 0.006851f
C1220 vdd.n252 gnd 0.003069f
C1221 vdd.n253 gnd 0.002899f
C1222 vdd.n254 gnd 0.005394f
C1223 vdd.n255 gnd 0.005394f
C1224 vdd.n256 gnd 0.002899f
C1225 vdd.n257 gnd 0.003069f
C1226 vdd.n258 gnd 0.006851f
C1227 vdd.n259 gnd 0.006851f
C1228 vdd.n260 gnd 0.016198f
C1229 vdd.n261 gnd 0.002984f
C1230 vdd.n262 gnd 0.002899f
C1231 vdd.n263 gnd 0.013942f
C1232 vdd.n264 gnd 0.009734f
C1233 vdd.t191 gnd 0.034101f
C1234 vdd.t216 gnd 0.034101f
C1235 vdd.n265 gnd 0.234366f
C1236 vdd.n266 gnd 0.184293f
C1237 vdd.t139 gnd 0.034101f
C1238 vdd.t189 gnd 0.034101f
C1239 vdd.n267 gnd 0.234366f
C1240 vdd.n268 gnd 0.148723f
C1241 vdd.t210 gnd 0.034101f
C1242 vdd.t134 gnd 0.034101f
C1243 vdd.n269 gnd 0.234366f
C1244 vdd.n270 gnd 0.148723f
C1245 vdd.t169 gnd 0.034101f
C1246 vdd.t171 gnd 0.034101f
C1247 vdd.n271 gnd 0.234366f
C1248 vdd.n272 gnd 0.148723f
C1249 vdd.t234 gnd 0.034101f
C1250 vdd.t164 gnd 0.034101f
C1251 vdd.n273 gnd 0.234366f
C1252 vdd.n274 gnd 0.148723f
C1253 vdd.t165 gnd 0.034101f
C1254 vdd.t232 gnd 0.034101f
C1255 vdd.n275 gnd 0.234366f
C1256 vdd.n276 gnd 0.148723f
C1257 vdd.t233 gnd 0.034101f
C1258 vdd.t144 gnd 0.034101f
C1259 vdd.n277 gnd 0.234366f
C1260 vdd.n278 gnd 0.148723f
C1261 vdd.n279 gnd 0.005813f
C1262 vdd.n280 gnd 0.005394f
C1263 vdd.n281 gnd 0.002984f
C1264 vdd.n282 gnd 0.006851f
C1265 vdd.n283 gnd 0.002899f
C1266 vdd.n284 gnd 0.003069f
C1267 vdd.n285 gnd 0.005394f
C1268 vdd.n286 gnd 0.002899f
C1269 vdd.n287 gnd 0.006851f
C1270 vdd.n288 gnd 0.003069f
C1271 vdd.n289 gnd 0.005394f
C1272 vdd.n290 gnd 0.002899f
C1273 vdd.n291 gnd 0.005138f
C1274 vdd.n292 gnd 0.005154f
C1275 vdd.t214 gnd 0.014719f
C1276 vdd.n293 gnd 0.03275f
C1277 vdd.n294 gnd 0.170439f
C1278 vdd.n295 gnd 0.002899f
C1279 vdd.n296 gnd 0.003069f
C1280 vdd.n297 gnd 0.006851f
C1281 vdd.n298 gnd 0.006851f
C1282 vdd.n299 gnd 0.003069f
C1283 vdd.n300 gnd 0.002899f
C1284 vdd.n301 gnd 0.005394f
C1285 vdd.n302 gnd 0.005394f
C1286 vdd.n303 gnd 0.002899f
C1287 vdd.n304 gnd 0.003069f
C1288 vdd.n305 gnd 0.006851f
C1289 vdd.n306 gnd 0.006851f
C1290 vdd.n307 gnd 0.003069f
C1291 vdd.n308 gnd 0.002899f
C1292 vdd.n309 gnd 0.005394f
C1293 vdd.n310 gnd 0.005394f
C1294 vdd.n311 gnd 0.002899f
C1295 vdd.n312 gnd 0.003069f
C1296 vdd.n313 gnd 0.006851f
C1297 vdd.n314 gnd 0.006851f
C1298 vdd.n315 gnd 0.016198f
C1299 vdd.n316 gnd 0.002984f
C1300 vdd.n317 gnd 0.002899f
C1301 vdd.n318 gnd 0.013942f
C1302 vdd.n319 gnd 0.009428f
C1303 vdd.n320 gnd 0.065826f
C1304 vdd.n321 gnd 0.26562f
C1305 vdd.n322 gnd 0.008141f
C1306 vdd.n323 gnd 0.010592f
C1307 vdd.n324 gnd 0.008525f
C1308 vdd.n325 gnd 0.008525f
C1309 vdd.n326 gnd 0.010592f
C1310 vdd.n327 gnd 0.010592f
C1311 vdd.n328 gnd 0.773951f
C1312 vdd.n329 gnd 0.010592f
C1313 vdd.n330 gnd 0.010592f
C1314 vdd.n331 gnd 0.010592f
C1315 vdd.n332 gnd 0.838898f
C1316 vdd.n333 gnd 0.010592f
C1317 vdd.n334 gnd 0.010592f
C1318 vdd.n335 gnd 0.010592f
C1319 vdd.n336 gnd 0.010592f
C1320 vdd.n337 gnd 0.008525f
C1321 vdd.n338 gnd 0.010592f
C1322 vdd.t150 gnd 0.541225f
C1323 vdd.n339 gnd 0.010592f
C1324 vdd.n340 gnd 0.010592f
C1325 vdd.n341 gnd 0.010592f
C1326 vdd.t176 gnd 0.541225f
C1327 vdd.n342 gnd 0.010592f
C1328 vdd.n343 gnd 0.010592f
C1329 vdd.n344 gnd 0.010592f
C1330 vdd.n345 gnd 0.010592f
C1331 vdd.n346 gnd 0.010592f
C1332 vdd.n347 gnd 0.008525f
C1333 vdd.n348 gnd 0.010592f
C1334 vdd.n349 gnd 0.611584f
C1335 vdd.n350 gnd 0.010592f
C1336 vdd.n351 gnd 0.010592f
C1337 vdd.n352 gnd 0.010592f
C1338 vdd.t128 gnd 0.541225f
C1339 vdd.n353 gnd 0.010592f
C1340 vdd.n354 gnd 0.010592f
C1341 vdd.n355 gnd 0.010592f
C1342 vdd.n356 gnd 0.010592f
C1343 vdd.n357 gnd 0.010592f
C1344 vdd.n358 gnd 0.008525f
C1345 vdd.n359 gnd 0.010592f
C1346 vdd.t135 gnd 0.541225f
C1347 vdd.n360 gnd 0.010592f
C1348 vdd.n361 gnd 0.010592f
C1349 vdd.n362 gnd 0.010592f
C1350 vdd.n363 gnd 0.91467f
C1351 vdd.n364 gnd 0.010592f
C1352 vdd.n365 gnd 0.010592f
C1353 vdd.n366 gnd 0.010592f
C1354 vdd.n367 gnd 0.010592f
C1355 vdd.n368 gnd 0.010592f
C1356 vdd.n369 gnd 0.007076f
C1357 vdd.n370 gnd 0.02412f
C1358 vdd.t9 gnd 0.541225f
C1359 vdd.n371 gnd 0.010592f
C1360 vdd.n372 gnd 0.02412f
C1361 vdd.n404 gnd 0.010592f
C1362 vdd.t11 gnd 0.130309f
C1363 vdd.t10 gnd 0.139265f
C1364 vdd.t8 gnd 0.170182f
C1365 vdd.n405 gnd 0.218149f
C1366 vdd.n406 gnd 0.184137f
C1367 vdd.n407 gnd 0.013981f
C1368 vdd.n408 gnd 0.010592f
C1369 vdd.n409 gnd 0.008525f
C1370 vdd.n410 gnd 0.010592f
C1371 vdd.n411 gnd 0.008525f
C1372 vdd.n412 gnd 0.010592f
C1373 vdd.n413 gnd 0.008525f
C1374 vdd.n414 gnd 0.010592f
C1375 vdd.n415 gnd 0.008525f
C1376 vdd.n416 gnd 0.010592f
C1377 vdd.n417 gnd 0.008525f
C1378 vdd.n418 gnd 0.010592f
C1379 vdd.t69 gnd 0.130309f
C1380 vdd.t68 gnd 0.139265f
C1381 vdd.t67 gnd 0.170182f
C1382 vdd.n419 gnd 0.218149f
C1383 vdd.n420 gnd 0.184137f
C1384 vdd.n421 gnd 0.008525f
C1385 vdd.n422 gnd 0.010592f
C1386 vdd.n423 gnd 0.008525f
C1387 vdd.n424 gnd 0.010592f
C1388 vdd.n425 gnd 0.008525f
C1389 vdd.n426 gnd 0.010592f
C1390 vdd.n427 gnd 0.008525f
C1391 vdd.n428 gnd 0.010592f
C1392 vdd.n429 gnd 0.008525f
C1393 vdd.n430 gnd 0.010592f
C1394 vdd.t75 gnd 0.130309f
C1395 vdd.t74 gnd 0.139265f
C1396 vdd.t73 gnd 0.170182f
C1397 vdd.n431 gnd 0.218149f
C1398 vdd.n432 gnd 0.184137f
C1399 vdd.n433 gnd 0.018244f
C1400 vdd.n434 gnd 0.010592f
C1401 vdd.n435 gnd 0.008525f
C1402 vdd.n436 gnd 0.010592f
C1403 vdd.n437 gnd 0.008525f
C1404 vdd.n438 gnd 0.010592f
C1405 vdd.n439 gnd 0.008525f
C1406 vdd.n440 gnd 0.010592f
C1407 vdd.n441 gnd 0.008525f
C1408 vdd.n442 gnd 0.010592f
C1409 vdd.n443 gnd 0.02412f
C1410 vdd.n444 gnd 0.024285f
C1411 vdd.n445 gnd 0.024285f
C1412 vdd.n446 gnd 0.007076f
C1413 vdd.n447 gnd 0.008525f
C1414 vdd.n448 gnd 0.010592f
C1415 vdd.n449 gnd 0.010592f
C1416 vdd.n450 gnd 0.008525f
C1417 vdd.n451 gnd 0.010592f
C1418 vdd.n452 gnd 0.010592f
C1419 vdd.n453 gnd 0.010592f
C1420 vdd.n454 gnd 0.010592f
C1421 vdd.n455 gnd 0.010592f
C1422 vdd.n456 gnd 0.008525f
C1423 vdd.n457 gnd 0.008525f
C1424 vdd.n458 gnd 0.010592f
C1425 vdd.n459 gnd 0.010592f
C1426 vdd.n460 gnd 0.008525f
C1427 vdd.n461 gnd 0.010592f
C1428 vdd.n462 gnd 0.010592f
C1429 vdd.n463 gnd 0.010592f
C1430 vdd.n464 gnd 0.010592f
C1431 vdd.n465 gnd 0.010592f
C1432 vdd.n466 gnd 0.008525f
C1433 vdd.n467 gnd 0.008525f
C1434 vdd.n468 gnd 0.010592f
C1435 vdd.n469 gnd 0.010592f
C1436 vdd.n470 gnd 0.008525f
C1437 vdd.n471 gnd 0.010592f
C1438 vdd.n472 gnd 0.010592f
C1439 vdd.n473 gnd 0.010592f
C1440 vdd.n474 gnd 0.010592f
C1441 vdd.n475 gnd 0.010592f
C1442 vdd.n476 gnd 0.008525f
C1443 vdd.n477 gnd 0.008525f
C1444 vdd.n478 gnd 0.010592f
C1445 vdd.n479 gnd 0.010592f
C1446 vdd.n480 gnd 0.008525f
C1447 vdd.n481 gnd 0.010592f
C1448 vdd.n482 gnd 0.010592f
C1449 vdd.n483 gnd 0.010592f
C1450 vdd.n484 gnd 0.010592f
C1451 vdd.n485 gnd 0.010592f
C1452 vdd.n486 gnd 0.008525f
C1453 vdd.n487 gnd 0.008525f
C1454 vdd.n488 gnd 0.010592f
C1455 vdd.n489 gnd 0.010592f
C1456 vdd.n490 gnd 0.007119f
C1457 vdd.n491 gnd 0.010592f
C1458 vdd.n492 gnd 0.010592f
C1459 vdd.n493 gnd 0.010592f
C1460 vdd.n494 gnd 0.010592f
C1461 vdd.n495 gnd 0.010592f
C1462 vdd.n496 gnd 0.007119f
C1463 vdd.n497 gnd 0.008525f
C1464 vdd.n498 gnd 0.010592f
C1465 vdd.n499 gnd 0.010592f
C1466 vdd.n500 gnd 0.008525f
C1467 vdd.n501 gnd 0.010592f
C1468 vdd.n502 gnd 0.010592f
C1469 vdd.n503 gnd 0.010592f
C1470 vdd.n504 gnd 0.010592f
C1471 vdd.n505 gnd 0.010592f
C1472 vdd.n506 gnd 0.008525f
C1473 vdd.n507 gnd 0.008525f
C1474 vdd.n508 gnd 0.010592f
C1475 vdd.n509 gnd 0.010592f
C1476 vdd.n510 gnd 0.008525f
C1477 vdd.n511 gnd 0.010592f
C1478 vdd.n512 gnd 0.010592f
C1479 vdd.n513 gnd 0.010592f
C1480 vdd.n514 gnd 0.010592f
C1481 vdd.n515 gnd 0.010592f
C1482 vdd.n516 gnd 0.008525f
C1483 vdd.n517 gnd 0.008525f
C1484 vdd.n518 gnd 0.010592f
C1485 vdd.n519 gnd 0.010592f
C1486 vdd.n520 gnd 0.008525f
C1487 vdd.n521 gnd 0.010592f
C1488 vdd.n522 gnd 0.010592f
C1489 vdd.n523 gnd 0.010592f
C1490 vdd.n524 gnd 0.010592f
C1491 vdd.n525 gnd 0.010592f
C1492 vdd.n526 gnd 0.008525f
C1493 vdd.n527 gnd 0.008525f
C1494 vdd.n528 gnd 0.010592f
C1495 vdd.n529 gnd 0.010592f
C1496 vdd.n530 gnd 0.008525f
C1497 vdd.n531 gnd 0.010592f
C1498 vdd.n532 gnd 0.010592f
C1499 vdd.n533 gnd 0.010592f
C1500 vdd.n534 gnd 0.010592f
C1501 vdd.n535 gnd 0.010592f
C1502 vdd.n536 gnd 0.008525f
C1503 vdd.n537 gnd 0.008525f
C1504 vdd.n538 gnd 0.010592f
C1505 vdd.n539 gnd 0.010592f
C1506 vdd.n540 gnd 0.008525f
C1507 vdd.n541 gnd 0.010592f
C1508 vdd.n542 gnd 0.010592f
C1509 vdd.n543 gnd 0.010592f
C1510 vdd.n544 gnd 0.010592f
C1511 vdd.n545 gnd 0.010592f
C1512 vdd.n546 gnd 0.005797f
C1513 vdd.n547 gnd 0.018244f
C1514 vdd.n548 gnd 0.010592f
C1515 vdd.n549 gnd 0.010592f
C1516 vdd.n550 gnd 0.00844f
C1517 vdd.n551 gnd 0.010592f
C1518 vdd.n552 gnd 0.010592f
C1519 vdd.n553 gnd 0.010592f
C1520 vdd.n554 gnd 0.010592f
C1521 vdd.n555 gnd 0.010592f
C1522 vdd.n556 gnd 0.008525f
C1523 vdd.n557 gnd 0.008525f
C1524 vdd.n558 gnd 0.010592f
C1525 vdd.n559 gnd 0.010592f
C1526 vdd.n560 gnd 0.008525f
C1527 vdd.n561 gnd 0.010592f
C1528 vdd.n562 gnd 0.010592f
C1529 vdd.n563 gnd 0.010592f
C1530 vdd.n564 gnd 0.010592f
C1531 vdd.n565 gnd 0.010592f
C1532 vdd.n566 gnd 0.008525f
C1533 vdd.n567 gnd 0.008525f
C1534 vdd.n568 gnd 0.010592f
C1535 vdd.n569 gnd 0.010592f
C1536 vdd.n570 gnd 0.008525f
C1537 vdd.n571 gnd 0.010592f
C1538 vdd.n572 gnd 0.010592f
C1539 vdd.n573 gnd 0.010592f
C1540 vdd.n574 gnd 0.010592f
C1541 vdd.n575 gnd 0.010592f
C1542 vdd.n576 gnd 0.008525f
C1543 vdd.n577 gnd 0.008525f
C1544 vdd.n578 gnd 0.010592f
C1545 vdd.n579 gnd 0.010592f
C1546 vdd.n580 gnd 0.008525f
C1547 vdd.n581 gnd 0.010592f
C1548 vdd.n582 gnd 0.010592f
C1549 vdd.n583 gnd 0.010592f
C1550 vdd.n584 gnd 0.010592f
C1551 vdd.n585 gnd 0.010592f
C1552 vdd.n586 gnd 0.008525f
C1553 vdd.n587 gnd 0.008525f
C1554 vdd.n588 gnd 0.010592f
C1555 vdd.n589 gnd 0.010592f
C1556 vdd.n590 gnd 0.008525f
C1557 vdd.n591 gnd 0.010592f
C1558 vdd.n592 gnd 0.010592f
C1559 vdd.n593 gnd 0.010592f
C1560 vdd.n594 gnd 0.010592f
C1561 vdd.n595 gnd 0.010592f
C1562 vdd.n596 gnd 0.008525f
C1563 vdd.n597 gnd 0.010592f
C1564 vdd.n598 gnd 0.008525f
C1565 vdd.n599 gnd 0.004476f
C1566 vdd.n600 gnd 0.010592f
C1567 vdd.n601 gnd 0.010592f
C1568 vdd.n602 gnd 0.008525f
C1569 vdd.n603 gnd 0.010592f
C1570 vdd.n604 gnd 0.008525f
C1571 vdd.n605 gnd 0.010592f
C1572 vdd.n606 gnd 0.008525f
C1573 vdd.n607 gnd 0.010592f
C1574 vdd.n608 gnd 0.008525f
C1575 vdd.n609 gnd 0.010592f
C1576 vdd.n610 gnd 0.008525f
C1577 vdd.n611 gnd 0.010592f
C1578 vdd.n612 gnd 0.010592f
C1579 vdd.n613 gnd 0.589935f
C1580 vdd.t155 gnd 0.541225f
C1581 vdd.n614 gnd 0.010592f
C1582 vdd.n615 gnd 0.008525f
C1583 vdd.n616 gnd 0.010592f
C1584 vdd.n617 gnd 0.008525f
C1585 vdd.n618 gnd 0.010592f
C1586 vdd.t200 gnd 0.541225f
C1587 vdd.n619 gnd 0.010592f
C1588 vdd.n620 gnd 0.008525f
C1589 vdd.n621 gnd 0.010592f
C1590 vdd.n622 gnd 0.008525f
C1591 vdd.n623 gnd 0.010592f
C1592 vdd.t145 gnd 0.541225f
C1593 vdd.n624 gnd 0.676531f
C1594 vdd.n625 gnd 0.010592f
C1595 vdd.n626 gnd 0.008525f
C1596 vdd.n627 gnd 0.010592f
C1597 vdd.n628 gnd 0.008525f
C1598 vdd.n629 gnd 0.010592f
C1599 vdd.t118 gnd 0.541225f
C1600 vdd.n630 gnd 0.010592f
C1601 vdd.n631 gnd 0.008525f
C1602 vdd.n632 gnd 0.010592f
C1603 vdd.n633 gnd 0.008525f
C1604 vdd.n634 gnd 0.010592f
C1605 vdd.n635 gnd 0.752302f
C1606 vdd.n636 gnd 0.898433f
C1607 vdd.t173 gnd 0.541225f
C1608 vdd.n637 gnd 0.010592f
C1609 vdd.n638 gnd 0.008525f
C1610 vdd.n639 gnd 0.010592f
C1611 vdd.n640 gnd 0.008525f
C1612 vdd.n641 gnd 0.010592f
C1613 vdd.n642 gnd 0.568286f
C1614 vdd.n643 gnd 0.010592f
C1615 vdd.n644 gnd 0.008525f
C1616 vdd.n645 gnd 0.010592f
C1617 vdd.n646 gnd 0.008525f
C1618 vdd.n647 gnd 0.010592f
C1619 vdd.n648 gnd 1.08245f
C1620 vdd.t112 gnd 0.541225f
C1621 vdd.n649 gnd 0.010592f
C1622 vdd.n650 gnd 0.008525f
C1623 vdd.n651 gnd 0.010592f
C1624 vdd.n652 gnd 0.008525f
C1625 vdd.n653 gnd 0.010592f
C1626 vdd.t5 gnd 0.541225f
C1627 vdd.n654 gnd 0.010592f
C1628 vdd.n655 gnd 0.008525f
C1629 vdd.n656 gnd 0.024285f
C1630 vdd.n657 gnd 0.024285f
C1631 vdd.n658 gnd 7.65292f
C1632 vdd.n659 gnd 0.600759f
C1633 vdd.n660 gnd 0.024285f
C1634 vdd.n661 gnd 0.009109f
C1635 vdd.n662 gnd 0.008525f
C1636 vdd.n667 gnd 0.006779f
C1637 vdd.n668 gnd 0.008525f
C1638 vdd.n669 gnd 0.010592f
C1639 vdd.n670 gnd 0.010592f
C1640 vdd.n671 gnd 0.010592f
C1641 vdd.n672 gnd 0.010592f
C1642 vdd.n673 gnd 0.010592f
C1643 vdd.n674 gnd 0.008525f
C1644 vdd.n675 gnd 0.010592f
C1645 vdd.n676 gnd 0.010592f
C1646 vdd.n677 gnd 0.010592f
C1647 vdd.n678 gnd 0.010592f
C1648 vdd.n679 gnd 0.010592f
C1649 vdd.n680 gnd 0.008525f
C1650 vdd.n681 gnd 0.010592f
C1651 vdd.n682 gnd 0.010592f
C1652 vdd.n683 gnd 0.010592f
C1653 vdd.n684 gnd 0.010592f
C1654 vdd.n685 gnd 0.010592f
C1655 vdd.t17 gnd 0.130309f
C1656 vdd.t18 gnd 0.139265f
C1657 vdd.t16 gnd 0.170182f
C1658 vdd.n686 gnd 0.218149f
C1659 vdd.n687 gnd 0.183285f
C1660 vdd.n688 gnd 0.017392f
C1661 vdd.n689 gnd 0.010592f
C1662 vdd.n690 gnd 0.010592f
C1663 vdd.n691 gnd 0.010592f
C1664 vdd.n692 gnd 0.010592f
C1665 vdd.n693 gnd 0.010592f
C1666 vdd.n694 gnd 0.008525f
C1667 vdd.n695 gnd 0.010592f
C1668 vdd.n696 gnd 0.010592f
C1669 vdd.n697 gnd 0.010592f
C1670 vdd.n698 gnd 0.010592f
C1671 vdd.n699 gnd 0.010592f
C1672 vdd.n700 gnd 0.008525f
C1673 vdd.n701 gnd 0.010592f
C1674 vdd.n702 gnd 0.010592f
C1675 vdd.n703 gnd 0.010592f
C1676 vdd.n704 gnd 0.010592f
C1677 vdd.n705 gnd 0.010592f
C1678 vdd.n706 gnd 0.008525f
C1679 vdd.n707 gnd 0.010592f
C1680 vdd.n708 gnd 0.010592f
C1681 vdd.n709 gnd 0.010592f
C1682 vdd.n710 gnd 0.010592f
C1683 vdd.n711 gnd 0.010592f
C1684 vdd.n712 gnd 0.008525f
C1685 vdd.n713 gnd 0.010592f
C1686 vdd.n714 gnd 0.010592f
C1687 vdd.n715 gnd 0.010592f
C1688 vdd.n716 gnd 0.010592f
C1689 vdd.n717 gnd 0.010592f
C1690 vdd.n718 gnd 0.008525f
C1691 vdd.n719 gnd 0.010592f
C1692 vdd.n720 gnd 0.010592f
C1693 vdd.n721 gnd 0.010592f
C1694 vdd.n722 gnd 0.00844f
C1695 vdd.t6 gnd 0.130309f
C1696 vdd.t7 gnd 0.139265f
C1697 vdd.t4 gnd 0.170182f
C1698 vdd.n723 gnd 0.218149f
C1699 vdd.n724 gnd 0.183285f
C1700 vdd.n725 gnd 0.010592f
C1701 vdd.n726 gnd 0.008525f
C1702 vdd.n728 gnd 0.010592f
C1703 vdd.n730 gnd 0.010592f
C1704 vdd.n731 gnd 0.010592f
C1705 vdd.n732 gnd 0.008525f
C1706 vdd.n733 gnd 0.010592f
C1707 vdd.n734 gnd 0.010592f
C1708 vdd.n735 gnd 0.010592f
C1709 vdd.n736 gnd 0.010592f
C1710 vdd.n737 gnd 0.010592f
C1711 vdd.n738 gnd 0.008525f
C1712 vdd.n739 gnd 0.010592f
C1713 vdd.n740 gnd 0.010592f
C1714 vdd.n741 gnd 0.010592f
C1715 vdd.n742 gnd 0.010592f
C1716 vdd.n743 gnd 0.010592f
C1717 vdd.n744 gnd 0.008525f
C1718 vdd.n745 gnd 0.010592f
C1719 vdd.n746 gnd 0.010592f
C1720 vdd.n747 gnd 0.010592f
C1721 vdd.n748 gnd 0.006779f
C1722 vdd.n753 gnd 0.007203f
C1723 vdd.n754 gnd 0.007203f
C1724 vdd.n755 gnd 0.007203f
C1725 vdd.n756 gnd 7.45808f
C1726 vdd.n757 gnd 0.007203f
C1727 vdd.n758 gnd 0.007203f
C1728 vdd.n759 gnd 0.007203f
C1729 vdd.n761 gnd 0.007203f
C1730 vdd.n762 gnd 0.007203f
C1731 vdd.n764 gnd 0.007203f
C1732 vdd.n765 gnd 0.005243f
C1733 vdd.n767 gnd 0.007203f
C1734 vdd.t53 gnd 0.291054f
C1735 vdd.t52 gnd 0.29793f
C1736 vdd.t51 gnd 0.190011f
C1737 vdd.n768 gnd 0.102691f
C1738 vdd.n769 gnd 0.058249f
C1739 vdd.n770 gnd 0.010294f
C1740 vdd.n771 gnd 0.016834f
C1741 vdd.n773 gnd 0.007203f
C1742 vdd.n774 gnd 0.736066f
C1743 vdd.n775 gnd 0.015957f
C1744 vdd.n776 gnd 0.015957f
C1745 vdd.n777 gnd 0.007203f
C1746 vdd.n778 gnd 0.01709f
C1747 vdd.n779 gnd 0.007203f
C1748 vdd.n780 gnd 0.007203f
C1749 vdd.n781 gnd 0.007203f
C1750 vdd.n782 gnd 0.007203f
C1751 vdd.n783 gnd 0.007203f
C1752 vdd.n785 gnd 0.007203f
C1753 vdd.n786 gnd 0.007203f
C1754 vdd.n788 gnd 0.007203f
C1755 vdd.n789 gnd 0.007203f
C1756 vdd.n791 gnd 0.007203f
C1757 vdd.n792 gnd 0.007203f
C1758 vdd.n794 gnd 0.007203f
C1759 vdd.n795 gnd 0.007203f
C1760 vdd.n797 gnd 0.007203f
C1761 vdd.n798 gnd 0.007203f
C1762 vdd.n800 gnd 0.007203f
C1763 vdd.n801 gnd 0.005243f
C1764 vdd.n803 gnd 0.007203f
C1765 vdd.t46 gnd 0.291054f
C1766 vdd.t45 gnd 0.29793f
C1767 vdd.t43 gnd 0.190011f
C1768 vdd.n804 gnd 0.102691f
C1769 vdd.n805 gnd 0.058249f
C1770 vdd.n806 gnd 0.010294f
C1771 vdd.n807 gnd 0.007203f
C1772 vdd.n808 gnd 0.007203f
C1773 vdd.t44 gnd 0.368033f
C1774 vdd.n809 gnd 0.007203f
C1775 vdd.n810 gnd 0.007203f
C1776 vdd.n811 gnd 0.007203f
C1777 vdd.n812 gnd 0.007203f
C1778 vdd.n813 gnd 0.007203f
C1779 vdd.n814 gnd 0.736066f
C1780 vdd.n815 gnd 0.007203f
C1781 vdd.n816 gnd 0.007203f
C1782 vdd.n817 gnd 0.644057f
C1783 vdd.n818 gnd 0.007203f
C1784 vdd.n819 gnd 0.007203f
C1785 vdd.n820 gnd 0.006355f
C1786 vdd.n821 gnd 0.007203f
C1787 vdd.n822 gnd 0.64947f
C1788 vdd.n823 gnd 0.007203f
C1789 vdd.n824 gnd 0.007203f
C1790 vdd.n825 gnd 0.007203f
C1791 vdd.n826 gnd 0.007203f
C1792 vdd.n827 gnd 0.007203f
C1793 vdd.n828 gnd 0.736066f
C1794 vdd.n829 gnd 0.007203f
C1795 vdd.n830 gnd 0.007203f
C1796 vdd.t27 gnd 0.330147f
C1797 vdd.t96 gnd 0.086596f
C1798 vdd.n831 gnd 0.007203f
C1799 vdd.n832 gnd 0.007203f
C1800 vdd.n833 gnd 0.007203f
C1801 vdd.t92 gnd 0.368033f
C1802 vdd.n834 gnd 0.007203f
C1803 vdd.n835 gnd 0.007203f
C1804 vdd.n836 gnd 0.007203f
C1805 vdd.n837 gnd 0.007203f
C1806 vdd.n838 gnd 0.007203f
C1807 vdd.t93 gnd 0.368033f
C1808 vdd.n839 gnd 0.007203f
C1809 vdd.n840 gnd 0.007203f
C1810 vdd.n841 gnd 0.611584f
C1811 vdd.n842 gnd 0.007203f
C1812 vdd.n843 gnd 0.007203f
C1813 vdd.n844 gnd 0.007203f
C1814 vdd.n845 gnd 0.449217f
C1815 vdd.n846 gnd 0.007203f
C1816 vdd.n847 gnd 0.007203f
C1817 vdd.t246 gnd 0.368033f
C1818 vdd.n848 gnd 0.007203f
C1819 vdd.n849 gnd 0.007203f
C1820 vdd.n850 gnd 0.007203f
C1821 vdd.n851 gnd 0.611584f
C1822 vdd.n852 gnd 0.007203f
C1823 vdd.n853 gnd 0.007203f
C1824 vdd.t97 gnd 0.31391f
C1825 vdd.t94 gnd 0.286849f
C1826 vdd.n854 gnd 0.007203f
C1827 vdd.n855 gnd 0.007203f
C1828 vdd.n856 gnd 0.007203f
C1829 vdd.t260 gnd 0.368033f
C1830 vdd.n857 gnd 0.007203f
C1831 vdd.n858 gnd 0.007203f
C1832 vdd.t109 gnd 0.368033f
C1833 vdd.n859 gnd 0.007203f
C1834 vdd.n860 gnd 0.007203f
C1835 vdd.n861 gnd 0.007203f
C1836 vdd.t104 gnd 0.270612f
C1837 vdd.n862 gnd 0.007203f
C1838 vdd.n863 gnd 0.007203f
C1839 vdd.n864 gnd 0.627821f
C1840 vdd.n865 gnd 0.007203f
C1841 vdd.n866 gnd 0.007203f
C1842 vdd.n867 gnd 0.007203f
C1843 vdd.n868 gnd 0.736066f
C1844 vdd.n869 gnd 0.007203f
C1845 vdd.n870 gnd 0.007203f
C1846 vdd.t240 gnd 0.330147f
C1847 vdd.n871 gnd 0.465453f
C1848 vdd.n872 gnd 0.007203f
C1849 vdd.n873 gnd 0.007203f
C1850 vdd.n874 gnd 0.007203f
C1851 vdd.t102 gnd 0.368033f
C1852 vdd.n875 gnd 0.007203f
C1853 vdd.n876 gnd 0.007203f
C1854 vdd.n877 gnd 0.007203f
C1855 vdd.n878 gnd 0.007203f
C1856 vdd.n879 gnd 0.007203f
C1857 vdd.t248 gnd 0.736066f
C1858 vdd.n880 gnd 0.007203f
C1859 vdd.n881 gnd 0.007203f
C1860 vdd.t48 gnd 0.368033f
C1861 vdd.n882 gnd 0.007203f
C1862 vdd.n883 gnd 0.01709f
C1863 vdd.n884 gnd 0.01709f
C1864 vdd.t250 gnd 0.692768f
C1865 vdd.n885 gnd 0.015957f
C1866 vdd.n886 gnd 0.015957f
C1867 vdd.n887 gnd 0.01709f
C1868 vdd.n888 gnd 0.007203f
C1869 vdd.n889 gnd 0.007203f
C1870 vdd.t258 gnd 0.692768f
C1871 vdd.n907 gnd 0.01709f
C1872 vdd.n925 gnd 0.015957f
C1873 vdd.n926 gnd 0.007203f
C1874 vdd.n927 gnd 0.015957f
C1875 vdd.t66 gnd 0.291054f
C1876 vdd.t65 gnd 0.29793f
C1877 vdd.t64 gnd 0.190011f
C1878 vdd.n928 gnd 0.102691f
C1879 vdd.n929 gnd 0.058249f
C1880 vdd.n930 gnd 0.016834f
C1881 vdd.n931 gnd 0.007203f
C1882 vdd.t262 gnd 0.736066f
C1883 vdd.n932 gnd 0.015957f
C1884 vdd.n933 gnd 0.007203f
C1885 vdd.n934 gnd 0.01709f
C1886 vdd.n935 gnd 0.007203f
C1887 vdd.t42 gnd 0.291054f
C1888 vdd.t41 gnd 0.29793f
C1889 vdd.t39 gnd 0.190011f
C1890 vdd.n936 gnd 0.102691f
C1891 vdd.n937 gnd 0.058249f
C1892 vdd.n938 gnd 0.010294f
C1893 vdd.n939 gnd 0.007203f
C1894 vdd.n940 gnd 0.007203f
C1895 vdd.t40 gnd 0.368033f
C1896 vdd.n941 gnd 0.007203f
C1897 vdd.n942 gnd 0.007203f
C1898 vdd.n943 gnd 0.007203f
C1899 vdd.n944 gnd 0.007203f
C1900 vdd.n945 gnd 0.007203f
C1901 vdd.n946 gnd 0.007203f
C1902 vdd.n947 gnd 0.736066f
C1903 vdd.n948 gnd 0.007203f
C1904 vdd.n949 gnd 0.007203f
C1905 vdd.t244 gnd 0.368033f
C1906 vdd.n950 gnd 0.007203f
C1907 vdd.n951 gnd 0.007203f
C1908 vdd.n952 gnd 0.007203f
C1909 vdd.n953 gnd 0.007203f
C1910 vdd.n954 gnd 0.465453f
C1911 vdd.n955 gnd 0.007203f
C1912 vdd.n956 gnd 0.007203f
C1913 vdd.n957 gnd 0.007203f
C1914 vdd.n958 gnd 0.007203f
C1915 vdd.n959 gnd 0.007203f
C1916 vdd.n960 gnd 0.627821f
C1917 vdd.n961 gnd 0.007203f
C1918 vdd.n962 gnd 0.007203f
C1919 vdd.t254 gnd 0.330147f
C1920 vdd.t98 gnd 0.270612f
C1921 vdd.n963 gnd 0.007203f
C1922 vdd.n964 gnd 0.007203f
C1923 vdd.n965 gnd 0.007203f
C1924 vdd.t108 gnd 0.368033f
C1925 vdd.n966 gnd 0.007203f
C1926 vdd.n967 gnd 0.007203f
C1927 vdd.t100 gnd 0.368033f
C1928 vdd.n968 gnd 0.007203f
C1929 vdd.n969 gnd 0.007203f
C1930 vdd.n970 gnd 0.007203f
C1931 vdd.t242 gnd 0.286849f
C1932 vdd.n971 gnd 0.007203f
C1933 vdd.n972 gnd 0.007203f
C1934 vdd.n973 gnd 0.611584f
C1935 vdd.n974 gnd 0.007203f
C1936 vdd.n975 gnd 0.007203f
C1937 vdd.n976 gnd 0.007203f
C1938 vdd.t256 gnd 0.368033f
C1939 vdd.n977 gnd 0.007203f
C1940 vdd.n978 gnd 0.007203f
C1941 vdd.t107 gnd 0.31391f
C1942 vdd.n979 gnd 0.449217f
C1943 vdd.n980 gnd 0.007203f
C1944 vdd.n981 gnd 0.007203f
C1945 vdd.n982 gnd 0.007203f
C1946 vdd.n983 gnd 0.611584f
C1947 vdd.n984 gnd 0.007203f
C1948 vdd.n985 gnd 0.007203f
C1949 vdd.t99 gnd 0.368033f
C1950 vdd.n986 gnd 0.007203f
C1951 vdd.n987 gnd 0.007203f
C1952 vdd.n988 gnd 0.007203f
C1953 vdd.n989 gnd 0.736066f
C1954 vdd.n990 gnd 0.007203f
C1955 vdd.n991 gnd 0.007203f
C1956 vdd.t106 gnd 0.368033f
C1957 vdd.n992 gnd 0.007203f
C1958 vdd.n993 gnd 0.007203f
C1959 vdd.n994 gnd 0.007203f
C1960 vdd.t105 gnd 0.086596f
C1961 vdd.n995 gnd 0.007203f
C1962 vdd.n996 gnd 0.007203f
C1963 vdd.n997 gnd 0.007203f
C1964 vdd.t59 gnd 0.29793f
C1965 vdd.t57 gnd 0.190011f
C1966 vdd.t60 gnd 0.29793f
C1967 vdd.n998 gnd 0.167449f
C1968 vdd.n999 gnd 0.007203f
C1969 vdd.n1000 gnd 0.007203f
C1970 vdd.n1001 gnd 0.736066f
C1971 vdd.n1002 gnd 0.007203f
C1972 vdd.n1003 gnd 0.007203f
C1973 vdd.t58 gnd 0.330147f
C1974 vdd.n1004 gnd 0.64947f
C1975 vdd.n1005 gnd 0.007203f
C1976 vdd.n1006 gnd 0.007203f
C1977 vdd.n1007 gnd 0.007203f
C1978 vdd.n1008 gnd 0.644057f
C1979 vdd.n1009 gnd 0.007203f
C1980 vdd.n1010 gnd 0.007203f
C1981 vdd.n1011 gnd 0.007203f
C1982 vdd.n1012 gnd 0.007203f
C1983 vdd.n1013 gnd 0.007203f
C1984 vdd.n1014 gnd 0.736066f
C1985 vdd.n1015 gnd 0.007203f
C1986 vdd.n1016 gnd 0.007203f
C1987 vdd.t1 gnd 0.368033f
C1988 vdd.n1017 gnd 0.007203f
C1989 vdd.n1018 gnd 0.01709f
C1990 vdd.n1019 gnd 0.01709f
C1991 vdd.n1020 gnd 7.45808f
C1992 vdd.n1021 gnd 0.015957f
C1993 vdd.n1022 gnd 0.015957f
C1994 vdd.n1023 gnd 0.01709f
C1995 vdd.n1024 gnd 0.007203f
C1996 vdd.n1025 gnd 0.007203f
C1997 vdd.n1026 gnd 0.007203f
C1998 vdd.n1027 gnd 0.007203f
C1999 vdd.n1028 gnd 0.007203f
C2000 vdd.n1029 gnd 0.007203f
C2001 vdd.n1030 gnd 0.007203f
C2002 vdd.n1031 gnd 0.007203f
C2003 vdd.n1033 gnd 0.007203f
C2004 vdd.n1034 gnd 0.007203f
C2005 vdd.n1035 gnd 0.006779f
C2006 vdd.n1038 gnd 0.024285f
C2007 vdd.n1039 gnd 0.008525f
C2008 vdd.n1040 gnd 0.010592f
C2009 vdd.n1042 gnd 0.010592f
C2010 vdd.n1043 gnd 0.007076f
C2011 vdd.n1044 gnd 0.600759f
C2012 vdd.n1045 gnd 7.65292f
C2013 vdd.n1046 gnd 0.010592f
C2014 vdd.n1047 gnd 0.024285f
C2015 vdd.n1048 gnd 0.008525f
C2016 vdd.n1049 gnd 0.010592f
C2017 vdd.n1050 gnd 0.008525f
C2018 vdd.n1051 gnd 0.010592f
C2019 vdd.n1052 gnd 1.08245f
C2020 vdd.n1053 gnd 0.010592f
C2021 vdd.n1054 gnd 0.008525f
C2022 vdd.n1055 gnd 0.008525f
C2023 vdd.n1056 gnd 0.010592f
C2024 vdd.n1057 gnd 0.008525f
C2025 vdd.n1058 gnd 0.010592f
C2026 vdd.t114 gnd 0.541225f
C2027 vdd.n1059 gnd 0.010592f
C2028 vdd.n1060 gnd 0.008525f
C2029 vdd.n1061 gnd 0.010592f
C2030 vdd.n1062 gnd 0.008525f
C2031 vdd.n1063 gnd 0.010592f
C2032 vdd.t217 gnd 0.541225f
C2033 vdd.n1064 gnd 0.010592f
C2034 vdd.n1065 gnd 0.008525f
C2035 vdd.n1066 gnd 0.010592f
C2036 vdd.n1067 gnd 0.008525f
C2037 vdd.n1068 gnd 0.010592f
C2038 vdd.t126 gnd 0.541225f
C2039 vdd.n1069 gnd 0.752302f
C2040 vdd.n1070 gnd 0.010592f
C2041 vdd.n1071 gnd 0.008525f
C2042 vdd.n1072 gnd 0.010592f
C2043 vdd.n1073 gnd 0.008525f
C2044 vdd.n1074 gnd 0.010592f
C2045 vdd.n1075 gnd 0.860547f
C2046 vdd.n1076 gnd 0.010592f
C2047 vdd.n1077 gnd 0.008525f
C2048 vdd.n1078 gnd 0.010592f
C2049 vdd.n1079 gnd 0.008525f
C2050 vdd.n1080 gnd 0.010592f
C2051 vdd.n1081 gnd 0.676531f
C2052 vdd.t147 gnd 0.541225f
C2053 vdd.n1082 gnd 0.010592f
C2054 vdd.n1083 gnd 0.008525f
C2055 vdd.n1084 gnd 0.010592f
C2056 vdd.n1085 gnd 0.008525f
C2057 vdd.n1086 gnd 0.010592f
C2058 vdd.t167 gnd 0.541225f
C2059 vdd.n1087 gnd 0.010592f
C2060 vdd.n1088 gnd 0.008525f
C2061 vdd.n1089 gnd 0.010592f
C2062 vdd.n1090 gnd 0.008525f
C2063 vdd.n1091 gnd 0.010592f
C2064 vdd.t196 gnd 0.541225f
C2065 vdd.n1092 gnd 0.589935f
C2066 vdd.n1093 gnd 0.010592f
C2067 vdd.n1094 gnd 0.008525f
C2068 vdd.n1095 gnd 0.010592f
C2069 vdd.n1096 gnd 0.008525f
C2070 vdd.n1097 gnd 0.010592f
C2071 vdd.t187 gnd 0.541225f
C2072 vdd.n1098 gnd 0.010592f
C2073 vdd.n1099 gnd 0.008525f
C2074 vdd.n1100 gnd 0.010592f
C2075 vdd.n1101 gnd 0.008525f
C2076 vdd.n1102 gnd 0.010592f
C2077 vdd.n1103 gnd 0.838898f
C2078 vdd.n1104 gnd 0.898433f
C2079 vdd.t124 gnd 0.541225f
C2080 vdd.n1105 gnd 0.010592f
C2081 vdd.n1106 gnd 0.008525f
C2082 vdd.n1107 gnd 0.010592f
C2083 vdd.n1108 gnd 0.008525f
C2084 vdd.n1109 gnd 0.010592f
C2085 vdd.n1110 gnd 0.654882f
C2086 vdd.n1111 gnd 0.010592f
C2087 vdd.n1112 gnd 0.008525f
C2088 vdd.n1113 gnd 0.010592f
C2089 vdd.n1114 gnd 0.008525f
C2090 vdd.n1115 gnd 0.010592f
C2091 vdd.t142 gnd 0.541225f
C2092 vdd.t132 gnd 0.541225f
C2093 vdd.n1116 gnd 0.010592f
C2094 vdd.n1117 gnd 0.008525f
C2095 vdd.n1118 gnd 0.010592f
C2096 vdd.n1119 gnd 0.008525f
C2097 vdd.n1120 gnd 0.010592f
C2098 vdd.t182 gnd 0.541225f
C2099 vdd.n1121 gnd 0.010592f
C2100 vdd.n1122 gnd 0.008525f
C2101 vdd.n1123 gnd 0.010592f
C2102 vdd.n1124 gnd 0.008525f
C2103 vdd.n1125 gnd 0.010592f
C2104 vdd.t184 gnd 0.541225f
C2105 vdd.n1126 gnd 0.7956f
C2106 vdd.n1127 gnd 0.010592f
C2107 vdd.n1128 gnd 0.008525f
C2108 vdd.n1129 gnd 0.010592f
C2109 vdd.n1130 gnd 0.008525f
C2110 vdd.n1131 gnd 0.010592f
C2111 vdd.n1132 gnd 1.08245f
C2112 vdd.n1133 gnd 0.010592f
C2113 vdd.n1134 gnd 0.008525f
C2114 vdd.n1135 gnd 0.010592f
C2115 vdd.n1136 gnd 0.008525f
C2116 vdd.n1137 gnd 0.010592f
C2117 vdd.n1138 gnd 0.91467f
C2118 vdd.n1139 gnd 0.010592f
C2119 vdd.n1140 gnd 0.008525f
C2120 vdd.n1141 gnd 0.02412f
C2121 vdd.n1142 gnd 0.007076f
C2122 vdd.n1143 gnd 0.02412f
C2123 vdd.n1144 gnd 1.42883f
C2124 vdd.n1145 gnd 0.02412f
C2125 vdd.n1146 gnd 0.007076f
C2126 vdd.n1147 gnd 0.010592f
C2127 vdd.t14 gnd 0.130309f
C2128 vdd.t15 gnd 0.139265f
C2129 vdd.t12 gnd 0.170182f
C2130 vdd.n1148 gnd 0.218149f
C2131 vdd.n1149 gnd 0.184137f
C2132 vdd.n1150 gnd 0.013981f
C2133 vdd.n1151 gnd 0.010592f
C2134 vdd.n1182 gnd 0.010592f
C2135 vdd.n1183 gnd 0.010592f
C2136 vdd.n1184 gnd 0.024285f
C2137 vdd.n1185 gnd 0.008525f
C2138 vdd.n1186 gnd 0.010592f
C2139 vdd.n1187 gnd 0.010592f
C2140 vdd.n1188 gnd 0.010592f
C2141 vdd.n1189 gnd 0.010592f
C2142 vdd.n1190 gnd 0.008525f
C2143 vdd.n1191 gnd 0.010592f
C2144 vdd.n1192 gnd 0.010592f
C2145 vdd.n1193 gnd 0.010592f
C2146 vdd.n1194 gnd 0.010592f
C2147 vdd.n1195 gnd 0.010592f
C2148 vdd.n1196 gnd 0.008525f
C2149 vdd.n1197 gnd 0.010592f
C2150 vdd.n1198 gnd 0.010592f
C2151 vdd.n1199 gnd 0.010592f
C2152 vdd.n1200 gnd 0.010592f
C2153 vdd.n1201 gnd 0.010592f
C2154 vdd.n1202 gnd 0.008525f
C2155 vdd.n1203 gnd 0.010592f
C2156 vdd.n1204 gnd 0.010592f
C2157 vdd.n1205 gnd 0.010592f
C2158 vdd.n1206 gnd 0.010592f
C2159 vdd.n1207 gnd 0.010592f
C2160 vdd.n1208 gnd 0.007119f
C2161 vdd.n1209 gnd 0.010592f
C2162 vdd.n1210 gnd 0.010592f
C2163 vdd.n1211 gnd 0.010592f
C2164 vdd.n1212 gnd 0.008525f
C2165 vdd.n1213 gnd 0.010592f
C2166 vdd.n1214 gnd 0.010592f
C2167 vdd.n1215 gnd 0.010592f
C2168 vdd.n1216 gnd 0.010592f
C2169 vdd.n1217 gnd 0.010592f
C2170 vdd.n1218 gnd 0.008525f
C2171 vdd.n1219 gnd 0.010592f
C2172 vdd.n1220 gnd 0.010592f
C2173 vdd.n1221 gnd 0.010592f
C2174 vdd.n1222 gnd 0.010592f
C2175 vdd.n1223 gnd 0.010592f
C2176 vdd.n1224 gnd 0.008525f
C2177 vdd.n1225 gnd 0.010592f
C2178 vdd.n1226 gnd 0.010592f
C2179 vdd.n1227 gnd 0.010592f
C2180 vdd.n1228 gnd 0.010592f
C2181 vdd.n1229 gnd 0.010592f
C2182 vdd.n1230 gnd 0.008525f
C2183 vdd.n1231 gnd 0.010592f
C2184 vdd.n1232 gnd 0.010592f
C2185 vdd.n1233 gnd 0.010592f
C2186 vdd.n1234 gnd 0.010592f
C2187 vdd.n1235 gnd 0.010592f
C2188 vdd.n1236 gnd 0.008525f
C2189 vdd.n1237 gnd 0.010592f
C2190 vdd.n1238 gnd 0.010592f
C2191 vdd.n1239 gnd 0.010592f
C2192 vdd.n1240 gnd 0.010592f
C2193 vdd.n1241 gnd 0.00844f
C2194 vdd.n1242 gnd 0.010592f
C2195 vdd.n1243 gnd 0.010592f
C2196 vdd.n1244 gnd 0.010592f
C2197 vdd.n1245 gnd 0.010592f
C2198 vdd.n1246 gnd 0.010592f
C2199 vdd.n1247 gnd 0.008525f
C2200 vdd.n1248 gnd 0.010592f
C2201 vdd.n1249 gnd 0.010592f
C2202 vdd.n1250 gnd 0.010592f
C2203 vdd.n1251 gnd 0.010592f
C2204 vdd.n1252 gnd 0.010592f
C2205 vdd.n1253 gnd 0.008525f
C2206 vdd.n1254 gnd 0.010592f
C2207 vdd.n1255 gnd 0.010592f
C2208 vdd.n1256 gnd 0.010592f
C2209 vdd.n1257 gnd 0.010592f
C2210 vdd.n1258 gnd 0.010592f
C2211 vdd.n1259 gnd 0.008525f
C2212 vdd.n1260 gnd 0.010592f
C2213 vdd.n1261 gnd 0.010592f
C2214 vdd.n1262 gnd 0.010592f
C2215 vdd.n1263 gnd 0.010592f
C2216 vdd.n1264 gnd 0.010592f
C2217 vdd.n1265 gnd 0.008525f
C2218 vdd.n1266 gnd 0.010592f
C2219 vdd.n1267 gnd 0.010592f
C2220 vdd.n1268 gnd 0.010592f
C2221 vdd.n1269 gnd 0.010592f
C2222 vdd.n1270 gnd 0.010592f
C2223 vdd.n1271 gnd 0.004476f
C2224 vdd.n1272 gnd 0.010592f
C2225 vdd.n1273 gnd 0.008525f
C2226 vdd.n1274 gnd 0.008525f
C2227 vdd.n1275 gnd 0.008525f
C2228 vdd.n1276 gnd 0.010592f
C2229 vdd.n1277 gnd 0.010592f
C2230 vdd.n1278 gnd 0.010592f
C2231 vdd.n1279 gnd 0.008525f
C2232 vdd.n1280 gnd 0.008525f
C2233 vdd.n1281 gnd 0.008525f
C2234 vdd.n1282 gnd 0.010592f
C2235 vdd.n1283 gnd 0.010592f
C2236 vdd.n1284 gnd 0.010592f
C2237 vdd.n1285 gnd 0.008525f
C2238 vdd.n1286 gnd 0.008525f
C2239 vdd.n1287 gnd 0.008525f
C2240 vdd.n1288 gnd 0.010592f
C2241 vdd.n1289 gnd 0.010592f
C2242 vdd.n1290 gnd 0.010592f
C2243 vdd.n1291 gnd 0.008525f
C2244 vdd.n1292 gnd 0.008525f
C2245 vdd.n1293 gnd 0.008525f
C2246 vdd.n1294 gnd 0.010592f
C2247 vdd.n1295 gnd 0.010592f
C2248 vdd.n1296 gnd 0.010592f
C2249 vdd.n1297 gnd 0.008525f
C2250 vdd.n1298 gnd 0.008525f
C2251 vdd.n1299 gnd 0.008525f
C2252 vdd.n1300 gnd 0.010592f
C2253 vdd.n1301 gnd 0.010592f
C2254 vdd.n1302 gnd 0.010592f
C2255 vdd.n1303 gnd 0.010592f
C2256 vdd.t24 gnd 0.130309f
C2257 vdd.t25 gnd 0.139265f
C2258 vdd.t23 gnd 0.170182f
C2259 vdd.n1304 gnd 0.218149f
C2260 vdd.n1305 gnd 0.184137f
C2261 vdd.n1306 gnd 0.018244f
C2262 vdd.n1307 gnd 0.005797f
C2263 vdd.n1308 gnd 0.008525f
C2264 vdd.n1309 gnd 0.010592f
C2265 vdd.n1310 gnd 0.010592f
C2266 vdd.n1311 gnd 0.010592f
C2267 vdd.n1312 gnd 0.008525f
C2268 vdd.n1313 gnd 0.008525f
C2269 vdd.n1314 gnd 0.008525f
C2270 vdd.n1315 gnd 0.010592f
C2271 vdd.n1316 gnd 0.010592f
C2272 vdd.n1317 gnd 0.010592f
C2273 vdd.n1318 gnd 0.008525f
C2274 vdd.n1319 gnd 0.008525f
C2275 vdd.n1320 gnd 0.008525f
C2276 vdd.n1321 gnd 0.010592f
C2277 vdd.n1322 gnd 0.010592f
C2278 vdd.n1323 gnd 0.010592f
C2279 vdd.n1324 gnd 0.008525f
C2280 vdd.n1325 gnd 0.008525f
C2281 vdd.n1326 gnd 0.008525f
C2282 vdd.n1327 gnd 0.010592f
C2283 vdd.n1328 gnd 0.010592f
C2284 vdd.n1329 gnd 0.010592f
C2285 vdd.n1330 gnd 0.008525f
C2286 vdd.n1331 gnd 0.008525f
C2287 vdd.n1332 gnd 0.008525f
C2288 vdd.n1333 gnd 0.010592f
C2289 vdd.n1334 gnd 0.010592f
C2290 vdd.n1335 gnd 0.010592f
C2291 vdd.n1336 gnd 0.008525f
C2292 vdd.n1337 gnd 0.007119f
C2293 vdd.n1338 gnd 0.010592f
C2294 vdd.n1339 gnd 0.010592f
C2295 vdd.t31 gnd 0.130309f
C2296 vdd.t32 gnd 0.139265f
C2297 vdd.t30 gnd 0.170182f
C2298 vdd.n1340 gnd 0.218149f
C2299 vdd.n1341 gnd 0.184137f
C2300 vdd.n1342 gnd 0.018244f
C2301 vdd.n1343 gnd 0.010592f
C2302 vdd.n1344 gnd 0.010592f
C2303 vdd.n1345 gnd 0.010592f
C2304 vdd.n1346 gnd 0.008525f
C2305 vdd.n1347 gnd 0.008525f
C2306 vdd.n1348 gnd 0.008525f
C2307 vdd.n1349 gnd 0.010592f
C2308 vdd.n1350 gnd 0.010592f
C2309 vdd.n1351 gnd 0.010592f
C2310 vdd.n1352 gnd 0.008525f
C2311 vdd.n1353 gnd 0.008525f
C2312 vdd.n1354 gnd 0.008525f
C2313 vdd.n1355 gnd 0.010592f
C2314 vdd.n1356 gnd 0.010592f
C2315 vdd.n1357 gnd 0.010592f
C2316 vdd.n1358 gnd 0.008525f
C2317 vdd.n1359 gnd 0.008525f
C2318 vdd.n1360 gnd 0.008525f
C2319 vdd.n1361 gnd 0.010592f
C2320 vdd.n1362 gnd 0.010592f
C2321 vdd.n1363 gnd 0.010592f
C2322 vdd.n1364 gnd 0.008525f
C2323 vdd.n1365 gnd 0.008525f
C2324 vdd.n1366 gnd 0.008525f
C2325 vdd.n1367 gnd 0.010592f
C2326 vdd.n1368 gnd 0.010592f
C2327 vdd.n1369 gnd 0.010592f
C2328 vdd.n1370 gnd 0.008525f
C2329 vdd.n1371 gnd 0.007076f
C2330 vdd.n1372 gnd 0.024285f
C2331 vdd.n1374 gnd 2.39221f
C2332 vdd.n1375 gnd 0.024285f
C2333 vdd.n1376 gnd 0.004049f
C2334 vdd.n1377 gnd 0.024285f
C2335 vdd.n1378 gnd 0.02412f
C2336 vdd.n1379 gnd 0.010592f
C2337 vdd.n1380 gnd 0.008525f
C2338 vdd.n1381 gnd 0.010592f
C2339 vdd.t13 gnd 0.541225f
C2340 vdd.n1382 gnd 0.709004f
C2341 vdd.n1383 gnd 0.010592f
C2342 vdd.n1384 gnd 0.008525f
C2343 vdd.n1385 gnd 0.010592f
C2344 vdd.n1386 gnd 0.010592f
C2345 vdd.n1387 gnd 0.010592f
C2346 vdd.n1388 gnd 0.008525f
C2347 vdd.n1389 gnd 0.010592f
C2348 vdd.n1390 gnd 1.08245f
C2349 vdd.n1391 gnd 0.010592f
C2350 vdd.n1392 gnd 0.008525f
C2351 vdd.n1393 gnd 0.010592f
C2352 vdd.n1394 gnd 0.010592f
C2353 vdd.n1395 gnd 0.010592f
C2354 vdd.n1396 gnd 0.008525f
C2355 vdd.n1397 gnd 0.010592f
C2356 vdd.n1398 gnd 0.898433f
C2357 vdd.t122 gnd 0.541225f
C2358 vdd.n1399 gnd 0.622408f
C2359 vdd.n1400 gnd 0.010592f
C2360 vdd.n1401 gnd 0.008525f
C2361 vdd.n1402 gnd 0.010592f
C2362 vdd.n1403 gnd 0.010592f
C2363 vdd.n1404 gnd 0.010592f
C2364 vdd.n1405 gnd 0.008525f
C2365 vdd.n1406 gnd 0.010592f
C2366 vdd.n1407 gnd 0.644057f
C2367 vdd.n1408 gnd 0.010592f
C2368 vdd.n1409 gnd 0.008525f
C2369 vdd.n1410 gnd 0.010592f
C2370 vdd.n1411 gnd 0.010592f
C2371 vdd.n1412 gnd 0.010592f
C2372 vdd.n1413 gnd 0.008525f
C2373 vdd.n1414 gnd 0.010592f
C2374 vdd.n1415 gnd 0.611584f
C2375 vdd.n1416 gnd 0.828074f
C2376 vdd.n1417 gnd 0.010592f
C2377 vdd.n1418 gnd 0.008525f
C2378 vdd.n1419 gnd 0.010592f
C2379 vdd.n1420 gnd 0.010592f
C2380 vdd.n1421 gnd 0.010592f
C2381 vdd.n1422 gnd 0.008525f
C2382 vdd.n1423 gnd 0.010592f
C2383 vdd.n1424 gnd 0.898433f
C2384 vdd.n1425 gnd 0.010592f
C2385 vdd.n1426 gnd 0.008525f
C2386 vdd.n1427 gnd 0.010592f
C2387 vdd.n1428 gnd 0.010592f
C2388 vdd.n1429 gnd 0.010592f
C2389 vdd.n1430 gnd 0.008525f
C2390 vdd.n1431 gnd 0.010592f
C2391 vdd.t160 gnd 0.541225f
C2392 vdd.n1432 gnd 0.784776f
C2393 vdd.n1433 gnd 0.010592f
C2394 vdd.n1434 gnd 0.008525f
C2395 vdd.n1435 gnd 0.010592f
C2396 vdd.n1436 gnd 0.010592f
C2397 vdd.n1437 gnd 0.010592f
C2398 vdd.n1438 gnd 0.008525f
C2399 vdd.n1439 gnd 0.010592f
C2400 vdd.n1440 gnd 0.600759f
C2401 vdd.n1441 gnd 0.010592f
C2402 vdd.n1442 gnd 0.008525f
C2403 vdd.n1443 gnd 0.010592f
C2404 vdd.n1444 gnd 0.010592f
C2405 vdd.n1445 gnd 0.010592f
C2406 vdd.n1446 gnd 0.008525f
C2407 vdd.n1447 gnd 0.010592f
C2408 vdd.n1448 gnd 0.773951f
C2409 vdd.n1449 gnd 0.665706f
C2410 vdd.n1450 gnd 0.010592f
C2411 vdd.n1451 gnd 0.008525f
C2412 vdd.n1452 gnd 0.008141f
C2413 vdd.n1453 gnd 0.005813f
C2414 vdd.n1454 gnd 0.005394f
C2415 vdd.n1455 gnd 0.002984f
C2416 vdd.n1456 gnd 0.006851f
C2417 vdd.n1457 gnd 0.002899f
C2418 vdd.n1458 gnd 0.003069f
C2419 vdd.n1459 gnd 0.005394f
C2420 vdd.n1460 gnd 0.002899f
C2421 vdd.n1461 gnd 0.006851f
C2422 vdd.n1462 gnd 0.003069f
C2423 vdd.n1463 gnd 0.005394f
C2424 vdd.n1464 gnd 0.002899f
C2425 vdd.n1465 gnd 0.005138f
C2426 vdd.n1466 gnd 0.005154f
C2427 vdd.t115 gnd 0.014719f
C2428 vdd.n1467 gnd 0.03275f
C2429 vdd.n1468 gnd 0.170439f
C2430 vdd.n1469 gnd 0.002899f
C2431 vdd.n1470 gnd 0.003069f
C2432 vdd.n1471 gnd 0.006851f
C2433 vdd.n1472 gnd 0.006851f
C2434 vdd.n1473 gnd 0.003069f
C2435 vdd.n1474 gnd 0.002899f
C2436 vdd.n1475 gnd 0.005394f
C2437 vdd.n1476 gnd 0.005394f
C2438 vdd.n1477 gnd 0.002899f
C2439 vdd.n1478 gnd 0.003069f
C2440 vdd.n1479 gnd 0.006851f
C2441 vdd.n1480 gnd 0.006851f
C2442 vdd.n1481 gnd 0.003069f
C2443 vdd.n1482 gnd 0.002899f
C2444 vdd.n1483 gnd 0.005394f
C2445 vdd.n1484 gnd 0.005394f
C2446 vdd.n1485 gnd 0.002899f
C2447 vdd.n1486 gnd 0.003069f
C2448 vdd.n1487 gnd 0.006851f
C2449 vdd.n1488 gnd 0.006851f
C2450 vdd.n1489 gnd 0.016198f
C2451 vdd.n1490 gnd 0.002984f
C2452 vdd.n1491 gnd 0.002899f
C2453 vdd.n1492 gnd 0.013942f
C2454 vdd.n1493 gnd 0.009734f
C2455 vdd.t175 gnd 0.034101f
C2456 vdd.t224 gnd 0.034101f
C2457 vdd.n1494 gnd 0.234366f
C2458 vdd.n1495 gnd 0.184293f
C2459 vdd.t148 gnd 0.034101f
C2460 vdd.t206 gnd 0.034101f
C2461 vdd.n1496 gnd 0.234366f
C2462 vdd.n1497 gnd 0.148723f
C2463 vdd.t168 gnd 0.034101f
C2464 vdd.t213 gnd 0.034101f
C2465 vdd.n1498 gnd 0.234366f
C2466 vdd.n1499 gnd 0.148723f
C2467 vdd.t188 gnd 0.034101f
C2468 vdd.t231 gnd 0.034101f
C2469 vdd.n1500 gnd 0.234366f
C2470 vdd.n1501 gnd 0.148723f
C2471 vdd.t161 gnd 0.034101f
C2472 vdd.t125 gnd 0.034101f
C2473 vdd.n1502 gnd 0.234366f
C2474 vdd.n1503 gnd 0.148723f
C2475 vdd.t178 gnd 0.034101f
C2476 vdd.t133 gnd 0.034101f
C2477 vdd.n1504 gnd 0.234366f
C2478 vdd.n1505 gnd 0.148723f
C2479 vdd.t220 gnd 0.034101f
C2480 vdd.t236 gnd 0.034101f
C2481 vdd.n1506 gnd 0.234366f
C2482 vdd.n1507 gnd 0.148723f
C2483 vdd.n1508 gnd 0.005813f
C2484 vdd.n1509 gnd 0.005394f
C2485 vdd.n1510 gnd 0.002984f
C2486 vdd.n1511 gnd 0.006851f
C2487 vdd.n1512 gnd 0.002899f
C2488 vdd.n1513 gnd 0.003069f
C2489 vdd.n1514 gnd 0.005394f
C2490 vdd.n1515 gnd 0.002899f
C2491 vdd.n1516 gnd 0.006851f
C2492 vdd.n1517 gnd 0.003069f
C2493 vdd.n1518 gnd 0.005394f
C2494 vdd.n1519 gnd 0.002899f
C2495 vdd.n1520 gnd 0.005138f
C2496 vdd.n1521 gnd 0.005154f
C2497 vdd.t137 gnd 0.014719f
C2498 vdd.n1522 gnd 0.03275f
C2499 vdd.n1523 gnd 0.170439f
C2500 vdd.n1524 gnd 0.002899f
C2501 vdd.n1525 gnd 0.003069f
C2502 vdd.n1526 gnd 0.006851f
C2503 vdd.n1527 gnd 0.006851f
C2504 vdd.n1528 gnd 0.003069f
C2505 vdd.n1529 gnd 0.002899f
C2506 vdd.n1530 gnd 0.005394f
C2507 vdd.n1531 gnd 0.005394f
C2508 vdd.n1532 gnd 0.002899f
C2509 vdd.n1533 gnd 0.003069f
C2510 vdd.n1534 gnd 0.006851f
C2511 vdd.n1535 gnd 0.006851f
C2512 vdd.n1536 gnd 0.003069f
C2513 vdd.n1537 gnd 0.002899f
C2514 vdd.n1538 gnd 0.005394f
C2515 vdd.n1539 gnd 0.005394f
C2516 vdd.n1540 gnd 0.002899f
C2517 vdd.n1541 gnd 0.003069f
C2518 vdd.n1542 gnd 0.006851f
C2519 vdd.n1543 gnd 0.006851f
C2520 vdd.n1544 gnd 0.016198f
C2521 vdd.n1545 gnd 0.002984f
C2522 vdd.n1546 gnd 0.002899f
C2523 vdd.n1547 gnd 0.013942f
C2524 vdd.n1548 gnd 0.009428f
C2525 vdd.n1549 gnd 0.110651f
C2526 vdd.n1550 gnd 0.005813f
C2527 vdd.n1551 gnd 0.005394f
C2528 vdd.n1552 gnd 0.002984f
C2529 vdd.n1553 gnd 0.006851f
C2530 vdd.n1554 gnd 0.002899f
C2531 vdd.n1555 gnd 0.003069f
C2532 vdd.n1556 gnd 0.005394f
C2533 vdd.n1557 gnd 0.002899f
C2534 vdd.n1558 gnd 0.006851f
C2535 vdd.n1559 gnd 0.003069f
C2536 vdd.n1560 gnd 0.005394f
C2537 vdd.n1561 gnd 0.002899f
C2538 vdd.n1562 gnd 0.005138f
C2539 vdd.n1563 gnd 0.005154f
C2540 vdd.t215 gnd 0.014719f
C2541 vdd.n1564 gnd 0.03275f
C2542 vdd.n1565 gnd 0.170439f
C2543 vdd.n1566 gnd 0.002899f
C2544 vdd.n1567 gnd 0.003069f
C2545 vdd.n1568 gnd 0.006851f
C2546 vdd.n1569 gnd 0.006851f
C2547 vdd.n1570 gnd 0.003069f
C2548 vdd.n1571 gnd 0.002899f
C2549 vdd.n1572 gnd 0.005394f
C2550 vdd.n1573 gnd 0.005394f
C2551 vdd.n1574 gnd 0.002899f
C2552 vdd.n1575 gnd 0.003069f
C2553 vdd.n1576 gnd 0.006851f
C2554 vdd.n1577 gnd 0.006851f
C2555 vdd.n1578 gnd 0.003069f
C2556 vdd.n1579 gnd 0.002899f
C2557 vdd.n1580 gnd 0.005394f
C2558 vdd.n1581 gnd 0.005394f
C2559 vdd.n1582 gnd 0.002899f
C2560 vdd.n1583 gnd 0.003069f
C2561 vdd.n1584 gnd 0.006851f
C2562 vdd.n1585 gnd 0.006851f
C2563 vdd.n1586 gnd 0.016198f
C2564 vdd.n1587 gnd 0.002984f
C2565 vdd.n1588 gnd 0.002899f
C2566 vdd.n1589 gnd 0.013942f
C2567 vdd.n1590 gnd 0.009734f
C2568 vdd.t127 gnd 0.034101f
C2569 vdd.t218 gnd 0.034101f
C2570 vdd.n1591 gnd 0.234366f
C2571 vdd.n1592 gnd 0.184293f
C2572 vdd.t211 gnd 0.034101f
C2573 vdd.t199 gnd 0.034101f
C2574 vdd.n1593 gnd 0.234366f
C2575 vdd.n1594 gnd 0.148723f
C2576 vdd.t170 gnd 0.034101f
C2577 vdd.t117 gnd 0.034101f
C2578 vdd.n1595 gnd 0.234366f
C2579 vdd.n1596 gnd 0.148723f
C2580 vdd.t227 gnd 0.034101f
C2581 vdd.t197 gnd 0.034101f
C2582 vdd.n1597 gnd 0.234366f
C2583 vdd.n1598 gnd 0.148723f
C2584 vdd.t194 gnd 0.034101f
C2585 vdd.t149 gnd 0.034101f
C2586 vdd.n1599 gnd 0.234366f
C2587 vdd.n1600 gnd 0.148723f
C2588 vdd.t143 gnd 0.034101f
C2589 vdd.t195 gnd 0.034101f
C2590 vdd.n1601 gnd 0.234366f
C2591 vdd.n1602 gnd 0.148723f
C2592 vdd.t185 gnd 0.034101f
C2593 vdd.t183 gnd 0.034101f
C2594 vdd.n1603 gnd 0.234366f
C2595 vdd.n1604 gnd 0.148723f
C2596 vdd.n1605 gnd 0.005813f
C2597 vdd.n1606 gnd 0.005394f
C2598 vdd.n1607 gnd 0.002984f
C2599 vdd.n1608 gnd 0.006851f
C2600 vdd.n1609 gnd 0.002899f
C2601 vdd.n1610 gnd 0.003069f
C2602 vdd.n1611 gnd 0.005394f
C2603 vdd.n1612 gnd 0.002899f
C2604 vdd.n1613 gnd 0.006851f
C2605 vdd.n1614 gnd 0.003069f
C2606 vdd.n1615 gnd 0.005394f
C2607 vdd.n1616 gnd 0.002899f
C2608 vdd.n1617 gnd 0.005138f
C2609 vdd.n1618 gnd 0.005154f
C2610 vdd.t123 gnd 0.014719f
C2611 vdd.n1619 gnd 0.03275f
C2612 vdd.n1620 gnd 0.170439f
C2613 vdd.n1621 gnd 0.002899f
C2614 vdd.n1622 gnd 0.003069f
C2615 vdd.n1623 gnd 0.006851f
C2616 vdd.n1624 gnd 0.006851f
C2617 vdd.n1625 gnd 0.003069f
C2618 vdd.n1626 gnd 0.002899f
C2619 vdd.n1627 gnd 0.005394f
C2620 vdd.n1628 gnd 0.005394f
C2621 vdd.n1629 gnd 0.002899f
C2622 vdd.n1630 gnd 0.003069f
C2623 vdd.n1631 gnd 0.006851f
C2624 vdd.n1632 gnd 0.006851f
C2625 vdd.n1633 gnd 0.003069f
C2626 vdd.n1634 gnd 0.002899f
C2627 vdd.n1635 gnd 0.005394f
C2628 vdd.n1636 gnd 0.005394f
C2629 vdd.n1637 gnd 0.002899f
C2630 vdd.n1638 gnd 0.003069f
C2631 vdd.n1639 gnd 0.006851f
C2632 vdd.n1640 gnd 0.006851f
C2633 vdd.n1641 gnd 0.016198f
C2634 vdd.n1642 gnd 0.002984f
C2635 vdd.n1643 gnd 0.002899f
C2636 vdd.n1644 gnd 0.013942f
C2637 vdd.n1645 gnd 0.009428f
C2638 vdd.n1646 gnd 0.065826f
C2639 vdd.n1647 gnd 0.237189f
C2640 vdd.n1648 gnd 0.005813f
C2641 vdd.n1649 gnd 0.005394f
C2642 vdd.n1650 gnd 0.002984f
C2643 vdd.n1651 gnd 0.006851f
C2644 vdd.n1652 gnd 0.002899f
C2645 vdd.n1653 gnd 0.003069f
C2646 vdd.n1654 gnd 0.005394f
C2647 vdd.n1655 gnd 0.002899f
C2648 vdd.n1656 gnd 0.006851f
C2649 vdd.n1657 gnd 0.003069f
C2650 vdd.n1658 gnd 0.005394f
C2651 vdd.n1659 gnd 0.002899f
C2652 vdd.n1660 gnd 0.005138f
C2653 vdd.n1661 gnd 0.005154f
C2654 vdd.t228 gnd 0.014719f
C2655 vdd.n1662 gnd 0.03275f
C2656 vdd.n1663 gnd 0.170439f
C2657 vdd.n1664 gnd 0.002899f
C2658 vdd.n1665 gnd 0.003069f
C2659 vdd.n1666 gnd 0.006851f
C2660 vdd.n1667 gnd 0.006851f
C2661 vdd.n1668 gnd 0.003069f
C2662 vdd.n1669 gnd 0.002899f
C2663 vdd.n1670 gnd 0.005394f
C2664 vdd.n1671 gnd 0.005394f
C2665 vdd.n1672 gnd 0.002899f
C2666 vdd.n1673 gnd 0.003069f
C2667 vdd.n1674 gnd 0.006851f
C2668 vdd.n1675 gnd 0.006851f
C2669 vdd.n1676 gnd 0.003069f
C2670 vdd.n1677 gnd 0.002899f
C2671 vdd.n1678 gnd 0.005394f
C2672 vdd.n1679 gnd 0.005394f
C2673 vdd.n1680 gnd 0.002899f
C2674 vdd.n1681 gnd 0.003069f
C2675 vdd.n1682 gnd 0.006851f
C2676 vdd.n1683 gnd 0.006851f
C2677 vdd.n1684 gnd 0.016198f
C2678 vdd.n1685 gnd 0.002984f
C2679 vdd.n1686 gnd 0.002899f
C2680 vdd.n1687 gnd 0.013942f
C2681 vdd.n1688 gnd 0.009734f
C2682 vdd.t141 gnd 0.034101f
C2683 vdd.t229 gnd 0.034101f
C2684 vdd.n1689 gnd 0.234366f
C2685 vdd.n1690 gnd 0.184293f
C2686 vdd.t226 gnd 0.034101f
C2687 vdd.t209 gnd 0.034101f
C2688 vdd.n1691 gnd 0.234366f
C2689 vdd.n1692 gnd 0.148723f
C2690 vdd.t186 gnd 0.034101f
C2691 vdd.t138 gnd 0.034101f
C2692 vdd.n1693 gnd 0.234366f
C2693 vdd.n1694 gnd 0.148723f
C2694 vdd.t237 gnd 0.034101f
C2695 vdd.t207 gnd 0.034101f
C2696 vdd.n1695 gnd 0.234366f
C2697 vdd.n1696 gnd 0.148723f
C2698 vdd.t204 gnd 0.034101f
C2699 vdd.t163 gnd 0.034101f
C2700 vdd.n1697 gnd 0.234366f
C2701 vdd.n1698 gnd 0.148723f
C2702 vdd.t162 gnd 0.034101f
C2703 vdd.t205 gnd 0.034101f
C2704 vdd.n1699 gnd 0.234366f
C2705 vdd.n1700 gnd 0.148723f
C2706 vdd.t193 gnd 0.034101f
C2707 vdd.t192 gnd 0.034101f
C2708 vdd.n1701 gnd 0.234366f
C2709 vdd.n1702 gnd 0.148723f
C2710 vdd.n1703 gnd 0.005813f
C2711 vdd.n1704 gnd 0.005394f
C2712 vdd.n1705 gnd 0.002984f
C2713 vdd.n1706 gnd 0.006851f
C2714 vdd.n1707 gnd 0.002899f
C2715 vdd.n1708 gnd 0.003069f
C2716 vdd.n1709 gnd 0.005394f
C2717 vdd.n1710 gnd 0.002899f
C2718 vdd.n1711 gnd 0.006851f
C2719 vdd.n1712 gnd 0.003069f
C2720 vdd.n1713 gnd 0.005394f
C2721 vdd.n1714 gnd 0.002899f
C2722 vdd.n1715 gnd 0.005138f
C2723 vdd.n1716 gnd 0.005154f
C2724 vdd.t140 gnd 0.014719f
C2725 vdd.n1717 gnd 0.03275f
C2726 vdd.n1718 gnd 0.170439f
C2727 vdd.n1719 gnd 0.002899f
C2728 vdd.n1720 gnd 0.003069f
C2729 vdd.n1721 gnd 0.006851f
C2730 vdd.n1722 gnd 0.006851f
C2731 vdd.n1723 gnd 0.003069f
C2732 vdd.n1724 gnd 0.002899f
C2733 vdd.n1725 gnd 0.005394f
C2734 vdd.n1726 gnd 0.005394f
C2735 vdd.n1727 gnd 0.002899f
C2736 vdd.n1728 gnd 0.003069f
C2737 vdd.n1729 gnd 0.006851f
C2738 vdd.n1730 gnd 0.006851f
C2739 vdd.n1731 gnd 0.003069f
C2740 vdd.n1732 gnd 0.002899f
C2741 vdd.n1733 gnd 0.005394f
C2742 vdd.n1734 gnd 0.005394f
C2743 vdd.n1735 gnd 0.002899f
C2744 vdd.n1736 gnd 0.003069f
C2745 vdd.n1737 gnd 0.006851f
C2746 vdd.n1738 gnd 0.006851f
C2747 vdd.n1739 gnd 0.016198f
C2748 vdd.n1740 gnd 0.002984f
C2749 vdd.n1741 gnd 0.002899f
C2750 vdd.n1742 gnd 0.013942f
C2751 vdd.n1743 gnd 0.009428f
C2752 vdd.n1744 gnd 0.065826f
C2753 vdd.n1745 gnd 0.26562f
C2754 vdd.n1746 gnd 2.53376f
C2755 vdd.n1747 gnd 0.624755f
C2756 vdd.n1748 gnd 0.008141f
C2757 vdd.n1749 gnd 0.010592f
C2758 vdd.n1750 gnd 0.008525f
C2759 vdd.n1751 gnd 0.010592f
C2760 vdd.n1752 gnd 0.849723f
C2761 vdd.n1753 gnd 0.010592f
C2762 vdd.n1754 gnd 0.008525f
C2763 vdd.n1755 gnd 0.010592f
C2764 vdd.n1756 gnd 0.010592f
C2765 vdd.n1757 gnd 0.010592f
C2766 vdd.n1758 gnd 0.008525f
C2767 vdd.n1759 gnd 0.010592f
C2768 vdd.t116 gnd 0.541225f
C2769 vdd.n1760 gnd 0.898433f
C2770 vdd.n1761 gnd 0.010592f
C2771 vdd.n1762 gnd 0.008525f
C2772 vdd.n1763 gnd 0.010592f
C2773 vdd.n1764 gnd 0.010592f
C2774 vdd.n1765 gnd 0.010592f
C2775 vdd.n1766 gnd 0.008525f
C2776 vdd.n1767 gnd 0.010592f
C2777 vdd.n1768 gnd 0.763127f
C2778 vdd.n1769 gnd 0.010592f
C2779 vdd.n1770 gnd 0.008525f
C2780 vdd.n1771 gnd 0.010592f
C2781 vdd.n1772 gnd 0.010592f
C2782 vdd.n1773 gnd 0.010592f
C2783 vdd.n1774 gnd 0.008525f
C2784 vdd.n1775 gnd 0.010592f
C2785 vdd.n1776 gnd 0.898433f
C2786 vdd.t198 gnd 0.541225f
C2787 vdd.n1777 gnd 0.57911f
C2788 vdd.n1778 gnd 0.010592f
C2789 vdd.n1779 gnd 0.008525f
C2790 vdd.n1780 gnd 0.010592f
C2791 vdd.n1781 gnd 0.010592f
C2792 vdd.n1782 gnd 0.010592f
C2793 vdd.n1783 gnd 0.008525f
C2794 vdd.n1784 gnd 0.010592f
C2795 vdd.n1785 gnd 0.687355f
C2796 vdd.n1786 gnd 0.010592f
C2797 vdd.n1787 gnd 0.008525f
C2798 vdd.n1788 gnd 0.010592f
C2799 vdd.n1789 gnd 0.010592f
C2800 vdd.n1790 gnd 0.010592f
C2801 vdd.n1791 gnd 0.008525f
C2802 vdd.n1792 gnd 0.010592f
C2803 vdd.n1793 gnd 0.568286f
C2804 vdd.n1794 gnd 0.871372f
C2805 vdd.n1795 gnd 0.010592f
C2806 vdd.n1796 gnd 0.008525f
C2807 vdd.n1797 gnd 0.010592f
C2808 vdd.n1798 gnd 0.010592f
C2809 vdd.n1799 gnd 0.010592f
C2810 vdd.n1800 gnd 0.008525f
C2811 vdd.n1801 gnd 0.010592f
C2812 vdd.n1802 gnd 1.05539f
C2813 vdd.n1803 gnd 0.010592f
C2814 vdd.n1804 gnd 0.008525f
C2815 vdd.n1805 gnd 0.010592f
C2816 vdd.n1806 gnd 0.010592f
C2817 vdd.n1807 gnd 0.02412f
C2818 vdd.n1808 gnd 0.010592f
C2819 vdd.n1809 gnd 0.010592f
C2820 vdd.n1810 gnd 0.008525f
C2821 vdd.n1811 gnd 0.010592f
C2822 vdd.t20 gnd 0.541225f
C2823 vdd.n1812 gnd 1.02291f
C2824 vdd.n1813 gnd 0.010592f
C2825 vdd.n1814 gnd 0.008525f
C2826 vdd.n1815 gnd 0.010592f
C2827 vdd.n1816 gnd 0.010592f
C2828 vdd.n1817 gnd 0.009109f
C2829 vdd.n1818 gnd 0.008525f
C2830 vdd.n1820 gnd 0.010592f
C2831 vdd.n1822 gnd 0.008525f
C2832 vdd.n1823 gnd 0.010592f
C2833 vdd.n1824 gnd 0.008525f
C2834 vdd.n1826 gnd 0.010592f
C2835 vdd.n1827 gnd 0.008525f
C2836 vdd.n1828 gnd 0.010592f
C2837 vdd.n1829 gnd 0.010592f
C2838 vdd.n1830 gnd 0.010592f
C2839 vdd.n1831 gnd 0.010592f
C2840 vdd.n1832 gnd 0.010592f
C2841 vdd.n1833 gnd 0.008525f
C2842 vdd.n1835 gnd 0.010592f
C2843 vdd.n1836 gnd 0.010592f
C2844 vdd.n1837 gnd 0.010592f
C2845 vdd.n1838 gnd 0.010592f
C2846 vdd.n1839 gnd 0.010592f
C2847 vdd.n1840 gnd 0.008525f
C2848 vdd.n1842 gnd 0.010592f
C2849 vdd.n1843 gnd 0.010592f
C2850 vdd.n1844 gnd 0.010592f
C2851 vdd.n1845 gnd 0.010592f
C2852 vdd.n1846 gnd 0.007119f
C2853 vdd.t38 gnd 0.130309f
C2854 vdd.t37 gnd 0.139265f
C2855 vdd.t36 gnd 0.170182f
C2856 vdd.n1847 gnd 0.218149f
C2857 vdd.n1848 gnd 0.183285f
C2858 vdd.n1850 gnd 0.010592f
C2859 vdd.n1851 gnd 0.010592f
C2860 vdd.n1852 gnd 0.008525f
C2861 vdd.n1853 gnd 0.010592f
C2862 vdd.n1855 gnd 0.010592f
C2863 vdd.n1856 gnd 0.010592f
C2864 vdd.n1857 gnd 0.010592f
C2865 vdd.n1858 gnd 0.010592f
C2866 vdd.n1859 gnd 0.008525f
C2867 vdd.n1861 gnd 0.010592f
C2868 vdd.n1862 gnd 0.010592f
C2869 vdd.n1863 gnd 0.010592f
C2870 vdd.n1864 gnd 0.010592f
C2871 vdd.n1865 gnd 0.010592f
C2872 vdd.n1866 gnd 0.008525f
C2873 vdd.n1868 gnd 0.010592f
C2874 vdd.n1869 gnd 0.010592f
C2875 vdd.n1870 gnd 0.010592f
C2876 vdd.n1871 gnd 0.010592f
C2877 vdd.n1872 gnd 0.010592f
C2878 vdd.n1873 gnd 0.008525f
C2879 vdd.n1875 gnd 0.010592f
C2880 vdd.n1876 gnd 0.010592f
C2881 vdd.n1877 gnd 0.010592f
C2882 vdd.n1878 gnd 0.010592f
C2883 vdd.n1879 gnd 0.010592f
C2884 vdd.n1880 gnd 0.008525f
C2885 vdd.n1882 gnd 0.010592f
C2886 vdd.n1883 gnd 0.010592f
C2887 vdd.n1884 gnd 0.010592f
C2888 vdd.n1885 gnd 0.010592f
C2889 vdd.n1886 gnd 0.00844f
C2890 vdd.t35 gnd 0.130309f
C2891 vdd.t34 gnd 0.139265f
C2892 vdd.t33 gnd 0.170182f
C2893 vdd.n1887 gnd 0.218149f
C2894 vdd.n1888 gnd 0.183285f
C2895 vdd.n1890 gnd 0.010592f
C2896 vdd.n1891 gnd 0.010592f
C2897 vdd.n1892 gnd 0.008525f
C2898 vdd.n1893 gnd 0.010592f
C2899 vdd.n1895 gnd 0.010592f
C2900 vdd.n1896 gnd 0.010592f
C2901 vdd.n1897 gnd 0.010592f
C2902 vdd.n1898 gnd 0.010592f
C2903 vdd.n1899 gnd 0.008525f
C2904 vdd.n1901 gnd 0.010592f
C2905 vdd.n1902 gnd 0.010592f
C2906 vdd.n1903 gnd 0.010592f
C2907 vdd.n1904 gnd 0.010592f
C2908 vdd.n1905 gnd 0.010592f
C2909 vdd.n1906 gnd 0.008525f
C2910 vdd.n1908 gnd 0.010592f
C2911 vdd.n1909 gnd 0.010592f
C2912 vdd.n1910 gnd 0.010592f
C2913 vdd.n1911 gnd 0.010592f
C2914 vdd.n1912 gnd 0.010592f
C2915 vdd.n1913 gnd 0.010592f
C2916 vdd.n1914 gnd 0.008525f
C2917 vdd.n1916 gnd 0.010592f
C2918 vdd.n1918 gnd 0.010592f
C2919 vdd.n1919 gnd 0.008525f
C2920 vdd.n1920 gnd 0.008525f
C2921 vdd.n1921 gnd 0.010592f
C2922 vdd.n1923 gnd 0.010592f
C2923 vdd.n1924 gnd 0.008525f
C2924 vdd.n1925 gnd 0.008525f
C2925 vdd.n1926 gnd 0.010592f
C2926 vdd.n1928 gnd 0.010592f
C2927 vdd.n1929 gnd 0.010592f
C2928 vdd.n1930 gnd 0.008525f
C2929 vdd.n1931 gnd 0.008525f
C2930 vdd.n1932 gnd 0.008525f
C2931 vdd.n1933 gnd 0.010592f
C2932 vdd.n1935 gnd 0.010592f
C2933 vdd.n1936 gnd 0.010592f
C2934 vdd.n1937 gnd 0.008525f
C2935 vdd.n1938 gnd 0.008525f
C2936 vdd.n1939 gnd 0.008525f
C2937 vdd.n1940 gnd 0.010592f
C2938 vdd.n1942 gnd 0.010592f
C2939 vdd.n1943 gnd 0.010592f
C2940 vdd.n1944 gnd 0.008525f
C2941 vdd.n1945 gnd 0.008525f
C2942 vdd.n1946 gnd 0.008525f
C2943 vdd.n1947 gnd 0.010592f
C2944 vdd.n1949 gnd 0.010592f
C2945 vdd.n1950 gnd 0.010592f
C2946 vdd.n1951 gnd 0.008525f
C2947 vdd.n1952 gnd 0.010592f
C2948 vdd.n1953 gnd 0.010592f
C2949 vdd.n1954 gnd 0.010592f
C2950 vdd.n1955 gnd 0.017392f
C2951 vdd.n1956 gnd 0.005797f
C2952 vdd.n1957 gnd 0.008525f
C2953 vdd.n1958 gnd 0.010592f
C2954 vdd.n1960 gnd 0.010592f
C2955 vdd.n1961 gnd 0.010592f
C2956 vdd.n1962 gnd 0.008525f
C2957 vdd.n1963 gnd 0.008525f
C2958 vdd.n1964 gnd 0.008525f
C2959 vdd.n1965 gnd 0.010592f
C2960 vdd.n1967 gnd 0.010592f
C2961 vdd.n1968 gnd 0.010592f
C2962 vdd.n1969 gnd 0.008525f
C2963 vdd.n1970 gnd 0.008525f
C2964 vdd.n1971 gnd 0.008525f
C2965 vdd.n1972 gnd 0.010592f
C2966 vdd.n1974 gnd 0.010592f
C2967 vdd.n1975 gnd 0.010592f
C2968 vdd.n1976 gnd 0.008525f
C2969 vdd.n1977 gnd 0.008525f
C2970 vdd.n1978 gnd 0.008525f
C2971 vdd.n1979 gnd 0.010592f
C2972 vdd.n1981 gnd 0.010592f
C2973 vdd.n1982 gnd 0.010592f
C2974 vdd.n1983 gnd 0.008525f
C2975 vdd.n1984 gnd 0.008525f
C2976 vdd.n1985 gnd 0.008525f
C2977 vdd.n1986 gnd 0.010592f
C2978 vdd.n1988 gnd 0.010592f
C2979 vdd.n1989 gnd 0.010592f
C2980 vdd.n1990 gnd 0.008525f
C2981 vdd.n1991 gnd 0.010592f
C2982 vdd.n1992 gnd 0.010592f
C2983 vdd.n1993 gnd 0.010592f
C2984 vdd.n1994 gnd 0.017392f
C2985 vdd.n1995 gnd 0.007119f
C2986 vdd.n1996 gnd 0.008525f
C2987 vdd.n1997 gnd 0.010592f
C2988 vdd.n1999 gnd 0.010592f
C2989 vdd.n2000 gnd 0.010592f
C2990 vdd.n2001 gnd 0.008525f
C2991 vdd.n2002 gnd 0.008525f
C2992 vdd.n2003 gnd 0.008525f
C2993 vdd.n2004 gnd 0.010592f
C2994 vdd.n2006 gnd 0.010592f
C2995 vdd.n2007 gnd 0.010592f
C2996 vdd.n2008 gnd 0.008525f
C2997 vdd.n2009 gnd 0.008525f
C2998 vdd.n2010 gnd 0.008525f
C2999 vdd.n2011 gnd 0.010592f
C3000 vdd.n2013 gnd 0.010592f
C3001 vdd.n2014 gnd 0.010592f
C3002 vdd.n2016 gnd 0.010592f
C3003 vdd.n2017 gnd 0.008525f
C3004 vdd.n2018 gnd 0.006779f
C3005 vdd.n2019 gnd 0.007203f
C3006 vdd.n2020 gnd 0.007203f
C3007 vdd.n2021 gnd 0.007203f
C3008 vdd.n2022 gnd 0.007203f
C3009 vdd.n2023 gnd 0.007203f
C3010 vdd.n2024 gnd 0.007203f
C3011 vdd.n2025 gnd 0.007203f
C3012 vdd.n2026 gnd 0.007203f
C3013 vdd.n2028 gnd 0.007203f
C3014 vdd.n2029 gnd 0.007203f
C3015 vdd.n2030 gnd 0.007203f
C3016 vdd.n2031 gnd 0.007203f
C3017 vdd.n2032 gnd 0.007203f
C3018 vdd.n2034 gnd 0.007203f
C3019 vdd.n2036 gnd 0.007203f
C3020 vdd.n2037 gnd 0.007203f
C3021 vdd.n2038 gnd 0.007203f
C3022 vdd.n2039 gnd 0.007203f
C3023 vdd.n2040 gnd 0.007203f
C3024 vdd.n2042 gnd 0.007203f
C3025 vdd.n2044 gnd 0.007203f
C3026 vdd.n2045 gnd 0.007203f
C3027 vdd.n2046 gnd 0.007203f
C3028 vdd.n2047 gnd 0.007203f
C3029 vdd.n2048 gnd 0.007203f
C3030 vdd.n2050 gnd 0.007203f
C3031 vdd.n2052 gnd 0.007203f
C3032 vdd.n2053 gnd 0.007203f
C3033 vdd.n2054 gnd 0.007203f
C3034 vdd.n2055 gnd 0.007203f
C3035 vdd.n2056 gnd 0.007203f
C3036 vdd.n2058 gnd 0.007203f
C3037 vdd.n2059 gnd 0.007203f
C3038 vdd.n2060 gnd 0.007203f
C3039 vdd.n2061 gnd 0.007203f
C3040 vdd.n2062 gnd 0.007203f
C3041 vdd.n2063 gnd 0.007203f
C3042 vdd.n2064 gnd 0.007203f
C3043 vdd.n2065 gnd 0.007203f
C3044 vdd.n2066 gnd 0.005243f
C3045 vdd.n2067 gnd 0.007203f
C3046 vdd.t2 gnd 0.291054f
C3047 vdd.t3 gnd 0.29793f
C3048 vdd.t0 gnd 0.190011f
C3049 vdd.n2068 gnd 0.102691f
C3050 vdd.n2069 gnd 0.058249f
C3051 vdd.n2070 gnd 0.010294f
C3052 vdd.n2071 gnd 0.007203f
C3053 vdd.n2072 gnd 0.007203f
C3054 vdd.n2073 gnd 0.438392f
C3055 vdd.n2074 gnd 0.007203f
C3056 vdd.n2075 gnd 0.007203f
C3057 vdd.n2076 gnd 0.007203f
C3058 vdd.n2077 gnd 0.007203f
C3059 vdd.n2078 gnd 0.007203f
C3060 vdd.n2079 gnd 0.007203f
C3061 vdd.n2080 gnd 0.007203f
C3062 vdd.n2081 gnd 0.007203f
C3063 vdd.n2082 gnd 0.007203f
C3064 vdd.n2083 gnd 0.007203f
C3065 vdd.n2084 gnd 0.007203f
C3066 vdd.n2085 gnd 0.007203f
C3067 vdd.n2086 gnd 0.007203f
C3068 vdd.n2087 gnd 0.007203f
C3069 vdd.n2088 gnd 0.007203f
C3070 vdd.n2089 gnd 0.007203f
C3071 vdd.n2090 gnd 0.007203f
C3072 vdd.n2091 gnd 0.007203f
C3073 vdd.n2092 gnd 0.007203f
C3074 vdd.n2093 gnd 0.007203f
C3075 vdd.t55 gnd 0.291054f
C3076 vdd.t56 gnd 0.29793f
C3077 vdd.t54 gnd 0.190011f
C3078 vdd.n2094 gnd 0.102691f
C3079 vdd.n2095 gnd 0.058249f
C3080 vdd.n2096 gnd 0.007203f
C3081 vdd.n2097 gnd 0.007203f
C3082 vdd.n2098 gnd 0.007203f
C3083 vdd.n2099 gnd 0.007203f
C3084 vdd.n2100 gnd 0.007203f
C3085 vdd.n2101 gnd 0.007203f
C3086 vdd.n2103 gnd 0.007203f
C3087 vdd.n2104 gnd 0.007203f
C3088 vdd.n2105 gnd 0.007203f
C3089 vdd.n2106 gnd 0.007203f
C3090 vdd.n2108 gnd 0.007203f
C3091 vdd.n2110 gnd 0.007203f
C3092 vdd.n2111 gnd 0.007203f
C3093 vdd.n2112 gnd 0.007203f
C3094 vdd.n2113 gnd 0.007203f
C3095 vdd.n2114 gnd 0.007203f
C3096 vdd.n2116 gnd 0.007203f
C3097 vdd.n2118 gnd 0.007203f
C3098 vdd.n2119 gnd 0.007203f
C3099 vdd.n2120 gnd 0.007203f
C3100 vdd.n2121 gnd 0.007203f
C3101 vdd.n2122 gnd 0.007203f
C3102 vdd.n2124 gnd 0.007203f
C3103 vdd.n2126 gnd 0.007203f
C3104 vdd.n2127 gnd 0.007203f
C3105 vdd.n2128 gnd 0.005243f
C3106 vdd.n2129 gnd 0.010294f
C3107 vdd.n2130 gnd 0.005561f
C3108 vdd.n2131 gnd 0.007203f
C3109 vdd.n2133 gnd 0.007203f
C3110 vdd.n2134 gnd 0.01709f
C3111 vdd.n2135 gnd 0.01709f
C3112 vdd.n2136 gnd 0.015957f
C3113 vdd.n2137 gnd 0.007203f
C3114 vdd.n2138 gnd 0.007203f
C3115 vdd.n2139 gnd 0.007203f
C3116 vdd.n2140 gnd 0.007203f
C3117 vdd.n2141 gnd 0.007203f
C3118 vdd.n2142 gnd 0.007203f
C3119 vdd.n2143 gnd 0.007203f
C3120 vdd.n2144 gnd 0.007203f
C3121 vdd.n2145 gnd 0.007203f
C3122 vdd.n2146 gnd 0.007203f
C3123 vdd.n2147 gnd 0.007203f
C3124 vdd.n2148 gnd 0.007203f
C3125 vdd.n2149 gnd 0.007203f
C3126 vdd.n2150 gnd 0.007203f
C3127 vdd.n2151 gnd 0.007203f
C3128 vdd.n2152 gnd 0.007203f
C3129 vdd.n2153 gnd 0.007203f
C3130 vdd.n2154 gnd 0.007203f
C3131 vdd.n2155 gnd 0.007203f
C3132 vdd.n2156 gnd 0.007203f
C3133 vdd.n2157 gnd 0.007203f
C3134 vdd.n2158 gnd 0.007203f
C3135 vdd.n2159 gnd 0.007203f
C3136 vdd.n2160 gnd 0.007203f
C3137 vdd.n2161 gnd 0.007203f
C3138 vdd.n2162 gnd 0.007203f
C3139 vdd.n2163 gnd 0.007203f
C3140 vdd.n2164 gnd 0.007203f
C3141 vdd.n2165 gnd 0.007203f
C3142 vdd.n2166 gnd 0.007203f
C3143 vdd.n2167 gnd 0.007203f
C3144 vdd.n2168 gnd 0.007203f
C3145 vdd.n2169 gnd 0.007203f
C3146 vdd.n2170 gnd 0.007203f
C3147 vdd.n2171 gnd 0.007203f
C3148 vdd.n2172 gnd 0.007203f
C3149 vdd.n2173 gnd 0.007203f
C3150 vdd.n2174 gnd 0.232727f
C3151 vdd.n2175 gnd 0.007203f
C3152 vdd.n2176 gnd 0.007203f
C3153 vdd.n2177 gnd 0.007203f
C3154 vdd.n2178 gnd 0.007203f
C3155 vdd.n2179 gnd 0.007203f
C3156 vdd.n2180 gnd 0.007203f
C3157 vdd.n2181 gnd 0.007203f
C3158 vdd.n2182 gnd 0.007203f
C3159 vdd.n2183 gnd 0.007203f
C3160 vdd.n2184 gnd 0.007203f
C3161 vdd.n2185 gnd 0.007203f
C3162 vdd.n2186 gnd 0.007203f
C3163 vdd.n2187 gnd 0.007203f
C3164 vdd.n2188 gnd 0.007203f
C3165 vdd.n2189 gnd 0.007203f
C3166 vdd.n2190 gnd 0.007203f
C3167 vdd.n2191 gnd 0.007203f
C3168 vdd.n2192 gnd 0.007203f
C3169 vdd.n2193 gnd 0.007203f
C3170 vdd.n2194 gnd 0.007203f
C3171 vdd.n2195 gnd 0.015957f
C3172 vdd.n2197 gnd 0.01709f
C3173 vdd.n2198 gnd 0.01709f
C3174 vdd.n2199 gnd 0.007203f
C3175 vdd.n2200 gnd 0.005561f
C3176 vdd.n2201 gnd 0.007203f
C3177 vdd.n2203 gnd 0.007203f
C3178 vdd.n2205 gnd 0.007203f
C3179 vdd.n2206 gnd 0.007203f
C3180 vdd.n2207 gnd 0.007203f
C3181 vdd.n2208 gnd 0.007203f
C3182 vdd.n2209 gnd 0.007203f
C3183 vdd.n2211 gnd 0.007203f
C3184 vdd.n2213 gnd 0.007203f
C3185 vdd.n2214 gnd 0.007203f
C3186 vdd.n2215 gnd 0.007203f
C3187 vdd.n2216 gnd 0.007203f
C3188 vdd.n2217 gnd 0.007203f
C3189 vdd.n2219 gnd 0.007203f
C3190 vdd.n2221 gnd 0.007203f
C3191 vdd.n2222 gnd 0.007203f
C3192 vdd.n2223 gnd 0.007203f
C3193 vdd.n2224 gnd 0.007203f
C3194 vdd.n2225 gnd 0.007203f
C3195 vdd.n2227 gnd 0.007203f
C3196 vdd.n2229 gnd 0.007203f
C3197 vdd.n2230 gnd 0.007203f
C3198 vdd.n2231 gnd 0.021484f
C3199 vdd.n2232 gnd 0.636868f
C3200 vdd.n2234 gnd 0.008525f
C3201 vdd.n2235 gnd 0.008525f
C3202 vdd.n2236 gnd 0.010592f
C3203 vdd.n2238 gnd 0.010592f
C3204 vdd.n2239 gnd 0.010592f
C3205 vdd.n2240 gnd 0.008525f
C3206 vdd.n2241 gnd 0.007076f
C3207 vdd.n2242 gnd 0.024285f
C3208 vdd.n2243 gnd 0.02412f
C3209 vdd.n2244 gnd 0.007076f
C3210 vdd.n2245 gnd 0.02412f
C3211 vdd.n2246 gnd 1.42883f
C3212 vdd.n2247 gnd 0.02412f
C3213 vdd.n2248 gnd 0.024285f
C3214 vdd.n2249 gnd 0.004049f
C3215 vdd.t22 gnd 0.130309f
C3216 vdd.t21 gnd 0.139265f
C3217 vdd.t19 gnd 0.170182f
C3218 vdd.n2250 gnd 0.218149f
C3219 vdd.n2251 gnd 0.183285f
C3220 vdd.n2252 gnd 0.013129f
C3221 vdd.n2253 gnd 0.004476f
C3222 vdd.n2254 gnd 0.009109f
C3223 vdd.n2255 gnd 0.636868f
C3224 vdd.n2256 gnd 0.021484f
C3225 vdd.n2257 gnd 0.007203f
C3226 vdd.n2258 gnd 0.007203f
C3227 vdd.n2259 gnd 0.007203f
C3228 vdd.n2261 gnd 0.007203f
C3229 vdd.n2263 gnd 0.007203f
C3230 vdd.n2264 gnd 0.007203f
C3231 vdd.n2265 gnd 0.007203f
C3232 vdd.n2266 gnd 0.007203f
C3233 vdd.n2267 gnd 0.007203f
C3234 vdd.n2269 gnd 0.007203f
C3235 vdd.n2271 gnd 0.007203f
C3236 vdd.n2272 gnd 0.007203f
C3237 vdd.n2273 gnd 0.007203f
C3238 vdd.n2274 gnd 0.007203f
C3239 vdd.n2275 gnd 0.007203f
C3240 vdd.n2277 gnd 0.007203f
C3241 vdd.n2279 gnd 0.007203f
C3242 vdd.n2280 gnd 0.007203f
C3243 vdd.n2281 gnd 0.007203f
C3244 vdd.n2282 gnd 0.007203f
C3245 vdd.n2283 gnd 0.007203f
C3246 vdd.n2285 gnd 0.007203f
C3247 vdd.n2287 gnd 0.007203f
C3248 vdd.n2288 gnd 0.007203f
C3249 vdd.n2289 gnd 0.01709f
C3250 vdd.n2290 gnd 0.015957f
C3251 vdd.n2291 gnd 0.015957f
C3252 vdd.n2292 gnd 1.0608f
C3253 vdd.n2293 gnd 0.015957f
C3254 vdd.n2294 gnd 0.015957f
C3255 vdd.n2295 gnd 0.007203f
C3256 vdd.n2296 gnd 0.007203f
C3257 vdd.n2297 gnd 0.007203f
C3258 vdd.n2298 gnd 0.460041f
C3259 vdd.n2299 gnd 0.007203f
C3260 vdd.n2300 gnd 0.007203f
C3261 vdd.n2301 gnd 0.007203f
C3262 vdd.n2302 gnd 0.007203f
C3263 vdd.n2303 gnd 0.007203f
C3264 vdd.n2304 gnd 0.736066f
C3265 vdd.n2305 gnd 0.007203f
C3266 vdd.n2306 gnd 0.007203f
C3267 vdd.n2307 gnd 0.007203f
C3268 vdd.n2308 gnd 0.007203f
C3269 vdd.n2309 gnd 0.007203f
C3270 vdd.n2310 gnd 0.736066f
C3271 vdd.n2311 gnd 0.007203f
C3272 vdd.n2312 gnd 0.007203f
C3273 vdd.n2313 gnd 0.006355f
C3274 vdd.n2314 gnd 0.020865f
C3275 vdd.n2315 gnd 0.004449f
C3276 vdd.n2316 gnd 0.007203f
C3277 vdd.n2317 gnd 0.405919f
C3278 vdd.n2318 gnd 0.007203f
C3279 vdd.n2319 gnd 0.007203f
C3280 vdd.n2320 gnd 0.007203f
C3281 vdd.n2321 gnd 0.007203f
C3282 vdd.n2322 gnd 0.007203f
C3283 vdd.n2323 gnd 0.492515f
C3284 vdd.n2324 gnd 0.007203f
C3285 vdd.n2325 gnd 0.007203f
C3286 vdd.n2326 gnd 0.007203f
C3287 vdd.n2327 gnd 0.007203f
C3288 vdd.n2328 gnd 0.007203f
C3289 vdd.n2329 gnd 0.654882f
C3290 vdd.n2330 gnd 0.007203f
C3291 vdd.n2331 gnd 0.007203f
C3292 vdd.n2332 gnd 0.007203f
C3293 vdd.n2333 gnd 0.007203f
C3294 vdd.n2334 gnd 0.007203f
C3295 vdd.n2335 gnd 0.584523f
C3296 vdd.n2336 gnd 0.007203f
C3297 vdd.n2337 gnd 0.007203f
C3298 vdd.n2338 gnd 0.007203f
C3299 vdd.n2339 gnd 0.007203f
C3300 vdd.n2340 gnd 0.007203f
C3301 vdd.n2341 gnd 0.422155f
C3302 vdd.n2342 gnd 0.007203f
C3303 vdd.n2343 gnd 0.007203f
C3304 vdd.n2344 gnd 0.007203f
C3305 vdd.n2345 gnd 0.007203f
C3306 vdd.n2346 gnd 0.007203f
C3307 vdd.n2347 gnd 0.232727f
C3308 vdd.n2348 gnd 0.007203f
C3309 vdd.n2349 gnd 0.007203f
C3310 vdd.n2350 gnd 0.007203f
C3311 vdd.n2351 gnd 0.007203f
C3312 vdd.n2352 gnd 0.007203f
C3313 vdd.n2353 gnd 0.405919f
C3314 vdd.n2354 gnd 0.007203f
C3315 vdd.n2355 gnd 0.007203f
C3316 vdd.n2356 gnd 0.007203f
C3317 vdd.n2357 gnd 0.007203f
C3318 vdd.n2358 gnd 0.007203f
C3319 vdd.n2359 gnd 0.736066f
C3320 vdd.n2360 gnd 0.007203f
C3321 vdd.n2361 gnd 0.007203f
C3322 vdd.n2362 gnd 0.007203f
C3323 vdd.n2363 gnd 0.007203f
C3324 vdd.n2364 gnd 0.007203f
C3325 vdd.n2365 gnd 0.007203f
C3326 vdd.n2366 gnd 0.007203f
C3327 vdd.n2367 gnd 0.573698f
C3328 vdd.n2368 gnd 0.007203f
C3329 vdd.n2369 gnd 0.007203f
C3330 vdd.n2370 gnd 0.007203f
C3331 vdd.n2371 gnd 0.007203f
C3332 vdd.n2372 gnd 0.007203f
C3333 vdd.n2373 gnd 0.007203f
C3334 vdd.n2374 gnd 0.460041f
C3335 vdd.n2375 gnd 0.007203f
C3336 vdd.n2376 gnd 0.007203f
C3337 vdd.n2377 gnd 0.007203f
C3338 vdd.n2378 gnd 0.016834f
C3339 vdd.n2379 gnd 0.016213f
C3340 vdd.n2380 gnd 0.007203f
C3341 vdd.n2381 gnd 0.007203f
C3342 vdd.n2382 gnd 0.005561f
C3343 vdd.n2383 gnd 0.007203f
C3344 vdd.n2384 gnd 0.007203f
C3345 vdd.n2385 gnd 0.005243f
C3346 vdd.n2386 gnd 0.007203f
C3347 vdd.n2387 gnd 0.007203f
C3348 vdd.n2388 gnd 0.007203f
C3349 vdd.n2389 gnd 0.007203f
C3350 vdd.n2390 gnd 0.007203f
C3351 vdd.n2391 gnd 0.007203f
C3352 vdd.n2392 gnd 0.007203f
C3353 vdd.n2393 gnd 0.007203f
C3354 vdd.n2394 gnd 0.007203f
C3355 vdd.n2395 gnd 0.007203f
C3356 vdd.n2396 gnd 0.007203f
C3357 vdd.n2397 gnd 0.007203f
C3358 vdd.n2398 gnd 0.007203f
C3359 vdd.n2399 gnd 0.007203f
C3360 vdd.n2400 gnd 0.007203f
C3361 vdd.n2401 gnd 0.007203f
C3362 vdd.n2402 gnd 0.007203f
C3363 vdd.n2403 gnd 0.007203f
C3364 vdd.n2404 gnd 0.007203f
C3365 vdd.n2405 gnd 0.007203f
C3366 vdd.n2406 gnd 0.007203f
C3367 vdd.n2407 gnd 0.007203f
C3368 vdd.n2408 gnd 0.007203f
C3369 vdd.n2409 gnd 0.007203f
C3370 vdd.n2410 gnd 0.007203f
C3371 vdd.n2411 gnd 0.007203f
C3372 vdd.n2412 gnd 0.007203f
C3373 vdd.n2413 gnd 0.007203f
C3374 vdd.n2414 gnd 0.007203f
C3375 vdd.n2415 gnd 0.007203f
C3376 vdd.n2416 gnd 0.007203f
C3377 vdd.n2417 gnd 0.007203f
C3378 vdd.n2418 gnd 0.007203f
C3379 vdd.n2419 gnd 0.007203f
C3380 vdd.n2420 gnd 0.007203f
C3381 vdd.n2421 gnd 0.007203f
C3382 vdd.n2422 gnd 0.007203f
C3383 vdd.n2423 gnd 0.007203f
C3384 vdd.n2424 gnd 0.007203f
C3385 vdd.n2425 gnd 0.007203f
C3386 vdd.n2426 gnd 0.007203f
C3387 vdd.n2427 gnd 0.007203f
C3388 vdd.n2428 gnd 0.007203f
C3389 vdd.n2429 gnd 0.007203f
C3390 vdd.n2430 gnd 0.007203f
C3391 vdd.n2431 gnd 0.007203f
C3392 vdd.n2432 gnd 0.007203f
C3393 vdd.n2433 gnd 0.007203f
C3394 vdd.n2434 gnd 0.007203f
C3395 vdd.n2435 gnd 0.007203f
C3396 vdd.n2436 gnd 0.007203f
C3397 vdd.n2437 gnd 0.007203f
C3398 vdd.n2438 gnd 0.007203f
C3399 vdd.n2439 gnd 0.007203f
C3400 vdd.n2440 gnd 0.007203f
C3401 vdd.n2441 gnd 0.007203f
C3402 vdd.n2442 gnd 0.007203f
C3403 vdd.n2443 gnd 0.007203f
C3404 vdd.n2444 gnd 0.007203f
C3405 vdd.n2445 gnd 0.007203f
C3406 vdd.n2446 gnd 0.01709f
C3407 vdd.n2447 gnd 0.015957f
C3408 vdd.n2448 gnd 0.015957f
C3409 vdd.n2449 gnd 0.898433f
C3410 vdd.n2450 gnd 0.015957f
C3411 vdd.n2451 gnd 0.01709f
C3412 vdd.n2452 gnd 0.016213f
C3413 vdd.n2453 gnd 0.007203f
C3414 vdd.n2454 gnd 0.007203f
C3415 vdd.n2455 gnd 0.007203f
C3416 vdd.n2456 gnd 0.005561f
C3417 vdd.n2457 gnd 0.010294f
C3418 vdd.n2458 gnd 0.005243f
C3419 vdd.n2459 gnd 0.007203f
C3420 vdd.n2460 gnd 0.007203f
C3421 vdd.n2461 gnd 0.007203f
C3422 vdd.n2462 gnd 0.007203f
C3423 vdd.n2463 gnd 0.007203f
C3424 vdd.n2464 gnd 0.007203f
C3425 vdd.n2465 gnd 0.007203f
C3426 vdd.n2466 gnd 0.007203f
C3427 vdd.n2467 gnd 0.007203f
C3428 vdd.n2468 gnd 0.007203f
C3429 vdd.n2469 gnd 0.007203f
C3430 vdd.n2470 gnd 0.007203f
C3431 vdd.n2471 gnd 0.007203f
C3432 vdd.n2472 gnd 0.007203f
C3433 vdd.n2473 gnd 0.007203f
C3434 vdd.n2474 gnd 0.007203f
C3435 vdd.n2475 gnd 0.007203f
C3436 vdd.n2476 gnd 0.007203f
C3437 vdd.n2477 gnd 0.007203f
C3438 vdd.n2478 gnd 0.007203f
C3439 vdd.n2479 gnd 0.007203f
C3440 vdd.n2480 gnd 0.007203f
C3441 vdd.n2481 gnd 0.007203f
C3442 vdd.n2482 gnd 0.007203f
C3443 vdd.n2483 gnd 0.007203f
C3444 vdd.n2484 gnd 0.007203f
C3445 vdd.n2485 gnd 0.007203f
C3446 vdd.n2486 gnd 0.007203f
C3447 vdd.n2487 gnd 0.007203f
C3448 vdd.n2488 gnd 0.007203f
C3449 vdd.n2489 gnd 0.007203f
C3450 vdd.n2490 gnd 0.007203f
C3451 vdd.n2491 gnd 0.007203f
C3452 vdd.n2492 gnd 0.007203f
C3453 vdd.n2493 gnd 0.007203f
C3454 vdd.n2494 gnd 0.007203f
C3455 vdd.n2495 gnd 0.007203f
C3456 vdd.n2496 gnd 0.007203f
C3457 vdd.n2497 gnd 0.007203f
C3458 vdd.n2498 gnd 0.007203f
C3459 vdd.n2499 gnd 0.007203f
C3460 vdd.n2500 gnd 0.007203f
C3461 vdd.n2501 gnd 0.007203f
C3462 vdd.n2502 gnd 0.007203f
C3463 vdd.n2503 gnd 0.007203f
C3464 vdd.n2504 gnd 0.007203f
C3465 vdd.n2505 gnd 0.007203f
C3466 vdd.n2506 gnd 0.007203f
C3467 vdd.n2507 gnd 0.007203f
C3468 vdd.n2508 gnd 0.007203f
C3469 vdd.n2509 gnd 0.007203f
C3470 vdd.n2510 gnd 0.007203f
C3471 vdd.n2511 gnd 0.007203f
C3472 vdd.n2512 gnd 0.007203f
C3473 vdd.n2513 gnd 0.007203f
C3474 vdd.n2514 gnd 0.007203f
C3475 vdd.n2515 gnd 0.007203f
C3476 vdd.n2516 gnd 0.007203f
C3477 vdd.n2517 gnd 0.007203f
C3478 vdd.n2518 gnd 0.007203f
C3479 vdd.n2519 gnd 0.01709f
C3480 vdd.n2520 gnd 0.01709f
C3481 vdd.n2521 gnd 0.898433f
C3482 vdd.t252 gnd 3.19323f
C3483 vdd.t238 gnd 3.19323f
C3484 vdd.n2554 gnd 0.01709f
C3485 vdd.n2555 gnd 0.007203f
C3486 vdd.t49 gnd 0.291054f
C3487 vdd.t50 gnd 0.29793f
C3488 vdd.t47 gnd 0.190011f
C3489 vdd.n2556 gnd 0.102691f
C3490 vdd.n2557 gnd 0.058249f
C3491 vdd.n2558 gnd 0.007203f
C3492 vdd.t62 gnd 0.291054f
C3493 vdd.t63 gnd 0.29793f
C3494 vdd.t61 gnd 0.190011f
C3495 vdd.n2559 gnd 0.102691f
C3496 vdd.n2560 gnd 0.058249f
C3497 vdd.n2561 gnd 0.010294f
C3498 vdd.n2562 gnd 0.007203f
C3499 vdd.n2563 gnd 0.007203f
C3500 vdd.n2564 gnd 0.007203f
C3501 vdd.n2565 gnd 0.007203f
C3502 vdd.n2566 gnd 0.007203f
C3503 vdd.n2567 gnd 0.007203f
C3504 vdd.n2568 gnd 0.007203f
C3505 vdd.n2569 gnd 0.007203f
C3506 vdd.n2570 gnd 0.007203f
C3507 vdd.n2571 gnd 0.007203f
C3508 vdd.n2572 gnd 0.007203f
C3509 vdd.n2573 gnd 0.007203f
C3510 vdd.n2574 gnd 0.007203f
C3511 vdd.n2575 gnd 0.007203f
C3512 vdd.n2576 gnd 0.007203f
C3513 vdd.n2577 gnd 0.007203f
C3514 vdd.n2578 gnd 0.007203f
C3515 vdd.n2579 gnd 0.007203f
C3516 vdd.n2580 gnd 0.007203f
C3517 vdd.n2581 gnd 0.007203f
C3518 vdd.n2582 gnd 0.007203f
C3519 vdd.n2583 gnd 0.007203f
C3520 vdd.n2584 gnd 0.007203f
C3521 vdd.n2585 gnd 0.007203f
C3522 vdd.n2586 gnd 0.007203f
C3523 vdd.n2587 gnd 0.007203f
C3524 vdd.n2588 gnd 0.007203f
C3525 vdd.n2589 gnd 0.007203f
C3526 vdd.n2590 gnd 0.007203f
C3527 vdd.n2591 gnd 0.007203f
C3528 vdd.n2592 gnd 0.007203f
C3529 vdd.n2593 gnd 0.007203f
C3530 vdd.n2594 gnd 0.007203f
C3531 vdd.n2595 gnd 0.007203f
C3532 vdd.n2596 gnd 0.007203f
C3533 vdd.n2597 gnd 0.007203f
C3534 vdd.n2598 gnd 0.007203f
C3535 vdd.n2599 gnd 0.007203f
C3536 vdd.n2600 gnd 0.007203f
C3537 vdd.n2601 gnd 0.007203f
C3538 vdd.n2602 gnd 0.007203f
C3539 vdd.n2603 gnd 0.007203f
C3540 vdd.n2604 gnd 0.007203f
C3541 vdd.n2605 gnd 0.007203f
C3542 vdd.n2606 gnd 0.007203f
C3543 vdd.n2607 gnd 0.007203f
C3544 vdd.n2608 gnd 0.007203f
C3545 vdd.n2609 gnd 0.007203f
C3546 vdd.n2610 gnd 0.007203f
C3547 vdd.n2611 gnd 0.007203f
C3548 vdd.n2612 gnd 0.007203f
C3549 vdd.n2613 gnd 0.007203f
C3550 vdd.n2614 gnd 0.007203f
C3551 vdd.n2615 gnd 0.007203f
C3552 vdd.n2616 gnd 0.007203f
C3553 vdd.n2617 gnd 0.007203f
C3554 vdd.n2618 gnd 0.005243f
C3555 vdd.n2619 gnd 0.007203f
C3556 vdd.n2620 gnd 0.007203f
C3557 vdd.n2621 gnd 0.005561f
C3558 vdd.n2622 gnd 0.007203f
C3559 vdd.n2623 gnd 0.007203f
C3560 vdd.n2624 gnd 0.01709f
C3561 vdd.n2625 gnd 0.015957f
C3562 vdd.n2626 gnd 0.007203f
C3563 vdd.n2627 gnd 0.007203f
C3564 vdd.n2628 gnd 0.007203f
C3565 vdd.n2629 gnd 0.007203f
C3566 vdd.n2630 gnd 0.007203f
C3567 vdd.n2631 gnd 0.007203f
C3568 vdd.n2632 gnd 0.007203f
C3569 vdd.n2633 gnd 0.007203f
C3570 vdd.n2634 gnd 0.007203f
C3571 vdd.n2635 gnd 0.007203f
C3572 vdd.n2636 gnd 0.007203f
C3573 vdd.n2637 gnd 0.007203f
C3574 vdd.n2638 gnd 0.007203f
C3575 vdd.n2639 gnd 0.007203f
C3576 vdd.n2640 gnd 0.007203f
C3577 vdd.n2641 gnd 0.007203f
C3578 vdd.n2642 gnd 0.007203f
C3579 vdd.n2643 gnd 0.007203f
C3580 vdd.n2644 gnd 0.007203f
C3581 vdd.n2645 gnd 0.007203f
C3582 vdd.n2646 gnd 0.007203f
C3583 vdd.n2647 gnd 0.007203f
C3584 vdd.n2648 gnd 0.007203f
C3585 vdd.n2649 gnd 0.007203f
C3586 vdd.n2650 gnd 0.007203f
C3587 vdd.n2651 gnd 0.007203f
C3588 vdd.n2652 gnd 0.007203f
C3589 vdd.n2653 gnd 0.007203f
C3590 vdd.n2654 gnd 0.007203f
C3591 vdd.n2655 gnd 0.007203f
C3592 vdd.n2656 gnd 0.007203f
C3593 vdd.n2657 gnd 0.007203f
C3594 vdd.n2658 gnd 0.007203f
C3595 vdd.n2659 gnd 0.007203f
C3596 vdd.n2660 gnd 0.007203f
C3597 vdd.n2661 gnd 0.007203f
C3598 vdd.n2662 gnd 0.007203f
C3599 vdd.n2663 gnd 0.007203f
C3600 vdd.n2664 gnd 0.007203f
C3601 vdd.n2665 gnd 0.007203f
C3602 vdd.n2666 gnd 0.007203f
C3603 vdd.n2667 gnd 0.007203f
C3604 vdd.n2668 gnd 0.007203f
C3605 vdd.n2669 gnd 0.007203f
C3606 vdd.n2670 gnd 0.007203f
C3607 vdd.n2671 gnd 0.007203f
C3608 vdd.n2672 gnd 0.007203f
C3609 vdd.n2673 gnd 0.007203f
C3610 vdd.n2674 gnd 0.007203f
C3611 vdd.n2675 gnd 0.007203f
C3612 vdd.n2676 gnd 0.007203f
C3613 vdd.n2677 gnd 0.232727f
C3614 vdd.n2678 gnd 0.007203f
C3615 vdd.n2679 gnd 0.007203f
C3616 vdd.n2680 gnd 0.007203f
C3617 vdd.n2681 gnd 0.007203f
C3618 vdd.n2682 gnd 0.007203f
C3619 vdd.n2683 gnd 0.007203f
C3620 vdd.n2684 gnd 0.007203f
C3621 vdd.n2685 gnd 0.007203f
C3622 vdd.n2686 gnd 0.007203f
C3623 vdd.n2687 gnd 0.007203f
C3624 vdd.n2688 gnd 0.007203f
C3625 vdd.n2689 gnd 0.007203f
C3626 vdd.n2690 gnd 0.007203f
C3627 vdd.n2691 gnd 0.007203f
C3628 vdd.n2692 gnd 0.007203f
C3629 vdd.n2693 gnd 0.007203f
C3630 vdd.n2694 gnd 0.007203f
C3631 vdd.n2695 gnd 0.007203f
C3632 vdd.n2696 gnd 0.007203f
C3633 vdd.n2697 gnd 0.007203f
C3634 vdd.n2698 gnd 0.438392f
C3635 vdd.n2699 gnd 0.007203f
C3636 vdd.n2700 gnd 0.007203f
C3637 vdd.n2701 gnd 0.007203f
C3638 vdd.n2702 gnd 0.007203f
C3639 vdd.n2703 gnd 0.007203f
C3640 vdd.n2704 gnd 0.015957f
C3641 vdd.n2705 gnd 0.01709f
C3642 vdd.n2706 gnd 0.01709f
C3643 vdd.n2707 gnd 0.007203f
C3644 vdd.n2708 gnd 0.007203f
C3645 vdd.n2709 gnd 0.007203f
C3646 vdd.n2710 gnd 0.005561f
C3647 vdd.n2711 gnd 0.010294f
C3648 vdd.n2712 gnd 0.005243f
C3649 vdd.n2713 gnd 0.007203f
C3650 vdd.n2714 gnd 0.007203f
C3651 vdd.n2715 gnd 0.007203f
C3652 vdd.n2716 gnd 0.007203f
C3653 vdd.n2717 gnd 0.007203f
C3654 vdd.n2718 gnd 0.007203f
C3655 vdd.n2719 gnd 0.007203f
C3656 vdd.n2720 gnd 0.007203f
C3657 vdd.n2721 gnd 0.007203f
C3658 vdd.n2722 gnd 0.007203f
C3659 vdd.n2723 gnd 0.007203f
C3660 vdd.n2724 gnd 0.007203f
C3661 vdd.n2725 gnd 0.007203f
C3662 vdd.n2726 gnd 0.007203f
C3663 vdd.n2727 gnd 0.007203f
C3664 vdd.n2728 gnd 0.007203f
C3665 vdd.n2729 gnd 0.007203f
C3666 vdd.n2730 gnd 0.007203f
C3667 vdd.n2731 gnd 0.007203f
C3668 vdd.n2732 gnd 0.007203f
C3669 vdd.n2733 gnd 0.007203f
C3670 vdd.n2734 gnd 0.007203f
C3671 vdd.n2735 gnd 0.007203f
C3672 vdd.n2736 gnd 0.007203f
C3673 vdd.n2737 gnd 0.007203f
C3674 vdd.n2738 gnd 0.007203f
C3675 vdd.n2739 gnd 0.007203f
C3676 vdd.n2740 gnd 0.007203f
C3677 vdd.n2741 gnd 0.007203f
C3678 vdd.n2742 gnd 0.007203f
C3679 vdd.n2743 gnd 0.007203f
C3680 vdd.n2744 gnd 0.007203f
C3681 vdd.n2745 gnd 0.007203f
C3682 vdd.n2746 gnd 0.007203f
C3683 vdd.n2747 gnd 0.007203f
C3684 vdd.n2748 gnd 0.007203f
C3685 vdd.n2749 gnd 0.007203f
C3686 vdd.n2750 gnd 0.007203f
C3687 vdd.n2751 gnd 0.007203f
C3688 vdd.n2752 gnd 0.007203f
C3689 vdd.n2753 gnd 0.007203f
C3690 vdd.n2754 gnd 0.007203f
C3691 vdd.n2755 gnd 0.007203f
C3692 vdd.n2756 gnd 0.007203f
C3693 vdd.n2757 gnd 0.007203f
C3694 vdd.n2758 gnd 0.007203f
C3695 vdd.n2759 gnd 0.007203f
C3696 vdd.n2760 gnd 0.007203f
C3697 vdd.n2761 gnd 0.007203f
C3698 vdd.n2762 gnd 0.007203f
C3699 vdd.n2763 gnd 0.007203f
C3700 vdd.n2764 gnd 0.007203f
C3701 vdd.n2765 gnd 0.007203f
C3702 vdd.n2766 gnd 0.007203f
C3703 vdd.n2767 gnd 0.007203f
C3704 vdd.n2768 gnd 0.007203f
C3705 vdd.n2769 gnd 0.007203f
C3706 vdd.n2770 gnd 0.007203f
C3707 vdd.n2771 gnd 0.007203f
C3708 vdd.n2772 gnd 0.007203f
C3709 vdd.n2774 gnd 0.898433f
C3710 vdd.n2776 gnd 0.007203f
C3711 vdd.n2777 gnd 0.007203f
C3712 vdd.n2778 gnd 0.01709f
C3713 vdd.n2779 gnd 0.015957f
C3714 vdd.n2780 gnd 0.015957f
C3715 vdd.n2781 gnd 0.898433f
C3716 vdd.n2782 gnd 0.015957f
C3717 vdd.n2783 gnd 0.015957f
C3718 vdd.n2784 gnd 0.007203f
C3719 vdd.n2785 gnd 0.007203f
C3720 vdd.n2786 gnd 0.007203f
C3721 vdd.n2787 gnd 0.460041f
C3722 vdd.n2788 gnd 0.007203f
C3723 vdd.n2789 gnd 0.007203f
C3724 vdd.n2790 gnd 0.007203f
C3725 vdd.n2791 gnd 0.007203f
C3726 vdd.n2792 gnd 0.007203f
C3727 vdd.n2793 gnd 0.573698f
C3728 vdd.n2794 gnd 0.007203f
C3729 vdd.n2795 gnd 0.007203f
C3730 vdd.n2796 gnd 0.007203f
C3731 vdd.n2797 gnd 0.007203f
C3732 vdd.n2798 gnd 0.007203f
C3733 vdd.n2799 gnd 0.736066f
C3734 vdd.n2800 gnd 0.007203f
C3735 vdd.n2801 gnd 0.007203f
C3736 vdd.n2802 gnd 0.007203f
C3737 vdd.n2803 gnd 0.007203f
C3738 vdd.n2804 gnd 0.007203f
C3739 vdd.n2805 gnd 0.405919f
C3740 vdd.n2806 gnd 0.007203f
C3741 vdd.n2807 gnd 0.007203f
C3742 vdd.n2808 gnd 0.007203f
C3743 vdd.n2809 gnd 0.007203f
C3744 vdd.n2810 gnd 0.007203f
C3745 vdd.n2811 gnd 0.232727f
C3746 vdd.n2812 gnd 0.007203f
C3747 vdd.n2813 gnd 0.007203f
C3748 vdd.n2814 gnd 0.007203f
C3749 vdd.n2815 gnd 0.007203f
C3750 vdd.n2816 gnd 0.007203f
C3751 vdd.n2817 gnd 0.422155f
C3752 vdd.n2818 gnd 0.007203f
C3753 vdd.n2819 gnd 0.007203f
C3754 vdd.n2820 gnd 0.007203f
C3755 vdd.n2821 gnd 0.007203f
C3756 vdd.n2822 gnd 0.007203f
C3757 vdd.n2823 gnd 0.584523f
C3758 vdd.n2824 gnd 0.007203f
C3759 vdd.n2825 gnd 0.007203f
C3760 vdd.n2826 gnd 0.007203f
C3761 vdd.n2827 gnd 0.007203f
C3762 vdd.n2828 gnd 0.007203f
C3763 vdd.n2829 gnd 0.654882f
C3764 vdd.n2830 gnd 0.007203f
C3765 vdd.n2831 gnd 0.007203f
C3766 vdd.n2832 gnd 0.007203f
C3767 vdd.n2833 gnd 0.007203f
C3768 vdd.n2834 gnd 0.007203f
C3769 vdd.n2835 gnd 0.492515f
C3770 vdd.n2836 gnd 0.007203f
C3771 vdd.n2837 gnd 0.007203f
C3772 vdd.n2838 gnd 0.007203f
C3773 vdd.t28 gnd 0.29793f
C3774 vdd.t26 gnd 0.190011f
C3775 vdd.t29 gnd 0.29793f
C3776 vdd.n2839 gnd 0.167449f
C3777 vdd.n2840 gnd 0.020865f
C3778 vdd.n2841 gnd 0.004449f
C3779 vdd.n2842 gnd 0.007203f
C3780 vdd.n2843 gnd 0.405919f
C3781 vdd.n2844 gnd 0.007203f
C3782 vdd.n2845 gnd 0.007203f
C3783 vdd.n2846 gnd 0.007203f
C3784 vdd.n2847 gnd 0.007203f
C3785 vdd.n2848 gnd 0.007203f
C3786 vdd.n2849 gnd 0.736066f
C3787 vdd.n2850 gnd 0.007203f
C3788 vdd.n2851 gnd 0.007203f
C3789 vdd.n2852 gnd 0.007203f
C3790 vdd.n2853 gnd 0.007203f
C3791 vdd.n2854 gnd 0.007203f
C3792 vdd.n2855 gnd 0.007203f
C3793 vdd.n2857 gnd 0.007203f
C3794 vdd.n2858 gnd 0.007203f
C3795 vdd.n2860 gnd 0.007203f
C3796 vdd.n2861 gnd 0.007203f
C3797 vdd.n2864 gnd 0.007203f
C3798 vdd.n2865 gnd 0.007203f
C3799 vdd.n2866 gnd 0.007203f
C3800 vdd.n2867 gnd 0.007203f
C3801 vdd.n2869 gnd 0.007203f
C3802 vdd.n2870 gnd 0.007203f
C3803 vdd.n2871 gnd 0.007203f
C3804 vdd.n2872 gnd 0.007203f
C3805 vdd.n2873 gnd 0.007203f
C3806 vdd.n2874 gnd 0.007203f
C3807 vdd.n2876 gnd 0.007203f
C3808 vdd.n2877 gnd 0.007203f
C3809 vdd.n2878 gnd 0.007203f
C3810 vdd.n2879 gnd 0.007203f
C3811 vdd.n2880 gnd 0.007203f
C3812 vdd.n2881 gnd 0.007203f
C3813 vdd.n2883 gnd 0.007203f
C3814 vdd.n2884 gnd 0.007203f
C3815 vdd.n2885 gnd 0.007203f
C3816 vdd.n2886 gnd 0.007203f
C3817 vdd.n2887 gnd 0.007203f
C3818 vdd.n2888 gnd 0.007203f
C3819 vdd.n2890 gnd 0.007203f
C3820 vdd.n2891 gnd 0.01709f
C3821 vdd.n2892 gnd 0.01709f
C3822 vdd.n2893 gnd 0.015957f
C3823 vdd.n2894 gnd 0.007203f
C3824 vdd.n2895 gnd 0.007203f
C3825 vdd.n2896 gnd 0.007203f
C3826 vdd.n2897 gnd 0.007203f
C3827 vdd.n2898 gnd 0.007203f
C3828 vdd.n2899 gnd 0.007203f
C3829 vdd.n2900 gnd 0.736066f
C3830 vdd.n2901 gnd 0.007203f
C3831 vdd.n2902 gnd 0.007203f
C3832 vdd.n2903 gnd 0.007203f
C3833 vdd.n2904 gnd 0.007203f
C3834 vdd.n2905 gnd 0.007203f
C3835 vdd.n2906 gnd 0.460041f
C3836 vdd.n2907 gnd 0.007203f
C3837 vdd.n2908 gnd 0.007203f
C3838 vdd.n2909 gnd 0.007203f
C3839 vdd.n2910 gnd 0.016834f
C3840 vdd.n2912 gnd 0.01709f
C3841 vdd.n2913 gnd 0.016213f
C3842 vdd.n2914 gnd 0.007203f
C3843 vdd.n2915 gnd 0.005561f
C3844 vdd.n2916 gnd 0.007203f
C3845 vdd.n2918 gnd 0.007203f
C3846 vdd.n2919 gnd 0.007203f
C3847 vdd.n2920 gnd 0.007203f
C3848 vdd.n2921 gnd 0.007203f
C3849 vdd.n2922 gnd 0.007203f
C3850 vdd.n2923 gnd 0.007203f
C3851 vdd.n2925 gnd 0.007203f
C3852 vdd.n2926 gnd 0.007203f
C3853 vdd.n2927 gnd 0.007203f
C3854 vdd.n2928 gnd 0.007203f
C3855 vdd.n2929 gnd 0.007203f
C3856 vdd.n2930 gnd 0.007203f
C3857 vdd.n2932 gnd 0.007203f
C3858 vdd.n2933 gnd 0.007203f
C3859 vdd.n2934 gnd 0.007203f
C3860 vdd.n2935 gnd 0.007203f
C3861 vdd.n2936 gnd 0.007203f
C3862 vdd.n2937 gnd 0.007203f
C3863 vdd.n2939 gnd 0.007203f
C3864 vdd.n2940 gnd 0.007203f
C3865 vdd.n2941 gnd 0.007203f
C3866 vdd.n2942 gnd 0.641044f
C3867 vdd.n2943 gnd 0.017308f
C3868 vdd.n2944 gnd 0.007203f
C3869 vdd.n2945 gnd 0.007203f
C3870 vdd.n2947 gnd 0.007203f
C3871 vdd.n2948 gnd 0.007203f
C3872 vdd.n2949 gnd 0.007203f
C3873 vdd.n2950 gnd 0.007203f
C3874 vdd.n2951 gnd 0.007203f
C3875 vdd.n2952 gnd 0.007203f
C3876 vdd.n2954 gnd 0.007203f
C3877 vdd.n2955 gnd 0.007203f
C3878 vdd.n2956 gnd 0.007203f
C3879 vdd.n2957 gnd 0.007203f
C3880 vdd.n2958 gnd 0.007203f
C3881 vdd.n2959 gnd 0.007203f
C3882 vdd.n2961 gnd 0.007203f
C3883 vdd.n2962 gnd 0.007203f
C3884 vdd.n2963 gnd 0.007203f
C3885 vdd.n2964 gnd 0.007203f
C3886 vdd.n2965 gnd 0.007203f
C3887 vdd.n2966 gnd 0.007203f
C3888 vdd.n2968 gnd 0.007203f
C3889 vdd.n2969 gnd 0.007203f
C3890 vdd.n2971 gnd 0.007203f
C3891 vdd.n2972 gnd 0.007203f
C3892 vdd.n2973 gnd 0.01709f
C3893 vdd.n2974 gnd 0.015957f
C3894 vdd.n2975 gnd 0.015957f
C3895 vdd.n2976 gnd 1.0608f
C3896 vdd.n2977 gnd 0.015957f
C3897 vdd.n2978 gnd 0.01709f
C3898 vdd.n2979 gnd 0.016213f
C3899 vdd.n2980 gnd 0.007203f
C3900 vdd.n2981 gnd 0.005561f
C3901 vdd.n2982 gnd 0.007203f
C3902 vdd.n2984 gnd 0.007203f
C3903 vdd.n2985 gnd 0.007203f
C3904 vdd.n2986 gnd 0.007203f
C3905 vdd.n2987 gnd 0.007203f
C3906 vdd.n2988 gnd 0.007203f
C3907 vdd.n2989 gnd 0.007203f
C3908 vdd.n2991 gnd 0.007203f
C3909 vdd.n2992 gnd 0.007203f
C3910 vdd.n2993 gnd 0.007203f
C3911 vdd.n2994 gnd 0.007203f
C3912 vdd.n2995 gnd 0.007203f
C3913 vdd.n2996 gnd 0.007203f
C3914 vdd.n2998 gnd 0.007203f
C3915 vdd.n2999 gnd 0.007203f
C3916 vdd.n3000 gnd 0.007203f
C3917 vdd.n3001 gnd 0.007203f
C3918 vdd.n3002 gnd 0.007203f
C3919 vdd.n3003 gnd 0.007203f
C3920 vdd.n3005 gnd 0.007203f
C3921 vdd.n3006 gnd 0.007203f
C3922 vdd.n3008 gnd 0.007203f
C3923 vdd.n3009 gnd 0.017308f
C3924 vdd.n3010 gnd 0.641044f
C3925 vdd.n3011 gnd 0.009109f
C3926 vdd.n3012 gnd 0.004049f
C3927 vdd.t71 gnd 0.130309f
C3928 vdd.t72 gnd 0.139265f
C3929 vdd.t70 gnd 0.170182f
C3930 vdd.n3013 gnd 0.218149f
C3931 vdd.n3014 gnd 0.183285f
C3932 vdd.n3015 gnd 0.013129f
C3933 vdd.n3016 gnd 0.010592f
C3934 vdd.n3017 gnd 0.004476f
C3935 vdd.n3018 gnd 0.008525f
C3936 vdd.n3019 gnd 0.010592f
C3937 vdd.n3020 gnd 0.010592f
C3938 vdd.n3021 gnd 0.008525f
C3939 vdd.n3022 gnd 0.008525f
C3940 vdd.n3023 gnd 0.010592f
C3941 vdd.n3025 gnd 0.010592f
C3942 vdd.n3026 gnd 0.008525f
C3943 vdd.n3027 gnd 0.008525f
C3944 vdd.n3028 gnd 0.008525f
C3945 vdd.n3029 gnd 0.010592f
C3946 vdd.n3031 gnd 0.010592f
C3947 vdd.n3033 gnd 0.010592f
C3948 vdd.n3034 gnd 0.008525f
C3949 vdd.n3035 gnd 0.008525f
C3950 vdd.n3036 gnd 0.008525f
C3951 vdd.n3037 gnd 0.010592f
C3952 vdd.n3039 gnd 0.010592f
C3953 vdd.n3041 gnd 0.010592f
C3954 vdd.n3042 gnd 0.008525f
C3955 vdd.n3043 gnd 0.008525f
C3956 vdd.n3044 gnd 0.008525f
C3957 vdd.n3045 gnd 0.010592f
C3958 vdd.n3047 gnd 0.010592f
C3959 vdd.n3048 gnd 0.010592f
C3960 vdd.n3049 gnd 0.008525f
C3961 vdd.n3050 gnd 0.008525f
C3962 vdd.n3051 gnd 0.010592f
C3963 vdd.n3052 gnd 0.010592f
C3964 vdd.n3054 gnd 0.010592f
C3965 vdd.n3055 gnd 0.008525f
C3966 vdd.n3056 gnd 0.010592f
C3967 vdd.n3057 gnd 0.010592f
C3968 vdd.n3058 gnd 0.010592f
C3969 vdd.n3059 gnd 0.017392f
C3970 vdd.n3060 gnd 0.005797f
C3971 vdd.n3061 gnd 0.010592f
C3972 vdd.n3063 gnd 0.010592f
C3973 vdd.n3065 gnd 0.010592f
C3974 vdd.n3066 gnd 0.008525f
C3975 vdd.n3067 gnd 0.008525f
C3976 vdd.n3068 gnd 0.008525f
C3977 vdd.n3069 gnd 0.010592f
C3978 vdd.n3071 gnd 0.010592f
C3979 vdd.n3073 gnd 0.010592f
C3980 vdd.n3074 gnd 0.008525f
C3981 vdd.n3075 gnd 0.008525f
C3982 vdd.n3076 gnd 0.008525f
C3983 vdd.n3077 gnd 0.010592f
C3984 vdd.n3079 gnd 0.010592f
C3985 vdd.n3081 gnd 0.010592f
C3986 vdd.n3082 gnd 0.008525f
C3987 vdd.n3083 gnd 0.008525f
C3988 vdd.n3084 gnd 0.008525f
C3989 vdd.n3085 gnd 0.010592f
C3990 vdd.n3087 gnd 0.010592f
C3991 vdd.n3089 gnd 0.010592f
C3992 vdd.n3090 gnd 0.008525f
C3993 vdd.n3091 gnd 0.008525f
C3994 vdd.n3092 gnd 0.008525f
C3995 vdd.n3093 gnd 0.010592f
C3996 vdd.n3095 gnd 0.010592f
C3997 vdd.n3097 gnd 0.010592f
C3998 vdd.n3098 gnd 0.008525f
C3999 vdd.n3099 gnd 0.008525f
C4000 vdd.n3100 gnd 0.007119f
C4001 vdd.n3101 gnd 0.010592f
C4002 vdd.n3103 gnd 0.010592f
C4003 vdd.n3105 gnd 0.010592f
C4004 vdd.n3106 gnd 0.007119f
C4005 vdd.n3107 gnd 0.008525f
C4006 vdd.n3108 gnd 0.008525f
C4007 vdd.n3109 gnd 0.010592f
C4008 vdd.n3111 gnd 0.010592f
C4009 vdd.n3113 gnd 0.010592f
C4010 vdd.n3114 gnd 0.008525f
C4011 vdd.n3115 gnd 0.008525f
C4012 vdd.n3116 gnd 0.008525f
C4013 vdd.n3117 gnd 0.010592f
C4014 vdd.n3119 gnd 0.010592f
C4015 vdd.n3121 gnd 0.010592f
C4016 vdd.n3122 gnd 0.008525f
C4017 vdd.n3123 gnd 0.008525f
C4018 vdd.n3124 gnd 0.008525f
C4019 vdd.n3125 gnd 0.010592f
C4020 vdd.n3127 gnd 0.010592f
C4021 vdd.n3128 gnd 0.010592f
C4022 vdd.n3129 gnd 0.008525f
C4023 vdd.n3130 gnd 0.008525f
C4024 vdd.n3131 gnd 0.010592f
C4025 vdd.n3132 gnd 0.010592f
C4026 vdd.n3133 gnd 0.008525f
C4027 vdd.n3134 gnd 0.008525f
C4028 vdd.n3135 gnd 0.010592f
C4029 vdd.n3136 gnd 0.010592f
C4030 vdd.n3138 gnd 0.010592f
C4031 vdd.n3139 gnd 0.008525f
C4032 vdd.n3140 gnd 0.007076f
C4033 vdd.n3141 gnd 0.024285f
C4034 vdd.n3142 gnd 0.02412f
C4035 vdd.n3143 gnd 0.007076f
C4036 vdd.n3144 gnd 0.02412f
C4037 vdd.n3145 gnd 1.42883f
C4038 vdd.n3146 gnd 0.02412f
C4039 vdd.n3147 gnd 0.007076f
C4040 vdd.n3148 gnd 0.02412f
C4041 vdd.n3149 gnd 0.010592f
C4042 vdd.n3150 gnd 0.010592f
C4043 vdd.n3151 gnd 0.008525f
C4044 vdd.n3152 gnd 0.010592f
C4045 vdd.n3153 gnd 1.02291f
C4046 vdd.n3154 gnd 0.010592f
C4047 vdd.n3155 gnd 0.008525f
C4048 vdd.n3156 gnd 0.010592f
C4049 vdd.n3157 gnd 0.010592f
C4050 vdd.n3158 gnd 0.010592f
C4051 vdd.n3159 gnd 0.008525f
C4052 vdd.n3160 gnd 0.010592f
C4053 vdd.n3161 gnd 1.05539f
C4054 vdd.n3162 gnd 0.010592f
C4055 vdd.n3163 gnd 0.008525f
C4056 vdd.n3164 gnd 0.010592f
C4057 vdd.n3165 gnd 0.010592f
C4058 vdd.n3166 gnd 0.010592f
C4059 vdd.n3167 gnd 0.008525f
C4060 vdd.n3168 gnd 0.010592f
C4061 vdd.t180 gnd 0.541225f
C4062 vdd.n3169 gnd 0.871372f
C4063 vdd.n3170 gnd 0.010592f
C4064 vdd.n3171 gnd 0.008525f
C4065 vdd.n3172 gnd 0.010592f
C4066 vdd.n3173 gnd 0.010592f
C4067 vdd.n3174 gnd 0.010592f
C4068 vdd.n3175 gnd 0.008525f
C4069 vdd.n3176 gnd 0.010592f
C4070 vdd.n3177 gnd 0.687355f
C4071 vdd.n3178 gnd 0.010592f
C4072 vdd.n3179 gnd 0.008525f
C4073 vdd.n3180 gnd 0.010592f
C4074 vdd.n3181 gnd 0.010592f
C4075 vdd.n3182 gnd 0.010592f
C4076 vdd.n3183 gnd 0.008525f
C4077 vdd.n3184 gnd 0.010592f
C4078 vdd.n3185 gnd 0.860547f
C4079 vdd.n3186 gnd 0.57911f
C4080 vdd.n3187 gnd 0.010592f
C4081 vdd.n3188 gnd 0.008525f
C4082 vdd.n3189 gnd 0.010592f
C4083 vdd.n3190 gnd 0.010592f
C4084 vdd.n3191 gnd 0.010592f
C4085 vdd.n3192 gnd 0.008525f
C4086 vdd.n3193 gnd 0.010592f
C4087 vdd.n3194 gnd 0.763127f
C4088 vdd.n3195 gnd 0.010592f
C4089 vdd.n3196 gnd 0.008525f
C4090 vdd.n3197 gnd 0.010592f
C4091 vdd.n3198 gnd 0.010592f
C4092 vdd.n3199 gnd 0.010592f
C4093 vdd.n3200 gnd 0.010592f
C4094 vdd.n3201 gnd 0.010592f
C4095 vdd.n3202 gnd 0.008525f
C4096 vdd.n3203 gnd 0.008525f
C4097 vdd.n3204 gnd 0.010592f
C4098 vdd.t110 gnd 0.541225f
C4099 vdd.n3205 gnd 0.898433f
C4100 vdd.n3206 gnd 0.010592f
C4101 vdd.n3207 gnd 0.008525f
C4102 vdd.n3208 gnd 0.010592f
C4103 vdd.n3209 gnd 0.010592f
C4104 vdd.n3210 gnd 0.010592f
C4105 vdd.n3211 gnd 0.008525f
C4106 vdd.n3212 gnd 0.010592f
C4107 vdd.n3213 gnd 0.849723f
C4108 vdd.n3214 gnd 0.010592f
C4109 vdd.n3215 gnd 0.010592f
C4110 vdd.n3216 gnd 0.008525f
C4111 vdd.n3217 gnd 0.008525f
C4112 vdd.n3218 gnd 0.008525f
C4113 vdd.n3219 gnd 0.010592f
C4114 vdd.n3220 gnd 0.010592f
C4115 vdd.n3221 gnd 0.010592f
C4116 vdd.n3222 gnd 0.010592f
C4117 vdd.n3223 gnd 0.008525f
C4118 vdd.n3224 gnd 0.008525f
C4119 vdd.n3225 gnd 0.008525f
C4120 vdd.n3226 gnd 0.010592f
C4121 vdd.n3227 gnd 0.010592f
C4122 vdd.n3228 gnd 0.010592f
C4123 vdd.n3229 gnd 0.010592f
C4124 vdd.n3230 gnd 0.008525f
C4125 vdd.n3231 gnd 0.008525f
C4126 vdd.n3232 gnd 0.008525f
C4127 vdd.n3233 gnd 0.010592f
C4128 vdd.n3234 gnd 0.010592f
C4129 vdd.n3235 gnd 0.010592f
C4130 vdd.n3236 gnd 0.898433f
C4131 vdd.n3237 gnd 0.010592f
C4132 vdd.n3238 gnd 0.008525f
C4133 vdd.n3239 gnd 0.008525f
C4134 vdd.n3240 gnd 0.008525f
C4135 vdd.n3241 gnd 0.010592f
C4136 vdd.n3242 gnd 0.010592f
C4137 vdd.n3243 gnd 0.010592f
C4138 vdd.n3244 gnd 0.010592f
C4139 vdd.n3245 gnd 0.008525f
C4140 vdd.n3246 gnd 0.008525f
C4141 vdd.n3247 gnd 0.007076f
C4142 vdd.n3248 gnd 0.02412f
C4143 vdd.n3249 gnd 0.024285f
C4144 vdd.n3250 gnd 0.004049f
C4145 vdd.n3251 gnd 0.024285f
C4146 vdd.n3253 gnd 2.39221f
C4147 vdd.n3254 gnd 1.42883f
C4148 vdd.n3255 gnd 0.709004f
C4149 vdd.n3256 gnd 0.010592f
C4150 vdd.n3257 gnd 0.008525f
C4151 vdd.n3258 gnd 0.008525f
C4152 vdd.n3259 gnd 0.008525f
C4153 vdd.n3260 gnd 0.010592f
C4154 vdd.n3261 gnd 1.08245f
C4155 vdd.n3262 gnd 1.08245f
C4156 vdd.n3263 gnd 0.622408f
C4157 vdd.n3264 gnd 0.010592f
C4158 vdd.n3265 gnd 0.008525f
C4159 vdd.n3266 gnd 0.008525f
C4160 vdd.n3267 gnd 0.008525f
C4161 vdd.n3268 gnd 0.010592f
C4162 vdd.n3269 gnd 0.644057f
C4163 vdd.n3270 gnd 0.7956f
C4164 vdd.t153 gnd 0.541225f
C4165 vdd.n3271 gnd 0.828074f
C4166 vdd.n3272 gnd 0.010592f
C4167 vdd.n3273 gnd 0.008525f
C4168 vdd.n3274 gnd 0.008525f
C4169 vdd.n3275 gnd 0.008525f
C4170 vdd.n3276 gnd 0.010592f
C4171 vdd.n3277 gnd 0.898433f
C4172 vdd.t130 gnd 0.541225f
C4173 vdd.n3278 gnd 0.654882f
C4174 vdd.n3279 gnd 0.784776f
C4175 vdd.n3280 gnd 0.010592f
C4176 vdd.n3281 gnd 0.008525f
C4177 vdd.n3282 gnd 0.008525f
C4178 vdd.n3283 gnd 0.008525f
C4179 vdd.n3284 gnd 0.010592f
C4180 vdd.n3285 gnd 0.600759f
C4181 vdd.t120 gnd 0.541225f
C4182 vdd.n3286 gnd 0.898433f
C4183 vdd.t157 gnd 0.541225f
C4184 vdd.n3287 gnd 0.665706f
C4185 vdd.n3288 gnd 0.010592f
C4186 vdd.n3289 gnd 0.008525f
C4187 vdd.n3290 gnd 0.008141f
C4188 vdd.n3291 gnd 0.624755f
C4189 vdd.n3292 gnd 2.5217f
C4190 a_n6972_8799.n0 gnd 2.71557f
C4191 a_n6972_8799.n1 gnd 1.6453f
C4192 a_n6972_8799.n2 gnd 3.76426f
C4193 a_n6972_8799.n3 gnd 0.205303f
C4194 a_n6972_8799.n4 gnd 0.28695f
C4195 a_n6972_8799.n5 gnd 0.205303f
C4196 a_n6972_8799.n6 gnd 0.205303f
C4197 a_n6972_8799.n7 gnd 0.205303f
C4198 a_n6972_8799.n8 gnd 0.270477f
C4199 a_n6972_8799.n9 gnd 0.205303f
C4200 a_n6972_8799.n10 gnd 0.28695f
C4201 a_n6972_8799.n11 gnd 0.205303f
C4202 a_n6972_8799.n12 gnd 0.205303f
C4203 a_n6972_8799.n13 gnd 0.205303f
C4204 a_n6972_8799.n14 gnd 0.270477f
C4205 a_n6972_8799.n15 gnd 0.205303f
C4206 a_n6972_8799.n16 gnd 0.449706f
C4207 a_n6972_8799.n17 gnd 0.205303f
C4208 a_n6972_8799.n18 gnd 0.205303f
C4209 a_n6972_8799.n19 gnd 0.205303f
C4210 a_n6972_8799.n20 gnd 0.270477f
C4211 a_n6972_8799.n21 gnd 0.321803f
C4212 a_n6972_8799.n22 gnd 0.205303f
C4213 a_n6972_8799.n23 gnd 0.205303f
C4214 a_n6972_8799.n24 gnd 0.205303f
C4215 a_n6972_8799.n25 gnd 0.205303f
C4216 a_n6972_8799.n26 gnd 0.235624f
C4217 a_n6972_8799.n27 gnd 0.321803f
C4218 a_n6972_8799.n28 gnd 0.205303f
C4219 a_n6972_8799.n29 gnd 0.205303f
C4220 a_n6972_8799.n30 gnd 0.205303f
C4221 a_n6972_8799.n31 gnd 0.205303f
C4222 a_n6972_8799.n32 gnd 0.235624f
C4223 a_n6972_8799.n33 gnd 0.321803f
C4224 a_n6972_8799.n34 gnd 0.205303f
C4225 a_n6972_8799.n35 gnd 0.205303f
C4226 a_n6972_8799.n36 gnd 0.205303f
C4227 a_n6972_8799.n37 gnd 0.205303f
C4228 a_n6972_8799.n38 gnd 0.39838f
C4229 a_n6972_8799.n39 gnd 2.80287f
C4230 a_n6972_8799.n40 gnd 3.91963f
C4231 a_n6972_8799.n41 gnd 0.008515f
C4232 a_n6972_8799.n42 gnd 0.001143f
C4233 a_n6972_8799.n44 gnd 0.007647f
C4234 a_n6972_8799.n45 gnd 0.011558f
C4235 a_n6972_8799.n46 gnd 0.007949f
C4236 a_n6972_8799.n48 gnd 3.97e-19
C4237 a_n6972_8799.n49 gnd 0.008238f
C4238 a_n6972_8799.n50 gnd 0.011378f
C4239 a_n6972_8799.n51 gnd 0.007331f
C4240 a_n6972_8799.n52 gnd 0.008515f
C4241 a_n6972_8799.n53 gnd 0.001143f
C4242 a_n6972_8799.n55 gnd 0.007647f
C4243 a_n6972_8799.n56 gnd 0.011558f
C4244 a_n6972_8799.n57 gnd 0.007949f
C4245 a_n6972_8799.n59 gnd 3.97e-19
C4246 a_n6972_8799.n60 gnd 0.008238f
C4247 a_n6972_8799.n61 gnd 0.011378f
C4248 a_n6972_8799.n62 gnd 0.007331f
C4249 a_n6972_8799.n63 gnd 0.008515f
C4250 a_n6972_8799.n64 gnd 0.001143f
C4251 a_n6972_8799.n66 gnd 0.007647f
C4252 a_n6972_8799.n67 gnd 0.011558f
C4253 a_n6972_8799.n68 gnd 0.007949f
C4254 a_n6972_8799.n70 gnd 3.97e-19
C4255 a_n6972_8799.n71 gnd 0.008238f
C4256 a_n6972_8799.n72 gnd 0.011378f
C4257 a_n6972_8799.n73 gnd 0.007331f
C4258 a_n6972_8799.n74 gnd 0.001143f
C4259 a_n6972_8799.n76 gnd 0.007647f
C4260 a_n6972_8799.n77 gnd 0.011558f
C4261 a_n6972_8799.n78 gnd 0.007949f
C4262 a_n6972_8799.n80 gnd 3.97e-19
C4263 a_n6972_8799.n81 gnd 0.008238f
C4264 a_n6972_8799.n82 gnd 0.011378f
C4265 a_n6972_8799.n83 gnd 0.007331f
C4266 a_n6972_8799.n84 gnd 0.247165f
C4267 a_n6972_8799.n85 gnd 0.001143f
C4268 a_n6972_8799.n87 gnd 0.007647f
C4269 a_n6972_8799.n88 gnd 0.011558f
C4270 a_n6972_8799.n89 gnd 0.007949f
C4271 a_n6972_8799.n91 gnd 3.97e-19
C4272 a_n6972_8799.n92 gnd 0.008238f
C4273 a_n6972_8799.n93 gnd 0.011378f
C4274 a_n6972_8799.n94 gnd 0.007331f
C4275 a_n6972_8799.n95 gnd 0.247165f
C4276 a_n6972_8799.n96 gnd 0.001143f
C4277 a_n6972_8799.n98 gnd 0.007647f
C4278 a_n6972_8799.n99 gnd 0.011558f
C4279 a_n6972_8799.n100 gnd 0.007949f
C4280 a_n6972_8799.n102 gnd 3.97e-19
C4281 a_n6972_8799.n103 gnd 0.008238f
C4282 a_n6972_8799.n104 gnd 0.011378f
C4283 a_n6972_8799.n105 gnd 0.007331f
C4284 a_n6972_8799.n106 gnd 0.247165f
C4285 a_n6972_8799.t26 gnd 0.1424f
C4286 a_n6972_8799.t5 gnd 0.1424f
C4287 a_n6972_8799.t25 gnd 0.1424f
C4288 a_n6972_8799.n107 gnd 1.12313f
C4289 a_n6972_8799.t22 gnd 0.1424f
C4290 a_n6972_8799.t27 gnd 0.1424f
C4291 a_n6972_8799.n108 gnd 1.12128f
C4292 a_n6972_8799.t24 gnd 0.1424f
C4293 a_n6972_8799.t16 gnd 0.1424f
C4294 a_n6972_8799.n109 gnd 1.12128f
C4295 a_n6972_8799.t15 gnd 0.110756f
C4296 a_n6972_8799.t6 gnd 0.110756f
C4297 a_n6972_8799.n110 gnd 0.981561f
C4298 a_n6972_8799.t8 gnd 0.110756f
C4299 a_n6972_8799.t10 gnd 0.110756f
C4300 a_n6972_8799.n111 gnd 0.978675f
C4301 a_n6972_8799.t13 gnd 0.110756f
C4302 a_n6972_8799.t0 gnd 0.110756f
C4303 a_n6972_8799.n112 gnd 0.981561f
C4304 a_n6972_8799.t19 gnd 0.110756f
C4305 a_n6972_8799.t14 gnd 0.110756f
C4306 a_n6972_8799.n113 gnd 0.978675f
C4307 a_n6972_8799.t9 gnd 0.110756f
C4308 a_n6972_8799.t17 gnd 0.110756f
C4309 a_n6972_8799.n114 gnd 0.981561f
C4310 a_n6972_8799.t18 gnd 0.110756f
C4311 a_n6972_8799.t11 gnd 0.110756f
C4312 a_n6972_8799.n115 gnd 0.978675f
C4313 a_n6972_8799.t4 gnd 0.110756f
C4314 a_n6972_8799.t7 gnd 0.110756f
C4315 a_n6972_8799.n116 gnd 0.978675f
C4316 a_n6972_8799.t12 gnd 0.110756f
C4317 a_n6972_8799.t1 gnd 0.110756f
C4318 a_n6972_8799.n117 gnd 0.978675f
C4319 a_n6972_8799.t105 gnd 0.590457f
C4320 a_n6972_8799.n118 gnd 0.263979f
C4321 a_n6972_8799.t39 gnd 0.590457f
C4322 a_n6972_8799.t57 gnd 0.590457f
C4323 a_n6972_8799.n119 gnd 0.267249f
C4324 a_n6972_8799.t74 gnd 0.590457f
C4325 a_n6972_8799.t91 gnd 0.590457f
C4326 a_n6972_8799.t92 gnd 0.590457f
C4327 a_n6972_8799.n120 gnd 0.269308f
C4328 a_n6972_8799.t59 gnd 0.590457f
C4329 a_n6972_8799.t68 gnd 0.590457f
C4330 a_n6972_8799.n121 gnd 0.262918f
C4331 a_n6972_8799.t106 gnd 0.601632f
C4332 a_n6972_8799.n122 gnd 0.247545f
C4333 a_n6972_8799.n123 gnd 0.011647f
C4334 a_n6972_8799.t69 gnd 0.590457f
C4335 a_n6972_8799.n124 gnd 0.263709f
C4336 a_n6972_8799.n125 gnd 0.267235f
C4337 a_n6972_8799.t60 gnd 0.590457f
C4338 a_n6972_8799.n126 gnd 0.263798f
C4339 a_n6972_8799.n127 gnd 0.258488f
C4340 a_n6972_8799.t28 gnd 0.590457f
C4341 a_n6972_8799.n128 gnd 0.263551f
C4342 a_n6972_8799.n129 gnd 0.269738f
C4343 a_n6972_8799.t108 gnd 0.590457f
C4344 a_n6972_8799.n130 gnd 0.267118f
C4345 a_n6972_8799.n131 gnd 0.263235f
C4346 a_n6972_8799.t55 gnd 0.590457f
C4347 a_n6972_8799.n132 gnd 0.258804f
C4348 a_n6972_8799.t36 gnd 0.590457f
C4349 a_n6972_8799.n133 gnd 0.267234f
C4350 a_n6972_8799.t37 gnd 0.601622f
C4351 a_n6972_8799.t115 gnd 0.590457f
C4352 a_n6972_8799.n134 gnd 0.263979f
C4353 a_n6972_8799.t53 gnd 0.590457f
C4354 a_n6972_8799.t65 gnd 0.590457f
C4355 a_n6972_8799.n135 gnd 0.267249f
C4356 a_n6972_8799.t85 gnd 0.590457f
C4357 a_n6972_8799.t100 gnd 0.590457f
C4358 a_n6972_8799.t104 gnd 0.590457f
C4359 a_n6972_8799.n136 gnd 0.269308f
C4360 a_n6972_8799.t66 gnd 0.590457f
C4361 a_n6972_8799.t75 gnd 0.590457f
C4362 a_n6972_8799.n137 gnd 0.262918f
C4363 a_n6972_8799.t117 gnd 0.601632f
C4364 a_n6972_8799.n138 gnd 0.247545f
C4365 a_n6972_8799.n139 gnd 0.011647f
C4366 a_n6972_8799.t76 gnd 0.590457f
C4367 a_n6972_8799.n140 gnd 0.263709f
C4368 a_n6972_8799.n141 gnd 0.267235f
C4369 a_n6972_8799.t67 gnd 0.590457f
C4370 a_n6972_8799.n142 gnd 0.263798f
C4371 a_n6972_8799.n143 gnd 0.258488f
C4372 a_n6972_8799.t38 gnd 0.590457f
C4373 a_n6972_8799.n144 gnd 0.263551f
C4374 a_n6972_8799.n145 gnd 0.269738f
C4375 a_n6972_8799.t120 gnd 0.590457f
C4376 a_n6972_8799.n146 gnd 0.267118f
C4377 a_n6972_8799.n147 gnd 0.263235f
C4378 a_n6972_8799.t64 gnd 0.590457f
C4379 a_n6972_8799.n148 gnd 0.258804f
C4380 a_n6972_8799.t47 gnd 0.590457f
C4381 a_n6972_8799.n149 gnd 0.267234f
C4382 a_n6972_8799.t49 gnd 0.601622f
C4383 a_n6972_8799.n150 gnd 0.889294f
C4384 a_n6972_8799.t81 gnd 0.590457f
C4385 a_n6972_8799.n151 gnd 0.263979f
C4386 a_n6972_8799.t101 gnd 0.590457f
C4387 a_n6972_8799.t34 gnd 0.590457f
C4388 a_n6972_8799.n152 gnd 0.267249f
C4389 a_n6972_8799.t87 gnd 0.590457f
C4390 a_n6972_8799.t116 gnd 0.590457f
C4391 a_n6972_8799.t79 gnd 0.590457f
C4392 a_n6972_8799.n153 gnd 0.269308f
C4393 a_n6972_8799.t112 gnd 0.590457f
C4394 a_n6972_8799.t45 gnd 0.590457f
C4395 a_n6972_8799.n154 gnd 0.262918f
C4396 a_n6972_8799.t109 gnd 0.601632f
C4397 a_n6972_8799.n155 gnd 0.247545f
C4398 a_n6972_8799.n156 gnd 0.011647f
C4399 a_n6972_8799.t29 gnd 0.590457f
C4400 a_n6972_8799.n157 gnd 0.263709f
C4401 a_n6972_8799.n158 gnd 0.267235f
C4402 a_n6972_8799.t93 gnd 0.590457f
C4403 a_n6972_8799.n159 gnd 0.263798f
C4404 a_n6972_8799.n160 gnd 0.258488f
C4405 a_n6972_8799.t73 gnd 0.590457f
C4406 a_n6972_8799.n161 gnd 0.263551f
C4407 a_n6972_8799.n162 gnd 0.269738f
C4408 a_n6972_8799.t51 gnd 0.590457f
C4409 a_n6972_8799.n163 gnd 0.267118f
C4410 a_n6972_8799.n164 gnd 0.263235f
C4411 a_n6972_8799.t58 gnd 0.590457f
C4412 a_n6972_8799.n165 gnd 0.258804f
C4413 a_n6972_8799.t41 gnd 0.590457f
C4414 a_n6972_8799.n166 gnd 0.267234f
C4415 a_n6972_8799.t121 gnd 0.601622f
C4416 a_n6972_8799.n167 gnd 1.43412f
C4417 a_n6972_8799.t71 gnd 0.590457f
C4418 a_n6972_8799.t70 gnd 0.590457f
C4419 a_n6972_8799.t48 gnd 0.590457f
C4420 a_n6972_8799.n168 gnd 0.266841f
C4421 a_n6972_8799.t107 gnd 0.590457f
C4422 a_n6972_8799.t72 gnd 0.590457f
C4423 a_n6972_8799.t54 gnd 0.590457f
C4424 a_n6972_8799.n169 gnd 0.263798f
C4425 a_n6972_8799.t111 gnd 0.590457f
C4426 a_n6972_8799.t86 gnd 0.590457f
C4427 a_n6972_8799.t84 gnd 0.590457f
C4428 a_n6972_8799.n170 gnd 0.267249f
C4429 a_n6972_8799.t31 gnd 0.590457f
C4430 a_n6972_8799.t90 gnd 0.590457f
C4431 a_n6972_8799.t89 gnd 0.590457f
C4432 a_n6972_8799.n171 gnd 0.263235f
C4433 a_n6972_8799.t33 gnd 0.590457f
C4434 a_n6972_8799.t32 gnd 0.590457f
C4435 a_n6972_8799.t103 gnd 0.590457f
C4436 a_n6972_8799.n172 gnd 0.267234f
C4437 a_n6972_8799.t50 gnd 0.601632f
C4438 a_n6972_8799.n173 gnd 0.247545f
C4439 a_n6972_8799.n174 gnd 0.263979f
C4440 a_n6972_8799.n175 gnd 0.258804f
C4441 a_n6972_8799.n176 gnd 0.267118f
C4442 a_n6972_8799.n177 gnd 0.269738f
C4443 a_n6972_8799.n178 gnd 0.263551f
C4444 a_n6972_8799.n179 gnd 0.258488f
C4445 a_n6972_8799.n180 gnd 0.267235f
C4446 a_n6972_8799.n181 gnd 0.269308f
C4447 a_n6972_8799.n182 gnd 0.262918f
C4448 a_n6972_8799.n183 gnd 0.25833f
C4449 a_n6972_8799.t78 gnd 0.590457f
C4450 a_n6972_8799.t77 gnd 0.590457f
C4451 a_n6972_8799.t61 gnd 0.590457f
C4452 a_n6972_8799.n184 gnd 0.266841f
C4453 a_n6972_8799.t119 gnd 0.590457f
C4454 a_n6972_8799.t83 gnd 0.590457f
C4455 a_n6972_8799.t63 gnd 0.590457f
C4456 a_n6972_8799.n185 gnd 0.263798f
C4457 a_n6972_8799.t123 gnd 0.590457f
C4458 a_n6972_8799.t96 gnd 0.590457f
C4459 a_n6972_8799.t95 gnd 0.590457f
C4460 a_n6972_8799.n186 gnd 0.267249f
C4461 a_n6972_8799.t40 gnd 0.590457f
C4462 a_n6972_8799.t99 gnd 0.590457f
C4463 a_n6972_8799.t98 gnd 0.590457f
C4464 a_n6972_8799.n187 gnd 0.263235f
C4465 a_n6972_8799.t44 gnd 0.590457f
C4466 a_n6972_8799.t43 gnd 0.590457f
C4467 a_n6972_8799.t114 gnd 0.590457f
C4468 a_n6972_8799.n188 gnd 0.267234f
C4469 a_n6972_8799.t62 gnd 0.601632f
C4470 a_n6972_8799.n189 gnd 0.247545f
C4471 a_n6972_8799.n190 gnd 0.263979f
C4472 a_n6972_8799.n191 gnd 0.258804f
C4473 a_n6972_8799.n192 gnd 0.267118f
C4474 a_n6972_8799.n193 gnd 0.269738f
C4475 a_n6972_8799.n194 gnd 0.263551f
C4476 a_n6972_8799.n195 gnd 0.258488f
C4477 a_n6972_8799.n196 gnd 0.267235f
C4478 a_n6972_8799.n197 gnd 0.269308f
C4479 a_n6972_8799.n198 gnd 0.262918f
C4480 a_n6972_8799.n199 gnd 0.25833f
C4481 a_n6972_8799.n200 gnd 0.889294f
C4482 a_n6972_8799.t122 gnd 0.590457f
C4483 a_n6972_8799.t42 gnd 0.590457f
C4484 a_n6972_8799.t82 gnd 0.590457f
C4485 a_n6972_8799.n201 gnd 0.266841f
C4486 a_n6972_8799.t30 gnd 0.590457f
C4487 a_n6972_8799.t102 gnd 0.590457f
C4488 a_n6972_8799.t52 gnd 0.590457f
C4489 a_n6972_8799.n202 gnd 0.263798f
C4490 a_n6972_8799.t88 gnd 0.590457f
C4491 a_n6972_8799.t35 gnd 0.590457f
C4492 a_n6972_8799.t56 gnd 0.590457f
C4493 a_n6972_8799.n203 gnd 0.267249f
C4494 a_n6972_8799.t118 gnd 0.590457f
C4495 a_n6972_8799.t94 gnd 0.590457f
C4496 a_n6972_8799.t113 gnd 0.590457f
C4497 a_n6972_8799.n204 gnd 0.263235f
C4498 a_n6972_8799.t80 gnd 0.590457f
C4499 a_n6972_8799.t97 gnd 0.590457f
C4500 a_n6972_8799.t46 gnd 0.590457f
C4501 a_n6972_8799.n205 gnd 0.267234f
C4502 a_n6972_8799.t110 gnd 0.601632f
C4503 a_n6972_8799.n206 gnd 0.247545f
C4504 a_n6972_8799.n207 gnd 0.263979f
C4505 a_n6972_8799.n208 gnd 0.258804f
C4506 a_n6972_8799.n209 gnd 0.267118f
C4507 a_n6972_8799.n210 gnd 0.269738f
C4508 a_n6972_8799.n211 gnd 0.263551f
C4509 a_n6972_8799.n212 gnd 0.258488f
C4510 a_n6972_8799.n213 gnd 0.267235f
C4511 a_n6972_8799.n214 gnd 0.269308f
C4512 a_n6972_8799.n215 gnd 0.262918f
C4513 a_n6972_8799.n216 gnd 0.25833f
C4514 a_n6972_8799.n217 gnd 1.12457f
C4515 a_n6972_8799.n218 gnd 12.0955f
C4516 a_n6972_8799.n219 gnd 4.32129f
C4517 a_n6972_8799.n220 gnd 5.6226f
C4518 a_n6972_8799.t20 gnd 0.1424f
C4519 a_n6972_8799.t21 gnd 0.1424f
C4520 a_n6972_8799.n221 gnd 1.12128f
C4521 a_n6972_8799.t23 gnd 0.1424f
C4522 a_n6972_8799.t3 gnd 0.1424f
C4523 a_n6972_8799.n222 gnd 1.12313f
C4524 a_n6972_8799.n223 gnd 1.12128f
C4525 a_n6972_8799.t2 gnd 0.1424f
C4526 CSoutput.n0 gnd 0.044795f
C4527 CSoutput.t194 gnd 0.296307f
C4528 CSoutput.n1 gnd 0.133797f
C4529 CSoutput.n2 gnd 0.044795f
C4530 CSoutput.t192 gnd 0.296307f
C4531 CSoutput.n3 gnd 0.035503f
C4532 CSoutput.n4 gnd 0.044795f
C4533 CSoutput.t185 gnd 0.296307f
C4534 CSoutput.n5 gnd 0.030615f
C4535 CSoutput.n6 gnd 0.044795f
C4536 CSoutput.t189 gnd 0.296307f
C4537 CSoutput.t178 gnd 0.296307f
C4538 CSoutput.n7 gnd 0.132339f
C4539 CSoutput.n8 gnd 0.044795f
C4540 CSoutput.t177 gnd 0.296307f
C4541 CSoutput.n9 gnd 0.02919f
C4542 CSoutput.n10 gnd 0.044795f
C4543 CSoutput.t186 gnd 0.296307f
C4544 CSoutput.t191 gnd 0.296307f
C4545 CSoutput.n11 gnd 0.132339f
C4546 CSoutput.n12 gnd 0.044795f
C4547 CSoutput.t197 gnd 0.296307f
C4548 CSoutput.n13 gnd 0.030615f
C4549 CSoutput.n14 gnd 0.044795f
C4550 CSoutput.t179 gnd 0.296307f
C4551 CSoutput.t188 gnd 0.296307f
C4552 CSoutput.n15 gnd 0.132339f
C4553 CSoutput.n16 gnd 0.044795f
C4554 CSoutput.t195 gnd 0.296307f
C4555 CSoutput.n17 gnd 0.032698f
C4556 CSoutput.t182 gnd 0.354094f
C4557 CSoutput.t193 gnd 0.296307f
C4558 CSoutput.n18 gnd 0.168946f
C4559 CSoutput.n19 gnd 0.163936f
C4560 CSoutput.n20 gnd 0.190185f
C4561 CSoutput.n21 gnd 0.044795f
C4562 CSoutput.n22 gnd 0.037386f
C4563 CSoutput.n23 gnd 0.132339f
C4564 CSoutput.n24 gnd 0.036039f
C4565 CSoutput.n25 gnd 0.035503f
C4566 CSoutput.n26 gnd 0.044795f
C4567 CSoutput.n27 gnd 0.044795f
C4568 CSoutput.n28 gnd 0.037099f
C4569 CSoutput.n29 gnd 0.031498f
C4570 CSoutput.n30 gnd 0.135285f
C4571 CSoutput.n31 gnd 0.031932f
C4572 CSoutput.n32 gnd 0.044795f
C4573 CSoutput.n33 gnd 0.044795f
C4574 CSoutput.n34 gnd 0.044795f
C4575 CSoutput.n35 gnd 0.036704f
C4576 CSoutput.n36 gnd 0.132339f
C4577 CSoutput.n37 gnd 0.035102f
C4578 CSoutput.n38 gnd 0.036441f
C4579 CSoutput.n39 gnd 0.044795f
C4580 CSoutput.n40 gnd 0.044795f
C4581 CSoutput.n41 gnd 0.037378f
C4582 CSoutput.n42 gnd 0.034164f
C4583 CSoutput.n43 gnd 0.132339f
C4584 CSoutput.n44 gnd 0.03503f
C4585 CSoutput.n45 gnd 0.044795f
C4586 CSoutput.n46 gnd 0.044795f
C4587 CSoutput.n47 gnd 0.044795f
C4588 CSoutput.n48 gnd 0.03503f
C4589 CSoutput.n49 gnd 0.132339f
C4590 CSoutput.n50 gnd 0.034164f
C4591 CSoutput.n51 gnd 0.037378f
C4592 CSoutput.n52 gnd 0.044795f
C4593 CSoutput.n53 gnd 0.044795f
C4594 CSoutput.n54 gnd 0.036441f
C4595 CSoutput.n55 gnd 0.035102f
C4596 CSoutput.n56 gnd 0.132339f
C4597 CSoutput.n57 gnd 0.036704f
C4598 CSoutput.n58 gnd 0.044795f
C4599 CSoutput.n59 gnd 0.044795f
C4600 CSoutput.n60 gnd 0.044795f
C4601 CSoutput.n61 gnd 0.031932f
C4602 CSoutput.n62 gnd 0.135285f
C4603 CSoutput.n63 gnd 0.031498f
C4604 CSoutput.t181 gnd 0.296307f
C4605 CSoutput.n64 gnd 0.132339f
C4606 CSoutput.n65 gnd 0.037099f
C4607 CSoutput.n66 gnd 0.044795f
C4608 CSoutput.n67 gnd 0.044795f
C4609 CSoutput.n68 gnd 0.044795f
C4610 CSoutput.n69 gnd 0.036039f
C4611 CSoutput.n70 gnd 0.132339f
C4612 CSoutput.n71 gnd 0.037386f
C4613 CSoutput.n72 gnd 0.032698f
C4614 CSoutput.n73 gnd 0.044795f
C4615 CSoutput.n74 gnd 0.044795f
C4616 CSoutput.n75 gnd 0.03391f
C4617 CSoutput.n76 gnd 0.020139f
C4618 CSoutput.t184 gnd 0.332922f
C4619 CSoutput.n77 gnd 0.165382f
C4620 CSoutput.n78 gnd 0.707655f
C4621 CSoutput.t167 gnd 0.055875f
C4622 CSoutput.t72 gnd 0.055875f
C4623 CSoutput.n79 gnd 0.432603f
C4624 CSoutput.t63 gnd 0.055875f
C4625 CSoutput.t14 gnd 0.055875f
C4626 CSoutput.n80 gnd 0.431831f
C4627 CSoutput.n81 gnd 0.438308f
C4628 CSoutput.t38 gnd 0.055875f
C4629 CSoutput.t61 gnd 0.055875f
C4630 CSoutput.n82 gnd 0.431831f
C4631 CSoutput.n83 gnd 0.21598f
C4632 CSoutput.t24 gnd 0.055875f
C4633 CSoutput.t21 gnd 0.055875f
C4634 CSoutput.n84 gnd 0.431831f
C4635 CSoutput.n85 gnd 0.21598f
C4636 CSoutput.t25 gnd 0.055875f
C4637 CSoutput.t73 gnd 0.055875f
C4638 CSoutput.n86 gnd 0.431831f
C4639 CSoutput.n87 gnd 0.21598f
C4640 CSoutput.t50 gnd 0.055875f
C4641 CSoutput.t58 gnd 0.055875f
C4642 CSoutput.n88 gnd 0.431831f
C4643 CSoutput.n89 gnd 0.21598f
C4644 CSoutput.t175 gnd 0.055875f
C4645 CSoutput.t2 gnd 0.055875f
C4646 CSoutput.n90 gnd 0.431831f
C4647 CSoutput.n91 gnd 0.21598f
C4648 CSoutput.t48 gnd 0.055875f
C4649 CSoutput.t71 gnd 0.055875f
C4650 CSoutput.n92 gnd 0.431831f
C4651 CSoutput.n93 gnd 0.396057f
C4652 CSoutput.t62 gnd 0.055875f
C4653 CSoutput.t18 gnd 0.055875f
C4654 CSoutput.n94 gnd 0.432603f
C4655 CSoutput.t29 gnd 0.055875f
C4656 CSoutput.t68 gnd 0.055875f
C4657 CSoutput.n95 gnd 0.431831f
C4658 CSoutput.n96 gnd 0.438308f
C4659 CSoutput.t34 gnd 0.055875f
C4660 CSoutput.t27 gnd 0.055875f
C4661 CSoutput.n97 gnd 0.431831f
C4662 CSoutput.n98 gnd 0.21598f
C4663 CSoutput.t8 gnd 0.055875f
C4664 CSoutput.t9 gnd 0.055875f
C4665 CSoutput.n99 gnd 0.431831f
C4666 CSoutput.n100 gnd 0.21598f
C4667 CSoutput.t11 gnd 0.055875f
C4668 CSoutput.t6 gnd 0.055875f
C4669 CSoutput.n101 gnd 0.431831f
C4670 CSoutput.n102 gnd 0.21598f
C4671 CSoutput.t65 gnd 0.055875f
C4672 CSoutput.t74 gnd 0.055875f
C4673 CSoutput.n103 gnd 0.431831f
C4674 CSoutput.n104 gnd 0.21598f
C4675 CSoutput.t46 gnd 0.055875f
C4676 CSoutput.t0 gnd 0.055875f
C4677 CSoutput.n105 gnd 0.431831f
C4678 CSoutput.n106 gnd 0.21598f
C4679 CSoutput.t164 gnd 0.055875f
C4680 CSoutput.t30 gnd 0.055875f
C4681 CSoutput.n107 gnd 0.431831f
C4682 CSoutput.n108 gnd 0.32208f
C4683 CSoutput.n109 gnd 0.406141f
C4684 CSoutput.t32 gnd 0.055875f
C4685 CSoutput.t33 gnd 0.055875f
C4686 CSoutput.n110 gnd 0.432603f
C4687 CSoutput.t31 gnd 0.055875f
C4688 CSoutput.t1 gnd 0.055875f
C4689 CSoutput.n111 gnd 0.431831f
C4690 CSoutput.n112 gnd 0.438308f
C4691 CSoutput.t16 gnd 0.055875f
C4692 CSoutput.t49 gnd 0.055875f
C4693 CSoutput.n113 gnd 0.431831f
C4694 CSoutput.n114 gnd 0.21598f
C4695 CSoutput.t40 gnd 0.055875f
C4696 CSoutput.t47 gnd 0.055875f
C4697 CSoutput.n115 gnd 0.431831f
C4698 CSoutput.n116 gnd 0.21598f
C4699 CSoutput.t172 gnd 0.055875f
C4700 CSoutput.t163 gnd 0.055875f
C4701 CSoutput.n117 gnd 0.431831f
C4702 CSoutput.n118 gnd 0.21598f
C4703 CSoutput.t17 gnd 0.055875f
C4704 CSoutput.t3 gnd 0.055875f
C4705 CSoutput.n119 gnd 0.431831f
C4706 CSoutput.n120 gnd 0.21598f
C4707 CSoutput.t168 gnd 0.055875f
C4708 CSoutput.t66 gnd 0.055875f
C4709 CSoutput.n121 gnd 0.431831f
C4710 CSoutput.n122 gnd 0.21598f
C4711 CSoutput.t166 gnd 0.055875f
C4712 CSoutput.t69 gnd 0.055875f
C4713 CSoutput.n123 gnd 0.431831f
C4714 CSoutput.n124 gnd 0.32208f
C4715 CSoutput.n125 gnd 0.453962f
C4716 CSoutput.n126 gnd 8.897231f
C4717 CSoutput.n128 gnd 0.792409f
C4718 CSoutput.n129 gnd 0.594307f
C4719 CSoutput.n130 gnd 0.792409f
C4720 CSoutput.n131 gnd 0.792409f
C4721 CSoutput.n132 gnd 2.13341f
C4722 CSoutput.n133 gnd 0.792409f
C4723 CSoutput.n134 gnd 0.792409f
C4724 CSoutput.t187 gnd 0.990511f
C4725 CSoutput.n135 gnd 0.792409f
C4726 CSoutput.n136 gnd 0.792409f
C4727 CSoutput.n140 gnd 0.792409f
C4728 CSoutput.n144 gnd 0.792409f
C4729 CSoutput.n145 gnd 0.792409f
C4730 CSoutput.n147 gnd 0.792409f
C4731 CSoutput.n152 gnd 0.792409f
C4732 CSoutput.n154 gnd 0.792409f
C4733 CSoutput.n155 gnd 0.792409f
C4734 CSoutput.n157 gnd 0.792409f
C4735 CSoutput.n158 gnd 0.792409f
C4736 CSoutput.n160 gnd 0.792409f
C4737 CSoutput.t180 gnd 13.241099f
C4738 CSoutput.n162 gnd 0.792409f
C4739 CSoutput.n163 gnd 0.594307f
C4740 CSoutput.n164 gnd 0.792409f
C4741 CSoutput.n165 gnd 0.792409f
C4742 CSoutput.n166 gnd 2.13341f
C4743 CSoutput.n167 gnd 0.792409f
C4744 CSoutput.n168 gnd 0.792409f
C4745 CSoutput.t196 gnd 0.990511f
C4746 CSoutput.n169 gnd 0.792409f
C4747 CSoutput.n170 gnd 0.792409f
C4748 CSoutput.n174 gnd 0.792409f
C4749 CSoutput.n178 gnd 0.792409f
C4750 CSoutput.n179 gnd 0.792409f
C4751 CSoutput.n181 gnd 0.792409f
C4752 CSoutput.n186 gnd 0.792409f
C4753 CSoutput.n188 gnd 0.792409f
C4754 CSoutput.n189 gnd 0.792409f
C4755 CSoutput.n191 gnd 0.792409f
C4756 CSoutput.n192 gnd 0.792409f
C4757 CSoutput.n194 gnd 0.792409f
C4758 CSoutput.n195 gnd 0.594307f
C4759 CSoutput.n197 gnd 0.792409f
C4760 CSoutput.n198 gnd 0.594307f
C4761 CSoutput.n199 gnd 0.792409f
C4762 CSoutput.n200 gnd 0.792409f
C4763 CSoutput.n201 gnd 2.13341f
C4764 CSoutput.n202 gnd 0.792409f
C4765 CSoutput.n203 gnd 0.792409f
C4766 CSoutput.t190 gnd 0.990511f
C4767 CSoutput.n204 gnd 0.792409f
C4768 CSoutput.n205 gnd 2.13341f
C4769 CSoutput.n207 gnd 0.792409f
C4770 CSoutput.n208 gnd 0.792409f
C4771 CSoutput.n210 gnd 0.792409f
C4772 CSoutput.n211 gnd 0.792409f
C4773 CSoutput.t176 gnd 13.0253f
C4774 CSoutput.t183 gnd 13.241099f
C4775 CSoutput.n217 gnd 2.4859f
C4776 CSoutput.n218 gnd 10.126699f
C4777 CSoutput.n219 gnd 10.5504f
C4778 CSoutput.n224 gnd 2.6929f
C4779 CSoutput.n230 gnd 0.792409f
C4780 CSoutput.n232 gnd 0.792409f
C4781 CSoutput.n234 gnd 0.792409f
C4782 CSoutput.n236 gnd 0.792409f
C4783 CSoutput.n238 gnd 0.792409f
C4784 CSoutput.n244 gnd 0.792409f
C4785 CSoutput.n251 gnd 1.45377f
C4786 CSoutput.n252 gnd 1.45377f
C4787 CSoutput.n253 gnd 0.792409f
C4788 CSoutput.n254 gnd 0.792409f
C4789 CSoutput.n256 gnd 0.594307f
C4790 CSoutput.n257 gnd 0.50897f
C4791 CSoutput.n259 gnd 0.594307f
C4792 CSoutput.n260 gnd 0.50897f
C4793 CSoutput.n261 gnd 0.594307f
C4794 CSoutput.n263 gnd 0.792409f
C4795 CSoutput.n265 gnd 2.13341f
C4796 CSoutput.n266 gnd 2.4859f
C4797 CSoutput.n267 gnd 9.31393f
C4798 CSoutput.n269 gnd 0.594307f
C4799 CSoutput.n270 gnd 1.52919f
C4800 CSoutput.n271 gnd 0.594307f
C4801 CSoutput.n273 gnd 0.792409f
C4802 CSoutput.n275 gnd 2.13341f
C4803 CSoutput.n276 gnd 4.64691f
C4804 CSoutput.t173 gnd 0.055875f
C4805 CSoutput.t20 gnd 0.055875f
C4806 CSoutput.n277 gnd 0.432603f
C4807 CSoutput.t7 gnd 0.055875f
C4808 CSoutput.t160 gnd 0.055875f
C4809 CSoutput.n278 gnd 0.431831f
C4810 CSoutput.n279 gnd 0.438308f
C4811 CSoutput.t44 gnd 0.055875f
C4812 CSoutput.t51 gnd 0.055875f
C4813 CSoutput.n280 gnd 0.431831f
C4814 CSoutput.n281 gnd 0.21598f
C4815 CSoutput.t36 gnd 0.055875f
C4816 CSoutput.t161 gnd 0.055875f
C4817 CSoutput.n282 gnd 0.431831f
C4818 CSoutput.n283 gnd 0.21598f
C4819 CSoutput.t41 gnd 0.055875f
C4820 CSoutput.t159 gnd 0.055875f
C4821 CSoutput.n284 gnd 0.431831f
C4822 CSoutput.n285 gnd 0.21598f
C4823 CSoutput.t37 gnd 0.055875f
C4824 CSoutput.t28 gnd 0.055875f
C4825 CSoutput.n286 gnd 0.431831f
C4826 CSoutput.n287 gnd 0.21598f
C4827 CSoutput.t42 gnd 0.055875f
C4828 CSoutput.t23 gnd 0.055875f
C4829 CSoutput.n288 gnd 0.431831f
C4830 CSoutput.n289 gnd 0.21598f
C4831 CSoutput.t165 gnd 0.055875f
C4832 CSoutput.t55 gnd 0.055875f
C4833 CSoutput.n290 gnd 0.431831f
C4834 CSoutput.n291 gnd 0.396057f
C4835 CSoutput.t162 gnd 0.055875f
C4836 CSoutput.t171 gnd 0.055875f
C4837 CSoutput.n292 gnd 0.432603f
C4838 CSoutput.t57 gnd 0.055875f
C4839 CSoutput.t67 gnd 0.055875f
C4840 CSoutput.n293 gnd 0.431831f
C4841 CSoutput.n294 gnd 0.438308f
C4842 CSoutput.t170 gnd 0.055875f
C4843 CSoutput.t45 gnd 0.055875f
C4844 CSoutput.n295 gnd 0.431831f
C4845 CSoutput.n296 gnd 0.21598f
C4846 CSoutput.t5 gnd 0.055875f
C4847 CSoutput.t77 gnd 0.055875f
C4848 CSoutput.n297 gnd 0.431831f
C4849 CSoutput.n298 gnd 0.21598f
C4850 CSoutput.t75 gnd 0.055875f
C4851 CSoutput.t60 gnd 0.055875f
C4852 CSoutput.n299 gnd 0.431831f
C4853 CSoutput.n300 gnd 0.21598f
C4854 CSoutput.t52 gnd 0.055875f
C4855 CSoutput.t13 gnd 0.055875f
C4856 CSoutput.n301 gnd 0.431831f
C4857 CSoutput.n302 gnd 0.21598f
C4858 CSoutput.t76 gnd 0.055875f
C4859 CSoutput.t10 gnd 0.055875f
C4860 CSoutput.n303 gnd 0.431831f
C4861 CSoutput.n304 gnd 0.21598f
C4862 CSoutput.t59 gnd 0.055875f
C4863 CSoutput.t35 gnd 0.055875f
C4864 CSoutput.n305 gnd 0.431831f
C4865 CSoutput.n306 gnd 0.32208f
C4866 CSoutput.n307 gnd 0.406141f
C4867 CSoutput.t19 gnd 0.055875f
C4868 CSoutput.t56 gnd 0.055875f
C4869 CSoutput.n308 gnd 0.432603f
C4870 CSoutput.t64 gnd 0.055875f
C4871 CSoutput.t54 gnd 0.055875f
C4872 CSoutput.n309 gnd 0.431831f
C4873 CSoutput.n310 gnd 0.438308f
C4874 CSoutput.t70 gnd 0.055875f
C4875 CSoutput.t22 gnd 0.055875f
C4876 CSoutput.n311 gnd 0.431831f
C4877 CSoutput.n312 gnd 0.21598f
C4878 CSoutput.t26 gnd 0.055875f
C4879 CSoutput.t43 gnd 0.055875f
C4880 CSoutput.n313 gnd 0.431831f
C4881 CSoutput.n314 gnd 0.21598f
C4882 CSoutput.t169 gnd 0.055875f
C4883 CSoutput.t174 gnd 0.055875f
C4884 CSoutput.n315 gnd 0.431831f
C4885 CSoutput.n316 gnd 0.21598f
C4886 CSoutput.t53 gnd 0.055875f
C4887 CSoutput.t12 gnd 0.055875f
C4888 CSoutput.n317 gnd 0.431831f
C4889 CSoutput.n318 gnd 0.21598f
C4890 CSoutput.t39 gnd 0.055875f
C4891 CSoutput.t15 gnd 0.055875f
C4892 CSoutput.n319 gnd 0.431831f
C4893 CSoutput.n320 gnd 0.21598f
C4894 CSoutput.t158 gnd 0.055875f
C4895 CSoutput.t4 gnd 0.055875f
C4896 CSoutput.n321 gnd 0.43183f
C4897 CSoutput.n322 gnd 0.322082f
C4898 CSoutput.n323 gnd 0.453962f
C4899 CSoutput.n324 gnd 12.459499f
C4900 CSoutput.t113 gnd 0.048891f
C4901 CSoutput.t133 gnd 0.048891f
C4902 CSoutput.n325 gnd 0.433461f
C4903 CSoutput.t89 gnd 0.048891f
C4904 CSoutput.t90 gnd 0.048891f
C4905 CSoutput.n326 gnd 0.432015f
C4906 CSoutput.n327 gnd 0.402557f
C4907 CSoutput.t123 gnd 0.048891f
C4908 CSoutput.t152 gnd 0.048891f
C4909 CSoutput.n328 gnd 0.432015f
C4910 CSoutput.n329 gnd 0.198442f
C4911 CSoutput.t81 gnd 0.048891f
C4912 CSoutput.t114 gnd 0.048891f
C4913 CSoutput.n330 gnd 0.432015f
C4914 CSoutput.n331 gnd 0.198442f
C4915 CSoutput.t104 gnd 0.048891f
C4916 CSoutput.t137 gnd 0.048891f
C4917 CSoutput.n332 gnd 0.432015f
C4918 CSoutput.n333 gnd 0.198442f
C4919 CSoutput.t107 gnd 0.048891f
C4920 CSoutput.t110 gnd 0.048891f
C4921 CSoutput.n334 gnd 0.432015f
C4922 CSoutput.n335 gnd 0.198442f
C4923 CSoutput.t128 gnd 0.048891f
C4924 CSoutput.t130 gnd 0.048891f
C4925 CSoutput.n336 gnd 0.432015f
C4926 CSoutput.n337 gnd 0.198442f
C4927 CSoutput.t103 gnd 0.048891f
C4928 CSoutput.t119 gnd 0.048891f
C4929 CSoutput.n338 gnd 0.432015f
C4930 CSoutput.n339 gnd 0.198442f
C4931 CSoutput.t138 gnd 0.048891f
C4932 CSoutput.t93 gnd 0.048891f
C4933 CSoutput.n340 gnd 0.432015f
C4934 CSoutput.n341 gnd 0.198442f
C4935 CSoutput.t80 gnd 0.048891f
C4936 CSoutput.t111 gnd 0.048891f
C4937 CSoutput.n342 gnd 0.432015f
C4938 CSoutput.n343 gnd 0.365966f
C4939 CSoutput.t96 gnd 0.048891f
C4940 CSoutput.t129 gnd 0.048891f
C4941 CSoutput.n344 gnd 0.433461f
C4942 CSoutput.t83 gnd 0.048891f
C4943 CSoutput.t86 gnd 0.048891f
C4944 CSoutput.n345 gnd 0.432015f
C4945 CSoutput.n346 gnd 0.402557f
C4946 CSoutput.t105 gnd 0.048891f
C4947 CSoutput.t121 gnd 0.048891f
C4948 CSoutput.n347 gnd 0.432015f
C4949 CSoutput.n348 gnd 0.198442f
C4950 CSoutput.t140 gnd 0.048891f
C4951 CSoutput.t99 gnd 0.048891f
C4952 CSoutput.n349 gnd 0.432015f
C4953 CSoutput.n350 gnd 0.198442f
C4954 CSoutput.t102 gnd 0.048891f
C4955 CSoutput.t117 gnd 0.048891f
C4956 CSoutput.n351 gnd 0.432015f
C4957 CSoutput.n352 gnd 0.198442f
C4958 CSoutput.t87 gnd 0.048891f
C4959 CSoutput.t98 gnd 0.048891f
C4960 CSoutput.n353 gnd 0.432015f
C4961 CSoutput.n354 gnd 0.198442f
C4962 CSoutput.t109 gnd 0.048891f
C4963 CSoutput.t127 gnd 0.048891f
C4964 CSoutput.n355 gnd 0.432015f
C4965 CSoutput.n356 gnd 0.198442f
C4966 CSoutput.t79 gnd 0.048891f
C4967 CSoutput.t97 gnd 0.048891f
C4968 CSoutput.n357 gnd 0.432015f
C4969 CSoutput.n358 gnd 0.198442f
C4970 CSoutput.t118 gnd 0.048891f
C4971 CSoutput.t146 gnd 0.048891f
C4972 CSoutput.n359 gnd 0.432015f
C4973 CSoutput.n360 gnd 0.198442f
C4974 CSoutput.t139 gnd 0.048891f
C4975 CSoutput.t95 gnd 0.048891f
C4976 CSoutput.n361 gnd 0.432015f
C4977 CSoutput.n362 gnd 0.301277f
C4978 CSoutput.n363 gnd 0.559795f
C4979 CSoutput.n364 gnd 13.2863f
C4980 CSoutput.t150 gnd 0.048891f
C4981 CSoutput.t156 gnd 0.048891f
C4982 CSoutput.n365 gnd 0.433461f
C4983 CSoutput.t120 gnd 0.048891f
C4984 CSoutput.t94 gnd 0.048891f
C4985 CSoutput.n366 gnd 0.432015f
C4986 CSoutput.n367 gnd 0.402557f
C4987 CSoutput.t84 gnd 0.048891f
C4988 CSoutput.t151 gnd 0.048891f
C4989 CSoutput.n368 gnd 0.432015f
C4990 CSoutput.n369 gnd 0.198442f
C4991 CSoutput.t157 gnd 0.048891f
C4992 CSoutput.t147 gnd 0.048891f
C4993 CSoutput.n370 gnd 0.432015f
C4994 CSoutput.n371 gnd 0.198442f
C4995 CSoutput.t143 gnd 0.048891f
C4996 CSoutput.t135 gnd 0.048891f
C4997 CSoutput.n372 gnd 0.432015f
C4998 CSoutput.n373 gnd 0.198442f
C4999 CSoutput.t125 gnd 0.048891f
C5000 CSoutput.t101 gnd 0.048891f
C5001 CSoutput.n374 gnd 0.432015f
C5002 CSoutput.n375 gnd 0.198442f
C5003 CSoutput.t148 gnd 0.048891f
C5004 CSoutput.t78 gnd 0.048891f
C5005 CSoutput.n376 gnd 0.432015f
C5006 CSoutput.n377 gnd 0.198442f
C5007 CSoutput.t134 gnd 0.048891f
C5008 CSoutput.t116 gnd 0.048891f
C5009 CSoutput.n378 gnd 0.432015f
C5010 CSoutput.n379 gnd 0.198442f
C5011 CSoutput.t82 gnd 0.048891f
C5012 CSoutput.t141 gnd 0.048891f
C5013 CSoutput.n380 gnd 0.432015f
C5014 CSoutput.n381 gnd 0.198442f
C5015 CSoutput.t124 gnd 0.048891f
C5016 CSoutput.t92 gnd 0.048891f
C5017 CSoutput.n382 gnd 0.432015f
C5018 CSoutput.n383 gnd 0.365966f
C5019 CSoutput.t155 gnd 0.048891f
C5020 CSoutput.t126 gnd 0.048891f
C5021 CSoutput.n384 gnd 0.433461f
C5022 CSoutput.t88 gnd 0.048891f
C5023 CSoutput.t149 gnd 0.048891f
C5024 CSoutput.n385 gnd 0.432015f
C5025 CSoutput.n386 gnd 0.402557f
C5026 CSoutput.t144 gnd 0.048891f
C5027 CSoutput.t136 gnd 0.048891f
C5028 CSoutput.n387 gnd 0.432015f
C5029 CSoutput.n388 gnd 0.198442f
C5030 CSoutput.t85 gnd 0.048891f
C5031 CSoutput.t153 gnd 0.048891f
C5032 CSoutput.n389 gnd 0.432015f
C5033 CSoutput.n390 gnd 0.198442f
C5034 CSoutput.t131 gnd 0.048891f
C5035 CSoutput.t115 gnd 0.048891f
C5036 CSoutput.n391 gnd 0.432015f
C5037 CSoutput.n392 gnd 0.198442f
C5038 CSoutput.t108 gnd 0.048891f
C5039 CSoutput.t91 gnd 0.048891f
C5040 CSoutput.n393 gnd 0.432015f
C5041 CSoutput.n394 gnd 0.198442f
C5042 CSoutput.t154 gnd 0.048891f
C5043 CSoutput.t122 gnd 0.048891f
C5044 CSoutput.n395 gnd 0.432015f
C5045 CSoutput.n396 gnd 0.198442f
C5046 CSoutput.t112 gnd 0.048891f
C5047 CSoutput.t100 gnd 0.048891f
C5048 CSoutput.n397 gnd 0.432015f
C5049 CSoutput.n398 gnd 0.198442f
C5050 CSoutput.t142 gnd 0.048891f
C5051 CSoutput.t132 gnd 0.048891f
C5052 CSoutput.n399 gnd 0.432015f
C5053 CSoutput.n400 gnd 0.198442f
C5054 CSoutput.t106 gnd 0.048891f
C5055 CSoutput.t145 gnd 0.048891f
C5056 CSoutput.n401 gnd 0.432015f
C5057 CSoutput.n402 gnd 0.301277f
C5058 CSoutput.n403 gnd 0.559795f
C5059 CSoutput.n404 gnd 7.87078f
C5060 CSoutput.n405 gnd 14.572201f
C5061 commonsourceibias.n0 gnd 0.010705f
C5062 commonsourceibias.t117 gnd 0.162096f
C5063 commonsourceibias.t135 gnd 0.149881f
C5064 commonsourceibias.n1 gnd 0.007808f
C5065 commonsourceibias.n2 gnd 0.008022f
C5066 commonsourceibias.t92 gnd 0.149881f
C5067 commonsourceibias.n3 gnd 0.010321f
C5068 commonsourceibias.n4 gnd 0.008022f
C5069 commonsourceibias.t90 gnd 0.149881f
C5070 commonsourceibias.n5 gnd 0.059802f
C5071 commonsourceibias.t127 gnd 0.149881f
C5072 commonsourceibias.n6 gnd 0.007564f
C5073 commonsourceibias.n7 gnd 0.008022f
C5074 commonsourceibias.t145 gnd 0.149881f
C5075 commonsourceibias.n8 gnd 0.010168f
C5076 commonsourceibias.n9 gnd 0.008022f
C5077 commonsourceibias.t83 gnd 0.149881f
C5078 commonsourceibias.n10 gnd 0.059802f
C5079 commonsourceibias.t116 gnd 0.149881f
C5080 commonsourceibias.n11 gnd 0.007348f
C5081 commonsourceibias.n12 gnd 0.008022f
C5082 commonsourceibias.t110 gnd 0.149881f
C5083 commonsourceibias.n13 gnd 0.009997f
C5084 commonsourceibias.n14 gnd 0.010705f
C5085 commonsourceibias.t32 gnd 0.162096f
C5086 commonsourceibias.t66 gnd 0.149881f
C5087 commonsourceibias.n15 gnd 0.007808f
C5088 commonsourceibias.n16 gnd 0.008022f
C5089 commonsourceibias.t40 gnd 0.149881f
C5090 commonsourceibias.n17 gnd 0.010321f
C5091 commonsourceibias.n18 gnd 0.008022f
C5092 commonsourceibias.t30 gnd 0.149881f
C5093 commonsourceibias.n19 gnd 0.059802f
C5094 commonsourceibias.t50 gnd 0.149881f
C5095 commonsourceibias.n20 gnd 0.007564f
C5096 commonsourceibias.n21 gnd 0.008022f
C5097 commonsourceibias.t36 gnd 0.149881f
C5098 commonsourceibias.n22 gnd 0.010168f
C5099 commonsourceibias.n23 gnd 0.008022f
C5100 commonsourceibias.t2 gnd 0.149881f
C5101 commonsourceibias.n24 gnd 0.059802f
C5102 commonsourceibias.t46 gnd 0.149881f
C5103 commonsourceibias.n25 gnd 0.007348f
C5104 commonsourceibias.n26 gnd 0.008022f
C5105 commonsourceibias.t34 gnd 0.149881f
C5106 commonsourceibias.n27 gnd 0.009997f
C5107 commonsourceibias.n28 gnd 0.008022f
C5108 commonsourceibias.t72 gnd 0.149881f
C5109 commonsourceibias.n29 gnd 0.059802f
C5110 commonsourceibias.t24 gnd 0.149881f
C5111 commonsourceibias.n30 gnd 0.007159f
C5112 commonsourceibias.n31 gnd 0.008022f
C5113 commonsourceibias.t4 gnd 0.149881f
C5114 commonsourceibias.n32 gnd 0.009806f
C5115 commonsourceibias.n33 gnd 0.008022f
C5116 commonsourceibias.t58 gnd 0.149881f
C5117 commonsourceibias.n34 gnd 0.059802f
C5118 commonsourceibias.t16 gnd 0.149881f
C5119 commonsourceibias.n35 gnd 0.006995f
C5120 commonsourceibias.n36 gnd 0.008022f
C5121 commonsourceibias.t74 gnd 0.149881f
C5122 commonsourceibias.n37 gnd 0.009595f
C5123 commonsourceibias.n38 gnd 0.008022f
C5124 commonsourceibias.t48 gnd 0.149881f
C5125 commonsourceibias.n39 gnd 0.059802f
C5126 commonsourceibias.t8 gnd 0.149881f
C5127 commonsourceibias.n40 gnd 0.006855f
C5128 commonsourceibias.n41 gnd 0.008022f
C5129 commonsourceibias.t70 gnd 0.149881f
C5130 commonsourceibias.n42 gnd 0.00936f
C5131 commonsourceibias.t20 gnd 0.16664f
C5132 commonsourceibias.t64 gnd 0.149881f
C5133 commonsourceibias.n43 gnd 0.065328f
C5134 commonsourceibias.n44 gnd 0.07169f
C5135 commonsourceibias.n45 gnd 0.033265f
C5136 commonsourceibias.n46 gnd 0.008022f
C5137 commonsourceibias.n47 gnd 0.007808f
C5138 commonsourceibias.n48 gnd 0.01119f
C5139 commonsourceibias.n49 gnd 0.059802f
C5140 commonsourceibias.n50 gnd 0.011182f
C5141 commonsourceibias.n51 gnd 0.008022f
C5142 commonsourceibias.n52 gnd 0.008022f
C5143 commonsourceibias.n53 gnd 0.008022f
C5144 commonsourceibias.n54 gnd 0.010321f
C5145 commonsourceibias.n55 gnd 0.059802f
C5146 commonsourceibias.n56 gnd 0.010563f
C5147 commonsourceibias.n57 gnd 0.010263f
C5148 commonsourceibias.n58 gnd 0.008022f
C5149 commonsourceibias.n59 gnd 0.008022f
C5150 commonsourceibias.n60 gnd 0.008022f
C5151 commonsourceibias.n61 gnd 0.007564f
C5152 commonsourceibias.n62 gnd 0.0112f
C5153 commonsourceibias.n63 gnd 0.059802f
C5154 commonsourceibias.n64 gnd 0.011196f
C5155 commonsourceibias.n65 gnd 0.008022f
C5156 commonsourceibias.n66 gnd 0.008022f
C5157 commonsourceibias.n67 gnd 0.008022f
C5158 commonsourceibias.n68 gnd 0.010168f
C5159 commonsourceibias.n69 gnd 0.059802f
C5160 commonsourceibias.n70 gnd 0.010488f
C5161 commonsourceibias.n71 gnd 0.010338f
C5162 commonsourceibias.n72 gnd 0.008022f
C5163 commonsourceibias.n73 gnd 0.008022f
C5164 commonsourceibias.n74 gnd 0.008022f
C5165 commonsourceibias.n75 gnd 0.007348f
C5166 commonsourceibias.n76 gnd 0.011204f
C5167 commonsourceibias.n77 gnd 0.059802f
C5168 commonsourceibias.n78 gnd 0.011203f
C5169 commonsourceibias.n79 gnd 0.008022f
C5170 commonsourceibias.n80 gnd 0.008022f
C5171 commonsourceibias.n81 gnd 0.008022f
C5172 commonsourceibias.n82 gnd 0.009997f
C5173 commonsourceibias.n83 gnd 0.059802f
C5174 commonsourceibias.n84 gnd 0.010413f
C5175 commonsourceibias.n85 gnd 0.010413f
C5176 commonsourceibias.n86 gnd 0.008022f
C5177 commonsourceibias.n87 gnd 0.008022f
C5178 commonsourceibias.n88 gnd 0.008022f
C5179 commonsourceibias.n89 gnd 0.007159f
C5180 commonsourceibias.n90 gnd 0.011203f
C5181 commonsourceibias.n91 gnd 0.059802f
C5182 commonsourceibias.n92 gnd 0.011204f
C5183 commonsourceibias.n93 gnd 0.008022f
C5184 commonsourceibias.n94 gnd 0.008022f
C5185 commonsourceibias.n95 gnd 0.008022f
C5186 commonsourceibias.n96 gnd 0.009806f
C5187 commonsourceibias.n97 gnd 0.059802f
C5188 commonsourceibias.n98 gnd 0.010338f
C5189 commonsourceibias.n99 gnd 0.010488f
C5190 commonsourceibias.n100 gnd 0.008022f
C5191 commonsourceibias.n101 gnd 0.008022f
C5192 commonsourceibias.n102 gnd 0.008022f
C5193 commonsourceibias.n103 gnd 0.006995f
C5194 commonsourceibias.n104 gnd 0.011196f
C5195 commonsourceibias.n105 gnd 0.059802f
C5196 commonsourceibias.n106 gnd 0.0112f
C5197 commonsourceibias.n107 gnd 0.008022f
C5198 commonsourceibias.n108 gnd 0.008022f
C5199 commonsourceibias.n109 gnd 0.008022f
C5200 commonsourceibias.n110 gnd 0.009595f
C5201 commonsourceibias.n111 gnd 0.059802f
C5202 commonsourceibias.n112 gnd 0.010263f
C5203 commonsourceibias.n113 gnd 0.010563f
C5204 commonsourceibias.n114 gnd 0.008022f
C5205 commonsourceibias.n115 gnd 0.008022f
C5206 commonsourceibias.n116 gnd 0.008022f
C5207 commonsourceibias.n117 gnd 0.006855f
C5208 commonsourceibias.n118 gnd 0.011182f
C5209 commonsourceibias.n119 gnd 0.059802f
C5210 commonsourceibias.n120 gnd 0.01119f
C5211 commonsourceibias.n121 gnd 0.008022f
C5212 commonsourceibias.n122 gnd 0.008022f
C5213 commonsourceibias.n123 gnd 0.008022f
C5214 commonsourceibias.n124 gnd 0.00936f
C5215 commonsourceibias.n125 gnd 0.059802f
C5216 commonsourceibias.n126 gnd 0.009843f
C5217 commonsourceibias.n127 gnd 0.071758f
C5218 commonsourceibias.n128 gnd 0.079928f
C5219 commonsourceibias.t33 gnd 0.017311f
C5220 commonsourceibias.t67 gnd 0.017311f
C5221 commonsourceibias.n129 gnd 0.152968f
C5222 commonsourceibias.n130 gnd 0.132319f
C5223 commonsourceibias.t41 gnd 0.017311f
C5224 commonsourceibias.t31 gnd 0.017311f
C5225 commonsourceibias.n131 gnd 0.152968f
C5226 commonsourceibias.n132 gnd 0.070264f
C5227 commonsourceibias.t51 gnd 0.017311f
C5228 commonsourceibias.t37 gnd 0.017311f
C5229 commonsourceibias.n133 gnd 0.152968f
C5230 commonsourceibias.n134 gnd 0.070264f
C5231 commonsourceibias.t3 gnd 0.017311f
C5232 commonsourceibias.t47 gnd 0.017311f
C5233 commonsourceibias.n135 gnd 0.152968f
C5234 commonsourceibias.n136 gnd 0.070264f
C5235 commonsourceibias.t35 gnd 0.017311f
C5236 commonsourceibias.t73 gnd 0.017311f
C5237 commonsourceibias.n137 gnd 0.152968f
C5238 commonsourceibias.n138 gnd 0.058702f
C5239 commonsourceibias.t65 gnd 0.017311f
C5240 commonsourceibias.t21 gnd 0.017311f
C5241 commonsourceibias.n139 gnd 0.15348f
C5242 commonsourceibias.t9 gnd 0.017311f
C5243 commonsourceibias.t71 gnd 0.017311f
C5244 commonsourceibias.n140 gnd 0.152968f
C5245 commonsourceibias.n141 gnd 0.142538f
C5246 commonsourceibias.t75 gnd 0.017311f
C5247 commonsourceibias.t49 gnd 0.017311f
C5248 commonsourceibias.n142 gnd 0.152968f
C5249 commonsourceibias.n143 gnd 0.070264f
C5250 commonsourceibias.t59 gnd 0.017311f
C5251 commonsourceibias.t17 gnd 0.017311f
C5252 commonsourceibias.n144 gnd 0.152968f
C5253 commonsourceibias.n145 gnd 0.070264f
C5254 commonsourceibias.t25 gnd 0.017311f
C5255 commonsourceibias.t5 gnd 0.017311f
C5256 commonsourceibias.n146 gnd 0.152968f
C5257 commonsourceibias.n147 gnd 0.058702f
C5258 commonsourceibias.n148 gnd 0.071082f
C5259 commonsourceibias.n149 gnd 0.05192f
C5260 commonsourceibias.t131 gnd 0.149881f
C5261 commonsourceibias.n150 gnd 0.059802f
C5262 commonsourceibias.t107 gnd 0.149881f
C5263 commonsourceibias.n151 gnd 0.059802f
C5264 commonsourceibias.n152 gnd 0.008022f
C5265 commonsourceibias.t103 gnd 0.149881f
C5266 commonsourceibias.n153 gnd 0.059802f
C5267 commonsourceibias.n154 gnd 0.008022f
C5268 commonsourceibias.t121 gnd 0.149881f
C5269 commonsourceibias.n155 gnd 0.059802f
C5270 commonsourceibias.n156 gnd 0.008022f
C5271 commonsourceibias.t138 gnd 0.149881f
C5272 commonsourceibias.n157 gnd 0.006995f
C5273 commonsourceibias.n158 gnd 0.008022f
C5274 commonsourceibias.t95 gnd 0.149881f
C5275 commonsourceibias.n159 gnd 0.009595f
C5276 commonsourceibias.n160 gnd 0.008022f
C5277 commonsourceibias.t111 gnd 0.149881f
C5278 commonsourceibias.n161 gnd 0.059802f
C5279 commonsourceibias.t130 gnd 0.149881f
C5280 commonsourceibias.n162 gnd 0.006855f
C5281 commonsourceibias.n163 gnd 0.008022f
C5282 commonsourceibias.t87 gnd 0.149881f
C5283 commonsourceibias.n164 gnd 0.00936f
C5284 commonsourceibias.t119 gnd 0.16664f
C5285 commonsourceibias.t84 gnd 0.149881f
C5286 commonsourceibias.n165 gnd 0.065328f
C5287 commonsourceibias.n166 gnd 0.07169f
C5288 commonsourceibias.n167 gnd 0.033265f
C5289 commonsourceibias.n168 gnd 0.008022f
C5290 commonsourceibias.n169 gnd 0.007808f
C5291 commonsourceibias.n170 gnd 0.01119f
C5292 commonsourceibias.n171 gnd 0.059802f
C5293 commonsourceibias.n172 gnd 0.011182f
C5294 commonsourceibias.n173 gnd 0.008022f
C5295 commonsourceibias.n174 gnd 0.008022f
C5296 commonsourceibias.n175 gnd 0.008022f
C5297 commonsourceibias.n176 gnd 0.010321f
C5298 commonsourceibias.n177 gnd 0.059802f
C5299 commonsourceibias.n178 gnd 0.010563f
C5300 commonsourceibias.n179 gnd 0.010263f
C5301 commonsourceibias.n180 gnd 0.008022f
C5302 commonsourceibias.n181 gnd 0.008022f
C5303 commonsourceibias.n182 gnd 0.008022f
C5304 commonsourceibias.n183 gnd 0.007564f
C5305 commonsourceibias.n184 gnd 0.0112f
C5306 commonsourceibias.n185 gnd 0.059802f
C5307 commonsourceibias.n186 gnd 0.011196f
C5308 commonsourceibias.n187 gnd 0.008022f
C5309 commonsourceibias.n188 gnd 0.008022f
C5310 commonsourceibias.n189 gnd 0.008022f
C5311 commonsourceibias.n190 gnd 0.010168f
C5312 commonsourceibias.n191 gnd 0.059802f
C5313 commonsourceibias.n192 gnd 0.010488f
C5314 commonsourceibias.n193 gnd 0.010338f
C5315 commonsourceibias.n194 gnd 0.008022f
C5316 commonsourceibias.n195 gnd 0.008022f
C5317 commonsourceibias.n196 gnd 0.009806f
C5318 commonsourceibias.n197 gnd 0.007348f
C5319 commonsourceibias.n198 gnd 0.011204f
C5320 commonsourceibias.n199 gnd 0.008022f
C5321 commonsourceibias.n200 gnd 0.008022f
C5322 commonsourceibias.n201 gnd 0.011203f
C5323 commonsourceibias.n202 gnd 0.007159f
C5324 commonsourceibias.n203 gnd 0.009997f
C5325 commonsourceibias.n204 gnd 0.008022f
C5326 commonsourceibias.n205 gnd 0.007008f
C5327 commonsourceibias.n206 gnd 0.010413f
C5328 commonsourceibias.n207 gnd 0.010413f
C5329 commonsourceibias.n208 gnd 0.007008f
C5330 commonsourceibias.n209 gnd 0.008022f
C5331 commonsourceibias.n210 gnd 0.008022f
C5332 commonsourceibias.n211 gnd 0.007159f
C5333 commonsourceibias.n212 gnd 0.011203f
C5334 commonsourceibias.n213 gnd 0.059802f
C5335 commonsourceibias.n214 gnd 0.011204f
C5336 commonsourceibias.n215 gnd 0.008022f
C5337 commonsourceibias.n216 gnd 0.008022f
C5338 commonsourceibias.n217 gnd 0.008022f
C5339 commonsourceibias.n218 gnd 0.009806f
C5340 commonsourceibias.n219 gnd 0.059802f
C5341 commonsourceibias.n220 gnd 0.010338f
C5342 commonsourceibias.n221 gnd 0.010488f
C5343 commonsourceibias.n222 gnd 0.008022f
C5344 commonsourceibias.n223 gnd 0.008022f
C5345 commonsourceibias.n224 gnd 0.008022f
C5346 commonsourceibias.n225 gnd 0.006995f
C5347 commonsourceibias.n226 gnd 0.011196f
C5348 commonsourceibias.n227 gnd 0.059802f
C5349 commonsourceibias.n228 gnd 0.0112f
C5350 commonsourceibias.n229 gnd 0.008022f
C5351 commonsourceibias.n230 gnd 0.008022f
C5352 commonsourceibias.n231 gnd 0.008022f
C5353 commonsourceibias.n232 gnd 0.009595f
C5354 commonsourceibias.n233 gnd 0.059802f
C5355 commonsourceibias.n234 gnd 0.010263f
C5356 commonsourceibias.n235 gnd 0.010563f
C5357 commonsourceibias.n236 gnd 0.008022f
C5358 commonsourceibias.n237 gnd 0.008022f
C5359 commonsourceibias.n238 gnd 0.008022f
C5360 commonsourceibias.n239 gnd 0.006855f
C5361 commonsourceibias.n240 gnd 0.011182f
C5362 commonsourceibias.n241 gnd 0.059802f
C5363 commonsourceibias.n242 gnd 0.01119f
C5364 commonsourceibias.n243 gnd 0.008022f
C5365 commonsourceibias.n244 gnd 0.008022f
C5366 commonsourceibias.n245 gnd 0.008022f
C5367 commonsourceibias.n246 gnd 0.00936f
C5368 commonsourceibias.n247 gnd 0.059802f
C5369 commonsourceibias.n248 gnd 0.009843f
C5370 commonsourceibias.n249 gnd 0.071758f
C5371 commonsourceibias.n250 gnd 0.046883f
C5372 commonsourceibias.n251 gnd 0.010705f
C5373 commonsourceibias.t120 gnd 0.149881f
C5374 commonsourceibias.n252 gnd 0.007808f
C5375 commonsourceibias.n253 gnd 0.008022f
C5376 commonsourceibias.t81 gnd 0.149881f
C5377 commonsourceibias.n254 gnd 0.010321f
C5378 commonsourceibias.n255 gnd 0.008022f
C5379 commonsourceibias.t159 gnd 0.149881f
C5380 commonsourceibias.n256 gnd 0.059802f
C5381 commonsourceibias.t109 gnd 0.149881f
C5382 commonsourceibias.n257 gnd 0.007564f
C5383 commonsourceibias.n258 gnd 0.008022f
C5384 commonsourceibias.t129 gnd 0.149881f
C5385 commonsourceibias.n259 gnd 0.010168f
C5386 commonsourceibias.n260 gnd 0.008022f
C5387 commonsourceibias.t151 gnd 0.149881f
C5388 commonsourceibias.n261 gnd 0.059802f
C5389 commonsourceibias.t100 gnd 0.149881f
C5390 commonsourceibias.n262 gnd 0.007348f
C5391 commonsourceibias.n263 gnd 0.008022f
C5392 commonsourceibias.t96 gnd 0.149881f
C5393 commonsourceibias.n264 gnd 0.009997f
C5394 commonsourceibias.n265 gnd 0.008022f
C5395 commonsourceibias.t113 gnd 0.149881f
C5396 commonsourceibias.n266 gnd 0.059802f
C5397 commonsourceibias.t94 gnd 0.149881f
C5398 commonsourceibias.n267 gnd 0.007159f
C5399 commonsourceibias.n268 gnd 0.008022f
C5400 commonsourceibias.t91 gnd 0.149881f
C5401 commonsourceibias.n269 gnd 0.009806f
C5402 commonsourceibias.n270 gnd 0.008022f
C5403 commonsourceibias.t104 gnd 0.149881f
C5404 commonsourceibias.n271 gnd 0.059802f
C5405 commonsourceibias.t122 gnd 0.149881f
C5406 commonsourceibias.n272 gnd 0.006995f
C5407 commonsourceibias.n273 gnd 0.008022f
C5408 commonsourceibias.t85 gnd 0.149881f
C5409 commonsourceibias.n274 gnd 0.009595f
C5410 commonsourceibias.n275 gnd 0.008022f
C5411 commonsourceibias.t97 gnd 0.149881f
C5412 commonsourceibias.n276 gnd 0.059802f
C5413 commonsourceibias.t112 gnd 0.149881f
C5414 commonsourceibias.n277 gnd 0.006855f
C5415 commonsourceibias.n278 gnd 0.008022f
C5416 commonsourceibias.t157 gnd 0.149881f
C5417 commonsourceibias.n279 gnd 0.00936f
C5418 commonsourceibias.t102 gnd 0.16664f
C5419 commonsourceibias.t152 gnd 0.149881f
C5420 commonsourceibias.n280 gnd 0.065328f
C5421 commonsourceibias.n281 gnd 0.07169f
C5422 commonsourceibias.n282 gnd 0.033265f
C5423 commonsourceibias.n283 gnd 0.008022f
C5424 commonsourceibias.n284 gnd 0.007808f
C5425 commonsourceibias.n285 gnd 0.01119f
C5426 commonsourceibias.n286 gnd 0.059802f
C5427 commonsourceibias.n287 gnd 0.011182f
C5428 commonsourceibias.n288 gnd 0.008022f
C5429 commonsourceibias.n289 gnd 0.008022f
C5430 commonsourceibias.n290 gnd 0.008022f
C5431 commonsourceibias.n291 gnd 0.010321f
C5432 commonsourceibias.n292 gnd 0.059802f
C5433 commonsourceibias.n293 gnd 0.010563f
C5434 commonsourceibias.n294 gnd 0.010263f
C5435 commonsourceibias.n295 gnd 0.008022f
C5436 commonsourceibias.n296 gnd 0.008022f
C5437 commonsourceibias.n297 gnd 0.008022f
C5438 commonsourceibias.n298 gnd 0.007564f
C5439 commonsourceibias.n299 gnd 0.0112f
C5440 commonsourceibias.n300 gnd 0.059802f
C5441 commonsourceibias.n301 gnd 0.011196f
C5442 commonsourceibias.n302 gnd 0.008022f
C5443 commonsourceibias.n303 gnd 0.008022f
C5444 commonsourceibias.n304 gnd 0.008022f
C5445 commonsourceibias.n305 gnd 0.010168f
C5446 commonsourceibias.n306 gnd 0.059802f
C5447 commonsourceibias.n307 gnd 0.010488f
C5448 commonsourceibias.n308 gnd 0.010338f
C5449 commonsourceibias.n309 gnd 0.008022f
C5450 commonsourceibias.n310 gnd 0.008022f
C5451 commonsourceibias.n311 gnd 0.008022f
C5452 commonsourceibias.n312 gnd 0.007348f
C5453 commonsourceibias.n313 gnd 0.011204f
C5454 commonsourceibias.n314 gnd 0.059802f
C5455 commonsourceibias.n315 gnd 0.011203f
C5456 commonsourceibias.n316 gnd 0.008022f
C5457 commonsourceibias.n317 gnd 0.008022f
C5458 commonsourceibias.n318 gnd 0.008022f
C5459 commonsourceibias.n319 gnd 0.009997f
C5460 commonsourceibias.n320 gnd 0.059802f
C5461 commonsourceibias.n321 gnd 0.010413f
C5462 commonsourceibias.n322 gnd 0.010413f
C5463 commonsourceibias.n323 gnd 0.008022f
C5464 commonsourceibias.n324 gnd 0.008022f
C5465 commonsourceibias.n325 gnd 0.008022f
C5466 commonsourceibias.n326 gnd 0.007159f
C5467 commonsourceibias.n327 gnd 0.011203f
C5468 commonsourceibias.n328 gnd 0.059802f
C5469 commonsourceibias.n329 gnd 0.011204f
C5470 commonsourceibias.n330 gnd 0.008022f
C5471 commonsourceibias.n331 gnd 0.008022f
C5472 commonsourceibias.n332 gnd 0.008022f
C5473 commonsourceibias.n333 gnd 0.009806f
C5474 commonsourceibias.n334 gnd 0.059802f
C5475 commonsourceibias.n335 gnd 0.010338f
C5476 commonsourceibias.n336 gnd 0.010488f
C5477 commonsourceibias.n337 gnd 0.008022f
C5478 commonsourceibias.n338 gnd 0.008022f
C5479 commonsourceibias.n339 gnd 0.008022f
C5480 commonsourceibias.n340 gnd 0.006995f
C5481 commonsourceibias.n341 gnd 0.011196f
C5482 commonsourceibias.n342 gnd 0.059802f
C5483 commonsourceibias.n343 gnd 0.0112f
C5484 commonsourceibias.n344 gnd 0.008022f
C5485 commonsourceibias.n345 gnd 0.008022f
C5486 commonsourceibias.n346 gnd 0.008022f
C5487 commonsourceibias.n347 gnd 0.009595f
C5488 commonsourceibias.n348 gnd 0.059802f
C5489 commonsourceibias.n349 gnd 0.010263f
C5490 commonsourceibias.n350 gnd 0.010563f
C5491 commonsourceibias.n351 gnd 0.008022f
C5492 commonsourceibias.n352 gnd 0.008022f
C5493 commonsourceibias.n353 gnd 0.008022f
C5494 commonsourceibias.n354 gnd 0.006855f
C5495 commonsourceibias.n355 gnd 0.011182f
C5496 commonsourceibias.n356 gnd 0.059802f
C5497 commonsourceibias.n357 gnd 0.01119f
C5498 commonsourceibias.n358 gnd 0.008022f
C5499 commonsourceibias.n359 gnd 0.008022f
C5500 commonsourceibias.n360 gnd 0.008022f
C5501 commonsourceibias.n361 gnd 0.00936f
C5502 commonsourceibias.n362 gnd 0.059802f
C5503 commonsourceibias.n363 gnd 0.009843f
C5504 commonsourceibias.t101 gnd 0.162096f
C5505 commonsourceibias.n364 gnd 0.071758f
C5506 commonsourceibias.n365 gnd 0.024957f
C5507 commonsourceibias.n366 gnd 0.404135f
C5508 commonsourceibias.n367 gnd 0.010705f
C5509 commonsourceibias.t140 gnd 0.162096f
C5510 commonsourceibias.t153 gnd 0.149881f
C5511 commonsourceibias.n368 gnd 0.007808f
C5512 commonsourceibias.n369 gnd 0.008022f
C5513 commonsourceibias.t86 gnd 0.149881f
C5514 commonsourceibias.n370 gnd 0.010321f
C5515 commonsourceibias.n371 gnd 0.008022f
C5516 commonsourceibias.t146 gnd 0.149881f
C5517 commonsourceibias.n372 gnd 0.007564f
C5518 commonsourceibias.n373 gnd 0.008022f
C5519 commonsourceibias.t80 gnd 0.149881f
C5520 commonsourceibias.n374 gnd 0.010168f
C5521 commonsourceibias.n375 gnd 0.008022f
C5522 commonsourceibias.t139 gnd 0.149881f
C5523 commonsourceibias.n376 gnd 0.007348f
C5524 commonsourceibias.n377 gnd 0.008022f
C5525 commonsourceibias.t133 gnd 0.149881f
C5526 commonsourceibias.n378 gnd 0.009997f
C5527 commonsourceibias.t57 gnd 0.017311f
C5528 commonsourceibias.t45 gnd 0.017311f
C5529 commonsourceibias.n379 gnd 0.15348f
C5530 commonsourceibias.t43 gnd 0.017311f
C5531 commonsourceibias.t79 gnd 0.017311f
C5532 commonsourceibias.n380 gnd 0.152968f
C5533 commonsourceibias.n381 gnd 0.142538f
C5534 commonsourceibias.t23 gnd 0.017311f
C5535 commonsourceibias.t55 gnd 0.017311f
C5536 commonsourceibias.n382 gnd 0.152968f
C5537 commonsourceibias.n383 gnd 0.070264f
C5538 commonsourceibias.t15 gnd 0.017311f
C5539 commonsourceibias.t39 gnd 0.017311f
C5540 commonsourceibias.n384 gnd 0.152968f
C5541 commonsourceibias.n385 gnd 0.070264f
C5542 commonsourceibias.t77 gnd 0.017311f
C5543 commonsourceibias.t69 gnd 0.017311f
C5544 commonsourceibias.n386 gnd 0.152968f
C5545 commonsourceibias.n387 gnd 0.058702f
C5546 commonsourceibias.n388 gnd 0.010705f
C5547 commonsourceibias.t52 gnd 0.149881f
C5548 commonsourceibias.n389 gnd 0.007808f
C5549 commonsourceibias.n390 gnd 0.008022f
C5550 commonsourceibias.t18 gnd 0.149881f
C5551 commonsourceibias.n391 gnd 0.010321f
C5552 commonsourceibias.n392 gnd 0.008022f
C5553 commonsourceibias.t28 gnd 0.149881f
C5554 commonsourceibias.n393 gnd 0.007564f
C5555 commonsourceibias.n394 gnd 0.008022f
C5556 commonsourceibias.t12 gnd 0.149881f
C5557 commonsourceibias.n395 gnd 0.010168f
C5558 commonsourceibias.n396 gnd 0.008022f
C5559 commonsourceibias.t26 gnd 0.149881f
C5560 commonsourceibias.n397 gnd 0.007348f
C5561 commonsourceibias.n398 gnd 0.008022f
C5562 commonsourceibias.t10 gnd 0.149881f
C5563 commonsourceibias.n399 gnd 0.009997f
C5564 commonsourceibias.n400 gnd 0.008022f
C5565 commonsourceibias.t68 gnd 0.149881f
C5566 commonsourceibias.n401 gnd 0.007159f
C5567 commonsourceibias.n402 gnd 0.008022f
C5568 commonsourceibias.t76 gnd 0.149881f
C5569 commonsourceibias.n403 gnd 0.009806f
C5570 commonsourceibias.n404 gnd 0.008022f
C5571 commonsourceibias.t14 gnd 0.149881f
C5572 commonsourceibias.n405 gnd 0.006995f
C5573 commonsourceibias.n406 gnd 0.008022f
C5574 commonsourceibias.t54 gnd 0.149881f
C5575 commonsourceibias.n407 gnd 0.009595f
C5576 commonsourceibias.n408 gnd 0.008022f
C5577 commonsourceibias.t78 gnd 0.149881f
C5578 commonsourceibias.n409 gnd 0.006855f
C5579 commonsourceibias.n410 gnd 0.008022f
C5580 commonsourceibias.t42 gnd 0.149881f
C5581 commonsourceibias.n411 gnd 0.00936f
C5582 commonsourceibias.t56 gnd 0.16664f
C5583 commonsourceibias.t44 gnd 0.149881f
C5584 commonsourceibias.n412 gnd 0.065328f
C5585 commonsourceibias.n413 gnd 0.07169f
C5586 commonsourceibias.n414 gnd 0.033265f
C5587 commonsourceibias.n415 gnd 0.008022f
C5588 commonsourceibias.n416 gnd 0.007808f
C5589 commonsourceibias.n417 gnd 0.01119f
C5590 commonsourceibias.n418 gnd 0.059802f
C5591 commonsourceibias.n419 gnd 0.011182f
C5592 commonsourceibias.n420 gnd 0.008022f
C5593 commonsourceibias.n421 gnd 0.008022f
C5594 commonsourceibias.n422 gnd 0.008022f
C5595 commonsourceibias.n423 gnd 0.010321f
C5596 commonsourceibias.n424 gnd 0.059802f
C5597 commonsourceibias.n425 gnd 0.010563f
C5598 commonsourceibias.t22 gnd 0.149881f
C5599 commonsourceibias.n426 gnd 0.059802f
C5600 commonsourceibias.n427 gnd 0.010263f
C5601 commonsourceibias.n428 gnd 0.008022f
C5602 commonsourceibias.n429 gnd 0.008022f
C5603 commonsourceibias.n430 gnd 0.008022f
C5604 commonsourceibias.n431 gnd 0.007564f
C5605 commonsourceibias.n432 gnd 0.0112f
C5606 commonsourceibias.n433 gnd 0.059802f
C5607 commonsourceibias.n434 gnd 0.011196f
C5608 commonsourceibias.n435 gnd 0.008022f
C5609 commonsourceibias.n436 gnd 0.008022f
C5610 commonsourceibias.n437 gnd 0.008022f
C5611 commonsourceibias.n438 gnd 0.010168f
C5612 commonsourceibias.n439 gnd 0.059802f
C5613 commonsourceibias.n440 gnd 0.010488f
C5614 commonsourceibias.t38 gnd 0.149881f
C5615 commonsourceibias.n441 gnd 0.059802f
C5616 commonsourceibias.n442 gnd 0.010338f
C5617 commonsourceibias.n443 gnd 0.008022f
C5618 commonsourceibias.n444 gnd 0.008022f
C5619 commonsourceibias.n445 gnd 0.008022f
C5620 commonsourceibias.n446 gnd 0.007348f
C5621 commonsourceibias.n447 gnd 0.011204f
C5622 commonsourceibias.n448 gnd 0.059802f
C5623 commonsourceibias.n449 gnd 0.011203f
C5624 commonsourceibias.n450 gnd 0.008022f
C5625 commonsourceibias.n451 gnd 0.008022f
C5626 commonsourceibias.n452 gnd 0.008022f
C5627 commonsourceibias.n453 gnd 0.009997f
C5628 commonsourceibias.n454 gnd 0.059802f
C5629 commonsourceibias.n455 gnd 0.010413f
C5630 commonsourceibias.t60 gnd 0.149881f
C5631 commonsourceibias.n456 gnd 0.059802f
C5632 commonsourceibias.n457 gnd 0.010413f
C5633 commonsourceibias.n458 gnd 0.008022f
C5634 commonsourceibias.n459 gnd 0.008022f
C5635 commonsourceibias.n460 gnd 0.008022f
C5636 commonsourceibias.n461 gnd 0.007159f
C5637 commonsourceibias.n462 gnd 0.011203f
C5638 commonsourceibias.n463 gnd 0.059802f
C5639 commonsourceibias.n464 gnd 0.011204f
C5640 commonsourceibias.n465 gnd 0.008022f
C5641 commonsourceibias.n466 gnd 0.008022f
C5642 commonsourceibias.n467 gnd 0.008022f
C5643 commonsourceibias.n468 gnd 0.009806f
C5644 commonsourceibias.n469 gnd 0.059802f
C5645 commonsourceibias.n470 gnd 0.010338f
C5646 commonsourceibias.t62 gnd 0.149881f
C5647 commonsourceibias.n471 gnd 0.059802f
C5648 commonsourceibias.n472 gnd 0.010488f
C5649 commonsourceibias.n473 gnd 0.008022f
C5650 commonsourceibias.n474 gnd 0.008022f
C5651 commonsourceibias.n475 gnd 0.008022f
C5652 commonsourceibias.n476 gnd 0.006995f
C5653 commonsourceibias.n477 gnd 0.011196f
C5654 commonsourceibias.n478 gnd 0.059802f
C5655 commonsourceibias.n479 gnd 0.0112f
C5656 commonsourceibias.n480 gnd 0.008022f
C5657 commonsourceibias.n481 gnd 0.008022f
C5658 commonsourceibias.n482 gnd 0.008022f
C5659 commonsourceibias.n483 gnd 0.009595f
C5660 commonsourceibias.n484 gnd 0.059802f
C5661 commonsourceibias.n485 gnd 0.010263f
C5662 commonsourceibias.t0 gnd 0.149881f
C5663 commonsourceibias.n486 gnd 0.059802f
C5664 commonsourceibias.n487 gnd 0.010563f
C5665 commonsourceibias.n488 gnd 0.008022f
C5666 commonsourceibias.n489 gnd 0.008022f
C5667 commonsourceibias.n490 gnd 0.008022f
C5668 commonsourceibias.n491 gnd 0.006855f
C5669 commonsourceibias.n492 gnd 0.011182f
C5670 commonsourceibias.n493 gnd 0.059802f
C5671 commonsourceibias.n494 gnd 0.01119f
C5672 commonsourceibias.n495 gnd 0.008022f
C5673 commonsourceibias.n496 gnd 0.008022f
C5674 commonsourceibias.n497 gnd 0.008022f
C5675 commonsourceibias.n498 gnd 0.00936f
C5676 commonsourceibias.n499 gnd 0.059802f
C5677 commonsourceibias.n500 gnd 0.009843f
C5678 commonsourceibias.t6 gnd 0.162096f
C5679 commonsourceibias.n501 gnd 0.071758f
C5680 commonsourceibias.n502 gnd 0.079928f
C5681 commonsourceibias.t53 gnd 0.017311f
C5682 commonsourceibias.t7 gnd 0.017311f
C5683 commonsourceibias.n503 gnd 0.152968f
C5684 commonsourceibias.n504 gnd 0.132319f
C5685 commonsourceibias.t1 gnd 0.017311f
C5686 commonsourceibias.t19 gnd 0.017311f
C5687 commonsourceibias.n505 gnd 0.152968f
C5688 commonsourceibias.n506 gnd 0.070264f
C5689 commonsourceibias.t13 gnd 0.017311f
C5690 commonsourceibias.t29 gnd 0.017311f
C5691 commonsourceibias.n507 gnd 0.152968f
C5692 commonsourceibias.n508 gnd 0.070264f
C5693 commonsourceibias.t27 gnd 0.017311f
C5694 commonsourceibias.t63 gnd 0.017311f
C5695 commonsourceibias.n509 gnd 0.152968f
C5696 commonsourceibias.n510 gnd 0.070264f
C5697 commonsourceibias.t61 gnd 0.017311f
C5698 commonsourceibias.t11 gnd 0.017311f
C5699 commonsourceibias.n511 gnd 0.152968f
C5700 commonsourceibias.n512 gnd 0.058702f
C5701 commonsourceibias.n513 gnd 0.071082f
C5702 commonsourceibias.n514 gnd 0.05192f
C5703 commonsourceibias.t98 gnd 0.149881f
C5704 commonsourceibias.n515 gnd 0.059802f
C5705 commonsourceibias.n516 gnd 0.008022f
C5706 commonsourceibias.t125 gnd 0.149881f
C5707 commonsourceibias.n517 gnd 0.059802f
C5708 commonsourceibias.n518 gnd 0.008022f
C5709 commonsourceibias.t142 gnd 0.149881f
C5710 commonsourceibias.n519 gnd 0.059802f
C5711 commonsourceibias.n520 gnd 0.008022f
C5712 commonsourceibias.t155 gnd 0.149881f
C5713 commonsourceibias.n521 gnd 0.006995f
C5714 commonsourceibias.n522 gnd 0.008022f
C5715 commonsourceibias.t114 gnd 0.149881f
C5716 commonsourceibias.n523 gnd 0.009595f
C5717 commonsourceibias.n524 gnd 0.008022f
C5718 commonsourceibias.t148 gnd 0.149881f
C5719 commonsourceibias.n525 gnd 0.006855f
C5720 commonsourceibias.n526 gnd 0.008022f
C5721 commonsourceibias.t82 gnd 0.149881f
C5722 commonsourceibias.n527 gnd 0.00936f
C5723 commonsourceibias.t126 gnd 0.16664f
C5724 commonsourceibias.t89 gnd 0.149881f
C5725 commonsourceibias.n528 gnd 0.065328f
C5726 commonsourceibias.n529 gnd 0.07169f
C5727 commonsourceibias.n530 gnd 0.033265f
C5728 commonsourceibias.n531 gnd 0.008022f
C5729 commonsourceibias.n532 gnd 0.007808f
C5730 commonsourceibias.n533 gnd 0.01119f
C5731 commonsourceibias.n534 gnd 0.059802f
C5732 commonsourceibias.n535 gnd 0.011182f
C5733 commonsourceibias.n536 gnd 0.008022f
C5734 commonsourceibias.n537 gnd 0.008022f
C5735 commonsourceibias.n538 gnd 0.008022f
C5736 commonsourceibias.n539 gnd 0.010321f
C5737 commonsourceibias.n540 gnd 0.059802f
C5738 commonsourceibias.n541 gnd 0.010563f
C5739 commonsourceibias.t134 gnd 0.149881f
C5740 commonsourceibias.n542 gnd 0.059802f
C5741 commonsourceibias.n543 gnd 0.010263f
C5742 commonsourceibias.n544 gnd 0.008022f
C5743 commonsourceibias.n545 gnd 0.008022f
C5744 commonsourceibias.n546 gnd 0.008022f
C5745 commonsourceibias.n547 gnd 0.007564f
C5746 commonsourceibias.n548 gnd 0.0112f
C5747 commonsourceibias.n549 gnd 0.059802f
C5748 commonsourceibias.n550 gnd 0.011196f
C5749 commonsourceibias.n551 gnd 0.008022f
C5750 commonsourceibias.n552 gnd 0.008022f
C5751 commonsourceibias.n553 gnd 0.008022f
C5752 commonsourceibias.n554 gnd 0.010168f
C5753 commonsourceibias.n555 gnd 0.059802f
C5754 commonsourceibias.n556 gnd 0.010488f
C5755 commonsourceibias.n557 gnd 0.010338f
C5756 commonsourceibias.n558 gnd 0.008022f
C5757 commonsourceibias.n559 gnd 0.008022f
C5758 commonsourceibias.n560 gnd 0.009806f
C5759 commonsourceibias.n561 gnd 0.007348f
C5760 commonsourceibias.n562 gnd 0.011204f
C5761 commonsourceibias.n563 gnd 0.008022f
C5762 commonsourceibias.n564 gnd 0.008022f
C5763 commonsourceibias.n565 gnd 0.011203f
C5764 commonsourceibias.n566 gnd 0.007159f
C5765 commonsourceibias.n567 gnd 0.009997f
C5766 commonsourceibias.n568 gnd 0.008022f
C5767 commonsourceibias.n569 gnd 0.007008f
C5768 commonsourceibias.n570 gnd 0.010413f
C5769 commonsourceibias.t149 gnd 0.149881f
C5770 commonsourceibias.n571 gnd 0.059802f
C5771 commonsourceibias.n572 gnd 0.010413f
C5772 commonsourceibias.n573 gnd 0.007008f
C5773 commonsourceibias.n574 gnd 0.008022f
C5774 commonsourceibias.n575 gnd 0.008022f
C5775 commonsourceibias.n576 gnd 0.007159f
C5776 commonsourceibias.n577 gnd 0.011203f
C5777 commonsourceibias.n578 gnd 0.059802f
C5778 commonsourceibias.n579 gnd 0.011204f
C5779 commonsourceibias.n580 gnd 0.008022f
C5780 commonsourceibias.n581 gnd 0.008022f
C5781 commonsourceibias.n582 gnd 0.008022f
C5782 commonsourceibias.n583 gnd 0.009806f
C5783 commonsourceibias.n584 gnd 0.059802f
C5784 commonsourceibias.n585 gnd 0.010338f
C5785 commonsourceibias.t156 gnd 0.149881f
C5786 commonsourceibias.n586 gnd 0.059802f
C5787 commonsourceibias.n587 gnd 0.010488f
C5788 commonsourceibias.n588 gnd 0.008022f
C5789 commonsourceibias.n589 gnd 0.008022f
C5790 commonsourceibias.n590 gnd 0.008022f
C5791 commonsourceibias.n591 gnd 0.006995f
C5792 commonsourceibias.n592 gnd 0.011196f
C5793 commonsourceibias.n593 gnd 0.059802f
C5794 commonsourceibias.n594 gnd 0.0112f
C5795 commonsourceibias.n595 gnd 0.008022f
C5796 commonsourceibias.n596 gnd 0.008022f
C5797 commonsourceibias.n597 gnd 0.008022f
C5798 commonsourceibias.n598 gnd 0.009595f
C5799 commonsourceibias.n599 gnd 0.059802f
C5800 commonsourceibias.n600 gnd 0.010263f
C5801 commonsourceibias.t105 gnd 0.149881f
C5802 commonsourceibias.n601 gnd 0.059802f
C5803 commonsourceibias.n602 gnd 0.010563f
C5804 commonsourceibias.n603 gnd 0.008022f
C5805 commonsourceibias.n604 gnd 0.008022f
C5806 commonsourceibias.n605 gnd 0.008022f
C5807 commonsourceibias.n606 gnd 0.006855f
C5808 commonsourceibias.n607 gnd 0.011182f
C5809 commonsourceibias.n608 gnd 0.059802f
C5810 commonsourceibias.n609 gnd 0.01119f
C5811 commonsourceibias.n610 gnd 0.008022f
C5812 commonsourceibias.n611 gnd 0.008022f
C5813 commonsourceibias.n612 gnd 0.008022f
C5814 commonsourceibias.n613 gnd 0.00936f
C5815 commonsourceibias.n614 gnd 0.059802f
C5816 commonsourceibias.n615 gnd 0.009843f
C5817 commonsourceibias.n616 gnd 0.071758f
C5818 commonsourceibias.n617 gnd 0.046883f
C5819 commonsourceibias.n618 gnd 0.010705f
C5820 commonsourceibias.t141 gnd 0.149881f
C5821 commonsourceibias.n619 gnd 0.007808f
C5822 commonsourceibias.n620 gnd 0.008022f
C5823 commonsourceibias.t154 gnd 0.149881f
C5824 commonsourceibias.n621 gnd 0.010321f
C5825 commonsourceibias.n622 gnd 0.008022f
C5826 commonsourceibias.t132 gnd 0.149881f
C5827 commonsourceibias.n623 gnd 0.007564f
C5828 commonsourceibias.n624 gnd 0.008022f
C5829 commonsourceibias.t147 gnd 0.149881f
C5830 commonsourceibias.n625 gnd 0.010168f
C5831 commonsourceibias.n626 gnd 0.008022f
C5832 commonsourceibias.t123 gnd 0.149881f
C5833 commonsourceibias.n627 gnd 0.007348f
C5834 commonsourceibias.n628 gnd 0.008022f
C5835 commonsourceibias.t115 gnd 0.149881f
C5836 commonsourceibias.n629 gnd 0.009997f
C5837 commonsourceibias.n630 gnd 0.008022f
C5838 commonsourceibias.t88 gnd 0.149881f
C5839 commonsourceibias.n631 gnd 0.007159f
C5840 commonsourceibias.n632 gnd 0.008022f
C5841 commonsourceibias.t106 gnd 0.149881f
C5842 commonsourceibias.n633 gnd 0.009806f
C5843 commonsourceibias.n634 gnd 0.008022f
C5844 commonsourceibias.t143 gnd 0.149881f
C5845 commonsourceibias.n635 gnd 0.006995f
C5846 commonsourceibias.n636 gnd 0.008022f
C5847 commonsourceibias.t99 gnd 0.149881f
C5848 commonsourceibias.n637 gnd 0.009595f
C5849 commonsourceibias.n638 gnd 0.008022f
C5850 commonsourceibias.t136 gnd 0.149881f
C5851 commonsourceibias.n639 gnd 0.006855f
C5852 commonsourceibias.n640 gnd 0.008022f
C5853 commonsourceibias.t150 gnd 0.149881f
C5854 commonsourceibias.n641 gnd 0.00936f
C5855 commonsourceibias.t108 gnd 0.16664f
C5856 commonsourceibias.t158 gnd 0.149881f
C5857 commonsourceibias.n642 gnd 0.065328f
C5858 commonsourceibias.n643 gnd 0.07169f
C5859 commonsourceibias.n644 gnd 0.033265f
C5860 commonsourceibias.n645 gnd 0.008022f
C5861 commonsourceibias.n646 gnd 0.007808f
C5862 commonsourceibias.n647 gnd 0.01119f
C5863 commonsourceibias.n648 gnd 0.059802f
C5864 commonsourceibias.n649 gnd 0.011182f
C5865 commonsourceibias.n650 gnd 0.008022f
C5866 commonsourceibias.n651 gnd 0.008022f
C5867 commonsourceibias.n652 gnd 0.008022f
C5868 commonsourceibias.n653 gnd 0.010321f
C5869 commonsourceibias.n654 gnd 0.059802f
C5870 commonsourceibias.n655 gnd 0.010563f
C5871 commonsourceibias.t118 gnd 0.149881f
C5872 commonsourceibias.n656 gnd 0.059802f
C5873 commonsourceibias.n657 gnd 0.010263f
C5874 commonsourceibias.n658 gnd 0.008022f
C5875 commonsourceibias.n659 gnd 0.008022f
C5876 commonsourceibias.n660 gnd 0.008022f
C5877 commonsourceibias.n661 gnd 0.007564f
C5878 commonsourceibias.n662 gnd 0.0112f
C5879 commonsourceibias.n663 gnd 0.059802f
C5880 commonsourceibias.n664 gnd 0.011196f
C5881 commonsourceibias.n665 gnd 0.008022f
C5882 commonsourceibias.n666 gnd 0.008022f
C5883 commonsourceibias.n667 gnd 0.008022f
C5884 commonsourceibias.n668 gnd 0.010168f
C5885 commonsourceibias.n669 gnd 0.059802f
C5886 commonsourceibias.n670 gnd 0.010488f
C5887 commonsourceibias.t128 gnd 0.149881f
C5888 commonsourceibias.n671 gnd 0.059802f
C5889 commonsourceibias.n672 gnd 0.010338f
C5890 commonsourceibias.n673 gnd 0.008022f
C5891 commonsourceibias.n674 gnd 0.008022f
C5892 commonsourceibias.n675 gnd 0.008022f
C5893 commonsourceibias.n676 gnd 0.007348f
C5894 commonsourceibias.n677 gnd 0.011204f
C5895 commonsourceibias.n678 gnd 0.059802f
C5896 commonsourceibias.n679 gnd 0.011203f
C5897 commonsourceibias.n680 gnd 0.008022f
C5898 commonsourceibias.n681 gnd 0.008022f
C5899 commonsourceibias.n682 gnd 0.008022f
C5900 commonsourceibias.n683 gnd 0.009997f
C5901 commonsourceibias.n684 gnd 0.059802f
C5902 commonsourceibias.n685 gnd 0.010413f
C5903 commonsourceibias.t137 gnd 0.149881f
C5904 commonsourceibias.n686 gnd 0.059802f
C5905 commonsourceibias.n687 gnd 0.010413f
C5906 commonsourceibias.n688 gnd 0.008022f
C5907 commonsourceibias.n689 gnd 0.008022f
C5908 commonsourceibias.n690 gnd 0.008022f
C5909 commonsourceibias.n691 gnd 0.007159f
C5910 commonsourceibias.n692 gnd 0.011203f
C5911 commonsourceibias.n693 gnd 0.059802f
C5912 commonsourceibias.n694 gnd 0.011204f
C5913 commonsourceibias.n695 gnd 0.008022f
C5914 commonsourceibias.n696 gnd 0.008022f
C5915 commonsourceibias.n697 gnd 0.008022f
C5916 commonsourceibias.n698 gnd 0.009806f
C5917 commonsourceibias.n699 gnd 0.059802f
C5918 commonsourceibias.n700 gnd 0.010338f
C5919 commonsourceibias.t144 gnd 0.149881f
C5920 commonsourceibias.n701 gnd 0.059802f
C5921 commonsourceibias.n702 gnd 0.010488f
C5922 commonsourceibias.n703 gnd 0.008022f
C5923 commonsourceibias.n704 gnd 0.008022f
C5924 commonsourceibias.n705 gnd 0.008022f
C5925 commonsourceibias.n706 gnd 0.006995f
C5926 commonsourceibias.n707 gnd 0.011196f
C5927 commonsourceibias.n708 gnd 0.059802f
C5928 commonsourceibias.n709 gnd 0.0112f
C5929 commonsourceibias.n710 gnd 0.008022f
C5930 commonsourceibias.n711 gnd 0.008022f
C5931 commonsourceibias.n712 gnd 0.008022f
C5932 commonsourceibias.n713 gnd 0.009595f
C5933 commonsourceibias.n714 gnd 0.059802f
C5934 commonsourceibias.n715 gnd 0.010263f
C5935 commonsourceibias.t93 gnd 0.149881f
C5936 commonsourceibias.n716 gnd 0.059802f
C5937 commonsourceibias.n717 gnd 0.010563f
C5938 commonsourceibias.n718 gnd 0.008022f
C5939 commonsourceibias.n719 gnd 0.008022f
C5940 commonsourceibias.n720 gnd 0.008022f
C5941 commonsourceibias.n721 gnd 0.006855f
C5942 commonsourceibias.n722 gnd 0.011182f
C5943 commonsourceibias.n723 gnd 0.059802f
C5944 commonsourceibias.n724 gnd 0.01119f
C5945 commonsourceibias.n725 gnd 0.008022f
C5946 commonsourceibias.n726 gnd 0.008022f
C5947 commonsourceibias.n727 gnd 0.008022f
C5948 commonsourceibias.n728 gnd 0.00936f
C5949 commonsourceibias.n729 gnd 0.059802f
C5950 commonsourceibias.n730 gnd 0.009843f
C5951 commonsourceibias.t124 gnd 0.162096f
C5952 commonsourceibias.n731 gnd 0.071758f
C5953 commonsourceibias.n732 gnd 0.024957f
C5954 commonsourceibias.n733 gnd 0.221543f
C5955 commonsourceibias.n734 gnd 4.49224f
.ends

