* NGSPICE file created from opamp31.ext - technology: sky130A

.subckt opamp31 gnd CSoutput output vdd plus minus commonsourceibias outputibias diffpairibias
X0 a_n8300_8799.t44 plus.t5 a_n2903_n3924.t45 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X1 a_n2804_13878.t24 a_n2982_13878.t19 a_n2982_13878.t20 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X2 CSoutput.t167 commonsourceibias.t64 gnd.t118 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X3 a_n2804_13878.t25 a_n2982_13878.t72 vdd.t56 vdd.t55 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 gnd.t320 gnd.t318 gnd.t319 gnd.t271 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X5 CSoutput.t168 a_n2982_8322.t37 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X6 vdd.t155 a_n8300_8799.t48 CSoutput.t71 vdd.t119 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X7 gnd.t119 commonsourceibias.t65 CSoutput.t166 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 gnd.t317 gnd.t315 minus.t4 gnd.t316 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X9 CSoutput.t165 commonsourceibias.t66 gnd.t111 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X10 CSoutput.t164 commonsourceibias.t67 gnd.t112 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X11 CSoutput.t70 a_n8300_8799.t49 vdd.t154 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X12 a_n2903_n3924.t48 plus.t6 a_n8300_8799.t43 gnd.t49 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X13 a_n2903_n3924.t18 minus.t5 a_n2982_13878.t63 gnd.t97 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X14 a_n2982_8322.t23 a_n2982_13878.t73 a_n8300_8799.t17 vdd.t53 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X15 vdd.t0 CSoutput.t169 output.t19 gnd.t65 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X16 CSoutput.t69 a_n8300_8799.t50 vdd.t153 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X17 CSoutput.t163 commonsourceibias.t68 gnd.t353 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X18 gnd.t354 commonsourceibias.t69 CSoutput.t162 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 CSoutput.t161 commonsourceibias.t70 gnd.t175 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 gnd.t176 commonsourceibias.t71 CSoutput.t160 gnd.t36 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X21 vdd.t152 a_n8300_8799.t51 CSoutput.t68 vdd.t112 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X22 CSoutput.t159 commonsourceibias.t72 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X23 CSoutput.t158 commonsourceibias.t73 gnd.t21 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X24 gnd.t57 commonsourceibias.t74 CSoutput.t157 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X25 a_n2982_13878.t4 minus.t6 a_n2903_n3924.t4 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X26 commonsourceibias.t63 commonsourceibias.t62 gnd.t130 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X27 CSoutput.t156 commonsourceibias.t75 gnd.t59 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X28 a_n8300_8799.t12 a_n2982_13878.t74 a_n2982_8322.t22 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X29 vdd.t151 a_n8300_8799.t52 CSoutput.t67 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X30 a_n2982_13878.t10 minus.t7 a_n2903_n3924.t10 gnd.t64 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X31 vdd.t150 a_n8300_8799.t53 CSoutput.t66 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X32 a_n8300_8799.t0 a_n2982_13878.t75 a_n2982_8322.t21 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X33 CSoutput.t170 a_n2982_8322.t36 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X34 CSoutput.t155 commonsourceibias.t76 gnd.t148 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 gnd.t149 commonsourceibias.t77 CSoutput.t154 gnd.t120 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X36 gnd.t314 gnd.t312 gnd.t313 gnd.t235 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X37 CSoutput.t153 commonsourceibias.t78 gnd.t22 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X38 CSoutput.t152 commonsourceibias.t79 gnd.t24 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X39 a_n2903_n3924.t2 minus.t8 a_n2982_13878.t2 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X40 gnd.t311 gnd.t309 gnd.t310 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X41 CSoutput.t151 commonsourceibias.t80 gnd.t342 gnd.t109 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X42 a_n2903_n3924.t53 diffpairibias.t16 gnd.t335 gnd.t334 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X43 CSoutput.t65 a_n8300_8799.t54 vdd.t149 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X44 gnd.t343 commonsourceibias.t81 CSoutput.t150 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X45 vdd.t148 a_n8300_8799.t55 CSoutput.t64 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X46 CSoutput.t149 commonsourceibias.t82 gnd.t131 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X47 gnd.t93 commonsourceibias.t60 commonsourceibias.t61 gnd.t92 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X48 CSoutput.t148 commonsourceibias.t83 gnd.t132 gnd.t109 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X49 output.t2 outputibias.t8 gnd.t43 gnd.t42 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X50 gnd.t150 commonsourceibias.t84 CSoutput.t147 gnd.t115 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X51 a_n2903_n3924.t41 plus.t7 a_n8300_8799.t42 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X52 a_n2804_13878.t23 a_n2982_13878.t51 a_n2982_13878.t52 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X53 CSoutput.t146 commonsourceibias.t85 gnd.t152 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X54 gnd.t361 commonsourceibias.t86 CSoutput.t145 gnd.t115 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X55 vdd.t242 CSoutput.t171 output.t18 gnd.t325 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X56 a_n8300_8799.t41 plus.t8 a_n2903_n3924.t37 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X57 a_n2982_13878.t40 a_n2982_13878.t39 a_n2804_13878.t22 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X58 CSoutput.t144 commonsourceibias.t87 gnd.t362 gnd.t78 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X59 gnd.t344 commonsourceibias.t88 CSoutput.t143 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X60 a_n8300_8799.t40 plus.t9 a_n2903_n3924.t40 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X61 CSoutput.t63 a_n8300_8799.t56 vdd.t147 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X62 vdd.t235 vdd.t233 vdd.t234 vdd.t210 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X63 gnd.t87 commonsourceibias.t58 commonsourceibias.t59 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X64 CSoutput.t142 commonsourceibias.t89 gnd.t345 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X65 gnd.t308 gnd.t305 gnd.t307 gnd.t306 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X66 vdd.t146 a_n8300_8799.t57 CSoutput.t62 vdd.t112 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X67 gnd.t304 gnd.t302 gnd.t303 gnd.t235 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X68 CSoutput.t141 commonsourceibias.t90 gnd.t153 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X69 diffpairibias.t15 diffpairibias.t14 gnd.t108 gnd.t107 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X70 a_n2903_n3924.t33 plus.t10 a_n8300_8799.t39 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X71 a_n2982_13878.t0 minus.t9 a_n2903_n3924.t0 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X72 a_n2982_13878.t36 a_n2982_13878.t35 a_n2804_13878.t21 vdd.t38 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X73 CSoutput.t140 commonsourceibias.t91 gnd.t154 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X74 CSoutput.t139 commonsourceibias.t92 gnd.t363 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X75 gnd.t364 commonsourceibias.t93 CSoutput.t138 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X76 gnd.t346 commonsourceibias.t94 CSoutput.t137 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X77 a_n8300_8799.t15 a_n2982_13878.t76 a_n2982_8322.t20 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X78 CSoutput.t61 a_n8300_8799.t58 vdd.t145 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X79 gnd.t347 commonsourceibias.t95 CSoutput.t136 gnd.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 gnd.t301 gnd.t299 plus.t3 gnd.t300 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X81 a_n2982_13878.t58 a_n2982_13878.t57 a_n2804_13878.t20 vdd.t54 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X82 vdd.t144 a_n8300_8799.t59 CSoutput.t60 vdd.t74 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 vdd.t143 a_n8300_8799.t60 CSoutput.t59 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X84 a_n8300_8799.t19 a_n2982_13878.t77 a_n2982_8322.t19 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X85 CSoutput.t135 commonsourceibias.t96 gnd.t53 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X86 diffpairibias.t13 diffpairibias.t12 gnd.t103 gnd.t102 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X87 CSoutput.t58 a_n8300_8799.t61 vdd.t142 vdd.t77 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X88 gnd.t174 commonsourceibias.t56 commonsourceibias.t57 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 gnd.t366 commonsourceibias.t97 CSoutput.t134 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X90 CSoutput.t133 commonsourceibias.t98 gnd.t177 gnd.t78 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 a_n8300_8799.t20 a_n2982_13878.t78 a_n2982_8322.t18 vdd.t46 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X92 gnd.t26 commonsourceibias.t99 CSoutput.t132 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X93 gnd.t298 gnd.t296 gnd.t297 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X94 CSoutput.t131 commonsourceibias.t100 gnd.t333 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X95 CSoutput.t130 commonsourceibias.t101 gnd.t133 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X96 a_n2982_8322.t17 a_n2982_13878.t79 a_n8300_8799.t46 vdd.t54 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X97 gnd.t126 commonsourceibias.t102 CSoutput.t129 gnd.t120 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X98 vdd.t232 vdd.t230 vdd.t231 vdd.t197 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X99 CSoutput.t57 a_n8300_8799.t62 vdd.t141 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X100 CSoutput.t172 a_n2982_8322.t35 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X101 gnd.t76 commonsourceibias.t54 commonsourceibias.t55 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X102 gnd.t295 gnd.t293 gnd.t294 gnd.t224 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X103 gnd.t292 gnd.t290 plus.t2 gnd.t291 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X104 output.t17 CSoutput.t173 vdd.t243 gnd.t326 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X105 a_n2903_n3924.t29 plus.t11 a_n8300_8799.t38 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X106 gnd.t60 commonsourceibias.t103 CSoutput.t128 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X107 a_n2903_n3924.t11 diffpairibias.t17 gnd.t69 gnd.t68 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X108 vdd.t140 a_n8300_8799.t63 CSoutput.t56 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X109 gnd.t289 gnd.t287 gnd.t288 gnd.t213 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X110 vdd.t139 a_n8300_8799.t64 CSoutput.t55 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X111 a_n2982_13878.t42 a_n2982_13878.t41 a_n2804_13878.t19 vdd.t53 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X112 vdd.t138 a_n8300_8799.t65 CSoutput.t54 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X113 gnd.t28 commonsourceibias.t104 CSoutput.t127 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X114 a_n8300_8799.t2 a_n2982_13878.t80 a_n2982_8322.t16 vdd.t42 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X115 a_n2982_13878.t24 a_n2982_13878.t23 a_n2804_13878.t18 vdd.t5 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X116 gnd.t286 gnd.t284 gnd.t285 gnd.t213 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X117 CSoutput.t126 commonsourceibias.t105 gnd.t29 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X118 gnd.t89 commonsourceibias.t106 CSoutput.t125 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X119 a_n2982_13878.t62 minus.t10 a_n2903_n3924.t17 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X120 output.t16 CSoutput.t174 vdd.t156 gnd.t98 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X121 vdd.t229 vdd.t227 vdd.t228 vdd.t217 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X122 gnd.t159 commonsourceibias.t52 commonsourceibias.t53 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X123 gnd.t367 commonsourceibias.t107 CSoutput.t124 gnd.t92 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X124 CSoutput.t53 a_n8300_8799.t66 vdd.t137 vdd.t77 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X125 vdd.t226 vdd.t223 vdd.t225 vdd.t224 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X126 output.t0 outputibias.t9 gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X127 a_n2804_13878.t17 a_n2982_13878.t45 a_n2982_13878.t46 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X128 a_n2903_n3924.t16 minus.t11 a_n2982_13878.t61 gnd.t95 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X129 CSoutput.t52 a_n8300_8799.t67 vdd.t136 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X130 CSoutput.t175 a_n2982_8322.t34 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X131 vdd.t135 a_n8300_8799.t68 CSoutput.t51 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X132 vdd.t52 a_n2982_13878.t81 a_n2982_8322.t31 vdd.t51 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X133 a_n2982_13878.t56 a_n2982_13878.t55 a_n2804_13878.t16 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X134 vdd.t222 vdd.t220 vdd.t221 vdd.t197 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X135 a_n2982_8322.t30 a_n2982_13878.t82 vdd.t50 vdd.t49 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X136 gnd.t94 commonsourceibias.t108 CSoutput.t123 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X137 a_n2903_n3924.t15 diffpairibias.t18 gnd.t91 gnd.t90 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X138 output.t15 CSoutput.t176 vdd.t157 gnd.t99 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X139 CSoutput.t50 a_n8300_8799.t69 vdd.t134 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X140 vdd.t158 CSoutput.t177 output.t14 gnd.t100 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X141 gnd.t180 commonsourceibias.t109 CSoutput.t122 gnd.t115 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X142 gnd.t193 commonsourceibias.t50 commonsourceibias.t51 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X143 CSoutput.t121 commonsourceibias.t110 gnd.t336 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X144 gnd.t113 commonsourceibias.t111 CSoutput.t120 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X145 CSoutput.t119 commonsourceibias.t112 gnd.t355 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X146 CSoutput.t118 commonsourceibias.t113 gnd.t55 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X147 a_n2903_n3924.t12 minus.t12 a_n2982_13878.t59 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X148 a_n2903_n3924.t1 minus.t13 a_n2982_13878.t1 gnd.t8 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X149 CSoutput.t178 a_n2982_8322.t33 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X150 vdd.t48 a_n2982_13878.t83 a_n2804_13878.t28 vdd.t47 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X151 a_n2982_13878.t7 minus.t14 a_n2903_n3924.t7 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X152 a_n2903_n3924.t34 plus.t12 a_n8300_8799.t37 gnd.t324 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X153 a_n2903_n3924.t36 plus.t13 a_n8300_8799.t36 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X154 vdd.t219 vdd.t216 vdd.t218 vdd.t217 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X155 a_n2982_13878.t6 minus.t15 a_n2903_n3924.t6 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X156 gnd.t283 gnd.t281 gnd.t282 gnd.t213 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X157 a_n2804_13878.t15 a_n2982_13878.t37 a_n2982_13878.t38 vdd.t46 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X158 vdd.t133 a_n8300_8799.t70 CSoutput.t49 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X159 vdd.t131 a_n8300_8799.t71 CSoutput.t48 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X160 a_n2982_8322.t15 a_n2982_13878.t84 a_n8300_8799.t16 vdd.t32 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X161 gnd.t280 gnd.t278 plus.t1 gnd.t279 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X162 a_n8300_8799.t35 plus.t14 a_n2903_n3924.t31 gnd.t323 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X163 a_n8300_8799.t34 plus.t15 a_n2903_n3924.t42 gnd.t164 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X164 vdd.t215 vdd.t213 vdd.t214 vdd.t179 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X165 vdd.t212 vdd.t209 vdd.t211 vdd.t210 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X166 a_n2982_8322.t29 a_n2982_13878.t85 vdd.t45 vdd.t44 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X167 a_n8300_8799.t13 a_n2982_13878.t86 a_n2982_8322.t14 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X168 CSoutput.t47 a_n8300_8799.t72 vdd.t130 vdd.t85 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X169 diffpairibias.t11 diffpairibias.t10 gnd.t71 gnd.t70 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X170 vdd.t129 a_n8300_8799.t73 CSoutput.t46 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X171 a_n2982_13878.t68 minus.t16 a_n2903_n3924.t26 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X172 a_n2982_13878.t26 a_n2982_13878.t25 a_n2804_13878.t14 vdd.t26 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X173 CSoutput.t117 commonsourceibias.t114 gnd.t196 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X174 a_n8300_8799.t11 a_n2982_13878.t87 a_n2982_8322.t13 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X175 commonsourceibias.t49 commonsourceibias.t48 gnd.t341 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X176 output.t13 CSoutput.t179 vdd.t159 gnd.t101 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X177 gnd.t160 commonsourceibias.t115 CSoutput.t116 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X178 a_n2804_13878.t13 a_n2982_13878.t53 a_n2982_13878.t54 vdd.t42 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X179 a_n2903_n3924.t3 minus.t17 a_n2982_13878.t3 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X180 gnd.t277 gnd.t274 gnd.t276 gnd.t275 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X181 CSoutput.t115 commonsourceibias.t116 gnd.t77 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X182 vdd.t208 vdd.t206 vdd.t207 vdd.t165 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X183 output.t12 CSoutput.t180 vdd.t57 gnd.t72 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X184 CSoutput.t45 a_n8300_8799.t74 vdd.t127 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X185 gnd.t273 gnd.t270 gnd.t272 gnd.t271 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X186 CSoutput.t114 commonsourceibias.t117 gnd.t327 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X187 gnd.t269 gnd.t267 gnd.t268 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X188 vdd.t41 a_n2982_13878.t88 a_n2982_8322.t28 vdd.t40 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X189 a_n2804_13878.t12 a_n2982_13878.t13 a_n2982_13878.t14 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X190 outputibias.t7 outputibias.t6 gnd.t179 gnd.t178 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X191 vdd.t126 a_n8300_8799.t75 CSoutput.t44 vdd.t119 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X192 a_n2982_13878.t44 a_n2982_13878.t43 a_n2804_13878.t11 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X193 gnd.t329 commonsourceibias.t118 CSoutput.t113 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X194 gnd.t121 commonsourceibias.t119 CSoutput.t112 gnd.t120 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X195 commonsourceibias.t47 commonsourceibias.t46 gnd.t360 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 minus.t3 gnd.t264 gnd.t266 gnd.t265 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X197 gnd.t166 commonsourceibias.t120 CSoutput.t111 gnd.t36 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X198 outputibias.t5 outputibias.t4 gnd.t10 gnd.t9 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X199 a_n2903_n3924.t32 plus.t16 a_n8300_8799.t33 gnd.t97 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X200 vdd.t125 a_n8300_8799.t76 CSoutput.t43 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X201 CSoutput.t110 commonsourceibias.t121 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X202 a_n2903_n3924.t14 diffpairibias.t19 gnd.t86 gnd.t85 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X203 gnd.t263 gnd.t260 gnd.t262 gnd.t261 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X204 a_n2903_n3924.t24 diffpairibias.t20 gnd.t173 gnd.t172 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X205 commonsourceibias.t45 commonsourceibias.t44 gnd.t145 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X206 vdd.t124 a_n8300_8799.t77 CSoutput.t42 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X207 a_n8300_8799.t32 plus.t17 a_n2903_n3924.t30 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X208 gnd.t259 gnd.t257 gnd.t258 gnd.t235 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X209 gnd.t256 gnd.t254 gnd.t255 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X210 vdd.t205 vdd.t203 vdd.t204 vdd.t179 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X211 vdd.t58 CSoutput.t181 output.t11 gnd.t73 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X212 CSoutput.t109 commonsourceibias.t122 gnd.t31 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X213 CSoutput.t108 commonsourceibias.t123 gnd.t167 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X214 a_n2804_13878.t10 a_n2982_13878.t29 a_n2982_13878.t30 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X215 a_n2982_8322.t12 a_n2982_13878.t89 a_n8300_8799.t5 vdd.t38 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X216 CSoutput.t41 a_n8300_8799.t78 vdd.t123 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X217 commonsourceibias.t43 commonsourceibias.t42 gnd.t110 gnd.t109 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X218 gnd.t116 commonsourceibias.t40 commonsourceibias.t41 gnd.t115 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X219 vdd.t59 CSoutput.t182 output.t10 gnd.t74 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X220 diffpairibias.t9 diffpairibias.t8 gnd.t67 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X221 a_n2804_13878.t29 a_n2982_13878.t90 vdd.t37 vdd.t36 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X222 vdd.t35 a_n2982_13878.t91 a_n2804_13878.t0 vdd.t34 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X223 CSoutput.t107 commonsourceibias.t124 gnd.t197 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X224 CSoutput.t106 commonsourceibias.t125 gnd.t155 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X225 CSoutput.t40 a_n8300_8799.t79 vdd.t122 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X226 gnd.t63 commonsourceibias.t38 commonsourceibias.t39 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X227 vdd.t120 a_n8300_8799.t80 CSoutput.t39 vdd.t119 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X228 vdd.t118 a_n8300_8799.t81 CSoutput.t38 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X229 commonsourceibias.t37 commonsourceibias.t36 gnd.t340 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X230 outputibias.t3 outputibias.t2 gnd.t137 gnd.t136 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X231 CSoutput.t37 a_n8300_8799.t82 vdd.t116 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X232 plus.t4 gnd.t251 gnd.t253 gnd.t252 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X233 a_n2804_13878.t9 a_n2982_13878.t15 a_n2982_13878.t16 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X234 a_n2903_n3924.t25 minus.t18 a_n2982_13878.t67 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X235 gnd.t161 commonsourceibias.t126 CSoutput.t105 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X236 commonsourceibias.t35 commonsourceibias.t34 gnd.t15 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X237 vdd.t115 a_n8300_8799.t83 CSoutput.t36 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X238 a_n2982_13878.t60 minus.t19 a_n2903_n3924.t13 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X239 gnd.t144 commonsourceibias.t32 commonsourceibias.t33 gnd.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X240 a_n2982_8322.t11 a_n2982_13878.t92 a_n8300_8799.t9 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X241 a_n2982_13878.t22 a_n2982_13878.t21 a_n2804_13878.t8 vdd.t32 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X242 CSoutput.t104 commonsourceibias.t127 gnd.t79 gnd.t78 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X243 CSoutput.t35 a_n8300_8799.t84 vdd.t114 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X244 diffpairibias.t7 diffpairibias.t6 gnd.t17 gnd.t16 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X245 vdd.t113 a_n8300_8799.t85 CSoutput.t34 vdd.t112 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X246 a_n2804_13878.t7 a_n2982_13878.t27 a_n2982_13878.t28 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X247 commonsourceibias.t31 commonsourceibias.t30 gnd.t185 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X248 a_n2982_13878.t64 minus.t20 a_n2903_n3924.t20 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X249 a_n2982_13878.t69 minus.t21 a_n2903_n3924.t27 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X250 vdd.t202 vdd.t200 vdd.t201 vdd.t183 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X251 vdd.t30 a_n2982_13878.t93 a_n2982_8322.t27 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X252 vdd.t111 a_n8300_8799.t86 CSoutput.t33 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X253 a_n2903_n3924.t23 minus.t22 a_n2982_13878.t66 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X254 a_n8300_8799.t31 plus.t18 a_n2903_n3924.t39 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X255 gnd.t33 commonsourceibias.t128 CSoutput.t103 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X256 a_n2903_n3924.t8 minus.t23 a_n2982_13878.t8 gnd.t49 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X257 CSoutput.t32 a_n8300_8799.t87 vdd.t109 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X258 gnd.t171 commonsourceibias.t28 commonsourceibias.t29 gnd.t120 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X259 CSoutput.t102 commonsourceibias.t129 gnd.t328 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X260 a_n2804_13878.t26 a_n2982_13878.t94 vdd.t28 vdd.t27 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X261 vdd.t199 vdd.t196 vdd.t198 vdd.t197 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X262 vdd.t195 vdd.t193 vdd.t194 vdd.t183 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X263 output.t9 CSoutput.t183 vdd.t239 gnd.t190 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X264 CSoutput.t31 a_n8300_8799.t88 vdd.t108 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X265 gnd.t250 gnd.t248 minus.t2 gnd.t249 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X266 gnd.t330 commonsourceibias.t130 CSoutput.t101 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X267 gnd.t247 gnd.t244 gnd.t246 gnd.t245 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X268 vdd.t192 vdd.t190 vdd.t191 vdd.t169 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X269 vdd.t107 a_n8300_8799.t89 CSoutput.t30 vdd.t94 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X270 a_n2903_n3924.t55 diffpairibias.t21 gnd.t352 gnd.t351 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X271 a_n2982_8322.t10 a_n2982_13878.t95 a_n8300_8799.t3 vdd.t26 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X272 vdd.t25 a_n2982_13878.t96 a_n2982_8322.t26 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X273 gnd.t339 commonsourceibias.t26 commonsourceibias.t27 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X274 a_n8300_8799.t30 plus.t19 a_n2903_n3924.t28 gnd.t64 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X275 output.t1 outputibias.t10 gnd.t41 gnd.t40 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X276 gnd.t243 gnd.t241 gnd.t242 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X277 gnd.t359 commonsourceibias.t24 commonsourceibias.t25 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 vdd.t189 vdd.t186 vdd.t188 vdd.t187 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X279 gnd.t240 gnd.t238 gnd.t239 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X280 CSoutput.t100 commonsourceibias.t131 gnd.t134 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X281 a_n2903_n3924.t50 plus.t20 a_n8300_8799.t29 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X282 vdd.t106 a_n8300_8799.t90 CSoutput.t29 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X283 vdd.t240 CSoutput.t184 output.t8 gnd.t191 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X284 CSoutput.t28 a_n8300_8799.t91 vdd.t105 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X285 CSoutput.t99 commonsourceibias.t132 gnd.t122 gnd.t109 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X286 output.t3 outputibias.t11 gnd.t182 gnd.t181 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X287 a_n2804_13878.t6 a_n2982_13878.t31 a_n2982_13878.t32 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X288 CSoutput.t27 a_n8300_8799.t92 vdd.t101 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X289 a_n2982_8322.t9 a_n2982_13878.t97 a_n8300_8799.t8 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X290 vdd.t185 vdd.t182 vdd.t184 vdd.t183 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X291 diffpairibias.t5 diffpairibias.t4 gnd.t195 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X292 gnd.t237 gnd.t234 gnd.t236 gnd.t235 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X293 CSoutput.t26 a_n8300_8799.t93 vdd.t103 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X294 CSoutput.t25 a_n8300_8799.t94 vdd.t100 vdd.t85 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X295 gnd.t143 commonsourceibias.t22 commonsourceibias.t23 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X296 output.t7 CSoutput.t185 vdd.t241 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X297 vdd.t181 vdd.t178 vdd.t180 vdd.t179 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X298 CSoutput.t98 commonsourceibias.t133 gnd.t356 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X299 a_n2982_8322.t25 a_n2982_13878.t98 vdd.t22 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X300 CSoutput.t24 a_n8300_8799.t95 vdd.t99 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X301 vdd.t95 a_n8300_8799.t96 CSoutput.t23 vdd.t94 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X302 gnd.t348 commonsourceibias.t134 CSoutput.t97 gnd.t92 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X303 CSoutput.t22 a_n8300_8799.t97 vdd.t97 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X304 vdd.t20 a_n2982_13878.t99 a_n2804_13878.t31 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X305 plus.t0 gnd.t231 gnd.t233 gnd.t232 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X306 vdd.t96 a_n8300_8799.t98 CSoutput.t21 vdd.t94 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X307 CSoutput.t20 a_n8300_8799.t99 vdd.t93 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X308 a_n2903_n3924.t47 plus.t21 a_n8300_8799.t28 gnd.t8 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X309 gnd.t139 commonsourceibias.t135 CSoutput.t96 gnd.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X310 gnd.t35 commonsourceibias.t136 CSoutput.t95 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X311 output.t6 CSoutput.t186 vdd.t236 gnd.t187 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X312 a_n2903_n3924.t52 minus.t24 a_n2982_13878.t70 gnd.t324 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X313 a_n2982_8322.t8 a_n2982_13878.t100 a_n8300_8799.t45 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X314 commonsourceibias.t21 commonsourceibias.t20 gnd.t104 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X315 vdd.t237 CSoutput.t187 output.t5 gnd.t188 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X316 a_n8300_8799.t10 a_n2982_13878.t101 a_n2982_8322.t7 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X317 a_n8300_8799.t27 plus.t22 a_n2903_n3924.t46 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X318 a_n2804_13878.t30 a_n2982_13878.t102 vdd.t17 vdd.t16 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X319 gnd.t168 commonsourceibias.t137 CSoutput.t94 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X320 vdd.t177 vdd.t175 vdd.t176 vdd.t161 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X321 vdd.t91 a_n8300_8799.t100 CSoutput.t19 vdd.t74 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X322 a_n2982_13878.t71 minus.t25 a_n2903_n3924.t54 gnd.t323 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X323 CSoutput.t18 a_n8300_8799.t101 vdd.t90 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X324 commonsourceibias.t19 commonsourceibias.t18 gnd.t114 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X325 a_n2982_13878.t12 a_n2982_13878.t11 a_n2804_13878.t5 vdd.t6 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X326 a_n8300_8799.t1 a_n2982_13878.t103 a_n2982_8322.t6 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X327 gnd.t230 gnd.t227 gnd.t229 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X328 a_n8300_8799.t4 a_n2982_13878.t104 a_n2982_8322.t5 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X329 gnd.t156 commonsourceibias.t138 CSoutput.t93 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 commonsourceibias.t17 commonsourceibias.t16 gnd.t338 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X331 a_n8300_8799.t26 plus.t23 a_n2903_n3924.t49 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X332 gnd.t226 gnd.t223 gnd.t225 gnd.t224 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X333 gnd.t222 gnd.t220 minus.t1 gnd.t221 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X334 a_n2982_8322.t4 a_n2982_13878.t105 a_n8300_8799.t18 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X335 gnd.t365 commonsourceibias.t139 CSoutput.t92 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X336 CSoutput.t91 commonsourceibias.t140 gnd.t349 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X337 a_n2903_n3924.t9 minus.t26 a_n2982_13878.t9 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X338 vdd.t88 a_n8300_8799.t102 CSoutput.t17 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X339 gnd.t13 commonsourceibias.t14 commonsourceibias.t15 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X340 CSoutput.t16 a_n8300_8799.t103 vdd.t86 vdd.t85 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X341 CSoutput.t15 a_n8300_8799.t104 vdd.t84 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X342 CSoutput.t14 a_n8300_8799.t105 vdd.t83 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X343 gnd.t219 gnd.t216 gnd.t218 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X344 a_n2804_13878.t4 a_n2982_13878.t49 a_n2982_13878.t50 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X345 a_n2903_n3924.t43 plus.t24 a_n8300_8799.t25 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X346 vdd.t82 a_n8300_8799.t106 CSoutput.t13 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X347 gnd.t142 commonsourceibias.t12 commonsourceibias.t13 gnd.t36 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X348 commonsourceibias.t11 commonsourceibias.t10 gnd.t184 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X349 gnd.t198 commonsourceibias.t141 CSoutput.t90 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X350 a_n2903_n3924.t19 diffpairibias.t22 gnd.t106 gnd.t105 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X351 gnd.t162 commonsourceibias.t142 CSoutput.t89 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X352 CSoutput.t88 commonsourceibias.t143 gnd.t80 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X353 vdd.t81 a_n8300_8799.t107 CSoutput.t12 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X354 gnd.t331 commonsourceibias.t144 CSoutput.t87 gnd.t92 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X355 CSoutput.t11 a_n8300_8799.t108 vdd.t80 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X356 CSoutput.t86 commonsourceibias.t145 gnd.t169 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X357 a_n2982_13878.t18 a_n2982_13878.t17 a_n2804_13878.t3 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X358 gnd.t215 gnd.t212 gnd.t214 gnd.t213 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X359 a_n8300_8799.t7 a_n2982_13878.t106 a_n2982_8322.t3 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X360 vdd.t238 CSoutput.t188 output.t4 gnd.t189 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X361 vdd.t79 a_n8300_8799.t109 CSoutput.t10 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X362 CSoutput.t9 a_n8300_8799.t110 vdd.t78 vdd.t77 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X363 a_n8300_8799.t24 plus.t25 a_n2903_n3924.t38 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X364 vdd.t174 vdd.t172 vdd.t173 vdd.t169 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X365 CSoutput.t85 commonsourceibias.t146 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X366 gnd.t37 commonsourceibias.t147 CSoutput.t84 gnd.t36 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X367 commonsourceibias.t9 commonsourceibias.t8 gnd.t51 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X368 diffpairibias.t3 diffpairibias.t2 gnd.t322 gnd.t321 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X369 CSoutput.t8 a_n8300_8799.t111 vdd.t76 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X370 CSoutput.t189 a_n2982_8322.t32 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X371 a_n2982_8322.t2 a_n2982_13878.t107 a_n8300_8799.t6 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X372 gnd.t170 commonsourceibias.t148 CSoutput.t83 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X373 a_n2903_n3924.t44 plus.t26 a_n8300_8799.t23 gnd.t95 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X374 vdd.t75 a_n8300_8799.t112 CSoutput.t7 vdd.t74 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X375 gnd.t211 gnd.t208 gnd.t210 gnd.t209 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X376 CSoutput.t6 a_n8300_8799.t113 vdd.t73 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X377 diffpairibias.t1 diffpairibias.t0 gnd.t147 gnd.t146 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X378 gnd.t199 commonsourceibias.t149 CSoutput.t82 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X379 commonsourceibias.t7 commonsourceibias.t6 gnd.t7 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X380 gnd.t157 commonsourceibias.t150 CSoutput.t81 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X381 a_n2903_n3924.t51 plus.t27 a_n8300_8799.t22 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X382 CSoutput.t80 commonsourceibias.t151 gnd.t163 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X383 vdd.t8 a_n2982_13878.t108 a_n2804_13878.t27 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X384 a_n8300_8799.t21 plus.t28 a_n2903_n3924.t35 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X385 CSoutput.t5 a_n8300_8799.t114 vdd.t71 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X386 a_n2903_n3924.t5 minus.t27 a_n2982_13878.t5 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X387 vdd.t69 a_n8300_8799.t115 CSoutput.t4 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X388 gnd.t337 commonsourceibias.t4 commonsourceibias.t5 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X389 gnd.t82 commonsourceibias.t152 CSoutput.t79 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X390 a_n2982_8322.t1 a_n2982_13878.t109 a_n8300_8799.t14 vdd.t6 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X391 a_n2982_13878.t65 minus.t28 a_n2903_n3924.t22 gnd.t164 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X392 commonsourceibias.t3 commonsourceibias.t2 gnd.t358 gnd.t78 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X393 gnd.t39 commonsourceibias.t153 CSoutput.t78 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X394 gnd.t207 gnd.t204 gnd.t206 gnd.t205 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X395 gnd.t332 commonsourceibias.t154 CSoutput.t77 gnd.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X396 a_n2982_8322.t0 a_n2982_13878.t110 a_n8300_8799.t47 vdd.t5 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X397 vdd.t67 a_n8300_8799.t116 CSoutput.t3 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X398 vdd.t65 a_n8300_8799.t117 CSoutput.t2 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X399 CSoutput.t1 a_n8300_8799.t118 vdd.t63 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X400 gnd.t135 commonsourceibias.t155 CSoutput.t76 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X401 vdd.t171 vdd.t168 vdd.t170 vdd.t169 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X402 a_n2982_8322.t24 a_n2982_13878.t111 vdd.t4 vdd.t3 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X403 gnd.t123 commonsourceibias.t156 CSoutput.t75 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X404 a_n2804_13878.t2 a_n2982_13878.t33 a_n2982_13878.t34 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X405 gnd.t357 commonsourceibias.t157 CSoutput.t74 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X406 CSoutput.t73 commonsourceibias.t158 gnd.t350 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X407 commonsourceibias.t1 commonsourceibias.t0 gnd.t141 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X408 CSoutput.t72 commonsourceibias.t159 gnd.t158 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X409 minus.t0 gnd.t201 gnd.t203 gnd.t202 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X410 outputibias.t1 outputibias.t0 gnd.t125 gnd.t124 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X411 vdd.t167 vdd.t164 vdd.t166 vdd.t165 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X412 a_n2903_n3924.t21 diffpairibias.t23 gnd.t128 gnd.t127 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X413 vdd.t163 vdd.t160 vdd.t162 vdd.t161 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X414 CSoutput.t0 a_n8300_8799.t119 vdd.t61 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X415 a_n2982_13878.t48 a_n2982_13878.t47 a_n2804_13878.t1 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 plus.n53 plus.t20 323.478
R1 plus.n11 plus.t15 323.478
R2 plus.n52 plus.t19 297.12
R3 plus.n56 plus.t26 297.12
R4 plus.n58 plus.t25 297.12
R5 plus.n62 plus.t27 297.12
R6 plus.n64 plus.t9 297.12
R7 plus.n68 plus.t7 297.12
R8 plus.n70 plus.t14 297.12
R9 plus.n74 plus.t12 297.12
R10 plus.n76 plus.t28 297.12
R11 plus.n80 plus.t10 297.12
R12 plus.n82 plus.t8 297.12
R13 plus.n40 plus.t21 297.12
R14 plus.n38 plus.t22 297.12
R15 plus.n2 plus.t16 297.12
R16 plus.n32 plus.t17 297.12
R17 plus.n4 plus.t11 297.12
R18 plus.n26 plus.t5 297.12
R19 plus.n6 plus.t6 297.12
R20 plus.n20 plus.t23 297.12
R21 plus.n8 plus.t24 297.12
R22 plus.n14 plus.t18 297.12
R23 plus.n10 plus.t13 297.12
R24 plus.n86 plus.t1 243.97
R25 plus.n86 plus.n85 223.454
R26 plus.n88 plus.n87 223.454
R27 plus.n83 plus.n82 161.3
R28 plus.n81 plus.n42 161.3
R29 plus.n80 plus.n79 161.3
R30 plus.n78 plus.n43 161.3
R31 plus.n77 plus.n76 161.3
R32 plus.n75 plus.n44 161.3
R33 plus.n74 plus.n73 161.3
R34 plus.n72 plus.n45 161.3
R35 plus.n71 plus.n70 161.3
R36 plus.n69 plus.n46 161.3
R37 plus.n68 plus.n67 161.3
R38 plus.n66 plus.n47 161.3
R39 plus.n65 plus.n64 161.3
R40 plus.n63 plus.n48 161.3
R41 plus.n62 plus.n61 161.3
R42 plus.n60 plus.n49 161.3
R43 plus.n59 plus.n58 161.3
R44 plus.n57 plus.n50 161.3
R45 plus.n56 plus.n55 161.3
R46 plus.n54 plus.n51 161.3
R47 plus.n13 plus.n12 161.3
R48 plus.n14 plus.n9 161.3
R49 plus.n16 plus.n15 161.3
R50 plus.n17 plus.n8 161.3
R51 plus.n19 plus.n18 161.3
R52 plus.n20 plus.n7 161.3
R53 plus.n22 plus.n21 161.3
R54 plus.n23 plus.n6 161.3
R55 plus.n25 plus.n24 161.3
R56 plus.n26 plus.n5 161.3
R57 plus.n28 plus.n27 161.3
R58 plus.n29 plus.n4 161.3
R59 plus.n31 plus.n30 161.3
R60 plus.n32 plus.n3 161.3
R61 plus.n34 plus.n33 161.3
R62 plus.n35 plus.n2 161.3
R63 plus.n37 plus.n36 161.3
R64 plus.n38 plus.n1 161.3
R65 plus.n39 plus.n0 161.3
R66 plus.n41 plus.n40 161.3
R67 plus.n82 plus.n81 46.0096
R68 plus.n40 plus.n39 46.0096
R69 plus.n54 plus.n53 45.0871
R70 plus.n12 plus.n11 45.0871
R71 plus.n52 plus.n51 41.6278
R72 plus.n80 plus.n43 41.6278
R73 plus.n38 plus.n37 41.6278
R74 plus.n13 plus.n10 41.6278
R75 plus.n57 plus.n56 37.246
R76 plus.n76 plus.n75 37.246
R77 plus.n33 plus.n2 37.246
R78 plus.n15 plus.n14 37.246
R79 plus.n84 plus.n83 33.1766
R80 plus.n58 plus.n49 32.8641
R81 plus.n74 plus.n45 32.8641
R82 plus.n32 plus.n31 32.8641
R83 plus.n19 plus.n8 32.8641
R84 plus.n63 plus.n62 28.4823
R85 plus.n70 plus.n69 28.4823
R86 plus.n27 plus.n4 28.4823
R87 plus.n21 plus.n20 28.4823
R88 plus.n64 plus.n47 24.1005
R89 plus.n68 plus.n47 24.1005
R90 plus.n26 plus.n25 24.1005
R91 plus.n25 plus.n6 24.1005
R92 plus.n85 plus.t2 19.8005
R93 plus.n85 plus.t4 19.8005
R94 plus.n87 plus.t3 19.8005
R95 plus.n87 plus.t0 19.8005
R96 plus.n64 plus.n63 19.7187
R97 plus.n69 plus.n68 19.7187
R98 plus.n27 plus.n26 19.7187
R99 plus.n21 plus.n6 19.7187
R100 plus.n62 plus.n49 15.3369
R101 plus.n70 plus.n45 15.3369
R102 plus.n31 plus.n4 15.3369
R103 plus.n20 plus.n19 15.3369
R104 plus plus.n89 14.5734
R105 plus.n53 plus.n52 14.1472
R106 plus.n11 plus.n10 14.1472
R107 plus.n84 plus.n41 11.8774
R108 plus.n58 plus.n57 10.955
R109 plus.n75 plus.n74 10.955
R110 plus.n33 plus.n32 10.955
R111 plus.n15 plus.n8 10.955
R112 plus.n56 plus.n51 6.57323
R113 plus.n76 plus.n43 6.57323
R114 plus.n37 plus.n2 6.57323
R115 plus.n14 plus.n13 6.57323
R116 plus.n89 plus.n88 5.40567
R117 plus.n81 plus.n80 2.19141
R118 plus.n39 plus.n38 2.19141
R119 plus.n89 plus.n84 1.188
R120 plus.n88 plus.n86 0.716017
R121 plus.n55 plus.n54 0.189894
R122 plus.n55 plus.n50 0.189894
R123 plus.n59 plus.n50 0.189894
R124 plus.n60 plus.n59 0.189894
R125 plus.n61 plus.n60 0.189894
R126 plus.n61 plus.n48 0.189894
R127 plus.n65 plus.n48 0.189894
R128 plus.n66 plus.n65 0.189894
R129 plus.n67 plus.n66 0.189894
R130 plus.n67 plus.n46 0.189894
R131 plus.n71 plus.n46 0.189894
R132 plus.n72 plus.n71 0.189894
R133 plus.n73 plus.n72 0.189894
R134 plus.n73 plus.n44 0.189894
R135 plus.n77 plus.n44 0.189894
R136 plus.n78 plus.n77 0.189894
R137 plus.n79 plus.n78 0.189894
R138 plus.n79 plus.n42 0.189894
R139 plus.n83 plus.n42 0.189894
R140 plus.n41 plus.n0 0.189894
R141 plus.n1 plus.n0 0.189894
R142 plus.n36 plus.n1 0.189894
R143 plus.n36 plus.n35 0.189894
R144 plus.n35 plus.n34 0.189894
R145 plus.n34 plus.n3 0.189894
R146 plus.n30 plus.n3 0.189894
R147 plus.n30 plus.n29 0.189894
R148 plus.n29 plus.n28 0.189894
R149 plus.n28 plus.n5 0.189894
R150 plus.n24 plus.n5 0.189894
R151 plus.n24 plus.n23 0.189894
R152 plus.n23 plus.n22 0.189894
R153 plus.n22 plus.n7 0.189894
R154 plus.n18 plus.n7 0.189894
R155 plus.n18 plus.n17 0.189894
R156 plus.n17 plus.n16 0.189894
R157 plus.n16 plus.n9 0.189894
R158 plus.n12 plus.n9 0.189894
R159 a_n2903_n3924.n11 a_n2903_n3924.t55 214.643
R160 a_n2903_n3924.n7 a_n2903_n3924.t15 214.321
R161 a_n2903_n3924.n7 a_n2903_n3924.t19 214.321
R162 a_n2903_n3924.n5 a_n2903_n3924.t24 214.321
R163 a_n2903_n3924.n5 a_n2903_n3924.t21 214.321
R164 a_n2903_n3924.n6 a_n2903_n3924.t14 214.321
R165 a_n2903_n3924.n6 a_n2903_n3924.t53 214.321
R166 a_n2903_n3924.n11 a_n2903_n3924.t11 214.321
R167 a_n2903_n3924.n1 a_n2903_n3924.t50 55.8337
R168 a_n2903_n3924.n1 a_n2903_n3924.t22 55.8337
R169 a_n2903_n3924.n10 a_n2903_n3924.t1 55.8337
R170 a_n2903_n3924.n0 a_n2903_n3924.t37 55.8335
R171 a_n2903_n3924.n8 a_n2903_n3924.t13 55.8335
R172 a_n2903_n3924.n4 a_n2903_n3924.t2 55.8335
R173 a_n2903_n3924.n4 a_n2903_n3924.t42 55.8335
R174 a_n2903_n3924.n3 a_n2903_n3924.t47 55.8335
R175 a_n2903_n3924.n0 a_n2903_n3924.n28 53.0052
R176 a_n2903_n3924.n0 a_n2903_n3924.n29 53.0052
R177 a_n2903_n3924.n0 a_n2903_n3924.n30 53.0052
R178 a_n2903_n3924.n1 a_n2903_n3924.n31 53.0052
R179 a_n2903_n3924.n1 a_n2903_n3924.n32 53.0052
R180 a_n2903_n3924.n1 a_n2903_n3924.n12 53.0052
R181 a_n2903_n3924.n9 a_n2903_n3924.n13 53.0052
R182 a_n2903_n3924.n9 a_n2903_n3924.n14 53.0052
R183 a_n2903_n3924.n10 a_n2903_n3924.n15 53.0052
R184 a_n2903_n3924.n8 a_n2903_n3924.n26 53.0051
R185 a_n2903_n3924.n2 a_n2903_n3924.n25 53.0051
R186 a_n2903_n3924.n2 a_n2903_n3924.n24 53.0051
R187 a_n2903_n3924.n2 a_n2903_n3924.n23 53.0051
R188 a_n2903_n3924.n2 a_n2903_n3924.n22 53.0051
R189 a_n2903_n3924.n4 a_n2903_n3924.n21 53.0051
R190 a_n2903_n3924.n4 a_n2903_n3924.n20 53.0051
R191 a_n2903_n3924.n4 a_n2903_n3924.n19 53.0051
R192 a_n2903_n3924.n3 a_n2903_n3924.n18 53.0051
R193 a_n2903_n3924.n3 a_n2903_n3924.n17 53.0051
R194 a_n2903_n3924.n33 a_n2903_n3924.n1 53.0051
R195 a_n2903_n3924.n16 a_n2903_n3924.n10 12.1986
R196 a_n2903_n3924.n0 a_n2903_n3924.n27 12.1986
R197 a_n2903_n3924.n3 a_n2903_n3924.n16 5.11903
R198 a_n2903_n3924.n27 a_n2903_n3924.n8 5.11903
R199 a_n2903_n3924.n28 a_n2903_n3924.t35 2.82907
R200 a_n2903_n3924.n28 a_n2903_n3924.t33 2.82907
R201 a_n2903_n3924.n29 a_n2903_n3924.t31 2.82907
R202 a_n2903_n3924.n29 a_n2903_n3924.t34 2.82907
R203 a_n2903_n3924.n30 a_n2903_n3924.t40 2.82907
R204 a_n2903_n3924.n30 a_n2903_n3924.t41 2.82907
R205 a_n2903_n3924.n31 a_n2903_n3924.t38 2.82907
R206 a_n2903_n3924.n31 a_n2903_n3924.t51 2.82907
R207 a_n2903_n3924.n32 a_n2903_n3924.t28 2.82907
R208 a_n2903_n3924.n32 a_n2903_n3924.t44 2.82907
R209 a_n2903_n3924.n12 a_n2903_n3924.t26 2.82907
R210 a_n2903_n3924.n12 a_n2903_n3924.t3 2.82907
R211 a_n2903_n3924.n13 a_n2903_n3924.t27 2.82907
R212 a_n2903_n3924.n13 a_n2903_n3924.t8 2.82907
R213 a_n2903_n3924.n14 a_n2903_n3924.t4 2.82907
R214 a_n2903_n3924.n14 a_n2903_n3924.t9 2.82907
R215 a_n2903_n3924.n15 a_n2903_n3924.t6 2.82907
R216 a_n2903_n3924.n15 a_n2903_n3924.t18 2.82907
R217 a_n2903_n3924.n26 a_n2903_n3924.t7 2.82907
R218 a_n2903_n3924.n26 a_n2903_n3924.t23 2.82907
R219 a_n2903_n3924.n25 a_n2903_n3924.t54 2.82907
R220 a_n2903_n3924.n25 a_n2903_n3924.t52 2.82907
R221 a_n2903_n3924.n24 a_n2903_n3924.t20 2.82907
R222 a_n2903_n3924.n24 a_n2903_n3924.t25 2.82907
R223 a_n2903_n3924.n23 a_n2903_n3924.t17 2.82907
R224 a_n2903_n3924.n23 a_n2903_n3924.t12 2.82907
R225 a_n2903_n3924.n22 a_n2903_n3924.t10 2.82907
R226 a_n2903_n3924.n22 a_n2903_n3924.t16 2.82907
R227 a_n2903_n3924.n21 a_n2903_n3924.t39 2.82907
R228 a_n2903_n3924.n21 a_n2903_n3924.t36 2.82907
R229 a_n2903_n3924.n20 a_n2903_n3924.t49 2.82907
R230 a_n2903_n3924.n20 a_n2903_n3924.t43 2.82907
R231 a_n2903_n3924.n19 a_n2903_n3924.t45 2.82907
R232 a_n2903_n3924.n19 a_n2903_n3924.t48 2.82907
R233 a_n2903_n3924.n18 a_n2903_n3924.t30 2.82907
R234 a_n2903_n3924.n18 a_n2903_n3924.t29 2.82907
R235 a_n2903_n3924.n17 a_n2903_n3924.t46 2.82907
R236 a_n2903_n3924.n17 a_n2903_n3924.t32 2.82907
R237 a_n2903_n3924.t0 a_n2903_n3924.n33 2.82907
R238 a_n2903_n3924.n33 a_n2903_n3924.t5 2.82907
R239 a_n2903_n3924.n1 a_n2903_n3924.n0 2.66429
R240 a_n2903_n3924.n27 a_n2903_n3924.n7 2.16406
R241 a_n2903_n3924.n2 a_n2903_n3924.n4 2.01128
R242 a_n2903_n3924.n16 a_n2903_n3924.n11 1.95694
R243 a_n2903_n3924.n4 a_n2903_n3924.n3 1.77636
R244 a_n2903_n3924.n8 a_n2903_n3924.n2 1.77636
R245 a_n2903_n3924.n11 a_n2903_n3924.n6 1.69309
R246 a_n2903_n3924.n9 a_n2903_n3924.n1 1.56731
R247 a_n2903_n3924.n5 a_n2903_n3924.n7 1.34352
R248 a_n2903_n3924.n6 a_n2903_n3924.n5 1.34352
R249 a_n2903_n3924.n10 a_n2903_n3924.n9 1.3324
R250 a_n8300_8799.n141 a_n8300_8799.t113 490.524
R251 a_n8300_8799.n175 a_n8300_8799.t49 490.524
R252 a_n8300_8799.n210 a_n8300_8799.t97 490.524
R253 a_n8300_8799.n35 a_n8300_8799.t89 490.524
R254 a_n8300_8799.n69 a_n8300_8799.t96 490.524
R255 a_n8300_8799.n104 a_n8300_8799.t98 490.524
R256 a_n8300_8799.n162 a_n8300_8799.t51 464.166
R257 a_n8300_8799.n160 a_n8300_8799.t50 464.166
R258 a_n8300_8799.n159 a_n8300_8799.t100 464.166
R259 a_n8300_8799.n133 a_n8300_8799.t61 464.166
R260 a_n8300_8799.n153 a_n8300_8799.t53 464.166
R261 a_n8300_8799.n152 a_n8300_8799.t104 464.166
R262 a_n8300_8799.n136 a_n8300_8799.t77 464.166
R263 a_n8300_8799.n147 a_n8300_8799.t62 464.166
R264 a_n8300_8799.n145 a_n8300_8799.t117 464.166
R265 a_n8300_8799.n139 a_n8300_8799.t88 464.166
R266 a_n8300_8799.n140 a_n8300_8799.t64 464.166
R267 a_n8300_8799.n196 a_n8300_8799.t57 464.166
R268 a_n8300_8799.n194 a_n8300_8799.t56 464.166
R269 a_n8300_8799.n193 a_n8300_8799.t112 464.166
R270 a_n8300_8799.n167 a_n8300_8799.t66 464.166
R271 a_n8300_8799.n187 a_n8300_8799.t60 464.166
R272 a_n8300_8799.n186 a_n8300_8799.t114 464.166
R273 a_n8300_8799.n170 a_n8300_8799.t86 464.166
R274 a_n8300_8799.n181 a_n8300_8799.t69 464.166
R275 a_n8300_8799.n179 a_n8300_8799.t52 464.166
R276 a_n8300_8799.n173 a_n8300_8799.t95 464.166
R277 a_n8300_8799.n174 a_n8300_8799.t70 464.166
R278 a_n8300_8799.n231 a_n8300_8799.t85 464.166
R279 a_n8300_8799.n229 a_n8300_8799.t99 464.166
R280 a_n8300_8799.n228 a_n8300_8799.t59 464.166
R281 a_n8300_8799.n202 a_n8300_8799.t110 464.166
R282 a_n8300_8799.n222 a_n8300_8799.t73 464.166
R283 a_n8300_8799.n221 a_n8300_8799.t105 464.166
R284 a_n8300_8799.n205 a_n8300_8799.t63 464.166
R285 a_n8300_8799.n216 a_n8300_8799.t91 464.166
R286 a_n8300_8799.n214 a_n8300_8799.t55 464.166
R287 a_n8300_8799.n208 a_n8300_8799.t82 464.166
R288 a_n8300_8799.n209 a_n8300_8799.t68 464.166
R289 a_n8300_8799.n34 a_n8300_8799.t111 464.166
R290 a_n8300_8799.n33 a_n8300_8799.t65 464.166
R291 a_n8300_8799.n39 a_n8300_8799.t87 464.166
R292 a_n8300_8799.n31 a_n8300_8799.t107 464.166
R293 a_n8300_8799.n44 a_n8300_8799.t108 464.166
R294 a_n8300_8799.n46 a_n8300_8799.t76 464.166
R295 a_n8300_8799.n29 a_n8300_8799.t94 464.166
R296 a_n8300_8799.n51 a_n8300_8799.t106 464.166
R297 a_n8300_8799.n27 a_n8300_8799.t74 464.166
R298 a_n8300_8799.n56 a_n8300_8799.t75 464.166
R299 a_n8300_8799.n58 a_n8300_8799.t92 464.166
R300 a_n8300_8799.n68 a_n8300_8799.t119 464.166
R301 a_n8300_8799.n67 a_n8300_8799.t71 464.166
R302 a_n8300_8799.n73 a_n8300_8799.t93 464.166
R303 a_n8300_8799.n65 a_n8300_8799.t116 464.166
R304 a_n8300_8799.n78 a_n8300_8799.t118 464.166
R305 a_n8300_8799.n80 a_n8300_8799.t83 464.166
R306 a_n8300_8799.n63 a_n8300_8799.t103 464.166
R307 a_n8300_8799.n85 a_n8300_8799.t115 464.166
R308 a_n8300_8799.n61 a_n8300_8799.t79 464.166
R309 a_n8300_8799.n90 a_n8300_8799.t80 464.166
R310 a_n8300_8799.n92 a_n8300_8799.t101 464.166
R311 a_n8300_8799.n103 a_n8300_8799.t67 464.166
R312 a_n8300_8799.n102 a_n8300_8799.t81 464.166
R313 a_n8300_8799.n108 a_n8300_8799.t54 464.166
R314 a_n8300_8799.n100 a_n8300_8799.t90 464.166
R315 a_n8300_8799.n113 a_n8300_8799.t78 464.166
R316 a_n8300_8799.n115 a_n8300_8799.t102 464.166
R317 a_n8300_8799.n98 a_n8300_8799.t72 464.166
R318 a_n8300_8799.n120 a_n8300_8799.t109 464.166
R319 a_n8300_8799.n96 a_n8300_8799.t58 464.166
R320 a_n8300_8799.n125 a_n8300_8799.t48 464.166
R321 a_n8300_8799.n127 a_n8300_8799.t84 464.166
R322 a_n8300_8799.n142 a_n8300_8799.n139 161.3
R323 a_n8300_8799.n144 a_n8300_8799.n143 161.3
R324 a_n8300_8799.n145 a_n8300_8799.n138 161.3
R325 a_n8300_8799.n146 a_n8300_8799.n137 161.3
R326 a_n8300_8799.n148 a_n8300_8799.n147 161.3
R327 a_n8300_8799.n149 a_n8300_8799.n136 161.3
R328 a_n8300_8799.n151 a_n8300_8799.n150 161.3
R329 a_n8300_8799.n152 a_n8300_8799.n135 161.3
R330 a_n8300_8799.n153 a_n8300_8799.n134 161.3
R331 a_n8300_8799.n155 a_n8300_8799.n154 161.3
R332 a_n8300_8799.n156 a_n8300_8799.n133 161.3
R333 a_n8300_8799.n158 a_n8300_8799.n157 161.3
R334 a_n8300_8799.n159 a_n8300_8799.n132 161.3
R335 a_n8300_8799.n160 a_n8300_8799.n131 161.3
R336 a_n8300_8799.n161 a_n8300_8799.n130 161.3
R337 a_n8300_8799.n163 a_n8300_8799.n162 161.3
R338 a_n8300_8799.n176 a_n8300_8799.n173 161.3
R339 a_n8300_8799.n178 a_n8300_8799.n177 161.3
R340 a_n8300_8799.n179 a_n8300_8799.n172 161.3
R341 a_n8300_8799.n180 a_n8300_8799.n171 161.3
R342 a_n8300_8799.n182 a_n8300_8799.n181 161.3
R343 a_n8300_8799.n183 a_n8300_8799.n170 161.3
R344 a_n8300_8799.n185 a_n8300_8799.n184 161.3
R345 a_n8300_8799.n186 a_n8300_8799.n169 161.3
R346 a_n8300_8799.n187 a_n8300_8799.n168 161.3
R347 a_n8300_8799.n189 a_n8300_8799.n188 161.3
R348 a_n8300_8799.n190 a_n8300_8799.n167 161.3
R349 a_n8300_8799.n192 a_n8300_8799.n191 161.3
R350 a_n8300_8799.n193 a_n8300_8799.n166 161.3
R351 a_n8300_8799.n194 a_n8300_8799.n165 161.3
R352 a_n8300_8799.n195 a_n8300_8799.n164 161.3
R353 a_n8300_8799.n197 a_n8300_8799.n196 161.3
R354 a_n8300_8799.n211 a_n8300_8799.n208 161.3
R355 a_n8300_8799.n213 a_n8300_8799.n212 161.3
R356 a_n8300_8799.n214 a_n8300_8799.n207 161.3
R357 a_n8300_8799.n215 a_n8300_8799.n206 161.3
R358 a_n8300_8799.n217 a_n8300_8799.n216 161.3
R359 a_n8300_8799.n218 a_n8300_8799.n205 161.3
R360 a_n8300_8799.n220 a_n8300_8799.n219 161.3
R361 a_n8300_8799.n221 a_n8300_8799.n204 161.3
R362 a_n8300_8799.n222 a_n8300_8799.n203 161.3
R363 a_n8300_8799.n224 a_n8300_8799.n223 161.3
R364 a_n8300_8799.n225 a_n8300_8799.n202 161.3
R365 a_n8300_8799.n227 a_n8300_8799.n226 161.3
R366 a_n8300_8799.n228 a_n8300_8799.n201 161.3
R367 a_n8300_8799.n229 a_n8300_8799.n200 161.3
R368 a_n8300_8799.n230 a_n8300_8799.n199 161.3
R369 a_n8300_8799.n232 a_n8300_8799.n231 161.3
R370 a_n8300_8799.n59 a_n8300_8799.n58 161.3
R371 a_n8300_8799.n57 a_n8300_8799.n26 161.3
R372 a_n8300_8799.n56 a_n8300_8799.n55 161.3
R373 a_n8300_8799.n54 a_n8300_8799.n27 161.3
R374 a_n8300_8799.n53 a_n8300_8799.n52 161.3
R375 a_n8300_8799.n51 a_n8300_8799.n28 161.3
R376 a_n8300_8799.n50 a_n8300_8799.n49 161.3
R377 a_n8300_8799.n48 a_n8300_8799.n29 161.3
R378 a_n8300_8799.n47 a_n8300_8799.n46 161.3
R379 a_n8300_8799.n45 a_n8300_8799.n30 161.3
R380 a_n8300_8799.n44 a_n8300_8799.n43 161.3
R381 a_n8300_8799.n42 a_n8300_8799.n31 161.3
R382 a_n8300_8799.n41 a_n8300_8799.n40 161.3
R383 a_n8300_8799.n39 a_n8300_8799.n32 161.3
R384 a_n8300_8799.n38 a_n8300_8799.n37 161.3
R385 a_n8300_8799.n36 a_n8300_8799.n33 161.3
R386 a_n8300_8799.n93 a_n8300_8799.n92 161.3
R387 a_n8300_8799.n91 a_n8300_8799.n60 161.3
R388 a_n8300_8799.n90 a_n8300_8799.n89 161.3
R389 a_n8300_8799.n88 a_n8300_8799.n61 161.3
R390 a_n8300_8799.n87 a_n8300_8799.n86 161.3
R391 a_n8300_8799.n85 a_n8300_8799.n62 161.3
R392 a_n8300_8799.n84 a_n8300_8799.n83 161.3
R393 a_n8300_8799.n82 a_n8300_8799.n63 161.3
R394 a_n8300_8799.n81 a_n8300_8799.n80 161.3
R395 a_n8300_8799.n79 a_n8300_8799.n64 161.3
R396 a_n8300_8799.n78 a_n8300_8799.n77 161.3
R397 a_n8300_8799.n76 a_n8300_8799.n65 161.3
R398 a_n8300_8799.n75 a_n8300_8799.n74 161.3
R399 a_n8300_8799.n73 a_n8300_8799.n66 161.3
R400 a_n8300_8799.n72 a_n8300_8799.n71 161.3
R401 a_n8300_8799.n70 a_n8300_8799.n67 161.3
R402 a_n8300_8799.n128 a_n8300_8799.n127 161.3
R403 a_n8300_8799.n126 a_n8300_8799.n95 161.3
R404 a_n8300_8799.n125 a_n8300_8799.n124 161.3
R405 a_n8300_8799.n123 a_n8300_8799.n96 161.3
R406 a_n8300_8799.n122 a_n8300_8799.n121 161.3
R407 a_n8300_8799.n120 a_n8300_8799.n97 161.3
R408 a_n8300_8799.n119 a_n8300_8799.n118 161.3
R409 a_n8300_8799.n117 a_n8300_8799.n98 161.3
R410 a_n8300_8799.n116 a_n8300_8799.n115 161.3
R411 a_n8300_8799.n114 a_n8300_8799.n99 161.3
R412 a_n8300_8799.n113 a_n8300_8799.n112 161.3
R413 a_n8300_8799.n111 a_n8300_8799.n100 161.3
R414 a_n8300_8799.n110 a_n8300_8799.n109 161.3
R415 a_n8300_8799.n108 a_n8300_8799.n101 161.3
R416 a_n8300_8799.n107 a_n8300_8799.n106 161.3
R417 a_n8300_8799.n105 a_n8300_8799.n102 161.3
R418 a_n8300_8799.n16 a_n8300_8799.n14 98.9633
R419 a_n8300_8799.n5 a_n8300_8799.n3 98.9631
R420 a_n8300_8799.n24 a_n8300_8799.n23 98.6055
R421 a_n8300_8799.n22 a_n8300_8799.n21 98.6055
R422 a_n8300_8799.n20 a_n8300_8799.n19 98.6055
R423 a_n8300_8799.n18 a_n8300_8799.n17 98.6055
R424 a_n8300_8799.n16 a_n8300_8799.n15 98.6055
R425 a_n8300_8799.n5 a_n8300_8799.n4 98.6055
R426 a_n8300_8799.n7 a_n8300_8799.n6 98.6055
R427 a_n8300_8799.n9 a_n8300_8799.n8 98.6055
R428 a_n8300_8799.n11 a_n8300_8799.n10 98.6055
R429 a_n8300_8799.n13 a_n8300_8799.n12 98.6055
R430 a_n8300_8799.n238 a_n8300_8799.n236 81.3764
R431 a_n8300_8799.n250 a_n8300_8799.n248 81.3764
R432 a_n8300_8799.n2 a_n8300_8799.n0 81.3764
R433 a_n8300_8799.n255 a_n8300_8799.n254 80.9326
R434 a_n8300_8799.n247 a_n8300_8799.n246 80.9324
R435 a_n8300_8799.n245 a_n8300_8799.n244 80.9324
R436 a_n8300_8799.n243 a_n8300_8799.n242 80.9324
R437 a_n8300_8799.n240 a_n8300_8799.n239 80.9324
R438 a_n8300_8799.n238 a_n8300_8799.n237 80.9324
R439 a_n8300_8799.n250 a_n8300_8799.n249 80.9324
R440 a_n8300_8799.n252 a_n8300_8799.n251 80.9324
R441 a_n8300_8799.n2 a_n8300_8799.n1 80.9324
R442 a_n8300_8799.n160 a_n8300_8799.n159 48.2005
R443 a_n8300_8799.n153 a_n8300_8799.n152 48.2005
R444 a_n8300_8799.n147 a_n8300_8799.n136 48.2005
R445 a_n8300_8799.n140 a_n8300_8799.n139 48.2005
R446 a_n8300_8799.n194 a_n8300_8799.n193 48.2005
R447 a_n8300_8799.n187 a_n8300_8799.n186 48.2005
R448 a_n8300_8799.n181 a_n8300_8799.n170 48.2005
R449 a_n8300_8799.n174 a_n8300_8799.n173 48.2005
R450 a_n8300_8799.n229 a_n8300_8799.n228 48.2005
R451 a_n8300_8799.n222 a_n8300_8799.n221 48.2005
R452 a_n8300_8799.n216 a_n8300_8799.n205 48.2005
R453 a_n8300_8799.n209 a_n8300_8799.n208 48.2005
R454 a_n8300_8799.n34 a_n8300_8799.n33 48.2005
R455 a_n8300_8799.n44 a_n8300_8799.n31 48.2005
R456 a_n8300_8799.n46 a_n8300_8799.n29 48.2005
R457 a_n8300_8799.n56 a_n8300_8799.n27 48.2005
R458 a_n8300_8799.n68 a_n8300_8799.n67 48.2005
R459 a_n8300_8799.n78 a_n8300_8799.n65 48.2005
R460 a_n8300_8799.n80 a_n8300_8799.n63 48.2005
R461 a_n8300_8799.n90 a_n8300_8799.n61 48.2005
R462 a_n8300_8799.n103 a_n8300_8799.n102 48.2005
R463 a_n8300_8799.n113 a_n8300_8799.n100 48.2005
R464 a_n8300_8799.n115 a_n8300_8799.n98 48.2005
R465 a_n8300_8799.n125 a_n8300_8799.n96 48.2005
R466 a_n8300_8799.n154 a_n8300_8799.n133 47.4702
R467 a_n8300_8799.n146 a_n8300_8799.n145 47.4702
R468 a_n8300_8799.n188 a_n8300_8799.n167 47.4702
R469 a_n8300_8799.n180 a_n8300_8799.n179 47.4702
R470 a_n8300_8799.n223 a_n8300_8799.n202 47.4702
R471 a_n8300_8799.n215 a_n8300_8799.n214 47.4702
R472 a_n8300_8799.n40 a_n8300_8799.n39 47.4702
R473 a_n8300_8799.n51 a_n8300_8799.n50 47.4702
R474 a_n8300_8799.n74 a_n8300_8799.n73 47.4702
R475 a_n8300_8799.n85 a_n8300_8799.n84 47.4702
R476 a_n8300_8799.n109 a_n8300_8799.n108 47.4702
R477 a_n8300_8799.n120 a_n8300_8799.n119 47.4702
R478 a_n8300_8799.n162 a_n8300_8799.n161 46.0096
R479 a_n8300_8799.n196 a_n8300_8799.n195 46.0096
R480 a_n8300_8799.n231 a_n8300_8799.n230 46.0096
R481 a_n8300_8799.n58 a_n8300_8799.n57 46.0096
R482 a_n8300_8799.n92 a_n8300_8799.n91 46.0096
R483 a_n8300_8799.n127 a_n8300_8799.n126 46.0096
R484 a_n8300_8799.n36 a_n8300_8799.n35 45.0871
R485 a_n8300_8799.n70 a_n8300_8799.n69 45.0871
R486 a_n8300_8799.n105 a_n8300_8799.n104 45.0871
R487 a_n8300_8799.n142 a_n8300_8799.n141 45.0871
R488 a_n8300_8799.n176 a_n8300_8799.n175 45.0871
R489 a_n8300_8799.n211 a_n8300_8799.n210 45.0871
R490 a_n8300_8799.n25 a_n8300_8799.n13 34.1553
R491 a_n8300_8799.n253 a_n8300_8799.n247 33.4185
R492 a_n8300_8799.n158 a_n8300_8799.n133 25.5611
R493 a_n8300_8799.n145 a_n8300_8799.n144 25.5611
R494 a_n8300_8799.n192 a_n8300_8799.n167 25.5611
R495 a_n8300_8799.n179 a_n8300_8799.n178 25.5611
R496 a_n8300_8799.n227 a_n8300_8799.n202 25.5611
R497 a_n8300_8799.n214 a_n8300_8799.n213 25.5611
R498 a_n8300_8799.n39 a_n8300_8799.n38 25.5611
R499 a_n8300_8799.n52 a_n8300_8799.n51 25.5611
R500 a_n8300_8799.n73 a_n8300_8799.n72 25.5611
R501 a_n8300_8799.n86 a_n8300_8799.n85 25.5611
R502 a_n8300_8799.n108 a_n8300_8799.n107 25.5611
R503 a_n8300_8799.n121 a_n8300_8799.n120 25.5611
R504 a_n8300_8799.n152 a_n8300_8799.n151 24.1005
R505 a_n8300_8799.n151 a_n8300_8799.n136 24.1005
R506 a_n8300_8799.n186 a_n8300_8799.n185 24.1005
R507 a_n8300_8799.n185 a_n8300_8799.n170 24.1005
R508 a_n8300_8799.n221 a_n8300_8799.n220 24.1005
R509 a_n8300_8799.n220 a_n8300_8799.n205 24.1005
R510 a_n8300_8799.n45 a_n8300_8799.n44 24.1005
R511 a_n8300_8799.n46 a_n8300_8799.n45 24.1005
R512 a_n8300_8799.n79 a_n8300_8799.n78 24.1005
R513 a_n8300_8799.n80 a_n8300_8799.n79 24.1005
R514 a_n8300_8799.n114 a_n8300_8799.n113 24.1005
R515 a_n8300_8799.n115 a_n8300_8799.n114 24.1005
R516 a_n8300_8799.n159 a_n8300_8799.n158 22.6399
R517 a_n8300_8799.n144 a_n8300_8799.n139 22.6399
R518 a_n8300_8799.n193 a_n8300_8799.n192 22.6399
R519 a_n8300_8799.n178 a_n8300_8799.n173 22.6399
R520 a_n8300_8799.n228 a_n8300_8799.n227 22.6399
R521 a_n8300_8799.n213 a_n8300_8799.n208 22.6399
R522 a_n8300_8799.n38 a_n8300_8799.n33 22.6399
R523 a_n8300_8799.n52 a_n8300_8799.n27 22.6399
R524 a_n8300_8799.n72 a_n8300_8799.n67 22.6399
R525 a_n8300_8799.n86 a_n8300_8799.n61 22.6399
R526 a_n8300_8799.n107 a_n8300_8799.n102 22.6399
R527 a_n8300_8799.n121 a_n8300_8799.n96 22.6399
R528 a_n8300_8799.n25 a_n8300_8799.n24 20.7339
R529 a_n8300_8799.n141 a_n8300_8799.n140 14.1472
R530 a_n8300_8799.n175 a_n8300_8799.n174 14.1472
R531 a_n8300_8799.n210 a_n8300_8799.n209 14.1472
R532 a_n8300_8799.n35 a_n8300_8799.n34 14.1472
R533 a_n8300_8799.n69 a_n8300_8799.n68 14.1472
R534 a_n8300_8799.n104 a_n8300_8799.n103 14.1472
R535 a_n8300_8799.n241 a_n8300_8799.n235 12.3339
R536 a_n8300_8799.n235 a_n8300_8799.n25 11.4887
R537 a_n8300_8799.n198 a_n8300_8799.n163 9.01755
R538 a_n8300_8799.n94 a_n8300_8799.n59 9.01755
R539 a_n8300_8799.n234 a_n8300_8799.n129 7.2142
R540 a_n8300_8799.n234 a_n8300_8799.n233 6.79277
R541 a_n8300_8799.n198 a_n8300_8799.n197 4.90959
R542 a_n8300_8799.n233 a_n8300_8799.n232 4.90959
R543 a_n8300_8799.n94 a_n8300_8799.n93 4.90959
R544 a_n8300_8799.n129 a_n8300_8799.n128 4.90959
R545 a_n8300_8799.n233 a_n8300_8799.n198 4.10845
R546 a_n8300_8799.n129 a_n8300_8799.n94 4.10845
R547 a_n8300_8799.n23 a_n8300_8799.t16 3.61217
R548 a_n8300_8799.n23 a_n8300_8799.t1 3.61217
R549 a_n8300_8799.n21 a_n8300_8799.t5 3.61217
R550 a_n8300_8799.n21 a_n8300_8799.t19 3.61217
R551 a_n8300_8799.n19 a_n8300_8799.t6 3.61217
R552 a_n8300_8799.n19 a_n8300_8799.t12 3.61217
R553 a_n8300_8799.n17 a_n8300_8799.t8 3.61217
R554 a_n8300_8799.n17 a_n8300_8799.t7 3.61217
R555 a_n8300_8799.n15 a_n8300_8799.t9 3.61217
R556 a_n8300_8799.n15 a_n8300_8799.t2 3.61217
R557 a_n8300_8799.n14 a_n8300_8799.t47 3.61217
R558 a_n8300_8799.n14 a_n8300_8799.t11 3.61217
R559 a_n8300_8799.n3 a_n8300_8799.t3 3.61217
R560 a_n8300_8799.n3 a_n8300_8799.t0 3.61217
R561 a_n8300_8799.n4 a_n8300_8799.t17 3.61217
R562 a_n8300_8799.n4 a_n8300_8799.t13 3.61217
R563 a_n8300_8799.n6 a_n8300_8799.t45 3.61217
R564 a_n8300_8799.n6 a_n8300_8799.t10 3.61217
R565 a_n8300_8799.n8 a_n8300_8799.t18 3.61217
R566 a_n8300_8799.n8 a_n8300_8799.t15 3.61217
R567 a_n8300_8799.n10 a_n8300_8799.t46 3.61217
R568 a_n8300_8799.n10 a_n8300_8799.t4 3.61217
R569 a_n8300_8799.n12 a_n8300_8799.t14 3.61217
R570 a_n8300_8799.n12 a_n8300_8799.t20 3.61217
R571 a_n8300_8799.n235 a_n8300_8799.n234 3.4105
R572 a_n8300_8799.n248 a_n8300_8799.t36 2.82907
R573 a_n8300_8799.n248 a_n8300_8799.t34 2.82907
R574 a_n8300_8799.n249 a_n8300_8799.t25 2.82907
R575 a_n8300_8799.n249 a_n8300_8799.t31 2.82907
R576 a_n8300_8799.n251 a_n8300_8799.t43 2.82907
R577 a_n8300_8799.n251 a_n8300_8799.t26 2.82907
R578 a_n8300_8799.n1 a_n8300_8799.t33 2.82907
R579 a_n8300_8799.n1 a_n8300_8799.t32 2.82907
R580 a_n8300_8799.n0 a_n8300_8799.t28 2.82907
R581 a_n8300_8799.n0 a_n8300_8799.t27 2.82907
R582 a_n8300_8799.n246 a_n8300_8799.t39 2.82907
R583 a_n8300_8799.n246 a_n8300_8799.t41 2.82907
R584 a_n8300_8799.n244 a_n8300_8799.t37 2.82907
R585 a_n8300_8799.n244 a_n8300_8799.t21 2.82907
R586 a_n8300_8799.n242 a_n8300_8799.t42 2.82907
R587 a_n8300_8799.n242 a_n8300_8799.t35 2.82907
R588 a_n8300_8799.n239 a_n8300_8799.t22 2.82907
R589 a_n8300_8799.n239 a_n8300_8799.t40 2.82907
R590 a_n8300_8799.n237 a_n8300_8799.t23 2.82907
R591 a_n8300_8799.n237 a_n8300_8799.t24 2.82907
R592 a_n8300_8799.n236 a_n8300_8799.t29 2.82907
R593 a_n8300_8799.n236 a_n8300_8799.t30 2.82907
R594 a_n8300_8799.n255 a_n8300_8799.t38 2.82907
R595 a_n8300_8799.t44 a_n8300_8799.n255 2.82907
R596 a_n8300_8799.n161 a_n8300_8799.n160 2.19141
R597 a_n8300_8799.n195 a_n8300_8799.n194 2.19141
R598 a_n8300_8799.n230 a_n8300_8799.n229 2.19141
R599 a_n8300_8799.n57 a_n8300_8799.n56 2.19141
R600 a_n8300_8799.n91 a_n8300_8799.n90 2.19141
R601 a_n8300_8799.n126 a_n8300_8799.n125 2.19141
R602 a_n8300_8799.n154 a_n8300_8799.n153 0.730803
R603 a_n8300_8799.n147 a_n8300_8799.n146 0.730803
R604 a_n8300_8799.n188 a_n8300_8799.n187 0.730803
R605 a_n8300_8799.n181 a_n8300_8799.n180 0.730803
R606 a_n8300_8799.n223 a_n8300_8799.n222 0.730803
R607 a_n8300_8799.n216 a_n8300_8799.n215 0.730803
R608 a_n8300_8799.n40 a_n8300_8799.n31 0.730803
R609 a_n8300_8799.n50 a_n8300_8799.n29 0.730803
R610 a_n8300_8799.n74 a_n8300_8799.n65 0.730803
R611 a_n8300_8799.n84 a_n8300_8799.n63 0.730803
R612 a_n8300_8799.n109 a_n8300_8799.n100 0.730803
R613 a_n8300_8799.n119 a_n8300_8799.n98 0.730803
R614 a_n8300_8799.n240 a_n8300_8799.n238 0.444466
R615 a_n8300_8799.n245 a_n8300_8799.n243 0.444466
R616 a_n8300_8799.n247 a_n8300_8799.n245 0.444466
R617 a_n8300_8799.n254 a_n8300_8799.n2 0.444466
R618 a_n8300_8799.n252 a_n8300_8799.n250 0.444466
R619 a_n8300_8799.n18 a_n8300_8799.n16 0.358259
R620 a_n8300_8799.n20 a_n8300_8799.n18 0.358259
R621 a_n8300_8799.n22 a_n8300_8799.n20 0.358259
R622 a_n8300_8799.n24 a_n8300_8799.n22 0.358259
R623 a_n8300_8799.n13 a_n8300_8799.n11 0.358259
R624 a_n8300_8799.n11 a_n8300_8799.n9 0.358259
R625 a_n8300_8799.n9 a_n8300_8799.n7 0.358259
R626 a_n8300_8799.n7 a_n8300_8799.n5 0.358259
R627 a_n8300_8799.n241 a_n8300_8799.n240 0.222483
R628 a_n8300_8799.n243 a_n8300_8799.n241 0.222483
R629 a_n8300_8799.n254 a_n8300_8799.n253 0.222483
R630 a_n8300_8799.n253 a_n8300_8799.n252 0.222483
R631 a_n8300_8799.n163 a_n8300_8799.n130 0.189894
R632 a_n8300_8799.n131 a_n8300_8799.n130 0.189894
R633 a_n8300_8799.n132 a_n8300_8799.n131 0.189894
R634 a_n8300_8799.n157 a_n8300_8799.n132 0.189894
R635 a_n8300_8799.n157 a_n8300_8799.n156 0.189894
R636 a_n8300_8799.n156 a_n8300_8799.n155 0.189894
R637 a_n8300_8799.n155 a_n8300_8799.n134 0.189894
R638 a_n8300_8799.n135 a_n8300_8799.n134 0.189894
R639 a_n8300_8799.n150 a_n8300_8799.n135 0.189894
R640 a_n8300_8799.n150 a_n8300_8799.n149 0.189894
R641 a_n8300_8799.n149 a_n8300_8799.n148 0.189894
R642 a_n8300_8799.n148 a_n8300_8799.n137 0.189894
R643 a_n8300_8799.n138 a_n8300_8799.n137 0.189894
R644 a_n8300_8799.n143 a_n8300_8799.n138 0.189894
R645 a_n8300_8799.n143 a_n8300_8799.n142 0.189894
R646 a_n8300_8799.n197 a_n8300_8799.n164 0.189894
R647 a_n8300_8799.n165 a_n8300_8799.n164 0.189894
R648 a_n8300_8799.n166 a_n8300_8799.n165 0.189894
R649 a_n8300_8799.n191 a_n8300_8799.n166 0.189894
R650 a_n8300_8799.n191 a_n8300_8799.n190 0.189894
R651 a_n8300_8799.n190 a_n8300_8799.n189 0.189894
R652 a_n8300_8799.n189 a_n8300_8799.n168 0.189894
R653 a_n8300_8799.n169 a_n8300_8799.n168 0.189894
R654 a_n8300_8799.n184 a_n8300_8799.n169 0.189894
R655 a_n8300_8799.n184 a_n8300_8799.n183 0.189894
R656 a_n8300_8799.n183 a_n8300_8799.n182 0.189894
R657 a_n8300_8799.n182 a_n8300_8799.n171 0.189894
R658 a_n8300_8799.n172 a_n8300_8799.n171 0.189894
R659 a_n8300_8799.n177 a_n8300_8799.n172 0.189894
R660 a_n8300_8799.n177 a_n8300_8799.n176 0.189894
R661 a_n8300_8799.n232 a_n8300_8799.n199 0.189894
R662 a_n8300_8799.n200 a_n8300_8799.n199 0.189894
R663 a_n8300_8799.n201 a_n8300_8799.n200 0.189894
R664 a_n8300_8799.n226 a_n8300_8799.n201 0.189894
R665 a_n8300_8799.n226 a_n8300_8799.n225 0.189894
R666 a_n8300_8799.n225 a_n8300_8799.n224 0.189894
R667 a_n8300_8799.n224 a_n8300_8799.n203 0.189894
R668 a_n8300_8799.n204 a_n8300_8799.n203 0.189894
R669 a_n8300_8799.n219 a_n8300_8799.n204 0.189894
R670 a_n8300_8799.n219 a_n8300_8799.n218 0.189894
R671 a_n8300_8799.n218 a_n8300_8799.n217 0.189894
R672 a_n8300_8799.n217 a_n8300_8799.n206 0.189894
R673 a_n8300_8799.n207 a_n8300_8799.n206 0.189894
R674 a_n8300_8799.n212 a_n8300_8799.n207 0.189894
R675 a_n8300_8799.n212 a_n8300_8799.n211 0.189894
R676 a_n8300_8799.n37 a_n8300_8799.n36 0.189894
R677 a_n8300_8799.n37 a_n8300_8799.n32 0.189894
R678 a_n8300_8799.n41 a_n8300_8799.n32 0.189894
R679 a_n8300_8799.n42 a_n8300_8799.n41 0.189894
R680 a_n8300_8799.n43 a_n8300_8799.n42 0.189894
R681 a_n8300_8799.n43 a_n8300_8799.n30 0.189894
R682 a_n8300_8799.n47 a_n8300_8799.n30 0.189894
R683 a_n8300_8799.n48 a_n8300_8799.n47 0.189894
R684 a_n8300_8799.n49 a_n8300_8799.n48 0.189894
R685 a_n8300_8799.n49 a_n8300_8799.n28 0.189894
R686 a_n8300_8799.n53 a_n8300_8799.n28 0.189894
R687 a_n8300_8799.n54 a_n8300_8799.n53 0.189894
R688 a_n8300_8799.n55 a_n8300_8799.n54 0.189894
R689 a_n8300_8799.n55 a_n8300_8799.n26 0.189894
R690 a_n8300_8799.n59 a_n8300_8799.n26 0.189894
R691 a_n8300_8799.n71 a_n8300_8799.n70 0.189894
R692 a_n8300_8799.n71 a_n8300_8799.n66 0.189894
R693 a_n8300_8799.n75 a_n8300_8799.n66 0.189894
R694 a_n8300_8799.n76 a_n8300_8799.n75 0.189894
R695 a_n8300_8799.n77 a_n8300_8799.n76 0.189894
R696 a_n8300_8799.n77 a_n8300_8799.n64 0.189894
R697 a_n8300_8799.n81 a_n8300_8799.n64 0.189894
R698 a_n8300_8799.n82 a_n8300_8799.n81 0.189894
R699 a_n8300_8799.n83 a_n8300_8799.n82 0.189894
R700 a_n8300_8799.n83 a_n8300_8799.n62 0.189894
R701 a_n8300_8799.n87 a_n8300_8799.n62 0.189894
R702 a_n8300_8799.n88 a_n8300_8799.n87 0.189894
R703 a_n8300_8799.n89 a_n8300_8799.n88 0.189894
R704 a_n8300_8799.n89 a_n8300_8799.n60 0.189894
R705 a_n8300_8799.n93 a_n8300_8799.n60 0.189894
R706 a_n8300_8799.n106 a_n8300_8799.n105 0.189894
R707 a_n8300_8799.n106 a_n8300_8799.n101 0.189894
R708 a_n8300_8799.n110 a_n8300_8799.n101 0.189894
R709 a_n8300_8799.n111 a_n8300_8799.n110 0.189894
R710 a_n8300_8799.n112 a_n8300_8799.n111 0.189894
R711 a_n8300_8799.n112 a_n8300_8799.n99 0.189894
R712 a_n8300_8799.n116 a_n8300_8799.n99 0.189894
R713 a_n8300_8799.n117 a_n8300_8799.n116 0.189894
R714 a_n8300_8799.n118 a_n8300_8799.n117 0.189894
R715 a_n8300_8799.n118 a_n8300_8799.n97 0.189894
R716 a_n8300_8799.n122 a_n8300_8799.n97 0.189894
R717 a_n8300_8799.n123 a_n8300_8799.n122 0.189894
R718 a_n8300_8799.n124 a_n8300_8799.n123 0.189894
R719 a_n8300_8799.n124 a_n8300_8799.n95 0.189894
R720 a_n8300_8799.n128 a_n8300_8799.n95 0.189894
R721 gnd.n7201 gnd.n525 1768.67
R722 gnd.n5165 gnd.n5164 939.716
R723 gnd.n7676 gnd.n208 795.207
R724 gnd.n348 gnd.n211 795.207
R725 gnd.n3903 gnd.n1620 795.207
R726 gnd.n3971 gnd.n1622 795.207
R727 gnd.n4907 gnd.n1372 795.207
R728 gnd.n3190 gnd.n1375 795.207
R729 gnd.n2606 gnd.n1067 795.207
R730 gnd.n2563 gnd.n2562 795.207
R731 gnd.n3178 gnd.n2387 771.183
R732 gnd.n4664 gnd.n1597 771.183
R733 gnd.n3200 gnd.n2398 771.183
R734 gnd.n4059 gnd.n1599 771.183
R735 gnd.n6547 gnd.n1026 766.379
R736 gnd.n6463 gnd.n1028 766.379
R737 gnd.n5675 gnd.n5574 766.379
R738 gnd.n5673 gnd.n5576 766.379
R739 gnd.n6544 gnd.n5167 756.769
R740 gnd.n6513 gnd.n1029 756.769
R741 gnd.n5807 gnd.n5536 756.769
R742 gnd.n5793 gnd.n5525 756.769
R743 gnd.n7674 gnd.n213 739.952
R744 gnd.n7565 gnd.n210 739.952
R745 gnd.n4423 gnd.n1619 739.952
R746 gnd.n4646 gnd.n1623 739.952
R747 gnd.n4905 gnd.n1377 739.952
R748 gnd.n3057 gnd.n1374 739.952
R749 gnd.n5042 gnd.n1140 739.952
R750 gnd.n5162 gnd.n1071 739.952
R751 gnd.n6748 gnd.n800 670.282
R752 gnd.n7202 gnd.n526 670.282
R753 gnd.n7415 gnd.n399 670.282
R754 gnd.n2654 gnd.n2648 670.282
R755 gnd.n6748 gnd.n6747 585
R756 gnd.n6749 gnd.n6748 585
R757 gnd.n6746 gnd.n802 585
R758 gnd.n802 gnd.n801 585
R759 gnd.n6745 gnd.n6744 585
R760 gnd.n6744 gnd.n6743 585
R761 gnd.n807 gnd.n806 585
R762 gnd.n6742 gnd.n807 585
R763 gnd.n6740 gnd.n6739 585
R764 gnd.n6741 gnd.n6740 585
R765 gnd.n6738 gnd.n809 585
R766 gnd.n809 gnd.n808 585
R767 gnd.n6737 gnd.n6736 585
R768 gnd.n6736 gnd.n6735 585
R769 gnd.n815 gnd.n814 585
R770 gnd.n6734 gnd.n815 585
R771 gnd.n6732 gnd.n6731 585
R772 gnd.n6733 gnd.n6732 585
R773 gnd.n6730 gnd.n817 585
R774 gnd.n817 gnd.n816 585
R775 gnd.n6729 gnd.n6728 585
R776 gnd.n6728 gnd.n6727 585
R777 gnd.n823 gnd.n822 585
R778 gnd.n6726 gnd.n823 585
R779 gnd.n6724 gnd.n6723 585
R780 gnd.n6725 gnd.n6724 585
R781 gnd.n6722 gnd.n825 585
R782 gnd.n825 gnd.n824 585
R783 gnd.n6721 gnd.n6720 585
R784 gnd.n6720 gnd.n6719 585
R785 gnd.n831 gnd.n830 585
R786 gnd.n6718 gnd.n831 585
R787 gnd.n6716 gnd.n6715 585
R788 gnd.n6717 gnd.n6716 585
R789 gnd.n6714 gnd.n833 585
R790 gnd.n833 gnd.n832 585
R791 gnd.n6713 gnd.n6712 585
R792 gnd.n6712 gnd.n6711 585
R793 gnd.n839 gnd.n838 585
R794 gnd.n6710 gnd.n839 585
R795 gnd.n6708 gnd.n6707 585
R796 gnd.n6709 gnd.n6708 585
R797 gnd.n6706 gnd.n841 585
R798 gnd.n841 gnd.n840 585
R799 gnd.n6705 gnd.n6704 585
R800 gnd.n6704 gnd.n6703 585
R801 gnd.n847 gnd.n846 585
R802 gnd.n6702 gnd.n847 585
R803 gnd.n6700 gnd.n6699 585
R804 gnd.n6701 gnd.n6700 585
R805 gnd.n6698 gnd.n849 585
R806 gnd.n849 gnd.n848 585
R807 gnd.n6697 gnd.n6696 585
R808 gnd.n6696 gnd.n6695 585
R809 gnd.n855 gnd.n854 585
R810 gnd.n6694 gnd.n855 585
R811 gnd.n6692 gnd.n6691 585
R812 gnd.n6693 gnd.n6692 585
R813 gnd.n6690 gnd.n857 585
R814 gnd.n857 gnd.n856 585
R815 gnd.n6689 gnd.n6688 585
R816 gnd.n6688 gnd.n6687 585
R817 gnd.n863 gnd.n862 585
R818 gnd.n6686 gnd.n863 585
R819 gnd.n6684 gnd.n6683 585
R820 gnd.n6685 gnd.n6684 585
R821 gnd.n6682 gnd.n865 585
R822 gnd.n865 gnd.n864 585
R823 gnd.n6681 gnd.n6680 585
R824 gnd.n6680 gnd.n6679 585
R825 gnd.n871 gnd.n870 585
R826 gnd.n6678 gnd.n871 585
R827 gnd.n6676 gnd.n6675 585
R828 gnd.n6677 gnd.n6676 585
R829 gnd.n6674 gnd.n873 585
R830 gnd.n873 gnd.n872 585
R831 gnd.n6673 gnd.n6672 585
R832 gnd.n6672 gnd.n6671 585
R833 gnd.n879 gnd.n878 585
R834 gnd.n6670 gnd.n879 585
R835 gnd.n6668 gnd.n6667 585
R836 gnd.n6669 gnd.n6668 585
R837 gnd.n6666 gnd.n881 585
R838 gnd.n881 gnd.n880 585
R839 gnd.n6665 gnd.n6664 585
R840 gnd.n6664 gnd.n6663 585
R841 gnd.n887 gnd.n886 585
R842 gnd.n6662 gnd.n887 585
R843 gnd.n6660 gnd.n6659 585
R844 gnd.n6661 gnd.n6660 585
R845 gnd.n6658 gnd.n889 585
R846 gnd.n889 gnd.n888 585
R847 gnd.n6657 gnd.n6656 585
R848 gnd.n6656 gnd.n6655 585
R849 gnd.n895 gnd.n894 585
R850 gnd.n6654 gnd.n895 585
R851 gnd.n6652 gnd.n6651 585
R852 gnd.n6653 gnd.n6652 585
R853 gnd.n6650 gnd.n897 585
R854 gnd.n897 gnd.n896 585
R855 gnd.n6649 gnd.n6648 585
R856 gnd.n6648 gnd.n6647 585
R857 gnd.n903 gnd.n902 585
R858 gnd.n6646 gnd.n903 585
R859 gnd.n6644 gnd.n6643 585
R860 gnd.n6645 gnd.n6644 585
R861 gnd.n6642 gnd.n905 585
R862 gnd.n905 gnd.n904 585
R863 gnd.n6641 gnd.n6640 585
R864 gnd.n6640 gnd.n6639 585
R865 gnd.n911 gnd.n910 585
R866 gnd.n6638 gnd.n911 585
R867 gnd.n6636 gnd.n6635 585
R868 gnd.n6637 gnd.n6636 585
R869 gnd.n6634 gnd.n913 585
R870 gnd.n913 gnd.n912 585
R871 gnd.n6633 gnd.n6632 585
R872 gnd.n6632 gnd.n6631 585
R873 gnd.n919 gnd.n918 585
R874 gnd.n6630 gnd.n919 585
R875 gnd.n6628 gnd.n6627 585
R876 gnd.n6629 gnd.n6628 585
R877 gnd.n6626 gnd.n921 585
R878 gnd.n921 gnd.n920 585
R879 gnd.n6625 gnd.n6624 585
R880 gnd.n6624 gnd.n6623 585
R881 gnd.n927 gnd.n926 585
R882 gnd.n6622 gnd.n927 585
R883 gnd.n6620 gnd.n6619 585
R884 gnd.n6621 gnd.n6620 585
R885 gnd.n6618 gnd.n929 585
R886 gnd.n929 gnd.n928 585
R887 gnd.n6617 gnd.n6616 585
R888 gnd.n6616 gnd.n6615 585
R889 gnd.n935 gnd.n934 585
R890 gnd.n6614 gnd.n935 585
R891 gnd.n6612 gnd.n6611 585
R892 gnd.n6613 gnd.n6612 585
R893 gnd.n6610 gnd.n937 585
R894 gnd.n937 gnd.n936 585
R895 gnd.n6609 gnd.n6608 585
R896 gnd.n6608 gnd.n6607 585
R897 gnd.n943 gnd.n942 585
R898 gnd.n6606 gnd.n943 585
R899 gnd.n6604 gnd.n6603 585
R900 gnd.n6605 gnd.n6604 585
R901 gnd.n6602 gnd.n945 585
R902 gnd.n945 gnd.n944 585
R903 gnd.n6601 gnd.n6600 585
R904 gnd.n6600 gnd.n6599 585
R905 gnd.n951 gnd.n950 585
R906 gnd.n6598 gnd.n951 585
R907 gnd.n6596 gnd.n6595 585
R908 gnd.n6597 gnd.n6596 585
R909 gnd.n6594 gnd.n953 585
R910 gnd.n953 gnd.n952 585
R911 gnd.n6593 gnd.n6592 585
R912 gnd.n6592 gnd.n6591 585
R913 gnd.n959 gnd.n958 585
R914 gnd.n6590 gnd.n959 585
R915 gnd.n6588 gnd.n6587 585
R916 gnd.n6589 gnd.n6588 585
R917 gnd.n6586 gnd.n961 585
R918 gnd.n961 gnd.n960 585
R919 gnd.n6585 gnd.n6584 585
R920 gnd.n6584 gnd.n6583 585
R921 gnd.n967 gnd.n966 585
R922 gnd.n6582 gnd.n967 585
R923 gnd.n800 gnd.n799 585
R924 gnd.n6750 gnd.n800 585
R925 gnd.n6753 gnd.n6752 585
R926 gnd.n6752 gnd.n6751 585
R927 gnd.n797 gnd.n796 585
R928 gnd.n796 gnd.n795 585
R929 gnd.n6758 gnd.n6757 585
R930 gnd.n6759 gnd.n6758 585
R931 gnd.n794 gnd.n793 585
R932 gnd.n6760 gnd.n794 585
R933 gnd.n6763 gnd.n6762 585
R934 gnd.n6762 gnd.n6761 585
R935 gnd.n791 gnd.n790 585
R936 gnd.n790 gnd.n789 585
R937 gnd.n6768 gnd.n6767 585
R938 gnd.n6769 gnd.n6768 585
R939 gnd.n788 gnd.n787 585
R940 gnd.n6770 gnd.n788 585
R941 gnd.n6773 gnd.n6772 585
R942 gnd.n6772 gnd.n6771 585
R943 gnd.n785 gnd.n784 585
R944 gnd.n784 gnd.n783 585
R945 gnd.n6778 gnd.n6777 585
R946 gnd.n6779 gnd.n6778 585
R947 gnd.n782 gnd.n781 585
R948 gnd.n6780 gnd.n782 585
R949 gnd.n6783 gnd.n6782 585
R950 gnd.n6782 gnd.n6781 585
R951 gnd.n779 gnd.n778 585
R952 gnd.n778 gnd.n777 585
R953 gnd.n6788 gnd.n6787 585
R954 gnd.n6789 gnd.n6788 585
R955 gnd.n776 gnd.n775 585
R956 gnd.n6790 gnd.n776 585
R957 gnd.n6793 gnd.n6792 585
R958 gnd.n6792 gnd.n6791 585
R959 gnd.n773 gnd.n772 585
R960 gnd.n772 gnd.n771 585
R961 gnd.n6798 gnd.n6797 585
R962 gnd.n6799 gnd.n6798 585
R963 gnd.n770 gnd.n769 585
R964 gnd.n6800 gnd.n770 585
R965 gnd.n6803 gnd.n6802 585
R966 gnd.n6802 gnd.n6801 585
R967 gnd.n767 gnd.n766 585
R968 gnd.n766 gnd.n765 585
R969 gnd.n6808 gnd.n6807 585
R970 gnd.n6809 gnd.n6808 585
R971 gnd.n764 gnd.n763 585
R972 gnd.n6810 gnd.n764 585
R973 gnd.n6813 gnd.n6812 585
R974 gnd.n6812 gnd.n6811 585
R975 gnd.n761 gnd.n760 585
R976 gnd.n760 gnd.n759 585
R977 gnd.n6818 gnd.n6817 585
R978 gnd.n6819 gnd.n6818 585
R979 gnd.n758 gnd.n757 585
R980 gnd.n6820 gnd.n758 585
R981 gnd.n6823 gnd.n6822 585
R982 gnd.n6822 gnd.n6821 585
R983 gnd.n755 gnd.n754 585
R984 gnd.n754 gnd.n753 585
R985 gnd.n6828 gnd.n6827 585
R986 gnd.n6829 gnd.n6828 585
R987 gnd.n752 gnd.n751 585
R988 gnd.n6830 gnd.n752 585
R989 gnd.n6833 gnd.n6832 585
R990 gnd.n6832 gnd.n6831 585
R991 gnd.n749 gnd.n748 585
R992 gnd.n748 gnd.n747 585
R993 gnd.n6838 gnd.n6837 585
R994 gnd.n6839 gnd.n6838 585
R995 gnd.n746 gnd.n745 585
R996 gnd.n6840 gnd.n746 585
R997 gnd.n6843 gnd.n6842 585
R998 gnd.n6842 gnd.n6841 585
R999 gnd.n743 gnd.n742 585
R1000 gnd.n742 gnd.n741 585
R1001 gnd.n6848 gnd.n6847 585
R1002 gnd.n6849 gnd.n6848 585
R1003 gnd.n740 gnd.n739 585
R1004 gnd.n6850 gnd.n740 585
R1005 gnd.n6853 gnd.n6852 585
R1006 gnd.n6852 gnd.n6851 585
R1007 gnd.n737 gnd.n736 585
R1008 gnd.n736 gnd.n735 585
R1009 gnd.n6858 gnd.n6857 585
R1010 gnd.n6859 gnd.n6858 585
R1011 gnd.n734 gnd.n733 585
R1012 gnd.n6860 gnd.n734 585
R1013 gnd.n6863 gnd.n6862 585
R1014 gnd.n6862 gnd.n6861 585
R1015 gnd.n731 gnd.n730 585
R1016 gnd.n730 gnd.n729 585
R1017 gnd.n6868 gnd.n6867 585
R1018 gnd.n6869 gnd.n6868 585
R1019 gnd.n728 gnd.n727 585
R1020 gnd.n6870 gnd.n728 585
R1021 gnd.n6873 gnd.n6872 585
R1022 gnd.n6872 gnd.n6871 585
R1023 gnd.n725 gnd.n724 585
R1024 gnd.n724 gnd.n723 585
R1025 gnd.n6878 gnd.n6877 585
R1026 gnd.n6879 gnd.n6878 585
R1027 gnd.n722 gnd.n721 585
R1028 gnd.n6880 gnd.n722 585
R1029 gnd.n6883 gnd.n6882 585
R1030 gnd.n6882 gnd.n6881 585
R1031 gnd.n719 gnd.n718 585
R1032 gnd.n718 gnd.n717 585
R1033 gnd.n6888 gnd.n6887 585
R1034 gnd.n6889 gnd.n6888 585
R1035 gnd.n716 gnd.n715 585
R1036 gnd.n6890 gnd.n716 585
R1037 gnd.n6893 gnd.n6892 585
R1038 gnd.n6892 gnd.n6891 585
R1039 gnd.n713 gnd.n712 585
R1040 gnd.n712 gnd.n711 585
R1041 gnd.n6898 gnd.n6897 585
R1042 gnd.n6899 gnd.n6898 585
R1043 gnd.n710 gnd.n709 585
R1044 gnd.n6900 gnd.n710 585
R1045 gnd.n6903 gnd.n6902 585
R1046 gnd.n6902 gnd.n6901 585
R1047 gnd.n707 gnd.n706 585
R1048 gnd.n706 gnd.n705 585
R1049 gnd.n6908 gnd.n6907 585
R1050 gnd.n6909 gnd.n6908 585
R1051 gnd.n704 gnd.n703 585
R1052 gnd.n6910 gnd.n704 585
R1053 gnd.n6913 gnd.n6912 585
R1054 gnd.n6912 gnd.n6911 585
R1055 gnd.n701 gnd.n700 585
R1056 gnd.n700 gnd.n699 585
R1057 gnd.n6918 gnd.n6917 585
R1058 gnd.n6919 gnd.n6918 585
R1059 gnd.n698 gnd.n697 585
R1060 gnd.n6920 gnd.n698 585
R1061 gnd.n6923 gnd.n6922 585
R1062 gnd.n6922 gnd.n6921 585
R1063 gnd.n695 gnd.n694 585
R1064 gnd.n694 gnd.n693 585
R1065 gnd.n6928 gnd.n6927 585
R1066 gnd.n6929 gnd.n6928 585
R1067 gnd.n692 gnd.n691 585
R1068 gnd.n6930 gnd.n692 585
R1069 gnd.n6933 gnd.n6932 585
R1070 gnd.n6932 gnd.n6931 585
R1071 gnd.n689 gnd.n688 585
R1072 gnd.n688 gnd.n687 585
R1073 gnd.n6938 gnd.n6937 585
R1074 gnd.n6939 gnd.n6938 585
R1075 gnd.n686 gnd.n685 585
R1076 gnd.n6940 gnd.n686 585
R1077 gnd.n6943 gnd.n6942 585
R1078 gnd.n6942 gnd.n6941 585
R1079 gnd.n683 gnd.n682 585
R1080 gnd.n682 gnd.n681 585
R1081 gnd.n6948 gnd.n6947 585
R1082 gnd.n6949 gnd.n6948 585
R1083 gnd.n680 gnd.n679 585
R1084 gnd.n6950 gnd.n680 585
R1085 gnd.n6953 gnd.n6952 585
R1086 gnd.n6952 gnd.n6951 585
R1087 gnd.n677 gnd.n676 585
R1088 gnd.n676 gnd.n675 585
R1089 gnd.n6958 gnd.n6957 585
R1090 gnd.n6959 gnd.n6958 585
R1091 gnd.n674 gnd.n673 585
R1092 gnd.n6960 gnd.n674 585
R1093 gnd.n6963 gnd.n6962 585
R1094 gnd.n6962 gnd.n6961 585
R1095 gnd.n671 gnd.n670 585
R1096 gnd.n670 gnd.n669 585
R1097 gnd.n6968 gnd.n6967 585
R1098 gnd.n6969 gnd.n6968 585
R1099 gnd.n668 gnd.n667 585
R1100 gnd.n6970 gnd.n668 585
R1101 gnd.n6973 gnd.n6972 585
R1102 gnd.n6972 gnd.n6971 585
R1103 gnd.n665 gnd.n664 585
R1104 gnd.n664 gnd.n663 585
R1105 gnd.n6978 gnd.n6977 585
R1106 gnd.n6979 gnd.n6978 585
R1107 gnd.n662 gnd.n661 585
R1108 gnd.n6980 gnd.n662 585
R1109 gnd.n6983 gnd.n6982 585
R1110 gnd.n6982 gnd.n6981 585
R1111 gnd.n659 gnd.n658 585
R1112 gnd.n658 gnd.n657 585
R1113 gnd.n6988 gnd.n6987 585
R1114 gnd.n6989 gnd.n6988 585
R1115 gnd.n656 gnd.n655 585
R1116 gnd.n6990 gnd.n656 585
R1117 gnd.n6993 gnd.n6992 585
R1118 gnd.n6992 gnd.n6991 585
R1119 gnd.n653 gnd.n652 585
R1120 gnd.n652 gnd.n651 585
R1121 gnd.n6998 gnd.n6997 585
R1122 gnd.n6999 gnd.n6998 585
R1123 gnd.n650 gnd.n649 585
R1124 gnd.n7000 gnd.n650 585
R1125 gnd.n7003 gnd.n7002 585
R1126 gnd.n7002 gnd.n7001 585
R1127 gnd.n647 gnd.n646 585
R1128 gnd.n646 gnd.n645 585
R1129 gnd.n7008 gnd.n7007 585
R1130 gnd.n7009 gnd.n7008 585
R1131 gnd.n644 gnd.n643 585
R1132 gnd.n7010 gnd.n644 585
R1133 gnd.n7013 gnd.n7012 585
R1134 gnd.n7012 gnd.n7011 585
R1135 gnd.n641 gnd.n640 585
R1136 gnd.n640 gnd.n639 585
R1137 gnd.n7018 gnd.n7017 585
R1138 gnd.n7019 gnd.n7018 585
R1139 gnd.n638 gnd.n637 585
R1140 gnd.n7020 gnd.n638 585
R1141 gnd.n7023 gnd.n7022 585
R1142 gnd.n7022 gnd.n7021 585
R1143 gnd.n635 gnd.n634 585
R1144 gnd.n634 gnd.n633 585
R1145 gnd.n7028 gnd.n7027 585
R1146 gnd.n7029 gnd.n7028 585
R1147 gnd.n632 gnd.n631 585
R1148 gnd.n7030 gnd.n632 585
R1149 gnd.n7033 gnd.n7032 585
R1150 gnd.n7032 gnd.n7031 585
R1151 gnd.n629 gnd.n628 585
R1152 gnd.n628 gnd.n627 585
R1153 gnd.n7038 gnd.n7037 585
R1154 gnd.n7039 gnd.n7038 585
R1155 gnd.n626 gnd.n625 585
R1156 gnd.n7040 gnd.n626 585
R1157 gnd.n7043 gnd.n7042 585
R1158 gnd.n7042 gnd.n7041 585
R1159 gnd.n623 gnd.n622 585
R1160 gnd.n622 gnd.n621 585
R1161 gnd.n7048 gnd.n7047 585
R1162 gnd.n7049 gnd.n7048 585
R1163 gnd.n620 gnd.n619 585
R1164 gnd.n7050 gnd.n620 585
R1165 gnd.n7053 gnd.n7052 585
R1166 gnd.n7052 gnd.n7051 585
R1167 gnd.n617 gnd.n616 585
R1168 gnd.n616 gnd.n615 585
R1169 gnd.n7058 gnd.n7057 585
R1170 gnd.n7059 gnd.n7058 585
R1171 gnd.n614 gnd.n613 585
R1172 gnd.n7060 gnd.n614 585
R1173 gnd.n7063 gnd.n7062 585
R1174 gnd.n7062 gnd.n7061 585
R1175 gnd.n611 gnd.n610 585
R1176 gnd.n610 gnd.n609 585
R1177 gnd.n7068 gnd.n7067 585
R1178 gnd.n7069 gnd.n7068 585
R1179 gnd.n608 gnd.n607 585
R1180 gnd.n7070 gnd.n608 585
R1181 gnd.n7073 gnd.n7072 585
R1182 gnd.n7072 gnd.n7071 585
R1183 gnd.n605 gnd.n604 585
R1184 gnd.n604 gnd.n603 585
R1185 gnd.n7078 gnd.n7077 585
R1186 gnd.n7079 gnd.n7078 585
R1187 gnd.n602 gnd.n601 585
R1188 gnd.n7080 gnd.n602 585
R1189 gnd.n7083 gnd.n7082 585
R1190 gnd.n7082 gnd.n7081 585
R1191 gnd.n599 gnd.n598 585
R1192 gnd.n598 gnd.n597 585
R1193 gnd.n7088 gnd.n7087 585
R1194 gnd.n7089 gnd.n7088 585
R1195 gnd.n596 gnd.n595 585
R1196 gnd.n7090 gnd.n596 585
R1197 gnd.n7093 gnd.n7092 585
R1198 gnd.n7092 gnd.n7091 585
R1199 gnd.n593 gnd.n592 585
R1200 gnd.n592 gnd.n591 585
R1201 gnd.n7098 gnd.n7097 585
R1202 gnd.n7099 gnd.n7098 585
R1203 gnd.n590 gnd.n589 585
R1204 gnd.n7100 gnd.n590 585
R1205 gnd.n7103 gnd.n7102 585
R1206 gnd.n7102 gnd.n7101 585
R1207 gnd.n587 gnd.n586 585
R1208 gnd.n586 gnd.n585 585
R1209 gnd.n7108 gnd.n7107 585
R1210 gnd.n7109 gnd.n7108 585
R1211 gnd.n584 gnd.n583 585
R1212 gnd.n7110 gnd.n584 585
R1213 gnd.n7113 gnd.n7112 585
R1214 gnd.n7112 gnd.n7111 585
R1215 gnd.n581 gnd.n580 585
R1216 gnd.n580 gnd.n579 585
R1217 gnd.n7118 gnd.n7117 585
R1218 gnd.n7119 gnd.n7118 585
R1219 gnd.n578 gnd.n577 585
R1220 gnd.n7120 gnd.n578 585
R1221 gnd.n7123 gnd.n7122 585
R1222 gnd.n7122 gnd.n7121 585
R1223 gnd.n575 gnd.n574 585
R1224 gnd.n574 gnd.n573 585
R1225 gnd.n7128 gnd.n7127 585
R1226 gnd.n7129 gnd.n7128 585
R1227 gnd.n572 gnd.n571 585
R1228 gnd.n7130 gnd.n572 585
R1229 gnd.n7133 gnd.n7132 585
R1230 gnd.n7132 gnd.n7131 585
R1231 gnd.n569 gnd.n568 585
R1232 gnd.n568 gnd.n567 585
R1233 gnd.n7138 gnd.n7137 585
R1234 gnd.n7139 gnd.n7138 585
R1235 gnd.n566 gnd.n565 585
R1236 gnd.n7140 gnd.n566 585
R1237 gnd.n7143 gnd.n7142 585
R1238 gnd.n7142 gnd.n7141 585
R1239 gnd.n563 gnd.n562 585
R1240 gnd.n562 gnd.n561 585
R1241 gnd.n7148 gnd.n7147 585
R1242 gnd.n7149 gnd.n7148 585
R1243 gnd.n560 gnd.n559 585
R1244 gnd.n7150 gnd.n560 585
R1245 gnd.n7153 gnd.n7152 585
R1246 gnd.n7152 gnd.n7151 585
R1247 gnd.n557 gnd.n556 585
R1248 gnd.n556 gnd.n555 585
R1249 gnd.n7158 gnd.n7157 585
R1250 gnd.n7159 gnd.n7158 585
R1251 gnd.n554 gnd.n553 585
R1252 gnd.n7160 gnd.n554 585
R1253 gnd.n7163 gnd.n7162 585
R1254 gnd.n7162 gnd.n7161 585
R1255 gnd.n551 gnd.n550 585
R1256 gnd.n550 gnd.n549 585
R1257 gnd.n7168 gnd.n7167 585
R1258 gnd.n7169 gnd.n7168 585
R1259 gnd.n548 gnd.n547 585
R1260 gnd.n7170 gnd.n548 585
R1261 gnd.n7173 gnd.n7172 585
R1262 gnd.n7172 gnd.n7171 585
R1263 gnd.n545 gnd.n544 585
R1264 gnd.n544 gnd.n543 585
R1265 gnd.n7178 gnd.n7177 585
R1266 gnd.n7179 gnd.n7178 585
R1267 gnd.n542 gnd.n541 585
R1268 gnd.n7180 gnd.n542 585
R1269 gnd.n7183 gnd.n7182 585
R1270 gnd.n7182 gnd.n7181 585
R1271 gnd.n539 gnd.n538 585
R1272 gnd.n538 gnd.n537 585
R1273 gnd.n7188 gnd.n7187 585
R1274 gnd.n7189 gnd.n7188 585
R1275 gnd.n536 gnd.n535 585
R1276 gnd.n7190 gnd.n536 585
R1277 gnd.n7193 gnd.n7192 585
R1278 gnd.n7192 gnd.n7191 585
R1279 gnd.n533 gnd.n532 585
R1280 gnd.n532 gnd.n531 585
R1281 gnd.n7198 gnd.n7197 585
R1282 gnd.n7199 gnd.n7198 585
R1283 gnd.n530 gnd.n529 585
R1284 gnd.n7200 gnd.n530 585
R1285 gnd.n7203 gnd.n7202 585
R1286 gnd.n7202 gnd.n7201 585
R1287 gnd.n7414 gnd.n403 585
R1288 gnd.n7414 gnd.n7413 585
R1289 gnd.n7408 gnd.n404 585
R1290 gnd.n7412 gnd.n404 585
R1291 gnd.n7410 gnd.n7409 585
R1292 gnd.n7411 gnd.n7410 585
R1293 gnd.n407 gnd.n406 585
R1294 gnd.n406 gnd.n405 585
R1295 gnd.n7403 gnd.n7402 585
R1296 gnd.n7402 gnd.n7401 585
R1297 gnd.n410 gnd.n409 585
R1298 gnd.n7400 gnd.n410 585
R1299 gnd.n7398 gnd.n7397 585
R1300 gnd.n7399 gnd.n7398 585
R1301 gnd.n413 gnd.n412 585
R1302 gnd.n412 gnd.n411 585
R1303 gnd.n7393 gnd.n7392 585
R1304 gnd.n7392 gnd.n7391 585
R1305 gnd.n416 gnd.n415 585
R1306 gnd.n7390 gnd.n416 585
R1307 gnd.n7388 gnd.n7387 585
R1308 gnd.n7389 gnd.n7388 585
R1309 gnd.n419 gnd.n418 585
R1310 gnd.n418 gnd.n417 585
R1311 gnd.n7383 gnd.n7382 585
R1312 gnd.n7382 gnd.n7381 585
R1313 gnd.n422 gnd.n421 585
R1314 gnd.n7380 gnd.n422 585
R1315 gnd.n7378 gnd.n7377 585
R1316 gnd.n7379 gnd.n7378 585
R1317 gnd.n425 gnd.n424 585
R1318 gnd.n424 gnd.n423 585
R1319 gnd.n7373 gnd.n7372 585
R1320 gnd.n7372 gnd.n7371 585
R1321 gnd.n428 gnd.n427 585
R1322 gnd.n7370 gnd.n428 585
R1323 gnd.n7368 gnd.n7367 585
R1324 gnd.n7369 gnd.n7368 585
R1325 gnd.n431 gnd.n430 585
R1326 gnd.n430 gnd.n429 585
R1327 gnd.n7363 gnd.n7362 585
R1328 gnd.n7362 gnd.n7361 585
R1329 gnd.n434 gnd.n433 585
R1330 gnd.n7360 gnd.n434 585
R1331 gnd.n7358 gnd.n7357 585
R1332 gnd.n7359 gnd.n7358 585
R1333 gnd.n437 gnd.n436 585
R1334 gnd.n436 gnd.n435 585
R1335 gnd.n7353 gnd.n7352 585
R1336 gnd.n7352 gnd.n7351 585
R1337 gnd.n440 gnd.n439 585
R1338 gnd.n7350 gnd.n440 585
R1339 gnd.n7348 gnd.n7347 585
R1340 gnd.n7349 gnd.n7348 585
R1341 gnd.n443 gnd.n442 585
R1342 gnd.n442 gnd.n441 585
R1343 gnd.n7343 gnd.n7342 585
R1344 gnd.n7342 gnd.n7341 585
R1345 gnd.n446 gnd.n445 585
R1346 gnd.n7340 gnd.n446 585
R1347 gnd.n7338 gnd.n7337 585
R1348 gnd.n7339 gnd.n7338 585
R1349 gnd.n449 gnd.n448 585
R1350 gnd.n448 gnd.n447 585
R1351 gnd.n7333 gnd.n7332 585
R1352 gnd.n7332 gnd.n7331 585
R1353 gnd.n452 gnd.n451 585
R1354 gnd.n7330 gnd.n452 585
R1355 gnd.n7328 gnd.n7327 585
R1356 gnd.n7329 gnd.n7328 585
R1357 gnd.n455 gnd.n454 585
R1358 gnd.n454 gnd.n453 585
R1359 gnd.n7323 gnd.n7322 585
R1360 gnd.n7322 gnd.n7321 585
R1361 gnd.n458 gnd.n457 585
R1362 gnd.n7320 gnd.n458 585
R1363 gnd.n7318 gnd.n7317 585
R1364 gnd.n7319 gnd.n7318 585
R1365 gnd.n461 gnd.n460 585
R1366 gnd.n460 gnd.n459 585
R1367 gnd.n7313 gnd.n7312 585
R1368 gnd.n7312 gnd.n7311 585
R1369 gnd.n464 gnd.n463 585
R1370 gnd.n7310 gnd.n464 585
R1371 gnd.n7308 gnd.n7307 585
R1372 gnd.n7309 gnd.n7308 585
R1373 gnd.n467 gnd.n466 585
R1374 gnd.n466 gnd.n465 585
R1375 gnd.n7303 gnd.n7302 585
R1376 gnd.n7302 gnd.n7301 585
R1377 gnd.n470 gnd.n469 585
R1378 gnd.n7300 gnd.n470 585
R1379 gnd.n7298 gnd.n7297 585
R1380 gnd.n7299 gnd.n7298 585
R1381 gnd.n473 gnd.n472 585
R1382 gnd.n472 gnd.n471 585
R1383 gnd.n7293 gnd.n7292 585
R1384 gnd.n7292 gnd.n7291 585
R1385 gnd.n476 gnd.n475 585
R1386 gnd.n7290 gnd.n476 585
R1387 gnd.n7288 gnd.n7287 585
R1388 gnd.n7289 gnd.n7288 585
R1389 gnd.n479 gnd.n478 585
R1390 gnd.n478 gnd.n477 585
R1391 gnd.n7283 gnd.n7282 585
R1392 gnd.n7282 gnd.n7281 585
R1393 gnd.n482 gnd.n481 585
R1394 gnd.n7280 gnd.n482 585
R1395 gnd.n7278 gnd.n7277 585
R1396 gnd.n7279 gnd.n7278 585
R1397 gnd.n485 gnd.n484 585
R1398 gnd.n484 gnd.n483 585
R1399 gnd.n7273 gnd.n7272 585
R1400 gnd.n7272 gnd.n7271 585
R1401 gnd.n488 gnd.n487 585
R1402 gnd.n7270 gnd.n488 585
R1403 gnd.n7268 gnd.n7267 585
R1404 gnd.n7269 gnd.n7268 585
R1405 gnd.n491 gnd.n490 585
R1406 gnd.n490 gnd.n489 585
R1407 gnd.n7263 gnd.n7262 585
R1408 gnd.n7262 gnd.n7261 585
R1409 gnd.n494 gnd.n493 585
R1410 gnd.n7260 gnd.n494 585
R1411 gnd.n7258 gnd.n7257 585
R1412 gnd.n7259 gnd.n7258 585
R1413 gnd.n497 gnd.n496 585
R1414 gnd.n496 gnd.n495 585
R1415 gnd.n7253 gnd.n7252 585
R1416 gnd.n7252 gnd.n7251 585
R1417 gnd.n500 gnd.n499 585
R1418 gnd.n7250 gnd.n500 585
R1419 gnd.n7248 gnd.n7247 585
R1420 gnd.n7249 gnd.n7248 585
R1421 gnd.n503 gnd.n502 585
R1422 gnd.n502 gnd.n501 585
R1423 gnd.n7243 gnd.n7242 585
R1424 gnd.n7242 gnd.n7241 585
R1425 gnd.n506 gnd.n505 585
R1426 gnd.n7240 gnd.n506 585
R1427 gnd.n7238 gnd.n7237 585
R1428 gnd.n7239 gnd.n7238 585
R1429 gnd.n509 gnd.n508 585
R1430 gnd.n508 gnd.n507 585
R1431 gnd.n7233 gnd.n7232 585
R1432 gnd.n7232 gnd.n7231 585
R1433 gnd.n512 gnd.n511 585
R1434 gnd.n7230 gnd.n512 585
R1435 gnd.n7228 gnd.n7227 585
R1436 gnd.n7229 gnd.n7228 585
R1437 gnd.n515 gnd.n514 585
R1438 gnd.n514 gnd.n513 585
R1439 gnd.n7223 gnd.n7222 585
R1440 gnd.n7222 gnd.n7221 585
R1441 gnd.n518 gnd.n517 585
R1442 gnd.n7220 gnd.n518 585
R1443 gnd.n7218 gnd.n7217 585
R1444 gnd.n7219 gnd.n7218 585
R1445 gnd.n521 gnd.n520 585
R1446 gnd.n520 gnd.n519 585
R1447 gnd.n7213 gnd.n7212 585
R1448 gnd.n7212 gnd.n7211 585
R1449 gnd.n524 gnd.n523 585
R1450 gnd.n7210 gnd.n524 585
R1451 gnd.n7208 gnd.n7207 585
R1452 gnd.n7209 gnd.n7208 585
R1453 gnd.n527 gnd.n526 585
R1454 gnd.n526 gnd.n525 585
R1455 gnd.n4908 gnd.n4907 585
R1456 gnd.n4907 gnd.n4906 585
R1457 gnd.n4909 gnd.n1368 585
R1458 gnd.n2883 gnd.n1368 585
R1459 gnd.n4911 gnd.n4910 585
R1460 gnd.n4912 gnd.n4911 585
R1461 gnd.n1352 gnd.n1351 585
R1462 gnd.n2876 gnd.n1352 585
R1463 gnd.n4920 gnd.n4919 585
R1464 gnd.n4919 gnd.n4918 585
R1465 gnd.n4921 gnd.n1347 585
R1466 gnd.n2871 gnd.n1347 585
R1467 gnd.n4923 gnd.n4922 585
R1468 gnd.n4924 gnd.n4923 585
R1469 gnd.n1332 gnd.n1331 585
R1470 gnd.n2898 gnd.n1332 585
R1471 gnd.n4932 gnd.n4931 585
R1472 gnd.n4931 gnd.n4930 585
R1473 gnd.n4933 gnd.n1327 585
R1474 gnd.n2864 gnd.n1327 585
R1475 gnd.n4935 gnd.n4934 585
R1476 gnd.n4936 gnd.n4935 585
R1477 gnd.n1312 gnd.n1311 585
R1478 gnd.n2856 gnd.n1312 585
R1479 gnd.n4944 gnd.n4943 585
R1480 gnd.n4943 gnd.n4942 585
R1481 gnd.n4945 gnd.n1307 585
R1482 gnd.n2849 gnd.n1307 585
R1483 gnd.n4947 gnd.n4946 585
R1484 gnd.n4948 gnd.n4947 585
R1485 gnd.n1292 gnd.n1291 585
R1486 gnd.n2841 gnd.n1292 585
R1487 gnd.n4956 gnd.n4955 585
R1488 gnd.n4955 gnd.n4954 585
R1489 gnd.n4957 gnd.n1287 585
R1490 gnd.n2788 gnd.n1287 585
R1491 gnd.n4959 gnd.n4958 585
R1492 gnd.n4960 gnd.n4959 585
R1493 gnd.n1273 gnd.n1272 585
R1494 gnd.n2779 gnd.n1273 585
R1495 gnd.n4968 gnd.n4967 585
R1496 gnd.n4967 gnd.n4966 585
R1497 gnd.n4969 gnd.n1267 585
R1498 gnd.n2773 gnd.n1267 585
R1499 gnd.n4971 gnd.n4970 585
R1500 gnd.n4972 gnd.n4971 585
R1501 gnd.n1268 gnd.n1266 585
R1502 gnd.n2802 gnd.n1266 585
R1503 gnd.n2768 gnd.n2767 585
R1504 gnd.n2767 gnd.n2766 585
R1505 gnd.n2473 gnd.n2472 585
R1506 gnd.n2761 gnd.n2473 585
R1507 gnd.n2743 gnd.n2742 585
R1508 gnd.n2742 gnd.n2741 585
R1509 gnd.n2744 gnd.n2485 585
R1510 gnd.n2752 gnd.n2485 585
R1511 gnd.n2746 gnd.n2745 585
R1512 gnd.n2747 gnd.n2746 585
R1513 gnd.n2492 gnd.n2491 585
R1514 gnd.n2715 gnd.n2491 585
R1515 gnd.n2721 gnd.n2720 585
R1516 gnd.n2723 gnd.n2721 585
R1517 gnd.n1244 gnd.n1243 585
R1518 gnd.n2503 gnd.n1244 585
R1519 gnd.n4982 gnd.n4981 585
R1520 gnd.n4981 gnd.n4980 585
R1521 gnd.n4983 gnd.n1239 585
R1522 gnd.n2704 gnd.n1239 585
R1523 gnd.n4985 gnd.n4984 585
R1524 gnd.n4986 gnd.n4985 585
R1525 gnd.n1223 gnd.n1222 585
R1526 gnd.n2697 gnd.n1223 585
R1527 gnd.n4994 gnd.n4993 585
R1528 gnd.n4993 gnd.n4992 585
R1529 gnd.n4995 gnd.n1218 585
R1530 gnd.n2688 gnd.n1218 585
R1531 gnd.n4997 gnd.n4996 585
R1532 gnd.n4998 gnd.n4997 585
R1533 gnd.n1203 gnd.n1202 585
R1534 gnd.n2682 gnd.n1203 585
R1535 gnd.n5006 gnd.n5005 585
R1536 gnd.n5005 gnd.n5004 585
R1537 gnd.n5007 gnd.n1198 585
R1538 gnd.n2635 gnd.n1198 585
R1539 gnd.n5009 gnd.n5008 585
R1540 gnd.n5010 gnd.n5009 585
R1541 gnd.n1183 gnd.n1182 585
R1542 gnd.n2629 gnd.n1183 585
R1543 gnd.n5018 gnd.n5017 585
R1544 gnd.n5017 gnd.n5016 585
R1545 gnd.n5019 gnd.n1178 585
R1546 gnd.n1178 gnd.n1177 585
R1547 gnd.n5021 gnd.n5020 585
R1548 gnd.n5022 gnd.n5021 585
R1549 gnd.n1164 gnd.n1163 585
R1550 gnd.n1167 gnd.n1164 585
R1551 gnd.n5030 gnd.n5029 585
R1552 gnd.n5029 gnd.n5028 585
R1553 gnd.n5031 gnd.n1157 585
R1554 gnd.n1157 gnd.n1155 585
R1555 gnd.n5033 gnd.n5032 585
R1556 gnd.n5034 gnd.n5033 585
R1557 gnd.n1159 gnd.n1156 585
R1558 gnd.n1156 gnd.n1152 585
R1559 gnd.n1158 gnd.n1143 585
R1560 gnd.n5040 gnd.n1143 585
R1561 gnd.n2562 gnd.n1137 585
R1562 gnd.n2562 gnd.n1068 585
R1563 gnd.n2564 gnd.n2563 585
R1564 gnd.n2566 gnd.n2565 585
R1565 gnd.n2568 gnd.n2567 585
R1566 gnd.n2572 gnd.n2560 585
R1567 gnd.n2574 gnd.n2573 585
R1568 gnd.n2576 gnd.n2575 585
R1569 gnd.n2578 gnd.n2577 585
R1570 gnd.n2582 gnd.n2558 585
R1571 gnd.n2584 gnd.n2583 585
R1572 gnd.n2586 gnd.n2585 585
R1573 gnd.n2588 gnd.n2587 585
R1574 gnd.n2592 gnd.n2556 585
R1575 gnd.n2594 gnd.n2593 585
R1576 gnd.n2596 gnd.n2595 585
R1577 gnd.n2598 gnd.n2597 585
R1578 gnd.n2553 gnd.n2552 585
R1579 gnd.n2602 gnd.n2554 585
R1580 gnd.n2603 gnd.n2549 585
R1581 gnd.n2604 gnd.n1067 585
R1582 gnd.n5164 gnd.n1067 585
R1583 gnd.n3191 gnd.n3190 585
R1584 gnd.n3188 gnd.n2406 585
R1585 gnd.n3187 gnd.n3186 585
R1586 gnd.n3118 gnd.n2408 585
R1587 gnd.n3127 gnd.n3119 585
R1588 gnd.n3128 gnd.n3116 585
R1589 gnd.n3115 gnd.n3108 585
R1590 gnd.n3135 gnd.n3107 585
R1591 gnd.n3136 gnd.n3106 585
R1592 gnd.n3104 gnd.n3096 585
R1593 gnd.n3143 gnd.n3095 585
R1594 gnd.n3144 gnd.n3093 585
R1595 gnd.n3092 gnd.n3085 585
R1596 gnd.n3151 gnd.n3084 585
R1597 gnd.n3152 gnd.n3083 585
R1598 gnd.n3081 gnd.n3073 585
R1599 gnd.n3159 gnd.n3072 585
R1600 gnd.n3160 gnd.n3070 585
R1601 gnd.n3069 gnd.n1372 585
R1602 gnd.n1381 gnd.n1372 585
R1603 gnd.n2885 gnd.n1375 585
R1604 gnd.n4906 gnd.n1375 585
R1605 gnd.n2886 gnd.n2884 585
R1606 gnd.n2884 gnd.n2883 585
R1607 gnd.n2437 gnd.n1366 585
R1608 gnd.n4912 gnd.n1366 585
R1609 gnd.n2890 gnd.n2436 585
R1610 gnd.n2876 gnd.n2436 585
R1611 gnd.n2891 gnd.n1355 585
R1612 gnd.n4918 gnd.n1355 585
R1613 gnd.n2892 gnd.n2435 585
R1614 gnd.n2871 gnd.n2435 585
R1615 gnd.n2432 gnd.n1345 585
R1616 gnd.n4924 gnd.n1345 585
R1617 gnd.n2897 gnd.n2896 585
R1618 gnd.n2898 gnd.n2897 585
R1619 gnd.n2431 gnd.n1335 585
R1620 gnd.n4930 gnd.n1335 585
R1621 gnd.n2863 gnd.n2862 585
R1622 gnd.n2864 gnd.n2863 585
R1623 gnd.n2440 gnd.n1325 585
R1624 gnd.n4936 gnd.n1325 585
R1625 gnd.n2858 gnd.n2857 585
R1626 gnd.n2857 gnd.n2856 585
R1627 gnd.n2442 gnd.n1315 585
R1628 gnd.n4942 gnd.n1315 585
R1629 gnd.n2848 gnd.n2847 585
R1630 gnd.n2849 gnd.n2848 585
R1631 gnd.n2445 gnd.n1305 585
R1632 gnd.n4948 gnd.n1305 585
R1633 gnd.n2843 gnd.n2842 585
R1634 gnd.n2842 gnd.n2841 585
R1635 gnd.n2447 gnd.n1295 585
R1636 gnd.n4954 gnd.n1295 585
R1637 gnd.n2790 gnd.n2789 585
R1638 gnd.n2789 gnd.n2788 585
R1639 gnd.n2469 gnd.n1285 585
R1640 gnd.n4960 gnd.n1285 585
R1641 gnd.n2794 gnd.n2468 585
R1642 gnd.n2779 gnd.n2468 585
R1643 gnd.n2795 gnd.n1276 585
R1644 gnd.n4966 gnd.n1276 585
R1645 gnd.n2796 gnd.n2467 585
R1646 gnd.n2773 gnd.n2467 585
R1647 gnd.n2464 gnd.n1264 585
R1648 gnd.n4972 gnd.n1264 585
R1649 gnd.n2801 gnd.n2800 585
R1650 gnd.n2802 gnd.n2801 585
R1651 gnd.n2463 gnd.n2462 585
R1652 gnd.n2766 gnd.n2462 585
R1653 gnd.n2760 gnd.n2759 585
R1654 gnd.n2761 gnd.n2760 585
R1655 gnd.n2479 gnd.n2478 585
R1656 gnd.n2741 gnd.n2478 585
R1657 gnd.n2754 gnd.n2753 585
R1658 gnd.n2753 gnd.n2752 585
R1659 gnd.n2482 gnd.n2481 585
R1660 gnd.n2747 gnd.n2482 585
R1661 gnd.n2714 gnd.n2713 585
R1662 gnd.n2715 gnd.n2714 585
R1663 gnd.n2515 gnd.n2505 585
R1664 gnd.n2723 gnd.n2505 585
R1665 gnd.n2709 gnd.n2708 585
R1666 gnd.n2708 gnd.n2503 585
R1667 gnd.n2707 gnd.n1247 585
R1668 gnd.n4980 gnd.n1247 585
R1669 gnd.n2706 gnd.n2705 585
R1670 gnd.n2705 gnd.n2704 585
R1671 gnd.n2517 gnd.n1237 585
R1672 gnd.n4986 gnd.n1237 585
R1673 gnd.n2696 gnd.n2695 585
R1674 gnd.n2697 gnd.n2696 585
R1675 gnd.n2521 gnd.n1226 585
R1676 gnd.n4992 gnd.n1226 585
R1677 gnd.n2690 gnd.n2689 585
R1678 gnd.n2689 gnd.n2688 585
R1679 gnd.n2523 gnd.n1216 585
R1680 gnd.n4998 gnd.n1216 585
R1681 gnd.n2642 gnd.n2641 585
R1682 gnd.n2682 gnd.n2642 585
R1683 gnd.n2526 gnd.n1206 585
R1684 gnd.n5004 gnd.n1206 585
R1685 gnd.n2637 gnd.n2636 585
R1686 gnd.n2636 gnd.n2635 585
R1687 gnd.n2528 gnd.n1196 585
R1688 gnd.n5010 gnd.n1196 585
R1689 gnd.n2628 gnd.n2627 585
R1690 gnd.n2629 gnd.n2628 585
R1691 gnd.n2543 gnd.n1186 585
R1692 gnd.n5016 gnd.n1186 585
R1693 gnd.n2623 gnd.n2622 585
R1694 gnd.n2622 gnd.n1177 585
R1695 gnd.n2621 gnd.n1176 585
R1696 gnd.n5022 gnd.n1176 585
R1697 gnd.n2620 gnd.n2619 585
R1698 gnd.n2619 gnd.n1167 585
R1699 gnd.n2545 gnd.n1166 585
R1700 gnd.n5028 gnd.n1166 585
R1701 gnd.n2615 gnd.n2614 585
R1702 gnd.n2614 gnd.n1155 585
R1703 gnd.n2613 gnd.n1154 585
R1704 gnd.n5034 gnd.n1154 585
R1705 gnd.n2612 gnd.n2611 585
R1706 gnd.n2611 gnd.n1152 585
R1707 gnd.n2547 gnd.n1142 585
R1708 gnd.n5040 gnd.n1142 585
R1709 gnd.n2607 gnd.n2606 585
R1710 gnd.n2606 gnd.n1068 585
R1711 gnd.n6548 gnd.n6547 585
R1712 gnd.n6547 gnd.n6546 585
R1713 gnd.n6549 gnd.n1021 585
R1714 gnd.n6456 gnd.n1021 585
R1715 gnd.n6551 gnd.n6550 585
R1716 gnd.n6552 gnd.n6551 585
R1717 gnd.n1022 gnd.n1020 585
R1718 gnd.n1020 gnd.n1016 585
R1719 gnd.n1001 gnd.n1000 585
R1720 gnd.n1005 gnd.n1001 585
R1721 gnd.n6562 gnd.n6561 585
R1722 gnd.n6561 gnd.n6560 585
R1723 gnd.n6563 gnd.n995 585
R1724 gnd.n6445 gnd.n995 585
R1725 gnd.n6565 gnd.n6564 585
R1726 gnd.n6566 gnd.n6565 585
R1727 gnd.n996 gnd.n994 585
R1728 gnd.n994 gnd.n990 585
R1729 gnd.n978 gnd.n977 585
R1730 gnd.n6438 gnd.n978 585
R1731 gnd.n6576 gnd.n6575 585
R1732 gnd.n6575 gnd.n6574 585
R1733 gnd.n6577 gnd.n972 585
R1734 gnd.n6101 gnd.n972 585
R1735 gnd.n6579 gnd.n6578 585
R1736 gnd.n6580 gnd.n6579 585
R1737 gnd.n973 gnd.n971 585
R1738 gnd.n5263 gnd.n971 585
R1739 gnd.n6139 gnd.n6138 585
R1740 gnd.n6138 gnd.n6137 585
R1741 gnd.n5261 gnd.n5260 585
R1742 gnd.n6121 gnd.n5261 585
R1743 gnd.n6113 gnd.n6112 585
R1744 gnd.n6112 gnd.n6111 585
R1745 gnd.n5275 gnd.n5274 585
R1746 gnd.n5283 gnd.n5275 585
R1747 gnd.n6087 gnd.n6086 585
R1748 gnd.n6088 gnd.n6087 585
R1749 gnd.n5286 gnd.n5285 585
R1750 gnd.n5293 gnd.n5285 585
R1751 gnd.n6061 gnd.n5305 585
R1752 gnd.n5305 gnd.n5292 585
R1753 gnd.n6063 gnd.n6062 585
R1754 gnd.n6064 gnd.n6063 585
R1755 gnd.n5306 gnd.n5304 585
R1756 gnd.n5304 gnd.n5300 585
R1757 gnd.n6050 gnd.n6049 585
R1758 gnd.n6049 gnd.n6048 585
R1759 gnd.n5311 gnd.n5310 585
R1760 gnd.n5321 gnd.n5311 585
R1761 gnd.n6039 gnd.n6038 585
R1762 gnd.n6038 gnd.n6037 585
R1763 gnd.n5318 gnd.n5317 585
R1764 gnd.n6025 gnd.n5318 585
R1765 gnd.n5999 gnd.n5403 585
R1766 gnd.n5403 gnd.n5328 585
R1767 gnd.n6001 gnd.n6000 585
R1768 gnd.n6002 gnd.n6001 585
R1769 gnd.n5404 gnd.n5402 585
R1770 gnd.n5412 gnd.n5402 585
R1771 gnd.n5977 gnd.n5424 585
R1772 gnd.n5424 gnd.n5411 585
R1773 gnd.n5979 gnd.n5978 585
R1774 gnd.n5980 gnd.n5979 585
R1775 gnd.n5425 gnd.n5423 585
R1776 gnd.n5423 gnd.n5419 585
R1777 gnd.n5965 gnd.n5964 585
R1778 gnd.n5964 gnd.n5963 585
R1779 gnd.n5430 gnd.n5429 585
R1780 gnd.n5439 gnd.n5430 585
R1781 gnd.n5954 gnd.n5953 585
R1782 gnd.n5953 gnd.n5952 585
R1783 gnd.n5437 gnd.n5436 585
R1784 gnd.n5940 gnd.n5437 585
R1785 gnd.n5912 gnd.n5911 585
R1786 gnd.n5911 gnd.n5446 585
R1787 gnd.n5913 gnd.n5457 585
R1788 gnd.n5904 gnd.n5457 585
R1789 gnd.n5915 gnd.n5914 585
R1790 gnd.n5916 gnd.n5915 585
R1791 gnd.n5458 gnd.n5456 585
R1792 gnd.n5472 gnd.n5456 585
R1793 gnd.n5896 gnd.n5895 585
R1794 gnd.n5895 gnd.n5894 585
R1795 gnd.n5469 gnd.n5468 585
R1796 gnd.n5879 gnd.n5469 585
R1797 gnd.n5866 gnd.n5489 585
R1798 gnd.n5489 gnd.n5479 585
R1799 gnd.n5868 gnd.n5867 585
R1800 gnd.n5869 gnd.n5868 585
R1801 gnd.n5490 gnd.n5488 585
R1802 gnd.n5498 gnd.n5488 585
R1803 gnd.n5842 gnd.n5510 585
R1804 gnd.n5510 gnd.n5497 585
R1805 gnd.n5844 gnd.n5843 585
R1806 gnd.n5845 gnd.n5844 585
R1807 gnd.n5511 gnd.n5509 585
R1808 gnd.n5509 gnd.n5505 585
R1809 gnd.n5830 gnd.n5829 585
R1810 gnd.n5829 gnd.n5828 585
R1811 gnd.n5516 gnd.n5515 585
R1812 gnd.n5520 gnd.n5516 585
R1813 gnd.n5814 gnd.n5813 585
R1814 gnd.n5815 gnd.n5814 585
R1815 gnd.n5531 gnd.n5530 585
R1816 gnd.n5530 gnd.n5526 585
R1817 gnd.n5804 gnd.n5803 585
R1818 gnd.n5805 gnd.n5804 585
R1819 gnd.n5540 gnd.n5539 585
R1820 gnd.n5539 gnd.n5537 585
R1821 gnd.n5798 gnd.n5797 585
R1822 gnd.n5797 gnd.n5796 585
R1823 gnd.n5544 gnd.n5543 585
R1824 gnd.n5552 gnd.n5544 585
R1825 gnd.n5705 gnd.n5704 585
R1826 gnd.n5706 gnd.n5705 585
R1827 gnd.n5554 gnd.n5553 585
R1828 gnd.n5553 gnd.n5551 585
R1829 gnd.n5700 gnd.n5699 585
R1830 gnd.n5699 gnd.n5698 585
R1831 gnd.n5557 gnd.n5556 585
R1832 gnd.n5558 gnd.n5557 585
R1833 gnd.n5689 gnd.n5688 585
R1834 gnd.n5690 gnd.n5689 585
R1835 gnd.n5566 gnd.n5565 585
R1836 gnd.n5565 gnd.n5564 585
R1837 gnd.n5684 gnd.n5683 585
R1838 gnd.n5683 gnd.n5682 585
R1839 gnd.n5569 gnd.n5568 585
R1840 gnd.n5570 gnd.n5569 585
R1841 gnd.n5673 gnd.n5672 585
R1842 gnd.n5674 gnd.n5673 585
R1843 gnd.n5669 gnd.n5576 585
R1844 gnd.n5668 gnd.n5667 585
R1845 gnd.n5665 gnd.n5578 585
R1846 gnd.n5665 gnd.n5575 585
R1847 gnd.n5664 gnd.n5663 585
R1848 gnd.n5662 gnd.n5661 585
R1849 gnd.n5660 gnd.n5583 585
R1850 gnd.n5658 gnd.n5657 585
R1851 gnd.n5656 gnd.n5584 585
R1852 gnd.n5655 gnd.n5654 585
R1853 gnd.n5652 gnd.n5589 585
R1854 gnd.n5650 gnd.n5649 585
R1855 gnd.n5648 gnd.n5590 585
R1856 gnd.n5647 gnd.n5646 585
R1857 gnd.n5644 gnd.n5595 585
R1858 gnd.n5642 gnd.n5641 585
R1859 gnd.n5640 gnd.n5596 585
R1860 gnd.n5639 gnd.n5638 585
R1861 gnd.n5636 gnd.n5601 585
R1862 gnd.n5634 gnd.n5633 585
R1863 gnd.n5632 gnd.n5602 585
R1864 gnd.n5631 gnd.n5630 585
R1865 gnd.n5628 gnd.n5607 585
R1866 gnd.n5626 gnd.n5625 585
R1867 gnd.n5623 gnd.n5608 585
R1868 gnd.n5622 gnd.n5621 585
R1869 gnd.n5619 gnd.n5617 585
R1870 gnd.n5615 gnd.n5574 585
R1871 gnd.n6464 gnd.n6463 585
R1872 gnd.n6465 gnd.n5244 585
R1873 gnd.n6467 gnd.n6466 585
R1874 gnd.n6469 gnd.n5243 585
R1875 gnd.n6471 gnd.n6470 585
R1876 gnd.n6472 gnd.n5234 585
R1877 gnd.n6474 gnd.n6473 585
R1878 gnd.n6476 gnd.n5232 585
R1879 gnd.n6478 gnd.n6477 585
R1880 gnd.n6479 gnd.n5227 585
R1881 gnd.n6481 gnd.n6480 585
R1882 gnd.n6483 gnd.n5225 585
R1883 gnd.n6485 gnd.n6484 585
R1884 gnd.n6486 gnd.n5220 585
R1885 gnd.n6488 gnd.n6487 585
R1886 gnd.n6490 gnd.n5218 585
R1887 gnd.n6492 gnd.n6491 585
R1888 gnd.n6493 gnd.n5213 585
R1889 gnd.n6495 gnd.n6494 585
R1890 gnd.n6497 gnd.n5211 585
R1891 gnd.n6499 gnd.n6498 585
R1892 gnd.n6500 gnd.n5206 585
R1893 gnd.n6502 gnd.n6501 585
R1894 gnd.n6504 gnd.n5204 585
R1895 gnd.n6506 gnd.n6505 585
R1896 gnd.n6507 gnd.n5202 585
R1897 gnd.n6508 gnd.n1026 585
R1898 gnd.n5165 gnd.n1026 585
R1899 gnd.n6459 gnd.n1028 585
R1900 gnd.n6546 gnd.n1028 585
R1901 gnd.n6458 gnd.n6457 585
R1902 gnd.n6457 gnd.n6456 585
R1903 gnd.n6455 gnd.n1018 585
R1904 gnd.n6552 gnd.n1018 585
R1905 gnd.n6449 gnd.n5249 585
R1906 gnd.n6449 gnd.n1016 585
R1907 gnd.n6451 gnd.n6450 585
R1908 gnd.n6450 gnd.n1005 585
R1909 gnd.n6448 gnd.n1003 585
R1910 gnd.n6560 gnd.n1003 585
R1911 gnd.n6447 gnd.n6446 585
R1912 gnd.n6446 gnd.n6445 585
R1913 gnd.n5251 gnd.n992 585
R1914 gnd.n6566 gnd.n992 585
R1915 gnd.n6441 gnd.n6440 585
R1916 gnd.n6440 gnd.n990 585
R1917 gnd.n6439 gnd.n5253 585
R1918 gnd.n6439 gnd.n6438 585
R1919 gnd.n6100 gnd.n980 585
R1920 gnd.n6574 gnd.n980 585
R1921 gnd.n6103 gnd.n6102 585
R1922 gnd.n6102 gnd.n6101 585
R1923 gnd.n6104 gnd.n969 585
R1924 gnd.n6580 gnd.n969 585
R1925 gnd.n6106 gnd.n6105 585
R1926 gnd.n6105 gnd.n5263 585
R1927 gnd.n6107 gnd.n5262 585
R1928 gnd.n6137 gnd.n5262 585
R1929 gnd.n6108 gnd.n5271 585
R1930 gnd.n6121 gnd.n5271 585
R1931 gnd.n6110 gnd.n6109 585
R1932 gnd.n6111 gnd.n6110 585
R1933 gnd.n5278 gnd.n5277 585
R1934 gnd.n5283 gnd.n5277 585
R1935 gnd.n6090 gnd.n6089 585
R1936 gnd.n6089 gnd.n6088 585
R1937 gnd.n5281 gnd.n5280 585
R1938 gnd.n5293 gnd.n5281 585
R1939 gnd.n6015 gnd.n6014 585
R1940 gnd.n6014 gnd.n5292 585
R1941 gnd.n6016 gnd.n5302 585
R1942 gnd.n6064 gnd.n5302 585
R1943 gnd.n6018 gnd.n6017 585
R1944 gnd.n6017 gnd.n5300 585
R1945 gnd.n6019 gnd.n5313 585
R1946 gnd.n6048 gnd.n5313 585
R1947 gnd.n6021 gnd.n6020 585
R1948 gnd.n6020 gnd.n5321 585
R1949 gnd.n6022 gnd.n5320 585
R1950 gnd.n6037 gnd.n5320 585
R1951 gnd.n6024 gnd.n6023 585
R1952 gnd.n6025 gnd.n6024 585
R1953 gnd.n5332 gnd.n5331 585
R1954 gnd.n5331 gnd.n5328 585
R1955 gnd.n6004 gnd.n6003 585
R1956 gnd.n6003 gnd.n6002 585
R1957 gnd.n5399 gnd.n5398 585
R1958 gnd.n5412 gnd.n5399 585
R1959 gnd.n5925 gnd.n5924 585
R1960 gnd.n5924 gnd.n5411 585
R1961 gnd.n5926 gnd.n5421 585
R1962 gnd.n5980 gnd.n5421 585
R1963 gnd.n5929 gnd.n5928 585
R1964 gnd.n5928 gnd.n5419 585
R1965 gnd.n5930 gnd.n5432 585
R1966 gnd.n5963 gnd.n5432 585
R1967 gnd.n5933 gnd.n5932 585
R1968 gnd.n5932 gnd.n5439 585
R1969 gnd.n5934 gnd.n5438 585
R1970 gnd.n5952 gnd.n5438 585
R1971 gnd.n5937 gnd.n5936 585
R1972 gnd.n5940 gnd.n5937 585
R1973 gnd.n5922 gnd.n5448 585
R1974 gnd.n5448 gnd.n5446 585
R1975 gnd.n5453 gnd.n5449 585
R1976 gnd.n5904 gnd.n5453 585
R1977 gnd.n5918 gnd.n5917 585
R1978 gnd.n5917 gnd.n5916 585
R1979 gnd.n5452 gnd.n5451 585
R1980 gnd.n5472 gnd.n5452 585
R1981 gnd.n5876 gnd.n5471 585
R1982 gnd.n5894 gnd.n5471 585
R1983 gnd.n5878 gnd.n5877 585
R1984 gnd.n5879 gnd.n5878 585
R1985 gnd.n5482 gnd.n5481 585
R1986 gnd.n5481 gnd.n5479 585
R1987 gnd.n5871 gnd.n5870 585
R1988 gnd.n5870 gnd.n5869 585
R1989 gnd.n5485 gnd.n5484 585
R1990 gnd.n5498 gnd.n5485 585
R1991 gnd.n5722 gnd.n5721 585
R1992 gnd.n5721 gnd.n5497 585
R1993 gnd.n5723 gnd.n5507 585
R1994 gnd.n5845 gnd.n5507 585
R1995 gnd.n5725 gnd.n5724 585
R1996 gnd.n5724 gnd.n5505 585
R1997 gnd.n5726 gnd.n5517 585
R1998 gnd.n5828 gnd.n5517 585
R1999 gnd.n5728 gnd.n5727 585
R2000 gnd.n5727 gnd.n5520 585
R2001 gnd.n5729 gnd.n5528 585
R2002 gnd.n5815 gnd.n5528 585
R2003 gnd.n5731 gnd.n5730 585
R2004 gnd.n5730 gnd.n5526 585
R2005 gnd.n5732 gnd.n5538 585
R2006 gnd.n5805 gnd.n5538 585
R2007 gnd.n5733 gnd.n5546 585
R2008 gnd.n5546 gnd.n5537 585
R2009 gnd.n5735 gnd.n5734 585
R2010 gnd.n5796 gnd.n5735 585
R2011 gnd.n5547 gnd.n5545 585
R2012 gnd.n5552 gnd.n5545 585
R2013 gnd.n5708 gnd.n5707 585
R2014 gnd.n5707 gnd.n5706 585
R2015 gnd.n5550 gnd.n5549 585
R2016 gnd.n5551 gnd.n5550 585
R2017 gnd.n5697 gnd.n5696 585
R2018 gnd.n5698 gnd.n5697 585
R2019 gnd.n5560 gnd.n5559 585
R2020 gnd.n5559 gnd.n5558 585
R2021 gnd.n5692 gnd.n5691 585
R2022 gnd.n5691 gnd.n5690 585
R2023 gnd.n5563 gnd.n5562 585
R2024 gnd.n5564 gnd.n5563 585
R2025 gnd.n5681 gnd.n5680 585
R2026 gnd.n5682 gnd.n5681 585
R2027 gnd.n5572 gnd.n5571 585
R2028 gnd.n5571 gnd.n5570 585
R2029 gnd.n5676 gnd.n5675 585
R2030 gnd.n5675 gnd.n5674 585
R2031 gnd.n7677 gnd.n7676 585
R2032 gnd.n7676 gnd.n7675 585
R2033 gnd.n7678 gnd.n204 585
R2034 gnd.n209 gnd.n204 585
R2035 gnd.n7680 gnd.n7679 585
R2036 gnd.n7681 gnd.n7680 585
R2037 gnd.n191 gnd.n190 585
R2038 gnd.n194 gnd.n191 585
R2039 gnd.n7689 gnd.n7688 585
R2040 gnd.n7688 gnd.n7687 585
R2041 gnd.n7690 gnd.n186 585
R2042 gnd.n186 gnd.n185 585
R2043 gnd.n7692 gnd.n7691 585
R2044 gnd.n7693 gnd.n7692 585
R2045 gnd.n171 gnd.n170 585
R2046 gnd.n175 gnd.n171 585
R2047 gnd.n7701 gnd.n7700 585
R2048 gnd.n7700 gnd.n7699 585
R2049 gnd.n7702 gnd.n166 585
R2050 gnd.n7510 gnd.n166 585
R2051 gnd.n7704 gnd.n7703 585
R2052 gnd.n7705 gnd.n7704 585
R2053 gnd.n152 gnd.n151 585
R2054 gnd.n7489 gnd.n152 585
R2055 gnd.n7713 gnd.n7712 585
R2056 gnd.n7712 gnd.n7711 585
R2057 gnd.n7714 gnd.n147 585
R2058 gnd.n7480 gnd.n147 585
R2059 gnd.n7716 gnd.n7715 585
R2060 gnd.n7717 gnd.n7716 585
R2061 gnd.n131 gnd.n130 585
R2062 gnd.n7474 gnd.n131 585
R2063 gnd.n7725 gnd.n7724 585
R2064 gnd.n7724 gnd.n7723 585
R2065 gnd.n7726 gnd.n126 585
R2066 gnd.n7466 gnd.n126 585
R2067 gnd.n7728 gnd.n7727 585
R2068 gnd.n7729 gnd.n7728 585
R2069 gnd.n113 gnd.n112 585
R2070 gnd.n7460 gnd.n113 585
R2071 gnd.n7737 gnd.n7736 585
R2072 gnd.n7736 gnd.n7735 585
R2073 gnd.n7738 gnd.n107 585
R2074 gnd.n7452 gnd.n107 585
R2075 gnd.n7740 gnd.n7739 585
R2076 gnd.n7741 gnd.n7740 585
R2077 gnd.n108 gnd.n106 585
R2078 gnd.n7446 gnd.n106 585
R2079 gnd.n4532 gnd.n4531 585
R2080 gnd.n4531 gnd.n381 585
R2081 gnd.n4533 gnd.n88 585
R2082 gnd.n7749 gnd.n88 585
R2083 gnd.n4535 gnd.n4534 585
R2084 gnd.n4536 gnd.n4535 585
R2085 gnd.n4526 gnd.n4525 585
R2086 gnd.n4525 gnd.n1751 585
R2087 gnd.n1739 gnd.n1738 585
R2088 gnd.n4572 gnd.n1739 585
R2089 gnd.n4577 gnd.n4576 585
R2090 gnd.n4576 gnd.n4575 585
R2091 gnd.n4578 gnd.n1734 585
R2092 gnd.n4557 gnd.n1734 585
R2093 gnd.n4580 gnd.n4579 585
R2094 gnd.n4581 gnd.n4580 585
R2095 gnd.n1722 gnd.n1721 585
R2096 gnd.n4546 gnd.n1722 585
R2097 gnd.n4589 gnd.n4588 585
R2098 gnd.n4588 gnd.n4587 585
R2099 gnd.n4590 gnd.n1717 585
R2100 gnd.n4516 gnd.n1717 585
R2101 gnd.n4592 gnd.n4591 585
R2102 gnd.n4593 gnd.n4592 585
R2103 gnd.n1701 gnd.n1700 585
R2104 gnd.n4475 gnd.n1701 585
R2105 gnd.n4601 gnd.n4600 585
R2106 gnd.n4600 gnd.n4599 585
R2107 gnd.n4602 gnd.n1696 585
R2108 gnd.n4468 gnd.n1696 585
R2109 gnd.n4604 gnd.n4603 585
R2110 gnd.n4605 gnd.n4604 585
R2111 gnd.n1682 gnd.n1681 585
R2112 gnd.n4463 gnd.n1682 585
R2113 gnd.n4613 gnd.n4612 585
R2114 gnd.n4612 gnd.n4611 585
R2115 gnd.n4614 gnd.n1677 585
R2116 gnd.n4492 gnd.n1677 585
R2117 gnd.n4616 gnd.n4615 585
R2118 gnd.n4617 gnd.n4616 585
R2119 gnd.n1661 gnd.n1660 585
R2120 gnd.n4456 gnd.n1661 585
R2121 gnd.n4625 gnd.n4624 585
R2122 gnd.n4624 gnd.n4623 585
R2123 gnd.n4626 gnd.n1656 585
R2124 gnd.n4448 gnd.n1656 585
R2125 gnd.n4628 gnd.n4627 585
R2126 gnd.n4629 gnd.n4628 585
R2127 gnd.n1641 gnd.n1640 585
R2128 gnd.n4442 gnd.n1641 585
R2129 gnd.n4637 gnd.n4636 585
R2130 gnd.n4636 gnd.n4635 585
R2131 gnd.n4638 gnd.n1635 585
R2132 gnd.n4434 gnd.n1635 585
R2133 gnd.n4640 gnd.n4639 585
R2134 gnd.n4641 gnd.n4640 585
R2135 gnd.n1636 gnd.n1634 585
R2136 gnd.n3886 gnd.n1634 585
R2137 gnd.n4427 gnd.n1622 585
R2138 gnd.n4647 gnd.n1622 585
R2139 gnd.n3972 gnd.n3971 585
R2140 gnd.n3936 gnd.n3935 585
R2141 gnd.n3986 gnd.n3985 585
R2142 gnd.n3988 gnd.n3934 585
R2143 gnd.n3991 gnd.n3990 585
R2144 gnd.n3927 gnd.n3926 585
R2145 gnd.n4005 gnd.n4004 585
R2146 gnd.n4007 gnd.n3925 585
R2147 gnd.n4010 gnd.n4009 585
R2148 gnd.n3918 gnd.n3917 585
R2149 gnd.n4024 gnd.n4023 585
R2150 gnd.n4026 gnd.n3916 585
R2151 gnd.n4029 gnd.n4028 585
R2152 gnd.n3909 gnd.n3908 585
R2153 gnd.n4044 gnd.n4043 585
R2154 gnd.n4046 gnd.n3907 585
R2155 gnd.n4049 gnd.n4048 585
R2156 gnd.n4050 gnd.n3904 585
R2157 gnd.n3903 gnd.n3902 585
R2158 gnd.n3903 gnd.n1610 585
R2159 gnd.n349 gnd.n348 585
R2160 gnd.n7531 gnd.n344 585
R2161 gnd.n7533 gnd.n7532 585
R2162 gnd.n7535 gnd.n342 585
R2163 gnd.n7537 gnd.n7536 585
R2164 gnd.n7538 gnd.n337 585
R2165 gnd.n7540 gnd.n7539 585
R2166 gnd.n7542 gnd.n335 585
R2167 gnd.n7544 gnd.n7543 585
R2168 gnd.n7545 gnd.n330 585
R2169 gnd.n7547 gnd.n7546 585
R2170 gnd.n7549 gnd.n328 585
R2171 gnd.n7551 gnd.n7550 585
R2172 gnd.n7552 gnd.n323 585
R2173 gnd.n7554 gnd.n7553 585
R2174 gnd.n7556 gnd.n321 585
R2175 gnd.n7558 gnd.n7557 585
R2176 gnd.n7559 gnd.n319 585
R2177 gnd.n7560 gnd.n208 585
R2178 gnd.n212 gnd.n208 585
R2179 gnd.n7527 gnd.n211 585
R2180 gnd.n7675 gnd.n211 585
R2181 gnd.n7526 gnd.n7525 585
R2182 gnd.n7525 gnd.n209 585
R2183 gnd.n7524 gnd.n203 585
R2184 gnd.n7681 gnd.n203 585
R2185 gnd.n354 gnd.n353 585
R2186 gnd.n353 gnd.n194 585
R2187 gnd.n7520 gnd.n193 585
R2188 gnd.n7687 gnd.n193 585
R2189 gnd.n7519 gnd.n7518 585
R2190 gnd.n7518 gnd.n185 585
R2191 gnd.n7517 gnd.n184 585
R2192 gnd.n7693 gnd.n184 585
R2193 gnd.n357 gnd.n356 585
R2194 gnd.n356 gnd.n175 585
R2195 gnd.n7513 gnd.n174 585
R2196 gnd.n7699 gnd.n174 585
R2197 gnd.n7512 gnd.n7511 585
R2198 gnd.n7511 gnd.n7510 585
R2199 gnd.n359 gnd.n165 585
R2200 gnd.n7705 gnd.n165 585
R2201 gnd.n7488 gnd.n7487 585
R2202 gnd.n7489 gnd.n7488 585
R2203 gnd.n363 gnd.n155 585
R2204 gnd.n7711 gnd.n155 585
R2205 gnd.n7482 gnd.n7481 585
R2206 gnd.n7481 gnd.n7480 585
R2207 gnd.n365 gnd.n145 585
R2208 gnd.n7717 gnd.n145 585
R2209 gnd.n7473 gnd.n7472 585
R2210 gnd.n7474 gnd.n7473 585
R2211 gnd.n368 gnd.n134 585
R2212 gnd.n7723 gnd.n134 585
R2213 gnd.n7468 gnd.n7467 585
R2214 gnd.n7467 gnd.n7466 585
R2215 gnd.n370 gnd.n125 585
R2216 gnd.n7729 gnd.n125 585
R2217 gnd.n7459 gnd.n7458 585
R2218 gnd.n7460 gnd.n7459 585
R2219 gnd.n375 gnd.n116 585
R2220 gnd.n7735 gnd.n116 585
R2221 gnd.n7454 gnd.n7453 585
R2222 gnd.n7453 gnd.n7452 585
R2223 gnd.n377 gnd.n104 585
R2224 gnd.n7741 gnd.n104 585
R2225 gnd.n7445 gnd.n7444 585
R2226 gnd.n7446 gnd.n7445 585
R2227 gnd.n84 gnd.n83 585
R2228 gnd.n381 gnd.n84 585
R2229 gnd.n7751 gnd.n7750 585
R2230 gnd.n7750 gnd.n7749 585
R2231 gnd.n7752 gnd.n82 585
R2232 gnd.n4536 gnd.n82 585
R2233 gnd.n1750 gnd.n81 585
R2234 gnd.n1751 gnd.n1750 585
R2235 gnd.n4551 gnd.n1749 585
R2236 gnd.n4572 gnd.n1749 585
R2237 gnd.n1758 gnd.n1742 585
R2238 gnd.n4575 gnd.n1742 585
R2239 gnd.n4556 gnd.n4555 585
R2240 gnd.n4557 gnd.n4556 585
R2241 gnd.n1757 gnd.n1733 585
R2242 gnd.n4581 gnd.n1733 585
R2243 gnd.n4548 gnd.n4547 585
R2244 gnd.n4547 gnd.n4546 585
R2245 gnd.n1760 gnd.n1724 585
R2246 gnd.n4587 gnd.n1724 585
R2247 gnd.n4478 gnd.n1762 585
R2248 gnd.n4516 gnd.n1762 585
R2249 gnd.n4479 gnd.n1715 585
R2250 gnd.n4593 gnd.n1715 585
R2251 gnd.n4480 gnd.n4476 585
R2252 gnd.n4476 gnd.n4475 585
R2253 gnd.n1781 gnd.n1704 585
R2254 gnd.n4599 gnd.n1704 585
R2255 gnd.n4484 gnd.n1780 585
R2256 gnd.n4468 gnd.n1780 585
R2257 gnd.n4485 gnd.n1695 585
R2258 gnd.n4605 gnd.n1695 585
R2259 gnd.n4486 gnd.n1779 585
R2260 gnd.n4463 gnd.n1779 585
R2261 gnd.n1776 gnd.n1684 585
R2262 gnd.n4611 gnd.n1684 585
R2263 gnd.n4491 gnd.n4490 585
R2264 gnd.n4492 gnd.n4491 585
R2265 gnd.n1775 gnd.n1675 585
R2266 gnd.n4617 gnd.n1675 585
R2267 gnd.n4455 gnd.n4454 585
R2268 gnd.n4456 gnd.n4455 585
R2269 gnd.n1785 gnd.n1664 585
R2270 gnd.n4623 gnd.n1664 585
R2271 gnd.n4450 gnd.n4449 585
R2272 gnd.n4449 gnd.n4448 585
R2273 gnd.n1787 gnd.n1655 585
R2274 gnd.n4629 gnd.n1655 585
R2275 gnd.n4441 gnd.n4440 585
R2276 gnd.n4442 gnd.n4441 585
R2277 gnd.n1822 gnd.n1644 585
R2278 gnd.n4635 gnd.n1644 585
R2279 gnd.n4436 gnd.n4435 585
R2280 gnd.n4435 gnd.n4434 585
R2281 gnd.n1824 gnd.n1632 585
R2282 gnd.n4641 gnd.n1632 585
R2283 gnd.n3888 gnd.n3887 585
R2284 gnd.n3887 gnd.n3886 585
R2285 gnd.n3889 gnd.n1620 585
R2286 gnd.n4647 gnd.n1620 585
R2287 gnd.n6544 gnd.n6543 585
R2288 gnd.n6545 gnd.n6544 585
R2289 gnd.n5168 gnd.n5166 585
R2290 gnd.n5166 gnd.n1027 585
R2291 gnd.n1015 gnd.n1014 585
R2292 gnd.n1019 gnd.n1015 585
R2293 gnd.n6555 gnd.n6554 585
R2294 gnd.n6554 gnd.n6553 585
R2295 gnd.n6556 gnd.n1007 585
R2296 gnd.n6426 gnd.n1007 585
R2297 gnd.n6558 gnd.n6557 585
R2298 gnd.n6559 gnd.n6558 585
R2299 gnd.n1008 gnd.n1006 585
R2300 gnd.n1006 gnd.n1002 585
R2301 gnd.n989 gnd.n988 585
R2302 gnd.n993 gnd.n989 585
R2303 gnd.n6569 gnd.n6568 585
R2304 gnd.n6568 gnd.n6567 585
R2305 gnd.n6570 gnd.n983 585
R2306 gnd.n6437 gnd.n983 585
R2307 gnd.n6572 gnd.n6571 585
R2308 gnd.n6573 gnd.n6572 585
R2309 gnd.n984 gnd.n982 585
R2310 gnd.n982 gnd.n979 585
R2311 gnd.n6132 gnd.n6131 585
R2312 gnd.n6131 gnd.n970 585
R2313 gnd.n6133 gnd.n5265 585
R2314 gnd.n5265 gnd.n968 585
R2315 gnd.n6135 gnd.n6134 585
R2316 gnd.n6136 gnd.n6135 585
R2317 gnd.n5266 gnd.n5264 585
R2318 gnd.n6120 gnd.n5264 585
R2319 gnd.n6124 gnd.n6123 585
R2320 gnd.n6123 gnd.n6122 585
R2321 gnd.n5269 gnd.n5268 585
R2322 gnd.n5276 gnd.n5269 585
R2323 gnd.n6074 gnd.n6073 585
R2324 gnd.n6073 gnd.n5284 585
R2325 gnd.n6075 gnd.n5295 585
R2326 gnd.n5295 gnd.n5282 585
R2327 gnd.n6077 gnd.n6076 585
R2328 gnd.n6078 gnd.n6077 585
R2329 gnd.n5296 gnd.n5294 585
R2330 gnd.n5303 gnd.n5294 585
R2331 gnd.n6067 gnd.n6066 585
R2332 gnd.n6066 gnd.n6065 585
R2333 gnd.n5299 gnd.n5298 585
R2334 gnd.n6047 gnd.n5299 585
R2335 gnd.n6033 gnd.n5323 585
R2336 gnd.n5323 gnd.n5312 585
R2337 gnd.n6035 gnd.n6034 585
R2338 gnd.n6036 gnd.n6035 585
R2339 gnd.n5324 gnd.n5322 585
R2340 gnd.n5322 gnd.n5319 585
R2341 gnd.n6028 gnd.n6027 585
R2342 gnd.n6027 gnd.n6026 585
R2343 gnd.n5327 gnd.n5326 585
R2344 gnd.n5401 gnd.n5327 585
R2345 gnd.n5988 gnd.n5414 585
R2346 gnd.n5414 gnd.n5400 585
R2347 gnd.n5990 gnd.n5989 585
R2348 gnd.n5991 gnd.n5990 585
R2349 gnd.n5415 gnd.n5413 585
R2350 gnd.n5422 gnd.n5413 585
R2351 gnd.n5983 gnd.n5982 585
R2352 gnd.n5982 gnd.n5981 585
R2353 gnd.n5418 gnd.n5417 585
R2354 gnd.n5962 gnd.n5418 585
R2355 gnd.n5948 gnd.n5441 585
R2356 gnd.n5441 gnd.n5431 585
R2357 gnd.n5950 gnd.n5949 585
R2358 gnd.n5951 gnd.n5950 585
R2359 gnd.n5442 gnd.n5440 585
R2360 gnd.n5939 gnd.n5440 585
R2361 gnd.n5943 gnd.n5942 585
R2362 gnd.n5942 gnd.n5941 585
R2363 gnd.n5445 gnd.n5444 585
R2364 gnd.n5905 gnd.n5445 585
R2365 gnd.n5889 gnd.n5888 585
R2366 gnd.n5888 gnd.n5455 585
R2367 gnd.n5890 gnd.n5474 585
R2368 gnd.n5474 gnd.n5454 585
R2369 gnd.n5892 gnd.n5891 585
R2370 gnd.n5893 gnd.n5892 585
R2371 gnd.n5475 gnd.n5473 585
R2372 gnd.n5473 gnd.n5470 585
R2373 gnd.n5882 gnd.n5881 585
R2374 gnd.n5881 gnd.n5880 585
R2375 gnd.n5478 gnd.n5477 585
R2376 gnd.n5487 gnd.n5478 585
R2377 gnd.n5853 gnd.n5500 585
R2378 gnd.n5500 gnd.n5486 585
R2379 gnd.n5855 gnd.n5854 585
R2380 gnd.n5856 gnd.n5855 585
R2381 gnd.n5501 gnd.n5499 585
R2382 gnd.n5508 gnd.n5499 585
R2383 gnd.n5848 gnd.n5847 585
R2384 gnd.n5847 gnd.n5846 585
R2385 gnd.n5504 gnd.n5503 585
R2386 gnd.n5827 gnd.n5504 585
R2387 gnd.n5823 gnd.n5822 585
R2388 gnd.n5824 gnd.n5823 585
R2389 gnd.n5522 gnd.n5521 585
R2390 gnd.n5529 gnd.n5521 585
R2391 gnd.n5818 gnd.n5817 585
R2392 gnd.n5817 gnd.n5816 585
R2393 gnd.n5525 gnd.n5524 585
R2394 gnd.n5806 gnd.n5525 585
R2395 gnd.n5793 gnd.n5792 585
R2396 gnd.n5791 gnd.n5744 585
R2397 gnd.n5790 gnd.n5743 585
R2398 gnd.n5795 gnd.n5743 585
R2399 gnd.n5789 gnd.n5788 585
R2400 gnd.n5787 gnd.n5786 585
R2401 gnd.n5785 gnd.n5784 585
R2402 gnd.n5783 gnd.n5782 585
R2403 gnd.n5781 gnd.n5780 585
R2404 gnd.n5779 gnd.n5778 585
R2405 gnd.n5777 gnd.n5776 585
R2406 gnd.n5775 gnd.n5774 585
R2407 gnd.n5773 gnd.n5772 585
R2408 gnd.n5771 gnd.n5770 585
R2409 gnd.n5769 gnd.n5768 585
R2410 gnd.n5767 gnd.n5766 585
R2411 gnd.n5765 gnd.n5764 585
R2412 gnd.n5760 gnd.n5536 585
R2413 gnd.n6513 gnd.n6512 585
R2414 gnd.n6515 gnd.n5197 585
R2415 gnd.n6517 gnd.n6516 585
R2416 gnd.n6518 gnd.n5190 585
R2417 gnd.n6520 gnd.n6519 585
R2418 gnd.n6522 gnd.n5188 585
R2419 gnd.n6524 gnd.n6523 585
R2420 gnd.n6525 gnd.n5183 585
R2421 gnd.n6527 gnd.n6526 585
R2422 gnd.n6529 gnd.n5181 585
R2423 gnd.n6531 gnd.n6530 585
R2424 gnd.n6532 gnd.n5176 585
R2425 gnd.n6534 gnd.n6533 585
R2426 gnd.n6536 gnd.n5174 585
R2427 gnd.n6538 gnd.n6537 585
R2428 gnd.n6539 gnd.n5172 585
R2429 gnd.n6540 gnd.n5167 585
R2430 gnd.n5167 gnd.n5165 585
R2431 gnd.n6420 gnd.n1029 585
R2432 gnd.n6545 gnd.n1029 585
R2433 gnd.n6422 gnd.n6421 585
R2434 gnd.n6422 gnd.n1027 585
R2435 gnd.n6424 gnd.n6423 585
R2436 gnd.n6423 gnd.n1019 585
R2437 gnd.n6425 gnd.n1017 585
R2438 gnd.n6553 gnd.n1017 585
R2439 gnd.n6428 gnd.n6427 585
R2440 gnd.n6427 gnd.n6426 585
R2441 gnd.n6429 gnd.n1004 585
R2442 gnd.n6559 gnd.n1004 585
R2443 gnd.n6431 gnd.n6430 585
R2444 gnd.n6431 gnd.n1002 585
R2445 gnd.n6433 gnd.n6432 585
R2446 gnd.n6432 gnd.n993 585
R2447 gnd.n6434 gnd.n991 585
R2448 gnd.n6567 gnd.n991 585
R2449 gnd.n6436 gnd.n6435 585
R2450 gnd.n6437 gnd.n6436 585
R2451 gnd.n6149 gnd.n981 585
R2452 gnd.n6573 gnd.n981 585
R2453 gnd.n6148 gnd.n6147 585
R2454 gnd.n6147 gnd.n979 585
R2455 gnd.n6146 gnd.n5255 585
R2456 gnd.n6146 gnd.n970 585
R2457 gnd.n6145 gnd.n6144 585
R2458 gnd.n6145 gnd.n968 585
R2459 gnd.n5258 gnd.n5257 585
R2460 gnd.n6136 gnd.n5257 585
R2461 gnd.n6119 gnd.n6118 585
R2462 gnd.n6120 gnd.n6119 585
R2463 gnd.n6117 gnd.n5270 585
R2464 gnd.n6122 gnd.n5270 585
R2465 gnd.n6081 gnd.n5272 585
R2466 gnd.n6081 gnd.n5276 585
R2467 gnd.n6083 gnd.n6082 585
R2468 gnd.n6082 gnd.n5284 585
R2469 gnd.n6080 gnd.n5289 585
R2470 gnd.n6080 gnd.n5282 585
R2471 gnd.n6079 gnd.n5291 585
R2472 gnd.n6079 gnd.n6078 585
R2473 gnd.n6056 gnd.n5290 585
R2474 gnd.n5303 gnd.n5290 585
R2475 gnd.n6055 gnd.n5301 585
R2476 gnd.n6065 gnd.n5301 585
R2477 gnd.n6046 gnd.n5308 585
R2478 gnd.n6047 gnd.n6046 585
R2479 gnd.n6045 gnd.n6044 585
R2480 gnd.n6045 gnd.n5312 585
R2481 gnd.n6043 gnd.n5314 585
R2482 gnd.n6036 gnd.n5314 585
R2483 gnd.n5329 gnd.n5315 585
R2484 gnd.n5329 gnd.n5319 585
R2485 gnd.n5996 gnd.n5330 585
R2486 gnd.n6026 gnd.n5330 585
R2487 gnd.n5995 gnd.n5994 585
R2488 gnd.n5994 gnd.n5401 585
R2489 gnd.n5993 gnd.n5408 585
R2490 gnd.n5993 gnd.n5400 585
R2491 gnd.n5992 gnd.n5410 585
R2492 gnd.n5992 gnd.n5991 585
R2493 gnd.n5971 gnd.n5409 585
R2494 gnd.n5422 gnd.n5409 585
R2495 gnd.n5970 gnd.n5420 585
R2496 gnd.n5981 gnd.n5420 585
R2497 gnd.n5961 gnd.n5427 585
R2498 gnd.n5962 gnd.n5961 585
R2499 gnd.n5960 gnd.n5959 585
R2500 gnd.n5960 gnd.n5431 585
R2501 gnd.n5958 gnd.n5433 585
R2502 gnd.n5951 gnd.n5433 585
R2503 gnd.n5938 gnd.n5434 585
R2504 gnd.n5939 gnd.n5938 585
R2505 gnd.n5908 gnd.n5447 585
R2506 gnd.n5941 gnd.n5447 585
R2507 gnd.n5907 gnd.n5906 585
R2508 gnd.n5906 gnd.n5905 585
R2509 gnd.n5903 gnd.n5464 585
R2510 gnd.n5903 gnd.n5455 585
R2511 gnd.n5902 gnd.n5901 585
R2512 gnd.n5902 gnd.n5454 585
R2513 gnd.n5466 gnd.n5465 585
R2514 gnd.n5893 gnd.n5465 585
R2515 gnd.n5862 gnd.n5861 585
R2516 gnd.n5861 gnd.n5470 585
R2517 gnd.n5863 gnd.n5480 585
R2518 gnd.n5880 gnd.n5480 585
R2519 gnd.n5860 gnd.n5859 585
R2520 gnd.n5859 gnd.n5487 585
R2521 gnd.n5858 gnd.n5494 585
R2522 gnd.n5858 gnd.n5486 585
R2523 gnd.n5857 gnd.n5496 585
R2524 gnd.n5857 gnd.n5856 585
R2525 gnd.n5836 gnd.n5495 585
R2526 gnd.n5508 gnd.n5495 585
R2527 gnd.n5835 gnd.n5506 585
R2528 gnd.n5846 gnd.n5506 585
R2529 gnd.n5826 gnd.n5513 585
R2530 gnd.n5827 gnd.n5826 585
R2531 gnd.n5825 gnd.n5519 585
R2532 gnd.n5825 gnd.n5824 585
R2533 gnd.n5810 gnd.n5518 585
R2534 gnd.n5529 gnd.n5518 585
R2535 gnd.n5809 gnd.n5527 585
R2536 gnd.n5816 gnd.n5527 585
R2537 gnd.n5808 gnd.n5807 585
R2538 gnd.n5807 gnd.n5806 585
R2539 gnd.n4178 gnd.n4177 585
R2540 gnd.n4179 gnd.n4178 585
R2541 gnd.n4092 gnd.n1903 585
R2542 gnd.n1910 gnd.n1903 585
R2543 gnd.n4091 gnd.n4090 585
R2544 gnd.n4090 gnd.n4089 585
R2545 gnd.n1906 gnd.n1905 585
R2546 gnd.n3860 gnd.n1906 585
R2547 gnd.n3849 gnd.n1953 585
R2548 gnd.n1953 gnd.n1947 585
R2549 gnd.n3851 gnd.n3850 585
R2550 gnd.n3852 gnd.n3851 585
R2551 gnd.n3848 gnd.n1952 585
R2552 gnd.n3842 gnd.n1952 585
R2553 gnd.n3847 gnd.n3846 585
R2554 gnd.n3846 gnd.n3845 585
R2555 gnd.n1955 gnd.n1954 585
R2556 gnd.n3829 gnd.n1955 585
R2557 gnd.n3804 gnd.n3803 585
R2558 gnd.n3803 gnd.n1966 585
R2559 gnd.n3805 gnd.n1975 585
R2560 gnd.n3818 gnd.n1975 585
R2561 gnd.n3806 gnd.n1985 585
R2562 gnd.n1985 gnd.n1974 585
R2563 gnd.n3808 gnd.n3807 585
R2564 gnd.n3809 gnd.n3808 585
R2565 gnd.n3802 gnd.n1984 585
R2566 gnd.n3797 gnd.n1984 585
R2567 gnd.n3801 gnd.n3800 585
R2568 gnd.n3800 gnd.n3799 585
R2569 gnd.n1987 gnd.n1986 585
R2570 gnd.n3784 gnd.n1987 585
R2571 gnd.n3773 gnd.n2002 585
R2572 gnd.n2002 gnd.n1996 585
R2573 gnd.n3775 gnd.n3774 585
R2574 gnd.n3776 gnd.n3775 585
R2575 gnd.n3772 gnd.n2001 585
R2576 gnd.n2008 gnd.n2001 585
R2577 gnd.n3771 gnd.n3770 585
R2578 gnd.n3770 gnd.n3769 585
R2579 gnd.n2004 gnd.n2003 585
R2580 gnd.n3650 gnd.n2004 585
R2581 gnd.n3757 gnd.n3756 585
R2582 gnd.n3758 gnd.n3757 585
R2583 gnd.n3755 gnd.n2020 585
R2584 gnd.n2020 gnd.n2016 585
R2585 gnd.n3754 gnd.n3753 585
R2586 gnd.n3753 gnd.n3752 585
R2587 gnd.n2022 gnd.n2021 585
R2588 gnd.n3660 gnd.n2022 585
R2589 gnd.n3726 gnd.n3725 585
R2590 gnd.n3727 gnd.n3726 585
R2591 gnd.n3724 gnd.n2033 585
R2592 gnd.n2033 gnd.n2030 585
R2593 gnd.n3723 gnd.n3722 585
R2594 gnd.n3722 gnd.n3721 585
R2595 gnd.n2035 gnd.n2034 585
R2596 gnd.n3667 gnd.n2035 585
R2597 gnd.n3707 gnd.n3706 585
R2598 gnd.n3708 gnd.n3707 585
R2599 gnd.n3705 gnd.n2046 585
R2600 gnd.n3700 gnd.n2046 585
R2601 gnd.n3704 gnd.n3703 585
R2602 gnd.n3703 gnd.n3702 585
R2603 gnd.n2048 gnd.n2047 585
R2604 gnd.n2060 gnd.n2048 585
R2605 gnd.n3636 gnd.n3635 585
R2606 gnd.n3636 gnd.n2059 585
R2607 gnd.n3640 gnd.n3639 585
R2608 gnd.n3639 gnd.n3638 585
R2609 gnd.n3641 gnd.n2066 585
R2610 gnd.n3680 gnd.n2066 585
R2611 gnd.n3642 gnd.n2075 585
R2612 gnd.n3566 gnd.n2075 585
R2613 gnd.n3644 gnd.n3643 585
R2614 gnd.n3645 gnd.n3644 585
R2615 gnd.n3634 gnd.n2074 585
R2616 gnd.n3629 gnd.n2074 585
R2617 gnd.n3633 gnd.n3632 585
R2618 gnd.n3632 gnd.n3631 585
R2619 gnd.n2077 gnd.n2076 585
R2620 gnd.n3618 gnd.n2077 585
R2621 gnd.n3608 gnd.n2095 585
R2622 gnd.n2095 gnd.n2086 585
R2623 gnd.n3610 gnd.n3609 585
R2624 gnd.n3611 gnd.n3610 585
R2625 gnd.n3607 gnd.n2094 585
R2626 gnd.n2099 gnd.n2094 585
R2627 gnd.n3606 gnd.n3605 585
R2628 gnd.n3605 gnd.n3604 585
R2629 gnd.n2097 gnd.n2096 585
R2630 gnd.n3558 gnd.n2097 585
R2631 gnd.n3592 gnd.n3591 585
R2632 gnd.n3593 gnd.n3592 585
R2633 gnd.n3590 gnd.n2110 585
R2634 gnd.n2110 gnd.n2106 585
R2635 gnd.n3589 gnd.n3588 585
R2636 gnd.n3588 gnd.n3587 585
R2637 gnd.n2112 gnd.n2111 585
R2638 gnd.n3548 gnd.n2112 585
R2639 gnd.n3533 gnd.n3532 585
R2640 gnd.n3532 gnd.n2122 585
R2641 gnd.n3534 gnd.n2132 585
R2642 gnd.n3517 gnd.n2132 585
R2643 gnd.n3536 gnd.n3535 585
R2644 gnd.n3537 gnd.n3536 585
R2645 gnd.n3531 gnd.n2131 585
R2646 gnd.n2131 gnd.n2128 585
R2647 gnd.n3530 gnd.n3529 585
R2648 gnd.n3529 gnd.n3528 585
R2649 gnd.n2134 gnd.n2133 585
R2650 gnd.n3508 gnd.n2134 585
R2651 gnd.n3493 gnd.n3492 585
R2652 gnd.n3492 gnd.n2145 585
R2653 gnd.n3494 gnd.n2155 585
R2654 gnd.n3481 gnd.n2155 585
R2655 gnd.n3496 gnd.n3495 585
R2656 gnd.n3497 gnd.n3496 585
R2657 gnd.n3491 gnd.n2154 585
R2658 gnd.n2154 gnd.n2151 585
R2659 gnd.n3490 gnd.n3489 585
R2660 gnd.n3489 gnd.n3488 585
R2661 gnd.n2157 gnd.n2156 585
R2662 gnd.n2170 gnd.n2157 585
R2663 gnd.n3466 gnd.n3465 585
R2664 gnd.n3467 gnd.n3466 585
R2665 gnd.n3464 gnd.n2172 585
R2666 gnd.n3459 gnd.n2172 585
R2667 gnd.n3463 gnd.n3462 585
R2668 gnd.n3462 gnd.n3461 585
R2669 gnd.n2174 gnd.n2173 585
R2670 gnd.n3445 gnd.n2174 585
R2671 gnd.n3433 gnd.n2192 585
R2672 gnd.n2192 gnd.n2184 585
R2673 gnd.n3435 gnd.n3434 585
R2674 gnd.n3436 gnd.n3435 585
R2675 gnd.n3432 gnd.n2191 585
R2676 gnd.n3377 gnd.n2191 585
R2677 gnd.n3431 gnd.n3430 585
R2678 gnd.n3430 gnd.n3429 585
R2679 gnd.n2194 gnd.n2193 585
R2680 gnd.n3403 gnd.n2194 585
R2681 gnd.n3416 gnd.n3415 585
R2682 gnd.n3417 gnd.n3416 585
R2683 gnd.n3414 gnd.n2205 585
R2684 gnd.n3409 gnd.n2205 585
R2685 gnd.n3413 gnd.n3412 585
R2686 gnd.n3412 gnd.n3411 585
R2687 gnd.n2207 gnd.n2206 585
R2688 gnd.n3398 gnd.n2207 585
R2689 gnd.n3350 gnd.n3347 585
R2690 gnd.n3350 gnd.n3349 585
R2691 gnd.n3351 gnd.n3346 585
R2692 gnd.n3351 gnd.n2221 585
R2693 gnd.n3353 gnd.n3352 585
R2694 gnd.n3352 gnd.n2220 585
R2695 gnd.n3354 gnd.n2232 585
R2696 gnd.n3334 gnd.n2232 585
R2697 gnd.n3356 gnd.n3355 585
R2698 gnd.n3357 gnd.n3356 585
R2699 gnd.n3345 gnd.n2231 585
R2700 gnd.n3340 gnd.n2231 585
R2701 gnd.n3344 gnd.n3343 585
R2702 gnd.n3343 gnd.n3342 585
R2703 gnd.n2234 gnd.n2233 585
R2704 gnd.n3325 gnd.n2234 585
R2705 gnd.n2257 gnd.n2256 585
R2706 gnd.n3300 gnd.n2257 585
R2707 gnd.n3304 gnd.n3303 585
R2708 gnd.n3303 gnd.n3302 585
R2709 gnd.n3305 gnd.n2246 585
R2710 gnd.n3316 gnd.n2246 585
R2711 gnd.n3306 gnd.n2254 585
R2712 gnd.n2258 gnd.n2254 585
R2713 gnd.n3308 gnd.n3307 585
R2714 gnd.n3309 gnd.n3308 585
R2715 gnd.n2255 gnd.n2253 585
R2716 gnd.n3282 gnd.n2253 585
R2717 gnd.n3275 gnd.n3274 585
R2718 gnd.n3276 gnd.n3275 585
R2719 gnd.n3273 gnd.n2268 585
R2720 gnd.n2268 gnd.n1504 585
R2721 gnd.n3272 gnd.n3271 585
R2722 gnd.n3271 gnd.n1502 585
R2723 gnd.n3270 gnd.n2269 585
R2724 gnd.n3270 gnd.n3269 585
R2725 gnd.n1490 gnd.n1489 585
R2726 gnd.n2349 gnd.n1490 585
R2727 gnd.n4783 gnd.n4782 585
R2728 gnd.n4782 gnd.n4781 585
R2729 gnd.n4784 gnd.n1468 585
R2730 gnd.n2355 gnd.n1468 585
R2731 gnd.n4849 gnd.n4848 585
R2732 gnd.n4847 gnd.n1467 585
R2733 gnd.n4846 gnd.n1466 585
R2734 gnd.n4851 gnd.n1466 585
R2735 gnd.n4845 gnd.n4844 585
R2736 gnd.n4843 gnd.n4842 585
R2737 gnd.n4841 gnd.n4840 585
R2738 gnd.n4839 gnd.n4838 585
R2739 gnd.n4837 gnd.n4836 585
R2740 gnd.n4835 gnd.n4834 585
R2741 gnd.n4833 gnd.n4832 585
R2742 gnd.n4831 gnd.n4830 585
R2743 gnd.n4829 gnd.n4828 585
R2744 gnd.n4827 gnd.n4826 585
R2745 gnd.n4825 gnd.n4824 585
R2746 gnd.n4823 gnd.n4822 585
R2747 gnd.n4821 gnd.n4820 585
R2748 gnd.n4819 gnd.n4818 585
R2749 gnd.n4817 gnd.n4816 585
R2750 gnd.n4815 gnd.n4814 585
R2751 gnd.n4813 gnd.n4812 585
R2752 gnd.n4811 gnd.n4810 585
R2753 gnd.n4809 gnd.n4808 585
R2754 gnd.n4807 gnd.n4806 585
R2755 gnd.n4805 gnd.n4804 585
R2756 gnd.n4803 gnd.n4802 585
R2757 gnd.n4801 gnd.n4800 585
R2758 gnd.n4799 gnd.n4798 585
R2759 gnd.n4797 gnd.n4796 585
R2760 gnd.n4795 gnd.n4794 585
R2761 gnd.n4793 gnd.n4792 585
R2762 gnd.n4791 gnd.n4790 585
R2763 gnd.n4789 gnd.n1430 585
R2764 gnd.n4854 gnd.n4853 585
R2765 gnd.n1432 gnd.n1429 585
R2766 gnd.n2282 gnd.n2281 585
R2767 gnd.n2284 gnd.n2283 585
R2768 gnd.n2287 gnd.n2286 585
R2769 gnd.n2289 gnd.n2288 585
R2770 gnd.n2291 gnd.n2290 585
R2771 gnd.n2293 gnd.n2292 585
R2772 gnd.n2295 gnd.n2294 585
R2773 gnd.n2297 gnd.n2296 585
R2774 gnd.n2299 gnd.n2298 585
R2775 gnd.n2301 gnd.n2300 585
R2776 gnd.n2303 gnd.n2302 585
R2777 gnd.n2305 gnd.n2304 585
R2778 gnd.n2307 gnd.n2306 585
R2779 gnd.n2309 gnd.n2308 585
R2780 gnd.n2311 gnd.n2310 585
R2781 gnd.n2313 gnd.n2312 585
R2782 gnd.n2315 gnd.n2314 585
R2783 gnd.n2317 gnd.n2316 585
R2784 gnd.n2319 gnd.n2318 585
R2785 gnd.n2321 gnd.n2320 585
R2786 gnd.n2323 gnd.n2322 585
R2787 gnd.n2325 gnd.n2324 585
R2788 gnd.n2327 gnd.n2326 585
R2789 gnd.n2329 gnd.n2328 585
R2790 gnd.n2331 gnd.n2330 585
R2791 gnd.n2333 gnd.n2332 585
R2792 gnd.n2335 gnd.n2334 585
R2793 gnd.n2337 gnd.n2336 585
R2794 gnd.n2339 gnd.n2338 585
R2795 gnd.n2341 gnd.n2340 585
R2796 gnd.n2342 gnd.n2278 585
R2797 gnd.n4182 gnd.n4181 585
R2798 gnd.n4184 gnd.n4183 585
R2799 gnd.n4186 gnd.n4185 585
R2800 gnd.n4188 gnd.n4187 585
R2801 gnd.n4190 gnd.n4189 585
R2802 gnd.n4192 gnd.n4191 585
R2803 gnd.n4194 gnd.n4193 585
R2804 gnd.n4196 gnd.n4195 585
R2805 gnd.n4198 gnd.n4197 585
R2806 gnd.n4200 gnd.n4199 585
R2807 gnd.n4202 gnd.n4201 585
R2808 gnd.n4204 gnd.n4203 585
R2809 gnd.n4206 gnd.n4205 585
R2810 gnd.n4208 gnd.n4207 585
R2811 gnd.n4210 gnd.n4209 585
R2812 gnd.n4212 gnd.n4211 585
R2813 gnd.n4214 gnd.n4213 585
R2814 gnd.n4216 gnd.n4215 585
R2815 gnd.n4218 gnd.n4217 585
R2816 gnd.n4220 gnd.n4219 585
R2817 gnd.n4222 gnd.n4221 585
R2818 gnd.n4224 gnd.n4223 585
R2819 gnd.n4226 gnd.n4225 585
R2820 gnd.n4228 gnd.n4227 585
R2821 gnd.n4230 gnd.n4229 585
R2822 gnd.n4232 gnd.n4231 585
R2823 gnd.n4234 gnd.n4233 585
R2824 gnd.n4236 gnd.n4235 585
R2825 gnd.n4238 gnd.n4237 585
R2826 gnd.n4240 gnd.n1897 585
R2827 gnd.n4242 gnd.n4241 585
R2828 gnd.n4244 gnd.n1861 585
R2829 gnd.n4246 gnd.n4245 585
R2830 gnd.n4249 gnd.n4248 585
R2831 gnd.n1864 gnd.n1862 585
R2832 gnd.n4115 gnd.n4114 585
R2833 gnd.n4117 gnd.n4116 585
R2834 gnd.n4120 gnd.n4119 585
R2835 gnd.n4122 gnd.n4121 585
R2836 gnd.n4124 gnd.n4123 585
R2837 gnd.n4126 gnd.n4125 585
R2838 gnd.n4128 gnd.n4127 585
R2839 gnd.n4130 gnd.n4129 585
R2840 gnd.n4132 gnd.n4131 585
R2841 gnd.n4134 gnd.n4133 585
R2842 gnd.n4136 gnd.n4135 585
R2843 gnd.n4138 gnd.n4137 585
R2844 gnd.n4140 gnd.n4139 585
R2845 gnd.n4142 gnd.n4141 585
R2846 gnd.n4144 gnd.n4143 585
R2847 gnd.n4146 gnd.n4145 585
R2848 gnd.n4148 gnd.n4147 585
R2849 gnd.n4150 gnd.n4149 585
R2850 gnd.n4152 gnd.n4151 585
R2851 gnd.n4154 gnd.n4153 585
R2852 gnd.n4156 gnd.n4155 585
R2853 gnd.n4158 gnd.n4157 585
R2854 gnd.n4160 gnd.n4159 585
R2855 gnd.n4162 gnd.n4161 585
R2856 gnd.n4164 gnd.n4163 585
R2857 gnd.n4166 gnd.n4165 585
R2858 gnd.n4168 gnd.n4167 585
R2859 gnd.n4170 gnd.n4169 585
R2860 gnd.n4172 gnd.n4171 585
R2861 gnd.n4174 gnd.n4173 585
R2862 gnd.n4175 gnd.n1904 585
R2863 gnd.n4180 gnd.n1900 585
R2864 gnd.n4180 gnd.n4179 585
R2865 gnd.n3856 gnd.n1901 585
R2866 gnd.n1910 gnd.n1901 585
R2867 gnd.n3857 gnd.n1908 585
R2868 gnd.n4089 gnd.n1908 585
R2869 gnd.n3859 gnd.n3858 585
R2870 gnd.n3860 gnd.n3859 585
R2871 gnd.n3855 gnd.n1948 585
R2872 gnd.n1948 gnd.n1947 585
R2873 gnd.n3854 gnd.n3853 585
R2874 gnd.n3853 gnd.n3852 585
R2875 gnd.n1950 gnd.n1949 585
R2876 gnd.n3842 gnd.n1950 585
R2877 gnd.n3813 gnd.n1957 585
R2878 gnd.n3845 gnd.n1957 585
R2879 gnd.n3814 gnd.n1967 585
R2880 gnd.n3829 gnd.n1967 585
R2881 gnd.n3815 gnd.n1978 585
R2882 gnd.n1978 gnd.n1966 585
R2883 gnd.n3817 gnd.n3816 585
R2884 gnd.n3818 gnd.n3817 585
R2885 gnd.n3812 gnd.n1977 585
R2886 gnd.n1977 gnd.n1974 585
R2887 gnd.n3811 gnd.n3810 585
R2888 gnd.n3810 gnd.n3809 585
R2889 gnd.n1980 gnd.n1979 585
R2890 gnd.n3797 gnd.n1980 585
R2891 gnd.n3780 gnd.n1988 585
R2892 gnd.n3799 gnd.n1988 585
R2893 gnd.n3782 gnd.n3781 585
R2894 gnd.n3784 gnd.n3782 585
R2895 gnd.n3779 gnd.n1998 585
R2896 gnd.n1998 gnd.n1996 585
R2897 gnd.n3778 gnd.n3777 585
R2898 gnd.n3777 gnd.n3776 585
R2899 gnd.n2000 gnd.n1999 585
R2900 gnd.n2008 gnd.n2000 585
R2901 gnd.n3649 gnd.n2006 585
R2902 gnd.n3769 gnd.n2006 585
R2903 gnd.n3652 gnd.n3651 585
R2904 gnd.n3651 gnd.n3650 585
R2905 gnd.n3653 gnd.n2018 585
R2906 gnd.n3758 gnd.n2018 585
R2907 gnd.n3655 gnd.n3654 585
R2908 gnd.n3654 gnd.n2016 585
R2909 gnd.n3656 gnd.n2023 585
R2910 gnd.n3752 gnd.n2023 585
R2911 gnd.n3662 gnd.n3661 585
R2912 gnd.n3661 gnd.n3660 585
R2913 gnd.n3663 gnd.n2031 585
R2914 gnd.n3727 gnd.n2031 585
R2915 gnd.n3665 gnd.n3664 585
R2916 gnd.n3664 gnd.n2030 585
R2917 gnd.n3666 gnd.n2037 585
R2918 gnd.n3721 gnd.n2037 585
R2919 gnd.n3669 gnd.n3668 585
R2920 gnd.n3668 gnd.n3667 585
R2921 gnd.n3670 gnd.n2044 585
R2922 gnd.n3708 gnd.n2044 585
R2923 gnd.n3671 gnd.n2051 585
R2924 gnd.n3700 gnd.n2051 585
R2925 gnd.n3672 gnd.n2050 585
R2926 gnd.n3702 gnd.n2050 585
R2927 gnd.n3674 gnd.n3673 585
R2928 gnd.n3674 gnd.n2060 585
R2929 gnd.n3676 gnd.n3675 585
R2930 gnd.n3675 gnd.n2059 585
R2931 gnd.n3677 gnd.n2069 585
R2932 gnd.n3638 gnd.n2069 585
R2933 gnd.n3679 gnd.n3678 585
R2934 gnd.n3680 gnd.n3679 585
R2935 gnd.n3648 gnd.n2068 585
R2936 gnd.n3566 gnd.n2068 585
R2937 gnd.n3647 gnd.n3646 585
R2938 gnd.n3646 gnd.n3645 585
R2939 gnd.n2071 gnd.n2070 585
R2940 gnd.n3629 gnd.n2071 585
R2941 gnd.n3615 gnd.n2079 585
R2942 gnd.n3631 gnd.n2079 585
R2943 gnd.n3617 gnd.n3616 585
R2944 gnd.n3618 gnd.n3617 585
R2945 gnd.n3614 gnd.n2088 585
R2946 gnd.n2088 gnd.n2086 585
R2947 gnd.n3613 gnd.n3612 585
R2948 gnd.n3612 gnd.n3611 585
R2949 gnd.n2090 gnd.n2089 585
R2950 gnd.n2099 gnd.n2090 585
R2951 gnd.n3555 gnd.n2098 585
R2952 gnd.n3604 gnd.n2098 585
R2953 gnd.n3557 gnd.n3556 585
R2954 gnd.n3558 gnd.n3557 585
R2955 gnd.n3554 gnd.n2108 585
R2956 gnd.n3593 gnd.n2108 585
R2957 gnd.n3553 gnd.n3552 585
R2958 gnd.n3552 gnd.n2106 585
R2959 gnd.n3551 gnd.n2114 585
R2960 gnd.n3587 gnd.n2114 585
R2961 gnd.n3550 gnd.n3549 585
R2962 gnd.n3549 gnd.n3548 585
R2963 gnd.n2121 gnd.n2120 585
R2964 gnd.n2122 gnd.n2121 585
R2965 gnd.n3516 gnd.n3515 585
R2966 gnd.n3517 gnd.n3516 585
R2967 gnd.n3514 gnd.n2129 585
R2968 gnd.n3537 gnd.n2129 585
R2969 gnd.n3513 gnd.n3512 585
R2970 gnd.n3512 gnd.n2128 585
R2971 gnd.n3511 gnd.n2136 585
R2972 gnd.n3528 gnd.n2136 585
R2973 gnd.n3510 gnd.n3509 585
R2974 gnd.n3509 gnd.n3508 585
R2975 gnd.n2144 gnd.n2143 585
R2976 gnd.n2145 gnd.n2144 585
R2977 gnd.n3483 gnd.n3482 585
R2978 gnd.n3482 gnd.n3481 585
R2979 gnd.n3484 gnd.n2152 585
R2980 gnd.n3497 gnd.n2152 585
R2981 gnd.n3485 gnd.n2160 585
R2982 gnd.n2160 gnd.n2151 585
R2983 gnd.n3487 gnd.n3486 585
R2984 gnd.n3488 gnd.n3487 585
R2985 gnd.n2161 gnd.n2159 585
R2986 gnd.n2170 gnd.n2159 585
R2987 gnd.n3440 gnd.n2169 585
R2988 gnd.n3467 gnd.n2169 585
R2989 gnd.n3441 gnd.n2177 585
R2990 gnd.n3459 gnd.n2177 585
R2991 gnd.n3442 gnd.n2176 585
R2992 gnd.n3461 gnd.n2176 585
R2993 gnd.n3444 gnd.n3443 585
R2994 gnd.n3445 gnd.n3444 585
R2995 gnd.n3439 gnd.n2186 585
R2996 gnd.n2186 gnd.n2184 585
R2997 gnd.n3438 gnd.n3437 585
R2998 gnd.n3437 gnd.n3436 585
R2999 gnd.n2188 gnd.n2187 585
R3000 gnd.n3377 gnd.n2188 585
R3001 gnd.n3402 gnd.n2196 585
R3002 gnd.n3429 gnd.n2196 585
R3003 gnd.n3405 gnd.n3404 585
R3004 gnd.n3404 gnd.n3403 585
R3005 gnd.n3406 gnd.n2203 585
R3006 gnd.n3417 gnd.n2203 585
R3007 gnd.n3408 gnd.n3407 585
R3008 gnd.n3409 gnd.n3408 585
R3009 gnd.n3401 gnd.n2209 585
R3010 gnd.n3411 gnd.n2209 585
R3011 gnd.n3400 gnd.n3399 585
R3012 gnd.n3399 gnd.n3398 585
R3013 gnd.n2212 gnd.n2211 585
R3014 gnd.n3349 gnd.n2212 585
R3015 gnd.n3331 gnd.n3330 585
R3016 gnd.n3331 gnd.n2221 585
R3017 gnd.n3332 gnd.n3329 585
R3018 gnd.n3332 gnd.n2220 585
R3019 gnd.n3336 gnd.n3335 585
R3020 gnd.n3335 gnd.n3334 585
R3021 gnd.n3337 gnd.n2229 585
R3022 gnd.n3357 gnd.n2229 585
R3023 gnd.n3339 gnd.n3338 585
R3024 gnd.n3340 gnd.n3339 585
R3025 gnd.n3328 gnd.n2236 585
R3026 gnd.n3342 gnd.n2236 585
R3027 gnd.n3327 gnd.n3326 585
R3028 gnd.n3326 gnd.n3325 585
R3029 gnd.n2238 gnd.n2237 585
R3030 gnd.n3300 gnd.n2238 585
R3031 gnd.n3313 gnd.n2248 585
R3032 gnd.n3302 gnd.n2248 585
R3033 gnd.n3315 gnd.n3314 585
R3034 gnd.n3316 gnd.n3315 585
R3035 gnd.n3312 gnd.n2247 585
R3036 gnd.n2258 gnd.n2247 585
R3037 gnd.n3311 gnd.n3310 585
R3038 gnd.n3310 gnd.n3309 585
R3039 gnd.n2250 gnd.n2249 585
R3040 gnd.n3282 gnd.n2250 585
R3041 gnd.n2343 gnd.n2267 585
R3042 gnd.n3276 gnd.n2267 585
R3043 gnd.n2345 gnd.n2344 585
R3044 gnd.n2345 gnd.n1504 585
R3045 gnd.n2347 gnd.n2346 585
R3046 gnd.n2346 gnd.n1502 585
R3047 gnd.n2348 gnd.n2271 585
R3048 gnd.n3269 gnd.n2271 585
R3049 gnd.n2351 gnd.n2350 585
R3050 gnd.n2350 gnd.n2349 585
R3051 gnd.n2352 gnd.n1492 585
R3052 gnd.n4781 gnd.n1492 585
R3053 gnd.n2354 gnd.n2353 585
R3054 gnd.n2355 gnd.n2354 585
R3055 gnd.n4905 gnd.n4904 585
R3056 gnd.n4906 gnd.n4905 585
R3057 gnd.n1363 gnd.n1362 585
R3058 gnd.n2883 gnd.n1363 585
R3059 gnd.n4914 gnd.n4913 585
R3060 gnd.n4913 gnd.n4912 585
R3061 gnd.n4915 gnd.n1357 585
R3062 gnd.n2876 gnd.n1357 585
R3063 gnd.n4917 gnd.n4916 585
R3064 gnd.n4918 gnd.n4917 585
R3065 gnd.n1343 gnd.n1342 585
R3066 gnd.n2871 gnd.n1343 585
R3067 gnd.n4926 gnd.n4925 585
R3068 gnd.n4925 gnd.n4924 585
R3069 gnd.n4927 gnd.n1337 585
R3070 gnd.n2898 gnd.n1337 585
R3071 gnd.n4929 gnd.n4928 585
R3072 gnd.n4930 gnd.n4929 585
R3073 gnd.n1322 gnd.n1321 585
R3074 gnd.n2864 gnd.n1322 585
R3075 gnd.n4938 gnd.n4937 585
R3076 gnd.n4937 gnd.n4936 585
R3077 gnd.n4939 gnd.n1316 585
R3078 gnd.n2856 gnd.n1316 585
R3079 gnd.n4941 gnd.n4940 585
R3080 gnd.n4942 gnd.n4941 585
R3081 gnd.n1303 gnd.n1302 585
R3082 gnd.n2849 gnd.n1303 585
R3083 gnd.n4950 gnd.n4949 585
R3084 gnd.n4949 gnd.n4948 585
R3085 gnd.n4951 gnd.n1297 585
R3086 gnd.n2841 gnd.n1297 585
R3087 gnd.n4953 gnd.n4952 585
R3088 gnd.n4954 gnd.n4953 585
R3089 gnd.n1282 gnd.n1281 585
R3090 gnd.n2788 gnd.n1282 585
R3091 gnd.n4962 gnd.n4961 585
R3092 gnd.n4961 gnd.n4960 585
R3093 gnd.n4963 gnd.n1277 585
R3094 gnd.n2779 gnd.n1277 585
R3095 gnd.n4965 gnd.n4964 585
R3096 gnd.n4966 gnd.n4965 585
R3097 gnd.n1262 gnd.n1260 585
R3098 gnd.n2773 gnd.n1262 585
R3099 gnd.n4974 gnd.n4973 585
R3100 gnd.n4973 gnd.n4972 585
R3101 gnd.n1261 gnd.n1259 585
R3102 gnd.n2802 gnd.n1261 585
R3103 gnd.n2765 gnd.n2764 585
R3104 gnd.n2766 gnd.n2765 585
R3105 gnd.n2763 gnd.n2762 585
R3106 gnd.n2762 gnd.n2761 585
R3107 gnd.n2749 gnd.n2476 585
R3108 gnd.n2741 gnd.n2476 585
R3109 gnd.n2751 gnd.n2750 585
R3110 gnd.n2752 gnd.n2751 585
R3111 gnd.n2748 gnd.n2487 585
R3112 gnd.n2748 gnd.n2747 585
R3113 gnd.n2486 gnd.n1258 585
R3114 gnd.n2715 gnd.n2486 585
R3115 gnd.n2722 gnd.n1252 585
R3116 gnd.n2723 gnd.n2722 585
R3117 gnd.n4977 gnd.n1249 585
R3118 gnd.n2503 gnd.n1249 585
R3119 gnd.n4979 gnd.n4978 585
R3120 gnd.n4980 gnd.n4979 585
R3121 gnd.n1234 gnd.n1233 585
R3122 gnd.n2704 gnd.n1234 585
R3123 gnd.n4988 gnd.n4987 585
R3124 gnd.n4987 gnd.n4986 585
R3125 gnd.n4989 gnd.n1228 585
R3126 gnd.n2697 gnd.n1228 585
R3127 gnd.n4991 gnd.n4990 585
R3128 gnd.n4992 gnd.n4991 585
R3129 gnd.n1214 gnd.n1213 585
R3130 gnd.n2688 gnd.n1214 585
R3131 gnd.n5000 gnd.n4999 585
R3132 gnd.n4999 gnd.n4998 585
R3133 gnd.n5001 gnd.n1208 585
R3134 gnd.n2682 gnd.n1208 585
R3135 gnd.n5003 gnd.n5002 585
R3136 gnd.n5004 gnd.n5003 585
R3137 gnd.n1193 gnd.n1192 585
R3138 gnd.n2635 gnd.n1193 585
R3139 gnd.n5012 gnd.n5011 585
R3140 gnd.n5011 gnd.n5010 585
R3141 gnd.n5013 gnd.n1187 585
R3142 gnd.n2629 gnd.n1187 585
R3143 gnd.n5015 gnd.n5014 585
R3144 gnd.n5016 gnd.n5015 585
R3145 gnd.n1174 gnd.n1173 585
R3146 gnd.n1177 gnd.n1174 585
R3147 gnd.n5024 gnd.n5023 585
R3148 gnd.n5023 gnd.n5022 585
R3149 gnd.n5025 gnd.n1168 585
R3150 gnd.n1168 gnd.n1167 585
R3151 gnd.n5027 gnd.n5026 585
R3152 gnd.n5028 gnd.n5027 585
R3153 gnd.n1151 gnd.n1150 585
R3154 gnd.n1155 gnd.n1151 585
R3155 gnd.n5036 gnd.n5035 585
R3156 gnd.n5035 gnd.n5034 585
R3157 gnd.n5037 gnd.n1144 585
R3158 gnd.n1152 gnd.n1144 585
R3159 gnd.n5039 gnd.n5038 585
R3160 gnd.n5040 gnd.n5039 585
R3161 gnd.n1145 gnd.n1071 585
R3162 gnd.n1071 gnd.n1068 585
R3163 gnd.n5162 gnd.n5161 585
R3164 gnd.n5160 gnd.n1070 585
R3165 gnd.n5159 gnd.n1069 585
R3166 gnd.n5164 gnd.n1069 585
R3167 gnd.n5158 gnd.n5157 585
R3168 gnd.n5156 gnd.n5155 585
R3169 gnd.n5154 gnd.n5153 585
R3170 gnd.n5152 gnd.n5151 585
R3171 gnd.n5150 gnd.n5149 585
R3172 gnd.n5148 gnd.n5147 585
R3173 gnd.n5146 gnd.n5145 585
R3174 gnd.n5144 gnd.n5143 585
R3175 gnd.n5142 gnd.n5141 585
R3176 gnd.n5140 gnd.n5139 585
R3177 gnd.n5138 gnd.n5137 585
R3178 gnd.n5136 gnd.n5135 585
R3179 gnd.n5134 gnd.n5133 585
R3180 gnd.n5132 gnd.n5131 585
R3181 gnd.n5130 gnd.n5129 585
R3182 gnd.n5127 gnd.n5126 585
R3183 gnd.n5125 gnd.n5124 585
R3184 gnd.n5123 gnd.n5122 585
R3185 gnd.n5121 gnd.n5120 585
R3186 gnd.n5119 gnd.n5118 585
R3187 gnd.n5117 gnd.n5116 585
R3188 gnd.n5115 gnd.n5114 585
R3189 gnd.n5113 gnd.n5112 585
R3190 gnd.n5111 gnd.n5110 585
R3191 gnd.n5109 gnd.n5108 585
R3192 gnd.n5107 gnd.n5106 585
R3193 gnd.n5105 gnd.n5104 585
R3194 gnd.n5103 gnd.n5102 585
R3195 gnd.n5101 gnd.n5100 585
R3196 gnd.n5099 gnd.n5098 585
R3197 gnd.n5097 gnd.n5096 585
R3198 gnd.n5095 gnd.n5094 585
R3199 gnd.n5093 gnd.n5092 585
R3200 gnd.n5091 gnd.n5090 585
R3201 gnd.n5089 gnd.n5088 585
R3202 gnd.n5087 gnd.n5086 585
R3203 gnd.n5085 gnd.n5084 585
R3204 gnd.n5083 gnd.n5082 585
R3205 gnd.n5081 gnd.n5080 585
R3206 gnd.n5079 gnd.n5078 585
R3207 gnd.n5077 gnd.n5076 585
R3208 gnd.n5075 gnd.n5074 585
R3209 gnd.n5073 gnd.n5072 585
R3210 gnd.n5071 gnd.n5070 585
R3211 gnd.n5069 gnd.n5068 585
R3212 gnd.n5067 gnd.n5066 585
R3213 gnd.n5065 gnd.n5064 585
R3214 gnd.n5063 gnd.n5062 585
R3215 gnd.n5061 gnd.n5060 585
R3216 gnd.n5059 gnd.n5058 585
R3217 gnd.n5057 gnd.n5056 585
R3218 gnd.n5055 gnd.n5054 585
R3219 gnd.n5053 gnd.n5052 585
R3220 gnd.n5051 gnd.n5050 585
R3221 gnd.n5049 gnd.n5048 585
R3222 gnd.n1140 gnd.n1133 585
R3223 gnd.n3058 gnd.n3057 585
R3224 gnd.n3055 gnd.n2951 585
R3225 gnd.n3054 gnd.n3053 585
R3226 gnd.n3047 gnd.n2953 585
R3227 gnd.n3049 gnd.n3048 585
R3228 gnd.n3045 gnd.n2955 585
R3229 gnd.n3044 gnd.n3043 585
R3230 gnd.n3037 gnd.n2957 585
R3231 gnd.n3039 gnd.n3038 585
R3232 gnd.n3035 gnd.n2959 585
R3233 gnd.n3034 gnd.n3033 585
R3234 gnd.n3027 gnd.n2961 585
R3235 gnd.n3029 gnd.n3028 585
R3236 gnd.n3025 gnd.n2963 585
R3237 gnd.n3024 gnd.n3023 585
R3238 gnd.n3017 gnd.n2965 585
R3239 gnd.n3019 gnd.n3018 585
R3240 gnd.n3015 gnd.n2967 585
R3241 gnd.n3014 gnd.n3013 585
R3242 gnd.n3007 gnd.n2969 585
R3243 gnd.n3009 gnd.n3008 585
R3244 gnd.n3005 gnd.n2973 585
R3245 gnd.n3004 gnd.n3003 585
R3246 gnd.n2997 gnd.n2975 585
R3247 gnd.n2999 gnd.n2998 585
R3248 gnd.n2995 gnd.n2977 585
R3249 gnd.n2994 gnd.n2993 585
R3250 gnd.n2987 gnd.n2979 585
R3251 gnd.n2989 gnd.n2988 585
R3252 gnd.n2985 gnd.n2982 585
R3253 gnd.n2984 gnd.n1425 585
R3254 gnd.n4856 gnd.n1421 585
R3255 gnd.n4858 gnd.n4857 585
R3256 gnd.n4860 gnd.n1419 585
R3257 gnd.n4862 gnd.n4861 585
R3258 gnd.n4863 gnd.n1414 585
R3259 gnd.n4865 gnd.n4864 585
R3260 gnd.n4867 gnd.n1412 585
R3261 gnd.n4869 gnd.n4868 585
R3262 gnd.n4871 gnd.n1405 585
R3263 gnd.n4873 gnd.n4872 585
R3264 gnd.n4875 gnd.n1403 585
R3265 gnd.n4877 gnd.n4876 585
R3266 gnd.n4878 gnd.n1398 585
R3267 gnd.n4880 gnd.n4879 585
R3268 gnd.n4882 gnd.n1396 585
R3269 gnd.n4884 gnd.n4883 585
R3270 gnd.n4885 gnd.n1391 585
R3271 gnd.n4887 gnd.n4886 585
R3272 gnd.n4889 gnd.n1389 585
R3273 gnd.n4891 gnd.n4890 585
R3274 gnd.n4892 gnd.n1383 585
R3275 gnd.n4894 gnd.n4893 585
R3276 gnd.n4896 gnd.n1382 585
R3277 gnd.n4897 gnd.n1380 585
R3278 gnd.n4900 gnd.n4899 585
R3279 gnd.n4901 gnd.n1377 585
R3280 gnd.n1381 gnd.n1377 585
R3281 gnd.n2880 gnd.n1374 585
R3282 gnd.n4906 gnd.n1374 585
R3283 gnd.n2882 gnd.n2881 585
R3284 gnd.n2883 gnd.n2882 585
R3285 gnd.n2879 gnd.n1365 585
R3286 gnd.n4912 gnd.n1365 585
R3287 gnd.n2878 gnd.n2877 585
R3288 gnd.n2877 gnd.n2876 585
R3289 gnd.n2874 gnd.n1354 585
R3290 gnd.n4918 gnd.n1354 585
R3291 gnd.n2873 gnd.n2872 585
R3292 gnd.n2872 gnd.n2871 585
R3293 gnd.n2870 gnd.n1344 585
R3294 gnd.n4924 gnd.n1344 585
R3295 gnd.n2869 gnd.n2430 585
R3296 gnd.n2898 gnd.n2430 585
R3297 gnd.n2867 gnd.n1334 585
R3298 gnd.n4930 gnd.n1334 585
R3299 gnd.n2866 gnd.n2865 585
R3300 gnd.n2865 gnd.n2864 585
R3301 gnd.n2439 gnd.n1324 585
R3302 gnd.n4936 gnd.n1324 585
R3303 gnd.n2855 gnd.n2854 585
R3304 gnd.n2856 gnd.n2855 585
R3305 gnd.n2852 gnd.n1314 585
R3306 gnd.n4942 gnd.n1314 585
R3307 gnd.n2851 gnd.n2850 585
R3308 gnd.n2850 gnd.n2849 585
R3309 gnd.n2444 gnd.n1304 585
R3310 gnd.n4948 gnd.n1304 585
R3311 gnd.n2784 gnd.n2448 585
R3312 gnd.n2841 gnd.n2448 585
R3313 gnd.n2785 gnd.n1294 585
R3314 gnd.n4954 gnd.n1294 585
R3315 gnd.n2787 gnd.n2786 585
R3316 gnd.n2788 gnd.n2787 585
R3317 gnd.n2782 gnd.n1284 585
R3318 gnd.n4960 gnd.n1284 585
R3319 gnd.n2781 gnd.n2780 585
R3320 gnd.n2780 gnd.n2779 585
R3321 gnd.n2776 gnd.n1275 585
R3322 gnd.n4966 gnd.n1275 585
R3323 gnd.n2775 gnd.n2774 585
R3324 gnd.n2774 gnd.n2773 585
R3325 gnd.n2772 gnd.n1263 585
R3326 gnd.n4972 gnd.n1263 585
R3327 gnd.n2771 gnd.n2461 585
R3328 gnd.n2802 gnd.n2461 585
R3329 gnd.n2475 gnd.n2470 585
R3330 gnd.n2766 gnd.n2475 585
R3331 gnd.n2511 gnd.n2477 585
R3332 gnd.n2761 gnd.n2477 585
R3333 gnd.n2512 gnd.n2496 585
R3334 gnd.n2741 gnd.n2496 585
R3335 gnd.n2513 gnd.n2483 585
R3336 gnd.n2752 gnd.n2483 585
R3337 gnd.n2514 gnd.n2489 585
R3338 gnd.n2747 gnd.n2489 585
R3339 gnd.n2717 gnd.n2716 585
R3340 gnd.n2716 gnd.n2715 585
R3341 gnd.n2718 gnd.n2504 585
R3342 gnd.n2723 gnd.n2504 585
R3343 gnd.n2510 gnd.n2509 585
R3344 gnd.n2509 gnd.n2503 585
R3345 gnd.n2701 gnd.n1246 585
R3346 gnd.n4980 gnd.n1246 585
R3347 gnd.n2703 gnd.n2702 585
R3348 gnd.n2704 gnd.n2703 585
R3349 gnd.n2700 gnd.n1236 585
R3350 gnd.n4986 gnd.n1236 585
R3351 gnd.n2699 gnd.n2698 585
R3352 gnd.n2698 gnd.n2697 585
R3353 gnd.n2519 gnd.n1225 585
R3354 gnd.n4992 gnd.n1225 585
R3355 gnd.n2687 gnd.n2686 585
R3356 gnd.n2688 gnd.n2687 585
R3357 gnd.n2685 gnd.n1215 585
R3358 gnd.n4998 gnd.n1215 585
R3359 gnd.n2684 gnd.n2683 585
R3360 gnd.n2683 gnd.n2682 585
R3361 gnd.n2524 gnd.n1205 585
R3362 gnd.n5004 gnd.n1205 585
R3363 gnd.n2634 gnd.n2633 585
R3364 gnd.n2635 gnd.n2634 585
R3365 gnd.n2632 gnd.n1195 585
R3366 gnd.n5010 gnd.n1195 585
R3367 gnd.n2631 gnd.n2630 585
R3368 gnd.n2630 gnd.n2629 585
R3369 gnd.n2541 gnd.n1185 585
R3370 gnd.n5016 gnd.n1185 585
R3371 gnd.n2540 gnd.n2539 585
R3372 gnd.n2539 gnd.n1177 585
R3373 gnd.n2538 gnd.n1175 585
R3374 gnd.n5022 gnd.n1175 585
R3375 gnd.n2537 gnd.n2536 585
R3376 gnd.n2536 gnd.n1167 585
R3377 gnd.n2534 gnd.n1165 585
R3378 gnd.n5028 gnd.n1165 585
R3379 gnd.n2533 gnd.n2532 585
R3380 gnd.n2532 gnd.n1155 585
R3381 gnd.n2531 gnd.n1153 585
R3382 gnd.n5034 gnd.n1153 585
R3383 gnd.n2530 gnd.n1141 585
R3384 gnd.n1152 gnd.n1141 585
R3385 gnd.n5041 gnd.n1139 585
R3386 gnd.n5041 gnd.n5040 585
R3387 gnd.n5043 gnd.n5042 585
R3388 gnd.n5042 gnd.n1068 585
R3389 gnd.n7674 gnd.n7673 585
R3390 gnd.n7675 gnd.n7674 585
R3391 gnd.n201 gnd.n200 585
R3392 gnd.n209 gnd.n201 585
R3393 gnd.n7683 gnd.n7682 585
R3394 gnd.n7682 gnd.n7681 585
R3395 gnd.n7684 gnd.n195 585
R3396 gnd.n195 gnd.n194 585
R3397 gnd.n7686 gnd.n7685 585
R3398 gnd.n7687 gnd.n7686 585
R3399 gnd.n182 gnd.n181 585
R3400 gnd.n185 gnd.n182 585
R3401 gnd.n7695 gnd.n7694 585
R3402 gnd.n7694 gnd.n7693 585
R3403 gnd.n7696 gnd.n176 585
R3404 gnd.n176 gnd.n175 585
R3405 gnd.n7698 gnd.n7697 585
R3406 gnd.n7699 gnd.n7698 585
R3407 gnd.n162 gnd.n161 585
R3408 gnd.n7510 gnd.n162 585
R3409 gnd.n7707 gnd.n7706 585
R3410 gnd.n7706 gnd.n7705 585
R3411 gnd.n7708 gnd.n156 585
R3412 gnd.n7489 gnd.n156 585
R3413 gnd.n7710 gnd.n7709 585
R3414 gnd.n7711 gnd.n7710 585
R3415 gnd.n142 gnd.n141 585
R3416 gnd.n7480 gnd.n142 585
R3417 gnd.n7719 gnd.n7718 585
R3418 gnd.n7718 gnd.n7717 585
R3419 gnd.n7720 gnd.n136 585
R3420 gnd.n7474 gnd.n136 585
R3421 gnd.n7722 gnd.n7721 585
R3422 gnd.n7723 gnd.n7722 585
R3423 gnd.n122 gnd.n121 585
R3424 gnd.n7466 gnd.n122 585
R3425 gnd.n7731 gnd.n7730 585
R3426 gnd.n7730 gnd.n7729 585
R3427 gnd.n7732 gnd.n117 585
R3428 gnd.n7460 gnd.n117 585
R3429 gnd.n7734 gnd.n7733 585
R3430 gnd.n7735 gnd.n7734 585
R3431 gnd.n101 gnd.n99 585
R3432 gnd.n7452 gnd.n101 585
R3433 gnd.n7743 gnd.n7742 585
R3434 gnd.n7742 gnd.n7741 585
R3435 gnd.n100 gnd.n92 585
R3436 gnd.n7446 gnd.n100 585
R3437 gnd.n7746 gnd.n90 585
R3438 gnd.n381 gnd.n90 585
R3439 gnd.n7748 gnd.n7747 585
R3440 gnd.n7749 gnd.n7748 585
R3441 gnd.n1744 gnd.n89 585
R3442 gnd.n4536 gnd.n89 585
R3443 gnd.n1746 gnd.n1745 585
R3444 gnd.n1751 gnd.n1746 585
R3445 gnd.n4573 gnd.n1747 585
R3446 gnd.n4573 gnd.n4572 585
R3447 gnd.n4574 gnd.n97 585
R3448 gnd.n4575 gnd.n4574 585
R3449 gnd.n1730 gnd.n1729 585
R3450 gnd.n4557 gnd.n1730 585
R3451 gnd.n4583 gnd.n4582 585
R3452 gnd.n4582 gnd.n4581 585
R3453 gnd.n4584 gnd.n1726 585
R3454 gnd.n4546 gnd.n1726 585
R3455 gnd.n4586 gnd.n4585 585
R3456 gnd.n4587 gnd.n4586 585
R3457 gnd.n1712 gnd.n1711 585
R3458 gnd.n4516 gnd.n1712 585
R3459 gnd.n4595 gnd.n4594 585
R3460 gnd.n4594 gnd.n4593 585
R3461 gnd.n4596 gnd.n1706 585
R3462 gnd.n4475 gnd.n1706 585
R3463 gnd.n4598 gnd.n4597 585
R3464 gnd.n4599 gnd.n4598 585
R3465 gnd.n1692 gnd.n1691 585
R3466 gnd.n4468 gnd.n1692 585
R3467 gnd.n4607 gnd.n4606 585
R3468 gnd.n4606 gnd.n4605 585
R3469 gnd.n4608 gnd.n1686 585
R3470 gnd.n4463 gnd.n1686 585
R3471 gnd.n4610 gnd.n4609 585
R3472 gnd.n4611 gnd.n4610 585
R3473 gnd.n1672 gnd.n1671 585
R3474 gnd.n4492 gnd.n1672 585
R3475 gnd.n4619 gnd.n4618 585
R3476 gnd.n4618 gnd.n4617 585
R3477 gnd.n4620 gnd.n1666 585
R3478 gnd.n4456 gnd.n1666 585
R3479 gnd.n4622 gnd.n4621 585
R3480 gnd.n4623 gnd.n4622 585
R3481 gnd.n1652 gnd.n1651 585
R3482 gnd.n4448 gnd.n1652 585
R3483 gnd.n4631 gnd.n4630 585
R3484 gnd.n4630 gnd.n4629 585
R3485 gnd.n4632 gnd.n1646 585
R3486 gnd.n4442 gnd.n1646 585
R3487 gnd.n4634 gnd.n4633 585
R3488 gnd.n4635 gnd.n4634 585
R3489 gnd.n1629 gnd.n1628 585
R3490 gnd.n4434 gnd.n1629 585
R3491 gnd.n4643 gnd.n4642 585
R3492 gnd.n4642 gnd.n4641 585
R3493 gnd.n4644 gnd.n1624 585
R3494 gnd.n3886 gnd.n1624 585
R3495 gnd.n4646 gnd.n4645 585
R3496 gnd.n4647 gnd.n4646 585
R3497 gnd.n4275 gnd.n1623 585
R3498 gnd.n4280 gnd.n4278 585
R3499 gnd.n4281 gnd.n4274 585
R3500 gnd.n4281 gnd.n1610 585
R3501 gnd.n4284 gnd.n4283 585
R3502 gnd.n4272 gnd.n4271 585
R3503 gnd.n4289 gnd.n4288 585
R3504 gnd.n4291 gnd.n4270 585
R3505 gnd.n4294 gnd.n4293 585
R3506 gnd.n4268 gnd.n4267 585
R3507 gnd.n4299 gnd.n4298 585
R3508 gnd.n4301 gnd.n4266 585
R3509 gnd.n4304 gnd.n4303 585
R3510 gnd.n4264 gnd.n4263 585
R3511 gnd.n4309 gnd.n4308 585
R3512 gnd.n4311 gnd.n4262 585
R3513 gnd.n4314 gnd.n4313 585
R3514 gnd.n4260 gnd.n4259 585
R3515 gnd.n4322 gnd.n4321 585
R3516 gnd.n4324 gnd.n4258 585
R3517 gnd.n4327 gnd.n4326 585
R3518 gnd.n4256 gnd.n4255 585
R3519 gnd.n4332 gnd.n4331 585
R3520 gnd.n4334 gnd.n4254 585
R3521 gnd.n4337 gnd.n4336 585
R3522 gnd.n4252 gnd.n4251 585
R3523 gnd.n4343 gnd.n4342 585
R3524 gnd.n4347 gnd.n1860 585
R3525 gnd.n4350 gnd.n4349 585
R3526 gnd.n1858 gnd.n1857 585
R3527 gnd.n4355 gnd.n4354 585
R3528 gnd.n4357 gnd.n1856 585
R3529 gnd.n4360 gnd.n4359 585
R3530 gnd.n1854 gnd.n1853 585
R3531 gnd.n4365 gnd.n4364 585
R3532 gnd.n4367 gnd.n1852 585
R3533 gnd.n4372 gnd.n4369 585
R3534 gnd.n1850 gnd.n1849 585
R3535 gnd.n4377 gnd.n4376 585
R3536 gnd.n4379 gnd.n1848 585
R3537 gnd.n4382 gnd.n4381 585
R3538 gnd.n1846 gnd.n1845 585
R3539 gnd.n4387 gnd.n4386 585
R3540 gnd.n4389 gnd.n1844 585
R3541 gnd.n4392 gnd.n4391 585
R3542 gnd.n1842 gnd.n1841 585
R3543 gnd.n4397 gnd.n4396 585
R3544 gnd.n4399 gnd.n1840 585
R3545 gnd.n4402 gnd.n4401 585
R3546 gnd.n1838 gnd.n1837 585
R3547 gnd.n4407 gnd.n4406 585
R3548 gnd.n4409 gnd.n1836 585
R3549 gnd.n4412 gnd.n4411 585
R3550 gnd.n1834 gnd.n1833 585
R3551 gnd.n4418 gnd.n4417 585
R3552 gnd.n4420 gnd.n1832 585
R3553 gnd.n4421 gnd.n1831 585
R3554 gnd.n4424 gnd.n4423 585
R3555 gnd.n7565 gnd.n7564 585
R3556 gnd.n7567 gnd.n315 585
R3557 gnd.n7569 gnd.n7568 585
R3558 gnd.n7570 gnd.n308 585
R3559 gnd.n7572 gnd.n7571 585
R3560 gnd.n7574 gnd.n306 585
R3561 gnd.n7576 gnd.n7575 585
R3562 gnd.n7577 gnd.n301 585
R3563 gnd.n7579 gnd.n7578 585
R3564 gnd.n7581 gnd.n299 585
R3565 gnd.n7583 gnd.n7582 585
R3566 gnd.n7584 gnd.n294 585
R3567 gnd.n7586 gnd.n7585 585
R3568 gnd.n7588 gnd.n292 585
R3569 gnd.n7590 gnd.n7589 585
R3570 gnd.n7591 gnd.n287 585
R3571 gnd.n7593 gnd.n7592 585
R3572 gnd.n7595 gnd.n286 585
R3573 gnd.n7596 gnd.n283 585
R3574 gnd.n7599 gnd.n7598 585
R3575 gnd.n285 gnd.n279 585
R3576 gnd.n7603 gnd.n276 585
R3577 gnd.n7605 gnd.n7604 585
R3578 gnd.n7607 gnd.n274 585
R3579 gnd.n7609 gnd.n7608 585
R3580 gnd.n7610 gnd.n269 585
R3581 gnd.n7612 gnd.n7611 585
R3582 gnd.n7614 gnd.n267 585
R3583 gnd.n7616 gnd.n7615 585
R3584 gnd.n7617 gnd.n262 585
R3585 gnd.n7619 gnd.n7618 585
R3586 gnd.n7621 gnd.n260 585
R3587 gnd.n7623 gnd.n7622 585
R3588 gnd.n7624 gnd.n255 585
R3589 gnd.n7626 gnd.n7625 585
R3590 gnd.n7628 gnd.n253 585
R3591 gnd.n7630 gnd.n7629 585
R3592 gnd.n7631 gnd.n248 585
R3593 gnd.n7633 gnd.n7632 585
R3594 gnd.n7635 gnd.n246 585
R3595 gnd.n7637 gnd.n7636 585
R3596 gnd.n7641 gnd.n241 585
R3597 gnd.n7643 gnd.n7642 585
R3598 gnd.n7645 gnd.n239 585
R3599 gnd.n7647 gnd.n7646 585
R3600 gnd.n7648 gnd.n234 585
R3601 gnd.n7650 gnd.n7649 585
R3602 gnd.n7652 gnd.n232 585
R3603 gnd.n7654 gnd.n7653 585
R3604 gnd.n7655 gnd.n227 585
R3605 gnd.n7657 gnd.n7656 585
R3606 gnd.n7659 gnd.n225 585
R3607 gnd.n7661 gnd.n7660 585
R3608 gnd.n7662 gnd.n220 585
R3609 gnd.n7664 gnd.n7663 585
R3610 gnd.n7666 gnd.n218 585
R3611 gnd.n7668 gnd.n7667 585
R3612 gnd.n7669 gnd.n216 585
R3613 gnd.n7670 gnd.n213 585
R3614 gnd.n213 gnd.n212 585
R3615 gnd.n7495 gnd.n210 585
R3616 gnd.n7675 gnd.n210 585
R3617 gnd.n7497 gnd.n7496 585
R3618 gnd.n7496 gnd.n209 585
R3619 gnd.n7498 gnd.n202 585
R3620 gnd.n7681 gnd.n202 585
R3621 gnd.n7500 gnd.n7499 585
R3622 gnd.n7499 gnd.n194 585
R3623 gnd.n7501 gnd.n192 585
R3624 gnd.n7687 gnd.n192 585
R3625 gnd.n7503 gnd.n7502 585
R3626 gnd.n7502 gnd.n185 585
R3627 gnd.n7504 gnd.n183 585
R3628 gnd.n7693 gnd.n183 585
R3629 gnd.n7506 gnd.n7505 585
R3630 gnd.n7505 gnd.n175 585
R3631 gnd.n7507 gnd.n173 585
R3632 gnd.n7699 gnd.n173 585
R3633 gnd.n7509 gnd.n7508 585
R3634 gnd.n7510 gnd.n7509 585
R3635 gnd.n7492 gnd.n164 585
R3636 gnd.n7705 gnd.n164 585
R3637 gnd.n7491 gnd.n7490 585
R3638 gnd.n7490 gnd.n7489 585
R3639 gnd.n360 gnd.n154 585
R3640 gnd.n7711 gnd.n154 585
R3641 gnd.n7479 gnd.n7478 585
R3642 gnd.n7480 gnd.n7479 585
R3643 gnd.n7477 gnd.n144 585
R3644 gnd.n7717 gnd.n144 585
R3645 gnd.n7476 gnd.n7475 585
R3646 gnd.n7475 gnd.n7474 585
R3647 gnd.n366 gnd.n133 585
R3648 gnd.n7723 gnd.n133 585
R3649 gnd.n7465 gnd.n7464 585
R3650 gnd.n7466 gnd.n7465 585
R3651 gnd.n7463 gnd.n124 585
R3652 gnd.n7729 gnd.n124 585
R3653 gnd.n7462 gnd.n7461 585
R3654 gnd.n7461 gnd.n7460 585
R3655 gnd.n372 gnd.n115 585
R3656 gnd.n7735 gnd.n115 585
R3657 gnd.n7451 gnd.n7450 585
R3658 gnd.n7452 gnd.n7451 585
R3659 gnd.n7449 gnd.n103 585
R3660 gnd.n7741 gnd.n103 585
R3661 gnd.n7448 gnd.n7447 585
R3662 gnd.n7447 gnd.n7446 585
R3663 gnd.n380 gnd.n378 585
R3664 gnd.n381 gnd.n380 585
R3665 gnd.n4528 gnd.n86 585
R3666 gnd.n7749 gnd.n86 585
R3667 gnd.n4537 gnd.n4523 585
R3668 gnd.n4537 gnd.n4536 585
R3669 gnd.n4539 gnd.n4538 585
R3670 gnd.n4538 gnd.n1751 585
R3671 gnd.n4540 gnd.n1748 585
R3672 gnd.n4572 gnd.n1748 585
R3673 gnd.n4541 gnd.n1741 585
R3674 gnd.n4575 gnd.n1741 585
R3675 gnd.n4542 gnd.n1756 585
R3676 gnd.n4557 gnd.n1756 585
R3677 gnd.n4543 gnd.n1732 585
R3678 gnd.n4581 gnd.n1732 585
R3679 gnd.n4545 gnd.n4544 585
R3680 gnd.n4546 gnd.n4545 585
R3681 gnd.n4519 gnd.n1723 585
R3682 gnd.n4587 gnd.n1723 585
R3683 gnd.n4518 gnd.n4517 585
R3684 gnd.n4517 gnd.n4516 585
R3685 gnd.n1761 gnd.n1714 585
R3686 gnd.n4593 gnd.n1714 585
R3687 gnd.n4474 gnd.n4473 585
R3688 gnd.n4475 gnd.n4474 585
R3689 gnd.n4471 gnd.n1703 585
R3690 gnd.n4599 gnd.n1703 585
R3691 gnd.n4470 gnd.n4469 585
R3692 gnd.n4469 gnd.n4468 585
R3693 gnd.n4466 gnd.n1694 585
R3694 gnd.n4605 gnd.n1694 585
R3695 gnd.n4465 gnd.n4464 585
R3696 gnd.n4464 gnd.n4463 585
R3697 gnd.n4461 gnd.n1683 585
R3698 gnd.n4611 gnd.n1683 585
R3699 gnd.n4460 gnd.n1774 585
R3700 gnd.n4492 gnd.n1774 585
R3701 gnd.n4459 gnd.n1674 585
R3702 gnd.n4617 gnd.n1674 585
R3703 gnd.n4458 gnd.n4457 585
R3704 gnd.n4457 gnd.n4456 585
R3705 gnd.n1783 gnd.n1663 585
R3706 gnd.n4623 gnd.n1663 585
R3707 gnd.n4447 gnd.n4446 585
R3708 gnd.n4448 gnd.n4447 585
R3709 gnd.n4445 gnd.n1654 585
R3710 gnd.n4629 gnd.n1654 585
R3711 gnd.n4444 gnd.n4443 585
R3712 gnd.n4443 gnd.n4442 585
R3713 gnd.n1820 gnd.n1643 585
R3714 gnd.n4635 gnd.n1643 585
R3715 gnd.n4433 gnd.n4432 585
R3716 gnd.n4434 gnd.n4433 585
R3717 gnd.n4431 gnd.n1631 585
R3718 gnd.n4641 gnd.n1631 585
R3719 gnd.n4430 gnd.n1826 585
R3720 gnd.n3886 gnd.n1826 585
R3721 gnd.n1825 gnd.n1619 585
R3722 gnd.n4647 gnd.n1619 585
R3723 gnd.n2650 gnd.n2648 585
R3724 gnd.n2648 gnd.n1184 585
R3725 gnd.n7416 gnd.n7415 585
R3726 gnd.n7415 gnd.n172 585
R3727 gnd.n7419 gnd.n399 585
R3728 gnd.n399 gnd.n163 585
R3729 gnd.n7421 gnd.n7420 585
R3730 gnd.n7421 gnd.n362 585
R3731 gnd.n7422 gnd.n398 585
R3732 gnd.n7422 gnd.n153 585
R3733 gnd.n7424 gnd.n7423 585
R3734 gnd.n7423 gnd.n146 585
R3735 gnd.n7425 gnd.n393 585
R3736 gnd.n393 gnd.n143 585
R3737 gnd.n7427 gnd.n7426 585
R3738 gnd.n7427 gnd.n135 585
R3739 gnd.n7428 gnd.n392 585
R3740 gnd.n7428 gnd.n132 585
R3741 gnd.n7430 gnd.n7429 585
R3742 gnd.n7429 gnd.n371 585
R3743 gnd.n7431 gnd.n387 585
R3744 gnd.n387 gnd.n123 585
R3745 gnd.n7433 gnd.n7432 585
R3746 gnd.n7433 gnd.n374 585
R3747 gnd.n7434 gnd.n386 585
R3748 gnd.n7434 gnd.n114 585
R3749 gnd.n7436 gnd.n7435 585
R3750 gnd.n7435 gnd.n105 585
R3751 gnd.n7437 gnd.n383 585
R3752 gnd.n383 gnd.n102 585
R3753 gnd.n7440 gnd.n7439 585
R3754 gnd.n7441 gnd.n7440 585
R3755 gnd.n384 gnd.n382 585
R3756 gnd.n382 gnd.n87 585
R3757 gnd.n4566 gnd.n4565 585
R3758 gnd.n4565 gnd.n85 585
R3759 gnd.n4567 gnd.n1753 585
R3760 gnd.n4524 gnd.n1753 585
R3761 gnd.n4570 gnd.n4569 585
R3762 gnd.n4571 gnd.n4570 585
R3763 gnd.n4563 gnd.n1752 585
R3764 gnd.n1752 gnd.n1743 585
R3765 gnd.n4561 gnd.n4560 585
R3766 gnd.n4560 gnd.n1740 585
R3767 gnd.n4559 gnd.n1754 585
R3768 gnd.n4559 gnd.n4558 585
R3769 gnd.n4511 gnd.n1755 585
R3770 gnd.n1755 gnd.n1731 585
R3771 gnd.n4512 gnd.n1764 585
R3772 gnd.n1764 gnd.n1725 585
R3773 gnd.n4514 gnd.n4513 585
R3774 gnd.n4515 gnd.n4514 585
R3775 gnd.n1765 gnd.n1763 585
R3776 gnd.n1763 gnd.n1716 585
R3777 gnd.n4505 gnd.n4504 585
R3778 gnd.n4504 gnd.n1713 585
R3779 gnd.n4503 gnd.n1767 585
R3780 gnd.n4503 gnd.n1705 585
R3781 gnd.n4502 gnd.n4501 585
R3782 gnd.n4502 gnd.n1702 585
R3783 gnd.n1769 gnd.n1768 585
R3784 gnd.n4467 gnd.n1768 585
R3785 gnd.n4497 gnd.n4496 585
R3786 gnd.n4496 gnd.n1693 585
R3787 gnd.n4495 gnd.n1771 585
R3788 gnd.n4495 gnd.n1685 585
R3789 gnd.n4494 gnd.n1773 585
R3790 gnd.n4494 gnd.n4493 585
R3791 gnd.n1811 gnd.n1772 585
R3792 gnd.n1772 gnd.n1676 585
R3793 gnd.n1813 gnd.n1812 585
R3794 gnd.n1813 gnd.n1673 585
R3795 gnd.n1815 gnd.n1814 585
R3796 gnd.n1814 gnd.n1665 585
R3797 gnd.n1816 gnd.n1789 585
R3798 gnd.n1789 gnd.n1662 585
R3799 gnd.n1818 gnd.n1817 585
R3800 gnd.n1819 gnd.n1818 585
R3801 gnd.n1790 gnd.n1788 585
R3802 gnd.n1788 gnd.n1653 585
R3803 gnd.n1802 gnd.n1801 585
R3804 gnd.n1801 gnd.n1645 585
R3805 gnd.n1800 gnd.n1792 585
R3806 gnd.n1800 gnd.n1642 585
R3807 gnd.n1799 gnd.n1798 585
R3808 gnd.n1799 gnd.n1633 585
R3809 gnd.n1794 gnd.n1793 585
R3810 gnd.n1793 gnd.n1630 585
R3811 gnd.n1617 gnd.n1616 585
R3812 gnd.n1621 gnd.n1617 585
R3813 gnd.n4650 gnd.n4649 585
R3814 gnd.n4649 gnd.n4648 585
R3815 gnd.n4651 gnd.n1611 585
R3816 gnd.n1618 gnd.n1611 585
R3817 gnd.n4653 gnd.n4652 585
R3818 gnd.n4654 gnd.n4653 585
R3819 gnd.n1608 gnd.n1607 585
R3820 gnd.n4655 gnd.n1608 585
R3821 gnd.n4658 gnd.n4657 585
R3822 gnd.n4657 gnd.n4656 585
R3823 gnd.n4659 gnd.n1602 585
R3824 gnd.n1602 gnd.n1600 585
R3825 gnd.n4661 gnd.n4660 585
R3826 gnd.n4662 gnd.n4661 585
R3827 gnd.n1603 gnd.n1601 585
R3828 gnd.n1601 gnd.n1598 585
R3829 gnd.n1933 gnd.n1932 585
R3830 gnd.n4067 gnd.n1933 585
R3831 gnd.n4071 gnd.n4070 585
R3832 gnd.n4070 gnd.n4069 585
R3833 gnd.n4072 gnd.n1923 585
R3834 gnd.n1934 gnd.n1923 585
R3835 gnd.n4074 gnd.n4073 585
R3836 gnd.n4075 gnd.n4074 585
R3837 gnd.n1924 gnd.n1918 585
R3838 gnd.n4078 gnd.n1918 585
R3839 gnd.n4081 gnd.n1917 585
R3840 gnd.n4081 gnd.n4080 585
R3841 gnd.n4083 gnd.n4082 585
R3842 gnd.n4082 gnd.n1865 585
R3843 gnd.n4084 gnd.n1912 585
R3844 gnd.n1912 gnd.n1902 585
R3845 gnd.n4086 gnd.n4085 585
R3846 gnd.n4087 gnd.n4086 585
R3847 gnd.n1913 gnd.n1911 585
R3848 gnd.n1911 gnd.n1907 585
R3849 gnd.n3838 gnd.n1961 585
R3850 gnd.n1961 gnd.n1960 585
R3851 gnd.n3840 gnd.n3839 585
R3852 gnd.n3841 gnd.n3840 585
R3853 gnd.n1962 gnd.n1959 585
R3854 gnd.n1959 gnd.n1956 585
R3855 gnd.n3832 gnd.n3831 585
R3856 gnd.n3831 gnd.n3830 585
R3857 gnd.n1965 gnd.n1964 585
R3858 gnd.n3818 gnd.n1965 585
R3859 gnd.n3793 gnd.n1991 585
R3860 gnd.n1991 gnd.n1983 585
R3861 gnd.n3795 gnd.n3794 585
R3862 gnd.n3796 gnd.n3795 585
R3863 gnd.n1992 gnd.n1990 585
R3864 gnd.n3783 gnd.n1990 585
R3865 gnd.n3788 gnd.n3787 585
R3866 gnd.n3787 gnd.n3786 585
R3867 gnd.n1995 gnd.n1994 585
R3868 gnd.n2007 gnd.n1995 585
R3869 gnd.n3767 gnd.n3766 585
R3870 gnd.n3768 gnd.n3767 585
R3871 gnd.n2012 gnd.n2011 585
R3872 gnd.n2019 gnd.n2011 585
R3873 gnd.n3762 gnd.n3761 585
R3874 gnd.n3761 gnd.n3760 585
R3875 gnd.n2015 gnd.n2014 585
R3876 gnd.n3657 gnd.n2015 585
R3877 gnd.n3716 gnd.n2039 585
R3878 gnd.n2039 gnd.n2032 585
R3879 gnd.n3718 gnd.n3717 585
R3880 gnd.n3719 gnd.n3718 585
R3881 gnd.n2040 gnd.n2038 585
R3882 gnd.n2038 gnd.n2036 585
R3883 gnd.n3711 gnd.n3710 585
R3884 gnd.n3710 gnd.n3709 585
R3885 gnd.n2043 gnd.n2042 585
R3886 gnd.n3701 gnd.n2043 585
R3887 gnd.n3687 gnd.n3686 585
R3888 gnd.n3688 gnd.n3687 585
R3889 gnd.n2062 gnd.n2061 585
R3890 gnd.n3637 gnd.n2061 585
R3891 gnd.n3682 gnd.n3681 585
R3892 gnd.n3681 gnd.n3680 585
R3893 gnd.n2065 gnd.n2064 585
R3894 gnd.n2073 gnd.n2065 585
R3895 gnd.n3627 gnd.n3626 585
R3896 gnd.n3628 gnd.n3627 585
R3897 gnd.n2082 gnd.n2081 585
R3898 gnd.n2081 gnd.n2078 585
R3899 gnd.n3622 gnd.n3621 585
R3900 gnd.n3621 gnd.n3620 585
R3901 gnd.n2085 gnd.n2084 585
R3902 gnd.n2091 gnd.n2085 585
R3903 gnd.n3602 gnd.n3601 585
R3904 gnd.n3603 gnd.n3602 585
R3905 gnd.n2102 gnd.n2101 585
R3906 gnd.n2109 gnd.n2101 585
R3907 gnd.n3597 gnd.n3596 585
R3908 gnd.n3596 gnd.n3595 585
R3909 gnd.n2105 gnd.n2104 585
R3910 gnd.n2113 gnd.n2105 585
R3911 gnd.n3545 gnd.n3544 585
R3912 gnd.n3546 gnd.n3545 585
R3913 gnd.n2124 gnd.n2123 585
R3914 gnd.n2142 gnd.n2123 585
R3915 gnd.n3540 gnd.n3539 585
R3916 gnd.n3539 gnd.n3538 585
R3917 gnd.n2127 gnd.n2126 585
R3918 gnd.n2135 gnd.n2127 585
R3919 gnd.n3505 gnd.n3504 585
R3920 gnd.n3506 gnd.n3505 585
R3921 gnd.n2147 gnd.n2146 585
R3922 gnd.n2162 gnd.n2146 585
R3923 gnd.n3500 gnd.n3499 585
R3924 gnd.n3499 gnd.n3498 585
R3925 gnd.n2150 gnd.n2149 585
R3926 gnd.n3488 gnd.n2150 585
R3927 gnd.n3455 gnd.n2179 585
R3928 gnd.n2179 gnd.n2171 585
R3929 gnd.n3457 gnd.n3456 585
R3930 gnd.n3458 gnd.n3457 585
R3931 gnd.n2180 gnd.n2178 585
R3932 gnd.n2178 gnd.n2175 585
R3933 gnd.n3450 gnd.n3449 585
R3934 gnd.n3449 gnd.n3448 585
R3935 gnd.n2183 gnd.n2182 585
R3936 gnd.n2189 gnd.n2183 585
R3937 gnd.n3427 gnd.n3426 585
R3938 gnd.n3428 gnd.n3427 585
R3939 gnd.n2198 gnd.n2197 585
R3940 gnd.n2204 gnd.n2197 585
R3941 gnd.n3422 gnd.n3421 585
R3942 gnd.n3421 gnd.n3420 585
R3943 gnd.n2201 gnd.n2200 585
R3944 gnd.n2208 gnd.n2201 585
R3945 gnd.n3365 gnd.n2223 585
R3946 gnd.n2223 gnd.n2213 585
R3947 gnd.n3367 gnd.n3366 585
R3948 gnd.n3368 gnd.n3367 585
R3949 gnd.n2224 gnd.n2222 585
R3950 gnd.n3333 gnd.n2222 585
R3951 gnd.n3360 gnd.n3359 585
R3952 gnd.n3359 gnd.n3358 585
R3953 gnd.n2227 gnd.n2226 585
R3954 gnd.n3341 gnd.n2227 585
R3955 gnd.n3323 gnd.n3322 585
R3956 gnd.n3324 gnd.n3323 585
R3957 gnd.n2242 gnd.n2241 585
R3958 gnd.n3301 gnd.n2241 585
R3959 gnd.n3318 gnd.n3317 585
R3960 gnd.n3317 gnd.n3316 585
R3961 gnd.n2245 gnd.n2244 585
R3962 gnd.n2252 gnd.n2245 585
R3963 gnd.n3280 gnd.n3279 585
R3964 gnd.n3281 gnd.n3280 585
R3965 gnd.n1501 gnd.n1500 585
R3966 gnd.n2266 gnd.n1501 585
R3967 gnd.n4776 gnd.n4775 585
R3968 gnd.n4775 gnd.n4774 585
R3969 gnd.n4777 gnd.n1495 585
R3970 gnd.n2270 gnd.n1495 585
R3971 gnd.n4779 gnd.n4778 585
R3972 gnd.n4780 gnd.n4779 585
R3973 gnd.n1496 gnd.n1494 585
R3974 gnd.n2356 gnd.n1494 585
R3975 gnd.n3242 gnd.n2367 585
R3976 gnd.n2367 gnd.n1465 585
R3977 gnd.n3244 gnd.n3243 585
R3978 gnd.n3245 gnd.n3244 585
R3979 gnd.n2368 gnd.n2366 585
R3980 gnd.n2366 gnd.n2364 585
R3981 gnd.n3236 gnd.n3235 585
R3982 gnd.n3235 gnd.n3234 585
R3983 gnd.n2371 gnd.n2370 585
R3984 gnd.n2380 gnd.n2371 585
R3985 gnd.n3209 gnd.n2392 585
R3986 gnd.n2392 gnd.n2379 585
R3987 gnd.n3211 gnd.n3210 585
R3988 gnd.n3212 gnd.n3211 585
R3989 gnd.n2393 gnd.n2391 585
R3990 gnd.n2391 gnd.n2388 585
R3991 gnd.n3204 gnd.n3203 585
R3992 gnd.n3203 gnd.n3202 585
R3993 gnd.n2396 gnd.n2395 585
R3994 gnd.n2397 gnd.n2396 585
R3995 gnd.n2925 gnd.n2924 585
R3996 gnd.n2926 gnd.n2925 585
R3997 gnd.n2418 gnd.n2417 585
R3998 gnd.n2417 gnd.n2416 585
R3999 gnd.n2920 gnd.n2919 585
R4000 gnd.n2919 gnd.n2918 585
R4001 gnd.n2917 gnd.n2420 585
R4002 gnd.n2917 gnd.n2916 585
R4003 gnd.n2915 gnd.n2914 585
R4004 gnd.n2915 gnd.n1376 585
R4005 gnd.n2422 gnd.n2421 585
R4006 gnd.n2421 gnd.n1373 585
R4007 gnd.n2910 gnd.n2909 585
R4008 gnd.n2909 gnd.n1367 585
R4009 gnd.n2908 gnd.n2424 585
R4010 gnd.n2908 gnd.n1364 585
R4011 gnd.n2907 gnd.n2906 585
R4012 gnd.n2907 gnd.n1356 585
R4013 gnd.n2426 gnd.n2425 585
R4014 gnd.n2425 gnd.n1353 585
R4015 gnd.n2902 gnd.n2901 585
R4016 gnd.n2901 gnd.n1346 585
R4017 gnd.n2900 gnd.n2428 585
R4018 gnd.n2900 gnd.n2899 585
R4019 gnd.n2828 gnd.n2429 585
R4020 gnd.n2429 gnd.n1336 585
R4021 gnd.n2830 gnd.n2829 585
R4022 gnd.n2829 gnd.n1333 585
R4023 gnd.n2831 gnd.n2822 585
R4024 gnd.n2822 gnd.n1326 585
R4025 gnd.n2833 gnd.n2832 585
R4026 gnd.n2833 gnd.n1323 585
R4027 gnd.n2834 gnd.n2821 585
R4028 gnd.n2834 gnd.n2443 585
R4029 gnd.n2836 gnd.n2835 585
R4030 gnd.n2835 gnd.n1313 585
R4031 gnd.n2837 gnd.n2450 585
R4032 gnd.n2450 gnd.n1306 585
R4033 gnd.n2839 gnd.n2838 585
R4034 gnd.n2840 gnd.n2839 585
R4035 gnd.n2451 gnd.n2449 585
R4036 gnd.n2449 gnd.n1296 585
R4037 gnd.n2815 gnd.n2814 585
R4038 gnd.n2814 gnd.n1293 585
R4039 gnd.n2813 gnd.n2453 585
R4040 gnd.n2813 gnd.n1286 585
R4041 gnd.n2812 gnd.n2811 585
R4042 gnd.n2812 gnd.n1283 585
R4043 gnd.n2455 gnd.n2454 585
R4044 gnd.n2778 gnd.n2454 585
R4045 gnd.n2807 gnd.n2806 585
R4046 gnd.n2806 gnd.n1274 585
R4047 gnd.n2805 gnd.n2456 585
R4048 gnd.n2805 gnd.n1265 585
R4049 gnd.n2804 gnd.n2459 585
R4050 gnd.n2804 gnd.n2803 585
R4051 gnd.n2735 gnd.n2457 585
R4052 gnd.n2460 gnd.n2457 585
R4053 gnd.n2737 gnd.n2498 585
R4054 gnd.n2498 gnd.n2474 585
R4055 gnd.n2739 gnd.n2738 585
R4056 gnd.n2740 gnd.n2739 585
R4057 gnd.n2733 gnd.n2497 585
R4058 gnd.n2497 gnd.n2484 585
R4059 gnd.n2732 gnd.n2731 585
R4060 gnd.n2731 gnd.n2490 585
R4061 gnd.n2730 gnd.n2729 585
R4062 gnd.n2730 gnd.n2488 585
R4063 gnd.n2728 gnd.n2500 585
R4064 gnd.n2506 gnd.n2500 585
R4065 gnd.n2726 gnd.n2725 585
R4066 gnd.n2725 gnd.n2724 585
R4067 gnd.n2502 gnd.n2501 585
R4068 gnd.n2502 gnd.n1248 585
R4069 gnd.n2671 gnd.n2670 585
R4070 gnd.n2670 gnd.n1245 585
R4071 gnd.n2672 gnd.n2664 585
R4072 gnd.n2664 gnd.n1238 585
R4073 gnd.n2674 gnd.n2673 585
R4074 gnd.n2674 gnd.n1235 585
R4075 gnd.n2675 gnd.n2663 585
R4076 gnd.n2675 gnd.n1227 585
R4077 gnd.n2677 gnd.n2676 585
R4078 gnd.n2676 gnd.n1224 585
R4079 gnd.n2678 gnd.n2644 585
R4080 gnd.n2644 gnd.n1217 585
R4081 gnd.n2680 gnd.n2679 585
R4082 gnd.n2681 gnd.n2680 585
R4083 gnd.n2645 gnd.n2643 585
R4084 gnd.n2643 gnd.n1207 585
R4085 gnd.n2657 gnd.n2656 585
R4086 gnd.n2656 gnd.n1204 585
R4087 gnd.n2655 gnd.n2647 585
R4088 gnd.n2655 gnd.n1197 585
R4089 gnd.n2654 gnd.n2653 585
R4090 gnd.n2654 gnd.n1194 585
R4091 gnd.n4665 gnd.n4664 585
R4092 gnd.n4664 gnd.n4663 585
R4093 gnd.n1596 gnd.n1594 585
R4094 gnd.n4066 gnd.n1596 585
R4095 gnd.n4669 gnd.n1593 585
R4096 gnd.n4068 gnd.n1593 585
R4097 gnd.n4670 gnd.n1592 585
R4098 gnd.n1935 gnd.n1592 585
R4099 gnd.n4671 gnd.n1591 585
R4100 gnd.n1922 gnd.n1591 585
R4101 gnd.n4076 gnd.n1589 585
R4102 gnd.n4077 gnd.n4076 585
R4103 gnd.n4675 gnd.n1588 585
R4104 gnd.n4079 gnd.n1588 585
R4105 gnd.n4676 gnd.n1587 585
R4106 gnd.n1919 gnd.n1587 585
R4107 gnd.n4677 gnd.n1586 585
R4108 gnd.n3871 gnd.n1586 585
R4109 gnd.n3868 gnd.n1584 585
R4110 gnd.n3869 gnd.n3868 585
R4111 gnd.n4681 gnd.n1583 585
R4112 gnd.n4088 gnd.n1583 585
R4113 gnd.n4682 gnd.n1582 585
R4114 gnd.n3861 gnd.n1582 585
R4115 gnd.n4683 gnd.n1581 585
R4116 gnd.n1951 gnd.n1581 585
R4117 gnd.n3843 gnd.n1579 585
R4118 gnd.n3844 gnd.n3843 585
R4119 gnd.n4687 gnd.n1578 585
R4120 gnd.n3828 gnd.n1578 585
R4121 gnd.n4688 gnd.n1577 585
R4122 gnd.n1976 gnd.n1577 585
R4123 gnd.n4689 gnd.n1576 585
R4124 gnd.n3819 gnd.n1576 585
R4125 gnd.n1981 gnd.n1574 585
R4126 gnd.n1982 gnd.n1981 585
R4127 gnd.n4693 gnd.n1573 585
R4128 gnd.n3798 gnd.n1573 585
R4129 gnd.n4694 gnd.n1572 585
R4130 gnd.n3785 gnd.n1572 585
R4131 gnd.n4695 gnd.n1571 585
R4132 gnd.n3736 gnd.n1571 585
R4133 gnd.n2009 gnd.n1569 585
R4134 gnd.n2010 gnd.n2009 585
R4135 gnd.n4699 gnd.n1568 585
R4136 gnd.n2005 gnd.n1568 585
R4137 gnd.n4700 gnd.n1567 585
R4138 gnd.n3759 gnd.n1567 585
R4139 gnd.n4701 gnd.n1566 585
R4140 gnd.n3751 gnd.n1566 585
R4141 gnd.n3658 gnd.n1564 585
R4142 gnd.n3659 gnd.n3658 585
R4143 gnd.n4705 gnd.n1563 585
R4144 gnd.n3728 gnd.n1563 585
R4145 gnd.n4706 gnd.n1562 585
R4146 gnd.n3720 gnd.n1562 585
R4147 gnd.n4707 gnd.n1561 585
R4148 gnd.n2045 gnd.n1561 585
R4149 gnd.n3698 gnd.n1559 585
R4150 gnd.n3699 gnd.n3698 585
R4151 gnd.n4711 gnd.n1558 585
R4152 gnd.n2049 gnd.n1558 585
R4153 gnd.n4712 gnd.n1557 585
R4154 gnd.n3689 gnd.n1557 585
R4155 gnd.n4713 gnd.n1556 585
R4156 gnd.n2067 gnd.n1556 585
R4157 gnd.n3567 gnd.n1554 585
R4158 gnd.n3568 gnd.n3567 585
R4159 gnd.n4717 gnd.n1553 585
R4160 gnd.n2072 gnd.n1553 585
R4161 gnd.n4718 gnd.n1552 585
R4162 gnd.n3630 gnd.n1552 585
R4163 gnd.n4719 gnd.n1551 585
R4164 gnd.n3619 gnd.n1551 585
R4165 gnd.n2092 gnd.n1549 585
R4166 gnd.n2093 gnd.n2092 585
R4167 gnd.n4723 gnd.n1548 585
R4168 gnd.n2100 gnd.n1548 585
R4169 gnd.n4724 gnd.n1547 585
R4170 gnd.n3559 gnd.n1547 585
R4171 gnd.n4725 gnd.n1546 585
R4172 gnd.n3594 gnd.n1546 585
R4173 gnd.n3585 gnd.n1544 585
R4174 gnd.n3586 gnd.n3585 585
R4175 gnd.n4729 gnd.n1543 585
R4176 gnd.n3547 gnd.n1543 585
R4177 gnd.n4730 gnd.n1542 585
R4178 gnd.n3518 gnd.n1542 585
R4179 gnd.n4731 gnd.n1541 585
R4180 gnd.n2130 gnd.n1541 585
R4181 gnd.n3526 gnd.n1539 585
R4182 gnd.n3527 gnd.n3526 585
R4183 gnd.n4735 gnd.n1538 585
R4184 gnd.n3507 gnd.n1538 585
R4185 gnd.n4736 gnd.n1537 585
R4186 gnd.n3480 gnd.n1537 585
R4187 gnd.n4737 gnd.n1536 585
R4188 gnd.n2153 gnd.n1536 585
R4189 gnd.n3471 gnd.n1534 585
R4190 gnd.n3472 gnd.n3471 585
R4191 gnd.n4741 gnd.n1533 585
R4192 gnd.n2158 gnd.n1533 585
R4193 gnd.n4742 gnd.n1532 585
R4194 gnd.n3468 gnd.n1532 585
R4195 gnd.n4743 gnd.n1531 585
R4196 gnd.n3460 gnd.n1531 585
R4197 gnd.n3446 gnd.n1529 585
R4198 gnd.n3447 gnd.n3446 585
R4199 gnd.n4747 gnd.n1528 585
R4200 gnd.n2190 gnd.n1528 585
R4201 gnd.n4748 gnd.n1527 585
R4202 gnd.n3378 gnd.n1527 585
R4203 gnd.n4749 gnd.n1526 585
R4204 gnd.n2195 gnd.n1526 585
R4205 gnd.n3418 gnd.n1524 585
R4206 gnd.n3419 gnd.n3418 585
R4207 gnd.n4753 gnd.n1523 585
R4208 gnd.n3410 gnd.n1523 585
R4209 gnd.n4754 gnd.n1522 585
R4210 gnd.n3397 gnd.n1522 585
R4211 gnd.n4755 gnd.n1521 585
R4212 gnd.n3348 gnd.n1521 585
R4213 gnd.n3369 gnd.n1519 585
R4214 gnd.n3370 gnd.n3369 585
R4215 gnd.n4759 gnd.n1518 585
R4216 gnd.n2230 gnd.n1518 585
R4217 gnd.n4760 gnd.n1517 585
R4218 gnd.n2228 gnd.n1517 585
R4219 gnd.n4761 gnd.n1516 585
R4220 gnd.n2235 gnd.n1516 585
R4221 gnd.n2239 gnd.n1514 585
R4222 gnd.n2240 gnd.n2239 585
R4223 gnd.n4765 gnd.n1513 585
R4224 gnd.n3299 gnd.n1513 585
R4225 gnd.n4766 gnd.n1512 585
R4226 gnd.n2259 gnd.n1512 585
R4227 gnd.n4767 gnd.n1511 585
R4228 gnd.n2251 gnd.n1511 585
R4229 gnd.n1508 gnd.n1506 585
R4230 gnd.n3283 gnd.n1506 585
R4231 gnd.n4772 gnd.n4771 585
R4232 gnd.n4773 gnd.n4772 585
R4233 gnd.n1507 gnd.n1505 585
R4234 gnd.n3268 gnd.n1505 585
R4235 gnd.n3252 gnd.n3251 585
R4236 gnd.n3251 gnd.n1493 585
R4237 gnd.n2360 gnd.n2358 585
R4238 gnd.n2358 gnd.n1491 585
R4239 gnd.n3257 gnd.n3256 585
R4240 gnd.n3258 gnd.n3257 585
R4241 gnd.n2359 gnd.n2357 585
R4242 gnd.n2357 gnd.n1433 585
R4243 gnd.n3248 gnd.n3247 585
R4244 gnd.n3247 gnd.n3246 585
R4245 gnd.n2363 gnd.n2362 585
R4246 gnd.n3233 gnd.n2363 585
R4247 gnd.n2384 gnd.n2382 585
R4248 gnd.n2382 gnd.n2372 585
R4249 gnd.n3221 gnd.n3220 585
R4250 gnd.n3222 gnd.n3221 585
R4251 gnd.n2383 gnd.n2381 585
R4252 gnd.n2390 gnd.n2381 585
R4253 gnd.n3215 gnd.n3214 585
R4254 gnd.n3214 gnd.n3213 585
R4255 gnd.n2387 gnd.n2386 585
R4256 gnd.n3201 gnd.n2387 585
R4257 gnd.n3178 gnd.n3177 585
R4258 gnd.n3176 gnd.n2940 585
R4259 gnd.n2942 gnd.n2939 585
R4260 gnd.n3180 gnd.n2939 585
R4261 gnd.n3172 gnd.n2944 585
R4262 gnd.n3171 gnd.n2945 585
R4263 gnd.n3170 gnd.n2946 585
R4264 gnd.n3062 gnd.n2947 585
R4265 gnd.n3165 gnd.n3063 585
R4266 gnd.n3164 gnd.n3064 585
R4267 gnd.n3163 gnd.n3065 585
R4268 gnd.n3075 gnd.n3066 585
R4269 gnd.n3156 gnd.n3076 585
R4270 gnd.n3155 gnd.n3077 585
R4271 gnd.n3079 gnd.n3078 585
R4272 gnd.n3148 gnd.n3087 585
R4273 gnd.n3147 gnd.n3088 585
R4274 gnd.n3098 gnd.n3089 585
R4275 gnd.n3140 gnd.n3099 585
R4276 gnd.n3139 gnd.n3100 585
R4277 gnd.n3102 gnd.n3101 585
R4278 gnd.n3132 gnd.n3110 585
R4279 gnd.n3131 gnd.n3111 585
R4280 gnd.n3121 gnd.n3112 585
R4281 gnd.n3124 gnd.n3122 585
R4282 gnd.n3123 gnd.n2414 585
R4283 gnd.n3183 gnd.n3182 585
R4284 gnd.n2415 gnd.n2401 585
R4285 gnd.n3194 gnd.n2402 585
R4286 gnd.n3195 gnd.n2398 585
R4287 gnd.n1938 gnd.n1599 585
R4288 gnd.n4663 gnd.n1599 585
R4289 gnd.n4065 gnd.n4064 585
R4290 gnd.n4066 gnd.n4065 585
R4291 gnd.n1937 gnd.n1936 585
R4292 gnd.n4068 gnd.n1936 585
R4293 gnd.n3882 gnd.n3881 585
R4294 gnd.n3881 gnd.n1935 585
R4295 gnd.n3880 gnd.n3879 585
R4296 gnd.n3880 gnd.n1922 585
R4297 gnd.n3878 gnd.n1921 585
R4298 gnd.n4077 gnd.n1921 585
R4299 gnd.n1940 gnd.n1920 585
R4300 gnd.n4079 gnd.n1920 585
R4301 gnd.n3874 gnd.n3873 585
R4302 gnd.n3873 gnd.n1919 585
R4303 gnd.n3872 gnd.n1942 585
R4304 gnd.n3872 gnd.n3871 585
R4305 gnd.n3870 gnd.n3867 585
R4306 gnd.n3870 gnd.n3869 585
R4307 gnd.n1943 gnd.n1909 585
R4308 gnd.n4088 gnd.n1909 585
R4309 gnd.n3863 gnd.n3862 585
R4310 gnd.n3862 gnd.n3861 585
R4311 gnd.n1946 gnd.n1945 585
R4312 gnd.n1951 gnd.n1946 585
R4313 gnd.n1970 gnd.n1958 585
R4314 gnd.n3844 gnd.n1958 585
R4315 gnd.n3827 gnd.n3826 585
R4316 gnd.n3828 gnd.n3827 585
R4317 gnd.n1969 gnd.n1968 585
R4318 gnd.n1976 gnd.n1968 585
R4319 gnd.n3821 gnd.n3820 585
R4320 gnd.n3820 gnd.n3819 585
R4321 gnd.n1973 gnd.n1972 585
R4322 gnd.n1982 gnd.n1973 585
R4323 gnd.n3739 gnd.n1989 585
R4324 gnd.n3798 gnd.n1989 585
R4325 gnd.n3738 gnd.n1997 585
R4326 gnd.n3785 gnd.n1997 585
R4327 gnd.n3743 gnd.n3737 585
R4328 gnd.n3737 gnd.n3736 585
R4329 gnd.n3744 gnd.n3735 585
R4330 gnd.n3735 gnd.n2010 585
R4331 gnd.n3745 gnd.n3734 585
R4332 gnd.n3734 gnd.n2005 585
R4333 gnd.n2026 gnd.n2017 585
R4334 gnd.n3759 gnd.n2017 585
R4335 gnd.n3750 gnd.n3749 585
R4336 gnd.n3751 gnd.n3750 585
R4337 gnd.n2025 gnd.n2024 585
R4338 gnd.n3659 gnd.n2024 585
R4339 gnd.n3730 gnd.n3729 585
R4340 gnd.n3729 gnd.n3728 585
R4341 gnd.n2029 gnd.n2028 585
R4342 gnd.n3720 gnd.n2029 585
R4343 gnd.n2055 gnd.n2053 585
R4344 gnd.n2053 gnd.n2045 585
R4345 gnd.n3697 gnd.n3696 585
R4346 gnd.n3699 gnd.n3697 585
R4347 gnd.n2054 gnd.n2052 585
R4348 gnd.n2052 gnd.n2049 585
R4349 gnd.n3691 gnd.n3690 585
R4350 gnd.n3690 gnd.n3689 585
R4351 gnd.n2058 gnd.n2057 585
R4352 gnd.n2067 gnd.n2058 585
R4353 gnd.n3571 gnd.n3569 585
R4354 gnd.n3569 gnd.n3568 585
R4355 gnd.n3572 gnd.n3565 585
R4356 gnd.n3565 gnd.n2072 585
R4357 gnd.n3573 gnd.n2080 585
R4358 gnd.n3630 gnd.n2080 585
R4359 gnd.n3563 gnd.n2087 585
R4360 gnd.n3619 gnd.n2087 585
R4361 gnd.n3577 gnd.n3562 585
R4362 gnd.n3562 gnd.n2093 585
R4363 gnd.n3578 gnd.n3561 585
R4364 gnd.n3561 gnd.n2100 585
R4365 gnd.n3579 gnd.n3560 585
R4366 gnd.n3560 gnd.n3559 585
R4367 gnd.n2117 gnd.n2107 585
R4368 gnd.n3594 gnd.n2107 585
R4369 gnd.n3584 gnd.n3583 585
R4370 gnd.n3586 gnd.n3584 585
R4371 gnd.n2116 gnd.n2115 585
R4372 gnd.n3547 gnd.n2115 585
R4373 gnd.n3520 gnd.n3519 585
R4374 gnd.n3519 gnd.n3518 585
R4375 gnd.n2140 gnd.n2138 585
R4376 gnd.n2138 gnd.n2130 585
R4377 gnd.n3525 gnd.n3524 585
R4378 gnd.n3527 gnd.n3525 585
R4379 gnd.n2139 gnd.n2137 585
R4380 gnd.n3507 gnd.n2137 585
R4381 gnd.n3479 gnd.n3478 585
R4382 gnd.n3480 gnd.n3479 585
R4383 gnd.n2164 gnd.n2163 585
R4384 gnd.n2163 gnd.n2153 585
R4385 gnd.n3474 gnd.n3473 585
R4386 gnd.n3473 gnd.n3472 585
R4387 gnd.n3470 gnd.n2166 585
R4388 gnd.n3470 gnd.n2158 585
R4389 gnd.n3469 gnd.n2168 585
R4390 gnd.n3469 gnd.n3468 585
R4391 gnd.n3384 gnd.n2167 585
R4392 gnd.n3460 gnd.n2167 585
R4393 gnd.n3385 gnd.n2185 585
R4394 gnd.n3447 gnd.n2185 585
R4395 gnd.n3381 gnd.n3380 585
R4396 gnd.n3380 gnd.n2190 585
R4397 gnd.n3389 gnd.n3379 585
R4398 gnd.n3379 gnd.n3378 585
R4399 gnd.n3390 gnd.n3376 585
R4400 gnd.n3376 gnd.n2195 585
R4401 gnd.n3391 gnd.n2202 585
R4402 gnd.n3419 gnd.n2202 585
R4403 gnd.n2216 gnd.n2210 585
R4404 gnd.n3410 gnd.n2210 585
R4405 gnd.n3396 gnd.n3395 585
R4406 gnd.n3397 gnd.n3396 585
R4407 gnd.n2215 gnd.n2214 585
R4408 gnd.n3348 gnd.n2214 585
R4409 gnd.n3372 gnd.n3371 585
R4410 gnd.n3371 gnd.n3370 585
R4411 gnd.n2219 gnd.n2218 585
R4412 gnd.n2230 gnd.n2219 585
R4413 gnd.n3292 gnd.n3291 585
R4414 gnd.n3291 gnd.n2228 585
R4415 gnd.n3293 gnd.n3290 585
R4416 gnd.n3290 gnd.n2235 585
R4417 gnd.n2263 gnd.n2261 585
R4418 gnd.n2261 gnd.n2240 585
R4419 gnd.n3298 gnd.n3297 585
R4420 gnd.n3299 gnd.n3298 585
R4421 gnd.n2262 gnd.n2260 585
R4422 gnd.n2260 gnd.n2259 585
R4423 gnd.n3286 gnd.n3285 585
R4424 gnd.n3285 gnd.n2251 585
R4425 gnd.n3284 gnd.n2265 585
R4426 gnd.n3284 gnd.n3283 585
R4427 gnd.n2274 gnd.n1503 585
R4428 gnd.n4773 gnd.n1503 585
R4429 gnd.n3267 gnd.n3266 585
R4430 gnd.n3268 gnd.n3267 585
R4431 gnd.n2273 gnd.n2272 585
R4432 gnd.n2272 gnd.n1493 585
R4433 gnd.n3261 gnd.n3260 585
R4434 gnd.n3260 gnd.n1491 585
R4435 gnd.n3259 gnd.n2276 585
R4436 gnd.n3259 gnd.n3258 585
R4437 gnd.n3227 gnd.n2277 585
R4438 gnd.n2277 gnd.n1433 585
R4439 gnd.n2375 gnd.n2365 585
R4440 gnd.n3246 gnd.n2365 585
R4441 gnd.n3232 gnd.n3231 585
R4442 gnd.n3233 gnd.n3232 585
R4443 gnd.n2374 gnd.n2373 585
R4444 gnd.n2373 gnd.n2372 585
R4445 gnd.n3224 gnd.n3223 585
R4446 gnd.n3223 gnd.n3222 585
R4447 gnd.n2378 gnd.n2377 585
R4448 gnd.n2390 gnd.n2378 585
R4449 gnd.n2399 gnd.n2389 585
R4450 gnd.n3213 gnd.n2389 585
R4451 gnd.n3200 gnd.n3199 585
R4452 gnd.n3201 gnd.n3200 585
R4453 gnd.n4039 gnd.n3894 585
R4454 gnd.n3894 gnd.n1609 585
R4455 gnd.n4040 gnd.n4037 585
R4456 gnd.n4035 gnd.n3912 585
R4457 gnd.n4034 gnd.n4033 585
R4458 gnd.n4018 gnd.n3914 585
R4459 gnd.n4020 gnd.n4019 585
R4460 gnd.n4016 gnd.n3921 585
R4461 gnd.n4015 gnd.n4014 585
R4462 gnd.n3999 gnd.n3923 585
R4463 gnd.n4001 gnd.n4000 585
R4464 gnd.n3997 gnd.n3930 585
R4465 gnd.n3996 gnd.n3995 585
R4466 gnd.n3980 gnd.n3932 585
R4467 gnd.n3982 gnd.n3981 585
R4468 gnd.n3978 gnd.n3939 585
R4469 gnd.n3977 gnd.n3976 585
R4470 gnd.n3965 gnd.n3941 585
R4471 gnd.n3967 gnd.n3966 585
R4472 gnd.n3963 gnd.n3942 585
R4473 gnd.n3962 gnd.n3961 585
R4474 gnd.n3954 gnd.n3944 585
R4475 gnd.n3956 gnd.n3955 585
R4476 gnd.n3952 gnd.n3946 585
R4477 gnd.n3951 gnd.n3950 585
R4478 gnd.n3948 gnd.n1597 585
R4479 gnd.n4060 gnd.n4059 585
R4480 gnd.n4057 gnd.n3892 585
R4481 gnd.n4056 gnd.n3893 585
R4482 gnd.n4054 gnd.n4053 585
R4483 gnd.n4178 gnd.n1904 482.89
R4484 gnd.n4181 gnd.n4180 482.89
R4485 gnd.n2354 gnd.n2278 482.89
R4486 gnd.n4849 gnd.n1468 482.89
R4487 gnd.n2279 gnd.t270 443.966
R4488 gnd.n1898 gnd.t293 443.966
R4489 gnd.n4786 gnd.t318 443.966
R4490 gnd.n4112 gnd.t223 443.966
R4491 gnd.n6750 gnd.n6749 434.747
R4492 gnd.n2411 gnd.t260 371.625
R4493 gnd.n3905 gnd.t287 371.625
R4494 gnd.n2404 gnd.t312 371.625
R4495 gnd.n4318 gnd.t284 371.625
R4496 gnd.n4370 gnd.t281 371.625
R4497 gnd.n1829 gnd.t212 371.625
R4498 gnd.n313 gnd.t309 371.625
R4499 gnd.n280 gnd.t227 371.625
R4500 gnd.n7638 gnd.t267 371.625
R4501 gnd.n350 gnd.t254 371.625
R4502 gnd.n1090 gnd.t241 371.625
R4503 gnd.n1112 gnd.t238 371.625
R4504 gnd.n1134 gnd.t216 371.625
R4505 gnd.n2550 gnd.t296 371.625
R4506 gnd.n1409 gnd.t302 371.625
R4507 gnd.n2949 gnd.t234 371.625
R4508 gnd.n2971 gnd.t257 371.625
R4509 gnd.n3895 gnd.t244 371.625
R4510 gnd.n5761 gnd.t274 323.425
R4511 gnd.n5195 gnd.t305 323.425
R4512 gnd.n6406 gnd.n6380 289.615
R4513 gnd.n6374 gnd.n6348 289.615
R4514 gnd.n6342 gnd.n6316 289.615
R4515 gnd.n6311 gnd.n6285 289.615
R4516 gnd.n6279 gnd.n6253 289.615
R4517 gnd.n6247 gnd.n6221 289.615
R4518 gnd.n6215 gnd.n6189 289.615
R4519 gnd.n6184 gnd.n6158 289.615
R4520 gnd.n5611 gnd.t208 279.217
R4521 gnd.n5239 gnd.t204 279.217
R4522 gnd.n1475 gnd.t301 260.649
R4523 gnd.n4104 gnd.t222 260.649
R4524 gnd.n4851 gnd.n4850 256.663
R4525 gnd.n4851 gnd.n1434 256.663
R4526 gnd.n4851 gnd.n1435 256.663
R4527 gnd.n4851 gnd.n1436 256.663
R4528 gnd.n4851 gnd.n1437 256.663
R4529 gnd.n4851 gnd.n1438 256.663
R4530 gnd.n4851 gnd.n1439 256.663
R4531 gnd.n4851 gnd.n1440 256.663
R4532 gnd.n4851 gnd.n1441 256.663
R4533 gnd.n4851 gnd.n1442 256.663
R4534 gnd.n4851 gnd.n1443 256.663
R4535 gnd.n4851 gnd.n1444 256.663
R4536 gnd.n4851 gnd.n1445 256.663
R4537 gnd.n4851 gnd.n1446 256.663
R4538 gnd.n4851 gnd.n1447 256.663
R4539 gnd.n4851 gnd.n1448 256.663
R4540 gnd.n4854 gnd.n1431 256.663
R4541 gnd.n4852 gnd.n4851 256.663
R4542 gnd.n4851 gnd.n1449 256.663
R4543 gnd.n4851 gnd.n1450 256.663
R4544 gnd.n4851 gnd.n1451 256.663
R4545 gnd.n4851 gnd.n1452 256.663
R4546 gnd.n4851 gnd.n1453 256.663
R4547 gnd.n4851 gnd.n1454 256.663
R4548 gnd.n4851 gnd.n1455 256.663
R4549 gnd.n4851 gnd.n1456 256.663
R4550 gnd.n4851 gnd.n1457 256.663
R4551 gnd.n4851 gnd.n1458 256.663
R4552 gnd.n4851 gnd.n1459 256.663
R4553 gnd.n4851 gnd.n1460 256.663
R4554 gnd.n4851 gnd.n1461 256.663
R4555 gnd.n4851 gnd.n1462 256.663
R4556 gnd.n4851 gnd.n1463 256.663
R4557 gnd.n4851 gnd.n1464 256.663
R4558 gnd.n4246 gnd.n1882 256.663
R4559 gnd.n4246 gnd.n1883 256.663
R4560 gnd.n4246 gnd.n1884 256.663
R4561 gnd.n4246 gnd.n1885 256.663
R4562 gnd.n4246 gnd.n1886 256.663
R4563 gnd.n4246 gnd.n1887 256.663
R4564 gnd.n4246 gnd.n1888 256.663
R4565 gnd.n4246 gnd.n1889 256.663
R4566 gnd.n4246 gnd.n1890 256.663
R4567 gnd.n4246 gnd.n1891 256.663
R4568 gnd.n4246 gnd.n1892 256.663
R4569 gnd.n4246 gnd.n1893 256.663
R4570 gnd.n4246 gnd.n1894 256.663
R4571 gnd.n4246 gnd.n1895 256.663
R4572 gnd.n4246 gnd.n1896 256.663
R4573 gnd.n4246 gnd.n4243 256.663
R4574 gnd.n4249 gnd.n1863 256.663
R4575 gnd.n4247 gnd.n4246 256.663
R4576 gnd.n4246 gnd.n1881 256.663
R4577 gnd.n4246 gnd.n1880 256.663
R4578 gnd.n4246 gnd.n1879 256.663
R4579 gnd.n4246 gnd.n1878 256.663
R4580 gnd.n4246 gnd.n1877 256.663
R4581 gnd.n4246 gnd.n1876 256.663
R4582 gnd.n4246 gnd.n1875 256.663
R4583 gnd.n4246 gnd.n1874 256.663
R4584 gnd.n4246 gnd.n1873 256.663
R4585 gnd.n4246 gnd.n1872 256.663
R4586 gnd.n4246 gnd.n1871 256.663
R4587 gnd.n4246 gnd.n1870 256.663
R4588 gnd.n4246 gnd.n1869 256.663
R4589 gnd.n4246 gnd.n1868 256.663
R4590 gnd.n4246 gnd.n1867 256.663
R4591 gnd.n4246 gnd.n1866 256.663
R4592 gnd.n5164 gnd.n1058 242.672
R4593 gnd.n5164 gnd.n1059 242.672
R4594 gnd.n5164 gnd.n1060 242.672
R4595 gnd.n5164 gnd.n1061 242.672
R4596 gnd.n5164 gnd.n1062 242.672
R4597 gnd.n5164 gnd.n1063 242.672
R4598 gnd.n5164 gnd.n1064 242.672
R4599 gnd.n5164 gnd.n1065 242.672
R4600 gnd.n5164 gnd.n1066 242.672
R4601 gnd.n3189 gnd.n1381 242.672
R4602 gnd.n2407 gnd.n1381 242.672
R4603 gnd.n3117 gnd.n1381 242.672
R4604 gnd.n3114 gnd.n1381 242.672
R4605 gnd.n3105 gnd.n1381 242.672
R4606 gnd.n3094 gnd.n1381 242.672
R4607 gnd.n3091 gnd.n1381 242.672
R4608 gnd.n3082 gnd.n1381 242.672
R4609 gnd.n3071 gnd.n1381 242.672
R4610 gnd.n5666 gnd.n5575 242.672
R4611 gnd.n5579 gnd.n5575 242.672
R4612 gnd.n5659 gnd.n5575 242.672
R4613 gnd.n5653 gnd.n5575 242.672
R4614 gnd.n5651 gnd.n5575 242.672
R4615 gnd.n5645 gnd.n5575 242.672
R4616 gnd.n5643 gnd.n5575 242.672
R4617 gnd.n5637 gnd.n5575 242.672
R4618 gnd.n5635 gnd.n5575 242.672
R4619 gnd.n5629 gnd.n5575 242.672
R4620 gnd.n5627 gnd.n5575 242.672
R4621 gnd.n5620 gnd.n5575 242.672
R4622 gnd.n5618 gnd.n5575 242.672
R4623 gnd.n6462 gnd.n5165 242.672
R4624 gnd.n6468 gnd.n5165 242.672
R4625 gnd.n5242 gnd.n5165 242.672
R4626 gnd.n6475 gnd.n5165 242.672
R4627 gnd.n5233 gnd.n5165 242.672
R4628 gnd.n6482 gnd.n5165 242.672
R4629 gnd.n5226 gnd.n5165 242.672
R4630 gnd.n6489 gnd.n5165 242.672
R4631 gnd.n5219 gnd.n5165 242.672
R4632 gnd.n6496 gnd.n5165 242.672
R4633 gnd.n5212 gnd.n5165 242.672
R4634 gnd.n6503 gnd.n5165 242.672
R4635 gnd.n5205 gnd.n5165 242.672
R4636 gnd.n3970 gnd.n1610 242.672
R4637 gnd.n3987 gnd.n1610 242.672
R4638 gnd.n3989 gnd.n1610 242.672
R4639 gnd.n4006 gnd.n1610 242.672
R4640 gnd.n4008 gnd.n1610 242.672
R4641 gnd.n4025 gnd.n1610 242.672
R4642 gnd.n4027 gnd.n1610 242.672
R4643 gnd.n4045 gnd.n1610 242.672
R4644 gnd.n4047 gnd.n1610 242.672
R4645 gnd.n347 gnd.n212 242.672
R4646 gnd.n7534 gnd.n212 242.672
R4647 gnd.n343 gnd.n212 242.672
R4648 gnd.n7541 gnd.n212 242.672
R4649 gnd.n336 gnd.n212 242.672
R4650 gnd.n7548 gnd.n212 242.672
R4651 gnd.n329 gnd.n212 242.672
R4652 gnd.n7555 gnd.n212 242.672
R4653 gnd.n322 gnd.n212 242.672
R4654 gnd.n5795 gnd.n5794 242.672
R4655 gnd.n5795 gnd.n5736 242.672
R4656 gnd.n5795 gnd.n5737 242.672
R4657 gnd.n5795 gnd.n5738 242.672
R4658 gnd.n5795 gnd.n5739 242.672
R4659 gnd.n5795 gnd.n5740 242.672
R4660 gnd.n5795 gnd.n5741 242.672
R4661 gnd.n5795 gnd.n5742 242.672
R4662 gnd.n6514 gnd.n5165 242.672
R4663 gnd.n5198 gnd.n5165 242.672
R4664 gnd.n6521 gnd.n5165 242.672
R4665 gnd.n5189 gnd.n5165 242.672
R4666 gnd.n6528 gnd.n5165 242.672
R4667 gnd.n5182 gnd.n5165 242.672
R4668 gnd.n6535 gnd.n5165 242.672
R4669 gnd.n5175 gnd.n5165 242.672
R4670 gnd.n5164 gnd.n5163 242.672
R4671 gnd.n5164 gnd.n1030 242.672
R4672 gnd.n5164 gnd.n1031 242.672
R4673 gnd.n5164 gnd.n1032 242.672
R4674 gnd.n5164 gnd.n1033 242.672
R4675 gnd.n5164 gnd.n1034 242.672
R4676 gnd.n5164 gnd.n1035 242.672
R4677 gnd.n5164 gnd.n1036 242.672
R4678 gnd.n5164 gnd.n1037 242.672
R4679 gnd.n5164 gnd.n1038 242.672
R4680 gnd.n5164 gnd.n1039 242.672
R4681 gnd.n5164 gnd.n1040 242.672
R4682 gnd.n5164 gnd.n1041 242.672
R4683 gnd.n5164 gnd.n1042 242.672
R4684 gnd.n5164 gnd.n1043 242.672
R4685 gnd.n5164 gnd.n1044 242.672
R4686 gnd.n5164 gnd.n1045 242.672
R4687 gnd.n5164 gnd.n1046 242.672
R4688 gnd.n5164 gnd.n1047 242.672
R4689 gnd.n5164 gnd.n1048 242.672
R4690 gnd.n5164 gnd.n1049 242.672
R4691 gnd.n5164 gnd.n1050 242.672
R4692 gnd.n5164 gnd.n1051 242.672
R4693 gnd.n5164 gnd.n1052 242.672
R4694 gnd.n5164 gnd.n1053 242.672
R4695 gnd.n5164 gnd.n1054 242.672
R4696 gnd.n5164 gnd.n1055 242.672
R4697 gnd.n5164 gnd.n1056 242.672
R4698 gnd.n5164 gnd.n1057 242.672
R4699 gnd.n3056 gnd.n1381 242.672
R4700 gnd.n2952 gnd.n1381 242.672
R4701 gnd.n3046 gnd.n1381 242.672
R4702 gnd.n2956 gnd.n1381 242.672
R4703 gnd.n3036 gnd.n1381 242.672
R4704 gnd.n2960 gnd.n1381 242.672
R4705 gnd.n3026 gnd.n1381 242.672
R4706 gnd.n2964 gnd.n1381 242.672
R4707 gnd.n3016 gnd.n1381 242.672
R4708 gnd.n2968 gnd.n1381 242.672
R4709 gnd.n3006 gnd.n1381 242.672
R4710 gnd.n2974 gnd.n1381 242.672
R4711 gnd.n2996 gnd.n1381 242.672
R4712 gnd.n2978 gnd.n1381 242.672
R4713 gnd.n2986 gnd.n1381 242.672
R4714 gnd.n2983 gnd.n1381 242.672
R4715 gnd.n4855 gnd.n1427 242.672
R4716 gnd.n1426 gnd.n1381 242.672
R4717 gnd.n4859 gnd.n1381 242.672
R4718 gnd.n1420 gnd.n1381 242.672
R4719 gnd.n4866 gnd.n1381 242.672
R4720 gnd.n1413 gnd.n1381 242.672
R4721 gnd.n4874 gnd.n1381 242.672
R4722 gnd.n1404 gnd.n1381 242.672
R4723 gnd.n4881 gnd.n1381 242.672
R4724 gnd.n1397 gnd.n1381 242.672
R4725 gnd.n4888 gnd.n1381 242.672
R4726 gnd.n1390 gnd.n1381 242.672
R4727 gnd.n4895 gnd.n1381 242.672
R4728 gnd.n4898 gnd.n1381 242.672
R4729 gnd.n4279 gnd.n1610 242.672
R4730 gnd.n4282 gnd.n1610 242.672
R4731 gnd.n4290 gnd.n1610 242.672
R4732 gnd.n4292 gnd.n1610 242.672
R4733 gnd.n4300 gnd.n1610 242.672
R4734 gnd.n4302 gnd.n1610 242.672
R4735 gnd.n4310 gnd.n1610 242.672
R4736 gnd.n4312 gnd.n1610 242.672
R4737 gnd.n4323 gnd.n1610 242.672
R4738 gnd.n4325 gnd.n1610 242.672
R4739 gnd.n4333 gnd.n1610 242.672
R4740 gnd.n4335 gnd.n1610 242.672
R4741 gnd.n4344 gnd.n1610 242.672
R4742 gnd.n4345 gnd.n4250 242.672
R4743 gnd.n4346 gnd.n1610 242.672
R4744 gnd.n4348 gnd.n1610 242.672
R4745 gnd.n4356 gnd.n1610 242.672
R4746 gnd.n4358 gnd.n1610 242.672
R4747 gnd.n4366 gnd.n1610 242.672
R4748 gnd.n4368 gnd.n1610 242.672
R4749 gnd.n4378 gnd.n1610 242.672
R4750 gnd.n4380 gnd.n1610 242.672
R4751 gnd.n4388 gnd.n1610 242.672
R4752 gnd.n4390 gnd.n1610 242.672
R4753 gnd.n4398 gnd.n1610 242.672
R4754 gnd.n4400 gnd.n1610 242.672
R4755 gnd.n4408 gnd.n1610 242.672
R4756 gnd.n4410 gnd.n1610 242.672
R4757 gnd.n4419 gnd.n1610 242.672
R4758 gnd.n4422 gnd.n1610 242.672
R4759 gnd.n7566 gnd.n212 242.672
R4760 gnd.n316 gnd.n212 242.672
R4761 gnd.n7573 gnd.n212 242.672
R4762 gnd.n307 gnd.n212 242.672
R4763 gnd.n7580 gnd.n212 242.672
R4764 gnd.n300 gnd.n212 242.672
R4765 gnd.n7587 gnd.n212 242.672
R4766 gnd.n293 gnd.n212 242.672
R4767 gnd.n7594 gnd.n212 242.672
R4768 gnd.n7597 gnd.n212 242.672
R4769 gnd.n284 gnd.n212 242.672
R4770 gnd.n7606 gnd.n212 242.672
R4771 gnd.n275 gnd.n212 242.672
R4772 gnd.n7613 gnd.n212 242.672
R4773 gnd.n268 gnd.n212 242.672
R4774 gnd.n7620 gnd.n212 242.672
R4775 gnd.n261 gnd.n212 242.672
R4776 gnd.n7627 gnd.n212 242.672
R4777 gnd.n254 gnd.n212 242.672
R4778 gnd.n7634 gnd.n212 242.672
R4779 gnd.n247 gnd.n212 242.672
R4780 gnd.n7644 gnd.n212 242.672
R4781 gnd.n240 gnd.n212 242.672
R4782 gnd.n7651 gnd.n212 242.672
R4783 gnd.n233 gnd.n212 242.672
R4784 gnd.n7658 gnd.n212 242.672
R4785 gnd.n226 gnd.n212 242.672
R4786 gnd.n7665 gnd.n212 242.672
R4787 gnd.n219 gnd.n212 242.672
R4788 gnd.n3180 gnd.n3179 242.672
R4789 gnd.n3180 gnd.n2927 242.672
R4790 gnd.n3180 gnd.n2928 242.672
R4791 gnd.n3180 gnd.n2929 242.672
R4792 gnd.n3180 gnd.n2930 242.672
R4793 gnd.n3180 gnd.n2931 242.672
R4794 gnd.n3180 gnd.n2932 242.672
R4795 gnd.n3180 gnd.n2933 242.672
R4796 gnd.n3180 gnd.n2934 242.672
R4797 gnd.n3180 gnd.n2935 242.672
R4798 gnd.n3180 gnd.n2936 242.672
R4799 gnd.n3180 gnd.n2937 242.672
R4800 gnd.n3181 gnd.n3180 242.672
R4801 gnd.n3180 gnd.n2938 242.672
R4802 gnd.n4036 gnd.n1609 242.672
R4803 gnd.n3913 gnd.n1609 242.672
R4804 gnd.n4017 gnd.n1609 242.672
R4805 gnd.n3922 gnd.n1609 242.672
R4806 gnd.n3998 gnd.n1609 242.672
R4807 gnd.n3931 gnd.n1609 242.672
R4808 gnd.n3979 gnd.n1609 242.672
R4809 gnd.n3940 gnd.n1609 242.672
R4810 gnd.n3964 gnd.n1609 242.672
R4811 gnd.n3943 gnd.n1609 242.672
R4812 gnd.n3953 gnd.n1609 242.672
R4813 gnd.n3947 gnd.n1609 242.672
R4814 gnd.n4058 gnd.n1609 242.672
R4815 gnd.n4055 gnd.n1609 242.672
R4816 gnd.n216 gnd.n213 240.244
R4817 gnd.n7667 gnd.n7666 240.244
R4818 gnd.n7664 gnd.n220 240.244
R4819 gnd.n7660 gnd.n7659 240.244
R4820 gnd.n7657 gnd.n227 240.244
R4821 gnd.n7653 gnd.n7652 240.244
R4822 gnd.n7650 gnd.n234 240.244
R4823 gnd.n7646 gnd.n7645 240.244
R4824 gnd.n7643 gnd.n241 240.244
R4825 gnd.n7636 gnd.n7635 240.244
R4826 gnd.n7633 gnd.n248 240.244
R4827 gnd.n7629 gnd.n7628 240.244
R4828 gnd.n7626 gnd.n255 240.244
R4829 gnd.n7622 gnd.n7621 240.244
R4830 gnd.n7619 gnd.n262 240.244
R4831 gnd.n7615 gnd.n7614 240.244
R4832 gnd.n7612 gnd.n269 240.244
R4833 gnd.n7608 gnd.n7607 240.244
R4834 gnd.n7605 gnd.n276 240.244
R4835 gnd.n7598 gnd.n285 240.244
R4836 gnd.n7596 gnd.n7595 240.244
R4837 gnd.n7593 gnd.n287 240.244
R4838 gnd.n7589 gnd.n7588 240.244
R4839 gnd.n7586 gnd.n294 240.244
R4840 gnd.n7582 gnd.n7581 240.244
R4841 gnd.n7579 gnd.n301 240.244
R4842 gnd.n7575 gnd.n7574 240.244
R4843 gnd.n7572 gnd.n308 240.244
R4844 gnd.n7568 gnd.n7567 240.244
R4845 gnd.n1826 gnd.n1619 240.244
R4846 gnd.n1826 gnd.n1631 240.244
R4847 gnd.n4433 gnd.n1631 240.244
R4848 gnd.n4433 gnd.n1643 240.244
R4849 gnd.n4443 gnd.n1643 240.244
R4850 gnd.n4443 gnd.n1654 240.244
R4851 gnd.n4447 gnd.n1654 240.244
R4852 gnd.n4447 gnd.n1663 240.244
R4853 gnd.n4457 gnd.n1663 240.244
R4854 gnd.n4457 gnd.n1674 240.244
R4855 gnd.n1774 gnd.n1674 240.244
R4856 gnd.n1774 gnd.n1683 240.244
R4857 gnd.n4464 gnd.n1683 240.244
R4858 gnd.n4464 gnd.n1694 240.244
R4859 gnd.n4469 gnd.n1694 240.244
R4860 gnd.n4469 gnd.n1703 240.244
R4861 gnd.n4474 gnd.n1703 240.244
R4862 gnd.n4474 gnd.n1714 240.244
R4863 gnd.n4517 gnd.n1714 240.244
R4864 gnd.n4517 gnd.n1723 240.244
R4865 gnd.n4545 gnd.n1723 240.244
R4866 gnd.n4545 gnd.n1732 240.244
R4867 gnd.n1756 gnd.n1732 240.244
R4868 gnd.n1756 gnd.n1741 240.244
R4869 gnd.n1748 gnd.n1741 240.244
R4870 gnd.n4538 gnd.n1748 240.244
R4871 gnd.n4538 gnd.n4537 240.244
R4872 gnd.n4537 gnd.n86 240.244
R4873 gnd.n380 gnd.n86 240.244
R4874 gnd.n7447 gnd.n380 240.244
R4875 gnd.n7447 gnd.n103 240.244
R4876 gnd.n7451 gnd.n103 240.244
R4877 gnd.n7451 gnd.n115 240.244
R4878 gnd.n7461 gnd.n115 240.244
R4879 gnd.n7461 gnd.n124 240.244
R4880 gnd.n7465 gnd.n124 240.244
R4881 gnd.n7465 gnd.n133 240.244
R4882 gnd.n7475 gnd.n133 240.244
R4883 gnd.n7475 gnd.n144 240.244
R4884 gnd.n7479 gnd.n144 240.244
R4885 gnd.n7479 gnd.n154 240.244
R4886 gnd.n7490 gnd.n154 240.244
R4887 gnd.n7490 gnd.n164 240.244
R4888 gnd.n7509 gnd.n164 240.244
R4889 gnd.n7509 gnd.n173 240.244
R4890 gnd.n7505 gnd.n173 240.244
R4891 gnd.n7505 gnd.n183 240.244
R4892 gnd.n7502 gnd.n183 240.244
R4893 gnd.n7502 gnd.n192 240.244
R4894 gnd.n7499 gnd.n192 240.244
R4895 gnd.n7499 gnd.n202 240.244
R4896 gnd.n7496 gnd.n202 240.244
R4897 gnd.n7496 gnd.n210 240.244
R4898 gnd.n4281 gnd.n4280 240.244
R4899 gnd.n4283 gnd.n4281 240.244
R4900 gnd.n4289 gnd.n4271 240.244
R4901 gnd.n4293 gnd.n4291 240.244
R4902 gnd.n4299 gnd.n4267 240.244
R4903 gnd.n4303 gnd.n4301 240.244
R4904 gnd.n4309 gnd.n4263 240.244
R4905 gnd.n4313 gnd.n4311 240.244
R4906 gnd.n4322 gnd.n4259 240.244
R4907 gnd.n4326 gnd.n4324 240.244
R4908 gnd.n4332 gnd.n4255 240.244
R4909 gnd.n4336 gnd.n4334 240.244
R4910 gnd.n4343 gnd.n4251 240.244
R4911 gnd.n4349 gnd.n4347 240.244
R4912 gnd.n4355 gnd.n1857 240.244
R4913 gnd.n4359 gnd.n4357 240.244
R4914 gnd.n4365 gnd.n1853 240.244
R4915 gnd.n4369 gnd.n4367 240.244
R4916 gnd.n4377 gnd.n1849 240.244
R4917 gnd.n4381 gnd.n4379 240.244
R4918 gnd.n4387 gnd.n1845 240.244
R4919 gnd.n4391 gnd.n4389 240.244
R4920 gnd.n4397 gnd.n1841 240.244
R4921 gnd.n4401 gnd.n4399 240.244
R4922 gnd.n4407 gnd.n1837 240.244
R4923 gnd.n4411 gnd.n4409 240.244
R4924 gnd.n4418 gnd.n1833 240.244
R4925 gnd.n4421 gnd.n4420 240.244
R4926 gnd.n4646 gnd.n1624 240.244
R4927 gnd.n4642 gnd.n1624 240.244
R4928 gnd.n4642 gnd.n1629 240.244
R4929 gnd.n4634 gnd.n1629 240.244
R4930 gnd.n4634 gnd.n1646 240.244
R4931 gnd.n4630 gnd.n1646 240.244
R4932 gnd.n4630 gnd.n1652 240.244
R4933 gnd.n4622 gnd.n1652 240.244
R4934 gnd.n4622 gnd.n1666 240.244
R4935 gnd.n4618 gnd.n1666 240.244
R4936 gnd.n4618 gnd.n1672 240.244
R4937 gnd.n4610 gnd.n1672 240.244
R4938 gnd.n4610 gnd.n1686 240.244
R4939 gnd.n4606 gnd.n1686 240.244
R4940 gnd.n4606 gnd.n1692 240.244
R4941 gnd.n4598 gnd.n1692 240.244
R4942 gnd.n4598 gnd.n1706 240.244
R4943 gnd.n4594 gnd.n1706 240.244
R4944 gnd.n4594 gnd.n1712 240.244
R4945 gnd.n4586 gnd.n1712 240.244
R4946 gnd.n4586 gnd.n1726 240.244
R4947 gnd.n4582 gnd.n1726 240.244
R4948 gnd.n4582 gnd.n1730 240.244
R4949 gnd.n4574 gnd.n1730 240.244
R4950 gnd.n4574 gnd.n4573 240.244
R4951 gnd.n4573 gnd.n1746 240.244
R4952 gnd.n1746 gnd.n89 240.244
R4953 gnd.n7748 gnd.n89 240.244
R4954 gnd.n7748 gnd.n90 240.244
R4955 gnd.n100 gnd.n90 240.244
R4956 gnd.n7742 gnd.n100 240.244
R4957 gnd.n7742 gnd.n101 240.244
R4958 gnd.n7734 gnd.n101 240.244
R4959 gnd.n7734 gnd.n117 240.244
R4960 gnd.n7730 gnd.n117 240.244
R4961 gnd.n7730 gnd.n122 240.244
R4962 gnd.n7722 gnd.n122 240.244
R4963 gnd.n7722 gnd.n136 240.244
R4964 gnd.n7718 gnd.n136 240.244
R4965 gnd.n7718 gnd.n142 240.244
R4966 gnd.n7710 gnd.n142 240.244
R4967 gnd.n7710 gnd.n156 240.244
R4968 gnd.n7706 gnd.n156 240.244
R4969 gnd.n7706 gnd.n162 240.244
R4970 gnd.n7698 gnd.n162 240.244
R4971 gnd.n7698 gnd.n176 240.244
R4972 gnd.n7694 gnd.n176 240.244
R4973 gnd.n7694 gnd.n182 240.244
R4974 gnd.n7686 gnd.n182 240.244
R4975 gnd.n7686 gnd.n195 240.244
R4976 gnd.n7682 gnd.n195 240.244
R4977 gnd.n7682 gnd.n201 240.244
R4978 gnd.n7674 gnd.n201 240.244
R4979 gnd.n4899 gnd.n1377 240.244
R4980 gnd.n4897 gnd.n4896 240.244
R4981 gnd.n4894 gnd.n1383 240.244
R4982 gnd.n4890 gnd.n4889 240.244
R4983 gnd.n4887 gnd.n1391 240.244
R4984 gnd.n4883 gnd.n4882 240.244
R4985 gnd.n4880 gnd.n1398 240.244
R4986 gnd.n4876 gnd.n4875 240.244
R4987 gnd.n4873 gnd.n1405 240.244
R4988 gnd.n4868 gnd.n4867 240.244
R4989 gnd.n4865 gnd.n1414 240.244
R4990 gnd.n4861 gnd.n4860 240.244
R4991 gnd.n4858 gnd.n1421 240.244
R4992 gnd.n2985 gnd.n2984 240.244
R4993 gnd.n2988 gnd.n2987 240.244
R4994 gnd.n2995 gnd.n2994 240.244
R4995 gnd.n2998 gnd.n2997 240.244
R4996 gnd.n3005 gnd.n3004 240.244
R4997 gnd.n3008 gnd.n3007 240.244
R4998 gnd.n3015 gnd.n3014 240.244
R4999 gnd.n3018 gnd.n3017 240.244
R5000 gnd.n3025 gnd.n3024 240.244
R5001 gnd.n3028 gnd.n3027 240.244
R5002 gnd.n3035 gnd.n3034 240.244
R5003 gnd.n3038 gnd.n3037 240.244
R5004 gnd.n3045 gnd.n3044 240.244
R5005 gnd.n3048 gnd.n3047 240.244
R5006 gnd.n3055 gnd.n3054 240.244
R5007 gnd.n5042 gnd.n5041 240.244
R5008 gnd.n5041 gnd.n1141 240.244
R5009 gnd.n1153 gnd.n1141 240.244
R5010 gnd.n2532 gnd.n1153 240.244
R5011 gnd.n2532 gnd.n1165 240.244
R5012 gnd.n2536 gnd.n1165 240.244
R5013 gnd.n2536 gnd.n1175 240.244
R5014 gnd.n2539 gnd.n1175 240.244
R5015 gnd.n2539 gnd.n1185 240.244
R5016 gnd.n2630 gnd.n1185 240.244
R5017 gnd.n2630 gnd.n1195 240.244
R5018 gnd.n2634 gnd.n1195 240.244
R5019 gnd.n2634 gnd.n1205 240.244
R5020 gnd.n2683 gnd.n1205 240.244
R5021 gnd.n2683 gnd.n1215 240.244
R5022 gnd.n2687 gnd.n1215 240.244
R5023 gnd.n2687 gnd.n1225 240.244
R5024 gnd.n2698 gnd.n1225 240.244
R5025 gnd.n2698 gnd.n1236 240.244
R5026 gnd.n2703 gnd.n1236 240.244
R5027 gnd.n2703 gnd.n1246 240.244
R5028 gnd.n2509 gnd.n1246 240.244
R5029 gnd.n2509 gnd.n2504 240.244
R5030 gnd.n2716 gnd.n2504 240.244
R5031 gnd.n2716 gnd.n2489 240.244
R5032 gnd.n2489 gnd.n2483 240.244
R5033 gnd.n2496 gnd.n2483 240.244
R5034 gnd.n2496 gnd.n2477 240.244
R5035 gnd.n2477 gnd.n2475 240.244
R5036 gnd.n2475 gnd.n2461 240.244
R5037 gnd.n2461 gnd.n1263 240.244
R5038 gnd.n2774 gnd.n1263 240.244
R5039 gnd.n2774 gnd.n1275 240.244
R5040 gnd.n2780 gnd.n1275 240.244
R5041 gnd.n2780 gnd.n1284 240.244
R5042 gnd.n2787 gnd.n1284 240.244
R5043 gnd.n2787 gnd.n1294 240.244
R5044 gnd.n2448 gnd.n1294 240.244
R5045 gnd.n2448 gnd.n1304 240.244
R5046 gnd.n2850 gnd.n1304 240.244
R5047 gnd.n2850 gnd.n1314 240.244
R5048 gnd.n2855 gnd.n1314 240.244
R5049 gnd.n2855 gnd.n1324 240.244
R5050 gnd.n2865 gnd.n1324 240.244
R5051 gnd.n2865 gnd.n1334 240.244
R5052 gnd.n2430 gnd.n1334 240.244
R5053 gnd.n2430 gnd.n1344 240.244
R5054 gnd.n2872 gnd.n1344 240.244
R5055 gnd.n2872 gnd.n1354 240.244
R5056 gnd.n2877 gnd.n1354 240.244
R5057 gnd.n2877 gnd.n1365 240.244
R5058 gnd.n2882 gnd.n1365 240.244
R5059 gnd.n2882 gnd.n1374 240.244
R5060 gnd.n1070 gnd.n1069 240.244
R5061 gnd.n5157 gnd.n1069 240.244
R5062 gnd.n5155 gnd.n5154 240.244
R5063 gnd.n5151 gnd.n5150 240.244
R5064 gnd.n5147 gnd.n5146 240.244
R5065 gnd.n5143 gnd.n5142 240.244
R5066 gnd.n5139 gnd.n5138 240.244
R5067 gnd.n5135 gnd.n5134 240.244
R5068 gnd.n5131 gnd.n5130 240.244
R5069 gnd.n5126 gnd.n5125 240.244
R5070 gnd.n5122 gnd.n5121 240.244
R5071 gnd.n5118 gnd.n5117 240.244
R5072 gnd.n5114 gnd.n5113 240.244
R5073 gnd.n5110 gnd.n5109 240.244
R5074 gnd.n5106 gnd.n5105 240.244
R5075 gnd.n5102 gnd.n5101 240.244
R5076 gnd.n5098 gnd.n5097 240.244
R5077 gnd.n5094 gnd.n5093 240.244
R5078 gnd.n5090 gnd.n5089 240.244
R5079 gnd.n5086 gnd.n5085 240.244
R5080 gnd.n5082 gnd.n5081 240.244
R5081 gnd.n5078 gnd.n5077 240.244
R5082 gnd.n5074 gnd.n5073 240.244
R5083 gnd.n5070 gnd.n5069 240.244
R5084 gnd.n5066 gnd.n5065 240.244
R5085 gnd.n5062 gnd.n5061 240.244
R5086 gnd.n5058 gnd.n5057 240.244
R5087 gnd.n5054 gnd.n5053 240.244
R5088 gnd.n5050 gnd.n5049 240.244
R5089 gnd.n5039 gnd.n1071 240.244
R5090 gnd.n5039 gnd.n1144 240.244
R5091 gnd.n5035 gnd.n1144 240.244
R5092 gnd.n5035 gnd.n1151 240.244
R5093 gnd.n5027 gnd.n1151 240.244
R5094 gnd.n5027 gnd.n1168 240.244
R5095 gnd.n5023 gnd.n1168 240.244
R5096 gnd.n5023 gnd.n1174 240.244
R5097 gnd.n5015 gnd.n1174 240.244
R5098 gnd.n5015 gnd.n1187 240.244
R5099 gnd.n5011 gnd.n1187 240.244
R5100 gnd.n5011 gnd.n1193 240.244
R5101 gnd.n5003 gnd.n1193 240.244
R5102 gnd.n5003 gnd.n1208 240.244
R5103 gnd.n4999 gnd.n1208 240.244
R5104 gnd.n4999 gnd.n1214 240.244
R5105 gnd.n4991 gnd.n1214 240.244
R5106 gnd.n4991 gnd.n1228 240.244
R5107 gnd.n4987 gnd.n1228 240.244
R5108 gnd.n4987 gnd.n1234 240.244
R5109 gnd.n4979 gnd.n1234 240.244
R5110 gnd.n4979 gnd.n1249 240.244
R5111 gnd.n2722 gnd.n1249 240.244
R5112 gnd.n2722 gnd.n2486 240.244
R5113 gnd.n2748 gnd.n2486 240.244
R5114 gnd.n2751 gnd.n2748 240.244
R5115 gnd.n2751 gnd.n2476 240.244
R5116 gnd.n2762 gnd.n2476 240.244
R5117 gnd.n2765 gnd.n2762 240.244
R5118 gnd.n2765 gnd.n1261 240.244
R5119 gnd.n4973 gnd.n1261 240.244
R5120 gnd.n4973 gnd.n1262 240.244
R5121 gnd.n4965 gnd.n1262 240.244
R5122 gnd.n4965 gnd.n1277 240.244
R5123 gnd.n4961 gnd.n1277 240.244
R5124 gnd.n4961 gnd.n1282 240.244
R5125 gnd.n4953 gnd.n1282 240.244
R5126 gnd.n4953 gnd.n1297 240.244
R5127 gnd.n4949 gnd.n1297 240.244
R5128 gnd.n4949 gnd.n1303 240.244
R5129 gnd.n4941 gnd.n1303 240.244
R5130 gnd.n4941 gnd.n1316 240.244
R5131 gnd.n4937 gnd.n1316 240.244
R5132 gnd.n4937 gnd.n1322 240.244
R5133 gnd.n4929 gnd.n1322 240.244
R5134 gnd.n4929 gnd.n1337 240.244
R5135 gnd.n4925 gnd.n1337 240.244
R5136 gnd.n4925 gnd.n1343 240.244
R5137 gnd.n4917 gnd.n1343 240.244
R5138 gnd.n4917 gnd.n1357 240.244
R5139 gnd.n4913 gnd.n1357 240.244
R5140 gnd.n4913 gnd.n1363 240.244
R5141 gnd.n4905 gnd.n1363 240.244
R5142 gnd.n5172 gnd.n5167 240.244
R5143 gnd.n6537 gnd.n6536 240.244
R5144 gnd.n6534 gnd.n5176 240.244
R5145 gnd.n6530 gnd.n6529 240.244
R5146 gnd.n6527 gnd.n5183 240.244
R5147 gnd.n6523 gnd.n6522 240.244
R5148 gnd.n6520 gnd.n5190 240.244
R5149 gnd.n6516 gnd.n6515 240.244
R5150 gnd.n5807 gnd.n5527 240.244
R5151 gnd.n5527 gnd.n5518 240.244
R5152 gnd.n5825 gnd.n5518 240.244
R5153 gnd.n5826 gnd.n5825 240.244
R5154 gnd.n5826 gnd.n5506 240.244
R5155 gnd.n5506 gnd.n5495 240.244
R5156 gnd.n5857 gnd.n5495 240.244
R5157 gnd.n5858 gnd.n5857 240.244
R5158 gnd.n5859 gnd.n5858 240.244
R5159 gnd.n5859 gnd.n5480 240.244
R5160 gnd.n5861 gnd.n5480 240.244
R5161 gnd.n5861 gnd.n5465 240.244
R5162 gnd.n5902 gnd.n5465 240.244
R5163 gnd.n5903 gnd.n5902 240.244
R5164 gnd.n5906 gnd.n5903 240.244
R5165 gnd.n5906 gnd.n5447 240.244
R5166 gnd.n5938 gnd.n5447 240.244
R5167 gnd.n5938 gnd.n5433 240.244
R5168 gnd.n5960 gnd.n5433 240.244
R5169 gnd.n5961 gnd.n5960 240.244
R5170 gnd.n5961 gnd.n5420 240.244
R5171 gnd.n5420 gnd.n5409 240.244
R5172 gnd.n5992 gnd.n5409 240.244
R5173 gnd.n5993 gnd.n5992 240.244
R5174 gnd.n5994 gnd.n5993 240.244
R5175 gnd.n5994 gnd.n5330 240.244
R5176 gnd.n5330 gnd.n5329 240.244
R5177 gnd.n5329 gnd.n5314 240.244
R5178 gnd.n6045 gnd.n5314 240.244
R5179 gnd.n6046 gnd.n6045 240.244
R5180 gnd.n6046 gnd.n5301 240.244
R5181 gnd.n5301 gnd.n5290 240.244
R5182 gnd.n6079 gnd.n5290 240.244
R5183 gnd.n6080 gnd.n6079 240.244
R5184 gnd.n6082 gnd.n6080 240.244
R5185 gnd.n6082 gnd.n6081 240.244
R5186 gnd.n6081 gnd.n5270 240.244
R5187 gnd.n6119 gnd.n5270 240.244
R5188 gnd.n6119 gnd.n5257 240.244
R5189 gnd.n6145 gnd.n5257 240.244
R5190 gnd.n6146 gnd.n6145 240.244
R5191 gnd.n6147 gnd.n6146 240.244
R5192 gnd.n6147 gnd.n981 240.244
R5193 gnd.n6436 gnd.n981 240.244
R5194 gnd.n6436 gnd.n991 240.244
R5195 gnd.n6432 gnd.n991 240.244
R5196 gnd.n6432 gnd.n6431 240.244
R5197 gnd.n6431 gnd.n1004 240.244
R5198 gnd.n6427 gnd.n1004 240.244
R5199 gnd.n6427 gnd.n1017 240.244
R5200 gnd.n6423 gnd.n1017 240.244
R5201 gnd.n6423 gnd.n6422 240.244
R5202 gnd.n6422 gnd.n1029 240.244
R5203 gnd.n5744 gnd.n5743 240.244
R5204 gnd.n5788 gnd.n5743 240.244
R5205 gnd.n5786 gnd.n5785 240.244
R5206 gnd.n5782 gnd.n5781 240.244
R5207 gnd.n5778 gnd.n5777 240.244
R5208 gnd.n5774 gnd.n5773 240.244
R5209 gnd.n5770 gnd.n5769 240.244
R5210 gnd.n5766 gnd.n5765 240.244
R5211 gnd.n5817 gnd.n5525 240.244
R5212 gnd.n5817 gnd.n5521 240.244
R5213 gnd.n5823 gnd.n5521 240.244
R5214 gnd.n5823 gnd.n5504 240.244
R5215 gnd.n5847 gnd.n5504 240.244
R5216 gnd.n5847 gnd.n5499 240.244
R5217 gnd.n5855 gnd.n5499 240.244
R5218 gnd.n5855 gnd.n5500 240.244
R5219 gnd.n5500 gnd.n5478 240.244
R5220 gnd.n5881 gnd.n5478 240.244
R5221 gnd.n5881 gnd.n5473 240.244
R5222 gnd.n5892 gnd.n5473 240.244
R5223 gnd.n5892 gnd.n5474 240.244
R5224 gnd.n5888 gnd.n5474 240.244
R5225 gnd.n5888 gnd.n5445 240.244
R5226 gnd.n5942 gnd.n5445 240.244
R5227 gnd.n5942 gnd.n5440 240.244
R5228 gnd.n5950 gnd.n5440 240.244
R5229 gnd.n5950 gnd.n5441 240.244
R5230 gnd.n5441 gnd.n5418 240.244
R5231 gnd.n5982 gnd.n5418 240.244
R5232 gnd.n5982 gnd.n5413 240.244
R5233 gnd.n5990 gnd.n5413 240.244
R5234 gnd.n5990 gnd.n5414 240.244
R5235 gnd.n5414 gnd.n5327 240.244
R5236 gnd.n6027 gnd.n5327 240.244
R5237 gnd.n6027 gnd.n5322 240.244
R5238 gnd.n6035 gnd.n5322 240.244
R5239 gnd.n6035 gnd.n5323 240.244
R5240 gnd.n5323 gnd.n5299 240.244
R5241 gnd.n6066 gnd.n5299 240.244
R5242 gnd.n6066 gnd.n5294 240.244
R5243 gnd.n6077 gnd.n5294 240.244
R5244 gnd.n6077 gnd.n5295 240.244
R5245 gnd.n6073 gnd.n5295 240.244
R5246 gnd.n6073 gnd.n5269 240.244
R5247 gnd.n6123 gnd.n5269 240.244
R5248 gnd.n6123 gnd.n5264 240.244
R5249 gnd.n6135 gnd.n5264 240.244
R5250 gnd.n6135 gnd.n5265 240.244
R5251 gnd.n6131 gnd.n5265 240.244
R5252 gnd.n6131 gnd.n982 240.244
R5253 gnd.n6572 gnd.n982 240.244
R5254 gnd.n6572 gnd.n983 240.244
R5255 gnd.n6568 gnd.n983 240.244
R5256 gnd.n6568 gnd.n989 240.244
R5257 gnd.n1006 gnd.n989 240.244
R5258 gnd.n6558 gnd.n1006 240.244
R5259 gnd.n6558 gnd.n1007 240.244
R5260 gnd.n6554 gnd.n1007 240.244
R5261 gnd.n6554 gnd.n1015 240.244
R5262 gnd.n5166 gnd.n1015 240.244
R5263 gnd.n6544 gnd.n5166 240.244
R5264 gnd.n319 gnd.n208 240.244
R5265 gnd.n7557 gnd.n7556 240.244
R5266 gnd.n7554 gnd.n323 240.244
R5267 gnd.n7550 gnd.n7549 240.244
R5268 gnd.n7547 gnd.n330 240.244
R5269 gnd.n7543 gnd.n7542 240.244
R5270 gnd.n7540 gnd.n337 240.244
R5271 gnd.n7536 gnd.n7535 240.244
R5272 gnd.n7533 gnd.n344 240.244
R5273 gnd.n3887 gnd.n1620 240.244
R5274 gnd.n3887 gnd.n1632 240.244
R5275 gnd.n4435 gnd.n1632 240.244
R5276 gnd.n4435 gnd.n1644 240.244
R5277 gnd.n4441 gnd.n1644 240.244
R5278 gnd.n4441 gnd.n1655 240.244
R5279 gnd.n4449 gnd.n1655 240.244
R5280 gnd.n4449 gnd.n1664 240.244
R5281 gnd.n4455 gnd.n1664 240.244
R5282 gnd.n4455 gnd.n1675 240.244
R5283 gnd.n4491 gnd.n1675 240.244
R5284 gnd.n4491 gnd.n1684 240.244
R5285 gnd.n1779 gnd.n1684 240.244
R5286 gnd.n1779 gnd.n1695 240.244
R5287 gnd.n1780 gnd.n1695 240.244
R5288 gnd.n1780 gnd.n1704 240.244
R5289 gnd.n4476 gnd.n1704 240.244
R5290 gnd.n4476 gnd.n1715 240.244
R5291 gnd.n1762 gnd.n1715 240.244
R5292 gnd.n1762 gnd.n1724 240.244
R5293 gnd.n4547 gnd.n1724 240.244
R5294 gnd.n4547 gnd.n1733 240.244
R5295 gnd.n4556 gnd.n1733 240.244
R5296 gnd.n4556 gnd.n1742 240.244
R5297 gnd.n1749 gnd.n1742 240.244
R5298 gnd.n1750 gnd.n1749 240.244
R5299 gnd.n1750 gnd.n82 240.244
R5300 gnd.n7750 gnd.n82 240.244
R5301 gnd.n7750 gnd.n84 240.244
R5302 gnd.n7445 gnd.n84 240.244
R5303 gnd.n7445 gnd.n104 240.244
R5304 gnd.n7453 gnd.n104 240.244
R5305 gnd.n7453 gnd.n116 240.244
R5306 gnd.n7459 gnd.n116 240.244
R5307 gnd.n7459 gnd.n125 240.244
R5308 gnd.n7467 gnd.n125 240.244
R5309 gnd.n7467 gnd.n134 240.244
R5310 gnd.n7473 gnd.n134 240.244
R5311 gnd.n7473 gnd.n145 240.244
R5312 gnd.n7481 gnd.n145 240.244
R5313 gnd.n7481 gnd.n155 240.244
R5314 gnd.n7488 gnd.n155 240.244
R5315 gnd.n7488 gnd.n165 240.244
R5316 gnd.n7511 gnd.n165 240.244
R5317 gnd.n7511 gnd.n174 240.244
R5318 gnd.n356 gnd.n174 240.244
R5319 gnd.n356 gnd.n184 240.244
R5320 gnd.n7518 gnd.n184 240.244
R5321 gnd.n7518 gnd.n193 240.244
R5322 gnd.n353 gnd.n193 240.244
R5323 gnd.n353 gnd.n203 240.244
R5324 gnd.n7525 gnd.n203 240.244
R5325 gnd.n7525 gnd.n211 240.244
R5326 gnd.n3986 gnd.n3935 240.244
R5327 gnd.n3990 gnd.n3988 240.244
R5328 gnd.n4005 gnd.n3926 240.244
R5329 gnd.n4009 gnd.n4007 240.244
R5330 gnd.n4024 gnd.n3917 240.244
R5331 gnd.n4028 gnd.n4026 240.244
R5332 gnd.n4044 gnd.n3908 240.244
R5333 gnd.n4048 gnd.n4046 240.244
R5334 gnd.n3904 gnd.n3903 240.244
R5335 gnd.n1634 gnd.n1622 240.244
R5336 gnd.n4640 gnd.n1634 240.244
R5337 gnd.n4640 gnd.n1635 240.244
R5338 gnd.n4636 gnd.n1635 240.244
R5339 gnd.n4636 gnd.n1641 240.244
R5340 gnd.n4628 gnd.n1641 240.244
R5341 gnd.n4628 gnd.n1656 240.244
R5342 gnd.n4624 gnd.n1656 240.244
R5343 gnd.n4624 gnd.n1661 240.244
R5344 gnd.n4616 gnd.n1661 240.244
R5345 gnd.n4616 gnd.n1677 240.244
R5346 gnd.n4612 gnd.n1677 240.244
R5347 gnd.n4612 gnd.n1682 240.244
R5348 gnd.n4604 gnd.n1682 240.244
R5349 gnd.n4604 gnd.n1696 240.244
R5350 gnd.n4600 gnd.n1696 240.244
R5351 gnd.n4600 gnd.n1701 240.244
R5352 gnd.n4592 gnd.n1701 240.244
R5353 gnd.n4592 gnd.n1717 240.244
R5354 gnd.n4588 gnd.n1717 240.244
R5355 gnd.n4588 gnd.n1722 240.244
R5356 gnd.n4580 gnd.n1722 240.244
R5357 gnd.n4580 gnd.n1734 240.244
R5358 gnd.n4576 gnd.n1734 240.244
R5359 gnd.n4576 gnd.n1739 240.244
R5360 gnd.n4525 gnd.n1739 240.244
R5361 gnd.n4535 gnd.n4525 240.244
R5362 gnd.n4535 gnd.n88 240.244
R5363 gnd.n4531 gnd.n88 240.244
R5364 gnd.n4531 gnd.n106 240.244
R5365 gnd.n7740 gnd.n106 240.244
R5366 gnd.n7740 gnd.n107 240.244
R5367 gnd.n7736 gnd.n107 240.244
R5368 gnd.n7736 gnd.n113 240.244
R5369 gnd.n7728 gnd.n113 240.244
R5370 gnd.n7728 gnd.n126 240.244
R5371 gnd.n7724 gnd.n126 240.244
R5372 gnd.n7724 gnd.n131 240.244
R5373 gnd.n7716 gnd.n131 240.244
R5374 gnd.n7716 gnd.n147 240.244
R5375 gnd.n7712 gnd.n147 240.244
R5376 gnd.n7712 gnd.n152 240.244
R5377 gnd.n7704 gnd.n152 240.244
R5378 gnd.n7704 gnd.n166 240.244
R5379 gnd.n7700 gnd.n166 240.244
R5380 gnd.n7700 gnd.n171 240.244
R5381 gnd.n7692 gnd.n171 240.244
R5382 gnd.n7692 gnd.n186 240.244
R5383 gnd.n7688 gnd.n186 240.244
R5384 gnd.n7688 gnd.n191 240.244
R5385 gnd.n7680 gnd.n191 240.244
R5386 gnd.n7680 gnd.n204 240.244
R5387 gnd.n7676 gnd.n204 240.244
R5388 gnd.n5202 gnd.n1026 240.244
R5389 gnd.n6505 gnd.n6504 240.244
R5390 gnd.n6502 gnd.n5206 240.244
R5391 gnd.n6498 gnd.n6497 240.244
R5392 gnd.n6495 gnd.n5213 240.244
R5393 gnd.n6491 gnd.n6490 240.244
R5394 gnd.n6488 gnd.n5220 240.244
R5395 gnd.n6484 gnd.n6483 240.244
R5396 gnd.n6481 gnd.n5227 240.244
R5397 gnd.n6477 gnd.n6476 240.244
R5398 gnd.n6474 gnd.n5234 240.244
R5399 gnd.n6470 gnd.n6469 240.244
R5400 gnd.n6467 gnd.n5244 240.244
R5401 gnd.n5675 gnd.n5571 240.244
R5402 gnd.n5681 gnd.n5571 240.244
R5403 gnd.n5681 gnd.n5563 240.244
R5404 gnd.n5691 gnd.n5563 240.244
R5405 gnd.n5691 gnd.n5559 240.244
R5406 gnd.n5697 gnd.n5559 240.244
R5407 gnd.n5697 gnd.n5550 240.244
R5408 gnd.n5707 gnd.n5550 240.244
R5409 gnd.n5707 gnd.n5545 240.244
R5410 gnd.n5735 gnd.n5545 240.244
R5411 gnd.n5735 gnd.n5546 240.244
R5412 gnd.n5546 gnd.n5538 240.244
R5413 gnd.n5730 gnd.n5538 240.244
R5414 gnd.n5730 gnd.n5528 240.244
R5415 gnd.n5727 gnd.n5528 240.244
R5416 gnd.n5727 gnd.n5517 240.244
R5417 gnd.n5724 gnd.n5517 240.244
R5418 gnd.n5724 gnd.n5507 240.244
R5419 gnd.n5721 gnd.n5507 240.244
R5420 gnd.n5721 gnd.n5485 240.244
R5421 gnd.n5870 gnd.n5485 240.244
R5422 gnd.n5870 gnd.n5481 240.244
R5423 gnd.n5878 gnd.n5481 240.244
R5424 gnd.n5878 gnd.n5471 240.244
R5425 gnd.n5471 gnd.n5452 240.244
R5426 gnd.n5917 gnd.n5452 240.244
R5427 gnd.n5917 gnd.n5453 240.244
R5428 gnd.n5453 gnd.n5448 240.244
R5429 gnd.n5937 gnd.n5448 240.244
R5430 gnd.n5937 gnd.n5438 240.244
R5431 gnd.n5932 gnd.n5438 240.244
R5432 gnd.n5932 gnd.n5432 240.244
R5433 gnd.n5928 gnd.n5432 240.244
R5434 gnd.n5928 gnd.n5421 240.244
R5435 gnd.n5924 gnd.n5421 240.244
R5436 gnd.n5924 gnd.n5399 240.244
R5437 gnd.n6003 gnd.n5399 240.244
R5438 gnd.n6003 gnd.n5331 240.244
R5439 gnd.n6024 gnd.n5331 240.244
R5440 gnd.n6024 gnd.n5320 240.244
R5441 gnd.n6020 gnd.n5320 240.244
R5442 gnd.n6020 gnd.n5313 240.244
R5443 gnd.n6017 gnd.n5313 240.244
R5444 gnd.n6017 gnd.n5302 240.244
R5445 gnd.n6014 gnd.n5302 240.244
R5446 gnd.n6014 gnd.n5281 240.244
R5447 gnd.n6089 gnd.n5281 240.244
R5448 gnd.n6089 gnd.n5277 240.244
R5449 gnd.n6110 gnd.n5277 240.244
R5450 gnd.n6110 gnd.n5271 240.244
R5451 gnd.n5271 gnd.n5262 240.244
R5452 gnd.n6105 gnd.n5262 240.244
R5453 gnd.n6105 gnd.n969 240.244
R5454 gnd.n6102 gnd.n969 240.244
R5455 gnd.n6102 gnd.n980 240.244
R5456 gnd.n6439 gnd.n980 240.244
R5457 gnd.n6440 gnd.n6439 240.244
R5458 gnd.n6440 gnd.n992 240.244
R5459 gnd.n6446 gnd.n992 240.244
R5460 gnd.n6446 gnd.n1003 240.244
R5461 gnd.n6450 gnd.n1003 240.244
R5462 gnd.n6450 gnd.n6449 240.244
R5463 gnd.n6449 gnd.n1018 240.244
R5464 gnd.n6457 gnd.n1018 240.244
R5465 gnd.n6457 gnd.n1028 240.244
R5466 gnd.n5667 gnd.n5665 240.244
R5467 gnd.n5665 gnd.n5664 240.244
R5468 gnd.n5661 gnd.n5660 240.244
R5469 gnd.n5658 gnd.n5584 240.244
R5470 gnd.n5654 gnd.n5652 240.244
R5471 gnd.n5650 gnd.n5590 240.244
R5472 gnd.n5646 gnd.n5644 240.244
R5473 gnd.n5642 gnd.n5596 240.244
R5474 gnd.n5638 gnd.n5636 240.244
R5475 gnd.n5634 gnd.n5602 240.244
R5476 gnd.n5630 gnd.n5628 240.244
R5477 gnd.n5626 gnd.n5608 240.244
R5478 gnd.n5621 gnd.n5619 240.244
R5479 gnd.n5673 gnd.n5569 240.244
R5480 gnd.n5683 gnd.n5569 240.244
R5481 gnd.n5683 gnd.n5565 240.244
R5482 gnd.n5689 gnd.n5565 240.244
R5483 gnd.n5689 gnd.n5557 240.244
R5484 gnd.n5699 gnd.n5557 240.244
R5485 gnd.n5699 gnd.n5553 240.244
R5486 gnd.n5705 gnd.n5553 240.244
R5487 gnd.n5705 gnd.n5544 240.244
R5488 gnd.n5797 gnd.n5544 240.244
R5489 gnd.n5797 gnd.n5539 240.244
R5490 gnd.n5804 gnd.n5539 240.244
R5491 gnd.n5804 gnd.n5530 240.244
R5492 gnd.n5814 gnd.n5530 240.244
R5493 gnd.n5814 gnd.n5516 240.244
R5494 gnd.n5829 gnd.n5516 240.244
R5495 gnd.n5829 gnd.n5509 240.244
R5496 gnd.n5844 gnd.n5509 240.244
R5497 gnd.n5844 gnd.n5510 240.244
R5498 gnd.n5510 gnd.n5488 240.244
R5499 gnd.n5868 gnd.n5488 240.244
R5500 gnd.n5868 gnd.n5489 240.244
R5501 gnd.n5489 gnd.n5469 240.244
R5502 gnd.n5895 gnd.n5469 240.244
R5503 gnd.n5895 gnd.n5456 240.244
R5504 gnd.n5915 gnd.n5456 240.244
R5505 gnd.n5915 gnd.n5457 240.244
R5506 gnd.n5911 gnd.n5457 240.244
R5507 gnd.n5911 gnd.n5437 240.244
R5508 gnd.n5953 gnd.n5437 240.244
R5509 gnd.n5953 gnd.n5430 240.244
R5510 gnd.n5964 gnd.n5430 240.244
R5511 gnd.n5964 gnd.n5423 240.244
R5512 gnd.n5979 gnd.n5423 240.244
R5513 gnd.n5979 gnd.n5424 240.244
R5514 gnd.n5424 gnd.n5402 240.244
R5515 gnd.n6001 gnd.n5402 240.244
R5516 gnd.n6001 gnd.n5403 240.244
R5517 gnd.n5403 gnd.n5318 240.244
R5518 gnd.n6038 gnd.n5318 240.244
R5519 gnd.n6038 gnd.n5311 240.244
R5520 gnd.n6049 gnd.n5311 240.244
R5521 gnd.n6049 gnd.n5304 240.244
R5522 gnd.n6063 gnd.n5304 240.244
R5523 gnd.n6063 gnd.n5305 240.244
R5524 gnd.n5305 gnd.n5285 240.244
R5525 gnd.n6087 gnd.n5285 240.244
R5526 gnd.n6087 gnd.n5275 240.244
R5527 gnd.n6112 gnd.n5275 240.244
R5528 gnd.n6112 gnd.n5261 240.244
R5529 gnd.n6138 gnd.n5261 240.244
R5530 gnd.n6138 gnd.n971 240.244
R5531 gnd.n6579 gnd.n971 240.244
R5532 gnd.n6579 gnd.n972 240.244
R5533 gnd.n6575 gnd.n972 240.244
R5534 gnd.n6575 gnd.n978 240.244
R5535 gnd.n994 gnd.n978 240.244
R5536 gnd.n6565 gnd.n994 240.244
R5537 gnd.n6565 gnd.n995 240.244
R5538 gnd.n6561 gnd.n995 240.244
R5539 gnd.n6561 gnd.n1001 240.244
R5540 gnd.n1020 gnd.n1001 240.244
R5541 gnd.n6551 gnd.n1020 240.244
R5542 gnd.n6551 gnd.n1021 240.244
R5543 gnd.n6547 gnd.n1021 240.244
R5544 gnd.n3070 gnd.n1372 240.244
R5545 gnd.n3081 gnd.n3072 240.244
R5546 gnd.n3084 gnd.n3083 240.244
R5547 gnd.n3093 gnd.n3092 240.244
R5548 gnd.n3104 gnd.n3095 240.244
R5549 gnd.n3107 gnd.n3106 240.244
R5550 gnd.n3116 gnd.n3115 240.244
R5551 gnd.n3119 gnd.n3118 240.244
R5552 gnd.n3188 gnd.n3187 240.244
R5553 gnd.n2606 gnd.n1142 240.244
R5554 gnd.n2611 gnd.n1142 240.244
R5555 gnd.n2611 gnd.n1154 240.244
R5556 gnd.n2614 gnd.n1154 240.244
R5557 gnd.n2614 gnd.n1166 240.244
R5558 gnd.n2619 gnd.n1166 240.244
R5559 gnd.n2619 gnd.n1176 240.244
R5560 gnd.n2622 gnd.n1176 240.244
R5561 gnd.n2622 gnd.n1186 240.244
R5562 gnd.n2628 gnd.n1186 240.244
R5563 gnd.n2628 gnd.n1196 240.244
R5564 gnd.n2636 gnd.n1196 240.244
R5565 gnd.n2636 gnd.n1206 240.244
R5566 gnd.n2642 gnd.n1206 240.244
R5567 gnd.n2642 gnd.n1216 240.244
R5568 gnd.n2689 gnd.n1216 240.244
R5569 gnd.n2689 gnd.n1226 240.244
R5570 gnd.n2696 gnd.n1226 240.244
R5571 gnd.n2696 gnd.n1237 240.244
R5572 gnd.n2705 gnd.n1237 240.244
R5573 gnd.n2705 gnd.n1247 240.244
R5574 gnd.n2708 gnd.n1247 240.244
R5575 gnd.n2708 gnd.n2505 240.244
R5576 gnd.n2714 gnd.n2505 240.244
R5577 gnd.n2714 gnd.n2482 240.244
R5578 gnd.n2753 gnd.n2482 240.244
R5579 gnd.n2753 gnd.n2478 240.244
R5580 gnd.n2760 gnd.n2478 240.244
R5581 gnd.n2760 gnd.n2462 240.244
R5582 gnd.n2801 gnd.n2462 240.244
R5583 gnd.n2801 gnd.n1264 240.244
R5584 gnd.n2467 gnd.n1264 240.244
R5585 gnd.n2467 gnd.n1276 240.244
R5586 gnd.n2468 gnd.n1276 240.244
R5587 gnd.n2468 gnd.n1285 240.244
R5588 gnd.n2789 gnd.n1285 240.244
R5589 gnd.n2789 gnd.n1295 240.244
R5590 gnd.n2842 gnd.n1295 240.244
R5591 gnd.n2842 gnd.n1305 240.244
R5592 gnd.n2848 gnd.n1305 240.244
R5593 gnd.n2848 gnd.n1315 240.244
R5594 gnd.n2857 gnd.n1315 240.244
R5595 gnd.n2857 gnd.n1325 240.244
R5596 gnd.n2863 gnd.n1325 240.244
R5597 gnd.n2863 gnd.n1335 240.244
R5598 gnd.n2897 gnd.n1335 240.244
R5599 gnd.n2897 gnd.n1345 240.244
R5600 gnd.n2435 gnd.n1345 240.244
R5601 gnd.n2435 gnd.n1355 240.244
R5602 gnd.n2436 gnd.n1355 240.244
R5603 gnd.n2436 gnd.n1366 240.244
R5604 gnd.n2884 gnd.n1366 240.244
R5605 gnd.n2884 gnd.n1375 240.244
R5606 gnd.n2567 gnd.n2566 240.244
R5607 gnd.n2573 gnd.n2572 240.244
R5608 gnd.n2577 gnd.n2576 240.244
R5609 gnd.n2583 gnd.n2582 240.244
R5610 gnd.n2587 gnd.n2586 240.244
R5611 gnd.n2593 gnd.n2592 240.244
R5612 gnd.n2597 gnd.n2596 240.244
R5613 gnd.n2554 gnd.n2553 240.244
R5614 gnd.n2549 gnd.n1067 240.244
R5615 gnd.n2562 gnd.n1143 240.244
R5616 gnd.n1156 gnd.n1143 240.244
R5617 gnd.n5033 gnd.n1156 240.244
R5618 gnd.n5033 gnd.n1157 240.244
R5619 gnd.n5029 gnd.n1157 240.244
R5620 gnd.n5029 gnd.n1164 240.244
R5621 gnd.n5021 gnd.n1164 240.244
R5622 gnd.n5021 gnd.n1178 240.244
R5623 gnd.n5017 gnd.n1178 240.244
R5624 gnd.n5017 gnd.n1183 240.244
R5625 gnd.n5009 gnd.n1183 240.244
R5626 gnd.n5009 gnd.n1198 240.244
R5627 gnd.n5005 gnd.n1198 240.244
R5628 gnd.n5005 gnd.n1203 240.244
R5629 gnd.n4997 gnd.n1203 240.244
R5630 gnd.n4997 gnd.n1218 240.244
R5631 gnd.n4993 gnd.n1218 240.244
R5632 gnd.n4993 gnd.n1223 240.244
R5633 gnd.n4985 gnd.n1223 240.244
R5634 gnd.n4985 gnd.n1239 240.244
R5635 gnd.n4981 gnd.n1239 240.244
R5636 gnd.n4981 gnd.n1244 240.244
R5637 gnd.n2721 gnd.n1244 240.244
R5638 gnd.n2721 gnd.n2491 240.244
R5639 gnd.n2746 gnd.n2491 240.244
R5640 gnd.n2746 gnd.n2485 240.244
R5641 gnd.n2742 gnd.n2485 240.244
R5642 gnd.n2742 gnd.n2473 240.244
R5643 gnd.n2767 gnd.n2473 240.244
R5644 gnd.n2767 gnd.n1266 240.244
R5645 gnd.n4971 gnd.n1266 240.244
R5646 gnd.n4971 gnd.n1267 240.244
R5647 gnd.n4967 gnd.n1267 240.244
R5648 gnd.n4967 gnd.n1273 240.244
R5649 gnd.n4959 gnd.n1273 240.244
R5650 gnd.n4959 gnd.n1287 240.244
R5651 gnd.n4955 gnd.n1287 240.244
R5652 gnd.n4955 gnd.n1292 240.244
R5653 gnd.n4947 gnd.n1292 240.244
R5654 gnd.n4947 gnd.n1307 240.244
R5655 gnd.n4943 gnd.n1307 240.244
R5656 gnd.n4943 gnd.n1312 240.244
R5657 gnd.n4935 gnd.n1312 240.244
R5658 gnd.n4935 gnd.n1327 240.244
R5659 gnd.n4931 gnd.n1327 240.244
R5660 gnd.n4931 gnd.n1332 240.244
R5661 gnd.n4923 gnd.n1332 240.244
R5662 gnd.n4923 gnd.n1347 240.244
R5663 gnd.n4919 gnd.n1347 240.244
R5664 gnd.n4919 gnd.n1352 240.244
R5665 gnd.n4911 gnd.n1352 240.244
R5666 gnd.n4911 gnd.n1368 240.244
R5667 gnd.n4907 gnd.n1368 240.244
R5668 gnd.n6752 gnd.n800 240.244
R5669 gnd.n6752 gnd.n796 240.244
R5670 gnd.n6758 gnd.n796 240.244
R5671 gnd.n6758 gnd.n794 240.244
R5672 gnd.n6762 gnd.n794 240.244
R5673 gnd.n6762 gnd.n790 240.244
R5674 gnd.n6768 gnd.n790 240.244
R5675 gnd.n6768 gnd.n788 240.244
R5676 gnd.n6772 gnd.n788 240.244
R5677 gnd.n6772 gnd.n784 240.244
R5678 gnd.n6778 gnd.n784 240.244
R5679 gnd.n6778 gnd.n782 240.244
R5680 gnd.n6782 gnd.n782 240.244
R5681 gnd.n6782 gnd.n778 240.244
R5682 gnd.n6788 gnd.n778 240.244
R5683 gnd.n6788 gnd.n776 240.244
R5684 gnd.n6792 gnd.n776 240.244
R5685 gnd.n6792 gnd.n772 240.244
R5686 gnd.n6798 gnd.n772 240.244
R5687 gnd.n6798 gnd.n770 240.244
R5688 gnd.n6802 gnd.n770 240.244
R5689 gnd.n6802 gnd.n766 240.244
R5690 gnd.n6808 gnd.n766 240.244
R5691 gnd.n6808 gnd.n764 240.244
R5692 gnd.n6812 gnd.n764 240.244
R5693 gnd.n6812 gnd.n760 240.244
R5694 gnd.n6818 gnd.n760 240.244
R5695 gnd.n6818 gnd.n758 240.244
R5696 gnd.n6822 gnd.n758 240.244
R5697 gnd.n6822 gnd.n754 240.244
R5698 gnd.n6828 gnd.n754 240.244
R5699 gnd.n6828 gnd.n752 240.244
R5700 gnd.n6832 gnd.n752 240.244
R5701 gnd.n6832 gnd.n748 240.244
R5702 gnd.n6838 gnd.n748 240.244
R5703 gnd.n6838 gnd.n746 240.244
R5704 gnd.n6842 gnd.n746 240.244
R5705 gnd.n6842 gnd.n742 240.244
R5706 gnd.n6848 gnd.n742 240.244
R5707 gnd.n6848 gnd.n740 240.244
R5708 gnd.n6852 gnd.n740 240.244
R5709 gnd.n6852 gnd.n736 240.244
R5710 gnd.n6858 gnd.n736 240.244
R5711 gnd.n6858 gnd.n734 240.244
R5712 gnd.n6862 gnd.n734 240.244
R5713 gnd.n6862 gnd.n730 240.244
R5714 gnd.n6868 gnd.n730 240.244
R5715 gnd.n6868 gnd.n728 240.244
R5716 gnd.n6872 gnd.n728 240.244
R5717 gnd.n6872 gnd.n724 240.244
R5718 gnd.n6878 gnd.n724 240.244
R5719 gnd.n6878 gnd.n722 240.244
R5720 gnd.n6882 gnd.n722 240.244
R5721 gnd.n6882 gnd.n718 240.244
R5722 gnd.n6888 gnd.n718 240.244
R5723 gnd.n6888 gnd.n716 240.244
R5724 gnd.n6892 gnd.n716 240.244
R5725 gnd.n6892 gnd.n712 240.244
R5726 gnd.n6898 gnd.n712 240.244
R5727 gnd.n6898 gnd.n710 240.244
R5728 gnd.n6902 gnd.n710 240.244
R5729 gnd.n6902 gnd.n706 240.244
R5730 gnd.n6908 gnd.n706 240.244
R5731 gnd.n6908 gnd.n704 240.244
R5732 gnd.n6912 gnd.n704 240.244
R5733 gnd.n6912 gnd.n700 240.244
R5734 gnd.n6918 gnd.n700 240.244
R5735 gnd.n6918 gnd.n698 240.244
R5736 gnd.n6922 gnd.n698 240.244
R5737 gnd.n6922 gnd.n694 240.244
R5738 gnd.n6928 gnd.n694 240.244
R5739 gnd.n6928 gnd.n692 240.244
R5740 gnd.n6932 gnd.n692 240.244
R5741 gnd.n6932 gnd.n688 240.244
R5742 gnd.n6938 gnd.n688 240.244
R5743 gnd.n6938 gnd.n686 240.244
R5744 gnd.n6942 gnd.n686 240.244
R5745 gnd.n6942 gnd.n682 240.244
R5746 gnd.n6948 gnd.n682 240.244
R5747 gnd.n6948 gnd.n680 240.244
R5748 gnd.n6952 gnd.n680 240.244
R5749 gnd.n6952 gnd.n676 240.244
R5750 gnd.n6958 gnd.n676 240.244
R5751 gnd.n6958 gnd.n674 240.244
R5752 gnd.n6962 gnd.n674 240.244
R5753 gnd.n6962 gnd.n670 240.244
R5754 gnd.n6968 gnd.n670 240.244
R5755 gnd.n6968 gnd.n668 240.244
R5756 gnd.n6972 gnd.n668 240.244
R5757 gnd.n6972 gnd.n664 240.244
R5758 gnd.n6978 gnd.n664 240.244
R5759 gnd.n6978 gnd.n662 240.244
R5760 gnd.n6982 gnd.n662 240.244
R5761 gnd.n6982 gnd.n658 240.244
R5762 gnd.n6988 gnd.n658 240.244
R5763 gnd.n6988 gnd.n656 240.244
R5764 gnd.n6992 gnd.n656 240.244
R5765 gnd.n6992 gnd.n652 240.244
R5766 gnd.n6998 gnd.n652 240.244
R5767 gnd.n6998 gnd.n650 240.244
R5768 gnd.n7002 gnd.n650 240.244
R5769 gnd.n7002 gnd.n646 240.244
R5770 gnd.n7008 gnd.n646 240.244
R5771 gnd.n7008 gnd.n644 240.244
R5772 gnd.n7012 gnd.n644 240.244
R5773 gnd.n7012 gnd.n640 240.244
R5774 gnd.n7018 gnd.n640 240.244
R5775 gnd.n7018 gnd.n638 240.244
R5776 gnd.n7022 gnd.n638 240.244
R5777 gnd.n7022 gnd.n634 240.244
R5778 gnd.n7028 gnd.n634 240.244
R5779 gnd.n7028 gnd.n632 240.244
R5780 gnd.n7032 gnd.n632 240.244
R5781 gnd.n7032 gnd.n628 240.244
R5782 gnd.n7038 gnd.n628 240.244
R5783 gnd.n7038 gnd.n626 240.244
R5784 gnd.n7042 gnd.n626 240.244
R5785 gnd.n7042 gnd.n622 240.244
R5786 gnd.n7048 gnd.n622 240.244
R5787 gnd.n7048 gnd.n620 240.244
R5788 gnd.n7052 gnd.n620 240.244
R5789 gnd.n7052 gnd.n616 240.244
R5790 gnd.n7058 gnd.n616 240.244
R5791 gnd.n7058 gnd.n614 240.244
R5792 gnd.n7062 gnd.n614 240.244
R5793 gnd.n7062 gnd.n610 240.244
R5794 gnd.n7068 gnd.n610 240.244
R5795 gnd.n7068 gnd.n608 240.244
R5796 gnd.n7072 gnd.n608 240.244
R5797 gnd.n7072 gnd.n604 240.244
R5798 gnd.n7078 gnd.n604 240.244
R5799 gnd.n7078 gnd.n602 240.244
R5800 gnd.n7082 gnd.n602 240.244
R5801 gnd.n7082 gnd.n598 240.244
R5802 gnd.n7088 gnd.n598 240.244
R5803 gnd.n7088 gnd.n596 240.244
R5804 gnd.n7092 gnd.n596 240.244
R5805 gnd.n7092 gnd.n592 240.244
R5806 gnd.n7098 gnd.n592 240.244
R5807 gnd.n7098 gnd.n590 240.244
R5808 gnd.n7102 gnd.n590 240.244
R5809 gnd.n7102 gnd.n586 240.244
R5810 gnd.n7108 gnd.n586 240.244
R5811 gnd.n7108 gnd.n584 240.244
R5812 gnd.n7112 gnd.n584 240.244
R5813 gnd.n7112 gnd.n580 240.244
R5814 gnd.n7118 gnd.n580 240.244
R5815 gnd.n7118 gnd.n578 240.244
R5816 gnd.n7122 gnd.n578 240.244
R5817 gnd.n7122 gnd.n574 240.244
R5818 gnd.n7128 gnd.n574 240.244
R5819 gnd.n7128 gnd.n572 240.244
R5820 gnd.n7132 gnd.n572 240.244
R5821 gnd.n7132 gnd.n568 240.244
R5822 gnd.n7138 gnd.n568 240.244
R5823 gnd.n7138 gnd.n566 240.244
R5824 gnd.n7142 gnd.n566 240.244
R5825 gnd.n7142 gnd.n562 240.244
R5826 gnd.n7148 gnd.n562 240.244
R5827 gnd.n7148 gnd.n560 240.244
R5828 gnd.n7152 gnd.n560 240.244
R5829 gnd.n7152 gnd.n556 240.244
R5830 gnd.n7158 gnd.n556 240.244
R5831 gnd.n7158 gnd.n554 240.244
R5832 gnd.n7162 gnd.n554 240.244
R5833 gnd.n7162 gnd.n550 240.244
R5834 gnd.n7168 gnd.n550 240.244
R5835 gnd.n7168 gnd.n548 240.244
R5836 gnd.n7172 gnd.n548 240.244
R5837 gnd.n7172 gnd.n544 240.244
R5838 gnd.n7178 gnd.n544 240.244
R5839 gnd.n7178 gnd.n542 240.244
R5840 gnd.n7182 gnd.n542 240.244
R5841 gnd.n7182 gnd.n538 240.244
R5842 gnd.n7188 gnd.n538 240.244
R5843 gnd.n7188 gnd.n536 240.244
R5844 gnd.n7192 gnd.n536 240.244
R5845 gnd.n7192 gnd.n532 240.244
R5846 gnd.n7198 gnd.n532 240.244
R5847 gnd.n7198 gnd.n530 240.244
R5848 gnd.n7202 gnd.n530 240.244
R5849 gnd.n7208 gnd.n526 240.244
R5850 gnd.n7208 gnd.n524 240.244
R5851 gnd.n7212 gnd.n524 240.244
R5852 gnd.n7212 gnd.n520 240.244
R5853 gnd.n7218 gnd.n520 240.244
R5854 gnd.n7218 gnd.n518 240.244
R5855 gnd.n7222 gnd.n518 240.244
R5856 gnd.n7222 gnd.n514 240.244
R5857 gnd.n7228 gnd.n514 240.244
R5858 gnd.n7228 gnd.n512 240.244
R5859 gnd.n7232 gnd.n512 240.244
R5860 gnd.n7232 gnd.n508 240.244
R5861 gnd.n7238 gnd.n508 240.244
R5862 gnd.n7238 gnd.n506 240.244
R5863 gnd.n7242 gnd.n506 240.244
R5864 gnd.n7242 gnd.n502 240.244
R5865 gnd.n7248 gnd.n502 240.244
R5866 gnd.n7248 gnd.n500 240.244
R5867 gnd.n7252 gnd.n500 240.244
R5868 gnd.n7252 gnd.n496 240.244
R5869 gnd.n7258 gnd.n496 240.244
R5870 gnd.n7258 gnd.n494 240.244
R5871 gnd.n7262 gnd.n494 240.244
R5872 gnd.n7262 gnd.n490 240.244
R5873 gnd.n7268 gnd.n490 240.244
R5874 gnd.n7268 gnd.n488 240.244
R5875 gnd.n7272 gnd.n488 240.244
R5876 gnd.n7272 gnd.n484 240.244
R5877 gnd.n7278 gnd.n484 240.244
R5878 gnd.n7278 gnd.n482 240.244
R5879 gnd.n7282 gnd.n482 240.244
R5880 gnd.n7282 gnd.n478 240.244
R5881 gnd.n7288 gnd.n478 240.244
R5882 gnd.n7288 gnd.n476 240.244
R5883 gnd.n7292 gnd.n476 240.244
R5884 gnd.n7292 gnd.n472 240.244
R5885 gnd.n7298 gnd.n472 240.244
R5886 gnd.n7298 gnd.n470 240.244
R5887 gnd.n7302 gnd.n470 240.244
R5888 gnd.n7302 gnd.n466 240.244
R5889 gnd.n7308 gnd.n466 240.244
R5890 gnd.n7308 gnd.n464 240.244
R5891 gnd.n7312 gnd.n464 240.244
R5892 gnd.n7312 gnd.n460 240.244
R5893 gnd.n7318 gnd.n460 240.244
R5894 gnd.n7318 gnd.n458 240.244
R5895 gnd.n7322 gnd.n458 240.244
R5896 gnd.n7322 gnd.n454 240.244
R5897 gnd.n7328 gnd.n454 240.244
R5898 gnd.n7328 gnd.n452 240.244
R5899 gnd.n7332 gnd.n452 240.244
R5900 gnd.n7332 gnd.n448 240.244
R5901 gnd.n7338 gnd.n448 240.244
R5902 gnd.n7338 gnd.n446 240.244
R5903 gnd.n7342 gnd.n446 240.244
R5904 gnd.n7342 gnd.n442 240.244
R5905 gnd.n7348 gnd.n442 240.244
R5906 gnd.n7348 gnd.n440 240.244
R5907 gnd.n7352 gnd.n440 240.244
R5908 gnd.n7352 gnd.n436 240.244
R5909 gnd.n7358 gnd.n436 240.244
R5910 gnd.n7358 gnd.n434 240.244
R5911 gnd.n7362 gnd.n434 240.244
R5912 gnd.n7362 gnd.n430 240.244
R5913 gnd.n7368 gnd.n430 240.244
R5914 gnd.n7368 gnd.n428 240.244
R5915 gnd.n7372 gnd.n428 240.244
R5916 gnd.n7372 gnd.n424 240.244
R5917 gnd.n7378 gnd.n424 240.244
R5918 gnd.n7378 gnd.n422 240.244
R5919 gnd.n7382 gnd.n422 240.244
R5920 gnd.n7382 gnd.n418 240.244
R5921 gnd.n7388 gnd.n418 240.244
R5922 gnd.n7388 gnd.n416 240.244
R5923 gnd.n7392 gnd.n416 240.244
R5924 gnd.n7392 gnd.n412 240.244
R5925 gnd.n7398 gnd.n412 240.244
R5926 gnd.n7398 gnd.n410 240.244
R5927 gnd.n7402 gnd.n410 240.244
R5928 gnd.n7402 gnd.n406 240.244
R5929 gnd.n7410 gnd.n406 240.244
R5930 gnd.n7410 gnd.n404 240.244
R5931 gnd.n7414 gnd.n404 240.244
R5932 gnd.n7415 gnd.n7414 240.244
R5933 gnd.n2655 gnd.n2654 240.244
R5934 gnd.n2656 gnd.n2655 240.244
R5935 gnd.n2656 gnd.n2643 240.244
R5936 gnd.n2680 gnd.n2643 240.244
R5937 gnd.n2680 gnd.n2644 240.244
R5938 gnd.n2676 gnd.n2644 240.244
R5939 gnd.n2676 gnd.n2675 240.244
R5940 gnd.n2675 gnd.n2674 240.244
R5941 gnd.n2674 gnd.n2664 240.244
R5942 gnd.n2670 gnd.n2664 240.244
R5943 gnd.n2670 gnd.n2502 240.244
R5944 gnd.n2725 gnd.n2502 240.244
R5945 gnd.n2725 gnd.n2500 240.244
R5946 gnd.n2730 gnd.n2500 240.244
R5947 gnd.n2731 gnd.n2730 240.244
R5948 gnd.n2731 gnd.n2497 240.244
R5949 gnd.n2739 gnd.n2497 240.244
R5950 gnd.n2739 gnd.n2498 240.244
R5951 gnd.n2498 gnd.n2457 240.244
R5952 gnd.n2804 gnd.n2457 240.244
R5953 gnd.n2805 gnd.n2804 240.244
R5954 gnd.n2806 gnd.n2805 240.244
R5955 gnd.n2806 gnd.n2454 240.244
R5956 gnd.n2812 gnd.n2454 240.244
R5957 gnd.n2813 gnd.n2812 240.244
R5958 gnd.n2814 gnd.n2813 240.244
R5959 gnd.n2814 gnd.n2449 240.244
R5960 gnd.n2839 gnd.n2449 240.244
R5961 gnd.n2839 gnd.n2450 240.244
R5962 gnd.n2835 gnd.n2450 240.244
R5963 gnd.n2835 gnd.n2834 240.244
R5964 gnd.n2834 gnd.n2833 240.244
R5965 gnd.n2833 gnd.n2822 240.244
R5966 gnd.n2829 gnd.n2822 240.244
R5967 gnd.n2829 gnd.n2429 240.244
R5968 gnd.n2900 gnd.n2429 240.244
R5969 gnd.n2901 gnd.n2900 240.244
R5970 gnd.n2901 gnd.n2425 240.244
R5971 gnd.n2907 gnd.n2425 240.244
R5972 gnd.n2908 gnd.n2907 240.244
R5973 gnd.n2909 gnd.n2908 240.244
R5974 gnd.n2909 gnd.n2421 240.244
R5975 gnd.n2915 gnd.n2421 240.244
R5976 gnd.n2917 gnd.n2915 240.244
R5977 gnd.n2919 gnd.n2917 240.244
R5978 gnd.n2919 gnd.n2417 240.244
R5979 gnd.n2925 gnd.n2417 240.244
R5980 gnd.n2925 gnd.n2396 240.244
R5981 gnd.n3203 gnd.n2396 240.244
R5982 gnd.n3203 gnd.n2391 240.244
R5983 gnd.n3211 gnd.n2391 240.244
R5984 gnd.n3211 gnd.n2392 240.244
R5985 gnd.n2392 gnd.n2371 240.244
R5986 gnd.n3235 gnd.n2371 240.244
R5987 gnd.n3235 gnd.n2366 240.244
R5988 gnd.n3244 gnd.n2366 240.244
R5989 gnd.n3244 gnd.n2367 240.244
R5990 gnd.n2367 gnd.n1494 240.244
R5991 gnd.n4779 gnd.n1494 240.244
R5992 gnd.n4779 gnd.n1495 240.244
R5993 gnd.n4775 gnd.n1495 240.244
R5994 gnd.n4775 gnd.n1501 240.244
R5995 gnd.n3280 gnd.n1501 240.244
R5996 gnd.n3280 gnd.n2245 240.244
R5997 gnd.n3317 gnd.n2245 240.244
R5998 gnd.n3317 gnd.n2241 240.244
R5999 gnd.n3323 gnd.n2241 240.244
R6000 gnd.n3323 gnd.n2227 240.244
R6001 gnd.n3359 gnd.n2227 240.244
R6002 gnd.n3359 gnd.n2222 240.244
R6003 gnd.n3367 gnd.n2222 240.244
R6004 gnd.n3367 gnd.n2223 240.244
R6005 gnd.n2223 gnd.n2201 240.244
R6006 gnd.n3421 gnd.n2201 240.244
R6007 gnd.n3421 gnd.n2197 240.244
R6008 gnd.n3427 gnd.n2197 240.244
R6009 gnd.n3427 gnd.n2183 240.244
R6010 gnd.n3449 gnd.n2183 240.244
R6011 gnd.n3449 gnd.n2178 240.244
R6012 gnd.n3457 gnd.n2178 240.244
R6013 gnd.n3457 gnd.n2179 240.244
R6014 gnd.n2179 gnd.n2150 240.244
R6015 gnd.n3499 gnd.n2150 240.244
R6016 gnd.n3499 gnd.n2146 240.244
R6017 gnd.n3505 gnd.n2146 240.244
R6018 gnd.n3505 gnd.n2127 240.244
R6019 gnd.n3539 gnd.n2127 240.244
R6020 gnd.n3539 gnd.n2123 240.244
R6021 gnd.n3545 gnd.n2123 240.244
R6022 gnd.n3545 gnd.n2105 240.244
R6023 gnd.n3596 gnd.n2105 240.244
R6024 gnd.n3596 gnd.n2101 240.244
R6025 gnd.n3602 gnd.n2101 240.244
R6026 gnd.n3602 gnd.n2085 240.244
R6027 gnd.n3621 gnd.n2085 240.244
R6028 gnd.n3621 gnd.n2081 240.244
R6029 gnd.n3627 gnd.n2081 240.244
R6030 gnd.n3627 gnd.n2065 240.244
R6031 gnd.n3681 gnd.n2065 240.244
R6032 gnd.n3681 gnd.n2061 240.244
R6033 gnd.n3687 gnd.n2061 240.244
R6034 gnd.n3687 gnd.n2043 240.244
R6035 gnd.n3710 gnd.n2043 240.244
R6036 gnd.n3710 gnd.n2038 240.244
R6037 gnd.n3718 gnd.n2038 240.244
R6038 gnd.n3718 gnd.n2039 240.244
R6039 gnd.n2039 gnd.n2015 240.244
R6040 gnd.n3761 gnd.n2015 240.244
R6041 gnd.n3761 gnd.n2011 240.244
R6042 gnd.n3767 gnd.n2011 240.244
R6043 gnd.n3767 gnd.n1995 240.244
R6044 gnd.n3787 gnd.n1995 240.244
R6045 gnd.n3787 gnd.n1990 240.244
R6046 gnd.n3795 gnd.n1990 240.244
R6047 gnd.n3795 gnd.n1991 240.244
R6048 gnd.n1991 gnd.n1965 240.244
R6049 gnd.n3831 gnd.n1965 240.244
R6050 gnd.n3831 gnd.n1959 240.244
R6051 gnd.n3840 gnd.n1959 240.244
R6052 gnd.n3840 gnd.n1961 240.244
R6053 gnd.n1961 gnd.n1911 240.244
R6054 gnd.n4086 gnd.n1911 240.244
R6055 gnd.n4086 gnd.n1912 240.244
R6056 gnd.n4082 gnd.n1912 240.244
R6057 gnd.n4082 gnd.n4081 240.244
R6058 gnd.n4081 gnd.n1918 240.244
R6059 gnd.n4074 gnd.n1918 240.244
R6060 gnd.n4074 gnd.n1923 240.244
R6061 gnd.n4070 gnd.n1923 240.244
R6062 gnd.n4070 gnd.n1933 240.244
R6063 gnd.n1933 gnd.n1601 240.244
R6064 gnd.n4661 gnd.n1601 240.244
R6065 gnd.n4661 gnd.n1602 240.244
R6066 gnd.n4657 gnd.n1602 240.244
R6067 gnd.n4657 gnd.n1608 240.244
R6068 gnd.n4653 gnd.n1608 240.244
R6069 gnd.n4653 gnd.n1611 240.244
R6070 gnd.n4649 gnd.n1611 240.244
R6071 gnd.n4649 gnd.n1617 240.244
R6072 gnd.n1793 gnd.n1617 240.244
R6073 gnd.n1799 gnd.n1793 240.244
R6074 gnd.n1800 gnd.n1799 240.244
R6075 gnd.n1801 gnd.n1800 240.244
R6076 gnd.n1801 gnd.n1788 240.244
R6077 gnd.n1818 gnd.n1788 240.244
R6078 gnd.n1818 gnd.n1789 240.244
R6079 gnd.n1814 gnd.n1789 240.244
R6080 gnd.n1814 gnd.n1813 240.244
R6081 gnd.n1813 gnd.n1772 240.244
R6082 gnd.n4494 gnd.n1772 240.244
R6083 gnd.n4495 gnd.n4494 240.244
R6084 gnd.n4496 gnd.n4495 240.244
R6085 gnd.n4496 gnd.n1768 240.244
R6086 gnd.n4502 gnd.n1768 240.244
R6087 gnd.n4503 gnd.n4502 240.244
R6088 gnd.n4504 gnd.n4503 240.244
R6089 gnd.n4504 gnd.n1763 240.244
R6090 gnd.n4514 gnd.n1763 240.244
R6091 gnd.n4514 gnd.n1764 240.244
R6092 gnd.n1764 gnd.n1755 240.244
R6093 gnd.n4559 gnd.n1755 240.244
R6094 gnd.n4560 gnd.n4559 240.244
R6095 gnd.n4560 gnd.n1752 240.244
R6096 gnd.n4570 gnd.n1752 240.244
R6097 gnd.n4570 gnd.n1753 240.244
R6098 gnd.n4565 gnd.n1753 240.244
R6099 gnd.n4565 gnd.n382 240.244
R6100 gnd.n7440 gnd.n382 240.244
R6101 gnd.n7440 gnd.n383 240.244
R6102 gnd.n7435 gnd.n383 240.244
R6103 gnd.n7435 gnd.n7434 240.244
R6104 gnd.n7434 gnd.n7433 240.244
R6105 gnd.n7433 gnd.n387 240.244
R6106 gnd.n7429 gnd.n387 240.244
R6107 gnd.n7429 gnd.n7428 240.244
R6108 gnd.n7428 gnd.n7427 240.244
R6109 gnd.n7427 gnd.n393 240.244
R6110 gnd.n7423 gnd.n393 240.244
R6111 gnd.n7423 gnd.n7422 240.244
R6112 gnd.n7422 gnd.n7421 240.244
R6113 gnd.n7421 gnd.n399 240.244
R6114 gnd.n6748 gnd.n802 240.244
R6115 gnd.n6744 gnd.n802 240.244
R6116 gnd.n6744 gnd.n807 240.244
R6117 gnd.n6740 gnd.n807 240.244
R6118 gnd.n6740 gnd.n809 240.244
R6119 gnd.n6736 gnd.n809 240.244
R6120 gnd.n6736 gnd.n815 240.244
R6121 gnd.n6732 gnd.n815 240.244
R6122 gnd.n6732 gnd.n817 240.244
R6123 gnd.n6728 gnd.n817 240.244
R6124 gnd.n6728 gnd.n823 240.244
R6125 gnd.n6724 gnd.n823 240.244
R6126 gnd.n6724 gnd.n825 240.244
R6127 gnd.n6720 gnd.n825 240.244
R6128 gnd.n6720 gnd.n831 240.244
R6129 gnd.n6716 gnd.n831 240.244
R6130 gnd.n6716 gnd.n833 240.244
R6131 gnd.n6712 gnd.n833 240.244
R6132 gnd.n6712 gnd.n839 240.244
R6133 gnd.n6708 gnd.n839 240.244
R6134 gnd.n6708 gnd.n841 240.244
R6135 gnd.n6704 gnd.n841 240.244
R6136 gnd.n6704 gnd.n847 240.244
R6137 gnd.n6700 gnd.n847 240.244
R6138 gnd.n6700 gnd.n849 240.244
R6139 gnd.n6696 gnd.n849 240.244
R6140 gnd.n6696 gnd.n855 240.244
R6141 gnd.n6692 gnd.n855 240.244
R6142 gnd.n6692 gnd.n857 240.244
R6143 gnd.n6688 gnd.n857 240.244
R6144 gnd.n6688 gnd.n863 240.244
R6145 gnd.n6684 gnd.n863 240.244
R6146 gnd.n6684 gnd.n865 240.244
R6147 gnd.n6680 gnd.n865 240.244
R6148 gnd.n6680 gnd.n871 240.244
R6149 gnd.n6676 gnd.n871 240.244
R6150 gnd.n6676 gnd.n873 240.244
R6151 gnd.n6672 gnd.n873 240.244
R6152 gnd.n6672 gnd.n879 240.244
R6153 gnd.n6668 gnd.n879 240.244
R6154 gnd.n6668 gnd.n881 240.244
R6155 gnd.n6664 gnd.n881 240.244
R6156 gnd.n6664 gnd.n887 240.244
R6157 gnd.n6660 gnd.n887 240.244
R6158 gnd.n6660 gnd.n889 240.244
R6159 gnd.n6656 gnd.n889 240.244
R6160 gnd.n6656 gnd.n895 240.244
R6161 gnd.n6652 gnd.n895 240.244
R6162 gnd.n6652 gnd.n897 240.244
R6163 gnd.n6648 gnd.n897 240.244
R6164 gnd.n6648 gnd.n903 240.244
R6165 gnd.n6644 gnd.n903 240.244
R6166 gnd.n6644 gnd.n905 240.244
R6167 gnd.n6640 gnd.n905 240.244
R6168 gnd.n6640 gnd.n911 240.244
R6169 gnd.n6636 gnd.n911 240.244
R6170 gnd.n6636 gnd.n913 240.244
R6171 gnd.n6632 gnd.n913 240.244
R6172 gnd.n6632 gnd.n919 240.244
R6173 gnd.n6628 gnd.n919 240.244
R6174 gnd.n6628 gnd.n921 240.244
R6175 gnd.n6624 gnd.n921 240.244
R6176 gnd.n6624 gnd.n927 240.244
R6177 gnd.n6620 gnd.n927 240.244
R6178 gnd.n6620 gnd.n929 240.244
R6179 gnd.n6616 gnd.n929 240.244
R6180 gnd.n6616 gnd.n935 240.244
R6181 gnd.n6612 gnd.n935 240.244
R6182 gnd.n6612 gnd.n937 240.244
R6183 gnd.n6608 gnd.n937 240.244
R6184 gnd.n6608 gnd.n943 240.244
R6185 gnd.n6604 gnd.n943 240.244
R6186 gnd.n6604 gnd.n945 240.244
R6187 gnd.n6600 gnd.n945 240.244
R6188 gnd.n6600 gnd.n951 240.244
R6189 gnd.n6596 gnd.n951 240.244
R6190 gnd.n6596 gnd.n953 240.244
R6191 gnd.n6592 gnd.n953 240.244
R6192 gnd.n6592 gnd.n959 240.244
R6193 gnd.n6588 gnd.n959 240.244
R6194 gnd.n6588 gnd.n961 240.244
R6195 gnd.n6584 gnd.n961 240.244
R6196 gnd.n6584 gnd.n967 240.244
R6197 gnd.n2648 gnd.n967 240.244
R6198 gnd.n3214 gnd.n2387 240.244
R6199 gnd.n3214 gnd.n2381 240.244
R6200 gnd.n3221 gnd.n2381 240.244
R6201 gnd.n3221 gnd.n2382 240.244
R6202 gnd.n2382 gnd.n2363 240.244
R6203 gnd.n3247 gnd.n2363 240.244
R6204 gnd.n3247 gnd.n2357 240.244
R6205 gnd.n3257 gnd.n2357 240.244
R6206 gnd.n3257 gnd.n2358 240.244
R6207 gnd.n3251 gnd.n2358 240.244
R6208 gnd.n3251 gnd.n1505 240.244
R6209 gnd.n4772 gnd.n1505 240.244
R6210 gnd.n4772 gnd.n1506 240.244
R6211 gnd.n1511 gnd.n1506 240.244
R6212 gnd.n1512 gnd.n1511 240.244
R6213 gnd.n1513 gnd.n1512 240.244
R6214 gnd.n2239 gnd.n1513 240.244
R6215 gnd.n2239 gnd.n1516 240.244
R6216 gnd.n1517 gnd.n1516 240.244
R6217 gnd.n1518 gnd.n1517 240.244
R6218 gnd.n3369 gnd.n1518 240.244
R6219 gnd.n3369 gnd.n1521 240.244
R6220 gnd.n1522 gnd.n1521 240.244
R6221 gnd.n1523 gnd.n1522 240.244
R6222 gnd.n3418 gnd.n1523 240.244
R6223 gnd.n3418 gnd.n1526 240.244
R6224 gnd.n1527 gnd.n1526 240.244
R6225 gnd.n1528 gnd.n1527 240.244
R6226 gnd.n3446 gnd.n1528 240.244
R6227 gnd.n3446 gnd.n1531 240.244
R6228 gnd.n1532 gnd.n1531 240.244
R6229 gnd.n1533 gnd.n1532 240.244
R6230 gnd.n3471 gnd.n1533 240.244
R6231 gnd.n3471 gnd.n1536 240.244
R6232 gnd.n1537 gnd.n1536 240.244
R6233 gnd.n1538 gnd.n1537 240.244
R6234 gnd.n3526 gnd.n1538 240.244
R6235 gnd.n3526 gnd.n1541 240.244
R6236 gnd.n1542 gnd.n1541 240.244
R6237 gnd.n1543 gnd.n1542 240.244
R6238 gnd.n3585 gnd.n1543 240.244
R6239 gnd.n3585 gnd.n1546 240.244
R6240 gnd.n1547 gnd.n1546 240.244
R6241 gnd.n1548 gnd.n1547 240.244
R6242 gnd.n2092 gnd.n1548 240.244
R6243 gnd.n2092 gnd.n1551 240.244
R6244 gnd.n1552 gnd.n1551 240.244
R6245 gnd.n1553 gnd.n1552 240.244
R6246 gnd.n3567 gnd.n1553 240.244
R6247 gnd.n3567 gnd.n1556 240.244
R6248 gnd.n1557 gnd.n1556 240.244
R6249 gnd.n1558 gnd.n1557 240.244
R6250 gnd.n3698 gnd.n1558 240.244
R6251 gnd.n3698 gnd.n1561 240.244
R6252 gnd.n1562 gnd.n1561 240.244
R6253 gnd.n1563 gnd.n1562 240.244
R6254 gnd.n3658 gnd.n1563 240.244
R6255 gnd.n3658 gnd.n1566 240.244
R6256 gnd.n1567 gnd.n1566 240.244
R6257 gnd.n1568 gnd.n1567 240.244
R6258 gnd.n2009 gnd.n1568 240.244
R6259 gnd.n2009 gnd.n1571 240.244
R6260 gnd.n1572 gnd.n1571 240.244
R6261 gnd.n1573 gnd.n1572 240.244
R6262 gnd.n1981 gnd.n1573 240.244
R6263 gnd.n1981 gnd.n1576 240.244
R6264 gnd.n1577 gnd.n1576 240.244
R6265 gnd.n1578 gnd.n1577 240.244
R6266 gnd.n3843 gnd.n1578 240.244
R6267 gnd.n3843 gnd.n1581 240.244
R6268 gnd.n1582 gnd.n1581 240.244
R6269 gnd.n1583 gnd.n1582 240.244
R6270 gnd.n3868 gnd.n1583 240.244
R6271 gnd.n3868 gnd.n1586 240.244
R6272 gnd.n1587 gnd.n1586 240.244
R6273 gnd.n1588 gnd.n1587 240.244
R6274 gnd.n4076 gnd.n1588 240.244
R6275 gnd.n4076 gnd.n1591 240.244
R6276 gnd.n1592 gnd.n1591 240.244
R6277 gnd.n1593 gnd.n1592 240.244
R6278 gnd.n1596 gnd.n1593 240.244
R6279 gnd.n4664 gnd.n1596 240.244
R6280 gnd.n2940 gnd.n2939 240.244
R6281 gnd.n2944 gnd.n2939 240.244
R6282 gnd.n2946 gnd.n2945 240.244
R6283 gnd.n3063 gnd.n3062 240.244
R6284 gnd.n3065 gnd.n3064 240.244
R6285 gnd.n3076 gnd.n3075 240.244
R6286 gnd.n3078 gnd.n3077 240.244
R6287 gnd.n3088 gnd.n3087 240.244
R6288 gnd.n3099 gnd.n3098 240.244
R6289 gnd.n3101 gnd.n3100 240.244
R6290 gnd.n3111 gnd.n3110 240.244
R6291 gnd.n3122 gnd.n3121 240.244
R6292 gnd.n3182 gnd.n2414 240.244
R6293 gnd.n2415 gnd.n2402 240.244
R6294 gnd.n3200 gnd.n2389 240.244
R6295 gnd.n2389 gnd.n2378 240.244
R6296 gnd.n3223 gnd.n2378 240.244
R6297 gnd.n3223 gnd.n2373 240.244
R6298 gnd.n3232 gnd.n2373 240.244
R6299 gnd.n3232 gnd.n2365 240.244
R6300 gnd.n2365 gnd.n2277 240.244
R6301 gnd.n3259 gnd.n2277 240.244
R6302 gnd.n3260 gnd.n3259 240.244
R6303 gnd.n3260 gnd.n2272 240.244
R6304 gnd.n3267 gnd.n2272 240.244
R6305 gnd.n3267 gnd.n1503 240.244
R6306 gnd.n3284 gnd.n1503 240.244
R6307 gnd.n3285 gnd.n3284 240.244
R6308 gnd.n3285 gnd.n2260 240.244
R6309 gnd.n3298 gnd.n2260 240.244
R6310 gnd.n3298 gnd.n2261 240.244
R6311 gnd.n3290 gnd.n2261 240.244
R6312 gnd.n3291 gnd.n3290 240.244
R6313 gnd.n3291 gnd.n2219 240.244
R6314 gnd.n3371 gnd.n2219 240.244
R6315 gnd.n3371 gnd.n2214 240.244
R6316 gnd.n3396 gnd.n2214 240.244
R6317 gnd.n3396 gnd.n2210 240.244
R6318 gnd.n2210 gnd.n2202 240.244
R6319 gnd.n3376 gnd.n2202 240.244
R6320 gnd.n3379 gnd.n3376 240.244
R6321 gnd.n3380 gnd.n3379 240.244
R6322 gnd.n3380 gnd.n2185 240.244
R6323 gnd.n2185 gnd.n2167 240.244
R6324 gnd.n3469 gnd.n2167 240.244
R6325 gnd.n3470 gnd.n3469 240.244
R6326 gnd.n3473 gnd.n3470 240.244
R6327 gnd.n3473 gnd.n2163 240.244
R6328 gnd.n3479 gnd.n2163 240.244
R6329 gnd.n3479 gnd.n2137 240.244
R6330 gnd.n3525 gnd.n2137 240.244
R6331 gnd.n3525 gnd.n2138 240.244
R6332 gnd.n3519 gnd.n2138 240.244
R6333 gnd.n3519 gnd.n2115 240.244
R6334 gnd.n3584 gnd.n2115 240.244
R6335 gnd.n3584 gnd.n2107 240.244
R6336 gnd.n3560 gnd.n2107 240.244
R6337 gnd.n3561 gnd.n3560 240.244
R6338 gnd.n3562 gnd.n3561 240.244
R6339 gnd.n3562 gnd.n2087 240.244
R6340 gnd.n2087 gnd.n2080 240.244
R6341 gnd.n3565 gnd.n2080 240.244
R6342 gnd.n3569 gnd.n3565 240.244
R6343 gnd.n3569 gnd.n2058 240.244
R6344 gnd.n3690 gnd.n2058 240.244
R6345 gnd.n3690 gnd.n2052 240.244
R6346 gnd.n3697 gnd.n2052 240.244
R6347 gnd.n3697 gnd.n2053 240.244
R6348 gnd.n2053 gnd.n2029 240.244
R6349 gnd.n3729 gnd.n2029 240.244
R6350 gnd.n3729 gnd.n2024 240.244
R6351 gnd.n3750 gnd.n2024 240.244
R6352 gnd.n3750 gnd.n2017 240.244
R6353 gnd.n3734 gnd.n2017 240.244
R6354 gnd.n3735 gnd.n3734 240.244
R6355 gnd.n3737 gnd.n3735 240.244
R6356 gnd.n3737 gnd.n1997 240.244
R6357 gnd.n1997 gnd.n1989 240.244
R6358 gnd.n1989 gnd.n1973 240.244
R6359 gnd.n3820 gnd.n1973 240.244
R6360 gnd.n3820 gnd.n1968 240.244
R6361 gnd.n3827 gnd.n1968 240.244
R6362 gnd.n3827 gnd.n1958 240.244
R6363 gnd.n1958 gnd.n1946 240.244
R6364 gnd.n3862 gnd.n1946 240.244
R6365 gnd.n3862 gnd.n1909 240.244
R6366 gnd.n3870 gnd.n1909 240.244
R6367 gnd.n3872 gnd.n3870 240.244
R6368 gnd.n3873 gnd.n3872 240.244
R6369 gnd.n3873 gnd.n1920 240.244
R6370 gnd.n1921 gnd.n1920 240.244
R6371 gnd.n3880 gnd.n1921 240.244
R6372 gnd.n3881 gnd.n3880 240.244
R6373 gnd.n3881 gnd.n1936 240.244
R6374 gnd.n4065 gnd.n1936 240.244
R6375 gnd.n4065 gnd.n1599 240.244
R6376 gnd.n3952 gnd.n3951 240.244
R6377 gnd.n3955 gnd.n3954 240.244
R6378 gnd.n3963 gnd.n3962 240.244
R6379 gnd.n3966 gnd.n3965 240.244
R6380 gnd.n3978 gnd.n3977 240.244
R6381 gnd.n3981 gnd.n3980 240.244
R6382 gnd.n3997 gnd.n3996 240.244
R6383 gnd.n4000 gnd.n3999 240.244
R6384 gnd.n4016 gnd.n4015 240.244
R6385 gnd.n4019 gnd.n4018 240.244
R6386 gnd.n4035 gnd.n4034 240.244
R6387 gnd.n4037 gnd.n3894 240.244
R6388 gnd.n4054 gnd.n3894 240.244
R6389 gnd.n4057 gnd.n4056 240.244
R6390 gnd.n1475 gnd.n1474 240.132
R6391 gnd.n4104 gnd.n4103 240.132
R6392 gnd.n6751 gnd.n6750 225.874
R6393 gnd.n6751 gnd.n795 225.874
R6394 gnd.n6759 gnd.n795 225.874
R6395 gnd.n6760 gnd.n6759 225.874
R6396 gnd.n6761 gnd.n6760 225.874
R6397 gnd.n6761 gnd.n789 225.874
R6398 gnd.n6769 gnd.n789 225.874
R6399 gnd.n6770 gnd.n6769 225.874
R6400 gnd.n6771 gnd.n6770 225.874
R6401 gnd.n6771 gnd.n783 225.874
R6402 gnd.n6779 gnd.n783 225.874
R6403 gnd.n6780 gnd.n6779 225.874
R6404 gnd.n6781 gnd.n6780 225.874
R6405 gnd.n6781 gnd.n777 225.874
R6406 gnd.n6789 gnd.n777 225.874
R6407 gnd.n6790 gnd.n6789 225.874
R6408 gnd.n6791 gnd.n6790 225.874
R6409 gnd.n6791 gnd.n771 225.874
R6410 gnd.n6799 gnd.n771 225.874
R6411 gnd.n6800 gnd.n6799 225.874
R6412 gnd.n6801 gnd.n6800 225.874
R6413 gnd.n6801 gnd.n765 225.874
R6414 gnd.n6809 gnd.n765 225.874
R6415 gnd.n6810 gnd.n6809 225.874
R6416 gnd.n6811 gnd.n6810 225.874
R6417 gnd.n6811 gnd.n759 225.874
R6418 gnd.n6819 gnd.n759 225.874
R6419 gnd.n6820 gnd.n6819 225.874
R6420 gnd.n6821 gnd.n6820 225.874
R6421 gnd.n6821 gnd.n753 225.874
R6422 gnd.n6829 gnd.n753 225.874
R6423 gnd.n6830 gnd.n6829 225.874
R6424 gnd.n6831 gnd.n6830 225.874
R6425 gnd.n6831 gnd.n747 225.874
R6426 gnd.n6839 gnd.n747 225.874
R6427 gnd.n6840 gnd.n6839 225.874
R6428 gnd.n6841 gnd.n6840 225.874
R6429 gnd.n6841 gnd.n741 225.874
R6430 gnd.n6849 gnd.n741 225.874
R6431 gnd.n6850 gnd.n6849 225.874
R6432 gnd.n6851 gnd.n6850 225.874
R6433 gnd.n6851 gnd.n735 225.874
R6434 gnd.n6859 gnd.n735 225.874
R6435 gnd.n6860 gnd.n6859 225.874
R6436 gnd.n6861 gnd.n6860 225.874
R6437 gnd.n6861 gnd.n729 225.874
R6438 gnd.n6869 gnd.n729 225.874
R6439 gnd.n6870 gnd.n6869 225.874
R6440 gnd.n6871 gnd.n6870 225.874
R6441 gnd.n6871 gnd.n723 225.874
R6442 gnd.n6879 gnd.n723 225.874
R6443 gnd.n6880 gnd.n6879 225.874
R6444 gnd.n6881 gnd.n6880 225.874
R6445 gnd.n6881 gnd.n717 225.874
R6446 gnd.n6889 gnd.n717 225.874
R6447 gnd.n6890 gnd.n6889 225.874
R6448 gnd.n6891 gnd.n6890 225.874
R6449 gnd.n6891 gnd.n711 225.874
R6450 gnd.n6899 gnd.n711 225.874
R6451 gnd.n6900 gnd.n6899 225.874
R6452 gnd.n6901 gnd.n6900 225.874
R6453 gnd.n6901 gnd.n705 225.874
R6454 gnd.n6909 gnd.n705 225.874
R6455 gnd.n6910 gnd.n6909 225.874
R6456 gnd.n6911 gnd.n6910 225.874
R6457 gnd.n6911 gnd.n699 225.874
R6458 gnd.n6919 gnd.n699 225.874
R6459 gnd.n6920 gnd.n6919 225.874
R6460 gnd.n6921 gnd.n6920 225.874
R6461 gnd.n6921 gnd.n693 225.874
R6462 gnd.n6929 gnd.n693 225.874
R6463 gnd.n6930 gnd.n6929 225.874
R6464 gnd.n6931 gnd.n6930 225.874
R6465 gnd.n6931 gnd.n687 225.874
R6466 gnd.n6939 gnd.n687 225.874
R6467 gnd.n6940 gnd.n6939 225.874
R6468 gnd.n6941 gnd.n6940 225.874
R6469 gnd.n6941 gnd.n681 225.874
R6470 gnd.n6949 gnd.n681 225.874
R6471 gnd.n6950 gnd.n6949 225.874
R6472 gnd.n6951 gnd.n6950 225.874
R6473 gnd.n6951 gnd.n675 225.874
R6474 gnd.n6959 gnd.n675 225.874
R6475 gnd.n6960 gnd.n6959 225.874
R6476 gnd.n6961 gnd.n6960 225.874
R6477 gnd.n6961 gnd.n669 225.874
R6478 gnd.n6969 gnd.n669 225.874
R6479 gnd.n6970 gnd.n6969 225.874
R6480 gnd.n6971 gnd.n6970 225.874
R6481 gnd.n6971 gnd.n663 225.874
R6482 gnd.n6979 gnd.n663 225.874
R6483 gnd.n6980 gnd.n6979 225.874
R6484 gnd.n6981 gnd.n6980 225.874
R6485 gnd.n6981 gnd.n657 225.874
R6486 gnd.n6989 gnd.n657 225.874
R6487 gnd.n6990 gnd.n6989 225.874
R6488 gnd.n6991 gnd.n6990 225.874
R6489 gnd.n6991 gnd.n651 225.874
R6490 gnd.n6999 gnd.n651 225.874
R6491 gnd.n7000 gnd.n6999 225.874
R6492 gnd.n7001 gnd.n7000 225.874
R6493 gnd.n7001 gnd.n645 225.874
R6494 gnd.n7009 gnd.n645 225.874
R6495 gnd.n7010 gnd.n7009 225.874
R6496 gnd.n7011 gnd.n7010 225.874
R6497 gnd.n7011 gnd.n639 225.874
R6498 gnd.n7019 gnd.n639 225.874
R6499 gnd.n7020 gnd.n7019 225.874
R6500 gnd.n7021 gnd.n7020 225.874
R6501 gnd.n7021 gnd.n633 225.874
R6502 gnd.n7029 gnd.n633 225.874
R6503 gnd.n7030 gnd.n7029 225.874
R6504 gnd.n7031 gnd.n7030 225.874
R6505 gnd.n7031 gnd.n627 225.874
R6506 gnd.n7039 gnd.n627 225.874
R6507 gnd.n7040 gnd.n7039 225.874
R6508 gnd.n7041 gnd.n7040 225.874
R6509 gnd.n7041 gnd.n621 225.874
R6510 gnd.n7049 gnd.n621 225.874
R6511 gnd.n7050 gnd.n7049 225.874
R6512 gnd.n7051 gnd.n7050 225.874
R6513 gnd.n7051 gnd.n615 225.874
R6514 gnd.n7059 gnd.n615 225.874
R6515 gnd.n7060 gnd.n7059 225.874
R6516 gnd.n7061 gnd.n7060 225.874
R6517 gnd.n7061 gnd.n609 225.874
R6518 gnd.n7069 gnd.n609 225.874
R6519 gnd.n7070 gnd.n7069 225.874
R6520 gnd.n7071 gnd.n7070 225.874
R6521 gnd.n7071 gnd.n603 225.874
R6522 gnd.n7079 gnd.n603 225.874
R6523 gnd.n7080 gnd.n7079 225.874
R6524 gnd.n7081 gnd.n7080 225.874
R6525 gnd.n7081 gnd.n597 225.874
R6526 gnd.n7089 gnd.n597 225.874
R6527 gnd.n7090 gnd.n7089 225.874
R6528 gnd.n7091 gnd.n7090 225.874
R6529 gnd.n7091 gnd.n591 225.874
R6530 gnd.n7099 gnd.n591 225.874
R6531 gnd.n7100 gnd.n7099 225.874
R6532 gnd.n7101 gnd.n7100 225.874
R6533 gnd.n7101 gnd.n585 225.874
R6534 gnd.n7109 gnd.n585 225.874
R6535 gnd.n7110 gnd.n7109 225.874
R6536 gnd.n7111 gnd.n7110 225.874
R6537 gnd.n7111 gnd.n579 225.874
R6538 gnd.n7119 gnd.n579 225.874
R6539 gnd.n7120 gnd.n7119 225.874
R6540 gnd.n7121 gnd.n7120 225.874
R6541 gnd.n7121 gnd.n573 225.874
R6542 gnd.n7129 gnd.n573 225.874
R6543 gnd.n7130 gnd.n7129 225.874
R6544 gnd.n7131 gnd.n7130 225.874
R6545 gnd.n7131 gnd.n567 225.874
R6546 gnd.n7139 gnd.n567 225.874
R6547 gnd.n7140 gnd.n7139 225.874
R6548 gnd.n7141 gnd.n7140 225.874
R6549 gnd.n7141 gnd.n561 225.874
R6550 gnd.n7149 gnd.n561 225.874
R6551 gnd.n7150 gnd.n7149 225.874
R6552 gnd.n7151 gnd.n7150 225.874
R6553 gnd.n7151 gnd.n555 225.874
R6554 gnd.n7159 gnd.n555 225.874
R6555 gnd.n7160 gnd.n7159 225.874
R6556 gnd.n7161 gnd.n7160 225.874
R6557 gnd.n7161 gnd.n549 225.874
R6558 gnd.n7169 gnd.n549 225.874
R6559 gnd.n7170 gnd.n7169 225.874
R6560 gnd.n7171 gnd.n7170 225.874
R6561 gnd.n7171 gnd.n543 225.874
R6562 gnd.n7179 gnd.n543 225.874
R6563 gnd.n7180 gnd.n7179 225.874
R6564 gnd.n7181 gnd.n7180 225.874
R6565 gnd.n7181 gnd.n537 225.874
R6566 gnd.n7189 gnd.n537 225.874
R6567 gnd.n7190 gnd.n7189 225.874
R6568 gnd.n7191 gnd.n7190 225.874
R6569 gnd.n7191 gnd.n531 225.874
R6570 gnd.n7199 gnd.n531 225.874
R6571 gnd.n7200 gnd.n7199 225.874
R6572 gnd.n7201 gnd.n7200 225.874
R6573 gnd.n5611 gnd.t211 224.174
R6574 gnd.n5239 gnd.t206 224.174
R6575 gnd.n4345 gnd.n4344 199.319
R6576 gnd.n4346 gnd.n4345 199.319
R6577 gnd.n1427 gnd.n1426 199.319
R6578 gnd.n2983 gnd.n1427 199.319
R6579 gnd.n1476 gnd.n1473 186.49
R6580 gnd.n4105 gnd.n4102 186.49
R6581 gnd.n6407 gnd.n6406 185
R6582 gnd.n6405 gnd.n6404 185
R6583 gnd.n6384 gnd.n6383 185
R6584 gnd.n6399 gnd.n6398 185
R6585 gnd.n6397 gnd.n6396 185
R6586 gnd.n6388 gnd.n6387 185
R6587 gnd.n6391 gnd.n6390 185
R6588 gnd.n6375 gnd.n6374 185
R6589 gnd.n6373 gnd.n6372 185
R6590 gnd.n6352 gnd.n6351 185
R6591 gnd.n6367 gnd.n6366 185
R6592 gnd.n6365 gnd.n6364 185
R6593 gnd.n6356 gnd.n6355 185
R6594 gnd.n6359 gnd.n6358 185
R6595 gnd.n6343 gnd.n6342 185
R6596 gnd.n6341 gnd.n6340 185
R6597 gnd.n6320 gnd.n6319 185
R6598 gnd.n6335 gnd.n6334 185
R6599 gnd.n6333 gnd.n6332 185
R6600 gnd.n6324 gnd.n6323 185
R6601 gnd.n6327 gnd.n6326 185
R6602 gnd.n6312 gnd.n6311 185
R6603 gnd.n6310 gnd.n6309 185
R6604 gnd.n6289 gnd.n6288 185
R6605 gnd.n6304 gnd.n6303 185
R6606 gnd.n6302 gnd.n6301 185
R6607 gnd.n6293 gnd.n6292 185
R6608 gnd.n6296 gnd.n6295 185
R6609 gnd.n6280 gnd.n6279 185
R6610 gnd.n6278 gnd.n6277 185
R6611 gnd.n6257 gnd.n6256 185
R6612 gnd.n6272 gnd.n6271 185
R6613 gnd.n6270 gnd.n6269 185
R6614 gnd.n6261 gnd.n6260 185
R6615 gnd.n6264 gnd.n6263 185
R6616 gnd.n6248 gnd.n6247 185
R6617 gnd.n6246 gnd.n6245 185
R6618 gnd.n6225 gnd.n6224 185
R6619 gnd.n6240 gnd.n6239 185
R6620 gnd.n6238 gnd.n6237 185
R6621 gnd.n6229 gnd.n6228 185
R6622 gnd.n6232 gnd.n6231 185
R6623 gnd.n6216 gnd.n6215 185
R6624 gnd.n6214 gnd.n6213 185
R6625 gnd.n6193 gnd.n6192 185
R6626 gnd.n6208 gnd.n6207 185
R6627 gnd.n6206 gnd.n6205 185
R6628 gnd.n6197 gnd.n6196 185
R6629 gnd.n6200 gnd.n6199 185
R6630 gnd.n6185 gnd.n6184 185
R6631 gnd.n6183 gnd.n6182 185
R6632 gnd.n6162 gnd.n6161 185
R6633 gnd.n6177 gnd.n6176 185
R6634 gnd.n6175 gnd.n6174 185
R6635 gnd.n6166 gnd.n6165 185
R6636 gnd.n6169 gnd.n6168 185
R6637 gnd.n5612 gnd.t210 178.987
R6638 gnd.n5240 gnd.t207 178.987
R6639 gnd.n7209 gnd.n525 173.845
R6640 gnd.n7210 gnd.n7209 173.845
R6641 gnd.n7211 gnd.n7210 173.845
R6642 gnd.n7211 gnd.n519 173.845
R6643 gnd.n7219 gnd.n519 173.845
R6644 gnd.n7220 gnd.n7219 173.845
R6645 gnd.n7221 gnd.n7220 173.845
R6646 gnd.n7221 gnd.n513 173.845
R6647 gnd.n7229 gnd.n513 173.845
R6648 gnd.n7230 gnd.n7229 173.845
R6649 gnd.n7231 gnd.n7230 173.845
R6650 gnd.n7231 gnd.n507 173.845
R6651 gnd.n7239 gnd.n507 173.845
R6652 gnd.n7240 gnd.n7239 173.845
R6653 gnd.n7241 gnd.n7240 173.845
R6654 gnd.n7241 gnd.n501 173.845
R6655 gnd.n7249 gnd.n501 173.845
R6656 gnd.n7250 gnd.n7249 173.845
R6657 gnd.n7251 gnd.n7250 173.845
R6658 gnd.n7251 gnd.n495 173.845
R6659 gnd.n7259 gnd.n495 173.845
R6660 gnd.n7260 gnd.n7259 173.845
R6661 gnd.n7261 gnd.n7260 173.845
R6662 gnd.n7261 gnd.n489 173.845
R6663 gnd.n7269 gnd.n489 173.845
R6664 gnd.n7270 gnd.n7269 173.845
R6665 gnd.n7271 gnd.n7270 173.845
R6666 gnd.n7271 gnd.n483 173.845
R6667 gnd.n7279 gnd.n483 173.845
R6668 gnd.n7280 gnd.n7279 173.845
R6669 gnd.n7281 gnd.n7280 173.845
R6670 gnd.n7281 gnd.n477 173.845
R6671 gnd.n7289 gnd.n477 173.845
R6672 gnd.n7290 gnd.n7289 173.845
R6673 gnd.n7291 gnd.n7290 173.845
R6674 gnd.n7291 gnd.n471 173.845
R6675 gnd.n7299 gnd.n471 173.845
R6676 gnd.n7300 gnd.n7299 173.845
R6677 gnd.n7301 gnd.n7300 173.845
R6678 gnd.n7301 gnd.n465 173.845
R6679 gnd.n7309 gnd.n465 173.845
R6680 gnd.n7310 gnd.n7309 173.845
R6681 gnd.n7311 gnd.n7310 173.845
R6682 gnd.n7311 gnd.n459 173.845
R6683 gnd.n7319 gnd.n459 173.845
R6684 gnd.n7320 gnd.n7319 173.845
R6685 gnd.n7321 gnd.n7320 173.845
R6686 gnd.n7321 gnd.n453 173.845
R6687 gnd.n7329 gnd.n453 173.845
R6688 gnd.n7330 gnd.n7329 173.845
R6689 gnd.n7331 gnd.n7330 173.845
R6690 gnd.n7331 gnd.n447 173.845
R6691 gnd.n7339 gnd.n447 173.845
R6692 gnd.n7340 gnd.n7339 173.845
R6693 gnd.n7341 gnd.n7340 173.845
R6694 gnd.n7341 gnd.n441 173.845
R6695 gnd.n7349 gnd.n441 173.845
R6696 gnd.n7350 gnd.n7349 173.845
R6697 gnd.n7351 gnd.n7350 173.845
R6698 gnd.n7351 gnd.n435 173.845
R6699 gnd.n7359 gnd.n435 173.845
R6700 gnd.n7360 gnd.n7359 173.845
R6701 gnd.n7361 gnd.n7360 173.845
R6702 gnd.n7361 gnd.n429 173.845
R6703 gnd.n7369 gnd.n429 173.845
R6704 gnd.n7370 gnd.n7369 173.845
R6705 gnd.n7371 gnd.n7370 173.845
R6706 gnd.n7371 gnd.n423 173.845
R6707 gnd.n7379 gnd.n423 173.845
R6708 gnd.n7380 gnd.n7379 173.845
R6709 gnd.n7381 gnd.n7380 173.845
R6710 gnd.n7381 gnd.n417 173.845
R6711 gnd.n7389 gnd.n417 173.845
R6712 gnd.n7390 gnd.n7389 173.845
R6713 gnd.n7391 gnd.n7390 173.845
R6714 gnd.n7391 gnd.n411 173.845
R6715 gnd.n7399 gnd.n411 173.845
R6716 gnd.n7400 gnd.n7399 173.845
R6717 gnd.n7401 gnd.n7400 173.845
R6718 gnd.n7401 gnd.n405 173.845
R6719 gnd.n7411 gnd.n405 173.845
R6720 gnd.n7412 gnd.n7411 173.845
R6721 gnd.n7413 gnd.n7412 173.845
R6722 gnd.n1 gnd.t352 170.774
R6723 gnd.n7 gnd.t91 170.103
R6724 gnd.n6 gnd.t106 170.103
R6725 gnd.n5 gnd.t173 170.103
R6726 gnd.n4 gnd.t128 170.103
R6727 gnd.n3 gnd.t86 170.103
R6728 gnd.n2 gnd.t335 170.103
R6729 gnd.n1 gnd.t69 170.103
R6730 gnd.n4173 gnd.n4172 163.367
R6731 gnd.n4169 gnd.n4168 163.367
R6732 gnd.n4165 gnd.n4164 163.367
R6733 gnd.n4161 gnd.n4160 163.367
R6734 gnd.n4157 gnd.n4156 163.367
R6735 gnd.n4153 gnd.n4152 163.367
R6736 gnd.n4149 gnd.n4148 163.367
R6737 gnd.n4145 gnd.n4144 163.367
R6738 gnd.n4141 gnd.n4140 163.367
R6739 gnd.n4137 gnd.n4136 163.367
R6740 gnd.n4133 gnd.n4132 163.367
R6741 gnd.n4129 gnd.n4128 163.367
R6742 gnd.n4125 gnd.n4124 163.367
R6743 gnd.n4121 gnd.n4120 163.367
R6744 gnd.n4116 gnd.n4115 163.367
R6745 gnd.n4248 gnd.n1864 163.367
R6746 gnd.n4245 gnd.n4244 163.367
R6747 gnd.n4242 gnd.n1897 163.367
R6748 gnd.n4237 gnd.n4236 163.367
R6749 gnd.n4233 gnd.n4232 163.367
R6750 gnd.n4229 gnd.n4228 163.367
R6751 gnd.n4225 gnd.n4224 163.367
R6752 gnd.n4221 gnd.n4220 163.367
R6753 gnd.n4217 gnd.n4216 163.367
R6754 gnd.n4213 gnd.n4212 163.367
R6755 gnd.n4209 gnd.n4208 163.367
R6756 gnd.n4205 gnd.n4204 163.367
R6757 gnd.n4201 gnd.n4200 163.367
R6758 gnd.n4197 gnd.n4196 163.367
R6759 gnd.n4193 gnd.n4192 163.367
R6760 gnd.n4189 gnd.n4188 163.367
R6761 gnd.n4185 gnd.n4184 163.367
R6762 gnd.n2354 gnd.n1492 163.367
R6763 gnd.n2350 gnd.n1492 163.367
R6764 gnd.n2350 gnd.n2271 163.367
R6765 gnd.n2346 gnd.n2271 163.367
R6766 gnd.n2346 gnd.n2345 163.367
R6767 gnd.n2345 gnd.n2267 163.367
R6768 gnd.n2267 gnd.n2250 163.367
R6769 gnd.n3310 gnd.n2250 163.367
R6770 gnd.n3310 gnd.n2247 163.367
R6771 gnd.n3315 gnd.n2247 163.367
R6772 gnd.n3315 gnd.n2248 163.367
R6773 gnd.n2248 gnd.n2238 163.367
R6774 gnd.n3326 gnd.n2238 163.367
R6775 gnd.n3326 gnd.n2236 163.367
R6776 gnd.n3339 gnd.n2236 163.367
R6777 gnd.n3339 gnd.n2229 163.367
R6778 gnd.n3335 gnd.n2229 163.367
R6779 gnd.n3335 gnd.n3332 163.367
R6780 gnd.n3332 gnd.n3331 163.367
R6781 gnd.n3331 gnd.n2212 163.367
R6782 gnd.n3399 gnd.n2212 163.367
R6783 gnd.n3399 gnd.n2209 163.367
R6784 gnd.n3408 gnd.n2209 163.367
R6785 gnd.n3408 gnd.n2203 163.367
R6786 gnd.n3404 gnd.n2203 163.367
R6787 gnd.n3404 gnd.n2196 163.367
R6788 gnd.n2196 gnd.n2188 163.367
R6789 gnd.n3437 gnd.n2188 163.367
R6790 gnd.n3437 gnd.n2186 163.367
R6791 gnd.n3444 gnd.n2186 163.367
R6792 gnd.n3444 gnd.n2176 163.367
R6793 gnd.n2177 gnd.n2176 163.367
R6794 gnd.n2177 gnd.n2169 163.367
R6795 gnd.n2169 gnd.n2159 163.367
R6796 gnd.n3487 gnd.n2159 163.367
R6797 gnd.n3487 gnd.n2160 163.367
R6798 gnd.n2160 gnd.n2152 163.367
R6799 gnd.n3482 gnd.n2152 163.367
R6800 gnd.n3482 gnd.n2144 163.367
R6801 gnd.n3509 gnd.n2144 163.367
R6802 gnd.n3509 gnd.n2136 163.367
R6803 gnd.n3512 gnd.n2136 163.367
R6804 gnd.n3512 gnd.n2129 163.367
R6805 gnd.n3516 gnd.n2129 163.367
R6806 gnd.n3516 gnd.n2121 163.367
R6807 gnd.n3549 gnd.n2121 163.367
R6808 gnd.n3549 gnd.n2114 163.367
R6809 gnd.n3552 gnd.n2114 163.367
R6810 gnd.n3552 gnd.n2108 163.367
R6811 gnd.n3557 gnd.n2108 163.367
R6812 gnd.n3557 gnd.n2098 163.367
R6813 gnd.n2098 gnd.n2090 163.367
R6814 gnd.n3612 gnd.n2090 163.367
R6815 gnd.n3612 gnd.n2088 163.367
R6816 gnd.n3617 gnd.n2088 163.367
R6817 gnd.n3617 gnd.n2079 163.367
R6818 gnd.n2079 gnd.n2071 163.367
R6819 gnd.n3646 gnd.n2071 163.367
R6820 gnd.n3646 gnd.n2068 163.367
R6821 gnd.n3679 gnd.n2068 163.367
R6822 gnd.n3679 gnd.n2069 163.367
R6823 gnd.n3675 gnd.n2069 163.367
R6824 gnd.n3675 gnd.n3674 163.367
R6825 gnd.n3674 gnd.n2050 163.367
R6826 gnd.n2051 gnd.n2050 163.367
R6827 gnd.n2051 gnd.n2044 163.367
R6828 gnd.n3668 gnd.n2044 163.367
R6829 gnd.n3668 gnd.n2037 163.367
R6830 gnd.n3664 gnd.n2037 163.367
R6831 gnd.n3664 gnd.n2031 163.367
R6832 gnd.n3661 gnd.n2031 163.367
R6833 gnd.n3661 gnd.n2023 163.367
R6834 gnd.n3654 gnd.n2023 163.367
R6835 gnd.n3654 gnd.n2018 163.367
R6836 gnd.n3651 gnd.n2018 163.367
R6837 gnd.n3651 gnd.n2006 163.367
R6838 gnd.n2006 gnd.n2000 163.367
R6839 gnd.n3777 gnd.n2000 163.367
R6840 gnd.n3777 gnd.n1998 163.367
R6841 gnd.n3782 gnd.n1998 163.367
R6842 gnd.n3782 gnd.n1988 163.367
R6843 gnd.n1988 gnd.n1980 163.367
R6844 gnd.n3810 gnd.n1980 163.367
R6845 gnd.n3810 gnd.n1977 163.367
R6846 gnd.n3817 gnd.n1977 163.367
R6847 gnd.n3817 gnd.n1978 163.367
R6848 gnd.n1978 gnd.n1967 163.367
R6849 gnd.n1967 gnd.n1957 163.367
R6850 gnd.n1957 gnd.n1950 163.367
R6851 gnd.n3853 gnd.n1950 163.367
R6852 gnd.n3853 gnd.n1948 163.367
R6853 gnd.n3859 gnd.n1948 163.367
R6854 gnd.n3859 gnd.n1908 163.367
R6855 gnd.n1908 gnd.n1901 163.367
R6856 gnd.n4180 gnd.n1901 163.367
R6857 gnd.n1467 gnd.n1466 163.367
R6858 gnd.n4844 gnd.n1466 163.367
R6859 gnd.n4842 gnd.n4841 163.367
R6860 gnd.n4838 gnd.n4837 163.367
R6861 gnd.n4834 gnd.n4833 163.367
R6862 gnd.n4830 gnd.n4829 163.367
R6863 gnd.n4826 gnd.n4825 163.367
R6864 gnd.n4822 gnd.n4821 163.367
R6865 gnd.n4818 gnd.n4817 163.367
R6866 gnd.n4814 gnd.n4813 163.367
R6867 gnd.n4810 gnd.n4809 163.367
R6868 gnd.n4806 gnd.n4805 163.367
R6869 gnd.n4802 gnd.n4801 163.367
R6870 gnd.n4798 gnd.n4797 163.367
R6871 gnd.n4794 gnd.n4793 163.367
R6872 gnd.n4790 gnd.n4789 163.367
R6873 gnd.n4853 gnd.n1432 163.367
R6874 gnd.n2283 gnd.n2282 163.367
R6875 gnd.n2288 gnd.n2287 163.367
R6876 gnd.n2292 gnd.n2291 163.367
R6877 gnd.n2296 gnd.n2295 163.367
R6878 gnd.n2300 gnd.n2299 163.367
R6879 gnd.n2304 gnd.n2303 163.367
R6880 gnd.n2308 gnd.n2307 163.367
R6881 gnd.n2312 gnd.n2311 163.367
R6882 gnd.n2316 gnd.n2315 163.367
R6883 gnd.n2320 gnd.n2319 163.367
R6884 gnd.n2324 gnd.n2323 163.367
R6885 gnd.n2328 gnd.n2327 163.367
R6886 gnd.n2332 gnd.n2331 163.367
R6887 gnd.n2336 gnd.n2335 163.367
R6888 gnd.n2340 gnd.n2339 163.367
R6889 gnd.n4782 gnd.n1468 163.367
R6890 gnd.n4782 gnd.n1490 163.367
R6891 gnd.n3270 gnd.n1490 163.367
R6892 gnd.n3271 gnd.n3270 163.367
R6893 gnd.n3271 gnd.n2268 163.367
R6894 gnd.n3275 gnd.n2268 163.367
R6895 gnd.n3275 gnd.n2253 163.367
R6896 gnd.n3308 gnd.n2253 163.367
R6897 gnd.n3308 gnd.n2254 163.367
R6898 gnd.n2254 gnd.n2246 163.367
R6899 gnd.n3303 gnd.n2246 163.367
R6900 gnd.n3303 gnd.n2257 163.367
R6901 gnd.n2257 gnd.n2234 163.367
R6902 gnd.n3343 gnd.n2234 163.367
R6903 gnd.n3343 gnd.n2231 163.367
R6904 gnd.n3356 gnd.n2231 163.367
R6905 gnd.n3356 gnd.n2232 163.367
R6906 gnd.n3352 gnd.n2232 163.367
R6907 gnd.n3352 gnd.n3351 163.367
R6908 gnd.n3351 gnd.n3350 163.367
R6909 gnd.n3350 gnd.n2207 163.367
R6910 gnd.n3412 gnd.n2207 163.367
R6911 gnd.n3412 gnd.n2205 163.367
R6912 gnd.n3416 gnd.n2205 163.367
R6913 gnd.n3416 gnd.n2194 163.367
R6914 gnd.n3430 gnd.n2194 163.367
R6915 gnd.n3430 gnd.n2191 163.367
R6916 gnd.n3435 gnd.n2191 163.367
R6917 gnd.n3435 gnd.n2192 163.367
R6918 gnd.n2192 gnd.n2174 163.367
R6919 gnd.n3462 gnd.n2174 163.367
R6920 gnd.n3462 gnd.n2172 163.367
R6921 gnd.n3466 gnd.n2172 163.367
R6922 gnd.n3466 gnd.n2157 163.367
R6923 gnd.n3489 gnd.n2157 163.367
R6924 gnd.n3489 gnd.n2154 163.367
R6925 gnd.n3496 gnd.n2154 163.367
R6926 gnd.n3496 gnd.n2155 163.367
R6927 gnd.n3492 gnd.n2155 163.367
R6928 gnd.n3492 gnd.n2134 163.367
R6929 gnd.n3529 gnd.n2134 163.367
R6930 gnd.n3529 gnd.n2131 163.367
R6931 gnd.n3536 gnd.n2131 163.367
R6932 gnd.n3536 gnd.n2132 163.367
R6933 gnd.n3532 gnd.n2132 163.367
R6934 gnd.n3532 gnd.n2112 163.367
R6935 gnd.n3588 gnd.n2112 163.367
R6936 gnd.n3588 gnd.n2110 163.367
R6937 gnd.n3592 gnd.n2110 163.367
R6938 gnd.n3592 gnd.n2097 163.367
R6939 gnd.n3605 gnd.n2097 163.367
R6940 gnd.n3605 gnd.n2094 163.367
R6941 gnd.n3610 gnd.n2094 163.367
R6942 gnd.n3610 gnd.n2095 163.367
R6943 gnd.n2095 gnd.n2077 163.367
R6944 gnd.n3632 gnd.n2077 163.367
R6945 gnd.n3632 gnd.n2074 163.367
R6946 gnd.n3644 gnd.n2074 163.367
R6947 gnd.n3644 gnd.n2075 163.367
R6948 gnd.n2075 gnd.n2066 163.367
R6949 gnd.n3639 gnd.n2066 163.367
R6950 gnd.n3639 gnd.n3636 163.367
R6951 gnd.n3636 gnd.n2048 163.367
R6952 gnd.n3703 gnd.n2048 163.367
R6953 gnd.n3703 gnd.n2046 163.367
R6954 gnd.n3707 gnd.n2046 163.367
R6955 gnd.n3707 gnd.n2035 163.367
R6956 gnd.n3722 gnd.n2035 163.367
R6957 gnd.n3722 gnd.n2033 163.367
R6958 gnd.n3726 gnd.n2033 163.367
R6959 gnd.n3726 gnd.n2022 163.367
R6960 gnd.n3753 gnd.n2022 163.367
R6961 gnd.n3753 gnd.n2020 163.367
R6962 gnd.n3757 gnd.n2020 163.367
R6963 gnd.n3757 gnd.n2004 163.367
R6964 gnd.n3770 gnd.n2004 163.367
R6965 gnd.n3770 gnd.n2001 163.367
R6966 gnd.n3775 gnd.n2001 163.367
R6967 gnd.n3775 gnd.n2002 163.367
R6968 gnd.n2002 gnd.n1987 163.367
R6969 gnd.n3800 gnd.n1987 163.367
R6970 gnd.n3800 gnd.n1984 163.367
R6971 gnd.n3808 gnd.n1984 163.367
R6972 gnd.n3808 gnd.n1985 163.367
R6973 gnd.n1985 gnd.n1975 163.367
R6974 gnd.n3803 gnd.n1975 163.367
R6975 gnd.n3803 gnd.n1955 163.367
R6976 gnd.n3846 gnd.n1955 163.367
R6977 gnd.n3846 gnd.n1952 163.367
R6978 gnd.n3851 gnd.n1952 163.367
R6979 gnd.n3851 gnd.n1953 163.367
R6980 gnd.n1953 gnd.n1906 163.367
R6981 gnd.n4090 gnd.n1906 163.367
R6982 gnd.n4090 gnd.n1903 163.367
R6983 gnd.n4178 gnd.n1903 163.367
R6984 gnd.n4111 gnd.n4110 156.462
R6985 gnd.n6347 gnd.n6315 153.042
R6986 gnd.n6411 gnd.n6410 152.079
R6987 gnd.n6379 gnd.n6378 152.079
R6988 gnd.n6347 gnd.n6346 152.079
R6989 gnd.n1481 gnd.n1480 152
R6990 gnd.n1482 gnd.n1471 152
R6991 gnd.n1484 gnd.n1483 152
R6992 gnd.n1486 gnd.n1469 152
R6993 gnd.n1488 gnd.n1487 152
R6994 gnd.n4109 gnd.n4093 152
R6995 gnd.n4101 gnd.n4094 152
R6996 gnd.n4100 gnd.n4099 152
R6997 gnd.n4098 gnd.n4095 152
R6998 gnd.n4096 gnd.t220 150.546
R6999 gnd.t41 gnd.n6389 147.661
R7000 gnd.t5 gnd.n6357 147.661
R7001 gnd.t43 gnd.n6325 147.661
R7002 gnd.t182 gnd.n6294 147.661
R7003 gnd.t179 gnd.n6262 147.661
R7004 gnd.t125 gnd.n6230 147.661
R7005 gnd.t137 gnd.n6198 147.661
R7006 gnd.t10 gnd.n6167 147.661
R7007 gnd.n4247 gnd.n1863 143.351
R7008 gnd.n1448 gnd.n1431 143.351
R7009 gnd.n4852 gnd.n1431 143.351
R7010 gnd.n7413 gnd.n212 132.349
R7011 gnd.n1478 gnd.t278 130.484
R7012 gnd.n1487 gnd.t299 126.766
R7013 gnd.n1485 gnd.t231 126.766
R7014 gnd.n1471 gnd.t290 126.766
R7015 gnd.n1479 gnd.t251 126.766
R7016 gnd.n4097 gnd.t201 126.766
R7017 gnd.n4099 gnd.t315 126.766
R7018 gnd.n4108 gnd.t264 126.766
R7019 gnd.n4110 gnd.t248 126.766
R7020 gnd.n6406 gnd.n6405 104.615
R7021 gnd.n6405 gnd.n6383 104.615
R7022 gnd.n6398 gnd.n6383 104.615
R7023 gnd.n6398 gnd.n6397 104.615
R7024 gnd.n6397 gnd.n6387 104.615
R7025 gnd.n6390 gnd.n6387 104.615
R7026 gnd.n6374 gnd.n6373 104.615
R7027 gnd.n6373 gnd.n6351 104.615
R7028 gnd.n6366 gnd.n6351 104.615
R7029 gnd.n6366 gnd.n6365 104.615
R7030 gnd.n6365 gnd.n6355 104.615
R7031 gnd.n6358 gnd.n6355 104.615
R7032 gnd.n6342 gnd.n6341 104.615
R7033 gnd.n6341 gnd.n6319 104.615
R7034 gnd.n6334 gnd.n6319 104.615
R7035 gnd.n6334 gnd.n6333 104.615
R7036 gnd.n6333 gnd.n6323 104.615
R7037 gnd.n6326 gnd.n6323 104.615
R7038 gnd.n6311 gnd.n6310 104.615
R7039 gnd.n6310 gnd.n6288 104.615
R7040 gnd.n6303 gnd.n6288 104.615
R7041 gnd.n6303 gnd.n6302 104.615
R7042 gnd.n6302 gnd.n6292 104.615
R7043 gnd.n6295 gnd.n6292 104.615
R7044 gnd.n6279 gnd.n6278 104.615
R7045 gnd.n6278 gnd.n6256 104.615
R7046 gnd.n6271 gnd.n6256 104.615
R7047 gnd.n6271 gnd.n6270 104.615
R7048 gnd.n6270 gnd.n6260 104.615
R7049 gnd.n6263 gnd.n6260 104.615
R7050 gnd.n6247 gnd.n6246 104.615
R7051 gnd.n6246 gnd.n6224 104.615
R7052 gnd.n6239 gnd.n6224 104.615
R7053 gnd.n6239 gnd.n6238 104.615
R7054 gnd.n6238 gnd.n6228 104.615
R7055 gnd.n6231 gnd.n6228 104.615
R7056 gnd.n6215 gnd.n6214 104.615
R7057 gnd.n6214 gnd.n6192 104.615
R7058 gnd.n6207 gnd.n6192 104.615
R7059 gnd.n6207 gnd.n6206 104.615
R7060 gnd.n6206 gnd.n6196 104.615
R7061 gnd.n6199 gnd.n6196 104.615
R7062 gnd.n6184 gnd.n6183 104.615
R7063 gnd.n6183 gnd.n6161 104.615
R7064 gnd.n6176 gnd.n6161 104.615
R7065 gnd.n6176 gnd.n6175 104.615
R7066 gnd.n6175 gnd.n6165 104.615
R7067 gnd.n6168 gnd.n6165 104.615
R7068 gnd.n5761 gnd.t277 100.632
R7069 gnd.n5195 gnd.t307 100.632
R7070 gnd.n7667 gnd.n219 99.6594
R7071 gnd.n7665 gnd.n7664 99.6594
R7072 gnd.n7660 gnd.n226 99.6594
R7073 gnd.n7658 gnd.n7657 99.6594
R7074 gnd.n7653 gnd.n233 99.6594
R7075 gnd.n7651 gnd.n7650 99.6594
R7076 gnd.n7646 gnd.n240 99.6594
R7077 gnd.n7644 gnd.n7643 99.6594
R7078 gnd.n7636 gnd.n247 99.6594
R7079 gnd.n7634 gnd.n7633 99.6594
R7080 gnd.n7629 gnd.n254 99.6594
R7081 gnd.n7627 gnd.n7626 99.6594
R7082 gnd.n7622 gnd.n261 99.6594
R7083 gnd.n7620 gnd.n7619 99.6594
R7084 gnd.n7615 gnd.n268 99.6594
R7085 gnd.n7613 gnd.n7612 99.6594
R7086 gnd.n7608 gnd.n275 99.6594
R7087 gnd.n7606 gnd.n7605 99.6594
R7088 gnd.n285 gnd.n284 99.6594
R7089 gnd.n7597 gnd.n7596 99.6594
R7090 gnd.n7594 gnd.n7593 99.6594
R7091 gnd.n7589 gnd.n293 99.6594
R7092 gnd.n7587 gnd.n7586 99.6594
R7093 gnd.n7582 gnd.n300 99.6594
R7094 gnd.n7580 gnd.n7579 99.6594
R7095 gnd.n7575 gnd.n307 99.6594
R7096 gnd.n7573 gnd.n7572 99.6594
R7097 gnd.n7568 gnd.n316 99.6594
R7098 gnd.n7566 gnd.n7565 99.6594
R7099 gnd.n4279 gnd.n1623 99.6594
R7100 gnd.n4283 gnd.n4282 99.6594
R7101 gnd.n4290 gnd.n4289 99.6594
R7102 gnd.n4293 gnd.n4292 99.6594
R7103 gnd.n4300 gnd.n4299 99.6594
R7104 gnd.n4303 gnd.n4302 99.6594
R7105 gnd.n4310 gnd.n4309 99.6594
R7106 gnd.n4313 gnd.n4312 99.6594
R7107 gnd.n4323 gnd.n4322 99.6594
R7108 gnd.n4326 gnd.n4325 99.6594
R7109 gnd.n4333 gnd.n4332 99.6594
R7110 gnd.n4336 gnd.n4335 99.6594
R7111 gnd.n4344 gnd.n4343 99.6594
R7112 gnd.n4349 gnd.n4348 99.6594
R7113 gnd.n4356 gnd.n4355 99.6594
R7114 gnd.n4359 gnd.n4358 99.6594
R7115 gnd.n4366 gnd.n4365 99.6594
R7116 gnd.n4369 gnd.n4368 99.6594
R7117 gnd.n4378 gnd.n4377 99.6594
R7118 gnd.n4381 gnd.n4380 99.6594
R7119 gnd.n4388 gnd.n4387 99.6594
R7120 gnd.n4391 gnd.n4390 99.6594
R7121 gnd.n4398 gnd.n4397 99.6594
R7122 gnd.n4401 gnd.n4400 99.6594
R7123 gnd.n4408 gnd.n4407 99.6594
R7124 gnd.n4411 gnd.n4410 99.6594
R7125 gnd.n4419 gnd.n4418 99.6594
R7126 gnd.n4422 gnd.n4421 99.6594
R7127 gnd.n4898 gnd.n4897 99.6594
R7128 gnd.n4895 gnd.n4894 99.6594
R7129 gnd.n4890 gnd.n1390 99.6594
R7130 gnd.n4888 gnd.n4887 99.6594
R7131 gnd.n4883 gnd.n1397 99.6594
R7132 gnd.n4881 gnd.n4880 99.6594
R7133 gnd.n4876 gnd.n1404 99.6594
R7134 gnd.n4874 gnd.n4873 99.6594
R7135 gnd.n4868 gnd.n1413 99.6594
R7136 gnd.n4866 gnd.n4865 99.6594
R7137 gnd.n4861 gnd.n1420 99.6594
R7138 gnd.n4859 gnd.n4858 99.6594
R7139 gnd.n2984 gnd.n2983 99.6594
R7140 gnd.n2988 gnd.n2986 99.6594
R7141 gnd.n2994 gnd.n2978 99.6594
R7142 gnd.n2998 gnd.n2996 99.6594
R7143 gnd.n3004 gnd.n2974 99.6594
R7144 gnd.n3008 gnd.n3006 99.6594
R7145 gnd.n3014 gnd.n2968 99.6594
R7146 gnd.n3018 gnd.n3016 99.6594
R7147 gnd.n3024 gnd.n2964 99.6594
R7148 gnd.n3028 gnd.n3026 99.6594
R7149 gnd.n3034 gnd.n2960 99.6594
R7150 gnd.n3038 gnd.n3036 99.6594
R7151 gnd.n3044 gnd.n2956 99.6594
R7152 gnd.n3048 gnd.n3046 99.6594
R7153 gnd.n3054 gnd.n2952 99.6594
R7154 gnd.n3057 gnd.n3056 99.6594
R7155 gnd.n5163 gnd.n5162 99.6594
R7156 gnd.n5157 gnd.n1030 99.6594
R7157 gnd.n5154 gnd.n1031 99.6594
R7158 gnd.n5150 gnd.n1032 99.6594
R7159 gnd.n5146 gnd.n1033 99.6594
R7160 gnd.n5142 gnd.n1034 99.6594
R7161 gnd.n5138 gnd.n1035 99.6594
R7162 gnd.n5134 gnd.n1036 99.6594
R7163 gnd.n5130 gnd.n1037 99.6594
R7164 gnd.n5125 gnd.n1038 99.6594
R7165 gnd.n5121 gnd.n1039 99.6594
R7166 gnd.n5117 gnd.n1040 99.6594
R7167 gnd.n5113 gnd.n1041 99.6594
R7168 gnd.n5109 gnd.n1042 99.6594
R7169 gnd.n5105 gnd.n1043 99.6594
R7170 gnd.n5101 gnd.n1044 99.6594
R7171 gnd.n5097 gnd.n1045 99.6594
R7172 gnd.n5093 gnd.n1046 99.6594
R7173 gnd.n5089 gnd.n1047 99.6594
R7174 gnd.n5085 gnd.n1048 99.6594
R7175 gnd.n5081 gnd.n1049 99.6594
R7176 gnd.n5077 gnd.n1050 99.6594
R7177 gnd.n5073 gnd.n1051 99.6594
R7178 gnd.n5069 gnd.n1052 99.6594
R7179 gnd.n5065 gnd.n1053 99.6594
R7180 gnd.n5061 gnd.n1054 99.6594
R7181 gnd.n5057 gnd.n1055 99.6594
R7182 gnd.n5053 gnd.n1056 99.6594
R7183 gnd.n5049 gnd.n1057 99.6594
R7184 gnd.n6537 gnd.n5175 99.6594
R7185 gnd.n6535 gnd.n6534 99.6594
R7186 gnd.n6530 gnd.n5182 99.6594
R7187 gnd.n6528 gnd.n6527 99.6594
R7188 gnd.n6523 gnd.n5189 99.6594
R7189 gnd.n6521 gnd.n6520 99.6594
R7190 gnd.n6516 gnd.n5198 99.6594
R7191 gnd.n6514 gnd.n6513 99.6594
R7192 gnd.n5794 gnd.n5793 99.6594
R7193 gnd.n5788 gnd.n5736 99.6594
R7194 gnd.n5785 gnd.n5737 99.6594
R7195 gnd.n5781 gnd.n5738 99.6594
R7196 gnd.n5777 gnd.n5739 99.6594
R7197 gnd.n5773 gnd.n5740 99.6594
R7198 gnd.n5769 gnd.n5741 99.6594
R7199 gnd.n5765 gnd.n5742 99.6594
R7200 gnd.n7557 gnd.n322 99.6594
R7201 gnd.n7555 gnd.n7554 99.6594
R7202 gnd.n7550 gnd.n329 99.6594
R7203 gnd.n7548 gnd.n7547 99.6594
R7204 gnd.n7543 gnd.n336 99.6594
R7205 gnd.n7541 gnd.n7540 99.6594
R7206 gnd.n7536 gnd.n343 99.6594
R7207 gnd.n7534 gnd.n7533 99.6594
R7208 gnd.n348 gnd.n347 99.6594
R7209 gnd.n3971 gnd.n3970 99.6594
R7210 gnd.n3987 gnd.n3986 99.6594
R7211 gnd.n3990 gnd.n3989 99.6594
R7212 gnd.n4006 gnd.n4005 99.6594
R7213 gnd.n4009 gnd.n4008 99.6594
R7214 gnd.n4025 gnd.n4024 99.6594
R7215 gnd.n4028 gnd.n4027 99.6594
R7216 gnd.n4045 gnd.n4044 99.6594
R7217 gnd.n4048 gnd.n4047 99.6594
R7218 gnd.n6505 gnd.n5205 99.6594
R7219 gnd.n6503 gnd.n6502 99.6594
R7220 gnd.n6498 gnd.n5212 99.6594
R7221 gnd.n6496 gnd.n6495 99.6594
R7222 gnd.n6491 gnd.n5219 99.6594
R7223 gnd.n6489 gnd.n6488 99.6594
R7224 gnd.n6484 gnd.n5226 99.6594
R7225 gnd.n6482 gnd.n6481 99.6594
R7226 gnd.n6477 gnd.n5233 99.6594
R7227 gnd.n6475 gnd.n6474 99.6594
R7228 gnd.n6470 gnd.n5242 99.6594
R7229 gnd.n6468 gnd.n6467 99.6594
R7230 gnd.n6463 gnd.n6462 99.6594
R7231 gnd.n5666 gnd.n5576 99.6594
R7232 gnd.n5664 gnd.n5579 99.6594
R7233 gnd.n5660 gnd.n5659 99.6594
R7234 gnd.n5653 gnd.n5584 99.6594
R7235 gnd.n5652 gnd.n5651 99.6594
R7236 gnd.n5645 gnd.n5590 99.6594
R7237 gnd.n5644 gnd.n5643 99.6594
R7238 gnd.n5637 gnd.n5596 99.6594
R7239 gnd.n5636 gnd.n5635 99.6594
R7240 gnd.n5629 gnd.n5602 99.6594
R7241 gnd.n5628 gnd.n5627 99.6594
R7242 gnd.n5620 gnd.n5608 99.6594
R7243 gnd.n5619 gnd.n5618 99.6594
R7244 gnd.n3072 gnd.n3071 99.6594
R7245 gnd.n3083 gnd.n3082 99.6594
R7246 gnd.n3092 gnd.n3091 99.6594
R7247 gnd.n3095 gnd.n3094 99.6594
R7248 gnd.n3106 gnd.n3105 99.6594
R7249 gnd.n3115 gnd.n3114 99.6594
R7250 gnd.n3119 gnd.n3117 99.6594
R7251 gnd.n3187 gnd.n2407 99.6594
R7252 gnd.n3190 gnd.n3189 99.6594
R7253 gnd.n2563 gnd.n1058 99.6594
R7254 gnd.n2567 gnd.n1059 99.6594
R7255 gnd.n2573 gnd.n1060 99.6594
R7256 gnd.n2577 gnd.n1061 99.6594
R7257 gnd.n2583 gnd.n1062 99.6594
R7258 gnd.n2587 gnd.n1063 99.6594
R7259 gnd.n2593 gnd.n1064 99.6594
R7260 gnd.n2597 gnd.n1065 99.6594
R7261 gnd.n2554 gnd.n1066 99.6594
R7262 gnd.n2566 gnd.n1058 99.6594
R7263 gnd.n2572 gnd.n1059 99.6594
R7264 gnd.n2576 gnd.n1060 99.6594
R7265 gnd.n2582 gnd.n1061 99.6594
R7266 gnd.n2586 gnd.n1062 99.6594
R7267 gnd.n2592 gnd.n1063 99.6594
R7268 gnd.n2596 gnd.n1064 99.6594
R7269 gnd.n2553 gnd.n1065 99.6594
R7270 gnd.n2549 gnd.n1066 99.6594
R7271 gnd.n3189 gnd.n3188 99.6594
R7272 gnd.n3118 gnd.n2407 99.6594
R7273 gnd.n3117 gnd.n3116 99.6594
R7274 gnd.n3114 gnd.n3107 99.6594
R7275 gnd.n3105 gnd.n3104 99.6594
R7276 gnd.n3094 gnd.n3093 99.6594
R7277 gnd.n3091 gnd.n3084 99.6594
R7278 gnd.n3082 gnd.n3081 99.6594
R7279 gnd.n3071 gnd.n3070 99.6594
R7280 gnd.n5667 gnd.n5666 99.6594
R7281 gnd.n5661 gnd.n5579 99.6594
R7282 gnd.n5659 gnd.n5658 99.6594
R7283 gnd.n5654 gnd.n5653 99.6594
R7284 gnd.n5651 gnd.n5650 99.6594
R7285 gnd.n5646 gnd.n5645 99.6594
R7286 gnd.n5643 gnd.n5642 99.6594
R7287 gnd.n5638 gnd.n5637 99.6594
R7288 gnd.n5635 gnd.n5634 99.6594
R7289 gnd.n5630 gnd.n5629 99.6594
R7290 gnd.n5627 gnd.n5626 99.6594
R7291 gnd.n5621 gnd.n5620 99.6594
R7292 gnd.n5618 gnd.n5574 99.6594
R7293 gnd.n6462 gnd.n5244 99.6594
R7294 gnd.n6469 gnd.n6468 99.6594
R7295 gnd.n5242 gnd.n5234 99.6594
R7296 gnd.n6476 gnd.n6475 99.6594
R7297 gnd.n5233 gnd.n5227 99.6594
R7298 gnd.n6483 gnd.n6482 99.6594
R7299 gnd.n5226 gnd.n5220 99.6594
R7300 gnd.n6490 gnd.n6489 99.6594
R7301 gnd.n5219 gnd.n5213 99.6594
R7302 gnd.n6497 gnd.n6496 99.6594
R7303 gnd.n5212 gnd.n5206 99.6594
R7304 gnd.n6504 gnd.n6503 99.6594
R7305 gnd.n5205 gnd.n5202 99.6594
R7306 gnd.n3970 gnd.n3935 99.6594
R7307 gnd.n3988 gnd.n3987 99.6594
R7308 gnd.n3989 gnd.n3926 99.6594
R7309 gnd.n4007 gnd.n4006 99.6594
R7310 gnd.n4008 gnd.n3917 99.6594
R7311 gnd.n4026 gnd.n4025 99.6594
R7312 gnd.n4027 gnd.n3908 99.6594
R7313 gnd.n4046 gnd.n4045 99.6594
R7314 gnd.n4047 gnd.n3904 99.6594
R7315 gnd.n347 gnd.n344 99.6594
R7316 gnd.n7535 gnd.n7534 99.6594
R7317 gnd.n343 gnd.n337 99.6594
R7318 gnd.n7542 gnd.n7541 99.6594
R7319 gnd.n336 gnd.n330 99.6594
R7320 gnd.n7549 gnd.n7548 99.6594
R7321 gnd.n329 gnd.n323 99.6594
R7322 gnd.n7556 gnd.n7555 99.6594
R7323 gnd.n322 gnd.n319 99.6594
R7324 gnd.n5794 gnd.n5744 99.6594
R7325 gnd.n5786 gnd.n5736 99.6594
R7326 gnd.n5782 gnd.n5737 99.6594
R7327 gnd.n5778 gnd.n5738 99.6594
R7328 gnd.n5774 gnd.n5739 99.6594
R7329 gnd.n5770 gnd.n5740 99.6594
R7330 gnd.n5766 gnd.n5741 99.6594
R7331 gnd.n5742 gnd.n5536 99.6594
R7332 gnd.n6515 gnd.n6514 99.6594
R7333 gnd.n5198 gnd.n5190 99.6594
R7334 gnd.n6522 gnd.n6521 99.6594
R7335 gnd.n5189 gnd.n5183 99.6594
R7336 gnd.n6529 gnd.n6528 99.6594
R7337 gnd.n5182 gnd.n5176 99.6594
R7338 gnd.n6536 gnd.n6535 99.6594
R7339 gnd.n5175 gnd.n5172 99.6594
R7340 gnd.n5163 gnd.n1070 99.6594
R7341 gnd.n5155 gnd.n1030 99.6594
R7342 gnd.n5151 gnd.n1031 99.6594
R7343 gnd.n5147 gnd.n1032 99.6594
R7344 gnd.n5143 gnd.n1033 99.6594
R7345 gnd.n5139 gnd.n1034 99.6594
R7346 gnd.n5135 gnd.n1035 99.6594
R7347 gnd.n5131 gnd.n1036 99.6594
R7348 gnd.n5126 gnd.n1037 99.6594
R7349 gnd.n5122 gnd.n1038 99.6594
R7350 gnd.n5118 gnd.n1039 99.6594
R7351 gnd.n5114 gnd.n1040 99.6594
R7352 gnd.n5110 gnd.n1041 99.6594
R7353 gnd.n5106 gnd.n1042 99.6594
R7354 gnd.n5102 gnd.n1043 99.6594
R7355 gnd.n5098 gnd.n1044 99.6594
R7356 gnd.n5094 gnd.n1045 99.6594
R7357 gnd.n5090 gnd.n1046 99.6594
R7358 gnd.n5086 gnd.n1047 99.6594
R7359 gnd.n5082 gnd.n1048 99.6594
R7360 gnd.n5078 gnd.n1049 99.6594
R7361 gnd.n5074 gnd.n1050 99.6594
R7362 gnd.n5070 gnd.n1051 99.6594
R7363 gnd.n5066 gnd.n1052 99.6594
R7364 gnd.n5062 gnd.n1053 99.6594
R7365 gnd.n5058 gnd.n1054 99.6594
R7366 gnd.n5054 gnd.n1055 99.6594
R7367 gnd.n5050 gnd.n1056 99.6594
R7368 gnd.n1140 gnd.n1057 99.6594
R7369 gnd.n3056 gnd.n3055 99.6594
R7370 gnd.n3047 gnd.n2952 99.6594
R7371 gnd.n3046 gnd.n3045 99.6594
R7372 gnd.n3037 gnd.n2956 99.6594
R7373 gnd.n3036 gnd.n3035 99.6594
R7374 gnd.n3027 gnd.n2960 99.6594
R7375 gnd.n3026 gnd.n3025 99.6594
R7376 gnd.n3017 gnd.n2964 99.6594
R7377 gnd.n3016 gnd.n3015 99.6594
R7378 gnd.n3007 gnd.n2968 99.6594
R7379 gnd.n3006 gnd.n3005 99.6594
R7380 gnd.n2997 gnd.n2974 99.6594
R7381 gnd.n2996 gnd.n2995 99.6594
R7382 gnd.n2987 gnd.n2978 99.6594
R7383 gnd.n2986 gnd.n2985 99.6594
R7384 gnd.n1426 gnd.n1421 99.6594
R7385 gnd.n4860 gnd.n4859 99.6594
R7386 gnd.n1420 gnd.n1414 99.6594
R7387 gnd.n4867 gnd.n4866 99.6594
R7388 gnd.n1413 gnd.n1405 99.6594
R7389 gnd.n4875 gnd.n4874 99.6594
R7390 gnd.n1404 gnd.n1398 99.6594
R7391 gnd.n4882 gnd.n4881 99.6594
R7392 gnd.n1397 gnd.n1391 99.6594
R7393 gnd.n4889 gnd.n4888 99.6594
R7394 gnd.n1390 gnd.n1383 99.6594
R7395 gnd.n4896 gnd.n4895 99.6594
R7396 gnd.n4899 gnd.n4898 99.6594
R7397 gnd.n4280 gnd.n4279 99.6594
R7398 gnd.n4282 gnd.n4271 99.6594
R7399 gnd.n4291 gnd.n4290 99.6594
R7400 gnd.n4292 gnd.n4267 99.6594
R7401 gnd.n4301 gnd.n4300 99.6594
R7402 gnd.n4302 gnd.n4263 99.6594
R7403 gnd.n4311 gnd.n4310 99.6594
R7404 gnd.n4312 gnd.n4259 99.6594
R7405 gnd.n4324 gnd.n4323 99.6594
R7406 gnd.n4325 gnd.n4255 99.6594
R7407 gnd.n4334 gnd.n4333 99.6594
R7408 gnd.n4335 gnd.n4251 99.6594
R7409 gnd.n4347 gnd.n4346 99.6594
R7410 gnd.n4348 gnd.n1857 99.6594
R7411 gnd.n4357 gnd.n4356 99.6594
R7412 gnd.n4358 gnd.n1853 99.6594
R7413 gnd.n4367 gnd.n4366 99.6594
R7414 gnd.n4368 gnd.n1849 99.6594
R7415 gnd.n4379 gnd.n4378 99.6594
R7416 gnd.n4380 gnd.n1845 99.6594
R7417 gnd.n4389 gnd.n4388 99.6594
R7418 gnd.n4390 gnd.n1841 99.6594
R7419 gnd.n4399 gnd.n4398 99.6594
R7420 gnd.n4400 gnd.n1837 99.6594
R7421 gnd.n4409 gnd.n4408 99.6594
R7422 gnd.n4410 gnd.n1833 99.6594
R7423 gnd.n4420 gnd.n4419 99.6594
R7424 gnd.n4423 gnd.n4422 99.6594
R7425 gnd.n7567 gnd.n7566 99.6594
R7426 gnd.n316 gnd.n308 99.6594
R7427 gnd.n7574 gnd.n7573 99.6594
R7428 gnd.n307 gnd.n301 99.6594
R7429 gnd.n7581 gnd.n7580 99.6594
R7430 gnd.n300 gnd.n294 99.6594
R7431 gnd.n7588 gnd.n7587 99.6594
R7432 gnd.n293 gnd.n287 99.6594
R7433 gnd.n7595 gnd.n7594 99.6594
R7434 gnd.n7598 gnd.n7597 99.6594
R7435 gnd.n284 gnd.n276 99.6594
R7436 gnd.n7607 gnd.n7606 99.6594
R7437 gnd.n275 gnd.n269 99.6594
R7438 gnd.n7614 gnd.n7613 99.6594
R7439 gnd.n268 gnd.n262 99.6594
R7440 gnd.n7621 gnd.n7620 99.6594
R7441 gnd.n261 gnd.n255 99.6594
R7442 gnd.n7628 gnd.n7627 99.6594
R7443 gnd.n254 gnd.n248 99.6594
R7444 gnd.n7635 gnd.n7634 99.6594
R7445 gnd.n247 gnd.n241 99.6594
R7446 gnd.n7645 gnd.n7644 99.6594
R7447 gnd.n240 gnd.n234 99.6594
R7448 gnd.n7652 gnd.n7651 99.6594
R7449 gnd.n233 gnd.n227 99.6594
R7450 gnd.n7659 gnd.n7658 99.6594
R7451 gnd.n226 gnd.n220 99.6594
R7452 gnd.n7666 gnd.n7665 99.6594
R7453 gnd.n219 gnd.n216 99.6594
R7454 gnd.n3179 gnd.n3178 99.6594
R7455 gnd.n2944 gnd.n2927 99.6594
R7456 gnd.n2946 gnd.n2928 99.6594
R7457 gnd.n3063 gnd.n2929 99.6594
R7458 gnd.n3065 gnd.n2930 99.6594
R7459 gnd.n3076 gnd.n2931 99.6594
R7460 gnd.n3078 gnd.n2932 99.6594
R7461 gnd.n3088 gnd.n2933 99.6594
R7462 gnd.n3099 gnd.n2934 99.6594
R7463 gnd.n3101 gnd.n2935 99.6594
R7464 gnd.n3111 gnd.n2936 99.6594
R7465 gnd.n3122 gnd.n2937 99.6594
R7466 gnd.n3182 gnd.n3181 99.6594
R7467 gnd.n2938 gnd.n2402 99.6594
R7468 gnd.n3179 gnd.n2940 99.6594
R7469 gnd.n2945 gnd.n2927 99.6594
R7470 gnd.n3062 gnd.n2928 99.6594
R7471 gnd.n3064 gnd.n2929 99.6594
R7472 gnd.n3075 gnd.n2930 99.6594
R7473 gnd.n3077 gnd.n2931 99.6594
R7474 gnd.n3087 gnd.n2932 99.6594
R7475 gnd.n3098 gnd.n2933 99.6594
R7476 gnd.n3100 gnd.n2934 99.6594
R7477 gnd.n3110 gnd.n2935 99.6594
R7478 gnd.n3121 gnd.n2936 99.6594
R7479 gnd.n2937 gnd.n2414 99.6594
R7480 gnd.n3181 gnd.n2415 99.6594
R7481 gnd.n2938 gnd.n2398 99.6594
R7482 gnd.n3951 gnd.n3947 99.6594
R7483 gnd.n3955 gnd.n3953 99.6594
R7484 gnd.n3962 gnd.n3943 99.6594
R7485 gnd.n3966 gnd.n3964 99.6594
R7486 gnd.n3977 gnd.n3940 99.6594
R7487 gnd.n3981 gnd.n3979 99.6594
R7488 gnd.n3996 gnd.n3931 99.6594
R7489 gnd.n4000 gnd.n3998 99.6594
R7490 gnd.n4015 gnd.n3922 99.6594
R7491 gnd.n4019 gnd.n4017 99.6594
R7492 gnd.n4034 gnd.n3913 99.6594
R7493 gnd.n4037 gnd.n4036 99.6594
R7494 gnd.n4055 gnd.n4054 99.6594
R7495 gnd.n4058 gnd.n4057 99.6594
R7496 gnd.n4036 gnd.n4035 99.6594
R7497 gnd.n4018 gnd.n3913 99.6594
R7498 gnd.n4017 gnd.n4016 99.6594
R7499 gnd.n3999 gnd.n3922 99.6594
R7500 gnd.n3998 gnd.n3997 99.6594
R7501 gnd.n3980 gnd.n3931 99.6594
R7502 gnd.n3979 gnd.n3978 99.6594
R7503 gnd.n3965 gnd.n3940 99.6594
R7504 gnd.n3964 gnd.n3963 99.6594
R7505 gnd.n3954 gnd.n3943 99.6594
R7506 gnd.n3953 gnd.n3952 99.6594
R7507 gnd.n3947 gnd.n1597 99.6594
R7508 gnd.n4059 gnd.n4058 99.6594
R7509 gnd.n4056 gnd.n4055 99.6594
R7510 gnd.n2411 gnd.t263 98.63
R7511 gnd.n3905 gnd.t289 98.63
R7512 gnd.n2404 gnd.t313 98.63
R7513 gnd.n4318 gnd.t286 98.63
R7514 gnd.n4370 gnd.t283 98.63
R7515 gnd.n1829 gnd.t215 98.63
R7516 gnd.n313 gnd.t310 98.63
R7517 gnd.n280 gnd.t229 98.63
R7518 gnd.n7638 gnd.t268 98.63
R7519 gnd.n350 gnd.t255 98.63
R7520 gnd.n1090 gnd.t243 98.63
R7521 gnd.n1112 gnd.t240 98.63
R7522 gnd.n1134 gnd.t219 98.63
R7523 gnd.n2550 gnd.t298 98.63
R7524 gnd.n1409 gnd.t303 98.63
R7525 gnd.n2949 gnd.t236 98.63
R7526 gnd.n2971 gnd.t258 98.63
R7527 gnd.n3895 gnd.t246 98.63
R7528 gnd.n2279 gnd.t273 92.8196
R7529 gnd.n1898 gnd.t294 92.8196
R7530 gnd.n4786 gnd.t320 92.8118
R7531 gnd.n4112 gnd.t225 92.8118
R7532 gnd.n1478 gnd.n1477 81.8399
R7533 gnd.n4250 gnd.n4249 78.9125
R7534 gnd.n4855 gnd.n4854 78.9125
R7535 gnd.n5762 gnd.t276 74.8376
R7536 gnd.n5196 gnd.t308 74.8376
R7537 gnd.n2280 gnd.t272 72.8438
R7538 gnd.n1899 gnd.t295 72.8438
R7539 gnd.n1479 gnd.n1472 72.8411
R7540 gnd.n1485 gnd.n1470 72.8411
R7541 gnd.n4108 gnd.n4107 72.8411
R7542 gnd.n2412 gnd.t262 72.836
R7543 gnd.n4787 gnd.t319 72.836
R7544 gnd.n4113 gnd.t226 72.836
R7545 gnd.n3906 gnd.t288 72.836
R7546 gnd.n2405 gnd.t314 72.836
R7547 gnd.n4319 gnd.t285 72.836
R7548 gnd.n4371 gnd.t282 72.836
R7549 gnd.n1830 gnd.t214 72.836
R7550 gnd.n314 gnd.t311 72.836
R7551 gnd.n281 gnd.t230 72.836
R7552 gnd.n7639 gnd.t269 72.836
R7553 gnd.n351 gnd.t256 72.836
R7554 gnd.n1091 gnd.t242 72.836
R7555 gnd.n1113 gnd.t239 72.836
R7556 gnd.n1135 gnd.t218 72.836
R7557 gnd.n2551 gnd.t297 72.836
R7558 gnd.n1410 gnd.t304 72.836
R7559 gnd.n2950 gnd.t237 72.836
R7560 gnd.n2972 gnd.t259 72.836
R7561 gnd.n3896 gnd.t247 72.836
R7562 gnd.n4173 gnd.n1866 71.676
R7563 gnd.n4169 gnd.n1867 71.676
R7564 gnd.n4165 gnd.n1868 71.676
R7565 gnd.n4161 gnd.n1869 71.676
R7566 gnd.n4157 gnd.n1870 71.676
R7567 gnd.n4153 gnd.n1871 71.676
R7568 gnd.n4149 gnd.n1872 71.676
R7569 gnd.n4145 gnd.n1873 71.676
R7570 gnd.n4141 gnd.n1874 71.676
R7571 gnd.n4137 gnd.n1875 71.676
R7572 gnd.n4133 gnd.n1876 71.676
R7573 gnd.n4129 gnd.n1877 71.676
R7574 gnd.n4125 gnd.n1878 71.676
R7575 gnd.n4121 gnd.n1879 71.676
R7576 gnd.n4116 gnd.n1880 71.676
R7577 gnd.n1881 gnd.n1864 71.676
R7578 gnd.n4245 gnd.n1863 71.676
R7579 gnd.n4243 gnd.n4242 71.676
R7580 gnd.n4237 gnd.n1896 71.676
R7581 gnd.n4233 gnd.n1895 71.676
R7582 gnd.n4229 gnd.n1894 71.676
R7583 gnd.n4225 gnd.n1893 71.676
R7584 gnd.n4221 gnd.n1892 71.676
R7585 gnd.n4217 gnd.n1891 71.676
R7586 gnd.n4213 gnd.n1890 71.676
R7587 gnd.n4209 gnd.n1889 71.676
R7588 gnd.n4205 gnd.n1888 71.676
R7589 gnd.n4201 gnd.n1887 71.676
R7590 gnd.n4197 gnd.n1886 71.676
R7591 gnd.n4193 gnd.n1885 71.676
R7592 gnd.n4189 gnd.n1884 71.676
R7593 gnd.n4185 gnd.n1883 71.676
R7594 gnd.n4181 gnd.n1882 71.676
R7595 gnd.n4850 gnd.n4849 71.676
R7596 gnd.n4844 gnd.n1434 71.676
R7597 gnd.n4841 gnd.n1435 71.676
R7598 gnd.n4837 gnd.n1436 71.676
R7599 gnd.n4833 gnd.n1437 71.676
R7600 gnd.n4829 gnd.n1438 71.676
R7601 gnd.n4825 gnd.n1439 71.676
R7602 gnd.n4821 gnd.n1440 71.676
R7603 gnd.n4817 gnd.n1441 71.676
R7604 gnd.n4813 gnd.n1442 71.676
R7605 gnd.n4809 gnd.n1443 71.676
R7606 gnd.n4805 gnd.n1444 71.676
R7607 gnd.n4801 gnd.n1445 71.676
R7608 gnd.n4797 gnd.n1446 71.676
R7609 gnd.n4793 gnd.n1447 71.676
R7610 gnd.n4789 gnd.n1448 71.676
R7611 gnd.n1449 gnd.n1432 71.676
R7612 gnd.n2283 gnd.n1450 71.676
R7613 gnd.n2288 gnd.n1451 71.676
R7614 gnd.n2292 gnd.n1452 71.676
R7615 gnd.n2296 gnd.n1453 71.676
R7616 gnd.n2300 gnd.n1454 71.676
R7617 gnd.n2304 gnd.n1455 71.676
R7618 gnd.n2308 gnd.n1456 71.676
R7619 gnd.n2312 gnd.n1457 71.676
R7620 gnd.n2316 gnd.n1458 71.676
R7621 gnd.n2320 gnd.n1459 71.676
R7622 gnd.n2324 gnd.n1460 71.676
R7623 gnd.n2328 gnd.n1461 71.676
R7624 gnd.n2332 gnd.n1462 71.676
R7625 gnd.n2336 gnd.n1463 71.676
R7626 gnd.n2340 gnd.n1464 71.676
R7627 gnd.n4850 gnd.n1467 71.676
R7628 gnd.n4842 gnd.n1434 71.676
R7629 gnd.n4838 gnd.n1435 71.676
R7630 gnd.n4834 gnd.n1436 71.676
R7631 gnd.n4830 gnd.n1437 71.676
R7632 gnd.n4826 gnd.n1438 71.676
R7633 gnd.n4822 gnd.n1439 71.676
R7634 gnd.n4818 gnd.n1440 71.676
R7635 gnd.n4814 gnd.n1441 71.676
R7636 gnd.n4810 gnd.n1442 71.676
R7637 gnd.n4806 gnd.n1443 71.676
R7638 gnd.n4802 gnd.n1444 71.676
R7639 gnd.n4798 gnd.n1445 71.676
R7640 gnd.n4794 gnd.n1446 71.676
R7641 gnd.n4790 gnd.n1447 71.676
R7642 gnd.n4853 gnd.n4852 71.676
R7643 gnd.n2282 gnd.n1449 71.676
R7644 gnd.n2287 gnd.n1450 71.676
R7645 gnd.n2291 gnd.n1451 71.676
R7646 gnd.n2295 gnd.n1452 71.676
R7647 gnd.n2299 gnd.n1453 71.676
R7648 gnd.n2303 gnd.n1454 71.676
R7649 gnd.n2307 gnd.n1455 71.676
R7650 gnd.n2311 gnd.n1456 71.676
R7651 gnd.n2315 gnd.n1457 71.676
R7652 gnd.n2319 gnd.n1458 71.676
R7653 gnd.n2323 gnd.n1459 71.676
R7654 gnd.n2327 gnd.n1460 71.676
R7655 gnd.n2331 gnd.n1461 71.676
R7656 gnd.n2335 gnd.n1462 71.676
R7657 gnd.n2339 gnd.n1463 71.676
R7658 gnd.n2278 gnd.n1464 71.676
R7659 gnd.n4184 gnd.n1882 71.676
R7660 gnd.n4188 gnd.n1883 71.676
R7661 gnd.n4192 gnd.n1884 71.676
R7662 gnd.n4196 gnd.n1885 71.676
R7663 gnd.n4200 gnd.n1886 71.676
R7664 gnd.n4204 gnd.n1887 71.676
R7665 gnd.n4208 gnd.n1888 71.676
R7666 gnd.n4212 gnd.n1889 71.676
R7667 gnd.n4216 gnd.n1890 71.676
R7668 gnd.n4220 gnd.n1891 71.676
R7669 gnd.n4224 gnd.n1892 71.676
R7670 gnd.n4228 gnd.n1893 71.676
R7671 gnd.n4232 gnd.n1894 71.676
R7672 gnd.n4236 gnd.n1895 71.676
R7673 gnd.n1897 gnd.n1896 71.676
R7674 gnd.n4244 gnd.n4243 71.676
R7675 gnd.n4248 gnd.n4247 71.676
R7676 gnd.n4115 gnd.n1881 71.676
R7677 gnd.n4120 gnd.n1880 71.676
R7678 gnd.n4124 gnd.n1879 71.676
R7679 gnd.n4128 gnd.n1878 71.676
R7680 gnd.n4132 gnd.n1877 71.676
R7681 gnd.n4136 gnd.n1876 71.676
R7682 gnd.n4140 gnd.n1875 71.676
R7683 gnd.n4144 gnd.n1874 71.676
R7684 gnd.n4148 gnd.n1873 71.676
R7685 gnd.n4152 gnd.n1872 71.676
R7686 gnd.n4156 gnd.n1871 71.676
R7687 gnd.n4160 gnd.n1870 71.676
R7688 gnd.n4164 gnd.n1869 71.676
R7689 gnd.n4168 gnd.n1868 71.676
R7690 gnd.n4172 gnd.n1867 71.676
R7691 gnd.n1904 gnd.n1866 71.676
R7692 gnd.n8 gnd.t108 69.1507
R7693 gnd.n14 gnd.t147 68.4792
R7694 gnd.n13 gnd.t67 68.4792
R7695 gnd.n12 gnd.t71 68.4792
R7696 gnd.n11 gnd.t17 68.4792
R7697 gnd.n10 gnd.t322 68.4792
R7698 gnd.n9 gnd.t103 68.4792
R7699 gnd.n8 gnd.t195 68.4792
R7700 gnd.n5674 gnd.n5575 64.369
R7701 gnd.n2285 gnd.n2280 59.5399
R7702 gnd.n4239 gnd.n1899 59.5399
R7703 gnd.n4788 gnd.n4787 59.5399
R7704 gnd.n4118 gnd.n4113 59.5399
R7705 gnd.n4785 gnd.n1488 59.1804
R7706 gnd.n6545 gnd.n5165 57.3586
R7707 gnd.n5164 gnd.n1068 57.3586
R7708 gnd.n7675 gnd.n212 57.3586
R7709 gnd.n5381 gnd.t15 56.407
R7710 gnd.n5334 gnd.t131 56.407
R7711 gnd.n5349 gnd.t163 56.407
R7712 gnd.n5365 gnd.t154 56.407
R7713 gnd.n64 gnd.t142 56.407
R7714 gnd.n17 gnd.t37 56.407
R7715 gnd.n32 gnd.t176 56.407
R7716 gnd.n48 gnd.t166 56.407
R7717 gnd.n5394 gnd.t143 55.8337
R7718 gnd.n5347 gnd.t57 55.8337
R7719 gnd.n5362 gnd.t366 55.8337
R7720 gnd.n5378 gnd.t94 55.8337
R7721 gnd.n77 gnd.t141 55.8337
R7722 gnd.n30 gnd.t349 55.8337
R7723 gnd.n45 gnd.t355 55.8337
R7724 gnd.n61 gnd.t328 55.8337
R7725 gnd.n1476 gnd.n1475 54.358
R7726 gnd.n4105 gnd.n4104 54.358
R7727 gnd.n5381 gnd.n5380 53.0052
R7728 gnd.n5383 gnd.n5382 53.0052
R7729 gnd.n5385 gnd.n5384 53.0052
R7730 gnd.n5387 gnd.n5386 53.0052
R7731 gnd.n5389 gnd.n5388 53.0052
R7732 gnd.n5391 gnd.n5390 53.0052
R7733 gnd.n5393 gnd.n5392 53.0052
R7734 gnd.n5334 gnd.n5333 53.0052
R7735 gnd.n5336 gnd.n5335 53.0052
R7736 gnd.n5338 gnd.n5337 53.0052
R7737 gnd.n5340 gnd.n5339 53.0052
R7738 gnd.n5342 gnd.n5341 53.0052
R7739 gnd.n5344 gnd.n5343 53.0052
R7740 gnd.n5346 gnd.n5345 53.0052
R7741 gnd.n5349 gnd.n5348 53.0052
R7742 gnd.n5351 gnd.n5350 53.0052
R7743 gnd.n5353 gnd.n5352 53.0052
R7744 gnd.n5355 gnd.n5354 53.0052
R7745 gnd.n5357 gnd.n5356 53.0052
R7746 gnd.n5359 gnd.n5358 53.0052
R7747 gnd.n5361 gnd.n5360 53.0052
R7748 gnd.n5365 gnd.n5364 53.0052
R7749 gnd.n5367 gnd.n5366 53.0052
R7750 gnd.n5369 gnd.n5368 53.0052
R7751 gnd.n5371 gnd.n5370 53.0052
R7752 gnd.n5373 gnd.n5372 53.0052
R7753 gnd.n5375 gnd.n5374 53.0052
R7754 gnd.n5377 gnd.n5376 53.0052
R7755 gnd.n76 gnd.n75 53.0052
R7756 gnd.n74 gnd.n73 53.0052
R7757 gnd.n72 gnd.n71 53.0052
R7758 gnd.n70 gnd.n69 53.0052
R7759 gnd.n68 gnd.n67 53.0052
R7760 gnd.n66 gnd.n65 53.0052
R7761 gnd.n64 gnd.n63 53.0052
R7762 gnd.n29 gnd.n28 53.0052
R7763 gnd.n27 gnd.n26 53.0052
R7764 gnd.n25 gnd.n24 53.0052
R7765 gnd.n23 gnd.n22 53.0052
R7766 gnd.n21 gnd.n20 53.0052
R7767 gnd.n19 gnd.n18 53.0052
R7768 gnd.n17 gnd.n16 53.0052
R7769 gnd.n44 gnd.n43 53.0052
R7770 gnd.n42 gnd.n41 53.0052
R7771 gnd.n40 gnd.n39 53.0052
R7772 gnd.n38 gnd.n37 53.0052
R7773 gnd.n36 gnd.n35 53.0052
R7774 gnd.n34 gnd.n33 53.0052
R7775 gnd.n32 gnd.n31 53.0052
R7776 gnd.n60 gnd.n59 53.0052
R7777 gnd.n58 gnd.n57 53.0052
R7778 gnd.n56 gnd.n55 53.0052
R7779 gnd.n54 gnd.n53 53.0052
R7780 gnd.n52 gnd.n51 53.0052
R7781 gnd.n50 gnd.n49 53.0052
R7782 gnd.n48 gnd.n47 53.0052
R7783 gnd.n4096 gnd.n4095 52.4801
R7784 gnd.n6390 gnd.t41 52.3082
R7785 gnd.n6358 gnd.t5 52.3082
R7786 gnd.n6326 gnd.t43 52.3082
R7787 gnd.n6295 gnd.t182 52.3082
R7788 gnd.n6263 gnd.t179 52.3082
R7789 gnd.n6231 gnd.t125 52.3082
R7790 gnd.n6199 gnd.t137 52.3082
R7791 gnd.n6168 gnd.t10 52.3082
R7792 gnd.n6220 gnd.n6188 51.4173
R7793 gnd.n6284 gnd.n6283 50.455
R7794 gnd.n6252 gnd.n6251 50.455
R7795 gnd.n6220 gnd.n6219 50.455
R7796 gnd.n5612 gnd.n5611 45.1884
R7797 gnd.n5240 gnd.n5239 45.1884
R7798 gnd.n4176 gnd.n4111 44.3322
R7799 gnd.n1479 gnd.n1478 44.3189
R7800 gnd.n2413 gnd.n2412 42.2793
R7801 gnd.n4050 gnd.n3906 42.2793
R7802 gnd.n5624 gnd.n5612 42.2793
R7803 gnd.n5241 gnd.n5240 42.2793
R7804 gnd.n5764 gnd.n5762 42.2793
R7805 gnd.n5197 gnd.n5196 42.2793
R7806 gnd.n2406 gnd.n2405 42.2793
R7807 gnd.n4320 gnd.n4319 42.2793
R7808 gnd.n4372 gnd.n4371 42.2793
R7809 gnd.n1831 gnd.n1830 42.2793
R7810 gnd.n315 gnd.n314 42.2793
R7811 gnd.n7603 gnd.n281 42.2793
R7812 gnd.n7640 gnd.n7639 42.2793
R7813 gnd.n7531 gnd.n351 42.2793
R7814 gnd.n5128 gnd.n1091 42.2793
R7815 gnd.n5088 gnd.n1113 42.2793
R7816 gnd.n5048 gnd.n1135 42.2793
R7817 gnd.n2603 gnd.n2551 42.2793
R7818 gnd.n4870 gnd.n1410 42.2793
R7819 gnd.n2951 gnd.n2950 42.2793
R7820 gnd.n2973 gnd.n2972 42.2793
R7821 gnd.n3897 gnd.n3896 42.2793
R7822 gnd.n1477 gnd.n1476 41.6274
R7823 gnd.n4106 gnd.n4105 41.6274
R7824 gnd.n1486 gnd.n1485 40.8975
R7825 gnd.n4109 gnd.n4108 40.8975
R7826 gnd.n6749 gnd.n801 39.6473
R7827 gnd.n6743 gnd.n801 39.6473
R7828 gnd.n6743 gnd.n6742 39.6473
R7829 gnd.n6742 gnd.n6741 39.6473
R7830 gnd.n6741 gnd.n808 39.6473
R7831 gnd.n6735 gnd.n808 39.6473
R7832 gnd.n6735 gnd.n6734 39.6473
R7833 gnd.n6734 gnd.n6733 39.6473
R7834 gnd.n6733 gnd.n816 39.6473
R7835 gnd.n6727 gnd.n816 39.6473
R7836 gnd.n6727 gnd.n6726 39.6473
R7837 gnd.n6726 gnd.n6725 39.6473
R7838 gnd.n6725 gnd.n824 39.6473
R7839 gnd.n6719 gnd.n824 39.6473
R7840 gnd.n6719 gnd.n6718 39.6473
R7841 gnd.n6718 gnd.n6717 39.6473
R7842 gnd.n6717 gnd.n832 39.6473
R7843 gnd.n6711 gnd.n832 39.6473
R7844 gnd.n6711 gnd.n6710 39.6473
R7845 gnd.n6710 gnd.n6709 39.6473
R7846 gnd.n6709 gnd.n840 39.6473
R7847 gnd.n6703 gnd.n840 39.6473
R7848 gnd.n6703 gnd.n6702 39.6473
R7849 gnd.n6702 gnd.n6701 39.6473
R7850 gnd.n6701 gnd.n848 39.6473
R7851 gnd.n6695 gnd.n848 39.6473
R7852 gnd.n6695 gnd.n6694 39.6473
R7853 gnd.n6694 gnd.n6693 39.6473
R7854 gnd.n6693 gnd.n856 39.6473
R7855 gnd.n6687 gnd.n856 39.6473
R7856 gnd.n6687 gnd.n6686 39.6473
R7857 gnd.n6686 gnd.n6685 39.6473
R7858 gnd.n6685 gnd.n864 39.6473
R7859 gnd.n6679 gnd.n864 39.6473
R7860 gnd.n6679 gnd.n6678 39.6473
R7861 gnd.n6678 gnd.n6677 39.6473
R7862 gnd.n6677 gnd.n872 39.6473
R7863 gnd.n6671 gnd.n872 39.6473
R7864 gnd.n6671 gnd.n6670 39.6473
R7865 gnd.n6670 gnd.n6669 39.6473
R7866 gnd.n6669 gnd.n880 39.6473
R7867 gnd.n6663 gnd.n880 39.6473
R7868 gnd.n6663 gnd.n6662 39.6473
R7869 gnd.n6662 gnd.n6661 39.6473
R7870 gnd.n6661 gnd.n888 39.6473
R7871 gnd.n6655 gnd.n888 39.6473
R7872 gnd.n6655 gnd.n6654 39.6473
R7873 gnd.n6654 gnd.n6653 39.6473
R7874 gnd.n6653 gnd.n896 39.6473
R7875 gnd.n6647 gnd.n896 39.6473
R7876 gnd.n6647 gnd.n6646 39.6473
R7877 gnd.n6646 gnd.n6645 39.6473
R7878 gnd.n6645 gnd.n904 39.6473
R7879 gnd.n6639 gnd.n904 39.6473
R7880 gnd.n6639 gnd.n6638 39.6473
R7881 gnd.n6638 gnd.n6637 39.6473
R7882 gnd.n6637 gnd.n912 39.6473
R7883 gnd.n6631 gnd.n912 39.6473
R7884 gnd.n6631 gnd.n6630 39.6473
R7885 gnd.n6630 gnd.n6629 39.6473
R7886 gnd.n6629 gnd.n920 39.6473
R7887 gnd.n6623 gnd.n920 39.6473
R7888 gnd.n6623 gnd.n6622 39.6473
R7889 gnd.n6622 gnd.n6621 39.6473
R7890 gnd.n6621 gnd.n928 39.6473
R7891 gnd.n6615 gnd.n928 39.6473
R7892 gnd.n6615 gnd.n6614 39.6473
R7893 gnd.n6614 gnd.n6613 39.6473
R7894 gnd.n6613 gnd.n936 39.6473
R7895 gnd.n6607 gnd.n936 39.6473
R7896 gnd.n6607 gnd.n6606 39.6473
R7897 gnd.n6606 gnd.n6605 39.6473
R7898 gnd.n6605 gnd.n944 39.6473
R7899 gnd.n6599 gnd.n944 39.6473
R7900 gnd.n6599 gnd.n6598 39.6473
R7901 gnd.n6598 gnd.n6597 39.6473
R7902 gnd.n6597 gnd.n952 39.6473
R7903 gnd.n6591 gnd.n952 39.6473
R7904 gnd.n6591 gnd.n6590 39.6473
R7905 gnd.n6590 gnd.n6589 39.6473
R7906 gnd.n6589 gnd.n960 39.6473
R7907 gnd.n6583 gnd.n960 39.6473
R7908 gnd.n6583 gnd.n6582 39.6473
R7909 gnd.n1485 gnd.n1484 35.055
R7910 gnd.n1480 gnd.n1479 35.055
R7911 gnd.n4098 gnd.n4097 35.055
R7912 gnd.n4108 gnd.n4094 35.055
R7913 gnd.n5674 gnd.n5570 31.8661
R7914 gnd.n5682 gnd.n5570 31.8661
R7915 gnd.n5690 gnd.n5564 31.8661
R7916 gnd.n5690 gnd.n5558 31.8661
R7917 gnd.n5698 gnd.n5558 31.8661
R7918 gnd.n5698 gnd.n5551 31.8661
R7919 gnd.n5706 gnd.n5551 31.8661
R7920 gnd.n5706 gnd.n5552 31.8661
R7921 gnd.n5805 gnd.n5537 31.8661
R7922 gnd.n5040 gnd.n1068 31.8661
R7923 gnd.n5034 gnd.n1152 31.8661
R7924 gnd.n5034 gnd.n1155 31.8661
R7925 gnd.n5028 gnd.n1155 31.8661
R7926 gnd.n5028 gnd.n1167 31.8661
R7927 gnd.n5022 gnd.n1177 31.8661
R7928 gnd.n2916 gnd.n1376 31.8661
R7929 gnd.n2918 gnd.n2416 31.8661
R7930 gnd.n2926 gnd.n2416 31.8661
R7931 gnd.n3202 gnd.n2397 31.8661
R7932 gnd.n4662 gnd.n1600 31.8661
R7933 gnd.n4656 gnd.n4655 31.8661
R7934 gnd.n4655 gnd.n4654 31.8661
R7935 gnd.n4648 gnd.n1618 31.8661
R7936 gnd.n7699 gnd.n175 31.8661
R7937 gnd.n7693 gnd.n185 31.8661
R7938 gnd.n7687 gnd.n185 31.8661
R7939 gnd.n7687 gnd.n194 31.8661
R7940 gnd.n7681 gnd.n194 31.8661
R7941 gnd.n7675 gnd.n209 31.8661
R7942 gnd.n4182 gnd.n1900 31.3761
R7943 gnd.n2353 gnd.n2342 31.3761
R7944 gnd.n5010 gnd.n1194 26.7676
R7945 gnd.n5004 gnd.n1204 26.7676
R7946 gnd.n2682 gnd.n1207 26.7676
R7947 gnd.n2688 gnd.n1217 26.7676
R7948 gnd.n4992 gnd.n1224 26.7676
R7949 gnd.n4986 gnd.n1235 26.7676
R7950 gnd.n4980 gnd.n1245 26.7676
R7951 gnd.n2503 gnd.n1248 26.7676
R7952 gnd.n2715 gnd.n2506 26.7676
R7953 gnd.n2747 gnd.n2488 26.7676
R7954 gnd.n2741 gnd.n2484 26.7676
R7955 gnd.n2766 gnd.n2474 26.7676
R7956 gnd.n2802 gnd.n2460 26.7676
R7957 gnd.n2773 gnd.n1265 26.7676
R7958 gnd.n4966 gnd.n1274 26.7676
R7959 gnd.n2779 gnd.n2778 26.7676
R7960 gnd.n4960 gnd.n1283 26.7676
R7961 gnd.n4954 gnd.n1293 26.7676
R7962 gnd.n2841 gnd.n1296 26.7676
R7963 gnd.n2849 gnd.n1306 26.7676
R7964 gnd.n4942 gnd.n1313 26.7676
R7965 gnd.n2856 gnd.n2443 26.7676
R7966 gnd.n4936 gnd.n1323 26.7676
R7967 gnd.n4930 gnd.n1333 26.7676
R7968 gnd.n2898 gnd.n1336 26.7676
R7969 gnd.n2871 gnd.n1346 26.7676
R7970 gnd.n4918 gnd.n1353 26.7676
R7971 gnd.n2876 gnd.n1356 26.7676
R7972 gnd.n4912 gnd.n1364 26.7676
R7973 gnd.n4906 gnd.n1373 26.7676
R7974 gnd.n4647 gnd.n1621 26.7676
R7975 gnd.n4641 gnd.n1633 26.7676
R7976 gnd.n4434 gnd.n1642 26.7676
R7977 gnd.n4635 gnd.n1645 26.7676
R7978 gnd.n4442 gnd.n1653 26.7676
R7979 gnd.n4448 gnd.n1662 26.7676
R7980 gnd.n4623 gnd.n1665 26.7676
R7981 gnd.n4617 gnd.n1676 26.7676
R7982 gnd.n4493 gnd.n4492 26.7676
R7983 gnd.n4611 gnd.n1685 26.7676
R7984 gnd.n4463 gnd.n1693 26.7676
R7985 gnd.n4468 gnd.n1702 26.7676
R7986 gnd.n4599 gnd.n1705 26.7676
R7987 gnd.n4593 gnd.n1716 26.7676
R7988 gnd.n4516 gnd.n4515 26.7676
R7989 gnd.n4587 gnd.n1725 26.7676
R7990 gnd.n4546 gnd.n1731 26.7676
R7991 gnd.n4557 gnd.n1740 26.7676
R7992 gnd.n4575 gnd.n1743 26.7676
R7993 gnd.n4524 gnd.n1751 26.7676
R7994 gnd.n7749 gnd.n87 26.7676
R7995 gnd.n7441 gnd.n381 26.7676
R7996 gnd.n7741 gnd.n105 26.7676
R7997 gnd.n7452 gnd.n114 26.7676
R7998 gnd.n7460 gnd.n123 26.7676
R7999 gnd.n7466 gnd.n132 26.7676
R8000 gnd.n7723 gnd.n135 26.7676
R8001 gnd.n7717 gnd.n146 26.7676
R8002 gnd.n7480 gnd.n153 26.7676
R8003 gnd.n7489 gnd.n163 26.7676
R8004 gnd.n2752 gnd.t18 26.4489
R8005 gnd.n4536 gnd.t12 26.4489
R8006 gnd.n2697 gnd.t38 25.8116
R8007 gnd.n7729 gnd.t52 25.8116
R8008 gnd.n2412 gnd.n2411 25.7944
R8009 gnd.n3906 gnd.n3905 25.7944
R8010 gnd.n5762 gnd.n5761 25.7944
R8011 gnd.n5196 gnd.n5195 25.7944
R8012 gnd.n2405 gnd.n2404 25.7944
R8013 gnd.n4319 gnd.n4318 25.7944
R8014 gnd.n4371 gnd.n4370 25.7944
R8015 gnd.n1830 gnd.n1829 25.7944
R8016 gnd.n314 gnd.n313 25.7944
R8017 gnd.n281 gnd.n280 25.7944
R8018 gnd.n7639 gnd.n7638 25.7944
R8019 gnd.n351 gnd.n350 25.7944
R8020 gnd.n1091 gnd.n1090 25.7944
R8021 gnd.n1113 gnd.n1112 25.7944
R8022 gnd.n1135 gnd.n1134 25.7944
R8023 gnd.n2551 gnd.n2550 25.7944
R8024 gnd.n1410 gnd.n1409 25.7944
R8025 gnd.n2950 gnd.n2949 25.7944
R8026 gnd.n2972 gnd.n2971 25.7944
R8027 gnd.n3896 gnd.n3895 25.7944
R8028 gnd.n2629 gnd.t129 25.1743
R8029 gnd.n7705 gnd.t81 25.1743
R8030 gnd.n5806 gnd.n5526 24.8557
R8031 gnd.n5529 gnd.n5520 24.8557
R8032 gnd.n5827 gnd.n5505 24.8557
R8033 gnd.n5846 gnd.n5845 24.8557
R8034 gnd.n5856 gnd.n5498 24.8557
R8035 gnd.n5869 gnd.n5486 24.8557
R8036 gnd.n5894 gnd.n5470 24.8557
R8037 gnd.n5893 gnd.n5472 24.8557
R8038 gnd.n5916 gnd.n5454 24.8557
R8039 gnd.n5905 gnd.n5446 24.8557
R8040 gnd.n5941 gnd.n5940 24.8557
R8041 gnd.n5951 gnd.n5439 24.8557
R8042 gnd.n5963 gnd.n5431 24.8557
R8043 gnd.n5962 gnd.n5419 24.8557
R8044 gnd.n5981 gnd.n5980 24.8557
R8045 gnd.n6002 gnd.n5400 24.8557
R8046 gnd.n6026 gnd.n6025 24.8557
R8047 gnd.n6037 gnd.n5319 24.8557
R8048 gnd.n6036 gnd.n5321 24.8557
R8049 gnd.n6048 gnd.n5312 24.8557
R8050 gnd.n6065 gnd.n6064 24.8557
R8051 gnd.n5303 gnd.n5292 24.8557
R8052 gnd.n6088 gnd.n5282 24.8557
R8053 gnd.n5284 gnd.n5283 24.8557
R8054 gnd.n6111 gnd.n5276 24.8557
R8055 gnd.n6122 gnd.n6121 24.8557
R8056 gnd.n6136 gnd.n5263 24.8557
R8057 gnd.n6574 gnd.n979 24.8557
R8058 gnd.n6437 gnd.n990 24.8557
R8059 gnd.n6567 gnd.n6566 24.8557
R8060 gnd.n6560 gnd.n1002 24.8557
R8061 gnd.n6559 gnd.n1005 24.8557
R8062 gnd.n6426 gnd.n1016 24.8557
R8063 gnd.n6546 gnd.n1027 24.8557
R8064 gnd.n6582 gnd.n6581 23.7886
R8065 gnd.n5824 gnd.t9 23.2624
R8066 gnd.n5816 gnd.t275 22.6251
R8067 gnd.n5040 gnd.t217 22.6251
R8068 gnd.t115 gnd.n1197 22.6251
R8069 gnd.n2883 gnd.t235 22.6251
R8070 gnd.n3886 gnd.t213 22.6251
R8071 gnd.n362 gnd.t23 22.6251
R8072 gnd.n209 gnd.t228 22.6251
R8073 gnd.t109 gnd.n1238 21.9878
R8074 gnd.n374 gnd.t88 21.9878
R8075 gnd.n5796 gnd.t181 21.3504
R8076 gnd.n2740 gnd.t27 21.3504
R8077 gnd.t2 gnd.n4571 21.3504
R8078 gnd.n6101 gnd.t73 20.7131
R8079 gnd.t50 gnd.n1286 20.7131
R8080 gnd.t34 gnd.n1713 20.7131
R8081 gnd.n2916 gnd.n1381 20.3945
R8082 gnd.n1618 gnd.n1610 20.3945
R8083 gnd.t101 gnd.n5293 20.0758
R8084 gnd.t92 gnd.n1326 20.0758
R8085 gnd.t58 gnd.n1673 20.0758
R8086 gnd.n2280 gnd.n2279 19.9763
R8087 gnd.n1899 gnd.n1898 19.9763
R8088 gnd.n4787 gnd.n4786 19.9763
R8089 gnd.n4113 gnd.n4112 19.9763
R8090 gnd.n1474 gnd.t233 19.8005
R8091 gnd.n1474 gnd.t292 19.8005
R8092 gnd.n1473 gnd.t253 19.8005
R8093 gnd.n1473 gnd.t280 19.8005
R8094 gnd.n4103 gnd.t203 19.8005
R8095 gnd.n4103 gnd.t317 19.8005
R8096 gnd.n4102 gnd.t266 19.8005
R8097 gnd.n4102 gnd.t250 19.8005
R8098 gnd.n1470 gnd.n1469 19.5087
R8099 gnd.n1483 gnd.n1470 19.5087
R8100 gnd.n1481 gnd.n1472 19.5087
R8101 gnd.n4107 gnd.n4101 19.5087
R8102 gnd.t65 gnd.n5328 19.4385
R8103 gnd.n3199 gnd.n2399 19.3944
R8104 gnd.n2399 gnd.n2377 19.3944
R8105 gnd.n3224 gnd.n2377 19.3944
R8106 gnd.n3224 gnd.n2374 19.3944
R8107 gnd.n3231 gnd.n2374 19.3944
R8108 gnd.n3231 gnd.n2375 19.3944
R8109 gnd.n3227 gnd.n2375 19.3944
R8110 gnd.n3227 gnd.n2276 19.3944
R8111 gnd.n3261 gnd.n2276 19.3944
R8112 gnd.n3261 gnd.n2273 19.3944
R8113 gnd.n3266 gnd.n2273 19.3944
R8114 gnd.n3266 gnd.n2274 19.3944
R8115 gnd.n2274 gnd.n2265 19.3944
R8116 gnd.n3286 gnd.n2265 19.3944
R8117 gnd.n3286 gnd.n2262 19.3944
R8118 gnd.n3297 gnd.n2262 19.3944
R8119 gnd.n3297 gnd.n2263 19.3944
R8120 gnd.n3293 gnd.n2263 19.3944
R8121 gnd.n3293 gnd.n3292 19.3944
R8122 gnd.n3292 gnd.n2218 19.3944
R8123 gnd.n3372 gnd.n2218 19.3944
R8124 gnd.n3372 gnd.n2215 19.3944
R8125 gnd.n3395 gnd.n2215 19.3944
R8126 gnd.n3395 gnd.n2216 19.3944
R8127 gnd.n3391 gnd.n2216 19.3944
R8128 gnd.n3391 gnd.n3390 19.3944
R8129 gnd.n3390 gnd.n3389 19.3944
R8130 gnd.n3389 gnd.n3381 19.3944
R8131 gnd.n3385 gnd.n3381 19.3944
R8132 gnd.n3385 gnd.n3384 19.3944
R8133 gnd.n3384 gnd.n2168 19.3944
R8134 gnd.n2168 gnd.n2166 19.3944
R8135 gnd.n3474 gnd.n2166 19.3944
R8136 gnd.n3474 gnd.n2164 19.3944
R8137 gnd.n3478 gnd.n2164 19.3944
R8138 gnd.n3478 gnd.n2139 19.3944
R8139 gnd.n3524 gnd.n2139 19.3944
R8140 gnd.n3524 gnd.n2140 19.3944
R8141 gnd.n3520 gnd.n2140 19.3944
R8142 gnd.n3520 gnd.n2116 19.3944
R8143 gnd.n3583 gnd.n2116 19.3944
R8144 gnd.n3583 gnd.n2117 19.3944
R8145 gnd.n3579 gnd.n2117 19.3944
R8146 gnd.n3579 gnd.n3578 19.3944
R8147 gnd.n3578 gnd.n3577 19.3944
R8148 gnd.n3577 gnd.n3563 19.3944
R8149 gnd.n3573 gnd.n3563 19.3944
R8150 gnd.n3573 gnd.n3572 19.3944
R8151 gnd.n3572 gnd.n3571 19.3944
R8152 gnd.n3571 gnd.n2057 19.3944
R8153 gnd.n3691 gnd.n2057 19.3944
R8154 gnd.n3691 gnd.n2054 19.3944
R8155 gnd.n3696 gnd.n2054 19.3944
R8156 gnd.n3696 gnd.n2055 19.3944
R8157 gnd.n2055 gnd.n2028 19.3944
R8158 gnd.n3730 gnd.n2028 19.3944
R8159 gnd.n3730 gnd.n2025 19.3944
R8160 gnd.n3749 gnd.n2025 19.3944
R8161 gnd.n3749 gnd.n2026 19.3944
R8162 gnd.n3745 gnd.n2026 19.3944
R8163 gnd.n3745 gnd.n3744 19.3944
R8164 gnd.n3744 gnd.n3743 19.3944
R8165 gnd.n3743 gnd.n3738 19.3944
R8166 gnd.n3739 gnd.n3738 19.3944
R8167 gnd.n3739 gnd.n1972 19.3944
R8168 gnd.n3821 gnd.n1972 19.3944
R8169 gnd.n3821 gnd.n1969 19.3944
R8170 gnd.n3826 gnd.n1969 19.3944
R8171 gnd.n3826 gnd.n1970 19.3944
R8172 gnd.n1970 gnd.n1945 19.3944
R8173 gnd.n3863 gnd.n1945 19.3944
R8174 gnd.n3863 gnd.n1943 19.3944
R8175 gnd.n3867 gnd.n1943 19.3944
R8176 gnd.n3867 gnd.n1942 19.3944
R8177 gnd.n3874 gnd.n1942 19.3944
R8178 gnd.n3874 gnd.n1940 19.3944
R8179 gnd.n3878 gnd.n1940 19.3944
R8180 gnd.n3879 gnd.n3878 19.3944
R8181 gnd.n3882 gnd.n3879 19.3944
R8182 gnd.n3882 gnd.n1937 19.3944
R8183 gnd.n4064 gnd.n1937 19.3944
R8184 gnd.n4064 gnd.n1938 19.3944
R8185 gnd.n3183 gnd.n2401 19.3944
R8186 gnd.n3194 gnd.n2401 19.3944
R8187 gnd.n3195 gnd.n3194 19.3944
R8188 gnd.n3177 gnd.n3176 19.3944
R8189 gnd.n3176 gnd.n2942 19.3944
R8190 gnd.n3172 gnd.n2942 19.3944
R8191 gnd.n3172 gnd.n3171 19.3944
R8192 gnd.n3171 gnd.n3170 19.3944
R8193 gnd.n3170 gnd.n2947 19.3944
R8194 gnd.n3165 gnd.n2947 19.3944
R8195 gnd.n3165 gnd.n3164 19.3944
R8196 gnd.n3164 gnd.n3163 19.3944
R8197 gnd.n3163 gnd.n3066 19.3944
R8198 gnd.n3156 gnd.n3066 19.3944
R8199 gnd.n3156 gnd.n3155 19.3944
R8200 gnd.n3155 gnd.n3079 19.3944
R8201 gnd.n3148 gnd.n3079 19.3944
R8202 gnd.n3148 gnd.n3147 19.3944
R8203 gnd.n3147 gnd.n3089 19.3944
R8204 gnd.n3140 gnd.n3089 19.3944
R8205 gnd.n3140 gnd.n3139 19.3944
R8206 gnd.n3139 gnd.n3102 19.3944
R8207 gnd.n3132 gnd.n3102 19.3944
R8208 gnd.n3132 gnd.n3131 19.3944
R8209 gnd.n3131 gnd.n3112 19.3944
R8210 gnd.n3124 gnd.n3112 19.3944
R8211 gnd.n3124 gnd.n3123 19.3944
R8212 gnd.n3972 gnd.n3936 19.3944
R8213 gnd.n3985 gnd.n3936 19.3944
R8214 gnd.n3985 gnd.n3934 19.3944
R8215 gnd.n3991 gnd.n3934 19.3944
R8216 gnd.n3991 gnd.n3927 19.3944
R8217 gnd.n4004 gnd.n3927 19.3944
R8218 gnd.n4004 gnd.n3925 19.3944
R8219 gnd.n4010 gnd.n3925 19.3944
R8220 gnd.n4010 gnd.n3918 19.3944
R8221 gnd.n4023 gnd.n3918 19.3944
R8222 gnd.n4023 gnd.n3916 19.3944
R8223 gnd.n4029 gnd.n3916 19.3944
R8224 gnd.n4029 gnd.n3909 19.3944
R8225 gnd.n4043 gnd.n3909 19.3944
R8226 gnd.n4043 gnd.n3907 19.3944
R8227 gnd.n4049 gnd.n3907 19.3944
R8228 gnd.n5669 gnd.n5668 19.3944
R8229 gnd.n5668 gnd.n5578 19.3944
R8230 gnd.n5663 gnd.n5578 19.3944
R8231 gnd.n5663 gnd.n5662 19.3944
R8232 gnd.n5662 gnd.n5583 19.3944
R8233 gnd.n5657 gnd.n5583 19.3944
R8234 gnd.n5657 gnd.n5656 19.3944
R8235 gnd.n5656 gnd.n5655 19.3944
R8236 gnd.n5655 gnd.n5589 19.3944
R8237 gnd.n5649 gnd.n5589 19.3944
R8238 gnd.n5649 gnd.n5648 19.3944
R8239 gnd.n5648 gnd.n5647 19.3944
R8240 gnd.n5647 gnd.n5595 19.3944
R8241 gnd.n5641 gnd.n5595 19.3944
R8242 gnd.n5641 gnd.n5640 19.3944
R8243 gnd.n5640 gnd.n5639 19.3944
R8244 gnd.n5639 gnd.n5601 19.3944
R8245 gnd.n5633 gnd.n5601 19.3944
R8246 gnd.n5633 gnd.n5632 19.3944
R8247 gnd.n5632 gnd.n5631 19.3944
R8248 gnd.n5631 gnd.n5607 19.3944
R8249 gnd.n5625 gnd.n5607 19.3944
R8250 gnd.n5623 gnd.n5622 19.3944
R8251 gnd.n5622 gnd.n5617 19.3944
R8252 gnd.n5617 gnd.n5615 19.3944
R8253 gnd.n6466 gnd.n5243 19.3944
R8254 gnd.n6466 gnd.n6465 19.3944
R8255 gnd.n6465 gnd.n6464 19.3944
R8256 gnd.n6508 gnd.n6507 19.3944
R8257 gnd.n6507 gnd.n6506 19.3944
R8258 gnd.n6506 gnd.n5204 19.3944
R8259 gnd.n6501 gnd.n5204 19.3944
R8260 gnd.n6501 gnd.n6500 19.3944
R8261 gnd.n6500 gnd.n6499 19.3944
R8262 gnd.n6499 gnd.n5211 19.3944
R8263 gnd.n6494 gnd.n5211 19.3944
R8264 gnd.n6494 gnd.n6493 19.3944
R8265 gnd.n6493 gnd.n6492 19.3944
R8266 gnd.n6492 gnd.n5218 19.3944
R8267 gnd.n6487 gnd.n5218 19.3944
R8268 gnd.n6487 gnd.n6486 19.3944
R8269 gnd.n6486 gnd.n6485 19.3944
R8270 gnd.n6485 gnd.n5225 19.3944
R8271 gnd.n6480 gnd.n5225 19.3944
R8272 gnd.n6480 gnd.n6479 19.3944
R8273 gnd.n6479 gnd.n6478 19.3944
R8274 gnd.n6478 gnd.n5232 19.3944
R8275 gnd.n6473 gnd.n5232 19.3944
R8276 gnd.n6473 gnd.n6472 19.3944
R8277 gnd.n6472 gnd.n6471 19.3944
R8278 gnd.n5809 gnd.n5808 19.3944
R8279 gnd.n5810 gnd.n5809 19.3944
R8280 gnd.n5810 gnd.n5519 19.3944
R8281 gnd.n5519 gnd.n5513 19.3944
R8282 gnd.n5835 gnd.n5513 19.3944
R8283 gnd.n5836 gnd.n5835 19.3944
R8284 gnd.n5836 gnd.n5496 19.3944
R8285 gnd.n5496 gnd.n5494 19.3944
R8286 gnd.n5860 gnd.n5494 19.3944
R8287 gnd.n5863 gnd.n5860 19.3944
R8288 gnd.n5863 gnd.n5862 19.3944
R8289 gnd.n5862 gnd.n5466 19.3944
R8290 gnd.n5901 gnd.n5466 19.3944
R8291 gnd.n5901 gnd.n5464 19.3944
R8292 gnd.n5907 gnd.n5464 19.3944
R8293 gnd.n5908 gnd.n5907 19.3944
R8294 gnd.n5908 gnd.n5434 19.3944
R8295 gnd.n5958 gnd.n5434 19.3944
R8296 gnd.n5959 gnd.n5958 19.3944
R8297 gnd.n5959 gnd.n5427 19.3944
R8298 gnd.n5970 gnd.n5427 19.3944
R8299 gnd.n5971 gnd.n5970 19.3944
R8300 gnd.n5971 gnd.n5410 19.3944
R8301 gnd.n5410 gnd.n5408 19.3944
R8302 gnd.n5995 gnd.n5408 19.3944
R8303 gnd.n5996 gnd.n5995 19.3944
R8304 gnd.n5996 gnd.n5315 19.3944
R8305 gnd.n6043 gnd.n5315 19.3944
R8306 gnd.n6044 gnd.n6043 19.3944
R8307 gnd.n6044 gnd.n5308 19.3944
R8308 gnd.n6055 gnd.n5308 19.3944
R8309 gnd.n6056 gnd.n6055 19.3944
R8310 gnd.n6056 gnd.n5291 19.3944
R8311 gnd.n5291 gnd.n5289 19.3944
R8312 gnd.n6083 gnd.n5289 19.3944
R8313 gnd.n6083 gnd.n5272 19.3944
R8314 gnd.n6117 gnd.n5272 19.3944
R8315 gnd.n6118 gnd.n6117 19.3944
R8316 gnd.n6118 gnd.n5258 19.3944
R8317 gnd.n6144 gnd.n5258 19.3944
R8318 gnd.n6144 gnd.n5255 19.3944
R8319 gnd.n6148 gnd.n5255 19.3944
R8320 gnd.n6149 gnd.n6148 19.3944
R8321 gnd.n6435 gnd.n6149 19.3944
R8322 gnd.n6435 gnd.n6434 19.3944
R8323 gnd.n6434 gnd.n6433 19.3944
R8324 gnd.n6433 gnd.n6430 19.3944
R8325 gnd.n6430 gnd.n6429 19.3944
R8326 gnd.n6429 gnd.n6428 19.3944
R8327 gnd.n6428 gnd.n6425 19.3944
R8328 gnd.n6425 gnd.n6424 19.3944
R8329 gnd.n6424 gnd.n6421 19.3944
R8330 gnd.n6421 gnd.n6420 19.3944
R8331 gnd.n5792 gnd.n5791 19.3944
R8332 gnd.n5791 gnd.n5790 19.3944
R8333 gnd.n5790 gnd.n5789 19.3944
R8334 gnd.n5789 gnd.n5787 19.3944
R8335 gnd.n5787 gnd.n5784 19.3944
R8336 gnd.n5784 gnd.n5783 19.3944
R8337 gnd.n5783 gnd.n5780 19.3944
R8338 gnd.n5780 gnd.n5779 19.3944
R8339 gnd.n5779 gnd.n5776 19.3944
R8340 gnd.n5776 gnd.n5775 19.3944
R8341 gnd.n5775 gnd.n5772 19.3944
R8342 gnd.n5772 gnd.n5771 19.3944
R8343 gnd.n5771 gnd.n5768 19.3944
R8344 gnd.n5768 gnd.n5767 19.3944
R8345 gnd.n5818 gnd.n5524 19.3944
R8346 gnd.n5818 gnd.n5522 19.3944
R8347 gnd.n5822 gnd.n5522 19.3944
R8348 gnd.n5822 gnd.n5503 19.3944
R8349 gnd.n5848 gnd.n5503 19.3944
R8350 gnd.n5848 gnd.n5501 19.3944
R8351 gnd.n5854 gnd.n5501 19.3944
R8352 gnd.n5854 gnd.n5853 19.3944
R8353 gnd.n5853 gnd.n5477 19.3944
R8354 gnd.n5882 gnd.n5477 19.3944
R8355 gnd.n5882 gnd.n5475 19.3944
R8356 gnd.n5891 gnd.n5475 19.3944
R8357 gnd.n5891 gnd.n5890 19.3944
R8358 gnd.n5890 gnd.n5889 19.3944
R8359 gnd.n5889 gnd.n5444 19.3944
R8360 gnd.n5943 gnd.n5444 19.3944
R8361 gnd.n5943 gnd.n5442 19.3944
R8362 gnd.n5949 gnd.n5442 19.3944
R8363 gnd.n5949 gnd.n5948 19.3944
R8364 gnd.n5948 gnd.n5417 19.3944
R8365 gnd.n5983 gnd.n5417 19.3944
R8366 gnd.n5983 gnd.n5415 19.3944
R8367 gnd.n5989 gnd.n5415 19.3944
R8368 gnd.n5989 gnd.n5988 19.3944
R8369 gnd.n5988 gnd.n5326 19.3944
R8370 gnd.n6028 gnd.n5326 19.3944
R8371 gnd.n6028 gnd.n5324 19.3944
R8372 gnd.n6034 gnd.n5324 19.3944
R8373 gnd.n6034 gnd.n6033 19.3944
R8374 gnd.n6033 gnd.n5298 19.3944
R8375 gnd.n6067 gnd.n5298 19.3944
R8376 gnd.n6067 gnd.n5296 19.3944
R8377 gnd.n6076 gnd.n5296 19.3944
R8378 gnd.n6076 gnd.n6075 19.3944
R8379 gnd.n6075 gnd.n6074 19.3944
R8380 gnd.n6074 gnd.n5268 19.3944
R8381 gnd.n6124 gnd.n5268 19.3944
R8382 gnd.n6124 gnd.n5266 19.3944
R8383 gnd.n6134 gnd.n5266 19.3944
R8384 gnd.n6134 gnd.n6133 19.3944
R8385 gnd.n6133 gnd.n6132 19.3944
R8386 gnd.n6132 gnd.n984 19.3944
R8387 gnd.n6571 gnd.n984 19.3944
R8388 gnd.n6571 gnd.n6570 19.3944
R8389 gnd.n6570 gnd.n6569 19.3944
R8390 gnd.n6569 gnd.n988 19.3944
R8391 gnd.n1008 gnd.n988 19.3944
R8392 gnd.n6557 gnd.n1008 19.3944
R8393 gnd.n6557 gnd.n6556 19.3944
R8394 gnd.n6556 gnd.n6555 19.3944
R8395 gnd.n6555 gnd.n1014 19.3944
R8396 gnd.n5168 gnd.n1014 19.3944
R8397 gnd.n6543 gnd.n5168 19.3944
R8398 gnd.n6540 gnd.n6539 19.3944
R8399 gnd.n6539 gnd.n6538 19.3944
R8400 gnd.n6538 gnd.n5174 19.3944
R8401 gnd.n6533 gnd.n5174 19.3944
R8402 gnd.n6533 gnd.n6532 19.3944
R8403 gnd.n6532 gnd.n6531 19.3944
R8404 gnd.n6531 gnd.n5181 19.3944
R8405 gnd.n6526 gnd.n5181 19.3944
R8406 gnd.n6526 gnd.n6525 19.3944
R8407 gnd.n6525 gnd.n6524 19.3944
R8408 gnd.n6524 gnd.n5188 19.3944
R8409 gnd.n6519 gnd.n5188 19.3944
R8410 gnd.n6519 gnd.n6518 19.3944
R8411 gnd.n6518 gnd.n6517 19.3944
R8412 gnd.n5676 gnd.n5572 19.3944
R8413 gnd.n5680 gnd.n5572 19.3944
R8414 gnd.n5680 gnd.n5562 19.3944
R8415 gnd.n5692 gnd.n5562 19.3944
R8416 gnd.n5692 gnd.n5560 19.3944
R8417 gnd.n5696 gnd.n5560 19.3944
R8418 gnd.n5696 gnd.n5549 19.3944
R8419 gnd.n5708 gnd.n5549 19.3944
R8420 gnd.n5708 gnd.n5547 19.3944
R8421 gnd.n5734 gnd.n5547 19.3944
R8422 gnd.n5734 gnd.n5733 19.3944
R8423 gnd.n5733 gnd.n5732 19.3944
R8424 gnd.n5732 gnd.n5731 19.3944
R8425 gnd.n5731 gnd.n5729 19.3944
R8426 gnd.n5729 gnd.n5728 19.3944
R8427 gnd.n5728 gnd.n5726 19.3944
R8428 gnd.n5726 gnd.n5725 19.3944
R8429 gnd.n5725 gnd.n5723 19.3944
R8430 gnd.n5723 gnd.n5722 19.3944
R8431 gnd.n5722 gnd.n5484 19.3944
R8432 gnd.n5871 gnd.n5484 19.3944
R8433 gnd.n5871 gnd.n5482 19.3944
R8434 gnd.n5877 gnd.n5482 19.3944
R8435 gnd.n5877 gnd.n5876 19.3944
R8436 gnd.n5876 gnd.n5451 19.3944
R8437 gnd.n5918 gnd.n5451 19.3944
R8438 gnd.n5918 gnd.n5449 19.3944
R8439 gnd.n5922 gnd.n5449 19.3944
R8440 gnd.n5936 gnd.n5922 19.3944
R8441 gnd.n5934 gnd.n5933 19.3944
R8442 gnd.n5930 gnd.n5929 19.3944
R8443 gnd.n5926 gnd.n5925 19.3944
R8444 gnd.n6004 gnd.n5398 19.3944
R8445 gnd.n6004 gnd.n5332 19.3944
R8446 gnd.n6023 gnd.n5332 19.3944
R8447 gnd.n6023 gnd.n6022 19.3944
R8448 gnd.n6022 gnd.n6021 19.3944
R8449 gnd.n6021 gnd.n6019 19.3944
R8450 gnd.n6019 gnd.n6018 19.3944
R8451 gnd.n6018 gnd.n6016 19.3944
R8452 gnd.n6016 gnd.n6015 19.3944
R8453 gnd.n6015 gnd.n5280 19.3944
R8454 gnd.n6090 gnd.n5280 19.3944
R8455 gnd.n6090 gnd.n5278 19.3944
R8456 gnd.n6109 gnd.n5278 19.3944
R8457 gnd.n6109 gnd.n6108 19.3944
R8458 gnd.n6108 gnd.n6107 19.3944
R8459 gnd.n6107 gnd.n6106 19.3944
R8460 gnd.n6106 gnd.n6104 19.3944
R8461 gnd.n6104 gnd.n6103 19.3944
R8462 gnd.n6103 gnd.n6100 19.3944
R8463 gnd.n6100 gnd.n5253 19.3944
R8464 gnd.n6441 gnd.n5253 19.3944
R8465 gnd.n6441 gnd.n5251 19.3944
R8466 gnd.n6447 gnd.n5251 19.3944
R8467 gnd.n6448 gnd.n6447 19.3944
R8468 gnd.n6451 gnd.n6448 19.3944
R8469 gnd.n6451 gnd.n5249 19.3944
R8470 gnd.n6455 gnd.n5249 19.3944
R8471 gnd.n6458 gnd.n6455 19.3944
R8472 gnd.n6459 gnd.n6458 19.3944
R8473 gnd.n5672 gnd.n5568 19.3944
R8474 gnd.n5684 gnd.n5568 19.3944
R8475 gnd.n5684 gnd.n5566 19.3944
R8476 gnd.n5688 gnd.n5566 19.3944
R8477 gnd.n5688 gnd.n5556 19.3944
R8478 gnd.n5700 gnd.n5556 19.3944
R8479 gnd.n5700 gnd.n5554 19.3944
R8480 gnd.n5704 gnd.n5554 19.3944
R8481 gnd.n5704 gnd.n5543 19.3944
R8482 gnd.n5798 gnd.n5543 19.3944
R8483 gnd.n5798 gnd.n5540 19.3944
R8484 gnd.n5803 gnd.n5540 19.3944
R8485 gnd.n5803 gnd.n5531 19.3944
R8486 gnd.n5813 gnd.n5531 19.3944
R8487 gnd.n5813 gnd.n5515 19.3944
R8488 gnd.n5830 gnd.n5515 19.3944
R8489 gnd.n5830 gnd.n5511 19.3944
R8490 gnd.n5843 gnd.n5511 19.3944
R8491 gnd.n5843 gnd.n5842 19.3944
R8492 gnd.n5842 gnd.n5490 19.3944
R8493 gnd.n5867 gnd.n5490 19.3944
R8494 gnd.n5867 gnd.n5866 19.3944
R8495 gnd.n5866 gnd.n5468 19.3944
R8496 gnd.n5896 gnd.n5468 19.3944
R8497 gnd.n5896 gnd.n5458 19.3944
R8498 gnd.n5914 gnd.n5458 19.3944
R8499 gnd.n5914 gnd.n5913 19.3944
R8500 gnd.n5913 gnd.n5912 19.3944
R8501 gnd.n5912 gnd.n5436 19.3944
R8502 gnd.n5954 gnd.n5436 19.3944
R8503 gnd.n5954 gnd.n5429 19.3944
R8504 gnd.n5965 gnd.n5429 19.3944
R8505 gnd.n5965 gnd.n5425 19.3944
R8506 gnd.n5978 gnd.n5425 19.3944
R8507 gnd.n5978 gnd.n5977 19.3944
R8508 gnd.n5977 gnd.n5404 19.3944
R8509 gnd.n6000 gnd.n5404 19.3944
R8510 gnd.n6000 gnd.n5999 19.3944
R8511 gnd.n5999 gnd.n5317 19.3944
R8512 gnd.n6039 gnd.n5317 19.3944
R8513 gnd.n6039 gnd.n5310 19.3944
R8514 gnd.n6050 gnd.n5310 19.3944
R8515 gnd.n6050 gnd.n5306 19.3944
R8516 gnd.n6062 gnd.n5306 19.3944
R8517 gnd.n6062 gnd.n6061 19.3944
R8518 gnd.n6061 gnd.n5286 19.3944
R8519 gnd.n6086 gnd.n5286 19.3944
R8520 gnd.n6086 gnd.n5274 19.3944
R8521 gnd.n6113 gnd.n5274 19.3944
R8522 gnd.n6113 gnd.n5260 19.3944
R8523 gnd.n6139 gnd.n5260 19.3944
R8524 gnd.n6139 gnd.n973 19.3944
R8525 gnd.n6578 gnd.n973 19.3944
R8526 gnd.n6578 gnd.n6577 19.3944
R8527 gnd.n6577 gnd.n6576 19.3944
R8528 gnd.n6576 gnd.n977 19.3944
R8529 gnd.n996 gnd.n977 19.3944
R8530 gnd.n6564 gnd.n996 19.3944
R8531 gnd.n6564 gnd.n6563 19.3944
R8532 gnd.n6563 gnd.n6562 19.3944
R8533 gnd.n6562 gnd.n1000 19.3944
R8534 gnd.n1022 gnd.n1000 19.3944
R8535 gnd.n6550 gnd.n1022 19.3944
R8536 gnd.n6550 gnd.n6549 19.3944
R8537 gnd.n6549 gnd.n6548 19.3944
R8538 gnd.n3160 gnd.n3069 19.3944
R8539 gnd.n3160 gnd.n3159 19.3944
R8540 gnd.n3159 gnd.n3073 19.3944
R8541 gnd.n3152 gnd.n3073 19.3944
R8542 gnd.n3152 gnd.n3151 19.3944
R8543 gnd.n3151 gnd.n3085 19.3944
R8544 gnd.n3144 gnd.n3085 19.3944
R8545 gnd.n3144 gnd.n3143 19.3944
R8546 gnd.n3143 gnd.n3096 19.3944
R8547 gnd.n3136 gnd.n3096 19.3944
R8548 gnd.n3136 gnd.n3135 19.3944
R8549 gnd.n3135 gnd.n3108 19.3944
R8550 gnd.n3128 gnd.n3108 19.3944
R8551 gnd.n3128 gnd.n3127 19.3944
R8552 gnd.n3127 gnd.n2408 19.3944
R8553 gnd.n3186 gnd.n2408 19.3944
R8554 gnd.n7207 gnd.n527 19.3944
R8555 gnd.n7207 gnd.n523 19.3944
R8556 gnd.n7213 gnd.n523 19.3944
R8557 gnd.n7213 gnd.n521 19.3944
R8558 gnd.n7217 gnd.n521 19.3944
R8559 gnd.n7217 gnd.n517 19.3944
R8560 gnd.n7223 gnd.n517 19.3944
R8561 gnd.n7223 gnd.n515 19.3944
R8562 gnd.n7227 gnd.n515 19.3944
R8563 gnd.n7227 gnd.n511 19.3944
R8564 gnd.n7233 gnd.n511 19.3944
R8565 gnd.n7233 gnd.n509 19.3944
R8566 gnd.n7237 gnd.n509 19.3944
R8567 gnd.n7237 gnd.n505 19.3944
R8568 gnd.n7243 gnd.n505 19.3944
R8569 gnd.n7243 gnd.n503 19.3944
R8570 gnd.n7247 gnd.n503 19.3944
R8571 gnd.n7247 gnd.n499 19.3944
R8572 gnd.n7253 gnd.n499 19.3944
R8573 gnd.n7253 gnd.n497 19.3944
R8574 gnd.n7257 gnd.n497 19.3944
R8575 gnd.n7257 gnd.n493 19.3944
R8576 gnd.n7263 gnd.n493 19.3944
R8577 gnd.n7263 gnd.n491 19.3944
R8578 gnd.n7267 gnd.n491 19.3944
R8579 gnd.n7267 gnd.n487 19.3944
R8580 gnd.n7273 gnd.n487 19.3944
R8581 gnd.n7273 gnd.n485 19.3944
R8582 gnd.n7277 gnd.n485 19.3944
R8583 gnd.n7277 gnd.n481 19.3944
R8584 gnd.n7283 gnd.n481 19.3944
R8585 gnd.n7283 gnd.n479 19.3944
R8586 gnd.n7287 gnd.n479 19.3944
R8587 gnd.n7287 gnd.n475 19.3944
R8588 gnd.n7293 gnd.n475 19.3944
R8589 gnd.n7293 gnd.n473 19.3944
R8590 gnd.n7297 gnd.n473 19.3944
R8591 gnd.n7297 gnd.n469 19.3944
R8592 gnd.n7303 gnd.n469 19.3944
R8593 gnd.n7303 gnd.n467 19.3944
R8594 gnd.n7307 gnd.n467 19.3944
R8595 gnd.n7307 gnd.n463 19.3944
R8596 gnd.n7313 gnd.n463 19.3944
R8597 gnd.n7313 gnd.n461 19.3944
R8598 gnd.n7317 gnd.n461 19.3944
R8599 gnd.n7317 gnd.n457 19.3944
R8600 gnd.n7323 gnd.n457 19.3944
R8601 gnd.n7323 gnd.n455 19.3944
R8602 gnd.n7327 gnd.n455 19.3944
R8603 gnd.n7327 gnd.n451 19.3944
R8604 gnd.n7333 gnd.n451 19.3944
R8605 gnd.n7333 gnd.n449 19.3944
R8606 gnd.n7337 gnd.n449 19.3944
R8607 gnd.n7337 gnd.n445 19.3944
R8608 gnd.n7343 gnd.n445 19.3944
R8609 gnd.n7343 gnd.n443 19.3944
R8610 gnd.n7347 gnd.n443 19.3944
R8611 gnd.n7347 gnd.n439 19.3944
R8612 gnd.n7353 gnd.n439 19.3944
R8613 gnd.n7353 gnd.n437 19.3944
R8614 gnd.n7357 gnd.n437 19.3944
R8615 gnd.n7357 gnd.n433 19.3944
R8616 gnd.n7363 gnd.n433 19.3944
R8617 gnd.n7363 gnd.n431 19.3944
R8618 gnd.n7367 gnd.n431 19.3944
R8619 gnd.n7367 gnd.n427 19.3944
R8620 gnd.n7373 gnd.n427 19.3944
R8621 gnd.n7373 gnd.n425 19.3944
R8622 gnd.n7377 gnd.n425 19.3944
R8623 gnd.n7377 gnd.n421 19.3944
R8624 gnd.n7383 gnd.n421 19.3944
R8625 gnd.n7383 gnd.n419 19.3944
R8626 gnd.n7387 gnd.n419 19.3944
R8627 gnd.n7387 gnd.n415 19.3944
R8628 gnd.n7393 gnd.n415 19.3944
R8629 gnd.n7393 gnd.n413 19.3944
R8630 gnd.n7397 gnd.n413 19.3944
R8631 gnd.n7397 gnd.n409 19.3944
R8632 gnd.n7403 gnd.n409 19.3944
R8633 gnd.n7403 gnd.n407 19.3944
R8634 gnd.n7409 gnd.n407 19.3944
R8635 gnd.n7409 gnd.n7408 19.3944
R8636 gnd.n7408 gnd.n403 19.3944
R8637 gnd.n7416 gnd.n403 19.3944
R8638 gnd.n6753 gnd.n799 19.3944
R8639 gnd.n6753 gnd.n797 19.3944
R8640 gnd.n6757 gnd.n797 19.3944
R8641 gnd.n6757 gnd.n793 19.3944
R8642 gnd.n6763 gnd.n793 19.3944
R8643 gnd.n6763 gnd.n791 19.3944
R8644 gnd.n6767 gnd.n791 19.3944
R8645 gnd.n6767 gnd.n787 19.3944
R8646 gnd.n6773 gnd.n787 19.3944
R8647 gnd.n6773 gnd.n785 19.3944
R8648 gnd.n6777 gnd.n785 19.3944
R8649 gnd.n6777 gnd.n781 19.3944
R8650 gnd.n6783 gnd.n781 19.3944
R8651 gnd.n6783 gnd.n779 19.3944
R8652 gnd.n6787 gnd.n779 19.3944
R8653 gnd.n6787 gnd.n775 19.3944
R8654 gnd.n6793 gnd.n775 19.3944
R8655 gnd.n6793 gnd.n773 19.3944
R8656 gnd.n6797 gnd.n773 19.3944
R8657 gnd.n6797 gnd.n769 19.3944
R8658 gnd.n6803 gnd.n769 19.3944
R8659 gnd.n6803 gnd.n767 19.3944
R8660 gnd.n6807 gnd.n767 19.3944
R8661 gnd.n6807 gnd.n763 19.3944
R8662 gnd.n6813 gnd.n763 19.3944
R8663 gnd.n6813 gnd.n761 19.3944
R8664 gnd.n6817 gnd.n761 19.3944
R8665 gnd.n6817 gnd.n757 19.3944
R8666 gnd.n6823 gnd.n757 19.3944
R8667 gnd.n6823 gnd.n755 19.3944
R8668 gnd.n6827 gnd.n755 19.3944
R8669 gnd.n6827 gnd.n751 19.3944
R8670 gnd.n6833 gnd.n751 19.3944
R8671 gnd.n6833 gnd.n749 19.3944
R8672 gnd.n6837 gnd.n749 19.3944
R8673 gnd.n6837 gnd.n745 19.3944
R8674 gnd.n6843 gnd.n745 19.3944
R8675 gnd.n6843 gnd.n743 19.3944
R8676 gnd.n6847 gnd.n743 19.3944
R8677 gnd.n6847 gnd.n739 19.3944
R8678 gnd.n6853 gnd.n739 19.3944
R8679 gnd.n6853 gnd.n737 19.3944
R8680 gnd.n6857 gnd.n737 19.3944
R8681 gnd.n6857 gnd.n733 19.3944
R8682 gnd.n6863 gnd.n733 19.3944
R8683 gnd.n6863 gnd.n731 19.3944
R8684 gnd.n6867 gnd.n731 19.3944
R8685 gnd.n6867 gnd.n727 19.3944
R8686 gnd.n6873 gnd.n727 19.3944
R8687 gnd.n6873 gnd.n725 19.3944
R8688 gnd.n6877 gnd.n725 19.3944
R8689 gnd.n6877 gnd.n721 19.3944
R8690 gnd.n6883 gnd.n721 19.3944
R8691 gnd.n6883 gnd.n719 19.3944
R8692 gnd.n6887 gnd.n719 19.3944
R8693 gnd.n6887 gnd.n715 19.3944
R8694 gnd.n6893 gnd.n715 19.3944
R8695 gnd.n6893 gnd.n713 19.3944
R8696 gnd.n6897 gnd.n713 19.3944
R8697 gnd.n6897 gnd.n709 19.3944
R8698 gnd.n6903 gnd.n709 19.3944
R8699 gnd.n6903 gnd.n707 19.3944
R8700 gnd.n6907 gnd.n707 19.3944
R8701 gnd.n6907 gnd.n703 19.3944
R8702 gnd.n6913 gnd.n703 19.3944
R8703 gnd.n6913 gnd.n701 19.3944
R8704 gnd.n6917 gnd.n701 19.3944
R8705 gnd.n6917 gnd.n697 19.3944
R8706 gnd.n6923 gnd.n697 19.3944
R8707 gnd.n6923 gnd.n695 19.3944
R8708 gnd.n6927 gnd.n695 19.3944
R8709 gnd.n6927 gnd.n691 19.3944
R8710 gnd.n6933 gnd.n691 19.3944
R8711 gnd.n6933 gnd.n689 19.3944
R8712 gnd.n6937 gnd.n689 19.3944
R8713 gnd.n6937 gnd.n685 19.3944
R8714 gnd.n6943 gnd.n685 19.3944
R8715 gnd.n6943 gnd.n683 19.3944
R8716 gnd.n6947 gnd.n683 19.3944
R8717 gnd.n6947 gnd.n679 19.3944
R8718 gnd.n6953 gnd.n679 19.3944
R8719 gnd.n6953 gnd.n677 19.3944
R8720 gnd.n6957 gnd.n677 19.3944
R8721 gnd.n6957 gnd.n673 19.3944
R8722 gnd.n6963 gnd.n673 19.3944
R8723 gnd.n6963 gnd.n671 19.3944
R8724 gnd.n6967 gnd.n671 19.3944
R8725 gnd.n6967 gnd.n667 19.3944
R8726 gnd.n6973 gnd.n667 19.3944
R8727 gnd.n6973 gnd.n665 19.3944
R8728 gnd.n6977 gnd.n665 19.3944
R8729 gnd.n6977 gnd.n661 19.3944
R8730 gnd.n6983 gnd.n661 19.3944
R8731 gnd.n6983 gnd.n659 19.3944
R8732 gnd.n6987 gnd.n659 19.3944
R8733 gnd.n6987 gnd.n655 19.3944
R8734 gnd.n6993 gnd.n655 19.3944
R8735 gnd.n6993 gnd.n653 19.3944
R8736 gnd.n6997 gnd.n653 19.3944
R8737 gnd.n6997 gnd.n649 19.3944
R8738 gnd.n7003 gnd.n649 19.3944
R8739 gnd.n7003 gnd.n647 19.3944
R8740 gnd.n7007 gnd.n647 19.3944
R8741 gnd.n7007 gnd.n643 19.3944
R8742 gnd.n7013 gnd.n643 19.3944
R8743 gnd.n7013 gnd.n641 19.3944
R8744 gnd.n7017 gnd.n641 19.3944
R8745 gnd.n7017 gnd.n637 19.3944
R8746 gnd.n7023 gnd.n637 19.3944
R8747 gnd.n7023 gnd.n635 19.3944
R8748 gnd.n7027 gnd.n635 19.3944
R8749 gnd.n7027 gnd.n631 19.3944
R8750 gnd.n7033 gnd.n631 19.3944
R8751 gnd.n7033 gnd.n629 19.3944
R8752 gnd.n7037 gnd.n629 19.3944
R8753 gnd.n7037 gnd.n625 19.3944
R8754 gnd.n7043 gnd.n625 19.3944
R8755 gnd.n7043 gnd.n623 19.3944
R8756 gnd.n7047 gnd.n623 19.3944
R8757 gnd.n7047 gnd.n619 19.3944
R8758 gnd.n7053 gnd.n619 19.3944
R8759 gnd.n7053 gnd.n617 19.3944
R8760 gnd.n7057 gnd.n617 19.3944
R8761 gnd.n7057 gnd.n613 19.3944
R8762 gnd.n7063 gnd.n613 19.3944
R8763 gnd.n7063 gnd.n611 19.3944
R8764 gnd.n7067 gnd.n611 19.3944
R8765 gnd.n7067 gnd.n607 19.3944
R8766 gnd.n7073 gnd.n607 19.3944
R8767 gnd.n7073 gnd.n605 19.3944
R8768 gnd.n7077 gnd.n605 19.3944
R8769 gnd.n7077 gnd.n601 19.3944
R8770 gnd.n7083 gnd.n601 19.3944
R8771 gnd.n7083 gnd.n599 19.3944
R8772 gnd.n7087 gnd.n599 19.3944
R8773 gnd.n7087 gnd.n595 19.3944
R8774 gnd.n7093 gnd.n595 19.3944
R8775 gnd.n7093 gnd.n593 19.3944
R8776 gnd.n7097 gnd.n593 19.3944
R8777 gnd.n7097 gnd.n589 19.3944
R8778 gnd.n7103 gnd.n589 19.3944
R8779 gnd.n7103 gnd.n587 19.3944
R8780 gnd.n7107 gnd.n587 19.3944
R8781 gnd.n7107 gnd.n583 19.3944
R8782 gnd.n7113 gnd.n583 19.3944
R8783 gnd.n7113 gnd.n581 19.3944
R8784 gnd.n7117 gnd.n581 19.3944
R8785 gnd.n7117 gnd.n577 19.3944
R8786 gnd.n7123 gnd.n577 19.3944
R8787 gnd.n7123 gnd.n575 19.3944
R8788 gnd.n7127 gnd.n575 19.3944
R8789 gnd.n7127 gnd.n571 19.3944
R8790 gnd.n7133 gnd.n571 19.3944
R8791 gnd.n7133 gnd.n569 19.3944
R8792 gnd.n7137 gnd.n569 19.3944
R8793 gnd.n7137 gnd.n565 19.3944
R8794 gnd.n7143 gnd.n565 19.3944
R8795 gnd.n7143 gnd.n563 19.3944
R8796 gnd.n7147 gnd.n563 19.3944
R8797 gnd.n7147 gnd.n559 19.3944
R8798 gnd.n7153 gnd.n559 19.3944
R8799 gnd.n7153 gnd.n557 19.3944
R8800 gnd.n7157 gnd.n557 19.3944
R8801 gnd.n7157 gnd.n553 19.3944
R8802 gnd.n7163 gnd.n553 19.3944
R8803 gnd.n7163 gnd.n551 19.3944
R8804 gnd.n7167 gnd.n551 19.3944
R8805 gnd.n7167 gnd.n547 19.3944
R8806 gnd.n7173 gnd.n547 19.3944
R8807 gnd.n7173 gnd.n545 19.3944
R8808 gnd.n7177 gnd.n545 19.3944
R8809 gnd.n7177 gnd.n541 19.3944
R8810 gnd.n7183 gnd.n541 19.3944
R8811 gnd.n7183 gnd.n539 19.3944
R8812 gnd.n7187 gnd.n539 19.3944
R8813 gnd.n7187 gnd.n535 19.3944
R8814 gnd.n7193 gnd.n535 19.3944
R8815 gnd.n7193 gnd.n533 19.3944
R8816 gnd.n7197 gnd.n533 19.3944
R8817 gnd.n7197 gnd.n529 19.3944
R8818 gnd.n7203 gnd.n529 19.3944
R8819 gnd.n4278 gnd.n4275 19.3944
R8820 gnd.n4278 gnd.n4274 19.3944
R8821 gnd.n4284 gnd.n4274 19.3944
R8822 gnd.n4284 gnd.n4272 19.3944
R8823 gnd.n4288 gnd.n4272 19.3944
R8824 gnd.n4288 gnd.n4270 19.3944
R8825 gnd.n4294 gnd.n4270 19.3944
R8826 gnd.n4294 gnd.n4268 19.3944
R8827 gnd.n4298 gnd.n4268 19.3944
R8828 gnd.n4298 gnd.n4266 19.3944
R8829 gnd.n4304 gnd.n4266 19.3944
R8830 gnd.n4304 gnd.n4264 19.3944
R8831 gnd.n4308 gnd.n4264 19.3944
R8832 gnd.n4308 gnd.n4262 19.3944
R8833 gnd.n4314 gnd.n4262 19.3944
R8834 gnd.n4314 gnd.n4260 19.3944
R8835 gnd.n4321 gnd.n4260 19.3944
R8836 gnd.n4327 gnd.n4258 19.3944
R8837 gnd.n4327 gnd.n4256 19.3944
R8838 gnd.n4331 gnd.n4256 19.3944
R8839 gnd.n4331 gnd.n4254 19.3944
R8840 gnd.n4337 gnd.n4254 19.3944
R8841 gnd.n4337 gnd.n4252 19.3944
R8842 gnd.n4342 gnd.n4252 19.3944
R8843 gnd.n4350 gnd.n1860 19.3944
R8844 gnd.n4350 gnd.n1858 19.3944
R8845 gnd.n4354 gnd.n1858 19.3944
R8846 gnd.n4354 gnd.n1856 19.3944
R8847 gnd.n4360 gnd.n1856 19.3944
R8848 gnd.n4360 gnd.n1854 19.3944
R8849 gnd.n4364 gnd.n1854 19.3944
R8850 gnd.n4364 gnd.n1852 19.3944
R8851 gnd.n4376 gnd.n1850 19.3944
R8852 gnd.n4376 gnd.n1848 19.3944
R8853 gnd.n4382 gnd.n1848 19.3944
R8854 gnd.n4382 gnd.n1846 19.3944
R8855 gnd.n4386 gnd.n1846 19.3944
R8856 gnd.n4386 gnd.n1844 19.3944
R8857 gnd.n4392 gnd.n1844 19.3944
R8858 gnd.n4392 gnd.n1842 19.3944
R8859 gnd.n4396 gnd.n1842 19.3944
R8860 gnd.n4396 gnd.n1840 19.3944
R8861 gnd.n4402 gnd.n1840 19.3944
R8862 gnd.n4402 gnd.n1838 19.3944
R8863 gnd.n4406 gnd.n1838 19.3944
R8864 gnd.n4406 gnd.n1836 19.3944
R8865 gnd.n4412 gnd.n1836 19.3944
R8866 gnd.n4412 gnd.n1834 19.3944
R8867 gnd.n4417 gnd.n1834 19.3944
R8868 gnd.n4417 gnd.n1832 19.3944
R8869 gnd.n4430 gnd.n1825 19.3944
R8870 gnd.n4431 gnd.n4430 19.3944
R8871 gnd.n4432 gnd.n4431 19.3944
R8872 gnd.n4432 gnd.n1820 19.3944
R8873 gnd.n4444 gnd.n1820 19.3944
R8874 gnd.n4445 gnd.n4444 19.3944
R8875 gnd.n4446 gnd.n4445 19.3944
R8876 gnd.n4446 gnd.n1783 19.3944
R8877 gnd.n4458 gnd.n1783 19.3944
R8878 gnd.n4459 gnd.n4458 19.3944
R8879 gnd.n4460 gnd.n4459 19.3944
R8880 gnd.n4461 gnd.n4460 19.3944
R8881 gnd.n4465 gnd.n4461 19.3944
R8882 gnd.n4466 gnd.n4465 19.3944
R8883 gnd.n4470 gnd.n4466 19.3944
R8884 gnd.n4471 gnd.n4470 19.3944
R8885 gnd.n4473 gnd.n4471 19.3944
R8886 gnd.n4473 gnd.n1761 19.3944
R8887 gnd.n4518 gnd.n1761 19.3944
R8888 gnd.n4519 gnd.n4518 19.3944
R8889 gnd.n4544 gnd.n4519 19.3944
R8890 gnd.n4544 gnd.n4543 19.3944
R8891 gnd.n4543 gnd.n4542 19.3944
R8892 gnd.n4542 gnd.n4541 19.3944
R8893 gnd.n4541 gnd.n4540 19.3944
R8894 gnd.n4540 gnd.n4539 19.3944
R8895 gnd.n4539 gnd.n4523 19.3944
R8896 gnd.n4528 gnd.n4523 19.3944
R8897 gnd.n4528 gnd.n378 19.3944
R8898 gnd.n7448 gnd.n378 19.3944
R8899 gnd.n7449 gnd.n7448 19.3944
R8900 gnd.n7450 gnd.n7449 19.3944
R8901 gnd.n7450 gnd.n372 19.3944
R8902 gnd.n7462 gnd.n372 19.3944
R8903 gnd.n7463 gnd.n7462 19.3944
R8904 gnd.n7464 gnd.n7463 19.3944
R8905 gnd.n7464 gnd.n366 19.3944
R8906 gnd.n7476 gnd.n366 19.3944
R8907 gnd.n7477 gnd.n7476 19.3944
R8908 gnd.n7478 gnd.n7477 19.3944
R8909 gnd.n7478 gnd.n360 19.3944
R8910 gnd.n7491 gnd.n360 19.3944
R8911 gnd.n7492 gnd.n7491 19.3944
R8912 gnd.n7508 gnd.n7492 19.3944
R8913 gnd.n7508 gnd.n7507 19.3944
R8914 gnd.n7507 gnd.n7506 19.3944
R8915 gnd.n7506 gnd.n7504 19.3944
R8916 gnd.n7504 gnd.n7503 19.3944
R8917 gnd.n7503 gnd.n7501 19.3944
R8918 gnd.n7501 gnd.n7500 19.3944
R8919 gnd.n7500 gnd.n7498 19.3944
R8920 gnd.n7498 gnd.n7497 19.3944
R8921 gnd.n7497 gnd.n7495 19.3944
R8922 gnd.n4427 gnd.n1636 19.3944
R8923 gnd.n4639 gnd.n1636 19.3944
R8924 gnd.n4639 gnd.n4638 19.3944
R8925 gnd.n4638 gnd.n4637 19.3944
R8926 gnd.n4637 gnd.n1640 19.3944
R8927 gnd.n4627 gnd.n1640 19.3944
R8928 gnd.n4627 gnd.n4626 19.3944
R8929 gnd.n4626 gnd.n4625 19.3944
R8930 gnd.n4625 gnd.n1660 19.3944
R8931 gnd.n4615 gnd.n1660 19.3944
R8932 gnd.n4615 gnd.n4614 19.3944
R8933 gnd.n4614 gnd.n4613 19.3944
R8934 gnd.n4613 gnd.n1681 19.3944
R8935 gnd.n4603 gnd.n1681 19.3944
R8936 gnd.n4603 gnd.n4602 19.3944
R8937 gnd.n4602 gnd.n4601 19.3944
R8938 gnd.n4601 gnd.n1700 19.3944
R8939 gnd.n4591 gnd.n1700 19.3944
R8940 gnd.n4591 gnd.n4590 19.3944
R8941 gnd.n4590 gnd.n4589 19.3944
R8942 gnd.n4589 gnd.n1721 19.3944
R8943 gnd.n4579 gnd.n1721 19.3944
R8944 gnd.n4579 gnd.n4578 19.3944
R8945 gnd.n4578 gnd.n4577 19.3944
R8946 gnd.n4577 gnd.n1738 19.3944
R8947 gnd.n4526 gnd.n1738 19.3944
R8948 gnd.n4534 gnd.n4526 19.3944
R8949 gnd.n4534 gnd.n4533 19.3944
R8950 gnd.n4533 gnd.n4532 19.3944
R8951 gnd.n4532 gnd.n108 19.3944
R8952 gnd.n7739 gnd.n108 19.3944
R8953 gnd.n7739 gnd.n7738 19.3944
R8954 gnd.n7738 gnd.n7737 19.3944
R8955 gnd.n7737 gnd.n112 19.3944
R8956 gnd.n7727 gnd.n112 19.3944
R8957 gnd.n7727 gnd.n7726 19.3944
R8958 gnd.n7726 gnd.n7725 19.3944
R8959 gnd.n7725 gnd.n130 19.3944
R8960 gnd.n7715 gnd.n130 19.3944
R8961 gnd.n7715 gnd.n7714 19.3944
R8962 gnd.n7714 gnd.n7713 19.3944
R8963 gnd.n7713 gnd.n151 19.3944
R8964 gnd.n7703 gnd.n151 19.3944
R8965 gnd.n7703 gnd.n7702 19.3944
R8966 gnd.n7702 gnd.n7701 19.3944
R8967 gnd.n7701 gnd.n170 19.3944
R8968 gnd.n7691 gnd.n170 19.3944
R8969 gnd.n7691 gnd.n7690 19.3944
R8970 gnd.n7690 gnd.n7689 19.3944
R8971 gnd.n7689 gnd.n190 19.3944
R8972 gnd.n7679 gnd.n190 19.3944
R8973 gnd.n7679 gnd.n7678 19.3944
R8974 gnd.n7678 gnd.n7677 19.3944
R8975 gnd.n7599 gnd.n279 19.3944
R8976 gnd.n7599 gnd.n283 19.3944
R8977 gnd.n286 gnd.n283 19.3944
R8978 gnd.n7592 gnd.n286 19.3944
R8979 gnd.n7592 gnd.n7591 19.3944
R8980 gnd.n7591 gnd.n7590 19.3944
R8981 gnd.n7590 gnd.n292 19.3944
R8982 gnd.n7585 gnd.n292 19.3944
R8983 gnd.n7585 gnd.n7584 19.3944
R8984 gnd.n7584 gnd.n7583 19.3944
R8985 gnd.n7583 gnd.n299 19.3944
R8986 gnd.n7578 gnd.n299 19.3944
R8987 gnd.n7578 gnd.n7577 19.3944
R8988 gnd.n7577 gnd.n7576 19.3944
R8989 gnd.n7576 gnd.n306 19.3944
R8990 gnd.n7571 gnd.n306 19.3944
R8991 gnd.n7571 gnd.n7570 19.3944
R8992 gnd.n7570 gnd.n7569 19.3944
R8993 gnd.n7637 gnd.n246 19.3944
R8994 gnd.n7632 gnd.n246 19.3944
R8995 gnd.n7632 gnd.n7631 19.3944
R8996 gnd.n7631 gnd.n7630 19.3944
R8997 gnd.n7630 gnd.n253 19.3944
R8998 gnd.n7625 gnd.n253 19.3944
R8999 gnd.n7625 gnd.n7624 19.3944
R9000 gnd.n7624 gnd.n7623 19.3944
R9001 gnd.n7623 gnd.n260 19.3944
R9002 gnd.n7618 gnd.n260 19.3944
R9003 gnd.n7618 gnd.n7617 19.3944
R9004 gnd.n7617 gnd.n7616 19.3944
R9005 gnd.n7616 gnd.n267 19.3944
R9006 gnd.n7611 gnd.n267 19.3944
R9007 gnd.n7611 gnd.n7610 19.3944
R9008 gnd.n7610 gnd.n7609 19.3944
R9009 gnd.n7609 gnd.n274 19.3944
R9010 gnd.n7604 gnd.n274 19.3944
R9011 gnd.n7670 gnd.n7669 19.3944
R9012 gnd.n7669 gnd.n7668 19.3944
R9013 gnd.n7668 gnd.n218 19.3944
R9014 gnd.n7663 gnd.n218 19.3944
R9015 gnd.n7663 gnd.n7662 19.3944
R9016 gnd.n7662 gnd.n7661 19.3944
R9017 gnd.n7661 gnd.n225 19.3944
R9018 gnd.n7656 gnd.n225 19.3944
R9019 gnd.n7656 gnd.n7655 19.3944
R9020 gnd.n7655 gnd.n7654 19.3944
R9021 gnd.n7654 gnd.n232 19.3944
R9022 gnd.n7649 gnd.n232 19.3944
R9023 gnd.n7649 gnd.n7648 19.3944
R9024 gnd.n7648 gnd.n7647 19.3944
R9025 gnd.n7647 gnd.n239 19.3944
R9026 gnd.n7642 gnd.n239 19.3944
R9027 gnd.n7642 gnd.n7641 19.3944
R9028 gnd.n7560 gnd.n7559 19.3944
R9029 gnd.n7559 gnd.n7558 19.3944
R9030 gnd.n7558 gnd.n321 19.3944
R9031 gnd.n7553 gnd.n321 19.3944
R9032 gnd.n7553 gnd.n7552 19.3944
R9033 gnd.n7552 gnd.n7551 19.3944
R9034 gnd.n7551 gnd.n328 19.3944
R9035 gnd.n7546 gnd.n328 19.3944
R9036 gnd.n7546 gnd.n7545 19.3944
R9037 gnd.n7545 gnd.n7544 19.3944
R9038 gnd.n7544 gnd.n335 19.3944
R9039 gnd.n7539 gnd.n335 19.3944
R9040 gnd.n7539 gnd.n7538 19.3944
R9041 gnd.n7538 gnd.n7537 19.3944
R9042 gnd.n7537 gnd.n342 19.3944
R9043 gnd.n7532 gnd.n342 19.3944
R9044 gnd.n3889 gnd.n3888 19.3944
R9045 gnd.n3888 gnd.n1824 19.3944
R9046 gnd.n4436 gnd.n1824 19.3944
R9047 gnd.n4436 gnd.n1822 19.3944
R9048 gnd.n4440 gnd.n1822 19.3944
R9049 gnd.n4440 gnd.n1787 19.3944
R9050 gnd.n4450 gnd.n1787 19.3944
R9051 gnd.n4450 gnd.n1785 19.3944
R9052 gnd.n4454 gnd.n1785 19.3944
R9053 gnd.n4454 gnd.n1775 19.3944
R9054 gnd.n4490 gnd.n1775 19.3944
R9055 gnd.n4490 gnd.n1776 19.3944
R9056 gnd.n4486 gnd.n1776 19.3944
R9057 gnd.n4486 gnd.n4485 19.3944
R9058 gnd.n4485 gnd.n4484 19.3944
R9059 gnd.n4484 gnd.n1781 19.3944
R9060 gnd.n4480 gnd.n1781 19.3944
R9061 gnd.n4480 gnd.n4479 19.3944
R9062 gnd.n4479 gnd.n4478 19.3944
R9063 gnd.n4478 gnd.n1760 19.3944
R9064 gnd.n4548 gnd.n1760 19.3944
R9065 gnd.n4548 gnd.n1757 19.3944
R9066 gnd.n4555 gnd.n1757 19.3944
R9067 gnd.n4555 gnd.n1758 19.3944
R9068 gnd.n4551 gnd.n1758 19.3944
R9069 gnd.n4551 gnd.n81 19.3944
R9070 gnd.n7752 gnd.n81 19.3944
R9071 gnd.n7752 gnd.n7751 19.3944
R9072 gnd.n7751 gnd.n83 19.3944
R9073 gnd.n7444 gnd.n83 19.3944
R9074 gnd.n7444 gnd.n377 19.3944
R9075 gnd.n7454 gnd.n377 19.3944
R9076 gnd.n7454 gnd.n375 19.3944
R9077 gnd.n7458 gnd.n375 19.3944
R9078 gnd.n7458 gnd.n370 19.3944
R9079 gnd.n7468 gnd.n370 19.3944
R9080 gnd.n7468 gnd.n368 19.3944
R9081 gnd.n7472 gnd.n368 19.3944
R9082 gnd.n7472 gnd.n365 19.3944
R9083 gnd.n7482 gnd.n365 19.3944
R9084 gnd.n7482 gnd.n363 19.3944
R9085 gnd.n7487 gnd.n363 19.3944
R9086 gnd.n7487 gnd.n359 19.3944
R9087 gnd.n7512 gnd.n359 19.3944
R9088 gnd.n7513 gnd.n7512 19.3944
R9089 gnd.n7513 gnd.n357 19.3944
R9090 gnd.n7517 gnd.n357 19.3944
R9091 gnd.n7519 gnd.n7517 19.3944
R9092 gnd.n7520 gnd.n7519 19.3944
R9093 gnd.n7520 gnd.n354 19.3944
R9094 gnd.n7524 gnd.n354 19.3944
R9095 gnd.n7526 gnd.n7524 19.3944
R9096 gnd.n7527 gnd.n7526 19.3944
R9097 gnd.n4645 gnd.n4644 19.3944
R9098 gnd.n4644 gnd.n4643 19.3944
R9099 gnd.n4643 gnd.n1628 19.3944
R9100 gnd.n4633 gnd.n1628 19.3944
R9101 gnd.n4633 gnd.n4632 19.3944
R9102 gnd.n4632 gnd.n4631 19.3944
R9103 gnd.n4631 gnd.n1651 19.3944
R9104 gnd.n4621 gnd.n1651 19.3944
R9105 gnd.n4621 gnd.n4620 19.3944
R9106 gnd.n4620 gnd.n4619 19.3944
R9107 gnd.n4619 gnd.n1671 19.3944
R9108 gnd.n4609 gnd.n1671 19.3944
R9109 gnd.n4609 gnd.n4608 19.3944
R9110 gnd.n4608 gnd.n4607 19.3944
R9111 gnd.n4607 gnd.n1691 19.3944
R9112 gnd.n4597 gnd.n1691 19.3944
R9113 gnd.n4597 gnd.n4596 19.3944
R9114 gnd.n4596 gnd.n4595 19.3944
R9115 gnd.n4595 gnd.n1711 19.3944
R9116 gnd.n4585 gnd.n1711 19.3944
R9117 gnd.n4585 gnd.n4584 19.3944
R9118 gnd.n4584 gnd.n4583 19.3944
R9119 gnd.n1729 gnd.n97 19.3944
R9120 gnd.n1747 gnd.n97 19.3944
R9121 gnd.n1745 gnd.n1744 19.3944
R9122 gnd.n7747 gnd.n7746 19.3944
R9123 gnd.n7743 gnd.n92 19.3944
R9124 gnd.n7743 gnd.n99 19.3944
R9125 gnd.n7733 gnd.n99 19.3944
R9126 gnd.n7733 gnd.n7732 19.3944
R9127 gnd.n7732 gnd.n7731 19.3944
R9128 gnd.n7731 gnd.n121 19.3944
R9129 gnd.n7721 gnd.n121 19.3944
R9130 gnd.n7721 gnd.n7720 19.3944
R9131 gnd.n7720 gnd.n7719 19.3944
R9132 gnd.n7719 gnd.n141 19.3944
R9133 gnd.n7709 gnd.n141 19.3944
R9134 gnd.n7709 gnd.n7708 19.3944
R9135 gnd.n7708 gnd.n7707 19.3944
R9136 gnd.n7707 gnd.n161 19.3944
R9137 gnd.n7697 gnd.n161 19.3944
R9138 gnd.n7697 gnd.n7696 19.3944
R9139 gnd.n7696 gnd.n7695 19.3944
R9140 gnd.n7695 gnd.n181 19.3944
R9141 gnd.n7685 gnd.n181 19.3944
R9142 gnd.n7685 gnd.n7684 19.3944
R9143 gnd.n7684 gnd.n7683 19.3944
R9144 gnd.n7683 gnd.n200 19.3944
R9145 gnd.n7673 gnd.n200 19.3944
R9146 gnd.n2653 gnd.n2647 19.3944
R9147 gnd.n2657 gnd.n2647 19.3944
R9148 gnd.n2657 gnd.n2645 19.3944
R9149 gnd.n2679 gnd.n2645 19.3944
R9150 gnd.n2679 gnd.n2678 19.3944
R9151 gnd.n2678 gnd.n2677 19.3944
R9152 gnd.n2677 gnd.n2663 19.3944
R9153 gnd.n2673 gnd.n2663 19.3944
R9154 gnd.n2673 gnd.n2672 19.3944
R9155 gnd.n2672 gnd.n2671 19.3944
R9156 gnd.n2671 gnd.n2501 19.3944
R9157 gnd.n2726 gnd.n2501 19.3944
R9158 gnd.n2729 gnd.n2728 19.3944
R9159 gnd.n2733 gnd.n2732 19.3944
R9160 gnd.n2738 gnd.n2737 19.3944
R9161 gnd.n2735 gnd.n2459 19.3944
R9162 gnd.n2807 gnd.n2456 19.3944
R9163 gnd.n2807 gnd.n2455 19.3944
R9164 gnd.n2811 gnd.n2455 19.3944
R9165 gnd.n2811 gnd.n2453 19.3944
R9166 gnd.n2815 gnd.n2453 19.3944
R9167 gnd.n2815 gnd.n2451 19.3944
R9168 gnd.n2838 gnd.n2451 19.3944
R9169 gnd.n2838 gnd.n2837 19.3944
R9170 gnd.n2837 gnd.n2836 19.3944
R9171 gnd.n2836 gnd.n2821 19.3944
R9172 gnd.n2832 gnd.n2821 19.3944
R9173 gnd.n2832 gnd.n2831 19.3944
R9174 gnd.n2831 gnd.n2830 19.3944
R9175 gnd.n2830 gnd.n2828 19.3944
R9176 gnd.n2828 gnd.n2428 19.3944
R9177 gnd.n2902 gnd.n2428 19.3944
R9178 gnd.n2902 gnd.n2426 19.3944
R9179 gnd.n2906 gnd.n2426 19.3944
R9180 gnd.n2906 gnd.n2424 19.3944
R9181 gnd.n2910 gnd.n2424 19.3944
R9182 gnd.n2910 gnd.n2422 19.3944
R9183 gnd.n2914 gnd.n2422 19.3944
R9184 gnd.n2914 gnd.n2420 19.3944
R9185 gnd.n2920 gnd.n2420 19.3944
R9186 gnd.n2920 gnd.n2418 19.3944
R9187 gnd.n2924 gnd.n2418 19.3944
R9188 gnd.n2924 gnd.n2395 19.3944
R9189 gnd.n3204 gnd.n2395 19.3944
R9190 gnd.n3204 gnd.n2393 19.3944
R9191 gnd.n3210 gnd.n2393 19.3944
R9192 gnd.n3210 gnd.n3209 19.3944
R9193 gnd.n3209 gnd.n2370 19.3944
R9194 gnd.n3236 gnd.n2370 19.3944
R9195 gnd.n3236 gnd.n2368 19.3944
R9196 gnd.n3243 gnd.n2368 19.3944
R9197 gnd.n3243 gnd.n3242 19.3944
R9198 gnd.n3242 gnd.n1496 19.3944
R9199 gnd.n4778 gnd.n1496 19.3944
R9200 gnd.n4778 gnd.n4777 19.3944
R9201 gnd.n4777 gnd.n4776 19.3944
R9202 gnd.n4776 gnd.n1500 19.3944
R9203 gnd.n3279 gnd.n1500 19.3944
R9204 gnd.n3279 gnd.n2244 19.3944
R9205 gnd.n3318 gnd.n2244 19.3944
R9206 gnd.n3318 gnd.n2242 19.3944
R9207 gnd.n3322 gnd.n2242 19.3944
R9208 gnd.n3322 gnd.n2226 19.3944
R9209 gnd.n3360 gnd.n2226 19.3944
R9210 gnd.n3360 gnd.n2224 19.3944
R9211 gnd.n3366 gnd.n2224 19.3944
R9212 gnd.n3366 gnd.n3365 19.3944
R9213 gnd.n3365 gnd.n2200 19.3944
R9214 gnd.n3422 gnd.n2200 19.3944
R9215 gnd.n3422 gnd.n2198 19.3944
R9216 gnd.n3426 gnd.n2198 19.3944
R9217 gnd.n3426 gnd.n2182 19.3944
R9218 gnd.n3450 gnd.n2182 19.3944
R9219 gnd.n3450 gnd.n2180 19.3944
R9220 gnd.n3456 gnd.n2180 19.3944
R9221 gnd.n3456 gnd.n3455 19.3944
R9222 gnd.n3455 gnd.n2149 19.3944
R9223 gnd.n3500 gnd.n2149 19.3944
R9224 gnd.n3500 gnd.n2147 19.3944
R9225 gnd.n3504 gnd.n2147 19.3944
R9226 gnd.n3504 gnd.n2126 19.3944
R9227 gnd.n3540 gnd.n2126 19.3944
R9228 gnd.n3540 gnd.n2124 19.3944
R9229 gnd.n3544 gnd.n2124 19.3944
R9230 gnd.n3544 gnd.n2104 19.3944
R9231 gnd.n3597 gnd.n2104 19.3944
R9232 gnd.n3597 gnd.n2102 19.3944
R9233 gnd.n3601 gnd.n2102 19.3944
R9234 gnd.n3601 gnd.n2084 19.3944
R9235 gnd.n3622 gnd.n2084 19.3944
R9236 gnd.n3622 gnd.n2082 19.3944
R9237 gnd.n3626 gnd.n2082 19.3944
R9238 gnd.n3626 gnd.n2064 19.3944
R9239 gnd.n3682 gnd.n2064 19.3944
R9240 gnd.n3682 gnd.n2062 19.3944
R9241 gnd.n3686 gnd.n2062 19.3944
R9242 gnd.n3686 gnd.n2042 19.3944
R9243 gnd.n3711 gnd.n2042 19.3944
R9244 gnd.n3711 gnd.n2040 19.3944
R9245 gnd.n3717 gnd.n2040 19.3944
R9246 gnd.n3717 gnd.n3716 19.3944
R9247 gnd.n3716 gnd.n2014 19.3944
R9248 gnd.n3762 gnd.n2014 19.3944
R9249 gnd.n3762 gnd.n2012 19.3944
R9250 gnd.n3766 gnd.n2012 19.3944
R9251 gnd.n3766 gnd.n1994 19.3944
R9252 gnd.n3788 gnd.n1994 19.3944
R9253 gnd.n3788 gnd.n1992 19.3944
R9254 gnd.n3794 gnd.n1992 19.3944
R9255 gnd.n3794 gnd.n3793 19.3944
R9256 gnd.n3793 gnd.n1964 19.3944
R9257 gnd.n3832 gnd.n1964 19.3944
R9258 gnd.n3832 gnd.n1962 19.3944
R9259 gnd.n3839 gnd.n1962 19.3944
R9260 gnd.n3839 gnd.n3838 19.3944
R9261 gnd.n3838 gnd.n1913 19.3944
R9262 gnd.n4085 gnd.n1913 19.3944
R9263 gnd.n4085 gnd.n4084 19.3944
R9264 gnd.n4084 gnd.n4083 19.3944
R9265 gnd.n4083 gnd.n1917 19.3944
R9266 gnd.n1924 gnd.n1917 19.3944
R9267 gnd.n4073 gnd.n1924 19.3944
R9268 gnd.n4073 gnd.n4072 19.3944
R9269 gnd.n4072 gnd.n4071 19.3944
R9270 gnd.n4071 gnd.n1932 19.3944
R9271 gnd.n1932 gnd.n1603 19.3944
R9272 gnd.n4660 gnd.n1603 19.3944
R9273 gnd.n4660 gnd.n4659 19.3944
R9274 gnd.n4659 gnd.n4658 19.3944
R9275 gnd.n4658 gnd.n1607 19.3944
R9276 gnd.n4652 gnd.n1607 19.3944
R9277 gnd.n4652 gnd.n4651 19.3944
R9278 gnd.n4651 gnd.n4650 19.3944
R9279 gnd.n4650 gnd.n1616 19.3944
R9280 gnd.n1794 gnd.n1616 19.3944
R9281 gnd.n1798 gnd.n1794 19.3944
R9282 gnd.n1798 gnd.n1792 19.3944
R9283 gnd.n1802 gnd.n1792 19.3944
R9284 gnd.n1802 gnd.n1790 19.3944
R9285 gnd.n1817 gnd.n1790 19.3944
R9286 gnd.n1817 gnd.n1816 19.3944
R9287 gnd.n1816 gnd.n1815 19.3944
R9288 gnd.n1815 gnd.n1812 19.3944
R9289 gnd.n1812 gnd.n1811 19.3944
R9290 gnd.n1811 gnd.n1773 19.3944
R9291 gnd.n1773 gnd.n1771 19.3944
R9292 gnd.n4497 gnd.n1771 19.3944
R9293 gnd.n4497 gnd.n1769 19.3944
R9294 gnd.n4501 gnd.n1769 19.3944
R9295 gnd.n4501 gnd.n1767 19.3944
R9296 gnd.n4505 gnd.n1767 19.3944
R9297 gnd.n4505 gnd.n1765 19.3944
R9298 gnd.n4513 gnd.n1765 19.3944
R9299 gnd.n4513 gnd.n4512 19.3944
R9300 gnd.n4512 gnd.n4511 19.3944
R9301 gnd.n4561 gnd.n1754 19.3944
R9302 gnd.n4569 gnd.n4563 19.3944
R9303 gnd.n4567 gnd.n4566 19.3944
R9304 gnd.n7439 gnd.n384 19.3944
R9305 gnd.n7437 gnd.n7436 19.3944
R9306 gnd.n7436 gnd.n386 19.3944
R9307 gnd.n7432 gnd.n386 19.3944
R9308 gnd.n7432 gnd.n7431 19.3944
R9309 gnd.n7431 gnd.n7430 19.3944
R9310 gnd.n7430 gnd.n392 19.3944
R9311 gnd.n7426 gnd.n392 19.3944
R9312 gnd.n7426 gnd.n7425 19.3944
R9313 gnd.n7425 gnd.n7424 19.3944
R9314 gnd.n7424 gnd.n398 19.3944
R9315 gnd.n7420 gnd.n398 19.3944
R9316 gnd.n7420 gnd.n7419 19.3944
R9317 gnd.n5161 gnd.n5160 19.3944
R9318 gnd.n5160 gnd.n5159 19.3944
R9319 gnd.n5159 gnd.n5158 19.3944
R9320 gnd.n5158 gnd.n5156 19.3944
R9321 gnd.n5156 gnd.n5153 19.3944
R9322 gnd.n5153 gnd.n5152 19.3944
R9323 gnd.n5152 gnd.n5149 19.3944
R9324 gnd.n5149 gnd.n5148 19.3944
R9325 gnd.n5148 gnd.n5145 19.3944
R9326 gnd.n5145 gnd.n5144 19.3944
R9327 gnd.n5144 gnd.n5141 19.3944
R9328 gnd.n5141 gnd.n5140 19.3944
R9329 gnd.n5140 gnd.n5137 19.3944
R9330 gnd.n5137 gnd.n5136 19.3944
R9331 gnd.n5136 gnd.n5133 19.3944
R9332 gnd.n5133 gnd.n5132 19.3944
R9333 gnd.n5132 gnd.n5129 19.3944
R9334 gnd.n5127 gnd.n5124 19.3944
R9335 gnd.n5124 gnd.n5123 19.3944
R9336 gnd.n5123 gnd.n5120 19.3944
R9337 gnd.n5120 gnd.n5119 19.3944
R9338 gnd.n5119 gnd.n5116 19.3944
R9339 gnd.n5116 gnd.n5115 19.3944
R9340 gnd.n5115 gnd.n5112 19.3944
R9341 gnd.n5112 gnd.n5111 19.3944
R9342 gnd.n5111 gnd.n5108 19.3944
R9343 gnd.n5108 gnd.n5107 19.3944
R9344 gnd.n5107 gnd.n5104 19.3944
R9345 gnd.n5104 gnd.n5103 19.3944
R9346 gnd.n5103 gnd.n5100 19.3944
R9347 gnd.n5100 gnd.n5099 19.3944
R9348 gnd.n5099 gnd.n5096 19.3944
R9349 gnd.n5096 gnd.n5095 19.3944
R9350 gnd.n5095 gnd.n5092 19.3944
R9351 gnd.n5092 gnd.n5091 19.3944
R9352 gnd.n5087 gnd.n5084 19.3944
R9353 gnd.n5084 gnd.n5083 19.3944
R9354 gnd.n5083 gnd.n5080 19.3944
R9355 gnd.n5080 gnd.n5079 19.3944
R9356 gnd.n5079 gnd.n5076 19.3944
R9357 gnd.n5076 gnd.n5075 19.3944
R9358 gnd.n5075 gnd.n5072 19.3944
R9359 gnd.n5072 gnd.n5071 19.3944
R9360 gnd.n5071 gnd.n5068 19.3944
R9361 gnd.n5068 gnd.n5067 19.3944
R9362 gnd.n5067 gnd.n5064 19.3944
R9363 gnd.n5064 gnd.n5063 19.3944
R9364 gnd.n5063 gnd.n5060 19.3944
R9365 gnd.n5060 gnd.n5059 19.3944
R9366 gnd.n5059 gnd.n5056 19.3944
R9367 gnd.n5056 gnd.n5055 19.3944
R9368 gnd.n5055 gnd.n5052 19.3944
R9369 gnd.n5052 gnd.n5051 19.3944
R9370 gnd.n2565 gnd.n2564 19.3944
R9371 gnd.n2568 gnd.n2565 19.3944
R9372 gnd.n2568 gnd.n2560 19.3944
R9373 gnd.n2574 gnd.n2560 19.3944
R9374 gnd.n2575 gnd.n2574 19.3944
R9375 gnd.n2578 gnd.n2575 19.3944
R9376 gnd.n2578 gnd.n2558 19.3944
R9377 gnd.n2584 gnd.n2558 19.3944
R9378 gnd.n2585 gnd.n2584 19.3944
R9379 gnd.n2588 gnd.n2585 19.3944
R9380 gnd.n2588 gnd.n2556 19.3944
R9381 gnd.n2594 gnd.n2556 19.3944
R9382 gnd.n2595 gnd.n2594 19.3944
R9383 gnd.n2598 gnd.n2595 19.3944
R9384 gnd.n2598 gnd.n2552 19.3944
R9385 gnd.n2602 gnd.n2552 19.3944
R9386 gnd.n2607 gnd.n2547 19.3944
R9387 gnd.n2612 gnd.n2547 19.3944
R9388 gnd.n2613 gnd.n2612 19.3944
R9389 gnd.n2615 gnd.n2613 19.3944
R9390 gnd.n2615 gnd.n2545 19.3944
R9391 gnd.n2620 gnd.n2545 19.3944
R9392 gnd.n2621 gnd.n2620 19.3944
R9393 gnd.n2623 gnd.n2621 19.3944
R9394 gnd.n2623 gnd.n2543 19.3944
R9395 gnd.n2627 gnd.n2543 19.3944
R9396 gnd.n2627 gnd.n2528 19.3944
R9397 gnd.n2637 gnd.n2528 19.3944
R9398 gnd.n2637 gnd.n2526 19.3944
R9399 gnd.n2641 gnd.n2526 19.3944
R9400 gnd.n2641 gnd.n2523 19.3944
R9401 gnd.n2690 gnd.n2523 19.3944
R9402 gnd.n2690 gnd.n2521 19.3944
R9403 gnd.n2695 gnd.n2521 19.3944
R9404 gnd.n2695 gnd.n2517 19.3944
R9405 gnd.n2706 gnd.n2517 19.3944
R9406 gnd.n2707 gnd.n2706 19.3944
R9407 gnd.n2709 gnd.n2707 19.3944
R9408 gnd.n2709 gnd.n2515 19.3944
R9409 gnd.n2713 gnd.n2515 19.3944
R9410 gnd.n2713 gnd.n2481 19.3944
R9411 gnd.n2754 gnd.n2481 19.3944
R9412 gnd.n2754 gnd.n2479 19.3944
R9413 gnd.n2759 gnd.n2479 19.3944
R9414 gnd.n2759 gnd.n2463 19.3944
R9415 gnd.n2800 gnd.n2463 19.3944
R9416 gnd.n2800 gnd.n2464 19.3944
R9417 gnd.n2796 gnd.n2464 19.3944
R9418 gnd.n2796 gnd.n2795 19.3944
R9419 gnd.n2795 gnd.n2794 19.3944
R9420 gnd.n2794 gnd.n2469 19.3944
R9421 gnd.n2790 gnd.n2469 19.3944
R9422 gnd.n2790 gnd.n2447 19.3944
R9423 gnd.n2843 gnd.n2447 19.3944
R9424 gnd.n2843 gnd.n2445 19.3944
R9425 gnd.n2847 gnd.n2445 19.3944
R9426 gnd.n2847 gnd.n2442 19.3944
R9427 gnd.n2858 gnd.n2442 19.3944
R9428 gnd.n2858 gnd.n2440 19.3944
R9429 gnd.n2862 gnd.n2440 19.3944
R9430 gnd.n2862 gnd.n2431 19.3944
R9431 gnd.n2896 gnd.n2431 19.3944
R9432 gnd.n2896 gnd.n2432 19.3944
R9433 gnd.n2892 gnd.n2432 19.3944
R9434 gnd.n2892 gnd.n2891 19.3944
R9435 gnd.n2891 gnd.n2890 19.3944
R9436 gnd.n2890 gnd.n2437 19.3944
R9437 gnd.n2886 gnd.n2437 19.3944
R9438 gnd.n2886 gnd.n2885 19.3944
R9439 gnd.n5043 gnd.n1139 19.3944
R9440 gnd.n2530 gnd.n1139 19.3944
R9441 gnd.n2531 gnd.n2530 19.3944
R9442 gnd.n2533 gnd.n2531 19.3944
R9443 gnd.n2534 gnd.n2533 19.3944
R9444 gnd.n2537 gnd.n2534 19.3944
R9445 gnd.n2538 gnd.n2537 19.3944
R9446 gnd.n2540 gnd.n2538 19.3944
R9447 gnd.n2541 gnd.n2540 19.3944
R9448 gnd.n2631 gnd.n2541 19.3944
R9449 gnd.n2632 gnd.n2631 19.3944
R9450 gnd.n2633 gnd.n2632 19.3944
R9451 gnd.n2633 gnd.n2524 19.3944
R9452 gnd.n2684 gnd.n2524 19.3944
R9453 gnd.n2685 gnd.n2684 19.3944
R9454 gnd.n2686 gnd.n2685 19.3944
R9455 gnd.n2686 gnd.n2519 19.3944
R9456 gnd.n2699 gnd.n2519 19.3944
R9457 gnd.n2700 gnd.n2699 19.3944
R9458 gnd.n2702 gnd.n2700 19.3944
R9459 gnd.n2702 gnd.n2701 19.3944
R9460 gnd.n2701 gnd.n2510 19.3944
R9461 gnd.n2718 gnd.n2510 19.3944
R9462 gnd.n2718 gnd.n2717 19.3944
R9463 gnd.n2717 gnd.n2514 19.3944
R9464 gnd.n2514 gnd.n2513 19.3944
R9465 gnd.n2513 gnd.n2512 19.3944
R9466 gnd.n2512 gnd.n2511 19.3944
R9467 gnd.n2511 gnd.n2470 19.3944
R9468 gnd.n2771 gnd.n2470 19.3944
R9469 gnd.n2772 gnd.n2771 19.3944
R9470 gnd.n2775 gnd.n2772 19.3944
R9471 gnd.n2776 gnd.n2775 19.3944
R9472 gnd.n2781 gnd.n2776 19.3944
R9473 gnd.n2782 gnd.n2781 19.3944
R9474 gnd.n2786 gnd.n2782 19.3944
R9475 gnd.n2786 gnd.n2785 19.3944
R9476 gnd.n2785 gnd.n2784 19.3944
R9477 gnd.n2784 gnd.n2444 19.3944
R9478 gnd.n2851 gnd.n2444 19.3944
R9479 gnd.n2852 gnd.n2851 19.3944
R9480 gnd.n2854 gnd.n2852 19.3944
R9481 gnd.n2854 gnd.n2439 19.3944
R9482 gnd.n2866 gnd.n2439 19.3944
R9483 gnd.n2867 gnd.n2866 19.3944
R9484 gnd.n2869 gnd.n2867 19.3944
R9485 gnd.n2870 gnd.n2869 19.3944
R9486 gnd.n2873 gnd.n2870 19.3944
R9487 gnd.n2874 gnd.n2873 19.3944
R9488 gnd.n2878 gnd.n2874 19.3944
R9489 gnd.n2879 gnd.n2878 19.3944
R9490 gnd.n2881 gnd.n2879 19.3944
R9491 gnd.n2881 gnd.n2880 19.3944
R9492 gnd.n1158 gnd.n1137 19.3944
R9493 gnd.n1159 gnd.n1158 19.3944
R9494 gnd.n5032 gnd.n1159 19.3944
R9495 gnd.n5032 gnd.n5031 19.3944
R9496 gnd.n5031 gnd.n5030 19.3944
R9497 gnd.n5030 gnd.n1163 19.3944
R9498 gnd.n5020 gnd.n1163 19.3944
R9499 gnd.n5020 gnd.n5019 19.3944
R9500 gnd.n5019 gnd.n5018 19.3944
R9501 gnd.n5018 gnd.n1182 19.3944
R9502 gnd.n5008 gnd.n1182 19.3944
R9503 gnd.n5008 gnd.n5007 19.3944
R9504 gnd.n5007 gnd.n5006 19.3944
R9505 gnd.n5006 gnd.n1202 19.3944
R9506 gnd.n4996 gnd.n1202 19.3944
R9507 gnd.n4996 gnd.n4995 19.3944
R9508 gnd.n4995 gnd.n4994 19.3944
R9509 gnd.n4994 gnd.n1222 19.3944
R9510 gnd.n4984 gnd.n1222 19.3944
R9511 gnd.n4984 gnd.n4983 19.3944
R9512 gnd.n4983 gnd.n4982 19.3944
R9513 gnd.n4982 gnd.n1243 19.3944
R9514 gnd.n2720 gnd.n1243 19.3944
R9515 gnd.n2720 gnd.n2492 19.3944
R9516 gnd.n2745 gnd.n2492 19.3944
R9517 gnd.n2745 gnd.n2744 19.3944
R9518 gnd.n2744 gnd.n2743 19.3944
R9519 gnd.n2743 gnd.n2472 19.3944
R9520 gnd.n2768 gnd.n2472 19.3944
R9521 gnd.n2768 gnd.n1268 19.3944
R9522 gnd.n4970 gnd.n1268 19.3944
R9523 gnd.n4970 gnd.n4969 19.3944
R9524 gnd.n4969 gnd.n4968 19.3944
R9525 gnd.n4968 gnd.n1272 19.3944
R9526 gnd.n4958 gnd.n1272 19.3944
R9527 gnd.n4958 gnd.n4957 19.3944
R9528 gnd.n4957 gnd.n4956 19.3944
R9529 gnd.n4956 gnd.n1291 19.3944
R9530 gnd.n4946 gnd.n1291 19.3944
R9531 gnd.n4946 gnd.n4945 19.3944
R9532 gnd.n4945 gnd.n4944 19.3944
R9533 gnd.n4944 gnd.n1311 19.3944
R9534 gnd.n4934 gnd.n1311 19.3944
R9535 gnd.n4934 gnd.n4933 19.3944
R9536 gnd.n4933 gnd.n4932 19.3944
R9537 gnd.n4932 gnd.n1331 19.3944
R9538 gnd.n4922 gnd.n1331 19.3944
R9539 gnd.n4922 gnd.n4921 19.3944
R9540 gnd.n4921 gnd.n4920 19.3944
R9541 gnd.n4920 gnd.n1351 19.3944
R9542 gnd.n4910 gnd.n1351 19.3944
R9543 gnd.n4910 gnd.n4909 19.3944
R9544 gnd.n4909 gnd.n4908 19.3944
R9545 gnd.n4901 gnd.n4900 19.3944
R9546 gnd.n4900 gnd.n1380 19.3944
R9547 gnd.n1382 gnd.n1380 19.3944
R9548 gnd.n4893 gnd.n1382 19.3944
R9549 gnd.n4893 gnd.n4892 19.3944
R9550 gnd.n4892 gnd.n4891 19.3944
R9551 gnd.n4891 gnd.n1389 19.3944
R9552 gnd.n4886 gnd.n1389 19.3944
R9553 gnd.n4886 gnd.n4885 19.3944
R9554 gnd.n4885 gnd.n4884 19.3944
R9555 gnd.n4884 gnd.n1396 19.3944
R9556 gnd.n4879 gnd.n1396 19.3944
R9557 gnd.n4879 gnd.n4878 19.3944
R9558 gnd.n4878 gnd.n4877 19.3944
R9559 gnd.n4877 gnd.n1403 19.3944
R9560 gnd.n4872 gnd.n1403 19.3944
R9561 gnd.n4872 gnd.n4871 19.3944
R9562 gnd.n3009 gnd.n2969 19.3944
R9563 gnd.n3013 gnd.n2969 19.3944
R9564 gnd.n3013 gnd.n2967 19.3944
R9565 gnd.n3019 gnd.n2967 19.3944
R9566 gnd.n3019 gnd.n2965 19.3944
R9567 gnd.n3023 gnd.n2965 19.3944
R9568 gnd.n3023 gnd.n2963 19.3944
R9569 gnd.n3029 gnd.n2963 19.3944
R9570 gnd.n3029 gnd.n2961 19.3944
R9571 gnd.n3033 gnd.n2961 19.3944
R9572 gnd.n3033 gnd.n2959 19.3944
R9573 gnd.n3039 gnd.n2959 19.3944
R9574 gnd.n3039 gnd.n2957 19.3944
R9575 gnd.n3043 gnd.n2957 19.3944
R9576 gnd.n3043 gnd.n2955 19.3944
R9577 gnd.n3049 gnd.n2955 19.3944
R9578 gnd.n3049 gnd.n2953 19.3944
R9579 gnd.n3053 gnd.n2953 19.3944
R9580 gnd.n2982 gnd.n1425 19.3944
R9581 gnd.n2989 gnd.n2982 19.3944
R9582 gnd.n2989 gnd.n2979 19.3944
R9583 gnd.n2993 gnd.n2979 19.3944
R9584 gnd.n2993 gnd.n2977 19.3944
R9585 gnd.n2999 gnd.n2977 19.3944
R9586 gnd.n2999 gnd.n2975 19.3944
R9587 gnd.n3003 gnd.n2975 19.3944
R9588 gnd.n4869 gnd.n1412 19.3944
R9589 gnd.n4864 gnd.n1412 19.3944
R9590 gnd.n4864 gnd.n4863 19.3944
R9591 gnd.n4863 gnd.n4862 19.3944
R9592 gnd.n4862 gnd.n1419 19.3944
R9593 gnd.n4857 gnd.n1419 19.3944
R9594 gnd.n4857 gnd.n4856 19.3944
R9595 gnd.n5038 gnd.n1145 19.3944
R9596 gnd.n5038 gnd.n5037 19.3944
R9597 gnd.n5037 gnd.n5036 19.3944
R9598 gnd.n5036 gnd.n1150 19.3944
R9599 gnd.n5026 gnd.n1150 19.3944
R9600 gnd.n5026 gnd.n5025 19.3944
R9601 gnd.n5025 gnd.n5024 19.3944
R9602 gnd.n5024 gnd.n1173 19.3944
R9603 gnd.n5014 gnd.n1173 19.3944
R9604 gnd.n5014 gnd.n5013 19.3944
R9605 gnd.n5013 gnd.n5012 19.3944
R9606 gnd.n5012 gnd.n1192 19.3944
R9607 gnd.n5002 gnd.n1192 19.3944
R9608 gnd.n5002 gnd.n5001 19.3944
R9609 gnd.n5001 gnd.n5000 19.3944
R9610 gnd.n5000 gnd.n1213 19.3944
R9611 gnd.n4990 gnd.n1213 19.3944
R9612 gnd.n4990 gnd.n4989 19.3944
R9613 gnd.n4989 gnd.n4988 19.3944
R9614 gnd.n4988 gnd.n1233 19.3944
R9615 gnd.n4978 gnd.n1233 19.3944
R9616 gnd.n4978 gnd.n4977 19.3944
R9617 gnd.n1258 gnd.n1252 19.3944
R9618 gnd.n2487 gnd.n1258 19.3944
R9619 gnd.n2750 gnd.n2749 19.3944
R9620 gnd.n2764 gnd.n2763 19.3944
R9621 gnd.n4974 gnd.n1259 19.3944
R9622 gnd.n4974 gnd.n1260 19.3944
R9623 gnd.n4964 gnd.n1260 19.3944
R9624 gnd.n4964 gnd.n4963 19.3944
R9625 gnd.n4963 gnd.n4962 19.3944
R9626 gnd.n4962 gnd.n1281 19.3944
R9627 gnd.n4952 gnd.n1281 19.3944
R9628 gnd.n4952 gnd.n4951 19.3944
R9629 gnd.n4951 gnd.n4950 19.3944
R9630 gnd.n4950 gnd.n1302 19.3944
R9631 gnd.n4940 gnd.n1302 19.3944
R9632 gnd.n4940 gnd.n4939 19.3944
R9633 gnd.n4939 gnd.n4938 19.3944
R9634 gnd.n4938 gnd.n1321 19.3944
R9635 gnd.n4928 gnd.n1321 19.3944
R9636 gnd.n4928 gnd.n4927 19.3944
R9637 gnd.n4927 gnd.n4926 19.3944
R9638 gnd.n4926 gnd.n1342 19.3944
R9639 gnd.n4916 gnd.n1342 19.3944
R9640 gnd.n4916 gnd.n4915 19.3944
R9641 gnd.n4915 gnd.n4914 19.3944
R9642 gnd.n4914 gnd.n1362 19.3944
R9643 gnd.n4904 gnd.n1362 19.3944
R9644 gnd.n6747 gnd.n6746 19.3944
R9645 gnd.n6746 gnd.n6745 19.3944
R9646 gnd.n6745 gnd.n806 19.3944
R9647 gnd.n6739 gnd.n806 19.3944
R9648 gnd.n6739 gnd.n6738 19.3944
R9649 gnd.n6738 gnd.n6737 19.3944
R9650 gnd.n6737 gnd.n814 19.3944
R9651 gnd.n6731 gnd.n814 19.3944
R9652 gnd.n6731 gnd.n6730 19.3944
R9653 gnd.n6730 gnd.n6729 19.3944
R9654 gnd.n6729 gnd.n822 19.3944
R9655 gnd.n6723 gnd.n822 19.3944
R9656 gnd.n6723 gnd.n6722 19.3944
R9657 gnd.n6722 gnd.n6721 19.3944
R9658 gnd.n6721 gnd.n830 19.3944
R9659 gnd.n6715 gnd.n830 19.3944
R9660 gnd.n6715 gnd.n6714 19.3944
R9661 gnd.n6714 gnd.n6713 19.3944
R9662 gnd.n6713 gnd.n838 19.3944
R9663 gnd.n6707 gnd.n838 19.3944
R9664 gnd.n6707 gnd.n6706 19.3944
R9665 gnd.n6706 gnd.n6705 19.3944
R9666 gnd.n6705 gnd.n846 19.3944
R9667 gnd.n6699 gnd.n846 19.3944
R9668 gnd.n6699 gnd.n6698 19.3944
R9669 gnd.n6698 gnd.n6697 19.3944
R9670 gnd.n6697 gnd.n854 19.3944
R9671 gnd.n6691 gnd.n854 19.3944
R9672 gnd.n6691 gnd.n6690 19.3944
R9673 gnd.n6690 gnd.n6689 19.3944
R9674 gnd.n6689 gnd.n862 19.3944
R9675 gnd.n6683 gnd.n862 19.3944
R9676 gnd.n6683 gnd.n6682 19.3944
R9677 gnd.n6682 gnd.n6681 19.3944
R9678 gnd.n6681 gnd.n870 19.3944
R9679 gnd.n6675 gnd.n870 19.3944
R9680 gnd.n6675 gnd.n6674 19.3944
R9681 gnd.n6674 gnd.n6673 19.3944
R9682 gnd.n6673 gnd.n878 19.3944
R9683 gnd.n6667 gnd.n878 19.3944
R9684 gnd.n6667 gnd.n6666 19.3944
R9685 gnd.n6666 gnd.n6665 19.3944
R9686 gnd.n6665 gnd.n886 19.3944
R9687 gnd.n6659 gnd.n886 19.3944
R9688 gnd.n6659 gnd.n6658 19.3944
R9689 gnd.n6658 gnd.n6657 19.3944
R9690 gnd.n6657 gnd.n894 19.3944
R9691 gnd.n6651 gnd.n894 19.3944
R9692 gnd.n6651 gnd.n6650 19.3944
R9693 gnd.n6650 gnd.n6649 19.3944
R9694 gnd.n6649 gnd.n902 19.3944
R9695 gnd.n6643 gnd.n902 19.3944
R9696 gnd.n6643 gnd.n6642 19.3944
R9697 gnd.n6642 gnd.n6641 19.3944
R9698 gnd.n6641 gnd.n910 19.3944
R9699 gnd.n6635 gnd.n910 19.3944
R9700 gnd.n6635 gnd.n6634 19.3944
R9701 gnd.n6634 gnd.n6633 19.3944
R9702 gnd.n6633 gnd.n918 19.3944
R9703 gnd.n6627 gnd.n918 19.3944
R9704 gnd.n6627 gnd.n6626 19.3944
R9705 gnd.n6626 gnd.n6625 19.3944
R9706 gnd.n6625 gnd.n926 19.3944
R9707 gnd.n6619 gnd.n926 19.3944
R9708 gnd.n6619 gnd.n6618 19.3944
R9709 gnd.n6618 gnd.n6617 19.3944
R9710 gnd.n6617 gnd.n934 19.3944
R9711 gnd.n6611 gnd.n934 19.3944
R9712 gnd.n6611 gnd.n6610 19.3944
R9713 gnd.n6610 gnd.n6609 19.3944
R9714 gnd.n6609 gnd.n942 19.3944
R9715 gnd.n6603 gnd.n942 19.3944
R9716 gnd.n6603 gnd.n6602 19.3944
R9717 gnd.n6602 gnd.n6601 19.3944
R9718 gnd.n6601 gnd.n950 19.3944
R9719 gnd.n6595 gnd.n950 19.3944
R9720 gnd.n6595 gnd.n6594 19.3944
R9721 gnd.n6594 gnd.n6593 19.3944
R9722 gnd.n6593 gnd.n958 19.3944
R9723 gnd.n6587 gnd.n958 19.3944
R9724 gnd.n6587 gnd.n6586 19.3944
R9725 gnd.n6586 gnd.n6585 19.3944
R9726 gnd.n6585 gnd.n966 19.3944
R9727 gnd.n2650 gnd.n966 19.3944
R9728 gnd.n3215 gnd.n2386 19.3944
R9729 gnd.n3215 gnd.n2383 19.3944
R9730 gnd.n3220 gnd.n2383 19.3944
R9731 gnd.n3220 gnd.n2384 19.3944
R9732 gnd.n2384 gnd.n2362 19.3944
R9733 gnd.n3248 gnd.n2362 19.3944
R9734 gnd.n3248 gnd.n2359 19.3944
R9735 gnd.n3256 gnd.n2359 19.3944
R9736 gnd.n3256 gnd.n2360 19.3944
R9737 gnd.n3252 gnd.n2360 19.3944
R9738 gnd.n3252 gnd.n1507 19.3944
R9739 gnd.n4771 gnd.n1507 19.3944
R9740 gnd.n4771 gnd.n1508 19.3944
R9741 gnd.n4767 gnd.n1508 19.3944
R9742 gnd.n4767 gnd.n4766 19.3944
R9743 gnd.n4766 gnd.n4765 19.3944
R9744 gnd.n4765 gnd.n1514 19.3944
R9745 gnd.n4761 gnd.n1514 19.3944
R9746 gnd.n4761 gnd.n4760 19.3944
R9747 gnd.n4760 gnd.n4759 19.3944
R9748 gnd.n4759 gnd.n1519 19.3944
R9749 gnd.n4755 gnd.n1519 19.3944
R9750 gnd.n4755 gnd.n4754 19.3944
R9751 gnd.n4754 gnd.n4753 19.3944
R9752 gnd.n4753 gnd.n1524 19.3944
R9753 gnd.n4749 gnd.n1524 19.3944
R9754 gnd.n4749 gnd.n4748 19.3944
R9755 gnd.n4748 gnd.n4747 19.3944
R9756 gnd.n4747 gnd.n1529 19.3944
R9757 gnd.n4743 gnd.n1529 19.3944
R9758 gnd.n4743 gnd.n4742 19.3944
R9759 gnd.n4742 gnd.n4741 19.3944
R9760 gnd.n4741 gnd.n1534 19.3944
R9761 gnd.n4737 gnd.n1534 19.3944
R9762 gnd.n4737 gnd.n4736 19.3944
R9763 gnd.n4736 gnd.n4735 19.3944
R9764 gnd.n4735 gnd.n1539 19.3944
R9765 gnd.n4731 gnd.n1539 19.3944
R9766 gnd.n4731 gnd.n4730 19.3944
R9767 gnd.n4730 gnd.n4729 19.3944
R9768 gnd.n4729 gnd.n1544 19.3944
R9769 gnd.n4725 gnd.n1544 19.3944
R9770 gnd.n4725 gnd.n4724 19.3944
R9771 gnd.n4724 gnd.n4723 19.3944
R9772 gnd.n4723 gnd.n1549 19.3944
R9773 gnd.n4719 gnd.n1549 19.3944
R9774 gnd.n4719 gnd.n4718 19.3944
R9775 gnd.n4718 gnd.n4717 19.3944
R9776 gnd.n4717 gnd.n1554 19.3944
R9777 gnd.n4713 gnd.n1554 19.3944
R9778 gnd.n4713 gnd.n4712 19.3944
R9779 gnd.n4712 gnd.n4711 19.3944
R9780 gnd.n4711 gnd.n1559 19.3944
R9781 gnd.n4707 gnd.n1559 19.3944
R9782 gnd.n4707 gnd.n4706 19.3944
R9783 gnd.n4706 gnd.n4705 19.3944
R9784 gnd.n4705 gnd.n1564 19.3944
R9785 gnd.n4701 gnd.n1564 19.3944
R9786 gnd.n4701 gnd.n4700 19.3944
R9787 gnd.n4700 gnd.n4699 19.3944
R9788 gnd.n4699 gnd.n1569 19.3944
R9789 gnd.n4695 gnd.n1569 19.3944
R9790 gnd.n4695 gnd.n4694 19.3944
R9791 gnd.n4694 gnd.n4693 19.3944
R9792 gnd.n4693 gnd.n1574 19.3944
R9793 gnd.n4689 gnd.n1574 19.3944
R9794 gnd.n4689 gnd.n4688 19.3944
R9795 gnd.n4688 gnd.n4687 19.3944
R9796 gnd.n4687 gnd.n1579 19.3944
R9797 gnd.n4683 gnd.n1579 19.3944
R9798 gnd.n4683 gnd.n4682 19.3944
R9799 gnd.n4682 gnd.n4681 19.3944
R9800 gnd.n4681 gnd.n1584 19.3944
R9801 gnd.n4677 gnd.n1584 19.3944
R9802 gnd.n4677 gnd.n4676 19.3944
R9803 gnd.n4676 gnd.n4675 19.3944
R9804 gnd.n4675 gnd.n1589 19.3944
R9805 gnd.n4671 gnd.n1589 19.3944
R9806 gnd.n4671 gnd.n4670 19.3944
R9807 gnd.n4670 gnd.n4669 19.3944
R9808 gnd.n4669 gnd.n1594 19.3944
R9809 gnd.n4665 gnd.n1594 19.3944
R9810 gnd.n3950 gnd.n3948 19.3944
R9811 gnd.n3950 gnd.n3946 19.3944
R9812 gnd.n3956 gnd.n3946 19.3944
R9813 gnd.n3956 gnd.n3944 19.3944
R9814 gnd.n3961 gnd.n3944 19.3944
R9815 gnd.n3961 gnd.n3942 19.3944
R9816 gnd.n3967 gnd.n3942 19.3944
R9817 gnd.n3967 gnd.n3941 19.3944
R9818 gnd.n3976 gnd.n3941 19.3944
R9819 gnd.n3976 gnd.n3939 19.3944
R9820 gnd.n3982 gnd.n3939 19.3944
R9821 gnd.n3982 gnd.n3932 19.3944
R9822 gnd.n3995 gnd.n3932 19.3944
R9823 gnd.n3995 gnd.n3930 19.3944
R9824 gnd.n4001 gnd.n3930 19.3944
R9825 gnd.n4001 gnd.n3923 19.3944
R9826 gnd.n4014 gnd.n3923 19.3944
R9827 gnd.n4014 gnd.n3921 19.3944
R9828 gnd.n4020 gnd.n3921 19.3944
R9829 gnd.n4020 gnd.n3914 19.3944
R9830 gnd.n4033 gnd.n3914 19.3944
R9831 gnd.n4033 gnd.n3912 19.3944
R9832 gnd.n4040 gnd.n3912 19.3944
R9833 gnd.n4040 gnd.n4039 19.3944
R9834 gnd.n4053 gnd.n3893 19.3944
R9835 gnd.n3893 gnd.n3892 19.3944
R9836 gnd.n4060 gnd.n3892 19.3944
R9837 gnd.n4785 gnd.n4784 19.2005
R9838 gnd.n4177 gnd.n4176 19.2005
R9839 gnd.n5952 gnd.t190 18.8012
R9840 gnd.n5991 gnd.t4 18.8012
R9841 gnd.n5795 gnd.n5537 18.4825
R9842 gnd.n6581 gnd.n968 18.4825
R9843 gnd.n4342 gnd.n4250 18.4247
R9844 gnd.n4856 gnd.n4855 18.4247
R9845 gnd.n4050 gnd.n4049 18.2308
R9846 gnd.n3186 gnd.n2406 18.2308
R9847 gnd.n7532 gnd.n7531 18.2308
R9848 gnd.n2603 gnd.n2602 18.2308
R9849 gnd.t74 gnd.n5479 18.1639
R9850 gnd.n1184 gnd.n1177 18.1639
R9851 gnd.n7699 gnd.n172 18.1639
R9852 gnd.n5508 gnd.t192 17.5266
R9853 gnd.t56 gnd.n1167 17.5266
R9854 gnd.n4924 gnd.t14 17.5266
R9855 gnd.n4629 gnd.t36 17.5266
R9856 gnd.n7693 gnd.t140 17.5266
R9857 gnd.t325 gnd.n5455 16.8893
R9858 gnd.n4948 gnd.t138 16.8893
R9859 gnd.n4605 gnd.t0 16.8893
R9860 gnd.n4372 gnd.n1852 16.6793
R9861 gnd.n7604 gnd.n7603 16.6793
R9862 gnd.n5091 gnd.n5088 16.6793
R9863 gnd.n3003 gnd.n2973 16.6793
R9864 gnd.t209 gnd.n5564 16.2519
R9865 gnd.n5422 gnd.t326 16.2519
R9866 gnd.n4972 gnd.t20 16.2519
R9867 gnd.n4581 gnd.t120 16.2519
R9868 gnd.n3180 gnd.n2926 15.9333
R9869 gnd.n3180 gnd.n2397 15.9333
R9870 gnd.n3202 gnd.n3201 15.9333
R9871 gnd.n3201 gnd.n2388 15.9333
R9872 gnd.n3213 gnd.n2388 15.9333
R9873 gnd.n3213 gnd.n3212 15.9333
R9874 gnd.n2390 gnd.n2379 15.9333
R9875 gnd.n3222 gnd.n2379 15.9333
R9876 gnd.n3222 gnd.n2380 15.9333
R9877 gnd.n2380 gnd.n2372 15.9333
R9878 gnd.n3234 gnd.n2372 15.9333
R9879 gnd.n3234 gnd.n3233 15.9333
R9880 gnd.n3233 gnd.n2364 15.9333
R9881 gnd.n3246 gnd.n2364 15.9333
R9882 gnd.n3245 gnd.n1433 15.9333
R9883 gnd.n3258 gnd.n1465 15.9333
R9884 gnd.n4780 gnd.n1493 15.9333
R9885 gnd.n3281 gnd.n2251 15.9333
R9886 gnd.n3324 gnd.n2240 15.9333
R9887 gnd.n3358 gnd.n2228 15.9333
R9888 gnd.n3370 gnd.n3368 15.9333
R9889 gnd.n3397 gnd.n2208 15.9333
R9890 gnd.n3488 gnd.n2158 15.9333
R9891 gnd.n3507 gnd.n2135 15.9333
R9892 gnd.n2142 gnd.n2130 15.9333
R9893 gnd.n3547 gnd.n2113 15.9333
R9894 gnd.n3595 gnd.n3594 15.9333
R9895 gnd.n3603 gnd.n2100 15.9333
R9896 gnd.n3620 gnd.n3619 15.9333
R9897 gnd.n3680 gnd.n2067 15.9333
R9898 gnd.n3760 gnd.n3759 15.9333
R9899 gnd.n3768 gnd.n2010 15.9333
R9900 gnd.n3786 gnd.n3785 15.9333
R9901 gnd.n3796 gnd.n1982 15.9333
R9902 gnd.n3818 gnd.n1976 15.9333
R9903 gnd.n4088 gnd.n4087 15.9333
R9904 gnd.n3871 gnd.n1902 15.9333
R9905 gnd.n3871 gnd.n1865 15.9333
R9906 gnd.n4080 gnd.n1919 15.9333
R9907 gnd.n4079 gnd.n4078 15.9333
R9908 gnd.n4078 gnd.n4077 15.9333
R9909 gnd.n4077 gnd.n4075 15.9333
R9910 gnd.n4075 gnd.n1922 15.9333
R9911 gnd.n1934 gnd.n1922 15.9333
R9912 gnd.n1935 gnd.n1934 15.9333
R9913 gnd.n4069 gnd.n1935 15.9333
R9914 gnd.n4069 gnd.n4068 15.9333
R9915 gnd.n4067 gnd.n4066 15.9333
R9916 gnd.n4066 gnd.n1598 15.9333
R9917 gnd.n4663 gnd.n1598 15.9333
R9918 gnd.n4663 gnd.n4662 15.9333
R9919 gnd.n1609 gnd.n1600 15.9333
R9920 gnd.n4656 gnd.n1609 15.9333
R9921 gnd.n6391 gnd.n6389 15.6674
R9922 gnd.n6359 gnd.n6357 15.6674
R9923 gnd.n6327 gnd.n6325 15.6674
R9924 gnd.n6296 gnd.n6294 15.6674
R9925 gnd.n6264 gnd.n6262 15.6674
R9926 gnd.n6232 gnd.n6230 15.6674
R9927 gnd.n6200 gnd.n6198 15.6674
R9928 gnd.n6169 gnd.n6167 15.6674
R9929 gnd.n5682 gnd.t209 15.6146
R9930 gnd.t205 gnd.n6552 15.6146
R9931 gnd.n6456 gnd.t306 15.6146
R9932 gnd.t25 gnd.n2723 15.6146
R9933 gnd.t261 gnd.n2390 15.6146
R9934 gnd.n4068 gnd.t245 15.6146
R9935 gnd.n7446 gnd.t54 15.6146
R9936 gnd.n4424 gnd.n1831 15.3217
R9937 gnd.n7564 gnd.n315 15.3217
R9938 gnd.n5048 gnd.n1133 15.3217
R9939 gnd.n3058 gnd.n2951 15.3217
R9940 gnd.n3398 gnd.n2213 15.296
R9941 gnd.n3417 gnd.n2204 15.296
R9942 gnd.n3378 gnd.t200 15.296
R9943 gnd.n3548 gnd.n3546 15.296
R9944 gnd.n3593 gnd.n2109 15.296
R9945 gnd.n3720 gnd.t183 15.296
R9946 gnd.n3660 gnd.n2032 15.296
R9947 gnd.n3758 gnd.n2019 15.296
R9948 gnd.n1960 gnd.t224 15.296
R9949 gnd.n4097 gnd.n4096 15.0827
R9950 gnd.n1477 gnd.n1472 15.0481
R9951 gnd.n4107 gnd.n4106 15.0481
R9952 gnd.n6120 gnd.t72 14.9773
R9953 gnd.n4998 gnd.t78 14.9773
R9954 gnd.n4851 gnd.n1433 14.9773
R9955 gnd.n7474 gnd.t75 14.9773
R9956 gnd.n3258 gnd.t300 14.6587
R9957 gnd.n3325 gnd.n2235 14.6587
R9958 gnd.n3460 gnd.n3459 14.6587
R9959 gnd.n2060 gnd.n2049 14.6587
R9960 gnd.n3798 gnd.n3797 14.6587
R9961 gnd.t221 gnd.n1956 14.6587
R9962 gnd.n3845 gnd.n3844 14.6587
R9963 gnd.n6573 gnd.t178 14.34
R9964 gnd.t188 gnd.n993 14.34
R9965 gnd.n5022 gnd.t56 14.34
R9966 gnd.t140 gnd.n175 14.34
R9967 gnd.n3283 gnd.t252 14.0214
R9968 gnd.n3333 gnd.n2220 14.0214
R9969 gnd.n3377 gnd.n2189 14.0214
R9970 gnd.n3538 gnd.n3537 14.0214
R9971 gnd.n2099 gnd.n2091 14.0214
R9972 gnd.n3721 gnd.n2036 14.0214
R9973 gnd.n2008 gnd.n2007 14.0214
R9974 gnd.n4089 gnd.n1907 14.0214
R9975 gnd.t42 gnd.n5879 13.7027
R9976 gnd.n5016 gnd.n1184 13.7027
R9977 gnd.n2162 gnd.t85 13.7027
R9978 gnd.n3628 gnd.t16 13.7027
R9979 gnd.n7510 gnd.n172 13.7027
R9980 gnd.n5764 gnd.n5760 13.5763
R9981 gnd.n6512 gnd.n5197 13.5763
R9982 gnd.n5796 gnd.n5795 13.384
R9983 gnd.n3268 gnd.n1502 13.384
R9984 gnd.n3357 gnd.n2230 13.384
R9985 gnd.n2190 gnd.n2184 13.384
R9986 gnd.t49 gnd.n3447 13.384
R9987 gnd.n3699 gnd.t117 13.384
R9988 gnd.n3708 gnd.n2045 13.384
R9989 gnd.n3736 gnd.n1996 13.384
R9990 gnd.n3861 gnd.n1947 13.384
R9991 gnd.n1488 gnd.n1469 13.1884
R9992 gnd.n1483 gnd.n1482 13.1884
R9993 gnd.n1482 gnd.n1481 13.1884
R9994 gnd.n4100 gnd.n4095 13.1884
R9995 gnd.n4101 gnd.n4100 13.1884
R9996 gnd.n1484 gnd.n1471 13.146
R9997 gnd.n1480 gnd.n1471 13.146
R9998 gnd.n4099 gnd.n4098 13.146
R9999 gnd.n4099 gnd.n4094 13.146
R10000 gnd.n3299 gnd.t68 13.0654
R10001 gnd.n3819 gnd.t66 13.0654
R10002 gnd.n6392 gnd.n6388 12.8005
R10003 gnd.n6360 gnd.n6356 12.8005
R10004 gnd.n6328 gnd.n6324 12.8005
R10005 gnd.n6297 gnd.n6293 12.8005
R10006 gnd.n6265 gnd.n6261 12.8005
R10007 gnd.n6233 gnd.n6229 12.8005
R10008 gnd.n6201 gnd.n6197 12.8005
R10009 gnd.n6170 gnd.n6166 12.8005
R10010 gnd.n2266 gnd.n1504 12.7467
R10011 gnd.n3316 gnd.t279 12.7467
R10012 gnd.n3341 gnd.n3340 12.7467
R10013 gnd.n3508 gnd.n3506 12.7467
R10014 gnd.n3618 gnd.n2078 12.7467
R10015 gnd.n3784 gnd.n3783 12.7467
R10016 gnd.n5767 gnd.n5764 12.4126
R10017 gnd.n6517 gnd.n5197 12.4126
R10018 gnd.n4848 gnd.n4785 12.1761
R10019 gnd.n4176 gnd.n4175 12.1761
R10020 gnd.n4781 gnd.n1491 12.1094
R10021 gnd.t232 gnd.n2270 12.1094
R10022 gnd.n3348 gnd.n2221 12.1094
R10023 gnd.n3429 gnd.n2195 12.1094
R10024 gnd.n3728 gnd.n2030 12.1094
R10025 gnd.n3769 gnd.n2005 12.1094
R10026 gnd.n3869 gnd.n1910 12.1094
R10027 gnd.n6396 gnd.n6395 12.0247
R10028 gnd.n6364 gnd.n6363 12.0247
R10029 gnd.n6332 gnd.n6331 12.0247
R10030 gnd.n6301 gnd.n6300 12.0247
R10031 gnd.n6269 gnd.n6268 12.0247
R10032 gnd.n6237 gnd.n6236 12.0247
R10033 gnd.n6205 gnd.n6204 12.0247
R10034 gnd.n6174 gnd.n6173 12.0247
R10035 gnd.n2681 gnd.t78 11.7908
R10036 gnd.t75 gnd.n143 11.7908
R10037 gnd.n2918 gnd.n1381 11.4721
R10038 gnd.n3309 gnd.n2252 11.4721
R10039 gnd.n3301 gnd.n3300 11.4721
R10040 gnd.n3468 gnd.t186 11.4721
R10041 gnd.n3467 gnd.n2171 11.4721
R10042 gnd.n3498 gnd.n3497 11.4721
R10043 gnd.n3645 gnd.n2073 11.4721
R10044 gnd.n3637 gnd.n2059 11.4721
R10045 gnd.n3689 gnd.t83 11.4721
R10046 gnd.n3809 gnd.n1983 11.4721
R10047 gnd.n3830 gnd.n3829 11.4721
R10048 gnd.n4654 gnd.n1610 11.4721
R10049 gnd.n6399 gnd.n6386 11.249
R10050 gnd.n6367 gnd.n6354 11.249
R10051 gnd.n6335 gnd.n6322 11.249
R10052 gnd.n6304 gnd.n6291 11.249
R10053 gnd.n6272 gnd.n6259 11.249
R10054 gnd.n6240 gnd.n6227 11.249
R10055 gnd.n6208 gnd.n6195 11.249
R10056 gnd.n6177 gnd.n6164 11.249
R10057 gnd.n5880 gnd.t42 11.1535
R10058 gnd.n2724 gnd.t25 11.1535
R10059 gnd.n3246 gnd.t351 11.1535
R10060 gnd.n3445 gnd.t102 11.1535
R10061 gnd.t172 gnd.n3700 11.1535
R10062 gnd.t146 gnd.n4079 11.1535
R10063 gnd.t54 gnd.n102 11.1535
R10064 gnd.n3411 gnd.n3410 10.8348
R10065 gnd.n3410 gnd.n3409 10.8348
R10066 gnd.n3587 gnd.n3586 10.8348
R10067 gnd.n3586 gnd.n2106 10.8348
R10068 gnd.n3752 gnd.n3751 10.8348
R10069 gnd.n3751 gnd.n2016 10.8348
R10070 gnd.n1832 gnd.n1831 10.6672
R10071 gnd.n7569 gnd.n315 10.6672
R10072 gnd.n5051 gnd.n5048 10.6672
R10073 gnd.n3053 gnd.n2951 10.6672
R10074 gnd.n4241 gnd.n1861 10.6151
R10075 gnd.n4241 gnd.n4240 10.6151
R10076 gnd.n4238 gnd.n4235 10.6151
R10077 gnd.n4235 gnd.n4234 10.6151
R10078 gnd.n4234 gnd.n4231 10.6151
R10079 gnd.n4231 gnd.n4230 10.6151
R10080 gnd.n4230 gnd.n4227 10.6151
R10081 gnd.n4227 gnd.n4226 10.6151
R10082 gnd.n4226 gnd.n4223 10.6151
R10083 gnd.n4223 gnd.n4222 10.6151
R10084 gnd.n4222 gnd.n4219 10.6151
R10085 gnd.n4219 gnd.n4218 10.6151
R10086 gnd.n4218 gnd.n4215 10.6151
R10087 gnd.n4215 gnd.n4214 10.6151
R10088 gnd.n4214 gnd.n4211 10.6151
R10089 gnd.n4211 gnd.n4210 10.6151
R10090 gnd.n4210 gnd.n4207 10.6151
R10091 gnd.n4207 gnd.n4206 10.6151
R10092 gnd.n4206 gnd.n4203 10.6151
R10093 gnd.n4203 gnd.n4202 10.6151
R10094 gnd.n4202 gnd.n4199 10.6151
R10095 gnd.n4199 gnd.n4198 10.6151
R10096 gnd.n4198 gnd.n4195 10.6151
R10097 gnd.n4195 gnd.n4194 10.6151
R10098 gnd.n4194 gnd.n4191 10.6151
R10099 gnd.n4191 gnd.n4190 10.6151
R10100 gnd.n4190 gnd.n4187 10.6151
R10101 gnd.n4187 gnd.n4186 10.6151
R10102 gnd.n4186 gnd.n4183 10.6151
R10103 gnd.n4183 gnd.n4182 10.6151
R10104 gnd.n2353 gnd.n2352 10.6151
R10105 gnd.n2352 gnd.n2351 10.6151
R10106 gnd.n2351 gnd.n2348 10.6151
R10107 gnd.n2348 gnd.n2347 10.6151
R10108 gnd.n2347 gnd.n2344 10.6151
R10109 gnd.n2344 gnd.n2343 10.6151
R10110 gnd.n2343 gnd.n2249 10.6151
R10111 gnd.n3311 gnd.n2249 10.6151
R10112 gnd.n3312 gnd.n3311 10.6151
R10113 gnd.n3314 gnd.n3312 10.6151
R10114 gnd.n3314 gnd.n3313 10.6151
R10115 gnd.n3313 gnd.n2237 10.6151
R10116 gnd.n3327 gnd.n2237 10.6151
R10117 gnd.n3328 gnd.n3327 10.6151
R10118 gnd.n3338 gnd.n3328 10.6151
R10119 gnd.n3338 gnd.n3337 10.6151
R10120 gnd.n3337 gnd.n3336 10.6151
R10121 gnd.n3336 gnd.n3329 10.6151
R10122 gnd.n3330 gnd.n3329 10.6151
R10123 gnd.n3330 gnd.n2211 10.6151
R10124 gnd.n3400 gnd.n2211 10.6151
R10125 gnd.n3401 gnd.n3400 10.6151
R10126 gnd.n3407 gnd.n3401 10.6151
R10127 gnd.n3407 gnd.n3406 10.6151
R10128 gnd.n3406 gnd.n3405 10.6151
R10129 gnd.n3405 gnd.n3402 10.6151
R10130 gnd.n3402 gnd.n2187 10.6151
R10131 gnd.n3438 gnd.n2187 10.6151
R10132 gnd.n3439 gnd.n3438 10.6151
R10133 gnd.n3443 gnd.n3439 10.6151
R10134 gnd.n3443 gnd.n3442 10.6151
R10135 gnd.n3442 gnd.n3441 10.6151
R10136 gnd.n3441 gnd.n3440 10.6151
R10137 gnd.n3440 gnd.n2161 10.6151
R10138 gnd.n3486 gnd.n2161 10.6151
R10139 gnd.n3486 gnd.n3485 10.6151
R10140 gnd.n3485 gnd.n3484 10.6151
R10141 gnd.n3484 gnd.n3483 10.6151
R10142 gnd.n3483 gnd.n2143 10.6151
R10143 gnd.n3510 gnd.n2143 10.6151
R10144 gnd.n3511 gnd.n3510 10.6151
R10145 gnd.n3513 gnd.n3511 10.6151
R10146 gnd.n3514 gnd.n3513 10.6151
R10147 gnd.n3515 gnd.n3514 10.6151
R10148 gnd.n3515 gnd.n2120 10.6151
R10149 gnd.n3550 gnd.n2120 10.6151
R10150 gnd.n3551 gnd.n3550 10.6151
R10151 gnd.n3553 gnd.n3551 10.6151
R10152 gnd.n3554 gnd.n3553 10.6151
R10153 gnd.n3556 gnd.n3554 10.6151
R10154 gnd.n3556 gnd.n3555 10.6151
R10155 gnd.n3555 gnd.n2089 10.6151
R10156 gnd.n3613 gnd.n2089 10.6151
R10157 gnd.n3614 gnd.n3613 10.6151
R10158 gnd.n3616 gnd.n3614 10.6151
R10159 gnd.n3616 gnd.n3615 10.6151
R10160 gnd.n3615 gnd.n2070 10.6151
R10161 gnd.n3647 gnd.n2070 10.6151
R10162 gnd.n3648 gnd.n3647 10.6151
R10163 gnd.n3678 gnd.n3648 10.6151
R10164 gnd.n3678 gnd.n3677 10.6151
R10165 gnd.n3677 gnd.n3676 10.6151
R10166 gnd.n3676 gnd.n3673 10.6151
R10167 gnd.n3673 gnd.n3672 10.6151
R10168 gnd.n3672 gnd.n3671 10.6151
R10169 gnd.n3671 gnd.n3670 10.6151
R10170 gnd.n3670 gnd.n3669 10.6151
R10171 gnd.n3669 gnd.n3666 10.6151
R10172 gnd.n3666 gnd.n3665 10.6151
R10173 gnd.n3665 gnd.n3663 10.6151
R10174 gnd.n3663 gnd.n3662 10.6151
R10175 gnd.n3662 gnd.n3656 10.6151
R10176 gnd.n3656 gnd.n3655 10.6151
R10177 gnd.n3655 gnd.n3653 10.6151
R10178 gnd.n3653 gnd.n3652 10.6151
R10179 gnd.n3652 gnd.n3649 10.6151
R10180 gnd.n3649 gnd.n1999 10.6151
R10181 gnd.n3778 gnd.n1999 10.6151
R10182 gnd.n3779 gnd.n3778 10.6151
R10183 gnd.n3781 gnd.n3779 10.6151
R10184 gnd.n3781 gnd.n3780 10.6151
R10185 gnd.n3780 gnd.n1979 10.6151
R10186 gnd.n3811 gnd.n1979 10.6151
R10187 gnd.n3812 gnd.n3811 10.6151
R10188 gnd.n3816 gnd.n3812 10.6151
R10189 gnd.n3816 gnd.n3815 10.6151
R10190 gnd.n3815 gnd.n3814 10.6151
R10191 gnd.n3814 gnd.n3813 10.6151
R10192 gnd.n3813 gnd.n1949 10.6151
R10193 gnd.n3854 gnd.n1949 10.6151
R10194 gnd.n3855 gnd.n3854 10.6151
R10195 gnd.n3858 gnd.n3855 10.6151
R10196 gnd.n3858 gnd.n3857 10.6151
R10197 gnd.n3857 gnd.n3856 10.6151
R10198 gnd.n3856 gnd.n1900 10.6151
R10199 gnd.n2281 gnd.n1429 10.6151
R10200 gnd.n2284 gnd.n2281 10.6151
R10201 gnd.n2289 gnd.n2286 10.6151
R10202 gnd.n2290 gnd.n2289 10.6151
R10203 gnd.n2293 gnd.n2290 10.6151
R10204 gnd.n2294 gnd.n2293 10.6151
R10205 gnd.n2297 gnd.n2294 10.6151
R10206 gnd.n2298 gnd.n2297 10.6151
R10207 gnd.n2301 gnd.n2298 10.6151
R10208 gnd.n2302 gnd.n2301 10.6151
R10209 gnd.n2305 gnd.n2302 10.6151
R10210 gnd.n2306 gnd.n2305 10.6151
R10211 gnd.n2309 gnd.n2306 10.6151
R10212 gnd.n2310 gnd.n2309 10.6151
R10213 gnd.n2313 gnd.n2310 10.6151
R10214 gnd.n2314 gnd.n2313 10.6151
R10215 gnd.n2317 gnd.n2314 10.6151
R10216 gnd.n2318 gnd.n2317 10.6151
R10217 gnd.n2321 gnd.n2318 10.6151
R10218 gnd.n2322 gnd.n2321 10.6151
R10219 gnd.n2325 gnd.n2322 10.6151
R10220 gnd.n2326 gnd.n2325 10.6151
R10221 gnd.n2329 gnd.n2326 10.6151
R10222 gnd.n2330 gnd.n2329 10.6151
R10223 gnd.n2333 gnd.n2330 10.6151
R10224 gnd.n2334 gnd.n2333 10.6151
R10225 gnd.n2337 gnd.n2334 10.6151
R10226 gnd.n2338 gnd.n2337 10.6151
R10227 gnd.n2341 gnd.n2338 10.6151
R10228 gnd.n2342 gnd.n2341 10.6151
R10229 gnd.n4848 gnd.n4847 10.6151
R10230 gnd.n4847 gnd.n4846 10.6151
R10231 gnd.n4846 gnd.n4845 10.6151
R10232 gnd.n4845 gnd.n4843 10.6151
R10233 gnd.n4843 gnd.n4840 10.6151
R10234 gnd.n4840 gnd.n4839 10.6151
R10235 gnd.n4839 gnd.n4836 10.6151
R10236 gnd.n4836 gnd.n4835 10.6151
R10237 gnd.n4835 gnd.n4832 10.6151
R10238 gnd.n4832 gnd.n4831 10.6151
R10239 gnd.n4831 gnd.n4828 10.6151
R10240 gnd.n4828 gnd.n4827 10.6151
R10241 gnd.n4827 gnd.n4824 10.6151
R10242 gnd.n4824 gnd.n4823 10.6151
R10243 gnd.n4823 gnd.n4820 10.6151
R10244 gnd.n4820 gnd.n4819 10.6151
R10245 gnd.n4819 gnd.n4816 10.6151
R10246 gnd.n4816 gnd.n4815 10.6151
R10247 gnd.n4815 gnd.n4812 10.6151
R10248 gnd.n4812 gnd.n4811 10.6151
R10249 gnd.n4811 gnd.n4808 10.6151
R10250 gnd.n4808 gnd.n4807 10.6151
R10251 gnd.n4807 gnd.n4804 10.6151
R10252 gnd.n4804 gnd.n4803 10.6151
R10253 gnd.n4803 gnd.n4800 10.6151
R10254 gnd.n4800 gnd.n4799 10.6151
R10255 gnd.n4799 gnd.n4796 10.6151
R10256 gnd.n4796 gnd.n4795 10.6151
R10257 gnd.n4792 gnd.n4791 10.6151
R10258 gnd.n4791 gnd.n1430 10.6151
R10259 gnd.n4175 gnd.n4174 10.6151
R10260 gnd.n4174 gnd.n4171 10.6151
R10261 gnd.n4171 gnd.n4170 10.6151
R10262 gnd.n4170 gnd.n4167 10.6151
R10263 gnd.n4167 gnd.n4166 10.6151
R10264 gnd.n4166 gnd.n4163 10.6151
R10265 gnd.n4163 gnd.n4162 10.6151
R10266 gnd.n4162 gnd.n4159 10.6151
R10267 gnd.n4159 gnd.n4158 10.6151
R10268 gnd.n4158 gnd.n4155 10.6151
R10269 gnd.n4155 gnd.n4154 10.6151
R10270 gnd.n4154 gnd.n4151 10.6151
R10271 gnd.n4151 gnd.n4150 10.6151
R10272 gnd.n4150 gnd.n4147 10.6151
R10273 gnd.n4147 gnd.n4146 10.6151
R10274 gnd.n4146 gnd.n4143 10.6151
R10275 gnd.n4143 gnd.n4142 10.6151
R10276 gnd.n4142 gnd.n4139 10.6151
R10277 gnd.n4139 gnd.n4138 10.6151
R10278 gnd.n4138 gnd.n4135 10.6151
R10279 gnd.n4135 gnd.n4134 10.6151
R10280 gnd.n4134 gnd.n4131 10.6151
R10281 gnd.n4131 gnd.n4130 10.6151
R10282 gnd.n4130 gnd.n4127 10.6151
R10283 gnd.n4127 gnd.n4126 10.6151
R10284 gnd.n4126 gnd.n4123 10.6151
R10285 gnd.n4123 gnd.n4122 10.6151
R10286 gnd.n4122 gnd.n4119 10.6151
R10287 gnd.n4117 gnd.n4114 10.6151
R10288 gnd.n4114 gnd.n1862 10.6151
R10289 gnd.n4784 gnd.n4783 10.6151
R10290 gnd.n4783 gnd.n1489 10.6151
R10291 gnd.n2269 gnd.n1489 10.6151
R10292 gnd.n3272 gnd.n2269 10.6151
R10293 gnd.n3273 gnd.n3272 10.6151
R10294 gnd.n3274 gnd.n3273 10.6151
R10295 gnd.n3274 gnd.n2255 10.6151
R10296 gnd.n3307 gnd.n2255 10.6151
R10297 gnd.n3307 gnd.n3306 10.6151
R10298 gnd.n3306 gnd.n3305 10.6151
R10299 gnd.n3305 gnd.n3304 10.6151
R10300 gnd.n3304 gnd.n2256 10.6151
R10301 gnd.n2256 gnd.n2233 10.6151
R10302 gnd.n3344 gnd.n2233 10.6151
R10303 gnd.n3345 gnd.n3344 10.6151
R10304 gnd.n3355 gnd.n3345 10.6151
R10305 gnd.n3355 gnd.n3354 10.6151
R10306 gnd.n3354 gnd.n3353 10.6151
R10307 gnd.n3353 gnd.n3346 10.6151
R10308 gnd.n3347 gnd.n3346 10.6151
R10309 gnd.n3347 gnd.n2206 10.6151
R10310 gnd.n3413 gnd.n2206 10.6151
R10311 gnd.n3414 gnd.n3413 10.6151
R10312 gnd.n3415 gnd.n3414 10.6151
R10313 gnd.n3415 gnd.n2193 10.6151
R10314 gnd.n3431 gnd.n2193 10.6151
R10315 gnd.n3432 gnd.n3431 10.6151
R10316 gnd.n3434 gnd.n3432 10.6151
R10317 gnd.n3434 gnd.n3433 10.6151
R10318 gnd.n3433 gnd.n2173 10.6151
R10319 gnd.n3463 gnd.n2173 10.6151
R10320 gnd.n3464 gnd.n3463 10.6151
R10321 gnd.n3465 gnd.n3464 10.6151
R10322 gnd.n3465 gnd.n2156 10.6151
R10323 gnd.n3490 gnd.n2156 10.6151
R10324 gnd.n3491 gnd.n3490 10.6151
R10325 gnd.n3495 gnd.n3491 10.6151
R10326 gnd.n3495 gnd.n3494 10.6151
R10327 gnd.n3494 gnd.n3493 10.6151
R10328 gnd.n3493 gnd.n2133 10.6151
R10329 gnd.n3530 gnd.n2133 10.6151
R10330 gnd.n3531 gnd.n3530 10.6151
R10331 gnd.n3535 gnd.n3531 10.6151
R10332 gnd.n3535 gnd.n3534 10.6151
R10333 gnd.n3534 gnd.n3533 10.6151
R10334 gnd.n3533 gnd.n2111 10.6151
R10335 gnd.n3589 gnd.n2111 10.6151
R10336 gnd.n3590 gnd.n3589 10.6151
R10337 gnd.n3591 gnd.n3590 10.6151
R10338 gnd.n3591 gnd.n2096 10.6151
R10339 gnd.n3606 gnd.n2096 10.6151
R10340 gnd.n3607 gnd.n3606 10.6151
R10341 gnd.n3609 gnd.n3607 10.6151
R10342 gnd.n3609 gnd.n3608 10.6151
R10343 gnd.n3608 gnd.n2076 10.6151
R10344 gnd.n3633 gnd.n2076 10.6151
R10345 gnd.n3634 gnd.n3633 10.6151
R10346 gnd.n3643 gnd.n3634 10.6151
R10347 gnd.n3643 gnd.n3642 10.6151
R10348 gnd.n3642 gnd.n3641 10.6151
R10349 gnd.n3641 gnd.n3640 10.6151
R10350 gnd.n3640 gnd.n3635 10.6151
R10351 gnd.n3635 gnd.n2047 10.6151
R10352 gnd.n3704 gnd.n2047 10.6151
R10353 gnd.n3705 gnd.n3704 10.6151
R10354 gnd.n3706 gnd.n3705 10.6151
R10355 gnd.n3706 gnd.n2034 10.6151
R10356 gnd.n3723 gnd.n2034 10.6151
R10357 gnd.n3724 gnd.n3723 10.6151
R10358 gnd.n3725 gnd.n3724 10.6151
R10359 gnd.n3725 gnd.n2021 10.6151
R10360 gnd.n3754 gnd.n2021 10.6151
R10361 gnd.n3755 gnd.n3754 10.6151
R10362 gnd.n3756 gnd.n3755 10.6151
R10363 gnd.n3756 gnd.n2003 10.6151
R10364 gnd.n3771 gnd.n2003 10.6151
R10365 gnd.n3772 gnd.n3771 10.6151
R10366 gnd.n3774 gnd.n3772 10.6151
R10367 gnd.n3774 gnd.n3773 10.6151
R10368 gnd.n3773 gnd.n1986 10.6151
R10369 gnd.n3801 gnd.n1986 10.6151
R10370 gnd.n3802 gnd.n3801 10.6151
R10371 gnd.n3807 gnd.n3802 10.6151
R10372 gnd.n3807 gnd.n3806 10.6151
R10373 gnd.n3806 gnd.n3805 10.6151
R10374 gnd.n3805 gnd.n3804 10.6151
R10375 gnd.n3804 gnd.n1954 10.6151
R10376 gnd.n3847 gnd.n1954 10.6151
R10377 gnd.n3848 gnd.n3847 10.6151
R10378 gnd.n3850 gnd.n3848 10.6151
R10379 gnd.n3850 gnd.n3849 10.6151
R10380 gnd.n3849 gnd.n1905 10.6151
R10381 gnd.n4091 gnd.n1905 10.6151
R10382 gnd.n4092 gnd.n4091 10.6151
R10383 gnd.n4177 gnd.n4092 10.6151
R10384 gnd.n5552 gnd.t181 10.5161
R10385 gnd.n6438 gnd.t178 10.5161
R10386 gnd.n6445 gnd.t188 10.5161
R10387 gnd.n2803 gnd.t20 10.5161
R10388 gnd.n3420 gnd.t334 10.5161
R10389 gnd.t70 gnd.n3657 10.5161
R10390 gnd.n4558 gnd.t120 10.5161
R10391 gnd.n6400 gnd.n6384 10.4732
R10392 gnd.n6368 gnd.n6352 10.4732
R10393 gnd.n6336 gnd.n6320 10.4732
R10394 gnd.n6305 gnd.n6289 10.4732
R10395 gnd.n6273 gnd.n6257 10.4732
R10396 gnd.n6241 gnd.n6225 10.4732
R10397 gnd.n6209 gnd.n6193 10.4732
R10398 gnd.n6178 gnd.n6162 10.4732
R10399 gnd.n2258 gnd.n2252 10.1975
R10400 gnd.n2171 gnd.n2170 10.1975
R10401 gnd.n3498 gnd.n2151 10.1975
R10402 gnd.n3566 gnd.n2073 10.1975
R10403 gnd.n3638 gnd.n3637 10.1975
R10404 gnd.n3830 gnd.n1966 10.1975
R10405 gnd.n1919 gnd.t249 10.1975
R10406 gnd.n6137 gnd.t72 9.87883
R10407 gnd.n2840 gnd.t138 9.87883
R10408 gnd.n4467 gnd.t0 9.87883
R10409 gnd.n6404 gnd.n6403 9.69747
R10410 gnd.n6372 gnd.n6371 9.69747
R10411 gnd.n6340 gnd.n6339 9.69747
R10412 gnd.n6309 gnd.n6308 9.69747
R10413 gnd.n6277 gnd.n6276 9.69747
R10414 gnd.n6245 gnd.n6244 9.69747
R10415 gnd.n6213 gnd.n6212 9.69747
R10416 gnd.n6182 gnd.n6181 9.69747
R10417 gnd.n2355 gnd.n1491 9.56018
R10418 gnd.n3349 gnd.n3348 9.56018
R10419 gnd.n3403 gnd.n2195 9.56018
R10420 gnd.n3472 gnd.t44 9.56018
R10421 gnd.n3518 gnd.n2122 9.56018
R10422 gnd.n3559 gnd.n3558 9.56018
R10423 gnd.n3568 gnd.t96 9.56018
R10424 gnd.n3728 gnd.n3727 9.56018
R10425 gnd.n3650 gnd.n2005 9.56018
R10426 gnd.n6410 gnd.n6409 9.45567
R10427 gnd.n6378 gnd.n6377 9.45567
R10428 gnd.n6346 gnd.n6345 9.45567
R10429 gnd.n6315 gnd.n6314 9.45567
R10430 gnd.n6283 gnd.n6282 9.45567
R10431 gnd.n6251 gnd.n6250 9.45567
R10432 gnd.n6219 gnd.n6218 9.45567
R10433 gnd.n6188 gnd.n6187 9.45567
R10434 gnd.n4372 gnd.n1850 9.30959
R10435 gnd.n7603 gnd.n279 9.30959
R10436 gnd.n5088 gnd.n5087 9.30959
R10437 gnd.n3009 gnd.n2973 9.30959
R10438 gnd.n6409 gnd.n6408 9.3005
R10439 gnd.n6382 gnd.n6381 9.3005
R10440 gnd.n6403 gnd.n6402 9.3005
R10441 gnd.n6401 gnd.n6400 9.3005
R10442 gnd.n6386 gnd.n6385 9.3005
R10443 gnd.n6395 gnd.n6394 9.3005
R10444 gnd.n6393 gnd.n6392 9.3005
R10445 gnd.n6377 gnd.n6376 9.3005
R10446 gnd.n6350 gnd.n6349 9.3005
R10447 gnd.n6371 gnd.n6370 9.3005
R10448 gnd.n6369 gnd.n6368 9.3005
R10449 gnd.n6354 gnd.n6353 9.3005
R10450 gnd.n6363 gnd.n6362 9.3005
R10451 gnd.n6361 gnd.n6360 9.3005
R10452 gnd.n6345 gnd.n6344 9.3005
R10453 gnd.n6318 gnd.n6317 9.3005
R10454 gnd.n6339 gnd.n6338 9.3005
R10455 gnd.n6337 gnd.n6336 9.3005
R10456 gnd.n6322 gnd.n6321 9.3005
R10457 gnd.n6331 gnd.n6330 9.3005
R10458 gnd.n6329 gnd.n6328 9.3005
R10459 gnd.n6314 gnd.n6313 9.3005
R10460 gnd.n6287 gnd.n6286 9.3005
R10461 gnd.n6308 gnd.n6307 9.3005
R10462 gnd.n6306 gnd.n6305 9.3005
R10463 gnd.n6291 gnd.n6290 9.3005
R10464 gnd.n6300 gnd.n6299 9.3005
R10465 gnd.n6298 gnd.n6297 9.3005
R10466 gnd.n6282 gnd.n6281 9.3005
R10467 gnd.n6255 gnd.n6254 9.3005
R10468 gnd.n6276 gnd.n6275 9.3005
R10469 gnd.n6274 gnd.n6273 9.3005
R10470 gnd.n6259 gnd.n6258 9.3005
R10471 gnd.n6268 gnd.n6267 9.3005
R10472 gnd.n6266 gnd.n6265 9.3005
R10473 gnd.n6250 gnd.n6249 9.3005
R10474 gnd.n6223 gnd.n6222 9.3005
R10475 gnd.n6244 gnd.n6243 9.3005
R10476 gnd.n6242 gnd.n6241 9.3005
R10477 gnd.n6227 gnd.n6226 9.3005
R10478 gnd.n6236 gnd.n6235 9.3005
R10479 gnd.n6234 gnd.n6233 9.3005
R10480 gnd.n6218 gnd.n6217 9.3005
R10481 gnd.n6191 gnd.n6190 9.3005
R10482 gnd.n6212 gnd.n6211 9.3005
R10483 gnd.n6210 gnd.n6209 9.3005
R10484 gnd.n6195 gnd.n6194 9.3005
R10485 gnd.n6204 gnd.n6203 9.3005
R10486 gnd.n6202 gnd.n6201 9.3005
R10487 gnd.n6187 gnd.n6186 9.3005
R10488 gnd.n6160 gnd.n6159 9.3005
R10489 gnd.n6181 gnd.n6180 9.3005
R10490 gnd.n6179 gnd.n6178 9.3005
R10491 gnd.n6164 gnd.n6163 9.3005
R10492 gnd.n6173 gnd.n6172 9.3005
R10493 gnd.n6171 gnd.n6170 9.3005
R10494 gnd.n6539 gnd.n5171 9.3005
R10495 gnd.n6538 gnd.n5173 9.3005
R10496 gnd.n5177 gnd.n5174 9.3005
R10497 gnd.n6533 gnd.n5178 9.3005
R10498 gnd.n6532 gnd.n5179 9.3005
R10499 gnd.n6531 gnd.n5180 9.3005
R10500 gnd.n5184 gnd.n5181 9.3005
R10501 gnd.n6526 gnd.n5185 9.3005
R10502 gnd.n6525 gnd.n5186 9.3005
R10503 gnd.n6524 gnd.n5187 9.3005
R10504 gnd.n5191 gnd.n5188 9.3005
R10505 gnd.n6519 gnd.n5192 9.3005
R10506 gnd.n6518 gnd.n5193 9.3005
R10507 gnd.n6517 gnd.n5194 9.3005
R10508 gnd.n5199 gnd.n5197 9.3005
R10509 gnd.n6512 gnd.n6511 9.3005
R10510 gnd.n6541 gnd.n6540 9.3005
R10511 gnd.n5819 gnd.n5818 9.3005
R10512 gnd.n5820 gnd.n5522 9.3005
R10513 gnd.n5822 gnd.n5821 9.3005
R10514 gnd.n5503 gnd.n5502 9.3005
R10515 gnd.n5849 gnd.n5848 9.3005
R10516 gnd.n5850 gnd.n5501 9.3005
R10517 gnd.n5854 gnd.n5851 9.3005
R10518 gnd.n5853 gnd.n5852 9.3005
R10519 gnd.n5477 gnd.n5476 9.3005
R10520 gnd.n5883 gnd.n5882 9.3005
R10521 gnd.n5884 gnd.n5475 9.3005
R10522 gnd.n5891 gnd.n5885 9.3005
R10523 gnd.n5890 gnd.n5886 9.3005
R10524 gnd.n5889 gnd.n5887 9.3005
R10525 gnd.n5444 gnd.n5443 9.3005
R10526 gnd.n5944 gnd.n5943 9.3005
R10527 gnd.n5945 gnd.n5442 9.3005
R10528 gnd.n5949 gnd.n5946 9.3005
R10529 gnd.n5948 gnd.n5947 9.3005
R10530 gnd.n5417 gnd.n5416 9.3005
R10531 gnd.n5984 gnd.n5983 9.3005
R10532 gnd.n5985 gnd.n5415 9.3005
R10533 gnd.n5989 gnd.n5986 9.3005
R10534 gnd.n5988 gnd.n5987 9.3005
R10535 gnd.n5326 gnd.n5325 9.3005
R10536 gnd.n6029 gnd.n6028 9.3005
R10537 gnd.n6030 gnd.n5324 9.3005
R10538 gnd.n6034 gnd.n6031 9.3005
R10539 gnd.n6033 gnd.n6032 9.3005
R10540 gnd.n5298 gnd.n5297 9.3005
R10541 gnd.n6068 gnd.n6067 9.3005
R10542 gnd.n6069 gnd.n5296 9.3005
R10543 gnd.n6076 gnd.n6070 9.3005
R10544 gnd.n6075 gnd.n6071 9.3005
R10545 gnd.n6074 gnd.n6072 9.3005
R10546 gnd.n5268 gnd.n5267 9.3005
R10547 gnd.n6125 gnd.n6124 9.3005
R10548 gnd.n6126 gnd.n5266 9.3005
R10549 gnd.n6134 gnd.n6127 9.3005
R10550 gnd.n6133 gnd.n6128 9.3005
R10551 gnd.n6132 gnd.n6130 9.3005
R10552 gnd.n6129 gnd.n984 9.3005
R10553 gnd.n6571 gnd.n985 9.3005
R10554 gnd.n6570 gnd.n986 9.3005
R10555 gnd.n6569 gnd.n987 9.3005
R10556 gnd.n1009 gnd.n988 9.3005
R10557 gnd.n1010 gnd.n1008 9.3005
R10558 gnd.n6557 gnd.n1011 9.3005
R10559 gnd.n6556 gnd.n1012 9.3005
R10560 gnd.n6555 gnd.n1013 9.3005
R10561 gnd.n5169 gnd.n1014 9.3005
R10562 gnd.n5170 gnd.n5168 9.3005
R10563 gnd.n6543 gnd.n6542 9.3005
R10564 gnd.n5524 gnd.n5523 9.3005
R10565 gnd.n5764 gnd.n5763 9.3005
R10566 gnd.n5767 gnd.n5759 9.3005
R10567 gnd.n5768 gnd.n5758 9.3005
R10568 gnd.n5771 gnd.n5757 9.3005
R10569 gnd.n5772 gnd.n5756 9.3005
R10570 gnd.n5775 gnd.n5755 9.3005
R10571 gnd.n5776 gnd.n5754 9.3005
R10572 gnd.n5779 gnd.n5753 9.3005
R10573 gnd.n5780 gnd.n5752 9.3005
R10574 gnd.n5783 gnd.n5751 9.3005
R10575 gnd.n5784 gnd.n5750 9.3005
R10576 gnd.n5787 gnd.n5749 9.3005
R10577 gnd.n5789 gnd.n5748 9.3005
R10578 gnd.n5790 gnd.n5747 9.3005
R10579 gnd.n5791 gnd.n5746 9.3005
R10580 gnd.n5792 gnd.n5745 9.3005
R10581 gnd.n5760 gnd.n5541 9.3005
R10582 gnd.n5809 gnd.n5532 9.3005
R10583 gnd.n5811 gnd.n5810 9.3005
R10584 gnd.n5519 gnd.n5514 9.3005
R10585 gnd.n5832 gnd.n5513 9.3005
R10586 gnd.n5835 gnd.n5834 9.3005
R10587 gnd.n5837 gnd.n5836 9.3005
R10588 gnd.n5840 gnd.n5496 9.3005
R10589 gnd.n5838 gnd.n5494 9.3005
R10590 gnd.n5860 gnd.n5492 9.3005
R10591 gnd.n5864 gnd.n5863 9.3005
R10592 gnd.n5862 gnd.n5467 9.3005
R10593 gnd.n5898 gnd.n5466 9.3005
R10594 gnd.n5901 gnd.n5900 9.3005
R10595 gnd.n5464 gnd.n5463 9.3005
R10596 gnd.n5907 gnd.n5461 9.3005
R10597 gnd.n5909 gnd.n5908 9.3005
R10598 gnd.n5435 gnd.n5434 9.3005
R10599 gnd.n5958 gnd.n5957 9.3005
R10600 gnd.n5959 gnd.n5428 9.3005
R10601 gnd.n5967 gnd.n5427 9.3005
R10602 gnd.n5970 gnd.n5969 9.3005
R10603 gnd.n5972 gnd.n5971 9.3005
R10604 gnd.n5975 gnd.n5410 9.3005
R10605 gnd.n5973 gnd.n5408 9.3005
R10606 gnd.n5995 gnd.n5406 9.3005
R10607 gnd.n5997 gnd.n5996 9.3005
R10608 gnd.n5316 gnd.n5315 9.3005
R10609 gnd.n6043 gnd.n6042 9.3005
R10610 gnd.n6044 gnd.n5309 9.3005
R10611 gnd.n6052 gnd.n5308 9.3005
R10612 gnd.n6055 gnd.n6054 9.3005
R10613 gnd.n6057 gnd.n6056 9.3005
R10614 gnd.n6059 gnd.n5291 9.3005
R10615 gnd.n5289 gnd.n5287 9.3005
R10616 gnd.n6084 gnd.n6083 9.3005
R10617 gnd.n5273 gnd.n5272 9.3005
R10618 gnd.n6117 gnd.n6116 9.3005
R10619 gnd.n6118 gnd.n5259 9.3005
R10620 gnd.n6141 gnd.n5258 9.3005
R10621 gnd.n6144 gnd.n6143 9.3005
R10622 gnd.n5255 gnd.n5254 9.3005
R10623 gnd.n6148 gnd.n5256 9.3005
R10624 gnd.n6150 gnd.n6149 9.3005
R10625 gnd.n6435 gnd.n6152 9.3005
R10626 gnd.n6434 gnd.n6154 9.3005
R10627 gnd.n6433 gnd.n6155 9.3005
R10628 gnd.n6430 gnd.n6156 9.3005
R10629 gnd.n6429 gnd.n6157 9.3005
R10630 gnd.n6428 gnd.n6415 9.3005
R10631 gnd.n6425 gnd.n6417 9.3005
R10632 gnd.n6424 gnd.n6418 9.3005
R10633 gnd.n6421 gnd.n6419 9.3005
R10634 gnd.n6420 gnd.n5200 9.3005
R10635 gnd.n5808 gnd.n5535 9.3005
R10636 gnd.n6507 gnd.n5201 9.3005
R10637 gnd.n6506 gnd.n5203 9.3005
R10638 gnd.n5207 gnd.n5204 9.3005
R10639 gnd.n6501 gnd.n5208 9.3005
R10640 gnd.n6500 gnd.n5209 9.3005
R10641 gnd.n6499 gnd.n5210 9.3005
R10642 gnd.n5214 gnd.n5211 9.3005
R10643 gnd.n6494 gnd.n5215 9.3005
R10644 gnd.n6493 gnd.n5216 9.3005
R10645 gnd.n6492 gnd.n5217 9.3005
R10646 gnd.n5221 gnd.n5218 9.3005
R10647 gnd.n6487 gnd.n5222 9.3005
R10648 gnd.n6486 gnd.n5223 9.3005
R10649 gnd.n6485 gnd.n5224 9.3005
R10650 gnd.n5228 gnd.n5225 9.3005
R10651 gnd.n6480 gnd.n5229 9.3005
R10652 gnd.n6479 gnd.n5230 9.3005
R10653 gnd.n6478 gnd.n5231 9.3005
R10654 gnd.n5235 gnd.n5232 9.3005
R10655 gnd.n6473 gnd.n5236 9.3005
R10656 gnd.n6472 gnd.n5237 9.3005
R10657 gnd.n6471 gnd.n5238 9.3005
R10658 gnd.n5245 gnd.n5243 9.3005
R10659 gnd.n6466 gnd.n5246 9.3005
R10660 gnd.n6465 gnd.n5247 9.3005
R10661 gnd.n6464 gnd.n6461 9.3005
R10662 gnd.n6509 gnd.n6508 9.3005
R10663 gnd.n6005 gnd.n6004 9.3005
R10664 gnd.n6006 gnd.n5332 9.3005
R10665 gnd.n6023 gnd.n6007 9.3005
R10666 gnd.n6022 gnd.n6008 9.3005
R10667 gnd.n6021 gnd.n6009 9.3005
R10668 gnd.n6019 gnd.n6010 9.3005
R10669 gnd.n6018 gnd.n6011 9.3005
R10670 gnd.n6016 gnd.n6012 9.3005
R10671 gnd.n6015 gnd.n6013 9.3005
R10672 gnd.n5280 gnd.n5279 9.3005
R10673 gnd.n6091 gnd.n6090 9.3005
R10674 gnd.n6092 gnd.n5278 9.3005
R10675 gnd.n6109 gnd.n6093 9.3005
R10676 gnd.n6108 gnd.n6094 9.3005
R10677 gnd.n6107 gnd.n6095 9.3005
R10678 gnd.n6106 gnd.n6096 9.3005
R10679 gnd.n6104 gnd.n6097 9.3005
R10680 gnd.n6103 gnd.n6098 9.3005
R10681 gnd.n6100 gnd.n6099 9.3005
R10682 gnd.n5253 gnd.n5252 9.3005
R10683 gnd.n6442 gnd.n6441 9.3005
R10684 gnd.n6443 gnd.n5251 9.3005
R10685 gnd.n6447 gnd.n6444 9.3005
R10686 gnd.n6448 gnd.n5250 9.3005
R10687 gnd.n6452 gnd.n6451 9.3005
R10688 gnd.n6453 gnd.n5249 9.3005
R10689 gnd.n6455 gnd.n6454 9.3005
R10690 gnd.n6458 gnd.n5248 9.3005
R10691 gnd.n6460 gnd.n6459 9.3005
R10692 gnd.n5678 gnd.n5572 9.3005
R10693 gnd.n5680 gnd.n5679 9.3005
R10694 gnd.n5562 gnd.n5561 9.3005
R10695 gnd.n5693 gnd.n5692 9.3005
R10696 gnd.n5694 gnd.n5560 9.3005
R10697 gnd.n5696 gnd.n5695 9.3005
R10698 gnd.n5549 gnd.n5548 9.3005
R10699 gnd.n5709 gnd.n5708 9.3005
R10700 gnd.n5710 gnd.n5547 9.3005
R10701 gnd.n5734 gnd.n5711 9.3005
R10702 gnd.n5733 gnd.n5712 9.3005
R10703 gnd.n5732 gnd.n5713 9.3005
R10704 gnd.n5731 gnd.n5714 9.3005
R10705 gnd.n5729 gnd.n5715 9.3005
R10706 gnd.n5728 gnd.n5716 9.3005
R10707 gnd.n5726 gnd.n5717 9.3005
R10708 gnd.n5725 gnd.n5718 9.3005
R10709 gnd.n5723 gnd.n5719 9.3005
R10710 gnd.n5722 gnd.n5720 9.3005
R10711 gnd.n5484 gnd.n5483 9.3005
R10712 gnd.n5872 gnd.n5871 9.3005
R10713 gnd.n5873 gnd.n5482 9.3005
R10714 gnd.n5877 gnd.n5874 9.3005
R10715 gnd.n5876 gnd.n5875 9.3005
R10716 gnd.n5451 gnd.n5450 9.3005
R10717 gnd.n5919 gnd.n5918 9.3005
R10718 gnd.n5920 gnd.n5449 9.3005
R10719 gnd.n5922 gnd.n5921 9.3005
R10720 gnd.n5677 gnd.n5676 9.3005
R10721 gnd.n5617 gnd.n5616 9.3005
R10722 gnd.n5622 gnd.n5614 9.3005
R10723 gnd.n5623 gnd.n5613 9.3005
R10724 gnd.n5625 gnd.n5610 9.3005
R10725 gnd.n5609 gnd.n5607 9.3005
R10726 gnd.n5631 gnd.n5606 9.3005
R10727 gnd.n5632 gnd.n5605 9.3005
R10728 gnd.n5633 gnd.n5604 9.3005
R10729 gnd.n5603 gnd.n5601 9.3005
R10730 gnd.n5639 gnd.n5600 9.3005
R10731 gnd.n5640 gnd.n5599 9.3005
R10732 gnd.n5641 gnd.n5598 9.3005
R10733 gnd.n5597 gnd.n5595 9.3005
R10734 gnd.n5647 gnd.n5594 9.3005
R10735 gnd.n5648 gnd.n5593 9.3005
R10736 gnd.n5649 gnd.n5592 9.3005
R10737 gnd.n5591 gnd.n5589 9.3005
R10738 gnd.n5655 gnd.n5588 9.3005
R10739 gnd.n5656 gnd.n5587 9.3005
R10740 gnd.n5657 gnd.n5586 9.3005
R10741 gnd.n5585 gnd.n5583 9.3005
R10742 gnd.n5662 gnd.n5582 9.3005
R10743 gnd.n5663 gnd.n5581 9.3005
R10744 gnd.n5580 gnd.n5578 9.3005
R10745 gnd.n5668 gnd.n5577 9.3005
R10746 gnd.n5670 gnd.n5669 9.3005
R10747 gnd.n5615 gnd.n5573 9.3005
R10748 gnd.n5568 gnd.n5567 9.3005
R10749 gnd.n5685 gnd.n5684 9.3005
R10750 gnd.n5686 gnd.n5566 9.3005
R10751 gnd.n5688 gnd.n5687 9.3005
R10752 gnd.n5556 gnd.n5555 9.3005
R10753 gnd.n5701 gnd.n5700 9.3005
R10754 gnd.n5702 gnd.n5554 9.3005
R10755 gnd.n5704 gnd.n5703 9.3005
R10756 gnd.n5543 gnd.n5542 9.3005
R10757 gnd.n5799 gnd.n5798 9.3005
R10758 gnd.n5801 gnd.n5540 9.3005
R10759 gnd.n5803 gnd.n5802 9.3005
R10760 gnd.n5534 gnd.n5531 9.3005
R10761 gnd.n5813 gnd.n5812 9.3005
R10762 gnd.n5533 gnd.n5515 9.3005
R10763 gnd.n5831 gnd.n5830 9.3005
R10764 gnd.n5833 gnd.n5511 9.3005
R10765 gnd.n5843 gnd.n5512 9.3005
R10766 gnd.n5842 gnd.n5841 9.3005
R10767 gnd.n5839 gnd.n5490 9.3005
R10768 gnd.n5867 gnd.n5491 9.3005
R10769 gnd.n5866 gnd.n5865 9.3005
R10770 gnd.n5493 gnd.n5468 9.3005
R10771 gnd.n5897 gnd.n5896 9.3005
R10772 gnd.n5899 gnd.n5458 9.3005
R10773 gnd.n5914 gnd.n5459 9.3005
R10774 gnd.n5913 gnd.n5460 9.3005
R10775 gnd.n5912 gnd.n5910 9.3005
R10776 gnd.n5462 gnd.n5436 9.3005
R10777 gnd.n5955 gnd.n5954 9.3005
R10778 gnd.n5956 gnd.n5429 9.3005
R10779 gnd.n5966 gnd.n5965 9.3005
R10780 gnd.n5968 gnd.n5425 9.3005
R10781 gnd.n5978 gnd.n5426 9.3005
R10782 gnd.n5977 gnd.n5976 9.3005
R10783 gnd.n5974 gnd.n5404 9.3005
R10784 gnd.n6000 gnd.n5405 9.3005
R10785 gnd.n5999 gnd.n5998 9.3005
R10786 gnd.n5407 gnd.n5317 9.3005
R10787 gnd.n6040 gnd.n6039 9.3005
R10788 gnd.n6041 gnd.n5310 9.3005
R10789 gnd.n6051 gnd.n6050 9.3005
R10790 gnd.n6053 gnd.n5306 9.3005
R10791 gnd.n6062 gnd.n5307 9.3005
R10792 gnd.n6061 gnd.n6060 9.3005
R10793 gnd.n6058 gnd.n5286 9.3005
R10794 gnd.n6086 gnd.n6085 9.3005
R10795 gnd.n5288 gnd.n5274 9.3005
R10796 gnd.n6114 gnd.n6113 9.3005
R10797 gnd.n6115 gnd.n5260 9.3005
R10798 gnd.n6140 gnd.n6139 9.3005
R10799 gnd.n6142 gnd.n973 9.3005
R10800 gnd.n6578 gnd.n974 9.3005
R10801 gnd.n6577 gnd.n975 9.3005
R10802 gnd.n6576 gnd.n976 9.3005
R10803 gnd.n6151 gnd.n977 9.3005
R10804 gnd.n6153 gnd.n996 9.3005
R10805 gnd.n6564 gnd.n997 9.3005
R10806 gnd.n6563 gnd.n998 9.3005
R10807 gnd.n6562 gnd.n999 9.3005
R10808 gnd.n6414 gnd.n1000 9.3005
R10809 gnd.n6416 gnd.n1022 9.3005
R10810 gnd.n6550 gnd.n1023 9.3005
R10811 gnd.n6549 gnd.n1024 9.3005
R10812 gnd.n6548 gnd.n1025 9.3005
R10813 gnd.n5672 gnd.n5671 9.3005
R10814 gnd.n799 gnd.n798 9.3005
R10815 gnd.n6754 gnd.n6753 9.3005
R10816 gnd.n6755 gnd.n797 9.3005
R10817 gnd.n6757 gnd.n6756 9.3005
R10818 gnd.n793 gnd.n792 9.3005
R10819 gnd.n6764 gnd.n6763 9.3005
R10820 gnd.n6765 gnd.n791 9.3005
R10821 gnd.n6767 gnd.n6766 9.3005
R10822 gnd.n787 gnd.n786 9.3005
R10823 gnd.n6774 gnd.n6773 9.3005
R10824 gnd.n6775 gnd.n785 9.3005
R10825 gnd.n6777 gnd.n6776 9.3005
R10826 gnd.n781 gnd.n780 9.3005
R10827 gnd.n6784 gnd.n6783 9.3005
R10828 gnd.n6785 gnd.n779 9.3005
R10829 gnd.n6787 gnd.n6786 9.3005
R10830 gnd.n775 gnd.n774 9.3005
R10831 gnd.n6794 gnd.n6793 9.3005
R10832 gnd.n6795 gnd.n773 9.3005
R10833 gnd.n6797 gnd.n6796 9.3005
R10834 gnd.n769 gnd.n768 9.3005
R10835 gnd.n6804 gnd.n6803 9.3005
R10836 gnd.n6805 gnd.n767 9.3005
R10837 gnd.n6807 gnd.n6806 9.3005
R10838 gnd.n763 gnd.n762 9.3005
R10839 gnd.n6814 gnd.n6813 9.3005
R10840 gnd.n6815 gnd.n761 9.3005
R10841 gnd.n6817 gnd.n6816 9.3005
R10842 gnd.n757 gnd.n756 9.3005
R10843 gnd.n6824 gnd.n6823 9.3005
R10844 gnd.n6825 gnd.n755 9.3005
R10845 gnd.n6827 gnd.n6826 9.3005
R10846 gnd.n751 gnd.n750 9.3005
R10847 gnd.n6834 gnd.n6833 9.3005
R10848 gnd.n6835 gnd.n749 9.3005
R10849 gnd.n6837 gnd.n6836 9.3005
R10850 gnd.n745 gnd.n744 9.3005
R10851 gnd.n6844 gnd.n6843 9.3005
R10852 gnd.n6845 gnd.n743 9.3005
R10853 gnd.n6847 gnd.n6846 9.3005
R10854 gnd.n739 gnd.n738 9.3005
R10855 gnd.n6854 gnd.n6853 9.3005
R10856 gnd.n6855 gnd.n737 9.3005
R10857 gnd.n6857 gnd.n6856 9.3005
R10858 gnd.n733 gnd.n732 9.3005
R10859 gnd.n6864 gnd.n6863 9.3005
R10860 gnd.n6865 gnd.n731 9.3005
R10861 gnd.n6867 gnd.n6866 9.3005
R10862 gnd.n727 gnd.n726 9.3005
R10863 gnd.n6874 gnd.n6873 9.3005
R10864 gnd.n6875 gnd.n725 9.3005
R10865 gnd.n6877 gnd.n6876 9.3005
R10866 gnd.n721 gnd.n720 9.3005
R10867 gnd.n6884 gnd.n6883 9.3005
R10868 gnd.n6885 gnd.n719 9.3005
R10869 gnd.n6887 gnd.n6886 9.3005
R10870 gnd.n715 gnd.n714 9.3005
R10871 gnd.n6894 gnd.n6893 9.3005
R10872 gnd.n6895 gnd.n713 9.3005
R10873 gnd.n6897 gnd.n6896 9.3005
R10874 gnd.n709 gnd.n708 9.3005
R10875 gnd.n6904 gnd.n6903 9.3005
R10876 gnd.n6905 gnd.n707 9.3005
R10877 gnd.n6907 gnd.n6906 9.3005
R10878 gnd.n703 gnd.n702 9.3005
R10879 gnd.n6914 gnd.n6913 9.3005
R10880 gnd.n6915 gnd.n701 9.3005
R10881 gnd.n6917 gnd.n6916 9.3005
R10882 gnd.n697 gnd.n696 9.3005
R10883 gnd.n6924 gnd.n6923 9.3005
R10884 gnd.n6925 gnd.n695 9.3005
R10885 gnd.n6927 gnd.n6926 9.3005
R10886 gnd.n691 gnd.n690 9.3005
R10887 gnd.n6934 gnd.n6933 9.3005
R10888 gnd.n6935 gnd.n689 9.3005
R10889 gnd.n6937 gnd.n6936 9.3005
R10890 gnd.n685 gnd.n684 9.3005
R10891 gnd.n6944 gnd.n6943 9.3005
R10892 gnd.n6945 gnd.n683 9.3005
R10893 gnd.n6947 gnd.n6946 9.3005
R10894 gnd.n679 gnd.n678 9.3005
R10895 gnd.n6954 gnd.n6953 9.3005
R10896 gnd.n6955 gnd.n677 9.3005
R10897 gnd.n6957 gnd.n6956 9.3005
R10898 gnd.n673 gnd.n672 9.3005
R10899 gnd.n6964 gnd.n6963 9.3005
R10900 gnd.n6965 gnd.n671 9.3005
R10901 gnd.n6967 gnd.n6966 9.3005
R10902 gnd.n667 gnd.n666 9.3005
R10903 gnd.n6974 gnd.n6973 9.3005
R10904 gnd.n6975 gnd.n665 9.3005
R10905 gnd.n6977 gnd.n6976 9.3005
R10906 gnd.n661 gnd.n660 9.3005
R10907 gnd.n6984 gnd.n6983 9.3005
R10908 gnd.n6985 gnd.n659 9.3005
R10909 gnd.n6987 gnd.n6986 9.3005
R10910 gnd.n655 gnd.n654 9.3005
R10911 gnd.n6994 gnd.n6993 9.3005
R10912 gnd.n6995 gnd.n653 9.3005
R10913 gnd.n6997 gnd.n6996 9.3005
R10914 gnd.n649 gnd.n648 9.3005
R10915 gnd.n7004 gnd.n7003 9.3005
R10916 gnd.n7005 gnd.n647 9.3005
R10917 gnd.n7007 gnd.n7006 9.3005
R10918 gnd.n643 gnd.n642 9.3005
R10919 gnd.n7014 gnd.n7013 9.3005
R10920 gnd.n7015 gnd.n641 9.3005
R10921 gnd.n7017 gnd.n7016 9.3005
R10922 gnd.n637 gnd.n636 9.3005
R10923 gnd.n7024 gnd.n7023 9.3005
R10924 gnd.n7025 gnd.n635 9.3005
R10925 gnd.n7027 gnd.n7026 9.3005
R10926 gnd.n631 gnd.n630 9.3005
R10927 gnd.n7034 gnd.n7033 9.3005
R10928 gnd.n7035 gnd.n629 9.3005
R10929 gnd.n7037 gnd.n7036 9.3005
R10930 gnd.n625 gnd.n624 9.3005
R10931 gnd.n7044 gnd.n7043 9.3005
R10932 gnd.n7045 gnd.n623 9.3005
R10933 gnd.n7047 gnd.n7046 9.3005
R10934 gnd.n619 gnd.n618 9.3005
R10935 gnd.n7054 gnd.n7053 9.3005
R10936 gnd.n7055 gnd.n617 9.3005
R10937 gnd.n7057 gnd.n7056 9.3005
R10938 gnd.n613 gnd.n612 9.3005
R10939 gnd.n7064 gnd.n7063 9.3005
R10940 gnd.n7065 gnd.n611 9.3005
R10941 gnd.n7067 gnd.n7066 9.3005
R10942 gnd.n607 gnd.n606 9.3005
R10943 gnd.n7074 gnd.n7073 9.3005
R10944 gnd.n7075 gnd.n605 9.3005
R10945 gnd.n7077 gnd.n7076 9.3005
R10946 gnd.n601 gnd.n600 9.3005
R10947 gnd.n7084 gnd.n7083 9.3005
R10948 gnd.n7085 gnd.n599 9.3005
R10949 gnd.n7087 gnd.n7086 9.3005
R10950 gnd.n595 gnd.n594 9.3005
R10951 gnd.n7094 gnd.n7093 9.3005
R10952 gnd.n7095 gnd.n593 9.3005
R10953 gnd.n7097 gnd.n7096 9.3005
R10954 gnd.n589 gnd.n588 9.3005
R10955 gnd.n7104 gnd.n7103 9.3005
R10956 gnd.n7105 gnd.n587 9.3005
R10957 gnd.n7107 gnd.n7106 9.3005
R10958 gnd.n583 gnd.n582 9.3005
R10959 gnd.n7114 gnd.n7113 9.3005
R10960 gnd.n7115 gnd.n581 9.3005
R10961 gnd.n7117 gnd.n7116 9.3005
R10962 gnd.n577 gnd.n576 9.3005
R10963 gnd.n7124 gnd.n7123 9.3005
R10964 gnd.n7125 gnd.n575 9.3005
R10965 gnd.n7127 gnd.n7126 9.3005
R10966 gnd.n571 gnd.n570 9.3005
R10967 gnd.n7134 gnd.n7133 9.3005
R10968 gnd.n7135 gnd.n569 9.3005
R10969 gnd.n7137 gnd.n7136 9.3005
R10970 gnd.n565 gnd.n564 9.3005
R10971 gnd.n7144 gnd.n7143 9.3005
R10972 gnd.n7145 gnd.n563 9.3005
R10973 gnd.n7147 gnd.n7146 9.3005
R10974 gnd.n559 gnd.n558 9.3005
R10975 gnd.n7154 gnd.n7153 9.3005
R10976 gnd.n7155 gnd.n557 9.3005
R10977 gnd.n7157 gnd.n7156 9.3005
R10978 gnd.n553 gnd.n552 9.3005
R10979 gnd.n7164 gnd.n7163 9.3005
R10980 gnd.n7165 gnd.n551 9.3005
R10981 gnd.n7167 gnd.n7166 9.3005
R10982 gnd.n547 gnd.n546 9.3005
R10983 gnd.n7174 gnd.n7173 9.3005
R10984 gnd.n7175 gnd.n545 9.3005
R10985 gnd.n7177 gnd.n7176 9.3005
R10986 gnd.n541 gnd.n540 9.3005
R10987 gnd.n7184 gnd.n7183 9.3005
R10988 gnd.n7185 gnd.n539 9.3005
R10989 gnd.n7187 gnd.n7186 9.3005
R10990 gnd.n535 gnd.n534 9.3005
R10991 gnd.n7194 gnd.n7193 9.3005
R10992 gnd.n7195 gnd.n533 9.3005
R10993 gnd.n7197 gnd.n7196 9.3005
R10994 gnd.n529 gnd.n528 9.3005
R10995 gnd.n7204 gnd.n7203 9.3005
R10996 gnd.n7207 gnd.n7206 9.3005
R10997 gnd.n523 gnd.n522 9.3005
R10998 gnd.n7214 gnd.n7213 9.3005
R10999 gnd.n7215 gnd.n521 9.3005
R11000 gnd.n7217 gnd.n7216 9.3005
R11001 gnd.n517 gnd.n516 9.3005
R11002 gnd.n7224 gnd.n7223 9.3005
R11003 gnd.n7225 gnd.n515 9.3005
R11004 gnd.n7227 gnd.n7226 9.3005
R11005 gnd.n511 gnd.n510 9.3005
R11006 gnd.n7234 gnd.n7233 9.3005
R11007 gnd.n7235 gnd.n509 9.3005
R11008 gnd.n7237 gnd.n7236 9.3005
R11009 gnd.n505 gnd.n504 9.3005
R11010 gnd.n7244 gnd.n7243 9.3005
R11011 gnd.n7245 gnd.n503 9.3005
R11012 gnd.n7247 gnd.n7246 9.3005
R11013 gnd.n499 gnd.n498 9.3005
R11014 gnd.n7254 gnd.n7253 9.3005
R11015 gnd.n7255 gnd.n497 9.3005
R11016 gnd.n7257 gnd.n7256 9.3005
R11017 gnd.n493 gnd.n492 9.3005
R11018 gnd.n7264 gnd.n7263 9.3005
R11019 gnd.n7265 gnd.n491 9.3005
R11020 gnd.n7267 gnd.n7266 9.3005
R11021 gnd.n487 gnd.n486 9.3005
R11022 gnd.n7274 gnd.n7273 9.3005
R11023 gnd.n7275 gnd.n485 9.3005
R11024 gnd.n7277 gnd.n7276 9.3005
R11025 gnd.n481 gnd.n480 9.3005
R11026 gnd.n7284 gnd.n7283 9.3005
R11027 gnd.n7285 gnd.n479 9.3005
R11028 gnd.n7287 gnd.n7286 9.3005
R11029 gnd.n475 gnd.n474 9.3005
R11030 gnd.n7294 gnd.n7293 9.3005
R11031 gnd.n7295 gnd.n473 9.3005
R11032 gnd.n7297 gnd.n7296 9.3005
R11033 gnd.n469 gnd.n468 9.3005
R11034 gnd.n7304 gnd.n7303 9.3005
R11035 gnd.n7305 gnd.n467 9.3005
R11036 gnd.n7307 gnd.n7306 9.3005
R11037 gnd.n463 gnd.n462 9.3005
R11038 gnd.n7314 gnd.n7313 9.3005
R11039 gnd.n7315 gnd.n461 9.3005
R11040 gnd.n7317 gnd.n7316 9.3005
R11041 gnd.n457 gnd.n456 9.3005
R11042 gnd.n7324 gnd.n7323 9.3005
R11043 gnd.n7325 gnd.n455 9.3005
R11044 gnd.n7327 gnd.n7326 9.3005
R11045 gnd.n451 gnd.n450 9.3005
R11046 gnd.n7334 gnd.n7333 9.3005
R11047 gnd.n7335 gnd.n449 9.3005
R11048 gnd.n7337 gnd.n7336 9.3005
R11049 gnd.n445 gnd.n444 9.3005
R11050 gnd.n7344 gnd.n7343 9.3005
R11051 gnd.n7345 gnd.n443 9.3005
R11052 gnd.n7347 gnd.n7346 9.3005
R11053 gnd.n439 gnd.n438 9.3005
R11054 gnd.n7354 gnd.n7353 9.3005
R11055 gnd.n7355 gnd.n437 9.3005
R11056 gnd.n7357 gnd.n7356 9.3005
R11057 gnd.n433 gnd.n432 9.3005
R11058 gnd.n7364 gnd.n7363 9.3005
R11059 gnd.n7365 gnd.n431 9.3005
R11060 gnd.n7367 gnd.n7366 9.3005
R11061 gnd.n427 gnd.n426 9.3005
R11062 gnd.n7374 gnd.n7373 9.3005
R11063 gnd.n7375 gnd.n425 9.3005
R11064 gnd.n7377 gnd.n7376 9.3005
R11065 gnd.n421 gnd.n420 9.3005
R11066 gnd.n7384 gnd.n7383 9.3005
R11067 gnd.n7385 gnd.n419 9.3005
R11068 gnd.n7387 gnd.n7386 9.3005
R11069 gnd.n415 gnd.n414 9.3005
R11070 gnd.n7394 gnd.n7393 9.3005
R11071 gnd.n7395 gnd.n413 9.3005
R11072 gnd.n7397 gnd.n7396 9.3005
R11073 gnd.n409 gnd.n408 9.3005
R11074 gnd.n7404 gnd.n7403 9.3005
R11075 gnd.n7405 gnd.n407 9.3005
R11076 gnd.n7409 gnd.n7406 9.3005
R11077 gnd.n7408 gnd.n7407 9.3005
R11078 gnd.n403 gnd.n402 9.3005
R11079 gnd.n7417 gnd.n7416 9.3005
R11080 gnd.n7205 gnd.n527 9.3005
R11081 gnd.n7753 gnd.n7752 9.3005
R11082 gnd.n7751 gnd.n80 9.3005
R11083 gnd.n7442 gnd.n83 9.3005
R11084 gnd.n7444 gnd.n7443 9.3005
R11085 gnd.n377 gnd.n376 9.3005
R11086 gnd.n7455 gnd.n7454 9.3005
R11087 gnd.n7456 gnd.n375 9.3005
R11088 gnd.n7458 gnd.n7457 9.3005
R11089 gnd.n370 gnd.n369 9.3005
R11090 gnd.n7469 gnd.n7468 9.3005
R11091 gnd.n7470 gnd.n368 9.3005
R11092 gnd.n7472 gnd.n7471 9.3005
R11093 gnd.n365 gnd.n364 9.3005
R11094 gnd.n7483 gnd.n7482 9.3005
R11095 gnd.n7484 gnd.n363 9.3005
R11096 gnd.n7487 gnd.n7486 9.3005
R11097 gnd.n7485 gnd.n359 9.3005
R11098 gnd.n7512 gnd.n358 9.3005
R11099 gnd.n7514 gnd.n7513 9.3005
R11100 gnd.n7515 gnd.n357 9.3005
R11101 gnd.n7517 gnd.n7516 9.3005
R11102 gnd.n7519 gnd.n355 9.3005
R11103 gnd.n7521 gnd.n7520 9.3005
R11104 gnd.n7522 gnd.n354 9.3005
R11105 gnd.n7524 gnd.n7523 9.3005
R11106 gnd.n7526 gnd.n352 9.3005
R11107 gnd.n7528 gnd.n7527 9.3005
R11108 gnd.n7559 gnd.n318 9.3005
R11109 gnd.n7558 gnd.n320 9.3005
R11110 gnd.n324 gnd.n321 9.3005
R11111 gnd.n7553 gnd.n325 9.3005
R11112 gnd.n7552 gnd.n326 9.3005
R11113 gnd.n7551 gnd.n327 9.3005
R11114 gnd.n331 gnd.n328 9.3005
R11115 gnd.n7546 gnd.n332 9.3005
R11116 gnd.n7545 gnd.n333 9.3005
R11117 gnd.n7544 gnd.n334 9.3005
R11118 gnd.n338 gnd.n335 9.3005
R11119 gnd.n7539 gnd.n339 9.3005
R11120 gnd.n7538 gnd.n340 9.3005
R11121 gnd.n7537 gnd.n341 9.3005
R11122 gnd.n345 gnd.n342 9.3005
R11123 gnd.n7532 gnd.n346 9.3005
R11124 gnd.n7531 gnd.n7530 9.3005
R11125 gnd.n7529 gnd.n349 9.3005
R11126 gnd.n7561 gnd.n7560 9.3005
R11127 gnd.n7669 gnd.n215 9.3005
R11128 gnd.n7668 gnd.n217 9.3005
R11129 gnd.n221 gnd.n218 9.3005
R11130 gnd.n7663 gnd.n222 9.3005
R11131 gnd.n7662 gnd.n223 9.3005
R11132 gnd.n7661 gnd.n224 9.3005
R11133 gnd.n228 gnd.n225 9.3005
R11134 gnd.n7656 gnd.n229 9.3005
R11135 gnd.n7655 gnd.n230 9.3005
R11136 gnd.n7654 gnd.n231 9.3005
R11137 gnd.n235 gnd.n232 9.3005
R11138 gnd.n7649 gnd.n236 9.3005
R11139 gnd.n7648 gnd.n237 9.3005
R11140 gnd.n7647 gnd.n238 9.3005
R11141 gnd.n242 gnd.n239 9.3005
R11142 gnd.n7642 gnd.n243 9.3005
R11143 gnd.n7641 gnd.n244 9.3005
R11144 gnd.n7637 gnd.n245 9.3005
R11145 gnd.n249 gnd.n246 9.3005
R11146 gnd.n7632 gnd.n250 9.3005
R11147 gnd.n7631 gnd.n251 9.3005
R11148 gnd.n7630 gnd.n252 9.3005
R11149 gnd.n256 gnd.n253 9.3005
R11150 gnd.n7625 gnd.n257 9.3005
R11151 gnd.n7624 gnd.n258 9.3005
R11152 gnd.n7623 gnd.n259 9.3005
R11153 gnd.n263 gnd.n260 9.3005
R11154 gnd.n7618 gnd.n264 9.3005
R11155 gnd.n7617 gnd.n265 9.3005
R11156 gnd.n7616 gnd.n266 9.3005
R11157 gnd.n270 gnd.n267 9.3005
R11158 gnd.n7611 gnd.n271 9.3005
R11159 gnd.n7610 gnd.n272 9.3005
R11160 gnd.n7609 gnd.n273 9.3005
R11161 gnd.n277 gnd.n274 9.3005
R11162 gnd.n7604 gnd.n278 9.3005
R11163 gnd.n7603 gnd.n7602 9.3005
R11164 gnd.n7601 gnd.n279 9.3005
R11165 gnd.n7600 gnd.n7599 9.3005
R11166 gnd.n283 gnd.n282 9.3005
R11167 gnd.n288 gnd.n286 9.3005
R11168 gnd.n7592 gnd.n289 9.3005
R11169 gnd.n7591 gnd.n290 9.3005
R11170 gnd.n7590 gnd.n291 9.3005
R11171 gnd.n295 gnd.n292 9.3005
R11172 gnd.n7585 gnd.n296 9.3005
R11173 gnd.n7584 gnd.n297 9.3005
R11174 gnd.n7583 gnd.n298 9.3005
R11175 gnd.n302 gnd.n299 9.3005
R11176 gnd.n7578 gnd.n303 9.3005
R11177 gnd.n7577 gnd.n304 9.3005
R11178 gnd.n7576 gnd.n305 9.3005
R11179 gnd.n309 gnd.n306 9.3005
R11180 gnd.n7571 gnd.n310 9.3005
R11181 gnd.n7570 gnd.n311 9.3005
R11182 gnd.n7569 gnd.n312 9.3005
R11183 gnd.n317 gnd.n315 9.3005
R11184 gnd.n7564 gnd.n7563 9.3005
R11185 gnd.n7671 gnd.n7670 9.3005
R11186 gnd.n4429 gnd.n1636 9.3005
R11187 gnd.n4639 gnd.n1637 9.3005
R11188 gnd.n4638 gnd.n1638 9.3005
R11189 gnd.n4637 gnd.n1639 9.3005
R11190 gnd.n1821 gnd.n1640 9.3005
R11191 gnd.n4627 gnd.n1657 9.3005
R11192 gnd.n4626 gnd.n1658 9.3005
R11193 gnd.n4625 gnd.n1659 9.3005
R11194 gnd.n1784 gnd.n1660 9.3005
R11195 gnd.n4615 gnd.n1678 9.3005
R11196 gnd.n4614 gnd.n1679 9.3005
R11197 gnd.n4613 gnd.n1680 9.3005
R11198 gnd.n4462 gnd.n1681 9.3005
R11199 gnd.n4603 gnd.n1697 9.3005
R11200 gnd.n4602 gnd.n1698 9.3005
R11201 gnd.n4601 gnd.n1699 9.3005
R11202 gnd.n4472 gnd.n1700 9.3005
R11203 gnd.n4591 gnd.n1718 9.3005
R11204 gnd.n4590 gnd.n1719 9.3005
R11205 gnd.n4589 gnd.n1720 9.3005
R11206 gnd.n4520 gnd.n1721 9.3005
R11207 gnd.n4579 gnd.n1735 9.3005
R11208 gnd.n4578 gnd.n1736 9.3005
R11209 gnd.n4577 gnd.n1737 9.3005
R11210 gnd.n4521 gnd.n1738 9.3005
R11211 gnd.n4526 gnd.n4522 9.3005
R11212 gnd.n4534 gnd.n4527 9.3005
R11213 gnd.n4533 gnd.n4529 9.3005
R11214 gnd.n4532 gnd.n4530 9.3005
R11215 gnd.n379 gnd.n108 9.3005
R11216 gnd.n7739 gnd.n109 9.3005
R11217 gnd.n7738 gnd.n110 9.3005
R11218 gnd.n7737 gnd.n111 9.3005
R11219 gnd.n373 gnd.n112 9.3005
R11220 gnd.n7727 gnd.n127 9.3005
R11221 gnd.n7726 gnd.n128 9.3005
R11222 gnd.n7725 gnd.n129 9.3005
R11223 gnd.n367 gnd.n130 9.3005
R11224 gnd.n7715 gnd.n148 9.3005
R11225 gnd.n7714 gnd.n149 9.3005
R11226 gnd.n7713 gnd.n150 9.3005
R11227 gnd.n361 gnd.n151 9.3005
R11228 gnd.n7703 gnd.n167 9.3005
R11229 gnd.n7702 gnd.n168 9.3005
R11230 gnd.n7701 gnd.n169 9.3005
R11231 gnd.n7493 gnd.n170 9.3005
R11232 gnd.n7691 gnd.n187 9.3005
R11233 gnd.n7690 gnd.n188 9.3005
R11234 gnd.n7689 gnd.n189 9.3005
R11235 gnd.n7494 gnd.n190 9.3005
R11236 gnd.n7679 gnd.n205 9.3005
R11237 gnd.n7678 gnd.n206 9.3005
R11238 gnd.n7677 gnd.n207 9.3005
R11239 gnd.n4428 gnd.n4427 9.3005
R11240 gnd.n4430 gnd.n4429 9.3005
R11241 gnd.n4431 gnd.n1637 9.3005
R11242 gnd.n4432 gnd.n1638 9.3005
R11243 gnd.n1820 gnd.n1639 9.3005
R11244 gnd.n4444 gnd.n1821 9.3005
R11245 gnd.n4445 gnd.n1657 9.3005
R11246 gnd.n4446 gnd.n1658 9.3005
R11247 gnd.n1783 gnd.n1659 9.3005
R11248 gnd.n4458 gnd.n1784 9.3005
R11249 gnd.n4459 gnd.n1678 9.3005
R11250 gnd.n4460 gnd.n1679 9.3005
R11251 gnd.n4461 gnd.n1680 9.3005
R11252 gnd.n4465 gnd.n4462 9.3005
R11253 gnd.n4466 gnd.n1697 9.3005
R11254 gnd.n4470 gnd.n1698 9.3005
R11255 gnd.n4471 gnd.n1699 9.3005
R11256 gnd.n4473 gnd.n4472 9.3005
R11257 gnd.n1761 gnd.n1718 9.3005
R11258 gnd.n4518 gnd.n1719 9.3005
R11259 gnd.n4519 gnd.n1720 9.3005
R11260 gnd.n4544 gnd.n4520 9.3005
R11261 gnd.n4543 gnd.n1735 9.3005
R11262 gnd.n4542 gnd.n1736 9.3005
R11263 gnd.n4541 gnd.n1737 9.3005
R11264 gnd.n4540 gnd.n4521 9.3005
R11265 gnd.n4539 gnd.n4522 9.3005
R11266 gnd.n4527 gnd.n4523 9.3005
R11267 gnd.n4529 gnd.n4528 9.3005
R11268 gnd.n4530 gnd.n378 9.3005
R11269 gnd.n7448 gnd.n379 9.3005
R11270 gnd.n7449 gnd.n109 9.3005
R11271 gnd.n7450 gnd.n110 9.3005
R11272 gnd.n372 gnd.n111 9.3005
R11273 gnd.n7462 gnd.n373 9.3005
R11274 gnd.n7463 gnd.n127 9.3005
R11275 gnd.n7464 gnd.n128 9.3005
R11276 gnd.n366 gnd.n129 9.3005
R11277 gnd.n7476 gnd.n367 9.3005
R11278 gnd.n7477 gnd.n148 9.3005
R11279 gnd.n7478 gnd.n149 9.3005
R11280 gnd.n360 gnd.n150 9.3005
R11281 gnd.n7491 gnd.n361 9.3005
R11282 gnd.n7492 gnd.n167 9.3005
R11283 gnd.n7508 gnd.n168 9.3005
R11284 gnd.n7507 gnd.n169 9.3005
R11285 gnd.n7506 gnd.n7493 9.3005
R11286 gnd.n7504 gnd.n187 9.3005
R11287 gnd.n7503 gnd.n188 9.3005
R11288 gnd.n7501 gnd.n189 9.3005
R11289 gnd.n7500 gnd.n7494 9.3005
R11290 gnd.n7498 gnd.n205 9.3005
R11291 gnd.n7497 gnd.n206 9.3005
R11292 gnd.n7495 gnd.n207 9.3005
R11293 gnd.n4428 gnd.n1825 9.3005
R11294 gnd.n1831 gnd.n1828 9.3005
R11295 gnd.n4415 gnd.n1832 9.3005
R11296 gnd.n4417 gnd.n4416 9.3005
R11297 gnd.n4414 gnd.n1834 9.3005
R11298 gnd.n4413 gnd.n4412 9.3005
R11299 gnd.n1836 gnd.n1835 9.3005
R11300 gnd.n4406 gnd.n4405 9.3005
R11301 gnd.n4404 gnd.n1838 9.3005
R11302 gnd.n4403 gnd.n4402 9.3005
R11303 gnd.n1840 gnd.n1839 9.3005
R11304 gnd.n4396 gnd.n4395 9.3005
R11305 gnd.n4394 gnd.n1842 9.3005
R11306 gnd.n4393 gnd.n4392 9.3005
R11307 gnd.n1844 gnd.n1843 9.3005
R11308 gnd.n4386 gnd.n4385 9.3005
R11309 gnd.n4384 gnd.n1846 9.3005
R11310 gnd.n4383 gnd.n4382 9.3005
R11311 gnd.n1848 gnd.n1847 9.3005
R11312 gnd.n4376 gnd.n4375 9.3005
R11313 gnd.n4374 gnd.n1850 9.3005
R11314 gnd.n1852 gnd.n1851 9.3005
R11315 gnd.n4364 gnd.n4363 9.3005
R11316 gnd.n4362 gnd.n1854 9.3005
R11317 gnd.n4361 gnd.n4360 9.3005
R11318 gnd.n1856 gnd.n1855 9.3005
R11319 gnd.n4354 gnd.n4353 9.3005
R11320 gnd.n4352 gnd.n1858 9.3005
R11321 gnd.n4351 gnd.n4350 9.3005
R11322 gnd.n1860 gnd.n1859 9.3005
R11323 gnd.n4342 gnd.n4341 9.3005
R11324 gnd.n4339 gnd.n4252 9.3005
R11325 gnd.n4338 gnd.n4337 9.3005
R11326 gnd.n4254 gnd.n4253 9.3005
R11327 gnd.n4331 gnd.n4330 9.3005
R11328 gnd.n4329 gnd.n4256 9.3005
R11329 gnd.n4328 gnd.n4327 9.3005
R11330 gnd.n4258 gnd.n4257 9.3005
R11331 gnd.n4321 gnd.n4317 9.3005
R11332 gnd.n4316 gnd.n4260 9.3005
R11333 gnd.n4315 gnd.n4314 9.3005
R11334 gnd.n4262 gnd.n4261 9.3005
R11335 gnd.n4308 gnd.n4307 9.3005
R11336 gnd.n4306 gnd.n4264 9.3005
R11337 gnd.n4305 gnd.n4304 9.3005
R11338 gnd.n4266 gnd.n4265 9.3005
R11339 gnd.n4298 gnd.n4297 9.3005
R11340 gnd.n4296 gnd.n4268 9.3005
R11341 gnd.n4295 gnd.n4294 9.3005
R11342 gnd.n4270 gnd.n4269 9.3005
R11343 gnd.n4288 gnd.n4287 9.3005
R11344 gnd.n4286 gnd.n4272 9.3005
R11345 gnd.n4285 gnd.n4284 9.3005
R11346 gnd.n4274 gnd.n4273 9.3005
R11347 gnd.n4278 gnd.n4277 9.3005
R11348 gnd.n4276 gnd.n4275 9.3005
R11349 gnd.n4373 gnd.n4372 9.3005
R11350 gnd.n4425 gnd.n4424 9.3005
R11351 gnd.n4644 gnd.n1626 9.3005
R11352 gnd.n4643 gnd.n1627 9.3005
R11353 gnd.n1647 gnd.n1628 9.3005
R11354 gnd.n4633 gnd.n1648 9.3005
R11355 gnd.n4632 gnd.n1649 9.3005
R11356 gnd.n4631 gnd.n1650 9.3005
R11357 gnd.n1667 gnd.n1651 9.3005
R11358 gnd.n4621 gnd.n1668 9.3005
R11359 gnd.n4620 gnd.n1669 9.3005
R11360 gnd.n4619 gnd.n1670 9.3005
R11361 gnd.n1687 gnd.n1671 9.3005
R11362 gnd.n4609 gnd.n1688 9.3005
R11363 gnd.n4608 gnd.n1689 9.3005
R11364 gnd.n4607 gnd.n1690 9.3005
R11365 gnd.n1707 gnd.n1691 9.3005
R11366 gnd.n4597 gnd.n1708 9.3005
R11367 gnd.n4596 gnd.n1709 9.3005
R11368 gnd.n4595 gnd.n1710 9.3005
R11369 gnd.n1727 gnd.n1711 9.3005
R11370 gnd.n4585 gnd.n1728 9.3005
R11371 gnd.n4584 gnd.n94 9.3005
R11372 gnd.n99 gnd.n93 9.3005
R11373 gnd.n7733 gnd.n118 9.3005
R11374 gnd.n7732 gnd.n119 9.3005
R11375 gnd.n7731 gnd.n120 9.3005
R11376 gnd.n137 gnd.n121 9.3005
R11377 gnd.n7721 gnd.n138 9.3005
R11378 gnd.n7720 gnd.n139 9.3005
R11379 gnd.n7719 gnd.n140 9.3005
R11380 gnd.n157 gnd.n141 9.3005
R11381 gnd.n7709 gnd.n158 9.3005
R11382 gnd.n7708 gnd.n159 9.3005
R11383 gnd.n7707 gnd.n160 9.3005
R11384 gnd.n177 gnd.n161 9.3005
R11385 gnd.n7697 gnd.n178 9.3005
R11386 gnd.n7696 gnd.n179 9.3005
R11387 gnd.n7695 gnd.n180 9.3005
R11388 gnd.n196 gnd.n181 9.3005
R11389 gnd.n7685 gnd.n197 9.3005
R11390 gnd.n7684 gnd.n198 9.3005
R11391 gnd.n7683 gnd.n199 9.3005
R11392 gnd.n214 gnd.n200 9.3005
R11393 gnd.n7673 gnd.n7672 9.3005
R11394 gnd.n4645 gnd.n1625 9.3005
R11395 gnd.n7744 gnd.n97 9.3005
R11396 gnd.n7744 gnd.n7743 9.3005
R11397 gnd.n2808 gnd.n2807 9.3005
R11398 gnd.n2809 gnd.n2455 9.3005
R11399 gnd.n2811 gnd.n2810 9.3005
R11400 gnd.n2453 gnd.n2452 9.3005
R11401 gnd.n2816 gnd.n2815 9.3005
R11402 gnd.n2817 gnd.n2451 9.3005
R11403 gnd.n2838 gnd.n2818 9.3005
R11404 gnd.n2837 gnd.n2819 9.3005
R11405 gnd.n2836 gnd.n2820 9.3005
R11406 gnd.n2823 gnd.n2821 9.3005
R11407 gnd.n2832 gnd.n2824 9.3005
R11408 gnd.n2831 gnd.n2825 9.3005
R11409 gnd.n2830 gnd.n2826 9.3005
R11410 gnd.n2828 gnd.n2827 9.3005
R11411 gnd.n2428 gnd.n2427 9.3005
R11412 gnd.n2903 gnd.n2902 9.3005
R11413 gnd.n2904 gnd.n2426 9.3005
R11414 gnd.n2906 gnd.n2905 9.3005
R11415 gnd.n2424 gnd.n2423 9.3005
R11416 gnd.n2911 gnd.n2910 9.3005
R11417 gnd.n2912 gnd.n2422 9.3005
R11418 gnd.n2914 gnd.n2913 9.3005
R11419 gnd.n2420 gnd.n2419 9.3005
R11420 gnd.n2921 gnd.n2920 9.3005
R11421 gnd.n2922 gnd.n2418 9.3005
R11422 gnd.n2924 gnd.n2923 9.3005
R11423 gnd.n2395 gnd.n2394 9.3005
R11424 gnd.n3205 gnd.n3204 9.3005
R11425 gnd.n3206 gnd.n2393 9.3005
R11426 gnd.n3210 gnd.n3207 9.3005
R11427 gnd.n3209 gnd.n3208 9.3005
R11428 gnd.n2370 gnd.n2369 9.3005
R11429 gnd.n3237 gnd.n3236 9.3005
R11430 gnd.n3238 gnd.n2368 9.3005
R11431 gnd.n3243 gnd.n3239 9.3005
R11432 gnd.n3242 gnd.n3241 9.3005
R11433 gnd.n3240 gnd.n1496 9.3005
R11434 gnd.n4778 gnd.n1497 9.3005
R11435 gnd.n4777 gnd.n1498 9.3005
R11436 gnd.n4776 gnd.n1499 9.3005
R11437 gnd.n3277 gnd.n1500 9.3005
R11438 gnd.n3279 gnd.n3278 9.3005
R11439 gnd.n2244 gnd.n2243 9.3005
R11440 gnd.n3319 gnd.n3318 9.3005
R11441 gnd.n3320 gnd.n2242 9.3005
R11442 gnd.n3322 gnd.n3321 9.3005
R11443 gnd.n2226 gnd.n2225 9.3005
R11444 gnd.n3361 gnd.n3360 9.3005
R11445 gnd.n3362 gnd.n2224 9.3005
R11446 gnd.n3366 gnd.n3363 9.3005
R11447 gnd.n3365 gnd.n3364 9.3005
R11448 gnd.n2200 gnd.n2199 9.3005
R11449 gnd.n3423 gnd.n3422 9.3005
R11450 gnd.n3424 gnd.n2198 9.3005
R11451 gnd.n3426 gnd.n3425 9.3005
R11452 gnd.n2182 gnd.n2181 9.3005
R11453 gnd.n3451 gnd.n3450 9.3005
R11454 gnd.n3452 gnd.n2180 9.3005
R11455 gnd.n3456 gnd.n3453 9.3005
R11456 gnd.n3455 gnd.n3454 9.3005
R11457 gnd.n2149 gnd.n2148 9.3005
R11458 gnd.n3501 gnd.n3500 9.3005
R11459 gnd.n3502 gnd.n2147 9.3005
R11460 gnd.n3504 gnd.n3503 9.3005
R11461 gnd.n2126 gnd.n2125 9.3005
R11462 gnd.n3541 gnd.n3540 9.3005
R11463 gnd.n3542 gnd.n2124 9.3005
R11464 gnd.n3544 gnd.n3543 9.3005
R11465 gnd.n2104 gnd.n2103 9.3005
R11466 gnd.n3598 gnd.n3597 9.3005
R11467 gnd.n3599 gnd.n2102 9.3005
R11468 gnd.n3601 gnd.n3600 9.3005
R11469 gnd.n2084 gnd.n2083 9.3005
R11470 gnd.n3623 gnd.n3622 9.3005
R11471 gnd.n3624 gnd.n2082 9.3005
R11472 gnd.n3626 gnd.n3625 9.3005
R11473 gnd.n2064 gnd.n2063 9.3005
R11474 gnd.n3683 gnd.n3682 9.3005
R11475 gnd.n3684 gnd.n2062 9.3005
R11476 gnd.n3686 gnd.n3685 9.3005
R11477 gnd.n2042 gnd.n2041 9.3005
R11478 gnd.n3712 gnd.n3711 9.3005
R11479 gnd.n3713 gnd.n2040 9.3005
R11480 gnd.n3717 gnd.n3714 9.3005
R11481 gnd.n3716 gnd.n3715 9.3005
R11482 gnd.n2014 gnd.n2013 9.3005
R11483 gnd.n3763 gnd.n3762 9.3005
R11484 gnd.n3764 gnd.n2012 9.3005
R11485 gnd.n3766 gnd.n3765 9.3005
R11486 gnd.n1994 gnd.n1993 9.3005
R11487 gnd.n3789 gnd.n3788 9.3005
R11488 gnd.n3790 gnd.n1992 9.3005
R11489 gnd.n3794 gnd.n3791 9.3005
R11490 gnd.n3793 gnd.n3792 9.3005
R11491 gnd.n1964 gnd.n1963 9.3005
R11492 gnd.n3833 gnd.n3832 9.3005
R11493 gnd.n3834 gnd.n1962 9.3005
R11494 gnd.n3839 gnd.n3835 9.3005
R11495 gnd.n3838 gnd.n3837 9.3005
R11496 gnd.n3836 gnd.n1913 9.3005
R11497 gnd.n4085 gnd.n1914 9.3005
R11498 gnd.n4084 gnd.n1915 9.3005
R11499 gnd.n4083 gnd.n1916 9.3005
R11500 gnd.n1925 gnd.n1917 9.3005
R11501 gnd.n1926 gnd.n1924 9.3005
R11502 gnd.n4073 gnd.n1927 9.3005
R11503 gnd.n4072 gnd.n1928 9.3005
R11504 gnd.n4071 gnd.n1929 9.3005
R11505 gnd.n1932 gnd.n1931 9.3005
R11506 gnd.n1930 gnd.n1603 9.3005
R11507 gnd.n4660 gnd.n1604 9.3005
R11508 gnd.n4659 gnd.n1605 9.3005
R11509 gnd.n4658 gnd.n1606 9.3005
R11510 gnd.n1612 gnd.n1607 9.3005
R11511 gnd.n4652 gnd.n1613 9.3005
R11512 gnd.n4651 gnd.n1614 9.3005
R11513 gnd.n4650 gnd.n1615 9.3005
R11514 gnd.n1795 gnd.n1616 9.3005
R11515 gnd.n1796 gnd.n1794 9.3005
R11516 gnd.n1798 gnd.n1797 9.3005
R11517 gnd.n1792 gnd.n1791 9.3005
R11518 gnd.n1803 gnd.n1802 9.3005
R11519 gnd.n1804 gnd.n1790 9.3005
R11520 gnd.n1817 gnd.n1805 9.3005
R11521 gnd.n1816 gnd.n1806 9.3005
R11522 gnd.n1815 gnd.n1807 9.3005
R11523 gnd.n1812 gnd.n1808 9.3005
R11524 gnd.n1811 gnd.n1810 9.3005
R11525 gnd.n1809 gnd.n1773 9.3005
R11526 gnd.n1771 gnd.n1770 9.3005
R11527 gnd.n4498 gnd.n4497 9.3005
R11528 gnd.n4499 gnd.n1769 9.3005
R11529 gnd.n4501 gnd.n4500 9.3005
R11530 gnd.n1767 gnd.n1766 9.3005
R11531 gnd.n4506 gnd.n4505 9.3005
R11532 gnd.n4507 gnd.n1765 9.3005
R11533 gnd.n4513 gnd.n4508 9.3005
R11534 gnd.n4512 gnd.n4509 9.3005
R11535 gnd.n7436 gnd.n385 9.3005
R11536 gnd.n388 gnd.n386 9.3005
R11537 gnd.n7432 gnd.n389 9.3005
R11538 gnd.n7431 gnd.n390 9.3005
R11539 gnd.n7430 gnd.n391 9.3005
R11540 gnd.n394 gnd.n392 9.3005
R11541 gnd.n7426 gnd.n395 9.3005
R11542 gnd.n7425 gnd.n396 9.3005
R11543 gnd.n7424 gnd.n397 9.3005
R11544 gnd.n400 gnd.n398 9.3005
R11545 gnd.n7420 gnd.n401 9.3005
R11546 gnd.n7419 gnd.n7418 9.3005
R11547 gnd.n2609 gnd.n2547 9.3005
R11548 gnd.n2612 gnd.n2610 9.3005
R11549 gnd.n2613 gnd.n2546 9.3005
R11550 gnd.n2616 gnd.n2615 9.3005
R11551 gnd.n2617 gnd.n2545 9.3005
R11552 gnd.n2620 gnd.n2618 9.3005
R11553 gnd.n2621 gnd.n2544 9.3005
R11554 gnd.n2624 gnd.n2623 9.3005
R11555 gnd.n2625 gnd.n2543 9.3005
R11556 gnd.n2627 gnd.n2626 9.3005
R11557 gnd.n2528 gnd.n2527 9.3005
R11558 gnd.n2638 gnd.n2637 9.3005
R11559 gnd.n2639 gnd.n2526 9.3005
R11560 gnd.n2641 gnd.n2640 9.3005
R11561 gnd.n2523 gnd.n2522 9.3005
R11562 gnd.n2691 gnd.n2690 9.3005
R11563 gnd.n2692 gnd.n2521 9.3005
R11564 gnd.n2695 gnd.n2694 9.3005
R11565 gnd.n2693 gnd.n2517 9.3005
R11566 gnd.n2706 gnd.n2518 9.3005
R11567 gnd.n2707 gnd.n2516 9.3005
R11568 gnd.n2710 gnd.n2709 9.3005
R11569 gnd.n2711 gnd.n2515 9.3005
R11570 gnd.n2713 gnd.n2712 9.3005
R11571 gnd.n2481 gnd.n2480 9.3005
R11572 gnd.n2755 gnd.n2754 9.3005
R11573 gnd.n2608 gnd.n2607 9.3005
R11574 gnd.n2602 gnd.n2601 9.3005
R11575 gnd.n2600 gnd.n2552 9.3005
R11576 gnd.n2599 gnd.n2598 9.3005
R11577 gnd.n2595 gnd.n2555 9.3005
R11578 gnd.n2594 gnd.n2591 9.3005
R11579 gnd.n2590 gnd.n2556 9.3005
R11580 gnd.n2589 gnd.n2588 9.3005
R11581 gnd.n2585 gnd.n2557 9.3005
R11582 gnd.n2584 gnd.n2581 9.3005
R11583 gnd.n2580 gnd.n2558 9.3005
R11584 gnd.n2579 gnd.n2578 9.3005
R11585 gnd.n2575 gnd.n2559 9.3005
R11586 gnd.n2574 gnd.n2571 9.3005
R11587 gnd.n2570 gnd.n2560 9.3005
R11588 gnd.n2569 gnd.n2568 9.3005
R11589 gnd.n2565 gnd.n2561 9.3005
R11590 gnd.n2564 gnd.n1136 9.3005
R11591 gnd.n2603 gnd.n2548 9.3005
R11592 gnd.n2605 gnd.n2604 9.3005
R11593 gnd.n4856 gnd.n1424 9.3005
R11594 gnd.n4857 gnd.n1423 9.3005
R11595 gnd.n1422 gnd.n1419 9.3005
R11596 gnd.n4862 gnd.n1418 9.3005
R11597 gnd.n4863 gnd.n1417 9.3005
R11598 gnd.n4864 gnd.n1416 9.3005
R11599 gnd.n1415 gnd.n1412 9.3005
R11600 gnd.n4869 gnd.n1411 9.3005
R11601 gnd.n4871 gnd.n1408 9.3005
R11602 gnd.n4872 gnd.n1407 9.3005
R11603 gnd.n1406 gnd.n1403 9.3005
R11604 gnd.n4877 gnd.n1402 9.3005
R11605 gnd.n4878 gnd.n1401 9.3005
R11606 gnd.n4879 gnd.n1400 9.3005
R11607 gnd.n1399 gnd.n1396 9.3005
R11608 gnd.n4884 gnd.n1395 9.3005
R11609 gnd.n4885 gnd.n1394 9.3005
R11610 gnd.n4886 gnd.n1393 9.3005
R11611 gnd.n1392 gnd.n1389 9.3005
R11612 gnd.n4891 gnd.n1388 9.3005
R11613 gnd.n4892 gnd.n1387 9.3005
R11614 gnd.n4893 gnd.n1386 9.3005
R11615 gnd.n1385 gnd.n1382 9.3005
R11616 gnd.n1384 gnd.n1380 9.3005
R11617 gnd.n4900 gnd.n1379 9.3005
R11618 gnd.n4902 gnd.n4901 9.3005
R11619 gnd.n2982 gnd.n2981 9.3005
R11620 gnd.n2990 gnd.n2989 9.3005
R11621 gnd.n2991 gnd.n2979 9.3005
R11622 gnd.n2993 gnd.n2992 9.3005
R11623 gnd.n2977 gnd.n2976 9.3005
R11624 gnd.n3000 gnd.n2999 9.3005
R11625 gnd.n3001 gnd.n2975 9.3005
R11626 gnd.n3003 gnd.n3002 9.3005
R11627 gnd.n2973 gnd.n2970 9.3005
R11628 gnd.n3010 gnd.n3009 9.3005
R11629 gnd.n3011 gnd.n2969 9.3005
R11630 gnd.n3013 gnd.n3012 9.3005
R11631 gnd.n2967 gnd.n2966 9.3005
R11632 gnd.n3020 gnd.n3019 9.3005
R11633 gnd.n3021 gnd.n2965 9.3005
R11634 gnd.n3023 gnd.n3022 9.3005
R11635 gnd.n2963 gnd.n2962 9.3005
R11636 gnd.n3030 gnd.n3029 9.3005
R11637 gnd.n3031 gnd.n2961 9.3005
R11638 gnd.n3033 gnd.n3032 9.3005
R11639 gnd.n2959 gnd.n2958 9.3005
R11640 gnd.n3040 gnd.n3039 9.3005
R11641 gnd.n3041 gnd.n2957 9.3005
R11642 gnd.n3043 gnd.n3042 9.3005
R11643 gnd.n2955 gnd.n2954 9.3005
R11644 gnd.n3050 gnd.n3049 9.3005
R11645 gnd.n3051 gnd.n2953 9.3005
R11646 gnd.n3053 gnd.n3052 9.3005
R11647 gnd.n2951 gnd.n2948 9.3005
R11648 gnd.n3059 gnd.n3058 9.3005
R11649 gnd.n2980 gnd.n1425 9.3005
R11650 gnd.n1158 gnd.n1138 9.3005
R11651 gnd.n2529 gnd.n1159 9.3005
R11652 gnd.n5032 gnd.n1160 9.3005
R11653 gnd.n5031 gnd.n1161 9.3005
R11654 gnd.n5030 gnd.n1162 9.3005
R11655 gnd.n2535 gnd.n1163 9.3005
R11656 gnd.n5020 gnd.n1179 9.3005
R11657 gnd.n5019 gnd.n1180 9.3005
R11658 gnd.n5018 gnd.n1181 9.3005
R11659 gnd.n2542 gnd.n1182 9.3005
R11660 gnd.n5008 gnd.n1199 9.3005
R11661 gnd.n5007 gnd.n1200 9.3005
R11662 gnd.n5006 gnd.n1201 9.3005
R11663 gnd.n2525 gnd.n1202 9.3005
R11664 gnd.n4996 gnd.n1219 9.3005
R11665 gnd.n4995 gnd.n1220 9.3005
R11666 gnd.n4994 gnd.n1221 9.3005
R11667 gnd.n2520 gnd.n1222 9.3005
R11668 gnd.n4984 gnd.n1240 9.3005
R11669 gnd.n4983 gnd.n1241 9.3005
R11670 gnd.n4982 gnd.n1242 9.3005
R11671 gnd.n2507 gnd.n1243 9.3005
R11672 gnd.n2720 gnd.n2719 9.3005
R11673 gnd.n2508 gnd.n2492 9.3005
R11674 gnd.n2745 gnd.n2493 9.3005
R11675 gnd.n2744 gnd.n2494 9.3005
R11676 gnd.n2743 gnd.n2495 9.3005
R11677 gnd.n2472 gnd.n2471 9.3005
R11678 gnd.n2769 gnd.n2768 9.3005
R11679 gnd.n2770 gnd.n1268 9.3005
R11680 gnd.n4970 gnd.n1269 9.3005
R11681 gnd.n4969 gnd.n1270 9.3005
R11682 gnd.n4968 gnd.n1271 9.3005
R11683 gnd.n2777 gnd.n1272 9.3005
R11684 gnd.n4958 gnd.n1288 9.3005
R11685 gnd.n4957 gnd.n1289 9.3005
R11686 gnd.n4956 gnd.n1290 9.3005
R11687 gnd.n2783 gnd.n1291 9.3005
R11688 gnd.n4946 gnd.n1308 9.3005
R11689 gnd.n4945 gnd.n1309 9.3005
R11690 gnd.n4944 gnd.n1310 9.3005
R11691 gnd.n2853 gnd.n1311 9.3005
R11692 gnd.n4934 gnd.n1328 9.3005
R11693 gnd.n4933 gnd.n1329 9.3005
R11694 gnd.n4932 gnd.n1330 9.3005
R11695 gnd.n2868 gnd.n1331 9.3005
R11696 gnd.n4922 gnd.n1348 9.3005
R11697 gnd.n4921 gnd.n1349 9.3005
R11698 gnd.n4920 gnd.n1350 9.3005
R11699 gnd.n2875 gnd.n1351 9.3005
R11700 gnd.n4910 gnd.n1369 9.3005
R11701 gnd.n4909 gnd.n1370 9.3005
R11702 gnd.n4908 gnd.n1371 9.3005
R11703 gnd.n5044 gnd.n1137 9.3005
R11704 gnd.n1139 gnd.n1138 9.3005
R11705 gnd.n2530 gnd.n2529 9.3005
R11706 gnd.n2531 gnd.n1160 9.3005
R11707 gnd.n2533 gnd.n1161 9.3005
R11708 gnd.n2534 gnd.n1162 9.3005
R11709 gnd.n2537 gnd.n2535 9.3005
R11710 gnd.n2538 gnd.n1179 9.3005
R11711 gnd.n2540 gnd.n1180 9.3005
R11712 gnd.n2541 gnd.n1181 9.3005
R11713 gnd.n2631 gnd.n2542 9.3005
R11714 gnd.n2632 gnd.n1199 9.3005
R11715 gnd.n2633 gnd.n1200 9.3005
R11716 gnd.n2524 gnd.n1201 9.3005
R11717 gnd.n2684 gnd.n2525 9.3005
R11718 gnd.n2685 gnd.n1219 9.3005
R11719 gnd.n2686 gnd.n1220 9.3005
R11720 gnd.n2519 gnd.n1221 9.3005
R11721 gnd.n2699 gnd.n2520 9.3005
R11722 gnd.n2700 gnd.n1240 9.3005
R11723 gnd.n2702 gnd.n1241 9.3005
R11724 gnd.n2701 gnd.n1242 9.3005
R11725 gnd.n2510 gnd.n2507 9.3005
R11726 gnd.n2719 gnd.n2718 9.3005
R11727 gnd.n2717 gnd.n2508 9.3005
R11728 gnd.n2514 gnd.n2493 9.3005
R11729 gnd.n2513 gnd.n2494 9.3005
R11730 gnd.n2512 gnd.n2495 9.3005
R11731 gnd.n2511 gnd.n2471 9.3005
R11732 gnd.n2769 gnd.n2470 9.3005
R11733 gnd.n2771 gnd.n2770 9.3005
R11734 gnd.n2772 gnd.n1269 9.3005
R11735 gnd.n2775 gnd.n1270 9.3005
R11736 gnd.n2776 gnd.n1271 9.3005
R11737 gnd.n2781 gnd.n2777 9.3005
R11738 gnd.n2782 gnd.n1288 9.3005
R11739 gnd.n2786 gnd.n1289 9.3005
R11740 gnd.n2785 gnd.n1290 9.3005
R11741 gnd.n2784 gnd.n2783 9.3005
R11742 gnd.n2444 gnd.n1308 9.3005
R11743 gnd.n2851 gnd.n1309 9.3005
R11744 gnd.n2852 gnd.n1310 9.3005
R11745 gnd.n2854 gnd.n2853 9.3005
R11746 gnd.n2439 gnd.n1328 9.3005
R11747 gnd.n2866 gnd.n1329 9.3005
R11748 gnd.n2867 gnd.n1330 9.3005
R11749 gnd.n2869 gnd.n2868 9.3005
R11750 gnd.n2870 gnd.n1348 9.3005
R11751 gnd.n2873 gnd.n1349 9.3005
R11752 gnd.n2874 gnd.n1350 9.3005
R11753 gnd.n2878 gnd.n2875 9.3005
R11754 gnd.n2879 gnd.n1369 9.3005
R11755 gnd.n2881 gnd.n1370 9.3005
R11756 gnd.n2880 gnd.n1371 9.3005
R11757 gnd.n5044 gnd.n5043 9.3005
R11758 gnd.n5048 gnd.n5047 9.3005
R11759 gnd.n5051 gnd.n1132 9.3005
R11760 gnd.n5052 gnd.n1131 9.3005
R11761 gnd.n5055 gnd.n1130 9.3005
R11762 gnd.n5056 gnd.n1129 9.3005
R11763 gnd.n5059 gnd.n1128 9.3005
R11764 gnd.n5060 gnd.n1127 9.3005
R11765 gnd.n5063 gnd.n1126 9.3005
R11766 gnd.n5064 gnd.n1125 9.3005
R11767 gnd.n5067 gnd.n1124 9.3005
R11768 gnd.n5068 gnd.n1123 9.3005
R11769 gnd.n5071 gnd.n1122 9.3005
R11770 gnd.n5072 gnd.n1121 9.3005
R11771 gnd.n5075 gnd.n1120 9.3005
R11772 gnd.n5076 gnd.n1119 9.3005
R11773 gnd.n5079 gnd.n1118 9.3005
R11774 gnd.n5080 gnd.n1117 9.3005
R11775 gnd.n5083 gnd.n1116 9.3005
R11776 gnd.n5084 gnd.n1115 9.3005
R11777 gnd.n5087 gnd.n1114 9.3005
R11778 gnd.n5091 gnd.n1110 9.3005
R11779 gnd.n5092 gnd.n1109 9.3005
R11780 gnd.n5095 gnd.n1108 9.3005
R11781 gnd.n5096 gnd.n1107 9.3005
R11782 gnd.n5099 gnd.n1106 9.3005
R11783 gnd.n5100 gnd.n1105 9.3005
R11784 gnd.n5103 gnd.n1104 9.3005
R11785 gnd.n5104 gnd.n1103 9.3005
R11786 gnd.n5107 gnd.n1102 9.3005
R11787 gnd.n5108 gnd.n1101 9.3005
R11788 gnd.n5111 gnd.n1100 9.3005
R11789 gnd.n5112 gnd.n1099 9.3005
R11790 gnd.n5115 gnd.n1098 9.3005
R11791 gnd.n5116 gnd.n1097 9.3005
R11792 gnd.n5119 gnd.n1096 9.3005
R11793 gnd.n5120 gnd.n1095 9.3005
R11794 gnd.n5123 gnd.n1094 9.3005
R11795 gnd.n5124 gnd.n1093 9.3005
R11796 gnd.n5127 gnd.n1092 9.3005
R11797 gnd.n5129 gnd.n1089 9.3005
R11798 gnd.n5132 gnd.n1088 9.3005
R11799 gnd.n5133 gnd.n1087 9.3005
R11800 gnd.n5136 gnd.n1086 9.3005
R11801 gnd.n5137 gnd.n1085 9.3005
R11802 gnd.n5140 gnd.n1084 9.3005
R11803 gnd.n5141 gnd.n1083 9.3005
R11804 gnd.n5144 gnd.n1082 9.3005
R11805 gnd.n5145 gnd.n1081 9.3005
R11806 gnd.n5148 gnd.n1080 9.3005
R11807 gnd.n5149 gnd.n1079 9.3005
R11808 gnd.n5152 gnd.n1078 9.3005
R11809 gnd.n5153 gnd.n1077 9.3005
R11810 gnd.n5156 gnd.n1076 9.3005
R11811 gnd.n5158 gnd.n1075 9.3005
R11812 gnd.n5159 gnd.n1074 9.3005
R11813 gnd.n5160 gnd.n1073 9.3005
R11814 gnd.n5161 gnd.n1072 9.3005
R11815 gnd.n5088 gnd.n1111 9.3005
R11816 gnd.n5046 gnd.n1133 9.3005
R11817 gnd.n5038 gnd.n1147 9.3005
R11818 gnd.n5037 gnd.n1148 9.3005
R11819 gnd.n5036 gnd.n1149 9.3005
R11820 gnd.n1169 gnd.n1150 9.3005
R11821 gnd.n5026 gnd.n1170 9.3005
R11822 gnd.n5025 gnd.n1171 9.3005
R11823 gnd.n5024 gnd.n1172 9.3005
R11824 gnd.n1188 gnd.n1173 9.3005
R11825 gnd.n5014 gnd.n1189 9.3005
R11826 gnd.n5013 gnd.n1190 9.3005
R11827 gnd.n5012 gnd.n1191 9.3005
R11828 gnd.n1209 gnd.n1192 9.3005
R11829 gnd.n5002 gnd.n1210 9.3005
R11830 gnd.n5001 gnd.n1211 9.3005
R11831 gnd.n5000 gnd.n1212 9.3005
R11832 gnd.n1229 gnd.n1213 9.3005
R11833 gnd.n4990 gnd.n1230 9.3005
R11834 gnd.n4989 gnd.n1231 9.3005
R11835 gnd.n4988 gnd.n1232 9.3005
R11836 gnd.n1250 gnd.n1233 9.3005
R11837 gnd.n4978 gnd.n1251 9.3005
R11838 gnd.n1260 gnd.n1253 9.3005
R11839 gnd.n4964 gnd.n1278 9.3005
R11840 gnd.n4963 gnd.n1279 9.3005
R11841 gnd.n4962 gnd.n1280 9.3005
R11842 gnd.n1298 gnd.n1281 9.3005
R11843 gnd.n4952 gnd.n1299 9.3005
R11844 gnd.n4951 gnd.n1300 9.3005
R11845 gnd.n4950 gnd.n1301 9.3005
R11846 gnd.n1317 gnd.n1302 9.3005
R11847 gnd.n4940 gnd.n1318 9.3005
R11848 gnd.n4939 gnd.n1319 9.3005
R11849 gnd.n4938 gnd.n1320 9.3005
R11850 gnd.n1338 gnd.n1321 9.3005
R11851 gnd.n4928 gnd.n1339 9.3005
R11852 gnd.n4927 gnd.n1340 9.3005
R11853 gnd.n4926 gnd.n1341 9.3005
R11854 gnd.n1358 gnd.n1342 9.3005
R11855 gnd.n4916 gnd.n1359 9.3005
R11856 gnd.n4915 gnd.n1360 9.3005
R11857 gnd.n4914 gnd.n1361 9.3005
R11858 gnd.n1378 gnd.n1362 9.3005
R11859 gnd.n4904 gnd.n4903 9.3005
R11860 gnd.n1146 gnd.n1145 9.3005
R11861 gnd.n4975 gnd.n1258 9.3005
R11862 gnd.n4975 gnd.n4974 9.3005
R11863 gnd.n2647 gnd.n2646 9.3005
R11864 gnd.n2658 gnd.n2657 9.3005
R11865 gnd.n2659 gnd.n2645 9.3005
R11866 gnd.n2679 gnd.n2660 9.3005
R11867 gnd.n2678 gnd.n2661 9.3005
R11868 gnd.n2677 gnd.n2662 9.3005
R11869 gnd.n2665 gnd.n2663 9.3005
R11870 gnd.n2673 gnd.n2666 9.3005
R11871 gnd.n2672 gnd.n2667 9.3005
R11872 gnd.n2671 gnd.n2669 9.3005
R11873 gnd.n2668 gnd.n2501 9.3005
R11874 gnd.n2653 gnd.n2652 9.3005
R11875 gnd.n2649 gnd.n966 9.3005
R11876 gnd.n6585 gnd.n965 9.3005
R11877 gnd.n6586 gnd.n964 9.3005
R11878 gnd.n6587 gnd.n963 9.3005
R11879 gnd.n962 gnd.n958 9.3005
R11880 gnd.n6593 gnd.n957 9.3005
R11881 gnd.n6594 gnd.n956 9.3005
R11882 gnd.n6595 gnd.n955 9.3005
R11883 gnd.n954 gnd.n950 9.3005
R11884 gnd.n6601 gnd.n949 9.3005
R11885 gnd.n6602 gnd.n948 9.3005
R11886 gnd.n6603 gnd.n947 9.3005
R11887 gnd.n946 gnd.n942 9.3005
R11888 gnd.n6609 gnd.n941 9.3005
R11889 gnd.n6610 gnd.n940 9.3005
R11890 gnd.n6611 gnd.n939 9.3005
R11891 gnd.n938 gnd.n934 9.3005
R11892 gnd.n6617 gnd.n933 9.3005
R11893 gnd.n6618 gnd.n932 9.3005
R11894 gnd.n6619 gnd.n931 9.3005
R11895 gnd.n930 gnd.n926 9.3005
R11896 gnd.n6625 gnd.n925 9.3005
R11897 gnd.n6626 gnd.n924 9.3005
R11898 gnd.n6627 gnd.n923 9.3005
R11899 gnd.n922 gnd.n918 9.3005
R11900 gnd.n6633 gnd.n917 9.3005
R11901 gnd.n6634 gnd.n916 9.3005
R11902 gnd.n6635 gnd.n915 9.3005
R11903 gnd.n914 gnd.n910 9.3005
R11904 gnd.n6641 gnd.n909 9.3005
R11905 gnd.n6642 gnd.n908 9.3005
R11906 gnd.n6643 gnd.n907 9.3005
R11907 gnd.n906 gnd.n902 9.3005
R11908 gnd.n6649 gnd.n901 9.3005
R11909 gnd.n6650 gnd.n900 9.3005
R11910 gnd.n6651 gnd.n899 9.3005
R11911 gnd.n898 gnd.n894 9.3005
R11912 gnd.n6657 gnd.n893 9.3005
R11913 gnd.n6658 gnd.n892 9.3005
R11914 gnd.n6659 gnd.n891 9.3005
R11915 gnd.n890 gnd.n886 9.3005
R11916 gnd.n6665 gnd.n885 9.3005
R11917 gnd.n6666 gnd.n884 9.3005
R11918 gnd.n6667 gnd.n883 9.3005
R11919 gnd.n882 gnd.n878 9.3005
R11920 gnd.n6673 gnd.n877 9.3005
R11921 gnd.n6674 gnd.n876 9.3005
R11922 gnd.n6675 gnd.n875 9.3005
R11923 gnd.n874 gnd.n870 9.3005
R11924 gnd.n6681 gnd.n869 9.3005
R11925 gnd.n6682 gnd.n868 9.3005
R11926 gnd.n6683 gnd.n867 9.3005
R11927 gnd.n866 gnd.n862 9.3005
R11928 gnd.n6689 gnd.n861 9.3005
R11929 gnd.n6690 gnd.n860 9.3005
R11930 gnd.n6691 gnd.n859 9.3005
R11931 gnd.n858 gnd.n854 9.3005
R11932 gnd.n6697 gnd.n853 9.3005
R11933 gnd.n6698 gnd.n852 9.3005
R11934 gnd.n6699 gnd.n851 9.3005
R11935 gnd.n850 gnd.n846 9.3005
R11936 gnd.n6705 gnd.n845 9.3005
R11937 gnd.n6706 gnd.n844 9.3005
R11938 gnd.n6707 gnd.n843 9.3005
R11939 gnd.n842 gnd.n838 9.3005
R11940 gnd.n6713 gnd.n837 9.3005
R11941 gnd.n6714 gnd.n836 9.3005
R11942 gnd.n6715 gnd.n835 9.3005
R11943 gnd.n834 gnd.n830 9.3005
R11944 gnd.n6721 gnd.n829 9.3005
R11945 gnd.n6722 gnd.n828 9.3005
R11946 gnd.n6723 gnd.n827 9.3005
R11947 gnd.n826 gnd.n822 9.3005
R11948 gnd.n6729 gnd.n821 9.3005
R11949 gnd.n6730 gnd.n820 9.3005
R11950 gnd.n6731 gnd.n819 9.3005
R11951 gnd.n818 gnd.n814 9.3005
R11952 gnd.n6737 gnd.n813 9.3005
R11953 gnd.n6738 gnd.n812 9.3005
R11954 gnd.n6739 gnd.n811 9.3005
R11955 gnd.n810 gnd.n806 9.3005
R11956 gnd.n6745 gnd.n805 9.3005
R11957 gnd.n6746 gnd.n804 9.3005
R11958 gnd.n6747 gnd.n803 9.3005
R11959 gnd.n2651 gnd.n2650 9.3005
R11960 gnd.n4061 gnd.n4060 9.3005
R11961 gnd.n3197 gnd.n2399 9.3005
R11962 gnd.n2377 gnd.n2376 9.3005
R11963 gnd.n3225 gnd.n3224 9.3005
R11964 gnd.n3226 gnd.n2374 9.3005
R11965 gnd.n3231 gnd.n3230 9.3005
R11966 gnd.n3229 gnd.n2375 9.3005
R11967 gnd.n3228 gnd.n3227 9.3005
R11968 gnd.n2276 gnd.n2275 9.3005
R11969 gnd.n3262 gnd.n3261 9.3005
R11970 gnd.n3263 gnd.n2273 9.3005
R11971 gnd.n3266 gnd.n3265 9.3005
R11972 gnd.n3264 gnd.n2274 9.3005
R11973 gnd.n2265 gnd.n2264 9.3005
R11974 gnd.n3287 gnd.n3286 9.3005
R11975 gnd.n3288 gnd.n2262 9.3005
R11976 gnd.n3297 gnd.n3296 9.3005
R11977 gnd.n3295 gnd.n2263 9.3005
R11978 gnd.n3294 gnd.n3293 9.3005
R11979 gnd.n3292 gnd.n3289 9.3005
R11980 gnd.n2218 gnd.n2217 9.3005
R11981 gnd.n3373 gnd.n3372 9.3005
R11982 gnd.n3374 gnd.n2215 9.3005
R11983 gnd.n3395 gnd.n3394 9.3005
R11984 gnd.n3393 gnd.n2216 9.3005
R11985 gnd.n3392 gnd.n3391 9.3005
R11986 gnd.n3390 gnd.n3375 9.3005
R11987 gnd.n3389 gnd.n3388 9.3005
R11988 gnd.n3387 gnd.n3381 9.3005
R11989 gnd.n3386 gnd.n3385 9.3005
R11990 gnd.n3384 gnd.n3383 9.3005
R11991 gnd.n3382 gnd.n2168 9.3005
R11992 gnd.n2166 gnd.n2165 9.3005
R11993 gnd.n3475 gnd.n3474 9.3005
R11994 gnd.n3476 gnd.n2164 9.3005
R11995 gnd.n3478 gnd.n3477 9.3005
R11996 gnd.n2141 gnd.n2139 9.3005
R11997 gnd.n3524 gnd.n3523 9.3005
R11998 gnd.n3522 gnd.n2140 9.3005
R11999 gnd.n3521 gnd.n3520 9.3005
R12000 gnd.n2118 gnd.n2116 9.3005
R12001 gnd.n3583 gnd.n3582 9.3005
R12002 gnd.n3581 gnd.n2117 9.3005
R12003 gnd.n3580 gnd.n3579 9.3005
R12004 gnd.n3578 gnd.n2119 9.3005
R12005 gnd.n3577 gnd.n3576 9.3005
R12006 gnd.n3575 gnd.n3563 9.3005
R12007 gnd.n3574 gnd.n3573 9.3005
R12008 gnd.n3572 gnd.n3564 9.3005
R12009 gnd.n3571 gnd.n3570 9.3005
R12010 gnd.n2057 gnd.n2056 9.3005
R12011 gnd.n3692 gnd.n3691 9.3005
R12012 gnd.n3693 gnd.n2054 9.3005
R12013 gnd.n3696 gnd.n3695 9.3005
R12014 gnd.n3694 gnd.n2055 9.3005
R12015 gnd.n2028 gnd.n2027 9.3005
R12016 gnd.n3731 gnd.n3730 9.3005
R12017 gnd.n3732 gnd.n2025 9.3005
R12018 gnd.n3749 gnd.n3748 9.3005
R12019 gnd.n3747 gnd.n2026 9.3005
R12020 gnd.n3746 gnd.n3745 9.3005
R12021 gnd.n3744 gnd.n3733 9.3005
R12022 gnd.n3743 gnd.n3742 9.3005
R12023 gnd.n3741 gnd.n3738 9.3005
R12024 gnd.n3740 gnd.n3739 9.3005
R12025 gnd.n1972 gnd.n1971 9.3005
R12026 gnd.n3822 gnd.n3821 9.3005
R12027 gnd.n3823 gnd.n1969 9.3005
R12028 gnd.n3826 gnd.n3825 9.3005
R12029 gnd.n3824 gnd.n1970 9.3005
R12030 gnd.n1945 gnd.n1944 9.3005
R12031 gnd.n3864 gnd.n3863 9.3005
R12032 gnd.n3865 gnd.n1943 9.3005
R12033 gnd.n3867 gnd.n3866 9.3005
R12034 gnd.n1942 gnd.n1941 9.3005
R12035 gnd.n3875 gnd.n3874 9.3005
R12036 gnd.n3876 gnd.n1940 9.3005
R12037 gnd.n3878 gnd.n3877 9.3005
R12038 gnd.n3879 gnd.n1939 9.3005
R12039 gnd.n3883 gnd.n3882 9.3005
R12040 gnd.n3884 gnd.n1937 9.3005
R12041 gnd.n4064 gnd.n4063 9.3005
R12042 gnd.n4062 gnd.n1938 9.3005
R12043 gnd.n3199 gnd.n3198 9.3005
R12044 gnd.n3196 gnd.n3195 9.3005
R12045 gnd.n2757 gnd.n2479 9.3005
R12046 gnd.n2759 gnd.n2758 9.3005
R12047 gnd.n2465 gnd.n2463 9.3005
R12048 gnd.n2800 gnd.n2799 9.3005
R12049 gnd.n2798 gnd.n2464 9.3005
R12050 gnd.n2797 gnd.n2796 9.3005
R12051 gnd.n2795 gnd.n2466 9.3005
R12052 gnd.n2794 gnd.n2793 9.3005
R12053 gnd.n2792 gnd.n2469 9.3005
R12054 gnd.n2791 gnd.n2790 9.3005
R12055 gnd.n2447 gnd.n2446 9.3005
R12056 gnd.n2844 gnd.n2843 9.3005
R12057 gnd.n2845 gnd.n2445 9.3005
R12058 gnd.n2847 gnd.n2846 9.3005
R12059 gnd.n2442 gnd.n2441 9.3005
R12060 gnd.n2859 gnd.n2858 9.3005
R12061 gnd.n2860 gnd.n2440 9.3005
R12062 gnd.n2862 gnd.n2861 9.3005
R12063 gnd.n2433 gnd.n2431 9.3005
R12064 gnd.n2896 gnd.n2895 9.3005
R12065 gnd.n2894 gnd.n2432 9.3005
R12066 gnd.n2893 gnd.n2892 9.3005
R12067 gnd.n2891 gnd.n2434 9.3005
R12068 gnd.n2890 gnd.n2889 9.3005
R12069 gnd.n2888 gnd.n2437 9.3005
R12070 gnd.n2887 gnd.n2886 9.3005
R12071 gnd.n2885 gnd.n2438 9.3005
R12072 gnd.n3161 gnd.n3160 9.3005
R12073 gnd.n3159 gnd.n3158 9.3005
R12074 gnd.n3074 gnd.n3073 9.3005
R12075 gnd.n3153 gnd.n3152 9.3005
R12076 gnd.n3151 gnd.n3150 9.3005
R12077 gnd.n3086 gnd.n3085 9.3005
R12078 gnd.n3145 gnd.n3144 9.3005
R12079 gnd.n3143 gnd.n3142 9.3005
R12080 gnd.n3097 gnd.n3096 9.3005
R12081 gnd.n3137 gnd.n3136 9.3005
R12082 gnd.n3135 gnd.n3134 9.3005
R12083 gnd.n3109 gnd.n3108 9.3005
R12084 gnd.n3129 gnd.n3128 9.3005
R12085 gnd.n3127 gnd.n3126 9.3005
R12086 gnd.n3120 gnd.n2408 9.3005
R12087 gnd.n3186 gnd.n3185 9.3005
R12088 gnd.n2410 gnd.n2406 9.3005
R12089 gnd.n3192 gnd.n3191 9.3005
R12090 gnd.n3069 gnd.n3067 9.3005
R12091 gnd.n3194 gnd.n3193 9.3005
R12092 gnd.n2403 gnd.n2401 9.3005
R12093 gnd.n3184 gnd.n3183 9.3005
R12094 gnd.n3123 gnd.n2409 9.3005
R12095 gnd.n3125 gnd.n3124 9.3005
R12096 gnd.n3113 gnd.n3112 9.3005
R12097 gnd.n3131 gnd.n3130 9.3005
R12098 gnd.n3133 gnd.n3132 9.3005
R12099 gnd.n3103 gnd.n3102 9.3005
R12100 gnd.n3139 gnd.n3138 9.3005
R12101 gnd.n3141 gnd.n3140 9.3005
R12102 gnd.n3090 gnd.n3089 9.3005
R12103 gnd.n3147 gnd.n3146 9.3005
R12104 gnd.n3149 gnd.n3148 9.3005
R12105 gnd.n3080 gnd.n3079 9.3005
R12106 gnd.n3155 gnd.n3154 9.3005
R12107 gnd.n3157 gnd.n3156 9.3005
R12108 gnd.n3068 gnd.n3066 9.3005
R12109 gnd.n3163 gnd.n3162 9.3005
R12110 gnd.n3164 gnd.n3061 9.3005
R12111 gnd.n3166 gnd.n3165 9.3005
R12112 gnd.n3168 gnd.n2947 9.3005
R12113 gnd.n3170 gnd.n3169 9.3005
R12114 gnd.n3171 gnd.n2943 9.3005
R12115 gnd.n3173 gnd.n3172 9.3005
R12116 gnd.n3174 gnd.n2942 9.3005
R12117 gnd.n3176 gnd.n3175 9.3005
R12118 gnd.n3177 gnd.n2941 9.3005
R12119 gnd.n3216 gnd.n3215 9.3005
R12120 gnd.n3217 gnd.n2383 9.3005
R12121 gnd.n3220 gnd.n3219 9.3005
R12122 gnd.n3218 gnd.n2384 9.3005
R12123 gnd.n2362 gnd.n2361 9.3005
R12124 gnd.n3249 gnd.n3248 9.3005
R12125 gnd.n3250 gnd.n2359 9.3005
R12126 gnd.n3256 gnd.n3255 9.3005
R12127 gnd.n3254 gnd.n2360 9.3005
R12128 gnd.n3253 gnd.n3252 9.3005
R12129 gnd.n1509 gnd.n1507 9.3005
R12130 gnd.n4771 gnd.n4770 9.3005
R12131 gnd.n4769 gnd.n1508 9.3005
R12132 gnd.n4768 gnd.n4767 9.3005
R12133 gnd.n4766 gnd.n1510 9.3005
R12134 gnd.n4765 gnd.n4764 9.3005
R12135 gnd.n4763 gnd.n1514 9.3005
R12136 gnd.n4762 gnd.n4761 9.3005
R12137 gnd.n4760 gnd.n1515 9.3005
R12138 gnd.n4759 gnd.n4758 9.3005
R12139 gnd.n4757 gnd.n1519 9.3005
R12140 gnd.n4756 gnd.n4755 9.3005
R12141 gnd.n4754 gnd.n1520 9.3005
R12142 gnd.n4753 gnd.n4752 9.3005
R12143 gnd.n4751 gnd.n1524 9.3005
R12144 gnd.n4750 gnd.n4749 9.3005
R12145 gnd.n4748 gnd.n1525 9.3005
R12146 gnd.n4747 gnd.n4746 9.3005
R12147 gnd.n4745 gnd.n1529 9.3005
R12148 gnd.n4744 gnd.n4743 9.3005
R12149 gnd.n4742 gnd.n1530 9.3005
R12150 gnd.n4741 gnd.n4740 9.3005
R12151 gnd.n4739 gnd.n1534 9.3005
R12152 gnd.n4738 gnd.n4737 9.3005
R12153 gnd.n4736 gnd.n1535 9.3005
R12154 gnd.n4735 gnd.n4734 9.3005
R12155 gnd.n4733 gnd.n1539 9.3005
R12156 gnd.n4732 gnd.n4731 9.3005
R12157 gnd.n4730 gnd.n1540 9.3005
R12158 gnd.n4729 gnd.n4728 9.3005
R12159 gnd.n4727 gnd.n1544 9.3005
R12160 gnd.n4726 gnd.n4725 9.3005
R12161 gnd.n4724 gnd.n1545 9.3005
R12162 gnd.n4723 gnd.n4722 9.3005
R12163 gnd.n4721 gnd.n1549 9.3005
R12164 gnd.n4720 gnd.n4719 9.3005
R12165 gnd.n4718 gnd.n1550 9.3005
R12166 gnd.n4717 gnd.n4716 9.3005
R12167 gnd.n4715 gnd.n1554 9.3005
R12168 gnd.n4714 gnd.n4713 9.3005
R12169 gnd.n4712 gnd.n1555 9.3005
R12170 gnd.n4711 gnd.n4710 9.3005
R12171 gnd.n4709 gnd.n1559 9.3005
R12172 gnd.n4708 gnd.n4707 9.3005
R12173 gnd.n4706 gnd.n1560 9.3005
R12174 gnd.n4705 gnd.n4704 9.3005
R12175 gnd.n4703 gnd.n1564 9.3005
R12176 gnd.n4702 gnd.n4701 9.3005
R12177 gnd.n4700 gnd.n1565 9.3005
R12178 gnd.n4699 gnd.n4698 9.3005
R12179 gnd.n4697 gnd.n1569 9.3005
R12180 gnd.n4696 gnd.n4695 9.3005
R12181 gnd.n4694 gnd.n1570 9.3005
R12182 gnd.n4693 gnd.n4692 9.3005
R12183 gnd.n4691 gnd.n1574 9.3005
R12184 gnd.n4690 gnd.n4689 9.3005
R12185 gnd.n4688 gnd.n1575 9.3005
R12186 gnd.n4687 gnd.n4686 9.3005
R12187 gnd.n4685 gnd.n1579 9.3005
R12188 gnd.n4684 gnd.n4683 9.3005
R12189 gnd.n4682 gnd.n1580 9.3005
R12190 gnd.n4681 gnd.n4680 9.3005
R12191 gnd.n4679 gnd.n1584 9.3005
R12192 gnd.n4678 gnd.n4677 9.3005
R12193 gnd.n4676 gnd.n1585 9.3005
R12194 gnd.n4675 gnd.n4674 9.3005
R12195 gnd.n4673 gnd.n1589 9.3005
R12196 gnd.n4672 gnd.n4671 9.3005
R12197 gnd.n4670 gnd.n1590 9.3005
R12198 gnd.n4669 gnd.n4668 9.3005
R12199 gnd.n4667 gnd.n1594 9.3005
R12200 gnd.n4666 gnd.n4665 9.3005
R12201 gnd.n2386 gnd.n2385 9.3005
R12202 gnd.n3950 gnd.n3949 9.3005
R12203 gnd.n3946 gnd.n3945 9.3005
R12204 gnd.n3957 gnd.n3956 9.3005
R12205 gnd.n3958 gnd.n3944 9.3005
R12206 gnd.n3961 gnd.n3960 9.3005
R12207 gnd.n3959 gnd.n3942 9.3005
R12208 gnd.n3948 gnd.n1595 9.3005
R12209 gnd.n4049 gnd.n3898 9.3005
R12210 gnd.n3911 gnd.n3907 9.3005
R12211 gnd.n4043 gnd.n4042 9.3005
R12212 gnd.n4031 gnd.n3909 9.3005
R12213 gnd.n4030 gnd.n4029 9.3005
R12214 gnd.n3920 gnd.n3916 9.3005
R12215 gnd.n4023 gnd.n4022 9.3005
R12216 gnd.n4012 gnd.n3918 9.3005
R12217 gnd.n4011 gnd.n4010 9.3005
R12218 gnd.n3929 gnd.n3925 9.3005
R12219 gnd.n4004 gnd.n4003 9.3005
R12220 gnd.n3993 gnd.n3927 9.3005
R12221 gnd.n3992 gnd.n3991 9.3005
R12222 gnd.n3938 gnd.n3934 9.3005
R12223 gnd.n3985 gnd.n3984 9.3005
R12224 gnd.n3974 gnd.n3936 9.3005
R12225 gnd.n3973 gnd.n3972 9.3005
R12226 gnd.n4051 gnd.n4050 9.3005
R12227 gnd.n3902 gnd.n3901 9.3005
R12228 gnd.n3968 gnd.n3967 9.3005
R12229 gnd.n3969 gnd.n3941 9.3005
R12230 gnd.n3976 gnd.n3975 9.3005
R12231 gnd.n3939 gnd.n3937 9.3005
R12232 gnd.n3983 gnd.n3982 9.3005
R12233 gnd.n3933 gnd.n3932 9.3005
R12234 gnd.n3995 gnd.n3994 9.3005
R12235 gnd.n3930 gnd.n3928 9.3005
R12236 gnd.n4002 gnd.n4001 9.3005
R12237 gnd.n3924 gnd.n3923 9.3005
R12238 gnd.n4014 gnd.n4013 9.3005
R12239 gnd.n3921 gnd.n3919 9.3005
R12240 gnd.n4021 gnd.n4020 9.3005
R12241 gnd.n3915 gnd.n3914 9.3005
R12242 gnd.n4033 gnd.n4032 9.3005
R12243 gnd.n3912 gnd.n3910 9.3005
R12244 gnd.n4041 gnd.n4040 9.3005
R12245 gnd.n4039 gnd.n4038 9.3005
R12246 gnd.n4053 gnd.n4052 9.3005
R12247 gnd.n3899 gnd.n3893 9.3005
R12248 gnd.n3900 gnd.n3892 9.3005
R12249 gnd.n3888 gnd.n3885 9.3005
R12250 gnd.n1824 gnd.n1823 9.3005
R12251 gnd.n4437 gnd.n4436 9.3005
R12252 gnd.n4438 gnd.n1822 9.3005
R12253 gnd.n4440 gnd.n4439 9.3005
R12254 gnd.n1787 gnd.n1786 9.3005
R12255 gnd.n4451 gnd.n4450 9.3005
R12256 gnd.n4452 gnd.n1785 9.3005
R12257 gnd.n4454 gnd.n4453 9.3005
R12258 gnd.n1777 gnd.n1775 9.3005
R12259 gnd.n4490 gnd.n4489 9.3005
R12260 gnd.n4488 gnd.n1776 9.3005
R12261 gnd.n4487 gnd.n4486 9.3005
R12262 gnd.n4485 gnd.n1778 9.3005
R12263 gnd.n4484 gnd.n4483 9.3005
R12264 gnd.n4482 gnd.n1781 9.3005
R12265 gnd.n4481 gnd.n4480 9.3005
R12266 gnd.n4479 gnd.n1782 9.3005
R12267 gnd.n4478 gnd.n4477 9.3005
R12268 gnd.n1760 gnd.n1759 9.3005
R12269 gnd.n4549 gnd.n4548 9.3005
R12270 gnd.n4550 gnd.n1757 9.3005
R12271 gnd.n4555 gnd.n4554 9.3005
R12272 gnd.n4553 gnd.n1758 9.3005
R12273 gnd.n4552 gnd.n4551 9.3005
R12274 gnd.n81 gnd.n79 9.3005
R12275 gnd.n3890 gnd.n3889 9.3005
R12276 gnd.t100 gnd.n5300 9.24152
R12277 gnd.n6553 gnd.t205 9.24152
R12278 gnd.t306 gnd.n1019 9.24152
R12279 gnd.n1152 gnd.t217 9.24152
R12280 gnd.n2899 gnd.t14 9.24152
R12281 gnd.n1819 gnd.t36 9.24152
R12282 gnd.n7681 gnd.t228 9.24152
R12283 gnd.t124 gnd.t100 8.92286
R12284 gnd.n4774 gnd.t291 8.92286
R12285 gnd.n3276 gnd.n2266 8.92286
R12286 gnd.t8 gnd.n3301 8.92286
R12287 gnd.n3461 gnd.n2175 8.92286
R12288 gnd.n3506 gnd.n2145 8.92286
R12289 gnd.n3631 gnd.n2078 8.92286
R12290 gnd.n3702 gnd.n3701 8.92286
R12291 gnd.n1983 gnd.t84 8.92286
R12292 gnd.n3842 gnd.n3841 8.92286
R12293 gnd.n4179 gnd.t265 8.92286
R12294 gnd.n6407 gnd.n6382 8.92171
R12295 gnd.n6375 gnd.n6350 8.92171
R12296 gnd.n6343 gnd.n6318 8.92171
R12297 gnd.n6312 gnd.n6287 8.92171
R12298 gnd.n6280 gnd.n6255 8.92171
R12299 gnd.n6248 gnd.n6223 8.92171
R12300 gnd.n6216 gnd.n6191 8.92171
R12301 gnd.n6185 gnd.n6160 8.92171
R12302 gnd.n4111 gnd.n4093 8.72777
R12303 gnd.t326 gnd.n5411 8.60421
R12304 gnd.n5363 gnd.n5347 8.43656
R12305 gnd.n46 gnd.n30 8.43656
R12306 gnd.n3436 gnd.n2190 8.28555
R12307 gnd.n3527 gnd.n2128 8.28555
R12308 gnd.n3611 gnd.n2093 8.28555
R12309 gnd.n3667 gnd.n2045 8.28555
R12310 gnd.n6408 gnd.n6380 8.14595
R12311 gnd.n6376 gnd.n6348 8.14595
R12312 gnd.n6344 gnd.n6316 8.14595
R12313 gnd.n6313 gnd.n6285 8.14595
R12314 gnd.n6281 gnd.n6253 8.14595
R12315 gnd.n6249 gnd.n6221 8.14595
R12316 gnd.n6217 gnd.n6189 8.14595
R12317 gnd.n6186 gnd.n6158 8.14595
R12318 gnd.n2756 gnd.n0 8.10675
R12319 gnd.n7755 gnd.n7754 8.10675
R12320 gnd.n6413 gnd.n6412 7.97301
R12321 gnd.n5904 gnd.t325 7.9669
R12322 gnd.n7755 gnd.n78 7.86902
R12323 gnd.n4050 gnd.n3902 7.75808
R12324 gnd.n3191 gnd.n2406 7.75808
R12325 gnd.n7531 gnd.n349 7.75808
R12326 gnd.n2604 gnd.n2603 7.75808
R12327 gnd.n3269 gnd.n2270 7.64824
R12328 gnd.n3436 gnd.n2189 7.64824
R12329 gnd.t6 gnd.n3480 7.64824
R12330 gnd.n3528 gnd.t46 7.64824
R12331 gnd.n3538 gnd.n2128 7.64824
R12332 gnd.n3611 gnd.n2091 7.64824
R12333 gnd.t64 gnd.n2086 7.64824
R12334 gnd.n3630 gnd.t95 7.64824
R12335 gnd.n3667 gnd.n2036 7.64824
R12336 gnd.n5396 gnd.n5395 7.53171
R12337 gnd.t192 gnd.n5497 7.32958
R12338 gnd.n3269 gnd.t107 7.32958
R12339 gnd.t90 gnd.n3860 7.32958
R12340 gnd.n1487 gnd.n1486 7.30353
R12341 gnd.n4110 gnd.n4109 7.30353
R12342 gnd.n5806 gnd.n5805 7.01093
R12343 gnd.n5816 gnd.n5526 7.01093
R12344 gnd.n5815 gnd.n5529 7.01093
R12345 gnd.n5824 gnd.n5520 7.01093
R12346 gnd.n5828 gnd.n5827 7.01093
R12347 gnd.n5846 gnd.n5505 7.01093
R12348 gnd.n5845 gnd.n5508 7.01093
R12349 gnd.n5856 gnd.n5497 7.01093
R12350 gnd.n5498 gnd.n5486 7.01093
R12351 gnd.n5869 gnd.n5487 7.01093
R12352 gnd.n5880 gnd.n5479 7.01093
R12353 gnd.n5879 gnd.n5470 7.01093
R12354 gnd.n5472 gnd.n5454 7.01093
R12355 gnd.n5916 gnd.n5455 7.01093
R12356 gnd.n5905 gnd.n5904 7.01093
R12357 gnd.n5941 gnd.n5446 7.01093
R12358 gnd.n5952 gnd.n5951 7.01093
R12359 gnd.n5439 gnd.n5431 7.01093
R12360 gnd.n5981 gnd.n5419 7.01093
R12361 gnd.n5980 gnd.n5422 7.01093
R12362 gnd.n5991 gnd.n5411 7.01093
R12363 gnd.n5412 gnd.n5400 7.01093
R12364 gnd.n6002 gnd.n5401 7.01093
R12365 gnd.n6026 gnd.n5328 7.01093
R12366 gnd.n6025 gnd.n5319 7.01093
R12367 gnd.n5321 gnd.n5312 7.01093
R12368 gnd.n6048 gnd.n6047 7.01093
R12369 gnd.n6065 gnd.n5300 7.01093
R12370 gnd.n6064 gnd.n5303 7.01093
R12371 gnd.n6078 gnd.n5292 7.01093
R12372 gnd.n5293 gnd.n5282 7.01093
R12373 gnd.n6088 gnd.n5284 7.01093
R12374 gnd.n6121 gnd.n6120 7.01093
R12375 gnd.n6137 gnd.n6136 7.01093
R12376 gnd.n5263 gnd.n968 7.01093
R12377 gnd.n6580 gnd.n970 7.01093
R12378 gnd.n6101 gnd.n979 7.01093
R12379 gnd.n6574 gnd.n6573 7.01093
R12380 gnd.n6567 gnd.n990 7.01093
R12381 gnd.n6566 gnd.n993 7.01093
R12382 gnd.n6445 gnd.n1002 7.01093
R12383 gnd.n6560 gnd.n6559 7.01093
R12384 gnd.n6426 gnd.n1005 7.01093
R12385 gnd.n6553 gnd.n1016 7.01093
R12386 gnd.n6552 gnd.n1019 7.01093
R12387 gnd.n6456 gnd.n1027 7.01093
R12388 gnd.n6546 gnd.n6545 7.01093
R12389 gnd.n3283 gnd.n3276 7.01093
R12390 gnd.n3342 gnd.n2235 7.01093
R12391 gnd.t47 gnd.n3341 7.01093
R12392 gnd.n3461 gnd.n3460 7.01093
R12393 gnd.n3481 gnd.t6 7.01093
R12394 gnd.n3480 gnd.n2145 7.01093
R12395 gnd.n3631 gnd.n3630 7.01093
R12396 gnd.t95 gnd.n3629 7.01093
R12397 gnd.n3702 gnd.n2049 7.01093
R12398 gnd.n3783 gnd.t165 7.01093
R12399 gnd.n3799 gnd.n3798 7.01093
R12400 gnd.n3844 gnd.n3842 7.01093
R12401 gnd.n5487 gnd.t74 6.69227
R12402 gnd.n6047 gnd.t124 6.69227
R12403 gnd.t98 gnd.n6437 6.69227
R12404 gnd.n5016 gnd.t129 6.69227
R12405 gnd.n2864 gnd.t92 6.69227
R12406 gnd.t194 gnd.n2230 6.69227
R12407 gnd.n3736 gnd.t105 6.69227
R12408 gnd.n4456 gnd.t58 6.69227
R12409 gnd.n7510 gnd.t81 6.69227
R12410 gnd.n4240 gnd.n4239 6.5566
R12411 gnd.n2285 gnd.n2284 6.5566
R12412 gnd.n4792 gnd.n4788 6.5566
R12413 gnd.n4118 gnd.n4117 6.5566
R12414 gnd.n6581 gnd.n6580 6.37362
R12415 gnd.n2356 gnd.n2355 6.37362
R12416 gnd.t291 gnd.t271 6.37362
R12417 gnd.n3403 gnd.n2204 6.37362
R12418 gnd.n3488 gnd.t44 6.37362
R12419 gnd.n3546 gnd.n2122 6.37362
R12420 gnd.n3558 gnd.n2109 6.37362
R12421 gnd.n3680 gnd.t96 6.37362
R12422 gnd.n3727 gnd.n2032 6.37362
R12423 gnd.n3841 gnd.t202 6.37362
R12424 gnd.n3852 gnd.t202 6.37362
R12425 gnd.n4179 gnd.n1902 6.37362
R12426 gnd.n3183 gnd.n2413 6.20656
R12427 gnd.n4053 gnd.n3897 6.20656
R12428 gnd.n5940 gnd.t136 6.05496
R12429 gnd.n5939 gnd.t190 6.05496
R12430 gnd.t4 gnd.n5412 6.05496
R12431 gnd.t189 gnd.n5276 6.05496
R12432 gnd.n2788 gnd.t50 6.05496
R12433 gnd.t164 gnd.t321 6.05496
R12434 gnd.t11 gnd.t127 6.05496
R12435 gnd.n4475 gnd.t34 6.05496
R12436 gnd.n6410 gnd.n6380 5.81868
R12437 gnd.n6378 gnd.n6348 5.81868
R12438 gnd.n6346 gnd.n6316 5.81868
R12439 gnd.n6315 gnd.n6285 5.81868
R12440 gnd.n6283 gnd.n6253 5.81868
R12441 gnd.n6251 gnd.n6221 5.81868
R12442 gnd.n6219 gnd.n6189 5.81868
R12443 gnd.n6188 gnd.n6158 5.81868
R12444 gnd.n2259 gnd.n2258 5.73631
R12445 gnd.n3302 gnd.n3299 5.73631
R12446 gnd.n2170 gnd.n2158 5.73631
R12447 gnd.n3472 gnd.n2151 5.73631
R12448 gnd.t46 gnd.n3527 5.73631
R12449 gnd.n2093 gnd.t64 5.73631
R12450 gnd.n3568 gnd.n3566 5.73631
R12451 gnd.n3638 gnd.n2067 5.73631
R12452 gnd.n3819 gnd.n1974 5.73631
R12453 gnd.n1976 gnd.n1966 5.73631
R12454 gnd.n4249 gnd.n1861 5.62001
R12455 gnd.n4854 gnd.n1429 5.62001
R12456 gnd.n4854 gnd.n1430 5.62001
R12457 gnd.n4249 gnd.n1862 5.62001
R12458 gnd.n5624 gnd.n5623 5.4308
R12459 gnd.n5243 gnd.n5241 5.4308
R12460 gnd.n5401 gnd.t65 5.41765
R12461 gnd.t187 gnd.n6036 5.41765
R12462 gnd.n6122 gnd.t40 5.41765
R12463 gnd.n2761 gnd.t27 5.41765
R12464 gnd.t334 gnd.n3419 5.41765
R12465 gnd.n3659 gnd.t70 5.41765
R12466 gnd.n4572 gnd.t2 5.41765
R12467 gnd.n2629 gnd.n1194 5.09899
R12468 gnd.n5010 gnd.n1197 5.09899
R12469 gnd.n2635 gnd.n1204 5.09899
R12470 gnd.n5004 gnd.n1207 5.09899
R12471 gnd.n2682 gnd.n2681 5.09899
R12472 gnd.n4998 gnd.n1217 5.09899
R12473 gnd.n2688 gnd.n1224 5.09899
R12474 gnd.n4992 gnd.n1227 5.09899
R12475 gnd.n2697 gnd.n1235 5.09899
R12476 gnd.n4986 gnd.n1238 5.09899
R12477 gnd.n2704 gnd.n1245 5.09899
R12478 gnd.n4980 gnd.n1248 5.09899
R12479 gnd.n2724 gnd.n2503 5.09899
R12480 gnd.n2723 gnd.n2506 5.09899
R12481 gnd.n2715 gnd.n2488 5.09899
R12482 gnd.n2747 gnd.n2490 5.09899
R12483 gnd.n2752 gnd.n2484 5.09899
R12484 gnd.n2741 gnd.n2740 5.09899
R12485 gnd.n2761 gnd.n2474 5.09899
R12486 gnd.n2766 gnd.n2460 5.09899
R12487 gnd.n2803 gnd.n2802 5.09899
R12488 gnd.n4972 gnd.n1265 5.09899
R12489 gnd.n2773 gnd.n1274 5.09899
R12490 gnd.n2779 gnd.n1283 5.09899
R12491 gnd.n4960 gnd.n1286 5.09899
R12492 gnd.n2788 gnd.n1293 5.09899
R12493 gnd.n4954 gnd.n1296 5.09899
R12494 gnd.n2841 gnd.n2840 5.09899
R12495 gnd.n4948 gnd.n1306 5.09899
R12496 gnd.n2849 gnd.n1313 5.09899
R12497 gnd.n2856 gnd.n1323 5.09899
R12498 gnd.n4936 gnd.n1326 5.09899
R12499 gnd.n2864 gnd.n1333 5.09899
R12500 gnd.n4930 gnd.n1336 5.09899
R12501 gnd.n2899 gnd.n2898 5.09899
R12502 gnd.n4924 gnd.n1346 5.09899
R12503 gnd.n2871 gnd.n1353 5.09899
R12504 gnd.n4918 gnd.n1356 5.09899
R12505 gnd.n2876 gnd.n1364 5.09899
R12506 gnd.n4912 gnd.n1367 5.09899
R12507 gnd.n2883 gnd.n1373 5.09899
R12508 gnd.n4906 gnd.n1376 5.09899
R12509 gnd.t97 gnd.n3333 5.09899
R12510 gnd.n3411 gnd.n2208 5.09899
R12511 gnd.n3587 gnd.n2113 5.09899
R12512 gnd.n3595 gnd.n2106 5.09899
R12513 gnd.n3760 gnd.n2016 5.09899
R12514 gnd.n2007 gnd.t48 5.09899
R12515 gnd.n4648 gnd.n4647 5.09899
R12516 gnd.n3886 gnd.n1621 5.09899
R12517 gnd.n4641 gnd.n1630 5.09899
R12518 gnd.n4434 gnd.n1633 5.09899
R12519 gnd.n4635 gnd.n1642 5.09899
R12520 gnd.n4442 gnd.n1645 5.09899
R12521 gnd.n4629 gnd.n1653 5.09899
R12522 gnd.n4448 gnd.n1819 5.09899
R12523 gnd.n4623 gnd.n1662 5.09899
R12524 gnd.n4456 gnd.n1665 5.09899
R12525 gnd.n4617 gnd.n1673 5.09899
R12526 gnd.n4492 gnd.n1676 5.09899
R12527 gnd.n4463 gnd.n1685 5.09899
R12528 gnd.n4605 gnd.n1693 5.09899
R12529 gnd.n4468 gnd.n4467 5.09899
R12530 gnd.n4599 gnd.n1702 5.09899
R12531 gnd.n4475 gnd.n1705 5.09899
R12532 gnd.n4593 gnd.n1713 5.09899
R12533 gnd.n4516 gnd.n1716 5.09899
R12534 gnd.n4546 gnd.n1725 5.09899
R12535 gnd.n4581 gnd.n1731 5.09899
R12536 gnd.n4558 gnd.n4557 5.09899
R12537 gnd.n4575 gnd.n1740 5.09899
R12538 gnd.n4572 gnd.n1743 5.09899
R12539 gnd.n4571 gnd.n1751 5.09899
R12540 gnd.n4536 gnd.n4524 5.09899
R12541 gnd.n7749 gnd.n85 5.09899
R12542 gnd.n381 gnd.n87 5.09899
R12543 gnd.n7446 gnd.n7441 5.09899
R12544 gnd.n7741 gnd.n102 5.09899
R12545 gnd.n7452 gnd.n105 5.09899
R12546 gnd.n7735 gnd.n114 5.09899
R12547 gnd.n7460 gnd.n374 5.09899
R12548 gnd.n7729 gnd.n123 5.09899
R12549 gnd.n7466 gnd.n371 5.09899
R12550 gnd.n7723 gnd.n132 5.09899
R12551 gnd.n7474 gnd.n135 5.09899
R12552 gnd.n7717 gnd.n143 5.09899
R12553 gnd.n7480 gnd.n146 5.09899
R12554 gnd.n7711 gnd.n153 5.09899
R12555 gnd.n7489 gnd.n362 5.09899
R12556 gnd.n7705 gnd.n163 5.09899
R12557 gnd.n6408 gnd.n6407 5.04292
R12558 gnd.n6376 gnd.n6375 5.04292
R12559 gnd.n6344 gnd.n6343 5.04292
R12560 gnd.n6313 gnd.n6312 5.04292
R12561 gnd.n6281 gnd.n6280 5.04292
R12562 gnd.n6249 gnd.n6248 5.04292
R12563 gnd.n6217 gnd.n6216 5.04292
R12564 gnd.n6186 gnd.n6185 5.04292
R12565 gnd.t191 gnd.n5962 4.78034
R12566 gnd.n6078 gnd.t101 4.78034
R12567 gnd.n2704 gnd.t109 4.78034
R12568 gnd.n4966 gnd.t62 4.78034
R12569 gnd.t351 gnd.n3245 4.78034
R12570 gnd.n4246 gnd.t249 4.78034
R12571 gnd.n4080 gnd.t146 4.78034
R12572 gnd.n4587 gnd.t151 4.78034
R12573 gnd.n7735 gnd.t88 4.78034
R12574 gnd.n5936 gnd.n5935 4.74817
R12575 gnd.n5931 gnd.n5930 4.74817
R12576 gnd.n5927 gnd.n5926 4.74817
R12577 gnd.n5923 gnd.n5398 4.74817
R12578 gnd.n5935 gnd.n5934 4.74817
R12579 gnd.n5933 gnd.n5931 4.74817
R12580 gnd.n5929 gnd.n5927 4.74817
R12581 gnd.n5925 gnd.n5923 4.74817
R12582 gnd.n4583 gnd.n98 4.74817
R12583 gnd.n1745 gnd.n96 4.74817
R12584 gnd.n7747 gnd.n91 4.74817
R12585 gnd.n7745 gnd.n92 4.74817
R12586 gnd.n1729 gnd.n98 4.74817
R12587 gnd.n1747 gnd.n96 4.74817
R12588 gnd.n1744 gnd.n91 4.74817
R12589 gnd.n7746 gnd.n7745 4.74817
R12590 gnd.n2727 gnd.n2726 4.74817
R12591 gnd.n2732 gnd.n2499 4.74817
R12592 gnd.n2738 gnd.n2734 4.74817
R12593 gnd.n2736 gnd.n2735 4.74817
R12594 gnd.n2458 gnd.n2456 4.74817
R12595 gnd.n4510 gnd.n1754 4.74817
R12596 gnd.n4563 gnd.n4562 4.74817
R12597 gnd.n4568 gnd.n4567 4.74817
R12598 gnd.n4564 gnd.n384 4.74817
R12599 gnd.n7438 gnd.n7437 4.74817
R12600 gnd.n4511 gnd.n4510 4.74817
R12601 gnd.n4562 gnd.n4561 4.74817
R12602 gnd.n4569 gnd.n4568 4.74817
R12603 gnd.n4566 gnd.n4564 4.74817
R12604 gnd.n7439 gnd.n7438 4.74817
R12605 gnd.n4977 gnd.n4976 4.74817
R12606 gnd.n2750 gnd.n1257 4.74817
R12607 gnd.n2763 gnd.n1256 4.74817
R12608 gnd.n1259 gnd.n1255 4.74817
R12609 gnd.n4976 gnd.n1252 4.74817
R12610 gnd.n2487 gnd.n1257 4.74817
R12611 gnd.n2749 gnd.n1256 4.74817
R12612 gnd.n2764 gnd.n1255 4.74817
R12613 gnd.n2728 gnd.n2727 4.74817
R12614 gnd.n2729 gnd.n2499 4.74817
R12615 gnd.n2734 gnd.n2733 4.74817
R12616 gnd.n2737 gnd.n2736 4.74817
R12617 gnd.n2459 gnd.n2458 4.74817
R12618 gnd.n5395 gnd.n5394 4.74296
R12619 gnd.n78 gnd.n77 4.74296
R12620 gnd.n5363 gnd.n5362 4.7074
R12621 gnd.n5379 gnd.n5378 4.7074
R12622 gnd.n46 gnd.n45 4.7074
R12623 gnd.n62 gnd.n61 4.7074
R12624 gnd.n5395 gnd.n5379 4.65959
R12625 gnd.n78 gnd.n62 4.65959
R12626 gnd.n4340 gnd.n4250 4.6132
R12627 gnd.n4855 gnd.n1428 4.6132
R12628 gnd.n3309 gnd.n2251 4.46168
R12629 gnd.n3300 gnd.n2240 4.46168
R12630 gnd.n3458 gnd.t186 4.46168
R12631 gnd.n3468 gnd.n3467 4.46168
R12632 gnd.n3497 gnd.n2153 4.46168
R12633 gnd.n3645 gnd.n2072 4.46168
R12634 gnd.n3689 gnd.n2059 4.46168
R12635 gnd.t83 gnd.n3688 4.46168
R12636 gnd.n3809 gnd.n1982 4.46168
R12637 gnd.n3829 gnd.n3828 4.46168
R12638 gnd.t316 gnd.n1907 4.46168
R12639 gnd.n4106 gnd.n4093 4.46111
R12640 gnd.n6393 gnd.n6389 4.38594
R12641 gnd.n6361 gnd.n6357 4.38594
R12642 gnd.n6329 gnd.n6325 4.38594
R12643 gnd.n6298 gnd.n6294 4.38594
R12644 gnd.n6266 gnd.n6262 4.38594
R12645 gnd.n6234 gnd.n6230 4.38594
R12646 gnd.n6202 gnd.n6198 4.38594
R12647 gnd.n6171 gnd.n6167 4.38594
R12648 gnd.n6404 gnd.n6382 4.26717
R12649 gnd.n6372 gnd.n6350 4.26717
R12650 gnd.n6340 gnd.n6318 4.26717
R12651 gnd.n6309 gnd.n6287 4.26717
R12652 gnd.n6277 gnd.n6255 4.26717
R12653 gnd.n6245 gnd.n6223 4.26717
R12654 gnd.n6213 gnd.n6191 4.26717
R12655 gnd.n6182 gnd.n6160 4.26717
R12656 gnd.t99 gnd.n5893 4.14303
R12657 gnd.t73 gnd.n970 4.14303
R12658 gnd.n2635 gnd.t115 4.14303
R12659 gnd.n4942 gnd.t30 4.14303
R12660 gnd.t235 gnd.n1367 4.14303
R12661 gnd.t213 gnd.n1630 4.14303
R12662 gnd.n4611 gnd.t32 4.14303
R12663 gnd.n7711 gnd.t23 4.14303
R12664 gnd.n6412 gnd.n6411 4.08274
R12665 gnd.n4239 gnd.n4238 4.05904
R12666 gnd.n2286 gnd.n2285 4.05904
R12667 gnd.n4795 gnd.n4788 4.05904
R12668 gnd.n4119 gnd.n4118 4.05904
R12669 gnd.n15 gnd.n7 3.99943
R12670 gnd.n4781 gnd.n4780 3.82437
R12671 gnd.n3368 gnd.n2221 3.82437
R12672 gnd.n3409 gnd.t61 3.82437
R12673 gnd.n3429 gnd.n3428 3.82437
R12674 gnd.n3517 gnd.n2142 3.82437
R12675 gnd.n3518 gnd.t164 3.82437
R12676 gnd.n3559 gnd.t11 3.82437
R12677 gnd.n3604 gnd.n3603 3.82437
R12678 gnd.n3719 gnd.n2030 3.82437
R12679 gnd.n3752 gnd.t323 3.82437
R12680 gnd.n3769 gnd.n3768 3.82437
R12681 gnd.n4087 gnd.n1910 3.82437
R12682 gnd.n5397 gnd.n5396 3.81325
R12683 gnd.n5379 gnd.n5363 3.72967
R12684 gnd.n62 gnd.n46 3.72967
R12685 gnd.n6412 gnd.n6284 3.70378
R12686 gnd.n15 gnd.n14 3.60163
R12687 gnd.n6403 gnd.n6384 3.49141
R12688 gnd.n6371 gnd.n6352 3.49141
R12689 gnd.n6339 gnd.n6320 3.49141
R12690 gnd.n6308 gnd.n6289 3.49141
R12691 gnd.n6276 gnd.n6257 3.49141
R12692 gnd.n6244 gnd.n6225 3.49141
R12693 gnd.n6212 gnd.n6193 3.49141
R12694 gnd.n6181 gnd.n6162 3.49141
R12695 gnd.n4321 gnd.n4320 3.29747
R12696 gnd.n4320 gnd.n4258 3.29747
R12697 gnd.n7640 gnd.n7637 3.29747
R12698 gnd.n7641 gnd.n7640 3.29747
R12699 gnd.n5129 gnd.n5128 3.29747
R12700 gnd.n5128 gnd.n5127 3.29747
R12701 gnd.n4871 gnd.n4870 3.29747
R12702 gnd.n4870 gnd.n4869 3.29747
R12703 gnd.n4773 gnd.n1504 3.18706
R12704 gnd.n2259 gnd.t279 3.18706
R12705 gnd.n3340 gnd.n2228 3.18706
R12706 gnd.n3349 gnd.t45 3.18706
R12707 gnd.t45 gnd.n2213 3.18706
R12708 gnd.n3447 gnd.n3445 3.18706
R12709 gnd.n3508 gnd.n3507 3.18706
R12710 gnd.n3619 gnd.n3618 3.18706
R12711 gnd.n3700 gnd.n3699 3.18706
R12712 gnd.t324 gnd.n2019 3.18706
R12713 gnd.n3650 gnd.t324 3.18706
R12714 gnd.n3785 gnd.n3784 3.18706
R12715 gnd.n3852 gnd.n1951 3.18706
R12716 gnd.n3860 gnd.t316 3.18706
R12717 gnd.n5894 gnd.t99 2.8684
R12718 gnd.n3316 gnd.t68 2.8684
R12719 gnd.t66 gnd.n3818 2.8684
R12720 gnd.n5380 gnd.t104 2.82907
R12721 gnd.n5380 gnd.t93 2.82907
R12722 gnd.n5382 gnd.t51 2.82907
R12723 gnd.n5382 gnd.t144 2.82907
R12724 gnd.n5384 gnd.t360 2.82907
R12725 gnd.n5384 gnd.t63 2.82907
R12726 gnd.n5386 gnd.t340 2.82907
R12727 gnd.n5386 gnd.t339 2.82907
R12728 gnd.n5388 gnd.t110 2.82907
R12729 gnd.n5388 gnd.t174 2.82907
R12730 gnd.n5390 gnd.t358 2.82907
R12731 gnd.n5390 gnd.t159 2.82907
R12732 gnd.n5392 gnd.t130 2.82907
R12733 gnd.n5392 gnd.t116 2.82907
R12734 gnd.n5333 gnd.t31 2.82907
R12735 gnd.n5333 gnd.t367 2.82907
R12736 gnd.n5335 gnd.t133 2.82907
R12737 gnd.n5335 gnd.t139 2.82907
R12738 gnd.n5337 gnd.t336 2.82907
R12739 gnd.n5337 gnd.t160 2.82907
R12740 gnd.n5339 gnd.t175 2.82907
R12741 gnd.n5339 gnd.t343 2.82907
R12742 gnd.n5341 gnd.t122 2.82907
R12743 gnd.n5341 gnd.t60 2.82907
R12744 gnd.n5343 gnd.t362 2.82907
R12745 gnd.n5343 gnd.t39 2.82907
R12746 gnd.n5345 gnd.t169 2.82907
R12747 gnd.n5345 gnd.t180 2.82907
R12748 gnd.n5348 gnd.t111 2.82907
R12749 gnd.n5348 gnd.t331 2.82907
R12750 gnd.n5350 gnd.t80 2.82907
R12751 gnd.n5350 gnd.t332 2.82907
R12752 gnd.n5352 gnd.t333 2.82907
R12753 gnd.n5352 gnd.t119 2.82907
R12754 gnd.n5354 gnd.t19 2.82907
R12755 gnd.n5354 gnd.t162 2.82907
R12756 gnd.n5356 gnd.t342 2.82907
R12757 gnd.n5356 gnd.t26 2.82907
R12758 gnd.n5358 gnd.t177 2.82907
R12759 gnd.n5358 gnd.t354 2.82907
R12760 gnd.n5360 gnd.t353 2.82907
R12761 gnd.n5360 gnd.t361 2.82907
R12762 gnd.n5364 gnd.t196 2.82907
R12763 gnd.n5364 gnd.t348 2.82907
R12764 gnd.n5366 gnd.t167 2.82907
R12765 gnd.n5366 gnd.t347 2.82907
R12766 gnd.n5368 gnd.t21 2.82907
R12767 gnd.n5368 gnd.t344 2.82907
R12768 gnd.n5370 gnd.t345 2.82907
R12769 gnd.n5370 gnd.t28 2.82907
R12770 gnd.n5372 gnd.t132 2.82907
R12771 gnd.n5372 gnd.t365 2.82907
R12772 gnd.n5374 gnd.t79 2.82907
R12773 gnd.n5374 gnd.t157 2.82907
R12774 gnd.n5376 gnd.t134 2.82907
R12775 gnd.n5376 gnd.t150 2.82907
R12776 gnd.n75 gnd.t114 2.82907
R12777 gnd.n75 gnd.t193 2.82907
R12778 gnd.n73 gnd.t185 2.82907
R12779 gnd.n73 gnd.t76 2.82907
R12780 gnd.n71 gnd.t145 2.82907
R12781 gnd.n71 gnd.t359 2.82907
R12782 gnd.n69 gnd.t7 2.82907
R12783 gnd.n69 gnd.t13 2.82907
R12784 gnd.n67 gnd.t338 2.82907
R12785 gnd.n67 gnd.t171 2.82907
R12786 gnd.n65 gnd.t184 2.82907
R12787 gnd.n65 gnd.t87 2.82907
R12788 gnd.n63 gnd.t341 2.82907
R12789 gnd.n63 gnd.t337 2.82907
R12790 gnd.n28 gnd.t24 2.82907
R12791 gnd.n28 gnd.t330 2.82907
R12792 gnd.n26 gnd.t356 2.82907
R12793 gnd.n26 gnd.t199 2.82907
R12794 gnd.n24 gnd.t118 2.82907
R12795 gnd.n24 gnd.t168 2.82907
R12796 gnd.n22 gnd.t3 2.82907
R12797 gnd.n22 gnd.t156 2.82907
R12798 gnd.n20 gnd.t153 2.82907
R12799 gnd.n20 gnd.t121 2.82907
R12800 gnd.n18 gnd.t197 2.82907
R12801 gnd.n18 gnd.t135 2.82907
R12802 gnd.n16 gnd.t59 2.82907
R12803 gnd.n16 gnd.t33 2.82907
R12804 gnd.n43 gnd.t29 2.82907
R12805 gnd.n43 gnd.t364 2.82907
R12806 gnd.n41 gnd.t363 2.82907
R12807 gnd.n41 gnd.t113 2.82907
R12808 gnd.n39 gnd.t55 2.82907
R12809 gnd.n39 gnd.t123 2.82907
R12810 gnd.n37 gnd.t350 2.82907
R12811 gnd.n37 gnd.t346 2.82907
R12812 gnd.n35 gnd.t152 2.82907
R12813 gnd.n35 gnd.t149 2.82907
R12814 gnd.n33 gnd.t22 2.82907
R12815 gnd.n33 gnd.t357 2.82907
R12816 gnd.n31 gnd.t158 2.82907
R12817 gnd.n31 gnd.t170 2.82907
R12818 gnd.n59 gnd.t77 2.82907
R12819 gnd.n59 gnd.t82 2.82907
R12820 gnd.n57 gnd.t53 2.82907
R12821 gnd.n57 gnd.t198 2.82907
R12822 gnd.n55 gnd.t148 2.82907
R12823 gnd.n55 gnd.t89 2.82907
R12824 gnd.n53 gnd.t155 2.82907
R12825 gnd.n53 gnd.t329 2.82907
R12826 gnd.n51 gnd.t327 2.82907
R12827 gnd.n51 gnd.t126 2.82907
R12828 gnd.n49 gnd.t1 2.82907
R12829 gnd.n49 gnd.t35 2.82907
R12830 gnd.n47 gnd.t112 2.82907
R12831 gnd.n47 gnd.t161 2.82907
R12832 gnd.n6400 gnd.n6399 2.71565
R12833 gnd.n6368 gnd.n6367 2.71565
R12834 gnd.n6336 gnd.n6335 2.71565
R12835 gnd.n6305 gnd.n6304 2.71565
R12836 gnd.n6273 gnd.n6272 2.71565
R12837 gnd.n6241 gnd.n6240 2.71565
R12838 gnd.n6209 gnd.n6208 2.71565
R12839 gnd.n6178 gnd.n6177 2.71565
R12840 gnd.n4774 gnd.n1502 2.54975
R12841 gnd.n3358 gnd.n3357 2.54975
R12842 gnd.n3334 gnd.t97 2.54975
R12843 gnd.n3448 gnd.n2184 2.54975
R12844 gnd.n3448 gnd.t49 2.54975
R12845 gnd.n3528 gnd.n2135 2.54975
R12846 gnd.n3620 gnd.n2086 2.54975
R12847 gnd.n3709 gnd.t117 2.54975
R12848 gnd.n3709 gnd.n3708 2.54975
R12849 gnd.n3776 gnd.t48 2.54975
R12850 gnd.n3786 gnd.n1996 2.54975
R12851 gnd.n1960 gnd.n1947 2.54975
R12852 gnd.n5935 gnd.n5397 2.27742
R12853 gnd.n5931 gnd.n5397 2.27742
R12854 gnd.n5927 gnd.n5397 2.27742
R12855 gnd.n5923 gnd.n5397 2.27742
R12856 gnd.n7744 gnd.n98 2.27742
R12857 gnd.n7744 gnd.n96 2.27742
R12858 gnd.n7744 gnd.n91 2.27742
R12859 gnd.n7745 gnd.n7744 2.27742
R12860 gnd.n4510 gnd.n95 2.27742
R12861 gnd.n4562 gnd.n95 2.27742
R12862 gnd.n4568 gnd.n95 2.27742
R12863 gnd.n4564 gnd.n95 2.27742
R12864 gnd.n7438 gnd.n95 2.27742
R12865 gnd.n4976 gnd.n4975 2.27742
R12866 gnd.n4975 gnd.n1257 2.27742
R12867 gnd.n4975 gnd.n1256 2.27742
R12868 gnd.n4975 gnd.n1255 2.27742
R12869 gnd.n2727 gnd.n1254 2.27742
R12870 gnd.n2499 gnd.n1254 2.27742
R12871 gnd.n2734 gnd.n1254 2.27742
R12872 gnd.n2736 gnd.n1254 2.27742
R12873 gnd.n2458 gnd.n1254 2.27742
R12874 gnd.t275 gnd.n5815 2.23109
R12875 gnd.n5963 gnd.t191 2.23109
R12876 gnd.t85 gnd.n2153 2.23109
R12877 gnd.t321 gnd.n3517 2.23109
R12878 gnd.n3604 gnd.t127 2.23109
R12879 gnd.t16 gnd.n2072 2.23109
R12880 gnd.n6396 gnd.n6386 1.93989
R12881 gnd.n6364 gnd.n6354 1.93989
R12882 gnd.n6332 gnd.n6322 1.93989
R12883 gnd.n6301 gnd.n6291 1.93989
R12884 gnd.n6269 gnd.n6259 1.93989
R12885 gnd.n6237 gnd.n6227 1.93989
R12886 gnd.n6205 gnd.n6195 1.93989
R12887 gnd.n6174 gnd.n6164 1.93989
R12888 gnd.n2349 gnd.n1493 1.91244
R12889 gnd.n2349 gnd.t232 1.91244
R12890 gnd.n3342 gnd.t47 1.91244
R12891 gnd.n3370 gnd.n2220 1.91244
R12892 gnd.n3378 gnd.n3377 1.91244
R12893 gnd.n3537 gnd.n2130 1.91244
R12894 gnd.n2100 gnd.n2099 1.91244
R12895 gnd.n3721 gnd.n3720 1.91244
R12896 gnd.n2010 gnd.n2008 1.91244
R12897 gnd.n3799 gnd.t165 1.91244
R12898 gnd.n4089 gnd.n4088 1.91244
R12899 gnd.n5828 gnd.t9 1.59378
R12900 gnd.n6037 gnd.t187 1.59378
R12901 gnd.n6111 gnd.t40 1.59378
R12902 gnd.n3334 gnd.t194 1.59378
R12903 gnd.t102 gnd.n2175 1.59378
R12904 gnd.n3701 gnd.t172 1.59378
R12905 gnd.n3776 gnd.t105 1.59378
R12906 gnd.t300 gnd.n2356 1.27512
R12907 gnd.n3282 gnd.n3281 1.27512
R12908 gnd.n3302 gnd.t8 1.27512
R12909 gnd.n3325 gnd.n3324 1.27512
R12910 gnd.n3420 gnd.t61 1.27512
R12911 gnd.n3459 gnd.n3458 1.27512
R12912 gnd.n3481 gnd.n2162 1.27512
R12913 gnd.n3629 gnd.n3628 1.27512
R12914 gnd.n3688 gnd.n2060 1.27512
R12915 gnd.n3657 gnd.t323 1.27512
R12916 gnd.n3797 gnd.n3796 1.27512
R12917 gnd.t84 gnd.n1974 1.27512
R12918 gnd.n3828 gnd.t221 1.27512
R12919 gnd.n3845 gnd.n1956 1.27512
R12920 gnd.n5625 gnd.n5624 1.16414
R12921 gnd.n6471 gnd.n5241 1.16414
R12922 gnd.n6395 gnd.n6388 1.16414
R12923 gnd.n6363 gnd.n6356 1.16414
R12924 gnd.n6331 gnd.n6324 1.16414
R12925 gnd.n6300 gnd.n6293 1.16414
R12926 gnd.n6268 gnd.n6261 1.16414
R12927 gnd.n6236 gnd.n6229 1.16414
R12928 gnd.n6204 gnd.n6197 1.16414
R12929 gnd.n6173 gnd.n6166 1.16414
R12930 gnd.n4250 gnd.n1860 0.970197
R12931 gnd.n4855 gnd.n1425 0.970197
R12932 gnd.n6379 gnd.n6347 0.962709
R12933 gnd.n6411 gnd.n6379 0.962709
R12934 gnd.n6252 gnd.n6220 0.962709
R12935 gnd.n6284 gnd.n6252 0.962709
R12936 gnd.t136 gnd.n5939 0.956468
R12937 gnd.n5283 gnd.t189 0.956468
R12938 gnd.t38 gnd.n1227 0.956468
R12939 gnd.n2443 gnd.t30 0.956468
R12940 gnd.n4851 gnd.n1465 0.956468
R12941 gnd.t107 gnd.n3268 0.956468
R12942 gnd.n3861 gnd.t90 0.956468
R12943 gnd.n4246 gnd.n1865 0.956468
R12944 gnd.n4493 gnd.t32 0.956468
R12945 gnd.n371 gnd.t52 0.956468
R12946 gnd.n2 gnd.n1 0.672012
R12947 gnd.n3 gnd.n2 0.672012
R12948 gnd.n4 gnd.n3 0.672012
R12949 gnd.n5 gnd.n4 0.672012
R12950 gnd.n6 gnd.n5 0.672012
R12951 gnd.n7 gnd.n6 0.672012
R12952 gnd.n9 gnd.n8 0.672012
R12953 gnd.n10 gnd.n9 0.672012
R12954 gnd.n11 gnd.n10 0.672012
R12955 gnd.n12 gnd.n11 0.672012
R12956 gnd.n13 gnd.n12 0.672012
R12957 gnd.n14 gnd.n13 0.672012
R12958 gnd.t271 gnd.n4773 0.637812
R12959 gnd.t252 gnd.n3282 0.637812
R12960 gnd.n3398 gnd.n3397 0.637812
R12961 gnd.n3419 gnd.n3417 0.637812
R12962 gnd.n3428 gnd.t200 0.637812
R12963 gnd.n3548 gnd.n3547 0.637812
R12964 gnd.n3594 gnd.n3593 0.637812
R12965 gnd.t183 gnd.n3719 0.637812
R12966 gnd.n3660 gnd.n3659 0.637812
R12967 gnd.n3759 gnd.n3758 0.637812
R12968 gnd.t224 gnd.n1951 0.637812
R12969 gnd.n3869 gnd.t265 0.637812
R12970 gnd gnd.n0 0.59317
R12971 gnd.n5394 gnd.n5393 0.573776
R12972 gnd.n5393 gnd.n5391 0.573776
R12973 gnd.n5391 gnd.n5389 0.573776
R12974 gnd.n5389 gnd.n5387 0.573776
R12975 gnd.n5387 gnd.n5385 0.573776
R12976 gnd.n5385 gnd.n5383 0.573776
R12977 gnd.n5383 gnd.n5381 0.573776
R12978 gnd.n5347 gnd.n5346 0.573776
R12979 gnd.n5346 gnd.n5344 0.573776
R12980 gnd.n5344 gnd.n5342 0.573776
R12981 gnd.n5342 gnd.n5340 0.573776
R12982 gnd.n5340 gnd.n5338 0.573776
R12983 gnd.n5338 gnd.n5336 0.573776
R12984 gnd.n5336 gnd.n5334 0.573776
R12985 gnd.n5362 gnd.n5361 0.573776
R12986 gnd.n5361 gnd.n5359 0.573776
R12987 gnd.n5359 gnd.n5357 0.573776
R12988 gnd.n5357 gnd.n5355 0.573776
R12989 gnd.n5355 gnd.n5353 0.573776
R12990 gnd.n5353 gnd.n5351 0.573776
R12991 gnd.n5351 gnd.n5349 0.573776
R12992 gnd.n5378 gnd.n5377 0.573776
R12993 gnd.n5377 gnd.n5375 0.573776
R12994 gnd.n5375 gnd.n5373 0.573776
R12995 gnd.n5373 gnd.n5371 0.573776
R12996 gnd.n5371 gnd.n5369 0.573776
R12997 gnd.n5369 gnd.n5367 0.573776
R12998 gnd.n5367 gnd.n5365 0.573776
R12999 gnd.n66 gnd.n64 0.573776
R13000 gnd.n68 gnd.n66 0.573776
R13001 gnd.n70 gnd.n68 0.573776
R13002 gnd.n72 gnd.n70 0.573776
R13003 gnd.n74 gnd.n72 0.573776
R13004 gnd.n76 gnd.n74 0.573776
R13005 gnd.n77 gnd.n76 0.573776
R13006 gnd.n19 gnd.n17 0.573776
R13007 gnd.n21 gnd.n19 0.573776
R13008 gnd.n23 gnd.n21 0.573776
R13009 gnd.n25 gnd.n23 0.573776
R13010 gnd.n27 gnd.n25 0.573776
R13011 gnd.n29 gnd.n27 0.573776
R13012 gnd.n30 gnd.n29 0.573776
R13013 gnd.n34 gnd.n32 0.573776
R13014 gnd.n36 gnd.n34 0.573776
R13015 gnd.n38 gnd.n36 0.573776
R13016 gnd.n40 gnd.n38 0.573776
R13017 gnd.n42 gnd.n40 0.573776
R13018 gnd.n44 gnd.n42 0.573776
R13019 gnd.n45 gnd.n44 0.573776
R13020 gnd.n50 gnd.n48 0.573776
R13021 gnd.n52 gnd.n50 0.573776
R13022 gnd.n54 gnd.n52 0.573776
R13023 gnd.n56 gnd.n54 0.573776
R13024 gnd.n58 gnd.n56 0.573776
R13025 gnd.n60 gnd.n58 0.573776
R13026 gnd.n61 gnd.n60 0.573776
R13027 gnd.n7756 gnd.n7755 0.553533
R13028 gnd.n7529 gnd.n7528 0.505073
R13029 gnd.n2608 gnd.n2605 0.505073
R13030 gnd.n4062 gnd.n4061 0.489829
R13031 gnd.n3198 gnd.n3196 0.489829
R13032 gnd.n2941 gnd.n2385 0.489829
R13033 gnd.n4666 gnd.n1595 0.489829
R13034 gnd.n6461 gnd.n6460 0.486781
R13035 gnd.n5677 gnd.n5573 0.48678
R13036 gnd.n6542 gnd.n6541 0.480683
R13037 gnd.n5745 gnd.n5523 0.480683
R13038 gnd.n7672 gnd.n7671 0.470012
R13039 gnd.n4276 gnd.n1625 0.470012
R13040 gnd.n4903 gnd.n4902 0.470012
R13041 gnd.n1146 gnd.n1072 0.470012
R13042 gnd.n803 gnd.n798 0.425805
R13043 gnd.n7205 gnd.n7204 0.425805
R13044 gnd.n7418 gnd.n7417 0.425805
R13045 gnd.n2652 gnd.n2651 0.425805
R13046 gnd.n7744 gnd.n95 0.4255
R13047 gnd.n4975 gnd.n1254 0.4255
R13048 gnd.n3123 gnd.n2413 0.388379
R13049 gnd.n6392 gnd.n6391 0.388379
R13050 gnd.n6360 gnd.n6359 0.388379
R13051 gnd.n6328 gnd.n6327 0.388379
R13052 gnd.n6297 gnd.n6296 0.388379
R13053 gnd.n6265 gnd.n6264 0.388379
R13054 gnd.n6233 gnd.n6232 0.388379
R13055 gnd.n6201 gnd.n6200 0.388379
R13056 gnd.n6170 gnd.n6169 0.388379
R13057 gnd.n4039 gnd.n3897 0.388379
R13058 gnd.n7756 gnd.n15 0.374463
R13059 gnd.n6438 gnd.t98 0.319156
R13060 gnd.n2490 gnd.t18 0.319156
R13061 gnd.n2778 gnd.t62 0.319156
R13062 gnd.n3212 gnd.t261 0.319156
R13063 gnd.t245 gnd.n4067 0.319156
R13064 gnd.n4515 gnd.t151 0.319156
R13065 gnd.t12 gnd.n85 0.319156
R13066 gnd.n5671 gnd.n5670 0.311721
R13067 gnd gnd.n7756 0.295112
R13068 gnd.n7562 gnd.n7561 0.293183
R13069 gnd.n5045 gnd.n1136 0.293183
R13070 gnd.n2438 gnd.n2400 0.27489
R13071 gnd.n3891 gnd.n3890 0.27489
R13072 gnd.n6511 gnd.n6510 0.268793
R13073 gnd.n7563 gnd.n7562 0.258122
R13074 gnd.n4426 gnd.n4425 0.258122
R13075 gnd.n3060 gnd.n3059 0.258122
R13076 gnd.n5046 gnd.n5045 0.258122
R13077 gnd.n6510 gnd.n6509 0.241354
R13078 gnd.n4341 gnd.n4340 0.229039
R13079 gnd.n4340 gnd.n1859 0.229039
R13080 gnd.n1428 gnd.n1424 0.229039
R13081 gnd.n2980 gnd.n1428 0.229039
R13082 gnd.n5800 gnd.n5541 0.206293
R13083 gnd.n5396 gnd.n0 0.169152
R13084 gnd.n6409 gnd.n6381 0.155672
R13085 gnd.n6402 gnd.n6381 0.155672
R13086 gnd.n6402 gnd.n6401 0.155672
R13087 gnd.n6401 gnd.n6385 0.155672
R13088 gnd.n6394 gnd.n6385 0.155672
R13089 gnd.n6394 gnd.n6393 0.155672
R13090 gnd.n6377 gnd.n6349 0.155672
R13091 gnd.n6370 gnd.n6349 0.155672
R13092 gnd.n6370 gnd.n6369 0.155672
R13093 gnd.n6369 gnd.n6353 0.155672
R13094 gnd.n6362 gnd.n6353 0.155672
R13095 gnd.n6362 gnd.n6361 0.155672
R13096 gnd.n6345 gnd.n6317 0.155672
R13097 gnd.n6338 gnd.n6317 0.155672
R13098 gnd.n6338 gnd.n6337 0.155672
R13099 gnd.n6337 gnd.n6321 0.155672
R13100 gnd.n6330 gnd.n6321 0.155672
R13101 gnd.n6330 gnd.n6329 0.155672
R13102 gnd.n6314 gnd.n6286 0.155672
R13103 gnd.n6307 gnd.n6286 0.155672
R13104 gnd.n6307 gnd.n6306 0.155672
R13105 gnd.n6306 gnd.n6290 0.155672
R13106 gnd.n6299 gnd.n6290 0.155672
R13107 gnd.n6299 gnd.n6298 0.155672
R13108 gnd.n6282 gnd.n6254 0.155672
R13109 gnd.n6275 gnd.n6254 0.155672
R13110 gnd.n6275 gnd.n6274 0.155672
R13111 gnd.n6274 gnd.n6258 0.155672
R13112 gnd.n6267 gnd.n6258 0.155672
R13113 gnd.n6267 gnd.n6266 0.155672
R13114 gnd.n6250 gnd.n6222 0.155672
R13115 gnd.n6243 gnd.n6222 0.155672
R13116 gnd.n6243 gnd.n6242 0.155672
R13117 gnd.n6242 gnd.n6226 0.155672
R13118 gnd.n6235 gnd.n6226 0.155672
R13119 gnd.n6235 gnd.n6234 0.155672
R13120 gnd.n6218 gnd.n6190 0.155672
R13121 gnd.n6211 gnd.n6190 0.155672
R13122 gnd.n6211 gnd.n6210 0.155672
R13123 gnd.n6210 gnd.n6194 0.155672
R13124 gnd.n6203 gnd.n6194 0.155672
R13125 gnd.n6203 gnd.n6202 0.155672
R13126 gnd.n6187 gnd.n6159 0.155672
R13127 gnd.n6180 gnd.n6159 0.155672
R13128 gnd.n6180 gnd.n6179 0.155672
R13129 gnd.n6179 gnd.n6163 0.155672
R13130 gnd.n6172 gnd.n6163 0.155672
R13131 gnd.n6172 gnd.n6171 0.155672
R13132 gnd.n6541 gnd.n5171 0.152939
R13133 gnd.n5173 gnd.n5171 0.152939
R13134 gnd.n5177 gnd.n5173 0.152939
R13135 gnd.n5178 gnd.n5177 0.152939
R13136 gnd.n5179 gnd.n5178 0.152939
R13137 gnd.n5180 gnd.n5179 0.152939
R13138 gnd.n5184 gnd.n5180 0.152939
R13139 gnd.n5185 gnd.n5184 0.152939
R13140 gnd.n5186 gnd.n5185 0.152939
R13141 gnd.n5187 gnd.n5186 0.152939
R13142 gnd.n5191 gnd.n5187 0.152939
R13143 gnd.n5192 gnd.n5191 0.152939
R13144 gnd.n5193 gnd.n5192 0.152939
R13145 gnd.n5194 gnd.n5193 0.152939
R13146 gnd.n5199 gnd.n5194 0.152939
R13147 gnd.n6511 gnd.n5199 0.152939
R13148 gnd.n5819 gnd.n5523 0.152939
R13149 gnd.n5820 gnd.n5819 0.152939
R13150 gnd.n5821 gnd.n5820 0.152939
R13151 gnd.n5821 gnd.n5502 0.152939
R13152 gnd.n5849 gnd.n5502 0.152939
R13153 gnd.n5850 gnd.n5849 0.152939
R13154 gnd.n5851 gnd.n5850 0.152939
R13155 gnd.n5852 gnd.n5851 0.152939
R13156 gnd.n5852 gnd.n5476 0.152939
R13157 gnd.n5883 gnd.n5476 0.152939
R13158 gnd.n5884 gnd.n5883 0.152939
R13159 gnd.n5885 gnd.n5884 0.152939
R13160 gnd.n5886 gnd.n5885 0.152939
R13161 gnd.n5887 gnd.n5886 0.152939
R13162 gnd.n5887 gnd.n5443 0.152939
R13163 gnd.n5944 gnd.n5443 0.152939
R13164 gnd.n5945 gnd.n5944 0.152939
R13165 gnd.n5946 gnd.n5945 0.152939
R13166 gnd.n5947 gnd.n5946 0.152939
R13167 gnd.n5947 gnd.n5416 0.152939
R13168 gnd.n5984 gnd.n5416 0.152939
R13169 gnd.n5985 gnd.n5984 0.152939
R13170 gnd.n5986 gnd.n5985 0.152939
R13171 gnd.n5987 gnd.n5986 0.152939
R13172 gnd.n5987 gnd.n5325 0.152939
R13173 gnd.n6029 gnd.n5325 0.152939
R13174 gnd.n6030 gnd.n6029 0.152939
R13175 gnd.n6031 gnd.n6030 0.152939
R13176 gnd.n6032 gnd.n6031 0.152939
R13177 gnd.n6032 gnd.n5297 0.152939
R13178 gnd.n6068 gnd.n5297 0.152939
R13179 gnd.n6069 gnd.n6068 0.152939
R13180 gnd.n6070 gnd.n6069 0.152939
R13181 gnd.n6071 gnd.n6070 0.152939
R13182 gnd.n6072 gnd.n6071 0.152939
R13183 gnd.n6072 gnd.n5267 0.152939
R13184 gnd.n6125 gnd.n5267 0.152939
R13185 gnd.n6126 gnd.n6125 0.152939
R13186 gnd.n6127 gnd.n6126 0.152939
R13187 gnd.n6128 gnd.n6127 0.152939
R13188 gnd.n6130 gnd.n6128 0.152939
R13189 gnd.n6130 gnd.n6129 0.152939
R13190 gnd.n6129 gnd.n985 0.152939
R13191 gnd.n986 gnd.n985 0.152939
R13192 gnd.n987 gnd.n986 0.152939
R13193 gnd.n1009 gnd.n987 0.152939
R13194 gnd.n1010 gnd.n1009 0.152939
R13195 gnd.n1011 gnd.n1010 0.152939
R13196 gnd.n1012 gnd.n1011 0.152939
R13197 gnd.n1013 gnd.n1012 0.152939
R13198 gnd.n5169 gnd.n1013 0.152939
R13199 gnd.n5170 gnd.n5169 0.152939
R13200 gnd.n6542 gnd.n5170 0.152939
R13201 gnd.n5746 gnd.n5745 0.152939
R13202 gnd.n5747 gnd.n5746 0.152939
R13203 gnd.n5748 gnd.n5747 0.152939
R13204 gnd.n5749 gnd.n5748 0.152939
R13205 gnd.n5750 gnd.n5749 0.152939
R13206 gnd.n5751 gnd.n5750 0.152939
R13207 gnd.n5752 gnd.n5751 0.152939
R13208 gnd.n5753 gnd.n5752 0.152939
R13209 gnd.n5754 gnd.n5753 0.152939
R13210 gnd.n5755 gnd.n5754 0.152939
R13211 gnd.n5756 gnd.n5755 0.152939
R13212 gnd.n5757 gnd.n5756 0.152939
R13213 gnd.n5758 gnd.n5757 0.152939
R13214 gnd.n5759 gnd.n5758 0.152939
R13215 gnd.n5763 gnd.n5759 0.152939
R13216 gnd.n5763 gnd.n5541 0.152939
R13217 gnd.n6509 gnd.n5201 0.152939
R13218 gnd.n5203 gnd.n5201 0.152939
R13219 gnd.n5207 gnd.n5203 0.152939
R13220 gnd.n5208 gnd.n5207 0.152939
R13221 gnd.n5209 gnd.n5208 0.152939
R13222 gnd.n5210 gnd.n5209 0.152939
R13223 gnd.n5214 gnd.n5210 0.152939
R13224 gnd.n5215 gnd.n5214 0.152939
R13225 gnd.n5216 gnd.n5215 0.152939
R13226 gnd.n5217 gnd.n5216 0.152939
R13227 gnd.n5221 gnd.n5217 0.152939
R13228 gnd.n5222 gnd.n5221 0.152939
R13229 gnd.n5223 gnd.n5222 0.152939
R13230 gnd.n5224 gnd.n5223 0.152939
R13231 gnd.n5228 gnd.n5224 0.152939
R13232 gnd.n5229 gnd.n5228 0.152939
R13233 gnd.n5230 gnd.n5229 0.152939
R13234 gnd.n5231 gnd.n5230 0.152939
R13235 gnd.n5235 gnd.n5231 0.152939
R13236 gnd.n5236 gnd.n5235 0.152939
R13237 gnd.n5237 gnd.n5236 0.152939
R13238 gnd.n5238 gnd.n5237 0.152939
R13239 gnd.n5245 gnd.n5238 0.152939
R13240 gnd.n5246 gnd.n5245 0.152939
R13241 gnd.n5247 gnd.n5246 0.152939
R13242 gnd.n6461 gnd.n5247 0.152939
R13243 gnd.n6006 gnd.n6005 0.152939
R13244 gnd.n6007 gnd.n6006 0.152939
R13245 gnd.n6008 gnd.n6007 0.152939
R13246 gnd.n6009 gnd.n6008 0.152939
R13247 gnd.n6010 gnd.n6009 0.152939
R13248 gnd.n6011 gnd.n6010 0.152939
R13249 gnd.n6012 gnd.n6011 0.152939
R13250 gnd.n6013 gnd.n6012 0.152939
R13251 gnd.n6013 gnd.n5279 0.152939
R13252 gnd.n6091 gnd.n5279 0.152939
R13253 gnd.n6092 gnd.n6091 0.152939
R13254 gnd.n6093 gnd.n6092 0.152939
R13255 gnd.n6094 gnd.n6093 0.152939
R13256 gnd.n6095 gnd.n6094 0.152939
R13257 gnd.n6096 gnd.n6095 0.152939
R13258 gnd.n6097 gnd.n6096 0.152939
R13259 gnd.n6098 gnd.n6097 0.152939
R13260 gnd.n6099 gnd.n6098 0.152939
R13261 gnd.n6099 gnd.n5252 0.152939
R13262 gnd.n6442 gnd.n5252 0.152939
R13263 gnd.n6443 gnd.n6442 0.152939
R13264 gnd.n6444 gnd.n6443 0.152939
R13265 gnd.n6444 gnd.n5250 0.152939
R13266 gnd.n6452 gnd.n5250 0.152939
R13267 gnd.n6453 gnd.n6452 0.152939
R13268 gnd.n6454 gnd.n6453 0.152939
R13269 gnd.n6454 gnd.n5248 0.152939
R13270 gnd.n6460 gnd.n5248 0.152939
R13271 gnd.n5678 gnd.n5677 0.152939
R13272 gnd.n5679 gnd.n5678 0.152939
R13273 gnd.n5679 gnd.n5561 0.152939
R13274 gnd.n5693 gnd.n5561 0.152939
R13275 gnd.n5694 gnd.n5693 0.152939
R13276 gnd.n5695 gnd.n5694 0.152939
R13277 gnd.n5695 gnd.n5548 0.152939
R13278 gnd.n5709 gnd.n5548 0.152939
R13279 gnd.n5710 gnd.n5709 0.152939
R13280 gnd.n5711 gnd.n5710 0.152939
R13281 gnd.n5712 gnd.n5711 0.152939
R13282 gnd.n5713 gnd.n5712 0.152939
R13283 gnd.n5714 gnd.n5713 0.152939
R13284 gnd.n5715 gnd.n5714 0.152939
R13285 gnd.n5716 gnd.n5715 0.152939
R13286 gnd.n5717 gnd.n5716 0.152939
R13287 gnd.n5718 gnd.n5717 0.152939
R13288 gnd.n5719 gnd.n5718 0.152939
R13289 gnd.n5720 gnd.n5719 0.152939
R13290 gnd.n5720 gnd.n5483 0.152939
R13291 gnd.n5872 gnd.n5483 0.152939
R13292 gnd.n5873 gnd.n5872 0.152939
R13293 gnd.n5874 gnd.n5873 0.152939
R13294 gnd.n5875 gnd.n5874 0.152939
R13295 gnd.n5875 gnd.n5450 0.152939
R13296 gnd.n5919 gnd.n5450 0.152939
R13297 gnd.n5920 gnd.n5919 0.152939
R13298 gnd.n5921 gnd.n5920 0.152939
R13299 gnd.n5670 gnd.n5577 0.152939
R13300 gnd.n5580 gnd.n5577 0.152939
R13301 gnd.n5581 gnd.n5580 0.152939
R13302 gnd.n5582 gnd.n5581 0.152939
R13303 gnd.n5585 gnd.n5582 0.152939
R13304 gnd.n5586 gnd.n5585 0.152939
R13305 gnd.n5587 gnd.n5586 0.152939
R13306 gnd.n5588 gnd.n5587 0.152939
R13307 gnd.n5591 gnd.n5588 0.152939
R13308 gnd.n5592 gnd.n5591 0.152939
R13309 gnd.n5593 gnd.n5592 0.152939
R13310 gnd.n5594 gnd.n5593 0.152939
R13311 gnd.n5597 gnd.n5594 0.152939
R13312 gnd.n5598 gnd.n5597 0.152939
R13313 gnd.n5599 gnd.n5598 0.152939
R13314 gnd.n5600 gnd.n5599 0.152939
R13315 gnd.n5603 gnd.n5600 0.152939
R13316 gnd.n5604 gnd.n5603 0.152939
R13317 gnd.n5605 gnd.n5604 0.152939
R13318 gnd.n5606 gnd.n5605 0.152939
R13319 gnd.n5609 gnd.n5606 0.152939
R13320 gnd.n5610 gnd.n5609 0.152939
R13321 gnd.n5613 gnd.n5610 0.152939
R13322 gnd.n5614 gnd.n5613 0.152939
R13323 gnd.n5616 gnd.n5614 0.152939
R13324 gnd.n5616 gnd.n5573 0.152939
R13325 gnd.n6754 gnd.n798 0.152939
R13326 gnd.n6755 gnd.n6754 0.152939
R13327 gnd.n6756 gnd.n6755 0.152939
R13328 gnd.n6756 gnd.n792 0.152939
R13329 gnd.n6764 gnd.n792 0.152939
R13330 gnd.n6765 gnd.n6764 0.152939
R13331 gnd.n6766 gnd.n6765 0.152939
R13332 gnd.n6766 gnd.n786 0.152939
R13333 gnd.n6774 gnd.n786 0.152939
R13334 gnd.n6775 gnd.n6774 0.152939
R13335 gnd.n6776 gnd.n6775 0.152939
R13336 gnd.n6776 gnd.n780 0.152939
R13337 gnd.n6784 gnd.n780 0.152939
R13338 gnd.n6785 gnd.n6784 0.152939
R13339 gnd.n6786 gnd.n6785 0.152939
R13340 gnd.n6786 gnd.n774 0.152939
R13341 gnd.n6794 gnd.n774 0.152939
R13342 gnd.n6795 gnd.n6794 0.152939
R13343 gnd.n6796 gnd.n6795 0.152939
R13344 gnd.n6796 gnd.n768 0.152939
R13345 gnd.n6804 gnd.n768 0.152939
R13346 gnd.n6805 gnd.n6804 0.152939
R13347 gnd.n6806 gnd.n6805 0.152939
R13348 gnd.n6806 gnd.n762 0.152939
R13349 gnd.n6814 gnd.n762 0.152939
R13350 gnd.n6815 gnd.n6814 0.152939
R13351 gnd.n6816 gnd.n6815 0.152939
R13352 gnd.n6816 gnd.n756 0.152939
R13353 gnd.n6824 gnd.n756 0.152939
R13354 gnd.n6825 gnd.n6824 0.152939
R13355 gnd.n6826 gnd.n6825 0.152939
R13356 gnd.n6826 gnd.n750 0.152939
R13357 gnd.n6834 gnd.n750 0.152939
R13358 gnd.n6835 gnd.n6834 0.152939
R13359 gnd.n6836 gnd.n6835 0.152939
R13360 gnd.n6836 gnd.n744 0.152939
R13361 gnd.n6844 gnd.n744 0.152939
R13362 gnd.n6845 gnd.n6844 0.152939
R13363 gnd.n6846 gnd.n6845 0.152939
R13364 gnd.n6846 gnd.n738 0.152939
R13365 gnd.n6854 gnd.n738 0.152939
R13366 gnd.n6855 gnd.n6854 0.152939
R13367 gnd.n6856 gnd.n6855 0.152939
R13368 gnd.n6856 gnd.n732 0.152939
R13369 gnd.n6864 gnd.n732 0.152939
R13370 gnd.n6865 gnd.n6864 0.152939
R13371 gnd.n6866 gnd.n6865 0.152939
R13372 gnd.n6866 gnd.n726 0.152939
R13373 gnd.n6874 gnd.n726 0.152939
R13374 gnd.n6875 gnd.n6874 0.152939
R13375 gnd.n6876 gnd.n6875 0.152939
R13376 gnd.n6876 gnd.n720 0.152939
R13377 gnd.n6884 gnd.n720 0.152939
R13378 gnd.n6885 gnd.n6884 0.152939
R13379 gnd.n6886 gnd.n6885 0.152939
R13380 gnd.n6886 gnd.n714 0.152939
R13381 gnd.n6894 gnd.n714 0.152939
R13382 gnd.n6895 gnd.n6894 0.152939
R13383 gnd.n6896 gnd.n6895 0.152939
R13384 gnd.n6896 gnd.n708 0.152939
R13385 gnd.n6904 gnd.n708 0.152939
R13386 gnd.n6905 gnd.n6904 0.152939
R13387 gnd.n6906 gnd.n6905 0.152939
R13388 gnd.n6906 gnd.n702 0.152939
R13389 gnd.n6914 gnd.n702 0.152939
R13390 gnd.n6915 gnd.n6914 0.152939
R13391 gnd.n6916 gnd.n6915 0.152939
R13392 gnd.n6916 gnd.n696 0.152939
R13393 gnd.n6924 gnd.n696 0.152939
R13394 gnd.n6925 gnd.n6924 0.152939
R13395 gnd.n6926 gnd.n6925 0.152939
R13396 gnd.n6926 gnd.n690 0.152939
R13397 gnd.n6934 gnd.n690 0.152939
R13398 gnd.n6935 gnd.n6934 0.152939
R13399 gnd.n6936 gnd.n6935 0.152939
R13400 gnd.n6936 gnd.n684 0.152939
R13401 gnd.n6944 gnd.n684 0.152939
R13402 gnd.n6945 gnd.n6944 0.152939
R13403 gnd.n6946 gnd.n6945 0.152939
R13404 gnd.n6946 gnd.n678 0.152939
R13405 gnd.n6954 gnd.n678 0.152939
R13406 gnd.n6955 gnd.n6954 0.152939
R13407 gnd.n6956 gnd.n6955 0.152939
R13408 gnd.n6956 gnd.n672 0.152939
R13409 gnd.n6964 gnd.n672 0.152939
R13410 gnd.n6965 gnd.n6964 0.152939
R13411 gnd.n6966 gnd.n6965 0.152939
R13412 gnd.n6966 gnd.n666 0.152939
R13413 gnd.n6974 gnd.n666 0.152939
R13414 gnd.n6975 gnd.n6974 0.152939
R13415 gnd.n6976 gnd.n6975 0.152939
R13416 gnd.n6976 gnd.n660 0.152939
R13417 gnd.n6984 gnd.n660 0.152939
R13418 gnd.n6985 gnd.n6984 0.152939
R13419 gnd.n6986 gnd.n6985 0.152939
R13420 gnd.n6986 gnd.n654 0.152939
R13421 gnd.n6994 gnd.n654 0.152939
R13422 gnd.n6995 gnd.n6994 0.152939
R13423 gnd.n6996 gnd.n6995 0.152939
R13424 gnd.n6996 gnd.n648 0.152939
R13425 gnd.n7004 gnd.n648 0.152939
R13426 gnd.n7005 gnd.n7004 0.152939
R13427 gnd.n7006 gnd.n7005 0.152939
R13428 gnd.n7006 gnd.n642 0.152939
R13429 gnd.n7014 gnd.n642 0.152939
R13430 gnd.n7015 gnd.n7014 0.152939
R13431 gnd.n7016 gnd.n7015 0.152939
R13432 gnd.n7016 gnd.n636 0.152939
R13433 gnd.n7024 gnd.n636 0.152939
R13434 gnd.n7025 gnd.n7024 0.152939
R13435 gnd.n7026 gnd.n7025 0.152939
R13436 gnd.n7026 gnd.n630 0.152939
R13437 gnd.n7034 gnd.n630 0.152939
R13438 gnd.n7035 gnd.n7034 0.152939
R13439 gnd.n7036 gnd.n7035 0.152939
R13440 gnd.n7036 gnd.n624 0.152939
R13441 gnd.n7044 gnd.n624 0.152939
R13442 gnd.n7045 gnd.n7044 0.152939
R13443 gnd.n7046 gnd.n7045 0.152939
R13444 gnd.n7046 gnd.n618 0.152939
R13445 gnd.n7054 gnd.n618 0.152939
R13446 gnd.n7055 gnd.n7054 0.152939
R13447 gnd.n7056 gnd.n7055 0.152939
R13448 gnd.n7056 gnd.n612 0.152939
R13449 gnd.n7064 gnd.n612 0.152939
R13450 gnd.n7065 gnd.n7064 0.152939
R13451 gnd.n7066 gnd.n7065 0.152939
R13452 gnd.n7066 gnd.n606 0.152939
R13453 gnd.n7074 gnd.n606 0.152939
R13454 gnd.n7075 gnd.n7074 0.152939
R13455 gnd.n7076 gnd.n7075 0.152939
R13456 gnd.n7076 gnd.n600 0.152939
R13457 gnd.n7084 gnd.n600 0.152939
R13458 gnd.n7085 gnd.n7084 0.152939
R13459 gnd.n7086 gnd.n7085 0.152939
R13460 gnd.n7086 gnd.n594 0.152939
R13461 gnd.n7094 gnd.n594 0.152939
R13462 gnd.n7095 gnd.n7094 0.152939
R13463 gnd.n7096 gnd.n7095 0.152939
R13464 gnd.n7096 gnd.n588 0.152939
R13465 gnd.n7104 gnd.n588 0.152939
R13466 gnd.n7105 gnd.n7104 0.152939
R13467 gnd.n7106 gnd.n7105 0.152939
R13468 gnd.n7106 gnd.n582 0.152939
R13469 gnd.n7114 gnd.n582 0.152939
R13470 gnd.n7115 gnd.n7114 0.152939
R13471 gnd.n7116 gnd.n7115 0.152939
R13472 gnd.n7116 gnd.n576 0.152939
R13473 gnd.n7124 gnd.n576 0.152939
R13474 gnd.n7125 gnd.n7124 0.152939
R13475 gnd.n7126 gnd.n7125 0.152939
R13476 gnd.n7126 gnd.n570 0.152939
R13477 gnd.n7134 gnd.n570 0.152939
R13478 gnd.n7135 gnd.n7134 0.152939
R13479 gnd.n7136 gnd.n7135 0.152939
R13480 gnd.n7136 gnd.n564 0.152939
R13481 gnd.n7144 gnd.n564 0.152939
R13482 gnd.n7145 gnd.n7144 0.152939
R13483 gnd.n7146 gnd.n7145 0.152939
R13484 gnd.n7146 gnd.n558 0.152939
R13485 gnd.n7154 gnd.n558 0.152939
R13486 gnd.n7155 gnd.n7154 0.152939
R13487 gnd.n7156 gnd.n7155 0.152939
R13488 gnd.n7156 gnd.n552 0.152939
R13489 gnd.n7164 gnd.n552 0.152939
R13490 gnd.n7165 gnd.n7164 0.152939
R13491 gnd.n7166 gnd.n7165 0.152939
R13492 gnd.n7166 gnd.n546 0.152939
R13493 gnd.n7174 gnd.n546 0.152939
R13494 gnd.n7175 gnd.n7174 0.152939
R13495 gnd.n7176 gnd.n7175 0.152939
R13496 gnd.n7176 gnd.n540 0.152939
R13497 gnd.n7184 gnd.n540 0.152939
R13498 gnd.n7185 gnd.n7184 0.152939
R13499 gnd.n7186 gnd.n7185 0.152939
R13500 gnd.n7186 gnd.n534 0.152939
R13501 gnd.n7194 gnd.n534 0.152939
R13502 gnd.n7195 gnd.n7194 0.152939
R13503 gnd.n7196 gnd.n7195 0.152939
R13504 gnd.n7196 gnd.n528 0.152939
R13505 gnd.n7204 gnd.n528 0.152939
R13506 gnd.n7206 gnd.n7205 0.152939
R13507 gnd.n7206 gnd.n522 0.152939
R13508 gnd.n7214 gnd.n522 0.152939
R13509 gnd.n7215 gnd.n7214 0.152939
R13510 gnd.n7216 gnd.n7215 0.152939
R13511 gnd.n7216 gnd.n516 0.152939
R13512 gnd.n7224 gnd.n516 0.152939
R13513 gnd.n7225 gnd.n7224 0.152939
R13514 gnd.n7226 gnd.n7225 0.152939
R13515 gnd.n7226 gnd.n510 0.152939
R13516 gnd.n7234 gnd.n510 0.152939
R13517 gnd.n7235 gnd.n7234 0.152939
R13518 gnd.n7236 gnd.n7235 0.152939
R13519 gnd.n7236 gnd.n504 0.152939
R13520 gnd.n7244 gnd.n504 0.152939
R13521 gnd.n7245 gnd.n7244 0.152939
R13522 gnd.n7246 gnd.n7245 0.152939
R13523 gnd.n7246 gnd.n498 0.152939
R13524 gnd.n7254 gnd.n498 0.152939
R13525 gnd.n7255 gnd.n7254 0.152939
R13526 gnd.n7256 gnd.n7255 0.152939
R13527 gnd.n7256 gnd.n492 0.152939
R13528 gnd.n7264 gnd.n492 0.152939
R13529 gnd.n7265 gnd.n7264 0.152939
R13530 gnd.n7266 gnd.n7265 0.152939
R13531 gnd.n7266 gnd.n486 0.152939
R13532 gnd.n7274 gnd.n486 0.152939
R13533 gnd.n7275 gnd.n7274 0.152939
R13534 gnd.n7276 gnd.n7275 0.152939
R13535 gnd.n7276 gnd.n480 0.152939
R13536 gnd.n7284 gnd.n480 0.152939
R13537 gnd.n7285 gnd.n7284 0.152939
R13538 gnd.n7286 gnd.n7285 0.152939
R13539 gnd.n7286 gnd.n474 0.152939
R13540 gnd.n7294 gnd.n474 0.152939
R13541 gnd.n7295 gnd.n7294 0.152939
R13542 gnd.n7296 gnd.n7295 0.152939
R13543 gnd.n7296 gnd.n468 0.152939
R13544 gnd.n7304 gnd.n468 0.152939
R13545 gnd.n7305 gnd.n7304 0.152939
R13546 gnd.n7306 gnd.n7305 0.152939
R13547 gnd.n7306 gnd.n462 0.152939
R13548 gnd.n7314 gnd.n462 0.152939
R13549 gnd.n7315 gnd.n7314 0.152939
R13550 gnd.n7316 gnd.n7315 0.152939
R13551 gnd.n7316 gnd.n456 0.152939
R13552 gnd.n7324 gnd.n456 0.152939
R13553 gnd.n7325 gnd.n7324 0.152939
R13554 gnd.n7326 gnd.n7325 0.152939
R13555 gnd.n7326 gnd.n450 0.152939
R13556 gnd.n7334 gnd.n450 0.152939
R13557 gnd.n7335 gnd.n7334 0.152939
R13558 gnd.n7336 gnd.n7335 0.152939
R13559 gnd.n7336 gnd.n444 0.152939
R13560 gnd.n7344 gnd.n444 0.152939
R13561 gnd.n7345 gnd.n7344 0.152939
R13562 gnd.n7346 gnd.n7345 0.152939
R13563 gnd.n7346 gnd.n438 0.152939
R13564 gnd.n7354 gnd.n438 0.152939
R13565 gnd.n7355 gnd.n7354 0.152939
R13566 gnd.n7356 gnd.n7355 0.152939
R13567 gnd.n7356 gnd.n432 0.152939
R13568 gnd.n7364 gnd.n432 0.152939
R13569 gnd.n7365 gnd.n7364 0.152939
R13570 gnd.n7366 gnd.n7365 0.152939
R13571 gnd.n7366 gnd.n426 0.152939
R13572 gnd.n7374 gnd.n426 0.152939
R13573 gnd.n7375 gnd.n7374 0.152939
R13574 gnd.n7376 gnd.n7375 0.152939
R13575 gnd.n7376 gnd.n420 0.152939
R13576 gnd.n7384 gnd.n420 0.152939
R13577 gnd.n7385 gnd.n7384 0.152939
R13578 gnd.n7386 gnd.n7385 0.152939
R13579 gnd.n7386 gnd.n414 0.152939
R13580 gnd.n7394 gnd.n414 0.152939
R13581 gnd.n7395 gnd.n7394 0.152939
R13582 gnd.n7396 gnd.n7395 0.152939
R13583 gnd.n7396 gnd.n408 0.152939
R13584 gnd.n7404 gnd.n408 0.152939
R13585 gnd.n7405 gnd.n7404 0.152939
R13586 gnd.n7406 gnd.n7405 0.152939
R13587 gnd.n7407 gnd.n7406 0.152939
R13588 gnd.n7407 gnd.n402 0.152939
R13589 gnd.n7417 gnd.n402 0.152939
R13590 gnd.n388 gnd.n385 0.152939
R13591 gnd.n389 gnd.n388 0.152939
R13592 gnd.n390 gnd.n389 0.152939
R13593 gnd.n391 gnd.n390 0.152939
R13594 gnd.n394 gnd.n391 0.152939
R13595 gnd.n395 gnd.n394 0.152939
R13596 gnd.n396 gnd.n395 0.152939
R13597 gnd.n397 gnd.n396 0.152939
R13598 gnd.n400 gnd.n397 0.152939
R13599 gnd.n401 gnd.n400 0.152939
R13600 gnd.n7418 gnd.n401 0.152939
R13601 gnd.n118 gnd.n93 0.152939
R13602 gnd.n119 gnd.n118 0.152939
R13603 gnd.n120 gnd.n119 0.152939
R13604 gnd.n137 gnd.n120 0.152939
R13605 gnd.n138 gnd.n137 0.152939
R13606 gnd.n139 gnd.n138 0.152939
R13607 gnd.n140 gnd.n139 0.152939
R13608 gnd.n157 gnd.n140 0.152939
R13609 gnd.n158 gnd.n157 0.152939
R13610 gnd.n159 gnd.n158 0.152939
R13611 gnd.n160 gnd.n159 0.152939
R13612 gnd.n177 gnd.n160 0.152939
R13613 gnd.n178 gnd.n177 0.152939
R13614 gnd.n179 gnd.n178 0.152939
R13615 gnd.n180 gnd.n179 0.152939
R13616 gnd.n196 gnd.n180 0.152939
R13617 gnd.n197 gnd.n196 0.152939
R13618 gnd.n198 gnd.n197 0.152939
R13619 gnd.n199 gnd.n198 0.152939
R13620 gnd.n214 gnd.n199 0.152939
R13621 gnd.n7672 gnd.n214 0.152939
R13622 gnd.n7753 gnd.n80 0.152939
R13623 gnd.n7442 gnd.n80 0.152939
R13624 gnd.n7443 gnd.n7442 0.152939
R13625 gnd.n7443 gnd.n376 0.152939
R13626 gnd.n7455 gnd.n376 0.152939
R13627 gnd.n7456 gnd.n7455 0.152939
R13628 gnd.n7457 gnd.n7456 0.152939
R13629 gnd.n7457 gnd.n369 0.152939
R13630 gnd.n7469 gnd.n369 0.152939
R13631 gnd.n7470 gnd.n7469 0.152939
R13632 gnd.n7471 gnd.n7470 0.152939
R13633 gnd.n7471 gnd.n364 0.152939
R13634 gnd.n7483 gnd.n364 0.152939
R13635 gnd.n7484 gnd.n7483 0.152939
R13636 gnd.n7486 gnd.n7484 0.152939
R13637 gnd.n7486 gnd.n7485 0.152939
R13638 gnd.n7485 gnd.n358 0.152939
R13639 gnd.n7514 gnd.n358 0.152939
R13640 gnd.n7515 gnd.n7514 0.152939
R13641 gnd.n7516 gnd.n7515 0.152939
R13642 gnd.n7516 gnd.n355 0.152939
R13643 gnd.n7521 gnd.n355 0.152939
R13644 gnd.n7522 gnd.n7521 0.152939
R13645 gnd.n7523 gnd.n7522 0.152939
R13646 gnd.n7523 gnd.n352 0.152939
R13647 gnd.n7528 gnd.n352 0.152939
R13648 gnd.n7561 gnd.n318 0.152939
R13649 gnd.n320 gnd.n318 0.152939
R13650 gnd.n324 gnd.n320 0.152939
R13651 gnd.n325 gnd.n324 0.152939
R13652 gnd.n326 gnd.n325 0.152939
R13653 gnd.n327 gnd.n326 0.152939
R13654 gnd.n331 gnd.n327 0.152939
R13655 gnd.n332 gnd.n331 0.152939
R13656 gnd.n333 gnd.n332 0.152939
R13657 gnd.n334 gnd.n333 0.152939
R13658 gnd.n338 gnd.n334 0.152939
R13659 gnd.n339 gnd.n338 0.152939
R13660 gnd.n340 gnd.n339 0.152939
R13661 gnd.n341 gnd.n340 0.152939
R13662 gnd.n345 gnd.n341 0.152939
R13663 gnd.n346 gnd.n345 0.152939
R13664 gnd.n7530 gnd.n346 0.152939
R13665 gnd.n7530 gnd.n7529 0.152939
R13666 gnd.n7671 gnd.n215 0.152939
R13667 gnd.n217 gnd.n215 0.152939
R13668 gnd.n221 gnd.n217 0.152939
R13669 gnd.n222 gnd.n221 0.152939
R13670 gnd.n223 gnd.n222 0.152939
R13671 gnd.n224 gnd.n223 0.152939
R13672 gnd.n228 gnd.n224 0.152939
R13673 gnd.n229 gnd.n228 0.152939
R13674 gnd.n230 gnd.n229 0.152939
R13675 gnd.n231 gnd.n230 0.152939
R13676 gnd.n235 gnd.n231 0.152939
R13677 gnd.n236 gnd.n235 0.152939
R13678 gnd.n237 gnd.n236 0.152939
R13679 gnd.n238 gnd.n237 0.152939
R13680 gnd.n242 gnd.n238 0.152939
R13681 gnd.n243 gnd.n242 0.152939
R13682 gnd.n244 gnd.n243 0.152939
R13683 gnd.n245 gnd.n244 0.152939
R13684 gnd.n249 gnd.n245 0.152939
R13685 gnd.n250 gnd.n249 0.152939
R13686 gnd.n251 gnd.n250 0.152939
R13687 gnd.n252 gnd.n251 0.152939
R13688 gnd.n256 gnd.n252 0.152939
R13689 gnd.n257 gnd.n256 0.152939
R13690 gnd.n258 gnd.n257 0.152939
R13691 gnd.n259 gnd.n258 0.152939
R13692 gnd.n263 gnd.n259 0.152939
R13693 gnd.n264 gnd.n263 0.152939
R13694 gnd.n265 gnd.n264 0.152939
R13695 gnd.n266 gnd.n265 0.152939
R13696 gnd.n270 gnd.n266 0.152939
R13697 gnd.n271 gnd.n270 0.152939
R13698 gnd.n272 gnd.n271 0.152939
R13699 gnd.n273 gnd.n272 0.152939
R13700 gnd.n277 gnd.n273 0.152939
R13701 gnd.n278 gnd.n277 0.152939
R13702 gnd.n7602 gnd.n278 0.152939
R13703 gnd.n7602 gnd.n7601 0.152939
R13704 gnd.n7601 gnd.n7600 0.152939
R13705 gnd.n7600 gnd.n282 0.152939
R13706 gnd.n288 gnd.n282 0.152939
R13707 gnd.n289 gnd.n288 0.152939
R13708 gnd.n290 gnd.n289 0.152939
R13709 gnd.n291 gnd.n290 0.152939
R13710 gnd.n295 gnd.n291 0.152939
R13711 gnd.n296 gnd.n295 0.152939
R13712 gnd.n297 gnd.n296 0.152939
R13713 gnd.n298 gnd.n297 0.152939
R13714 gnd.n302 gnd.n298 0.152939
R13715 gnd.n303 gnd.n302 0.152939
R13716 gnd.n304 gnd.n303 0.152939
R13717 gnd.n305 gnd.n304 0.152939
R13718 gnd.n309 gnd.n305 0.152939
R13719 gnd.n310 gnd.n309 0.152939
R13720 gnd.n311 gnd.n310 0.152939
R13721 gnd.n312 gnd.n311 0.152939
R13722 gnd.n317 gnd.n312 0.152939
R13723 gnd.n7563 gnd.n317 0.152939
R13724 gnd.n4277 gnd.n4276 0.152939
R13725 gnd.n4277 gnd.n4273 0.152939
R13726 gnd.n4285 gnd.n4273 0.152939
R13727 gnd.n4286 gnd.n4285 0.152939
R13728 gnd.n4287 gnd.n4286 0.152939
R13729 gnd.n4287 gnd.n4269 0.152939
R13730 gnd.n4295 gnd.n4269 0.152939
R13731 gnd.n4296 gnd.n4295 0.152939
R13732 gnd.n4297 gnd.n4296 0.152939
R13733 gnd.n4297 gnd.n4265 0.152939
R13734 gnd.n4305 gnd.n4265 0.152939
R13735 gnd.n4306 gnd.n4305 0.152939
R13736 gnd.n4307 gnd.n4306 0.152939
R13737 gnd.n4307 gnd.n4261 0.152939
R13738 gnd.n4315 gnd.n4261 0.152939
R13739 gnd.n4316 gnd.n4315 0.152939
R13740 gnd.n4317 gnd.n4316 0.152939
R13741 gnd.n4317 gnd.n4257 0.152939
R13742 gnd.n4328 gnd.n4257 0.152939
R13743 gnd.n4329 gnd.n4328 0.152939
R13744 gnd.n4330 gnd.n4329 0.152939
R13745 gnd.n4330 gnd.n4253 0.152939
R13746 gnd.n4338 gnd.n4253 0.152939
R13747 gnd.n4339 gnd.n4338 0.152939
R13748 gnd.n4341 gnd.n4339 0.152939
R13749 gnd.n4351 gnd.n1859 0.152939
R13750 gnd.n4352 gnd.n4351 0.152939
R13751 gnd.n4353 gnd.n4352 0.152939
R13752 gnd.n4353 gnd.n1855 0.152939
R13753 gnd.n4361 gnd.n1855 0.152939
R13754 gnd.n4362 gnd.n4361 0.152939
R13755 gnd.n4363 gnd.n4362 0.152939
R13756 gnd.n4363 gnd.n1851 0.152939
R13757 gnd.n4373 gnd.n1851 0.152939
R13758 gnd.n4374 gnd.n4373 0.152939
R13759 gnd.n4375 gnd.n4374 0.152939
R13760 gnd.n4375 gnd.n1847 0.152939
R13761 gnd.n4383 gnd.n1847 0.152939
R13762 gnd.n4384 gnd.n4383 0.152939
R13763 gnd.n4385 gnd.n4384 0.152939
R13764 gnd.n4385 gnd.n1843 0.152939
R13765 gnd.n4393 gnd.n1843 0.152939
R13766 gnd.n4394 gnd.n4393 0.152939
R13767 gnd.n4395 gnd.n4394 0.152939
R13768 gnd.n4395 gnd.n1839 0.152939
R13769 gnd.n4403 gnd.n1839 0.152939
R13770 gnd.n4404 gnd.n4403 0.152939
R13771 gnd.n4405 gnd.n4404 0.152939
R13772 gnd.n4405 gnd.n1835 0.152939
R13773 gnd.n4413 gnd.n1835 0.152939
R13774 gnd.n4414 gnd.n4413 0.152939
R13775 gnd.n4416 gnd.n4414 0.152939
R13776 gnd.n4416 gnd.n4415 0.152939
R13777 gnd.n4415 gnd.n1828 0.152939
R13778 gnd.n4425 gnd.n1828 0.152939
R13779 gnd.n1626 gnd.n1625 0.152939
R13780 gnd.n1627 gnd.n1626 0.152939
R13781 gnd.n1647 gnd.n1627 0.152939
R13782 gnd.n1648 gnd.n1647 0.152939
R13783 gnd.n1649 gnd.n1648 0.152939
R13784 gnd.n1650 gnd.n1649 0.152939
R13785 gnd.n1667 gnd.n1650 0.152939
R13786 gnd.n1668 gnd.n1667 0.152939
R13787 gnd.n1669 gnd.n1668 0.152939
R13788 gnd.n1670 gnd.n1669 0.152939
R13789 gnd.n1687 gnd.n1670 0.152939
R13790 gnd.n1688 gnd.n1687 0.152939
R13791 gnd.n1689 gnd.n1688 0.152939
R13792 gnd.n1690 gnd.n1689 0.152939
R13793 gnd.n1707 gnd.n1690 0.152939
R13794 gnd.n1708 gnd.n1707 0.152939
R13795 gnd.n1709 gnd.n1708 0.152939
R13796 gnd.n1710 gnd.n1709 0.152939
R13797 gnd.n1727 gnd.n1710 0.152939
R13798 gnd.n1728 gnd.n1727 0.152939
R13799 gnd.n1728 gnd.n94 0.152939
R13800 gnd.n2809 gnd.n2808 0.152939
R13801 gnd.n2810 gnd.n2809 0.152939
R13802 gnd.n2810 gnd.n2452 0.152939
R13803 gnd.n2816 gnd.n2452 0.152939
R13804 gnd.n2817 gnd.n2816 0.152939
R13805 gnd.n2818 gnd.n2817 0.152939
R13806 gnd.n2819 gnd.n2818 0.152939
R13807 gnd.n2820 gnd.n2819 0.152939
R13808 gnd.n2823 gnd.n2820 0.152939
R13809 gnd.n2824 gnd.n2823 0.152939
R13810 gnd.n2825 gnd.n2824 0.152939
R13811 gnd.n2826 gnd.n2825 0.152939
R13812 gnd.n2827 gnd.n2826 0.152939
R13813 gnd.n2827 gnd.n2427 0.152939
R13814 gnd.n2903 gnd.n2427 0.152939
R13815 gnd.n2904 gnd.n2903 0.152939
R13816 gnd.n2905 gnd.n2904 0.152939
R13817 gnd.n2905 gnd.n2423 0.152939
R13818 gnd.n2911 gnd.n2423 0.152939
R13819 gnd.n2912 gnd.n2911 0.152939
R13820 gnd.n2913 gnd.n2912 0.152939
R13821 gnd.n2913 gnd.n2419 0.152939
R13822 gnd.n2921 gnd.n2419 0.152939
R13823 gnd.n2922 gnd.n2921 0.152939
R13824 gnd.n2923 gnd.n2922 0.152939
R13825 gnd.n2923 gnd.n2394 0.152939
R13826 gnd.n3205 gnd.n2394 0.152939
R13827 gnd.n3206 gnd.n3205 0.152939
R13828 gnd.n3207 gnd.n3206 0.152939
R13829 gnd.n3208 gnd.n3207 0.152939
R13830 gnd.n3208 gnd.n2369 0.152939
R13831 gnd.n3237 gnd.n2369 0.152939
R13832 gnd.n3238 gnd.n3237 0.152939
R13833 gnd.n3239 gnd.n3238 0.152939
R13834 gnd.n3241 gnd.n3239 0.152939
R13835 gnd.n3241 gnd.n3240 0.152939
R13836 gnd.n3240 gnd.n1497 0.152939
R13837 gnd.n1498 gnd.n1497 0.152939
R13838 gnd.n1499 gnd.n1498 0.152939
R13839 gnd.n3277 gnd.n1499 0.152939
R13840 gnd.n3278 gnd.n3277 0.152939
R13841 gnd.n3278 gnd.n2243 0.152939
R13842 gnd.n3319 gnd.n2243 0.152939
R13843 gnd.n3320 gnd.n3319 0.152939
R13844 gnd.n3321 gnd.n3320 0.152939
R13845 gnd.n3321 gnd.n2225 0.152939
R13846 gnd.n3361 gnd.n2225 0.152939
R13847 gnd.n3362 gnd.n3361 0.152939
R13848 gnd.n3363 gnd.n3362 0.152939
R13849 gnd.n3364 gnd.n3363 0.152939
R13850 gnd.n3364 gnd.n2199 0.152939
R13851 gnd.n3423 gnd.n2199 0.152939
R13852 gnd.n3424 gnd.n3423 0.152939
R13853 gnd.n3425 gnd.n3424 0.152939
R13854 gnd.n3425 gnd.n2181 0.152939
R13855 gnd.n3451 gnd.n2181 0.152939
R13856 gnd.n3452 gnd.n3451 0.152939
R13857 gnd.n3453 gnd.n3452 0.152939
R13858 gnd.n3454 gnd.n3453 0.152939
R13859 gnd.n3454 gnd.n2148 0.152939
R13860 gnd.n3501 gnd.n2148 0.152939
R13861 gnd.n3502 gnd.n3501 0.152939
R13862 gnd.n3503 gnd.n3502 0.152939
R13863 gnd.n3503 gnd.n2125 0.152939
R13864 gnd.n3541 gnd.n2125 0.152939
R13865 gnd.n3542 gnd.n3541 0.152939
R13866 gnd.n3543 gnd.n3542 0.152939
R13867 gnd.n3543 gnd.n2103 0.152939
R13868 gnd.n3598 gnd.n2103 0.152939
R13869 gnd.n3599 gnd.n3598 0.152939
R13870 gnd.n3600 gnd.n3599 0.152939
R13871 gnd.n3600 gnd.n2083 0.152939
R13872 gnd.n3623 gnd.n2083 0.152939
R13873 gnd.n3624 gnd.n3623 0.152939
R13874 gnd.n3625 gnd.n3624 0.152939
R13875 gnd.n3625 gnd.n2063 0.152939
R13876 gnd.n3683 gnd.n2063 0.152939
R13877 gnd.n3684 gnd.n3683 0.152939
R13878 gnd.n3685 gnd.n3684 0.152939
R13879 gnd.n3685 gnd.n2041 0.152939
R13880 gnd.n3712 gnd.n2041 0.152939
R13881 gnd.n3713 gnd.n3712 0.152939
R13882 gnd.n3714 gnd.n3713 0.152939
R13883 gnd.n3715 gnd.n3714 0.152939
R13884 gnd.n3715 gnd.n2013 0.152939
R13885 gnd.n3763 gnd.n2013 0.152939
R13886 gnd.n3764 gnd.n3763 0.152939
R13887 gnd.n3765 gnd.n3764 0.152939
R13888 gnd.n3765 gnd.n1993 0.152939
R13889 gnd.n3789 gnd.n1993 0.152939
R13890 gnd.n3790 gnd.n3789 0.152939
R13891 gnd.n3791 gnd.n3790 0.152939
R13892 gnd.n3792 gnd.n3791 0.152939
R13893 gnd.n3792 gnd.n1963 0.152939
R13894 gnd.n3833 gnd.n1963 0.152939
R13895 gnd.n3834 gnd.n3833 0.152939
R13896 gnd.n3835 gnd.n3834 0.152939
R13897 gnd.n3837 gnd.n3835 0.152939
R13898 gnd.n3837 gnd.n3836 0.152939
R13899 gnd.n3836 gnd.n1914 0.152939
R13900 gnd.n1915 gnd.n1914 0.152939
R13901 gnd.n1916 gnd.n1915 0.152939
R13902 gnd.n1925 gnd.n1916 0.152939
R13903 gnd.n1926 gnd.n1925 0.152939
R13904 gnd.n1927 gnd.n1926 0.152939
R13905 gnd.n1928 gnd.n1927 0.152939
R13906 gnd.n1929 gnd.n1928 0.152939
R13907 gnd.n1931 gnd.n1929 0.152939
R13908 gnd.n1931 gnd.n1930 0.152939
R13909 gnd.n1930 gnd.n1604 0.152939
R13910 gnd.n1605 gnd.n1604 0.152939
R13911 gnd.n1606 gnd.n1605 0.152939
R13912 gnd.n1612 gnd.n1606 0.152939
R13913 gnd.n1613 gnd.n1612 0.152939
R13914 gnd.n1614 gnd.n1613 0.152939
R13915 gnd.n1615 gnd.n1614 0.152939
R13916 gnd.n1795 gnd.n1615 0.152939
R13917 gnd.n1796 gnd.n1795 0.152939
R13918 gnd.n1797 gnd.n1796 0.152939
R13919 gnd.n1797 gnd.n1791 0.152939
R13920 gnd.n1803 gnd.n1791 0.152939
R13921 gnd.n1804 gnd.n1803 0.152939
R13922 gnd.n1805 gnd.n1804 0.152939
R13923 gnd.n1806 gnd.n1805 0.152939
R13924 gnd.n1807 gnd.n1806 0.152939
R13925 gnd.n1808 gnd.n1807 0.152939
R13926 gnd.n1810 gnd.n1808 0.152939
R13927 gnd.n1810 gnd.n1809 0.152939
R13928 gnd.n1809 gnd.n1770 0.152939
R13929 gnd.n4498 gnd.n1770 0.152939
R13930 gnd.n4499 gnd.n4498 0.152939
R13931 gnd.n4500 gnd.n4499 0.152939
R13932 gnd.n4500 gnd.n1766 0.152939
R13933 gnd.n4506 gnd.n1766 0.152939
R13934 gnd.n4507 gnd.n4506 0.152939
R13935 gnd.n4508 gnd.n4507 0.152939
R13936 gnd.n4509 gnd.n4508 0.152939
R13937 gnd.n2609 gnd.n2608 0.152939
R13938 gnd.n2610 gnd.n2609 0.152939
R13939 gnd.n2610 gnd.n2546 0.152939
R13940 gnd.n2616 gnd.n2546 0.152939
R13941 gnd.n2617 gnd.n2616 0.152939
R13942 gnd.n2618 gnd.n2617 0.152939
R13943 gnd.n2618 gnd.n2544 0.152939
R13944 gnd.n2624 gnd.n2544 0.152939
R13945 gnd.n2625 gnd.n2624 0.152939
R13946 gnd.n2626 gnd.n2625 0.152939
R13947 gnd.n2626 gnd.n2527 0.152939
R13948 gnd.n2638 gnd.n2527 0.152939
R13949 gnd.n2639 gnd.n2638 0.152939
R13950 gnd.n2640 gnd.n2639 0.152939
R13951 gnd.n2640 gnd.n2522 0.152939
R13952 gnd.n2691 gnd.n2522 0.152939
R13953 gnd.n2692 gnd.n2691 0.152939
R13954 gnd.n2694 gnd.n2692 0.152939
R13955 gnd.n2694 gnd.n2693 0.152939
R13956 gnd.n2693 gnd.n2518 0.152939
R13957 gnd.n2518 gnd.n2516 0.152939
R13958 gnd.n2710 gnd.n2516 0.152939
R13959 gnd.n2711 gnd.n2710 0.152939
R13960 gnd.n2712 gnd.n2711 0.152939
R13961 gnd.n2712 gnd.n2480 0.152939
R13962 gnd.n2755 gnd.n2480 0.152939
R13963 gnd.n2561 gnd.n1136 0.152939
R13964 gnd.n2569 gnd.n2561 0.152939
R13965 gnd.n2570 gnd.n2569 0.152939
R13966 gnd.n2571 gnd.n2570 0.152939
R13967 gnd.n2571 gnd.n2559 0.152939
R13968 gnd.n2579 gnd.n2559 0.152939
R13969 gnd.n2580 gnd.n2579 0.152939
R13970 gnd.n2581 gnd.n2580 0.152939
R13971 gnd.n2581 gnd.n2557 0.152939
R13972 gnd.n2589 gnd.n2557 0.152939
R13973 gnd.n2590 gnd.n2589 0.152939
R13974 gnd.n2591 gnd.n2590 0.152939
R13975 gnd.n2591 gnd.n2555 0.152939
R13976 gnd.n2599 gnd.n2555 0.152939
R13977 gnd.n2600 gnd.n2599 0.152939
R13978 gnd.n2601 gnd.n2600 0.152939
R13979 gnd.n2601 gnd.n2548 0.152939
R13980 gnd.n2605 gnd.n2548 0.152939
R13981 gnd.n1278 gnd.n1253 0.152939
R13982 gnd.n1279 gnd.n1278 0.152939
R13983 gnd.n1280 gnd.n1279 0.152939
R13984 gnd.n1298 gnd.n1280 0.152939
R13985 gnd.n1299 gnd.n1298 0.152939
R13986 gnd.n1300 gnd.n1299 0.152939
R13987 gnd.n1301 gnd.n1300 0.152939
R13988 gnd.n1317 gnd.n1301 0.152939
R13989 gnd.n1318 gnd.n1317 0.152939
R13990 gnd.n1319 gnd.n1318 0.152939
R13991 gnd.n1320 gnd.n1319 0.152939
R13992 gnd.n1338 gnd.n1320 0.152939
R13993 gnd.n1339 gnd.n1338 0.152939
R13994 gnd.n1340 gnd.n1339 0.152939
R13995 gnd.n1341 gnd.n1340 0.152939
R13996 gnd.n1358 gnd.n1341 0.152939
R13997 gnd.n1359 gnd.n1358 0.152939
R13998 gnd.n1360 gnd.n1359 0.152939
R13999 gnd.n1361 gnd.n1360 0.152939
R14000 gnd.n1378 gnd.n1361 0.152939
R14001 gnd.n4903 gnd.n1378 0.152939
R14002 gnd.n4902 gnd.n1379 0.152939
R14003 gnd.n1384 gnd.n1379 0.152939
R14004 gnd.n1385 gnd.n1384 0.152939
R14005 gnd.n1386 gnd.n1385 0.152939
R14006 gnd.n1387 gnd.n1386 0.152939
R14007 gnd.n1388 gnd.n1387 0.152939
R14008 gnd.n1392 gnd.n1388 0.152939
R14009 gnd.n1393 gnd.n1392 0.152939
R14010 gnd.n1394 gnd.n1393 0.152939
R14011 gnd.n1395 gnd.n1394 0.152939
R14012 gnd.n1399 gnd.n1395 0.152939
R14013 gnd.n1400 gnd.n1399 0.152939
R14014 gnd.n1401 gnd.n1400 0.152939
R14015 gnd.n1402 gnd.n1401 0.152939
R14016 gnd.n1406 gnd.n1402 0.152939
R14017 gnd.n1407 gnd.n1406 0.152939
R14018 gnd.n1408 gnd.n1407 0.152939
R14019 gnd.n1411 gnd.n1408 0.152939
R14020 gnd.n1415 gnd.n1411 0.152939
R14021 gnd.n1416 gnd.n1415 0.152939
R14022 gnd.n1417 gnd.n1416 0.152939
R14023 gnd.n1418 gnd.n1417 0.152939
R14024 gnd.n1422 gnd.n1418 0.152939
R14025 gnd.n1423 gnd.n1422 0.152939
R14026 gnd.n1424 gnd.n1423 0.152939
R14027 gnd.n2981 gnd.n2980 0.152939
R14028 gnd.n2990 gnd.n2981 0.152939
R14029 gnd.n2991 gnd.n2990 0.152939
R14030 gnd.n2992 gnd.n2991 0.152939
R14031 gnd.n2992 gnd.n2976 0.152939
R14032 gnd.n3000 gnd.n2976 0.152939
R14033 gnd.n3001 gnd.n3000 0.152939
R14034 gnd.n3002 gnd.n3001 0.152939
R14035 gnd.n3002 gnd.n2970 0.152939
R14036 gnd.n3010 gnd.n2970 0.152939
R14037 gnd.n3011 gnd.n3010 0.152939
R14038 gnd.n3012 gnd.n3011 0.152939
R14039 gnd.n3012 gnd.n2966 0.152939
R14040 gnd.n3020 gnd.n2966 0.152939
R14041 gnd.n3021 gnd.n3020 0.152939
R14042 gnd.n3022 gnd.n3021 0.152939
R14043 gnd.n3022 gnd.n2962 0.152939
R14044 gnd.n3030 gnd.n2962 0.152939
R14045 gnd.n3031 gnd.n3030 0.152939
R14046 gnd.n3032 gnd.n3031 0.152939
R14047 gnd.n3032 gnd.n2958 0.152939
R14048 gnd.n3040 gnd.n2958 0.152939
R14049 gnd.n3041 gnd.n3040 0.152939
R14050 gnd.n3042 gnd.n3041 0.152939
R14051 gnd.n3042 gnd.n2954 0.152939
R14052 gnd.n3050 gnd.n2954 0.152939
R14053 gnd.n3051 gnd.n3050 0.152939
R14054 gnd.n3052 gnd.n3051 0.152939
R14055 gnd.n3052 gnd.n2948 0.152939
R14056 gnd.n3059 gnd.n2948 0.152939
R14057 gnd.n1073 gnd.n1072 0.152939
R14058 gnd.n1074 gnd.n1073 0.152939
R14059 gnd.n1075 gnd.n1074 0.152939
R14060 gnd.n1076 gnd.n1075 0.152939
R14061 gnd.n1077 gnd.n1076 0.152939
R14062 gnd.n1078 gnd.n1077 0.152939
R14063 gnd.n1079 gnd.n1078 0.152939
R14064 gnd.n1080 gnd.n1079 0.152939
R14065 gnd.n1081 gnd.n1080 0.152939
R14066 gnd.n1082 gnd.n1081 0.152939
R14067 gnd.n1083 gnd.n1082 0.152939
R14068 gnd.n1084 gnd.n1083 0.152939
R14069 gnd.n1085 gnd.n1084 0.152939
R14070 gnd.n1086 gnd.n1085 0.152939
R14071 gnd.n1087 gnd.n1086 0.152939
R14072 gnd.n1088 gnd.n1087 0.152939
R14073 gnd.n1089 gnd.n1088 0.152939
R14074 gnd.n1092 gnd.n1089 0.152939
R14075 gnd.n1093 gnd.n1092 0.152939
R14076 gnd.n1094 gnd.n1093 0.152939
R14077 gnd.n1095 gnd.n1094 0.152939
R14078 gnd.n1096 gnd.n1095 0.152939
R14079 gnd.n1097 gnd.n1096 0.152939
R14080 gnd.n1098 gnd.n1097 0.152939
R14081 gnd.n1099 gnd.n1098 0.152939
R14082 gnd.n1100 gnd.n1099 0.152939
R14083 gnd.n1101 gnd.n1100 0.152939
R14084 gnd.n1102 gnd.n1101 0.152939
R14085 gnd.n1103 gnd.n1102 0.152939
R14086 gnd.n1104 gnd.n1103 0.152939
R14087 gnd.n1105 gnd.n1104 0.152939
R14088 gnd.n1106 gnd.n1105 0.152939
R14089 gnd.n1107 gnd.n1106 0.152939
R14090 gnd.n1108 gnd.n1107 0.152939
R14091 gnd.n1109 gnd.n1108 0.152939
R14092 gnd.n1110 gnd.n1109 0.152939
R14093 gnd.n1111 gnd.n1110 0.152939
R14094 gnd.n1114 gnd.n1111 0.152939
R14095 gnd.n1115 gnd.n1114 0.152939
R14096 gnd.n1116 gnd.n1115 0.152939
R14097 gnd.n1117 gnd.n1116 0.152939
R14098 gnd.n1118 gnd.n1117 0.152939
R14099 gnd.n1119 gnd.n1118 0.152939
R14100 gnd.n1120 gnd.n1119 0.152939
R14101 gnd.n1121 gnd.n1120 0.152939
R14102 gnd.n1122 gnd.n1121 0.152939
R14103 gnd.n1123 gnd.n1122 0.152939
R14104 gnd.n1124 gnd.n1123 0.152939
R14105 gnd.n1125 gnd.n1124 0.152939
R14106 gnd.n1126 gnd.n1125 0.152939
R14107 gnd.n1127 gnd.n1126 0.152939
R14108 gnd.n1128 gnd.n1127 0.152939
R14109 gnd.n1129 gnd.n1128 0.152939
R14110 gnd.n1130 gnd.n1129 0.152939
R14111 gnd.n1131 gnd.n1130 0.152939
R14112 gnd.n1132 gnd.n1131 0.152939
R14113 gnd.n5047 gnd.n1132 0.152939
R14114 gnd.n5047 gnd.n5046 0.152939
R14115 gnd.n1147 gnd.n1146 0.152939
R14116 gnd.n1148 gnd.n1147 0.152939
R14117 gnd.n1149 gnd.n1148 0.152939
R14118 gnd.n1169 gnd.n1149 0.152939
R14119 gnd.n1170 gnd.n1169 0.152939
R14120 gnd.n1171 gnd.n1170 0.152939
R14121 gnd.n1172 gnd.n1171 0.152939
R14122 gnd.n1188 gnd.n1172 0.152939
R14123 gnd.n1189 gnd.n1188 0.152939
R14124 gnd.n1190 gnd.n1189 0.152939
R14125 gnd.n1191 gnd.n1190 0.152939
R14126 gnd.n1209 gnd.n1191 0.152939
R14127 gnd.n1210 gnd.n1209 0.152939
R14128 gnd.n1211 gnd.n1210 0.152939
R14129 gnd.n1212 gnd.n1211 0.152939
R14130 gnd.n1229 gnd.n1212 0.152939
R14131 gnd.n1230 gnd.n1229 0.152939
R14132 gnd.n1231 gnd.n1230 0.152939
R14133 gnd.n1232 gnd.n1231 0.152939
R14134 gnd.n1250 gnd.n1232 0.152939
R14135 gnd.n1251 gnd.n1250 0.152939
R14136 gnd.n2652 gnd.n2646 0.152939
R14137 gnd.n2658 gnd.n2646 0.152939
R14138 gnd.n2659 gnd.n2658 0.152939
R14139 gnd.n2660 gnd.n2659 0.152939
R14140 gnd.n2661 gnd.n2660 0.152939
R14141 gnd.n2662 gnd.n2661 0.152939
R14142 gnd.n2665 gnd.n2662 0.152939
R14143 gnd.n2666 gnd.n2665 0.152939
R14144 gnd.n2667 gnd.n2666 0.152939
R14145 gnd.n2669 gnd.n2667 0.152939
R14146 gnd.n2669 gnd.n2668 0.152939
R14147 gnd.n804 gnd.n803 0.152939
R14148 gnd.n805 gnd.n804 0.152939
R14149 gnd.n810 gnd.n805 0.152939
R14150 gnd.n811 gnd.n810 0.152939
R14151 gnd.n812 gnd.n811 0.152939
R14152 gnd.n813 gnd.n812 0.152939
R14153 gnd.n818 gnd.n813 0.152939
R14154 gnd.n819 gnd.n818 0.152939
R14155 gnd.n820 gnd.n819 0.152939
R14156 gnd.n821 gnd.n820 0.152939
R14157 gnd.n826 gnd.n821 0.152939
R14158 gnd.n827 gnd.n826 0.152939
R14159 gnd.n828 gnd.n827 0.152939
R14160 gnd.n829 gnd.n828 0.152939
R14161 gnd.n834 gnd.n829 0.152939
R14162 gnd.n835 gnd.n834 0.152939
R14163 gnd.n836 gnd.n835 0.152939
R14164 gnd.n837 gnd.n836 0.152939
R14165 gnd.n842 gnd.n837 0.152939
R14166 gnd.n843 gnd.n842 0.152939
R14167 gnd.n844 gnd.n843 0.152939
R14168 gnd.n845 gnd.n844 0.152939
R14169 gnd.n850 gnd.n845 0.152939
R14170 gnd.n851 gnd.n850 0.152939
R14171 gnd.n852 gnd.n851 0.152939
R14172 gnd.n853 gnd.n852 0.152939
R14173 gnd.n858 gnd.n853 0.152939
R14174 gnd.n859 gnd.n858 0.152939
R14175 gnd.n860 gnd.n859 0.152939
R14176 gnd.n861 gnd.n860 0.152939
R14177 gnd.n866 gnd.n861 0.152939
R14178 gnd.n867 gnd.n866 0.152939
R14179 gnd.n868 gnd.n867 0.152939
R14180 gnd.n869 gnd.n868 0.152939
R14181 gnd.n874 gnd.n869 0.152939
R14182 gnd.n875 gnd.n874 0.152939
R14183 gnd.n876 gnd.n875 0.152939
R14184 gnd.n877 gnd.n876 0.152939
R14185 gnd.n882 gnd.n877 0.152939
R14186 gnd.n883 gnd.n882 0.152939
R14187 gnd.n884 gnd.n883 0.152939
R14188 gnd.n885 gnd.n884 0.152939
R14189 gnd.n890 gnd.n885 0.152939
R14190 gnd.n891 gnd.n890 0.152939
R14191 gnd.n892 gnd.n891 0.152939
R14192 gnd.n893 gnd.n892 0.152939
R14193 gnd.n898 gnd.n893 0.152939
R14194 gnd.n899 gnd.n898 0.152939
R14195 gnd.n900 gnd.n899 0.152939
R14196 gnd.n901 gnd.n900 0.152939
R14197 gnd.n906 gnd.n901 0.152939
R14198 gnd.n907 gnd.n906 0.152939
R14199 gnd.n908 gnd.n907 0.152939
R14200 gnd.n909 gnd.n908 0.152939
R14201 gnd.n914 gnd.n909 0.152939
R14202 gnd.n915 gnd.n914 0.152939
R14203 gnd.n916 gnd.n915 0.152939
R14204 gnd.n917 gnd.n916 0.152939
R14205 gnd.n922 gnd.n917 0.152939
R14206 gnd.n923 gnd.n922 0.152939
R14207 gnd.n924 gnd.n923 0.152939
R14208 gnd.n925 gnd.n924 0.152939
R14209 gnd.n930 gnd.n925 0.152939
R14210 gnd.n931 gnd.n930 0.152939
R14211 gnd.n932 gnd.n931 0.152939
R14212 gnd.n933 gnd.n932 0.152939
R14213 gnd.n938 gnd.n933 0.152939
R14214 gnd.n939 gnd.n938 0.152939
R14215 gnd.n940 gnd.n939 0.152939
R14216 gnd.n941 gnd.n940 0.152939
R14217 gnd.n946 gnd.n941 0.152939
R14218 gnd.n947 gnd.n946 0.152939
R14219 gnd.n948 gnd.n947 0.152939
R14220 gnd.n949 gnd.n948 0.152939
R14221 gnd.n954 gnd.n949 0.152939
R14222 gnd.n955 gnd.n954 0.152939
R14223 gnd.n956 gnd.n955 0.152939
R14224 gnd.n957 gnd.n956 0.152939
R14225 gnd.n962 gnd.n957 0.152939
R14226 gnd.n963 gnd.n962 0.152939
R14227 gnd.n964 gnd.n963 0.152939
R14228 gnd.n965 gnd.n964 0.152939
R14229 gnd.n2649 gnd.n965 0.152939
R14230 gnd.n2651 gnd.n2649 0.152939
R14231 gnd.n3198 gnd.n3197 0.152939
R14232 gnd.n3197 gnd.n2376 0.152939
R14233 gnd.n3225 gnd.n2376 0.152939
R14234 gnd.n3226 gnd.n3225 0.152939
R14235 gnd.n3230 gnd.n3226 0.152939
R14236 gnd.n3230 gnd.n3229 0.152939
R14237 gnd.n3229 gnd.n3228 0.152939
R14238 gnd.n3228 gnd.n2275 0.152939
R14239 gnd.n3262 gnd.n2275 0.152939
R14240 gnd.n3263 gnd.n3262 0.152939
R14241 gnd.n3265 gnd.n3263 0.152939
R14242 gnd.n3265 gnd.n3264 0.152939
R14243 gnd.n3264 gnd.n2264 0.152939
R14244 gnd.n3287 gnd.n2264 0.152939
R14245 gnd.n3288 gnd.n3287 0.152939
R14246 gnd.n3296 gnd.n3288 0.152939
R14247 gnd.n3296 gnd.n3295 0.152939
R14248 gnd.n3295 gnd.n3294 0.152939
R14249 gnd.n3294 gnd.n3289 0.152939
R14250 gnd.n3289 gnd.n2217 0.152939
R14251 gnd.n3373 gnd.n2217 0.152939
R14252 gnd.n3374 gnd.n3373 0.152939
R14253 gnd.n3394 gnd.n3374 0.152939
R14254 gnd.n3394 gnd.n3393 0.152939
R14255 gnd.n3393 gnd.n3392 0.152939
R14256 gnd.n3392 gnd.n3375 0.152939
R14257 gnd.n3388 gnd.n3375 0.152939
R14258 gnd.n3388 gnd.n3387 0.152939
R14259 gnd.n3387 gnd.n3386 0.152939
R14260 gnd.n3386 gnd.n3383 0.152939
R14261 gnd.n3383 gnd.n3382 0.152939
R14262 gnd.n3382 gnd.n2165 0.152939
R14263 gnd.n3475 gnd.n2165 0.152939
R14264 gnd.n3476 gnd.n3475 0.152939
R14265 gnd.n3477 gnd.n3476 0.152939
R14266 gnd.n3477 gnd.n2141 0.152939
R14267 gnd.n3523 gnd.n2141 0.152939
R14268 gnd.n3523 gnd.n3522 0.152939
R14269 gnd.n3522 gnd.n3521 0.152939
R14270 gnd.n3521 gnd.n2118 0.152939
R14271 gnd.n3582 gnd.n2118 0.152939
R14272 gnd.n3582 gnd.n3581 0.152939
R14273 gnd.n3581 gnd.n3580 0.152939
R14274 gnd.n3580 gnd.n2119 0.152939
R14275 gnd.n3576 gnd.n2119 0.152939
R14276 gnd.n3576 gnd.n3575 0.152939
R14277 gnd.n3575 gnd.n3574 0.152939
R14278 gnd.n3574 gnd.n3564 0.152939
R14279 gnd.n3570 gnd.n3564 0.152939
R14280 gnd.n3570 gnd.n2056 0.152939
R14281 gnd.n3692 gnd.n2056 0.152939
R14282 gnd.n3693 gnd.n3692 0.152939
R14283 gnd.n3695 gnd.n3693 0.152939
R14284 gnd.n3695 gnd.n3694 0.152939
R14285 gnd.n3694 gnd.n2027 0.152939
R14286 gnd.n3731 gnd.n2027 0.152939
R14287 gnd.n3732 gnd.n3731 0.152939
R14288 gnd.n3748 gnd.n3732 0.152939
R14289 gnd.n3748 gnd.n3747 0.152939
R14290 gnd.n3747 gnd.n3746 0.152939
R14291 gnd.n3746 gnd.n3733 0.152939
R14292 gnd.n3742 gnd.n3733 0.152939
R14293 gnd.n3742 gnd.n3741 0.152939
R14294 gnd.n3741 gnd.n3740 0.152939
R14295 gnd.n3740 gnd.n1971 0.152939
R14296 gnd.n3822 gnd.n1971 0.152939
R14297 gnd.n3823 gnd.n3822 0.152939
R14298 gnd.n3825 gnd.n3823 0.152939
R14299 gnd.n3825 gnd.n3824 0.152939
R14300 gnd.n3824 gnd.n1944 0.152939
R14301 gnd.n3864 gnd.n1944 0.152939
R14302 gnd.n3865 gnd.n3864 0.152939
R14303 gnd.n3866 gnd.n3865 0.152939
R14304 gnd.n3866 gnd.n1941 0.152939
R14305 gnd.n3875 gnd.n1941 0.152939
R14306 gnd.n3876 gnd.n3875 0.152939
R14307 gnd.n3877 gnd.n3876 0.152939
R14308 gnd.n3877 gnd.n1939 0.152939
R14309 gnd.n3883 gnd.n1939 0.152939
R14310 gnd.n3884 gnd.n3883 0.152939
R14311 gnd.n4063 gnd.n3884 0.152939
R14312 gnd.n4063 gnd.n4062 0.152939
R14313 gnd.n2758 gnd.n2757 0.152939
R14314 gnd.n2758 gnd.n2465 0.152939
R14315 gnd.n2799 gnd.n2465 0.152939
R14316 gnd.n2799 gnd.n2798 0.152939
R14317 gnd.n2798 gnd.n2797 0.152939
R14318 gnd.n2797 gnd.n2466 0.152939
R14319 gnd.n2793 gnd.n2466 0.152939
R14320 gnd.n2793 gnd.n2792 0.152939
R14321 gnd.n2792 gnd.n2791 0.152939
R14322 gnd.n2791 gnd.n2446 0.152939
R14323 gnd.n2844 gnd.n2446 0.152939
R14324 gnd.n2845 gnd.n2844 0.152939
R14325 gnd.n2846 gnd.n2845 0.152939
R14326 gnd.n2846 gnd.n2441 0.152939
R14327 gnd.n2859 gnd.n2441 0.152939
R14328 gnd.n2860 gnd.n2859 0.152939
R14329 gnd.n2861 gnd.n2860 0.152939
R14330 gnd.n2861 gnd.n2433 0.152939
R14331 gnd.n2895 gnd.n2433 0.152939
R14332 gnd.n2895 gnd.n2894 0.152939
R14333 gnd.n2894 gnd.n2893 0.152939
R14334 gnd.n2893 gnd.n2434 0.152939
R14335 gnd.n2889 gnd.n2434 0.152939
R14336 gnd.n2889 gnd.n2888 0.152939
R14337 gnd.n2888 gnd.n2887 0.152939
R14338 gnd.n2887 gnd.n2438 0.152939
R14339 gnd.n3175 gnd.n2941 0.152939
R14340 gnd.n3175 gnd.n3174 0.152939
R14341 gnd.n3174 gnd.n3173 0.152939
R14342 gnd.n3173 gnd.n2943 0.152939
R14343 gnd.n3169 gnd.n2943 0.152939
R14344 gnd.n3169 gnd.n3168 0.152939
R14345 gnd.n3216 gnd.n2385 0.152939
R14346 gnd.n3217 gnd.n3216 0.152939
R14347 gnd.n3219 gnd.n3217 0.152939
R14348 gnd.n3219 gnd.n3218 0.152939
R14349 gnd.n3218 gnd.n2361 0.152939
R14350 gnd.n3249 gnd.n2361 0.152939
R14351 gnd.n3250 gnd.n3249 0.152939
R14352 gnd.n3255 gnd.n3250 0.152939
R14353 gnd.n3255 gnd.n3254 0.152939
R14354 gnd.n3254 gnd.n3253 0.152939
R14355 gnd.n3253 gnd.n1509 0.152939
R14356 gnd.n4770 gnd.n1509 0.152939
R14357 gnd.n4770 gnd.n4769 0.152939
R14358 gnd.n4769 gnd.n4768 0.152939
R14359 gnd.n4768 gnd.n1510 0.152939
R14360 gnd.n4764 gnd.n1510 0.152939
R14361 gnd.n4764 gnd.n4763 0.152939
R14362 gnd.n4763 gnd.n4762 0.152939
R14363 gnd.n4762 gnd.n1515 0.152939
R14364 gnd.n4758 gnd.n1515 0.152939
R14365 gnd.n4758 gnd.n4757 0.152939
R14366 gnd.n4757 gnd.n4756 0.152939
R14367 gnd.n4756 gnd.n1520 0.152939
R14368 gnd.n4752 gnd.n1520 0.152939
R14369 gnd.n4752 gnd.n4751 0.152939
R14370 gnd.n4751 gnd.n4750 0.152939
R14371 gnd.n4750 gnd.n1525 0.152939
R14372 gnd.n4746 gnd.n1525 0.152939
R14373 gnd.n4746 gnd.n4745 0.152939
R14374 gnd.n4745 gnd.n4744 0.152939
R14375 gnd.n4744 gnd.n1530 0.152939
R14376 gnd.n4740 gnd.n1530 0.152939
R14377 gnd.n4740 gnd.n4739 0.152939
R14378 gnd.n4739 gnd.n4738 0.152939
R14379 gnd.n4738 gnd.n1535 0.152939
R14380 gnd.n4734 gnd.n1535 0.152939
R14381 gnd.n4734 gnd.n4733 0.152939
R14382 gnd.n4733 gnd.n4732 0.152939
R14383 gnd.n4732 gnd.n1540 0.152939
R14384 gnd.n4728 gnd.n1540 0.152939
R14385 gnd.n4728 gnd.n4727 0.152939
R14386 gnd.n4727 gnd.n4726 0.152939
R14387 gnd.n4726 gnd.n1545 0.152939
R14388 gnd.n4722 gnd.n1545 0.152939
R14389 gnd.n4722 gnd.n4721 0.152939
R14390 gnd.n4721 gnd.n4720 0.152939
R14391 gnd.n4720 gnd.n1550 0.152939
R14392 gnd.n4716 gnd.n1550 0.152939
R14393 gnd.n4716 gnd.n4715 0.152939
R14394 gnd.n4715 gnd.n4714 0.152939
R14395 gnd.n4714 gnd.n1555 0.152939
R14396 gnd.n4710 gnd.n1555 0.152939
R14397 gnd.n4710 gnd.n4709 0.152939
R14398 gnd.n4709 gnd.n4708 0.152939
R14399 gnd.n4708 gnd.n1560 0.152939
R14400 gnd.n4704 gnd.n1560 0.152939
R14401 gnd.n4704 gnd.n4703 0.152939
R14402 gnd.n4703 gnd.n4702 0.152939
R14403 gnd.n4702 gnd.n1565 0.152939
R14404 gnd.n4698 gnd.n1565 0.152939
R14405 gnd.n4698 gnd.n4697 0.152939
R14406 gnd.n4697 gnd.n4696 0.152939
R14407 gnd.n4696 gnd.n1570 0.152939
R14408 gnd.n4692 gnd.n1570 0.152939
R14409 gnd.n4692 gnd.n4691 0.152939
R14410 gnd.n4691 gnd.n4690 0.152939
R14411 gnd.n4690 gnd.n1575 0.152939
R14412 gnd.n4686 gnd.n1575 0.152939
R14413 gnd.n4686 gnd.n4685 0.152939
R14414 gnd.n4685 gnd.n4684 0.152939
R14415 gnd.n4684 gnd.n1580 0.152939
R14416 gnd.n4680 gnd.n1580 0.152939
R14417 gnd.n4680 gnd.n4679 0.152939
R14418 gnd.n4679 gnd.n4678 0.152939
R14419 gnd.n4678 gnd.n1585 0.152939
R14420 gnd.n4674 gnd.n1585 0.152939
R14421 gnd.n4674 gnd.n4673 0.152939
R14422 gnd.n4673 gnd.n4672 0.152939
R14423 gnd.n4672 gnd.n1590 0.152939
R14424 gnd.n4668 gnd.n1590 0.152939
R14425 gnd.n4668 gnd.n4667 0.152939
R14426 gnd.n4667 gnd.n4666 0.152939
R14427 gnd.n3949 gnd.n1595 0.152939
R14428 gnd.n3949 gnd.n3945 0.152939
R14429 gnd.n3957 gnd.n3945 0.152939
R14430 gnd.n3958 gnd.n3957 0.152939
R14431 gnd.n3960 gnd.n3958 0.152939
R14432 gnd.n3960 gnd.n3959 0.152939
R14433 gnd.n3890 gnd.n3885 0.152939
R14434 gnd.n3885 gnd.n1823 0.152939
R14435 gnd.n4437 gnd.n1823 0.152939
R14436 gnd.n4438 gnd.n4437 0.152939
R14437 gnd.n4439 gnd.n4438 0.152939
R14438 gnd.n4439 gnd.n1786 0.152939
R14439 gnd.n4451 gnd.n1786 0.152939
R14440 gnd.n4452 gnd.n4451 0.152939
R14441 gnd.n4453 gnd.n4452 0.152939
R14442 gnd.n4453 gnd.n1777 0.152939
R14443 gnd.n4489 gnd.n1777 0.152939
R14444 gnd.n4489 gnd.n4488 0.152939
R14445 gnd.n4488 gnd.n4487 0.152939
R14446 gnd.n4487 gnd.n1778 0.152939
R14447 gnd.n4483 gnd.n1778 0.152939
R14448 gnd.n4483 gnd.n4482 0.152939
R14449 gnd.n4482 gnd.n4481 0.152939
R14450 gnd.n4481 gnd.n1782 0.152939
R14451 gnd.n4477 gnd.n1782 0.152939
R14452 gnd.n4477 gnd.n1759 0.152939
R14453 gnd.n4549 gnd.n1759 0.152939
R14454 gnd.n4550 gnd.n4549 0.152939
R14455 gnd.n4554 gnd.n4550 0.152939
R14456 gnd.n4554 gnd.n4553 0.152939
R14457 gnd.n4553 gnd.n4552 0.152939
R14458 gnd.n4552 gnd.n79 0.152939
R14459 gnd.n3168 gnd.n3167 0.128549
R14460 gnd.n3959 gnd.n1827 0.128549
R14461 gnd.n2808 gnd.n1254 0.10111
R14462 gnd.n4509 gnd.n95 0.10111
R14463 gnd.n6005 gnd.n5397 0.0767195
R14464 gnd.n5921 gnd.n5397 0.0767195
R14465 gnd.n7744 gnd.n93 0.0767195
R14466 gnd.n7744 gnd.n94 0.0767195
R14467 gnd.n4975 gnd.n1253 0.0767195
R14468 gnd.n4975 gnd.n1251 0.0767195
R14469 gnd.n7754 gnd.n7753 0.0695946
R14470 gnd.n2756 gnd.n2755 0.0695946
R14471 gnd.n2757 gnd.n2756 0.0695946
R14472 gnd.n7754 gnd.n79 0.0695946
R14473 gnd.n3167 gnd.n3060 0.063
R14474 gnd.n4426 gnd.n1827 0.063
R14475 gnd.n385 gnd.n95 0.0523293
R14476 gnd.n2668 gnd.n1254 0.0523293
R14477 gnd.n6510 gnd.n5200 0.0477147
R14478 gnd.n4428 gnd.n4426 0.0477147
R14479 gnd.n7562 gnd.n207 0.0477147
R14480 gnd.n5045 gnd.n5044 0.0477147
R14481 gnd.n3060 gnd.n1371 0.0477147
R14482 gnd.n5671 gnd.n5567 0.0442063
R14483 gnd.n5685 gnd.n5567 0.0442063
R14484 gnd.n5686 gnd.n5685 0.0442063
R14485 gnd.n5687 gnd.n5686 0.0442063
R14486 gnd.n5687 gnd.n5555 0.0442063
R14487 gnd.n5701 gnd.n5555 0.0442063
R14488 gnd.n5702 gnd.n5701 0.0442063
R14489 gnd.n5703 gnd.n5702 0.0442063
R14490 gnd.n5703 gnd.n5542 0.0442063
R14491 gnd.n5799 gnd.n5542 0.0442063
R14492 gnd.n5802 gnd.n5801 0.0344674
R14493 gnd.n4429 gnd.n4428 0.0344674
R14494 gnd.n4429 gnd.n1637 0.0344674
R14495 gnd.n1638 gnd.n1637 0.0344674
R14496 gnd.n1639 gnd.n1638 0.0344674
R14497 gnd.n1821 gnd.n1639 0.0344674
R14498 gnd.n1821 gnd.n1657 0.0344674
R14499 gnd.n1658 gnd.n1657 0.0344674
R14500 gnd.n1659 gnd.n1658 0.0344674
R14501 gnd.n1784 gnd.n1659 0.0344674
R14502 gnd.n1784 gnd.n1678 0.0344674
R14503 gnd.n1679 gnd.n1678 0.0344674
R14504 gnd.n1680 gnd.n1679 0.0344674
R14505 gnd.n4462 gnd.n1680 0.0344674
R14506 gnd.n4462 gnd.n1697 0.0344674
R14507 gnd.n1698 gnd.n1697 0.0344674
R14508 gnd.n1699 gnd.n1698 0.0344674
R14509 gnd.n4472 gnd.n1699 0.0344674
R14510 gnd.n4472 gnd.n1718 0.0344674
R14511 gnd.n1719 gnd.n1718 0.0344674
R14512 gnd.n1720 gnd.n1719 0.0344674
R14513 gnd.n4520 gnd.n1720 0.0344674
R14514 gnd.n4520 gnd.n1735 0.0344674
R14515 gnd.n1736 gnd.n1735 0.0344674
R14516 gnd.n1737 gnd.n1736 0.0344674
R14517 gnd.n4521 gnd.n1737 0.0344674
R14518 gnd.n4522 gnd.n4521 0.0344674
R14519 gnd.n4527 gnd.n4522 0.0344674
R14520 gnd.n4529 gnd.n4527 0.0344674
R14521 gnd.n4530 gnd.n4529 0.0344674
R14522 gnd.n4530 gnd.n379 0.0344674
R14523 gnd.n379 gnd.n109 0.0344674
R14524 gnd.n110 gnd.n109 0.0344674
R14525 gnd.n111 gnd.n110 0.0344674
R14526 gnd.n373 gnd.n111 0.0344674
R14527 gnd.n373 gnd.n127 0.0344674
R14528 gnd.n128 gnd.n127 0.0344674
R14529 gnd.n129 gnd.n128 0.0344674
R14530 gnd.n367 gnd.n129 0.0344674
R14531 gnd.n367 gnd.n148 0.0344674
R14532 gnd.n149 gnd.n148 0.0344674
R14533 gnd.n150 gnd.n149 0.0344674
R14534 gnd.n361 gnd.n150 0.0344674
R14535 gnd.n361 gnd.n167 0.0344674
R14536 gnd.n168 gnd.n167 0.0344674
R14537 gnd.n169 gnd.n168 0.0344674
R14538 gnd.n7493 gnd.n169 0.0344674
R14539 gnd.n7493 gnd.n187 0.0344674
R14540 gnd.n188 gnd.n187 0.0344674
R14541 gnd.n189 gnd.n188 0.0344674
R14542 gnd.n7494 gnd.n189 0.0344674
R14543 gnd.n7494 gnd.n205 0.0344674
R14544 gnd.n206 gnd.n205 0.0344674
R14545 gnd.n207 gnd.n206 0.0344674
R14546 gnd.n5044 gnd.n1138 0.0344674
R14547 gnd.n2529 gnd.n1138 0.0344674
R14548 gnd.n2529 gnd.n1160 0.0344674
R14549 gnd.n1161 gnd.n1160 0.0344674
R14550 gnd.n1162 gnd.n1161 0.0344674
R14551 gnd.n2535 gnd.n1162 0.0344674
R14552 gnd.n2535 gnd.n1179 0.0344674
R14553 gnd.n1180 gnd.n1179 0.0344674
R14554 gnd.n1181 gnd.n1180 0.0344674
R14555 gnd.n2542 gnd.n1181 0.0344674
R14556 gnd.n2542 gnd.n1199 0.0344674
R14557 gnd.n1200 gnd.n1199 0.0344674
R14558 gnd.n1201 gnd.n1200 0.0344674
R14559 gnd.n2525 gnd.n1201 0.0344674
R14560 gnd.n2525 gnd.n1219 0.0344674
R14561 gnd.n1220 gnd.n1219 0.0344674
R14562 gnd.n1221 gnd.n1220 0.0344674
R14563 gnd.n2520 gnd.n1221 0.0344674
R14564 gnd.n2520 gnd.n1240 0.0344674
R14565 gnd.n1241 gnd.n1240 0.0344674
R14566 gnd.n1242 gnd.n1241 0.0344674
R14567 gnd.n2507 gnd.n1242 0.0344674
R14568 gnd.n2719 gnd.n2507 0.0344674
R14569 gnd.n2719 gnd.n2508 0.0344674
R14570 gnd.n2508 gnd.n2493 0.0344674
R14571 gnd.n2494 gnd.n2493 0.0344674
R14572 gnd.n2495 gnd.n2494 0.0344674
R14573 gnd.n2495 gnd.n2471 0.0344674
R14574 gnd.n2769 gnd.n2471 0.0344674
R14575 gnd.n2770 gnd.n2769 0.0344674
R14576 gnd.n2770 gnd.n1269 0.0344674
R14577 gnd.n1270 gnd.n1269 0.0344674
R14578 gnd.n1271 gnd.n1270 0.0344674
R14579 gnd.n2777 gnd.n1271 0.0344674
R14580 gnd.n2777 gnd.n1288 0.0344674
R14581 gnd.n1289 gnd.n1288 0.0344674
R14582 gnd.n1290 gnd.n1289 0.0344674
R14583 gnd.n2783 gnd.n1290 0.0344674
R14584 gnd.n2783 gnd.n1308 0.0344674
R14585 gnd.n1309 gnd.n1308 0.0344674
R14586 gnd.n1310 gnd.n1309 0.0344674
R14587 gnd.n2853 gnd.n1310 0.0344674
R14588 gnd.n2853 gnd.n1328 0.0344674
R14589 gnd.n1329 gnd.n1328 0.0344674
R14590 gnd.n1330 gnd.n1329 0.0344674
R14591 gnd.n2868 gnd.n1330 0.0344674
R14592 gnd.n2868 gnd.n1348 0.0344674
R14593 gnd.n1349 gnd.n1348 0.0344674
R14594 gnd.n1350 gnd.n1349 0.0344674
R14595 gnd.n2875 gnd.n1350 0.0344674
R14596 gnd.n2875 gnd.n1369 0.0344674
R14597 gnd.n1370 gnd.n1369 0.0344674
R14598 gnd.n1371 gnd.n1370 0.0344674
R14599 gnd.n3166 gnd.n3061 0.0344674
R14600 gnd.n3969 gnd.n3968 0.0344674
R14601 gnd.n3193 gnd.n2400 0.029712
R14602 gnd.n3900 gnd.n3891 0.029712
R14603 gnd.n5535 gnd.n5534 0.0269946
R14604 gnd.n5812 gnd.n5532 0.0269946
R14605 gnd.n5811 gnd.n5533 0.0269946
R14606 gnd.n5831 gnd.n5514 0.0269946
R14607 gnd.n5833 gnd.n5832 0.0269946
R14608 gnd.n5834 gnd.n5512 0.0269946
R14609 gnd.n5841 gnd.n5837 0.0269946
R14610 gnd.n5840 gnd.n5839 0.0269946
R14611 gnd.n5838 gnd.n5491 0.0269946
R14612 gnd.n5865 gnd.n5492 0.0269946
R14613 gnd.n5864 gnd.n5493 0.0269946
R14614 gnd.n5897 gnd.n5467 0.0269946
R14615 gnd.n5899 gnd.n5898 0.0269946
R14616 gnd.n5900 gnd.n5459 0.0269946
R14617 gnd.n5463 gnd.n5460 0.0269946
R14618 gnd.n5910 gnd.n5461 0.0269946
R14619 gnd.n5909 gnd.n5462 0.0269946
R14620 gnd.n5955 gnd.n5435 0.0269946
R14621 gnd.n5957 gnd.n5956 0.0269946
R14622 gnd.n5966 gnd.n5428 0.0269946
R14623 gnd.n5968 gnd.n5967 0.0269946
R14624 gnd.n5969 gnd.n5426 0.0269946
R14625 gnd.n5976 gnd.n5972 0.0269946
R14626 gnd.n5975 gnd.n5974 0.0269946
R14627 gnd.n5973 gnd.n5405 0.0269946
R14628 gnd.n5998 gnd.n5406 0.0269946
R14629 gnd.n5997 gnd.n5407 0.0269946
R14630 gnd.n6040 gnd.n5316 0.0269946
R14631 gnd.n6042 gnd.n6041 0.0269946
R14632 gnd.n6051 gnd.n5309 0.0269946
R14633 gnd.n6053 gnd.n6052 0.0269946
R14634 gnd.n6054 gnd.n5307 0.0269946
R14635 gnd.n6060 gnd.n6057 0.0269946
R14636 gnd.n6059 gnd.n6058 0.0269946
R14637 gnd.n6085 gnd.n5287 0.0269946
R14638 gnd.n6084 gnd.n5288 0.0269946
R14639 gnd.n6114 gnd.n5273 0.0269946
R14640 gnd.n6116 gnd.n6115 0.0269946
R14641 gnd.n6140 gnd.n5259 0.0269946
R14642 gnd.n6142 gnd.n6141 0.0269946
R14643 gnd.n6143 gnd.n974 0.0269946
R14644 gnd.n5254 gnd.n975 0.0269946
R14645 gnd.n5256 gnd.n976 0.0269946
R14646 gnd.n6151 gnd.n6150 0.0269946
R14647 gnd.n6153 gnd.n6152 0.0269946
R14648 gnd.n6154 gnd.n997 0.0269946
R14649 gnd.n6155 gnd.n998 0.0269946
R14650 gnd.n6156 gnd.n999 0.0269946
R14651 gnd.n6416 gnd.n6415 0.0269946
R14652 gnd.n6417 gnd.n1023 0.0269946
R14653 gnd.n6418 gnd.n1024 0.0269946
R14654 gnd.n6419 gnd.n1025 0.0269946
R14655 gnd.n3162 gnd.n3067 0.0225788
R14656 gnd.n3161 gnd.n3068 0.0225788
R14657 gnd.n3158 gnd.n3157 0.0225788
R14658 gnd.n3154 gnd.n3074 0.0225788
R14659 gnd.n3153 gnd.n3080 0.0225788
R14660 gnd.n3150 gnd.n3149 0.0225788
R14661 gnd.n3146 gnd.n3086 0.0225788
R14662 gnd.n3145 gnd.n3090 0.0225788
R14663 gnd.n3142 gnd.n3141 0.0225788
R14664 gnd.n3138 gnd.n3097 0.0225788
R14665 gnd.n3137 gnd.n3103 0.0225788
R14666 gnd.n3134 gnd.n3133 0.0225788
R14667 gnd.n3130 gnd.n3109 0.0225788
R14668 gnd.n3129 gnd.n3113 0.0225788
R14669 gnd.n3126 gnd.n3125 0.0225788
R14670 gnd.n3120 gnd.n2409 0.0225788
R14671 gnd.n3185 gnd.n3184 0.0225788
R14672 gnd.n2410 gnd.n2403 0.0225788
R14673 gnd.n3193 gnd.n3192 0.0225788
R14674 gnd.n3975 gnd.n3973 0.0225788
R14675 gnd.n3974 gnd.n3937 0.0225788
R14676 gnd.n3984 gnd.n3983 0.0225788
R14677 gnd.n3938 gnd.n3933 0.0225788
R14678 gnd.n3994 gnd.n3992 0.0225788
R14679 gnd.n3993 gnd.n3928 0.0225788
R14680 gnd.n4003 gnd.n4002 0.0225788
R14681 gnd.n3929 gnd.n3924 0.0225788
R14682 gnd.n4013 gnd.n4011 0.0225788
R14683 gnd.n4012 gnd.n3919 0.0225788
R14684 gnd.n4022 gnd.n4021 0.0225788
R14685 gnd.n3920 gnd.n3915 0.0225788
R14686 gnd.n4032 gnd.n4030 0.0225788
R14687 gnd.n4031 gnd.n3910 0.0225788
R14688 gnd.n4042 gnd.n4041 0.0225788
R14689 gnd.n4038 gnd.n3911 0.0225788
R14690 gnd.n4052 gnd.n3898 0.0225788
R14691 gnd.n4051 gnd.n3899 0.0225788
R14692 gnd.n3901 gnd.n3900 0.0225788
R14693 gnd.n4061 gnd.n3891 0.0218415
R14694 gnd.n3196 gnd.n2400 0.0218415
R14695 gnd.n5801 gnd.n5800 0.0202011
R14696 gnd.n5800 gnd.n5799 0.0148637
R14697 gnd.n6413 gnd.n6157 0.0144266
R14698 gnd.n6414 gnd.n6413 0.0130679
R14699 gnd.n3067 gnd.n3061 0.0123886
R14700 gnd.n3162 gnd.n3161 0.0123886
R14701 gnd.n3158 gnd.n3068 0.0123886
R14702 gnd.n3157 gnd.n3074 0.0123886
R14703 gnd.n3154 gnd.n3153 0.0123886
R14704 gnd.n3150 gnd.n3080 0.0123886
R14705 gnd.n3149 gnd.n3086 0.0123886
R14706 gnd.n3146 gnd.n3145 0.0123886
R14707 gnd.n3142 gnd.n3090 0.0123886
R14708 gnd.n3141 gnd.n3097 0.0123886
R14709 gnd.n3138 gnd.n3137 0.0123886
R14710 gnd.n3134 gnd.n3103 0.0123886
R14711 gnd.n3133 gnd.n3109 0.0123886
R14712 gnd.n3130 gnd.n3129 0.0123886
R14713 gnd.n3126 gnd.n3113 0.0123886
R14714 gnd.n3125 gnd.n3120 0.0123886
R14715 gnd.n3185 gnd.n2409 0.0123886
R14716 gnd.n3184 gnd.n2410 0.0123886
R14717 gnd.n3192 gnd.n2403 0.0123886
R14718 gnd.n3973 gnd.n3969 0.0123886
R14719 gnd.n3975 gnd.n3974 0.0123886
R14720 gnd.n3984 gnd.n3937 0.0123886
R14721 gnd.n3983 gnd.n3938 0.0123886
R14722 gnd.n3992 gnd.n3933 0.0123886
R14723 gnd.n3994 gnd.n3993 0.0123886
R14724 gnd.n4003 gnd.n3928 0.0123886
R14725 gnd.n4002 gnd.n3929 0.0123886
R14726 gnd.n4011 gnd.n3924 0.0123886
R14727 gnd.n4013 gnd.n4012 0.0123886
R14728 gnd.n4022 gnd.n3919 0.0123886
R14729 gnd.n4021 gnd.n3920 0.0123886
R14730 gnd.n4030 gnd.n3915 0.0123886
R14731 gnd.n4032 gnd.n4031 0.0123886
R14732 gnd.n4042 gnd.n3910 0.0123886
R14733 gnd.n4041 gnd.n3911 0.0123886
R14734 gnd.n4038 gnd.n3898 0.0123886
R14735 gnd.n4052 gnd.n4051 0.0123886
R14736 gnd.n3901 gnd.n3899 0.0123886
R14737 gnd.n5802 gnd.n5535 0.00797283
R14738 gnd.n5534 gnd.n5532 0.00797283
R14739 gnd.n5812 gnd.n5811 0.00797283
R14740 gnd.n5533 gnd.n5514 0.00797283
R14741 gnd.n5832 gnd.n5831 0.00797283
R14742 gnd.n5834 gnd.n5833 0.00797283
R14743 gnd.n5837 gnd.n5512 0.00797283
R14744 gnd.n5841 gnd.n5840 0.00797283
R14745 gnd.n5839 gnd.n5838 0.00797283
R14746 gnd.n5492 gnd.n5491 0.00797283
R14747 gnd.n5865 gnd.n5864 0.00797283
R14748 gnd.n5493 gnd.n5467 0.00797283
R14749 gnd.n5898 gnd.n5897 0.00797283
R14750 gnd.n5900 gnd.n5899 0.00797283
R14751 gnd.n5463 gnd.n5459 0.00797283
R14752 gnd.n5461 gnd.n5460 0.00797283
R14753 gnd.n5910 gnd.n5909 0.00797283
R14754 gnd.n5462 gnd.n5435 0.00797283
R14755 gnd.n5957 gnd.n5955 0.00797283
R14756 gnd.n5956 gnd.n5428 0.00797283
R14757 gnd.n5967 gnd.n5966 0.00797283
R14758 gnd.n5969 gnd.n5968 0.00797283
R14759 gnd.n5972 gnd.n5426 0.00797283
R14760 gnd.n5976 gnd.n5975 0.00797283
R14761 gnd.n5974 gnd.n5973 0.00797283
R14762 gnd.n5406 gnd.n5405 0.00797283
R14763 gnd.n5998 gnd.n5997 0.00797283
R14764 gnd.n5407 gnd.n5316 0.00797283
R14765 gnd.n6042 gnd.n6040 0.00797283
R14766 gnd.n6041 gnd.n5309 0.00797283
R14767 gnd.n6052 gnd.n6051 0.00797283
R14768 gnd.n6054 gnd.n6053 0.00797283
R14769 gnd.n6057 gnd.n5307 0.00797283
R14770 gnd.n6060 gnd.n6059 0.00797283
R14771 gnd.n6058 gnd.n5287 0.00797283
R14772 gnd.n6085 gnd.n6084 0.00797283
R14773 gnd.n5288 gnd.n5273 0.00797283
R14774 gnd.n6116 gnd.n6114 0.00797283
R14775 gnd.n6115 gnd.n5259 0.00797283
R14776 gnd.n6141 gnd.n6140 0.00797283
R14777 gnd.n6143 gnd.n6142 0.00797283
R14778 gnd.n5254 gnd.n974 0.00797283
R14779 gnd.n5256 gnd.n975 0.00797283
R14780 gnd.n6150 gnd.n976 0.00797283
R14781 gnd.n6152 gnd.n6151 0.00797283
R14782 gnd.n6154 gnd.n6153 0.00797283
R14783 gnd.n6155 gnd.n997 0.00797283
R14784 gnd.n6156 gnd.n998 0.00797283
R14785 gnd.n6157 gnd.n999 0.00797283
R14786 gnd.n6415 gnd.n6414 0.00797283
R14787 gnd.n6417 gnd.n6416 0.00797283
R14788 gnd.n6418 gnd.n1023 0.00797283
R14789 gnd.n6419 gnd.n1024 0.00797283
R14790 gnd.n5200 gnd.n1025 0.00797283
R14791 gnd.n3167 gnd.n3166 0.00593478
R14792 gnd.n3968 gnd.n1827 0.00593478
R14793 a_n2982_13878.n125 a_n2982_13878.t94 512.366
R14794 a_n2982_13878.n115 a_n2982_13878.t83 512.366
R14795 a_n2982_13878.n126 a_n2982_13878.t72 512.366
R14796 a_n2982_13878.n123 a_n2982_13878.t102 512.366
R14797 a_n2982_13878.n116 a_n2982_13878.t91 512.366
R14798 a_n2982_13878.n124 a_n2982_13878.t90 512.366
R14799 a_n2982_13878.n121 a_n2982_13878.t98 512.366
R14800 a_n2982_13878.n117 a_n2982_13878.t81 512.366
R14801 a_n2982_13878.n122 a_n2982_13878.t82 512.366
R14802 a_n2982_13878.n119 a_n2982_13878.t85 512.366
R14803 a_n2982_13878.n118 a_n2982_13878.t96 512.366
R14804 a_n2982_13878.n120 a_n2982_13878.t111 512.366
R14805 a_n2982_13878.n31 a_n2982_13878.t110 538.698
R14806 a_n2982_13878.n134 a_n2982_13878.t87 512.366
R14807 a_n2982_13878.n133 a_n2982_13878.t92 512.366
R14808 a_n2982_13878.n86 a_n2982_13878.t80 512.366
R14809 a_n2982_13878.n132 a_n2982_13878.t97 512.366
R14810 a_n2982_13878.n131 a_n2982_13878.t106 512.366
R14811 a_n2982_13878.n87 a_n2982_13878.t107 512.366
R14812 a_n2982_13878.n130 a_n2982_13878.t74 512.366
R14813 a_n2982_13878.n129 a_n2982_13878.t89 512.366
R14814 a_n2982_13878.n88 a_n2982_13878.t77 512.366
R14815 a_n2982_13878.n128 a_n2982_13878.t84 512.366
R14816 a_n2982_13878.n33 a_n2982_13878.t33 538.699
R14817 a_n2982_13878.n135 a_n2982_13878.t25 512.366
R14818 a_n2982_13878.n83 a_n2982_13878.t49 512.366
R14819 a_n2982_13878.n38 a_n2982_13878.t11 538.698
R14820 a_n2982_13878.n153 a_n2982_13878.t37 512.366
R14821 a_n2982_13878.n152 a_n2982_13878.t57 512.366
R14822 a_n2982_13878.n84 a_n2982_13878.t29 512.366
R14823 a_n2982_13878.n151 a_n2982_13878.t55 512.366
R14824 a_n2982_13878.n150 a_n2982_13878.t15 512.366
R14825 a_n2982_13878.n85 a_n2982_13878.t17 512.366
R14826 a_n2982_13878.n149 a_n2982_13878.t31 512.366
R14827 a_n2982_13878.n148 a_n2982_13878.t41 512.366
R14828 a_n2982_13878.n19 a_n2982_13878.t23 538.698
R14829 a_n2982_13878.n108 a_n2982_13878.t19 512.366
R14830 a_n2982_13878.n97 a_n2982_13878.t47 512.366
R14831 a_n2982_13878.n109 a_n2982_13878.t53 512.366
R14832 a_n2982_13878.n96 a_n2982_13878.t39 512.366
R14833 a_n2982_13878.n110 a_n2982_13878.t51 512.366
R14834 a_n2982_13878.n111 a_n2982_13878.t43 512.366
R14835 a_n2982_13878.n95 a_n2982_13878.t13 512.366
R14836 a_n2982_13878.n112 a_n2982_13878.t35 512.366
R14837 a_n2982_13878.n94 a_n2982_13878.t27 512.366
R14838 a_n2982_13878.n113 a_n2982_13878.t21 512.366
R14839 a_n2982_13878.n25 a_n2982_13878.t109 538.698
R14840 a_n2982_13878.n102 a_n2982_13878.t78 512.366
R14841 a_n2982_13878.n101 a_n2982_13878.t79 512.366
R14842 a_n2982_13878.n103 a_n2982_13878.t104 512.366
R14843 a_n2982_13878.n100 a_n2982_13878.t105 512.366
R14844 a_n2982_13878.n104 a_n2982_13878.t76 512.366
R14845 a_n2982_13878.n105 a_n2982_13878.t100 512.366
R14846 a_n2982_13878.n99 a_n2982_13878.t101 512.366
R14847 a_n2982_13878.n106 a_n2982_13878.t73 512.366
R14848 a_n2982_13878.n98 a_n2982_13878.t86 512.366
R14849 a_n2982_13878.n107 a_n2982_13878.t95 512.366
R14850 a_n2982_13878.n5 a_n2982_13878.n82 70.1674
R14851 a_n2982_13878.n7 a_n2982_13878.n80 70.1674
R14852 a_n2982_13878.n9 a_n2982_13878.n78 70.1674
R14853 a_n2982_13878.n12 a_n2982_13878.n76 70.1674
R14854 a_n2982_13878.n58 a_n2982_13878.n26 70.5844
R14855 a_n2982_13878.n50 a_n2982_13878.n32 44.5605
R14856 a_n2982_13878.n148 a_n2982_13878.n50 21.3688
R14857 a_n2982_13878.n49 a_n2982_13878.n34 80.4688
R14858 a_n2982_13878.n49 a_n2982_13878.n149 0.365327
R14859 a_n2982_13878.n35 a_n2982_13878.n48 75.0448
R14860 a_n2982_13878.n47 a_n2982_13878.n35 70.1674
R14861 a_n2982_13878.n151 a_n2982_13878.n47 20.9683
R14862 a_n2982_13878.n37 a_n2982_13878.n46 70.3058
R14863 a_n2982_13878.n46 a_n2982_13878.n84 20.6913
R14864 a_n2982_13878.n45 a_n2982_13878.n37 75.3623
R14865 a_n2982_13878.n152 a_n2982_13878.n45 10.5784
R14866 a_n2982_13878.n36 a_n2982_13878.n38 44.7878
R14867 a_n2982_13878.n33 a_n2982_13878.n32 44.7878
R14868 a_n2982_13878.n33 a_n2982_13878.n135 14.1664
R14869 a_n2982_13878.n26 a_n2982_13878.n57 70.1674
R14870 a_n2982_13878.n57 a_n2982_13878.n88 20.9683
R14871 a_n2982_13878.n56 a_n2982_13878.n27 74.73
R14872 a_n2982_13878.n129 a_n2982_13878.n56 11.843
R14873 a_n2982_13878.n55 a_n2982_13878.n27 80.4688
R14874 a_n2982_13878.n55 a_n2982_13878.n130 0.365327
R14875 a_n2982_13878.n28 a_n2982_13878.n54 75.0448
R14876 a_n2982_13878.n53 a_n2982_13878.n28 70.1674
R14877 a_n2982_13878.n132 a_n2982_13878.n53 20.9683
R14878 a_n2982_13878.n30 a_n2982_13878.n52 70.3058
R14879 a_n2982_13878.n52 a_n2982_13878.n86 20.6913
R14880 a_n2982_13878.n51 a_n2982_13878.n30 75.3623
R14881 a_n2982_13878.n133 a_n2982_13878.n51 10.5784
R14882 a_n2982_13878.n29 a_n2982_13878.n31 44.7878
R14883 a_n2982_13878.n15 a_n2982_13878.n74 70.5844
R14884 a_n2982_13878.n21 a_n2982_13878.n66 70.5844
R14885 a_n2982_13878.n65 a_n2982_13878.n21 70.1674
R14886 a_n2982_13878.n65 a_n2982_13878.n98 20.9683
R14887 a_n2982_13878.n20 a_n2982_13878.n64 74.73
R14888 a_n2982_13878.n106 a_n2982_13878.n64 11.843
R14889 a_n2982_13878.n63 a_n2982_13878.n20 80.4688
R14890 a_n2982_13878.n63 a_n2982_13878.n99 0.365327
R14891 a_n2982_13878.n22 a_n2982_13878.n62 75.0448
R14892 a_n2982_13878.n61 a_n2982_13878.n22 70.1674
R14893 a_n2982_13878.n61 a_n2982_13878.n100 20.9683
R14894 a_n2982_13878.n23 a_n2982_13878.n60 70.3058
R14895 a_n2982_13878.n103 a_n2982_13878.n60 20.6913
R14896 a_n2982_13878.n59 a_n2982_13878.n23 75.3623
R14897 a_n2982_13878.n59 a_n2982_13878.n101 10.5784
R14898 a_n2982_13878.n25 a_n2982_13878.n24 44.7878
R14899 a_n2982_13878.n73 a_n2982_13878.n15 70.1674
R14900 a_n2982_13878.n73 a_n2982_13878.n94 20.9683
R14901 a_n2982_13878.n14 a_n2982_13878.n72 74.73
R14902 a_n2982_13878.n112 a_n2982_13878.n72 11.843
R14903 a_n2982_13878.n71 a_n2982_13878.n14 80.4688
R14904 a_n2982_13878.n71 a_n2982_13878.n95 0.365327
R14905 a_n2982_13878.n16 a_n2982_13878.n70 75.0448
R14906 a_n2982_13878.n69 a_n2982_13878.n16 70.1674
R14907 a_n2982_13878.n69 a_n2982_13878.n96 20.9683
R14908 a_n2982_13878.n17 a_n2982_13878.n68 70.3058
R14909 a_n2982_13878.n109 a_n2982_13878.n68 20.6913
R14910 a_n2982_13878.n67 a_n2982_13878.n17 75.3623
R14911 a_n2982_13878.n67 a_n2982_13878.n97 10.5784
R14912 a_n2982_13878.n19 a_n2982_13878.n18 44.7878
R14913 a_n2982_13878.n120 a_n2982_13878.n76 20.9683
R14914 a_n2982_13878.n75 a_n2982_13878.n13 75.0448
R14915 a_n2982_13878.n75 a_n2982_13878.n118 11.2134
R14916 a_n2982_13878.n13 a_n2982_13878.n119 161.3
R14917 a_n2982_13878.n122 a_n2982_13878.n78 20.9683
R14918 a_n2982_13878.n77 a_n2982_13878.n10 75.0448
R14919 a_n2982_13878.n77 a_n2982_13878.n117 11.2134
R14920 a_n2982_13878.n10 a_n2982_13878.n121 161.3
R14921 a_n2982_13878.n124 a_n2982_13878.n80 20.9683
R14922 a_n2982_13878.n79 a_n2982_13878.n8 75.0448
R14923 a_n2982_13878.n79 a_n2982_13878.n116 11.2134
R14924 a_n2982_13878.n8 a_n2982_13878.n123 161.3
R14925 a_n2982_13878.n126 a_n2982_13878.n82 20.9683
R14926 a_n2982_13878.n81 a_n2982_13878.n6 75.0448
R14927 a_n2982_13878.n81 a_n2982_13878.n115 11.2134
R14928 a_n2982_13878.n6 a_n2982_13878.n125 161.3
R14929 a_n2982_13878.n3 a_n2982_13878.n145 81.3764
R14930 a_n2982_13878.n4 a_n2982_13878.n139 81.3764
R14931 a_n2982_13878.n0 a_n2982_13878.n136 81.3764
R14932 a_n2982_13878.n3 a_n2982_13878.n146 80.9324
R14933 a_n2982_13878.n2 a_n2982_13878.n147 80.9324
R14934 a_n2982_13878.n2 a_n2982_13878.n144 80.9324
R14935 a_n2982_13878.n2 a_n2982_13878.n143 80.9324
R14936 a_n2982_13878.n1 a_n2982_13878.n142 80.9324
R14937 a_n2982_13878.n4 a_n2982_13878.n140 80.9324
R14938 a_n2982_13878.n0 a_n2982_13878.n141 80.9324
R14939 a_n2982_13878.n0 a_n2982_13878.n138 80.9324
R14940 a_n2982_13878.n0 a_n2982_13878.n137 80.9324
R14941 a_n2982_13878.n44 a_n2982_13878.t34 74.6477
R14942 a_n2982_13878.n39 a_n2982_13878.t24 74.6477
R14943 a_n2982_13878.t12 a_n2982_13878.n43 74.2899
R14944 a_n2982_13878.n41 a_n2982_13878.t46 74.2897
R14945 a_n2982_13878.n44 a_n2982_13878.n155 70.6783
R14946 a_n2982_13878.n44 a_n2982_13878.n156 70.6783
R14947 a_n2982_13878.n42 a_n2982_13878.n157 70.6783
R14948 a_n2982_13878.n42 a_n2982_13878.n158 70.6783
R14949 a_n2982_13878.n43 a_n2982_13878.n159 70.6783
R14950 a_n2982_13878.n41 a_n2982_13878.n93 70.6783
R14951 a_n2982_13878.n40 a_n2982_13878.n92 70.6783
R14952 a_n2982_13878.n40 a_n2982_13878.n91 70.6783
R14953 a_n2982_13878.n39 a_n2982_13878.n90 70.6783
R14954 a_n2982_13878.n39 a_n2982_13878.n89 70.6783
R14955 a_n2982_13878.n125 a_n2982_13878.n115 48.2005
R14956 a_n2982_13878.t99 a_n2982_13878.n82 533.335
R14957 a_n2982_13878.n123 a_n2982_13878.n116 48.2005
R14958 a_n2982_13878.t108 a_n2982_13878.n80 533.335
R14959 a_n2982_13878.n121 a_n2982_13878.n117 48.2005
R14960 a_n2982_13878.t93 a_n2982_13878.n78 533.335
R14961 a_n2982_13878.n119 a_n2982_13878.n118 48.2005
R14962 a_n2982_13878.t88 a_n2982_13878.n76 533.335
R14963 a_n2982_13878.n134 a_n2982_13878.n133 48.2005
R14964 a_n2982_13878.n53 a_n2982_13878.n131 20.9683
R14965 a_n2982_13878.n130 a_n2982_13878.n87 48.2005
R14966 a_n2982_13878.n128 a_n2982_13878.n57 20.9683
R14967 a_n2982_13878.n135 a_n2982_13878.n83 48.2005
R14968 a_n2982_13878.n153 a_n2982_13878.n152 48.2005
R14969 a_n2982_13878.n47 a_n2982_13878.n150 20.9683
R14970 a_n2982_13878.n149 a_n2982_13878.n85 48.2005
R14971 a_n2982_13878.n108 a_n2982_13878.n97 48.2005
R14972 a_n2982_13878.n110 a_n2982_13878.n69 20.9683
R14973 a_n2982_13878.n111 a_n2982_13878.n95 48.2005
R14974 a_n2982_13878.n113 a_n2982_13878.n73 20.9683
R14975 a_n2982_13878.n102 a_n2982_13878.n101 48.2005
R14976 a_n2982_13878.n104 a_n2982_13878.n61 20.9683
R14977 a_n2982_13878.n105 a_n2982_13878.n99 48.2005
R14978 a_n2982_13878.n107 a_n2982_13878.n65 20.9683
R14979 a_n2982_13878.n132 a_n2982_13878.n52 21.4216
R14980 a_n2982_13878.n151 a_n2982_13878.n46 21.4216
R14981 a_n2982_13878.n96 a_n2982_13878.n68 21.4216
R14982 a_n2982_13878.n100 a_n2982_13878.n60 21.4216
R14983 a_n2982_13878.n58 a_n2982_13878.t103 532.5
R14984 a_n2982_13878.t45 a_n2982_13878.n74 532.5
R14985 a_n2982_13878.t75 a_n2982_13878.n66 532.5
R14986 a_n2982_13878.n1 a_n2982_13878.n0 32.6799
R14987 a_n2982_13878.n56 a_n2982_13878.n88 34.4824
R14988 a_n2982_13878.n50 a_n2982_13878.n83 20.5623
R14989 a_n2982_13878.n94 a_n2982_13878.n72 34.4824
R14990 a_n2982_13878.n98 a_n2982_13878.n64 34.4824
R14991 a_n2982_13878.n126 a_n2982_13878.n81 35.3134
R14992 a_n2982_13878.n124 a_n2982_13878.n79 35.3134
R14993 a_n2982_13878.n122 a_n2982_13878.n77 35.3134
R14994 a_n2982_13878.n120 a_n2982_13878.n75 35.3134
R14995 a_n2982_13878.n131 a_n2982_13878.n54 35.3134
R14996 a_n2982_13878.n54 a_n2982_13878.n87 11.2134
R14997 a_n2982_13878.n150 a_n2982_13878.n48 35.3134
R14998 a_n2982_13878.n48 a_n2982_13878.n85 11.2134
R14999 a_n2982_13878.n70 a_n2982_13878.n110 35.3134
R15000 a_n2982_13878.n111 a_n2982_13878.n70 11.2134
R15001 a_n2982_13878.n62 a_n2982_13878.n104 35.3134
R15002 a_n2982_13878.n105 a_n2982_13878.n62 11.2134
R15003 a_n2982_13878.n32 a_n2982_13878.n2 23.891
R15004 a_n2982_13878.n51 a_n2982_13878.n86 36.139
R15005 a_n2982_13878.n45 a_n2982_13878.n84 36.139
R15006 a_n2982_13878.n109 a_n2982_13878.n67 36.139
R15007 a_n2982_13878.n103 a_n2982_13878.n59 36.139
R15008 a_n2982_13878.n24 a_n2982_13878.n11 13.9285
R15009 a_n2982_13878.n26 a_n2982_13878.n127 13.724
R15010 a_n2982_13878.n154 a_n2982_13878.n36 12.4191
R15011 a_n2982_13878.n127 a_n2982_13878.n5 11.2486
R15012 a_n2982_13878.n13 a_n2982_13878.n11 11.2486
R15013 a_n2982_13878.n114 a_n2982_13878.n41 10.5745
R15014 a_n2982_13878.n114 a_n2982_13878.n15 8.58383
R15015 a_n2982_13878.n43 a_n2982_13878.n154 6.7311
R15016 a_n2982_13878.n127 a_n2982_13878.n114 5.3452
R15017 a_n2982_13878.n32 a_n2982_13878.n29 3.94368
R15018 a_n2982_13878.n18 a_n2982_13878.n21 3.94368
R15019 a_n2982_13878.n155 a_n2982_13878.t50 3.61217
R15020 a_n2982_13878.n155 a_n2982_13878.t26 3.61217
R15021 a_n2982_13878.n156 a_n2982_13878.t32 3.61217
R15022 a_n2982_13878.n156 a_n2982_13878.t42 3.61217
R15023 a_n2982_13878.n157 a_n2982_13878.t16 3.61217
R15024 a_n2982_13878.n157 a_n2982_13878.t18 3.61217
R15025 a_n2982_13878.n158 a_n2982_13878.t30 3.61217
R15026 a_n2982_13878.n158 a_n2982_13878.t56 3.61217
R15027 a_n2982_13878.n159 a_n2982_13878.t38 3.61217
R15028 a_n2982_13878.n159 a_n2982_13878.t58 3.61217
R15029 a_n2982_13878.n93 a_n2982_13878.t28 3.61217
R15030 a_n2982_13878.n93 a_n2982_13878.t22 3.61217
R15031 a_n2982_13878.n92 a_n2982_13878.t14 3.61217
R15032 a_n2982_13878.n92 a_n2982_13878.t36 3.61217
R15033 a_n2982_13878.n91 a_n2982_13878.t52 3.61217
R15034 a_n2982_13878.n91 a_n2982_13878.t44 3.61217
R15035 a_n2982_13878.n90 a_n2982_13878.t54 3.61217
R15036 a_n2982_13878.n90 a_n2982_13878.t40 3.61217
R15037 a_n2982_13878.n89 a_n2982_13878.t20 3.61217
R15038 a_n2982_13878.n89 a_n2982_13878.t48 3.61217
R15039 a_n2982_13878.n145 a_n2982_13878.t5 2.82907
R15040 a_n2982_13878.n145 a_n2982_13878.t65 2.82907
R15041 a_n2982_13878.n146 a_n2982_13878.t3 2.82907
R15042 a_n2982_13878.n146 a_n2982_13878.t0 2.82907
R15043 a_n2982_13878.n147 a_n2982_13878.t8 2.82907
R15044 a_n2982_13878.n147 a_n2982_13878.t68 2.82907
R15045 a_n2982_13878.n144 a_n2982_13878.t9 2.82907
R15046 a_n2982_13878.n144 a_n2982_13878.t69 2.82907
R15047 a_n2982_13878.n143 a_n2982_13878.t63 2.82907
R15048 a_n2982_13878.n143 a_n2982_13878.t4 2.82907
R15049 a_n2982_13878.n142 a_n2982_13878.t1 2.82907
R15050 a_n2982_13878.n142 a_n2982_13878.t6 2.82907
R15051 a_n2982_13878.n139 a_n2982_13878.t66 2.82907
R15052 a_n2982_13878.n139 a_n2982_13878.t60 2.82907
R15053 a_n2982_13878.n140 a_n2982_13878.t70 2.82907
R15054 a_n2982_13878.n140 a_n2982_13878.t7 2.82907
R15055 a_n2982_13878.n141 a_n2982_13878.t67 2.82907
R15056 a_n2982_13878.n141 a_n2982_13878.t71 2.82907
R15057 a_n2982_13878.n138 a_n2982_13878.t59 2.82907
R15058 a_n2982_13878.n138 a_n2982_13878.t64 2.82907
R15059 a_n2982_13878.n137 a_n2982_13878.t61 2.82907
R15060 a_n2982_13878.n137 a_n2982_13878.t62 2.82907
R15061 a_n2982_13878.n136 a_n2982_13878.t2 2.82907
R15062 a_n2982_13878.n136 a_n2982_13878.t10 2.82907
R15063 a_n2982_13878.n31 a_n2982_13878.n134 14.1668
R15064 a_n2982_13878.n128 a_n2982_13878.n58 22.3251
R15065 a_n2982_13878.n38 a_n2982_13878.n153 14.1668
R15066 a_n2982_13878.n108 a_n2982_13878.n19 14.1668
R15067 a_n2982_13878.n74 a_n2982_13878.n113 22.3251
R15068 a_n2982_13878.n102 a_n2982_13878.n25 14.1668
R15069 a_n2982_13878.n66 a_n2982_13878.n107 22.3251
R15070 a_n2982_13878.n154 a_n2982_13878.n11 1.30542
R15071 a_n2982_13878.n8 a_n2982_13878.n9 1.04595
R15072 a_n2982_13878.n55 a_n2982_13878.n129 47.835
R15073 a_n2982_13878.n49 a_n2982_13878.n148 47.835
R15074 a_n2982_13878.n112 a_n2982_13878.n71 47.835
R15075 a_n2982_13878.n106 a_n2982_13878.n63 47.835
R15076 a_n2982_13878.n0 a_n2982_13878.n4 1.3324
R15077 a_n2982_13878.n27 a_n2982_13878.n26 1.13686
R15078 a_n2982_13878.n21 a_n2982_13878.n20 1.13686
R15079 a_n2982_13878.n15 a_n2982_13878.n14 1.13686
R15080 a_n2982_13878.n32 a_n2982_13878.n34 1.09898
R15081 a_n2982_13878.n43 a_n2982_13878.n42 1.07378
R15082 a_n2982_13878.n40 a_n2982_13878.n39 1.07378
R15083 a_n2982_13878.n2 a_n2982_13878.n3 0.888431
R15084 a_n2982_13878.n2 a_n2982_13878.n1 0.888431
R15085 a_n2982_13878.n37 a_n2982_13878.n36 0.758076
R15086 a_n2982_13878.n37 a_n2982_13878.n35 0.758076
R15087 a_n2982_13878.n35 a_n2982_13878.n34 0.758076
R15088 a_n2982_13878.n30 a_n2982_13878.n29 0.758076
R15089 a_n2982_13878.n30 a_n2982_13878.n28 0.758076
R15090 a_n2982_13878.n28 a_n2982_13878.n27 0.758076
R15091 a_n2982_13878.n23 a_n2982_13878.n24 0.758076
R15092 a_n2982_13878.n22 a_n2982_13878.n23 0.758076
R15093 a_n2982_13878.n20 a_n2982_13878.n22 0.758076
R15094 a_n2982_13878.n17 a_n2982_13878.n18 0.758076
R15095 a_n2982_13878.n16 a_n2982_13878.n17 0.758076
R15096 a_n2982_13878.n14 a_n2982_13878.n16 0.758076
R15097 a_n2982_13878.n13 a_n2982_13878.n12 0.758076
R15098 a_n2982_13878.n10 a_n2982_13878.n9 0.758076
R15099 a_n2982_13878.n8 a_n2982_13878.n7 0.758076
R15100 a_n2982_13878.n6 a_n2982_13878.n5 0.758076
R15101 a_n2982_13878.n42 a_n2982_13878.n44 0.716017
R15102 a_n2982_13878.n41 a_n2982_13878.n40 0.716017
R15103 a_n2982_13878.n10 a_n2982_13878.n12 0.67853
R15104 a_n2982_13878.n6 a_n2982_13878.n7 0.67853
R15105 a_n2804_13878.n29 a_n2804_13878.n28 98.9632
R15106 a_n2804_13878.n2 a_n2804_13878.n0 98.7517
R15107 a_n2804_13878.n22 a_n2804_13878.n21 98.6055
R15108 a_n2804_13878.n24 a_n2804_13878.n23 98.6055
R15109 a_n2804_13878.n26 a_n2804_13878.n25 98.6055
R15110 a_n2804_13878.n28 a_n2804_13878.n27 98.6055
R15111 a_n2804_13878.n10 a_n2804_13878.n9 98.6055
R15112 a_n2804_13878.n8 a_n2804_13878.n7 98.6055
R15113 a_n2804_13878.n6 a_n2804_13878.n5 98.6055
R15114 a_n2804_13878.n4 a_n2804_13878.n3 98.6055
R15115 a_n2804_13878.n2 a_n2804_13878.n1 98.6055
R15116 a_n2804_13878.n20 a_n2804_13878.n19 98.6054
R15117 a_n2804_13878.n12 a_n2804_13878.t30 74.6477
R15118 a_n2804_13878.n17 a_n2804_13878.t31 74.2899
R15119 a_n2804_13878.n14 a_n2804_13878.t26 74.2899
R15120 a_n2804_13878.n13 a_n2804_13878.t27 74.2899
R15121 a_n2804_13878.n16 a_n2804_13878.n15 70.6783
R15122 a_n2804_13878.n12 a_n2804_13878.n11 70.6783
R15123 a_n2804_13878.n18 a_n2804_13878.n10 15.7159
R15124 a_n2804_13878.n20 a_n2804_13878.n18 12.6495
R15125 a_n2804_13878.n18 a_n2804_13878.n17 8.38735
R15126 a_n2804_13878.n19 a_n2804_13878.t8 3.61217
R15127 a_n2804_13878.n19 a_n2804_13878.t17 3.61217
R15128 a_n2804_13878.n21 a_n2804_13878.t21 3.61217
R15129 a_n2804_13878.n21 a_n2804_13878.t7 3.61217
R15130 a_n2804_13878.n23 a_n2804_13878.t11 3.61217
R15131 a_n2804_13878.n23 a_n2804_13878.t12 3.61217
R15132 a_n2804_13878.n25 a_n2804_13878.t22 3.61217
R15133 a_n2804_13878.n25 a_n2804_13878.t23 3.61217
R15134 a_n2804_13878.n27 a_n2804_13878.t1 3.61217
R15135 a_n2804_13878.n27 a_n2804_13878.t13 3.61217
R15136 a_n2804_13878.n15 a_n2804_13878.t28 3.61217
R15137 a_n2804_13878.n15 a_n2804_13878.t25 3.61217
R15138 a_n2804_13878.n11 a_n2804_13878.t0 3.61217
R15139 a_n2804_13878.n11 a_n2804_13878.t29 3.61217
R15140 a_n2804_13878.n9 a_n2804_13878.t14 3.61217
R15141 a_n2804_13878.n9 a_n2804_13878.t2 3.61217
R15142 a_n2804_13878.n7 a_n2804_13878.t19 3.61217
R15143 a_n2804_13878.n7 a_n2804_13878.t4 3.61217
R15144 a_n2804_13878.n5 a_n2804_13878.t3 3.61217
R15145 a_n2804_13878.n5 a_n2804_13878.t6 3.61217
R15146 a_n2804_13878.n3 a_n2804_13878.t16 3.61217
R15147 a_n2804_13878.n3 a_n2804_13878.t9 3.61217
R15148 a_n2804_13878.n1 a_n2804_13878.t20 3.61217
R15149 a_n2804_13878.n1 a_n2804_13878.t10 3.61217
R15150 a_n2804_13878.n0 a_n2804_13878.t5 3.61217
R15151 a_n2804_13878.n0 a_n2804_13878.t15 3.61217
R15152 a_n2804_13878.n29 a_n2804_13878.t18 3.61217
R15153 a_n2804_13878.t24 a_n2804_13878.n29 3.61217
R15154 a_n2804_13878.n13 a_n2804_13878.n12 0.358259
R15155 a_n2804_13878.n16 a_n2804_13878.n14 0.358259
R15156 a_n2804_13878.n17 a_n2804_13878.n16 0.358259
R15157 a_n2804_13878.n28 a_n2804_13878.n26 0.358259
R15158 a_n2804_13878.n26 a_n2804_13878.n24 0.358259
R15159 a_n2804_13878.n24 a_n2804_13878.n22 0.358259
R15160 a_n2804_13878.n22 a_n2804_13878.n20 0.358259
R15161 a_n2804_13878.n4 a_n2804_13878.n2 0.146627
R15162 a_n2804_13878.n6 a_n2804_13878.n4 0.146627
R15163 a_n2804_13878.n8 a_n2804_13878.n6 0.146627
R15164 a_n2804_13878.n10 a_n2804_13878.n8 0.146627
R15165 a_n2804_13878.n14 a_n2804_13878.n13 0.101793
R15166 vdd.n303 vdd.n267 756.745
R15167 vdd.n252 vdd.n216 756.745
R15168 vdd.n209 vdd.n173 756.745
R15169 vdd.n158 vdd.n122 756.745
R15170 vdd.n116 vdd.n80 756.745
R15171 vdd.n65 vdd.n29 756.745
R15172 vdd.n1953 vdd.n1917 756.745
R15173 vdd.n2004 vdd.n1968 756.745
R15174 vdd.n1859 vdd.n1823 756.745
R15175 vdd.n1910 vdd.n1874 756.745
R15176 vdd.n1766 vdd.n1730 756.745
R15177 vdd.n1817 vdd.n1781 756.745
R15178 vdd.n1143 vdd.t164 640.208
R15179 vdd.n838 vdd.t209 640.208
R15180 vdd.n1147 vdd.t206 640.208
R15181 vdd.n829 vdd.t233 640.208
R15182 vdd.n724 vdd.t186 640.208
R15183 vdd.n2535 vdd.t227 640.208
R15184 vdd.n661 vdd.t175 640.208
R15185 vdd.n2532 vdd.t216 640.208
R15186 vdd.n625 vdd.t160 640.208
R15187 vdd.n899 vdd.t223 640.208
R15188 vdd.n1565 vdd.t196 592.009
R15189 vdd.n1602 vdd.t220 592.009
R15190 vdd.n1476 vdd.t230 592.009
R15191 vdd.n2074 vdd.t190 592.009
R15192 vdd.n1076 vdd.t168 592.009
R15193 vdd.n1036 vdd.t172 592.009
R15194 vdd.n3293 vdd.t193 592.009
R15195 vdd.n427 vdd.t182 592.009
R15196 vdd.n387 vdd.t200 592.009
R15197 vdd.n580 vdd.t203 592.009
R15198 vdd.n543 vdd.t213 592.009
R15199 vdd.n3080 vdd.t178 592.009
R15200 vdd.n304 vdd.n303 585
R15201 vdd.n302 vdd.n269 585
R15202 vdd.n301 vdd.n300 585
R15203 vdd.n272 vdd.n270 585
R15204 vdd.n295 vdd.n294 585
R15205 vdd.n293 vdd.n292 585
R15206 vdd.n276 vdd.n275 585
R15207 vdd.n287 vdd.n286 585
R15208 vdd.n285 vdd.n284 585
R15209 vdd.n280 vdd.n279 585
R15210 vdd.n253 vdd.n252 585
R15211 vdd.n251 vdd.n218 585
R15212 vdd.n250 vdd.n249 585
R15213 vdd.n221 vdd.n219 585
R15214 vdd.n244 vdd.n243 585
R15215 vdd.n242 vdd.n241 585
R15216 vdd.n225 vdd.n224 585
R15217 vdd.n236 vdd.n235 585
R15218 vdd.n234 vdd.n233 585
R15219 vdd.n229 vdd.n228 585
R15220 vdd.n210 vdd.n209 585
R15221 vdd.n208 vdd.n175 585
R15222 vdd.n207 vdd.n206 585
R15223 vdd.n178 vdd.n176 585
R15224 vdd.n201 vdd.n200 585
R15225 vdd.n199 vdd.n198 585
R15226 vdd.n182 vdd.n181 585
R15227 vdd.n193 vdd.n192 585
R15228 vdd.n191 vdd.n190 585
R15229 vdd.n186 vdd.n185 585
R15230 vdd.n159 vdd.n158 585
R15231 vdd.n157 vdd.n124 585
R15232 vdd.n156 vdd.n155 585
R15233 vdd.n127 vdd.n125 585
R15234 vdd.n150 vdd.n149 585
R15235 vdd.n148 vdd.n147 585
R15236 vdd.n131 vdd.n130 585
R15237 vdd.n142 vdd.n141 585
R15238 vdd.n140 vdd.n139 585
R15239 vdd.n135 vdd.n134 585
R15240 vdd.n117 vdd.n116 585
R15241 vdd.n115 vdd.n82 585
R15242 vdd.n114 vdd.n113 585
R15243 vdd.n85 vdd.n83 585
R15244 vdd.n108 vdd.n107 585
R15245 vdd.n106 vdd.n105 585
R15246 vdd.n89 vdd.n88 585
R15247 vdd.n100 vdd.n99 585
R15248 vdd.n98 vdd.n97 585
R15249 vdd.n93 vdd.n92 585
R15250 vdd.n66 vdd.n65 585
R15251 vdd.n64 vdd.n31 585
R15252 vdd.n63 vdd.n62 585
R15253 vdd.n34 vdd.n32 585
R15254 vdd.n57 vdd.n56 585
R15255 vdd.n55 vdd.n54 585
R15256 vdd.n38 vdd.n37 585
R15257 vdd.n49 vdd.n48 585
R15258 vdd.n47 vdd.n46 585
R15259 vdd.n42 vdd.n41 585
R15260 vdd.n1954 vdd.n1953 585
R15261 vdd.n1952 vdd.n1919 585
R15262 vdd.n1951 vdd.n1950 585
R15263 vdd.n1922 vdd.n1920 585
R15264 vdd.n1945 vdd.n1944 585
R15265 vdd.n1943 vdd.n1942 585
R15266 vdd.n1926 vdd.n1925 585
R15267 vdd.n1937 vdd.n1936 585
R15268 vdd.n1935 vdd.n1934 585
R15269 vdd.n1930 vdd.n1929 585
R15270 vdd.n2005 vdd.n2004 585
R15271 vdd.n2003 vdd.n1970 585
R15272 vdd.n2002 vdd.n2001 585
R15273 vdd.n1973 vdd.n1971 585
R15274 vdd.n1996 vdd.n1995 585
R15275 vdd.n1994 vdd.n1993 585
R15276 vdd.n1977 vdd.n1976 585
R15277 vdd.n1988 vdd.n1987 585
R15278 vdd.n1986 vdd.n1985 585
R15279 vdd.n1981 vdd.n1980 585
R15280 vdd.n1860 vdd.n1859 585
R15281 vdd.n1858 vdd.n1825 585
R15282 vdd.n1857 vdd.n1856 585
R15283 vdd.n1828 vdd.n1826 585
R15284 vdd.n1851 vdd.n1850 585
R15285 vdd.n1849 vdd.n1848 585
R15286 vdd.n1832 vdd.n1831 585
R15287 vdd.n1843 vdd.n1842 585
R15288 vdd.n1841 vdd.n1840 585
R15289 vdd.n1836 vdd.n1835 585
R15290 vdd.n1911 vdd.n1910 585
R15291 vdd.n1909 vdd.n1876 585
R15292 vdd.n1908 vdd.n1907 585
R15293 vdd.n1879 vdd.n1877 585
R15294 vdd.n1902 vdd.n1901 585
R15295 vdd.n1900 vdd.n1899 585
R15296 vdd.n1883 vdd.n1882 585
R15297 vdd.n1894 vdd.n1893 585
R15298 vdd.n1892 vdd.n1891 585
R15299 vdd.n1887 vdd.n1886 585
R15300 vdd.n1767 vdd.n1766 585
R15301 vdd.n1765 vdd.n1732 585
R15302 vdd.n1764 vdd.n1763 585
R15303 vdd.n1735 vdd.n1733 585
R15304 vdd.n1758 vdd.n1757 585
R15305 vdd.n1756 vdd.n1755 585
R15306 vdd.n1739 vdd.n1738 585
R15307 vdd.n1750 vdd.n1749 585
R15308 vdd.n1748 vdd.n1747 585
R15309 vdd.n1743 vdd.n1742 585
R15310 vdd.n1818 vdd.n1817 585
R15311 vdd.n1816 vdd.n1783 585
R15312 vdd.n1815 vdd.n1814 585
R15313 vdd.n1786 vdd.n1784 585
R15314 vdd.n1809 vdd.n1808 585
R15315 vdd.n1807 vdd.n1806 585
R15316 vdd.n1790 vdd.n1789 585
R15317 vdd.n1801 vdd.n1800 585
R15318 vdd.n1799 vdd.n1798 585
R15319 vdd.n1794 vdd.n1793 585
R15320 vdd.n3409 vdd.n352 488.781
R15321 vdd.n3291 vdd.n350 488.781
R15322 vdd.n3213 vdd.n515 488.781
R15323 vdd.n3211 vdd.n517 488.781
R15324 vdd.n2069 vdd.n1358 488.781
R15325 vdd.n2072 vdd.n2071 488.781
R15326 vdd.n1671 vdd.n1436 488.781
R15327 vdd.n1669 vdd.n1439 488.781
R15328 vdd.n281 vdd.t73 329.043
R15329 vdd.n230 vdd.t152 329.043
R15330 vdd.n187 vdd.t154 329.043
R15331 vdd.n136 vdd.t146 329.043
R15332 vdd.n94 vdd.t97 329.043
R15333 vdd.n43 vdd.t113 329.043
R15334 vdd.n1931 vdd.t101 329.043
R15335 vdd.n1982 vdd.t107 329.043
R15336 vdd.n1837 vdd.t90 329.043
R15337 vdd.n1888 vdd.t95 329.043
R15338 vdd.n1744 vdd.t114 329.043
R15339 vdd.n1795 vdd.t96 329.043
R15340 vdd.n1565 vdd.t199 319.788
R15341 vdd.n1602 vdd.t222 319.788
R15342 vdd.n1476 vdd.t232 319.788
R15343 vdd.n2074 vdd.t191 319.788
R15344 vdd.n1076 vdd.t170 319.788
R15345 vdd.n1036 vdd.t173 319.788
R15346 vdd.n3293 vdd.t194 319.788
R15347 vdd.n427 vdd.t184 319.788
R15348 vdd.n387 vdd.t201 319.788
R15349 vdd.n580 vdd.t205 319.788
R15350 vdd.n543 vdd.t215 319.788
R15351 vdd.n3080 vdd.t181 319.788
R15352 vdd.n1566 vdd.t198 303.69
R15353 vdd.n1603 vdd.t221 303.69
R15354 vdd.n1477 vdd.t231 303.69
R15355 vdd.n2075 vdd.t192 303.69
R15356 vdd.n1077 vdd.t171 303.69
R15357 vdd.n1037 vdd.t174 303.69
R15358 vdd.n3294 vdd.t195 303.69
R15359 vdd.n428 vdd.t185 303.69
R15360 vdd.n388 vdd.t202 303.69
R15361 vdd.n581 vdd.t204 303.69
R15362 vdd.n544 vdd.t214 303.69
R15363 vdd.n3081 vdd.t180 303.69
R15364 vdd.n2802 vdd.n788 279.512
R15365 vdd.n3042 vdd.n635 279.512
R15366 vdd.n2979 vdd.n632 279.512
R15367 vdd.n2734 vdd.n2733 279.512
R15368 vdd.n2495 vdd.n826 279.512
R15369 vdd.n2426 vdd.n2425 279.512
R15370 vdd.n1183 vdd.n1182 279.512
R15371 vdd.n2220 vdd.n966 279.512
R15372 vdd.n2958 vdd.n633 279.512
R15373 vdd.n3045 vdd.n3044 279.512
R15374 vdd.n2607 vdd.n2530 279.512
R15375 vdd.n2538 vdd.n784 279.512
R15376 vdd.n2423 vdd.n836 279.512
R15377 vdd.n834 vdd.n808 279.512
R15378 vdd.n1308 vdd.n1003 279.512
R15379 vdd.n1108 vdd.n961 279.512
R15380 vdd.n2218 vdd.n969 254.619
R15381 vdd.n613 vdd.n516 254.619
R15382 vdd.n2960 vdd.n633 185
R15383 vdd.n3043 vdd.n633 185
R15384 vdd.n2962 vdd.n2961 185
R15385 vdd.n2961 vdd.n631 185
R15386 vdd.n2963 vdd.n667 185
R15387 vdd.n2973 vdd.n667 185
R15388 vdd.n2964 vdd.n676 185
R15389 vdd.n676 vdd.n674 185
R15390 vdd.n2966 vdd.n2965 185
R15391 vdd.n2967 vdd.n2966 185
R15392 vdd.n2919 vdd.n675 185
R15393 vdd.n675 vdd.n671 185
R15394 vdd.n2918 vdd.n2917 185
R15395 vdd.n2917 vdd.n2916 185
R15396 vdd.n678 vdd.n677 185
R15397 vdd.n679 vdd.n678 185
R15398 vdd.n2909 vdd.n2908 185
R15399 vdd.n2910 vdd.n2909 185
R15400 vdd.n2907 vdd.n687 185
R15401 vdd.n692 vdd.n687 185
R15402 vdd.n2906 vdd.n2905 185
R15403 vdd.n2905 vdd.n2904 185
R15404 vdd.n689 vdd.n688 185
R15405 vdd.n698 vdd.n689 185
R15406 vdd.n2897 vdd.n2896 185
R15407 vdd.n2898 vdd.n2897 185
R15408 vdd.n2895 vdd.n699 185
R15409 vdd.n705 vdd.n699 185
R15410 vdd.n2894 vdd.n2893 185
R15411 vdd.n2893 vdd.n2892 185
R15412 vdd.n701 vdd.n700 185
R15413 vdd.n702 vdd.n701 185
R15414 vdd.n2885 vdd.n2884 185
R15415 vdd.n2886 vdd.n2885 185
R15416 vdd.n2883 vdd.n712 185
R15417 vdd.n712 vdd.n709 185
R15418 vdd.n2882 vdd.n2881 185
R15419 vdd.n2881 vdd.n2880 185
R15420 vdd.n714 vdd.n713 185
R15421 vdd.n715 vdd.n714 185
R15422 vdd.n2873 vdd.n2872 185
R15423 vdd.n2874 vdd.n2873 185
R15424 vdd.n2871 vdd.n723 185
R15425 vdd.n729 vdd.n723 185
R15426 vdd.n2870 vdd.n2869 185
R15427 vdd.n2869 vdd.n2868 185
R15428 vdd.n2859 vdd.n726 185
R15429 vdd.n736 vdd.n726 185
R15430 vdd.n2861 vdd.n2860 185
R15431 vdd.n2862 vdd.n2861 185
R15432 vdd.n2858 vdd.n737 185
R15433 vdd.n737 vdd.n733 185
R15434 vdd.n2857 vdd.n2856 185
R15435 vdd.n2856 vdd.n2855 185
R15436 vdd.n739 vdd.n738 185
R15437 vdd.n740 vdd.n739 185
R15438 vdd.n2848 vdd.n2847 185
R15439 vdd.n2849 vdd.n2848 185
R15440 vdd.n2846 vdd.n748 185
R15441 vdd.n753 vdd.n748 185
R15442 vdd.n2845 vdd.n2844 185
R15443 vdd.n2844 vdd.n2843 185
R15444 vdd.n750 vdd.n749 185
R15445 vdd.n759 vdd.n750 185
R15446 vdd.n2836 vdd.n2835 185
R15447 vdd.n2837 vdd.n2836 185
R15448 vdd.n2834 vdd.n760 185
R15449 vdd.n2710 vdd.n760 185
R15450 vdd.n2833 vdd.n2832 185
R15451 vdd.n2832 vdd.n2831 185
R15452 vdd.n762 vdd.n761 185
R15453 vdd.n2716 vdd.n762 185
R15454 vdd.n2824 vdd.n2823 185
R15455 vdd.n2825 vdd.n2824 185
R15456 vdd.n2822 vdd.n771 185
R15457 vdd.n771 vdd.n768 185
R15458 vdd.n2821 vdd.n2820 185
R15459 vdd.n2820 vdd.n2819 185
R15460 vdd.n773 vdd.n772 185
R15461 vdd.n774 vdd.n773 185
R15462 vdd.n2812 vdd.n2811 185
R15463 vdd.n2813 vdd.n2812 185
R15464 vdd.n2810 vdd.n782 185
R15465 vdd.n2728 vdd.n782 185
R15466 vdd.n2809 vdd.n2808 185
R15467 vdd.n2808 vdd.n2807 185
R15468 vdd.n784 vdd.n783 185
R15469 vdd.n785 vdd.n784 185
R15470 vdd.n2539 vdd.n2538 185
R15471 vdd.n2541 vdd.n2540 185
R15472 vdd.n2543 vdd.n2542 185
R15473 vdd.n2545 vdd.n2544 185
R15474 vdd.n2547 vdd.n2546 185
R15475 vdd.n2549 vdd.n2548 185
R15476 vdd.n2551 vdd.n2550 185
R15477 vdd.n2553 vdd.n2552 185
R15478 vdd.n2555 vdd.n2554 185
R15479 vdd.n2557 vdd.n2556 185
R15480 vdd.n2559 vdd.n2558 185
R15481 vdd.n2561 vdd.n2560 185
R15482 vdd.n2563 vdd.n2562 185
R15483 vdd.n2565 vdd.n2564 185
R15484 vdd.n2567 vdd.n2566 185
R15485 vdd.n2569 vdd.n2568 185
R15486 vdd.n2571 vdd.n2570 185
R15487 vdd.n2573 vdd.n2572 185
R15488 vdd.n2575 vdd.n2574 185
R15489 vdd.n2577 vdd.n2576 185
R15490 vdd.n2579 vdd.n2578 185
R15491 vdd.n2581 vdd.n2580 185
R15492 vdd.n2583 vdd.n2582 185
R15493 vdd.n2585 vdd.n2584 185
R15494 vdd.n2587 vdd.n2586 185
R15495 vdd.n2589 vdd.n2588 185
R15496 vdd.n2591 vdd.n2590 185
R15497 vdd.n2593 vdd.n2592 185
R15498 vdd.n2595 vdd.n2594 185
R15499 vdd.n2597 vdd.n2596 185
R15500 vdd.n2599 vdd.n2598 185
R15501 vdd.n2601 vdd.n2600 185
R15502 vdd.n2603 vdd.n2602 185
R15503 vdd.n2605 vdd.n2604 185
R15504 vdd.n2606 vdd.n2530 185
R15505 vdd.n2800 vdd.n2530 185
R15506 vdd.n3046 vdd.n3045 185
R15507 vdd.n3047 vdd.n624 185
R15508 vdd.n3049 vdd.n3048 185
R15509 vdd.n3051 vdd.n622 185
R15510 vdd.n3053 vdd.n3052 185
R15511 vdd.n3054 vdd.n621 185
R15512 vdd.n3056 vdd.n3055 185
R15513 vdd.n3058 vdd.n619 185
R15514 vdd.n3060 vdd.n3059 185
R15515 vdd.n3061 vdd.n618 185
R15516 vdd.n3063 vdd.n3062 185
R15517 vdd.n3065 vdd.n616 185
R15518 vdd.n3067 vdd.n3066 185
R15519 vdd.n3068 vdd.n615 185
R15520 vdd.n3070 vdd.n3069 185
R15521 vdd.n3072 vdd.n614 185
R15522 vdd.n3073 vdd.n611 185
R15523 vdd.n3076 vdd.n3075 185
R15524 vdd.n612 vdd.n610 185
R15525 vdd.n2932 vdd.n2931 185
R15526 vdd.n2934 vdd.n2933 185
R15527 vdd.n2936 vdd.n2928 185
R15528 vdd.n2938 vdd.n2937 185
R15529 vdd.n2939 vdd.n2927 185
R15530 vdd.n2941 vdd.n2940 185
R15531 vdd.n2943 vdd.n2925 185
R15532 vdd.n2945 vdd.n2944 185
R15533 vdd.n2946 vdd.n2924 185
R15534 vdd.n2948 vdd.n2947 185
R15535 vdd.n2950 vdd.n2922 185
R15536 vdd.n2952 vdd.n2951 185
R15537 vdd.n2953 vdd.n2921 185
R15538 vdd.n2955 vdd.n2954 185
R15539 vdd.n2957 vdd.n2920 185
R15540 vdd.n2959 vdd.n2958 185
R15541 vdd.n2958 vdd.n613 185
R15542 vdd.n3044 vdd.n628 185
R15543 vdd.n3044 vdd.n3043 185
R15544 vdd.n2661 vdd.n630 185
R15545 vdd.n631 vdd.n630 185
R15546 vdd.n2662 vdd.n666 185
R15547 vdd.n2973 vdd.n666 185
R15548 vdd.n2664 vdd.n2663 185
R15549 vdd.n2663 vdd.n674 185
R15550 vdd.n2665 vdd.n673 185
R15551 vdd.n2967 vdd.n673 185
R15552 vdd.n2667 vdd.n2666 185
R15553 vdd.n2666 vdd.n671 185
R15554 vdd.n2668 vdd.n681 185
R15555 vdd.n2916 vdd.n681 185
R15556 vdd.n2670 vdd.n2669 185
R15557 vdd.n2669 vdd.n679 185
R15558 vdd.n2671 vdd.n686 185
R15559 vdd.n2910 vdd.n686 185
R15560 vdd.n2673 vdd.n2672 185
R15561 vdd.n2672 vdd.n692 185
R15562 vdd.n2674 vdd.n691 185
R15563 vdd.n2904 vdd.n691 185
R15564 vdd.n2676 vdd.n2675 185
R15565 vdd.n2675 vdd.n698 185
R15566 vdd.n2677 vdd.n697 185
R15567 vdd.n2898 vdd.n697 185
R15568 vdd.n2679 vdd.n2678 185
R15569 vdd.n2678 vdd.n705 185
R15570 vdd.n2680 vdd.n704 185
R15571 vdd.n2892 vdd.n704 185
R15572 vdd.n2682 vdd.n2681 185
R15573 vdd.n2681 vdd.n702 185
R15574 vdd.n2683 vdd.n711 185
R15575 vdd.n2886 vdd.n711 185
R15576 vdd.n2685 vdd.n2684 185
R15577 vdd.n2684 vdd.n709 185
R15578 vdd.n2686 vdd.n717 185
R15579 vdd.n2880 vdd.n717 185
R15580 vdd.n2688 vdd.n2687 185
R15581 vdd.n2687 vdd.n715 185
R15582 vdd.n2689 vdd.n722 185
R15583 vdd.n2874 vdd.n722 185
R15584 vdd.n2691 vdd.n2690 185
R15585 vdd.n2690 vdd.n729 185
R15586 vdd.n2692 vdd.n728 185
R15587 vdd.n2868 vdd.n728 185
R15588 vdd.n2694 vdd.n2693 185
R15589 vdd.n2693 vdd.n736 185
R15590 vdd.n2695 vdd.n735 185
R15591 vdd.n2862 vdd.n735 185
R15592 vdd.n2697 vdd.n2696 185
R15593 vdd.n2696 vdd.n733 185
R15594 vdd.n2698 vdd.n742 185
R15595 vdd.n2855 vdd.n742 185
R15596 vdd.n2700 vdd.n2699 185
R15597 vdd.n2699 vdd.n740 185
R15598 vdd.n2701 vdd.n747 185
R15599 vdd.n2849 vdd.n747 185
R15600 vdd.n2703 vdd.n2702 185
R15601 vdd.n2702 vdd.n753 185
R15602 vdd.n2704 vdd.n752 185
R15603 vdd.n2843 vdd.n752 185
R15604 vdd.n2706 vdd.n2705 185
R15605 vdd.n2705 vdd.n759 185
R15606 vdd.n2707 vdd.n758 185
R15607 vdd.n2837 vdd.n758 185
R15608 vdd.n2709 vdd.n2708 185
R15609 vdd.n2710 vdd.n2709 185
R15610 vdd.n2610 vdd.n764 185
R15611 vdd.n2831 vdd.n764 185
R15612 vdd.n2718 vdd.n2717 185
R15613 vdd.n2717 vdd.n2716 185
R15614 vdd.n2719 vdd.n770 185
R15615 vdd.n2825 vdd.n770 185
R15616 vdd.n2721 vdd.n2720 185
R15617 vdd.n2720 vdd.n768 185
R15618 vdd.n2722 vdd.n776 185
R15619 vdd.n2819 vdd.n776 185
R15620 vdd.n2724 vdd.n2723 185
R15621 vdd.n2723 vdd.n774 185
R15622 vdd.n2725 vdd.n781 185
R15623 vdd.n2813 vdd.n781 185
R15624 vdd.n2727 vdd.n2726 185
R15625 vdd.n2728 vdd.n2727 185
R15626 vdd.n2609 vdd.n787 185
R15627 vdd.n2807 vdd.n787 185
R15628 vdd.n2608 vdd.n2607 185
R15629 vdd.n2607 vdd.n785 185
R15630 vdd.n2069 vdd.n2068 185
R15631 vdd.n2070 vdd.n2069 185
R15632 vdd.n1359 vdd.n1357 185
R15633 vdd.n2061 vdd.n1357 185
R15634 vdd.n2064 vdd.n2063 185
R15635 vdd.n2063 vdd.n2062 185
R15636 vdd.n1362 vdd.n1361 185
R15637 vdd.n1363 vdd.n1362 185
R15638 vdd.n2050 vdd.n2049 185
R15639 vdd.n2051 vdd.n2050 185
R15640 vdd.n1371 vdd.n1370 185
R15641 vdd.n2042 vdd.n1370 185
R15642 vdd.n2045 vdd.n2044 185
R15643 vdd.n2044 vdd.n2043 185
R15644 vdd.n1374 vdd.n1373 185
R15645 vdd.n1380 vdd.n1374 185
R15646 vdd.n2033 vdd.n2032 185
R15647 vdd.n2034 vdd.n2033 185
R15648 vdd.n1382 vdd.n1381 185
R15649 vdd.n2025 vdd.n1381 185
R15650 vdd.n2028 vdd.n2027 185
R15651 vdd.n2027 vdd.n2026 185
R15652 vdd.n1385 vdd.n1384 185
R15653 vdd.n1386 vdd.n1385 185
R15654 vdd.n2016 vdd.n2015 185
R15655 vdd.n2017 vdd.n2016 185
R15656 vdd.n1394 vdd.n1393 185
R15657 vdd.n1393 vdd.n1392 185
R15658 vdd.n1729 vdd.n1728 185
R15659 vdd.n1728 vdd.n1727 185
R15660 vdd.n1397 vdd.n1396 185
R15661 vdd.n1403 vdd.n1397 185
R15662 vdd.n1718 vdd.n1717 185
R15663 vdd.n1719 vdd.n1718 185
R15664 vdd.n1405 vdd.n1404 185
R15665 vdd.n1710 vdd.n1404 185
R15666 vdd.n1713 vdd.n1712 185
R15667 vdd.n1712 vdd.n1711 185
R15668 vdd.n1408 vdd.n1407 185
R15669 vdd.n1415 vdd.n1408 185
R15670 vdd.n1701 vdd.n1700 185
R15671 vdd.n1702 vdd.n1701 185
R15672 vdd.n1417 vdd.n1416 185
R15673 vdd.n1416 vdd.n1414 185
R15674 vdd.n1696 vdd.n1695 185
R15675 vdd.n1695 vdd.n1694 185
R15676 vdd.n1420 vdd.n1419 185
R15677 vdd.n1421 vdd.n1420 185
R15678 vdd.n1685 vdd.n1684 185
R15679 vdd.n1686 vdd.n1685 185
R15680 vdd.n1429 vdd.n1428 185
R15681 vdd.n1428 vdd.n1427 185
R15682 vdd.n1680 vdd.n1679 185
R15683 vdd.n1679 vdd.n1678 185
R15684 vdd.n1432 vdd.n1431 185
R15685 vdd.n1438 vdd.n1432 185
R15686 vdd.n1669 vdd.n1668 185
R15687 vdd.n1670 vdd.n1669 185
R15688 vdd.n1665 vdd.n1439 185
R15689 vdd.n1664 vdd.n1442 185
R15690 vdd.n1663 vdd.n1443 185
R15691 vdd.n1443 vdd.n1437 185
R15692 vdd.n1446 vdd.n1444 185
R15693 vdd.n1659 vdd.n1448 185
R15694 vdd.n1658 vdd.n1449 185
R15695 vdd.n1657 vdd.n1451 185
R15696 vdd.n1454 vdd.n1452 185
R15697 vdd.n1653 vdd.n1456 185
R15698 vdd.n1652 vdd.n1457 185
R15699 vdd.n1651 vdd.n1459 185
R15700 vdd.n1462 vdd.n1460 185
R15701 vdd.n1647 vdd.n1464 185
R15702 vdd.n1646 vdd.n1465 185
R15703 vdd.n1645 vdd.n1467 185
R15704 vdd.n1470 vdd.n1468 185
R15705 vdd.n1641 vdd.n1472 185
R15706 vdd.n1640 vdd.n1473 185
R15707 vdd.n1639 vdd.n1475 185
R15708 vdd.n1480 vdd.n1478 185
R15709 vdd.n1635 vdd.n1482 185
R15710 vdd.n1634 vdd.n1483 185
R15711 vdd.n1633 vdd.n1485 185
R15712 vdd.n1488 vdd.n1486 185
R15713 vdd.n1629 vdd.n1490 185
R15714 vdd.n1628 vdd.n1491 185
R15715 vdd.n1627 vdd.n1493 185
R15716 vdd.n1496 vdd.n1494 185
R15717 vdd.n1623 vdd.n1498 185
R15718 vdd.n1622 vdd.n1499 185
R15719 vdd.n1621 vdd.n1501 185
R15720 vdd.n1504 vdd.n1502 185
R15721 vdd.n1617 vdd.n1506 185
R15722 vdd.n1616 vdd.n1507 185
R15723 vdd.n1615 vdd.n1509 185
R15724 vdd.n1512 vdd.n1510 185
R15725 vdd.n1611 vdd.n1514 185
R15726 vdd.n1610 vdd.n1515 185
R15727 vdd.n1609 vdd.n1517 185
R15728 vdd.n1520 vdd.n1518 185
R15729 vdd.n1605 vdd.n1522 185
R15730 vdd.n1604 vdd.n1601 185
R15731 vdd.n1599 vdd.n1523 185
R15732 vdd.n1598 vdd.n1597 185
R15733 vdd.n1528 vdd.n1525 185
R15734 vdd.n1593 vdd.n1529 185
R15735 vdd.n1592 vdd.n1531 185
R15736 vdd.n1591 vdd.n1532 185
R15737 vdd.n1536 vdd.n1533 185
R15738 vdd.n1587 vdd.n1537 185
R15739 vdd.n1586 vdd.n1539 185
R15740 vdd.n1585 vdd.n1540 185
R15741 vdd.n1544 vdd.n1541 185
R15742 vdd.n1581 vdd.n1545 185
R15743 vdd.n1580 vdd.n1547 185
R15744 vdd.n1579 vdd.n1548 185
R15745 vdd.n1552 vdd.n1549 185
R15746 vdd.n1575 vdd.n1553 185
R15747 vdd.n1574 vdd.n1555 185
R15748 vdd.n1573 vdd.n1556 185
R15749 vdd.n1560 vdd.n1557 185
R15750 vdd.n1569 vdd.n1561 185
R15751 vdd.n1568 vdd.n1563 185
R15752 vdd.n1564 vdd.n1436 185
R15753 vdd.n1437 vdd.n1436 185
R15754 vdd.n2073 vdd.n2072 185
R15755 vdd.n2077 vdd.n1353 185
R15756 vdd.n1352 vdd.n1346 185
R15757 vdd.n1350 vdd.n1349 185
R15758 vdd.n1348 vdd.n1107 185
R15759 vdd.n2081 vdd.n1104 185
R15760 vdd.n2083 vdd.n2082 185
R15761 vdd.n2085 vdd.n1102 185
R15762 vdd.n2087 vdd.n2086 185
R15763 vdd.n2088 vdd.n1097 185
R15764 vdd.n2090 vdd.n2089 185
R15765 vdd.n2092 vdd.n1095 185
R15766 vdd.n2094 vdd.n2093 185
R15767 vdd.n2095 vdd.n1090 185
R15768 vdd.n2097 vdd.n2096 185
R15769 vdd.n2099 vdd.n1088 185
R15770 vdd.n2101 vdd.n2100 185
R15771 vdd.n2102 vdd.n1084 185
R15772 vdd.n2104 vdd.n2103 185
R15773 vdd.n2106 vdd.n1081 185
R15774 vdd.n2108 vdd.n2107 185
R15775 vdd.n1082 vdd.n1075 185
R15776 vdd.n2112 vdd.n1079 185
R15777 vdd.n2113 vdd.n1071 185
R15778 vdd.n2115 vdd.n2114 185
R15779 vdd.n2117 vdd.n1069 185
R15780 vdd.n2119 vdd.n2118 185
R15781 vdd.n2120 vdd.n1064 185
R15782 vdd.n2122 vdd.n2121 185
R15783 vdd.n2124 vdd.n1062 185
R15784 vdd.n2126 vdd.n2125 185
R15785 vdd.n2127 vdd.n1057 185
R15786 vdd.n2129 vdd.n2128 185
R15787 vdd.n2131 vdd.n1055 185
R15788 vdd.n2133 vdd.n2132 185
R15789 vdd.n2134 vdd.n1050 185
R15790 vdd.n2136 vdd.n2135 185
R15791 vdd.n2138 vdd.n1048 185
R15792 vdd.n2140 vdd.n2139 185
R15793 vdd.n2141 vdd.n1044 185
R15794 vdd.n2143 vdd.n2142 185
R15795 vdd.n2145 vdd.n1041 185
R15796 vdd.n2147 vdd.n2146 185
R15797 vdd.n1042 vdd.n1035 185
R15798 vdd.n2151 vdd.n1039 185
R15799 vdd.n2152 vdd.n1031 185
R15800 vdd.n2154 vdd.n2153 185
R15801 vdd.n2156 vdd.n1029 185
R15802 vdd.n2158 vdd.n2157 185
R15803 vdd.n2159 vdd.n1024 185
R15804 vdd.n2161 vdd.n2160 185
R15805 vdd.n2163 vdd.n1022 185
R15806 vdd.n2165 vdd.n2164 185
R15807 vdd.n2166 vdd.n1017 185
R15808 vdd.n2168 vdd.n2167 185
R15809 vdd.n2170 vdd.n1015 185
R15810 vdd.n2172 vdd.n2171 185
R15811 vdd.n2173 vdd.n1013 185
R15812 vdd.n2175 vdd.n2174 185
R15813 vdd.n2178 vdd.n2177 185
R15814 vdd.n2180 vdd.n2179 185
R15815 vdd.n2182 vdd.n1011 185
R15816 vdd.n2184 vdd.n2183 185
R15817 vdd.n1358 vdd.n1010 185
R15818 vdd.n2071 vdd.n1356 185
R15819 vdd.n2071 vdd.n2070 185
R15820 vdd.n1366 vdd.n1355 185
R15821 vdd.n2061 vdd.n1355 185
R15822 vdd.n2060 vdd.n2059 185
R15823 vdd.n2062 vdd.n2060 185
R15824 vdd.n1365 vdd.n1364 185
R15825 vdd.n1364 vdd.n1363 185
R15826 vdd.n2053 vdd.n2052 185
R15827 vdd.n2052 vdd.n2051 185
R15828 vdd.n1369 vdd.n1368 185
R15829 vdd.n2042 vdd.n1369 185
R15830 vdd.n2041 vdd.n2040 185
R15831 vdd.n2043 vdd.n2041 185
R15832 vdd.n1376 vdd.n1375 185
R15833 vdd.n1380 vdd.n1375 185
R15834 vdd.n2036 vdd.n2035 185
R15835 vdd.n2035 vdd.n2034 185
R15836 vdd.n1379 vdd.n1378 185
R15837 vdd.n2025 vdd.n1379 185
R15838 vdd.n2024 vdd.n2023 185
R15839 vdd.n2026 vdd.n2024 185
R15840 vdd.n1388 vdd.n1387 185
R15841 vdd.n1387 vdd.n1386 185
R15842 vdd.n2019 vdd.n2018 185
R15843 vdd.n2018 vdd.n2017 185
R15844 vdd.n1391 vdd.n1390 185
R15845 vdd.n1392 vdd.n1391 185
R15846 vdd.n1726 vdd.n1725 185
R15847 vdd.n1727 vdd.n1726 185
R15848 vdd.n1399 vdd.n1398 185
R15849 vdd.n1403 vdd.n1398 185
R15850 vdd.n1721 vdd.n1720 185
R15851 vdd.n1720 vdd.n1719 185
R15852 vdd.n1402 vdd.n1401 185
R15853 vdd.n1710 vdd.n1402 185
R15854 vdd.n1709 vdd.n1708 185
R15855 vdd.n1711 vdd.n1709 185
R15856 vdd.n1410 vdd.n1409 185
R15857 vdd.n1415 vdd.n1409 185
R15858 vdd.n1704 vdd.n1703 185
R15859 vdd.n1703 vdd.n1702 185
R15860 vdd.n1413 vdd.n1412 185
R15861 vdd.n1414 vdd.n1413 185
R15862 vdd.n1693 vdd.n1692 185
R15863 vdd.n1694 vdd.n1693 185
R15864 vdd.n1423 vdd.n1422 185
R15865 vdd.n1422 vdd.n1421 185
R15866 vdd.n1688 vdd.n1687 185
R15867 vdd.n1687 vdd.n1686 185
R15868 vdd.n1426 vdd.n1425 185
R15869 vdd.n1427 vdd.n1426 185
R15870 vdd.n1677 vdd.n1676 185
R15871 vdd.n1678 vdd.n1677 185
R15872 vdd.n1434 vdd.n1433 185
R15873 vdd.n1438 vdd.n1433 185
R15874 vdd.n1672 vdd.n1671 185
R15875 vdd.n1671 vdd.n1670 185
R15876 vdd.n828 vdd.n826 185
R15877 vdd.n2424 vdd.n826 185
R15878 vdd.n2346 vdd.n846 185
R15879 vdd.n846 vdd.n833 185
R15880 vdd.n2348 vdd.n2347 185
R15881 vdd.n2349 vdd.n2348 185
R15882 vdd.n2345 vdd.n845 185
R15883 vdd.n1227 vdd.n845 185
R15884 vdd.n2344 vdd.n2343 185
R15885 vdd.n2343 vdd.n2342 185
R15886 vdd.n848 vdd.n847 185
R15887 vdd.n849 vdd.n848 185
R15888 vdd.n2333 vdd.n2332 185
R15889 vdd.n2334 vdd.n2333 185
R15890 vdd.n2331 vdd.n859 185
R15891 vdd.n859 vdd.n856 185
R15892 vdd.n2330 vdd.n2329 185
R15893 vdd.n2329 vdd.n2328 185
R15894 vdd.n861 vdd.n860 185
R15895 vdd.n1253 vdd.n861 185
R15896 vdd.n2321 vdd.n2320 185
R15897 vdd.n2322 vdd.n2321 185
R15898 vdd.n2319 vdd.n869 185
R15899 vdd.n874 vdd.n869 185
R15900 vdd.n2318 vdd.n2317 185
R15901 vdd.n2317 vdd.n2316 185
R15902 vdd.n871 vdd.n870 185
R15903 vdd.n880 vdd.n871 185
R15904 vdd.n2309 vdd.n2308 185
R15905 vdd.n2310 vdd.n2309 185
R15906 vdd.n2307 vdd.n881 185
R15907 vdd.n1265 vdd.n881 185
R15908 vdd.n2306 vdd.n2305 185
R15909 vdd.n2305 vdd.n2304 185
R15910 vdd.n883 vdd.n882 185
R15911 vdd.n884 vdd.n883 185
R15912 vdd.n2297 vdd.n2296 185
R15913 vdd.n2298 vdd.n2297 185
R15914 vdd.n2295 vdd.n893 185
R15915 vdd.n893 vdd.n890 185
R15916 vdd.n2294 vdd.n2293 185
R15917 vdd.n2293 vdd.n2292 185
R15918 vdd.n895 vdd.n894 185
R15919 vdd.n904 vdd.n895 185
R15920 vdd.n2284 vdd.n2283 185
R15921 vdd.n2285 vdd.n2284 185
R15922 vdd.n2282 vdd.n905 185
R15923 vdd.n911 vdd.n905 185
R15924 vdd.n2281 vdd.n2280 185
R15925 vdd.n2280 vdd.n2279 185
R15926 vdd.n907 vdd.n906 185
R15927 vdd.n908 vdd.n907 185
R15928 vdd.n2272 vdd.n2271 185
R15929 vdd.n2273 vdd.n2272 185
R15930 vdd.n2270 vdd.n918 185
R15931 vdd.n918 vdd.n915 185
R15932 vdd.n2269 vdd.n2268 185
R15933 vdd.n2268 vdd.n2267 185
R15934 vdd.n920 vdd.n919 185
R15935 vdd.n921 vdd.n920 185
R15936 vdd.n2260 vdd.n2259 185
R15937 vdd.n2261 vdd.n2260 185
R15938 vdd.n2258 vdd.n929 185
R15939 vdd.n934 vdd.n929 185
R15940 vdd.n2257 vdd.n2256 185
R15941 vdd.n2256 vdd.n2255 185
R15942 vdd.n931 vdd.n930 185
R15943 vdd.n940 vdd.n931 185
R15944 vdd.n2248 vdd.n2247 185
R15945 vdd.n2249 vdd.n2248 185
R15946 vdd.n2246 vdd.n941 185
R15947 vdd.n947 vdd.n941 185
R15948 vdd.n2245 vdd.n2244 185
R15949 vdd.n2244 vdd.n2243 185
R15950 vdd.n943 vdd.n942 185
R15951 vdd.n944 vdd.n943 185
R15952 vdd.n2236 vdd.n2235 185
R15953 vdd.n2237 vdd.n2236 185
R15954 vdd.n2234 vdd.n954 185
R15955 vdd.n954 vdd.n951 185
R15956 vdd.n2233 vdd.n2232 185
R15957 vdd.n2232 vdd.n2231 185
R15958 vdd.n956 vdd.n955 185
R15959 vdd.n965 vdd.n956 185
R15960 vdd.n2224 vdd.n2223 185
R15961 vdd.n2225 vdd.n2224 185
R15962 vdd.n2222 vdd.n966 185
R15963 vdd.n966 vdd.n962 185
R15964 vdd.n2221 vdd.n2220 185
R15965 vdd.n968 vdd.n967 185
R15966 vdd.n2217 vdd.n2216 185
R15967 vdd.n2218 vdd.n2217 185
R15968 vdd.n2215 vdd.n1004 185
R15969 vdd.n2214 vdd.n2213 185
R15970 vdd.n2212 vdd.n2211 185
R15971 vdd.n2210 vdd.n2209 185
R15972 vdd.n2208 vdd.n2207 185
R15973 vdd.n2206 vdd.n2205 185
R15974 vdd.n2204 vdd.n2203 185
R15975 vdd.n2202 vdd.n2201 185
R15976 vdd.n2200 vdd.n2199 185
R15977 vdd.n2198 vdd.n2197 185
R15978 vdd.n2196 vdd.n2195 185
R15979 vdd.n2194 vdd.n2193 185
R15980 vdd.n2192 vdd.n2191 185
R15981 vdd.n2190 vdd.n2189 185
R15982 vdd.n2188 vdd.n2187 185
R15983 vdd.n1149 vdd.n1005 185
R15984 vdd.n1151 vdd.n1150 185
R15985 vdd.n1153 vdd.n1152 185
R15986 vdd.n1155 vdd.n1154 185
R15987 vdd.n1157 vdd.n1156 185
R15988 vdd.n1159 vdd.n1158 185
R15989 vdd.n1161 vdd.n1160 185
R15990 vdd.n1163 vdd.n1162 185
R15991 vdd.n1165 vdd.n1164 185
R15992 vdd.n1167 vdd.n1166 185
R15993 vdd.n1169 vdd.n1168 185
R15994 vdd.n1171 vdd.n1170 185
R15995 vdd.n1173 vdd.n1172 185
R15996 vdd.n1175 vdd.n1174 185
R15997 vdd.n1178 vdd.n1177 185
R15998 vdd.n1180 vdd.n1179 185
R15999 vdd.n1182 vdd.n1181 185
R16000 vdd.n2427 vdd.n2426 185
R16001 vdd.n2429 vdd.n2428 185
R16002 vdd.n2431 vdd.n2430 185
R16003 vdd.n2434 vdd.n2433 185
R16004 vdd.n2436 vdd.n2435 185
R16005 vdd.n2438 vdd.n2437 185
R16006 vdd.n2440 vdd.n2439 185
R16007 vdd.n2442 vdd.n2441 185
R16008 vdd.n2444 vdd.n2443 185
R16009 vdd.n2446 vdd.n2445 185
R16010 vdd.n2448 vdd.n2447 185
R16011 vdd.n2450 vdd.n2449 185
R16012 vdd.n2452 vdd.n2451 185
R16013 vdd.n2454 vdd.n2453 185
R16014 vdd.n2456 vdd.n2455 185
R16015 vdd.n2458 vdd.n2457 185
R16016 vdd.n2460 vdd.n2459 185
R16017 vdd.n2462 vdd.n2461 185
R16018 vdd.n2464 vdd.n2463 185
R16019 vdd.n2466 vdd.n2465 185
R16020 vdd.n2468 vdd.n2467 185
R16021 vdd.n2470 vdd.n2469 185
R16022 vdd.n2472 vdd.n2471 185
R16023 vdd.n2474 vdd.n2473 185
R16024 vdd.n2476 vdd.n2475 185
R16025 vdd.n2478 vdd.n2477 185
R16026 vdd.n2480 vdd.n2479 185
R16027 vdd.n2482 vdd.n2481 185
R16028 vdd.n2484 vdd.n2483 185
R16029 vdd.n2486 vdd.n2485 185
R16030 vdd.n2488 vdd.n2487 185
R16031 vdd.n2490 vdd.n2489 185
R16032 vdd.n2492 vdd.n2491 185
R16033 vdd.n2493 vdd.n827 185
R16034 vdd.n2495 vdd.n2494 185
R16035 vdd.n2496 vdd.n2495 185
R16036 vdd.n2425 vdd.n831 185
R16037 vdd.n2425 vdd.n2424 185
R16038 vdd.n1225 vdd.n832 185
R16039 vdd.n833 vdd.n832 185
R16040 vdd.n1226 vdd.n843 185
R16041 vdd.n2349 vdd.n843 185
R16042 vdd.n1229 vdd.n1228 185
R16043 vdd.n1228 vdd.n1227 185
R16044 vdd.n1230 vdd.n850 185
R16045 vdd.n2342 vdd.n850 185
R16046 vdd.n1232 vdd.n1231 185
R16047 vdd.n1231 vdd.n849 185
R16048 vdd.n1233 vdd.n857 185
R16049 vdd.n2334 vdd.n857 185
R16050 vdd.n1235 vdd.n1234 185
R16051 vdd.n1234 vdd.n856 185
R16052 vdd.n1236 vdd.n862 185
R16053 vdd.n2328 vdd.n862 185
R16054 vdd.n1255 vdd.n1254 185
R16055 vdd.n1254 vdd.n1253 185
R16056 vdd.n1256 vdd.n867 185
R16057 vdd.n2322 vdd.n867 185
R16058 vdd.n1258 vdd.n1257 185
R16059 vdd.n1257 vdd.n874 185
R16060 vdd.n1259 vdd.n872 185
R16061 vdd.n2316 vdd.n872 185
R16062 vdd.n1261 vdd.n1260 185
R16063 vdd.n1260 vdd.n880 185
R16064 vdd.n1262 vdd.n878 185
R16065 vdd.n2310 vdd.n878 185
R16066 vdd.n1264 vdd.n1263 185
R16067 vdd.n1265 vdd.n1264 185
R16068 vdd.n1224 vdd.n885 185
R16069 vdd.n2304 vdd.n885 185
R16070 vdd.n1223 vdd.n1222 185
R16071 vdd.n1222 vdd.n884 185
R16072 vdd.n1221 vdd.n891 185
R16073 vdd.n2298 vdd.n891 185
R16074 vdd.n1220 vdd.n1219 185
R16075 vdd.n1219 vdd.n890 185
R16076 vdd.n1218 vdd.n896 185
R16077 vdd.n2292 vdd.n896 185
R16078 vdd.n1217 vdd.n1216 185
R16079 vdd.n1216 vdd.n904 185
R16080 vdd.n1215 vdd.n902 185
R16081 vdd.n2285 vdd.n902 185
R16082 vdd.n1214 vdd.n1213 185
R16083 vdd.n1213 vdd.n911 185
R16084 vdd.n1212 vdd.n909 185
R16085 vdd.n2279 vdd.n909 185
R16086 vdd.n1211 vdd.n1210 185
R16087 vdd.n1210 vdd.n908 185
R16088 vdd.n1209 vdd.n916 185
R16089 vdd.n2273 vdd.n916 185
R16090 vdd.n1208 vdd.n1207 185
R16091 vdd.n1207 vdd.n915 185
R16092 vdd.n1206 vdd.n922 185
R16093 vdd.n2267 vdd.n922 185
R16094 vdd.n1205 vdd.n1204 185
R16095 vdd.n1204 vdd.n921 185
R16096 vdd.n1203 vdd.n927 185
R16097 vdd.n2261 vdd.n927 185
R16098 vdd.n1202 vdd.n1201 185
R16099 vdd.n1201 vdd.n934 185
R16100 vdd.n1200 vdd.n932 185
R16101 vdd.n2255 vdd.n932 185
R16102 vdd.n1199 vdd.n1198 185
R16103 vdd.n1198 vdd.n940 185
R16104 vdd.n1197 vdd.n938 185
R16105 vdd.n2249 vdd.n938 185
R16106 vdd.n1196 vdd.n1195 185
R16107 vdd.n1195 vdd.n947 185
R16108 vdd.n1194 vdd.n945 185
R16109 vdd.n2243 vdd.n945 185
R16110 vdd.n1193 vdd.n1192 185
R16111 vdd.n1192 vdd.n944 185
R16112 vdd.n1191 vdd.n952 185
R16113 vdd.n2237 vdd.n952 185
R16114 vdd.n1190 vdd.n1189 185
R16115 vdd.n1189 vdd.n951 185
R16116 vdd.n1188 vdd.n957 185
R16117 vdd.n2231 vdd.n957 185
R16118 vdd.n1187 vdd.n1186 185
R16119 vdd.n1186 vdd.n965 185
R16120 vdd.n1185 vdd.n963 185
R16121 vdd.n2225 vdd.n963 185
R16122 vdd.n1184 vdd.n1183 185
R16123 vdd.n1183 vdd.n962 185
R16124 vdd.n3409 vdd.n3408 185
R16125 vdd.n3410 vdd.n3409 185
R16126 vdd.n347 vdd.n346 185
R16127 vdd.n3411 vdd.n347 185
R16128 vdd.n3414 vdd.n3413 185
R16129 vdd.n3413 vdd.n3412 185
R16130 vdd.n3415 vdd.n341 185
R16131 vdd.n341 vdd.n340 185
R16132 vdd.n3417 vdd.n3416 185
R16133 vdd.n3418 vdd.n3417 185
R16134 vdd.n336 vdd.n335 185
R16135 vdd.n3419 vdd.n336 185
R16136 vdd.n3422 vdd.n3421 185
R16137 vdd.n3421 vdd.n3420 185
R16138 vdd.n3423 vdd.n330 185
R16139 vdd.n330 vdd.n329 185
R16140 vdd.n3425 vdd.n3424 185
R16141 vdd.n3426 vdd.n3425 185
R16142 vdd.n324 vdd.n323 185
R16143 vdd.n3427 vdd.n324 185
R16144 vdd.n3430 vdd.n3429 185
R16145 vdd.n3429 vdd.n3428 185
R16146 vdd.n3431 vdd.n319 185
R16147 vdd.n325 vdd.n319 185
R16148 vdd.n3433 vdd.n3432 185
R16149 vdd.n3434 vdd.n3433 185
R16150 vdd.n315 vdd.n313 185
R16151 vdd.n3435 vdd.n315 185
R16152 vdd.n3438 vdd.n3437 185
R16153 vdd.n3437 vdd.n3436 185
R16154 vdd.n314 vdd.n312 185
R16155 vdd.n481 vdd.n314 185
R16156 vdd.n3260 vdd.n3259 185
R16157 vdd.n3261 vdd.n3260 185
R16158 vdd.n483 vdd.n482 185
R16159 vdd.n3252 vdd.n482 185
R16160 vdd.n3255 vdd.n3254 185
R16161 vdd.n3254 vdd.n3253 185
R16162 vdd.n486 vdd.n485 185
R16163 vdd.n493 vdd.n486 185
R16164 vdd.n3243 vdd.n3242 185
R16165 vdd.n3244 vdd.n3243 185
R16166 vdd.n495 vdd.n494 185
R16167 vdd.n494 vdd.n492 185
R16168 vdd.n3238 vdd.n3237 185
R16169 vdd.n3237 vdd.n3236 185
R16170 vdd.n498 vdd.n497 185
R16171 vdd.n499 vdd.n498 185
R16172 vdd.n3227 vdd.n3226 185
R16173 vdd.n3228 vdd.n3227 185
R16174 vdd.n507 vdd.n506 185
R16175 vdd.n506 vdd.n505 185
R16176 vdd.n3222 vdd.n3221 185
R16177 vdd.n3221 vdd.n3220 185
R16178 vdd.n510 vdd.n509 185
R16179 vdd.n511 vdd.n510 185
R16180 vdd.n3211 vdd.n3210 185
R16181 vdd.n3212 vdd.n3211 185
R16182 vdd.n3207 vdd.n517 185
R16183 vdd.n3206 vdd.n3205 185
R16184 vdd.n3203 vdd.n519 185
R16185 vdd.n3203 vdd.n516 185
R16186 vdd.n3202 vdd.n3201 185
R16187 vdd.n3200 vdd.n3199 185
R16188 vdd.n3198 vdd.n3197 185
R16189 vdd.n3196 vdd.n3195 185
R16190 vdd.n3194 vdd.n525 185
R16191 vdd.n3192 vdd.n3191 185
R16192 vdd.n3190 vdd.n526 185
R16193 vdd.n3189 vdd.n3188 185
R16194 vdd.n3186 vdd.n531 185
R16195 vdd.n3184 vdd.n3183 185
R16196 vdd.n3182 vdd.n532 185
R16197 vdd.n3181 vdd.n3180 185
R16198 vdd.n3178 vdd.n537 185
R16199 vdd.n3176 vdd.n3175 185
R16200 vdd.n3174 vdd.n538 185
R16201 vdd.n3173 vdd.n3172 185
R16202 vdd.n3170 vdd.n545 185
R16203 vdd.n3168 vdd.n3167 185
R16204 vdd.n3166 vdd.n546 185
R16205 vdd.n3165 vdd.n3164 185
R16206 vdd.n3162 vdd.n551 185
R16207 vdd.n3160 vdd.n3159 185
R16208 vdd.n3158 vdd.n552 185
R16209 vdd.n3157 vdd.n3156 185
R16210 vdd.n3154 vdd.n557 185
R16211 vdd.n3152 vdd.n3151 185
R16212 vdd.n3150 vdd.n558 185
R16213 vdd.n3149 vdd.n3148 185
R16214 vdd.n3146 vdd.n563 185
R16215 vdd.n3144 vdd.n3143 185
R16216 vdd.n3142 vdd.n564 185
R16217 vdd.n3141 vdd.n3140 185
R16218 vdd.n3138 vdd.n569 185
R16219 vdd.n3136 vdd.n3135 185
R16220 vdd.n3134 vdd.n570 185
R16221 vdd.n3133 vdd.n3132 185
R16222 vdd.n3130 vdd.n575 185
R16223 vdd.n3128 vdd.n3127 185
R16224 vdd.n3126 vdd.n576 185
R16225 vdd.n585 vdd.n579 185
R16226 vdd.n3122 vdd.n3121 185
R16227 vdd.n3119 vdd.n583 185
R16228 vdd.n3118 vdd.n3117 185
R16229 vdd.n3116 vdd.n3115 185
R16230 vdd.n3114 vdd.n589 185
R16231 vdd.n3112 vdd.n3111 185
R16232 vdd.n3110 vdd.n590 185
R16233 vdd.n3109 vdd.n3108 185
R16234 vdd.n3106 vdd.n595 185
R16235 vdd.n3104 vdd.n3103 185
R16236 vdd.n3102 vdd.n596 185
R16237 vdd.n3101 vdd.n3100 185
R16238 vdd.n3098 vdd.n601 185
R16239 vdd.n3096 vdd.n3095 185
R16240 vdd.n3094 vdd.n602 185
R16241 vdd.n3093 vdd.n3092 185
R16242 vdd.n3090 vdd.n3089 185
R16243 vdd.n3088 vdd.n3087 185
R16244 vdd.n3086 vdd.n3085 185
R16245 vdd.n3084 vdd.n3083 185
R16246 vdd.n3079 vdd.n515 185
R16247 vdd.n516 vdd.n515 185
R16248 vdd.n3292 vdd.n3291 185
R16249 vdd.n3296 vdd.n462 185
R16250 vdd.n3298 vdd.n3297 185
R16251 vdd.n3300 vdd.n460 185
R16252 vdd.n3302 vdd.n3301 185
R16253 vdd.n3303 vdd.n455 185
R16254 vdd.n3305 vdd.n3304 185
R16255 vdd.n3307 vdd.n453 185
R16256 vdd.n3309 vdd.n3308 185
R16257 vdd.n3310 vdd.n448 185
R16258 vdd.n3312 vdd.n3311 185
R16259 vdd.n3314 vdd.n446 185
R16260 vdd.n3316 vdd.n3315 185
R16261 vdd.n3317 vdd.n441 185
R16262 vdd.n3319 vdd.n3318 185
R16263 vdd.n3321 vdd.n439 185
R16264 vdd.n3323 vdd.n3322 185
R16265 vdd.n3324 vdd.n435 185
R16266 vdd.n3326 vdd.n3325 185
R16267 vdd.n3328 vdd.n432 185
R16268 vdd.n3330 vdd.n3329 185
R16269 vdd.n433 vdd.n426 185
R16270 vdd.n3334 vdd.n430 185
R16271 vdd.n3335 vdd.n422 185
R16272 vdd.n3337 vdd.n3336 185
R16273 vdd.n3339 vdd.n420 185
R16274 vdd.n3341 vdd.n3340 185
R16275 vdd.n3342 vdd.n415 185
R16276 vdd.n3344 vdd.n3343 185
R16277 vdd.n3346 vdd.n413 185
R16278 vdd.n3348 vdd.n3347 185
R16279 vdd.n3349 vdd.n408 185
R16280 vdd.n3351 vdd.n3350 185
R16281 vdd.n3353 vdd.n406 185
R16282 vdd.n3355 vdd.n3354 185
R16283 vdd.n3356 vdd.n401 185
R16284 vdd.n3358 vdd.n3357 185
R16285 vdd.n3360 vdd.n399 185
R16286 vdd.n3362 vdd.n3361 185
R16287 vdd.n3363 vdd.n395 185
R16288 vdd.n3365 vdd.n3364 185
R16289 vdd.n3367 vdd.n392 185
R16290 vdd.n3369 vdd.n3368 185
R16291 vdd.n393 vdd.n386 185
R16292 vdd.n3373 vdd.n390 185
R16293 vdd.n3374 vdd.n382 185
R16294 vdd.n3376 vdd.n3375 185
R16295 vdd.n3378 vdd.n380 185
R16296 vdd.n3380 vdd.n3379 185
R16297 vdd.n3381 vdd.n375 185
R16298 vdd.n3383 vdd.n3382 185
R16299 vdd.n3385 vdd.n373 185
R16300 vdd.n3387 vdd.n3386 185
R16301 vdd.n3388 vdd.n368 185
R16302 vdd.n3390 vdd.n3389 185
R16303 vdd.n3392 vdd.n366 185
R16304 vdd.n3394 vdd.n3393 185
R16305 vdd.n3395 vdd.n360 185
R16306 vdd.n3397 vdd.n3396 185
R16307 vdd.n3399 vdd.n359 185
R16308 vdd.n3400 vdd.n358 185
R16309 vdd.n3403 vdd.n3402 185
R16310 vdd.n3404 vdd.n356 185
R16311 vdd.n3405 vdd.n352 185
R16312 vdd.n3287 vdd.n350 185
R16313 vdd.n3410 vdd.n350 185
R16314 vdd.n3286 vdd.n349 185
R16315 vdd.n3411 vdd.n349 185
R16316 vdd.n3285 vdd.n348 185
R16317 vdd.n3412 vdd.n348 185
R16318 vdd.n468 vdd.n467 185
R16319 vdd.n467 vdd.n340 185
R16320 vdd.n3281 vdd.n339 185
R16321 vdd.n3418 vdd.n339 185
R16322 vdd.n3280 vdd.n338 185
R16323 vdd.n3419 vdd.n338 185
R16324 vdd.n3279 vdd.n337 185
R16325 vdd.n3420 vdd.n337 185
R16326 vdd.n471 vdd.n470 185
R16327 vdd.n470 vdd.n329 185
R16328 vdd.n3275 vdd.n328 185
R16329 vdd.n3426 vdd.n328 185
R16330 vdd.n3274 vdd.n327 185
R16331 vdd.n3427 vdd.n327 185
R16332 vdd.n3273 vdd.n326 185
R16333 vdd.n3428 vdd.n326 185
R16334 vdd.n474 vdd.n473 185
R16335 vdd.n473 vdd.n325 185
R16336 vdd.n3269 vdd.n318 185
R16337 vdd.n3434 vdd.n318 185
R16338 vdd.n3268 vdd.n317 185
R16339 vdd.n3435 vdd.n317 185
R16340 vdd.n3267 vdd.n316 185
R16341 vdd.n3436 vdd.n316 185
R16342 vdd.n480 vdd.n476 185
R16343 vdd.n481 vdd.n480 185
R16344 vdd.n3263 vdd.n3262 185
R16345 vdd.n3262 vdd.n3261 185
R16346 vdd.n479 vdd.n478 185
R16347 vdd.n3252 vdd.n479 185
R16348 vdd.n3251 vdd.n3250 185
R16349 vdd.n3253 vdd.n3251 185
R16350 vdd.n488 vdd.n487 185
R16351 vdd.n493 vdd.n487 185
R16352 vdd.n3246 vdd.n3245 185
R16353 vdd.n3245 vdd.n3244 185
R16354 vdd.n491 vdd.n490 185
R16355 vdd.n492 vdd.n491 185
R16356 vdd.n3235 vdd.n3234 185
R16357 vdd.n3236 vdd.n3235 185
R16358 vdd.n501 vdd.n500 185
R16359 vdd.n500 vdd.n499 185
R16360 vdd.n3230 vdd.n3229 185
R16361 vdd.n3229 vdd.n3228 185
R16362 vdd.n504 vdd.n503 185
R16363 vdd.n505 vdd.n504 185
R16364 vdd.n3219 vdd.n3218 185
R16365 vdd.n3220 vdd.n3219 185
R16366 vdd.n513 vdd.n512 185
R16367 vdd.n512 vdd.n511 185
R16368 vdd.n3214 vdd.n3213 185
R16369 vdd.n3213 vdd.n3212 185
R16370 vdd.n2803 vdd.n2802 185
R16371 vdd.n790 vdd.n789 185
R16372 vdd.n2799 vdd.n2798 185
R16373 vdd.n2800 vdd.n2799 185
R16374 vdd.n2797 vdd.n2531 185
R16375 vdd.n2796 vdd.n2795 185
R16376 vdd.n2794 vdd.n2793 185
R16377 vdd.n2792 vdd.n2791 185
R16378 vdd.n2790 vdd.n2789 185
R16379 vdd.n2788 vdd.n2787 185
R16380 vdd.n2786 vdd.n2785 185
R16381 vdd.n2784 vdd.n2783 185
R16382 vdd.n2782 vdd.n2781 185
R16383 vdd.n2780 vdd.n2779 185
R16384 vdd.n2778 vdd.n2777 185
R16385 vdd.n2776 vdd.n2775 185
R16386 vdd.n2774 vdd.n2773 185
R16387 vdd.n2772 vdd.n2771 185
R16388 vdd.n2770 vdd.n2769 185
R16389 vdd.n2768 vdd.n2767 185
R16390 vdd.n2766 vdd.n2765 185
R16391 vdd.n2764 vdd.n2763 185
R16392 vdd.n2762 vdd.n2761 185
R16393 vdd.n2760 vdd.n2759 185
R16394 vdd.n2758 vdd.n2757 185
R16395 vdd.n2756 vdd.n2755 185
R16396 vdd.n2754 vdd.n2753 185
R16397 vdd.n2752 vdd.n2751 185
R16398 vdd.n2750 vdd.n2749 185
R16399 vdd.n2748 vdd.n2747 185
R16400 vdd.n2746 vdd.n2745 185
R16401 vdd.n2744 vdd.n2743 185
R16402 vdd.n2742 vdd.n2741 185
R16403 vdd.n2739 vdd.n2738 185
R16404 vdd.n2737 vdd.n2736 185
R16405 vdd.n2735 vdd.n2734 185
R16406 vdd.n2980 vdd.n2979 185
R16407 vdd.n2981 vdd.n660 185
R16408 vdd.n2983 vdd.n2982 185
R16409 vdd.n2985 vdd.n658 185
R16410 vdd.n2987 vdd.n2986 185
R16411 vdd.n2988 vdd.n657 185
R16412 vdd.n2990 vdd.n2989 185
R16413 vdd.n2992 vdd.n655 185
R16414 vdd.n2994 vdd.n2993 185
R16415 vdd.n2995 vdd.n654 185
R16416 vdd.n2997 vdd.n2996 185
R16417 vdd.n2999 vdd.n652 185
R16418 vdd.n3001 vdd.n3000 185
R16419 vdd.n3002 vdd.n651 185
R16420 vdd.n3004 vdd.n3003 185
R16421 vdd.n3006 vdd.n649 185
R16422 vdd.n3008 vdd.n3007 185
R16423 vdd.n3010 vdd.n648 185
R16424 vdd.n3012 vdd.n3011 185
R16425 vdd.n3014 vdd.n646 185
R16426 vdd.n3016 vdd.n3015 185
R16427 vdd.n3017 vdd.n645 185
R16428 vdd.n3019 vdd.n3018 185
R16429 vdd.n3021 vdd.n643 185
R16430 vdd.n3023 vdd.n3022 185
R16431 vdd.n3024 vdd.n642 185
R16432 vdd.n3026 vdd.n3025 185
R16433 vdd.n3028 vdd.n640 185
R16434 vdd.n3030 vdd.n3029 185
R16435 vdd.n3031 vdd.n639 185
R16436 vdd.n3033 vdd.n3032 185
R16437 vdd.n3035 vdd.n638 185
R16438 vdd.n3036 vdd.n637 185
R16439 vdd.n3039 vdd.n3038 185
R16440 vdd.n3040 vdd.n635 185
R16441 vdd.n635 vdd.n613 185
R16442 vdd.n2977 vdd.n632 185
R16443 vdd.n3043 vdd.n632 185
R16444 vdd.n2976 vdd.n2975 185
R16445 vdd.n2975 vdd.n631 185
R16446 vdd.n2974 vdd.n664 185
R16447 vdd.n2974 vdd.n2973 185
R16448 vdd.n2617 vdd.n665 185
R16449 vdd.n674 vdd.n665 185
R16450 vdd.n2618 vdd.n672 185
R16451 vdd.n2967 vdd.n672 185
R16452 vdd.n2620 vdd.n2619 185
R16453 vdd.n2619 vdd.n671 185
R16454 vdd.n2621 vdd.n680 185
R16455 vdd.n2916 vdd.n680 185
R16456 vdd.n2623 vdd.n2622 185
R16457 vdd.n2622 vdd.n679 185
R16458 vdd.n2624 vdd.n685 185
R16459 vdd.n2910 vdd.n685 185
R16460 vdd.n2626 vdd.n2625 185
R16461 vdd.n2625 vdd.n692 185
R16462 vdd.n2627 vdd.n690 185
R16463 vdd.n2904 vdd.n690 185
R16464 vdd.n2629 vdd.n2628 185
R16465 vdd.n2628 vdd.n698 185
R16466 vdd.n2630 vdd.n696 185
R16467 vdd.n2898 vdd.n696 185
R16468 vdd.n2632 vdd.n2631 185
R16469 vdd.n2631 vdd.n705 185
R16470 vdd.n2633 vdd.n703 185
R16471 vdd.n2892 vdd.n703 185
R16472 vdd.n2635 vdd.n2634 185
R16473 vdd.n2634 vdd.n702 185
R16474 vdd.n2636 vdd.n710 185
R16475 vdd.n2886 vdd.n710 185
R16476 vdd.n2638 vdd.n2637 185
R16477 vdd.n2637 vdd.n709 185
R16478 vdd.n2639 vdd.n716 185
R16479 vdd.n2880 vdd.n716 185
R16480 vdd.n2641 vdd.n2640 185
R16481 vdd.n2640 vdd.n715 185
R16482 vdd.n2642 vdd.n721 185
R16483 vdd.n2874 vdd.n721 185
R16484 vdd.n2644 vdd.n2643 185
R16485 vdd.n2643 vdd.n729 185
R16486 vdd.n2645 vdd.n727 185
R16487 vdd.n2868 vdd.n727 185
R16488 vdd.n2647 vdd.n2646 185
R16489 vdd.n2646 vdd.n736 185
R16490 vdd.n2648 vdd.n734 185
R16491 vdd.n2862 vdd.n734 185
R16492 vdd.n2650 vdd.n2649 185
R16493 vdd.n2649 vdd.n733 185
R16494 vdd.n2651 vdd.n741 185
R16495 vdd.n2855 vdd.n741 185
R16496 vdd.n2653 vdd.n2652 185
R16497 vdd.n2652 vdd.n740 185
R16498 vdd.n2654 vdd.n746 185
R16499 vdd.n2849 vdd.n746 185
R16500 vdd.n2656 vdd.n2655 185
R16501 vdd.n2655 vdd.n753 185
R16502 vdd.n2657 vdd.n751 185
R16503 vdd.n2843 vdd.n751 185
R16504 vdd.n2659 vdd.n2658 185
R16505 vdd.n2658 vdd.n759 185
R16506 vdd.n2660 vdd.n757 185
R16507 vdd.n2837 vdd.n757 185
R16508 vdd.n2712 vdd.n2711 185
R16509 vdd.n2711 vdd.n2710 185
R16510 vdd.n2713 vdd.n763 185
R16511 vdd.n2831 vdd.n763 185
R16512 vdd.n2715 vdd.n2714 185
R16513 vdd.n2716 vdd.n2715 185
R16514 vdd.n2616 vdd.n769 185
R16515 vdd.n2825 vdd.n769 185
R16516 vdd.n2615 vdd.n2614 185
R16517 vdd.n2614 vdd.n768 185
R16518 vdd.n2613 vdd.n775 185
R16519 vdd.n2819 vdd.n775 185
R16520 vdd.n2612 vdd.n2611 185
R16521 vdd.n2611 vdd.n774 185
R16522 vdd.n2534 vdd.n780 185
R16523 vdd.n2813 vdd.n780 185
R16524 vdd.n2730 vdd.n2729 185
R16525 vdd.n2729 vdd.n2728 185
R16526 vdd.n2731 vdd.n786 185
R16527 vdd.n2807 vdd.n786 185
R16528 vdd.n2733 vdd.n2732 185
R16529 vdd.n2733 vdd.n785 185
R16530 vdd.n2804 vdd.n788 185
R16531 vdd.n788 vdd.n785 185
R16532 vdd.n2806 vdd.n2805 185
R16533 vdd.n2807 vdd.n2806 185
R16534 vdd.n779 vdd.n778 185
R16535 vdd.n2728 vdd.n779 185
R16536 vdd.n2815 vdd.n2814 185
R16537 vdd.n2814 vdd.n2813 185
R16538 vdd.n2816 vdd.n777 185
R16539 vdd.n777 vdd.n774 185
R16540 vdd.n2818 vdd.n2817 185
R16541 vdd.n2819 vdd.n2818 185
R16542 vdd.n767 vdd.n766 185
R16543 vdd.n768 vdd.n767 185
R16544 vdd.n2827 vdd.n2826 185
R16545 vdd.n2826 vdd.n2825 185
R16546 vdd.n2828 vdd.n765 185
R16547 vdd.n2716 vdd.n765 185
R16548 vdd.n2830 vdd.n2829 185
R16549 vdd.n2831 vdd.n2830 185
R16550 vdd.n756 vdd.n755 185
R16551 vdd.n2710 vdd.n756 185
R16552 vdd.n2839 vdd.n2838 185
R16553 vdd.n2838 vdd.n2837 185
R16554 vdd.n2840 vdd.n754 185
R16555 vdd.n759 vdd.n754 185
R16556 vdd.n2842 vdd.n2841 185
R16557 vdd.n2843 vdd.n2842 185
R16558 vdd.n745 vdd.n744 185
R16559 vdd.n753 vdd.n745 185
R16560 vdd.n2851 vdd.n2850 185
R16561 vdd.n2850 vdd.n2849 185
R16562 vdd.n2852 vdd.n743 185
R16563 vdd.n743 vdd.n740 185
R16564 vdd.n2854 vdd.n2853 185
R16565 vdd.n2855 vdd.n2854 185
R16566 vdd.n732 vdd.n731 185
R16567 vdd.n733 vdd.n732 185
R16568 vdd.n2864 vdd.n2863 185
R16569 vdd.n2863 vdd.n2862 185
R16570 vdd.n2865 vdd.n730 185
R16571 vdd.n736 vdd.n730 185
R16572 vdd.n2867 vdd.n2866 185
R16573 vdd.n2868 vdd.n2867 185
R16574 vdd.n720 vdd.n719 185
R16575 vdd.n729 vdd.n720 185
R16576 vdd.n2876 vdd.n2875 185
R16577 vdd.n2875 vdd.n2874 185
R16578 vdd.n2877 vdd.n718 185
R16579 vdd.n718 vdd.n715 185
R16580 vdd.n2879 vdd.n2878 185
R16581 vdd.n2880 vdd.n2879 185
R16582 vdd.n708 vdd.n707 185
R16583 vdd.n709 vdd.n708 185
R16584 vdd.n2888 vdd.n2887 185
R16585 vdd.n2887 vdd.n2886 185
R16586 vdd.n2889 vdd.n706 185
R16587 vdd.n706 vdd.n702 185
R16588 vdd.n2891 vdd.n2890 185
R16589 vdd.n2892 vdd.n2891 185
R16590 vdd.n695 vdd.n694 185
R16591 vdd.n705 vdd.n695 185
R16592 vdd.n2900 vdd.n2899 185
R16593 vdd.n2899 vdd.n2898 185
R16594 vdd.n2901 vdd.n693 185
R16595 vdd.n698 vdd.n693 185
R16596 vdd.n2903 vdd.n2902 185
R16597 vdd.n2904 vdd.n2903 185
R16598 vdd.n684 vdd.n683 185
R16599 vdd.n692 vdd.n684 185
R16600 vdd.n2912 vdd.n2911 185
R16601 vdd.n2911 vdd.n2910 185
R16602 vdd.n2913 vdd.n682 185
R16603 vdd.n682 vdd.n679 185
R16604 vdd.n2915 vdd.n2914 185
R16605 vdd.n2916 vdd.n2915 185
R16606 vdd.n670 vdd.n669 185
R16607 vdd.n671 vdd.n670 185
R16608 vdd.n2969 vdd.n2968 185
R16609 vdd.n2968 vdd.n2967 185
R16610 vdd.n2970 vdd.n668 185
R16611 vdd.n674 vdd.n668 185
R16612 vdd.n2972 vdd.n2971 185
R16613 vdd.n2973 vdd.n2972 185
R16614 vdd.n636 vdd.n634 185
R16615 vdd.n634 vdd.n631 185
R16616 vdd.n3042 vdd.n3041 185
R16617 vdd.n3043 vdd.n3042 185
R16618 vdd.n2423 vdd.n2422 185
R16619 vdd.n2424 vdd.n2423 185
R16620 vdd.n837 vdd.n835 185
R16621 vdd.n835 vdd.n833 185
R16622 vdd.n2338 vdd.n844 185
R16623 vdd.n2349 vdd.n844 185
R16624 vdd.n2339 vdd.n853 185
R16625 vdd.n1227 vdd.n853 185
R16626 vdd.n2341 vdd.n2340 185
R16627 vdd.n2342 vdd.n2341 185
R16628 vdd.n2337 vdd.n852 185
R16629 vdd.n852 vdd.n849 185
R16630 vdd.n2336 vdd.n2335 185
R16631 vdd.n2335 vdd.n2334 185
R16632 vdd.n855 vdd.n854 185
R16633 vdd.n856 vdd.n855 185
R16634 vdd.n2327 vdd.n2326 185
R16635 vdd.n2328 vdd.n2327 185
R16636 vdd.n2325 vdd.n864 185
R16637 vdd.n1253 vdd.n864 185
R16638 vdd.n2324 vdd.n2323 185
R16639 vdd.n2323 vdd.n2322 185
R16640 vdd.n866 vdd.n865 185
R16641 vdd.n874 vdd.n866 185
R16642 vdd.n2315 vdd.n2314 185
R16643 vdd.n2316 vdd.n2315 185
R16644 vdd.n2313 vdd.n875 185
R16645 vdd.n880 vdd.n875 185
R16646 vdd.n2312 vdd.n2311 185
R16647 vdd.n2311 vdd.n2310 185
R16648 vdd.n877 vdd.n876 185
R16649 vdd.n1265 vdd.n877 185
R16650 vdd.n2303 vdd.n2302 185
R16651 vdd.n2304 vdd.n2303 185
R16652 vdd.n2301 vdd.n887 185
R16653 vdd.n887 vdd.n884 185
R16654 vdd.n2300 vdd.n2299 185
R16655 vdd.n2299 vdd.n2298 185
R16656 vdd.n889 vdd.n888 185
R16657 vdd.n890 vdd.n889 185
R16658 vdd.n2291 vdd.n2290 185
R16659 vdd.n2292 vdd.n2291 185
R16660 vdd.n2288 vdd.n898 185
R16661 vdd.n904 vdd.n898 185
R16662 vdd.n2287 vdd.n2286 185
R16663 vdd.n2286 vdd.n2285 185
R16664 vdd.n901 vdd.n900 185
R16665 vdd.n911 vdd.n901 185
R16666 vdd.n2278 vdd.n2277 185
R16667 vdd.n2279 vdd.n2278 185
R16668 vdd.n2276 vdd.n912 185
R16669 vdd.n912 vdd.n908 185
R16670 vdd.n2275 vdd.n2274 185
R16671 vdd.n2274 vdd.n2273 185
R16672 vdd.n914 vdd.n913 185
R16673 vdd.n915 vdd.n914 185
R16674 vdd.n2266 vdd.n2265 185
R16675 vdd.n2267 vdd.n2266 185
R16676 vdd.n2264 vdd.n924 185
R16677 vdd.n924 vdd.n921 185
R16678 vdd.n2263 vdd.n2262 185
R16679 vdd.n2262 vdd.n2261 185
R16680 vdd.n926 vdd.n925 185
R16681 vdd.n934 vdd.n926 185
R16682 vdd.n2254 vdd.n2253 185
R16683 vdd.n2255 vdd.n2254 185
R16684 vdd.n2252 vdd.n935 185
R16685 vdd.n940 vdd.n935 185
R16686 vdd.n2251 vdd.n2250 185
R16687 vdd.n2250 vdd.n2249 185
R16688 vdd.n937 vdd.n936 185
R16689 vdd.n947 vdd.n937 185
R16690 vdd.n2242 vdd.n2241 185
R16691 vdd.n2243 vdd.n2242 185
R16692 vdd.n2240 vdd.n948 185
R16693 vdd.n948 vdd.n944 185
R16694 vdd.n2239 vdd.n2238 185
R16695 vdd.n2238 vdd.n2237 185
R16696 vdd.n950 vdd.n949 185
R16697 vdd.n951 vdd.n950 185
R16698 vdd.n2230 vdd.n2229 185
R16699 vdd.n2231 vdd.n2230 185
R16700 vdd.n2228 vdd.n959 185
R16701 vdd.n965 vdd.n959 185
R16702 vdd.n2227 vdd.n2226 185
R16703 vdd.n2226 vdd.n2225 185
R16704 vdd.n961 vdd.n960 185
R16705 vdd.n962 vdd.n961 185
R16706 vdd.n2354 vdd.n808 185
R16707 vdd.n2496 vdd.n808 185
R16708 vdd.n2356 vdd.n2355 185
R16709 vdd.n2358 vdd.n2357 185
R16710 vdd.n2360 vdd.n2359 185
R16711 vdd.n2362 vdd.n2361 185
R16712 vdd.n2364 vdd.n2363 185
R16713 vdd.n2366 vdd.n2365 185
R16714 vdd.n2368 vdd.n2367 185
R16715 vdd.n2370 vdd.n2369 185
R16716 vdd.n2372 vdd.n2371 185
R16717 vdd.n2374 vdd.n2373 185
R16718 vdd.n2376 vdd.n2375 185
R16719 vdd.n2378 vdd.n2377 185
R16720 vdd.n2380 vdd.n2379 185
R16721 vdd.n2382 vdd.n2381 185
R16722 vdd.n2384 vdd.n2383 185
R16723 vdd.n2386 vdd.n2385 185
R16724 vdd.n2388 vdd.n2387 185
R16725 vdd.n2390 vdd.n2389 185
R16726 vdd.n2392 vdd.n2391 185
R16727 vdd.n2394 vdd.n2393 185
R16728 vdd.n2396 vdd.n2395 185
R16729 vdd.n2398 vdd.n2397 185
R16730 vdd.n2400 vdd.n2399 185
R16731 vdd.n2402 vdd.n2401 185
R16732 vdd.n2404 vdd.n2403 185
R16733 vdd.n2406 vdd.n2405 185
R16734 vdd.n2408 vdd.n2407 185
R16735 vdd.n2410 vdd.n2409 185
R16736 vdd.n2412 vdd.n2411 185
R16737 vdd.n2414 vdd.n2413 185
R16738 vdd.n2416 vdd.n2415 185
R16739 vdd.n2418 vdd.n2417 185
R16740 vdd.n2420 vdd.n2419 185
R16741 vdd.n2421 vdd.n836 185
R16742 vdd.n2353 vdd.n834 185
R16743 vdd.n2424 vdd.n834 185
R16744 vdd.n2352 vdd.n2351 185
R16745 vdd.n2351 vdd.n833 185
R16746 vdd.n2350 vdd.n841 185
R16747 vdd.n2350 vdd.n2349 185
R16748 vdd.n1243 vdd.n842 185
R16749 vdd.n1227 vdd.n842 185
R16750 vdd.n1244 vdd.n851 185
R16751 vdd.n2342 vdd.n851 185
R16752 vdd.n1246 vdd.n1245 185
R16753 vdd.n1245 vdd.n849 185
R16754 vdd.n1247 vdd.n858 185
R16755 vdd.n2334 vdd.n858 185
R16756 vdd.n1249 vdd.n1248 185
R16757 vdd.n1248 vdd.n856 185
R16758 vdd.n1250 vdd.n863 185
R16759 vdd.n2328 vdd.n863 185
R16760 vdd.n1252 vdd.n1251 185
R16761 vdd.n1253 vdd.n1252 185
R16762 vdd.n1242 vdd.n868 185
R16763 vdd.n2322 vdd.n868 185
R16764 vdd.n1241 vdd.n1240 185
R16765 vdd.n1240 vdd.n874 185
R16766 vdd.n1239 vdd.n873 185
R16767 vdd.n2316 vdd.n873 185
R16768 vdd.n1238 vdd.n1237 185
R16769 vdd.n1237 vdd.n880 185
R16770 vdd.n1146 vdd.n879 185
R16771 vdd.n2310 vdd.n879 185
R16772 vdd.n1267 vdd.n1266 185
R16773 vdd.n1266 vdd.n1265 185
R16774 vdd.n1268 vdd.n886 185
R16775 vdd.n2304 vdd.n886 185
R16776 vdd.n1270 vdd.n1269 185
R16777 vdd.n1269 vdd.n884 185
R16778 vdd.n1271 vdd.n892 185
R16779 vdd.n2298 vdd.n892 185
R16780 vdd.n1273 vdd.n1272 185
R16781 vdd.n1272 vdd.n890 185
R16782 vdd.n1274 vdd.n897 185
R16783 vdd.n2292 vdd.n897 185
R16784 vdd.n1276 vdd.n1275 185
R16785 vdd.n1275 vdd.n904 185
R16786 vdd.n1277 vdd.n903 185
R16787 vdd.n2285 vdd.n903 185
R16788 vdd.n1279 vdd.n1278 185
R16789 vdd.n1278 vdd.n911 185
R16790 vdd.n1280 vdd.n910 185
R16791 vdd.n2279 vdd.n910 185
R16792 vdd.n1282 vdd.n1281 185
R16793 vdd.n1281 vdd.n908 185
R16794 vdd.n1283 vdd.n917 185
R16795 vdd.n2273 vdd.n917 185
R16796 vdd.n1285 vdd.n1284 185
R16797 vdd.n1284 vdd.n915 185
R16798 vdd.n1286 vdd.n923 185
R16799 vdd.n2267 vdd.n923 185
R16800 vdd.n1288 vdd.n1287 185
R16801 vdd.n1287 vdd.n921 185
R16802 vdd.n1289 vdd.n928 185
R16803 vdd.n2261 vdd.n928 185
R16804 vdd.n1291 vdd.n1290 185
R16805 vdd.n1290 vdd.n934 185
R16806 vdd.n1292 vdd.n933 185
R16807 vdd.n2255 vdd.n933 185
R16808 vdd.n1294 vdd.n1293 185
R16809 vdd.n1293 vdd.n940 185
R16810 vdd.n1295 vdd.n939 185
R16811 vdd.n2249 vdd.n939 185
R16812 vdd.n1297 vdd.n1296 185
R16813 vdd.n1296 vdd.n947 185
R16814 vdd.n1298 vdd.n946 185
R16815 vdd.n2243 vdd.n946 185
R16816 vdd.n1300 vdd.n1299 185
R16817 vdd.n1299 vdd.n944 185
R16818 vdd.n1301 vdd.n953 185
R16819 vdd.n2237 vdd.n953 185
R16820 vdd.n1303 vdd.n1302 185
R16821 vdd.n1302 vdd.n951 185
R16822 vdd.n1304 vdd.n958 185
R16823 vdd.n2231 vdd.n958 185
R16824 vdd.n1306 vdd.n1305 185
R16825 vdd.n1305 vdd.n965 185
R16826 vdd.n1307 vdd.n964 185
R16827 vdd.n2225 vdd.n964 185
R16828 vdd.n1309 vdd.n1308 185
R16829 vdd.n1308 vdd.n962 185
R16830 vdd.n1109 vdd.n1108 185
R16831 vdd.n1111 vdd.n1110 185
R16832 vdd.n1113 vdd.n1112 185
R16833 vdd.n1115 vdd.n1114 185
R16834 vdd.n1117 vdd.n1116 185
R16835 vdd.n1119 vdd.n1118 185
R16836 vdd.n1121 vdd.n1120 185
R16837 vdd.n1123 vdd.n1122 185
R16838 vdd.n1125 vdd.n1124 185
R16839 vdd.n1127 vdd.n1126 185
R16840 vdd.n1129 vdd.n1128 185
R16841 vdd.n1131 vdd.n1130 185
R16842 vdd.n1133 vdd.n1132 185
R16843 vdd.n1135 vdd.n1134 185
R16844 vdd.n1137 vdd.n1136 185
R16845 vdd.n1139 vdd.n1138 185
R16846 vdd.n1141 vdd.n1140 185
R16847 vdd.n1343 vdd.n1142 185
R16848 vdd.n1342 vdd.n1341 185
R16849 vdd.n1340 vdd.n1339 185
R16850 vdd.n1338 vdd.n1337 185
R16851 vdd.n1336 vdd.n1335 185
R16852 vdd.n1334 vdd.n1333 185
R16853 vdd.n1332 vdd.n1331 185
R16854 vdd.n1330 vdd.n1329 185
R16855 vdd.n1328 vdd.n1327 185
R16856 vdd.n1326 vdd.n1325 185
R16857 vdd.n1324 vdd.n1323 185
R16858 vdd.n1322 vdd.n1321 185
R16859 vdd.n1320 vdd.n1319 185
R16860 vdd.n1318 vdd.n1317 185
R16861 vdd.n1316 vdd.n1315 185
R16862 vdd.n1314 vdd.n1313 185
R16863 vdd.n1312 vdd.n1311 185
R16864 vdd.n1310 vdd.n1003 185
R16865 vdd.n2218 vdd.n1003 185
R16866 vdd.n303 vdd.n302 171.744
R16867 vdd.n302 vdd.n301 171.744
R16868 vdd.n301 vdd.n270 171.744
R16869 vdd.n294 vdd.n270 171.744
R16870 vdd.n294 vdd.n293 171.744
R16871 vdd.n293 vdd.n275 171.744
R16872 vdd.n286 vdd.n275 171.744
R16873 vdd.n286 vdd.n285 171.744
R16874 vdd.n285 vdd.n279 171.744
R16875 vdd.n252 vdd.n251 171.744
R16876 vdd.n251 vdd.n250 171.744
R16877 vdd.n250 vdd.n219 171.744
R16878 vdd.n243 vdd.n219 171.744
R16879 vdd.n243 vdd.n242 171.744
R16880 vdd.n242 vdd.n224 171.744
R16881 vdd.n235 vdd.n224 171.744
R16882 vdd.n235 vdd.n234 171.744
R16883 vdd.n234 vdd.n228 171.744
R16884 vdd.n209 vdd.n208 171.744
R16885 vdd.n208 vdd.n207 171.744
R16886 vdd.n207 vdd.n176 171.744
R16887 vdd.n200 vdd.n176 171.744
R16888 vdd.n200 vdd.n199 171.744
R16889 vdd.n199 vdd.n181 171.744
R16890 vdd.n192 vdd.n181 171.744
R16891 vdd.n192 vdd.n191 171.744
R16892 vdd.n191 vdd.n185 171.744
R16893 vdd.n158 vdd.n157 171.744
R16894 vdd.n157 vdd.n156 171.744
R16895 vdd.n156 vdd.n125 171.744
R16896 vdd.n149 vdd.n125 171.744
R16897 vdd.n149 vdd.n148 171.744
R16898 vdd.n148 vdd.n130 171.744
R16899 vdd.n141 vdd.n130 171.744
R16900 vdd.n141 vdd.n140 171.744
R16901 vdd.n140 vdd.n134 171.744
R16902 vdd.n116 vdd.n115 171.744
R16903 vdd.n115 vdd.n114 171.744
R16904 vdd.n114 vdd.n83 171.744
R16905 vdd.n107 vdd.n83 171.744
R16906 vdd.n107 vdd.n106 171.744
R16907 vdd.n106 vdd.n88 171.744
R16908 vdd.n99 vdd.n88 171.744
R16909 vdd.n99 vdd.n98 171.744
R16910 vdd.n98 vdd.n92 171.744
R16911 vdd.n65 vdd.n64 171.744
R16912 vdd.n64 vdd.n63 171.744
R16913 vdd.n63 vdd.n32 171.744
R16914 vdd.n56 vdd.n32 171.744
R16915 vdd.n56 vdd.n55 171.744
R16916 vdd.n55 vdd.n37 171.744
R16917 vdd.n48 vdd.n37 171.744
R16918 vdd.n48 vdd.n47 171.744
R16919 vdd.n47 vdd.n41 171.744
R16920 vdd.n1953 vdd.n1952 171.744
R16921 vdd.n1952 vdd.n1951 171.744
R16922 vdd.n1951 vdd.n1920 171.744
R16923 vdd.n1944 vdd.n1920 171.744
R16924 vdd.n1944 vdd.n1943 171.744
R16925 vdd.n1943 vdd.n1925 171.744
R16926 vdd.n1936 vdd.n1925 171.744
R16927 vdd.n1936 vdd.n1935 171.744
R16928 vdd.n1935 vdd.n1929 171.744
R16929 vdd.n2004 vdd.n2003 171.744
R16930 vdd.n2003 vdd.n2002 171.744
R16931 vdd.n2002 vdd.n1971 171.744
R16932 vdd.n1995 vdd.n1971 171.744
R16933 vdd.n1995 vdd.n1994 171.744
R16934 vdd.n1994 vdd.n1976 171.744
R16935 vdd.n1987 vdd.n1976 171.744
R16936 vdd.n1987 vdd.n1986 171.744
R16937 vdd.n1986 vdd.n1980 171.744
R16938 vdd.n1859 vdd.n1858 171.744
R16939 vdd.n1858 vdd.n1857 171.744
R16940 vdd.n1857 vdd.n1826 171.744
R16941 vdd.n1850 vdd.n1826 171.744
R16942 vdd.n1850 vdd.n1849 171.744
R16943 vdd.n1849 vdd.n1831 171.744
R16944 vdd.n1842 vdd.n1831 171.744
R16945 vdd.n1842 vdd.n1841 171.744
R16946 vdd.n1841 vdd.n1835 171.744
R16947 vdd.n1910 vdd.n1909 171.744
R16948 vdd.n1909 vdd.n1908 171.744
R16949 vdd.n1908 vdd.n1877 171.744
R16950 vdd.n1901 vdd.n1877 171.744
R16951 vdd.n1901 vdd.n1900 171.744
R16952 vdd.n1900 vdd.n1882 171.744
R16953 vdd.n1893 vdd.n1882 171.744
R16954 vdd.n1893 vdd.n1892 171.744
R16955 vdd.n1892 vdd.n1886 171.744
R16956 vdd.n1766 vdd.n1765 171.744
R16957 vdd.n1765 vdd.n1764 171.744
R16958 vdd.n1764 vdd.n1733 171.744
R16959 vdd.n1757 vdd.n1733 171.744
R16960 vdd.n1757 vdd.n1756 171.744
R16961 vdd.n1756 vdd.n1738 171.744
R16962 vdd.n1749 vdd.n1738 171.744
R16963 vdd.n1749 vdd.n1748 171.744
R16964 vdd.n1748 vdd.n1742 171.744
R16965 vdd.n1817 vdd.n1816 171.744
R16966 vdd.n1816 vdd.n1815 171.744
R16967 vdd.n1815 vdd.n1784 171.744
R16968 vdd.n1808 vdd.n1784 171.744
R16969 vdd.n1808 vdd.n1807 171.744
R16970 vdd.n1807 vdd.n1789 171.744
R16971 vdd.n1800 vdd.n1789 171.744
R16972 vdd.n1800 vdd.n1799 171.744
R16973 vdd.n1799 vdd.n1793 171.744
R16974 vdd.n3402 vdd.n356 146.341
R16975 vdd.n3400 vdd.n3399 146.341
R16976 vdd.n3397 vdd.n360 146.341
R16977 vdd.n3393 vdd.n3392 146.341
R16978 vdd.n3390 vdd.n368 146.341
R16979 vdd.n3386 vdd.n3385 146.341
R16980 vdd.n3383 vdd.n375 146.341
R16981 vdd.n3379 vdd.n3378 146.341
R16982 vdd.n3376 vdd.n382 146.341
R16983 vdd.n393 vdd.n390 146.341
R16984 vdd.n3368 vdd.n3367 146.341
R16985 vdd.n3365 vdd.n395 146.341
R16986 vdd.n3361 vdd.n3360 146.341
R16987 vdd.n3358 vdd.n401 146.341
R16988 vdd.n3354 vdd.n3353 146.341
R16989 vdd.n3351 vdd.n408 146.341
R16990 vdd.n3347 vdd.n3346 146.341
R16991 vdd.n3344 vdd.n415 146.341
R16992 vdd.n3340 vdd.n3339 146.341
R16993 vdd.n3337 vdd.n422 146.341
R16994 vdd.n433 vdd.n430 146.341
R16995 vdd.n3329 vdd.n3328 146.341
R16996 vdd.n3326 vdd.n435 146.341
R16997 vdd.n3322 vdd.n3321 146.341
R16998 vdd.n3319 vdd.n441 146.341
R16999 vdd.n3315 vdd.n3314 146.341
R17000 vdd.n3312 vdd.n448 146.341
R17001 vdd.n3308 vdd.n3307 146.341
R17002 vdd.n3305 vdd.n455 146.341
R17003 vdd.n3301 vdd.n3300 146.341
R17004 vdd.n3298 vdd.n462 146.341
R17005 vdd.n3213 vdd.n512 146.341
R17006 vdd.n3219 vdd.n512 146.341
R17007 vdd.n3219 vdd.n504 146.341
R17008 vdd.n3229 vdd.n504 146.341
R17009 vdd.n3229 vdd.n500 146.341
R17010 vdd.n3235 vdd.n500 146.341
R17011 vdd.n3235 vdd.n491 146.341
R17012 vdd.n3245 vdd.n491 146.341
R17013 vdd.n3245 vdd.n487 146.341
R17014 vdd.n3251 vdd.n487 146.341
R17015 vdd.n3251 vdd.n479 146.341
R17016 vdd.n3262 vdd.n479 146.341
R17017 vdd.n3262 vdd.n480 146.341
R17018 vdd.n480 vdd.n316 146.341
R17019 vdd.n317 vdd.n316 146.341
R17020 vdd.n318 vdd.n317 146.341
R17021 vdd.n473 vdd.n318 146.341
R17022 vdd.n473 vdd.n326 146.341
R17023 vdd.n327 vdd.n326 146.341
R17024 vdd.n328 vdd.n327 146.341
R17025 vdd.n470 vdd.n328 146.341
R17026 vdd.n470 vdd.n337 146.341
R17027 vdd.n338 vdd.n337 146.341
R17028 vdd.n339 vdd.n338 146.341
R17029 vdd.n467 vdd.n339 146.341
R17030 vdd.n467 vdd.n348 146.341
R17031 vdd.n349 vdd.n348 146.341
R17032 vdd.n350 vdd.n349 146.341
R17033 vdd.n3205 vdd.n3203 146.341
R17034 vdd.n3203 vdd.n3202 146.341
R17035 vdd.n3199 vdd.n3198 146.341
R17036 vdd.n3195 vdd.n3194 146.341
R17037 vdd.n3192 vdd.n526 146.341
R17038 vdd.n3188 vdd.n3186 146.341
R17039 vdd.n3184 vdd.n532 146.341
R17040 vdd.n3180 vdd.n3178 146.341
R17041 vdd.n3176 vdd.n538 146.341
R17042 vdd.n3172 vdd.n3170 146.341
R17043 vdd.n3168 vdd.n546 146.341
R17044 vdd.n3164 vdd.n3162 146.341
R17045 vdd.n3160 vdd.n552 146.341
R17046 vdd.n3156 vdd.n3154 146.341
R17047 vdd.n3152 vdd.n558 146.341
R17048 vdd.n3148 vdd.n3146 146.341
R17049 vdd.n3144 vdd.n564 146.341
R17050 vdd.n3140 vdd.n3138 146.341
R17051 vdd.n3136 vdd.n570 146.341
R17052 vdd.n3132 vdd.n3130 146.341
R17053 vdd.n3128 vdd.n576 146.341
R17054 vdd.n3121 vdd.n585 146.341
R17055 vdd.n3119 vdd.n3118 146.341
R17056 vdd.n3115 vdd.n3114 146.341
R17057 vdd.n3112 vdd.n590 146.341
R17058 vdd.n3108 vdd.n3106 146.341
R17059 vdd.n3104 vdd.n596 146.341
R17060 vdd.n3100 vdd.n3098 146.341
R17061 vdd.n3096 vdd.n602 146.341
R17062 vdd.n3092 vdd.n3090 146.341
R17063 vdd.n3087 vdd.n3086 146.341
R17064 vdd.n3083 vdd.n515 146.341
R17065 vdd.n3211 vdd.n510 146.341
R17066 vdd.n3221 vdd.n510 146.341
R17067 vdd.n3221 vdd.n506 146.341
R17068 vdd.n3227 vdd.n506 146.341
R17069 vdd.n3227 vdd.n498 146.341
R17070 vdd.n3237 vdd.n498 146.341
R17071 vdd.n3237 vdd.n494 146.341
R17072 vdd.n3243 vdd.n494 146.341
R17073 vdd.n3243 vdd.n486 146.341
R17074 vdd.n3254 vdd.n486 146.341
R17075 vdd.n3254 vdd.n482 146.341
R17076 vdd.n3260 vdd.n482 146.341
R17077 vdd.n3260 vdd.n314 146.341
R17078 vdd.n3437 vdd.n314 146.341
R17079 vdd.n3437 vdd.n315 146.341
R17080 vdd.n3433 vdd.n315 146.341
R17081 vdd.n3433 vdd.n319 146.341
R17082 vdd.n3429 vdd.n319 146.341
R17083 vdd.n3429 vdd.n324 146.341
R17084 vdd.n3425 vdd.n324 146.341
R17085 vdd.n3425 vdd.n330 146.341
R17086 vdd.n3421 vdd.n330 146.341
R17087 vdd.n3421 vdd.n336 146.341
R17088 vdd.n3417 vdd.n336 146.341
R17089 vdd.n3417 vdd.n341 146.341
R17090 vdd.n3413 vdd.n341 146.341
R17091 vdd.n3413 vdd.n347 146.341
R17092 vdd.n3409 vdd.n347 146.341
R17093 vdd.n2183 vdd.n2182 146.341
R17094 vdd.n2180 vdd.n2177 146.341
R17095 vdd.n2175 vdd.n1013 146.341
R17096 vdd.n2171 vdd.n2170 146.341
R17097 vdd.n2168 vdd.n1017 146.341
R17098 vdd.n2164 vdd.n2163 146.341
R17099 vdd.n2161 vdd.n1024 146.341
R17100 vdd.n2157 vdd.n2156 146.341
R17101 vdd.n2154 vdd.n1031 146.341
R17102 vdd.n1042 vdd.n1039 146.341
R17103 vdd.n2146 vdd.n2145 146.341
R17104 vdd.n2143 vdd.n1044 146.341
R17105 vdd.n2139 vdd.n2138 146.341
R17106 vdd.n2136 vdd.n1050 146.341
R17107 vdd.n2132 vdd.n2131 146.341
R17108 vdd.n2129 vdd.n1057 146.341
R17109 vdd.n2125 vdd.n2124 146.341
R17110 vdd.n2122 vdd.n1064 146.341
R17111 vdd.n2118 vdd.n2117 146.341
R17112 vdd.n2115 vdd.n1071 146.341
R17113 vdd.n1082 vdd.n1079 146.341
R17114 vdd.n2107 vdd.n2106 146.341
R17115 vdd.n2104 vdd.n1084 146.341
R17116 vdd.n2100 vdd.n2099 146.341
R17117 vdd.n2097 vdd.n1090 146.341
R17118 vdd.n2093 vdd.n2092 146.341
R17119 vdd.n2090 vdd.n1097 146.341
R17120 vdd.n2086 vdd.n2085 146.341
R17121 vdd.n2083 vdd.n1104 146.341
R17122 vdd.n1350 vdd.n1348 146.341
R17123 vdd.n1353 vdd.n1352 146.341
R17124 vdd.n1671 vdd.n1433 146.341
R17125 vdd.n1677 vdd.n1433 146.341
R17126 vdd.n1677 vdd.n1426 146.341
R17127 vdd.n1687 vdd.n1426 146.341
R17128 vdd.n1687 vdd.n1422 146.341
R17129 vdd.n1693 vdd.n1422 146.341
R17130 vdd.n1693 vdd.n1413 146.341
R17131 vdd.n1703 vdd.n1413 146.341
R17132 vdd.n1703 vdd.n1409 146.341
R17133 vdd.n1709 vdd.n1409 146.341
R17134 vdd.n1709 vdd.n1402 146.341
R17135 vdd.n1720 vdd.n1402 146.341
R17136 vdd.n1720 vdd.n1398 146.341
R17137 vdd.n1726 vdd.n1398 146.341
R17138 vdd.n1726 vdd.n1391 146.341
R17139 vdd.n2018 vdd.n1391 146.341
R17140 vdd.n2018 vdd.n1387 146.341
R17141 vdd.n2024 vdd.n1387 146.341
R17142 vdd.n2024 vdd.n1379 146.341
R17143 vdd.n2035 vdd.n1379 146.341
R17144 vdd.n2035 vdd.n1375 146.341
R17145 vdd.n2041 vdd.n1375 146.341
R17146 vdd.n2041 vdd.n1369 146.341
R17147 vdd.n2052 vdd.n1369 146.341
R17148 vdd.n2052 vdd.n1364 146.341
R17149 vdd.n2060 vdd.n1364 146.341
R17150 vdd.n2060 vdd.n1355 146.341
R17151 vdd.n2071 vdd.n1355 146.341
R17152 vdd.n1443 vdd.n1442 146.341
R17153 vdd.n1446 vdd.n1443 146.341
R17154 vdd.n1449 vdd.n1448 146.341
R17155 vdd.n1454 vdd.n1451 146.341
R17156 vdd.n1457 vdd.n1456 146.341
R17157 vdd.n1462 vdd.n1459 146.341
R17158 vdd.n1465 vdd.n1464 146.341
R17159 vdd.n1470 vdd.n1467 146.341
R17160 vdd.n1473 vdd.n1472 146.341
R17161 vdd.n1480 vdd.n1475 146.341
R17162 vdd.n1483 vdd.n1482 146.341
R17163 vdd.n1488 vdd.n1485 146.341
R17164 vdd.n1491 vdd.n1490 146.341
R17165 vdd.n1496 vdd.n1493 146.341
R17166 vdd.n1499 vdd.n1498 146.341
R17167 vdd.n1504 vdd.n1501 146.341
R17168 vdd.n1507 vdd.n1506 146.341
R17169 vdd.n1512 vdd.n1509 146.341
R17170 vdd.n1515 vdd.n1514 146.341
R17171 vdd.n1520 vdd.n1517 146.341
R17172 vdd.n1601 vdd.n1522 146.341
R17173 vdd.n1599 vdd.n1598 146.341
R17174 vdd.n1529 vdd.n1528 146.341
R17175 vdd.n1532 vdd.n1531 146.341
R17176 vdd.n1537 vdd.n1536 146.341
R17177 vdd.n1540 vdd.n1539 146.341
R17178 vdd.n1545 vdd.n1544 146.341
R17179 vdd.n1548 vdd.n1547 146.341
R17180 vdd.n1553 vdd.n1552 146.341
R17181 vdd.n1556 vdd.n1555 146.341
R17182 vdd.n1561 vdd.n1560 146.341
R17183 vdd.n1563 vdd.n1436 146.341
R17184 vdd.n1669 vdd.n1432 146.341
R17185 vdd.n1679 vdd.n1432 146.341
R17186 vdd.n1679 vdd.n1428 146.341
R17187 vdd.n1685 vdd.n1428 146.341
R17188 vdd.n1685 vdd.n1420 146.341
R17189 vdd.n1695 vdd.n1420 146.341
R17190 vdd.n1695 vdd.n1416 146.341
R17191 vdd.n1701 vdd.n1416 146.341
R17192 vdd.n1701 vdd.n1408 146.341
R17193 vdd.n1712 vdd.n1408 146.341
R17194 vdd.n1712 vdd.n1404 146.341
R17195 vdd.n1718 vdd.n1404 146.341
R17196 vdd.n1718 vdd.n1397 146.341
R17197 vdd.n1728 vdd.n1397 146.341
R17198 vdd.n1728 vdd.n1393 146.341
R17199 vdd.n2016 vdd.n1393 146.341
R17200 vdd.n2016 vdd.n1385 146.341
R17201 vdd.n2027 vdd.n1385 146.341
R17202 vdd.n2027 vdd.n1381 146.341
R17203 vdd.n2033 vdd.n1381 146.341
R17204 vdd.n2033 vdd.n1374 146.341
R17205 vdd.n2044 vdd.n1374 146.341
R17206 vdd.n2044 vdd.n1370 146.341
R17207 vdd.n2050 vdd.n1370 146.341
R17208 vdd.n2050 vdd.n1362 146.341
R17209 vdd.n2063 vdd.n1362 146.341
R17210 vdd.n2063 vdd.n1357 146.341
R17211 vdd.n2069 vdd.n1357 146.341
R17212 vdd.n1143 vdd.t167 127.284
R17213 vdd.n838 vdd.t211 127.284
R17214 vdd.n1147 vdd.t208 127.284
R17215 vdd.n829 vdd.t234 127.284
R17216 vdd.n724 vdd.t188 127.284
R17217 vdd.n724 vdd.t189 127.284
R17218 vdd.n2535 vdd.t229 127.284
R17219 vdd.n661 vdd.t176 127.284
R17220 vdd.n2532 vdd.t219 127.284
R17221 vdd.n625 vdd.t162 127.284
R17222 vdd.n899 vdd.t225 127.284
R17223 vdd.n899 vdd.t226 127.284
R17224 vdd.n22 vdd.n20 117.314
R17225 vdd.n17 vdd.n15 117.314
R17226 vdd.n27 vdd.n26 116.927
R17227 vdd.n24 vdd.n23 116.927
R17228 vdd.n22 vdd.n21 116.927
R17229 vdd.n17 vdd.n16 116.927
R17230 vdd.n19 vdd.n18 116.927
R17231 vdd.n27 vdd.n25 116.927
R17232 vdd.n1144 vdd.t166 111.188
R17233 vdd.n839 vdd.t212 111.188
R17234 vdd.n1148 vdd.t207 111.188
R17235 vdd.n830 vdd.t235 111.188
R17236 vdd.n2536 vdd.t228 111.188
R17237 vdd.n662 vdd.t177 111.188
R17238 vdd.n2533 vdd.t218 111.188
R17239 vdd.n626 vdd.t163 111.188
R17240 vdd.n2806 vdd.n788 99.5127
R17241 vdd.n2806 vdd.n779 99.5127
R17242 vdd.n2814 vdd.n779 99.5127
R17243 vdd.n2814 vdd.n777 99.5127
R17244 vdd.n2818 vdd.n777 99.5127
R17245 vdd.n2818 vdd.n767 99.5127
R17246 vdd.n2826 vdd.n767 99.5127
R17247 vdd.n2826 vdd.n765 99.5127
R17248 vdd.n2830 vdd.n765 99.5127
R17249 vdd.n2830 vdd.n756 99.5127
R17250 vdd.n2838 vdd.n756 99.5127
R17251 vdd.n2838 vdd.n754 99.5127
R17252 vdd.n2842 vdd.n754 99.5127
R17253 vdd.n2842 vdd.n745 99.5127
R17254 vdd.n2850 vdd.n745 99.5127
R17255 vdd.n2850 vdd.n743 99.5127
R17256 vdd.n2854 vdd.n743 99.5127
R17257 vdd.n2854 vdd.n732 99.5127
R17258 vdd.n2863 vdd.n732 99.5127
R17259 vdd.n2863 vdd.n730 99.5127
R17260 vdd.n2867 vdd.n730 99.5127
R17261 vdd.n2867 vdd.n720 99.5127
R17262 vdd.n2875 vdd.n720 99.5127
R17263 vdd.n2875 vdd.n718 99.5127
R17264 vdd.n2879 vdd.n718 99.5127
R17265 vdd.n2879 vdd.n708 99.5127
R17266 vdd.n2887 vdd.n708 99.5127
R17267 vdd.n2887 vdd.n706 99.5127
R17268 vdd.n2891 vdd.n706 99.5127
R17269 vdd.n2891 vdd.n695 99.5127
R17270 vdd.n2899 vdd.n695 99.5127
R17271 vdd.n2899 vdd.n693 99.5127
R17272 vdd.n2903 vdd.n693 99.5127
R17273 vdd.n2903 vdd.n684 99.5127
R17274 vdd.n2911 vdd.n684 99.5127
R17275 vdd.n2911 vdd.n682 99.5127
R17276 vdd.n2915 vdd.n682 99.5127
R17277 vdd.n2915 vdd.n670 99.5127
R17278 vdd.n2968 vdd.n670 99.5127
R17279 vdd.n2968 vdd.n668 99.5127
R17280 vdd.n2972 vdd.n668 99.5127
R17281 vdd.n2972 vdd.n634 99.5127
R17282 vdd.n3042 vdd.n634 99.5127
R17283 vdd.n3038 vdd.n635 99.5127
R17284 vdd.n3036 vdd.n3035 99.5127
R17285 vdd.n3033 vdd.n639 99.5127
R17286 vdd.n3029 vdd.n3028 99.5127
R17287 vdd.n3026 vdd.n642 99.5127
R17288 vdd.n3022 vdd.n3021 99.5127
R17289 vdd.n3019 vdd.n645 99.5127
R17290 vdd.n3015 vdd.n3014 99.5127
R17291 vdd.n3012 vdd.n648 99.5127
R17292 vdd.n3007 vdd.n3006 99.5127
R17293 vdd.n3004 vdd.n651 99.5127
R17294 vdd.n3000 vdd.n2999 99.5127
R17295 vdd.n2997 vdd.n654 99.5127
R17296 vdd.n2993 vdd.n2992 99.5127
R17297 vdd.n2990 vdd.n657 99.5127
R17298 vdd.n2986 vdd.n2985 99.5127
R17299 vdd.n2983 vdd.n660 99.5127
R17300 vdd.n2733 vdd.n786 99.5127
R17301 vdd.n2729 vdd.n786 99.5127
R17302 vdd.n2729 vdd.n780 99.5127
R17303 vdd.n2611 vdd.n780 99.5127
R17304 vdd.n2611 vdd.n775 99.5127
R17305 vdd.n2614 vdd.n775 99.5127
R17306 vdd.n2614 vdd.n769 99.5127
R17307 vdd.n2715 vdd.n769 99.5127
R17308 vdd.n2715 vdd.n763 99.5127
R17309 vdd.n2711 vdd.n763 99.5127
R17310 vdd.n2711 vdd.n757 99.5127
R17311 vdd.n2658 vdd.n757 99.5127
R17312 vdd.n2658 vdd.n751 99.5127
R17313 vdd.n2655 vdd.n751 99.5127
R17314 vdd.n2655 vdd.n746 99.5127
R17315 vdd.n2652 vdd.n746 99.5127
R17316 vdd.n2652 vdd.n741 99.5127
R17317 vdd.n2649 vdd.n741 99.5127
R17318 vdd.n2649 vdd.n734 99.5127
R17319 vdd.n2646 vdd.n734 99.5127
R17320 vdd.n2646 vdd.n727 99.5127
R17321 vdd.n2643 vdd.n727 99.5127
R17322 vdd.n2643 vdd.n721 99.5127
R17323 vdd.n2640 vdd.n721 99.5127
R17324 vdd.n2640 vdd.n716 99.5127
R17325 vdd.n2637 vdd.n716 99.5127
R17326 vdd.n2637 vdd.n710 99.5127
R17327 vdd.n2634 vdd.n710 99.5127
R17328 vdd.n2634 vdd.n703 99.5127
R17329 vdd.n2631 vdd.n703 99.5127
R17330 vdd.n2631 vdd.n696 99.5127
R17331 vdd.n2628 vdd.n696 99.5127
R17332 vdd.n2628 vdd.n690 99.5127
R17333 vdd.n2625 vdd.n690 99.5127
R17334 vdd.n2625 vdd.n685 99.5127
R17335 vdd.n2622 vdd.n685 99.5127
R17336 vdd.n2622 vdd.n680 99.5127
R17337 vdd.n2619 vdd.n680 99.5127
R17338 vdd.n2619 vdd.n672 99.5127
R17339 vdd.n672 vdd.n665 99.5127
R17340 vdd.n2974 vdd.n665 99.5127
R17341 vdd.n2975 vdd.n2974 99.5127
R17342 vdd.n2975 vdd.n632 99.5127
R17343 vdd.n2799 vdd.n790 99.5127
R17344 vdd.n2799 vdd.n2531 99.5127
R17345 vdd.n2795 vdd.n2794 99.5127
R17346 vdd.n2791 vdd.n2790 99.5127
R17347 vdd.n2787 vdd.n2786 99.5127
R17348 vdd.n2783 vdd.n2782 99.5127
R17349 vdd.n2779 vdd.n2778 99.5127
R17350 vdd.n2775 vdd.n2774 99.5127
R17351 vdd.n2771 vdd.n2770 99.5127
R17352 vdd.n2767 vdd.n2766 99.5127
R17353 vdd.n2763 vdd.n2762 99.5127
R17354 vdd.n2759 vdd.n2758 99.5127
R17355 vdd.n2755 vdd.n2754 99.5127
R17356 vdd.n2751 vdd.n2750 99.5127
R17357 vdd.n2747 vdd.n2746 99.5127
R17358 vdd.n2743 vdd.n2742 99.5127
R17359 vdd.n2738 vdd.n2737 99.5127
R17360 vdd.n2495 vdd.n827 99.5127
R17361 vdd.n2491 vdd.n2490 99.5127
R17362 vdd.n2487 vdd.n2486 99.5127
R17363 vdd.n2483 vdd.n2482 99.5127
R17364 vdd.n2479 vdd.n2478 99.5127
R17365 vdd.n2475 vdd.n2474 99.5127
R17366 vdd.n2471 vdd.n2470 99.5127
R17367 vdd.n2467 vdd.n2466 99.5127
R17368 vdd.n2463 vdd.n2462 99.5127
R17369 vdd.n2459 vdd.n2458 99.5127
R17370 vdd.n2455 vdd.n2454 99.5127
R17371 vdd.n2451 vdd.n2450 99.5127
R17372 vdd.n2447 vdd.n2446 99.5127
R17373 vdd.n2443 vdd.n2442 99.5127
R17374 vdd.n2439 vdd.n2438 99.5127
R17375 vdd.n2435 vdd.n2434 99.5127
R17376 vdd.n2430 vdd.n2429 99.5127
R17377 vdd.n1183 vdd.n963 99.5127
R17378 vdd.n1186 vdd.n963 99.5127
R17379 vdd.n1186 vdd.n957 99.5127
R17380 vdd.n1189 vdd.n957 99.5127
R17381 vdd.n1189 vdd.n952 99.5127
R17382 vdd.n1192 vdd.n952 99.5127
R17383 vdd.n1192 vdd.n945 99.5127
R17384 vdd.n1195 vdd.n945 99.5127
R17385 vdd.n1195 vdd.n938 99.5127
R17386 vdd.n1198 vdd.n938 99.5127
R17387 vdd.n1198 vdd.n932 99.5127
R17388 vdd.n1201 vdd.n932 99.5127
R17389 vdd.n1201 vdd.n927 99.5127
R17390 vdd.n1204 vdd.n927 99.5127
R17391 vdd.n1204 vdd.n922 99.5127
R17392 vdd.n1207 vdd.n922 99.5127
R17393 vdd.n1207 vdd.n916 99.5127
R17394 vdd.n1210 vdd.n916 99.5127
R17395 vdd.n1210 vdd.n909 99.5127
R17396 vdd.n1213 vdd.n909 99.5127
R17397 vdd.n1213 vdd.n902 99.5127
R17398 vdd.n1216 vdd.n902 99.5127
R17399 vdd.n1216 vdd.n896 99.5127
R17400 vdd.n1219 vdd.n896 99.5127
R17401 vdd.n1219 vdd.n891 99.5127
R17402 vdd.n1222 vdd.n891 99.5127
R17403 vdd.n1222 vdd.n885 99.5127
R17404 vdd.n1264 vdd.n885 99.5127
R17405 vdd.n1264 vdd.n878 99.5127
R17406 vdd.n1260 vdd.n878 99.5127
R17407 vdd.n1260 vdd.n872 99.5127
R17408 vdd.n1257 vdd.n872 99.5127
R17409 vdd.n1257 vdd.n867 99.5127
R17410 vdd.n1254 vdd.n867 99.5127
R17411 vdd.n1254 vdd.n862 99.5127
R17412 vdd.n1234 vdd.n862 99.5127
R17413 vdd.n1234 vdd.n857 99.5127
R17414 vdd.n1231 vdd.n857 99.5127
R17415 vdd.n1231 vdd.n850 99.5127
R17416 vdd.n1228 vdd.n850 99.5127
R17417 vdd.n1228 vdd.n843 99.5127
R17418 vdd.n843 vdd.n832 99.5127
R17419 vdd.n2425 vdd.n832 99.5127
R17420 vdd.n2217 vdd.n968 99.5127
R17421 vdd.n2217 vdd.n1004 99.5127
R17422 vdd.n2213 vdd.n2212 99.5127
R17423 vdd.n2209 vdd.n2208 99.5127
R17424 vdd.n2205 vdd.n2204 99.5127
R17425 vdd.n2201 vdd.n2200 99.5127
R17426 vdd.n2197 vdd.n2196 99.5127
R17427 vdd.n2193 vdd.n2192 99.5127
R17428 vdd.n2189 vdd.n2188 99.5127
R17429 vdd.n1150 vdd.n1149 99.5127
R17430 vdd.n1154 vdd.n1153 99.5127
R17431 vdd.n1158 vdd.n1157 99.5127
R17432 vdd.n1162 vdd.n1161 99.5127
R17433 vdd.n1166 vdd.n1165 99.5127
R17434 vdd.n1170 vdd.n1169 99.5127
R17435 vdd.n1174 vdd.n1173 99.5127
R17436 vdd.n1179 vdd.n1178 99.5127
R17437 vdd.n2224 vdd.n966 99.5127
R17438 vdd.n2224 vdd.n956 99.5127
R17439 vdd.n2232 vdd.n956 99.5127
R17440 vdd.n2232 vdd.n954 99.5127
R17441 vdd.n2236 vdd.n954 99.5127
R17442 vdd.n2236 vdd.n943 99.5127
R17443 vdd.n2244 vdd.n943 99.5127
R17444 vdd.n2244 vdd.n941 99.5127
R17445 vdd.n2248 vdd.n941 99.5127
R17446 vdd.n2248 vdd.n931 99.5127
R17447 vdd.n2256 vdd.n931 99.5127
R17448 vdd.n2256 vdd.n929 99.5127
R17449 vdd.n2260 vdd.n929 99.5127
R17450 vdd.n2260 vdd.n920 99.5127
R17451 vdd.n2268 vdd.n920 99.5127
R17452 vdd.n2268 vdd.n918 99.5127
R17453 vdd.n2272 vdd.n918 99.5127
R17454 vdd.n2272 vdd.n907 99.5127
R17455 vdd.n2280 vdd.n907 99.5127
R17456 vdd.n2280 vdd.n905 99.5127
R17457 vdd.n2284 vdd.n905 99.5127
R17458 vdd.n2284 vdd.n895 99.5127
R17459 vdd.n2293 vdd.n895 99.5127
R17460 vdd.n2293 vdd.n893 99.5127
R17461 vdd.n2297 vdd.n893 99.5127
R17462 vdd.n2297 vdd.n883 99.5127
R17463 vdd.n2305 vdd.n883 99.5127
R17464 vdd.n2305 vdd.n881 99.5127
R17465 vdd.n2309 vdd.n881 99.5127
R17466 vdd.n2309 vdd.n871 99.5127
R17467 vdd.n2317 vdd.n871 99.5127
R17468 vdd.n2317 vdd.n869 99.5127
R17469 vdd.n2321 vdd.n869 99.5127
R17470 vdd.n2321 vdd.n861 99.5127
R17471 vdd.n2329 vdd.n861 99.5127
R17472 vdd.n2329 vdd.n859 99.5127
R17473 vdd.n2333 vdd.n859 99.5127
R17474 vdd.n2333 vdd.n848 99.5127
R17475 vdd.n2343 vdd.n848 99.5127
R17476 vdd.n2343 vdd.n845 99.5127
R17477 vdd.n2348 vdd.n845 99.5127
R17478 vdd.n2348 vdd.n846 99.5127
R17479 vdd.n846 vdd.n826 99.5127
R17480 vdd.n2958 vdd.n2957 99.5127
R17481 vdd.n2955 vdd.n2921 99.5127
R17482 vdd.n2951 vdd.n2950 99.5127
R17483 vdd.n2948 vdd.n2924 99.5127
R17484 vdd.n2944 vdd.n2943 99.5127
R17485 vdd.n2941 vdd.n2927 99.5127
R17486 vdd.n2937 vdd.n2936 99.5127
R17487 vdd.n2934 vdd.n2931 99.5127
R17488 vdd.n3075 vdd.n612 99.5127
R17489 vdd.n3073 vdd.n3072 99.5127
R17490 vdd.n3070 vdd.n615 99.5127
R17491 vdd.n3066 vdd.n3065 99.5127
R17492 vdd.n3063 vdd.n618 99.5127
R17493 vdd.n3059 vdd.n3058 99.5127
R17494 vdd.n3056 vdd.n621 99.5127
R17495 vdd.n3052 vdd.n3051 99.5127
R17496 vdd.n3049 vdd.n624 99.5127
R17497 vdd.n2607 vdd.n787 99.5127
R17498 vdd.n2727 vdd.n787 99.5127
R17499 vdd.n2727 vdd.n781 99.5127
R17500 vdd.n2723 vdd.n781 99.5127
R17501 vdd.n2723 vdd.n776 99.5127
R17502 vdd.n2720 vdd.n776 99.5127
R17503 vdd.n2720 vdd.n770 99.5127
R17504 vdd.n2717 vdd.n770 99.5127
R17505 vdd.n2717 vdd.n764 99.5127
R17506 vdd.n2709 vdd.n764 99.5127
R17507 vdd.n2709 vdd.n758 99.5127
R17508 vdd.n2705 vdd.n758 99.5127
R17509 vdd.n2705 vdd.n752 99.5127
R17510 vdd.n2702 vdd.n752 99.5127
R17511 vdd.n2702 vdd.n747 99.5127
R17512 vdd.n2699 vdd.n747 99.5127
R17513 vdd.n2699 vdd.n742 99.5127
R17514 vdd.n2696 vdd.n742 99.5127
R17515 vdd.n2696 vdd.n735 99.5127
R17516 vdd.n2693 vdd.n735 99.5127
R17517 vdd.n2693 vdd.n728 99.5127
R17518 vdd.n2690 vdd.n728 99.5127
R17519 vdd.n2690 vdd.n722 99.5127
R17520 vdd.n2687 vdd.n722 99.5127
R17521 vdd.n2687 vdd.n717 99.5127
R17522 vdd.n2684 vdd.n717 99.5127
R17523 vdd.n2684 vdd.n711 99.5127
R17524 vdd.n2681 vdd.n711 99.5127
R17525 vdd.n2681 vdd.n704 99.5127
R17526 vdd.n2678 vdd.n704 99.5127
R17527 vdd.n2678 vdd.n697 99.5127
R17528 vdd.n2675 vdd.n697 99.5127
R17529 vdd.n2675 vdd.n691 99.5127
R17530 vdd.n2672 vdd.n691 99.5127
R17531 vdd.n2672 vdd.n686 99.5127
R17532 vdd.n2669 vdd.n686 99.5127
R17533 vdd.n2669 vdd.n681 99.5127
R17534 vdd.n2666 vdd.n681 99.5127
R17535 vdd.n2666 vdd.n673 99.5127
R17536 vdd.n2663 vdd.n673 99.5127
R17537 vdd.n2663 vdd.n666 99.5127
R17538 vdd.n666 vdd.n630 99.5127
R17539 vdd.n3044 vdd.n630 99.5127
R17540 vdd.n2542 vdd.n2541 99.5127
R17541 vdd.n2546 vdd.n2545 99.5127
R17542 vdd.n2550 vdd.n2549 99.5127
R17543 vdd.n2554 vdd.n2553 99.5127
R17544 vdd.n2558 vdd.n2557 99.5127
R17545 vdd.n2562 vdd.n2561 99.5127
R17546 vdd.n2566 vdd.n2565 99.5127
R17547 vdd.n2570 vdd.n2569 99.5127
R17548 vdd.n2574 vdd.n2573 99.5127
R17549 vdd.n2578 vdd.n2577 99.5127
R17550 vdd.n2582 vdd.n2581 99.5127
R17551 vdd.n2586 vdd.n2585 99.5127
R17552 vdd.n2590 vdd.n2589 99.5127
R17553 vdd.n2594 vdd.n2593 99.5127
R17554 vdd.n2598 vdd.n2597 99.5127
R17555 vdd.n2602 vdd.n2601 99.5127
R17556 vdd.n2604 vdd.n2530 99.5127
R17557 vdd.n2808 vdd.n784 99.5127
R17558 vdd.n2808 vdd.n782 99.5127
R17559 vdd.n2812 vdd.n782 99.5127
R17560 vdd.n2812 vdd.n773 99.5127
R17561 vdd.n2820 vdd.n773 99.5127
R17562 vdd.n2820 vdd.n771 99.5127
R17563 vdd.n2824 vdd.n771 99.5127
R17564 vdd.n2824 vdd.n762 99.5127
R17565 vdd.n2832 vdd.n762 99.5127
R17566 vdd.n2832 vdd.n760 99.5127
R17567 vdd.n2836 vdd.n760 99.5127
R17568 vdd.n2836 vdd.n750 99.5127
R17569 vdd.n2844 vdd.n750 99.5127
R17570 vdd.n2844 vdd.n748 99.5127
R17571 vdd.n2848 vdd.n748 99.5127
R17572 vdd.n2848 vdd.n739 99.5127
R17573 vdd.n2856 vdd.n739 99.5127
R17574 vdd.n2856 vdd.n737 99.5127
R17575 vdd.n2861 vdd.n737 99.5127
R17576 vdd.n2861 vdd.n726 99.5127
R17577 vdd.n2869 vdd.n726 99.5127
R17578 vdd.n2869 vdd.n723 99.5127
R17579 vdd.n2873 vdd.n723 99.5127
R17580 vdd.n2873 vdd.n714 99.5127
R17581 vdd.n2881 vdd.n714 99.5127
R17582 vdd.n2881 vdd.n712 99.5127
R17583 vdd.n2885 vdd.n712 99.5127
R17584 vdd.n2885 vdd.n701 99.5127
R17585 vdd.n2893 vdd.n701 99.5127
R17586 vdd.n2893 vdd.n699 99.5127
R17587 vdd.n2897 vdd.n699 99.5127
R17588 vdd.n2897 vdd.n689 99.5127
R17589 vdd.n2905 vdd.n689 99.5127
R17590 vdd.n2905 vdd.n687 99.5127
R17591 vdd.n2909 vdd.n687 99.5127
R17592 vdd.n2909 vdd.n678 99.5127
R17593 vdd.n2917 vdd.n678 99.5127
R17594 vdd.n2917 vdd.n675 99.5127
R17595 vdd.n2966 vdd.n675 99.5127
R17596 vdd.n2966 vdd.n676 99.5127
R17597 vdd.n676 vdd.n667 99.5127
R17598 vdd.n2961 vdd.n667 99.5127
R17599 vdd.n2961 vdd.n633 99.5127
R17600 vdd.n2419 vdd.n2418 99.5127
R17601 vdd.n2415 vdd.n2414 99.5127
R17602 vdd.n2411 vdd.n2410 99.5127
R17603 vdd.n2407 vdd.n2406 99.5127
R17604 vdd.n2403 vdd.n2402 99.5127
R17605 vdd.n2399 vdd.n2398 99.5127
R17606 vdd.n2395 vdd.n2394 99.5127
R17607 vdd.n2391 vdd.n2390 99.5127
R17608 vdd.n2387 vdd.n2386 99.5127
R17609 vdd.n2383 vdd.n2382 99.5127
R17610 vdd.n2379 vdd.n2378 99.5127
R17611 vdd.n2375 vdd.n2374 99.5127
R17612 vdd.n2371 vdd.n2370 99.5127
R17613 vdd.n2367 vdd.n2366 99.5127
R17614 vdd.n2363 vdd.n2362 99.5127
R17615 vdd.n2359 vdd.n2358 99.5127
R17616 vdd.n2355 vdd.n808 99.5127
R17617 vdd.n1308 vdd.n964 99.5127
R17618 vdd.n1305 vdd.n964 99.5127
R17619 vdd.n1305 vdd.n958 99.5127
R17620 vdd.n1302 vdd.n958 99.5127
R17621 vdd.n1302 vdd.n953 99.5127
R17622 vdd.n1299 vdd.n953 99.5127
R17623 vdd.n1299 vdd.n946 99.5127
R17624 vdd.n1296 vdd.n946 99.5127
R17625 vdd.n1296 vdd.n939 99.5127
R17626 vdd.n1293 vdd.n939 99.5127
R17627 vdd.n1293 vdd.n933 99.5127
R17628 vdd.n1290 vdd.n933 99.5127
R17629 vdd.n1290 vdd.n928 99.5127
R17630 vdd.n1287 vdd.n928 99.5127
R17631 vdd.n1287 vdd.n923 99.5127
R17632 vdd.n1284 vdd.n923 99.5127
R17633 vdd.n1284 vdd.n917 99.5127
R17634 vdd.n1281 vdd.n917 99.5127
R17635 vdd.n1281 vdd.n910 99.5127
R17636 vdd.n1278 vdd.n910 99.5127
R17637 vdd.n1278 vdd.n903 99.5127
R17638 vdd.n1275 vdd.n903 99.5127
R17639 vdd.n1275 vdd.n897 99.5127
R17640 vdd.n1272 vdd.n897 99.5127
R17641 vdd.n1272 vdd.n892 99.5127
R17642 vdd.n1269 vdd.n892 99.5127
R17643 vdd.n1269 vdd.n886 99.5127
R17644 vdd.n1266 vdd.n886 99.5127
R17645 vdd.n1266 vdd.n879 99.5127
R17646 vdd.n1237 vdd.n879 99.5127
R17647 vdd.n1237 vdd.n873 99.5127
R17648 vdd.n1240 vdd.n873 99.5127
R17649 vdd.n1240 vdd.n868 99.5127
R17650 vdd.n1252 vdd.n868 99.5127
R17651 vdd.n1252 vdd.n863 99.5127
R17652 vdd.n1248 vdd.n863 99.5127
R17653 vdd.n1248 vdd.n858 99.5127
R17654 vdd.n1245 vdd.n858 99.5127
R17655 vdd.n1245 vdd.n851 99.5127
R17656 vdd.n851 vdd.n842 99.5127
R17657 vdd.n2350 vdd.n842 99.5127
R17658 vdd.n2351 vdd.n2350 99.5127
R17659 vdd.n2351 vdd.n834 99.5127
R17660 vdd.n1112 vdd.n1111 99.5127
R17661 vdd.n1116 vdd.n1115 99.5127
R17662 vdd.n1120 vdd.n1119 99.5127
R17663 vdd.n1124 vdd.n1123 99.5127
R17664 vdd.n1128 vdd.n1127 99.5127
R17665 vdd.n1132 vdd.n1131 99.5127
R17666 vdd.n1136 vdd.n1135 99.5127
R17667 vdd.n1140 vdd.n1139 99.5127
R17668 vdd.n1341 vdd.n1142 99.5127
R17669 vdd.n1339 vdd.n1338 99.5127
R17670 vdd.n1335 vdd.n1334 99.5127
R17671 vdd.n1331 vdd.n1330 99.5127
R17672 vdd.n1327 vdd.n1326 99.5127
R17673 vdd.n1323 vdd.n1322 99.5127
R17674 vdd.n1319 vdd.n1318 99.5127
R17675 vdd.n1315 vdd.n1314 99.5127
R17676 vdd.n1311 vdd.n1003 99.5127
R17677 vdd.n2226 vdd.n961 99.5127
R17678 vdd.n2226 vdd.n959 99.5127
R17679 vdd.n2230 vdd.n959 99.5127
R17680 vdd.n2230 vdd.n950 99.5127
R17681 vdd.n2238 vdd.n950 99.5127
R17682 vdd.n2238 vdd.n948 99.5127
R17683 vdd.n2242 vdd.n948 99.5127
R17684 vdd.n2242 vdd.n937 99.5127
R17685 vdd.n2250 vdd.n937 99.5127
R17686 vdd.n2250 vdd.n935 99.5127
R17687 vdd.n2254 vdd.n935 99.5127
R17688 vdd.n2254 vdd.n926 99.5127
R17689 vdd.n2262 vdd.n926 99.5127
R17690 vdd.n2262 vdd.n924 99.5127
R17691 vdd.n2266 vdd.n924 99.5127
R17692 vdd.n2266 vdd.n914 99.5127
R17693 vdd.n2274 vdd.n914 99.5127
R17694 vdd.n2274 vdd.n912 99.5127
R17695 vdd.n2278 vdd.n912 99.5127
R17696 vdd.n2278 vdd.n901 99.5127
R17697 vdd.n2286 vdd.n901 99.5127
R17698 vdd.n2286 vdd.n898 99.5127
R17699 vdd.n2291 vdd.n898 99.5127
R17700 vdd.n2291 vdd.n889 99.5127
R17701 vdd.n2299 vdd.n889 99.5127
R17702 vdd.n2299 vdd.n887 99.5127
R17703 vdd.n2303 vdd.n887 99.5127
R17704 vdd.n2303 vdd.n877 99.5127
R17705 vdd.n2311 vdd.n877 99.5127
R17706 vdd.n2311 vdd.n875 99.5127
R17707 vdd.n2315 vdd.n875 99.5127
R17708 vdd.n2315 vdd.n866 99.5127
R17709 vdd.n2323 vdd.n866 99.5127
R17710 vdd.n2323 vdd.n864 99.5127
R17711 vdd.n2327 vdd.n864 99.5127
R17712 vdd.n2327 vdd.n855 99.5127
R17713 vdd.n2335 vdd.n855 99.5127
R17714 vdd.n2335 vdd.n852 99.5127
R17715 vdd.n2341 vdd.n852 99.5127
R17716 vdd.n2341 vdd.n853 99.5127
R17717 vdd.n853 vdd.n844 99.5127
R17718 vdd.n844 vdd.n835 99.5127
R17719 vdd.n2423 vdd.n835 99.5127
R17720 vdd.n9 vdd.n7 98.9633
R17721 vdd.n2 vdd.n0 98.9633
R17722 vdd.n9 vdd.n8 98.6055
R17723 vdd.n11 vdd.n10 98.6055
R17724 vdd.n13 vdd.n12 98.6055
R17725 vdd.n6 vdd.n5 98.6055
R17726 vdd.n4 vdd.n3 98.6055
R17727 vdd.n2 vdd.n1 98.6055
R17728 vdd.t73 vdd.n279 85.8723
R17729 vdd.t152 vdd.n228 85.8723
R17730 vdd.t154 vdd.n185 85.8723
R17731 vdd.t146 vdd.n134 85.8723
R17732 vdd.t97 vdd.n92 85.8723
R17733 vdd.t113 vdd.n41 85.8723
R17734 vdd.t101 vdd.n1929 85.8723
R17735 vdd.t107 vdd.n1980 85.8723
R17736 vdd.t90 vdd.n1835 85.8723
R17737 vdd.t95 vdd.n1886 85.8723
R17738 vdd.t114 vdd.n1742 85.8723
R17739 vdd.t96 vdd.n1793 85.8723
R17740 vdd.n725 vdd.n724 78.546
R17741 vdd.n2289 vdd.n899 78.546
R17742 vdd.n266 vdd.n265 75.1835
R17743 vdd.n264 vdd.n263 75.1835
R17744 vdd.n262 vdd.n261 75.1835
R17745 vdd.n260 vdd.n259 75.1835
R17746 vdd.n258 vdd.n257 75.1835
R17747 vdd.n172 vdd.n171 75.1835
R17748 vdd.n170 vdd.n169 75.1835
R17749 vdd.n168 vdd.n167 75.1835
R17750 vdd.n166 vdd.n165 75.1835
R17751 vdd.n164 vdd.n163 75.1835
R17752 vdd.n79 vdd.n78 75.1835
R17753 vdd.n77 vdd.n76 75.1835
R17754 vdd.n75 vdd.n74 75.1835
R17755 vdd.n73 vdd.n72 75.1835
R17756 vdd.n71 vdd.n70 75.1835
R17757 vdd.n1959 vdd.n1958 75.1835
R17758 vdd.n1961 vdd.n1960 75.1835
R17759 vdd.n1963 vdd.n1962 75.1835
R17760 vdd.n1965 vdd.n1964 75.1835
R17761 vdd.n1967 vdd.n1966 75.1835
R17762 vdd.n1865 vdd.n1864 75.1835
R17763 vdd.n1867 vdd.n1866 75.1835
R17764 vdd.n1869 vdd.n1868 75.1835
R17765 vdd.n1871 vdd.n1870 75.1835
R17766 vdd.n1873 vdd.n1872 75.1835
R17767 vdd.n1772 vdd.n1771 75.1835
R17768 vdd.n1774 vdd.n1773 75.1835
R17769 vdd.n1776 vdd.n1775 75.1835
R17770 vdd.n1778 vdd.n1777 75.1835
R17771 vdd.n1780 vdd.n1779 75.1835
R17772 vdd.n2800 vdd.n2513 72.8958
R17773 vdd.n2800 vdd.n2514 72.8958
R17774 vdd.n2800 vdd.n2515 72.8958
R17775 vdd.n2800 vdd.n2516 72.8958
R17776 vdd.n2800 vdd.n2517 72.8958
R17777 vdd.n2800 vdd.n2518 72.8958
R17778 vdd.n2800 vdd.n2519 72.8958
R17779 vdd.n2800 vdd.n2520 72.8958
R17780 vdd.n2800 vdd.n2521 72.8958
R17781 vdd.n2800 vdd.n2522 72.8958
R17782 vdd.n2800 vdd.n2523 72.8958
R17783 vdd.n2800 vdd.n2524 72.8958
R17784 vdd.n2800 vdd.n2525 72.8958
R17785 vdd.n2800 vdd.n2526 72.8958
R17786 vdd.n2800 vdd.n2527 72.8958
R17787 vdd.n2800 vdd.n2528 72.8958
R17788 vdd.n2800 vdd.n2529 72.8958
R17789 vdd.n629 vdd.n613 72.8958
R17790 vdd.n3050 vdd.n613 72.8958
R17791 vdd.n623 vdd.n613 72.8958
R17792 vdd.n3057 vdd.n613 72.8958
R17793 vdd.n620 vdd.n613 72.8958
R17794 vdd.n3064 vdd.n613 72.8958
R17795 vdd.n617 vdd.n613 72.8958
R17796 vdd.n3071 vdd.n613 72.8958
R17797 vdd.n3074 vdd.n613 72.8958
R17798 vdd.n2930 vdd.n613 72.8958
R17799 vdd.n2935 vdd.n613 72.8958
R17800 vdd.n2929 vdd.n613 72.8958
R17801 vdd.n2942 vdd.n613 72.8958
R17802 vdd.n2926 vdd.n613 72.8958
R17803 vdd.n2949 vdd.n613 72.8958
R17804 vdd.n2923 vdd.n613 72.8958
R17805 vdd.n2956 vdd.n613 72.8958
R17806 vdd.n2219 vdd.n2218 72.8958
R17807 vdd.n2218 vdd.n970 72.8958
R17808 vdd.n2218 vdd.n971 72.8958
R17809 vdd.n2218 vdd.n972 72.8958
R17810 vdd.n2218 vdd.n973 72.8958
R17811 vdd.n2218 vdd.n974 72.8958
R17812 vdd.n2218 vdd.n975 72.8958
R17813 vdd.n2218 vdd.n976 72.8958
R17814 vdd.n2218 vdd.n977 72.8958
R17815 vdd.n2218 vdd.n978 72.8958
R17816 vdd.n2218 vdd.n979 72.8958
R17817 vdd.n2218 vdd.n980 72.8958
R17818 vdd.n2218 vdd.n981 72.8958
R17819 vdd.n2218 vdd.n982 72.8958
R17820 vdd.n2218 vdd.n983 72.8958
R17821 vdd.n2218 vdd.n984 72.8958
R17822 vdd.n2218 vdd.n985 72.8958
R17823 vdd.n2496 vdd.n809 72.8958
R17824 vdd.n2496 vdd.n810 72.8958
R17825 vdd.n2496 vdd.n811 72.8958
R17826 vdd.n2496 vdd.n812 72.8958
R17827 vdd.n2496 vdd.n813 72.8958
R17828 vdd.n2496 vdd.n814 72.8958
R17829 vdd.n2496 vdd.n815 72.8958
R17830 vdd.n2496 vdd.n816 72.8958
R17831 vdd.n2496 vdd.n817 72.8958
R17832 vdd.n2496 vdd.n818 72.8958
R17833 vdd.n2496 vdd.n819 72.8958
R17834 vdd.n2496 vdd.n820 72.8958
R17835 vdd.n2496 vdd.n821 72.8958
R17836 vdd.n2496 vdd.n822 72.8958
R17837 vdd.n2496 vdd.n823 72.8958
R17838 vdd.n2496 vdd.n824 72.8958
R17839 vdd.n2496 vdd.n825 72.8958
R17840 vdd.n2801 vdd.n2800 72.8958
R17841 vdd.n2800 vdd.n2497 72.8958
R17842 vdd.n2800 vdd.n2498 72.8958
R17843 vdd.n2800 vdd.n2499 72.8958
R17844 vdd.n2800 vdd.n2500 72.8958
R17845 vdd.n2800 vdd.n2501 72.8958
R17846 vdd.n2800 vdd.n2502 72.8958
R17847 vdd.n2800 vdd.n2503 72.8958
R17848 vdd.n2800 vdd.n2504 72.8958
R17849 vdd.n2800 vdd.n2505 72.8958
R17850 vdd.n2800 vdd.n2506 72.8958
R17851 vdd.n2800 vdd.n2507 72.8958
R17852 vdd.n2800 vdd.n2508 72.8958
R17853 vdd.n2800 vdd.n2509 72.8958
R17854 vdd.n2800 vdd.n2510 72.8958
R17855 vdd.n2800 vdd.n2511 72.8958
R17856 vdd.n2800 vdd.n2512 72.8958
R17857 vdd.n2978 vdd.n613 72.8958
R17858 vdd.n2984 vdd.n613 72.8958
R17859 vdd.n659 vdd.n613 72.8958
R17860 vdd.n2991 vdd.n613 72.8958
R17861 vdd.n656 vdd.n613 72.8958
R17862 vdd.n2998 vdd.n613 72.8958
R17863 vdd.n653 vdd.n613 72.8958
R17864 vdd.n3005 vdd.n613 72.8958
R17865 vdd.n650 vdd.n613 72.8958
R17866 vdd.n3013 vdd.n613 72.8958
R17867 vdd.n647 vdd.n613 72.8958
R17868 vdd.n3020 vdd.n613 72.8958
R17869 vdd.n644 vdd.n613 72.8958
R17870 vdd.n3027 vdd.n613 72.8958
R17871 vdd.n641 vdd.n613 72.8958
R17872 vdd.n3034 vdd.n613 72.8958
R17873 vdd.n3037 vdd.n613 72.8958
R17874 vdd.n2496 vdd.n807 72.8958
R17875 vdd.n2496 vdd.n806 72.8958
R17876 vdd.n2496 vdd.n805 72.8958
R17877 vdd.n2496 vdd.n804 72.8958
R17878 vdd.n2496 vdd.n803 72.8958
R17879 vdd.n2496 vdd.n802 72.8958
R17880 vdd.n2496 vdd.n801 72.8958
R17881 vdd.n2496 vdd.n800 72.8958
R17882 vdd.n2496 vdd.n799 72.8958
R17883 vdd.n2496 vdd.n798 72.8958
R17884 vdd.n2496 vdd.n797 72.8958
R17885 vdd.n2496 vdd.n796 72.8958
R17886 vdd.n2496 vdd.n795 72.8958
R17887 vdd.n2496 vdd.n794 72.8958
R17888 vdd.n2496 vdd.n793 72.8958
R17889 vdd.n2496 vdd.n792 72.8958
R17890 vdd.n2496 vdd.n791 72.8958
R17891 vdd.n2218 vdd.n986 72.8958
R17892 vdd.n2218 vdd.n987 72.8958
R17893 vdd.n2218 vdd.n988 72.8958
R17894 vdd.n2218 vdd.n989 72.8958
R17895 vdd.n2218 vdd.n990 72.8958
R17896 vdd.n2218 vdd.n991 72.8958
R17897 vdd.n2218 vdd.n992 72.8958
R17898 vdd.n2218 vdd.n993 72.8958
R17899 vdd.n2218 vdd.n994 72.8958
R17900 vdd.n2218 vdd.n995 72.8958
R17901 vdd.n2218 vdd.n996 72.8958
R17902 vdd.n2218 vdd.n997 72.8958
R17903 vdd.n2218 vdd.n998 72.8958
R17904 vdd.n2218 vdd.n999 72.8958
R17905 vdd.n2218 vdd.n1000 72.8958
R17906 vdd.n2218 vdd.n1001 72.8958
R17907 vdd.n2218 vdd.n1002 72.8958
R17908 vdd.n1441 vdd.n1437 66.2847
R17909 vdd.n1447 vdd.n1437 66.2847
R17910 vdd.n1450 vdd.n1437 66.2847
R17911 vdd.n1455 vdd.n1437 66.2847
R17912 vdd.n1458 vdd.n1437 66.2847
R17913 vdd.n1463 vdd.n1437 66.2847
R17914 vdd.n1466 vdd.n1437 66.2847
R17915 vdd.n1471 vdd.n1437 66.2847
R17916 vdd.n1474 vdd.n1437 66.2847
R17917 vdd.n1481 vdd.n1437 66.2847
R17918 vdd.n1484 vdd.n1437 66.2847
R17919 vdd.n1489 vdd.n1437 66.2847
R17920 vdd.n1492 vdd.n1437 66.2847
R17921 vdd.n1497 vdd.n1437 66.2847
R17922 vdd.n1500 vdd.n1437 66.2847
R17923 vdd.n1505 vdd.n1437 66.2847
R17924 vdd.n1508 vdd.n1437 66.2847
R17925 vdd.n1513 vdd.n1437 66.2847
R17926 vdd.n1516 vdd.n1437 66.2847
R17927 vdd.n1521 vdd.n1437 66.2847
R17928 vdd.n1600 vdd.n1437 66.2847
R17929 vdd.n1524 vdd.n1437 66.2847
R17930 vdd.n1530 vdd.n1437 66.2847
R17931 vdd.n1535 vdd.n1437 66.2847
R17932 vdd.n1538 vdd.n1437 66.2847
R17933 vdd.n1543 vdd.n1437 66.2847
R17934 vdd.n1546 vdd.n1437 66.2847
R17935 vdd.n1551 vdd.n1437 66.2847
R17936 vdd.n1554 vdd.n1437 66.2847
R17937 vdd.n1559 vdd.n1437 66.2847
R17938 vdd.n1562 vdd.n1437 66.2847
R17939 vdd.n1354 vdd.n969 66.2847
R17940 vdd.n1351 vdd.n969 66.2847
R17941 vdd.n1347 vdd.n969 66.2847
R17942 vdd.n2084 vdd.n969 66.2847
R17943 vdd.n1103 vdd.n969 66.2847
R17944 vdd.n2091 vdd.n969 66.2847
R17945 vdd.n1096 vdd.n969 66.2847
R17946 vdd.n2098 vdd.n969 66.2847
R17947 vdd.n1089 vdd.n969 66.2847
R17948 vdd.n2105 vdd.n969 66.2847
R17949 vdd.n1083 vdd.n969 66.2847
R17950 vdd.n1078 vdd.n969 66.2847
R17951 vdd.n2116 vdd.n969 66.2847
R17952 vdd.n1070 vdd.n969 66.2847
R17953 vdd.n2123 vdd.n969 66.2847
R17954 vdd.n1063 vdd.n969 66.2847
R17955 vdd.n2130 vdd.n969 66.2847
R17956 vdd.n1056 vdd.n969 66.2847
R17957 vdd.n2137 vdd.n969 66.2847
R17958 vdd.n1049 vdd.n969 66.2847
R17959 vdd.n2144 vdd.n969 66.2847
R17960 vdd.n1043 vdd.n969 66.2847
R17961 vdd.n1038 vdd.n969 66.2847
R17962 vdd.n2155 vdd.n969 66.2847
R17963 vdd.n1030 vdd.n969 66.2847
R17964 vdd.n2162 vdd.n969 66.2847
R17965 vdd.n1023 vdd.n969 66.2847
R17966 vdd.n2169 vdd.n969 66.2847
R17967 vdd.n1016 vdd.n969 66.2847
R17968 vdd.n2176 vdd.n969 66.2847
R17969 vdd.n2181 vdd.n969 66.2847
R17970 vdd.n1012 vdd.n969 66.2847
R17971 vdd.n3204 vdd.n516 66.2847
R17972 vdd.n520 vdd.n516 66.2847
R17973 vdd.n523 vdd.n516 66.2847
R17974 vdd.n3193 vdd.n516 66.2847
R17975 vdd.n3187 vdd.n516 66.2847
R17976 vdd.n3185 vdd.n516 66.2847
R17977 vdd.n3179 vdd.n516 66.2847
R17978 vdd.n3177 vdd.n516 66.2847
R17979 vdd.n3171 vdd.n516 66.2847
R17980 vdd.n3169 vdd.n516 66.2847
R17981 vdd.n3163 vdd.n516 66.2847
R17982 vdd.n3161 vdd.n516 66.2847
R17983 vdd.n3155 vdd.n516 66.2847
R17984 vdd.n3153 vdd.n516 66.2847
R17985 vdd.n3147 vdd.n516 66.2847
R17986 vdd.n3145 vdd.n516 66.2847
R17987 vdd.n3139 vdd.n516 66.2847
R17988 vdd.n3137 vdd.n516 66.2847
R17989 vdd.n3131 vdd.n516 66.2847
R17990 vdd.n3129 vdd.n516 66.2847
R17991 vdd.n584 vdd.n516 66.2847
R17992 vdd.n3120 vdd.n516 66.2847
R17993 vdd.n586 vdd.n516 66.2847
R17994 vdd.n3113 vdd.n516 66.2847
R17995 vdd.n3107 vdd.n516 66.2847
R17996 vdd.n3105 vdd.n516 66.2847
R17997 vdd.n3099 vdd.n516 66.2847
R17998 vdd.n3097 vdd.n516 66.2847
R17999 vdd.n3091 vdd.n516 66.2847
R18000 vdd.n607 vdd.n516 66.2847
R18001 vdd.n609 vdd.n516 66.2847
R18002 vdd.n3290 vdd.n351 66.2847
R18003 vdd.n3299 vdd.n351 66.2847
R18004 vdd.n461 vdd.n351 66.2847
R18005 vdd.n3306 vdd.n351 66.2847
R18006 vdd.n454 vdd.n351 66.2847
R18007 vdd.n3313 vdd.n351 66.2847
R18008 vdd.n447 vdd.n351 66.2847
R18009 vdd.n3320 vdd.n351 66.2847
R18010 vdd.n440 vdd.n351 66.2847
R18011 vdd.n3327 vdd.n351 66.2847
R18012 vdd.n434 vdd.n351 66.2847
R18013 vdd.n429 vdd.n351 66.2847
R18014 vdd.n3338 vdd.n351 66.2847
R18015 vdd.n421 vdd.n351 66.2847
R18016 vdd.n3345 vdd.n351 66.2847
R18017 vdd.n414 vdd.n351 66.2847
R18018 vdd.n3352 vdd.n351 66.2847
R18019 vdd.n407 vdd.n351 66.2847
R18020 vdd.n3359 vdd.n351 66.2847
R18021 vdd.n400 vdd.n351 66.2847
R18022 vdd.n3366 vdd.n351 66.2847
R18023 vdd.n394 vdd.n351 66.2847
R18024 vdd.n389 vdd.n351 66.2847
R18025 vdd.n3377 vdd.n351 66.2847
R18026 vdd.n381 vdd.n351 66.2847
R18027 vdd.n3384 vdd.n351 66.2847
R18028 vdd.n374 vdd.n351 66.2847
R18029 vdd.n3391 vdd.n351 66.2847
R18030 vdd.n367 vdd.n351 66.2847
R18031 vdd.n3398 vdd.n351 66.2847
R18032 vdd.n3401 vdd.n351 66.2847
R18033 vdd.n355 vdd.n351 66.2847
R18034 vdd.n356 vdd.n355 52.4337
R18035 vdd.n3401 vdd.n3400 52.4337
R18036 vdd.n3398 vdd.n3397 52.4337
R18037 vdd.n3393 vdd.n367 52.4337
R18038 vdd.n3391 vdd.n3390 52.4337
R18039 vdd.n3386 vdd.n374 52.4337
R18040 vdd.n3384 vdd.n3383 52.4337
R18041 vdd.n3379 vdd.n381 52.4337
R18042 vdd.n3377 vdd.n3376 52.4337
R18043 vdd.n390 vdd.n389 52.4337
R18044 vdd.n3368 vdd.n394 52.4337
R18045 vdd.n3366 vdd.n3365 52.4337
R18046 vdd.n3361 vdd.n400 52.4337
R18047 vdd.n3359 vdd.n3358 52.4337
R18048 vdd.n3354 vdd.n407 52.4337
R18049 vdd.n3352 vdd.n3351 52.4337
R18050 vdd.n3347 vdd.n414 52.4337
R18051 vdd.n3345 vdd.n3344 52.4337
R18052 vdd.n3340 vdd.n421 52.4337
R18053 vdd.n3338 vdd.n3337 52.4337
R18054 vdd.n430 vdd.n429 52.4337
R18055 vdd.n3329 vdd.n434 52.4337
R18056 vdd.n3327 vdd.n3326 52.4337
R18057 vdd.n3322 vdd.n440 52.4337
R18058 vdd.n3320 vdd.n3319 52.4337
R18059 vdd.n3315 vdd.n447 52.4337
R18060 vdd.n3313 vdd.n3312 52.4337
R18061 vdd.n3308 vdd.n454 52.4337
R18062 vdd.n3306 vdd.n3305 52.4337
R18063 vdd.n3301 vdd.n461 52.4337
R18064 vdd.n3299 vdd.n3298 52.4337
R18065 vdd.n3291 vdd.n3290 52.4337
R18066 vdd.n3204 vdd.n517 52.4337
R18067 vdd.n3202 vdd.n520 52.4337
R18068 vdd.n3198 vdd.n523 52.4337
R18069 vdd.n3194 vdd.n3193 52.4337
R18070 vdd.n3187 vdd.n526 52.4337
R18071 vdd.n3186 vdd.n3185 52.4337
R18072 vdd.n3179 vdd.n532 52.4337
R18073 vdd.n3178 vdd.n3177 52.4337
R18074 vdd.n3171 vdd.n538 52.4337
R18075 vdd.n3170 vdd.n3169 52.4337
R18076 vdd.n3163 vdd.n546 52.4337
R18077 vdd.n3162 vdd.n3161 52.4337
R18078 vdd.n3155 vdd.n552 52.4337
R18079 vdd.n3154 vdd.n3153 52.4337
R18080 vdd.n3147 vdd.n558 52.4337
R18081 vdd.n3146 vdd.n3145 52.4337
R18082 vdd.n3139 vdd.n564 52.4337
R18083 vdd.n3138 vdd.n3137 52.4337
R18084 vdd.n3131 vdd.n570 52.4337
R18085 vdd.n3130 vdd.n3129 52.4337
R18086 vdd.n584 vdd.n576 52.4337
R18087 vdd.n3121 vdd.n3120 52.4337
R18088 vdd.n3118 vdd.n586 52.4337
R18089 vdd.n3114 vdd.n3113 52.4337
R18090 vdd.n3107 vdd.n590 52.4337
R18091 vdd.n3106 vdd.n3105 52.4337
R18092 vdd.n3099 vdd.n596 52.4337
R18093 vdd.n3098 vdd.n3097 52.4337
R18094 vdd.n3091 vdd.n602 52.4337
R18095 vdd.n3090 vdd.n607 52.4337
R18096 vdd.n3086 vdd.n609 52.4337
R18097 vdd.n2183 vdd.n1012 52.4337
R18098 vdd.n2181 vdd.n2180 52.4337
R18099 vdd.n2176 vdd.n2175 52.4337
R18100 vdd.n2171 vdd.n1016 52.4337
R18101 vdd.n2169 vdd.n2168 52.4337
R18102 vdd.n2164 vdd.n1023 52.4337
R18103 vdd.n2162 vdd.n2161 52.4337
R18104 vdd.n2157 vdd.n1030 52.4337
R18105 vdd.n2155 vdd.n2154 52.4337
R18106 vdd.n1039 vdd.n1038 52.4337
R18107 vdd.n2146 vdd.n1043 52.4337
R18108 vdd.n2144 vdd.n2143 52.4337
R18109 vdd.n2139 vdd.n1049 52.4337
R18110 vdd.n2137 vdd.n2136 52.4337
R18111 vdd.n2132 vdd.n1056 52.4337
R18112 vdd.n2130 vdd.n2129 52.4337
R18113 vdd.n2125 vdd.n1063 52.4337
R18114 vdd.n2123 vdd.n2122 52.4337
R18115 vdd.n2118 vdd.n1070 52.4337
R18116 vdd.n2116 vdd.n2115 52.4337
R18117 vdd.n1079 vdd.n1078 52.4337
R18118 vdd.n2107 vdd.n1083 52.4337
R18119 vdd.n2105 vdd.n2104 52.4337
R18120 vdd.n2100 vdd.n1089 52.4337
R18121 vdd.n2098 vdd.n2097 52.4337
R18122 vdd.n2093 vdd.n1096 52.4337
R18123 vdd.n2091 vdd.n2090 52.4337
R18124 vdd.n2086 vdd.n1103 52.4337
R18125 vdd.n2084 vdd.n2083 52.4337
R18126 vdd.n1348 vdd.n1347 52.4337
R18127 vdd.n1352 vdd.n1351 52.4337
R18128 vdd.n2072 vdd.n1354 52.4337
R18129 vdd.n1441 vdd.n1439 52.4337
R18130 vdd.n1447 vdd.n1446 52.4337
R18131 vdd.n1450 vdd.n1449 52.4337
R18132 vdd.n1455 vdd.n1454 52.4337
R18133 vdd.n1458 vdd.n1457 52.4337
R18134 vdd.n1463 vdd.n1462 52.4337
R18135 vdd.n1466 vdd.n1465 52.4337
R18136 vdd.n1471 vdd.n1470 52.4337
R18137 vdd.n1474 vdd.n1473 52.4337
R18138 vdd.n1481 vdd.n1480 52.4337
R18139 vdd.n1484 vdd.n1483 52.4337
R18140 vdd.n1489 vdd.n1488 52.4337
R18141 vdd.n1492 vdd.n1491 52.4337
R18142 vdd.n1497 vdd.n1496 52.4337
R18143 vdd.n1500 vdd.n1499 52.4337
R18144 vdd.n1505 vdd.n1504 52.4337
R18145 vdd.n1508 vdd.n1507 52.4337
R18146 vdd.n1513 vdd.n1512 52.4337
R18147 vdd.n1516 vdd.n1515 52.4337
R18148 vdd.n1521 vdd.n1520 52.4337
R18149 vdd.n1601 vdd.n1600 52.4337
R18150 vdd.n1598 vdd.n1524 52.4337
R18151 vdd.n1530 vdd.n1529 52.4337
R18152 vdd.n1535 vdd.n1532 52.4337
R18153 vdd.n1538 vdd.n1537 52.4337
R18154 vdd.n1543 vdd.n1540 52.4337
R18155 vdd.n1546 vdd.n1545 52.4337
R18156 vdd.n1551 vdd.n1548 52.4337
R18157 vdd.n1554 vdd.n1553 52.4337
R18158 vdd.n1559 vdd.n1556 52.4337
R18159 vdd.n1562 vdd.n1561 52.4337
R18160 vdd.n1442 vdd.n1441 52.4337
R18161 vdd.n1448 vdd.n1447 52.4337
R18162 vdd.n1451 vdd.n1450 52.4337
R18163 vdd.n1456 vdd.n1455 52.4337
R18164 vdd.n1459 vdd.n1458 52.4337
R18165 vdd.n1464 vdd.n1463 52.4337
R18166 vdd.n1467 vdd.n1466 52.4337
R18167 vdd.n1472 vdd.n1471 52.4337
R18168 vdd.n1475 vdd.n1474 52.4337
R18169 vdd.n1482 vdd.n1481 52.4337
R18170 vdd.n1485 vdd.n1484 52.4337
R18171 vdd.n1490 vdd.n1489 52.4337
R18172 vdd.n1493 vdd.n1492 52.4337
R18173 vdd.n1498 vdd.n1497 52.4337
R18174 vdd.n1501 vdd.n1500 52.4337
R18175 vdd.n1506 vdd.n1505 52.4337
R18176 vdd.n1509 vdd.n1508 52.4337
R18177 vdd.n1514 vdd.n1513 52.4337
R18178 vdd.n1517 vdd.n1516 52.4337
R18179 vdd.n1522 vdd.n1521 52.4337
R18180 vdd.n1600 vdd.n1599 52.4337
R18181 vdd.n1528 vdd.n1524 52.4337
R18182 vdd.n1531 vdd.n1530 52.4337
R18183 vdd.n1536 vdd.n1535 52.4337
R18184 vdd.n1539 vdd.n1538 52.4337
R18185 vdd.n1544 vdd.n1543 52.4337
R18186 vdd.n1547 vdd.n1546 52.4337
R18187 vdd.n1552 vdd.n1551 52.4337
R18188 vdd.n1555 vdd.n1554 52.4337
R18189 vdd.n1560 vdd.n1559 52.4337
R18190 vdd.n1563 vdd.n1562 52.4337
R18191 vdd.n1354 vdd.n1353 52.4337
R18192 vdd.n1351 vdd.n1350 52.4337
R18193 vdd.n1347 vdd.n1104 52.4337
R18194 vdd.n2085 vdd.n2084 52.4337
R18195 vdd.n1103 vdd.n1097 52.4337
R18196 vdd.n2092 vdd.n2091 52.4337
R18197 vdd.n1096 vdd.n1090 52.4337
R18198 vdd.n2099 vdd.n2098 52.4337
R18199 vdd.n1089 vdd.n1084 52.4337
R18200 vdd.n2106 vdd.n2105 52.4337
R18201 vdd.n1083 vdd.n1082 52.4337
R18202 vdd.n1078 vdd.n1071 52.4337
R18203 vdd.n2117 vdd.n2116 52.4337
R18204 vdd.n1070 vdd.n1064 52.4337
R18205 vdd.n2124 vdd.n2123 52.4337
R18206 vdd.n1063 vdd.n1057 52.4337
R18207 vdd.n2131 vdd.n2130 52.4337
R18208 vdd.n1056 vdd.n1050 52.4337
R18209 vdd.n2138 vdd.n2137 52.4337
R18210 vdd.n1049 vdd.n1044 52.4337
R18211 vdd.n2145 vdd.n2144 52.4337
R18212 vdd.n1043 vdd.n1042 52.4337
R18213 vdd.n1038 vdd.n1031 52.4337
R18214 vdd.n2156 vdd.n2155 52.4337
R18215 vdd.n1030 vdd.n1024 52.4337
R18216 vdd.n2163 vdd.n2162 52.4337
R18217 vdd.n1023 vdd.n1017 52.4337
R18218 vdd.n2170 vdd.n2169 52.4337
R18219 vdd.n1016 vdd.n1013 52.4337
R18220 vdd.n2177 vdd.n2176 52.4337
R18221 vdd.n2182 vdd.n2181 52.4337
R18222 vdd.n1358 vdd.n1012 52.4337
R18223 vdd.n3205 vdd.n3204 52.4337
R18224 vdd.n3199 vdd.n520 52.4337
R18225 vdd.n3195 vdd.n523 52.4337
R18226 vdd.n3193 vdd.n3192 52.4337
R18227 vdd.n3188 vdd.n3187 52.4337
R18228 vdd.n3185 vdd.n3184 52.4337
R18229 vdd.n3180 vdd.n3179 52.4337
R18230 vdd.n3177 vdd.n3176 52.4337
R18231 vdd.n3172 vdd.n3171 52.4337
R18232 vdd.n3169 vdd.n3168 52.4337
R18233 vdd.n3164 vdd.n3163 52.4337
R18234 vdd.n3161 vdd.n3160 52.4337
R18235 vdd.n3156 vdd.n3155 52.4337
R18236 vdd.n3153 vdd.n3152 52.4337
R18237 vdd.n3148 vdd.n3147 52.4337
R18238 vdd.n3145 vdd.n3144 52.4337
R18239 vdd.n3140 vdd.n3139 52.4337
R18240 vdd.n3137 vdd.n3136 52.4337
R18241 vdd.n3132 vdd.n3131 52.4337
R18242 vdd.n3129 vdd.n3128 52.4337
R18243 vdd.n585 vdd.n584 52.4337
R18244 vdd.n3120 vdd.n3119 52.4337
R18245 vdd.n3115 vdd.n586 52.4337
R18246 vdd.n3113 vdd.n3112 52.4337
R18247 vdd.n3108 vdd.n3107 52.4337
R18248 vdd.n3105 vdd.n3104 52.4337
R18249 vdd.n3100 vdd.n3099 52.4337
R18250 vdd.n3097 vdd.n3096 52.4337
R18251 vdd.n3092 vdd.n3091 52.4337
R18252 vdd.n3087 vdd.n607 52.4337
R18253 vdd.n3083 vdd.n609 52.4337
R18254 vdd.n3290 vdd.n462 52.4337
R18255 vdd.n3300 vdd.n3299 52.4337
R18256 vdd.n461 vdd.n455 52.4337
R18257 vdd.n3307 vdd.n3306 52.4337
R18258 vdd.n454 vdd.n448 52.4337
R18259 vdd.n3314 vdd.n3313 52.4337
R18260 vdd.n447 vdd.n441 52.4337
R18261 vdd.n3321 vdd.n3320 52.4337
R18262 vdd.n440 vdd.n435 52.4337
R18263 vdd.n3328 vdd.n3327 52.4337
R18264 vdd.n434 vdd.n433 52.4337
R18265 vdd.n429 vdd.n422 52.4337
R18266 vdd.n3339 vdd.n3338 52.4337
R18267 vdd.n421 vdd.n415 52.4337
R18268 vdd.n3346 vdd.n3345 52.4337
R18269 vdd.n414 vdd.n408 52.4337
R18270 vdd.n3353 vdd.n3352 52.4337
R18271 vdd.n407 vdd.n401 52.4337
R18272 vdd.n3360 vdd.n3359 52.4337
R18273 vdd.n400 vdd.n395 52.4337
R18274 vdd.n3367 vdd.n3366 52.4337
R18275 vdd.n394 vdd.n393 52.4337
R18276 vdd.n389 vdd.n382 52.4337
R18277 vdd.n3378 vdd.n3377 52.4337
R18278 vdd.n381 vdd.n375 52.4337
R18279 vdd.n3385 vdd.n3384 52.4337
R18280 vdd.n374 vdd.n368 52.4337
R18281 vdd.n3392 vdd.n3391 52.4337
R18282 vdd.n367 vdd.n360 52.4337
R18283 vdd.n3399 vdd.n3398 52.4337
R18284 vdd.n3402 vdd.n3401 52.4337
R18285 vdd.n355 vdd.n352 52.4337
R18286 vdd.t16 vdd.t29 51.4683
R18287 vdd.n258 vdd.n256 42.0461
R18288 vdd.n164 vdd.n162 42.0461
R18289 vdd.n71 vdd.n69 42.0461
R18290 vdd.n1959 vdd.n1957 42.0461
R18291 vdd.n1865 vdd.n1863 42.0461
R18292 vdd.n1772 vdd.n1770 42.0461
R18293 vdd.n308 vdd.n307 41.6884
R18294 vdd.n214 vdd.n213 41.6884
R18295 vdd.n121 vdd.n120 41.6884
R18296 vdd.n2009 vdd.n2008 41.6884
R18297 vdd.n1915 vdd.n1914 41.6884
R18298 vdd.n1822 vdd.n1821 41.6884
R18299 vdd.n1567 vdd.n1566 41.1157
R18300 vdd.n1604 vdd.n1603 41.1157
R18301 vdd.n1478 vdd.n1477 41.1157
R18302 vdd.n3295 vdd.n3294 41.1157
R18303 vdd.n3334 vdd.n428 41.1157
R18304 vdd.n3373 vdd.n388 41.1157
R18305 vdd.n3037 vdd.n3036 39.2114
R18306 vdd.n3034 vdd.n3033 39.2114
R18307 vdd.n3029 vdd.n641 39.2114
R18308 vdd.n3027 vdd.n3026 39.2114
R18309 vdd.n3022 vdd.n644 39.2114
R18310 vdd.n3020 vdd.n3019 39.2114
R18311 vdd.n3015 vdd.n647 39.2114
R18312 vdd.n3013 vdd.n3012 39.2114
R18313 vdd.n3007 vdd.n650 39.2114
R18314 vdd.n3005 vdd.n3004 39.2114
R18315 vdd.n3000 vdd.n653 39.2114
R18316 vdd.n2998 vdd.n2997 39.2114
R18317 vdd.n2993 vdd.n656 39.2114
R18318 vdd.n2991 vdd.n2990 39.2114
R18319 vdd.n2986 vdd.n659 39.2114
R18320 vdd.n2984 vdd.n2983 39.2114
R18321 vdd.n2979 vdd.n2978 39.2114
R18322 vdd.n2802 vdd.n2801 39.2114
R18323 vdd.n2531 vdd.n2497 39.2114
R18324 vdd.n2794 vdd.n2498 39.2114
R18325 vdd.n2790 vdd.n2499 39.2114
R18326 vdd.n2786 vdd.n2500 39.2114
R18327 vdd.n2782 vdd.n2501 39.2114
R18328 vdd.n2778 vdd.n2502 39.2114
R18329 vdd.n2774 vdd.n2503 39.2114
R18330 vdd.n2770 vdd.n2504 39.2114
R18331 vdd.n2766 vdd.n2505 39.2114
R18332 vdd.n2762 vdd.n2506 39.2114
R18333 vdd.n2758 vdd.n2507 39.2114
R18334 vdd.n2754 vdd.n2508 39.2114
R18335 vdd.n2750 vdd.n2509 39.2114
R18336 vdd.n2746 vdd.n2510 39.2114
R18337 vdd.n2742 vdd.n2511 39.2114
R18338 vdd.n2737 vdd.n2512 39.2114
R18339 vdd.n2491 vdd.n825 39.2114
R18340 vdd.n2487 vdd.n824 39.2114
R18341 vdd.n2483 vdd.n823 39.2114
R18342 vdd.n2479 vdd.n822 39.2114
R18343 vdd.n2475 vdd.n821 39.2114
R18344 vdd.n2471 vdd.n820 39.2114
R18345 vdd.n2467 vdd.n819 39.2114
R18346 vdd.n2463 vdd.n818 39.2114
R18347 vdd.n2459 vdd.n817 39.2114
R18348 vdd.n2455 vdd.n816 39.2114
R18349 vdd.n2451 vdd.n815 39.2114
R18350 vdd.n2447 vdd.n814 39.2114
R18351 vdd.n2443 vdd.n813 39.2114
R18352 vdd.n2439 vdd.n812 39.2114
R18353 vdd.n2435 vdd.n811 39.2114
R18354 vdd.n2430 vdd.n810 39.2114
R18355 vdd.n2426 vdd.n809 39.2114
R18356 vdd.n2220 vdd.n2219 39.2114
R18357 vdd.n1004 vdd.n970 39.2114
R18358 vdd.n2212 vdd.n971 39.2114
R18359 vdd.n2208 vdd.n972 39.2114
R18360 vdd.n2204 vdd.n973 39.2114
R18361 vdd.n2200 vdd.n974 39.2114
R18362 vdd.n2196 vdd.n975 39.2114
R18363 vdd.n2192 vdd.n976 39.2114
R18364 vdd.n2188 vdd.n977 39.2114
R18365 vdd.n1150 vdd.n978 39.2114
R18366 vdd.n1154 vdd.n979 39.2114
R18367 vdd.n1158 vdd.n980 39.2114
R18368 vdd.n1162 vdd.n981 39.2114
R18369 vdd.n1166 vdd.n982 39.2114
R18370 vdd.n1170 vdd.n983 39.2114
R18371 vdd.n1174 vdd.n984 39.2114
R18372 vdd.n1179 vdd.n985 39.2114
R18373 vdd.n2956 vdd.n2955 39.2114
R18374 vdd.n2951 vdd.n2923 39.2114
R18375 vdd.n2949 vdd.n2948 39.2114
R18376 vdd.n2944 vdd.n2926 39.2114
R18377 vdd.n2942 vdd.n2941 39.2114
R18378 vdd.n2937 vdd.n2929 39.2114
R18379 vdd.n2935 vdd.n2934 39.2114
R18380 vdd.n2930 vdd.n612 39.2114
R18381 vdd.n3074 vdd.n3073 39.2114
R18382 vdd.n3071 vdd.n3070 39.2114
R18383 vdd.n3066 vdd.n617 39.2114
R18384 vdd.n3064 vdd.n3063 39.2114
R18385 vdd.n3059 vdd.n620 39.2114
R18386 vdd.n3057 vdd.n3056 39.2114
R18387 vdd.n3052 vdd.n623 39.2114
R18388 vdd.n3050 vdd.n3049 39.2114
R18389 vdd.n3045 vdd.n629 39.2114
R18390 vdd.n2538 vdd.n2513 39.2114
R18391 vdd.n2542 vdd.n2514 39.2114
R18392 vdd.n2546 vdd.n2515 39.2114
R18393 vdd.n2550 vdd.n2516 39.2114
R18394 vdd.n2554 vdd.n2517 39.2114
R18395 vdd.n2558 vdd.n2518 39.2114
R18396 vdd.n2562 vdd.n2519 39.2114
R18397 vdd.n2566 vdd.n2520 39.2114
R18398 vdd.n2570 vdd.n2521 39.2114
R18399 vdd.n2574 vdd.n2522 39.2114
R18400 vdd.n2578 vdd.n2523 39.2114
R18401 vdd.n2582 vdd.n2524 39.2114
R18402 vdd.n2586 vdd.n2525 39.2114
R18403 vdd.n2590 vdd.n2526 39.2114
R18404 vdd.n2594 vdd.n2527 39.2114
R18405 vdd.n2598 vdd.n2528 39.2114
R18406 vdd.n2602 vdd.n2529 39.2114
R18407 vdd.n2541 vdd.n2513 39.2114
R18408 vdd.n2545 vdd.n2514 39.2114
R18409 vdd.n2549 vdd.n2515 39.2114
R18410 vdd.n2553 vdd.n2516 39.2114
R18411 vdd.n2557 vdd.n2517 39.2114
R18412 vdd.n2561 vdd.n2518 39.2114
R18413 vdd.n2565 vdd.n2519 39.2114
R18414 vdd.n2569 vdd.n2520 39.2114
R18415 vdd.n2573 vdd.n2521 39.2114
R18416 vdd.n2577 vdd.n2522 39.2114
R18417 vdd.n2581 vdd.n2523 39.2114
R18418 vdd.n2585 vdd.n2524 39.2114
R18419 vdd.n2589 vdd.n2525 39.2114
R18420 vdd.n2593 vdd.n2526 39.2114
R18421 vdd.n2597 vdd.n2527 39.2114
R18422 vdd.n2601 vdd.n2528 39.2114
R18423 vdd.n2604 vdd.n2529 39.2114
R18424 vdd.n629 vdd.n624 39.2114
R18425 vdd.n3051 vdd.n3050 39.2114
R18426 vdd.n623 vdd.n621 39.2114
R18427 vdd.n3058 vdd.n3057 39.2114
R18428 vdd.n620 vdd.n618 39.2114
R18429 vdd.n3065 vdd.n3064 39.2114
R18430 vdd.n617 vdd.n615 39.2114
R18431 vdd.n3072 vdd.n3071 39.2114
R18432 vdd.n3075 vdd.n3074 39.2114
R18433 vdd.n2931 vdd.n2930 39.2114
R18434 vdd.n2936 vdd.n2935 39.2114
R18435 vdd.n2929 vdd.n2927 39.2114
R18436 vdd.n2943 vdd.n2942 39.2114
R18437 vdd.n2926 vdd.n2924 39.2114
R18438 vdd.n2950 vdd.n2949 39.2114
R18439 vdd.n2923 vdd.n2921 39.2114
R18440 vdd.n2957 vdd.n2956 39.2114
R18441 vdd.n2219 vdd.n968 39.2114
R18442 vdd.n2213 vdd.n970 39.2114
R18443 vdd.n2209 vdd.n971 39.2114
R18444 vdd.n2205 vdd.n972 39.2114
R18445 vdd.n2201 vdd.n973 39.2114
R18446 vdd.n2197 vdd.n974 39.2114
R18447 vdd.n2193 vdd.n975 39.2114
R18448 vdd.n2189 vdd.n976 39.2114
R18449 vdd.n1149 vdd.n977 39.2114
R18450 vdd.n1153 vdd.n978 39.2114
R18451 vdd.n1157 vdd.n979 39.2114
R18452 vdd.n1161 vdd.n980 39.2114
R18453 vdd.n1165 vdd.n981 39.2114
R18454 vdd.n1169 vdd.n982 39.2114
R18455 vdd.n1173 vdd.n983 39.2114
R18456 vdd.n1178 vdd.n984 39.2114
R18457 vdd.n1182 vdd.n985 39.2114
R18458 vdd.n2429 vdd.n809 39.2114
R18459 vdd.n2434 vdd.n810 39.2114
R18460 vdd.n2438 vdd.n811 39.2114
R18461 vdd.n2442 vdd.n812 39.2114
R18462 vdd.n2446 vdd.n813 39.2114
R18463 vdd.n2450 vdd.n814 39.2114
R18464 vdd.n2454 vdd.n815 39.2114
R18465 vdd.n2458 vdd.n816 39.2114
R18466 vdd.n2462 vdd.n817 39.2114
R18467 vdd.n2466 vdd.n818 39.2114
R18468 vdd.n2470 vdd.n819 39.2114
R18469 vdd.n2474 vdd.n820 39.2114
R18470 vdd.n2478 vdd.n821 39.2114
R18471 vdd.n2482 vdd.n822 39.2114
R18472 vdd.n2486 vdd.n823 39.2114
R18473 vdd.n2490 vdd.n824 39.2114
R18474 vdd.n827 vdd.n825 39.2114
R18475 vdd.n2801 vdd.n790 39.2114
R18476 vdd.n2795 vdd.n2497 39.2114
R18477 vdd.n2791 vdd.n2498 39.2114
R18478 vdd.n2787 vdd.n2499 39.2114
R18479 vdd.n2783 vdd.n2500 39.2114
R18480 vdd.n2779 vdd.n2501 39.2114
R18481 vdd.n2775 vdd.n2502 39.2114
R18482 vdd.n2771 vdd.n2503 39.2114
R18483 vdd.n2767 vdd.n2504 39.2114
R18484 vdd.n2763 vdd.n2505 39.2114
R18485 vdd.n2759 vdd.n2506 39.2114
R18486 vdd.n2755 vdd.n2507 39.2114
R18487 vdd.n2751 vdd.n2508 39.2114
R18488 vdd.n2747 vdd.n2509 39.2114
R18489 vdd.n2743 vdd.n2510 39.2114
R18490 vdd.n2738 vdd.n2511 39.2114
R18491 vdd.n2734 vdd.n2512 39.2114
R18492 vdd.n2978 vdd.n660 39.2114
R18493 vdd.n2985 vdd.n2984 39.2114
R18494 vdd.n659 vdd.n657 39.2114
R18495 vdd.n2992 vdd.n2991 39.2114
R18496 vdd.n656 vdd.n654 39.2114
R18497 vdd.n2999 vdd.n2998 39.2114
R18498 vdd.n653 vdd.n651 39.2114
R18499 vdd.n3006 vdd.n3005 39.2114
R18500 vdd.n650 vdd.n648 39.2114
R18501 vdd.n3014 vdd.n3013 39.2114
R18502 vdd.n647 vdd.n645 39.2114
R18503 vdd.n3021 vdd.n3020 39.2114
R18504 vdd.n644 vdd.n642 39.2114
R18505 vdd.n3028 vdd.n3027 39.2114
R18506 vdd.n641 vdd.n639 39.2114
R18507 vdd.n3035 vdd.n3034 39.2114
R18508 vdd.n3038 vdd.n3037 39.2114
R18509 vdd.n836 vdd.n791 39.2114
R18510 vdd.n2418 vdd.n792 39.2114
R18511 vdd.n2414 vdd.n793 39.2114
R18512 vdd.n2410 vdd.n794 39.2114
R18513 vdd.n2406 vdd.n795 39.2114
R18514 vdd.n2402 vdd.n796 39.2114
R18515 vdd.n2398 vdd.n797 39.2114
R18516 vdd.n2394 vdd.n798 39.2114
R18517 vdd.n2390 vdd.n799 39.2114
R18518 vdd.n2386 vdd.n800 39.2114
R18519 vdd.n2382 vdd.n801 39.2114
R18520 vdd.n2378 vdd.n802 39.2114
R18521 vdd.n2374 vdd.n803 39.2114
R18522 vdd.n2370 vdd.n804 39.2114
R18523 vdd.n2366 vdd.n805 39.2114
R18524 vdd.n2362 vdd.n806 39.2114
R18525 vdd.n2358 vdd.n807 39.2114
R18526 vdd.n1108 vdd.n986 39.2114
R18527 vdd.n1112 vdd.n987 39.2114
R18528 vdd.n1116 vdd.n988 39.2114
R18529 vdd.n1120 vdd.n989 39.2114
R18530 vdd.n1124 vdd.n990 39.2114
R18531 vdd.n1128 vdd.n991 39.2114
R18532 vdd.n1132 vdd.n992 39.2114
R18533 vdd.n1136 vdd.n993 39.2114
R18534 vdd.n1140 vdd.n994 39.2114
R18535 vdd.n1341 vdd.n995 39.2114
R18536 vdd.n1338 vdd.n996 39.2114
R18537 vdd.n1334 vdd.n997 39.2114
R18538 vdd.n1330 vdd.n998 39.2114
R18539 vdd.n1326 vdd.n999 39.2114
R18540 vdd.n1322 vdd.n1000 39.2114
R18541 vdd.n1318 vdd.n1001 39.2114
R18542 vdd.n1314 vdd.n1002 39.2114
R18543 vdd.n2355 vdd.n807 39.2114
R18544 vdd.n2359 vdd.n806 39.2114
R18545 vdd.n2363 vdd.n805 39.2114
R18546 vdd.n2367 vdd.n804 39.2114
R18547 vdd.n2371 vdd.n803 39.2114
R18548 vdd.n2375 vdd.n802 39.2114
R18549 vdd.n2379 vdd.n801 39.2114
R18550 vdd.n2383 vdd.n800 39.2114
R18551 vdd.n2387 vdd.n799 39.2114
R18552 vdd.n2391 vdd.n798 39.2114
R18553 vdd.n2395 vdd.n797 39.2114
R18554 vdd.n2399 vdd.n796 39.2114
R18555 vdd.n2403 vdd.n795 39.2114
R18556 vdd.n2407 vdd.n794 39.2114
R18557 vdd.n2411 vdd.n793 39.2114
R18558 vdd.n2415 vdd.n792 39.2114
R18559 vdd.n2419 vdd.n791 39.2114
R18560 vdd.n1111 vdd.n986 39.2114
R18561 vdd.n1115 vdd.n987 39.2114
R18562 vdd.n1119 vdd.n988 39.2114
R18563 vdd.n1123 vdd.n989 39.2114
R18564 vdd.n1127 vdd.n990 39.2114
R18565 vdd.n1131 vdd.n991 39.2114
R18566 vdd.n1135 vdd.n992 39.2114
R18567 vdd.n1139 vdd.n993 39.2114
R18568 vdd.n1142 vdd.n994 39.2114
R18569 vdd.n1339 vdd.n995 39.2114
R18570 vdd.n1335 vdd.n996 39.2114
R18571 vdd.n1331 vdd.n997 39.2114
R18572 vdd.n1327 vdd.n998 39.2114
R18573 vdd.n1323 vdd.n999 39.2114
R18574 vdd.n1319 vdd.n1000 39.2114
R18575 vdd.n1315 vdd.n1001 39.2114
R18576 vdd.n1311 vdd.n1002 39.2114
R18577 vdd.n2076 vdd.n2075 37.2369
R18578 vdd.n2112 vdd.n1077 37.2369
R18579 vdd.n2151 vdd.n1037 37.2369
R18580 vdd.n3126 vdd.n581 37.2369
R18581 vdd.n545 vdd.n544 37.2369
R18582 vdd.n3082 vdd.n3081 37.2369
R18583 vdd.n1145 vdd.n1144 30.449
R18584 vdd.n840 vdd.n839 30.449
R18585 vdd.n1176 vdd.n1148 30.449
R18586 vdd.n2432 vdd.n830 30.449
R18587 vdd.n2537 vdd.n2536 30.449
R18588 vdd.n663 vdd.n662 30.449
R18589 vdd.n2740 vdd.n2533 30.449
R18590 vdd.n627 vdd.n626 30.449
R18591 vdd.n2222 vdd.n2221 29.8151
R18592 vdd.n2494 vdd.n828 29.8151
R18593 vdd.n2427 vdd.n831 29.8151
R18594 vdd.n1184 vdd.n1181 29.8151
R18595 vdd.n2735 vdd.n2732 29.8151
R18596 vdd.n2980 vdd.n2977 29.8151
R18597 vdd.n2804 vdd.n2803 29.8151
R18598 vdd.n3041 vdd.n3040 29.8151
R18599 vdd.n2960 vdd.n2959 29.8151
R18600 vdd.n3046 vdd.n628 29.8151
R18601 vdd.n2608 vdd.n2606 29.8151
R18602 vdd.n2539 vdd.n783 29.8151
R18603 vdd.n1109 vdd.n960 29.8151
R18604 vdd.n2422 vdd.n2421 29.8151
R18605 vdd.n2354 vdd.n2353 29.8151
R18606 vdd.n1310 vdd.n1309 29.8151
R18607 vdd.n1670 vdd.n1437 20.633
R18608 vdd.n2070 vdd.n969 20.633
R18609 vdd.n3212 vdd.n516 20.633
R18610 vdd.n3410 vdd.n351 20.633
R18611 vdd.n1672 vdd.n1434 19.3944
R18612 vdd.n1676 vdd.n1434 19.3944
R18613 vdd.n1676 vdd.n1425 19.3944
R18614 vdd.n1688 vdd.n1425 19.3944
R18615 vdd.n1688 vdd.n1423 19.3944
R18616 vdd.n1692 vdd.n1423 19.3944
R18617 vdd.n1692 vdd.n1412 19.3944
R18618 vdd.n1704 vdd.n1412 19.3944
R18619 vdd.n1704 vdd.n1410 19.3944
R18620 vdd.n1708 vdd.n1410 19.3944
R18621 vdd.n1708 vdd.n1401 19.3944
R18622 vdd.n1721 vdd.n1401 19.3944
R18623 vdd.n1721 vdd.n1399 19.3944
R18624 vdd.n1725 vdd.n1399 19.3944
R18625 vdd.n1725 vdd.n1390 19.3944
R18626 vdd.n2019 vdd.n1390 19.3944
R18627 vdd.n2019 vdd.n1388 19.3944
R18628 vdd.n2023 vdd.n1388 19.3944
R18629 vdd.n2023 vdd.n1378 19.3944
R18630 vdd.n2036 vdd.n1378 19.3944
R18631 vdd.n2036 vdd.n1376 19.3944
R18632 vdd.n2040 vdd.n1376 19.3944
R18633 vdd.n2040 vdd.n1368 19.3944
R18634 vdd.n2053 vdd.n1368 19.3944
R18635 vdd.n2053 vdd.n1365 19.3944
R18636 vdd.n2059 vdd.n1365 19.3944
R18637 vdd.n2059 vdd.n1366 19.3944
R18638 vdd.n1366 vdd.n1356 19.3944
R18639 vdd.n1597 vdd.n1523 19.3944
R18640 vdd.n1597 vdd.n1525 19.3944
R18641 vdd.n1593 vdd.n1525 19.3944
R18642 vdd.n1593 vdd.n1592 19.3944
R18643 vdd.n1592 vdd.n1591 19.3944
R18644 vdd.n1591 vdd.n1533 19.3944
R18645 vdd.n1587 vdd.n1533 19.3944
R18646 vdd.n1587 vdd.n1586 19.3944
R18647 vdd.n1586 vdd.n1585 19.3944
R18648 vdd.n1585 vdd.n1541 19.3944
R18649 vdd.n1581 vdd.n1541 19.3944
R18650 vdd.n1581 vdd.n1580 19.3944
R18651 vdd.n1580 vdd.n1579 19.3944
R18652 vdd.n1579 vdd.n1549 19.3944
R18653 vdd.n1575 vdd.n1549 19.3944
R18654 vdd.n1575 vdd.n1574 19.3944
R18655 vdd.n1574 vdd.n1573 19.3944
R18656 vdd.n1573 vdd.n1557 19.3944
R18657 vdd.n1569 vdd.n1557 19.3944
R18658 vdd.n1569 vdd.n1568 19.3944
R18659 vdd.n1635 vdd.n1634 19.3944
R18660 vdd.n1634 vdd.n1633 19.3944
R18661 vdd.n1633 vdd.n1486 19.3944
R18662 vdd.n1629 vdd.n1486 19.3944
R18663 vdd.n1629 vdd.n1628 19.3944
R18664 vdd.n1628 vdd.n1627 19.3944
R18665 vdd.n1627 vdd.n1494 19.3944
R18666 vdd.n1623 vdd.n1494 19.3944
R18667 vdd.n1623 vdd.n1622 19.3944
R18668 vdd.n1622 vdd.n1621 19.3944
R18669 vdd.n1621 vdd.n1502 19.3944
R18670 vdd.n1617 vdd.n1502 19.3944
R18671 vdd.n1617 vdd.n1616 19.3944
R18672 vdd.n1616 vdd.n1615 19.3944
R18673 vdd.n1615 vdd.n1510 19.3944
R18674 vdd.n1611 vdd.n1510 19.3944
R18675 vdd.n1611 vdd.n1610 19.3944
R18676 vdd.n1610 vdd.n1609 19.3944
R18677 vdd.n1609 vdd.n1518 19.3944
R18678 vdd.n1605 vdd.n1518 19.3944
R18679 vdd.n1665 vdd.n1664 19.3944
R18680 vdd.n1664 vdd.n1663 19.3944
R18681 vdd.n1663 vdd.n1444 19.3944
R18682 vdd.n1659 vdd.n1444 19.3944
R18683 vdd.n1659 vdd.n1658 19.3944
R18684 vdd.n1658 vdd.n1657 19.3944
R18685 vdd.n1657 vdd.n1452 19.3944
R18686 vdd.n1653 vdd.n1452 19.3944
R18687 vdd.n1653 vdd.n1652 19.3944
R18688 vdd.n1652 vdd.n1651 19.3944
R18689 vdd.n1651 vdd.n1460 19.3944
R18690 vdd.n1647 vdd.n1460 19.3944
R18691 vdd.n1647 vdd.n1646 19.3944
R18692 vdd.n1646 vdd.n1645 19.3944
R18693 vdd.n1645 vdd.n1468 19.3944
R18694 vdd.n1641 vdd.n1468 19.3944
R18695 vdd.n1641 vdd.n1640 19.3944
R18696 vdd.n1640 vdd.n1639 19.3944
R18697 vdd.n2108 vdd.n1075 19.3944
R18698 vdd.n2108 vdd.n1081 19.3944
R18699 vdd.n2103 vdd.n1081 19.3944
R18700 vdd.n2103 vdd.n2102 19.3944
R18701 vdd.n2102 vdd.n2101 19.3944
R18702 vdd.n2101 vdd.n1088 19.3944
R18703 vdd.n2096 vdd.n1088 19.3944
R18704 vdd.n2096 vdd.n2095 19.3944
R18705 vdd.n2095 vdd.n2094 19.3944
R18706 vdd.n2094 vdd.n1095 19.3944
R18707 vdd.n2089 vdd.n1095 19.3944
R18708 vdd.n2089 vdd.n2088 19.3944
R18709 vdd.n2088 vdd.n2087 19.3944
R18710 vdd.n2087 vdd.n1102 19.3944
R18711 vdd.n2082 vdd.n1102 19.3944
R18712 vdd.n2082 vdd.n2081 19.3944
R18713 vdd.n1349 vdd.n1107 19.3944
R18714 vdd.n2077 vdd.n1346 19.3944
R18715 vdd.n2147 vdd.n1035 19.3944
R18716 vdd.n2147 vdd.n1041 19.3944
R18717 vdd.n2142 vdd.n1041 19.3944
R18718 vdd.n2142 vdd.n2141 19.3944
R18719 vdd.n2141 vdd.n2140 19.3944
R18720 vdd.n2140 vdd.n1048 19.3944
R18721 vdd.n2135 vdd.n1048 19.3944
R18722 vdd.n2135 vdd.n2134 19.3944
R18723 vdd.n2134 vdd.n2133 19.3944
R18724 vdd.n2133 vdd.n1055 19.3944
R18725 vdd.n2128 vdd.n1055 19.3944
R18726 vdd.n2128 vdd.n2127 19.3944
R18727 vdd.n2127 vdd.n2126 19.3944
R18728 vdd.n2126 vdd.n1062 19.3944
R18729 vdd.n2121 vdd.n1062 19.3944
R18730 vdd.n2121 vdd.n2120 19.3944
R18731 vdd.n2120 vdd.n2119 19.3944
R18732 vdd.n2119 vdd.n1069 19.3944
R18733 vdd.n2114 vdd.n1069 19.3944
R18734 vdd.n2114 vdd.n2113 19.3944
R18735 vdd.n2184 vdd.n1010 19.3944
R18736 vdd.n2184 vdd.n1011 19.3944
R18737 vdd.n2179 vdd.n2178 19.3944
R18738 vdd.n2174 vdd.n2173 19.3944
R18739 vdd.n2173 vdd.n2172 19.3944
R18740 vdd.n2172 vdd.n1015 19.3944
R18741 vdd.n2167 vdd.n1015 19.3944
R18742 vdd.n2167 vdd.n2166 19.3944
R18743 vdd.n2166 vdd.n2165 19.3944
R18744 vdd.n2165 vdd.n1022 19.3944
R18745 vdd.n2160 vdd.n1022 19.3944
R18746 vdd.n2160 vdd.n2159 19.3944
R18747 vdd.n2159 vdd.n2158 19.3944
R18748 vdd.n2158 vdd.n1029 19.3944
R18749 vdd.n2153 vdd.n1029 19.3944
R18750 vdd.n2153 vdd.n2152 19.3944
R18751 vdd.n1668 vdd.n1431 19.3944
R18752 vdd.n1680 vdd.n1431 19.3944
R18753 vdd.n1680 vdd.n1429 19.3944
R18754 vdd.n1684 vdd.n1429 19.3944
R18755 vdd.n1684 vdd.n1419 19.3944
R18756 vdd.n1696 vdd.n1419 19.3944
R18757 vdd.n1696 vdd.n1417 19.3944
R18758 vdd.n1700 vdd.n1417 19.3944
R18759 vdd.n1700 vdd.n1407 19.3944
R18760 vdd.n1713 vdd.n1407 19.3944
R18761 vdd.n1713 vdd.n1405 19.3944
R18762 vdd.n1717 vdd.n1405 19.3944
R18763 vdd.n1717 vdd.n1396 19.3944
R18764 vdd.n1729 vdd.n1396 19.3944
R18765 vdd.n1729 vdd.n1394 19.3944
R18766 vdd.n2015 vdd.n1394 19.3944
R18767 vdd.n2015 vdd.n1384 19.3944
R18768 vdd.n2028 vdd.n1384 19.3944
R18769 vdd.n2028 vdd.n1382 19.3944
R18770 vdd.n2032 vdd.n1382 19.3944
R18771 vdd.n2032 vdd.n1373 19.3944
R18772 vdd.n2045 vdd.n1373 19.3944
R18773 vdd.n2045 vdd.n1371 19.3944
R18774 vdd.n2049 vdd.n1371 19.3944
R18775 vdd.n2049 vdd.n1361 19.3944
R18776 vdd.n2064 vdd.n1361 19.3944
R18777 vdd.n2064 vdd.n1359 19.3944
R18778 vdd.n2068 vdd.n1359 19.3944
R18779 vdd.n3214 vdd.n513 19.3944
R18780 vdd.n3218 vdd.n513 19.3944
R18781 vdd.n3218 vdd.n503 19.3944
R18782 vdd.n3230 vdd.n503 19.3944
R18783 vdd.n3230 vdd.n501 19.3944
R18784 vdd.n3234 vdd.n501 19.3944
R18785 vdd.n3234 vdd.n490 19.3944
R18786 vdd.n3246 vdd.n490 19.3944
R18787 vdd.n3246 vdd.n488 19.3944
R18788 vdd.n3250 vdd.n488 19.3944
R18789 vdd.n3250 vdd.n478 19.3944
R18790 vdd.n3263 vdd.n478 19.3944
R18791 vdd.n3263 vdd.n476 19.3944
R18792 vdd.n3267 vdd.n476 19.3944
R18793 vdd.n3268 vdd.n3267 19.3944
R18794 vdd.n3269 vdd.n3268 19.3944
R18795 vdd.n3269 vdd.n474 19.3944
R18796 vdd.n3273 vdd.n474 19.3944
R18797 vdd.n3274 vdd.n3273 19.3944
R18798 vdd.n3275 vdd.n3274 19.3944
R18799 vdd.n3275 vdd.n471 19.3944
R18800 vdd.n3279 vdd.n471 19.3944
R18801 vdd.n3280 vdd.n3279 19.3944
R18802 vdd.n3281 vdd.n3280 19.3944
R18803 vdd.n3281 vdd.n468 19.3944
R18804 vdd.n3285 vdd.n468 19.3944
R18805 vdd.n3286 vdd.n3285 19.3944
R18806 vdd.n3287 vdd.n3286 19.3944
R18807 vdd.n3330 vdd.n426 19.3944
R18808 vdd.n3330 vdd.n432 19.3944
R18809 vdd.n3325 vdd.n432 19.3944
R18810 vdd.n3325 vdd.n3324 19.3944
R18811 vdd.n3324 vdd.n3323 19.3944
R18812 vdd.n3323 vdd.n439 19.3944
R18813 vdd.n3318 vdd.n439 19.3944
R18814 vdd.n3318 vdd.n3317 19.3944
R18815 vdd.n3317 vdd.n3316 19.3944
R18816 vdd.n3316 vdd.n446 19.3944
R18817 vdd.n3311 vdd.n446 19.3944
R18818 vdd.n3311 vdd.n3310 19.3944
R18819 vdd.n3310 vdd.n3309 19.3944
R18820 vdd.n3309 vdd.n453 19.3944
R18821 vdd.n3304 vdd.n453 19.3944
R18822 vdd.n3304 vdd.n3303 19.3944
R18823 vdd.n3303 vdd.n3302 19.3944
R18824 vdd.n3302 vdd.n460 19.3944
R18825 vdd.n3297 vdd.n460 19.3944
R18826 vdd.n3297 vdd.n3296 19.3944
R18827 vdd.n3369 vdd.n386 19.3944
R18828 vdd.n3369 vdd.n392 19.3944
R18829 vdd.n3364 vdd.n392 19.3944
R18830 vdd.n3364 vdd.n3363 19.3944
R18831 vdd.n3363 vdd.n3362 19.3944
R18832 vdd.n3362 vdd.n399 19.3944
R18833 vdd.n3357 vdd.n399 19.3944
R18834 vdd.n3357 vdd.n3356 19.3944
R18835 vdd.n3356 vdd.n3355 19.3944
R18836 vdd.n3355 vdd.n406 19.3944
R18837 vdd.n3350 vdd.n406 19.3944
R18838 vdd.n3350 vdd.n3349 19.3944
R18839 vdd.n3349 vdd.n3348 19.3944
R18840 vdd.n3348 vdd.n413 19.3944
R18841 vdd.n3343 vdd.n413 19.3944
R18842 vdd.n3343 vdd.n3342 19.3944
R18843 vdd.n3342 vdd.n3341 19.3944
R18844 vdd.n3341 vdd.n420 19.3944
R18845 vdd.n3336 vdd.n420 19.3944
R18846 vdd.n3336 vdd.n3335 19.3944
R18847 vdd.n3405 vdd.n3404 19.3944
R18848 vdd.n3404 vdd.n3403 19.3944
R18849 vdd.n3403 vdd.n358 19.3944
R18850 vdd.n359 vdd.n358 19.3944
R18851 vdd.n3396 vdd.n359 19.3944
R18852 vdd.n3396 vdd.n3395 19.3944
R18853 vdd.n3395 vdd.n3394 19.3944
R18854 vdd.n3394 vdd.n366 19.3944
R18855 vdd.n3389 vdd.n366 19.3944
R18856 vdd.n3389 vdd.n3388 19.3944
R18857 vdd.n3388 vdd.n3387 19.3944
R18858 vdd.n3387 vdd.n373 19.3944
R18859 vdd.n3382 vdd.n373 19.3944
R18860 vdd.n3382 vdd.n3381 19.3944
R18861 vdd.n3381 vdd.n3380 19.3944
R18862 vdd.n3380 vdd.n380 19.3944
R18863 vdd.n3375 vdd.n380 19.3944
R18864 vdd.n3375 vdd.n3374 19.3944
R18865 vdd.n3210 vdd.n509 19.3944
R18866 vdd.n3222 vdd.n509 19.3944
R18867 vdd.n3222 vdd.n507 19.3944
R18868 vdd.n3226 vdd.n507 19.3944
R18869 vdd.n3226 vdd.n497 19.3944
R18870 vdd.n3238 vdd.n497 19.3944
R18871 vdd.n3238 vdd.n495 19.3944
R18872 vdd.n3242 vdd.n495 19.3944
R18873 vdd.n3242 vdd.n485 19.3944
R18874 vdd.n3255 vdd.n485 19.3944
R18875 vdd.n3255 vdd.n483 19.3944
R18876 vdd.n3259 vdd.n483 19.3944
R18877 vdd.n3259 vdd.n312 19.3944
R18878 vdd.n3438 vdd.n312 19.3944
R18879 vdd.n3438 vdd.n313 19.3944
R18880 vdd.n3432 vdd.n313 19.3944
R18881 vdd.n3432 vdd.n3431 19.3944
R18882 vdd.n3431 vdd.n3430 19.3944
R18883 vdd.n3430 vdd.n323 19.3944
R18884 vdd.n3424 vdd.n323 19.3944
R18885 vdd.n3424 vdd.n3423 19.3944
R18886 vdd.n3423 vdd.n3422 19.3944
R18887 vdd.n3422 vdd.n335 19.3944
R18888 vdd.n3416 vdd.n335 19.3944
R18889 vdd.n3416 vdd.n3415 19.3944
R18890 vdd.n3415 vdd.n3414 19.3944
R18891 vdd.n3414 vdd.n346 19.3944
R18892 vdd.n3408 vdd.n346 19.3944
R18893 vdd.n3167 vdd.n3166 19.3944
R18894 vdd.n3166 vdd.n3165 19.3944
R18895 vdd.n3165 vdd.n551 19.3944
R18896 vdd.n3159 vdd.n551 19.3944
R18897 vdd.n3159 vdd.n3158 19.3944
R18898 vdd.n3158 vdd.n3157 19.3944
R18899 vdd.n3157 vdd.n557 19.3944
R18900 vdd.n3151 vdd.n557 19.3944
R18901 vdd.n3151 vdd.n3150 19.3944
R18902 vdd.n3150 vdd.n3149 19.3944
R18903 vdd.n3149 vdd.n563 19.3944
R18904 vdd.n3143 vdd.n563 19.3944
R18905 vdd.n3143 vdd.n3142 19.3944
R18906 vdd.n3142 vdd.n3141 19.3944
R18907 vdd.n3141 vdd.n569 19.3944
R18908 vdd.n3135 vdd.n569 19.3944
R18909 vdd.n3135 vdd.n3134 19.3944
R18910 vdd.n3134 vdd.n3133 19.3944
R18911 vdd.n3133 vdd.n575 19.3944
R18912 vdd.n3127 vdd.n575 19.3944
R18913 vdd.n3207 vdd.n3206 19.3944
R18914 vdd.n3206 vdd.n519 19.3944
R18915 vdd.n3201 vdd.n3200 19.3944
R18916 vdd.n3197 vdd.n3196 19.3944
R18917 vdd.n3196 vdd.n525 19.3944
R18918 vdd.n3191 vdd.n525 19.3944
R18919 vdd.n3191 vdd.n3190 19.3944
R18920 vdd.n3190 vdd.n3189 19.3944
R18921 vdd.n3189 vdd.n531 19.3944
R18922 vdd.n3183 vdd.n531 19.3944
R18923 vdd.n3183 vdd.n3182 19.3944
R18924 vdd.n3182 vdd.n3181 19.3944
R18925 vdd.n3181 vdd.n537 19.3944
R18926 vdd.n3175 vdd.n537 19.3944
R18927 vdd.n3175 vdd.n3174 19.3944
R18928 vdd.n3174 vdd.n3173 19.3944
R18929 vdd.n3122 vdd.n579 19.3944
R18930 vdd.n3122 vdd.n583 19.3944
R18931 vdd.n3117 vdd.n583 19.3944
R18932 vdd.n3117 vdd.n3116 19.3944
R18933 vdd.n3116 vdd.n589 19.3944
R18934 vdd.n3111 vdd.n589 19.3944
R18935 vdd.n3111 vdd.n3110 19.3944
R18936 vdd.n3110 vdd.n3109 19.3944
R18937 vdd.n3109 vdd.n595 19.3944
R18938 vdd.n3103 vdd.n595 19.3944
R18939 vdd.n3103 vdd.n3102 19.3944
R18940 vdd.n3102 vdd.n3101 19.3944
R18941 vdd.n3101 vdd.n601 19.3944
R18942 vdd.n3095 vdd.n601 19.3944
R18943 vdd.n3095 vdd.n3094 19.3944
R18944 vdd.n3094 vdd.n3093 19.3944
R18945 vdd.n3089 vdd.n3088 19.3944
R18946 vdd.n3085 vdd.n3084 19.3944
R18947 vdd.n1604 vdd.n1523 19.0066
R18948 vdd.n2112 vdd.n1075 19.0066
R18949 vdd.n3334 vdd.n426 19.0066
R18950 vdd.n3126 vdd.n579 19.0066
R18951 vdd.n1144 vdd.n1143 16.0975
R18952 vdd.n839 vdd.n838 16.0975
R18953 vdd.n1566 vdd.n1565 16.0975
R18954 vdd.n1603 vdd.n1602 16.0975
R18955 vdd.n1477 vdd.n1476 16.0975
R18956 vdd.n2075 vdd.n2074 16.0975
R18957 vdd.n1077 vdd.n1076 16.0975
R18958 vdd.n1037 vdd.n1036 16.0975
R18959 vdd.n1148 vdd.n1147 16.0975
R18960 vdd.n830 vdd.n829 16.0975
R18961 vdd.n2536 vdd.n2535 16.0975
R18962 vdd.n3294 vdd.n3293 16.0975
R18963 vdd.n428 vdd.n427 16.0975
R18964 vdd.n388 vdd.n387 16.0975
R18965 vdd.n581 vdd.n580 16.0975
R18966 vdd.n544 vdd.n543 16.0975
R18967 vdd.n662 vdd.n661 16.0975
R18968 vdd.n2533 vdd.n2532 16.0975
R18969 vdd.n3081 vdd.n3080 16.0975
R18970 vdd.n626 vdd.n625 16.0975
R18971 vdd.t29 vdd.n2496 15.4182
R18972 vdd.n2800 vdd.t16 15.4182
R18973 vdd.n28 vdd.n27 14.5674
R18974 vdd.n304 vdd.n269 13.1884
R18975 vdd.n253 vdd.n218 13.1884
R18976 vdd.n210 vdd.n175 13.1884
R18977 vdd.n159 vdd.n124 13.1884
R18978 vdd.n117 vdd.n82 13.1884
R18979 vdd.n66 vdd.n31 13.1884
R18980 vdd.n1954 vdd.n1919 13.1884
R18981 vdd.n2005 vdd.n1970 13.1884
R18982 vdd.n1860 vdd.n1825 13.1884
R18983 vdd.n1911 vdd.n1876 13.1884
R18984 vdd.n1767 vdd.n1732 13.1884
R18985 vdd.n1818 vdd.n1783 13.1884
R18986 vdd.n2218 vdd.n962 13.1509
R18987 vdd.n3043 vdd.n613 13.1509
R18988 vdd.n1635 vdd.n1478 12.9944
R18989 vdd.n1639 vdd.n1478 12.9944
R18990 vdd.n2151 vdd.n1035 12.9944
R18991 vdd.n2152 vdd.n2151 12.9944
R18992 vdd.n3373 vdd.n386 12.9944
R18993 vdd.n3374 vdd.n3373 12.9944
R18994 vdd.n3167 vdd.n545 12.9944
R18995 vdd.n3173 vdd.n545 12.9944
R18996 vdd.n305 vdd.n267 12.8005
R18997 vdd.n300 vdd.n271 12.8005
R18998 vdd.n254 vdd.n216 12.8005
R18999 vdd.n249 vdd.n220 12.8005
R19000 vdd.n211 vdd.n173 12.8005
R19001 vdd.n206 vdd.n177 12.8005
R19002 vdd.n160 vdd.n122 12.8005
R19003 vdd.n155 vdd.n126 12.8005
R19004 vdd.n118 vdd.n80 12.8005
R19005 vdd.n113 vdd.n84 12.8005
R19006 vdd.n67 vdd.n29 12.8005
R19007 vdd.n62 vdd.n33 12.8005
R19008 vdd.n1955 vdd.n1917 12.8005
R19009 vdd.n1950 vdd.n1921 12.8005
R19010 vdd.n2006 vdd.n1968 12.8005
R19011 vdd.n2001 vdd.n1972 12.8005
R19012 vdd.n1861 vdd.n1823 12.8005
R19013 vdd.n1856 vdd.n1827 12.8005
R19014 vdd.n1912 vdd.n1874 12.8005
R19015 vdd.n1907 vdd.n1878 12.8005
R19016 vdd.n1768 vdd.n1730 12.8005
R19017 vdd.n1763 vdd.n1734 12.8005
R19018 vdd.n1819 vdd.n1781 12.8005
R19019 vdd.n1814 vdd.n1785 12.8005
R19020 vdd.n299 vdd.n272 12.0247
R19021 vdd.n248 vdd.n221 12.0247
R19022 vdd.n205 vdd.n178 12.0247
R19023 vdd.n154 vdd.n127 12.0247
R19024 vdd.n112 vdd.n85 12.0247
R19025 vdd.n61 vdd.n34 12.0247
R19026 vdd.n1949 vdd.n1922 12.0247
R19027 vdd.n2000 vdd.n1973 12.0247
R19028 vdd.n1855 vdd.n1828 12.0247
R19029 vdd.n1906 vdd.n1879 12.0247
R19030 vdd.n1762 vdd.n1735 12.0247
R19031 vdd.n1813 vdd.n1786 12.0247
R19032 vdd.n1670 vdd.n1438 11.337
R19033 vdd.n1678 vdd.n1427 11.337
R19034 vdd.n1686 vdd.n1427 11.337
R19035 vdd.n1694 vdd.n1421 11.337
R19036 vdd.n1702 vdd.n1414 11.337
R19037 vdd.n1711 vdd.n1710 11.337
R19038 vdd.n1719 vdd.n1403 11.337
R19039 vdd.n2017 vdd.n1392 11.337
R19040 vdd.n2026 vdd.n1386 11.337
R19041 vdd.n2034 vdd.n1380 11.337
R19042 vdd.n2043 vdd.n2042 11.337
R19043 vdd.n2051 vdd.n1363 11.337
R19044 vdd.n2062 vdd.n1363 11.337
R19045 vdd.n2062 vdd.n2061 11.337
R19046 vdd.n3220 vdd.n511 11.337
R19047 vdd.n3220 vdd.n505 11.337
R19048 vdd.n3228 vdd.n505 11.337
R19049 vdd.n3236 vdd.n499 11.337
R19050 vdd.n3244 vdd.n492 11.337
R19051 vdd.n3253 vdd.n3252 11.337
R19052 vdd.n3261 vdd.n481 11.337
R19053 vdd.n3435 vdd.n3434 11.337
R19054 vdd.n3428 vdd.n325 11.337
R19055 vdd.n3426 vdd.n329 11.337
R19056 vdd.n3420 vdd.n3419 11.337
R19057 vdd.n3418 vdd.n340 11.337
R19058 vdd.n3412 vdd.n340 11.337
R19059 vdd.n3411 vdd.n3410 11.337
R19060 vdd.n296 vdd.n295 11.249
R19061 vdd.n245 vdd.n244 11.249
R19062 vdd.n202 vdd.n201 11.249
R19063 vdd.n151 vdd.n150 11.249
R19064 vdd.n109 vdd.n108 11.249
R19065 vdd.n58 vdd.n57 11.249
R19066 vdd.n1946 vdd.n1945 11.249
R19067 vdd.n1997 vdd.n1996 11.249
R19068 vdd.n1852 vdd.n1851 11.249
R19069 vdd.n1903 vdd.n1902 11.249
R19070 vdd.n1759 vdd.n1758 11.249
R19071 vdd.n1810 vdd.n1809 11.249
R19072 vdd.n1686 vdd.t94 10.9969
R19073 vdd.t72 vdd.n3418 10.9969
R19074 vdd.n1415 vdd.t102 10.7702
R19075 vdd.t64 vdd.n3427 10.7702
R19076 vdd.n281 vdd.n280 10.7238
R19077 vdd.n230 vdd.n229 10.7238
R19078 vdd.n187 vdd.n186 10.7238
R19079 vdd.n136 vdd.n135 10.7238
R19080 vdd.n94 vdd.n93 10.7238
R19081 vdd.n43 vdd.n42 10.7238
R19082 vdd.n1931 vdd.n1930 10.7238
R19083 vdd.n1982 vdd.n1981 10.7238
R19084 vdd.n1837 vdd.n1836 10.7238
R19085 vdd.n1888 vdd.n1887 10.7238
R19086 vdd.n1744 vdd.n1743 10.7238
R19087 vdd.n1795 vdd.n1794 10.7238
R19088 vdd.n2223 vdd.n2222 10.6151
R19089 vdd.n2223 vdd.n955 10.6151
R19090 vdd.n2233 vdd.n955 10.6151
R19091 vdd.n2234 vdd.n2233 10.6151
R19092 vdd.n2235 vdd.n2234 10.6151
R19093 vdd.n2235 vdd.n942 10.6151
R19094 vdd.n2245 vdd.n942 10.6151
R19095 vdd.n2246 vdd.n2245 10.6151
R19096 vdd.n2247 vdd.n2246 10.6151
R19097 vdd.n2247 vdd.n930 10.6151
R19098 vdd.n2257 vdd.n930 10.6151
R19099 vdd.n2258 vdd.n2257 10.6151
R19100 vdd.n2259 vdd.n2258 10.6151
R19101 vdd.n2259 vdd.n919 10.6151
R19102 vdd.n2269 vdd.n919 10.6151
R19103 vdd.n2270 vdd.n2269 10.6151
R19104 vdd.n2271 vdd.n2270 10.6151
R19105 vdd.n2271 vdd.n906 10.6151
R19106 vdd.n2281 vdd.n906 10.6151
R19107 vdd.n2282 vdd.n2281 10.6151
R19108 vdd.n2283 vdd.n2282 10.6151
R19109 vdd.n2283 vdd.n894 10.6151
R19110 vdd.n2294 vdd.n894 10.6151
R19111 vdd.n2295 vdd.n2294 10.6151
R19112 vdd.n2296 vdd.n2295 10.6151
R19113 vdd.n2296 vdd.n882 10.6151
R19114 vdd.n2306 vdd.n882 10.6151
R19115 vdd.n2307 vdd.n2306 10.6151
R19116 vdd.n2308 vdd.n2307 10.6151
R19117 vdd.n2308 vdd.n870 10.6151
R19118 vdd.n2318 vdd.n870 10.6151
R19119 vdd.n2319 vdd.n2318 10.6151
R19120 vdd.n2320 vdd.n2319 10.6151
R19121 vdd.n2320 vdd.n860 10.6151
R19122 vdd.n2330 vdd.n860 10.6151
R19123 vdd.n2331 vdd.n2330 10.6151
R19124 vdd.n2332 vdd.n2331 10.6151
R19125 vdd.n2332 vdd.n847 10.6151
R19126 vdd.n2344 vdd.n847 10.6151
R19127 vdd.n2345 vdd.n2344 10.6151
R19128 vdd.n2347 vdd.n2345 10.6151
R19129 vdd.n2347 vdd.n2346 10.6151
R19130 vdd.n2346 vdd.n828 10.6151
R19131 vdd.n2494 vdd.n2493 10.6151
R19132 vdd.n2493 vdd.n2492 10.6151
R19133 vdd.n2492 vdd.n2489 10.6151
R19134 vdd.n2489 vdd.n2488 10.6151
R19135 vdd.n2488 vdd.n2485 10.6151
R19136 vdd.n2485 vdd.n2484 10.6151
R19137 vdd.n2484 vdd.n2481 10.6151
R19138 vdd.n2481 vdd.n2480 10.6151
R19139 vdd.n2480 vdd.n2477 10.6151
R19140 vdd.n2477 vdd.n2476 10.6151
R19141 vdd.n2476 vdd.n2473 10.6151
R19142 vdd.n2473 vdd.n2472 10.6151
R19143 vdd.n2472 vdd.n2469 10.6151
R19144 vdd.n2469 vdd.n2468 10.6151
R19145 vdd.n2468 vdd.n2465 10.6151
R19146 vdd.n2465 vdd.n2464 10.6151
R19147 vdd.n2464 vdd.n2461 10.6151
R19148 vdd.n2461 vdd.n2460 10.6151
R19149 vdd.n2460 vdd.n2457 10.6151
R19150 vdd.n2457 vdd.n2456 10.6151
R19151 vdd.n2456 vdd.n2453 10.6151
R19152 vdd.n2453 vdd.n2452 10.6151
R19153 vdd.n2452 vdd.n2449 10.6151
R19154 vdd.n2449 vdd.n2448 10.6151
R19155 vdd.n2448 vdd.n2445 10.6151
R19156 vdd.n2445 vdd.n2444 10.6151
R19157 vdd.n2444 vdd.n2441 10.6151
R19158 vdd.n2441 vdd.n2440 10.6151
R19159 vdd.n2440 vdd.n2437 10.6151
R19160 vdd.n2437 vdd.n2436 10.6151
R19161 vdd.n2436 vdd.n2433 10.6151
R19162 vdd.n2431 vdd.n2428 10.6151
R19163 vdd.n2428 vdd.n2427 10.6151
R19164 vdd.n1185 vdd.n1184 10.6151
R19165 vdd.n1187 vdd.n1185 10.6151
R19166 vdd.n1188 vdd.n1187 10.6151
R19167 vdd.n1190 vdd.n1188 10.6151
R19168 vdd.n1191 vdd.n1190 10.6151
R19169 vdd.n1193 vdd.n1191 10.6151
R19170 vdd.n1194 vdd.n1193 10.6151
R19171 vdd.n1196 vdd.n1194 10.6151
R19172 vdd.n1197 vdd.n1196 10.6151
R19173 vdd.n1199 vdd.n1197 10.6151
R19174 vdd.n1200 vdd.n1199 10.6151
R19175 vdd.n1202 vdd.n1200 10.6151
R19176 vdd.n1203 vdd.n1202 10.6151
R19177 vdd.n1205 vdd.n1203 10.6151
R19178 vdd.n1206 vdd.n1205 10.6151
R19179 vdd.n1208 vdd.n1206 10.6151
R19180 vdd.n1209 vdd.n1208 10.6151
R19181 vdd.n1211 vdd.n1209 10.6151
R19182 vdd.n1212 vdd.n1211 10.6151
R19183 vdd.n1214 vdd.n1212 10.6151
R19184 vdd.n1215 vdd.n1214 10.6151
R19185 vdd.n1217 vdd.n1215 10.6151
R19186 vdd.n1218 vdd.n1217 10.6151
R19187 vdd.n1220 vdd.n1218 10.6151
R19188 vdd.n1221 vdd.n1220 10.6151
R19189 vdd.n1223 vdd.n1221 10.6151
R19190 vdd.n1224 vdd.n1223 10.6151
R19191 vdd.n1263 vdd.n1224 10.6151
R19192 vdd.n1263 vdd.n1262 10.6151
R19193 vdd.n1262 vdd.n1261 10.6151
R19194 vdd.n1261 vdd.n1259 10.6151
R19195 vdd.n1259 vdd.n1258 10.6151
R19196 vdd.n1258 vdd.n1256 10.6151
R19197 vdd.n1256 vdd.n1255 10.6151
R19198 vdd.n1255 vdd.n1236 10.6151
R19199 vdd.n1236 vdd.n1235 10.6151
R19200 vdd.n1235 vdd.n1233 10.6151
R19201 vdd.n1233 vdd.n1232 10.6151
R19202 vdd.n1232 vdd.n1230 10.6151
R19203 vdd.n1230 vdd.n1229 10.6151
R19204 vdd.n1229 vdd.n1226 10.6151
R19205 vdd.n1226 vdd.n1225 10.6151
R19206 vdd.n1225 vdd.n831 10.6151
R19207 vdd.n2221 vdd.n967 10.6151
R19208 vdd.n2216 vdd.n967 10.6151
R19209 vdd.n2216 vdd.n2215 10.6151
R19210 vdd.n2215 vdd.n2214 10.6151
R19211 vdd.n2214 vdd.n2211 10.6151
R19212 vdd.n2211 vdd.n2210 10.6151
R19213 vdd.n2210 vdd.n2207 10.6151
R19214 vdd.n2207 vdd.n2206 10.6151
R19215 vdd.n2206 vdd.n2203 10.6151
R19216 vdd.n2203 vdd.n2202 10.6151
R19217 vdd.n2202 vdd.n2199 10.6151
R19218 vdd.n2199 vdd.n2198 10.6151
R19219 vdd.n2198 vdd.n2195 10.6151
R19220 vdd.n2195 vdd.n2194 10.6151
R19221 vdd.n2194 vdd.n2191 10.6151
R19222 vdd.n2191 vdd.n2190 10.6151
R19223 vdd.n2190 vdd.n2187 10.6151
R19224 vdd.n2187 vdd.n1005 10.6151
R19225 vdd.n1151 vdd.n1005 10.6151
R19226 vdd.n1152 vdd.n1151 10.6151
R19227 vdd.n1155 vdd.n1152 10.6151
R19228 vdd.n1156 vdd.n1155 10.6151
R19229 vdd.n1159 vdd.n1156 10.6151
R19230 vdd.n1160 vdd.n1159 10.6151
R19231 vdd.n1163 vdd.n1160 10.6151
R19232 vdd.n1164 vdd.n1163 10.6151
R19233 vdd.n1167 vdd.n1164 10.6151
R19234 vdd.n1168 vdd.n1167 10.6151
R19235 vdd.n1171 vdd.n1168 10.6151
R19236 vdd.n1172 vdd.n1171 10.6151
R19237 vdd.n1175 vdd.n1172 10.6151
R19238 vdd.n1180 vdd.n1177 10.6151
R19239 vdd.n1181 vdd.n1180 10.6151
R19240 vdd.n2732 vdd.n2731 10.6151
R19241 vdd.n2731 vdd.n2730 10.6151
R19242 vdd.n2730 vdd.n2534 10.6151
R19243 vdd.n2612 vdd.n2534 10.6151
R19244 vdd.n2613 vdd.n2612 10.6151
R19245 vdd.n2615 vdd.n2613 10.6151
R19246 vdd.n2616 vdd.n2615 10.6151
R19247 vdd.n2714 vdd.n2616 10.6151
R19248 vdd.n2714 vdd.n2713 10.6151
R19249 vdd.n2713 vdd.n2712 10.6151
R19250 vdd.n2712 vdd.n2660 10.6151
R19251 vdd.n2660 vdd.n2659 10.6151
R19252 vdd.n2659 vdd.n2657 10.6151
R19253 vdd.n2657 vdd.n2656 10.6151
R19254 vdd.n2656 vdd.n2654 10.6151
R19255 vdd.n2654 vdd.n2653 10.6151
R19256 vdd.n2653 vdd.n2651 10.6151
R19257 vdd.n2651 vdd.n2650 10.6151
R19258 vdd.n2650 vdd.n2648 10.6151
R19259 vdd.n2648 vdd.n2647 10.6151
R19260 vdd.n2647 vdd.n2645 10.6151
R19261 vdd.n2645 vdd.n2644 10.6151
R19262 vdd.n2644 vdd.n2642 10.6151
R19263 vdd.n2642 vdd.n2641 10.6151
R19264 vdd.n2641 vdd.n2639 10.6151
R19265 vdd.n2639 vdd.n2638 10.6151
R19266 vdd.n2638 vdd.n2636 10.6151
R19267 vdd.n2636 vdd.n2635 10.6151
R19268 vdd.n2635 vdd.n2633 10.6151
R19269 vdd.n2633 vdd.n2632 10.6151
R19270 vdd.n2632 vdd.n2630 10.6151
R19271 vdd.n2630 vdd.n2629 10.6151
R19272 vdd.n2629 vdd.n2627 10.6151
R19273 vdd.n2627 vdd.n2626 10.6151
R19274 vdd.n2626 vdd.n2624 10.6151
R19275 vdd.n2624 vdd.n2623 10.6151
R19276 vdd.n2623 vdd.n2621 10.6151
R19277 vdd.n2621 vdd.n2620 10.6151
R19278 vdd.n2620 vdd.n2618 10.6151
R19279 vdd.n2618 vdd.n2617 10.6151
R19280 vdd.n2617 vdd.n664 10.6151
R19281 vdd.n2976 vdd.n664 10.6151
R19282 vdd.n2977 vdd.n2976 10.6151
R19283 vdd.n2803 vdd.n789 10.6151
R19284 vdd.n2798 vdd.n789 10.6151
R19285 vdd.n2798 vdd.n2797 10.6151
R19286 vdd.n2797 vdd.n2796 10.6151
R19287 vdd.n2796 vdd.n2793 10.6151
R19288 vdd.n2793 vdd.n2792 10.6151
R19289 vdd.n2792 vdd.n2789 10.6151
R19290 vdd.n2789 vdd.n2788 10.6151
R19291 vdd.n2788 vdd.n2785 10.6151
R19292 vdd.n2785 vdd.n2784 10.6151
R19293 vdd.n2784 vdd.n2781 10.6151
R19294 vdd.n2781 vdd.n2780 10.6151
R19295 vdd.n2780 vdd.n2777 10.6151
R19296 vdd.n2777 vdd.n2776 10.6151
R19297 vdd.n2776 vdd.n2773 10.6151
R19298 vdd.n2773 vdd.n2772 10.6151
R19299 vdd.n2772 vdd.n2769 10.6151
R19300 vdd.n2769 vdd.n2768 10.6151
R19301 vdd.n2768 vdd.n2765 10.6151
R19302 vdd.n2765 vdd.n2764 10.6151
R19303 vdd.n2764 vdd.n2761 10.6151
R19304 vdd.n2761 vdd.n2760 10.6151
R19305 vdd.n2760 vdd.n2757 10.6151
R19306 vdd.n2757 vdd.n2756 10.6151
R19307 vdd.n2756 vdd.n2753 10.6151
R19308 vdd.n2753 vdd.n2752 10.6151
R19309 vdd.n2752 vdd.n2749 10.6151
R19310 vdd.n2749 vdd.n2748 10.6151
R19311 vdd.n2748 vdd.n2745 10.6151
R19312 vdd.n2745 vdd.n2744 10.6151
R19313 vdd.n2744 vdd.n2741 10.6151
R19314 vdd.n2739 vdd.n2736 10.6151
R19315 vdd.n2736 vdd.n2735 10.6151
R19316 vdd.n2805 vdd.n2804 10.6151
R19317 vdd.n2805 vdd.n778 10.6151
R19318 vdd.n2815 vdd.n778 10.6151
R19319 vdd.n2816 vdd.n2815 10.6151
R19320 vdd.n2817 vdd.n2816 10.6151
R19321 vdd.n2817 vdd.n766 10.6151
R19322 vdd.n2827 vdd.n766 10.6151
R19323 vdd.n2828 vdd.n2827 10.6151
R19324 vdd.n2829 vdd.n2828 10.6151
R19325 vdd.n2829 vdd.n755 10.6151
R19326 vdd.n2839 vdd.n755 10.6151
R19327 vdd.n2840 vdd.n2839 10.6151
R19328 vdd.n2841 vdd.n2840 10.6151
R19329 vdd.n2841 vdd.n744 10.6151
R19330 vdd.n2851 vdd.n744 10.6151
R19331 vdd.n2852 vdd.n2851 10.6151
R19332 vdd.n2853 vdd.n2852 10.6151
R19333 vdd.n2853 vdd.n731 10.6151
R19334 vdd.n2864 vdd.n731 10.6151
R19335 vdd.n2865 vdd.n2864 10.6151
R19336 vdd.n2866 vdd.n2865 10.6151
R19337 vdd.n2866 vdd.n719 10.6151
R19338 vdd.n2876 vdd.n719 10.6151
R19339 vdd.n2877 vdd.n2876 10.6151
R19340 vdd.n2878 vdd.n2877 10.6151
R19341 vdd.n2878 vdd.n707 10.6151
R19342 vdd.n2888 vdd.n707 10.6151
R19343 vdd.n2889 vdd.n2888 10.6151
R19344 vdd.n2890 vdd.n2889 10.6151
R19345 vdd.n2890 vdd.n694 10.6151
R19346 vdd.n2900 vdd.n694 10.6151
R19347 vdd.n2901 vdd.n2900 10.6151
R19348 vdd.n2902 vdd.n2901 10.6151
R19349 vdd.n2902 vdd.n683 10.6151
R19350 vdd.n2912 vdd.n683 10.6151
R19351 vdd.n2913 vdd.n2912 10.6151
R19352 vdd.n2914 vdd.n2913 10.6151
R19353 vdd.n2914 vdd.n669 10.6151
R19354 vdd.n2969 vdd.n669 10.6151
R19355 vdd.n2970 vdd.n2969 10.6151
R19356 vdd.n2971 vdd.n2970 10.6151
R19357 vdd.n2971 vdd.n636 10.6151
R19358 vdd.n3041 vdd.n636 10.6151
R19359 vdd.n3040 vdd.n3039 10.6151
R19360 vdd.n3039 vdd.n637 10.6151
R19361 vdd.n638 vdd.n637 10.6151
R19362 vdd.n3032 vdd.n638 10.6151
R19363 vdd.n3032 vdd.n3031 10.6151
R19364 vdd.n3031 vdd.n3030 10.6151
R19365 vdd.n3030 vdd.n640 10.6151
R19366 vdd.n3025 vdd.n640 10.6151
R19367 vdd.n3025 vdd.n3024 10.6151
R19368 vdd.n3024 vdd.n3023 10.6151
R19369 vdd.n3023 vdd.n643 10.6151
R19370 vdd.n3018 vdd.n643 10.6151
R19371 vdd.n3018 vdd.n3017 10.6151
R19372 vdd.n3017 vdd.n3016 10.6151
R19373 vdd.n3016 vdd.n646 10.6151
R19374 vdd.n3011 vdd.n646 10.6151
R19375 vdd.n3011 vdd.n3010 10.6151
R19376 vdd.n3010 vdd.n3008 10.6151
R19377 vdd.n3008 vdd.n649 10.6151
R19378 vdd.n3003 vdd.n649 10.6151
R19379 vdd.n3003 vdd.n3002 10.6151
R19380 vdd.n3002 vdd.n3001 10.6151
R19381 vdd.n3001 vdd.n652 10.6151
R19382 vdd.n2996 vdd.n652 10.6151
R19383 vdd.n2996 vdd.n2995 10.6151
R19384 vdd.n2995 vdd.n2994 10.6151
R19385 vdd.n2994 vdd.n655 10.6151
R19386 vdd.n2989 vdd.n655 10.6151
R19387 vdd.n2989 vdd.n2988 10.6151
R19388 vdd.n2988 vdd.n2987 10.6151
R19389 vdd.n2987 vdd.n658 10.6151
R19390 vdd.n2982 vdd.n2981 10.6151
R19391 vdd.n2981 vdd.n2980 10.6151
R19392 vdd.n2959 vdd.n2920 10.6151
R19393 vdd.n2954 vdd.n2920 10.6151
R19394 vdd.n2954 vdd.n2953 10.6151
R19395 vdd.n2953 vdd.n2952 10.6151
R19396 vdd.n2952 vdd.n2922 10.6151
R19397 vdd.n2947 vdd.n2922 10.6151
R19398 vdd.n2947 vdd.n2946 10.6151
R19399 vdd.n2946 vdd.n2945 10.6151
R19400 vdd.n2945 vdd.n2925 10.6151
R19401 vdd.n2940 vdd.n2925 10.6151
R19402 vdd.n2940 vdd.n2939 10.6151
R19403 vdd.n2939 vdd.n2938 10.6151
R19404 vdd.n2938 vdd.n2928 10.6151
R19405 vdd.n2933 vdd.n2928 10.6151
R19406 vdd.n2933 vdd.n2932 10.6151
R19407 vdd.n2932 vdd.n610 10.6151
R19408 vdd.n3076 vdd.n610 10.6151
R19409 vdd.n3076 vdd.n611 10.6151
R19410 vdd.n614 vdd.n611 10.6151
R19411 vdd.n3069 vdd.n614 10.6151
R19412 vdd.n3069 vdd.n3068 10.6151
R19413 vdd.n3068 vdd.n3067 10.6151
R19414 vdd.n3067 vdd.n616 10.6151
R19415 vdd.n3062 vdd.n616 10.6151
R19416 vdd.n3062 vdd.n3061 10.6151
R19417 vdd.n3061 vdd.n3060 10.6151
R19418 vdd.n3060 vdd.n619 10.6151
R19419 vdd.n3055 vdd.n619 10.6151
R19420 vdd.n3055 vdd.n3054 10.6151
R19421 vdd.n3054 vdd.n3053 10.6151
R19422 vdd.n3053 vdd.n622 10.6151
R19423 vdd.n3048 vdd.n3047 10.6151
R19424 vdd.n3047 vdd.n3046 10.6151
R19425 vdd.n2609 vdd.n2608 10.6151
R19426 vdd.n2726 vdd.n2609 10.6151
R19427 vdd.n2726 vdd.n2725 10.6151
R19428 vdd.n2725 vdd.n2724 10.6151
R19429 vdd.n2724 vdd.n2722 10.6151
R19430 vdd.n2722 vdd.n2721 10.6151
R19431 vdd.n2721 vdd.n2719 10.6151
R19432 vdd.n2719 vdd.n2718 10.6151
R19433 vdd.n2718 vdd.n2610 10.6151
R19434 vdd.n2708 vdd.n2610 10.6151
R19435 vdd.n2708 vdd.n2707 10.6151
R19436 vdd.n2707 vdd.n2706 10.6151
R19437 vdd.n2706 vdd.n2704 10.6151
R19438 vdd.n2704 vdd.n2703 10.6151
R19439 vdd.n2703 vdd.n2701 10.6151
R19440 vdd.n2701 vdd.n2700 10.6151
R19441 vdd.n2700 vdd.n2698 10.6151
R19442 vdd.n2698 vdd.n2697 10.6151
R19443 vdd.n2697 vdd.n2695 10.6151
R19444 vdd.n2695 vdd.n2694 10.6151
R19445 vdd.n2694 vdd.n2692 10.6151
R19446 vdd.n2692 vdd.n2691 10.6151
R19447 vdd.n2691 vdd.n2689 10.6151
R19448 vdd.n2689 vdd.n2688 10.6151
R19449 vdd.n2688 vdd.n2686 10.6151
R19450 vdd.n2686 vdd.n2685 10.6151
R19451 vdd.n2685 vdd.n2683 10.6151
R19452 vdd.n2683 vdd.n2682 10.6151
R19453 vdd.n2682 vdd.n2680 10.6151
R19454 vdd.n2680 vdd.n2679 10.6151
R19455 vdd.n2679 vdd.n2677 10.6151
R19456 vdd.n2677 vdd.n2676 10.6151
R19457 vdd.n2676 vdd.n2674 10.6151
R19458 vdd.n2674 vdd.n2673 10.6151
R19459 vdd.n2673 vdd.n2671 10.6151
R19460 vdd.n2671 vdd.n2670 10.6151
R19461 vdd.n2670 vdd.n2668 10.6151
R19462 vdd.n2668 vdd.n2667 10.6151
R19463 vdd.n2667 vdd.n2665 10.6151
R19464 vdd.n2665 vdd.n2664 10.6151
R19465 vdd.n2664 vdd.n2662 10.6151
R19466 vdd.n2662 vdd.n2661 10.6151
R19467 vdd.n2661 vdd.n628 10.6151
R19468 vdd.n2540 vdd.n2539 10.6151
R19469 vdd.n2543 vdd.n2540 10.6151
R19470 vdd.n2544 vdd.n2543 10.6151
R19471 vdd.n2547 vdd.n2544 10.6151
R19472 vdd.n2548 vdd.n2547 10.6151
R19473 vdd.n2551 vdd.n2548 10.6151
R19474 vdd.n2552 vdd.n2551 10.6151
R19475 vdd.n2555 vdd.n2552 10.6151
R19476 vdd.n2556 vdd.n2555 10.6151
R19477 vdd.n2559 vdd.n2556 10.6151
R19478 vdd.n2560 vdd.n2559 10.6151
R19479 vdd.n2563 vdd.n2560 10.6151
R19480 vdd.n2564 vdd.n2563 10.6151
R19481 vdd.n2567 vdd.n2564 10.6151
R19482 vdd.n2568 vdd.n2567 10.6151
R19483 vdd.n2571 vdd.n2568 10.6151
R19484 vdd.n2572 vdd.n2571 10.6151
R19485 vdd.n2575 vdd.n2572 10.6151
R19486 vdd.n2576 vdd.n2575 10.6151
R19487 vdd.n2579 vdd.n2576 10.6151
R19488 vdd.n2580 vdd.n2579 10.6151
R19489 vdd.n2583 vdd.n2580 10.6151
R19490 vdd.n2584 vdd.n2583 10.6151
R19491 vdd.n2587 vdd.n2584 10.6151
R19492 vdd.n2588 vdd.n2587 10.6151
R19493 vdd.n2591 vdd.n2588 10.6151
R19494 vdd.n2592 vdd.n2591 10.6151
R19495 vdd.n2595 vdd.n2592 10.6151
R19496 vdd.n2596 vdd.n2595 10.6151
R19497 vdd.n2599 vdd.n2596 10.6151
R19498 vdd.n2600 vdd.n2599 10.6151
R19499 vdd.n2605 vdd.n2603 10.6151
R19500 vdd.n2606 vdd.n2605 10.6151
R19501 vdd.n2809 vdd.n783 10.6151
R19502 vdd.n2810 vdd.n2809 10.6151
R19503 vdd.n2811 vdd.n2810 10.6151
R19504 vdd.n2811 vdd.n772 10.6151
R19505 vdd.n2821 vdd.n772 10.6151
R19506 vdd.n2822 vdd.n2821 10.6151
R19507 vdd.n2823 vdd.n2822 10.6151
R19508 vdd.n2823 vdd.n761 10.6151
R19509 vdd.n2833 vdd.n761 10.6151
R19510 vdd.n2834 vdd.n2833 10.6151
R19511 vdd.n2835 vdd.n2834 10.6151
R19512 vdd.n2835 vdd.n749 10.6151
R19513 vdd.n2845 vdd.n749 10.6151
R19514 vdd.n2846 vdd.n2845 10.6151
R19515 vdd.n2847 vdd.n2846 10.6151
R19516 vdd.n2847 vdd.n738 10.6151
R19517 vdd.n2857 vdd.n738 10.6151
R19518 vdd.n2858 vdd.n2857 10.6151
R19519 vdd.n2860 vdd.n2858 10.6151
R19520 vdd.n2860 vdd.n2859 10.6151
R19521 vdd.n2871 vdd.n2870 10.6151
R19522 vdd.n2872 vdd.n2871 10.6151
R19523 vdd.n2872 vdd.n713 10.6151
R19524 vdd.n2882 vdd.n713 10.6151
R19525 vdd.n2883 vdd.n2882 10.6151
R19526 vdd.n2884 vdd.n2883 10.6151
R19527 vdd.n2884 vdd.n700 10.6151
R19528 vdd.n2894 vdd.n700 10.6151
R19529 vdd.n2895 vdd.n2894 10.6151
R19530 vdd.n2896 vdd.n2895 10.6151
R19531 vdd.n2896 vdd.n688 10.6151
R19532 vdd.n2906 vdd.n688 10.6151
R19533 vdd.n2907 vdd.n2906 10.6151
R19534 vdd.n2908 vdd.n2907 10.6151
R19535 vdd.n2908 vdd.n677 10.6151
R19536 vdd.n2918 vdd.n677 10.6151
R19537 vdd.n2919 vdd.n2918 10.6151
R19538 vdd.n2965 vdd.n2919 10.6151
R19539 vdd.n2965 vdd.n2964 10.6151
R19540 vdd.n2964 vdd.n2963 10.6151
R19541 vdd.n2963 vdd.n2962 10.6151
R19542 vdd.n2962 vdd.n2960 10.6151
R19543 vdd.n2227 vdd.n960 10.6151
R19544 vdd.n2228 vdd.n2227 10.6151
R19545 vdd.n2229 vdd.n2228 10.6151
R19546 vdd.n2229 vdd.n949 10.6151
R19547 vdd.n2239 vdd.n949 10.6151
R19548 vdd.n2240 vdd.n2239 10.6151
R19549 vdd.n2241 vdd.n2240 10.6151
R19550 vdd.n2241 vdd.n936 10.6151
R19551 vdd.n2251 vdd.n936 10.6151
R19552 vdd.n2252 vdd.n2251 10.6151
R19553 vdd.n2253 vdd.n2252 10.6151
R19554 vdd.n2253 vdd.n925 10.6151
R19555 vdd.n2263 vdd.n925 10.6151
R19556 vdd.n2264 vdd.n2263 10.6151
R19557 vdd.n2265 vdd.n2264 10.6151
R19558 vdd.n2265 vdd.n913 10.6151
R19559 vdd.n2275 vdd.n913 10.6151
R19560 vdd.n2276 vdd.n2275 10.6151
R19561 vdd.n2277 vdd.n2276 10.6151
R19562 vdd.n2277 vdd.n900 10.6151
R19563 vdd.n2287 vdd.n900 10.6151
R19564 vdd.n2288 vdd.n2287 10.6151
R19565 vdd.n2290 vdd.n888 10.6151
R19566 vdd.n2300 vdd.n888 10.6151
R19567 vdd.n2301 vdd.n2300 10.6151
R19568 vdd.n2302 vdd.n2301 10.6151
R19569 vdd.n2302 vdd.n876 10.6151
R19570 vdd.n2312 vdd.n876 10.6151
R19571 vdd.n2313 vdd.n2312 10.6151
R19572 vdd.n2314 vdd.n2313 10.6151
R19573 vdd.n2314 vdd.n865 10.6151
R19574 vdd.n2324 vdd.n865 10.6151
R19575 vdd.n2325 vdd.n2324 10.6151
R19576 vdd.n2326 vdd.n2325 10.6151
R19577 vdd.n2326 vdd.n854 10.6151
R19578 vdd.n2336 vdd.n854 10.6151
R19579 vdd.n2337 vdd.n2336 10.6151
R19580 vdd.n2340 vdd.n2337 10.6151
R19581 vdd.n2340 vdd.n2339 10.6151
R19582 vdd.n2339 vdd.n2338 10.6151
R19583 vdd.n2338 vdd.n837 10.6151
R19584 vdd.n2422 vdd.n837 10.6151
R19585 vdd.n2421 vdd.n2420 10.6151
R19586 vdd.n2420 vdd.n2417 10.6151
R19587 vdd.n2417 vdd.n2416 10.6151
R19588 vdd.n2416 vdd.n2413 10.6151
R19589 vdd.n2413 vdd.n2412 10.6151
R19590 vdd.n2412 vdd.n2409 10.6151
R19591 vdd.n2409 vdd.n2408 10.6151
R19592 vdd.n2408 vdd.n2405 10.6151
R19593 vdd.n2405 vdd.n2404 10.6151
R19594 vdd.n2404 vdd.n2401 10.6151
R19595 vdd.n2401 vdd.n2400 10.6151
R19596 vdd.n2400 vdd.n2397 10.6151
R19597 vdd.n2397 vdd.n2396 10.6151
R19598 vdd.n2396 vdd.n2393 10.6151
R19599 vdd.n2393 vdd.n2392 10.6151
R19600 vdd.n2392 vdd.n2389 10.6151
R19601 vdd.n2389 vdd.n2388 10.6151
R19602 vdd.n2388 vdd.n2385 10.6151
R19603 vdd.n2385 vdd.n2384 10.6151
R19604 vdd.n2384 vdd.n2381 10.6151
R19605 vdd.n2381 vdd.n2380 10.6151
R19606 vdd.n2380 vdd.n2377 10.6151
R19607 vdd.n2377 vdd.n2376 10.6151
R19608 vdd.n2376 vdd.n2373 10.6151
R19609 vdd.n2373 vdd.n2372 10.6151
R19610 vdd.n2372 vdd.n2369 10.6151
R19611 vdd.n2369 vdd.n2368 10.6151
R19612 vdd.n2368 vdd.n2365 10.6151
R19613 vdd.n2365 vdd.n2364 10.6151
R19614 vdd.n2364 vdd.n2361 10.6151
R19615 vdd.n2361 vdd.n2360 10.6151
R19616 vdd.n2357 vdd.n2356 10.6151
R19617 vdd.n2356 vdd.n2354 10.6151
R19618 vdd.n1309 vdd.n1307 10.6151
R19619 vdd.n1307 vdd.n1306 10.6151
R19620 vdd.n1306 vdd.n1304 10.6151
R19621 vdd.n1304 vdd.n1303 10.6151
R19622 vdd.n1303 vdd.n1301 10.6151
R19623 vdd.n1301 vdd.n1300 10.6151
R19624 vdd.n1300 vdd.n1298 10.6151
R19625 vdd.n1298 vdd.n1297 10.6151
R19626 vdd.n1297 vdd.n1295 10.6151
R19627 vdd.n1295 vdd.n1294 10.6151
R19628 vdd.n1294 vdd.n1292 10.6151
R19629 vdd.n1292 vdd.n1291 10.6151
R19630 vdd.n1291 vdd.n1289 10.6151
R19631 vdd.n1289 vdd.n1288 10.6151
R19632 vdd.n1288 vdd.n1286 10.6151
R19633 vdd.n1286 vdd.n1285 10.6151
R19634 vdd.n1285 vdd.n1283 10.6151
R19635 vdd.n1283 vdd.n1282 10.6151
R19636 vdd.n1282 vdd.n1280 10.6151
R19637 vdd.n1280 vdd.n1279 10.6151
R19638 vdd.n1279 vdd.n1277 10.6151
R19639 vdd.n1277 vdd.n1276 10.6151
R19640 vdd.n1276 vdd.n1274 10.6151
R19641 vdd.n1274 vdd.n1273 10.6151
R19642 vdd.n1273 vdd.n1271 10.6151
R19643 vdd.n1271 vdd.n1270 10.6151
R19644 vdd.n1270 vdd.n1268 10.6151
R19645 vdd.n1268 vdd.n1267 10.6151
R19646 vdd.n1267 vdd.n1146 10.6151
R19647 vdd.n1238 vdd.n1146 10.6151
R19648 vdd.n1239 vdd.n1238 10.6151
R19649 vdd.n1241 vdd.n1239 10.6151
R19650 vdd.n1242 vdd.n1241 10.6151
R19651 vdd.n1251 vdd.n1242 10.6151
R19652 vdd.n1251 vdd.n1250 10.6151
R19653 vdd.n1250 vdd.n1249 10.6151
R19654 vdd.n1249 vdd.n1247 10.6151
R19655 vdd.n1247 vdd.n1246 10.6151
R19656 vdd.n1246 vdd.n1244 10.6151
R19657 vdd.n1244 vdd.n1243 10.6151
R19658 vdd.n1243 vdd.n841 10.6151
R19659 vdd.n2352 vdd.n841 10.6151
R19660 vdd.n2353 vdd.n2352 10.6151
R19661 vdd.n1110 vdd.n1109 10.6151
R19662 vdd.n1113 vdd.n1110 10.6151
R19663 vdd.n1114 vdd.n1113 10.6151
R19664 vdd.n1117 vdd.n1114 10.6151
R19665 vdd.n1118 vdd.n1117 10.6151
R19666 vdd.n1121 vdd.n1118 10.6151
R19667 vdd.n1122 vdd.n1121 10.6151
R19668 vdd.n1125 vdd.n1122 10.6151
R19669 vdd.n1126 vdd.n1125 10.6151
R19670 vdd.n1129 vdd.n1126 10.6151
R19671 vdd.n1130 vdd.n1129 10.6151
R19672 vdd.n1133 vdd.n1130 10.6151
R19673 vdd.n1134 vdd.n1133 10.6151
R19674 vdd.n1137 vdd.n1134 10.6151
R19675 vdd.n1138 vdd.n1137 10.6151
R19676 vdd.n1141 vdd.n1138 10.6151
R19677 vdd.n1343 vdd.n1141 10.6151
R19678 vdd.n1343 vdd.n1342 10.6151
R19679 vdd.n1342 vdd.n1340 10.6151
R19680 vdd.n1340 vdd.n1337 10.6151
R19681 vdd.n1337 vdd.n1336 10.6151
R19682 vdd.n1336 vdd.n1333 10.6151
R19683 vdd.n1333 vdd.n1332 10.6151
R19684 vdd.n1332 vdd.n1329 10.6151
R19685 vdd.n1329 vdd.n1328 10.6151
R19686 vdd.n1328 vdd.n1325 10.6151
R19687 vdd.n1325 vdd.n1324 10.6151
R19688 vdd.n1324 vdd.n1321 10.6151
R19689 vdd.n1321 vdd.n1320 10.6151
R19690 vdd.n1320 vdd.n1317 10.6151
R19691 vdd.n1317 vdd.n1316 10.6151
R19692 vdd.n1313 vdd.n1312 10.6151
R19693 vdd.n1312 vdd.n1310 10.6151
R19694 vdd.n1727 vdd.t87 10.5435
R19695 vdd.n2070 vdd.t169 10.5435
R19696 vdd.n3212 vdd.t179 10.5435
R19697 vdd.n3436 vdd.t70 10.5435
R19698 vdd.n292 vdd.n274 10.4732
R19699 vdd.n241 vdd.n223 10.4732
R19700 vdd.n198 vdd.n180 10.4732
R19701 vdd.n147 vdd.n129 10.4732
R19702 vdd.n105 vdd.n87 10.4732
R19703 vdd.n54 vdd.n36 10.4732
R19704 vdd.n1942 vdd.n1924 10.4732
R19705 vdd.n1993 vdd.n1975 10.4732
R19706 vdd.n1848 vdd.n1830 10.4732
R19707 vdd.n1899 vdd.n1881 10.4732
R19708 vdd.n1755 vdd.n1737 10.4732
R19709 vdd.n1806 vdd.n1788 10.4732
R19710 vdd.n2025 vdd.t121 10.3167
R19711 vdd.t74 vdd.n493 10.3167
R19712 vdd.n2187 vdd.n2186 9.98956
R19713 vdd.n3010 vdd.n3009 9.98956
R19714 vdd.n3077 vdd.n3076 9.98956
R19715 vdd.n2079 vdd.n1343 9.98956
R19716 vdd.n1678 vdd.t197 9.86327
R19717 vdd.n3412 vdd.t183 9.86327
R19718 vdd.n2424 vdd.t49 9.7499
R19719 vdd.t34 vdd.n785 9.7499
R19720 vdd.n291 vdd.n276 9.69747
R19721 vdd.n240 vdd.n225 9.69747
R19722 vdd.n197 vdd.n182 9.69747
R19723 vdd.n146 vdd.n131 9.69747
R19724 vdd.n104 vdd.n89 9.69747
R19725 vdd.n53 vdd.n38 9.69747
R19726 vdd.n1941 vdd.n1926 9.69747
R19727 vdd.n1992 vdd.n1977 9.69747
R19728 vdd.n1847 vdd.n1832 9.69747
R19729 vdd.n1898 vdd.n1883 9.69747
R19730 vdd.n1754 vdd.n1739 9.69747
R19731 vdd.n1805 vdd.n1790 9.69747
R19732 vdd.n307 vdd.n306 9.45567
R19733 vdd.n256 vdd.n255 9.45567
R19734 vdd.n213 vdd.n212 9.45567
R19735 vdd.n162 vdd.n161 9.45567
R19736 vdd.n120 vdd.n119 9.45567
R19737 vdd.n69 vdd.n68 9.45567
R19738 vdd.n1957 vdd.n1956 9.45567
R19739 vdd.n2008 vdd.n2007 9.45567
R19740 vdd.n1863 vdd.n1862 9.45567
R19741 vdd.n1914 vdd.n1913 9.45567
R19742 vdd.n1770 vdd.n1769 9.45567
R19743 vdd.n1821 vdd.n1820 9.45567
R19744 vdd.n2149 vdd.n1035 9.3005
R19745 vdd.n2148 vdd.n2147 9.3005
R19746 vdd.n1041 vdd.n1040 9.3005
R19747 vdd.n2142 vdd.n1045 9.3005
R19748 vdd.n2141 vdd.n1046 9.3005
R19749 vdd.n2140 vdd.n1047 9.3005
R19750 vdd.n1051 vdd.n1048 9.3005
R19751 vdd.n2135 vdd.n1052 9.3005
R19752 vdd.n2134 vdd.n1053 9.3005
R19753 vdd.n2133 vdd.n1054 9.3005
R19754 vdd.n1058 vdd.n1055 9.3005
R19755 vdd.n2128 vdd.n1059 9.3005
R19756 vdd.n2127 vdd.n1060 9.3005
R19757 vdd.n2126 vdd.n1061 9.3005
R19758 vdd.n1065 vdd.n1062 9.3005
R19759 vdd.n2121 vdd.n1066 9.3005
R19760 vdd.n2120 vdd.n1067 9.3005
R19761 vdd.n2119 vdd.n1068 9.3005
R19762 vdd.n1072 vdd.n1069 9.3005
R19763 vdd.n2114 vdd.n1073 9.3005
R19764 vdd.n2113 vdd.n1074 9.3005
R19765 vdd.n2112 vdd.n2111 9.3005
R19766 vdd.n2110 vdd.n1075 9.3005
R19767 vdd.n2109 vdd.n2108 9.3005
R19768 vdd.n1081 vdd.n1080 9.3005
R19769 vdd.n2103 vdd.n1085 9.3005
R19770 vdd.n2102 vdd.n1086 9.3005
R19771 vdd.n2101 vdd.n1087 9.3005
R19772 vdd.n1091 vdd.n1088 9.3005
R19773 vdd.n2096 vdd.n1092 9.3005
R19774 vdd.n2095 vdd.n1093 9.3005
R19775 vdd.n2094 vdd.n1094 9.3005
R19776 vdd.n1098 vdd.n1095 9.3005
R19777 vdd.n2089 vdd.n1099 9.3005
R19778 vdd.n2088 vdd.n1100 9.3005
R19779 vdd.n2087 vdd.n1101 9.3005
R19780 vdd.n1105 vdd.n1102 9.3005
R19781 vdd.n2082 vdd.n1106 9.3005
R19782 vdd.n2151 vdd.n2150 9.3005
R19783 vdd.n2173 vdd.n1006 9.3005
R19784 vdd.n2172 vdd.n1014 9.3005
R19785 vdd.n1018 vdd.n1015 9.3005
R19786 vdd.n2167 vdd.n1019 9.3005
R19787 vdd.n2166 vdd.n1020 9.3005
R19788 vdd.n2165 vdd.n1021 9.3005
R19789 vdd.n1025 vdd.n1022 9.3005
R19790 vdd.n2160 vdd.n1026 9.3005
R19791 vdd.n2159 vdd.n1027 9.3005
R19792 vdd.n2158 vdd.n1028 9.3005
R19793 vdd.n1032 vdd.n1029 9.3005
R19794 vdd.n2153 vdd.n1033 9.3005
R19795 vdd.n2152 vdd.n1034 9.3005
R19796 vdd.n2185 vdd.n2184 9.3005
R19797 vdd.n1010 vdd.n1009 9.3005
R19798 vdd.n2013 vdd.n1394 9.3005
R19799 vdd.n2015 vdd.n2014 9.3005
R19800 vdd.n1384 vdd.n1383 9.3005
R19801 vdd.n2029 vdd.n2028 9.3005
R19802 vdd.n2030 vdd.n1382 9.3005
R19803 vdd.n2032 vdd.n2031 9.3005
R19804 vdd.n1373 vdd.n1372 9.3005
R19805 vdd.n2046 vdd.n2045 9.3005
R19806 vdd.n2047 vdd.n1371 9.3005
R19807 vdd.n2049 vdd.n2048 9.3005
R19808 vdd.n1361 vdd.n1360 9.3005
R19809 vdd.n2065 vdd.n2064 9.3005
R19810 vdd.n2066 vdd.n1359 9.3005
R19811 vdd.n2068 vdd.n2067 9.3005
R19812 vdd.n283 vdd.n282 9.3005
R19813 vdd.n278 vdd.n277 9.3005
R19814 vdd.n289 vdd.n288 9.3005
R19815 vdd.n291 vdd.n290 9.3005
R19816 vdd.n274 vdd.n273 9.3005
R19817 vdd.n297 vdd.n296 9.3005
R19818 vdd.n299 vdd.n298 9.3005
R19819 vdd.n271 vdd.n268 9.3005
R19820 vdd.n306 vdd.n305 9.3005
R19821 vdd.n232 vdd.n231 9.3005
R19822 vdd.n227 vdd.n226 9.3005
R19823 vdd.n238 vdd.n237 9.3005
R19824 vdd.n240 vdd.n239 9.3005
R19825 vdd.n223 vdd.n222 9.3005
R19826 vdd.n246 vdd.n245 9.3005
R19827 vdd.n248 vdd.n247 9.3005
R19828 vdd.n220 vdd.n217 9.3005
R19829 vdd.n255 vdd.n254 9.3005
R19830 vdd.n189 vdd.n188 9.3005
R19831 vdd.n184 vdd.n183 9.3005
R19832 vdd.n195 vdd.n194 9.3005
R19833 vdd.n197 vdd.n196 9.3005
R19834 vdd.n180 vdd.n179 9.3005
R19835 vdd.n203 vdd.n202 9.3005
R19836 vdd.n205 vdd.n204 9.3005
R19837 vdd.n177 vdd.n174 9.3005
R19838 vdd.n212 vdd.n211 9.3005
R19839 vdd.n138 vdd.n137 9.3005
R19840 vdd.n133 vdd.n132 9.3005
R19841 vdd.n144 vdd.n143 9.3005
R19842 vdd.n146 vdd.n145 9.3005
R19843 vdd.n129 vdd.n128 9.3005
R19844 vdd.n152 vdd.n151 9.3005
R19845 vdd.n154 vdd.n153 9.3005
R19846 vdd.n126 vdd.n123 9.3005
R19847 vdd.n161 vdd.n160 9.3005
R19848 vdd.n96 vdd.n95 9.3005
R19849 vdd.n91 vdd.n90 9.3005
R19850 vdd.n102 vdd.n101 9.3005
R19851 vdd.n104 vdd.n103 9.3005
R19852 vdd.n87 vdd.n86 9.3005
R19853 vdd.n110 vdd.n109 9.3005
R19854 vdd.n112 vdd.n111 9.3005
R19855 vdd.n84 vdd.n81 9.3005
R19856 vdd.n119 vdd.n118 9.3005
R19857 vdd.n45 vdd.n44 9.3005
R19858 vdd.n40 vdd.n39 9.3005
R19859 vdd.n51 vdd.n50 9.3005
R19860 vdd.n53 vdd.n52 9.3005
R19861 vdd.n36 vdd.n35 9.3005
R19862 vdd.n59 vdd.n58 9.3005
R19863 vdd.n61 vdd.n60 9.3005
R19864 vdd.n33 vdd.n30 9.3005
R19865 vdd.n68 vdd.n67 9.3005
R19866 vdd.n3126 vdd.n3125 9.3005
R19867 vdd.n3127 vdd.n578 9.3005
R19868 vdd.n577 vdd.n575 9.3005
R19869 vdd.n3133 vdd.n574 9.3005
R19870 vdd.n3134 vdd.n573 9.3005
R19871 vdd.n3135 vdd.n572 9.3005
R19872 vdd.n571 vdd.n569 9.3005
R19873 vdd.n3141 vdd.n568 9.3005
R19874 vdd.n3142 vdd.n567 9.3005
R19875 vdd.n3143 vdd.n566 9.3005
R19876 vdd.n565 vdd.n563 9.3005
R19877 vdd.n3149 vdd.n562 9.3005
R19878 vdd.n3150 vdd.n561 9.3005
R19879 vdd.n3151 vdd.n560 9.3005
R19880 vdd.n559 vdd.n557 9.3005
R19881 vdd.n3157 vdd.n556 9.3005
R19882 vdd.n3158 vdd.n555 9.3005
R19883 vdd.n3159 vdd.n554 9.3005
R19884 vdd.n553 vdd.n551 9.3005
R19885 vdd.n3165 vdd.n550 9.3005
R19886 vdd.n3166 vdd.n549 9.3005
R19887 vdd.n3167 vdd.n548 9.3005
R19888 vdd.n547 vdd.n545 9.3005
R19889 vdd.n3173 vdd.n542 9.3005
R19890 vdd.n3174 vdd.n541 9.3005
R19891 vdd.n3175 vdd.n540 9.3005
R19892 vdd.n539 vdd.n537 9.3005
R19893 vdd.n3181 vdd.n536 9.3005
R19894 vdd.n3182 vdd.n535 9.3005
R19895 vdd.n3183 vdd.n534 9.3005
R19896 vdd.n533 vdd.n531 9.3005
R19897 vdd.n3189 vdd.n530 9.3005
R19898 vdd.n3190 vdd.n529 9.3005
R19899 vdd.n3191 vdd.n528 9.3005
R19900 vdd.n527 vdd.n525 9.3005
R19901 vdd.n3196 vdd.n524 9.3005
R19902 vdd.n3206 vdd.n518 9.3005
R19903 vdd.n3208 vdd.n3207 9.3005
R19904 vdd.n509 vdd.n508 9.3005
R19905 vdd.n3223 vdd.n3222 9.3005
R19906 vdd.n3224 vdd.n507 9.3005
R19907 vdd.n3226 vdd.n3225 9.3005
R19908 vdd.n497 vdd.n496 9.3005
R19909 vdd.n3239 vdd.n3238 9.3005
R19910 vdd.n3240 vdd.n495 9.3005
R19911 vdd.n3242 vdd.n3241 9.3005
R19912 vdd.n485 vdd.n484 9.3005
R19913 vdd.n3256 vdd.n3255 9.3005
R19914 vdd.n3257 vdd.n483 9.3005
R19915 vdd.n3259 vdd.n3258 9.3005
R19916 vdd.n312 vdd.n310 9.3005
R19917 vdd.n3210 vdd.n3209 9.3005
R19918 vdd.n3439 vdd.n3438 9.3005
R19919 vdd.n313 vdd.n311 9.3005
R19920 vdd.n3432 vdd.n320 9.3005
R19921 vdd.n3431 vdd.n321 9.3005
R19922 vdd.n3430 vdd.n322 9.3005
R19923 vdd.n331 vdd.n323 9.3005
R19924 vdd.n3424 vdd.n332 9.3005
R19925 vdd.n3423 vdd.n333 9.3005
R19926 vdd.n3422 vdd.n334 9.3005
R19927 vdd.n342 vdd.n335 9.3005
R19928 vdd.n3416 vdd.n343 9.3005
R19929 vdd.n3415 vdd.n344 9.3005
R19930 vdd.n3414 vdd.n345 9.3005
R19931 vdd.n353 vdd.n346 9.3005
R19932 vdd.n3408 vdd.n3407 9.3005
R19933 vdd.n3404 vdd.n354 9.3005
R19934 vdd.n3403 vdd.n357 9.3005
R19935 vdd.n361 vdd.n358 9.3005
R19936 vdd.n362 vdd.n359 9.3005
R19937 vdd.n3396 vdd.n363 9.3005
R19938 vdd.n3395 vdd.n364 9.3005
R19939 vdd.n3394 vdd.n365 9.3005
R19940 vdd.n369 vdd.n366 9.3005
R19941 vdd.n3389 vdd.n370 9.3005
R19942 vdd.n3388 vdd.n371 9.3005
R19943 vdd.n3387 vdd.n372 9.3005
R19944 vdd.n376 vdd.n373 9.3005
R19945 vdd.n3382 vdd.n377 9.3005
R19946 vdd.n3381 vdd.n378 9.3005
R19947 vdd.n3380 vdd.n379 9.3005
R19948 vdd.n383 vdd.n380 9.3005
R19949 vdd.n3375 vdd.n384 9.3005
R19950 vdd.n3374 vdd.n385 9.3005
R19951 vdd.n3373 vdd.n3372 9.3005
R19952 vdd.n3371 vdd.n386 9.3005
R19953 vdd.n3370 vdd.n3369 9.3005
R19954 vdd.n392 vdd.n391 9.3005
R19955 vdd.n3364 vdd.n396 9.3005
R19956 vdd.n3363 vdd.n397 9.3005
R19957 vdd.n3362 vdd.n398 9.3005
R19958 vdd.n402 vdd.n399 9.3005
R19959 vdd.n3357 vdd.n403 9.3005
R19960 vdd.n3356 vdd.n404 9.3005
R19961 vdd.n3355 vdd.n405 9.3005
R19962 vdd.n409 vdd.n406 9.3005
R19963 vdd.n3350 vdd.n410 9.3005
R19964 vdd.n3349 vdd.n411 9.3005
R19965 vdd.n3348 vdd.n412 9.3005
R19966 vdd.n416 vdd.n413 9.3005
R19967 vdd.n3343 vdd.n417 9.3005
R19968 vdd.n3342 vdd.n418 9.3005
R19969 vdd.n3341 vdd.n419 9.3005
R19970 vdd.n423 vdd.n420 9.3005
R19971 vdd.n3336 vdd.n424 9.3005
R19972 vdd.n3335 vdd.n425 9.3005
R19973 vdd.n3334 vdd.n3333 9.3005
R19974 vdd.n3332 vdd.n426 9.3005
R19975 vdd.n3331 vdd.n3330 9.3005
R19976 vdd.n432 vdd.n431 9.3005
R19977 vdd.n3325 vdd.n436 9.3005
R19978 vdd.n3324 vdd.n437 9.3005
R19979 vdd.n3323 vdd.n438 9.3005
R19980 vdd.n442 vdd.n439 9.3005
R19981 vdd.n3318 vdd.n443 9.3005
R19982 vdd.n3317 vdd.n444 9.3005
R19983 vdd.n3316 vdd.n445 9.3005
R19984 vdd.n449 vdd.n446 9.3005
R19985 vdd.n3311 vdd.n450 9.3005
R19986 vdd.n3310 vdd.n451 9.3005
R19987 vdd.n3309 vdd.n452 9.3005
R19988 vdd.n456 vdd.n453 9.3005
R19989 vdd.n3304 vdd.n457 9.3005
R19990 vdd.n3303 vdd.n458 9.3005
R19991 vdd.n3302 vdd.n459 9.3005
R19992 vdd.n463 vdd.n460 9.3005
R19993 vdd.n3297 vdd.n464 9.3005
R19994 vdd.n3296 vdd.n465 9.3005
R19995 vdd.n3292 vdd.n3289 9.3005
R19996 vdd.n3406 vdd.n3405 9.3005
R19997 vdd.n3216 vdd.n513 9.3005
R19998 vdd.n3218 vdd.n3217 9.3005
R19999 vdd.n503 vdd.n502 9.3005
R20000 vdd.n3231 vdd.n3230 9.3005
R20001 vdd.n3232 vdd.n501 9.3005
R20002 vdd.n3234 vdd.n3233 9.3005
R20003 vdd.n490 vdd.n489 9.3005
R20004 vdd.n3247 vdd.n3246 9.3005
R20005 vdd.n3248 vdd.n488 9.3005
R20006 vdd.n3250 vdd.n3249 9.3005
R20007 vdd.n478 vdd.n477 9.3005
R20008 vdd.n3264 vdd.n3263 9.3005
R20009 vdd.n3265 vdd.n476 9.3005
R20010 vdd.n3267 vdd.n3266 9.3005
R20011 vdd.n3268 vdd.n475 9.3005
R20012 vdd.n3270 vdd.n3269 9.3005
R20013 vdd.n3271 vdd.n474 9.3005
R20014 vdd.n3273 vdd.n3272 9.3005
R20015 vdd.n3274 vdd.n472 9.3005
R20016 vdd.n3276 vdd.n3275 9.3005
R20017 vdd.n3277 vdd.n471 9.3005
R20018 vdd.n3279 vdd.n3278 9.3005
R20019 vdd.n3280 vdd.n469 9.3005
R20020 vdd.n3282 vdd.n3281 9.3005
R20021 vdd.n3283 vdd.n468 9.3005
R20022 vdd.n3285 vdd.n3284 9.3005
R20023 vdd.n3286 vdd.n466 9.3005
R20024 vdd.n3288 vdd.n3287 9.3005
R20025 vdd.n3215 vdd.n3214 9.3005
R20026 vdd.n3079 vdd.n514 9.3005
R20027 vdd.n3084 vdd.n3078 9.3005
R20028 vdd.n3094 vdd.n605 9.3005
R20029 vdd.n3095 vdd.n604 9.3005
R20030 vdd.n603 vdd.n601 9.3005
R20031 vdd.n3101 vdd.n600 9.3005
R20032 vdd.n3102 vdd.n599 9.3005
R20033 vdd.n3103 vdd.n598 9.3005
R20034 vdd.n597 vdd.n595 9.3005
R20035 vdd.n3109 vdd.n594 9.3005
R20036 vdd.n3110 vdd.n593 9.3005
R20037 vdd.n3111 vdd.n592 9.3005
R20038 vdd.n591 vdd.n589 9.3005
R20039 vdd.n3116 vdd.n588 9.3005
R20040 vdd.n3117 vdd.n587 9.3005
R20041 vdd.n583 vdd.n582 9.3005
R20042 vdd.n3123 vdd.n3122 9.3005
R20043 vdd.n3124 vdd.n579 9.3005
R20044 vdd.n2078 vdd.n2077 9.3005
R20045 vdd.n2073 vdd.n1345 9.3005
R20046 vdd.n1674 vdd.n1434 9.3005
R20047 vdd.n1676 vdd.n1675 9.3005
R20048 vdd.n1425 vdd.n1424 9.3005
R20049 vdd.n1689 vdd.n1688 9.3005
R20050 vdd.n1690 vdd.n1423 9.3005
R20051 vdd.n1692 vdd.n1691 9.3005
R20052 vdd.n1412 vdd.n1411 9.3005
R20053 vdd.n1705 vdd.n1704 9.3005
R20054 vdd.n1706 vdd.n1410 9.3005
R20055 vdd.n1708 vdd.n1707 9.3005
R20056 vdd.n1401 vdd.n1400 9.3005
R20057 vdd.n1722 vdd.n1721 9.3005
R20058 vdd.n1723 vdd.n1399 9.3005
R20059 vdd.n1725 vdd.n1724 9.3005
R20060 vdd.n1390 vdd.n1389 9.3005
R20061 vdd.n2020 vdd.n2019 9.3005
R20062 vdd.n2021 vdd.n1388 9.3005
R20063 vdd.n2023 vdd.n2022 9.3005
R20064 vdd.n1378 vdd.n1377 9.3005
R20065 vdd.n2037 vdd.n2036 9.3005
R20066 vdd.n2038 vdd.n1376 9.3005
R20067 vdd.n2040 vdd.n2039 9.3005
R20068 vdd.n1368 vdd.n1367 9.3005
R20069 vdd.n2054 vdd.n2053 9.3005
R20070 vdd.n2055 vdd.n1365 9.3005
R20071 vdd.n2059 vdd.n2058 9.3005
R20072 vdd.n2057 vdd.n1366 9.3005
R20073 vdd.n2056 vdd.n1356 9.3005
R20074 vdd.n1673 vdd.n1672 9.3005
R20075 vdd.n1568 vdd.n1558 9.3005
R20076 vdd.n1570 vdd.n1569 9.3005
R20077 vdd.n1571 vdd.n1557 9.3005
R20078 vdd.n1573 vdd.n1572 9.3005
R20079 vdd.n1574 vdd.n1550 9.3005
R20080 vdd.n1576 vdd.n1575 9.3005
R20081 vdd.n1577 vdd.n1549 9.3005
R20082 vdd.n1579 vdd.n1578 9.3005
R20083 vdd.n1580 vdd.n1542 9.3005
R20084 vdd.n1582 vdd.n1581 9.3005
R20085 vdd.n1583 vdd.n1541 9.3005
R20086 vdd.n1585 vdd.n1584 9.3005
R20087 vdd.n1586 vdd.n1534 9.3005
R20088 vdd.n1588 vdd.n1587 9.3005
R20089 vdd.n1589 vdd.n1533 9.3005
R20090 vdd.n1591 vdd.n1590 9.3005
R20091 vdd.n1592 vdd.n1527 9.3005
R20092 vdd.n1594 vdd.n1593 9.3005
R20093 vdd.n1595 vdd.n1525 9.3005
R20094 vdd.n1597 vdd.n1596 9.3005
R20095 vdd.n1526 vdd.n1523 9.3005
R20096 vdd.n1604 vdd.n1519 9.3005
R20097 vdd.n1606 vdd.n1605 9.3005
R20098 vdd.n1607 vdd.n1518 9.3005
R20099 vdd.n1609 vdd.n1608 9.3005
R20100 vdd.n1610 vdd.n1511 9.3005
R20101 vdd.n1612 vdd.n1611 9.3005
R20102 vdd.n1613 vdd.n1510 9.3005
R20103 vdd.n1615 vdd.n1614 9.3005
R20104 vdd.n1616 vdd.n1503 9.3005
R20105 vdd.n1618 vdd.n1617 9.3005
R20106 vdd.n1619 vdd.n1502 9.3005
R20107 vdd.n1621 vdd.n1620 9.3005
R20108 vdd.n1622 vdd.n1495 9.3005
R20109 vdd.n1624 vdd.n1623 9.3005
R20110 vdd.n1625 vdd.n1494 9.3005
R20111 vdd.n1627 vdd.n1626 9.3005
R20112 vdd.n1628 vdd.n1487 9.3005
R20113 vdd.n1630 vdd.n1629 9.3005
R20114 vdd.n1631 vdd.n1486 9.3005
R20115 vdd.n1633 vdd.n1632 9.3005
R20116 vdd.n1634 vdd.n1479 9.3005
R20117 vdd.n1636 vdd.n1635 9.3005
R20118 vdd.n1637 vdd.n1478 9.3005
R20119 vdd.n1639 vdd.n1638 9.3005
R20120 vdd.n1640 vdd.n1469 9.3005
R20121 vdd.n1642 vdd.n1641 9.3005
R20122 vdd.n1643 vdd.n1468 9.3005
R20123 vdd.n1645 vdd.n1644 9.3005
R20124 vdd.n1646 vdd.n1461 9.3005
R20125 vdd.n1648 vdd.n1647 9.3005
R20126 vdd.n1649 vdd.n1460 9.3005
R20127 vdd.n1651 vdd.n1650 9.3005
R20128 vdd.n1652 vdd.n1453 9.3005
R20129 vdd.n1654 vdd.n1653 9.3005
R20130 vdd.n1655 vdd.n1452 9.3005
R20131 vdd.n1657 vdd.n1656 9.3005
R20132 vdd.n1658 vdd.n1445 9.3005
R20133 vdd.n1660 vdd.n1659 9.3005
R20134 vdd.n1661 vdd.n1444 9.3005
R20135 vdd.n1663 vdd.n1662 9.3005
R20136 vdd.n1664 vdd.n1440 9.3005
R20137 vdd.n1666 vdd.n1665 9.3005
R20138 vdd.n1564 vdd.n1435 9.3005
R20139 vdd.n1431 vdd.n1430 9.3005
R20140 vdd.n1681 vdd.n1680 9.3005
R20141 vdd.n1682 vdd.n1429 9.3005
R20142 vdd.n1684 vdd.n1683 9.3005
R20143 vdd.n1419 vdd.n1418 9.3005
R20144 vdd.n1697 vdd.n1696 9.3005
R20145 vdd.n1698 vdd.n1417 9.3005
R20146 vdd.n1700 vdd.n1699 9.3005
R20147 vdd.n1407 vdd.n1406 9.3005
R20148 vdd.n1714 vdd.n1713 9.3005
R20149 vdd.n1715 vdd.n1405 9.3005
R20150 vdd.n1717 vdd.n1716 9.3005
R20151 vdd.n1396 vdd.n1395 9.3005
R20152 vdd.n1668 vdd.n1667 9.3005
R20153 vdd.n2012 vdd.n1729 9.3005
R20154 vdd.n1933 vdd.n1932 9.3005
R20155 vdd.n1928 vdd.n1927 9.3005
R20156 vdd.n1939 vdd.n1938 9.3005
R20157 vdd.n1941 vdd.n1940 9.3005
R20158 vdd.n1924 vdd.n1923 9.3005
R20159 vdd.n1947 vdd.n1946 9.3005
R20160 vdd.n1949 vdd.n1948 9.3005
R20161 vdd.n1921 vdd.n1918 9.3005
R20162 vdd.n1956 vdd.n1955 9.3005
R20163 vdd.n1984 vdd.n1983 9.3005
R20164 vdd.n1979 vdd.n1978 9.3005
R20165 vdd.n1990 vdd.n1989 9.3005
R20166 vdd.n1992 vdd.n1991 9.3005
R20167 vdd.n1975 vdd.n1974 9.3005
R20168 vdd.n1998 vdd.n1997 9.3005
R20169 vdd.n2000 vdd.n1999 9.3005
R20170 vdd.n1972 vdd.n1969 9.3005
R20171 vdd.n2007 vdd.n2006 9.3005
R20172 vdd.n1839 vdd.n1838 9.3005
R20173 vdd.n1834 vdd.n1833 9.3005
R20174 vdd.n1845 vdd.n1844 9.3005
R20175 vdd.n1847 vdd.n1846 9.3005
R20176 vdd.n1830 vdd.n1829 9.3005
R20177 vdd.n1853 vdd.n1852 9.3005
R20178 vdd.n1855 vdd.n1854 9.3005
R20179 vdd.n1827 vdd.n1824 9.3005
R20180 vdd.n1862 vdd.n1861 9.3005
R20181 vdd.n1890 vdd.n1889 9.3005
R20182 vdd.n1885 vdd.n1884 9.3005
R20183 vdd.n1896 vdd.n1895 9.3005
R20184 vdd.n1898 vdd.n1897 9.3005
R20185 vdd.n1881 vdd.n1880 9.3005
R20186 vdd.n1904 vdd.n1903 9.3005
R20187 vdd.n1906 vdd.n1905 9.3005
R20188 vdd.n1878 vdd.n1875 9.3005
R20189 vdd.n1913 vdd.n1912 9.3005
R20190 vdd.n1746 vdd.n1745 9.3005
R20191 vdd.n1741 vdd.n1740 9.3005
R20192 vdd.n1752 vdd.n1751 9.3005
R20193 vdd.n1754 vdd.n1753 9.3005
R20194 vdd.n1737 vdd.n1736 9.3005
R20195 vdd.n1760 vdd.n1759 9.3005
R20196 vdd.n1762 vdd.n1761 9.3005
R20197 vdd.n1734 vdd.n1731 9.3005
R20198 vdd.n1769 vdd.n1768 9.3005
R20199 vdd.n1797 vdd.n1796 9.3005
R20200 vdd.n1792 vdd.n1791 9.3005
R20201 vdd.n1803 vdd.n1802 9.3005
R20202 vdd.n1805 vdd.n1804 9.3005
R20203 vdd.n1788 vdd.n1787 9.3005
R20204 vdd.n1811 vdd.n1810 9.3005
R20205 vdd.n1813 vdd.n1812 9.3005
R20206 vdd.n1785 vdd.n1782 9.3005
R20207 vdd.n1820 vdd.n1819 9.3005
R20208 vdd.n288 vdd.n287 8.92171
R20209 vdd.n237 vdd.n236 8.92171
R20210 vdd.n194 vdd.n193 8.92171
R20211 vdd.n143 vdd.n142 8.92171
R20212 vdd.n101 vdd.n100 8.92171
R20213 vdd.n50 vdd.n49 8.92171
R20214 vdd.n1938 vdd.n1937 8.92171
R20215 vdd.n1989 vdd.n1988 8.92171
R20216 vdd.n1844 vdd.n1843 8.92171
R20217 vdd.n1895 vdd.n1894 8.92171
R20218 vdd.n1751 vdd.n1750 8.92171
R20219 vdd.n1802 vdd.n1801 8.92171
R20220 vdd.n215 vdd.n121 8.81535
R20221 vdd.n1916 vdd.n1822 8.81535
R20222 vdd.n2051 vdd.t89 8.72962
R20223 vdd.n3228 vdd.t112 8.72962
R20224 vdd.t68 vdd.n2025 8.50289
R20225 vdd.n493 vdd.t77 8.50289
R20226 vdd.n28 vdd.n14 8.42249
R20227 vdd.n1727 vdd.t62 8.27616
R20228 vdd.n3436 vdd.t110 8.27616
R20229 vdd.n3440 vdd.n3439 8.16225
R20230 vdd.n2012 vdd.n2011 8.16225
R20231 vdd.n284 vdd.n278 8.14595
R20232 vdd.n233 vdd.n227 8.14595
R20233 vdd.n190 vdd.n184 8.14595
R20234 vdd.n139 vdd.n133 8.14595
R20235 vdd.n97 vdd.n91 8.14595
R20236 vdd.n46 vdd.n40 8.14595
R20237 vdd.n1934 vdd.n1928 8.14595
R20238 vdd.n1985 vdd.n1979 8.14595
R20239 vdd.n1840 vdd.n1834 8.14595
R20240 vdd.n1891 vdd.n1885 8.14595
R20241 vdd.n1747 vdd.n1741 8.14595
R20242 vdd.n1798 vdd.n1792 8.14595
R20243 vdd.t117 vdd.n1415 8.04943
R20244 vdd.n3427 vdd.t98 8.04943
R20245 vdd.n2225 vdd.n962 7.70933
R20246 vdd.n2225 vdd.n965 7.70933
R20247 vdd.n2231 vdd.n951 7.70933
R20248 vdd.n2237 vdd.n951 7.70933
R20249 vdd.n2237 vdd.n944 7.70933
R20250 vdd.n2243 vdd.n944 7.70933
R20251 vdd.n2243 vdd.n947 7.70933
R20252 vdd.n2249 vdd.n940 7.70933
R20253 vdd.n2255 vdd.n934 7.70933
R20254 vdd.n2261 vdd.n921 7.70933
R20255 vdd.n2267 vdd.n921 7.70933
R20256 vdd.n2273 vdd.n915 7.70933
R20257 vdd.n2279 vdd.n908 7.70933
R20258 vdd.n2279 vdd.n911 7.70933
R20259 vdd.n2285 vdd.n904 7.70933
R20260 vdd.n2292 vdd.n890 7.70933
R20261 vdd.n2298 vdd.n890 7.70933
R20262 vdd.n2304 vdd.n884 7.70933
R20263 vdd.n2310 vdd.n880 7.70933
R20264 vdd.n2316 vdd.n874 7.70933
R20265 vdd.n2334 vdd.n856 7.70933
R20266 vdd.n2334 vdd.n849 7.70933
R20267 vdd.n2342 vdd.n849 7.70933
R20268 vdd.n2424 vdd.n833 7.70933
R20269 vdd.n2807 vdd.n785 7.70933
R20270 vdd.n2819 vdd.n774 7.70933
R20271 vdd.n2819 vdd.n768 7.70933
R20272 vdd.n2825 vdd.n768 7.70933
R20273 vdd.n2837 vdd.n759 7.70933
R20274 vdd.n2843 vdd.n753 7.70933
R20275 vdd.n2855 vdd.n740 7.70933
R20276 vdd.n2862 vdd.n733 7.70933
R20277 vdd.n2862 vdd.n736 7.70933
R20278 vdd.n2868 vdd.n729 7.70933
R20279 vdd.n2874 vdd.n715 7.70933
R20280 vdd.n2880 vdd.n715 7.70933
R20281 vdd.n2886 vdd.n709 7.70933
R20282 vdd.n2892 vdd.n702 7.70933
R20283 vdd.n2892 vdd.n705 7.70933
R20284 vdd.n2898 vdd.n698 7.70933
R20285 vdd.n2904 vdd.n692 7.70933
R20286 vdd.n2910 vdd.n679 7.70933
R20287 vdd.n2916 vdd.n679 7.70933
R20288 vdd.n2916 vdd.n671 7.70933
R20289 vdd.n2967 vdd.n671 7.70933
R20290 vdd.n2967 vdd.n674 7.70933
R20291 vdd.n2973 vdd.n631 7.70933
R20292 vdd.n3043 vdd.n631 7.70933
R20293 vdd.n283 vdd.n280 7.3702
R20294 vdd.n232 vdd.n229 7.3702
R20295 vdd.n189 vdd.n186 7.3702
R20296 vdd.n138 vdd.n135 7.3702
R20297 vdd.n96 vdd.n93 7.3702
R20298 vdd.n45 vdd.n42 7.3702
R20299 vdd.n1933 vdd.n1930 7.3702
R20300 vdd.n1984 vdd.n1981 7.3702
R20301 vdd.n1839 vdd.n1836 7.3702
R20302 vdd.n1890 vdd.n1887 7.3702
R20303 vdd.n1746 vdd.n1743 7.3702
R20304 vdd.n1797 vdd.n1794 7.3702
R20305 vdd.n934 vdd.t54 7.36923
R20306 vdd.n2898 vdd.t31 7.36923
R20307 vdd.n1694 vdd.t60 7.1425
R20308 vdd.n2249 vdd.t6 7.1425
R20309 vdd.n1253 vdd.t2 7.1425
R20310 vdd.n2831 vdd.t5 7.1425
R20311 vdd.n692 vdd.t15 7.1425
R20312 vdd.n3420 vdd.t132 7.1425
R20313 vdd.n1605 vdd.n1604 6.98232
R20314 vdd.n2113 vdd.n2112 6.98232
R20315 vdd.n3335 vdd.n3334 6.98232
R20316 vdd.n3127 vdd.n3126 6.98232
R20317 vdd.n1710 vdd.t66 6.91577
R20318 vdd.n325 vdd.t104 6.91577
R20319 vdd.n1253 vdd.t3 6.80241
R20320 vdd.n2831 vdd.t47 6.80241
R20321 vdd.n2017 vdd.t85 6.68904
R20322 vdd.n3261 vdd.t128 6.68904
R20323 vdd.n1380 vdd.t119 6.46231
R20324 vdd.n2273 vdd.t13 6.46231
R20325 vdd.t18 vdd.n884 6.46231
R20326 vdd.n2855 vdd.t23 6.46231
R20327 vdd.t39 vdd.n709 6.46231
R20328 vdd.t92 vdd.n492 6.46231
R20329 vdd.n2349 vdd.t51 6.34895
R20330 vdd.n2728 vdd.t36 6.34895
R20331 vdd.n3440 vdd.n309 6.27748
R20332 vdd.n2011 vdd.n2010 6.27748
R20333 vdd.n2870 vdd.n725 6.2444
R20334 vdd.n2289 vdd.n2288 6.2444
R20335 vdd.n2310 vdd.t44 5.89549
R20336 vdd.n753 vdd.t19 5.89549
R20337 vdd.n284 vdd.n283 5.81868
R20338 vdd.n233 vdd.n232 5.81868
R20339 vdd.n190 vdd.n189 5.81868
R20340 vdd.n139 vdd.n138 5.81868
R20341 vdd.n97 vdd.n96 5.81868
R20342 vdd.n46 vdd.n45 5.81868
R20343 vdd.n1934 vdd.n1933 5.81868
R20344 vdd.n1985 vdd.n1984 5.81868
R20345 vdd.n1840 vdd.n1839 5.81868
R20346 vdd.n1891 vdd.n1890 5.81868
R20347 vdd.n1747 vdd.n1746 5.81868
R20348 vdd.n1798 vdd.n1797 5.81868
R20349 vdd.n2432 vdd.n2431 5.77611
R20350 vdd.n1177 vdd.n1176 5.77611
R20351 vdd.n2740 vdd.n2739 5.77611
R20352 vdd.n2982 vdd.n663 5.77611
R20353 vdd.n3048 vdd.n627 5.77611
R20354 vdd.n2603 vdd.n2537 5.77611
R20355 vdd.n2357 vdd.n840 5.77611
R20356 vdd.n1313 vdd.n1145 5.77611
R20357 vdd.n1567 vdd.n1564 5.62474
R20358 vdd.n2076 vdd.n2073 5.62474
R20359 vdd.n3295 vdd.n3292 5.62474
R20360 vdd.n3082 vdd.n3079 5.62474
R20361 vdd.n2285 vdd.t33 5.55539
R20362 vdd.n729 vdd.t9 5.55539
R20363 vdd.n287 vdd.n278 5.04292
R20364 vdd.n236 vdd.n227 5.04292
R20365 vdd.n193 vdd.n184 5.04292
R20366 vdd.n142 vdd.n133 5.04292
R20367 vdd.n100 vdd.n91 5.04292
R20368 vdd.n49 vdd.n40 5.04292
R20369 vdd.n1937 vdd.n1928 5.04292
R20370 vdd.n1988 vdd.n1979 5.04292
R20371 vdd.n1843 vdd.n1834 5.04292
R20372 vdd.n1894 vdd.n1885 5.04292
R20373 vdd.n1750 vdd.n1741 5.04292
R20374 vdd.n1801 vdd.n1792 5.04292
R20375 vdd.n2043 vdd.t119 4.8752
R20376 vdd.t12 vdd.t24 4.8752
R20377 vdd.t55 vdd.t1 4.8752
R20378 vdd.n3236 vdd.t92 4.8752
R20379 vdd.n2433 vdd.n2432 4.83952
R20380 vdd.n1176 vdd.n1175 4.83952
R20381 vdd.n2741 vdd.n2740 4.83952
R20382 vdd.n663 vdd.n658 4.83952
R20383 vdd.n627 vdd.n622 4.83952
R20384 vdd.n2600 vdd.n2537 4.83952
R20385 vdd.n2360 vdd.n840 4.83952
R20386 vdd.n1316 vdd.n1145 4.83952
R20387 vdd.n1227 vdd.t21 4.76184
R20388 vdd.n2813 vdd.t7 4.76184
R20389 vdd.n2081 vdd.n2080 4.74817
R20390 vdd.n1349 vdd.n1344 4.74817
R20391 vdd.n1011 vdd.n1008 4.74817
R20392 vdd.n2174 vdd.n1007 4.74817
R20393 vdd.n2179 vdd.n1008 4.74817
R20394 vdd.n2178 vdd.n1007 4.74817
R20395 vdd.n521 vdd.n519 4.74817
R20396 vdd.n3197 vdd.n522 4.74817
R20397 vdd.n3200 vdd.n522 4.74817
R20398 vdd.n3201 vdd.n521 4.74817
R20399 vdd.n3089 vdd.n606 4.74817
R20400 vdd.n3085 vdd.n608 4.74817
R20401 vdd.n3088 vdd.n608 4.74817
R20402 vdd.n3093 vdd.n606 4.74817
R20403 vdd.n2080 vdd.n1107 4.74817
R20404 vdd.n1346 vdd.n1344 4.74817
R20405 vdd.n309 vdd.n308 4.7074
R20406 vdd.n215 vdd.n214 4.7074
R20407 vdd.n2010 vdd.n2009 4.7074
R20408 vdd.n1916 vdd.n1915 4.7074
R20409 vdd.t85 vdd.n1386 4.64847
R20410 vdd.t14 vdd.n915 4.64847
R20411 vdd.n2304 vdd.t53 4.64847
R20412 vdd.t42 vdd.n740 4.64847
R20413 vdd.n2886 vdd.t38 4.64847
R20414 vdd.n3252 vdd.t128 4.64847
R20415 vdd.n904 vdd.t224 4.53511
R20416 vdd.n2868 vdd.t187 4.53511
R20417 vdd.n1719 vdd.t66 4.42174
R20418 vdd.n2231 vdd.t165 4.42174
R20419 vdd.n1227 vdd.t210 4.42174
R20420 vdd.n2813 vdd.t217 4.42174
R20421 vdd.n674 vdd.t161 4.42174
R20422 vdd.n3434 vdd.t104 4.42174
R20423 vdd.n2859 vdd.n725 4.37123
R20424 vdd.n2290 vdd.n2289 4.37123
R20425 vdd.n2328 vdd.t40 4.30838
R20426 vdd.n2716 vdd.t27 4.30838
R20427 vdd.n288 vdd.n276 4.26717
R20428 vdd.n237 vdd.n225 4.26717
R20429 vdd.n194 vdd.n182 4.26717
R20430 vdd.n143 vdd.n131 4.26717
R20431 vdd.n101 vdd.n89 4.26717
R20432 vdd.n50 vdd.n38 4.26717
R20433 vdd.n1938 vdd.n1926 4.26717
R20434 vdd.n1989 vdd.n1977 4.26717
R20435 vdd.n1844 vdd.n1832 4.26717
R20436 vdd.n1895 vdd.n1883 4.26717
R20437 vdd.n1751 vdd.n1739 4.26717
R20438 vdd.n1802 vdd.n1790 4.26717
R20439 vdd.t60 vdd.n1414 4.19501
R20440 vdd.t132 vdd.n329 4.19501
R20441 vdd.n309 vdd.n215 4.10845
R20442 vdd.n2010 vdd.n1916 4.10845
R20443 vdd.n265 vdd.t108 4.06363
R20444 vdd.n265 vdd.t139 4.06363
R20445 vdd.n263 vdd.t141 4.06363
R20446 vdd.n263 vdd.t65 4.06363
R20447 vdd.n261 vdd.t84 4.06363
R20448 vdd.n261 vdd.t124 4.06363
R20449 vdd.n259 vdd.t142 4.06363
R20450 vdd.n259 vdd.t150 4.06363
R20451 vdd.n257 vdd.t153 4.06363
R20452 vdd.n257 vdd.t91 4.06363
R20453 vdd.n171 vdd.t99 4.06363
R20454 vdd.n171 vdd.t133 4.06363
R20455 vdd.n169 vdd.t134 4.06363
R20456 vdd.n169 vdd.t151 4.06363
R20457 vdd.n167 vdd.t71 4.06363
R20458 vdd.n167 vdd.t111 4.06363
R20459 vdd.n165 vdd.t137 4.06363
R20460 vdd.n165 vdd.t143 4.06363
R20461 vdd.n163 vdd.t147 4.06363
R20462 vdd.n163 vdd.t75 4.06363
R20463 vdd.n78 vdd.t116 4.06363
R20464 vdd.n78 vdd.t135 4.06363
R20465 vdd.n76 vdd.t105 4.06363
R20466 vdd.n76 vdd.t148 4.06363
R20467 vdd.n74 vdd.t83 4.06363
R20468 vdd.n74 vdd.t140 4.06363
R20469 vdd.n72 vdd.t78 4.06363
R20470 vdd.n72 vdd.t129 4.06363
R20471 vdd.n70 vdd.t93 4.06363
R20472 vdd.n70 vdd.t144 4.06363
R20473 vdd.n1958 vdd.t127 4.06363
R20474 vdd.n1958 vdd.t126 4.06363
R20475 vdd.n1960 vdd.t100 4.06363
R20476 vdd.n1960 vdd.t82 4.06363
R20477 vdd.n1962 vdd.t80 4.06363
R20478 vdd.n1962 vdd.t125 4.06363
R20479 vdd.n1964 vdd.t109 4.06363
R20480 vdd.n1964 vdd.t81 4.06363
R20481 vdd.n1966 vdd.t76 4.06363
R20482 vdd.n1966 vdd.t138 4.06363
R20483 vdd.n1864 vdd.t122 4.06363
R20484 vdd.n1864 vdd.t120 4.06363
R20485 vdd.n1866 vdd.t86 4.06363
R20486 vdd.n1866 vdd.t69 4.06363
R20487 vdd.n1868 vdd.t63 4.06363
R20488 vdd.n1868 vdd.t115 4.06363
R20489 vdd.n1870 vdd.t103 4.06363
R20490 vdd.n1870 vdd.t67 4.06363
R20491 vdd.n1872 vdd.t61 4.06363
R20492 vdd.n1872 vdd.t131 4.06363
R20493 vdd.n1771 vdd.t145 4.06363
R20494 vdd.n1771 vdd.t155 4.06363
R20495 vdd.n1773 vdd.t130 4.06363
R20496 vdd.n1773 vdd.t79 4.06363
R20497 vdd.n1775 vdd.t123 4.06363
R20498 vdd.n1775 vdd.t88 4.06363
R20499 vdd.n1777 vdd.t149 4.06363
R20500 vdd.n1777 vdd.t106 4.06363
R20501 vdd.n1779 vdd.t136 4.06363
R20502 vdd.n1779 vdd.t118 4.06363
R20503 vdd.n940 vdd.t46 3.96828
R20504 vdd.n2322 vdd.t26 3.96828
R20505 vdd.n2710 vdd.t43 3.96828
R20506 vdd.n2904 vdd.t32 3.96828
R20507 vdd.n26 vdd.t236 3.9605
R20508 vdd.n26 vdd.t158 3.9605
R20509 vdd.n23 vdd.t239 3.9605
R20510 vdd.n23 vdd.t240 3.9605
R20511 vdd.n21 vdd.t157 3.9605
R20512 vdd.n21 vdd.t242 3.9605
R20513 vdd.n20 vdd.t241 3.9605
R20514 vdd.n20 vdd.t59 3.9605
R20515 vdd.n15 vdd.t156 3.9605
R20516 vdd.n15 vdd.t237 3.9605
R20517 vdd.n16 vdd.t57 3.9605
R20518 vdd.n16 vdd.t58 3.9605
R20519 vdd.n18 vdd.t159 3.9605
R20520 vdd.n18 vdd.t238 3.9605
R20521 vdd.n25 vdd.t243 3.9605
R20522 vdd.n25 vdd.t0 3.9605
R20523 vdd.n2255 vdd.t46 3.74155
R20524 vdd.n874 vdd.t26 3.74155
R20525 vdd.n2837 vdd.t43 3.74155
R20526 vdd.n698 vdd.t32 3.74155
R20527 vdd.n7 vdd.t56 3.61217
R20528 vdd.n7 vdd.t20 3.61217
R20529 vdd.n8 vdd.t28 3.61217
R20530 vdd.n8 vdd.t48 3.61217
R20531 vdd.n10 vdd.t37 3.61217
R20532 vdd.n10 vdd.t8 3.61217
R20533 vdd.n12 vdd.t17 3.61217
R20534 vdd.n12 vdd.t35 3.61217
R20535 vdd.n5 vdd.t50 3.61217
R20536 vdd.n5 vdd.t30 3.61217
R20537 vdd.n3 vdd.t22 3.61217
R20538 vdd.n3 vdd.t52 3.61217
R20539 vdd.n1 vdd.t4 3.61217
R20540 vdd.n1 vdd.t41 3.61217
R20541 vdd.n0 vdd.t45 3.61217
R20542 vdd.n0 vdd.t25 3.61217
R20543 vdd.n292 vdd.n291 3.49141
R20544 vdd.n241 vdd.n240 3.49141
R20545 vdd.n198 vdd.n197 3.49141
R20546 vdd.n147 vdd.n146 3.49141
R20547 vdd.n105 vdd.n104 3.49141
R20548 vdd.n54 vdd.n53 3.49141
R20549 vdd.n1942 vdd.n1941 3.49141
R20550 vdd.n1993 vdd.n1992 3.49141
R20551 vdd.n1848 vdd.n1847 3.49141
R20552 vdd.n1899 vdd.n1898 3.49141
R20553 vdd.n1755 vdd.n1754 3.49141
R20554 vdd.n1806 vdd.n1805 3.49141
R20555 vdd.t40 vdd.n856 3.40145
R20556 vdd.n2496 vdd.t49 3.40145
R20557 vdd.n2800 vdd.t34 3.40145
R20558 vdd.n2825 vdd.t27 3.40145
R20559 vdd.n1702 vdd.t117 3.28809
R20560 vdd.n965 vdd.t165 3.28809
R20561 vdd.n2349 vdd.t210 3.28809
R20562 vdd.n2728 vdd.t217 3.28809
R20563 vdd.n2973 vdd.t161 3.28809
R20564 vdd.t98 vdd.n3426 3.28809
R20565 vdd.n1403 vdd.t62 3.06136
R20566 vdd.n2267 vdd.t14 3.06136
R20567 vdd.n1265 vdd.t53 3.06136
R20568 vdd.n2849 vdd.t42 3.06136
R20569 vdd.t38 vdd.n702 3.06136
R20570 vdd.t110 vdd.n3435 3.06136
R20571 vdd.n2342 vdd.t21 2.94799
R20572 vdd.t7 vdd.n774 2.94799
R20573 vdd.n2026 vdd.t68 2.83463
R20574 vdd.n3253 vdd.t77 2.83463
R20575 vdd.n295 vdd.n274 2.71565
R20576 vdd.n244 vdd.n223 2.71565
R20577 vdd.n201 vdd.n180 2.71565
R20578 vdd.n150 vdd.n129 2.71565
R20579 vdd.n108 vdd.n87 2.71565
R20580 vdd.n57 vdd.n36 2.71565
R20581 vdd.n1945 vdd.n1924 2.71565
R20582 vdd.n1996 vdd.n1975 2.71565
R20583 vdd.n1851 vdd.n1830 2.71565
R20584 vdd.n1902 vdd.n1881 2.71565
R20585 vdd.n1758 vdd.n1737 2.71565
R20586 vdd.n1809 vdd.n1788 2.71565
R20587 vdd.n2042 vdd.t89 2.6079
R20588 vdd.t112 vdd.n499 2.6079
R20589 vdd.n2316 vdd.t24 2.49453
R20590 vdd.n759 vdd.t55 2.49453
R20591 vdd.n282 vdd.n281 2.4129
R20592 vdd.n231 vdd.n230 2.4129
R20593 vdd.n188 vdd.n187 2.4129
R20594 vdd.n137 vdd.n136 2.4129
R20595 vdd.n95 vdd.n94 2.4129
R20596 vdd.n44 vdd.n43 2.4129
R20597 vdd.n1932 vdd.n1931 2.4129
R20598 vdd.n1983 vdd.n1982 2.4129
R20599 vdd.n1838 vdd.n1837 2.4129
R20600 vdd.n1889 vdd.n1888 2.4129
R20601 vdd.n1745 vdd.n1744 2.4129
R20602 vdd.n1796 vdd.n1795 2.4129
R20603 vdd.n2186 vdd.n1008 2.27742
R20604 vdd.n2186 vdd.n1007 2.27742
R20605 vdd.n3009 vdd.n522 2.27742
R20606 vdd.n3009 vdd.n521 2.27742
R20607 vdd.n3077 vdd.n608 2.27742
R20608 vdd.n3077 vdd.n606 2.27742
R20609 vdd.n2080 vdd.n2079 2.27742
R20610 vdd.n2079 vdd.n1344 2.27742
R20611 vdd.n911 vdd.t33 2.15444
R20612 vdd.n2292 vdd.t11 2.15444
R20613 vdd.n736 vdd.t10 2.15444
R20614 vdd.n2874 vdd.t9 2.15444
R20615 vdd.n296 vdd.n272 1.93989
R20616 vdd.n245 vdd.n221 1.93989
R20617 vdd.n202 vdd.n178 1.93989
R20618 vdd.n151 vdd.n127 1.93989
R20619 vdd.n109 vdd.n85 1.93989
R20620 vdd.n58 vdd.n34 1.93989
R20621 vdd.n1946 vdd.n1922 1.93989
R20622 vdd.n1997 vdd.n1973 1.93989
R20623 vdd.n1852 vdd.n1828 1.93989
R20624 vdd.n1903 vdd.n1879 1.93989
R20625 vdd.n1759 vdd.n1735 1.93989
R20626 vdd.n1810 vdd.n1786 1.93989
R20627 vdd.n1265 vdd.t44 1.81434
R20628 vdd.n2849 vdd.t19 1.81434
R20629 vdd.n1438 vdd.t197 1.47425
R20630 vdd.t183 vdd.n3411 1.47425
R20631 vdd.t51 vdd.n833 1.36088
R20632 vdd.n2807 vdd.t36 1.36088
R20633 vdd.t13 vdd.n908 1.24752
R20634 vdd.n2298 vdd.t18 1.24752
R20635 vdd.t23 vdd.n733 1.24752
R20636 vdd.n2880 vdd.t39 1.24752
R20637 vdd.n307 vdd.n267 1.16414
R20638 vdd.n300 vdd.n299 1.16414
R20639 vdd.n256 vdd.n216 1.16414
R20640 vdd.n249 vdd.n248 1.16414
R20641 vdd.n213 vdd.n173 1.16414
R20642 vdd.n206 vdd.n205 1.16414
R20643 vdd.n162 vdd.n122 1.16414
R20644 vdd.n155 vdd.n154 1.16414
R20645 vdd.n120 vdd.n80 1.16414
R20646 vdd.n113 vdd.n112 1.16414
R20647 vdd.n69 vdd.n29 1.16414
R20648 vdd.n62 vdd.n61 1.16414
R20649 vdd.n1957 vdd.n1917 1.16414
R20650 vdd.n1950 vdd.n1949 1.16414
R20651 vdd.n2008 vdd.n1968 1.16414
R20652 vdd.n2001 vdd.n2000 1.16414
R20653 vdd.n1863 vdd.n1823 1.16414
R20654 vdd.n1856 vdd.n1855 1.16414
R20655 vdd.n1914 vdd.n1874 1.16414
R20656 vdd.n1907 vdd.n1906 1.16414
R20657 vdd.n1770 vdd.n1730 1.16414
R20658 vdd.n1763 vdd.n1762 1.16414
R20659 vdd.n1821 vdd.n1781 1.16414
R20660 vdd.n1814 vdd.n1813 1.16414
R20661 vdd.n2011 vdd.n28 1.11236
R20662 vdd vdd.n3440 1.10453
R20663 vdd.n2034 vdd.t121 1.02079
R20664 vdd.t224 vdd.t11 1.02079
R20665 vdd.t10 vdd.t187 1.02079
R20666 vdd.n3244 vdd.t74 1.02079
R20667 vdd.n1568 vdd.n1567 0.970197
R20668 vdd.n2077 vdd.n2076 0.970197
R20669 vdd.n3296 vdd.n3295 0.970197
R20670 vdd.n3084 vdd.n3082 0.970197
R20671 vdd.n2322 vdd.t3 0.907421
R20672 vdd.n2710 vdd.t47 0.907421
R20673 vdd.t87 vdd.n1392 0.794056
R20674 vdd.n2061 vdd.t169 0.794056
R20675 vdd.t179 vdd.n511 0.794056
R20676 vdd.n481 vdd.t70 0.794056
R20677 vdd.n1711 vdd.t102 0.567326
R20678 vdd.n947 vdd.t6 0.567326
R20679 vdd.n2328 vdd.t2 0.567326
R20680 vdd.n2716 vdd.t5 0.567326
R20681 vdd.n2910 vdd.t15 0.567326
R20682 vdd.n3428 vdd.t64 0.567326
R20683 vdd.n2067 vdd.n1009 0.509646
R20684 vdd.n3209 vdd.n3208 0.509646
R20685 vdd.n3407 vdd.n3406 0.509646
R20686 vdd.n3289 vdd.n3288 0.509646
R20687 vdd.n3215 vdd.n514 0.509646
R20688 vdd.n2056 vdd.n1345 0.509646
R20689 vdd.n1673 vdd.n1435 0.509646
R20690 vdd.n1667 vdd.n1666 0.509646
R20691 vdd.n4 vdd.n2 0.459552
R20692 vdd.n11 vdd.n9 0.459552
R20693 vdd.n305 vdd.n304 0.388379
R20694 vdd.n271 vdd.n269 0.388379
R20695 vdd.n254 vdd.n253 0.388379
R20696 vdd.n220 vdd.n218 0.388379
R20697 vdd.n211 vdd.n210 0.388379
R20698 vdd.n177 vdd.n175 0.388379
R20699 vdd.n160 vdd.n159 0.388379
R20700 vdd.n126 vdd.n124 0.388379
R20701 vdd.n118 vdd.n117 0.388379
R20702 vdd.n84 vdd.n82 0.388379
R20703 vdd.n67 vdd.n66 0.388379
R20704 vdd.n33 vdd.n31 0.388379
R20705 vdd.n1955 vdd.n1954 0.388379
R20706 vdd.n1921 vdd.n1919 0.388379
R20707 vdd.n2006 vdd.n2005 0.388379
R20708 vdd.n1972 vdd.n1970 0.388379
R20709 vdd.n1861 vdd.n1860 0.388379
R20710 vdd.n1827 vdd.n1825 0.388379
R20711 vdd.n1912 vdd.n1911 0.388379
R20712 vdd.n1878 vdd.n1876 0.388379
R20713 vdd.n1768 vdd.n1767 0.388379
R20714 vdd.n1734 vdd.n1732 0.388379
R20715 vdd.n1819 vdd.n1818 0.388379
R20716 vdd.n1785 vdd.n1783 0.388379
R20717 vdd.n19 vdd.n17 0.387128
R20718 vdd.n24 vdd.n22 0.387128
R20719 vdd.n6 vdd.n4 0.358259
R20720 vdd.n13 vdd.n11 0.358259
R20721 vdd.n260 vdd.n258 0.358259
R20722 vdd.n262 vdd.n260 0.358259
R20723 vdd.n264 vdd.n262 0.358259
R20724 vdd.n266 vdd.n264 0.358259
R20725 vdd.n308 vdd.n266 0.358259
R20726 vdd.n166 vdd.n164 0.358259
R20727 vdd.n168 vdd.n166 0.358259
R20728 vdd.n170 vdd.n168 0.358259
R20729 vdd.n172 vdd.n170 0.358259
R20730 vdd.n214 vdd.n172 0.358259
R20731 vdd.n73 vdd.n71 0.358259
R20732 vdd.n75 vdd.n73 0.358259
R20733 vdd.n77 vdd.n75 0.358259
R20734 vdd.n79 vdd.n77 0.358259
R20735 vdd.n121 vdd.n79 0.358259
R20736 vdd.n2009 vdd.n1967 0.358259
R20737 vdd.n1967 vdd.n1965 0.358259
R20738 vdd.n1965 vdd.n1963 0.358259
R20739 vdd.n1963 vdd.n1961 0.358259
R20740 vdd.n1961 vdd.n1959 0.358259
R20741 vdd.n1915 vdd.n1873 0.358259
R20742 vdd.n1873 vdd.n1871 0.358259
R20743 vdd.n1871 vdd.n1869 0.358259
R20744 vdd.n1869 vdd.n1867 0.358259
R20745 vdd.n1867 vdd.n1865 0.358259
R20746 vdd.n1822 vdd.n1780 0.358259
R20747 vdd.n1780 vdd.n1778 0.358259
R20748 vdd.n1778 vdd.n1776 0.358259
R20749 vdd.n1776 vdd.n1774 0.358259
R20750 vdd.n1774 vdd.n1772 0.358259
R20751 vdd.t94 vdd.n1421 0.340595
R20752 vdd.n2261 vdd.t54 0.340595
R20753 vdd.n880 vdd.t12 0.340595
R20754 vdd.n2843 vdd.t1 0.340595
R20755 vdd.n705 vdd.t31 0.340595
R20756 vdd.n3419 vdd.t72 0.340595
R20757 vdd.n14 vdd.n6 0.334552
R20758 vdd.n14 vdd.n13 0.334552
R20759 vdd.n27 vdd.n19 0.21707
R20760 vdd.n27 vdd.n24 0.21707
R20761 vdd.n306 vdd.n268 0.155672
R20762 vdd.n298 vdd.n268 0.155672
R20763 vdd.n298 vdd.n297 0.155672
R20764 vdd.n297 vdd.n273 0.155672
R20765 vdd.n290 vdd.n273 0.155672
R20766 vdd.n290 vdd.n289 0.155672
R20767 vdd.n289 vdd.n277 0.155672
R20768 vdd.n282 vdd.n277 0.155672
R20769 vdd.n255 vdd.n217 0.155672
R20770 vdd.n247 vdd.n217 0.155672
R20771 vdd.n247 vdd.n246 0.155672
R20772 vdd.n246 vdd.n222 0.155672
R20773 vdd.n239 vdd.n222 0.155672
R20774 vdd.n239 vdd.n238 0.155672
R20775 vdd.n238 vdd.n226 0.155672
R20776 vdd.n231 vdd.n226 0.155672
R20777 vdd.n212 vdd.n174 0.155672
R20778 vdd.n204 vdd.n174 0.155672
R20779 vdd.n204 vdd.n203 0.155672
R20780 vdd.n203 vdd.n179 0.155672
R20781 vdd.n196 vdd.n179 0.155672
R20782 vdd.n196 vdd.n195 0.155672
R20783 vdd.n195 vdd.n183 0.155672
R20784 vdd.n188 vdd.n183 0.155672
R20785 vdd.n161 vdd.n123 0.155672
R20786 vdd.n153 vdd.n123 0.155672
R20787 vdd.n153 vdd.n152 0.155672
R20788 vdd.n152 vdd.n128 0.155672
R20789 vdd.n145 vdd.n128 0.155672
R20790 vdd.n145 vdd.n144 0.155672
R20791 vdd.n144 vdd.n132 0.155672
R20792 vdd.n137 vdd.n132 0.155672
R20793 vdd.n119 vdd.n81 0.155672
R20794 vdd.n111 vdd.n81 0.155672
R20795 vdd.n111 vdd.n110 0.155672
R20796 vdd.n110 vdd.n86 0.155672
R20797 vdd.n103 vdd.n86 0.155672
R20798 vdd.n103 vdd.n102 0.155672
R20799 vdd.n102 vdd.n90 0.155672
R20800 vdd.n95 vdd.n90 0.155672
R20801 vdd.n68 vdd.n30 0.155672
R20802 vdd.n60 vdd.n30 0.155672
R20803 vdd.n60 vdd.n59 0.155672
R20804 vdd.n59 vdd.n35 0.155672
R20805 vdd.n52 vdd.n35 0.155672
R20806 vdd.n52 vdd.n51 0.155672
R20807 vdd.n51 vdd.n39 0.155672
R20808 vdd.n44 vdd.n39 0.155672
R20809 vdd.n1956 vdd.n1918 0.155672
R20810 vdd.n1948 vdd.n1918 0.155672
R20811 vdd.n1948 vdd.n1947 0.155672
R20812 vdd.n1947 vdd.n1923 0.155672
R20813 vdd.n1940 vdd.n1923 0.155672
R20814 vdd.n1940 vdd.n1939 0.155672
R20815 vdd.n1939 vdd.n1927 0.155672
R20816 vdd.n1932 vdd.n1927 0.155672
R20817 vdd.n2007 vdd.n1969 0.155672
R20818 vdd.n1999 vdd.n1969 0.155672
R20819 vdd.n1999 vdd.n1998 0.155672
R20820 vdd.n1998 vdd.n1974 0.155672
R20821 vdd.n1991 vdd.n1974 0.155672
R20822 vdd.n1991 vdd.n1990 0.155672
R20823 vdd.n1990 vdd.n1978 0.155672
R20824 vdd.n1983 vdd.n1978 0.155672
R20825 vdd.n1862 vdd.n1824 0.155672
R20826 vdd.n1854 vdd.n1824 0.155672
R20827 vdd.n1854 vdd.n1853 0.155672
R20828 vdd.n1853 vdd.n1829 0.155672
R20829 vdd.n1846 vdd.n1829 0.155672
R20830 vdd.n1846 vdd.n1845 0.155672
R20831 vdd.n1845 vdd.n1833 0.155672
R20832 vdd.n1838 vdd.n1833 0.155672
R20833 vdd.n1913 vdd.n1875 0.155672
R20834 vdd.n1905 vdd.n1875 0.155672
R20835 vdd.n1905 vdd.n1904 0.155672
R20836 vdd.n1904 vdd.n1880 0.155672
R20837 vdd.n1897 vdd.n1880 0.155672
R20838 vdd.n1897 vdd.n1896 0.155672
R20839 vdd.n1896 vdd.n1884 0.155672
R20840 vdd.n1889 vdd.n1884 0.155672
R20841 vdd.n1769 vdd.n1731 0.155672
R20842 vdd.n1761 vdd.n1731 0.155672
R20843 vdd.n1761 vdd.n1760 0.155672
R20844 vdd.n1760 vdd.n1736 0.155672
R20845 vdd.n1753 vdd.n1736 0.155672
R20846 vdd.n1753 vdd.n1752 0.155672
R20847 vdd.n1752 vdd.n1740 0.155672
R20848 vdd.n1745 vdd.n1740 0.155672
R20849 vdd.n1820 vdd.n1782 0.155672
R20850 vdd.n1812 vdd.n1782 0.155672
R20851 vdd.n1812 vdd.n1811 0.155672
R20852 vdd.n1811 vdd.n1787 0.155672
R20853 vdd.n1804 vdd.n1787 0.155672
R20854 vdd.n1804 vdd.n1803 0.155672
R20855 vdd.n1803 vdd.n1791 0.155672
R20856 vdd.n1796 vdd.n1791 0.155672
R20857 vdd.n1014 vdd.n1006 0.152939
R20858 vdd.n1018 vdd.n1014 0.152939
R20859 vdd.n1019 vdd.n1018 0.152939
R20860 vdd.n1020 vdd.n1019 0.152939
R20861 vdd.n1021 vdd.n1020 0.152939
R20862 vdd.n1025 vdd.n1021 0.152939
R20863 vdd.n1026 vdd.n1025 0.152939
R20864 vdd.n1027 vdd.n1026 0.152939
R20865 vdd.n1028 vdd.n1027 0.152939
R20866 vdd.n1032 vdd.n1028 0.152939
R20867 vdd.n1033 vdd.n1032 0.152939
R20868 vdd.n1034 vdd.n1033 0.152939
R20869 vdd.n2150 vdd.n1034 0.152939
R20870 vdd.n2150 vdd.n2149 0.152939
R20871 vdd.n2149 vdd.n2148 0.152939
R20872 vdd.n2148 vdd.n1040 0.152939
R20873 vdd.n1045 vdd.n1040 0.152939
R20874 vdd.n1046 vdd.n1045 0.152939
R20875 vdd.n1047 vdd.n1046 0.152939
R20876 vdd.n1051 vdd.n1047 0.152939
R20877 vdd.n1052 vdd.n1051 0.152939
R20878 vdd.n1053 vdd.n1052 0.152939
R20879 vdd.n1054 vdd.n1053 0.152939
R20880 vdd.n1058 vdd.n1054 0.152939
R20881 vdd.n1059 vdd.n1058 0.152939
R20882 vdd.n1060 vdd.n1059 0.152939
R20883 vdd.n1061 vdd.n1060 0.152939
R20884 vdd.n1065 vdd.n1061 0.152939
R20885 vdd.n1066 vdd.n1065 0.152939
R20886 vdd.n1067 vdd.n1066 0.152939
R20887 vdd.n1068 vdd.n1067 0.152939
R20888 vdd.n1072 vdd.n1068 0.152939
R20889 vdd.n1073 vdd.n1072 0.152939
R20890 vdd.n1074 vdd.n1073 0.152939
R20891 vdd.n2111 vdd.n1074 0.152939
R20892 vdd.n2111 vdd.n2110 0.152939
R20893 vdd.n2110 vdd.n2109 0.152939
R20894 vdd.n2109 vdd.n1080 0.152939
R20895 vdd.n1085 vdd.n1080 0.152939
R20896 vdd.n1086 vdd.n1085 0.152939
R20897 vdd.n1087 vdd.n1086 0.152939
R20898 vdd.n1091 vdd.n1087 0.152939
R20899 vdd.n1092 vdd.n1091 0.152939
R20900 vdd.n1093 vdd.n1092 0.152939
R20901 vdd.n1094 vdd.n1093 0.152939
R20902 vdd.n1098 vdd.n1094 0.152939
R20903 vdd.n1099 vdd.n1098 0.152939
R20904 vdd.n1100 vdd.n1099 0.152939
R20905 vdd.n1101 vdd.n1100 0.152939
R20906 vdd.n1105 vdd.n1101 0.152939
R20907 vdd.n1106 vdd.n1105 0.152939
R20908 vdd.n2185 vdd.n1009 0.152939
R20909 vdd.n2014 vdd.n2013 0.152939
R20910 vdd.n2014 vdd.n1383 0.152939
R20911 vdd.n2029 vdd.n1383 0.152939
R20912 vdd.n2030 vdd.n2029 0.152939
R20913 vdd.n2031 vdd.n2030 0.152939
R20914 vdd.n2031 vdd.n1372 0.152939
R20915 vdd.n2046 vdd.n1372 0.152939
R20916 vdd.n2047 vdd.n2046 0.152939
R20917 vdd.n2048 vdd.n2047 0.152939
R20918 vdd.n2048 vdd.n1360 0.152939
R20919 vdd.n2065 vdd.n1360 0.152939
R20920 vdd.n2066 vdd.n2065 0.152939
R20921 vdd.n2067 vdd.n2066 0.152939
R20922 vdd.n527 vdd.n524 0.152939
R20923 vdd.n528 vdd.n527 0.152939
R20924 vdd.n529 vdd.n528 0.152939
R20925 vdd.n530 vdd.n529 0.152939
R20926 vdd.n533 vdd.n530 0.152939
R20927 vdd.n534 vdd.n533 0.152939
R20928 vdd.n535 vdd.n534 0.152939
R20929 vdd.n536 vdd.n535 0.152939
R20930 vdd.n539 vdd.n536 0.152939
R20931 vdd.n540 vdd.n539 0.152939
R20932 vdd.n541 vdd.n540 0.152939
R20933 vdd.n542 vdd.n541 0.152939
R20934 vdd.n547 vdd.n542 0.152939
R20935 vdd.n548 vdd.n547 0.152939
R20936 vdd.n549 vdd.n548 0.152939
R20937 vdd.n550 vdd.n549 0.152939
R20938 vdd.n553 vdd.n550 0.152939
R20939 vdd.n554 vdd.n553 0.152939
R20940 vdd.n555 vdd.n554 0.152939
R20941 vdd.n556 vdd.n555 0.152939
R20942 vdd.n559 vdd.n556 0.152939
R20943 vdd.n560 vdd.n559 0.152939
R20944 vdd.n561 vdd.n560 0.152939
R20945 vdd.n562 vdd.n561 0.152939
R20946 vdd.n565 vdd.n562 0.152939
R20947 vdd.n566 vdd.n565 0.152939
R20948 vdd.n567 vdd.n566 0.152939
R20949 vdd.n568 vdd.n567 0.152939
R20950 vdd.n571 vdd.n568 0.152939
R20951 vdd.n572 vdd.n571 0.152939
R20952 vdd.n573 vdd.n572 0.152939
R20953 vdd.n574 vdd.n573 0.152939
R20954 vdd.n577 vdd.n574 0.152939
R20955 vdd.n578 vdd.n577 0.152939
R20956 vdd.n3125 vdd.n578 0.152939
R20957 vdd.n3125 vdd.n3124 0.152939
R20958 vdd.n3124 vdd.n3123 0.152939
R20959 vdd.n3123 vdd.n582 0.152939
R20960 vdd.n587 vdd.n582 0.152939
R20961 vdd.n588 vdd.n587 0.152939
R20962 vdd.n591 vdd.n588 0.152939
R20963 vdd.n592 vdd.n591 0.152939
R20964 vdd.n593 vdd.n592 0.152939
R20965 vdd.n594 vdd.n593 0.152939
R20966 vdd.n597 vdd.n594 0.152939
R20967 vdd.n598 vdd.n597 0.152939
R20968 vdd.n599 vdd.n598 0.152939
R20969 vdd.n600 vdd.n599 0.152939
R20970 vdd.n603 vdd.n600 0.152939
R20971 vdd.n604 vdd.n603 0.152939
R20972 vdd.n605 vdd.n604 0.152939
R20973 vdd.n3208 vdd.n518 0.152939
R20974 vdd.n3209 vdd.n508 0.152939
R20975 vdd.n3223 vdd.n508 0.152939
R20976 vdd.n3224 vdd.n3223 0.152939
R20977 vdd.n3225 vdd.n3224 0.152939
R20978 vdd.n3225 vdd.n496 0.152939
R20979 vdd.n3239 vdd.n496 0.152939
R20980 vdd.n3240 vdd.n3239 0.152939
R20981 vdd.n3241 vdd.n3240 0.152939
R20982 vdd.n3241 vdd.n484 0.152939
R20983 vdd.n3256 vdd.n484 0.152939
R20984 vdd.n3257 vdd.n3256 0.152939
R20985 vdd.n3258 vdd.n3257 0.152939
R20986 vdd.n3258 vdd.n310 0.152939
R20987 vdd.n320 vdd.n311 0.152939
R20988 vdd.n321 vdd.n320 0.152939
R20989 vdd.n322 vdd.n321 0.152939
R20990 vdd.n331 vdd.n322 0.152939
R20991 vdd.n332 vdd.n331 0.152939
R20992 vdd.n333 vdd.n332 0.152939
R20993 vdd.n334 vdd.n333 0.152939
R20994 vdd.n342 vdd.n334 0.152939
R20995 vdd.n343 vdd.n342 0.152939
R20996 vdd.n344 vdd.n343 0.152939
R20997 vdd.n345 vdd.n344 0.152939
R20998 vdd.n353 vdd.n345 0.152939
R20999 vdd.n3407 vdd.n353 0.152939
R21000 vdd.n3406 vdd.n354 0.152939
R21001 vdd.n357 vdd.n354 0.152939
R21002 vdd.n361 vdd.n357 0.152939
R21003 vdd.n362 vdd.n361 0.152939
R21004 vdd.n363 vdd.n362 0.152939
R21005 vdd.n364 vdd.n363 0.152939
R21006 vdd.n365 vdd.n364 0.152939
R21007 vdd.n369 vdd.n365 0.152939
R21008 vdd.n370 vdd.n369 0.152939
R21009 vdd.n371 vdd.n370 0.152939
R21010 vdd.n372 vdd.n371 0.152939
R21011 vdd.n376 vdd.n372 0.152939
R21012 vdd.n377 vdd.n376 0.152939
R21013 vdd.n378 vdd.n377 0.152939
R21014 vdd.n379 vdd.n378 0.152939
R21015 vdd.n383 vdd.n379 0.152939
R21016 vdd.n384 vdd.n383 0.152939
R21017 vdd.n385 vdd.n384 0.152939
R21018 vdd.n3372 vdd.n385 0.152939
R21019 vdd.n3372 vdd.n3371 0.152939
R21020 vdd.n3371 vdd.n3370 0.152939
R21021 vdd.n3370 vdd.n391 0.152939
R21022 vdd.n396 vdd.n391 0.152939
R21023 vdd.n397 vdd.n396 0.152939
R21024 vdd.n398 vdd.n397 0.152939
R21025 vdd.n402 vdd.n398 0.152939
R21026 vdd.n403 vdd.n402 0.152939
R21027 vdd.n404 vdd.n403 0.152939
R21028 vdd.n405 vdd.n404 0.152939
R21029 vdd.n409 vdd.n405 0.152939
R21030 vdd.n410 vdd.n409 0.152939
R21031 vdd.n411 vdd.n410 0.152939
R21032 vdd.n412 vdd.n411 0.152939
R21033 vdd.n416 vdd.n412 0.152939
R21034 vdd.n417 vdd.n416 0.152939
R21035 vdd.n418 vdd.n417 0.152939
R21036 vdd.n419 vdd.n418 0.152939
R21037 vdd.n423 vdd.n419 0.152939
R21038 vdd.n424 vdd.n423 0.152939
R21039 vdd.n425 vdd.n424 0.152939
R21040 vdd.n3333 vdd.n425 0.152939
R21041 vdd.n3333 vdd.n3332 0.152939
R21042 vdd.n3332 vdd.n3331 0.152939
R21043 vdd.n3331 vdd.n431 0.152939
R21044 vdd.n436 vdd.n431 0.152939
R21045 vdd.n437 vdd.n436 0.152939
R21046 vdd.n438 vdd.n437 0.152939
R21047 vdd.n442 vdd.n438 0.152939
R21048 vdd.n443 vdd.n442 0.152939
R21049 vdd.n444 vdd.n443 0.152939
R21050 vdd.n445 vdd.n444 0.152939
R21051 vdd.n449 vdd.n445 0.152939
R21052 vdd.n450 vdd.n449 0.152939
R21053 vdd.n451 vdd.n450 0.152939
R21054 vdd.n452 vdd.n451 0.152939
R21055 vdd.n456 vdd.n452 0.152939
R21056 vdd.n457 vdd.n456 0.152939
R21057 vdd.n458 vdd.n457 0.152939
R21058 vdd.n459 vdd.n458 0.152939
R21059 vdd.n463 vdd.n459 0.152939
R21060 vdd.n464 vdd.n463 0.152939
R21061 vdd.n465 vdd.n464 0.152939
R21062 vdd.n3289 vdd.n465 0.152939
R21063 vdd.n3216 vdd.n3215 0.152939
R21064 vdd.n3217 vdd.n3216 0.152939
R21065 vdd.n3217 vdd.n502 0.152939
R21066 vdd.n3231 vdd.n502 0.152939
R21067 vdd.n3232 vdd.n3231 0.152939
R21068 vdd.n3233 vdd.n3232 0.152939
R21069 vdd.n3233 vdd.n489 0.152939
R21070 vdd.n3247 vdd.n489 0.152939
R21071 vdd.n3248 vdd.n3247 0.152939
R21072 vdd.n3249 vdd.n3248 0.152939
R21073 vdd.n3249 vdd.n477 0.152939
R21074 vdd.n3264 vdd.n477 0.152939
R21075 vdd.n3265 vdd.n3264 0.152939
R21076 vdd.n3266 vdd.n3265 0.152939
R21077 vdd.n3266 vdd.n475 0.152939
R21078 vdd.n3270 vdd.n475 0.152939
R21079 vdd.n3271 vdd.n3270 0.152939
R21080 vdd.n3272 vdd.n3271 0.152939
R21081 vdd.n3272 vdd.n472 0.152939
R21082 vdd.n3276 vdd.n472 0.152939
R21083 vdd.n3277 vdd.n3276 0.152939
R21084 vdd.n3278 vdd.n3277 0.152939
R21085 vdd.n3278 vdd.n469 0.152939
R21086 vdd.n3282 vdd.n469 0.152939
R21087 vdd.n3283 vdd.n3282 0.152939
R21088 vdd.n3284 vdd.n3283 0.152939
R21089 vdd.n3284 vdd.n466 0.152939
R21090 vdd.n3288 vdd.n466 0.152939
R21091 vdd.n3078 vdd.n514 0.152939
R21092 vdd.n2078 vdd.n1345 0.152939
R21093 vdd.n1674 vdd.n1673 0.152939
R21094 vdd.n1675 vdd.n1674 0.152939
R21095 vdd.n1675 vdd.n1424 0.152939
R21096 vdd.n1689 vdd.n1424 0.152939
R21097 vdd.n1690 vdd.n1689 0.152939
R21098 vdd.n1691 vdd.n1690 0.152939
R21099 vdd.n1691 vdd.n1411 0.152939
R21100 vdd.n1705 vdd.n1411 0.152939
R21101 vdd.n1706 vdd.n1705 0.152939
R21102 vdd.n1707 vdd.n1706 0.152939
R21103 vdd.n1707 vdd.n1400 0.152939
R21104 vdd.n1722 vdd.n1400 0.152939
R21105 vdd.n1723 vdd.n1722 0.152939
R21106 vdd.n1724 vdd.n1723 0.152939
R21107 vdd.n1724 vdd.n1389 0.152939
R21108 vdd.n2020 vdd.n1389 0.152939
R21109 vdd.n2021 vdd.n2020 0.152939
R21110 vdd.n2022 vdd.n2021 0.152939
R21111 vdd.n2022 vdd.n1377 0.152939
R21112 vdd.n2037 vdd.n1377 0.152939
R21113 vdd.n2038 vdd.n2037 0.152939
R21114 vdd.n2039 vdd.n2038 0.152939
R21115 vdd.n2039 vdd.n1367 0.152939
R21116 vdd.n2054 vdd.n1367 0.152939
R21117 vdd.n2055 vdd.n2054 0.152939
R21118 vdd.n2058 vdd.n2055 0.152939
R21119 vdd.n2058 vdd.n2057 0.152939
R21120 vdd.n2057 vdd.n2056 0.152939
R21121 vdd.n1666 vdd.n1440 0.152939
R21122 vdd.n1662 vdd.n1440 0.152939
R21123 vdd.n1662 vdd.n1661 0.152939
R21124 vdd.n1661 vdd.n1660 0.152939
R21125 vdd.n1660 vdd.n1445 0.152939
R21126 vdd.n1656 vdd.n1445 0.152939
R21127 vdd.n1656 vdd.n1655 0.152939
R21128 vdd.n1655 vdd.n1654 0.152939
R21129 vdd.n1654 vdd.n1453 0.152939
R21130 vdd.n1650 vdd.n1453 0.152939
R21131 vdd.n1650 vdd.n1649 0.152939
R21132 vdd.n1649 vdd.n1648 0.152939
R21133 vdd.n1648 vdd.n1461 0.152939
R21134 vdd.n1644 vdd.n1461 0.152939
R21135 vdd.n1644 vdd.n1643 0.152939
R21136 vdd.n1643 vdd.n1642 0.152939
R21137 vdd.n1642 vdd.n1469 0.152939
R21138 vdd.n1638 vdd.n1469 0.152939
R21139 vdd.n1638 vdd.n1637 0.152939
R21140 vdd.n1637 vdd.n1636 0.152939
R21141 vdd.n1636 vdd.n1479 0.152939
R21142 vdd.n1632 vdd.n1479 0.152939
R21143 vdd.n1632 vdd.n1631 0.152939
R21144 vdd.n1631 vdd.n1630 0.152939
R21145 vdd.n1630 vdd.n1487 0.152939
R21146 vdd.n1626 vdd.n1487 0.152939
R21147 vdd.n1626 vdd.n1625 0.152939
R21148 vdd.n1625 vdd.n1624 0.152939
R21149 vdd.n1624 vdd.n1495 0.152939
R21150 vdd.n1620 vdd.n1495 0.152939
R21151 vdd.n1620 vdd.n1619 0.152939
R21152 vdd.n1619 vdd.n1618 0.152939
R21153 vdd.n1618 vdd.n1503 0.152939
R21154 vdd.n1614 vdd.n1503 0.152939
R21155 vdd.n1614 vdd.n1613 0.152939
R21156 vdd.n1613 vdd.n1612 0.152939
R21157 vdd.n1612 vdd.n1511 0.152939
R21158 vdd.n1608 vdd.n1511 0.152939
R21159 vdd.n1608 vdd.n1607 0.152939
R21160 vdd.n1607 vdd.n1606 0.152939
R21161 vdd.n1606 vdd.n1519 0.152939
R21162 vdd.n1526 vdd.n1519 0.152939
R21163 vdd.n1596 vdd.n1526 0.152939
R21164 vdd.n1596 vdd.n1595 0.152939
R21165 vdd.n1595 vdd.n1594 0.152939
R21166 vdd.n1594 vdd.n1527 0.152939
R21167 vdd.n1590 vdd.n1527 0.152939
R21168 vdd.n1590 vdd.n1589 0.152939
R21169 vdd.n1589 vdd.n1588 0.152939
R21170 vdd.n1588 vdd.n1534 0.152939
R21171 vdd.n1584 vdd.n1534 0.152939
R21172 vdd.n1584 vdd.n1583 0.152939
R21173 vdd.n1583 vdd.n1582 0.152939
R21174 vdd.n1582 vdd.n1542 0.152939
R21175 vdd.n1578 vdd.n1542 0.152939
R21176 vdd.n1578 vdd.n1577 0.152939
R21177 vdd.n1577 vdd.n1576 0.152939
R21178 vdd.n1576 vdd.n1550 0.152939
R21179 vdd.n1572 vdd.n1550 0.152939
R21180 vdd.n1572 vdd.n1571 0.152939
R21181 vdd.n1571 vdd.n1570 0.152939
R21182 vdd.n1570 vdd.n1558 0.152939
R21183 vdd.n1558 vdd.n1435 0.152939
R21184 vdd.n1667 vdd.n1430 0.152939
R21185 vdd.n1681 vdd.n1430 0.152939
R21186 vdd.n1682 vdd.n1681 0.152939
R21187 vdd.n1683 vdd.n1682 0.152939
R21188 vdd.n1683 vdd.n1418 0.152939
R21189 vdd.n1697 vdd.n1418 0.152939
R21190 vdd.n1698 vdd.n1697 0.152939
R21191 vdd.n1699 vdd.n1698 0.152939
R21192 vdd.n1699 vdd.n1406 0.152939
R21193 vdd.n1714 vdd.n1406 0.152939
R21194 vdd.n1715 vdd.n1714 0.152939
R21195 vdd.n1716 vdd.n1715 0.152939
R21196 vdd.n1716 vdd.n1395 0.152939
R21197 vdd.n2013 vdd.n2012 0.145814
R21198 vdd.n3439 vdd.n310 0.145814
R21199 vdd.n3439 vdd.n311 0.145814
R21200 vdd.n2012 vdd.n1395 0.145814
R21201 vdd.n2186 vdd.n2185 0.110256
R21202 vdd.n3009 vdd.n518 0.110256
R21203 vdd.n3078 vdd.n3077 0.110256
R21204 vdd.n2079 vdd.n2078 0.110256
R21205 vdd.n2186 vdd.n1006 0.0431829
R21206 vdd.n2079 vdd.n1106 0.0431829
R21207 vdd.n3009 vdd.n524 0.0431829
R21208 vdd.n3077 vdd.n605 0.0431829
R21209 vdd vdd.n28 0.00833333
R21210 commonsourceibias.n35 commonsourceibias.t0 223.028
R21211 commonsourceibias.n128 commonsourceibias.t129 223.028
R21212 commonsourceibias.n307 commonsourceibias.t140 223.028
R21213 commonsourceibias.n217 commonsourceibias.t112 223.028
R21214 commonsourceibias.n454 commonsourceibias.t22 223.028
R21215 commonsourceibias.n395 commonsourceibias.t108 223.028
R21216 commonsourceibias.n679 commonsourceibias.t74 223.028
R21217 commonsourceibias.n589 commonsourceibias.t97 223.028
R21218 commonsourceibias.n99 commonsourceibias.t12 207.983
R21219 commonsourceibias.n192 commonsourceibias.t120 207.983
R21220 commonsourceibias.n371 commonsourceibias.t147 207.983
R21221 commonsourceibias.n281 commonsourceibias.t71 207.983
R21222 commonsourceibias.n520 commonsourceibias.t34 207.983
R21223 commonsourceibias.n566 commonsourceibias.t91 207.983
R21224 commonsourceibias.n745 commonsourceibias.t82 207.983
R21225 commonsourceibias.n655 commonsourceibias.t151 207.983
R21226 commonsourceibias.n97 commonsourceibias.t48 168.701
R21227 commonsourceibias.n91 commonsourceibias.t4 168.701
R21228 commonsourceibias.n17 commonsourceibias.t10 168.701
R21229 commonsourceibias.n83 commonsourceibias.t58 168.701
R21230 commonsourceibias.n77 commonsourceibias.t16 168.701
R21231 commonsourceibias.n22 commonsourceibias.t28 168.701
R21232 commonsourceibias.n69 commonsourceibias.t6 168.701
R21233 commonsourceibias.n63 commonsourceibias.t14 168.701
R21234 commonsourceibias.n25 commonsourceibias.t44 168.701
R21235 commonsourceibias.n27 commonsourceibias.t24 168.701
R21236 commonsourceibias.n29 commonsourceibias.t30 168.701
R21237 commonsourceibias.n46 commonsourceibias.t54 168.701
R21238 commonsourceibias.n40 commonsourceibias.t18 168.701
R21239 commonsourceibias.n34 commonsourceibias.t50 168.701
R21240 commonsourceibias.n190 commonsourceibias.t67 168.701
R21241 commonsourceibias.n184 commonsourceibias.t126 168.701
R21242 commonsourceibias.n5 commonsourceibias.t121 168.701
R21243 commonsourceibias.n176 commonsourceibias.t136 168.701
R21244 commonsourceibias.n170 commonsourceibias.t117 168.701
R21245 commonsourceibias.n10 commonsourceibias.t102 168.701
R21246 commonsourceibias.n162 commonsourceibias.t125 168.701
R21247 commonsourceibias.n156 commonsourceibias.t118 168.701
R21248 commonsourceibias.n118 commonsourceibias.t76 168.701
R21249 commonsourceibias.n120 commonsourceibias.t106 168.701
R21250 commonsourceibias.n122 commonsourceibias.t96 168.701
R21251 commonsourceibias.n139 commonsourceibias.t141 168.701
R21252 commonsourceibias.n133 commonsourceibias.t116 168.701
R21253 commonsourceibias.n127 commonsourceibias.t152 168.701
R21254 commonsourceibias.n306 commonsourceibias.t130 168.701
R21255 commonsourceibias.n312 commonsourceibias.t79 168.701
R21256 commonsourceibias.n318 commonsourceibias.t149 168.701
R21257 commonsourceibias.n301 commonsourceibias.t133 168.701
R21258 commonsourceibias.n299 commonsourceibias.t137 168.701
R21259 commonsourceibias.n297 commonsourceibias.t64 168.701
R21260 commonsourceibias.n335 commonsourceibias.t138 168.701
R21261 commonsourceibias.n341 commonsourceibias.t146 168.701
R21262 commonsourceibias.n294 commonsourceibias.t119 168.701
R21263 commonsourceibias.n349 commonsourceibias.t90 168.701
R21264 commonsourceibias.n355 commonsourceibias.t155 168.701
R21265 commonsourceibias.n289 commonsourceibias.t124 168.701
R21266 commonsourceibias.n363 commonsourceibias.t128 168.701
R21267 commonsourceibias.n369 commonsourceibias.t75 168.701
R21268 commonsourceibias.n279 commonsourceibias.t159 168.701
R21269 commonsourceibias.n273 commonsourceibias.t148 168.701
R21270 commonsourceibias.n199 commonsourceibias.t78 168.701
R21271 commonsourceibias.n265 commonsourceibias.t157 168.701
R21272 commonsourceibias.n259 commonsourceibias.t85 168.701
R21273 commonsourceibias.n204 commonsourceibias.t77 168.701
R21274 commonsourceibias.n251 commonsourceibias.t158 168.701
R21275 commonsourceibias.n245 commonsourceibias.t94 168.701
R21276 commonsourceibias.n207 commonsourceibias.t113 168.701
R21277 commonsourceibias.n209 commonsourceibias.t156 168.701
R21278 commonsourceibias.n211 commonsourceibias.t92 168.701
R21279 commonsourceibias.n228 commonsourceibias.t111 168.701
R21280 commonsourceibias.n222 commonsourceibias.t105 168.701
R21281 commonsourceibias.n216 commonsourceibias.t93 168.701
R21282 commonsourceibias.n453 commonsourceibias.t62 168.701
R21283 commonsourceibias.n459 commonsourceibias.t40 168.701
R21284 commonsourceibias.n465 commonsourceibias.t2 168.701
R21285 commonsourceibias.n448 commonsourceibias.t52 168.701
R21286 commonsourceibias.n446 commonsourceibias.t42 168.701
R21287 commonsourceibias.n444 commonsourceibias.t56 168.701
R21288 commonsourceibias.n482 commonsourceibias.t36 168.701
R21289 commonsourceibias.n488 commonsourceibias.t26 168.701
R21290 commonsourceibias.n490 commonsourceibias.t46 168.701
R21291 commonsourceibias.n497 commonsourceibias.t38 168.701
R21292 commonsourceibias.n503 commonsourceibias.t8 168.701
R21293 commonsourceibias.n505 commonsourceibias.t32 168.701
R21294 commonsourceibias.n512 commonsourceibias.t20 168.701
R21295 commonsourceibias.n518 commonsourceibias.t60 168.701
R21296 commonsourceibias.n564 commonsourceibias.t134 168.701
R21297 commonsourceibias.n558 commonsourceibias.t114 168.701
R21298 commonsourceibias.n551 commonsourceibias.t95 168.701
R21299 commonsourceibias.n549 commonsourceibias.t123 168.701
R21300 commonsourceibias.n543 commonsourceibias.t88 168.701
R21301 commonsourceibias.n536 commonsourceibias.t73 168.701
R21302 commonsourceibias.n534 commonsourceibias.t104 168.701
R21303 commonsourceibias.n394 commonsourceibias.t131 168.701
R21304 commonsourceibias.n400 commonsourceibias.t84 168.701
R21305 commonsourceibias.n406 commonsourceibias.t127 168.701
R21306 commonsourceibias.n389 commonsourceibias.t150 168.701
R21307 commonsourceibias.n387 commonsourceibias.t83 168.701
R21308 commonsourceibias.n385 commonsourceibias.t139 168.701
R21309 commonsourceibias.n423 commonsourceibias.t89 168.701
R21310 commonsourceibias.n678 commonsourceibias.t145 168.701
R21311 commonsourceibias.n684 commonsourceibias.t109 168.701
R21312 commonsourceibias.n690 commonsourceibias.t87 168.701
R21313 commonsourceibias.n673 commonsourceibias.t153 168.701
R21314 commonsourceibias.n671 commonsourceibias.t132 168.701
R21315 commonsourceibias.n669 commonsourceibias.t103 168.701
R21316 commonsourceibias.n707 commonsourceibias.t70 168.701
R21317 commonsourceibias.n713 commonsourceibias.t81 168.701
R21318 commonsourceibias.n715 commonsourceibias.t110 168.701
R21319 commonsourceibias.n722 commonsourceibias.t115 168.701
R21320 commonsourceibias.n728 commonsourceibias.t101 168.701
R21321 commonsourceibias.n730 commonsourceibias.t135 168.701
R21322 commonsourceibias.n737 commonsourceibias.t122 168.701
R21323 commonsourceibias.n743 commonsourceibias.t107 168.701
R21324 commonsourceibias.n588 commonsourceibias.t68 168.701
R21325 commonsourceibias.n594 commonsourceibias.t86 168.701
R21326 commonsourceibias.n600 commonsourceibias.t98 168.701
R21327 commonsourceibias.n583 commonsourceibias.t69 168.701
R21328 commonsourceibias.n581 commonsourceibias.t80 168.701
R21329 commonsourceibias.n579 commonsourceibias.t99 168.701
R21330 commonsourceibias.n617 commonsourceibias.t72 168.701
R21331 commonsourceibias.n623 commonsourceibias.t142 168.701
R21332 commonsourceibias.n625 commonsourceibias.t100 168.701
R21333 commonsourceibias.n632 commonsourceibias.t65 168.701
R21334 commonsourceibias.n638 commonsourceibias.t143 168.701
R21335 commonsourceibias.n640 commonsourceibias.t154 168.701
R21336 commonsourceibias.n647 commonsourceibias.t66 168.701
R21337 commonsourceibias.n653 commonsourceibias.t144 168.701
R21338 commonsourceibias.n36 commonsourceibias.n33 161.3
R21339 commonsourceibias.n38 commonsourceibias.n37 161.3
R21340 commonsourceibias.n39 commonsourceibias.n32 161.3
R21341 commonsourceibias.n42 commonsourceibias.n41 161.3
R21342 commonsourceibias.n43 commonsourceibias.n31 161.3
R21343 commonsourceibias.n45 commonsourceibias.n44 161.3
R21344 commonsourceibias.n47 commonsourceibias.n30 161.3
R21345 commonsourceibias.n49 commonsourceibias.n48 161.3
R21346 commonsourceibias.n51 commonsourceibias.n50 161.3
R21347 commonsourceibias.n52 commonsourceibias.n28 161.3
R21348 commonsourceibias.n54 commonsourceibias.n53 161.3
R21349 commonsourceibias.n56 commonsourceibias.n55 161.3
R21350 commonsourceibias.n57 commonsourceibias.n26 161.3
R21351 commonsourceibias.n59 commonsourceibias.n58 161.3
R21352 commonsourceibias.n61 commonsourceibias.n60 161.3
R21353 commonsourceibias.n62 commonsourceibias.n24 161.3
R21354 commonsourceibias.n65 commonsourceibias.n64 161.3
R21355 commonsourceibias.n66 commonsourceibias.n23 161.3
R21356 commonsourceibias.n68 commonsourceibias.n67 161.3
R21357 commonsourceibias.n70 commonsourceibias.n21 161.3
R21358 commonsourceibias.n72 commonsourceibias.n71 161.3
R21359 commonsourceibias.n73 commonsourceibias.n20 161.3
R21360 commonsourceibias.n75 commonsourceibias.n74 161.3
R21361 commonsourceibias.n76 commonsourceibias.n19 161.3
R21362 commonsourceibias.n79 commonsourceibias.n78 161.3
R21363 commonsourceibias.n80 commonsourceibias.n18 161.3
R21364 commonsourceibias.n82 commonsourceibias.n81 161.3
R21365 commonsourceibias.n84 commonsourceibias.n16 161.3
R21366 commonsourceibias.n86 commonsourceibias.n85 161.3
R21367 commonsourceibias.n87 commonsourceibias.n15 161.3
R21368 commonsourceibias.n89 commonsourceibias.n88 161.3
R21369 commonsourceibias.n90 commonsourceibias.n14 161.3
R21370 commonsourceibias.n93 commonsourceibias.n92 161.3
R21371 commonsourceibias.n94 commonsourceibias.n13 161.3
R21372 commonsourceibias.n96 commonsourceibias.n95 161.3
R21373 commonsourceibias.n98 commonsourceibias.n12 161.3
R21374 commonsourceibias.n129 commonsourceibias.n126 161.3
R21375 commonsourceibias.n131 commonsourceibias.n130 161.3
R21376 commonsourceibias.n132 commonsourceibias.n125 161.3
R21377 commonsourceibias.n135 commonsourceibias.n134 161.3
R21378 commonsourceibias.n136 commonsourceibias.n124 161.3
R21379 commonsourceibias.n138 commonsourceibias.n137 161.3
R21380 commonsourceibias.n140 commonsourceibias.n123 161.3
R21381 commonsourceibias.n142 commonsourceibias.n141 161.3
R21382 commonsourceibias.n144 commonsourceibias.n143 161.3
R21383 commonsourceibias.n145 commonsourceibias.n121 161.3
R21384 commonsourceibias.n147 commonsourceibias.n146 161.3
R21385 commonsourceibias.n149 commonsourceibias.n148 161.3
R21386 commonsourceibias.n150 commonsourceibias.n119 161.3
R21387 commonsourceibias.n152 commonsourceibias.n151 161.3
R21388 commonsourceibias.n154 commonsourceibias.n153 161.3
R21389 commonsourceibias.n155 commonsourceibias.n117 161.3
R21390 commonsourceibias.n158 commonsourceibias.n157 161.3
R21391 commonsourceibias.n159 commonsourceibias.n11 161.3
R21392 commonsourceibias.n161 commonsourceibias.n160 161.3
R21393 commonsourceibias.n163 commonsourceibias.n9 161.3
R21394 commonsourceibias.n165 commonsourceibias.n164 161.3
R21395 commonsourceibias.n166 commonsourceibias.n8 161.3
R21396 commonsourceibias.n168 commonsourceibias.n167 161.3
R21397 commonsourceibias.n169 commonsourceibias.n7 161.3
R21398 commonsourceibias.n172 commonsourceibias.n171 161.3
R21399 commonsourceibias.n173 commonsourceibias.n6 161.3
R21400 commonsourceibias.n175 commonsourceibias.n174 161.3
R21401 commonsourceibias.n177 commonsourceibias.n4 161.3
R21402 commonsourceibias.n179 commonsourceibias.n178 161.3
R21403 commonsourceibias.n180 commonsourceibias.n3 161.3
R21404 commonsourceibias.n182 commonsourceibias.n181 161.3
R21405 commonsourceibias.n183 commonsourceibias.n2 161.3
R21406 commonsourceibias.n186 commonsourceibias.n185 161.3
R21407 commonsourceibias.n187 commonsourceibias.n1 161.3
R21408 commonsourceibias.n189 commonsourceibias.n188 161.3
R21409 commonsourceibias.n191 commonsourceibias.n0 161.3
R21410 commonsourceibias.n370 commonsourceibias.n284 161.3
R21411 commonsourceibias.n368 commonsourceibias.n367 161.3
R21412 commonsourceibias.n366 commonsourceibias.n285 161.3
R21413 commonsourceibias.n365 commonsourceibias.n364 161.3
R21414 commonsourceibias.n362 commonsourceibias.n286 161.3
R21415 commonsourceibias.n361 commonsourceibias.n360 161.3
R21416 commonsourceibias.n359 commonsourceibias.n287 161.3
R21417 commonsourceibias.n358 commonsourceibias.n357 161.3
R21418 commonsourceibias.n356 commonsourceibias.n288 161.3
R21419 commonsourceibias.n354 commonsourceibias.n353 161.3
R21420 commonsourceibias.n352 commonsourceibias.n290 161.3
R21421 commonsourceibias.n351 commonsourceibias.n350 161.3
R21422 commonsourceibias.n348 commonsourceibias.n291 161.3
R21423 commonsourceibias.n347 commonsourceibias.n346 161.3
R21424 commonsourceibias.n345 commonsourceibias.n292 161.3
R21425 commonsourceibias.n344 commonsourceibias.n343 161.3
R21426 commonsourceibias.n342 commonsourceibias.n293 161.3
R21427 commonsourceibias.n340 commonsourceibias.n339 161.3
R21428 commonsourceibias.n338 commonsourceibias.n295 161.3
R21429 commonsourceibias.n337 commonsourceibias.n336 161.3
R21430 commonsourceibias.n334 commonsourceibias.n296 161.3
R21431 commonsourceibias.n333 commonsourceibias.n332 161.3
R21432 commonsourceibias.n331 commonsourceibias.n330 161.3
R21433 commonsourceibias.n329 commonsourceibias.n298 161.3
R21434 commonsourceibias.n328 commonsourceibias.n327 161.3
R21435 commonsourceibias.n326 commonsourceibias.n325 161.3
R21436 commonsourceibias.n324 commonsourceibias.n300 161.3
R21437 commonsourceibias.n323 commonsourceibias.n322 161.3
R21438 commonsourceibias.n321 commonsourceibias.n320 161.3
R21439 commonsourceibias.n319 commonsourceibias.n302 161.3
R21440 commonsourceibias.n317 commonsourceibias.n316 161.3
R21441 commonsourceibias.n315 commonsourceibias.n303 161.3
R21442 commonsourceibias.n314 commonsourceibias.n313 161.3
R21443 commonsourceibias.n311 commonsourceibias.n304 161.3
R21444 commonsourceibias.n310 commonsourceibias.n309 161.3
R21445 commonsourceibias.n308 commonsourceibias.n305 161.3
R21446 commonsourceibias.n218 commonsourceibias.n215 161.3
R21447 commonsourceibias.n220 commonsourceibias.n219 161.3
R21448 commonsourceibias.n221 commonsourceibias.n214 161.3
R21449 commonsourceibias.n224 commonsourceibias.n223 161.3
R21450 commonsourceibias.n225 commonsourceibias.n213 161.3
R21451 commonsourceibias.n227 commonsourceibias.n226 161.3
R21452 commonsourceibias.n229 commonsourceibias.n212 161.3
R21453 commonsourceibias.n231 commonsourceibias.n230 161.3
R21454 commonsourceibias.n233 commonsourceibias.n232 161.3
R21455 commonsourceibias.n234 commonsourceibias.n210 161.3
R21456 commonsourceibias.n236 commonsourceibias.n235 161.3
R21457 commonsourceibias.n238 commonsourceibias.n237 161.3
R21458 commonsourceibias.n239 commonsourceibias.n208 161.3
R21459 commonsourceibias.n241 commonsourceibias.n240 161.3
R21460 commonsourceibias.n243 commonsourceibias.n242 161.3
R21461 commonsourceibias.n244 commonsourceibias.n206 161.3
R21462 commonsourceibias.n247 commonsourceibias.n246 161.3
R21463 commonsourceibias.n248 commonsourceibias.n205 161.3
R21464 commonsourceibias.n250 commonsourceibias.n249 161.3
R21465 commonsourceibias.n252 commonsourceibias.n203 161.3
R21466 commonsourceibias.n254 commonsourceibias.n253 161.3
R21467 commonsourceibias.n255 commonsourceibias.n202 161.3
R21468 commonsourceibias.n257 commonsourceibias.n256 161.3
R21469 commonsourceibias.n258 commonsourceibias.n201 161.3
R21470 commonsourceibias.n261 commonsourceibias.n260 161.3
R21471 commonsourceibias.n262 commonsourceibias.n200 161.3
R21472 commonsourceibias.n264 commonsourceibias.n263 161.3
R21473 commonsourceibias.n266 commonsourceibias.n198 161.3
R21474 commonsourceibias.n268 commonsourceibias.n267 161.3
R21475 commonsourceibias.n269 commonsourceibias.n197 161.3
R21476 commonsourceibias.n271 commonsourceibias.n270 161.3
R21477 commonsourceibias.n272 commonsourceibias.n196 161.3
R21478 commonsourceibias.n275 commonsourceibias.n274 161.3
R21479 commonsourceibias.n276 commonsourceibias.n195 161.3
R21480 commonsourceibias.n278 commonsourceibias.n277 161.3
R21481 commonsourceibias.n280 commonsourceibias.n194 161.3
R21482 commonsourceibias.n519 commonsourceibias.n433 161.3
R21483 commonsourceibias.n517 commonsourceibias.n516 161.3
R21484 commonsourceibias.n515 commonsourceibias.n434 161.3
R21485 commonsourceibias.n514 commonsourceibias.n513 161.3
R21486 commonsourceibias.n511 commonsourceibias.n435 161.3
R21487 commonsourceibias.n510 commonsourceibias.n509 161.3
R21488 commonsourceibias.n508 commonsourceibias.n436 161.3
R21489 commonsourceibias.n507 commonsourceibias.n506 161.3
R21490 commonsourceibias.n504 commonsourceibias.n437 161.3
R21491 commonsourceibias.n502 commonsourceibias.n501 161.3
R21492 commonsourceibias.n500 commonsourceibias.n438 161.3
R21493 commonsourceibias.n499 commonsourceibias.n498 161.3
R21494 commonsourceibias.n496 commonsourceibias.n439 161.3
R21495 commonsourceibias.n495 commonsourceibias.n494 161.3
R21496 commonsourceibias.n493 commonsourceibias.n440 161.3
R21497 commonsourceibias.n492 commonsourceibias.n491 161.3
R21498 commonsourceibias.n489 commonsourceibias.n441 161.3
R21499 commonsourceibias.n487 commonsourceibias.n486 161.3
R21500 commonsourceibias.n485 commonsourceibias.n442 161.3
R21501 commonsourceibias.n484 commonsourceibias.n483 161.3
R21502 commonsourceibias.n481 commonsourceibias.n443 161.3
R21503 commonsourceibias.n480 commonsourceibias.n479 161.3
R21504 commonsourceibias.n478 commonsourceibias.n477 161.3
R21505 commonsourceibias.n476 commonsourceibias.n445 161.3
R21506 commonsourceibias.n475 commonsourceibias.n474 161.3
R21507 commonsourceibias.n473 commonsourceibias.n472 161.3
R21508 commonsourceibias.n471 commonsourceibias.n447 161.3
R21509 commonsourceibias.n470 commonsourceibias.n469 161.3
R21510 commonsourceibias.n468 commonsourceibias.n467 161.3
R21511 commonsourceibias.n466 commonsourceibias.n449 161.3
R21512 commonsourceibias.n464 commonsourceibias.n463 161.3
R21513 commonsourceibias.n462 commonsourceibias.n450 161.3
R21514 commonsourceibias.n461 commonsourceibias.n460 161.3
R21515 commonsourceibias.n458 commonsourceibias.n451 161.3
R21516 commonsourceibias.n457 commonsourceibias.n456 161.3
R21517 commonsourceibias.n455 commonsourceibias.n452 161.3
R21518 commonsourceibias.n425 commonsourceibias.n424 161.3
R21519 commonsourceibias.n422 commonsourceibias.n384 161.3
R21520 commonsourceibias.n421 commonsourceibias.n420 161.3
R21521 commonsourceibias.n419 commonsourceibias.n418 161.3
R21522 commonsourceibias.n417 commonsourceibias.n386 161.3
R21523 commonsourceibias.n416 commonsourceibias.n415 161.3
R21524 commonsourceibias.n414 commonsourceibias.n413 161.3
R21525 commonsourceibias.n412 commonsourceibias.n388 161.3
R21526 commonsourceibias.n411 commonsourceibias.n410 161.3
R21527 commonsourceibias.n409 commonsourceibias.n408 161.3
R21528 commonsourceibias.n407 commonsourceibias.n390 161.3
R21529 commonsourceibias.n405 commonsourceibias.n404 161.3
R21530 commonsourceibias.n403 commonsourceibias.n391 161.3
R21531 commonsourceibias.n402 commonsourceibias.n401 161.3
R21532 commonsourceibias.n399 commonsourceibias.n392 161.3
R21533 commonsourceibias.n398 commonsourceibias.n397 161.3
R21534 commonsourceibias.n396 commonsourceibias.n393 161.3
R21535 commonsourceibias.n531 commonsourceibias.n383 161.3
R21536 commonsourceibias.n565 commonsourceibias.n374 161.3
R21537 commonsourceibias.n563 commonsourceibias.n562 161.3
R21538 commonsourceibias.n561 commonsourceibias.n375 161.3
R21539 commonsourceibias.n560 commonsourceibias.n559 161.3
R21540 commonsourceibias.n557 commonsourceibias.n376 161.3
R21541 commonsourceibias.n556 commonsourceibias.n555 161.3
R21542 commonsourceibias.n554 commonsourceibias.n377 161.3
R21543 commonsourceibias.n553 commonsourceibias.n552 161.3
R21544 commonsourceibias.n550 commonsourceibias.n378 161.3
R21545 commonsourceibias.n548 commonsourceibias.n547 161.3
R21546 commonsourceibias.n546 commonsourceibias.n379 161.3
R21547 commonsourceibias.n545 commonsourceibias.n544 161.3
R21548 commonsourceibias.n542 commonsourceibias.n380 161.3
R21549 commonsourceibias.n541 commonsourceibias.n540 161.3
R21550 commonsourceibias.n539 commonsourceibias.n381 161.3
R21551 commonsourceibias.n538 commonsourceibias.n537 161.3
R21552 commonsourceibias.n535 commonsourceibias.n382 161.3
R21553 commonsourceibias.n533 commonsourceibias.n532 161.3
R21554 commonsourceibias.n744 commonsourceibias.n658 161.3
R21555 commonsourceibias.n742 commonsourceibias.n741 161.3
R21556 commonsourceibias.n740 commonsourceibias.n659 161.3
R21557 commonsourceibias.n739 commonsourceibias.n738 161.3
R21558 commonsourceibias.n736 commonsourceibias.n660 161.3
R21559 commonsourceibias.n735 commonsourceibias.n734 161.3
R21560 commonsourceibias.n733 commonsourceibias.n661 161.3
R21561 commonsourceibias.n732 commonsourceibias.n731 161.3
R21562 commonsourceibias.n729 commonsourceibias.n662 161.3
R21563 commonsourceibias.n727 commonsourceibias.n726 161.3
R21564 commonsourceibias.n725 commonsourceibias.n663 161.3
R21565 commonsourceibias.n724 commonsourceibias.n723 161.3
R21566 commonsourceibias.n721 commonsourceibias.n664 161.3
R21567 commonsourceibias.n720 commonsourceibias.n719 161.3
R21568 commonsourceibias.n718 commonsourceibias.n665 161.3
R21569 commonsourceibias.n717 commonsourceibias.n716 161.3
R21570 commonsourceibias.n714 commonsourceibias.n666 161.3
R21571 commonsourceibias.n712 commonsourceibias.n711 161.3
R21572 commonsourceibias.n710 commonsourceibias.n667 161.3
R21573 commonsourceibias.n709 commonsourceibias.n708 161.3
R21574 commonsourceibias.n706 commonsourceibias.n668 161.3
R21575 commonsourceibias.n705 commonsourceibias.n704 161.3
R21576 commonsourceibias.n703 commonsourceibias.n702 161.3
R21577 commonsourceibias.n701 commonsourceibias.n670 161.3
R21578 commonsourceibias.n700 commonsourceibias.n699 161.3
R21579 commonsourceibias.n698 commonsourceibias.n697 161.3
R21580 commonsourceibias.n696 commonsourceibias.n672 161.3
R21581 commonsourceibias.n695 commonsourceibias.n694 161.3
R21582 commonsourceibias.n693 commonsourceibias.n692 161.3
R21583 commonsourceibias.n691 commonsourceibias.n674 161.3
R21584 commonsourceibias.n689 commonsourceibias.n688 161.3
R21585 commonsourceibias.n687 commonsourceibias.n675 161.3
R21586 commonsourceibias.n686 commonsourceibias.n685 161.3
R21587 commonsourceibias.n683 commonsourceibias.n676 161.3
R21588 commonsourceibias.n682 commonsourceibias.n681 161.3
R21589 commonsourceibias.n680 commonsourceibias.n677 161.3
R21590 commonsourceibias.n654 commonsourceibias.n568 161.3
R21591 commonsourceibias.n652 commonsourceibias.n651 161.3
R21592 commonsourceibias.n650 commonsourceibias.n569 161.3
R21593 commonsourceibias.n649 commonsourceibias.n648 161.3
R21594 commonsourceibias.n646 commonsourceibias.n570 161.3
R21595 commonsourceibias.n645 commonsourceibias.n644 161.3
R21596 commonsourceibias.n643 commonsourceibias.n571 161.3
R21597 commonsourceibias.n642 commonsourceibias.n641 161.3
R21598 commonsourceibias.n639 commonsourceibias.n572 161.3
R21599 commonsourceibias.n637 commonsourceibias.n636 161.3
R21600 commonsourceibias.n635 commonsourceibias.n573 161.3
R21601 commonsourceibias.n634 commonsourceibias.n633 161.3
R21602 commonsourceibias.n631 commonsourceibias.n574 161.3
R21603 commonsourceibias.n630 commonsourceibias.n629 161.3
R21604 commonsourceibias.n628 commonsourceibias.n575 161.3
R21605 commonsourceibias.n627 commonsourceibias.n626 161.3
R21606 commonsourceibias.n624 commonsourceibias.n576 161.3
R21607 commonsourceibias.n622 commonsourceibias.n621 161.3
R21608 commonsourceibias.n620 commonsourceibias.n577 161.3
R21609 commonsourceibias.n619 commonsourceibias.n618 161.3
R21610 commonsourceibias.n616 commonsourceibias.n578 161.3
R21611 commonsourceibias.n615 commonsourceibias.n614 161.3
R21612 commonsourceibias.n613 commonsourceibias.n612 161.3
R21613 commonsourceibias.n611 commonsourceibias.n580 161.3
R21614 commonsourceibias.n610 commonsourceibias.n609 161.3
R21615 commonsourceibias.n608 commonsourceibias.n607 161.3
R21616 commonsourceibias.n606 commonsourceibias.n582 161.3
R21617 commonsourceibias.n605 commonsourceibias.n604 161.3
R21618 commonsourceibias.n603 commonsourceibias.n602 161.3
R21619 commonsourceibias.n601 commonsourceibias.n584 161.3
R21620 commonsourceibias.n599 commonsourceibias.n598 161.3
R21621 commonsourceibias.n597 commonsourceibias.n585 161.3
R21622 commonsourceibias.n596 commonsourceibias.n595 161.3
R21623 commonsourceibias.n593 commonsourceibias.n586 161.3
R21624 commonsourceibias.n592 commonsourceibias.n591 161.3
R21625 commonsourceibias.n590 commonsourceibias.n587 161.3
R21626 commonsourceibias.n111 commonsourceibias.n109 81.5057
R21627 commonsourceibias.n428 commonsourceibias.n426 81.5057
R21628 commonsourceibias.n111 commonsourceibias.n110 80.9324
R21629 commonsourceibias.n113 commonsourceibias.n112 80.9324
R21630 commonsourceibias.n115 commonsourceibias.n114 80.9324
R21631 commonsourceibias.n108 commonsourceibias.n107 80.9324
R21632 commonsourceibias.n106 commonsourceibias.n105 80.9324
R21633 commonsourceibias.n104 commonsourceibias.n103 80.9324
R21634 commonsourceibias.n102 commonsourceibias.n101 80.9324
R21635 commonsourceibias.n523 commonsourceibias.n522 80.9324
R21636 commonsourceibias.n525 commonsourceibias.n524 80.9324
R21637 commonsourceibias.n527 commonsourceibias.n526 80.9324
R21638 commonsourceibias.n529 commonsourceibias.n528 80.9324
R21639 commonsourceibias.n432 commonsourceibias.n431 80.9324
R21640 commonsourceibias.n430 commonsourceibias.n429 80.9324
R21641 commonsourceibias.n428 commonsourceibias.n427 80.9324
R21642 commonsourceibias.n100 commonsourceibias.n99 80.6037
R21643 commonsourceibias.n193 commonsourceibias.n192 80.6037
R21644 commonsourceibias.n372 commonsourceibias.n371 80.6037
R21645 commonsourceibias.n282 commonsourceibias.n281 80.6037
R21646 commonsourceibias.n521 commonsourceibias.n520 80.6037
R21647 commonsourceibias.n567 commonsourceibias.n566 80.6037
R21648 commonsourceibias.n746 commonsourceibias.n745 80.6037
R21649 commonsourceibias.n656 commonsourceibias.n655 80.6037
R21650 commonsourceibias.n85 commonsourceibias.n84 56.5617
R21651 commonsourceibias.n71 commonsourceibias.n70 56.5617
R21652 commonsourceibias.n62 commonsourceibias.n61 56.5617
R21653 commonsourceibias.n48 commonsourceibias.n47 56.5617
R21654 commonsourceibias.n178 commonsourceibias.n177 56.5617
R21655 commonsourceibias.n164 commonsourceibias.n163 56.5617
R21656 commonsourceibias.n155 commonsourceibias.n154 56.5617
R21657 commonsourceibias.n141 commonsourceibias.n140 56.5617
R21658 commonsourceibias.n320 commonsourceibias.n319 56.5617
R21659 commonsourceibias.n334 commonsourceibias.n333 56.5617
R21660 commonsourceibias.n343 commonsourceibias.n342 56.5617
R21661 commonsourceibias.n357 commonsourceibias.n356 56.5617
R21662 commonsourceibias.n267 commonsourceibias.n266 56.5617
R21663 commonsourceibias.n253 commonsourceibias.n252 56.5617
R21664 commonsourceibias.n244 commonsourceibias.n243 56.5617
R21665 commonsourceibias.n230 commonsourceibias.n229 56.5617
R21666 commonsourceibias.n467 commonsourceibias.n466 56.5617
R21667 commonsourceibias.n481 commonsourceibias.n480 56.5617
R21668 commonsourceibias.n491 commonsourceibias.n489 56.5617
R21669 commonsourceibias.n506 commonsourceibias.n504 56.5617
R21670 commonsourceibias.n552 commonsourceibias.n550 56.5617
R21671 commonsourceibias.n537 commonsourceibias.n535 56.5617
R21672 commonsourceibias.n408 commonsourceibias.n407 56.5617
R21673 commonsourceibias.n422 commonsourceibias.n421 56.5617
R21674 commonsourceibias.n692 commonsourceibias.n691 56.5617
R21675 commonsourceibias.n706 commonsourceibias.n705 56.5617
R21676 commonsourceibias.n716 commonsourceibias.n714 56.5617
R21677 commonsourceibias.n731 commonsourceibias.n729 56.5617
R21678 commonsourceibias.n602 commonsourceibias.n601 56.5617
R21679 commonsourceibias.n616 commonsourceibias.n615 56.5617
R21680 commonsourceibias.n626 commonsourceibias.n624 56.5617
R21681 commonsourceibias.n641 commonsourceibias.n639 56.5617
R21682 commonsourceibias.n76 commonsourceibias.n75 56.0773
R21683 commonsourceibias.n57 commonsourceibias.n56 56.0773
R21684 commonsourceibias.n169 commonsourceibias.n168 56.0773
R21685 commonsourceibias.n150 commonsourceibias.n149 56.0773
R21686 commonsourceibias.n329 commonsourceibias.n328 56.0773
R21687 commonsourceibias.n348 commonsourceibias.n347 56.0773
R21688 commonsourceibias.n258 commonsourceibias.n257 56.0773
R21689 commonsourceibias.n239 commonsourceibias.n238 56.0773
R21690 commonsourceibias.n476 commonsourceibias.n475 56.0773
R21691 commonsourceibias.n496 commonsourceibias.n495 56.0773
R21692 commonsourceibias.n542 commonsourceibias.n541 56.0773
R21693 commonsourceibias.n417 commonsourceibias.n416 56.0773
R21694 commonsourceibias.n701 commonsourceibias.n700 56.0773
R21695 commonsourceibias.n721 commonsourceibias.n720 56.0773
R21696 commonsourceibias.n611 commonsourceibias.n610 56.0773
R21697 commonsourceibias.n631 commonsourceibias.n630 56.0773
R21698 commonsourceibias.n99 commonsourceibias.n98 55.3321
R21699 commonsourceibias.n192 commonsourceibias.n191 55.3321
R21700 commonsourceibias.n371 commonsourceibias.n370 55.3321
R21701 commonsourceibias.n281 commonsourceibias.n280 55.3321
R21702 commonsourceibias.n520 commonsourceibias.n519 55.3321
R21703 commonsourceibias.n566 commonsourceibias.n565 55.3321
R21704 commonsourceibias.n745 commonsourceibias.n744 55.3321
R21705 commonsourceibias.n655 commonsourceibias.n654 55.3321
R21706 commonsourceibias.n90 commonsourceibias.n89 55.1086
R21707 commonsourceibias.n41 commonsourceibias.n31 55.1086
R21708 commonsourceibias.n183 commonsourceibias.n182 55.1086
R21709 commonsourceibias.n134 commonsourceibias.n124 55.1086
R21710 commonsourceibias.n313 commonsourceibias.n303 55.1086
R21711 commonsourceibias.n362 commonsourceibias.n361 55.1086
R21712 commonsourceibias.n272 commonsourceibias.n271 55.1086
R21713 commonsourceibias.n223 commonsourceibias.n213 55.1086
R21714 commonsourceibias.n460 commonsourceibias.n450 55.1086
R21715 commonsourceibias.n511 commonsourceibias.n510 55.1086
R21716 commonsourceibias.n557 commonsourceibias.n556 55.1086
R21717 commonsourceibias.n401 commonsourceibias.n391 55.1086
R21718 commonsourceibias.n685 commonsourceibias.n675 55.1086
R21719 commonsourceibias.n736 commonsourceibias.n735 55.1086
R21720 commonsourceibias.n595 commonsourceibias.n585 55.1086
R21721 commonsourceibias.n646 commonsourceibias.n645 55.1086
R21722 commonsourceibias.n35 commonsourceibias.n34 47.4592
R21723 commonsourceibias.n128 commonsourceibias.n127 47.4592
R21724 commonsourceibias.n307 commonsourceibias.n306 47.4592
R21725 commonsourceibias.n217 commonsourceibias.n216 47.4592
R21726 commonsourceibias.n454 commonsourceibias.n453 47.4592
R21727 commonsourceibias.n395 commonsourceibias.n394 47.4592
R21728 commonsourceibias.n679 commonsourceibias.n678 47.4592
R21729 commonsourceibias.n589 commonsourceibias.n588 47.4592
R21730 commonsourceibias.n308 commonsourceibias.n307 44.0436
R21731 commonsourceibias.n455 commonsourceibias.n454 44.0436
R21732 commonsourceibias.n396 commonsourceibias.n395 44.0436
R21733 commonsourceibias.n680 commonsourceibias.n679 44.0436
R21734 commonsourceibias.n590 commonsourceibias.n589 44.0436
R21735 commonsourceibias.n36 commonsourceibias.n35 44.0436
R21736 commonsourceibias.n129 commonsourceibias.n128 44.0436
R21737 commonsourceibias.n218 commonsourceibias.n217 44.0436
R21738 commonsourceibias.n92 commonsourceibias.n13 42.5146
R21739 commonsourceibias.n39 commonsourceibias.n38 42.5146
R21740 commonsourceibias.n185 commonsourceibias.n1 42.5146
R21741 commonsourceibias.n132 commonsourceibias.n131 42.5146
R21742 commonsourceibias.n311 commonsourceibias.n310 42.5146
R21743 commonsourceibias.n364 commonsourceibias.n285 42.5146
R21744 commonsourceibias.n274 commonsourceibias.n195 42.5146
R21745 commonsourceibias.n221 commonsourceibias.n220 42.5146
R21746 commonsourceibias.n458 commonsourceibias.n457 42.5146
R21747 commonsourceibias.n513 commonsourceibias.n434 42.5146
R21748 commonsourceibias.n559 commonsourceibias.n375 42.5146
R21749 commonsourceibias.n399 commonsourceibias.n398 42.5146
R21750 commonsourceibias.n683 commonsourceibias.n682 42.5146
R21751 commonsourceibias.n738 commonsourceibias.n659 42.5146
R21752 commonsourceibias.n593 commonsourceibias.n592 42.5146
R21753 commonsourceibias.n648 commonsourceibias.n569 42.5146
R21754 commonsourceibias.n78 commonsourceibias.n18 41.5458
R21755 commonsourceibias.n53 commonsourceibias.n52 41.5458
R21756 commonsourceibias.n171 commonsourceibias.n6 41.5458
R21757 commonsourceibias.n146 commonsourceibias.n145 41.5458
R21758 commonsourceibias.n325 commonsourceibias.n324 41.5458
R21759 commonsourceibias.n350 commonsourceibias.n290 41.5458
R21760 commonsourceibias.n260 commonsourceibias.n200 41.5458
R21761 commonsourceibias.n235 commonsourceibias.n234 41.5458
R21762 commonsourceibias.n472 commonsourceibias.n471 41.5458
R21763 commonsourceibias.n498 commonsourceibias.n438 41.5458
R21764 commonsourceibias.n544 commonsourceibias.n379 41.5458
R21765 commonsourceibias.n413 commonsourceibias.n412 41.5458
R21766 commonsourceibias.n697 commonsourceibias.n696 41.5458
R21767 commonsourceibias.n723 commonsourceibias.n663 41.5458
R21768 commonsourceibias.n607 commonsourceibias.n606 41.5458
R21769 commonsourceibias.n633 commonsourceibias.n573 41.5458
R21770 commonsourceibias.n68 commonsourceibias.n23 40.577
R21771 commonsourceibias.n64 commonsourceibias.n23 40.577
R21772 commonsourceibias.n161 commonsourceibias.n11 40.577
R21773 commonsourceibias.n157 commonsourceibias.n11 40.577
R21774 commonsourceibias.n336 commonsourceibias.n295 40.577
R21775 commonsourceibias.n340 commonsourceibias.n295 40.577
R21776 commonsourceibias.n250 commonsourceibias.n205 40.577
R21777 commonsourceibias.n246 commonsourceibias.n205 40.577
R21778 commonsourceibias.n483 commonsourceibias.n442 40.577
R21779 commonsourceibias.n487 commonsourceibias.n442 40.577
R21780 commonsourceibias.n533 commonsourceibias.n383 40.577
R21781 commonsourceibias.n424 commonsourceibias.n383 40.577
R21782 commonsourceibias.n708 commonsourceibias.n667 40.577
R21783 commonsourceibias.n712 commonsourceibias.n667 40.577
R21784 commonsourceibias.n618 commonsourceibias.n577 40.577
R21785 commonsourceibias.n622 commonsourceibias.n577 40.577
R21786 commonsourceibias.n82 commonsourceibias.n18 39.6083
R21787 commonsourceibias.n52 commonsourceibias.n51 39.6083
R21788 commonsourceibias.n175 commonsourceibias.n6 39.6083
R21789 commonsourceibias.n145 commonsourceibias.n144 39.6083
R21790 commonsourceibias.n324 commonsourceibias.n323 39.6083
R21791 commonsourceibias.n354 commonsourceibias.n290 39.6083
R21792 commonsourceibias.n264 commonsourceibias.n200 39.6083
R21793 commonsourceibias.n234 commonsourceibias.n233 39.6083
R21794 commonsourceibias.n471 commonsourceibias.n470 39.6083
R21795 commonsourceibias.n502 commonsourceibias.n438 39.6083
R21796 commonsourceibias.n548 commonsourceibias.n379 39.6083
R21797 commonsourceibias.n412 commonsourceibias.n411 39.6083
R21798 commonsourceibias.n696 commonsourceibias.n695 39.6083
R21799 commonsourceibias.n727 commonsourceibias.n663 39.6083
R21800 commonsourceibias.n606 commonsourceibias.n605 39.6083
R21801 commonsourceibias.n637 commonsourceibias.n573 39.6083
R21802 commonsourceibias.n96 commonsourceibias.n13 38.6395
R21803 commonsourceibias.n38 commonsourceibias.n33 38.6395
R21804 commonsourceibias.n189 commonsourceibias.n1 38.6395
R21805 commonsourceibias.n131 commonsourceibias.n126 38.6395
R21806 commonsourceibias.n310 commonsourceibias.n305 38.6395
R21807 commonsourceibias.n368 commonsourceibias.n285 38.6395
R21808 commonsourceibias.n278 commonsourceibias.n195 38.6395
R21809 commonsourceibias.n220 commonsourceibias.n215 38.6395
R21810 commonsourceibias.n457 commonsourceibias.n452 38.6395
R21811 commonsourceibias.n517 commonsourceibias.n434 38.6395
R21812 commonsourceibias.n563 commonsourceibias.n375 38.6395
R21813 commonsourceibias.n398 commonsourceibias.n393 38.6395
R21814 commonsourceibias.n682 commonsourceibias.n677 38.6395
R21815 commonsourceibias.n742 commonsourceibias.n659 38.6395
R21816 commonsourceibias.n592 commonsourceibias.n587 38.6395
R21817 commonsourceibias.n652 commonsourceibias.n569 38.6395
R21818 commonsourceibias.n89 commonsourceibias.n15 26.0455
R21819 commonsourceibias.n45 commonsourceibias.n31 26.0455
R21820 commonsourceibias.n182 commonsourceibias.n3 26.0455
R21821 commonsourceibias.n138 commonsourceibias.n124 26.0455
R21822 commonsourceibias.n317 commonsourceibias.n303 26.0455
R21823 commonsourceibias.n361 commonsourceibias.n287 26.0455
R21824 commonsourceibias.n271 commonsourceibias.n197 26.0455
R21825 commonsourceibias.n227 commonsourceibias.n213 26.0455
R21826 commonsourceibias.n464 commonsourceibias.n450 26.0455
R21827 commonsourceibias.n510 commonsourceibias.n436 26.0455
R21828 commonsourceibias.n556 commonsourceibias.n377 26.0455
R21829 commonsourceibias.n405 commonsourceibias.n391 26.0455
R21830 commonsourceibias.n689 commonsourceibias.n675 26.0455
R21831 commonsourceibias.n735 commonsourceibias.n661 26.0455
R21832 commonsourceibias.n599 commonsourceibias.n585 26.0455
R21833 commonsourceibias.n645 commonsourceibias.n571 26.0455
R21834 commonsourceibias.n75 commonsourceibias.n20 25.0767
R21835 commonsourceibias.n58 commonsourceibias.n57 25.0767
R21836 commonsourceibias.n168 commonsourceibias.n8 25.0767
R21837 commonsourceibias.n151 commonsourceibias.n150 25.0767
R21838 commonsourceibias.n330 commonsourceibias.n329 25.0767
R21839 commonsourceibias.n347 commonsourceibias.n292 25.0767
R21840 commonsourceibias.n257 commonsourceibias.n202 25.0767
R21841 commonsourceibias.n240 commonsourceibias.n239 25.0767
R21842 commonsourceibias.n477 commonsourceibias.n476 25.0767
R21843 commonsourceibias.n495 commonsourceibias.n440 25.0767
R21844 commonsourceibias.n541 commonsourceibias.n381 25.0767
R21845 commonsourceibias.n418 commonsourceibias.n417 25.0767
R21846 commonsourceibias.n702 commonsourceibias.n701 25.0767
R21847 commonsourceibias.n720 commonsourceibias.n665 25.0767
R21848 commonsourceibias.n612 commonsourceibias.n611 25.0767
R21849 commonsourceibias.n630 commonsourceibias.n575 25.0767
R21850 commonsourceibias.n71 commonsourceibias.n22 24.3464
R21851 commonsourceibias.n61 commonsourceibias.n25 24.3464
R21852 commonsourceibias.n164 commonsourceibias.n10 24.3464
R21853 commonsourceibias.n154 commonsourceibias.n118 24.3464
R21854 commonsourceibias.n333 commonsourceibias.n297 24.3464
R21855 commonsourceibias.n343 commonsourceibias.n294 24.3464
R21856 commonsourceibias.n253 commonsourceibias.n204 24.3464
R21857 commonsourceibias.n243 commonsourceibias.n207 24.3464
R21858 commonsourceibias.n480 commonsourceibias.n444 24.3464
R21859 commonsourceibias.n491 commonsourceibias.n490 24.3464
R21860 commonsourceibias.n537 commonsourceibias.n536 24.3464
R21861 commonsourceibias.n421 commonsourceibias.n385 24.3464
R21862 commonsourceibias.n705 commonsourceibias.n669 24.3464
R21863 commonsourceibias.n716 commonsourceibias.n715 24.3464
R21864 commonsourceibias.n615 commonsourceibias.n579 24.3464
R21865 commonsourceibias.n626 commonsourceibias.n625 24.3464
R21866 commonsourceibias.n85 commonsourceibias.n17 23.8546
R21867 commonsourceibias.n47 commonsourceibias.n46 23.8546
R21868 commonsourceibias.n178 commonsourceibias.n5 23.8546
R21869 commonsourceibias.n140 commonsourceibias.n139 23.8546
R21870 commonsourceibias.n319 commonsourceibias.n318 23.8546
R21871 commonsourceibias.n357 commonsourceibias.n289 23.8546
R21872 commonsourceibias.n267 commonsourceibias.n199 23.8546
R21873 commonsourceibias.n229 commonsourceibias.n228 23.8546
R21874 commonsourceibias.n466 commonsourceibias.n465 23.8546
R21875 commonsourceibias.n506 commonsourceibias.n505 23.8546
R21876 commonsourceibias.n552 commonsourceibias.n551 23.8546
R21877 commonsourceibias.n407 commonsourceibias.n406 23.8546
R21878 commonsourceibias.n691 commonsourceibias.n690 23.8546
R21879 commonsourceibias.n731 commonsourceibias.n730 23.8546
R21880 commonsourceibias.n601 commonsourceibias.n600 23.8546
R21881 commonsourceibias.n641 commonsourceibias.n640 23.8546
R21882 commonsourceibias.n98 commonsourceibias.n97 17.4607
R21883 commonsourceibias.n191 commonsourceibias.n190 17.4607
R21884 commonsourceibias.n370 commonsourceibias.n369 17.4607
R21885 commonsourceibias.n280 commonsourceibias.n279 17.4607
R21886 commonsourceibias.n519 commonsourceibias.n518 17.4607
R21887 commonsourceibias.n565 commonsourceibias.n564 17.4607
R21888 commonsourceibias.n744 commonsourceibias.n743 17.4607
R21889 commonsourceibias.n654 commonsourceibias.n653 17.4607
R21890 commonsourceibias.n84 commonsourceibias.n83 16.9689
R21891 commonsourceibias.n48 commonsourceibias.n29 16.9689
R21892 commonsourceibias.n177 commonsourceibias.n176 16.9689
R21893 commonsourceibias.n141 commonsourceibias.n122 16.9689
R21894 commonsourceibias.n320 commonsourceibias.n301 16.9689
R21895 commonsourceibias.n356 commonsourceibias.n355 16.9689
R21896 commonsourceibias.n266 commonsourceibias.n265 16.9689
R21897 commonsourceibias.n230 commonsourceibias.n211 16.9689
R21898 commonsourceibias.n467 commonsourceibias.n448 16.9689
R21899 commonsourceibias.n504 commonsourceibias.n503 16.9689
R21900 commonsourceibias.n550 commonsourceibias.n549 16.9689
R21901 commonsourceibias.n408 commonsourceibias.n389 16.9689
R21902 commonsourceibias.n692 commonsourceibias.n673 16.9689
R21903 commonsourceibias.n729 commonsourceibias.n728 16.9689
R21904 commonsourceibias.n602 commonsourceibias.n583 16.9689
R21905 commonsourceibias.n639 commonsourceibias.n638 16.9689
R21906 commonsourceibias.n70 commonsourceibias.n69 16.477
R21907 commonsourceibias.n63 commonsourceibias.n62 16.477
R21908 commonsourceibias.n163 commonsourceibias.n162 16.477
R21909 commonsourceibias.n156 commonsourceibias.n155 16.477
R21910 commonsourceibias.n335 commonsourceibias.n334 16.477
R21911 commonsourceibias.n342 commonsourceibias.n341 16.477
R21912 commonsourceibias.n252 commonsourceibias.n251 16.477
R21913 commonsourceibias.n245 commonsourceibias.n244 16.477
R21914 commonsourceibias.n482 commonsourceibias.n481 16.477
R21915 commonsourceibias.n489 commonsourceibias.n488 16.477
R21916 commonsourceibias.n535 commonsourceibias.n534 16.477
R21917 commonsourceibias.n423 commonsourceibias.n422 16.477
R21918 commonsourceibias.n707 commonsourceibias.n706 16.477
R21919 commonsourceibias.n714 commonsourceibias.n713 16.477
R21920 commonsourceibias.n617 commonsourceibias.n616 16.477
R21921 commonsourceibias.n624 commonsourceibias.n623 16.477
R21922 commonsourceibias.n77 commonsourceibias.n76 15.9852
R21923 commonsourceibias.n56 commonsourceibias.n27 15.9852
R21924 commonsourceibias.n170 commonsourceibias.n169 15.9852
R21925 commonsourceibias.n149 commonsourceibias.n120 15.9852
R21926 commonsourceibias.n328 commonsourceibias.n299 15.9852
R21927 commonsourceibias.n349 commonsourceibias.n348 15.9852
R21928 commonsourceibias.n259 commonsourceibias.n258 15.9852
R21929 commonsourceibias.n238 commonsourceibias.n209 15.9852
R21930 commonsourceibias.n475 commonsourceibias.n446 15.9852
R21931 commonsourceibias.n497 commonsourceibias.n496 15.9852
R21932 commonsourceibias.n543 commonsourceibias.n542 15.9852
R21933 commonsourceibias.n416 commonsourceibias.n387 15.9852
R21934 commonsourceibias.n700 commonsourceibias.n671 15.9852
R21935 commonsourceibias.n722 commonsourceibias.n721 15.9852
R21936 commonsourceibias.n610 commonsourceibias.n581 15.9852
R21937 commonsourceibias.n632 commonsourceibias.n631 15.9852
R21938 commonsourceibias.n91 commonsourceibias.n90 15.4934
R21939 commonsourceibias.n41 commonsourceibias.n40 15.4934
R21940 commonsourceibias.n184 commonsourceibias.n183 15.4934
R21941 commonsourceibias.n134 commonsourceibias.n133 15.4934
R21942 commonsourceibias.n313 commonsourceibias.n312 15.4934
R21943 commonsourceibias.n363 commonsourceibias.n362 15.4934
R21944 commonsourceibias.n273 commonsourceibias.n272 15.4934
R21945 commonsourceibias.n223 commonsourceibias.n222 15.4934
R21946 commonsourceibias.n460 commonsourceibias.n459 15.4934
R21947 commonsourceibias.n512 commonsourceibias.n511 15.4934
R21948 commonsourceibias.n558 commonsourceibias.n557 15.4934
R21949 commonsourceibias.n401 commonsourceibias.n400 15.4934
R21950 commonsourceibias.n685 commonsourceibias.n684 15.4934
R21951 commonsourceibias.n737 commonsourceibias.n736 15.4934
R21952 commonsourceibias.n595 commonsourceibias.n594 15.4934
R21953 commonsourceibias.n647 commonsourceibias.n646 15.4934
R21954 commonsourceibias.n102 commonsourceibias.n100 13.2663
R21955 commonsourceibias.n523 commonsourceibias.n521 13.2663
R21956 commonsourceibias.n748 commonsourceibias.n373 10.122
R21957 commonsourceibias.n159 commonsourceibias.n116 9.50363
R21958 commonsourceibias.n531 commonsourceibias.n530 9.50363
R21959 commonsourceibias.n92 commonsourceibias.n91 9.09948
R21960 commonsourceibias.n40 commonsourceibias.n39 9.09948
R21961 commonsourceibias.n185 commonsourceibias.n184 9.09948
R21962 commonsourceibias.n133 commonsourceibias.n132 9.09948
R21963 commonsourceibias.n312 commonsourceibias.n311 9.09948
R21964 commonsourceibias.n364 commonsourceibias.n363 9.09948
R21965 commonsourceibias.n274 commonsourceibias.n273 9.09948
R21966 commonsourceibias.n222 commonsourceibias.n221 9.09948
R21967 commonsourceibias.n459 commonsourceibias.n458 9.09948
R21968 commonsourceibias.n513 commonsourceibias.n512 9.09948
R21969 commonsourceibias.n559 commonsourceibias.n558 9.09948
R21970 commonsourceibias.n400 commonsourceibias.n399 9.09948
R21971 commonsourceibias.n684 commonsourceibias.n683 9.09948
R21972 commonsourceibias.n738 commonsourceibias.n737 9.09948
R21973 commonsourceibias.n594 commonsourceibias.n593 9.09948
R21974 commonsourceibias.n648 commonsourceibias.n647 9.09948
R21975 commonsourceibias.n283 commonsourceibias.n193 8.79451
R21976 commonsourceibias.n657 commonsourceibias.n567 8.79451
R21977 commonsourceibias.n78 commonsourceibias.n77 8.60764
R21978 commonsourceibias.n53 commonsourceibias.n27 8.60764
R21979 commonsourceibias.n171 commonsourceibias.n170 8.60764
R21980 commonsourceibias.n146 commonsourceibias.n120 8.60764
R21981 commonsourceibias.n325 commonsourceibias.n299 8.60764
R21982 commonsourceibias.n350 commonsourceibias.n349 8.60764
R21983 commonsourceibias.n260 commonsourceibias.n259 8.60764
R21984 commonsourceibias.n235 commonsourceibias.n209 8.60764
R21985 commonsourceibias.n472 commonsourceibias.n446 8.60764
R21986 commonsourceibias.n498 commonsourceibias.n497 8.60764
R21987 commonsourceibias.n544 commonsourceibias.n543 8.60764
R21988 commonsourceibias.n413 commonsourceibias.n387 8.60764
R21989 commonsourceibias.n697 commonsourceibias.n671 8.60764
R21990 commonsourceibias.n723 commonsourceibias.n722 8.60764
R21991 commonsourceibias.n607 commonsourceibias.n581 8.60764
R21992 commonsourceibias.n633 commonsourceibias.n632 8.60764
R21993 commonsourceibias.n748 commonsourceibias.n747 8.46921
R21994 commonsourceibias.n69 commonsourceibias.n68 8.11581
R21995 commonsourceibias.n64 commonsourceibias.n63 8.11581
R21996 commonsourceibias.n162 commonsourceibias.n161 8.11581
R21997 commonsourceibias.n157 commonsourceibias.n156 8.11581
R21998 commonsourceibias.n336 commonsourceibias.n335 8.11581
R21999 commonsourceibias.n341 commonsourceibias.n340 8.11581
R22000 commonsourceibias.n251 commonsourceibias.n250 8.11581
R22001 commonsourceibias.n246 commonsourceibias.n245 8.11581
R22002 commonsourceibias.n483 commonsourceibias.n482 8.11581
R22003 commonsourceibias.n488 commonsourceibias.n487 8.11581
R22004 commonsourceibias.n534 commonsourceibias.n533 8.11581
R22005 commonsourceibias.n424 commonsourceibias.n423 8.11581
R22006 commonsourceibias.n708 commonsourceibias.n707 8.11581
R22007 commonsourceibias.n713 commonsourceibias.n712 8.11581
R22008 commonsourceibias.n618 commonsourceibias.n617 8.11581
R22009 commonsourceibias.n623 commonsourceibias.n622 8.11581
R22010 commonsourceibias.n83 commonsourceibias.n82 7.62397
R22011 commonsourceibias.n51 commonsourceibias.n29 7.62397
R22012 commonsourceibias.n176 commonsourceibias.n175 7.62397
R22013 commonsourceibias.n144 commonsourceibias.n122 7.62397
R22014 commonsourceibias.n323 commonsourceibias.n301 7.62397
R22015 commonsourceibias.n355 commonsourceibias.n354 7.62397
R22016 commonsourceibias.n265 commonsourceibias.n264 7.62397
R22017 commonsourceibias.n233 commonsourceibias.n211 7.62397
R22018 commonsourceibias.n470 commonsourceibias.n448 7.62397
R22019 commonsourceibias.n503 commonsourceibias.n502 7.62397
R22020 commonsourceibias.n549 commonsourceibias.n548 7.62397
R22021 commonsourceibias.n411 commonsourceibias.n389 7.62397
R22022 commonsourceibias.n695 commonsourceibias.n673 7.62397
R22023 commonsourceibias.n728 commonsourceibias.n727 7.62397
R22024 commonsourceibias.n605 commonsourceibias.n583 7.62397
R22025 commonsourceibias.n638 commonsourceibias.n637 7.62397
R22026 commonsourceibias.n97 commonsourceibias.n96 7.13213
R22027 commonsourceibias.n34 commonsourceibias.n33 7.13213
R22028 commonsourceibias.n190 commonsourceibias.n189 7.13213
R22029 commonsourceibias.n127 commonsourceibias.n126 7.13213
R22030 commonsourceibias.n306 commonsourceibias.n305 7.13213
R22031 commonsourceibias.n369 commonsourceibias.n368 7.13213
R22032 commonsourceibias.n279 commonsourceibias.n278 7.13213
R22033 commonsourceibias.n216 commonsourceibias.n215 7.13213
R22034 commonsourceibias.n453 commonsourceibias.n452 7.13213
R22035 commonsourceibias.n518 commonsourceibias.n517 7.13213
R22036 commonsourceibias.n564 commonsourceibias.n563 7.13213
R22037 commonsourceibias.n394 commonsourceibias.n393 7.13213
R22038 commonsourceibias.n678 commonsourceibias.n677 7.13213
R22039 commonsourceibias.n743 commonsourceibias.n742 7.13213
R22040 commonsourceibias.n588 commonsourceibias.n587 7.13213
R22041 commonsourceibias.n653 commonsourceibias.n652 7.13213
R22042 commonsourceibias.n373 commonsourceibias.n372 5.06534
R22043 commonsourceibias.n283 commonsourceibias.n282 5.06534
R22044 commonsourceibias.n747 commonsourceibias.n746 5.06534
R22045 commonsourceibias.n657 commonsourceibias.n656 5.06534
R22046 commonsourceibias commonsourceibias.n748 4.04308
R22047 commonsourceibias.n373 commonsourceibias.n283 3.72967
R22048 commonsourceibias.n747 commonsourceibias.n657 3.72967
R22049 commonsourceibias.n109 commonsourceibias.t51 2.82907
R22050 commonsourceibias.n109 commonsourceibias.t1 2.82907
R22051 commonsourceibias.n110 commonsourceibias.t55 2.82907
R22052 commonsourceibias.n110 commonsourceibias.t19 2.82907
R22053 commonsourceibias.n112 commonsourceibias.t25 2.82907
R22054 commonsourceibias.n112 commonsourceibias.t31 2.82907
R22055 commonsourceibias.n114 commonsourceibias.t15 2.82907
R22056 commonsourceibias.n114 commonsourceibias.t45 2.82907
R22057 commonsourceibias.n107 commonsourceibias.t29 2.82907
R22058 commonsourceibias.n107 commonsourceibias.t7 2.82907
R22059 commonsourceibias.n105 commonsourceibias.t59 2.82907
R22060 commonsourceibias.n105 commonsourceibias.t17 2.82907
R22061 commonsourceibias.n103 commonsourceibias.t5 2.82907
R22062 commonsourceibias.n103 commonsourceibias.t11 2.82907
R22063 commonsourceibias.n101 commonsourceibias.t13 2.82907
R22064 commonsourceibias.n101 commonsourceibias.t49 2.82907
R22065 commonsourceibias.n522 commonsourceibias.t61 2.82907
R22066 commonsourceibias.n522 commonsourceibias.t35 2.82907
R22067 commonsourceibias.n524 commonsourceibias.t33 2.82907
R22068 commonsourceibias.n524 commonsourceibias.t21 2.82907
R22069 commonsourceibias.n526 commonsourceibias.t39 2.82907
R22070 commonsourceibias.n526 commonsourceibias.t9 2.82907
R22071 commonsourceibias.n528 commonsourceibias.t27 2.82907
R22072 commonsourceibias.n528 commonsourceibias.t47 2.82907
R22073 commonsourceibias.n431 commonsourceibias.t57 2.82907
R22074 commonsourceibias.n431 commonsourceibias.t37 2.82907
R22075 commonsourceibias.n429 commonsourceibias.t53 2.82907
R22076 commonsourceibias.n429 commonsourceibias.t43 2.82907
R22077 commonsourceibias.n427 commonsourceibias.t41 2.82907
R22078 commonsourceibias.n427 commonsourceibias.t3 2.82907
R22079 commonsourceibias.n426 commonsourceibias.t23 2.82907
R22080 commonsourceibias.n426 commonsourceibias.t63 2.82907
R22081 commonsourceibias.n17 commonsourceibias.n15 0.738255
R22082 commonsourceibias.n46 commonsourceibias.n45 0.738255
R22083 commonsourceibias.n5 commonsourceibias.n3 0.738255
R22084 commonsourceibias.n139 commonsourceibias.n138 0.738255
R22085 commonsourceibias.n318 commonsourceibias.n317 0.738255
R22086 commonsourceibias.n289 commonsourceibias.n287 0.738255
R22087 commonsourceibias.n199 commonsourceibias.n197 0.738255
R22088 commonsourceibias.n228 commonsourceibias.n227 0.738255
R22089 commonsourceibias.n465 commonsourceibias.n464 0.738255
R22090 commonsourceibias.n505 commonsourceibias.n436 0.738255
R22091 commonsourceibias.n551 commonsourceibias.n377 0.738255
R22092 commonsourceibias.n406 commonsourceibias.n405 0.738255
R22093 commonsourceibias.n690 commonsourceibias.n689 0.738255
R22094 commonsourceibias.n730 commonsourceibias.n661 0.738255
R22095 commonsourceibias.n600 commonsourceibias.n599 0.738255
R22096 commonsourceibias.n640 commonsourceibias.n571 0.738255
R22097 commonsourceibias.n104 commonsourceibias.n102 0.573776
R22098 commonsourceibias.n106 commonsourceibias.n104 0.573776
R22099 commonsourceibias.n108 commonsourceibias.n106 0.573776
R22100 commonsourceibias.n115 commonsourceibias.n113 0.573776
R22101 commonsourceibias.n113 commonsourceibias.n111 0.573776
R22102 commonsourceibias.n430 commonsourceibias.n428 0.573776
R22103 commonsourceibias.n432 commonsourceibias.n430 0.573776
R22104 commonsourceibias.n529 commonsourceibias.n527 0.573776
R22105 commonsourceibias.n527 commonsourceibias.n525 0.573776
R22106 commonsourceibias.n525 commonsourceibias.n523 0.573776
R22107 commonsourceibias.n116 commonsourceibias.n108 0.287138
R22108 commonsourceibias.n116 commonsourceibias.n115 0.287138
R22109 commonsourceibias.n530 commonsourceibias.n432 0.287138
R22110 commonsourceibias.n530 commonsourceibias.n529 0.287138
R22111 commonsourceibias.n100 commonsourceibias.n12 0.285035
R22112 commonsourceibias.n193 commonsourceibias.n0 0.285035
R22113 commonsourceibias.n372 commonsourceibias.n284 0.285035
R22114 commonsourceibias.n282 commonsourceibias.n194 0.285035
R22115 commonsourceibias.n521 commonsourceibias.n433 0.285035
R22116 commonsourceibias.n567 commonsourceibias.n374 0.285035
R22117 commonsourceibias.n746 commonsourceibias.n658 0.285035
R22118 commonsourceibias.n656 commonsourceibias.n568 0.285035
R22119 commonsourceibias.n22 commonsourceibias.n20 0.246418
R22120 commonsourceibias.n58 commonsourceibias.n25 0.246418
R22121 commonsourceibias.n10 commonsourceibias.n8 0.246418
R22122 commonsourceibias.n151 commonsourceibias.n118 0.246418
R22123 commonsourceibias.n330 commonsourceibias.n297 0.246418
R22124 commonsourceibias.n294 commonsourceibias.n292 0.246418
R22125 commonsourceibias.n204 commonsourceibias.n202 0.246418
R22126 commonsourceibias.n240 commonsourceibias.n207 0.246418
R22127 commonsourceibias.n477 commonsourceibias.n444 0.246418
R22128 commonsourceibias.n490 commonsourceibias.n440 0.246418
R22129 commonsourceibias.n536 commonsourceibias.n381 0.246418
R22130 commonsourceibias.n418 commonsourceibias.n385 0.246418
R22131 commonsourceibias.n702 commonsourceibias.n669 0.246418
R22132 commonsourceibias.n715 commonsourceibias.n665 0.246418
R22133 commonsourceibias.n612 commonsourceibias.n579 0.246418
R22134 commonsourceibias.n625 commonsourceibias.n575 0.246418
R22135 commonsourceibias.n95 commonsourceibias.n12 0.189894
R22136 commonsourceibias.n95 commonsourceibias.n94 0.189894
R22137 commonsourceibias.n94 commonsourceibias.n93 0.189894
R22138 commonsourceibias.n93 commonsourceibias.n14 0.189894
R22139 commonsourceibias.n88 commonsourceibias.n14 0.189894
R22140 commonsourceibias.n88 commonsourceibias.n87 0.189894
R22141 commonsourceibias.n87 commonsourceibias.n86 0.189894
R22142 commonsourceibias.n86 commonsourceibias.n16 0.189894
R22143 commonsourceibias.n81 commonsourceibias.n16 0.189894
R22144 commonsourceibias.n81 commonsourceibias.n80 0.189894
R22145 commonsourceibias.n80 commonsourceibias.n79 0.189894
R22146 commonsourceibias.n79 commonsourceibias.n19 0.189894
R22147 commonsourceibias.n74 commonsourceibias.n19 0.189894
R22148 commonsourceibias.n74 commonsourceibias.n73 0.189894
R22149 commonsourceibias.n73 commonsourceibias.n72 0.189894
R22150 commonsourceibias.n72 commonsourceibias.n21 0.189894
R22151 commonsourceibias.n67 commonsourceibias.n21 0.189894
R22152 commonsourceibias.n67 commonsourceibias.n66 0.189894
R22153 commonsourceibias.n66 commonsourceibias.n65 0.189894
R22154 commonsourceibias.n65 commonsourceibias.n24 0.189894
R22155 commonsourceibias.n60 commonsourceibias.n24 0.189894
R22156 commonsourceibias.n60 commonsourceibias.n59 0.189894
R22157 commonsourceibias.n59 commonsourceibias.n26 0.189894
R22158 commonsourceibias.n55 commonsourceibias.n26 0.189894
R22159 commonsourceibias.n55 commonsourceibias.n54 0.189894
R22160 commonsourceibias.n54 commonsourceibias.n28 0.189894
R22161 commonsourceibias.n50 commonsourceibias.n28 0.189894
R22162 commonsourceibias.n50 commonsourceibias.n49 0.189894
R22163 commonsourceibias.n49 commonsourceibias.n30 0.189894
R22164 commonsourceibias.n44 commonsourceibias.n30 0.189894
R22165 commonsourceibias.n44 commonsourceibias.n43 0.189894
R22166 commonsourceibias.n43 commonsourceibias.n42 0.189894
R22167 commonsourceibias.n42 commonsourceibias.n32 0.189894
R22168 commonsourceibias.n37 commonsourceibias.n32 0.189894
R22169 commonsourceibias.n37 commonsourceibias.n36 0.189894
R22170 commonsourceibias.n158 commonsourceibias.n117 0.189894
R22171 commonsourceibias.n153 commonsourceibias.n117 0.189894
R22172 commonsourceibias.n153 commonsourceibias.n152 0.189894
R22173 commonsourceibias.n152 commonsourceibias.n119 0.189894
R22174 commonsourceibias.n148 commonsourceibias.n119 0.189894
R22175 commonsourceibias.n148 commonsourceibias.n147 0.189894
R22176 commonsourceibias.n147 commonsourceibias.n121 0.189894
R22177 commonsourceibias.n143 commonsourceibias.n121 0.189894
R22178 commonsourceibias.n143 commonsourceibias.n142 0.189894
R22179 commonsourceibias.n142 commonsourceibias.n123 0.189894
R22180 commonsourceibias.n137 commonsourceibias.n123 0.189894
R22181 commonsourceibias.n137 commonsourceibias.n136 0.189894
R22182 commonsourceibias.n136 commonsourceibias.n135 0.189894
R22183 commonsourceibias.n135 commonsourceibias.n125 0.189894
R22184 commonsourceibias.n130 commonsourceibias.n125 0.189894
R22185 commonsourceibias.n130 commonsourceibias.n129 0.189894
R22186 commonsourceibias.n188 commonsourceibias.n0 0.189894
R22187 commonsourceibias.n188 commonsourceibias.n187 0.189894
R22188 commonsourceibias.n187 commonsourceibias.n186 0.189894
R22189 commonsourceibias.n186 commonsourceibias.n2 0.189894
R22190 commonsourceibias.n181 commonsourceibias.n2 0.189894
R22191 commonsourceibias.n181 commonsourceibias.n180 0.189894
R22192 commonsourceibias.n180 commonsourceibias.n179 0.189894
R22193 commonsourceibias.n179 commonsourceibias.n4 0.189894
R22194 commonsourceibias.n174 commonsourceibias.n4 0.189894
R22195 commonsourceibias.n174 commonsourceibias.n173 0.189894
R22196 commonsourceibias.n173 commonsourceibias.n172 0.189894
R22197 commonsourceibias.n172 commonsourceibias.n7 0.189894
R22198 commonsourceibias.n167 commonsourceibias.n7 0.189894
R22199 commonsourceibias.n167 commonsourceibias.n166 0.189894
R22200 commonsourceibias.n166 commonsourceibias.n165 0.189894
R22201 commonsourceibias.n165 commonsourceibias.n9 0.189894
R22202 commonsourceibias.n160 commonsourceibias.n9 0.189894
R22203 commonsourceibias.n367 commonsourceibias.n284 0.189894
R22204 commonsourceibias.n367 commonsourceibias.n366 0.189894
R22205 commonsourceibias.n366 commonsourceibias.n365 0.189894
R22206 commonsourceibias.n365 commonsourceibias.n286 0.189894
R22207 commonsourceibias.n360 commonsourceibias.n286 0.189894
R22208 commonsourceibias.n360 commonsourceibias.n359 0.189894
R22209 commonsourceibias.n359 commonsourceibias.n358 0.189894
R22210 commonsourceibias.n358 commonsourceibias.n288 0.189894
R22211 commonsourceibias.n353 commonsourceibias.n288 0.189894
R22212 commonsourceibias.n353 commonsourceibias.n352 0.189894
R22213 commonsourceibias.n352 commonsourceibias.n351 0.189894
R22214 commonsourceibias.n351 commonsourceibias.n291 0.189894
R22215 commonsourceibias.n346 commonsourceibias.n291 0.189894
R22216 commonsourceibias.n346 commonsourceibias.n345 0.189894
R22217 commonsourceibias.n345 commonsourceibias.n344 0.189894
R22218 commonsourceibias.n344 commonsourceibias.n293 0.189894
R22219 commonsourceibias.n339 commonsourceibias.n293 0.189894
R22220 commonsourceibias.n339 commonsourceibias.n338 0.189894
R22221 commonsourceibias.n338 commonsourceibias.n337 0.189894
R22222 commonsourceibias.n337 commonsourceibias.n296 0.189894
R22223 commonsourceibias.n332 commonsourceibias.n296 0.189894
R22224 commonsourceibias.n332 commonsourceibias.n331 0.189894
R22225 commonsourceibias.n331 commonsourceibias.n298 0.189894
R22226 commonsourceibias.n327 commonsourceibias.n298 0.189894
R22227 commonsourceibias.n327 commonsourceibias.n326 0.189894
R22228 commonsourceibias.n326 commonsourceibias.n300 0.189894
R22229 commonsourceibias.n322 commonsourceibias.n300 0.189894
R22230 commonsourceibias.n322 commonsourceibias.n321 0.189894
R22231 commonsourceibias.n321 commonsourceibias.n302 0.189894
R22232 commonsourceibias.n316 commonsourceibias.n302 0.189894
R22233 commonsourceibias.n316 commonsourceibias.n315 0.189894
R22234 commonsourceibias.n315 commonsourceibias.n314 0.189894
R22235 commonsourceibias.n314 commonsourceibias.n304 0.189894
R22236 commonsourceibias.n309 commonsourceibias.n304 0.189894
R22237 commonsourceibias.n309 commonsourceibias.n308 0.189894
R22238 commonsourceibias.n277 commonsourceibias.n194 0.189894
R22239 commonsourceibias.n277 commonsourceibias.n276 0.189894
R22240 commonsourceibias.n276 commonsourceibias.n275 0.189894
R22241 commonsourceibias.n275 commonsourceibias.n196 0.189894
R22242 commonsourceibias.n270 commonsourceibias.n196 0.189894
R22243 commonsourceibias.n270 commonsourceibias.n269 0.189894
R22244 commonsourceibias.n269 commonsourceibias.n268 0.189894
R22245 commonsourceibias.n268 commonsourceibias.n198 0.189894
R22246 commonsourceibias.n263 commonsourceibias.n198 0.189894
R22247 commonsourceibias.n263 commonsourceibias.n262 0.189894
R22248 commonsourceibias.n262 commonsourceibias.n261 0.189894
R22249 commonsourceibias.n261 commonsourceibias.n201 0.189894
R22250 commonsourceibias.n256 commonsourceibias.n201 0.189894
R22251 commonsourceibias.n256 commonsourceibias.n255 0.189894
R22252 commonsourceibias.n255 commonsourceibias.n254 0.189894
R22253 commonsourceibias.n254 commonsourceibias.n203 0.189894
R22254 commonsourceibias.n249 commonsourceibias.n203 0.189894
R22255 commonsourceibias.n249 commonsourceibias.n248 0.189894
R22256 commonsourceibias.n248 commonsourceibias.n247 0.189894
R22257 commonsourceibias.n247 commonsourceibias.n206 0.189894
R22258 commonsourceibias.n242 commonsourceibias.n206 0.189894
R22259 commonsourceibias.n242 commonsourceibias.n241 0.189894
R22260 commonsourceibias.n241 commonsourceibias.n208 0.189894
R22261 commonsourceibias.n237 commonsourceibias.n208 0.189894
R22262 commonsourceibias.n237 commonsourceibias.n236 0.189894
R22263 commonsourceibias.n236 commonsourceibias.n210 0.189894
R22264 commonsourceibias.n232 commonsourceibias.n210 0.189894
R22265 commonsourceibias.n232 commonsourceibias.n231 0.189894
R22266 commonsourceibias.n231 commonsourceibias.n212 0.189894
R22267 commonsourceibias.n226 commonsourceibias.n212 0.189894
R22268 commonsourceibias.n226 commonsourceibias.n225 0.189894
R22269 commonsourceibias.n225 commonsourceibias.n224 0.189894
R22270 commonsourceibias.n224 commonsourceibias.n214 0.189894
R22271 commonsourceibias.n219 commonsourceibias.n214 0.189894
R22272 commonsourceibias.n219 commonsourceibias.n218 0.189894
R22273 commonsourceibias.n456 commonsourceibias.n455 0.189894
R22274 commonsourceibias.n456 commonsourceibias.n451 0.189894
R22275 commonsourceibias.n461 commonsourceibias.n451 0.189894
R22276 commonsourceibias.n462 commonsourceibias.n461 0.189894
R22277 commonsourceibias.n463 commonsourceibias.n462 0.189894
R22278 commonsourceibias.n463 commonsourceibias.n449 0.189894
R22279 commonsourceibias.n468 commonsourceibias.n449 0.189894
R22280 commonsourceibias.n469 commonsourceibias.n468 0.189894
R22281 commonsourceibias.n469 commonsourceibias.n447 0.189894
R22282 commonsourceibias.n473 commonsourceibias.n447 0.189894
R22283 commonsourceibias.n474 commonsourceibias.n473 0.189894
R22284 commonsourceibias.n474 commonsourceibias.n445 0.189894
R22285 commonsourceibias.n478 commonsourceibias.n445 0.189894
R22286 commonsourceibias.n479 commonsourceibias.n478 0.189894
R22287 commonsourceibias.n479 commonsourceibias.n443 0.189894
R22288 commonsourceibias.n484 commonsourceibias.n443 0.189894
R22289 commonsourceibias.n485 commonsourceibias.n484 0.189894
R22290 commonsourceibias.n486 commonsourceibias.n485 0.189894
R22291 commonsourceibias.n486 commonsourceibias.n441 0.189894
R22292 commonsourceibias.n492 commonsourceibias.n441 0.189894
R22293 commonsourceibias.n493 commonsourceibias.n492 0.189894
R22294 commonsourceibias.n494 commonsourceibias.n493 0.189894
R22295 commonsourceibias.n494 commonsourceibias.n439 0.189894
R22296 commonsourceibias.n499 commonsourceibias.n439 0.189894
R22297 commonsourceibias.n500 commonsourceibias.n499 0.189894
R22298 commonsourceibias.n501 commonsourceibias.n500 0.189894
R22299 commonsourceibias.n501 commonsourceibias.n437 0.189894
R22300 commonsourceibias.n507 commonsourceibias.n437 0.189894
R22301 commonsourceibias.n508 commonsourceibias.n507 0.189894
R22302 commonsourceibias.n509 commonsourceibias.n508 0.189894
R22303 commonsourceibias.n509 commonsourceibias.n435 0.189894
R22304 commonsourceibias.n514 commonsourceibias.n435 0.189894
R22305 commonsourceibias.n515 commonsourceibias.n514 0.189894
R22306 commonsourceibias.n516 commonsourceibias.n515 0.189894
R22307 commonsourceibias.n516 commonsourceibias.n433 0.189894
R22308 commonsourceibias.n397 commonsourceibias.n396 0.189894
R22309 commonsourceibias.n397 commonsourceibias.n392 0.189894
R22310 commonsourceibias.n402 commonsourceibias.n392 0.189894
R22311 commonsourceibias.n403 commonsourceibias.n402 0.189894
R22312 commonsourceibias.n404 commonsourceibias.n403 0.189894
R22313 commonsourceibias.n404 commonsourceibias.n390 0.189894
R22314 commonsourceibias.n409 commonsourceibias.n390 0.189894
R22315 commonsourceibias.n410 commonsourceibias.n409 0.189894
R22316 commonsourceibias.n410 commonsourceibias.n388 0.189894
R22317 commonsourceibias.n414 commonsourceibias.n388 0.189894
R22318 commonsourceibias.n415 commonsourceibias.n414 0.189894
R22319 commonsourceibias.n415 commonsourceibias.n386 0.189894
R22320 commonsourceibias.n419 commonsourceibias.n386 0.189894
R22321 commonsourceibias.n420 commonsourceibias.n419 0.189894
R22322 commonsourceibias.n420 commonsourceibias.n384 0.189894
R22323 commonsourceibias.n425 commonsourceibias.n384 0.189894
R22324 commonsourceibias.n532 commonsourceibias.n382 0.189894
R22325 commonsourceibias.n538 commonsourceibias.n382 0.189894
R22326 commonsourceibias.n539 commonsourceibias.n538 0.189894
R22327 commonsourceibias.n540 commonsourceibias.n539 0.189894
R22328 commonsourceibias.n540 commonsourceibias.n380 0.189894
R22329 commonsourceibias.n545 commonsourceibias.n380 0.189894
R22330 commonsourceibias.n546 commonsourceibias.n545 0.189894
R22331 commonsourceibias.n547 commonsourceibias.n546 0.189894
R22332 commonsourceibias.n547 commonsourceibias.n378 0.189894
R22333 commonsourceibias.n553 commonsourceibias.n378 0.189894
R22334 commonsourceibias.n554 commonsourceibias.n553 0.189894
R22335 commonsourceibias.n555 commonsourceibias.n554 0.189894
R22336 commonsourceibias.n555 commonsourceibias.n376 0.189894
R22337 commonsourceibias.n560 commonsourceibias.n376 0.189894
R22338 commonsourceibias.n561 commonsourceibias.n560 0.189894
R22339 commonsourceibias.n562 commonsourceibias.n561 0.189894
R22340 commonsourceibias.n562 commonsourceibias.n374 0.189894
R22341 commonsourceibias.n681 commonsourceibias.n680 0.189894
R22342 commonsourceibias.n681 commonsourceibias.n676 0.189894
R22343 commonsourceibias.n686 commonsourceibias.n676 0.189894
R22344 commonsourceibias.n687 commonsourceibias.n686 0.189894
R22345 commonsourceibias.n688 commonsourceibias.n687 0.189894
R22346 commonsourceibias.n688 commonsourceibias.n674 0.189894
R22347 commonsourceibias.n693 commonsourceibias.n674 0.189894
R22348 commonsourceibias.n694 commonsourceibias.n693 0.189894
R22349 commonsourceibias.n694 commonsourceibias.n672 0.189894
R22350 commonsourceibias.n698 commonsourceibias.n672 0.189894
R22351 commonsourceibias.n699 commonsourceibias.n698 0.189894
R22352 commonsourceibias.n699 commonsourceibias.n670 0.189894
R22353 commonsourceibias.n703 commonsourceibias.n670 0.189894
R22354 commonsourceibias.n704 commonsourceibias.n703 0.189894
R22355 commonsourceibias.n704 commonsourceibias.n668 0.189894
R22356 commonsourceibias.n709 commonsourceibias.n668 0.189894
R22357 commonsourceibias.n710 commonsourceibias.n709 0.189894
R22358 commonsourceibias.n711 commonsourceibias.n710 0.189894
R22359 commonsourceibias.n711 commonsourceibias.n666 0.189894
R22360 commonsourceibias.n717 commonsourceibias.n666 0.189894
R22361 commonsourceibias.n718 commonsourceibias.n717 0.189894
R22362 commonsourceibias.n719 commonsourceibias.n718 0.189894
R22363 commonsourceibias.n719 commonsourceibias.n664 0.189894
R22364 commonsourceibias.n724 commonsourceibias.n664 0.189894
R22365 commonsourceibias.n725 commonsourceibias.n724 0.189894
R22366 commonsourceibias.n726 commonsourceibias.n725 0.189894
R22367 commonsourceibias.n726 commonsourceibias.n662 0.189894
R22368 commonsourceibias.n732 commonsourceibias.n662 0.189894
R22369 commonsourceibias.n733 commonsourceibias.n732 0.189894
R22370 commonsourceibias.n734 commonsourceibias.n733 0.189894
R22371 commonsourceibias.n734 commonsourceibias.n660 0.189894
R22372 commonsourceibias.n739 commonsourceibias.n660 0.189894
R22373 commonsourceibias.n740 commonsourceibias.n739 0.189894
R22374 commonsourceibias.n741 commonsourceibias.n740 0.189894
R22375 commonsourceibias.n741 commonsourceibias.n658 0.189894
R22376 commonsourceibias.n591 commonsourceibias.n590 0.189894
R22377 commonsourceibias.n591 commonsourceibias.n586 0.189894
R22378 commonsourceibias.n596 commonsourceibias.n586 0.189894
R22379 commonsourceibias.n597 commonsourceibias.n596 0.189894
R22380 commonsourceibias.n598 commonsourceibias.n597 0.189894
R22381 commonsourceibias.n598 commonsourceibias.n584 0.189894
R22382 commonsourceibias.n603 commonsourceibias.n584 0.189894
R22383 commonsourceibias.n604 commonsourceibias.n603 0.189894
R22384 commonsourceibias.n604 commonsourceibias.n582 0.189894
R22385 commonsourceibias.n608 commonsourceibias.n582 0.189894
R22386 commonsourceibias.n609 commonsourceibias.n608 0.189894
R22387 commonsourceibias.n609 commonsourceibias.n580 0.189894
R22388 commonsourceibias.n613 commonsourceibias.n580 0.189894
R22389 commonsourceibias.n614 commonsourceibias.n613 0.189894
R22390 commonsourceibias.n614 commonsourceibias.n578 0.189894
R22391 commonsourceibias.n619 commonsourceibias.n578 0.189894
R22392 commonsourceibias.n620 commonsourceibias.n619 0.189894
R22393 commonsourceibias.n621 commonsourceibias.n620 0.189894
R22394 commonsourceibias.n621 commonsourceibias.n576 0.189894
R22395 commonsourceibias.n627 commonsourceibias.n576 0.189894
R22396 commonsourceibias.n628 commonsourceibias.n627 0.189894
R22397 commonsourceibias.n629 commonsourceibias.n628 0.189894
R22398 commonsourceibias.n629 commonsourceibias.n574 0.189894
R22399 commonsourceibias.n634 commonsourceibias.n574 0.189894
R22400 commonsourceibias.n635 commonsourceibias.n634 0.189894
R22401 commonsourceibias.n636 commonsourceibias.n635 0.189894
R22402 commonsourceibias.n636 commonsourceibias.n572 0.189894
R22403 commonsourceibias.n642 commonsourceibias.n572 0.189894
R22404 commonsourceibias.n643 commonsourceibias.n642 0.189894
R22405 commonsourceibias.n644 commonsourceibias.n643 0.189894
R22406 commonsourceibias.n644 commonsourceibias.n570 0.189894
R22407 commonsourceibias.n649 commonsourceibias.n570 0.189894
R22408 commonsourceibias.n650 commonsourceibias.n649 0.189894
R22409 commonsourceibias.n651 commonsourceibias.n650 0.189894
R22410 commonsourceibias.n651 commonsourceibias.n568 0.189894
R22411 commonsourceibias.n159 commonsourceibias.n158 0.170955
R22412 commonsourceibias.n160 commonsourceibias.n159 0.170955
R22413 commonsourceibias.n531 commonsourceibias.n425 0.170955
R22414 commonsourceibias.n532 commonsourceibias.n531 0.170955
R22415 CSoutput.n19 CSoutput.t185 184.661
R22416 CSoutput.n78 CSoutput.n77 165.8
R22417 CSoutput.n76 CSoutput.n0 165.8
R22418 CSoutput.n75 CSoutput.n74 165.8
R22419 CSoutput.n73 CSoutput.n72 165.8
R22420 CSoutput.n71 CSoutput.n2 165.8
R22421 CSoutput.n69 CSoutput.n68 165.8
R22422 CSoutput.n67 CSoutput.n3 165.8
R22423 CSoutput.n66 CSoutput.n65 165.8
R22424 CSoutput.n63 CSoutput.n4 165.8
R22425 CSoutput.n61 CSoutput.n60 165.8
R22426 CSoutput.n59 CSoutput.n5 165.8
R22427 CSoutput.n58 CSoutput.n57 165.8
R22428 CSoutput.n55 CSoutput.n6 165.8
R22429 CSoutput.n54 CSoutput.n53 165.8
R22430 CSoutput.n52 CSoutput.n51 165.8
R22431 CSoutput.n50 CSoutput.n8 165.8
R22432 CSoutput.n48 CSoutput.n47 165.8
R22433 CSoutput.n46 CSoutput.n9 165.8
R22434 CSoutput.n45 CSoutput.n44 165.8
R22435 CSoutput.n42 CSoutput.n10 165.8
R22436 CSoutput.n41 CSoutput.n40 165.8
R22437 CSoutput.n39 CSoutput.n38 165.8
R22438 CSoutput.n37 CSoutput.n12 165.8
R22439 CSoutput.n35 CSoutput.n34 165.8
R22440 CSoutput.n33 CSoutput.n13 165.8
R22441 CSoutput.n32 CSoutput.n31 165.8
R22442 CSoutput.n29 CSoutput.n14 165.8
R22443 CSoutput.n28 CSoutput.n27 165.8
R22444 CSoutput.n26 CSoutput.n25 165.8
R22445 CSoutput.n24 CSoutput.n16 165.8
R22446 CSoutput.n22 CSoutput.n21 165.8
R22447 CSoutput.n20 CSoutput.n17 165.8
R22448 CSoutput.n77 CSoutput.t187 162.194
R22449 CSoutput.n18 CSoutput.t182 120.501
R22450 CSoutput.n23 CSoutput.t176 120.501
R22451 CSoutput.n15 CSoutput.t171 120.501
R22452 CSoutput.n30 CSoutput.t183 120.501
R22453 CSoutput.n36 CSoutput.t184 120.501
R22454 CSoutput.n11 CSoutput.t173 120.501
R22455 CSoutput.n43 CSoutput.t169 120.501
R22456 CSoutput.n49 CSoutput.t186 120.501
R22457 CSoutput.n7 CSoutput.t177 120.501
R22458 CSoutput.n56 CSoutput.t179 120.501
R22459 CSoutput.n62 CSoutput.t188 120.501
R22460 CSoutput.n64 CSoutput.t180 120.501
R22461 CSoutput.n70 CSoutput.t181 120.501
R22462 CSoutput.n1 CSoutput.t174 120.501
R22463 CSoutput.n290 CSoutput.n288 103.469
R22464 CSoutput.n278 CSoutput.n276 103.469
R22465 CSoutput.n267 CSoutput.n265 103.469
R22466 CSoutput.n104 CSoutput.n102 103.469
R22467 CSoutput.n92 CSoutput.n90 103.469
R22468 CSoutput.n81 CSoutput.n79 103.469
R22469 CSoutput.n296 CSoutput.n295 103.111
R22470 CSoutput.n294 CSoutput.n293 103.111
R22471 CSoutput.n292 CSoutput.n291 103.111
R22472 CSoutput.n290 CSoutput.n289 103.111
R22473 CSoutput.n286 CSoutput.n285 103.111
R22474 CSoutput.n284 CSoutput.n283 103.111
R22475 CSoutput.n282 CSoutput.n281 103.111
R22476 CSoutput.n280 CSoutput.n279 103.111
R22477 CSoutput.n278 CSoutput.n277 103.111
R22478 CSoutput.n275 CSoutput.n274 103.111
R22479 CSoutput.n273 CSoutput.n272 103.111
R22480 CSoutput.n271 CSoutput.n270 103.111
R22481 CSoutput.n269 CSoutput.n268 103.111
R22482 CSoutput.n267 CSoutput.n266 103.111
R22483 CSoutput.n104 CSoutput.n103 103.111
R22484 CSoutput.n106 CSoutput.n105 103.111
R22485 CSoutput.n108 CSoutput.n107 103.111
R22486 CSoutput.n110 CSoutput.n109 103.111
R22487 CSoutput.n112 CSoutput.n111 103.111
R22488 CSoutput.n92 CSoutput.n91 103.111
R22489 CSoutput.n94 CSoutput.n93 103.111
R22490 CSoutput.n96 CSoutput.n95 103.111
R22491 CSoutput.n98 CSoutput.n97 103.111
R22492 CSoutput.n100 CSoutput.n99 103.111
R22493 CSoutput.n81 CSoutput.n80 103.111
R22494 CSoutput.n83 CSoutput.n82 103.111
R22495 CSoutput.n85 CSoutput.n84 103.111
R22496 CSoutput.n87 CSoutput.n86 103.111
R22497 CSoutput.n89 CSoutput.n88 103.111
R22498 CSoutput.n298 CSoutput.n297 103.111
R22499 CSoutput.n334 CSoutput.n332 81.5057
R22500 CSoutput.n318 CSoutput.n316 81.5057
R22501 CSoutput.n303 CSoutput.n301 81.5057
R22502 CSoutput.n382 CSoutput.n380 81.5057
R22503 CSoutput.n366 CSoutput.n364 81.5057
R22504 CSoutput.n351 CSoutput.n349 81.5057
R22505 CSoutput.n346 CSoutput.n345 80.9324
R22506 CSoutput.n344 CSoutput.n343 80.9324
R22507 CSoutput.n342 CSoutput.n341 80.9324
R22508 CSoutput.n340 CSoutput.n339 80.9324
R22509 CSoutput.n338 CSoutput.n337 80.9324
R22510 CSoutput.n336 CSoutput.n335 80.9324
R22511 CSoutput.n334 CSoutput.n333 80.9324
R22512 CSoutput.n330 CSoutput.n329 80.9324
R22513 CSoutput.n328 CSoutput.n327 80.9324
R22514 CSoutput.n326 CSoutput.n325 80.9324
R22515 CSoutput.n324 CSoutput.n323 80.9324
R22516 CSoutput.n322 CSoutput.n321 80.9324
R22517 CSoutput.n320 CSoutput.n319 80.9324
R22518 CSoutput.n318 CSoutput.n317 80.9324
R22519 CSoutput.n315 CSoutput.n314 80.9324
R22520 CSoutput.n313 CSoutput.n312 80.9324
R22521 CSoutput.n311 CSoutput.n310 80.9324
R22522 CSoutput.n309 CSoutput.n308 80.9324
R22523 CSoutput.n307 CSoutput.n306 80.9324
R22524 CSoutput.n305 CSoutput.n304 80.9324
R22525 CSoutput.n303 CSoutput.n302 80.9324
R22526 CSoutput.n382 CSoutput.n381 80.9324
R22527 CSoutput.n384 CSoutput.n383 80.9324
R22528 CSoutput.n386 CSoutput.n385 80.9324
R22529 CSoutput.n388 CSoutput.n387 80.9324
R22530 CSoutput.n390 CSoutput.n389 80.9324
R22531 CSoutput.n392 CSoutput.n391 80.9324
R22532 CSoutput.n394 CSoutput.n393 80.9324
R22533 CSoutput.n366 CSoutput.n365 80.9324
R22534 CSoutput.n368 CSoutput.n367 80.9324
R22535 CSoutput.n370 CSoutput.n369 80.9324
R22536 CSoutput.n372 CSoutput.n371 80.9324
R22537 CSoutput.n374 CSoutput.n373 80.9324
R22538 CSoutput.n376 CSoutput.n375 80.9324
R22539 CSoutput.n378 CSoutput.n377 80.9324
R22540 CSoutput.n351 CSoutput.n350 80.9324
R22541 CSoutput.n353 CSoutput.n352 80.9324
R22542 CSoutput.n355 CSoutput.n354 80.9324
R22543 CSoutput.n357 CSoutput.n356 80.9324
R22544 CSoutput.n359 CSoutput.n358 80.9324
R22545 CSoutput.n361 CSoutput.n360 80.9324
R22546 CSoutput.n363 CSoutput.n362 80.9324
R22547 CSoutput.n25 CSoutput.n24 48.1486
R22548 CSoutput.n69 CSoutput.n3 48.1486
R22549 CSoutput.n38 CSoutput.n37 48.1486
R22550 CSoutput.n42 CSoutput.n41 48.1486
R22551 CSoutput.n51 CSoutput.n50 48.1486
R22552 CSoutput.n55 CSoutput.n54 48.1486
R22553 CSoutput.n22 CSoutput.n17 46.462
R22554 CSoutput.n72 CSoutput.n71 46.462
R22555 CSoutput.n20 CSoutput.n19 44.9055
R22556 CSoutput.n29 CSoutput.n28 43.7635
R22557 CSoutput.n65 CSoutput.n63 43.7635
R22558 CSoutput.n35 CSoutput.n13 41.7396
R22559 CSoutput.n57 CSoutput.n5 41.7396
R22560 CSoutput.n44 CSoutput.n9 37.0171
R22561 CSoutput.n48 CSoutput.n9 37.0171
R22562 CSoutput.n76 CSoutput.n75 34.9932
R22563 CSoutput.n31 CSoutput.n13 32.2947
R22564 CSoutput.n61 CSoutput.n5 32.2947
R22565 CSoutput.n30 CSoutput.n29 29.6014
R22566 CSoutput.n63 CSoutput.n62 29.6014
R22567 CSoutput.n19 CSoutput.n18 28.4085
R22568 CSoutput.n18 CSoutput.n17 25.1176
R22569 CSoutput.n72 CSoutput.n1 25.1176
R22570 CSoutput.n43 CSoutput.n42 22.0922
R22571 CSoutput.n50 CSoutput.n49 22.0922
R22572 CSoutput.n77 CSoutput.n76 21.8586
R22573 CSoutput.n37 CSoutput.n36 18.9681
R22574 CSoutput.n56 CSoutput.n55 18.9681
R22575 CSoutput.n25 CSoutput.n15 17.6292
R22576 CSoutput.n64 CSoutput.n3 17.6292
R22577 CSoutput.n24 CSoutput.n23 15.844
R22578 CSoutput.n70 CSoutput.n69 15.844
R22579 CSoutput.n38 CSoutput.n11 14.5051
R22580 CSoutput.n54 CSoutput.n7 14.5051
R22581 CSoutput.n397 CSoutput.n78 11.4982
R22582 CSoutput.n41 CSoutput.n11 11.3811
R22583 CSoutput.n51 CSoutput.n7 11.3811
R22584 CSoutput.n23 CSoutput.n22 10.0422
R22585 CSoutput.n71 CSoutput.n70 10.0422
R22586 CSoutput.n287 CSoutput.n275 9.25285
R22587 CSoutput.n101 CSoutput.n89 9.25285
R22588 CSoutput.n331 CSoutput.n315 8.98182
R22589 CSoutput.n379 CSoutput.n363 8.98182
R22590 CSoutput.n348 CSoutput.n300 8.67888
R22591 CSoutput.n28 CSoutput.n15 8.25698
R22592 CSoutput.n65 CSoutput.n64 8.25698
R22593 CSoutput.n300 CSoutput.n299 7.12641
R22594 CSoutput.n114 CSoutput.n113 7.12641
R22595 CSoutput.n36 CSoutput.n35 6.91809
R22596 CSoutput.n57 CSoutput.n56 6.91809
R22597 CSoutput.n348 CSoutput.n347 6.02792
R22598 CSoutput.n396 CSoutput.n395 6.02792
R22599 CSoutput.n347 CSoutput.n346 5.25266
R22600 CSoutput.n331 CSoutput.n330 5.25266
R22601 CSoutput.n395 CSoutput.n394 5.25266
R22602 CSoutput.n379 CSoutput.n378 5.25266
R22603 CSoutput.n299 CSoutput.n298 5.1449
R22604 CSoutput.n287 CSoutput.n286 5.1449
R22605 CSoutput.n113 CSoutput.n112 5.1449
R22606 CSoutput.n101 CSoutput.n100 5.1449
R22607 CSoutput.n397 CSoutput.n114 5.08644
R22608 CSoutput.n205 CSoutput.n158 4.5005
R22609 CSoutput.n174 CSoutput.n158 4.5005
R22610 CSoutput.n169 CSoutput.n153 4.5005
R22611 CSoutput.n169 CSoutput.n155 4.5005
R22612 CSoutput.n169 CSoutput.n152 4.5005
R22613 CSoutput.n169 CSoutput.n156 4.5005
R22614 CSoutput.n169 CSoutput.n151 4.5005
R22615 CSoutput.n169 CSoutput.t189 4.5005
R22616 CSoutput.n169 CSoutput.n150 4.5005
R22617 CSoutput.n169 CSoutput.n157 4.5005
R22618 CSoutput.n169 CSoutput.n158 4.5005
R22619 CSoutput.n167 CSoutput.n153 4.5005
R22620 CSoutput.n167 CSoutput.n155 4.5005
R22621 CSoutput.n167 CSoutput.n152 4.5005
R22622 CSoutput.n167 CSoutput.n156 4.5005
R22623 CSoutput.n167 CSoutput.n151 4.5005
R22624 CSoutput.n167 CSoutput.t189 4.5005
R22625 CSoutput.n167 CSoutput.n150 4.5005
R22626 CSoutput.n167 CSoutput.n157 4.5005
R22627 CSoutput.n167 CSoutput.n158 4.5005
R22628 CSoutput.n166 CSoutput.n153 4.5005
R22629 CSoutput.n166 CSoutput.n155 4.5005
R22630 CSoutput.n166 CSoutput.n152 4.5005
R22631 CSoutput.n166 CSoutput.n156 4.5005
R22632 CSoutput.n166 CSoutput.n151 4.5005
R22633 CSoutput.n166 CSoutput.t189 4.5005
R22634 CSoutput.n166 CSoutput.n150 4.5005
R22635 CSoutput.n166 CSoutput.n157 4.5005
R22636 CSoutput.n166 CSoutput.n158 4.5005
R22637 CSoutput.n251 CSoutput.n153 4.5005
R22638 CSoutput.n251 CSoutput.n155 4.5005
R22639 CSoutput.n251 CSoutput.n152 4.5005
R22640 CSoutput.n251 CSoutput.n156 4.5005
R22641 CSoutput.n251 CSoutput.n151 4.5005
R22642 CSoutput.n251 CSoutput.t189 4.5005
R22643 CSoutput.n251 CSoutput.n150 4.5005
R22644 CSoutput.n251 CSoutput.n157 4.5005
R22645 CSoutput.n251 CSoutput.n158 4.5005
R22646 CSoutput.n249 CSoutput.n153 4.5005
R22647 CSoutput.n249 CSoutput.n155 4.5005
R22648 CSoutput.n249 CSoutput.n152 4.5005
R22649 CSoutput.n249 CSoutput.n156 4.5005
R22650 CSoutput.n249 CSoutput.n151 4.5005
R22651 CSoutput.n249 CSoutput.t189 4.5005
R22652 CSoutput.n249 CSoutput.n150 4.5005
R22653 CSoutput.n249 CSoutput.n157 4.5005
R22654 CSoutput.n247 CSoutput.n153 4.5005
R22655 CSoutput.n247 CSoutput.n155 4.5005
R22656 CSoutput.n247 CSoutput.n152 4.5005
R22657 CSoutput.n247 CSoutput.n156 4.5005
R22658 CSoutput.n247 CSoutput.n151 4.5005
R22659 CSoutput.n247 CSoutput.t189 4.5005
R22660 CSoutput.n247 CSoutput.n150 4.5005
R22661 CSoutput.n247 CSoutput.n157 4.5005
R22662 CSoutput.n177 CSoutput.n153 4.5005
R22663 CSoutput.n177 CSoutput.n155 4.5005
R22664 CSoutput.n177 CSoutput.n152 4.5005
R22665 CSoutput.n177 CSoutput.n156 4.5005
R22666 CSoutput.n177 CSoutput.n151 4.5005
R22667 CSoutput.n177 CSoutput.t189 4.5005
R22668 CSoutput.n177 CSoutput.n150 4.5005
R22669 CSoutput.n177 CSoutput.n157 4.5005
R22670 CSoutput.n177 CSoutput.n158 4.5005
R22671 CSoutput.n176 CSoutput.n153 4.5005
R22672 CSoutput.n176 CSoutput.n155 4.5005
R22673 CSoutput.n176 CSoutput.n152 4.5005
R22674 CSoutput.n176 CSoutput.n156 4.5005
R22675 CSoutput.n176 CSoutput.n151 4.5005
R22676 CSoutput.n176 CSoutput.t189 4.5005
R22677 CSoutput.n176 CSoutput.n150 4.5005
R22678 CSoutput.n176 CSoutput.n157 4.5005
R22679 CSoutput.n176 CSoutput.n158 4.5005
R22680 CSoutput.n180 CSoutput.n153 4.5005
R22681 CSoutput.n180 CSoutput.n155 4.5005
R22682 CSoutput.n180 CSoutput.n152 4.5005
R22683 CSoutput.n180 CSoutput.n156 4.5005
R22684 CSoutput.n180 CSoutput.n151 4.5005
R22685 CSoutput.n180 CSoutput.t189 4.5005
R22686 CSoutput.n180 CSoutput.n150 4.5005
R22687 CSoutput.n180 CSoutput.n157 4.5005
R22688 CSoutput.n180 CSoutput.n158 4.5005
R22689 CSoutput.n179 CSoutput.n153 4.5005
R22690 CSoutput.n179 CSoutput.n155 4.5005
R22691 CSoutput.n179 CSoutput.n152 4.5005
R22692 CSoutput.n179 CSoutput.n156 4.5005
R22693 CSoutput.n179 CSoutput.n151 4.5005
R22694 CSoutput.n179 CSoutput.t189 4.5005
R22695 CSoutput.n179 CSoutput.n150 4.5005
R22696 CSoutput.n179 CSoutput.n157 4.5005
R22697 CSoutput.n179 CSoutput.n158 4.5005
R22698 CSoutput.n162 CSoutput.n153 4.5005
R22699 CSoutput.n162 CSoutput.n155 4.5005
R22700 CSoutput.n162 CSoutput.n152 4.5005
R22701 CSoutput.n162 CSoutput.n156 4.5005
R22702 CSoutput.n162 CSoutput.n151 4.5005
R22703 CSoutput.n162 CSoutput.t189 4.5005
R22704 CSoutput.n162 CSoutput.n150 4.5005
R22705 CSoutput.n162 CSoutput.n157 4.5005
R22706 CSoutput.n162 CSoutput.n158 4.5005
R22707 CSoutput.n254 CSoutput.n153 4.5005
R22708 CSoutput.n254 CSoutput.n155 4.5005
R22709 CSoutput.n254 CSoutput.n152 4.5005
R22710 CSoutput.n254 CSoutput.n156 4.5005
R22711 CSoutput.n254 CSoutput.n151 4.5005
R22712 CSoutput.n254 CSoutput.t189 4.5005
R22713 CSoutput.n254 CSoutput.n150 4.5005
R22714 CSoutput.n254 CSoutput.n157 4.5005
R22715 CSoutput.n254 CSoutput.n158 4.5005
R22716 CSoutput.n241 CSoutput.n212 4.5005
R22717 CSoutput.n241 CSoutput.n218 4.5005
R22718 CSoutput.n199 CSoutput.n188 4.5005
R22719 CSoutput.n199 CSoutput.n190 4.5005
R22720 CSoutput.n199 CSoutput.n187 4.5005
R22721 CSoutput.n199 CSoutput.n191 4.5005
R22722 CSoutput.n199 CSoutput.n186 4.5005
R22723 CSoutput.n199 CSoutput.t168 4.5005
R22724 CSoutput.n199 CSoutput.n185 4.5005
R22725 CSoutput.n199 CSoutput.n192 4.5005
R22726 CSoutput.n241 CSoutput.n199 4.5005
R22727 CSoutput.n220 CSoutput.n188 4.5005
R22728 CSoutput.n220 CSoutput.n190 4.5005
R22729 CSoutput.n220 CSoutput.n187 4.5005
R22730 CSoutput.n220 CSoutput.n191 4.5005
R22731 CSoutput.n220 CSoutput.n186 4.5005
R22732 CSoutput.n220 CSoutput.t168 4.5005
R22733 CSoutput.n220 CSoutput.n185 4.5005
R22734 CSoutput.n220 CSoutput.n192 4.5005
R22735 CSoutput.n241 CSoutput.n220 4.5005
R22736 CSoutput.n198 CSoutput.n188 4.5005
R22737 CSoutput.n198 CSoutput.n190 4.5005
R22738 CSoutput.n198 CSoutput.n187 4.5005
R22739 CSoutput.n198 CSoutput.n191 4.5005
R22740 CSoutput.n198 CSoutput.n186 4.5005
R22741 CSoutput.n198 CSoutput.t168 4.5005
R22742 CSoutput.n198 CSoutput.n185 4.5005
R22743 CSoutput.n198 CSoutput.n192 4.5005
R22744 CSoutput.n241 CSoutput.n198 4.5005
R22745 CSoutput.n222 CSoutput.n188 4.5005
R22746 CSoutput.n222 CSoutput.n190 4.5005
R22747 CSoutput.n222 CSoutput.n187 4.5005
R22748 CSoutput.n222 CSoutput.n191 4.5005
R22749 CSoutput.n222 CSoutput.n186 4.5005
R22750 CSoutput.n222 CSoutput.t168 4.5005
R22751 CSoutput.n222 CSoutput.n185 4.5005
R22752 CSoutput.n222 CSoutput.n192 4.5005
R22753 CSoutput.n241 CSoutput.n222 4.5005
R22754 CSoutput.n188 CSoutput.n183 4.5005
R22755 CSoutput.n190 CSoutput.n183 4.5005
R22756 CSoutput.n187 CSoutput.n183 4.5005
R22757 CSoutput.n191 CSoutput.n183 4.5005
R22758 CSoutput.n186 CSoutput.n183 4.5005
R22759 CSoutput.t168 CSoutput.n183 4.5005
R22760 CSoutput.n185 CSoutput.n183 4.5005
R22761 CSoutput.n192 CSoutput.n183 4.5005
R22762 CSoutput.n244 CSoutput.n188 4.5005
R22763 CSoutput.n244 CSoutput.n190 4.5005
R22764 CSoutput.n244 CSoutput.n187 4.5005
R22765 CSoutput.n244 CSoutput.n191 4.5005
R22766 CSoutput.n244 CSoutput.n186 4.5005
R22767 CSoutput.n244 CSoutput.t168 4.5005
R22768 CSoutput.n244 CSoutput.n185 4.5005
R22769 CSoutput.n244 CSoutput.n192 4.5005
R22770 CSoutput.n242 CSoutput.n188 4.5005
R22771 CSoutput.n242 CSoutput.n190 4.5005
R22772 CSoutput.n242 CSoutput.n187 4.5005
R22773 CSoutput.n242 CSoutput.n191 4.5005
R22774 CSoutput.n242 CSoutput.n186 4.5005
R22775 CSoutput.n242 CSoutput.t168 4.5005
R22776 CSoutput.n242 CSoutput.n185 4.5005
R22777 CSoutput.n242 CSoutput.n192 4.5005
R22778 CSoutput.n242 CSoutput.n241 4.5005
R22779 CSoutput.n224 CSoutput.n188 4.5005
R22780 CSoutput.n224 CSoutput.n190 4.5005
R22781 CSoutput.n224 CSoutput.n187 4.5005
R22782 CSoutput.n224 CSoutput.n191 4.5005
R22783 CSoutput.n224 CSoutput.n186 4.5005
R22784 CSoutput.n224 CSoutput.t168 4.5005
R22785 CSoutput.n224 CSoutput.n185 4.5005
R22786 CSoutput.n224 CSoutput.n192 4.5005
R22787 CSoutput.n241 CSoutput.n224 4.5005
R22788 CSoutput.n196 CSoutput.n188 4.5005
R22789 CSoutput.n196 CSoutput.n190 4.5005
R22790 CSoutput.n196 CSoutput.n187 4.5005
R22791 CSoutput.n196 CSoutput.n191 4.5005
R22792 CSoutput.n196 CSoutput.n186 4.5005
R22793 CSoutput.n196 CSoutput.t168 4.5005
R22794 CSoutput.n196 CSoutput.n185 4.5005
R22795 CSoutput.n196 CSoutput.n192 4.5005
R22796 CSoutput.n241 CSoutput.n196 4.5005
R22797 CSoutput.n226 CSoutput.n188 4.5005
R22798 CSoutput.n226 CSoutput.n190 4.5005
R22799 CSoutput.n226 CSoutput.n187 4.5005
R22800 CSoutput.n226 CSoutput.n191 4.5005
R22801 CSoutput.n226 CSoutput.n186 4.5005
R22802 CSoutput.n226 CSoutput.t168 4.5005
R22803 CSoutput.n226 CSoutput.n185 4.5005
R22804 CSoutput.n226 CSoutput.n192 4.5005
R22805 CSoutput.n241 CSoutput.n226 4.5005
R22806 CSoutput.n195 CSoutput.n188 4.5005
R22807 CSoutput.n195 CSoutput.n190 4.5005
R22808 CSoutput.n195 CSoutput.n187 4.5005
R22809 CSoutput.n195 CSoutput.n191 4.5005
R22810 CSoutput.n195 CSoutput.n186 4.5005
R22811 CSoutput.n195 CSoutput.t168 4.5005
R22812 CSoutput.n195 CSoutput.n185 4.5005
R22813 CSoutput.n195 CSoutput.n192 4.5005
R22814 CSoutput.n241 CSoutput.n195 4.5005
R22815 CSoutput.n240 CSoutput.n188 4.5005
R22816 CSoutput.n240 CSoutput.n190 4.5005
R22817 CSoutput.n240 CSoutput.n187 4.5005
R22818 CSoutput.n240 CSoutput.n191 4.5005
R22819 CSoutput.n240 CSoutput.n186 4.5005
R22820 CSoutput.n240 CSoutput.t168 4.5005
R22821 CSoutput.n240 CSoutput.n185 4.5005
R22822 CSoutput.n240 CSoutput.n192 4.5005
R22823 CSoutput.n241 CSoutput.n240 4.5005
R22824 CSoutput.n239 CSoutput.n124 4.5005
R22825 CSoutput.n140 CSoutput.n124 4.5005
R22826 CSoutput.n135 CSoutput.n119 4.5005
R22827 CSoutput.n135 CSoutput.n121 4.5005
R22828 CSoutput.n135 CSoutput.n118 4.5005
R22829 CSoutput.n135 CSoutput.n122 4.5005
R22830 CSoutput.n135 CSoutput.n117 4.5005
R22831 CSoutput.n135 CSoutput.t175 4.5005
R22832 CSoutput.n135 CSoutput.n116 4.5005
R22833 CSoutput.n135 CSoutput.n123 4.5005
R22834 CSoutput.n135 CSoutput.n124 4.5005
R22835 CSoutput.n133 CSoutput.n119 4.5005
R22836 CSoutput.n133 CSoutput.n121 4.5005
R22837 CSoutput.n133 CSoutput.n118 4.5005
R22838 CSoutput.n133 CSoutput.n122 4.5005
R22839 CSoutput.n133 CSoutput.n117 4.5005
R22840 CSoutput.n133 CSoutput.t175 4.5005
R22841 CSoutput.n133 CSoutput.n116 4.5005
R22842 CSoutput.n133 CSoutput.n123 4.5005
R22843 CSoutput.n133 CSoutput.n124 4.5005
R22844 CSoutput.n132 CSoutput.n119 4.5005
R22845 CSoutput.n132 CSoutput.n121 4.5005
R22846 CSoutput.n132 CSoutput.n118 4.5005
R22847 CSoutput.n132 CSoutput.n122 4.5005
R22848 CSoutput.n132 CSoutput.n117 4.5005
R22849 CSoutput.n132 CSoutput.t175 4.5005
R22850 CSoutput.n132 CSoutput.n116 4.5005
R22851 CSoutput.n132 CSoutput.n123 4.5005
R22852 CSoutput.n132 CSoutput.n124 4.5005
R22853 CSoutput.n261 CSoutput.n119 4.5005
R22854 CSoutput.n261 CSoutput.n121 4.5005
R22855 CSoutput.n261 CSoutput.n118 4.5005
R22856 CSoutput.n261 CSoutput.n122 4.5005
R22857 CSoutput.n261 CSoutput.n117 4.5005
R22858 CSoutput.n261 CSoutput.t175 4.5005
R22859 CSoutput.n261 CSoutput.n116 4.5005
R22860 CSoutput.n261 CSoutput.n123 4.5005
R22861 CSoutput.n261 CSoutput.n124 4.5005
R22862 CSoutput.n259 CSoutput.n119 4.5005
R22863 CSoutput.n259 CSoutput.n121 4.5005
R22864 CSoutput.n259 CSoutput.n118 4.5005
R22865 CSoutput.n259 CSoutput.n122 4.5005
R22866 CSoutput.n259 CSoutput.n117 4.5005
R22867 CSoutput.n259 CSoutput.t175 4.5005
R22868 CSoutput.n259 CSoutput.n116 4.5005
R22869 CSoutput.n259 CSoutput.n123 4.5005
R22870 CSoutput.n257 CSoutput.n119 4.5005
R22871 CSoutput.n257 CSoutput.n121 4.5005
R22872 CSoutput.n257 CSoutput.n118 4.5005
R22873 CSoutput.n257 CSoutput.n122 4.5005
R22874 CSoutput.n257 CSoutput.n117 4.5005
R22875 CSoutput.n257 CSoutput.t175 4.5005
R22876 CSoutput.n257 CSoutput.n116 4.5005
R22877 CSoutput.n257 CSoutput.n123 4.5005
R22878 CSoutput.n143 CSoutput.n119 4.5005
R22879 CSoutput.n143 CSoutput.n121 4.5005
R22880 CSoutput.n143 CSoutput.n118 4.5005
R22881 CSoutput.n143 CSoutput.n122 4.5005
R22882 CSoutput.n143 CSoutput.n117 4.5005
R22883 CSoutput.n143 CSoutput.t175 4.5005
R22884 CSoutput.n143 CSoutput.n116 4.5005
R22885 CSoutput.n143 CSoutput.n123 4.5005
R22886 CSoutput.n143 CSoutput.n124 4.5005
R22887 CSoutput.n142 CSoutput.n119 4.5005
R22888 CSoutput.n142 CSoutput.n121 4.5005
R22889 CSoutput.n142 CSoutput.n118 4.5005
R22890 CSoutput.n142 CSoutput.n122 4.5005
R22891 CSoutput.n142 CSoutput.n117 4.5005
R22892 CSoutput.n142 CSoutput.t175 4.5005
R22893 CSoutput.n142 CSoutput.n116 4.5005
R22894 CSoutput.n142 CSoutput.n123 4.5005
R22895 CSoutput.n142 CSoutput.n124 4.5005
R22896 CSoutput.n146 CSoutput.n119 4.5005
R22897 CSoutput.n146 CSoutput.n121 4.5005
R22898 CSoutput.n146 CSoutput.n118 4.5005
R22899 CSoutput.n146 CSoutput.n122 4.5005
R22900 CSoutput.n146 CSoutput.n117 4.5005
R22901 CSoutput.n146 CSoutput.t175 4.5005
R22902 CSoutput.n146 CSoutput.n116 4.5005
R22903 CSoutput.n146 CSoutput.n123 4.5005
R22904 CSoutput.n146 CSoutput.n124 4.5005
R22905 CSoutput.n145 CSoutput.n119 4.5005
R22906 CSoutput.n145 CSoutput.n121 4.5005
R22907 CSoutput.n145 CSoutput.n118 4.5005
R22908 CSoutput.n145 CSoutput.n122 4.5005
R22909 CSoutput.n145 CSoutput.n117 4.5005
R22910 CSoutput.n145 CSoutput.t175 4.5005
R22911 CSoutput.n145 CSoutput.n116 4.5005
R22912 CSoutput.n145 CSoutput.n123 4.5005
R22913 CSoutput.n145 CSoutput.n124 4.5005
R22914 CSoutput.n128 CSoutput.n119 4.5005
R22915 CSoutput.n128 CSoutput.n121 4.5005
R22916 CSoutput.n128 CSoutput.n118 4.5005
R22917 CSoutput.n128 CSoutput.n122 4.5005
R22918 CSoutput.n128 CSoutput.n117 4.5005
R22919 CSoutput.n128 CSoutput.t175 4.5005
R22920 CSoutput.n128 CSoutput.n116 4.5005
R22921 CSoutput.n128 CSoutput.n123 4.5005
R22922 CSoutput.n128 CSoutput.n124 4.5005
R22923 CSoutput.n264 CSoutput.n119 4.5005
R22924 CSoutput.n264 CSoutput.n121 4.5005
R22925 CSoutput.n264 CSoutput.n118 4.5005
R22926 CSoutput.n264 CSoutput.n122 4.5005
R22927 CSoutput.n264 CSoutput.n117 4.5005
R22928 CSoutput.n264 CSoutput.t175 4.5005
R22929 CSoutput.n264 CSoutput.n116 4.5005
R22930 CSoutput.n264 CSoutput.n123 4.5005
R22931 CSoutput.n264 CSoutput.n124 4.5005
R22932 CSoutput.n299 CSoutput.n287 4.10845
R22933 CSoutput.n113 CSoutput.n101 4.10845
R22934 CSoutput.n297 CSoutput.t55 4.06363
R22935 CSoutput.n297 CSoutput.t6 4.06363
R22936 CSoutput.n295 CSoutput.t2 4.06363
R22937 CSoutput.n295 CSoutput.t31 4.06363
R22938 CSoutput.n293 CSoutput.t42 4.06363
R22939 CSoutput.n293 CSoutput.t57 4.06363
R22940 CSoutput.n291 CSoutput.t66 4.06363
R22941 CSoutput.n291 CSoutput.t15 4.06363
R22942 CSoutput.n289 CSoutput.t19 4.06363
R22943 CSoutput.n289 CSoutput.t58 4.06363
R22944 CSoutput.n288 CSoutput.t68 4.06363
R22945 CSoutput.n288 CSoutput.t69 4.06363
R22946 CSoutput.n285 CSoutput.t49 4.06363
R22947 CSoutput.n285 CSoutput.t70 4.06363
R22948 CSoutput.n283 CSoutput.t67 4.06363
R22949 CSoutput.n283 CSoutput.t24 4.06363
R22950 CSoutput.n281 CSoutput.t33 4.06363
R22951 CSoutput.n281 CSoutput.t50 4.06363
R22952 CSoutput.n279 CSoutput.t59 4.06363
R22953 CSoutput.n279 CSoutput.t5 4.06363
R22954 CSoutput.n277 CSoutput.t7 4.06363
R22955 CSoutput.n277 CSoutput.t53 4.06363
R22956 CSoutput.n276 CSoutput.t62 4.06363
R22957 CSoutput.n276 CSoutput.t63 4.06363
R22958 CSoutput.n274 CSoutput.t51 4.06363
R22959 CSoutput.n274 CSoutput.t22 4.06363
R22960 CSoutput.n272 CSoutput.t64 4.06363
R22961 CSoutput.n272 CSoutput.t37 4.06363
R22962 CSoutput.n270 CSoutput.t56 4.06363
R22963 CSoutput.n270 CSoutput.t28 4.06363
R22964 CSoutput.n268 CSoutput.t46 4.06363
R22965 CSoutput.n268 CSoutput.t14 4.06363
R22966 CSoutput.n266 CSoutput.t60 4.06363
R22967 CSoutput.n266 CSoutput.t9 4.06363
R22968 CSoutput.n265 CSoutput.t34 4.06363
R22969 CSoutput.n265 CSoutput.t20 4.06363
R22970 CSoutput.n102 CSoutput.t44 4.06363
R22971 CSoutput.n102 CSoutput.t27 4.06363
R22972 CSoutput.n103 CSoutput.t13 4.06363
R22973 CSoutput.n103 CSoutput.t45 4.06363
R22974 CSoutput.n105 CSoutput.t43 4.06363
R22975 CSoutput.n105 CSoutput.t25 4.06363
R22976 CSoutput.n107 CSoutput.t12 4.06363
R22977 CSoutput.n107 CSoutput.t11 4.06363
R22978 CSoutput.n109 CSoutput.t54 4.06363
R22979 CSoutput.n109 CSoutput.t32 4.06363
R22980 CSoutput.n111 CSoutput.t30 4.06363
R22981 CSoutput.n111 CSoutput.t8 4.06363
R22982 CSoutput.n90 CSoutput.t39 4.06363
R22983 CSoutput.n90 CSoutput.t18 4.06363
R22984 CSoutput.n91 CSoutput.t4 4.06363
R22985 CSoutput.n91 CSoutput.t40 4.06363
R22986 CSoutput.n93 CSoutput.t36 4.06363
R22987 CSoutput.n93 CSoutput.t16 4.06363
R22988 CSoutput.n95 CSoutput.t3 4.06363
R22989 CSoutput.n95 CSoutput.t1 4.06363
R22990 CSoutput.n97 CSoutput.t48 4.06363
R22991 CSoutput.n97 CSoutput.t26 4.06363
R22992 CSoutput.n99 CSoutput.t23 4.06363
R22993 CSoutput.n99 CSoutput.t0 4.06363
R22994 CSoutput.n79 CSoutput.t71 4.06363
R22995 CSoutput.n79 CSoutput.t35 4.06363
R22996 CSoutput.n80 CSoutput.t10 4.06363
R22997 CSoutput.n80 CSoutput.t61 4.06363
R22998 CSoutput.n82 CSoutput.t17 4.06363
R22999 CSoutput.n82 CSoutput.t47 4.06363
R23000 CSoutput.n84 CSoutput.t29 4.06363
R23001 CSoutput.n84 CSoutput.t41 4.06363
R23002 CSoutput.n86 CSoutput.t38 4.06363
R23003 CSoutput.n86 CSoutput.t65 4.06363
R23004 CSoutput.n88 CSoutput.t21 4.06363
R23005 CSoutput.n88 CSoutput.t52 4.06363
R23006 CSoutput.n44 CSoutput.n43 3.79402
R23007 CSoutput.n49 CSoutput.n48 3.79402
R23008 CSoutput.n347 CSoutput.n331 3.72967
R23009 CSoutput.n395 CSoutput.n379 3.72967
R23010 CSoutput.n397 CSoutput.n396 3.57343
R23011 CSoutput.n396 CSoutput.n348 3.08965
R23012 CSoutput.n345 CSoutput.t101 2.82907
R23013 CSoutput.n345 CSoutput.t91 2.82907
R23014 CSoutput.n343 CSoutput.t82 2.82907
R23015 CSoutput.n343 CSoutput.t152 2.82907
R23016 CSoutput.n341 CSoutput.t94 2.82907
R23017 CSoutput.n341 CSoutput.t98 2.82907
R23018 CSoutput.n339 CSoutput.t93 2.82907
R23019 CSoutput.n339 CSoutput.t167 2.82907
R23020 CSoutput.n337 CSoutput.t112 2.82907
R23021 CSoutput.n337 CSoutput.t85 2.82907
R23022 CSoutput.n335 CSoutput.t76 2.82907
R23023 CSoutput.n335 CSoutput.t141 2.82907
R23024 CSoutput.n333 CSoutput.t103 2.82907
R23025 CSoutput.n333 CSoutput.t107 2.82907
R23026 CSoutput.n332 CSoutput.t84 2.82907
R23027 CSoutput.n332 CSoutput.t156 2.82907
R23028 CSoutput.n329 CSoutput.t138 2.82907
R23029 CSoutput.n329 CSoutput.t119 2.82907
R23030 CSoutput.n327 CSoutput.t120 2.82907
R23031 CSoutput.n327 CSoutput.t126 2.82907
R23032 CSoutput.n325 CSoutput.t75 2.82907
R23033 CSoutput.n325 CSoutput.t139 2.82907
R23034 CSoutput.n323 CSoutput.t137 2.82907
R23035 CSoutput.n323 CSoutput.t118 2.82907
R23036 CSoutput.n321 CSoutput.t154 2.82907
R23037 CSoutput.n321 CSoutput.t73 2.82907
R23038 CSoutput.n319 CSoutput.t74 2.82907
R23039 CSoutput.n319 CSoutput.t146 2.82907
R23040 CSoutput.n317 CSoutput.t83 2.82907
R23041 CSoutput.n317 CSoutput.t153 2.82907
R23042 CSoutput.n316 CSoutput.t160 2.82907
R23043 CSoutput.n316 CSoutput.t72 2.82907
R23044 CSoutput.n314 CSoutput.t79 2.82907
R23045 CSoutput.n314 CSoutput.t102 2.82907
R23046 CSoutput.n312 CSoutput.t90 2.82907
R23047 CSoutput.n312 CSoutput.t115 2.82907
R23048 CSoutput.n310 CSoutput.t125 2.82907
R23049 CSoutput.n310 CSoutput.t135 2.82907
R23050 CSoutput.n308 CSoutput.t113 2.82907
R23051 CSoutput.n308 CSoutput.t155 2.82907
R23052 CSoutput.n306 CSoutput.t129 2.82907
R23053 CSoutput.n306 CSoutput.t106 2.82907
R23054 CSoutput.n304 CSoutput.t95 2.82907
R23055 CSoutput.n304 CSoutput.t114 2.82907
R23056 CSoutput.n302 CSoutput.t105 2.82907
R23057 CSoutput.n302 CSoutput.t110 2.82907
R23058 CSoutput.n301 CSoutput.t111 2.82907
R23059 CSoutput.n301 CSoutput.t164 2.82907
R23060 CSoutput.n380 CSoutput.t124 2.82907
R23061 CSoutput.n380 CSoutput.t149 2.82907
R23062 CSoutput.n381 CSoutput.t96 2.82907
R23063 CSoutput.n381 CSoutput.t109 2.82907
R23064 CSoutput.n383 CSoutput.t116 2.82907
R23065 CSoutput.n383 CSoutput.t130 2.82907
R23066 CSoutput.n385 CSoutput.t150 2.82907
R23067 CSoutput.n385 CSoutput.t121 2.82907
R23068 CSoutput.n387 CSoutput.t128 2.82907
R23069 CSoutput.n387 CSoutput.t161 2.82907
R23070 CSoutput.n389 CSoutput.t78 2.82907
R23071 CSoutput.n389 CSoutput.t99 2.82907
R23072 CSoutput.n391 CSoutput.t122 2.82907
R23073 CSoutput.n391 CSoutput.t144 2.82907
R23074 CSoutput.n393 CSoutput.t157 2.82907
R23075 CSoutput.n393 CSoutput.t86 2.82907
R23076 CSoutput.n364 CSoutput.t87 2.82907
R23077 CSoutput.n364 CSoutput.t80 2.82907
R23078 CSoutput.n365 CSoutput.t77 2.82907
R23079 CSoutput.n365 CSoutput.t165 2.82907
R23080 CSoutput.n367 CSoutput.t166 2.82907
R23081 CSoutput.n367 CSoutput.t88 2.82907
R23082 CSoutput.n369 CSoutput.t89 2.82907
R23083 CSoutput.n369 CSoutput.t131 2.82907
R23084 CSoutput.n371 CSoutput.t132 2.82907
R23085 CSoutput.n371 CSoutput.t159 2.82907
R23086 CSoutput.n373 CSoutput.t162 2.82907
R23087 CSoutput.n373 CSoutput.t151 2.82907
R23088 CSoutput.n375 CSoutput.t145 2.82907
R23089 CSoutput.n375 CSoutput.t133 2.82907
R23090 CSoutput.n377 CSoutput.t134 2.82907
R23091 CSoutput.n377 CSoutput.t163 2.82907
R23092 CSoutput.n349 CSoutput.t97 2.82907
R23093 CSoutput.n349 CSoutput.t140 2.82907
R23094 CSoutput.n350 CSoutput.t136 2.82907
R23095 CSoutput.n350 CSoutput.t117 2.82907
R23096 CSoutput.n352 CSoutput.t143 2.82907
R23097 CSoutput.n352 CSoutput.t108 2.82907
R23098 CSoutput.n354 CSoutput.t127 2.82907
R23099 CSoutput.n354 CSoutput.t158 2.82907
R23100 CSoutput.n356 CSoutput.t92 2.82907
R23101 CSoutput.n356 CSoutput.t142 2.82907
R23102 CSoutput.n358 CSoutput.t81 2.82907
R23103 CSoutput.n358 CSoutput.t148 2.82907
R23104 CSoutput.n360 CSoutput.t147 2.82907
R23105 CSoutput.n360 CSoutput.t104 2.82907
R23106 CSoutput.n362 CSoutput.t123 2.82907
R23107 CSoutput.n362 CSoutput.t100 2.82907
R23108 CSoutput.n300 CSoutput.n114 2.78353
R23109 CSoutput.n75 CSoutput.n1 2.45513
R23110 CSoutput.n205 CSoutput.n203 2.251
R23111 CSoutput.n205 CSoutput.n202 2.251
R23112 CSoutput.n205 CSoutput.n201 2.251
R23113 CSoutput.n205 CSoutput.n200 2.251
R23114 CSoutput.n174 CSoutput.n173 2.251
R23115 CSoutput.n174 CSoutput.n172 2.251
R23116 CSoutput.n174 CSoutput.n171 2.251
R23117 CSoutput.n174 CSoutput.n170 2.251
R23118 CSoutput.n247 CSoutput.n246 2.251
R23119 CSoutput.n212 CSoutput.n210 2.251
R23120 CSoutput.n212 CSoutput.n209 2.251
R23121 CSoutput.n212 CSoutput.n208 2.251
R23122 CSoutput.n230 CSoutput.n212 2.251
R23123 CSoutput.n218 CSoutput.n217 2.251
R23124 CSoutput.n218 CSoutput.n216 2.251
R23125 CSoutput.n218 CSoutput.n215 2.251
R23126 CSoutput.n218 CSoutput.n214 2.251
R23127 CSoutput.n244 CSoutput.n184 2.251
R23128 CSoutput.n239 CSoutput.n237 2.251
R23129 CSoutput.n239 CSoutput.n236 2.251
R23130 CSoutput.n239 CSoutput.n235 2.251
R23131 CSoutput.n239 CSoutput.n234 2.251
R23132 CSoutput.n140 CSoutput.n139 2.251
R23133 CSoutput.n140 CSoutput.n138 2.251
R23134 CSoutput.n140 CSoutput.n137 2.251
R23135 CSoutput.n140 CSoutput.n136 2.251
R23136 CSoutput.n257 CSoutput.n256 2.251
R23137 CSoutput.n174 CSoutput.n154 2.2505
R23138 CSoutput.n169 CSoutput.n154 2.2505
R23139 CSoutput.n167 CSoutput.n154 2.2505
R23140 CSoutput.n166 CSoutput.n154 2.2505
R23141 CSoutput.n251 CSoutput.n154 2.2505
R23142 CSoutput.n249 CSoutput.n154 2.2505
R23143 CSoutput.n247 CSoutput.n154 2.2505
R23144 CSoutput.n177 CSoutput.n154 2.2505
R23145 CSoutput.n176 CSoutput.n154 2.2505
R23146 CSoutput.n180 CSoutput.n154 2.2505
R23147 CSoutput.n179 CSoutput.n154 2.2505
R23148 CSoutput.n162 CSoutput.n154 2.2505
R23149 CSoutput.n254 CSoutput.n154 2.2505
R23150 CSoutput.n254 CSoutput.n253 2.2505
R23151 CSoutput.n218 CSoutput.n189 2.2505
R23152 CSoutput.n199 CSoutput.n189 2.2505
R23153 CSoutput.n220 CSoutput.n189 2.2505
R23154 CSoutput.n198 CSoutput.n189 2.2505
R23155 CSoutput.n222 CSoutput.n189 2.2505
R23156 CSoutput.n189 CSoutput.n183 2.2505
R23157 CSoutput.n244 CSoutput.n189 2.2505
R23158 CSoutput.n242 CSoutput.n189 2.2505
R23159 CSoutput.n224 CSoutput.n189 2.2505
R23160 CSoutput.n196 CSoutput.n189 2.2505
R23161 CSoutput.n226 CSoutput.n189 2.2505
R23162 CSoutput.n195 CSoutput.n189 2.2505
R23163 CSoutput.n240 CSoutput.n189 2.2505
R23164 CSoutput.n240 CSoutput.n193 2.2505
R23165 CSoutput.n140 CSoutput.n120 2.2505
R23166 CSoutput.n135 CSoutput.n120 2.2505
R23167 CSoutput.n133 CSoutput.n120 2.2505
R23168 CSoutput.n132 CSoutput.n120 2.2505
R23169 CSoutput.n261 CSoutput.n120 2.2505
R23170 CSoutput.n259 CSoutput.n120 2.2505
R23171 CSoutput.n257 CSoutput.n120 2.2505
R23172 CSoutput.n143 CSoutput.n120 2.2505
R23173 CSoutput.n142 CSoutput.n120 2.2505
R23174 CSoutput.n146 CSoutput.n120 2.2505
R23175 CSoutput.n145 CSoutput.n120 2.2505
R23176 CSoutput.n128 CSoutput.n120 2.2505
R23177 CSoutput.n264 CSoutput.n120 2.2505
R23178 CSoutput.n264 CSoutput.n263 2.2505
R23179 CSoutput.n182 CSoutput.n175 2.25024
R23180 CSoutput.n182 CSoutput.n168 2.25024
R23181 CSoutput.n250 CSoutput.n182 2.25024
R23182 CSoutput.n182 CSoutput.n178 2.25024
R23183 CSoutput.n182 CSoutput.n181 2.25024
R23184 CSoutput.n182 CSoutput.n149 2.25024
R23185 CSoutput.n232 CSoutput.n229 2.25024
R23186 CSoutput.n232 CSoutput.n228 2.25024
R23187 CSoutput.n232 CSoutput.n227 2.25024
R23188 CSoutput.n232 CSoutput.n194 2.25024
R23189 CSoutput.n232 CSoutput.n231 2.25024
R23190 CSoutput.n233 CSoutput.n232 2.25024
R23191 CSoutput.n148 CSoutput.n141 2.25024
R23192 CSoutput.n148 CSoutput.n134 2.25024
R23193 CSoutput.n260 CSoutput.n148 2.25024
R23194 CSoutput.n148 CSoutput.n144 2.25024
R23195 CSoutput.n148 CSoutput.n147 2.25024
R23196 CSoutput.n148 CSoutput.n115 2.25024
R23197 CSoutput.n249 CSoutput.n159 1.50111
R23198 CSoutput.n197 CSoutput.n183 1.50111
R23199 CSoutput.n259 CSoutput.n125 1.50111
R23200 CSoutput.n205 CSoutput.n204 1.501
R23201 CSoutput.n212 CSoutput.n211 1.501
R23202 CSoutput.n239 CSoutput.n238 1.501
R23203 CSoutput.n253 CSoutput.n164 1.12536
R23204 CSoutput.n253 CSoutput.n165 1.12536
R23205 CSoutput.n253 CSoutput.n252 1.12536
R23206 CSoutput.n213 CSoutput.n193 1.12536
R23207 CSoutput.n219 CSoutput.n193 1.12536
R23208 CSoutput.n221 CSoutput.n193 1.12536
R23209 CSoutput.n263 CSoutput.n130 1.12536
R23210 CSoutput.n263 CSoutput.n131 1.12536
R23211 CSoutput.n263 CSoutput.n262 1.12536
R23212 CSoutput.n253 CSoutput.n160 1.12536
R23213 CSoutput.n253 CSoutput.n161 1.12536
R23214 CSoutput.n253 CSoutput.n163 1.12536
R23215 CSoutput.n243 CSoutput.n193 1.12536
R23216 CSoutput.n223 CSoutput.n193 1.12536
R23217 CSoutput.n225 CSoutput.n193 1.12536
R23218 CSoutput.n263 CSoutput.n126 1.12536
R23219 CSoutput.n263 CSoutput.n127 1.12536
R23220 CSoutput.n263 CSoutput.n129 1.12536
R23221 CSoutput.n31 CSoutput.n30 0.669944
R23222 CSoutput.n62 CSoutput.n61 0.669944
R23223 CSoutput.n336 CSoutput.n334 0.573776
R23224 CSoutput.n338 CSoutput.n336 0.573776
R23225 CSoutput.n340 CSoutput.n338 0.573776
R23226 CSoutput.n342 CSoutput.n340 0.573776
R23227 CSoutput.n344 CSoutput.n342 0.573776
R23228 CSoutput.n346 CSoutput.n344 0.573776
R23229 CSoutput.n320 CSoutput.n318 0.573776
R23230 CSoutput.n322 CSoutput.n320 0.573776
R23231 CSoutput.n324 CSoutput.n322 0.573776
R23232 CSoutput.n326 CSoutput.n324 0.573776
R23233 CSoutput.n328 CSoutput.n326 0.573776
R23234 CSoutput.n330 CSoutput.n328 0.573776
R23235 CSoutput.n305 CSoutput.n303 0.573776
R23236 CSoutput.n307 CSoutput.n305 0.573776
R23237 CSoutput.n309 CSoutput.n307 0.573776
R23238 CSoutput.n311 CSoutput.n309 0.573776
R23239 CSoutput.n313 CSoutput.n311 0.573776
R23240 CSoutput.n315 CSoutput.n313 0.573776
R23241 CSoutput.n394 CSoutput.n392 0.573776
R23242 CSoutput.n392 CSoutput.n390 0.573776
R23243 CSoutput.n390 CSoutput.n388 0.573776
R23244 CSoutput.n388 CSoutput.n386 0.573776
R23245 CSoutput.n386 CSoutput.n384 0.573776
R23246 CSoutput.n384 CSoutput.n382 0.573776
R23247 CSoutput.n378 CSoutput.n376 0.573776
R23248 CSoutput.n376 CSoutput.n374 0.573776
R23249 CSoutput.n374 CSoutput.n372 0.573776
R23250 CSoutput.n372 CSoutput.n370 0.573776
R23251 CSoutput.n370 CSoutput.n368 0.573776
R23252 CSoutput.n368 CSoutput.n366 0.573776
R23253 CSoutput.n363 CSoutput.n361 0.573776
R23254 CSoutput.n361 CSoutput.n359 0.573776
R23255 CSoutput.n359 CSoutput.n357 0.573776
R23256 CSoutput.n357 CSoutput.n355 0.573776
R23257 CSoutput.n355 CSoutput.n353 0.573776
R23258 CSoutput.n353 CSoutput.n351 0.573776
R23259 CSoutput.n397 CSoutput.n264 0.53442
R23260 CSoutput.n292 CSoutput.n290 0.358259
R23261 CSoutput.n294 CSoutput.n292 0.358259
R23262 CSoutput.n296 CSoutput.n294 0.358259
R23263 CSoutput.n298 CSoutput.n296 0.358259
R23264 CSoutput.n280 CSoutput.n278 0.358259
R23265 CSoutput.n282 CSoutput.n280 0.358259
R23266 CSoutput.n284 CSoutput.n282 0.358259
R23267 CSoutput.n286 CSoutput.n284 0.358259
R23268 CSoutput.n269 CSoutput.n267 0.358259
R23269 CSoutput.n271 CSoutput.n269 0.358259
R23270 CSoutput.n273 CSoutput.n271 0.358259
R23271 CSoutput.n275 CSoutput.n273 0.358259
R23272 CSoutput.n112 CSoutput.n110 0.358259
R23273 CSoutput.n110 CSoutput.n108 0.358259
R23274 CSoutput.n108 CSoutput.n106 0.358259
R23275 CSoutput.n106 CSoutput.n104 0.358259
R23276 CSoutput.n100 CSoutput.n98 0.358259
R23277 CSoutput.n98 CSoutput.n96 0.358259
R23278 CSoutput.n96 CSoutput.n94 0.358259
R23279 CSoutput.n94 CSoutput.n92 0.358259
R23280 CSoutput.n89 CSoutput.n87 0.358259
R23281 CSoutput.n87 CSoutput.n85 0.358259
R23282 CSoutput.n85 CSoutput.n83 0.358259
R23283 CSoutput.n83 CSoutput.n81 0.358259
R23284 CSoutput.n21 CSoutput.n20 0.169105
R23285 CSoutput.n21 CSoutput.n16 0.169105
R23286 CSoutput.n26 CSoutput.n16 0.169105
R23287 CSoutput.n27 CSoutput.n26 0.169105
R23288 CSoutput.n27 CSoutput.n14 0.169105
R23289 CSoutput.n32 CSoutput.n14 0.169105
R23290 CSoutput.n33 CSoutput.n32 0.169105
R23291 CSoutput.n34 CSoutput.n33 0.169105
R23292 CSoutput.n34 CSoutput.n12 0.169105
R23293 CSoutput.n39 CSoutput.n12 0.169105
R23294 CSoutput.n40 CSoutput.n39 0.169105
R23295 CSoutput.n40 CSoutput.n10 0.169105
R23296 CSoutput.n45 CSoutput.n10 0.169105
R23297 CSoutput.n46 CSoutput.n45 0.169105
R23298 CSoutput.n47 CSoutput.n46 0.169105
R23299 CSoutput.n47 CSoutput.n8 0.169105
R23300 CSoutput.n52 CSoutput.n8 0.169105
R23301 CSoutput.n53 CSoutput.n52 0.169105
R23302 CSoutput.n53 CSoutput.n6 0.169105
R23303 CSoutput.n58 CSoutput.n6 0.169105
R23304 CSoutput.n59 CSoutput.n58 0.169105
R23305 CSoutput.n60 CSoutput.n59 0.169105
R23306 CSoutput.n60 CSoutput.n4 0.169105
R23307 CSoutput.n66 CSoutput.n4 0.169105
R23308 CSoutput.n67 CSoutput.n66 0.169105
R23309 CSoutput.n68 CSoutput.n67 0.169105
R23310 CSoutput.n68 CSoutput.n2 0.169105
R23311 CSoutput.n73 CSoutput.n2 0.169105
R23312 CSoutput.n74 CSoutput.n73 0.169105
R23313 CSoutput.n74 CSoutput.n0 0.169105
R23314 CSoutput.n78 CSoutput.n0 0.169105
R23315 CSoutput.n207 CSoutput.n206 0.0910737
R23316 CSoutput.n258 CSoutput.n255 0.0723685
R23317 CSoutput.n212 CSoutput.n207 0.0522944
R23318 CSoutput.n255 CSoutput.n254 0.0499135
R23319 CSoutput.n206 CSoutput.n205 0.0499135
R23320 CSoutput.n240 CSoutput.n239 0.0464294
R23321 CSoutput.n248 CSoutput.n245 0.0391444
R23322 CSoutput.n207 CSoutput.t178 0.023435
R23323 CSoutput.n255 CSoutput.t170 0.02262
R23324 CSoutput.n206 CSoutput.t172 0.02262
R23325 CSoutput CSoutput.n397 0.0052
R23326 CSoutput.n177 CSoutput.n160 0.00365111
R23327 CSoutput.n180 CSoutput.n161 0.00365111
R23328 CSoutput.n163 CSoutput.n162 0.00365111
R23329 CSoutput.n205 CSoutput.n164 0.00365111
R23330 CSoutput.n169 CSoutput.n165 0.00365111
R23331 CSoutput.n252 CSoutput.n166 0.00365111
R23332 CSoutput.n243 CSoutput.n242 0.00365111
R23333 CSoutput.n223 CSoutput.n196 0.00365111
R23334 CSoutput.n225 CSoutput.n195 0.00365111
R23335 CSoutput.n213 CSoutput.n212 0.00365111
R23336 CSoutput.n219 CSoutput.n199 0.00365111
R23337 CSoutput.n221 CSoutput.n198 0.00365111
R23338 CSoutput.n143 CSoutput.n126 0.00365111
R23339 CSoutput.n146 CSoutput.n127 0.00365111
R23340 CSoutput.n129 CSoutput.n128 0.00365111
R23341 CSoutput.n239 CSoutput.n130 0.00365111
R23342 CSoutput.n135 CSoutput.n131 0.00365111
R23343 CSoutput.n262 CSoutput.n132 0.00365111
R23344 CSoutput.n174 CSoutput.n164 0.00340054
R23345 CSoutput.n167 CSoutput.n165 0.00340054
R23346 CSoutput.n252 CSoutput.n251 0.00340054
R23347 CSoutput.n247 CSoutput.n160 0.00340054
R23348 CSoutput.n176 CSoutput.n161 0.00340054
R23349 CSoutput.n179 CSoutput.n163 0.00340054
R23350 CSoutput.n218 CSoutput.n213 0.00340054
R23351 CSoutput.n220 CSoutput.n219 0.00340054
R23352 CSoutput.n222 CSoutput.n221 0.00340054
R23353 CSoutput.n244 CSoutput.n243 0.00340054
R23354 CSoutput.n224 CSoutput.n223 0.00340054
R23355 CSoutput.n226 CSoutput.n225 0.00340054
R23356 CSoutput.n140 CSoutput.n130 0.00340054
R23357 CSoutput.n133 CSoutput.n131 0.00340054
R23358 CSoutput.n262 CSoutput.n261 0.00340054
R23359 CSoutput.n257 CSoutput.n126 0.00340054
R23360 CSoutput.n142 CSoutput.n127 0.00340054
R23361 CSoutput.n145 CSoutput.n129 0.00340054
R23362 CSoutput.n175 CSoutput.n169 0.00252698
R23363 CSoutput.n168 CSoutput.n166 0.00252698
R23364 CSoutput.n250 CSoutput.n249 0.00252698
R23365 CSoutput.n178 CSoutput.n176 0.00252698
R23366 CSoutput.n181 CSoutput.n179 0.00252698
R23367 CSoutput.n254 CSoutput.n149 0.00252698
R23368 CSoutput.n175 CSoutput.n174 0.00252698
R23369 CSoutput.n168 CSoutput.n167 0.00252698
R23370 CSoutput.n251 CSoutput.n250 0.00252698
R23371 CSoutput.n178 CSoutput.n177 0.00252698
R23372 CSoutput.n181 CSoutput.n180 0.00252698
R23373 CSoutput.n162 CSoutput.n149 0.00252698
R23374 CSoutput.n229 CSoutput.n199 0.00252698
R23375 CSoutput.n228 CSoutput.n198 0.00252698
R23376 CSoutput.n227 CSoutput.n183 0.00252698
R23377 CSoutput.n224 CSoutput.n194 0.00252698
R23378 CSoutput.n231 CSoutput.n226 0.00252698
R23379 CSoutput.n240 CSoutput.n233 0.00252698
R23380 CSoutput.n229 CSoutput.n218 0.00252698
R23381 CSoutput.n228 CSoutput.n220 0.00252698
R23382 CSoutput.n227 CSoutput.n222 0.00252698
R23383 CSoutput.n242 CSoutput.n194 0.00252698
R23384 CSoutput.n231 CSoutput.n196 0.00252698
R23385 CSoutput.n233 CSoutput.n195 0.00252698
R23386 CSoutput.n141 CSoutput.n135 0.00252698
R23387 CSoutput.n134 CSoutput.n132 0.00252698
R23388 CSoutput.n260 CSoutput.n259 0.00252698
R23389 CSoutput.n144 CSoutput.n142 0.00252698
R23390 CSoutput.n147 CSoutput.n145 0.00252698
R23391 CSoutput.n264 CSoutput.n115 0.00252698
R23392 CSoutput.n141 CSoutput.n140 0.00252698
R23393 CSoutput.n134 CSoutput.n133 0.00252698
R23394 CSoutput.n261 CSoutput.n260 0.00252698
R23395 CSoutput.n144 CSoutput.n143 0.00252698
R23396 CSoutput.n147 CSoutput.n146 0.00252698
R23397 CSoutput.n128 CSoutput.n115 0.00252698
R23398 CSoutput.n249 CSoutput.n248 0.0020275
R23399 CSoutput.n248 CSoutput.n247 0.0020275
R23400 CSoutput.n245 CSoutput.n183 0.0020275
R23401 CSoutput.n245 CSoutput.n244 0.0020275
R23402 CSoutput.n259 CSoutput.n258 0.0020275
R23403 CSoutput.n258 CSoutput.n257 0.0020275
R23404 CSoutput.n159 CSoutput.n158 0.00166668
R23405 CSoutput.n241 CSoutput.n197 0.00166668
R23406 CSoutput.n125 CSoutput.n124 0.00166668
R23407 CSoutput.n263 CSoutput.n125 0.00133328
R23408 CSoutput.n197 CSoutput.n193 0.00133328
R23409 CSoutput.n253 CSoutput.n159 0.00133328
R23410 CSoutput.n256 CSoutput.n148 0.001
R23411 CSoutput.n234 CSoutput.n148 0.001
R23412 CSoutput.n136 CSoutput.n116 0.001
R23413 CSoutput.n235 CSoutput.n116 0.001
R23414 CSoutput.n137 CSoutput.n117 0.001
R23415 CSoutput.n236 CSoutput.n117 0.001
R23416 CSoutput.n138 CSoutput.n118 0.001
R23417 CSoutput.n237 CSoutput.n118 0.001
R23418 CSoutput.n139 CSoutput.n119 0.001
R23419 CSoutput.n238 CSoutput.n119 0.001
R23420 CSoutput.n232 CSoutput.n184 0.001
R23421 CSoutput.n232 CSoutput.n230 0.001
R23422 CSoutput.n214 CSoutput.n185 0.001
R23423 CSoutput.n208 CSoutput.n185 0.001
R23424 CSoutput.n215 CSoutput.n186 0.001
R23425 CSoutput.n209 CSoutput.n186 0.001
R23426 CSoutput.n216 CSoutput.n187 0.001
R23427 CSoutput.n210 CSoutput.n187 0.001
R23428 CSoutput.n217 CSoutput.n188 0.001
R23429 CSoutput.n211 CSoutput.n188 0.001
R23430 CSoutput.n246 CSoutput.n182 0.001
R23431 CSoutput.n200 CSoutput.n182 0.001
R23432 CSoutput.n170 CSoutput.n150 0.001
R23433 CSoutput.n201 CSoutput.n150 0.001
R23434 CSoutput.n171 CSoutput.n151 0.001
R23435 CSoutput.n202 CSoutput.n151 0.001
R23436 CSoutput.n172 CSoutput.n152 0.001
R23437 CSoutput.n203 CSoutput.n152 0.001
R23438 CSoutput.n173 CSoutput.n153 0.001
R23439 CSoutput.n204 CSoutput.n153 0.001
R23440 CSoutput.n204 CSoutput.n154 0.001
R23441 CSoutput.n203 CSoutput.n155 0.001
R23442 CSoutput.n202 CSoutput.n156 0.001
R23443 CSoutput.n201 CSoutput.t189 0.001
R23444 CSoutput.n200 CSoutput.n157 0.001
R23445 CSoutput.n173 CSoutput.n155 0.001
R23446 CSoutput.n172 CSoutput.n156 0.001
R23447 CSoutput.n171 CSoutput.t189 0.001
R23448 CSoutput.n170 CSoutput.n157 0.001
R23449 CSoutput.n246 CSoutput.n158 0.001
R23450 CSoutput.n211 CSoutput.n189 0.001
R23451 CSoutput.n210 CSoutput.n190 0.001
R23452 CSoutput.n209 CSoutput.n191 0.001
R23453 CSoutput.n208 CSoutput.t168 0.001
R23454 CSoutput.n230 CSoutput.n192 0.001
R23455 CSoutput.n217 CSoutput.n190 0.001
R23456 CSoutput.n216 CSoutput.n191 0.001
R23457 CSoutput.n215 CSoutput.t168 0.001
R23458 CSoutput.n214 CSoutput.n192 0.001
R23459 CSoutput.n241 CSoutput.n184 0.001
R23460 CSoutput.n238 CSoutput.n120 0.001
R23461 CSoutput.n237 CSoutput.n121 0.001
R23462 CSoutput.n236 CSoutput.n122 0.001
R23463 CSoutput.n235 CSoutput.t175 0.001
R23464 CSoutput.n234 CSoutput.n123 0.001
R23465 CSoutput.n139 CSoutput.n121 0.001
R23466 CSoutput.n138 CSoutput.n122 0.001
R23467 CSoutput.n137 CSoutput.t175 0.001
R23468 CSoutput.n136 CSoutput.n123 0.001
R23469 CSoutput.n256 CSoutput.n124 0.001
R23470 a_n2982_8322.n12 a_n2982_8322.t27 74.6477
R23471 a_n2982_8322.n1 a_n2982_8322.t6 74.6477
R23472 a_n2982_8322.n28 a_n2982_8322.t21 74.6474
R23473 a_n2982_8322.n20 a_n2982_8322.t1 74.2899
R23474 a_n2982_8322.n13 a_n2982_8322.t25 74.2899
R23475 a_n2982_8322.n14 a_n2982_8322.t28 74.2899
R23476 a_n2982_8322.n17 a_n2982_8322.t29 74.2899
R23477 a_n2982_8322.n10 a_n2982_8322.t0 74.2899
R23478 a_n2982_8322.n28 a_n2982_8322.n27 70.6783
R23479 a_n2982_8322.n26 a_n2982_8322.n25 70.6783
R23480 a_n2982_8322.n24 a_n2982_8322.n23 70.6783
R23481 a_n2982_8322.n22 a_n2982_8322.n21 70.6783
R23482 a_n2982_8322.n12 a_n2982_8322.n11 70.6783
R23483 a_n2982_8322.n16 a_n2982_8322.n15 70.6783
R23484 a_n2982_8322.n1 a_n2982_8322.n0 70.6783
R23485 a_n2982_8322.n3 a_n2982_8322.n2 70.6783
R23486 a_n2982_8322.n5 a_n2982_8322.n4 70.6783
R23487 a_n2982_8322.n7 a_n2982_8322.n6 70.6783
R23488 a_n2982_8322.n9 a_n2982_8322.n8 70.6783
R23489 a_n2982_8322.n30 a_n2982_8322.n29 70.6782
R23490 a_n2982_8322.n18 a_n2982_8322.n10 24.9022
R23491 a_n2982_8322.n19 a_n2982_8322.t33 9.65181
R23492 a_n2982_8322.n18 a_n2982_8322.n17 8.38735
R23493 a_n2982_8322.n20 a_n2982_8322.n19 6.90998
R23494 a_n2982_8322.n19 a_n2982_8322.n18 5.3452
R23495 a_n2982_8322.n27 a_n2982_8322.t14 3.61217
R23496 a_n2982_8322.n27 a_n2982_8322.t10 3.61217
R23497 a_n2982_8322.n25 a_n2982_8322.t20 3.61217
R23498 a_n2982_8322.n25 a_n2982_8322.t8 3.61217
R23499 a_n2982_8322.n23 a_n2982_8322.t5 3.61217
R23500 a_n2982_8322.n23 a_n2982_8322.t4 3.61217
R23501 a_n2982_8322.n21 a_n2982_8322.t18 3.61217
R23502 a_n2982_8322.n21 a_n2982_8322.t17 3.61217
R23503 a_n2982_8322.n11 a_n2982_8322.t31 3.61217
R23504 a_n2982_8322.n11 a_n2982_8322.t30 3.61217
R23505 a_n2982_8322.n15 a_n2982_8322.t26 3.61217
R23506 a_n2982_8322.n15 a_n2982_8322.t24 3.61217
R23507 a_n2982_8322.n0 a_n2982_8322.t19 3.61217
R23508 a_n2982_8322.n0 a_n2982_8322.t15 3.61217
R23509 a_n2982_8322.n2 a_n2982_8322.t22 3.61217
R23510 a_n2982_8322.n2 a_n2982_8322.t12 3.61217
R23511 a_n2982_8322.n4 a_n2982_8322.t3 3.61217
R23512 a_n2982_8322.n4 a_n2982_8322.t2 3.61217
R23513 a_n2982_8322.n6 a_n2982_8322.t16 3.61217
R23514 a_n2982_8322.n6 a_n2982_8322.t9 3.61217
R23515 a_n2982_8322.n8 a_n2982_8322.t13 3.61217
R23516 a_n2982_8322.n8 a_n2982_8322.t11 3.61217
R23517 a_n2982_8322.n30 a_n2982_8322.t7 3.61217
R23518 a_n2982_8322.t23 a_n2982_8322.n30 3.61217
R23519 a_n2982_8322.n17 a_n2982_8322.n16 0.358259
R23520 a_n2982_8322.n16 a_n2982_8322.n14 0.358259
R23521 a_n2982_8322.n13 a_n2982_8322.n12 0.358259
R23522 a_n2982_8322.n10 a_n2982_8322.n9 0.358259
R23523 a_n2982_8322.n9 a_n2982_8322.n7 0.358259
R23524 a_n2982_8322.n7 a_n2982_8322.n5 0.358259
R23525 a_n2982_8322.n5 a_n2982_8322.n3 0.358259
R23526 a_n2982_8322.n3 a_n2982_8322.n1 0.358259
R23527 a_n2982_8322.n22 a_n2982_8322.n20 0.358259
R23528 a_n2982_8322.n24 a_n2982_8322.n22 0.358259
R23529 a_n2982_8322.n26 a_n2982_8322.n24 0.358259
R23530 a_n2982_8322.n29 a_n2982_8322.n26 0.358259
R23531 a_n2982_8322.n29 a_n2982_8322.n28 0.358259
R23532 a_n2982_8322.n14 a_n2982_8322.n13 0.101793
R23533 a_n2982_8322.t36 a_n2982_8322.t34 0.0788333
R23534 a_n2982_8322.t32 a_n2982_8322.t37 0.0788333
R23535 a_n2982_8322.t33 a_n2982_8322.t35 0.0788333
R23536 a_n2982_8322.t32 a_n2982_8322.t36 0.0318333
R23537 a_n2982_8322.t33 a_n2982_8322.t37 0.0318333
R23538 a_n2982_8322.t34 a_n2982_8322.t37 0.0318333
R23539 a_n2982_8322.t35 a_n2982_8322.t32 0.0318333
R23540 minus.n53 minus.t28 323.478
R23541 minus.n11 minus.t8 323.478
R23542 minus.n82 minus.t13 297.12
R23543 minus.n80 minus.t15 297.12
R23544 minus.n44 minus.t5 297.12
R23545 minus.n74 minus.t6 297.12
R23546 minus.n46 minus.t26 297.12
R23547 minus.n68 minus.t21 297.12
R23548 minus.n48 minus.t23 297.12
R23549 minus.n62 minus.t16 297.12
R23550 minus.n50 minus.t17 297.12
R23551 minus.n56 minus.t9 297.12
R23552 minus.n52 minus.t27 297.12
R23553 minus.n10 minus.t7 297.12
R23554 minus.n14 minus.t11 297.12
R23555 minus.n16 minus.t10 297.12
R23556 minus.n20 minus.t12 297.12
R23557 minus.n22 minus.t20 297.12
R23558 minus.n26 minus.t18 297.12
R23559 minus.n28 minus.t25 297.12
R23560 minus.n32 minus.t24 297.12
R23561 minus.n34 minus.t14 297.12
R23562 minus.n38 minus.t22 297.12
R23563 minus.n40 minus.t19 297.12
R23564 minus.n88 minus.t2 243.255
R23565 minus.n87 minus.n85 224.169
R23566 minus.n87 minus.n86 223.454
R23567 minus.n55 minus.n54 161.3
R23568 minus.n56 minus.n51 161.3
R23569 minus.n58 minus.n57 161.3
R23570 minus.n59 minus.n50 161.3
R23571 minus.n61 minus.n60 161.3
R23572 minus.n62 minus.n49 161.3
R23573 minus.n64 minus.n63 161.3
R23574 minus.n65 minus.n48 161.3
R23575 minus.n67 minus.n66 161.3
R23576 minus.n68 minus.n47 161.3
R23577 minus.n70 minus.n69 161.3
R23578 minus.n71 minus.n46 161.3
R23579 minus.n73 minus.n72 161.3
R23580 minus.n74 minus.n45 161.3
R23581 minus.n76 minus.n75 161.3
R23582 minus.n77 minus.n44 161.3
R23583 minus.n79 minus.n78 161.3
R23584 minus.n80 minus.n43 161.3
R23585 minus.n81 minus.n42 161.3
R23586 minus.n83 minus.n82 161.3
R23587 minus.n41 minus.n40 161.3
R23588 minus.n39 minus.n0 161.3
R23589 minus.n38 minus.n37 161.3
R23590 minus.n36 minus.n1 161.3
R23591 minus.n35 minus.n34 161.3
R23592 minus.n33 minus.n2 161.3
R23593 minus.n32 minus.n31 161.3
R23594 minus.n30 minus.n3 161.3
R23595 minus.n29 minus.n28 161.3
R23596 minus.n27 minus.n4 161.3
R23597 minus.n26 minus.n25 161.3
R23598 minus.n24 minus.n5 161.3
R23599 minus.n23 minus.n22 161.3
R23600 minus.n21 minus.n6 161.3
R23601 minus.n20 minus.n19 161.3
R23602 minus.n18 minus.n7 161.3
R23603 minus.n17 minus.n16 161.3
R23604 minus.n15 minus.n8 161.3
R23605 minus.n14 minus.n13 161.3
R23606 minus.n12 minus.n9 161.3
R23607 minus.n82 minus.n81 46.0096
R23608 minus.n40 minus.n39 46.0096
R23609 minus.n12 minus.n11 45.0871
R23610 minus.n54 minus.n53 45.0871
R23611 minus.n80 minus.n79 41.6278
R23612 minus.n55 minus.n52 41.6278
R23613 minus.n10 minus.n9 41.6278
R23614 minus.n38 minus.n1 41.6278
R23615 minus.n75 minus.n44 37.246
R23616 minus.n57 minus.n56 37.246
R23617 minus.n15 minus.n14 37.246
R23618 minus.n34 minus.n33 37.246
R23619 minus.n84 minus.n83 33.3925
R23620 minus.n74 minus.n73 32.8641
R23621 minus.n61 minus.n50 32.8641
R23622 minus.n16 minus.n7 32.8641
R23623 minus.n32 minus.n3 32.8641
R23624 minus.n69 minus.n46 28.4823
R23625 minus.n63 minus.n62 28.4823
R23626 minus.n21 minus.n20 28.4823
R23627 minus.n28 minus.n27 28.4823
R23628 minus.n68 minus.n67 24.1005
R23629 minus.n67 minus.n48 24.1005
R23630 minus.n22 minus.n5 24.1005
R23631 minus.n26 minus.n5 24.1005
R23632 minus.n86 minus.t4 19.8005
R23633 minus.n86 minus.t3 19.8005
R23634 minus.n85 minus.t1 19.8005
R23635 minus.n85 minus.t0 19.8005
R23636 minus.n69 minus.n68 19.7187
R23637 minus.n63 minus.n48 19.7187
R23638 minus.n22 minus.n21 19.7187
R23639 minus.n27 minus.n26 19.7187
R23640 minus.n73 minus.n46 15.3369
R23641 minus.n62 minus.n61 15.3369
R23642 minus.n20 minus.n7 15.3369
R23643 minus.n28 minus.n3 15.3369
R23644 minus.n53 minus.n52 14.1472
R23645 minus.n11 minus.n10 14.1472
R23646 minus.n84 minus.n41 12.0933
R23647 minus minus.n89 11.4112
R23648 minus.n75 minus.n74 10.955
R23649 minus.n57 minus.n50 10.955
R23650 minus.n16 minus.n15 10.955
R23651 minus.n33 minus.n32 10.955
R23652 minus.n79 minus.n44 6.57323
R23653 minus.n56 minus.n55 6.57323
R23654 minus.n14 minus.n9 6.57323
R23655 minus.n34 minus.n1 6.57323
R23656 minus.n89 minus.n88 4.80222
R23657 minus.n81 minus.n80 2.19141
R23658 minus.n39 minus.n38 2.19141
R23659 minus.n89 minus.n84 0.972091
R23660 minus.n88 minus.n87 0.716017
R23661 minus.n83 minus.n42 0.189894
R23662 minus.n43 minus.n42 0.189894
R23663 minus.n78 minus.n43 0.189894
R23664 minus.n78 minus.n77 0.189894
R23665 minus.n77 minus.n76 0.189894
R23666 minus.n76 minus.n45 0.189894
R23667 minus.n72 minus.n45 0.189894
R23668 minus.n72 minus.n71 0.189894
R23669 minus.n71 minus.n70 0.189894
R23670 minus.n70 minus.n47 0.189894
R23671 minus.n66 minus.n47 0.189894
R23672 minus.n66 minus.n65 0.189894
R23673 minus.n65 minus.n64 0.189894
R23674 minus.n64 minus.n49 0.189894
R23675 minus.n60 minus.n49 0.189894
R23676 minus.n60 minus.n59 0.189894
R23677 minus.n59 minus.n58 0.189894
R23678 minus.n58 minus.n51 0.189894
R23679 minus.n54 minus.n51 0.189894
R23680 minus.n13 minus.n12 0.189894
R23681 minus.n13 minus.n8 0.189894
R23682 minus.n17 minus.n8 0.189894
R23683 minus.n18 minus.n17 0.189894
R23684 minus.n19 minus.n18 0.189894
R23685 minus.n19 minus.n6 0.189894
R23686 minus.n23 minus.n6 0.189894
R23687 minus.n24 minus.n23 0.189894
R23688 minus.n25 minus.n24 0.189894
R23689 minus.n25 minus.n4 0.189894
R23690 minus.n29 minus.n4 0.189894
R23691 minus.n30 minus.n29 0.189894
R23692 minus.n31 minus.n30 0.189894
R23693 minus.n31 minus.n2 0.189894
R23694 minus.n35 minus.n2 0.189894
R23695 minus.n36 minus.n35 0.189894
R23696 minus.n37 minus.n36 0.189894
R23697 minus.n37 minus.n0 0.189894
R23698 minus.n41 minus.n0 0.189894
R23699 output.n41 output.n15 289.615
R23700 output.n72 output.n46 289.615
R23701 output.n104 output.n78 289.615
R23702 output.n136 output.n110 289.615
R23703 output.n77 output.n45 197.26
R23704 output.n77 output.n76 196.298
R23705 output.n109 output.n108 196.298
R23706 output.n141 output.n140 196.298
R23707 output.n42 output.n41 185
R23708 output.n40 output.n39 185
R23709 output.n19 output.n18 185
R23710 output.n34 output.n33 185
R23711 output.n32 output.n31 185
R23712 output.n23 output.n22 185
R23713 output.n26 output.n25 185
R23714 output.n73 output.n72 185
R23715 output.n71 output.n70 185
R23716 output.n50 output.n49 185
R23717 output.n65 output.n64 185
R23718 output.n63 output.n62 185
R23719 output.n54 output.n53 185
R23720 output.n57 output.n56 185
R23721 output.n105 output.n104 185
R23722 output.n103 output.n102 185
R23723 output.n82 output.n81 185
R23724 output.n97 output.n96 185
R23725 output.n95 output.n94 185
R23726 output.n86 output.n85 185
R23727 output.n89 output.n88 185
R23728 output.n137 output.n136 185
R23729 output.n135 output.n134 185
R23730 output.n114 output.n113 185
R23731 output.n129 output.n128 185
R23732 output.n127 output.n126 185
R23733 output.n118 output.n117 185
R23734 output.n121 output.n120 185
R23735 output.t1 output.n24 147.661
R23736 output.t0 output.n55 147.661
R23737 output.t2 output.n87 147.661
R23738 output.t3 output.n119 147.661
R23739 output.n41 output.n40 104.615
R23740 output.n40 output.n18 104.615
R23741 output.n33 output.n18 104.615
R23742 output.n33 output.n32 104.615
R23743 output.n32 output.n22 104.615
R23744 output.n25 output.n22 104.615
R23745 output.n72 output.n71 104.615
R23746 output.n71 output.n49 104.615
R23747 output.n64 output.n49 104.615
R23748 output.n64 output.n63 104.615
R23749 output.n63 output.n53 104.615
R23750 output.n56 output.n53 104.615
R23751 output.n104 output.n103 104.615
R23752 output.n103 output.n81 104.615
R23753 output.n96 output.n81 104.615
R23754 output.n96 output.n95 104.615
R23755 output.n95 output.n85 104.615
R23756 output.n88 output.n85 104.615
R23757 output.n136 output.n135 104.615
R23758 output.n135 output.n113 104.615
R23759 output.n128 output.n113 104.615
R23760 output.n128 output.n127 104.615
R23761 output.n127 output.n117 104.615
R23762 output.n120 output.n117 104.615
R23763 output.n1 output.t5 77.056
R23764 output.n14 output.t7 76.6694
R23765 output.n1 output.n0 72.7095
R23766 output.n3 output.n2 72.7095
R23767 output.n5 output.n4 72.7095
R23768 output.n7 output.n6 72.7095
R23769 output.n9 output.n8 72.7095
R23770 output.n11 output.n10 72.7095
R23771 output.n13 output.n12 72.7095
R23772 output.n25 output.t1 52.3082
R23773 output.n56 output.t0 52.3082
R23774 output.n88 output.t2 52.3082
R23775 output.n120 output.t3 52.3082
R23776 output.n26 output.n24 15.6674
R23777 output.n57 output.n55 15.6674
R23778 output.n89 output.n87 15.6674
R23779 output.n121 output.n119 15.6674
R23780 output.n27 output.n23 12.8005
R23781 output.n58 output.n54 12.8005
R23782 output.n90 output.n86 12.8005
R23783 output.n122 output.n118 12.8005
R23784 output.n31 output.n30 12.0247
R23785 output.n62 output.n61 12.0247
R23786 output.n94 output.n93 12.0247
R23787 output.n126 output.n125 12.0247
R23788 output.n34 output.n21 11.249
R23789 output.n65 output.n52 11.249
R23790 output.n97 output.n84 11.249
R23791 output.n129 output.n116 11.249
R23792 output.n35 output.n19 10.4732
R23793 output.n66 output.n50 10.4732
R23794 output.n98 output.n82 10.4732
R23795 output.n130 output.n114 10.4732
R23796 output.n39 output.n38 9.69747
R23797 output.n70 output.n69 9.69747
R23798 output.n102 output.n101 9.69747
R23799 output.n134 output.n133 9.69747
R23800 output.n45 output.n44 9.45567
R23801 output.n76 output.n75 9.45567
R23802 output.n108 output.n107 9.45567
R23803 output.n140 output.n139 9.45567
R23804 output.n44 output.n43 9.3005
R23805 output.n17 output.n16 9.3005
R23806 output.n38 output.n37 9.3005
R23807 output.n36 output.n35 9.3005
R23808 output.n21 output.n20 9.3005
R23809 output.n30 output.n29 9.3005
R23810 output.n28 output.n27 9.3005
R23811 output.n75 output.n74 9.3005
R23812 output.n48 output.n47 9.3005
R23813 output.n69 output.n68 9.3005
R23814 output.n67 output.n66 9.3005
R23815 output.n52 output.n51 9.3005
R23816 output.n61 output.n60 9.3005
R23817 output.n59 output.n58 9.3005
R23818 output.n107 output.n106 9.3005
R23819 output.n80 output.n79 9.3005
R23820 output.n101 output.n100 9.3005
R23821 output.n99 output.n98 9.3005
R23822 output.n84 output.n83 9.3005
R23823 output.n93 output.n92 9.3005
R23824 output.n91 output.n90 9.3005
R23825 output.n139 output.n138 9.3005
R23826 output.n112 output.n111 9.3005
R23827 output.n133 output.n132 9.3005
R23828 output.n131 output.n130 9.3005
R23829 output.n116 output.n115 9.3005
R23830 output.n125 output.n124 9.3005
R23831 output.n123 output.n122 9.3005
R23832 output.n42 output.n17 8.92171
R23833 output.n73 output.n48 8.92171
R23834 output.n105 output.n80 8.92171
R23835 output.n137 output.n112 8.92171
R23836 output output.n141 8.15037
R23837 output.n43 output.n15 8.14595
R23838 output.n74 output.n46 8.14595
R23839 output.n106 output.n78 8.14595
R23840 output.n138 output.n110 8.14595
R23841 output.n45 output.n15 5.81868
R23842 output.n76 output.n46 5.81868
R23843 output.n108 output.n78 5.81868
R23844 output.n140 output.n110 5.81868
R23845 output.n43 output.n42 5.04292
R23846 output.n74 output.n73 5.04292
R23847 output.n106 output.n105 5.04292
R23848 output.n138 output.n137 5.04292
R23849 output.n28 output.n24 4.38594
R23850 output.n59 output.n55 4.38594
R23851 output.n91 output.n87 4.38594
R23852 output.n123 output.n119 4.38594
R23853 output.n39 output.n17 4.26717
R23854 output.n70 output.n48 4.26717
R23855 output.n102 output.n80 4.26717
R23856 output.n134 output.n112 4.26717
R23857 output.n0 output.t11 3.9605
R23858 output.n0 output.t16 3.9605
R23859 output.n2 output.t4 3.9605
R23860 output.n2 output.t12 3.9605
R23861 output.n4 output.t14 3.9605
R23862 output.n4 output.t13 3.9605
R23863 output.n6 output.t19 3.9605
R23864 output.n6 output.t6 3.9605
R23865 output.n8 output.t8 3.9605
R23866 output.n8 output.t17 3.9605
R23867 output.n10 output.t18 3.9605
R23868 output.n10 output.t9 3.9605
R23869 output.n12 output.t10 3.9605
R23870 output.n12 output.t15 3.9605
R23871 output.n38 output.n19 3.49141
R23872 output.n69 output.n50 3.49141
R23873 output.n101 output.n82 3.49141
R23874 output.n133 output.n114 3.49141
R23875 output.n35 output.n34 2.71565
R23876 output.n66 output.n65 2.71565
R23877 output.n98 output.n97 2.71565
R23878 output.n130 output.n129 2.71565
R23879 output.n31 output.n21 1.93989
R23880 output.n62 output.n52 1.93989
R23881 output.n94 output.n84 1.93989
R23882 output.n126 output.n116 1.93989
R23883 output.n30 output.n23 1.16414
R23884 output.n61 output.n54 1.16414
R23885 output.n93 output.n86 1.16414
R23886 output.n125 output.n118 1.16414
R23887 output.n141 output.n109 0.962709
R23888 output.n109 output.n77 0.962709
R23889 output.n27 output.n26 0.388379
R23890 output.n58 output.n57 0.388379
R23891 output.n90 output.n89 0.388379
R23892 output.n122 output.n121 0.388379
R23893 output.n14 output.n13 0.387128
R23894 output.n13 output.n11 0.387128
R23895 output.n11 output.n9 0.387128
R23896 output.n9 output.n7 0.387128
R23897 output.n7 output.n5 0.387128
R23898 output.n5 output.n3 0.387128
R23899 output.n3 output.n1 0.387128
R23900 output.n44 output.n16 0.155672
R23901 output.n37 output.n16 0.155672
R23902 output.n37 output.n36 0.155672
R23903 output.n36 output.n20 0.155672
R23904 output.n29 output.n20 0.155672
R23905 output.n29 output.n28 0.155672
R23906 output.n75 output.n47 0.155672
R23907 output.n68 output.n47 0.155672
R23908 output.n68 output.n67 0.155672
R23909 output.n67 output.n51 0.155672
R23910 output.n60 output.n51 0.155672
R23911 output.n60 output.n59 0.155672
R23912 output.n107 output.n79 0.155672
R23913 output.n100 output.n79 0.155672
R23914 output.n100 output.n99 0.155672
R23915 output.n99 output.n83 0.155672
R23916 output.n92 output.n83 0.155672
R23917 output.n92 output.n91 0.155672
R23918 output.n139 output.n111 0.155672
R23919 output.n132 output.n111 0.155672
R23920 output.n132 output.n131 0.155672
R23921 output.n131 output.n115 0.155672
R23922 output.n124 output.n115 0.155672
R23923 output.n124 output.n123 0.155672
R23924 output output.n14 0.126227
R23925 diffpairibias.n0 diffpairibias.t18 436.822
R23926 diffpairibias.n21 diffpairibias.t19 435.479
R23927 diffpairibias.n20 diffpairibias.t16 435.479
R23928 diffpairibias.n19 diffpairibias.t17 435.479
R23929 diffpairibias.n18 diffpairibias.t21 435.479
R23930 diffpairibias.n0 diffpairibias.t22 435.479
R23931 diffpairibias.n1 diffpairibias.t20 435.479
R23932 diffpairibias.n2 diffpairibias.t23 435.479
R23933 diffpairibias.n10 diffpairibias.t0 377.536
R23934 diffpairibias.n10 diffpairibias.t8 376.193
R23935 diffpairibias.n11 diffpairibias.t10 376.193
R23936 diffpairibias.n12 diffpairibias.t6 376.193
R23937 diffpairibias.n13 diffpairibias.t2 376.193
R23938 diffpairibias.n14 diffpairibias.t12 376.193
R23939 diffpairibias.n15 diffpairibias.t4 376.193
R23940 diffpairibias.n16 diffpairibias.t14 376.193
R23941 diffpairibias.n3 diffpairibias.t1 113.368
R23942 diffpairibias.n3 diffpairibias.t9 112.698
R23943 diffpairibias.n4 diffpairibias.t11 112.698
R23944 diffpairibias.n5 diffpairibias.t7 112.698
R23945 diffpairibias.n6 diffpairibias.t3 112.698
R23946 diffpairibias.n7 diffpairibias.t13 112.698
R23947 diffpairibias.n8 diffpairibias.t5 112.698
R23948 diffpairibias.n9 diffpairibias.t15 112.698
R23949 diffpairibias.n17 diffpairibias.n16 4.77242
R23950 diffpairibias.n17 diffpairibias.n9 4.30807
R23951 diffpairibias.n18 diffpairibias.n17 4.13945
R23952 diffpairibias.n16 diffpairibias.n15 1.34352
R23953 diffpairibias.n15 diffpairibias.n14 1.34352
R23954 diffpairibias.n14 diffpairibias.n13 1.34352
R23955 diffpairibias.n13 diffpairibias.n12 1.34352
R23956 diffpairibias.n12 diffpairibias.n11 1.34352
R23957 diffpairibias.n11 diffpairibias.n10 1.34352
R23958 diffpairibias.n2 diffpairibias.n1 1.34352
R23959 diffpairibias.n1 diffpairibias.n0 1.34352
R23960 diffpairibias.n19 diffpairibias.n18 1.34352
R23961 diffpairibias.n20 diffpairibias.n19 1.34352
R23962 diffpairibias.n21 diffpairibias.n20 1.34352
R23963 diffpairibias.n22 diffpairibias.n21 0.862419
R23964 diffpairibias diffpairibias.n22 0.684875
R23965 diffpairibias.n9 diffpairibias.n8 0.672012
R23966 diffpairibias.n8 diffpairibias.n7 0.672012
R23967 diffpairibias.n7 diffpairibias.n6 0.672012
R23968 diffpairibias.n6 diffpairibias.n5 0.672012
R23969 diffpairibias.n5 diffpairibias.n4 0.672012
R23970 diffpairibias.n4 diffpairibias.n3 0.672012
R23971 diffpairibias.n22 diffpairibias.n2 0.190907
R23972 outputibias.n27 outputibias.n1 289.615
R23973 outputibias.n58 outputibias.n32 289.615
R23974 outputibias.n90 outputibias.n64 289.615
R23975 outputibias.n122 outputibias.n96 289.615
R23976 outputibias.n28 outputibias.n27 185
R23977 outputibias.n26 outputibias.n25 185
R23978 outputibias.n5 outputibias.n4 185
R23979 outputibias.n20 outputibias.n19 185
R23980 outputibias.n18 outputibias.n17 185
R23981 outputibias.n9 outputibias.n8 185
R23982 outputibias.n12 outputibias.n11 185
R23983 outputibias.n59 outputibias.n58 185
R23984 outputibias.n57 outputibias.n56 185
R23985 outputibias.n36 outputibias.n35 185
R23986 outputibias.n51 outputibias.n50 185
R23987 outputibias.n49 outputibias.n48 185
R23988 outputibias.n40 outputibias.n39 185
R23989 outputibias.n43 outputibias.n42 185
R23990 outputibias.n91 outputibias.n90 185
R23991 outputibias.n89 outputibias.n88 185
R23992 outputibias.n68 outputibias.n67 185
R23993 outputibias.n83 outputibias.n82 185
R23994 outputibias.n81 outputibias.n80 185
R23995 outputibias.n72 outputibias.n71 185
R23996 outputibias.n75 outputibias.n74 185
R23997 outputibias.n123 outputibias.n122 185
R23998 outputibias.n121 outputibias.n120 185
R23999 outputibias.n100 outputibias.n99 185
R24000 outputibias.n115 outputibias.n114 185
R24001 outputibias.n113 outputibias.n112 185
R24002 outputibias.n104 outputibias.n103 185
R24003 outputibias.n107 outputibias.n106 185
R24004 outputibias.n0 outputibias.t10 178.945
R24005 outputibias.n133 outputibias.t8 177.018
R24006 outputibias.n132 outputibias.t11 177.018
R24007 outputibias.n0 outputibias.t9 177.018
R24008 outputibias.t7 outputibias.n10 147.661
R24009 outputibias.t1 outputibias.n41 147.661
R24010 outputibias.t3 outputibias.n73 147.661
R24011 outputibias.t5 outputibias.n105 147.661
R24012 outputibias.n128 outputibias.t6 132.363
R24013 outputibias.n128 outputibias.t0 130.436
R24014 outputibias.n129 outputibias.t2 130.436
R24015 outputibias.n130 outputibias.t4 130.436
R24016 outputibias.n27 outputibias.n26 104.615
R24017 outputibias.n26 outputibias.n4 104.615
R24018 outputibias.n19 outputibias.n4 104.615
R24019 outputibias.n19 outputibias.n18 104.615
R24020 outputibias.n18 outputibias.n8 104.615
R24021 outputibias.n11 outputibias.n8 104.615
R24022 outputibias.n58 outputibias.n57 104.615
R24023 outputibias.n57 outputibias.n35 104.615
R24024 outputibias.n50 outputibias.n35 104.615
R24025 outputibias.n50 outputibias.n49 104.615
R24026 outputibias.n49 outputibias.n39 104.615
R24027 outputibias.n42 outputibias.n39 104.615
R24028 outputibias.n90 outputibias.n89 104.615
R24029 outputibias.n89 outputibias.n67 104.615
R24030 outputibias.n82 outputibias.n67 104.615
R24031 outputibias.n82 outputibias.n81 104.615
R24032 outputibias.n81 outputibias.n71 104.615
R24033 outputibias.n74 outputibias.n71 104.615
R24034 outputibias.n122 outputibias.n121 104.615
R24035 outputibias.n121 outputibias.n99 104.615
R24036 outputibias.n114 outputibias.n99 104.615
R24037 outputibias.n114 outputibias.n113 104.615
R24038 outputibias.n113 outputibias.n103 104.615
R24039 outputibias.n106 outputibias.n103 104.615
R24040 outputibias.n63 outputibias.n31 95.6354
R24041 outputibias.n63 outputibias.n62 94.6732
R24042 outputibias.n95 outputibias.n94 94.6732
R24043 outputibias.n127 outputibias.n126 94.6732
R24044 outputibias.n11 outputibias.t7 52.3082
R24045 outputibias.n42 outputibias.t1 52.3082
R24046 outputibias.n74 outputibias.t3 52.3082
R24047 outputibias.n106 outputibias.t5 52.3082
R24048 outputibias.n12 outputibias.n10 15.6674
R24049 outputibias.n43 outputibias.n41 15.6674
R24050 outputibias.n75 outputibias.n73 15.6674
R24051 outputibias.n107 outputibias.n105 15.6674
R24052 outputibias.n13 outputibias.n9 12.8005
R24053 outputibias.n44 outputibias.n40 12.8005
R24054 outputibias.n76 outputibias.n72 12.8005
R24055 outputibias.n108 outputibias.n104 12.8005
R24056 outputibias.n17 outputibias.n16 12.0247
R24057 outputibias.n48 outputibias.n47 12.0247
R24058 outputibias.n80 outputibias.n79 12.0247
R24059 outputibias.n112 outputibias.n111 12.0247
R24060 outputibias.n20 outputibias.n7 11.249
R24061 outputibias.n51 outputibias.n38 11.249
R24062 outputibias.n83 outputibias.n70 11.249
R24063 outputibias.n115 outputibias.n102 11.249
R24064 outputibias.n21 outputibias.n5 10.4732
R24065 outputibias.n52 outputibias.n36 10.4732
R24066 outputibias.n84 outputibias.n68 10.4732
R24067 outputibias.n116 outputibias.n100 10.4732
R24068 outputibias.n25 outputibias.n24 9.69747
R24069 outputibias.n56 outputibias.n55 9.69747
R24070 outputibias.n88 outputibias.n87 9.69747
R24071 outputibias.n120 outputibias.n119 9.69747
R24072 outputibias.n31 outputibias.n30 9.45567
R24073 outputibias.n62 outputibias.n61 9.45567
R24074 outputibias.n94 outputibias.n93 9.45567
R24075 outputibias.n126 outputibias.n125 9.45567
R24076 outputibias.n30 outputibias.n29 9.3005
R24077 outputibias.n3 outputibias.n2 9.3005
R24078 outputibias.n24 outputibias.n23 9.3005
R24079 outputibias.n22 outputibias.n21 9.3005
R24080 outputibias.n7 outputibias.n6 9.3005
R24081 outputibias.n16 outputibias.n15 9.3005
R24082 outputibias.n14 outputibias.n13 9.3005
R24083 outputibias.n61 outputibias.n60 9.3005
R24084 outputibias.n34 outputibias.n33 9.3005
R24085 outputibias.n55 outputibias.n54 9.3005
R24086 outputibias.n53 outputibias.n52 9.3005
R24087 outputibias.n38 outputibias.n37 9.3005
R24088 outputibias.n47 outputibias.n46 9.3005
R24089 outputibias.n45 outputibias.n44 9.3005
R24090 outputibias.n93 outputibias.n92 9.3005
R24091 outputibias.n66 outputibias.n65 9.3005
R24092 outputibias.n87 outputibias.n86 9.3005
R24093 outputibias.n85 outputibias.n84 9.3005
R24094 outputibias.n70 outputibias.n69 9.3005
R24095 outputibias.n79 outputibias.n78 9.3005
R24096 outputibias.n77 outputibias.n76 9.3005
R24097 outputibias.n125 outputibias.n124 9.3005
R24098 outputibias.n98 outputibias.n97 9.3005
R24099 outputibias.n119 outputibias.n118 9.3005
R24100 outputibias.n117 outputibias.n116 9.3005
R24101 outputibias.n102 outputibias.n101 9.3005
R24102 outputibias.n111 outputibias.n110 9.3005
R24103 outputibias.n109 outputibias.n108 9.3005
R24104 outputibias.n28 outputibias.n3 8.92171
R24105 outputibias.n59 outputibias.n34 8.92171
R24106 outputibias.n91 outputibias.n66 8.92171
R24107 outputibias.n123 outputibias.n98 8.92171
R24108 outputibias.n29 outputibias.n1 8.14595
R24109 outputibias.n60 outputibias.n32 8.14595
R24110 outputibias.n92 outputibias.n64 8.14595
R24111 outputibias.n124 outputibias.n96 8.14595
R24112 outputibias.n31 outputibias.n1 5.81868
R24113 outputibias.n62 outputibias.n32 5.81868
R24114 outputibias.n94 outputibias.n64 5.81868
R24115 outputibias.n126 outputibias.n96 5.81868
R24116 outputibias.n131 outputibias.n130 5.20947
R24117 outputibias.n29 outputibias.n28 5.04292
R24118 outputibias.n60 outputibias.n59 5.04292
R24119 outputibias.n92 outputibias.n91 5.04292
R24120 outputibias.n124 outputibias.n123 5.04292
R24121 outputibias.n131 outputibias.n127 4.42209
R24122 outputibias.n14 outputibias.n10 4.38594
R24123 outputibias.n45 outputibias.n41 4.38594
R24124 outputibias.n77 outputibias.n73 4.38594
R24125 outputibias.n109 outputibias.n105 4.38594
R24126 outputibias.n132 outputibias.n131 4.28454
R24127 outputibias.n25 outputibias.n3 4.26717
R24128 outputibias.n56 outputibias.n34 4.26717
R24129 outputibias.n88 outputibias.n66 4.26717
R24130 outputibias.n120 outputibias.n98 4.26717
R24131 outputibias.n24 outputibias.n5 3.49141
R24132 outputibias.n55 outputibias.n36 3.49141
R24133 outputibias.n87 outputibias.n68 3.49141
R24134 outputibias.n119 outputibias.n100 3.49141
R24135 outputibias.n21 outputibias.n20 2.71565
R24136 outputibias.n52 outputibias.n51 2.71565
R24137 outputibias.n84 outputibias.n83 2.71565
R24138 outputibias.n116 outputibias.n115 2.71565
R24139 outputibias.n17 outputibias.n7 1.93989
R24140 outputibias.n48 outputibias.n38 1.93989
R24141 outputibias.n80 outputibias.n70 1.93989
R24142 outputibias.n112 outputibias.n102 1.93989
R24143 outputibias.n130 outputibias.n129 1.9266
R24144 outputibias.n129 outputibias.n128 1.9266
R24145 outputibias.n133 outputibias.n132 1.92658
R24146 outputibias.n134 outputibias.n133 1.29913
R24147 outputibias.n16 outputibias.n9 1.16414
R24148 outputibias.n47 outputibias.n40 1.16414
R24149 outputibias.n79 outputibias.n72 1.16414
R24150 outputibias.n111 outputibias.n104 1.16414
R24151 outputibias.n127 outputibias.n95 0.962709
R24152 outputibias.n95 outputibias.n63 0.962709
R24153 outputibias.n13 outputibias.n12 0.388379
R24154 outputibias.n44 outputibias.n43 0.388379
R24155 outputibias.n76 outputibias.n75 0.388379
R24156 outputibias.n108 outputibias.n107 0.388379
R24157 outputibias.n134 outputibias.n0 0.337251
R24158 outputibias outputibias.n134 0.302375
R24159 outputibias.n30 outputibias.n2 0.155672
R24160 outputibias.n23 outputibias.n2 0.155672
R24161 outputibias.n23 outputibias.n22 0.155672
R24162 outputibias.n22 outputibias.n6 0.155672
R24163 outputibias.n15 outputibias.n6 0.155672
R24164 outputibias.n15 outputibias.n14 0.155672
R24165 outputibias.n61 outputibias.n33 0.155672
R24166 outputibias.n54 outputibias.n33 0.155672
R24167 outputibias.n54 outputibias.n53 0.155672
R24168 outputibias.n53 outputibias.n37 0.155672
R24169 outputibias.n46 outputibias.n37 0.155672
R24170 outputibias.n46 outputibias.n45 0.155672
R24171 outputibias.n93 outputibias.n65 0.155672
R24172 outputibias.n86 outputibias.n65 0.155672
R24173 outputibias.n86 outputibias.n85 0.155672
R24174 outputibias.n85 outputibias.n69 0.155672
R24175 outputibias.n78 outputibias.n69 0.155672
R24176 outputibias.n78 outputibias.n77 0.155672
R24177 outputibias.n125 outputibias.n97 0.155672
R24178 outputibias.n118 outputibias.n97 0.155672
R24179 outputibias.n118 outputibias.n117 0.155672
R24180 outputibias.n117 outputibias.n101 0.155672
R24181 outputibias.n110 outputibias.n101 0.155672
R24182 outputibias.n110 outputibias.n109 0.155672
C0 minus diffpairibias 4.33e-19
C1 commonsourceibias output 0.006808f
C2 CSoutput minus 2.6584f
C3 vdd plus 0.0878f
C4 commonsourceibias outputibias 0.003832f
C5 plus diffpairibias 4.56e-19
C6 vdd commonsourceibias 0.004218f
C7 CSoutput plus 0.874787f
C8 commonsourceibias diffpairibias 0.06482f
C9 CSoutput commonsourceibias 54.0646f
C10 minus plus 9.59292f
C11 minus commonsourceibias 0.460231f
C12 plus commonsourceibias 0.415048f
C13 output outputibias 2.34152f
C14 vdd output 7.23429f
C15 CSoutput output 6.13881f
C16 CSoutput outputibias 0.032386f
C17 vdd CSoutput 92.9043f
C18 diffpairibias gnd 48.980137f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.183172p
C22 plus gnd 35.947304f
C23 minus gnd 28.75732f
C24 CSoutput gnd 0.124778p
C25 vdd gnd 0.479896p
C26 outputibias.t9 gnd 0.11477f
C27 outputibias.t10 gnd 0.115567f
C28 outputibias.n0 gnd 0.130108f
C29 outputibias.n1 gnd 0.001372f
C30 outputibias.n2 gnd 9.76e-19
C31 outputibias.n3 gnd 5.24e-19
C32 outputibias.n4 gnd 0.001239f
C33 outputibias.n5 gnd 5.55e-19
C34 outputibias.n6 gnd 9.76e-19
C35 outputibias.n7 gnd 5.24e-19
C36 outputibias.n8 gnd 0.001239f
C37 outputibias.n9 gnd 5.55e-19
C38 outputibias.n10 gnd 0.004176f
C39 outputibias.t7 gnd 0.00202f
C40 outputibias.n11 gnd 9.3e-19
C41 outputibias.n12 gnd 7.32e-19
C42 outputibias.n13 gnd 5.24e-19
C43 outputibias.n14 gnd 0.02322f
C44 outputibias.n15 gnd 9.76e-19
C45 outputibias.n16 gnd 5.24e-19
C46 outputibias.n17 gnd 5.55e-19
C47 outputibias.n18 gnd 0.001239f
C48 outputibias.n19 gnd 0.001239f
C49 outputibias.n20 gnd 5.55e-19
C50 outputibias.n21 gnd 5.24e-19
C51 outputibias.n22 gnd 9.76e-19
C52 outputibias.n23 gnd 9.76e-19
C53 outputibias.n24 gnd 5.24e-19
C54 outputibias.n25 gnd 5.55e-19
C55 outputibias.n26 gnd 0.001239f
C56 outputibias.n27 gnd 0.002683f
C57 outputibias.n28 gnd 5.55e-19
C58 outputibias.n29 gnd 5.24e-19
C59 outputibias.n30 gnd 0.002256f
C60 outputibias.n31 gnd 0.005781f
C61 outputibias.n32 gnd 0.001372f
C62 outputibias.n33 gnd 9.76e-19
C63 outputibias.n34 gnd 5.24e-19
C64 outputibias.n35 gnd 0.001239f
C65 outputibias.n36 gnd 5.55e-19
C66 outputibias.n37 gnd 9.76e-19
C67 outputibias.n38 gnd 5.24e-19
C68 outputibias.n39 gnd 0.001239f
C69 outputibias.n40 gnd 5.55e-19
C70 outputibias.n41 gnd 0.004176f
C71 outputibias.t1 gnd 0.00202f
C72 outputibias.n42 gnd 9.3e-19
C73 outputibias.n43 gnd 7.32e-19
C74 outputibias.n44 gnd 5.24e-19
C75 outputibias.n45 gnd 0.02322f
C76 outputibias.n46 gnd 9.76e-19
C77 outputibias.n47 gnd 5.24e-19
C78 outputibias.n48 gnd 5.55e-19
C79 outputibias.n49 gnd 0.001239f
C80 outputibias.n50 gnd 0.001239f
C81 outputibias.n51 gnd 5.55e-19
C82 outputibias.n52 gnd 5.24e-19
C83 outputibias.n53 gnd 9.76e-19
C84 outputibias.n54 gnd 9.76e-19
C85 outputibias.n55 gnd 5.24e-19
C86 outputibias.n56 gnd 5.55e-19
C87 outputibias.n57 gnd 0.001239f
C88 outputibias.n58 gnd 0.002683f
C89 outputibias.n59 gnd 5.55e-19
C90 outputibias.n60 gnd 5.24e-19
C91 outputibias.n61 gnd 0.002256f
C92 outputibias.n62 gnd 0.005197f
C93 outputibias.n63 gnd 0.121892f
C94 outputibias.n64 gnd 0.001372f
C95 outputibias.n65 gnd 9.76e-19
C96 outputibias.n66 gnd 5.24e-19
C97 outputibias.n67 gnd 0.001239f
C98 outputibias.n68 gnd 5.55e-19
C99 outputibias.n69 gnd 9.76e-19
C100 outputibias.n70 gnd 5.24e-19
C101 outputibias.n71 gnd 0.001239f
C102 outputibias.n72 gnd 5.55e-19
C103 outputibias.n73 gnd 0.004176f
C104 outputibias.t3 gnd 0.00202f
C105 outputibias.n74 gnd 9.3e-19
C106 outputibias.n75 gnd 7.32e-19
C107 outputibias.n76 gnd 5.24e-19
C108 outputibias.n77 gnd 0.02322f
C109 outputibias.n78 gnd 9.76e-19
C110 outputibias.n79 gnd 5.24e-19
C111 outputibias.n80 gnd 5.55e-19
C112 outputibias.n81 gnd 0.001239f
C113 outputibias.n82 gnd 0.001239f
C114 outputibias.n83 gnd 5.55e-19
C115 outputibias.n84 gnd 5.24e-19
C116 outputibias.n85 gnd 9.76e-19
C117 outputibias.n86 gnd 9.76e-19
C118 outputibias.n87 gnd 5.24e-19
C119 outputibias.n88 gnd 5.55e-19
C120 outputibias.n89 gnd 0.001239f
C121 outputibias.n90 gnd 0.002683f
C122 outputibias.n91 gnd 5.55e-19
C123 outputibias.n92 gnd 5.24e-19
C124 outputibias.n93 gnd 0.002256f
C125 outputibias.n94 gnd 0.005197f
C126 outputibias.n95 gnd 0.064513f
C127 outputibias.n96 gnd 0.001372f
C128 outputibias.n97 gnd 9.76e-19
C129 outputibias.n98 gnd 5.24e-19
C130 outputibias.n99 gnd 0.001239f
C131 outputibias.n100 gnd 5.55e-19
C132 outputibias.n101 gnd 9.76e-19
C133 outputibias.n102 gnd 5.24e-19
C134 outputibias.n103 gnd 0.001239f
C135 outputibias.n104 gnd 5.55e-19
C136 outputibias.n105 gnd 0.004176f
C137 outputibias.t5 gnd 0.00202f
C138 outputibias.n106 gnd 9.3e-19
C139 outputibias.n107 gnd 7.32e-19
C140 outputibias.n108 gnd 5.24e-19
C141 outputibias.n109 gnd 0.02322f
C142 outputibias.n110 gnd 9.76e-19
C143 outputibias.n111 gnd 5.24e-19
C144 outputibias.n112 gnd 5.55e-19
C145 outputibias.n113 gnd 0.001239f
C146 outputibias.n114 gnd 0.001239f
C147 outputibias.n115 gnd 5.55e-19
C148 outputibias.n116 gnd 5.24e-19
C149 outputibias.n117 gnd 9.76e-19
C150 outputibias.n118 gnd 9.76e-19
C151 outputibias.n119 gnd 5.24e-19
C152 outputibias.n120 gnd 5.55e-19
C153 outputibias.n121 gnd 0.001239f
C154 outputibias.n122 gnd 0.002683f
C155 outputibias.n123 gnd 5.55e-19
C156 outputibias.n124 gnd 5.24e-19
C157 outputibias.n125 gnd 0.002256f
C158 outputibias.n126 gnd 0.005197f
C159 outputibias.n127 gnd 0.084814f
C160 outputibias.t4 gnd 0.108319f
C161 outputibias.t2 gnd 0.108319f
C162 outputibias.t0 gnd 0.108319f
C163 outputibias.t6 gnd 0.109238f
C164 outputibias.n128 gnd 0.134674f
C165 outputibias.n129 gnd 0.07244f
C166 outputibias.n130 gnd 0.079818f
C167 outputibias.n131 gnd 0.164901f
C168 outputibias.t11 gnd 0.11477f
C169 outputibias.n132 gnd 0.067481f
C170 outputibias.t8 gnd 0.11477f
C171 outputibias.n133 gnd 0.065115f
C172 outputibias.n134 gnd 0.029159f
C173 diffpairibias.t18 gnd 0.087401f
C174 diffpairibias.t22 gnd 0.087239f
C175 diffpairibias.n0 gnd 0.102784f
C176 diffpairibias.t20 gnd 0.087239f
C177 diffpairibias.n1 gnd 0.050171f
C178 diffpairibias.t23 gnd 0.087239f
C179 diffpairibias.n2 gnd 0.039841f
C180 diffpairibias.t1 gnd 0.083757f
C181 diffpairibias.t9 gnd 0.083392f
C182 diffpairibias.n3 gnd 0.131682f
C183 diffpairibias.t11 gnd 0.083392f
C184 diffpairibias.n4 gnd 0.07027f
C185 diffpairibias.t7 gnd 0.083392f
C186 diffpairibias.n5 gnd 0.07027f
C187 diffpairibias.t3 gnd 0.083392f
C188 diffpairibias.n6 gnd 0.07027f
C189 diffpairibias.t13 gnd 0.083392f
C190 diffpairibias.n7 gnd 0.07027f
C191 diffpairibias.t5 gnd 0.083392f
C192 diffpairibias.n8 gnd 0.07027f
C193 diffpairibias.t15 gnd 0.083392f
C194 diffpairibias.n9 gnd 0.099771f
C195 diffpairibias.t0 gnd 0.08427f
C196 diffpairibias.t8 gnd 0.084123f
C197 diffpairibias.n10 gnd 0.091784f
C198 diffpairibias.t10 gnd 0.084123f
C199 diffpairibias.n11 gnd 0.050681f
C200 diffpairibias.t6 gnd 0.084123f
C201 diffpairibias.n12 gnd 0.050681f
C202 diffpairibias.t2 gnd 0.084123f
C203 diffpairibias.n13 gnd 0.050681f
C204 diffpairibias.t12 gnd 0.084123f
C205 diffpairibias.n14 gnd 0.050681f
C206 diffpairibias.t4 gnd 0.084123f
C207 diffpairibias.n15 gnd 0.050681f
C208 diffpairibias.t14 gnd 0.084123f
C209 diffpairibias.n16 gnd 0.059977f
C210 diffpairibias.n17 gnd 0.226448f
C211 diffpairibias.t21 gnd 0.087239f
C212 diffpairibias.n18 gnd 0.050181f
C213 diffpairibias.t17 gnd 0.087239f
C214 diffpairibias.n19 gnd 0.050171f
C215 diffpairibias.t16 gnd 0.087239f
C216 diffpairibias.n20 gnd 0.050171f
C217 diffpairibias.t19 gnd 0.087239f
C218 diffpairibias.n21 gnd 0.045859f
C219 diffpairibias.n22 gnd 0.046268f
C220 output.t5 gnd 0.464308f
C221 output.t11 gnd 0.044422f
C222 output.t16 gnd 0.044422f
C223 output.n0 gnd 0.364624f
C224 output.n1 gnd 0.614102f
C225 output.t4 gnd 0.044422f
C226 output.t12 gnd 0.044422f
C227 output.n2 gnd 0.364624f
C228 output.n3 gnd 0.350265f
C229 output.t14 gnd 0.044422f
C230 output.t13 gnd 0.044422f
C231 output.n4 gnd 0.364624f
C232 output.n5 gnd 0.350265f
C233 output.t19 gnd 0.044422f
C234 output.t6 gnd 0.044422f
C235 output.n6 gnd 0.364624f
C236 output.n7 gnd 0.350265f
C237 output.t8 gnd 0.044422f
C238 output.t17 gnd 0.044422f
C239 output.n8 gnd 0.364624f
C240 output.n9 gnd 0.350265f
C241 output.t18 gnd 0.044422f
C242 output.t9 gnd 0.044422f
C243 output.n10 gnd 0.364624f
C244 output.n11 gnd 0.350265f
C245 output.t10 gnd 0.044422f
C246 output.t15 gnd 0.044422f
C247 output.n12 gnd 0.364624f
C248 output.n13 gnd 0.350265f
C249 output.t7 gnd 0.462979f
C250 output.n14 gnd 0.28994f
C251 output.n15 gnd 0.015803f
C252 output.n16 gnd 0.011243f
C253 output.n17 gnd 0.006041f
C254 output.n18 gnd 0.01428f
C255 output.n19 gnd 0.006397f
C256 output.n20 gnd 0.011243f
C257 output.n21 gnd 0.006041f
C258 output.n22 gnd 0.01428f
C259 output.n23 gnd 0.006397f
C260 output.n24 gnd 0.048111f
C261 output.t1 gnd 0.023274f
C262 output.n25 gnd 0.01071f
C263 output.n26 gnd 0.008435f
C264 output.n27 gnd 0.006041f
C265 output.n28 gnd 0.267512f
C266 output.n29 gnd 0.011243f
C267 output.n30 gnd 0.006041f
C268 output.n31 gnd 0.006397f
C269 output.n32 gnd 0.01428f
C270 output.n33 gnd 0.01428f
C271 output.n34 gnd 0.006397f
C272 output.n35 gnd 0.006041f
C273 output.n36 gnd 0.011243f
C274 output.n37 gnd 0.011243f
C275 output.n38 gnd 0.006041f
C276 output.n39 gnd 0.006397f
C277 output.n40 gnd 0.01428f
C278 output.n41 gnd 0.030913f
C279 output.n42 gnd 0.006397f
C280 output.n43 gnd 0.006041f
C281 output.n44 gnd 0.025987f
C282 output.n45 gnd 0.097665f
C283 output.n46 gnd 0.015803f
C284 output.n47 gnd 0.011243f
C285 output.n48 gnd 0.006041f
C286 output.n49 gnd 0.01428f
C287 output.n50 gnd 0.006397f
C288 output.n51 gnd 0.011243f
C289 output.n52 gnd 0.006041f
C290 output.n53 gnd 0.01428f
C291 output.n54 gnd 0.006397f
C292 output.n55 gnd 0.048111f
C293 output.t0 gnd 0.023274f
C294 output.n56 gnd 0.01071f
C295 output.n57 gnd 0.008435f
C296 output.n58 gnd 0.006041f
C297 output.n59 gnd 0.267512f
C298 output.n60 gnd 0.011243f
C299 output.n61 gnd 0.006041f
C300 output.n62 gnd 0.006397f
C301 output.n63 gnd 0.01428f
C302 output.n64 gnd 0.01428f
C303 output.n65 gnd 0.006397f
C304 output.n66 gnd 0.006041f
C305 output.n67 gnd 0.011243f
C306 output.n68 gnd 0.011243f
C307 output.n69 gnd 0.006041f
C308 output.n70 gnd 0.006397f
C309 output.n71 gnd 0.01428f
C310 output.n72 gnd 0.030913f
C311 output.n73 gnd 0.006397f
C312 output.n74 gnd 0.006041f
C313 output.n75 gnd 0.025987f
C314 output.n76 gnd 0.09306f
C315 output.n77 gnd 1.65264f
C316 output.n78 gnd 0.015803f
C317 output.n79 gnd 0.011243f
C318 output.n80 gnd 0.006041f
C319 output.n81 gnd 0.01428f
C320 output.n82 gnd 0.006397f
C321 output.n83 gnd 0.011243f
C322 output.n84 gnd 0.006041f
C323 output.n85 gnd 0.01428f
C324 output.n86 gnd 0.006397f
C325 output.n87 gnd 0.048111f
C326 output.t2 gnd 0.023274f
C327 output.n88 gnd 0.01071f
C328 output.n89 gnd 0.008435f
C329 output.n90 gnd 0.006041f
C330 output.n91 gnd 0.267512f
C331 output.n92 gnd 0.011243f
C332 output.n93 gnd 0.006041f
C333 output.n94 gnd 0.006397f
C334 output.n95 gnd 0.01428f
C335 output.n96 gnd 0.01428f
C336 output.n97 gnd 0.006397f
C337 output.n98 gnd 0.006041f
C338 output.n99 gnd 0.011243f
C339 output.n100 gnd 0.011243f
C340 output.n101 gnd 0.006041f
C341 output.n102 gnd 0.006397f
C342 output.n103 gnd 0.01428f
C343 output.n104 gnd 0.030913f
C344 output.n105 gnd 0.006397f
C345 output.n106 gnd 0.006041f
C346 output.n107 gnd 0.025987f
C347 output.n108 gnd 0.09306f
C348 output.n109 gnd 0.713089f
C349 output.n110 gnd 0.015803f
C350 output.n111 gnd 0.011243f
C351 output.n112 gnd 0.006041f
C352 output.n113 gnd 0.01428f
C353 output.n114 gnd 0.006397f
C354 output.n115 gnd 0.011243f
C355 output.n116 gnd 0.006041f
C356 output.n117 gnd 0.01428f
C357 output.n118 gnd 0.006397f
C358 output.n119 gnd 0.048111f
C359 output.t3 gnd 0.023274f
C360 output.n120 gnd 0.01071f
C361 output.n121 gnd 0.008435f
C362 output.n122 gnd 0.006041f
C363 output.n123 gnd 0.267512f
C364 output.n124 gnd 0.011243f
C365 output.n125 gnd 0.006041f
C366 output.n126 gnd 0.006397f
C367 output.n127 gnd 0.01428f
C368 output.n128 gnd 0.01428f
C369 output.n129 gnd 0.006397f
C370 output.n130 gnd 0.006041f
C371 output.n131 gnd 0.011243f
C372 output.n132 gnd 0.011243f
C373 output.n133 gnd 0.006041f
C374 output.n134 gnd 0.006397f
C375 output.n135 gnd 0.01428f
C376 output.n136 gnd 0.030913f
C377 output.n137 gnd 0.006397f
C378 output.n138 gnd 0.006041f
C379 output.n139 gnd 0.025987f
C380 output.n140 gnd 0.09306f
C381 output.n141 gnd 1.67353f
C382 minus.n0 gnd 0.032421f
C383 minus.n1 gnd 0.007357f
C384 minus.n2 gnd 0.032421f
C385 minus.n3 gnd 0.007357f
C386 minus.n4 gnd 0.032421f
C387 minus.n5 gnd 0.007357f
C388 minus.n6 gnd 0.032421f
C389 minus.n7 gnd 0.007357f
C390 minus.n8 gnd 0.032421f
C391 minus.n9 gnd 0.007357f
C392 minus.t8 gnd 0.47521f
C393 minus.t7 gnd 0.458565f
C394 minus.n10 gnd 0.210344f
C395 minus.n11 gnd 0.18879f
C396 minus.n12 gnd 0.139574f
C397 minus.n13 gnd 0.032421f
C398 minus.t11 gnd 0.458565f
C399 minus.n14 gnd 0.203709f
C400 minus.n15 gnd 0.007357f
C401 minus.t10 gnd 0.458565f
C402 minus.n16 gnd 0.203709f
C403 minus.n17 gnd 0.032421f
C404 minus.n18 gnd 0.032421f
C405 minus.n19 gnd 0.032421f
C406 minus.t12 gnd 0.458565f
C407 minus.n20 gnd 0.203709f
C408 minus.n21 gnd 0.007357f
C409 minus.t20 gnd 0.458565f
C410 minus.n22 gnd 0.203709f
C411 minus.n23 gnd 0.032421f
C412 minus.n24 gnd 0.032421f
C413 minus.n25 gnd 0.032421f
C414 minus.t18 gnd 0.458565f
C415 minus.n26 gnd 0.203709f
C416 minus.n27 gnd 0.007357f
C417 minus.t25 gnd 0.458565f
C418 minus.n28 gnd 0.203709f
C419 minus.n29 gnd 0.032421f
C420 minus.n30 gnd 0.032421f
C421 minus.n31 gnd 0.032421f
C422 minus.t24 gnd 0.458565f
C423 minus.n32 gnd 0.203709f
C424 minus.n33 gnd 0.007357f
C425 minus.t14 gnd 0.458565f
C426 minus.n34 gnd 0.203709f
C427 minus.n35 gnd 0.032421f
C428 minus.n36 gnd 0.032421f
C429 minus.n37 gnd 0.032421f
C430 minus.t22 gnd 0.458565f
C431 minus.n38 gnd 0.203709f
C432 minus.n39 gnd 0.007357f
C433 minus.t19 gnd 0.458565f
C434 minus.n40 gnd 0.204009f
C435 minus.n41 gnd 0.375467f
C436 minus.n42 gnd 0.032421f
C437 minus.t13 gnd 0.458565f
C438 minus.t15 gnd 0.458565f
C439 minus.n43 gnd 0.032421f
C440 minus.t5 gnd 0.458565f
C441 minus.n44 gnd 0.203709f
C442 minus.n45 gnd 0.032421f
C443 minus.t6 gnd 0.458565f
C444 minus.t26 gnd 0.458565f
C445 minus.n46 gnd 0.203709f
C446 minus.n47 gnd 0.032421f
C447 minus.t21 gnd 0.458565f
C448 minus.t23 gnd 0.458565f
C449 minus.n48 gnd 0.203709f
C450 minus.n49 gnd 0.032421f
C451 minus.t16 gnd 0.458565f
C452 minus.t17 gnd 0.458565f
C453 minus.n50 gnd 0.203709f
C454 minus.n51 gnd 0.032421f
C455 minus.t9 gnd 0.458565f
C456 minus.t27 gnd 0.458565f
C457 minus.n52 gnd 0.210344f
C458 minus.t28 gnd 0.47521f
C459 minus.n53 gnd 0.18879f
C460 minus.n54 gnd 0.139574f
C461 minus.n55 gnd 0.007357f
C462 minus.n56 gnd 0.203709f
C463 minus.n57 gnd 0.007357f
C464 minus.n58 gnd 0.032421f
C465 minus.n59 gnd 0.032421f
C466 minus.n60 gnd 0.032421f
C467 minus.n61 gnd 0.007357f
C468 minus.n62 gnd 0.203709f
C469 minus.n63 gnd 0.007357f
C470 minus.n64 gnd 0.032421f
C471 minus.n65 gnd 0.032421f
C472 minus.n66 gnd 0.032421f
C473 minus.n67 gnd 0.007357f
C474 minus.n68 gnd 0.203709f
C475 minus.n69 gnd 0.007357f
C476 minus.n70 gnd 0.032421f
C477 minus.n71 gnd 0.032421f
C478 minus.n72 gnd 0.032421f
C479 minus.n73 gnd 0.007357f
C480 minus.n74 gnd 0.203709f
C481 minus.n75 gnd 0.007357f
C482 minus.n76 gnd 0.032421f
C483 minus.n77 gnd 0.032421f
C484 minus.n78 gnd 0.032421f
C485 minus.n79 gnd 0.007357f
C486 minus.n80 gnd 0.203709f
C487 minus.n81 gnd 0.007357f
C488 minus.n82 gnd 0.204009f
C489 minus.n83 gnd 1.08613f
C490 minus.n84 gnd 1.61832f
C491 minus.t1 gnd 0.009994f
C492 minus.t0 gnd 0.009994f
C493 minus.n85 gnd 0.032864f
C494 minus.t4 gnd 0.009994f
C495 minus.t3 gnd 0.009994f
C496 minus.n86 gnd 0.032414f
C497 minus.n87 gnd 0.276636f
C498 minus.t2 gnd 0.055628f
C499 minus.n88 gnd 0.150958f
C500 minus.n89 gnd 1.94905f
C501 a_n2982_8322.t7 gnd 0.100195f
C502 a_n2982_8322.t37 gnd 20.7864f
C503 a_n2982_8322.t34 gnd 20.640598f
C504 a_n2982_8322.t36 gnd 20.640598f
C505 a_n2982_8322.t32 gnd 20.7864f
C506 a_n2982_8322.t35 gnd 20.640598f
C507 a_n2982_8322.t33 gnd 28.793001f
C508 a_n2982_8322.t6 gnd 0.938175f
C509 a_n2982_8322.t19 gnd 0.100195f
C510 a_n2982_8322.t15 gnd 0.100195f
C511 a_n2982_8322.n0 gnd 0.705774f
C512 a_n2982_8322.n1 gnd 0.788598f
C513 a_n2982_8322.t22 gnd 0.100195f
C514 a_n2982_8322.t12 gnd 0.100195f
C515 a_n2982_8322.n2 gnd 0.705774f
C516 a_n2982_8322.n3 gnd 0.400677f
C517 a_n2982_8322.t3 gnd 0.100195f
C518 a_n2982_8322.t2 gnd 0.100195f
C519 a_n2982_8322.n4 gnd 0.705774f
C520 a_n2982_8322.n5 gnd 0.400677f
C521 a_n2982_8322.t16 gnd 0.100195f
C522 a_n2982_8322.t9 gnd 0.100195f
C523 a_n2982_8322.n6 gnd 0.705774f
C524 a_n2982_8322.n7 gnd 0.400677f
C525 a_n2982_8322.t13 gnd 0.100195f
C526 a_n2982_8322.t11 gnd 0.100195f
C527 a_n2982_8322.n8 gnd 0.705774f
C528 a_n2982_8322.n9 gnd 0.400677f
C529 a_n2982_8322.t0 gnd 0.936307f
C530 a_n2982_8322.n10 gnd 1.87205f
C531 a_n2982_8322.t27 gnd 0.938175f
C532 a_n2982_8322.t31 gnd 0.100195f
C533 a_n2982_8322.t30 gnd 0.100195f
C534 a_n2982_8322.n11 gnd 0.705774f
C535 a_n2982_8322.n12 gnd 0.788598f
C536 a_n2982_8322.t25 gnd 0.936307f
C537 a_n2982_8322.n13 gnd 0.396834f
C538 a_n2982_8322.t28 gnd 0.936307f
C539 a_n2982_8322.n14 gnd 0.396834f
C540 a_n2982_8322.t26 gnd 0.100195f
C541 a_n2982_8322.t24 gnd 0.100195f
C542 a_n2982_8322.n15 gnd 0.705774f
C543 a_n2982_8322.n16 gnd 0.400677f
C544 a_n2982_8322.t29 gnd 0.936307f
C545 a_n2982_8322.n17 gnd 1.47193f
C546 a_n2982_8322.n18 gnd 2.35218f
C547 a_n2982_8322.n19 gnd 3.2687f
C548 a_n2982_8322.t1 gnd 0.936307f
C549 a_n2982_8322.n20 gnd 1.11185f
C550 a_n2982_8322.t18 gnd 0.100195f
C551 a_n2982_8322.t17 gnd 0.100195f
C552 a_n2982_8322.n21 gnd 0.705774f
C553 a_n2982_8322.n22 gnd 0.400677f
C554 a_n2982_8322.t5 gnd 0.100195f
C555 a_n2982_8322.t4 gnd 0.100195f
C556 a_n2982_8322.n23 gnd 0.705774f
C557 a_n2982_8322.n24 gnd 0.400677f
C558 a_n2982_8322.t20 gnd 0.100195f
C559 a_n2982_8322.t8 gnd 0.100195f
C560 a_n2982_8322.n25 gnd 0.705774f
C561 a_n2982_8322.n26 gnd 0.400677f
C562 a_n2982_8322.t21 gnd 0.938173f
C563 a_n2982_8322.t14 gnd 0.100195f
C564 a_n2982_8322.t10 gnd 0.100195f
C565 a_n2982_8322.n27 gnd 0.705774f
C566 a_n2982_8322.n28 gnd 0.7886f
C567 a_n2982_8322.n29 gnd 0.400675f
C568 a_n2982_8322.n30 gnd 0.705776f
C569 a_n2982_8322.t23 gnd 0.100195f
C570 CSoutput.n0 gnd 0.041891f
C571 CSoutput.t174 gnd 0.277101f
C572 CSoutput.n1 gnd 0.125125f
C573 CSoutput.n2 gnd 0.041891f
C574 CSoutput.t181 gnd 0.277101f
C575 CSoutput.n3 gnd 0.033202f
C576 CSoutput.n4 gnd 0.041891f
C577 CSoutput.t188 gnd 0.277101f
C578 CSoutput.n5 gnd 0.028631f
C579 CSoutput.n6 gnd 0.041891f
C580 CSoutput.t179 gnd 0.277101f
C581 CSoutput.t177 gnd 0.277101f
C582 CSoutput.n7 gnd 0.123761f
C583 CSoutput.n8 gnd 0.041891f
C584 CSoutput.t186 gnd 0.277101f
C585 CSoutput.n9 gnd 0.027298f
C586 CSoutput.n10 gnd 0.041891f
C587 CSoutput.t169 gnd 0.277101f
C588 CSoutput.t173 gnd 0.277101f
C589 CSoutput.n11 gnd 0.123761f
C590 CSoutput.n12 gnd 0.041891f
C591 CSoutput.t184 gnd 0.277101f
C592 CSoutput.n13 gnd 0.028631f
C593 CSoutput.n14 gnd 0.041891f
C594 CSoutput.t183 gnd 0.277101f
C595 CSoutput.t171 gnd 0.277101f
C596 CSoutput.n15 gnd 0.123761f
C597 CSoutput.n16 gnd 0.041891f
C598 CSoutput.t176 gnd 0.277101f
C599 CSoutput.n17 gnd 0.030579f
C600 CSoutput.t185 gnd 0.331143f
C601 CSoutput.t182 gnd 0.277101f
C602 CSoutput.n18 gnd 0.157995f
C603 CSoutput.n19 gnd 0.15331f
C604 CSoutput.n20 gnd 0.177858f
C605 CSoutput.n21 gnd 0.041891f
C606 CSoutput.n22 gnd 0.034963f
C607 CSoutput.n23 gnd 0.123761f
C608 CSoutput.n24 gnd 0.033703f
C609 CSoutput.n25 gnd 0.033202f
C610 CSoutput.n26 gnd 0.041891f
C611 CSoutput.n27 gnd 0.041891f
C612 CSoutput.n28 gnd 0.034694f
C613 CSoutput.n29 gnd 0.029456f
C614 CSoutput.n30 gnd 0.126516f
C615 CSoutput.n31 gnd 0.029862f
C616 CSoutput.n32 gnd 0.041891f
C617 CSoutput.n33 gnd 0.041891f
C618 CSoutput.n34 gnd 0.041891f
C619 CSoutput.n35 gnd 0.034325f
C620 CSoutput.n36 gnd 0.123761f
C621 CSoutput.n37 gnd 0.032826f
C622 CSoutput.n38 gnd 0.034079f
C623 CSoutput.n39 gnd 0.041891f
C624 CSoutput.n40 gnd 0.041891f
C625 CSoutput.n41 gnd 0.034956f
C626 CSoutput.n42 gnd 0.03195f
C627 CSoutput.n43 gnd 0.123761f
C628 CSoutput.n44 gnd 0.03276f
C629 CSoutput.n45 gnd 0.041891f
C630 CSoutput.n46 gnd 0.041891f
C631 CSoutput.n47 gnd 0.041891f
C632 CSoutput.n48 gnd 0.03276f
C633 CSoutput.n49 gnd 0.123761f
C634 CSoutput.n50 gnd 0.03195f
C635 CSoutput.n51 gnd 0.034956f
C636 CSoutput.n52 gnd 0.041891f
C637 CSoutput.n53 gnd 0.041891f
C638 CSoutput.n54 gnd 0.034079f
C639 CSoutput.n55 gnd 0.032826f
C640 CSoutput.n56 gnd 0.123761f
C641 CSoutput.n57 gnd 0.034325f
C642 CSoutput.n58 gnd 0.041891f
C643 CSoutput.n59 gnd 0.041891f
C644 CSoutput.n60 gnd 0.041891f
C645 CSoutput.n61 gnd 0.029862f
C646 CSoutput.n62 gnd 0.126516f
C647 CSoutput.n63 gnd 0.029456f
C648 CSoutput.t180 gnd 0.277101f
C649 CSoutput.n64 gnd 0.123761f
C650 CSoutput.n65 gnd 0.034694f
C651 CSoutput.n66 gnd 0.041891f
C652 CSoutput.n67 gnd 0.041891f
C653 CSoutput.n68 gnd 0.041891f
C654 CSoutput.n69 gnd 0.033703f
C655 CSoutput.n70 gnd 0.123761f
C656 CSoutput.n71 gnd 0.034963f
C657 CSoutput.n72 gnd 0.030579f
C658 CSoutput.n73 gnd 0.041891f
C659 CSoutput.n74 gnd 0.041891f
C660 CSoutput.n75 gnd 0.031712f
C661 CSoutput.n76 gnd 0.018834f
C662 CSoutput.t187 gnd 0.311343f
C663 CSoutput.n77 gnd 0.154663f
C664 CSoutput.n78 gnd 0.632717f
C665 CSoutput.t71 gnd 0.052253f
C666 CSoutput.t35 gnd 0.052253f
C667 CSoutput.n79 gnd 0.404563f
C668 CSoutput.t10 gnd 0.052253f
C669 CSoutput.t61 gnd 0.052253f
C670 CSoutput.n80 gnd 0.403842f
C671 CSoutput.n81 gnd 0.409899f
C672 CSoutput.t17 gnd 0.052253f
C673 CSoutput.t47 gnd 0.052253f
C674 CSoutput.n82 gnd 0.403842f
C675 CSoutput.n83 gnd 0.201981f
C676 CSoutput.t29 gnd 0.052253f
C677 CSoutput.t41 gnd 0.052253f
C678 CSoutput.n84 gnd 0.403842f
C679 CSoutput.n85 gnd 0.201981f
C680 CSoutput.t38 gnd 0.052253f
C681 CSoutput.t65 gnd 0.052253f
C682 CSoutput.n86 gnd 0.403842f
C683 CSoutput.n87 gnd 0.201981f
C684 CSoutput.t21 gnd 0.052253f
C685 CSoutput.t52 gnd 0.052253f
C686 CSoutput.n88 gnd 0.403842f
C687 CSoutput.n89 gnd 0.370386f
C688 CSoutput.t39 gnd 0.052253f
C689 CSoutput.t18 gnd 0.052253f
C690 CSoutput.n90 gnd 0.404563f
C691 CSoutput.t4 gnd 0.052253f
C692 CSoutput.t40 gnd 0.052253f
C693 CSoutput.n91 gnd 0.403842f
C694 CSoutput.n92 gnd 0.409899f
C695 CSoutput.t36 gnd 0.052253f
C696 CSoutput.t16 gnd 0.052253f
C697 CSoutput.n93 gnd 0.403842f
C698 CSoutput.n94 gnd 0.201981f
C699 CSoutput.t3 gnd 0.052253f
C700 CSoutput.t1 gnd 0.052253f
C701 CSoutput.n95 gnd 0.403842f
C702 CSoutput.n96 gnd 0.201981f
C703 CSoutput.t48 gnd 0.052253f
C704 CSoutput.t26 gnd 0.052253f
C705 CSoutput.n97 gnd 0.403842f
C706 CSoutput.n98 gnd 0.201981f
C707 CSoutput.t23 gnd 0.052253f
C708 CSoutput.t0 gnd 0.052253f
C709 CSoutput.n99 gnd 0.403842f
C710 CSoutput.n100 gnd 0.301204f
C711 CSoutput.n101 gnd 0.379816f
C712 CSoutput.t44 gnd 0.052253f
C713 CSoutput.t27 gnd 0.052253f
C714 CSoutput.n102 gnd 0.404563f
C715 CSoutput.t13 gnd 0.052253f
C716 CSoutput.t45 gnd 0.052253f
C717 CSoutput.n103 gnd 0.403842f
C718 CSoutput.n104 gnd 0.409899f
C719 CSoutput.t43 gnd 0.052253f
C720 CSoutput.t25 gnd 0.052253f
C721 CSoutput.n105 gnd 0.403842f
C722 CSoutput.n106 gnd 0.201981f
C723 CSoutput.t12 gnd 0.052253f
C724 CSoutput.t11 gnd 0.052253f
C725 CSoutput.n107 gnd 0.403842f
C726 CSoutput.n108 gnd 0.201981f
C727 CSoutput.t54 gnd 0.052253f
C728 CSoutput.t32 gnd 0.052253f
C729 CSoutput.n109 gnd 0.403842f
C730 CSoutput.n110 gnd 0.201981f
C731 CSoutput.t30 gnd 0.052253f
C732 CSoutput.t8 gnd 0.052253f
C733 CSoutput.n111 gnd 0.403842f
C734 CSoutput.n112 gnd 0.301204f
C735 CSoutput.n113 gnd 0.424538f
C736 CSoutput.n114 gnd 7.90743f
C737 CSoutput.n116 gnd 0.741048f
C738 CSoutput.n117 gnd 0.555786f
C739 CSoutput.n118 gnd 0.741048f
C740 CSoutput.n119 gnd 0.741048f
C741 CSoutput.n120 gnd 1.99513f
C742 CSoutput.n121 gnd 0.741048f
C743 CSoutput.n122 gnd 0.741048f
C744 CSoutput.t175 gnd 0.92631f
C745 CSoutput.n123 gnd 0.741048f
C746 CSoutput.n124 gnd 0.741048f
C747 CSoutput.n128 gnd 0.741048f
C748 CSoutput.n132 gnd 0.741048f
C749 CSoutput.n133 gnd 0.741048f
C750 CSoutput.n135 gnd 0.741048f
C751 CSoutput.n140 gnd 0.741048f
C752 CSoutput.n142 gnd 0.741048f
C753 CSoutput.n143 gnd 0.741048f
C754 CSoutput.n145 gnd 0.741048f
C755 CSoutput.n146 gnd 0.741048f
C756 CSoutput.n148 gnd 0.741048f
C757 CSoutput.t170 gnd 12.3828f
C758 CSoutput.n150 gnd 0.741048f
C759 CSoutput.n151 gnd 0.555786f
C760 CSoutput.n152 gnd 0.741048f
C761 CSoutput.n153 gnd 0.741048f
C762 CSoutput.n154 gnd 1.99513f
C763 CSoutput.n155 gnd 0.741048f
C764 CSoutput.n156 gnd 0.741048f
C765 CSoutput.t189 gnd 0.92631f
C766 CSoutput.n157 gnd 0.741048f
C767 CSoutput.n158 gnd 0.741048f
C768 CSoutput.n162 gnd 0.741048f
C769 CSoutput.n166 gnd 0.741048f
C770 CSoutput.n167 gnd 0.741048f
C771 CSoutput.n169 gnd 0.741048f
C772 CSoutput.n174 gnd 0.741048f
C773 CSoutput.n176 gnd 0.741048f
C774 CSoutput.n177 gnd 0.741048f
C775 CSoutput.n179 gnd 0.741048f
C776 CSoutput.n180 gnd 0.741048f
C777 CSoutput.n182 gnd 0.741048f
C778 CSoutput.n183 gnd 0.555786f
C779 CSoutput.n185 gnd 0.741048f
C780 CSoutput.n186 gnd 0.555786f
C781 CSoutput.n187 gnd 0.741048f
C782 CSoutput.n188 gnd 0.741048f
C783 CSoutput.n189 gnd 1.99513f
C784 CSoutput.n190 gnd 0.741048f
C785 CSoutput.n191 gnd 0.741048f
C786 CSoutput.t168 gnd 0.92631f
C787 CSoutput.n192 gnd 0.741048f
C788 CSoutput.n193 gnd 1.99513f
C789 CSoutput.n195 gnd 0.741048f
C790 CSoutput.n196 gnd 0.741048f
C791 CSoutput.n198 gnd 0.741048f
C792 CSoutput.n199 gnd 0.741048f
C793 CSoutput.t178 gnd 12.181001f
C794 CSoutput.t172 gnd 12.3828f
C795 CSoutput.n205 gnd 2.32478f
C796 CSoutput.n206 gnd 9.47029f
C797 CSoutput.n207 gnd 9.86657f
C798 CSoutput.n212 gnd 2.51836f
C799 CSoutput.n218 gnd 0.741048f
C800 CSoutput.n220 gnd 0.741048f
C801 CSoutput.n222 gnd 0.741048f
C802 CSoutput.n224 gnd 0.741048f
C803 CSoutput.n226 gnd 0.741048f
C804 CSoutput.n232 gnd 0.741048f
C805 CSoutput.n239 gnd 1.35954f
C806 CSoutput.n240 gnd 1.35954f
C807 CSoutput.n241 gnd 0.741048f
C808 CSoutput.n242 gnd 0.741048f
C809 CSoutput.n244 gnd 0.555786f
C810 CSoutput.n245 gnd 0.475981f
C811 CSoutput.n247 gnd 0.555786f
C812 CSoutput.n248 gnd 0.475981f
C813 CSoutput.n249 gnd 0.555786f
C814 CSoutput.n251 gnd 0.741048f
C815 CSoutput.n253 gnd 1.99513f
C816 CSoutput.n254 gnd 2.32478f
C817 CSoutput.n255 gnd 8.710231f
C818 CSoutput.n257 gnd 0.555786f
C819 CSoutput.n258 gnd 1.43007f
C820 CSoutput.n259 gnd 0.555786f
C821 CSoutput.n261 gnd 0.741048f
C822 CSoutput.n263 gnd 1.99513f
C823 CSoutput.n264 gnd 4.34571f
C824 CSoutput.t34 gnd 0.052253f
C825 CSoutput.t20 gnd 0.052253f
C826 CSoutput.n265 gnd 0.404563f
C827 CSoutput.t60 gnd 0.052253f
C828 CSoutput.t9 gnd 0.052253f
C829 CSoutput.n266 gnd 0.403842f
C830 CSoutput.n267 gnd 0.409899f
C831 CSoutput.t46 gnd 0.052253f
C832 CSoutput.t14 gnd 0.052253f
C833 CSoutput.n268 gnd 0.403842f
C834 CSoutput.n269 gnd 0.201981f
C835 CSoutput.t56 gnd 0.052253f
C836 CSoutput.t28 gnd 0.052253f
C837 CSoutput.n270 gnd 0.403842f
C838 CSoutput.n271 gnd 0.201981f
C839 CSoutput.t64 gnd 0.052253f
C840 CSoutput.t37 gnd 0.052253f
C841 CSoutput.n272 gnd 0.403842f
C842 CSoutput.n273 gnd 0.201981f
C843 CSoutput.t51 gnd 0.052253f
C844 CSoutput.t22 gnd 0.052253f
C845 CSoutput.n274 gnd 0.403842f
C846 CSoutput.n275 gnd 0.370386f
C847 CSoutput.t62 gnd 0.052253f
C848 CSoutput.t63 gnd 0.052253f
C849 CSoutput.n276 gnd 0.404563f
C850 CSoutput.t7 gnd 0.052253f
C851 CSoutput.t53 gnd 0.052253f
C852 CSoutput.n277 gnd 0.403842f
C853 CSoutput.n278 gnd 0.409899f
C854 CSoutput.t59 gnd 0.052253f
C855 CSoutput.t5 gnd 0.052253f
C856 CSoutput.n279 gnd 0.403842f
C857 CSoutput.n280 gnd 0.201981f
C858 CSoutput.t33 gnd 0.052253f
C859 CSoutput.t50 gnd 0.052253f
C860 CSoutput.n281 gnd 0.403842f
C861 CSoutput.n282 gnd 0.201981f
C862 CSoutput.t67 gnd 0.052253f
C863 CSoutput.t24 gnd 0.052253f
C864 CSoutput.n283 gnd 0.403842f
C865 CSoutput.n284 gnd 0.201981f
C866 CSoutput.t49 gnd 0.052253f
C867 CSoutput.t70 gnd 0.052253f
C868 CSoutput.n285 gnd 0.403842f
C869 CSoutput.n286 gnd 0.301204f
C870 CSoutput.n287 gnd 0.379816f
C871 CSoutput.t68 gnd 0.052253f
C872 CSoutput.t69 gnd 0.052253f
C873 CSoutput.n288 gnd 0.404563f
C874 CSoutput.t19 gnd 0.052253f
C875 CSoutput.t58 gnd 0.052253f
C876 CSoutput.n289 gnd 0.403842f
C877 CSoutput.n290 gnd 0.409899f
C878 CSoutput.t66 gnd 0.052253f
C879 CSoutput.t15 gnd 0.052253f
C880 CSoutput.n291 gnd 0.403842f
C881 CSoutput.n292 gnd 0.201981f
C882 CSoutput.t42 gnd 0.052253f
C883 CSoutput.t57 gnd 0.052253f
C884 CSoutput.n293 gnd 0.403842f
C885 CSoutput.n294 gnd 0.201981f
C886 CSoutput.t2 gnd 0.052253f
C887 CSoutput.t31 gnd 0.052253f
C888 CSoutput.n295 gnd 0.403842f
C889 CSoutput.n296 gnd 0.201981f
C890 CSoutput.t55 gnd 0.052253f
C891 CSoutput.t6 gnd 0.052253f
C892 CSoutput.n297 gnd 0.40384f
C893 CSoutput.n298 gnd 0.301206f
C894 CSoutput.n299 gnd 0.424538f
C895 CSoutput.n300 gnd 11.292099f
C896 CSoutput.t111 gnd 0.045722f
C897 CSoutput.t164 gnd 0.045722f
C898 CSoutput.n301 gnd 0.405365f
C899 CSoutput.t105 gnd 0.045722f
C900 CSoutput.t110 gnd 0.045722f
C901 CSoutput.n302 gnd 0.404013f
C902 CSoutput.n303 gnd 0.376465f
C903 CSoutput.t95 gnd 0.045722f
C904 CSoutput.t114 gnd 0.045722f
C905 CSoutput.n304 gnd 0.404013f
C906 CSoutput.n305 gnd 0.185579f
C907 CSoutput.t129 gnd 0.045722f
C908 CSoutput.t106 gnd 0.045722f
C909 CSoutput.n306 gnd 0.404013f
C910 CSoutput.n307 gnd 0.185579f
C911 CSoutput.t113 gnd 0.045722f
C912 CSoutput.t155 gnd 0.045722f
C913 CSoutput.n308 gnd 0.404013f
C914 CSoutput.n309 gnd 0.185579f
C915 CSoutput.t125 gnd 0.045722f
C916 CSoutput.t135 gnd 0.045722f
C917 CSoutput.n310 gnd 0.404013f
C918 CSoutput.n311 gnd 0.185579f
C919 CSoutput.t90 gnd 0.045722f
C920 CSoutput.t115 gnd 0.045722f
C921 CSoutput.n312 gnd 0.404013f
C922 CSoutput.n313 gnd 0.185579f
C923 CSoutput.t79 gnd 0.045722f
C924 CSoutput.t102 gnd 0.045722f
C925 CSoutput.n314 gnd 0.404013f
C926 CSoutput.n315 gnd 0.342291f
C927 CSoutput.t160 gnd 0.045722f
C928 CSoutput.t72 gnd 0.045722f
C929 CSoutput.n316 gnd 0.405365f
C930 CSoutput.t83 gnd 0.045722f
C931 CSoutput.t153 gnd 0.045722f
C932 CSoutput.n317 gnd 0.404013f
C933 CSoutput.n318 gnd 0.376465f
C934 CSoutput.t74 gnd 0.045722f
C935 CSoutput.t146 gnd 0.045722f
C936 CSoutput.n319 gnd 0.404013f
C937 CSoutput.n320 gnd 0.185579f
C938 CSoutput.t154 gnd 0.045722f
C939 CSoutput.t73 gnd 0.045722f
C940 CSoutput.n321 gnd 0.404013f
C941 CSoutput.n322 gnd 0.185579f
C942 CSoutput.t137 gnd 0.045722f
C943 CSoutput.t118 gnd 0.045722f
C944 CSoutput.n323 gnd 0.404013f
C945 CSoutput.n324 gnd 0.185579f
C946 CSoutput.t75 gnd 0.045722f
C947 CSoutput.t139 gnd 0.045722f
C948 CSoutput.n325 gnd 0.404013f
C949 CSoutput.n326 gnd 0.185579f
C950 CSoutput.t120 gnd 0.045722f
C951 CSoutput.t126 gnd 0.045722f
C952 CSoutput.n327 gnd 0.404013f
C953 CSoutput.n328 gnd 0.185579f
C954 CSoutput.t138 gnd 0.045722f
C955 CSoutput.t119 gnd 0.045722f
C956 CSoutput.n329 gnd 0.404013f
C957 CSoutput.n330 gnd 0.281749f
C958 CSoutput.n331 gnd 0.355373f
C959 CSoutput.t84 gnd 0.045722f
C960 CSoutput.t156 gnd 0.045722f
C961 CSoutput.n332 gnd 0.405365f
C962 CSoutput.t103 gnd 0.045722f
C963 CSoutput.t107 gnd 0.045722f
C964 CSoutput.n333 gnd 0.404013f
C965 CSoutput.n334 gnd 0.376465f
C966 CSoutput.t76 gnd 0.045722f
C967 CSoutput.t141 gnd 0.045722f
C968 CSoutput.n335 gnd 0.404013f
C969 CSoutput.n336 gnd 0.185579f
C970 CSoutput.t112 gnd 0.045722f
C971 CSoutput.t85 gnd 0.045722f
C972 CSoutput.n337 gnd 0.404013f
C973 CSoutput.n338 gnd 0.185579f
C974 CSoutput.t93 gnd 0.045722f
C975 CSoutput.t167 gnd 0.045722f
C976 CSoutput.n339 gnd 0.404013f
C977 CSoutput.n340 gnd 0.185579f
C978 CSoutput.t94 gnd 0.045722f
C979 CSoutput.t98 gnd 0.045722f
C980 CSoutput.n341 gnd 0.404013f
C981 CSoutput.n342 gnd 0.185579f
C982 CSoutput.t82 gnd 0.045722f
C983 CSoutput.t152 gnd 0.045722f
C984 CSoutput.n343 gnd 0.404013f
C985 CSoutput.n344 gnd 0.185579f
C986 CSoutput.t101 gnd 0.045722f
C987 CSoutput.t91 gnd 0.045722f
C988 CSoutput.n345 gnd 0.404013f
C989 CSoutput.n346 gnd 0.281749f
C990 CSoutput.n347 gnd 0.381615f
C991 CSoutput.n348 gnd 11.4493f
C992 CSoutput.t97 gnd 0.045722f
C993 CSoutput.t140 gnd 0.045722f
C994 CSoutput.n349 gnd 0.405365f
C995 CSoutput.t136 gnd 0.045722f
C996 CSoutput.t117 gnd 0.045722f
C997 CSoutput.n350 gnd 0.404013f
C998 CSoutput.n351 gnd 0.376465f
C999 CSoutput.t143 gnd 0.045722f
C1000 CSoutput.t108 gnd 0.045722f
C1001 CSoutput.n352 gnd 0.404013f
C1002 CSoutput.n353 gnd 0.185579f
C1003 CSoutput.t127 gnd 0.045722f
C1004 CSoutput.t158 gnd 0.045722f
C1005 CSoutput.n354 gnd 0.404013f
C1006 CSoutput.n355 gnd 0.185579f
C1007 CSoutput.t92 gnd 0.045722f
C1008 CSoutput.t142 gnd 0.045722f
C1009 CSoutput.n356 gnd 0.404013f
C1010 CSoutput.n357 gnd 0.185579f
C1011 CSoutput.t81 gnd 0.045722f
C1012 CSoutput.t148 gnd 0.045722f
C1013 CSoutput.n358 gnd 0.404013f
C1014 CSoutput.n359 gnd 0.185579f
C1015 CSoutput.t147 gnd 0.045722f
C1016 CSoutput.t104 gnd 0.045722f
C1017 CSoutput.n360 gnd 0.404013f
C1018 CSoutput.n361 gnd 0.185579f
C1019 CSoutput.t123 gnd 0.045722f
C1020 CSoutput.t100 gnd 0.045722f
C1021 CSoutput.n362 gnd 0.404013f
C1022 CSoutput.n363 gnd 0.342291f
C1023 CSoutput.t87 gnd 0.045722f
C1024 CSoutput.t80 gnd 0.045722f
C1025 CSoutput.n364 gnd 0.405365f
C1026 CSoutput.t77 gnd 0.045722f
C1027 CSoutput.t165 gnd 0.045722f
C1028 CSoutput.n365 gnd 0.404013f
C1029 CSoutput.n366 gnd 0.376465f
C1030 CSoutput.t166 gnd 0.045722f
C1031 CSoutput.t88 gnd 0.045722f
C1032 CSoutput.n367 gnd 0.404013f
C1033 CSoutput.n368 gnd 0.185579f
C1034 CSoutput.t89 gnd 0.045722f
C1035 CSoutput.t131 gnd 0.045722f
C1036 CSoutput.n369 gnd 0.404013f
C1037 CSoutput.n370 gnd 0.185579f
C1038 CSoutput.t132 gnd 0.045722f
C1039 CSoutput.t159 gnd 0.045722f
C1040 CSoutput.n371 gnd 0.404013f
C1041 CSoutput.n372 gnd 0.185579f
C1042 CSoutput.t162 gnd 0.045722f
C1043 CSoutput.t151 gnd 0.045722f
C1044 CSoutput.n373 gnd 0.404013f
C1045 CSoutput.n374 gnd 0.185579f
C1046 CSoutput.t145 gnd 0.045722f
C1047 CSoutput.t133 gnd 0.045722f
C1048 CSoutput.n375 gnd 0.404013f
C1049 CSoutput.n376 gnd 0.185579f
C1050 CSoutput.t134 gnd 0.045722f
C1051 CSoutput.t163 gnd 0.045722f
C1052 CSoutput.n377 gnd 0.404013f
C1053 CSoutput.n378 gnd 0.281749f
C1054 CSoutput.n379 gnd 0.355373f
C1055 CSoutput.t124 gnd 0.045722f
C1056 CSoutput.t149 gnd 0.045722f
C1057 CSoutput.n380 gnd 0.405365f
C1058 CSoutput.t96 gnd 0.045722f
C1059 CSoutput.t109 gnd 0.045722f
C1060 CSoutput.n381 gnd 0.404013f
C1061 CSoutput.n382 gnd 0.376465f
C1062 CSoutput.t116 gnd 0.045722f
C1063 CSoutput.t130 gnd 0.045722f
C1064 CSoutput.n383 gnd 0.404013f
C1065 CSoutput.n384 gnd 0.185579f
C1066 CSoutput.t150 gnd 0.045722f
C1067 CSoutput.t121 gnd 0.045722f
C1068 CSoutput.n385 gnd 0.404013f
C1069 CSoutput.n386 gnd 0.185579f
C1070 CSoutput.t128 gnd 0.045722f
C1071 CSoutput.t161 gnd 0.045722f
C1072 CSoutput.n387 gnd 0.404013f
C1073 CSoutput.n388 gnd 0.185579f
C1074 CSoutput.t78 gnd 0.045722f
C1075 CSoutput.t99 gnd 0.045722f
C1076 CSoutput.n389 gnd 0.404013f
C1077 CSoutput.n390 gnd 0.185579f
C1078 CSoutput.t122 gnd 0.045722f
C1079 CSoutput.t144 gnd 0.045722f
C1080 CSoutput.n391 gnd 0.404013f
C1081 CSoutput.n392 gnd 0.185579f
C1082 CSoutput.t157 gnd 0.045722f
C1083 CSoutput.t86 gnd 0.045722f
C1084 CSoutput.n393 gnd 0.404013f
C1085 CSoutput.n394 gnd 0.281749f
C1086 CSoutput.n395 gnd 0.381615f
C1087 CSoutput.n396 gnd 6.65687f
C1088 CSoutput.n397 gnd 12.6582f
C1089 commonsourceibias.n0 gnd 0.012624f
C1090 commonsourceibias.t120 gnd 0.191163f
C1091 commonsourceibias.t67 gnd 0.176757f
C1092 commonsourceibias.n1 gnd 0.00769f
C1093 commonsourceibias.n2 gnd 0.009461f
C1094 commonsourceibias.t126 gnd 0.176757f
C1095 commonsourceibias.n3 gnd 0.009597f
C1096 commonsourceibias.n4 gnd 0.009461f
C1097 commonsourceibias.t121 gnd 0.176757f
C1098 commonsourceibias.n5 gnd 0.070526f
C1099 commonsourceibias.t136 gnd 0.176757f
C1100 commonsourceibias.n6 gnd 0.007653f
C1101 commonsourceibias.n7 gnd 0.009461f
C1102 commonsourceibias.t117 gnd 0.176757f
C1103 commonsourceibias.n8 gnd 0.009134f
C1104 commonsourceibias.n9 gnd 0.009461f
C1105 commonsourceibias.t102 gnd 0.176757f
C1106 commonsourceibias.n10 gnd 0.070526f
C1107 commonsourceibias.t125 gnd 0.176757f
C1108 commonsourceibias.n11 gnd 0.007641f
C1109 commonsourceibias.n12 gnd 0.012624f
C1110 commonsourceibias.t12 gnd 0.191163f
C1111 commonsourceibias.t48 gnd 0.176757f
C1112 commonsourceibias.n13 gnd 0.00769f
C1113 commonsourceibias.n14 gnd 0.009461f
C1114 commonsourceibias.t4 gnd 0.176757f
C1115 commonsourceibias.n15 gnd 0.009597f
C1116 commonsourceibias.n16 gnd 0.009461f
C1117 commonsourceibias.t10 gnd 0.176757f
C1118 commonsourceibias.n17 gnd 0.070526f
C1119 commonsourceibias.t58 gnd 0.176757f
C1120 commonsourceibias.n18 gnd 0.007653f
C1121 commonsourceibias.n19 gnd 0.009461f
C1122 commonsourceibias.t16 gnd 0.176757f
C1123 commonsourceibias.n20 gnd 0.009134f
C1124 commonsourceibias.n21 gnd 0.009461f
C1125 commonsourceibias.t28 gnd 0.176757f
C1126 commonsourceibias.n22 gnd 0.070526f
C1127 commonsourceibias.t6 gnd 0.176757f
C1128 commonsourceibias.n23 gnd 0.007641f
C1129 commonsourceibias.n24 gnd 0.009461f
C1130 commonsourceibias.t14 gnd 0.176757f
C1131 commonsourceibias.t44 gnd 0.176757f
C1132 commonsourceibias.n25 gnd 0.070526f
C1133 commonsourceibias.n26 gnd 0.009461f
C1134 commonsourceibias.t24 gnd 0.176757f
C1135 commonsourceibias.n27 gnd 0.070526f
C1136 commonsourceibias.n28 gnd 0.009461f
C1137 commonsourceibias.t30 gnd 0.176757f
C1138 commonsourceibias.n29 gnd 0.070526f
C1139 commonsourceibias.n30 gnd 0.009461f
C1140 commonsourceibias.t54 gnd 0.176757f
C1141 commonsourceibias.n31 gnd 0.010754f
C1142 commonsourceibias.n32 gnd 0.009461f
C1143 commonsourceibias.t18 gnd 0.176757f
C1144 commonsourceibias.n33 gnd 0.012717f
C1145 commonsourceibias.t0 gnd 0.196904f
C1146 commonsourceibias.t50 gnd 0.176757f
C1147 commonsourceibias.n34 gnd 0.078584f
C1148 commonsourceibias.n35 gnd 0.084191f
C1149 commonsourceibias.n36 gnd 0.04027f
C1150 commonsourceibias.n37 gnd 0.009461f
C1151 commonsourceibias.n38 gnd 0.00769f
C1152 commonsourceibias.n39 gnd 0.013037f
C1153 commonsourceibias.n40 gnd 0.070526f
C1154 commonsourceibias.n41 gnd 0.013093f
C1155 commonsourceibias.n42 gnd 0.009461f
C1156 commonsourceibias.n43 gnd 0.009461f
C1157 commonsourceibias.n44 gnd 0.009461f
C1158 commonsourceibias.n45 gnd 0.009597f
C1159 commonsourceibias.n46 gnd 0.070526f
C1160 commonsourceibias.n47 gnd 0.011661f
C1161 commonsourceibias.n48 gnd 0.0129f
C1162 commonsourceibias.n49 gnd 0.009461f
C1163 commonsourceibias.n50 gnd 0.009461f
C1164 commonsourceibias.n51 gnd 0.012816f
C1165 commonsourceibias.n52 gnd 0.007653f
C1166 commonsourceibias.n53 gnd 0.012975f
C1167 commonsourceibias.n54 gnd 0.009461f
C1168 commonsourceibias.n55 gnd 0.009461f
C1169 commonsourceibias.n56 gnd 0.013054f
C1170 commonsourceibias.n57 gnd 0.011256f
C1171 commonsourceibias.n58 gnd 0.009134f
C1172 commonsourceibias.n59 gnd 0.009461f
C1173 commonsourceibias.n60 gnd 0.009461f
C1174 commonsourceibias.n61 gnd 0.011572f
C1175 commonsourceibias.n62 gnd 0.012989f
C1176 commonsourceibias.n63 gnd 0.070526f
C1177 commonsourceibias.n64 gnd 0.012901f
C1178 commonsourceibias.n65 gnd 0.009461f
C1179 commonsourceibias.n66 gnd 0.009461f
C1180 commonsourceibias.n67 gnd 0.009461f
C1181 commonsourceibias.n68 gnd 0.012901f
C1182 commonsourceibias.n69 gnd 0.070526f
C1183 commonsourceibias.n70 gnd 0.012989f
C1184 commonsourceibias.n71 gnd 0.011572f
C1185 commonsourceibias.n72 gnd 0.009461f
C1186 commonsourceibias.n73 gnd 0.009461f
C1187 commonsourceibias.n74 gnd 0.009461f
C1188 commonsourceibias.n75 gnd 0.011256f
C1189 commonsourceibias.n76 gnd 0.013054f
C1190 commonsourceibias.n77 gnd 0.070526f
C1191 commonsourceibias.n78 gnd 0.012975f
C1192 commonsourceibias.n79 gnd 0.009461f
C1193 commonsourceibias.n80 gnd 0.009461f
C1194 commonsourceibias.n81 gnd 0.009461f
C1195 commonsourceibias.n82 gnd 0.012816f
C1196 commonsourceibias.n83 gnd 0.070526f
C1197 commonsourceibias.n84 gnd 0.0129f
C1198 commonsourceibias.n85 gnd 0.011661f
C1199 commonsourceibias.n86 gnd 0.009461f
C1200 commonsourceibias.n87 gnd 0.009461f
C1201 commonsourceibias.n88 gnd 0.009461f
C1202 commonsourceibias.n89 gnd 0.010754f
C1203 commonsourceibias.n90 gnd 0.013093f
C1204 commonsourceibias.n91 gnd 0.070526f
C1205 commonsourceibias.n92 gnd 0.013037f
C1206 commonsourceibias.n93 gnd 0.009461f
C1207 commonsourceibias.n94 gnd 0.009461f
C1208 commonsourceibias.n95 gnd 0.009461f
C1209 commonsourceibias.n96 gnd 0.012717f
C1210 commonsourceibias.n97 gnd 0.070526f
C1211 commonsourceibias.n98 gnd 0.012748f
C1212 commonsourceibias.n99 gnd 0.085044f
C1213 commonsourceibias.n100 gnd 0.095092f
C1214 commonsourceibias.t13 gnd 0.020415f
C1215 commonsourceibias.t49 gnd 0.020415f
C1216 commonsourceibias.n101 gnd 0.180398f
C1217 commonsourceibias.n102 gnd 0.156264f
C1218 commonsourceibias.t5 gnd 0.020415f
C1219 commonsourceibias.t11 gnd 0.020415f
C1220 commonsourceibias.n103 gnd 0.180398f
C1221 commonsourceibias.n104 gnd 0.082864f
C1222 commonsourceibias.t59 gnd 0.020415f
C1223 commonsourceibias.t17 gnd 0.020415f
C1224 commonsourceibias.n105 gnd 0.180398f
C1225 commonsourceibias.n106 gnd 0.082864f
C1226 commonsourceibias.t29 gnd 0.020415f
C1227 commonsourceibias.t7 gnd 0.020415f
C1228 commonsourceibias.n107 gnd 0.180398f
C1229 commonsourceibias.n108 gnd 0.069229f
C1230 commonsourceibias.t51 gnd 0.020415f
C1231 commonsourceibias.t1 gnd 0.020415f
C1232 commonsourceibias.n109 gnd 0.181002f
C1233 commonsourceibias.t55 gnd 0.020415f
C1234 commonsourceibias.t19 gnd 0.020415f
C1235 commonsourceibias.n110 gnd 0.180398f
C1236 commonsourceibias.n111 gnd 0.168097f
C1237 commonsourceibias.t25 gnd 0.020415f
C1238 commonsourceibias.t31 gnd 0.020415f
C1239 commonsourceibias.n112 gnd 0.180398f
C1240 commonsourceibias.n113 gnd 0.082864f
C1241 commonsourceibias.t15 gnd 0.020415f
C1242 commonsourceibias.t45 gnd 0.020415f
C1243 commonsourceibias.n114 gnd 0.180398f
C1244 commonsourceibias.n115 gnd 0.069229f
C1245 commonsourceibias.n116 gnd 0.083829f
C1246 commonsourceibias.n117 gnd 0.009461f
C1247 commonsourceibias.t118 gnd 0.176757f
C1248 commonsourceibias.t76 gnd 0.176757f
C1249 commonsourceibias.n118 gnd 0.070526f
C1250 commonsourceibias.n119 gnd 0.009461f
C1251 commonsourceibias.t106 gnd 0.176757f
C1252 commonsourceibias.n120 gnd 0.070526f
C1253 commonsourceibias.n121 gnd 0.009461f
C1254 commonsourceibias.t96 gnd 0.176757f
C1255 commonsourceibias.n122 gnd 0.070526f
C1256 commonsourceibias.n123 gnd 0.009461f
C1257 commonsourceibias.t141 gnd 0.176757f
C1258 commonsourceibias.n124 gnd 0.010754f
C1259 commonsourceibias.n125 gnd 0.009461f
C1260 commonsourceibias.t116 gnd 0.176757f
C1261 commonsourceibias.n126 gnd 0.012717f
C1262 commonsourceibias.t129 gnd 0.196904f
C1263 commonsourceibias.t152 gnd 0.176757f
C1264 commonsourceibias.n127 gnd 0.078584f
C1265 commonsourceibias.n128 gnd 0.084191f
C1266 commonsourceibias.n129 gnd 0.04027f
C1267 commonsourceibias.n130 gnd 0.009461f
C1268 commonsourceibias.n131 gnd 0.00769f
C1269 commonsourceibias.n132 gnd 0.013037f
C1270 commonsourceibias.n133 gnd 0.070526f
C1271 commonsourceibias.n134 gnd 0.013093f
C1272 commonsourceibias.n135 gnd 0.009461f
C1273 commonsourceibias.n136 gnd 0.009461f
C1274 commonsourceibias.n137 gnd 0.009461f
C1275 commonsourceibias.n138 gnd 0.009597f
C1276 commonsourceibias.n139 gnd 0.070526f
C1277 commonsourceibias.n140 gnd 0.011661f
C1278 commonsourceibias.n141 gnd 0.0129f
C1279 commonsourceibias.n142 gnd 0.009461f
C1280 commonsourceibias.n143 gnd 0.009461f
C1281 commonsourceibias.n144 gnd 0.012816f
C1282 commonsourceibias.n145 gnd 0.007653f
C1283 commonsourceibias.n146 gnd 0.012975f
C1284 commonsourceibias.n147 gnd 0.009461f
C1285 commonsourceibias.n148 gnd 0.009461f
C1286 commonsourceibias.n149 gnd 0.013054f
C1287 commonsourceibias.n150 gnd 0.011256f
C1288 commonsourceibias.n151 gnd 0.009134f
C1289 commonsourceibias.n152 gnd 0.009461f
C1290 commonsourceibias.n153 gnd 0.009461f
C1291 commonsourceibias.n154 gnd 0.011572f
C1292 commonsourceibias.n155 gnd 0.012989f
C1293 commonsourceibias.n156 gnd 0.070526f
C1294 commonsourceibias.n157 gnd 0.012901f
C1295 commonsourceibias.n158 gnd 0.009415f
C1296 commonsourceibias.n159 gnd 0.06839f
C1297 commonsourceibias.n160 gnd 0.009415f
C1298 commonsourceibias.n161 gnd 0.012901f
C1299 commonsourceibias.n162 gnd 0.070526f
C1300 commonsourceibias.n163 gnd 0.012989f
C1301 commonsourceibias.n164 gnd 0.011572f
C1302 commonsourceibias.n165 gnd 0.009461f
C1303 commonsourceibias.n166 gnd 0.009461f
C1304 commonsourceibias.n167 gnd 0.009461f
C1305 commonsourceibias.n168 gnd 0.011256f
C1306 commonsourceibias.n169 gnd 0.013054f
C1307 commonsourceibias.n170 gnd 0.070526f
C1308 commonsourceibias.n171 gnd 0.012975f
C1309 commonsourceibias.n172 gnd 0.009461f
C1310 commonsourceibias.n173 gnd 0.009461f
C1311 commonsourceibias.n174 gnd 0.009461f
C1312 commonsourceibias.n175 gnd 0.012816f
C1313 commonsourceibias.n176 gnd 0.070526f
C1314 commonsourceibias.n177 gnd 0.0129f
C1315 commonsourceibias.n178 gnd 0.011661f
C1316 commonsourceibias.n179 gnd 0.009461f
C1317 commonsourceibias.n180 gnd 0.009461f
C1318 commonsourceibias.n181 gnd 0.009461f
C1319 commonsourceibias.n182 gnd 0.010754f
C1320 commonsourceibias.n183 gnd 0.013093f
C1321 commonsourceibias.n184 gnd 0.070526f
C1322 commonsourceibias.n185 gnd 0.013037f
C1323 commonsourceibias.n186 gnd 0.009461f
C1324 commonsourceibias.n187 gnd 0.009461f
C1325 commonsourceibias.n188 gnd 0.009461f
C1326 commonsourceibias.n189 gnd 0.012717f
C1327 commonsourceibias.n190 gnd 0.070526f
C1328 commonsourceibias.n191 gnd 0.012748f
C1329 commonsourceibias.n192 gnd 0.085044f
C1330 commonsourceibias.n193 gnd 0.056182f
C1331 commonsourceibias.n194 gnd 0.012624f
C1332 commonsourceibias.t71 gnd 0.191163f
C1333 commonsourceibias.t159 gnd 0.176757f
C1334 commonsourceibias.n195 gnd 0.00769f
C1335 commonsourceibias.n196 gnd 0.009461f
C1336 commonsourceibias.t148 gnd 0.176757f
C1337 commonsourceibias.n197 gnd 0.009597f
C1338 commonsourceibias.n198 gnd 0.009461f
C1339 commonsourceibias.t78 gnd 0.176757f
C1340 commonsourceibias.n199 gnd 0.070526f
C1341 commonsourceibias.t157 gnd 0.176757f
C1342 commonsourceibias.n200 gnd 0.007653f
C1343 commonsourceibias.n201 gnd 0.009461f
C1344 commonsourceibias.t85 gnd 0.176757f
C1345 commonsourceibias.n202 gnd 0.009134f
C1346 commonsourceibias.n203 gnd 0.009461f
C1347 commonsourceibias.t77 gnd 0.176757f
C1348 commonsourceibias.n204 gnd 0.070526f
C1349 commonsourceibias.t158 gnd 0.176757f
C1350 commonsourceibias.n205 gnd 0.007641f
C1351 commonsourceibias.n206 gnd 0.009461f
C1352 commonsourceibias.t94 gnd 0.176757f
C1353 commonsourceibias.t113 gnd 0.176757f
C1354 commonsourceibias.n207 gnd 0.070526f
C1355 commonsourceibias.n208 gnd 0.009461f
C1356 commonsourceibias.t156 gnd 0.176757f
C1357 commonsourceibias.n209 gnd 0.070526f
C1358 commonsourceibias.n210 gnd 0.009461f
C1359 commonsourceibias.t92 gnd 0.176757f
C1360 commonsourceibias.n211 gnd 0.070526f
C1361 commonsourceibias.n212 gnd 0.009461f
C1362 commonsourceibias.t111 gnd 0.176757f
C1363 commonsourceibias.n213 gnd 0.010754f
C1364 commonsourceibias.n214 gnd 0.009461f
C1365 commonsourceibias.t105 gnd 0.176757f
C1366 commonsourceibias.n215 gnd 0.012717f
C1367 commonsourceibias.t112 gnd 0.196904f
C1368 commonsourceibias.t93 gnd 0.176757f
C1369 commonsourceibias.n216 gnd 0.078584f
C1370 commonsourceibias.n217 gnd 0.084191f
C1371 commonsourceibias.n218 gnd 0.04027f
C1372 commonsourceibias.n219 gnd 0.009461f
C1373 commonsourceibias.n220 gnd 0.00769f
C1374 commonsourceibias.n221 gnd 0.013037f
C1375 commonsourceibias.n222 gnd 0.070526f
C1376 commonsourceibias.n223 gnd 0.013093f
C1377 commonsourceibias.n224 gnd 0.009461f
C1378 commonsourceibias.n225 gnd 0.009461f
C1379 commonsourceibias.n226 gnd 0.009461f
C1380 commonsourceibias.n227 gnd 0.009597f
C1381 commonsourceibias.n228 gnd 0.070526f
C1382 commonsourceibias.n229 gnd 0.011661f
C1383 commonsourceibias.n230 gnd 0.0129f
C1384 commonsourceibias.n231 gnd 0.009461f
C1385 commonsourceibias.n232 gnd 0.009461f
C1386 commonsourceibias.n233 gnd 0.012816f
C1387 commonsourceibias.n234 gnd 0.007653f
C1388 commonsourceibias.n235 gnd 0.012975f
C1389 commonsourceibias.n236 gnd 0.009461f
C1390 commonsourceibias.n237 gnd 0.009461f
C1391 commonsourceibias.n238 gnd 0.013054f
C1392 commonsourceibias.n239 gnd 0.011256f
C1393 commonsourceibias.n240 gnd 0.009134f
C1394 commonsourceibias.n241 gnd 0.009461f
C1395 commonsourceibias.n242 gnd 0.009461f
C1396 commonsourceibias.n243 gnd 0.011572f
C1397 commonsourceibias.n244 gnd 0.012989f
C1398 commonsourceibias.n245 gnd 0.070526f
C1399 commonsourceibias.n246 gnd 0.012901f
C1400 commonsourceibias.n247 gnd 0.009461f
C1401 commonsourceibias.n248 gnd 0.009461f
C1402 commonsourceibias.n249 gnd 0.009461f
C1403 commonsourceibias.n250 gnd 0.012901f
C1404 commonsourceibias.n251 gnd 0.070526f
C1405 commonsourceibias.n252 gnd 0.012989f
C1406 commonsourceibias.n253 gnd 0.011572f
C1407 commonsourceibias.n254 gnd 0.009461f
C1408 commonsourceibias.n255 gnd 0.009461f
C1409 commonsourceibias.n256 gnd 0.009461f
C1410 commonsourceibias.n257 gnd 0.011256f
C1411 commonsourceibias.n258 gnd 0.013054f
C1412 commonsourceibias.n259 gnd 0.070526f
C1413 commonsourceibias.n260 gnd 0.012975f
C1414 commonsourceibias.n261 gnd 0.009461f
C1415 commonsourceibias.n262 gnd 0.009461f
C1416 commonsourceibias.n263 gnd 0.009461f
C1417 commonsourceibias.n264 gnd 0.012816f
C1418 commonsourceibias.n265 gnd 0.070526f
C1419 commonsourceibias.n266 gnd 0.0129f
C1420 commonsourceibias.n267 gnd 0.011661f
C1421 commonsourceibias.n268 gnd 0.009461f
C1422 commonsourceibias.n269 gnd 0.009461f
C1423 commonsourceibias.n270 gnd 0.009461f
C1424 commonsourceibias.n271 gnd 0.010754f
C1425 commonsourceibias.n272 gnd 0.013093f
C1426 commonsourceibias.n273 gnd 0.070526f
C1427 commonsourceibias.n274 gnd 0.013037f
C1428 commonsourceibias.n275 gnd 0.009461f
C1429 commonsourceibias.n276 gnd 0.009461f
C1430 commonsourceibias.n277 gnd 0.009461f
C1431 commonsourceibias.n278 gnd 0.012717f
C1432 commonsourceibias.n279 gnd 0.070526f
C1433 commonsourceibias.n280 gnd 0.012748f
C1434 commonsourceibias.n281 gnd 0.085044f
C1435 commonsourceibias.n282 gnd 0.030348f
C1436 commonsourceibias.n283 gnd 0.15151f
C1437 commonsourceibias.n284 gnd 0.012624f
C1438 commonsourceibias.t75 gnd 0.176757f
C1439 commonsourceibias.n285 gnd 0.00769f
C1440 commonsourceibias.n286 gnd 0.009461f
C1441 commonsourceibias.t128 gnd 0.176757f
C1442 commonsourceibias.n287 gnd 0.009597f
C1443 commonsourceibias.n288 gnd 0.009461f
C1444 commonsourceibias.t124 gnd 0.176757f
C1445 commonsourceibias.n289 gnd 0.070526f
C1446 commonsourceibias.t155 gnd 0.176757f
C1447 commonsourceibias.n290 gnd 0.007653f
C1448 commonsourceibias.n291 gnd 0.009461f
C1449 commonsourceibias.t90 gnd 0.176757f
C1450 commonsourceibias.n292 gnd 0.009134f
C1451 commonsourceibias.n293 gnd 0.009461f
C1452 commonsourceibias.t119 gnd 0.176757f
C1453 commonsourceibias.n294 gnd 0.070526f
C1454 commonsourceibias.t146 gnd 0.176757f
C1455 commonsourceibias.n295 gnd 0.007641f
C1456 commonsourceibias.n296 gnd 0.009461f
C1457 commonsourceibias.t138 gnd 0.176757f
C1458 commonsourceibias.t64 gnd 0.176757f
C1459 commonsourceibias.n297 gnd 0.070526f
C1460 commonsourceibias.n298 gnd 0.009461f
C1461 commonsourceibias.t137 gnd 0.176757f
C1462 commonsourceibias.n299 gnd 0.070526f
C1463 commonsourceibias.n300 gnd 0.009461f
C1464 commonsourceibias.t133 gnd 0.176757f
C1465 commonsourceibias.n301 gnd 0.070526f
C1466 commonsourceibias.n302 gnd 0.009461f
C1467 commonsourceibias.t149 gnd 0.176757f
C1468 commonsourceibias.n303 gnd 0.010754f
C1469 commonsourceibias.n304 gnd 0.009461f
C1470 commonsourceibias.t79 gnd 0.176757f
C1471 commonsourceibias.n305 gnd 0.012717f
C1472 commonsourceibias.t140 gnd 0.196904f
C1473 commonsourceibias.t130 gnd 0.176757f
C1474 commonsourceibias.n306 gnd 0.078584f
C1475 commonsourceibias.n307 gnd 0.084191f
C1476 commonsourceibias.n308 gnd 0.04027f
C1477 commonsourceibias.n309 gnd 0.009461f
C1478 commonsourceibias.n310 gnd 0.00769f
C1479 commonsourceibias.n311 gnd 0.013037f
C1480 commonsourceibias.n312 gnd 0.070526f
C1481 commonsourceibias.n313 gnd 0.013093f
C1482 commonsourceibias.n314 gnd 0.009461f
C1483 commonsourceibias.n315 gnd 0.009461f
C1484 commonsourceibias.n316 gnd 0.009461f
C1485 commonsourceibias.n317 gnd 0.009597f
C1486 commonsourceibias.n318 gnd 0.070526f
C1487 commonsourceibias.n319 gnd 0.011661f
C1488 commonsourceibias.n320 gnd 0.0129f
C1489 commonsourceibias.n321 gnd 0.009461f
C1490 commonsourceibias.n322 gnd 0.009461f
C1491 commonsourceibias.n323 gnd 0.012816f
C1492 commonsourceibias.n324 gnd 0.007653f
C1493 commonsourceibias.n325 gnd 0.012975f
C1494 commonsourceibias.n326 gnd 0.009461f
C1495 commonsourceibias.n327 gnd 0.009461f
C1496 commonsourceibias.n328 gnd 0.013054f
C1497 commonsourceibias.n329 gnd 0.011256f
C1498 commonsourceibias.n330 gnd 0.009134f
C1499 commonsourceibias.n331 gnd 0.009461f
C1500 commonsourceibias.n332 gnd 0.009461f
C1501 commonsourceibias.n333 gnd 0.011572f
C1502 commonsourceibias.n334 gnd 0.012989f
C1503 commonsourceibias.n335 gnd 0.070526f
C1504 commonsourceibias.n336 gnd 0.012901f
C1505 commonsourceibias.n337 gnd 0.009461f
C1506 commonsourceibias.n338 gnd 0.009461f
C1507 commonsourceibias.n339 gnd 0.009461f
C1508 commonsourceibias.n340 gnd 0.012901f
C1509 commonsourceibias.n341 gnd 0.070526f
C1510 commonsourceibias.n342 gnd 0.012989f
C1511 commonsourceibias.n343 gnd 0.011572f
C1512 commonsourceibias.n344 gnd 0.009461f
C1513 commonsourceibias.n345 gnd 0.009461f
C1514 commonsourceibias.n346 gnd 0.009461f
C1515 commonsourceibias.n347 gnd 0.011256f
C1516 commonsourceibias.n348 gnd 0.013054f
C1517 commonsourceibias.n349 gnd 0.070526f
C1518 commonsourceibias.n350 gnd 0.012975f
C1519 commonsourceibias.n351 gnd 0.009461f
C1520 commonsourceibias.n352 gnd 0.009461f
C1521 commonsourceibias.n353 gnd 0.009461f
C1522 commonsourceibias.n354 gnd 0.012816f
C1523 commonsourceibias.n355 gnd 0.070526f
C1524 commonsourceibias.n356 gnd 0.0129f
C1525 commonsourceibias.n357 gnd 0.011661f
C1526 commonsourceibias.n358 gnd 0.009461f
C1527 commonsourceibias.n359 gnd 0.009461f
C1528 commonsourceibias.n360 gnd 0.009461f
C1529 commonsourceibias.n361 gnd 0.010754f
C1530 commonsourceibias.n362 gnd 0.013093f
C1531 commonsourceibias.n363 gnd 0.070526f
C1532 commonsourceibias.n364 gnd 0.013037f
C1533 commonsourceibias.n365 gnd 0.009461f
C1534 commonsourceibias.n366 gnd 0.009461f
C1535 commonsourceibias.n367 gnd 0.009461f
C1536 commonsourceibias.n368 gnd 0.012717f
C1537 commonsourceibias.n369 gnd 0.070526f
C1538 commonsourceibias.n370 gnd 0.012748f
C1539 commonsourceibias.t147 gnd 0.191163f
C1540 commonsourceibias.n371 gnd 0.085044f
C1541 commonsourceibias.n372 gnd 0.030348f
C1542 commonsourceibias.n373 gnd 0.449685f
C1543 commonsourceibias.n374 gnd 0.012624f
C1544 commonsourceibias.t91 gnd 0.191163f
C1545 commonsourceibias.t134 gnd 0.176757f
C1546 commonsourceibias.n375 gnd 0.00769f
C1547 commonsourceibias.n376 gnd 0.009461f
C1548 commonsourceibias.t114 gnd 0.176757f
C1549 commonsourceibias.n377 gnd 0.009597f
C1550 commonsourceibias.n378 gnd 0.009461f
C1551 commonsourceibias.t123 gnd 0.176757f
C1552 commonsourceibias.n379 gnd 0.007653f
C1553 commonsourceibias.n380 gnd 0.009461f
C1554 commonsourceibias.t88 gnd 0.176757f
C1555 commonsourceibias.n381 gnd 0.009134f
C1556 commonsourceibias.n382 gnd 0.009461f
C1557 commonsourceibias.t104 gnd 0.176757f
C1558 commonsourceibias.n383 gnd 0.007641f
C1559 commonsourceibias.n384 gnd 0.009461f
C1560 commonsourceibias.t89 gnd 0.176757f
C1561 commonsourceibias.t139 gnd 0.176757f
C1562 commonsourceibias.n385 gnd 0.070526f
C1563 commonsourceibias.n386 gnd 0.009461f
C1564 commonsourceibias.t83 gnd 0.176757f
C1565 commonsourceibias.n387 gnd 0.070526f
C1566 commonsourceibias.n388 gnd 0.009461f
C1567 commonsourceibias.t150 gnd 0.176757f
C1568 commonsourceibias.n389 gnd 0.070526f
C1569 commonsourceibias.n390 gnd 0.009461f
C1570 commonsourceibias.t127 gnd 0.176757f
C1571 commonsourceibias.n391 gnd 0.010754f
C1572 commonsourceibias.n392 gnd 0.009461f
C1573 commonsourceibias.t84 gnd 0.176757f
C1574 commonsourceibias.n393 gnd 0.012717f
C1575 commonsourceibias.t108 gnd 0.196904f
C1576 commonsourceibias.t131 gnd 0.176757f
C1577 commonsourceibias.n394 gnd 0.078584f
C1578 commonsourceibias.n395 gnd 0.084191f
C1579 commonsourceibias.n396 gnd 0.04027f
C1580 commonsourceibias.n397 gnd 0.009461f
C1581 commonsourceibias.n398 gnd 0.00769f
C1582 commonsourceibias.n399 gnd 0.013037f
C1583 commonsourceibias.n400 gnd 0.070526f
C1584 commonsourceibias.n401 gnd 0.013093f
C1585 commonsourceibias.n402 gnd 0.009461f
C1586 commonsourceibias.n403 gnd 0.009461f
C1587 commonsourceibias.n404 gnd 0.009461f
C1588 commonsourceibias.n405 gnd 0.009597f
C1589 commonsourceibias.n406 gnd 0.070526f
C1590 commonsourceibias.n407 gnd 0.011661f
C1591 commonsourceibias.n408 gnd 0.0129f
C1592 commonsourceibias.n409 gnd 0.009461f
C1593 commonsourceibias.n410 gnd 0.009461f
C1594 commonsourceibias.n411 gnd 0.012816f
C1595 commonsourceibias.n412 gnd 0.007653f
C1596 commonsourceibias.n413 gnd 0.012975f
C1597 commonsourceibias.n414 gnd 0.009461f
C1598 commonsourceibias.n415 gnd 0.009461f
C1599 commonsourceibias.n416 gnd 0.013054f
C1600 commonsourceibias.n417 gnd 0.011256f
C1601 commonsourceibias.n418 gnd 0.009134f
C1602 commonsourceibias.n419 gnd 0.009461f
C1603 commonsourceibias.n420 gnd 0.009461f
C1604 commonsourceibias.n421 gnd 0.011572f
C1605 commonsourceibias.n422 gnd 0.012989f
C1606 commonsourceibias.n423 gnd 0.070526f
C1607 commonsourceibias.n424 gnd 0.012901f
C1608 commonsourceibias.n425 gnd 0.009415f
C1609 commonsourceibias.t23 gnd 0.020415f
C1610 commonsourceibias.t63 gnd 0.020415f
C1611 commonsourceibias.n426 gnd 0.181002f
C1612 commonsourceibias.t41 gnd 0.020415f
C1613 commonsourceibias.t3 gnd 0.020415f
C1614 commonsourceibias.n427 gnd 0.180398f
C1615 commonsourceibias.n428 gnd 0.168097f
C1616 commonsourceibias.t53 gnd 0.020415f
C1617 commonsourceibias.t43 gnd 0.020415f
C1618 commonsourceibias.n429 gnd 0.180398f
C1619 commonsourceibias.n430 gnd 0.082864f
C1620 commonsourceibias.t57 gnd 0.020415f
C1621 commonsourceibias.t37 gnd 0.020415f
C1622 commonsourceibias.n431 gnd 0.180398f
C1623 commonsourceibias.n432 gnd 0.069229f
C1624 commonsourceibias.n433 gnd 0.012624f
C1625 commonsourceibias.t60 gnd 0.176757f
C1626 commonsourceibias.n434 gnd 0.00769f
C1627 commonsourceibias.n435 gnd 0.009461f
C1628 commonsourceibias.t20 gnd 0.176757f
C1629 commonsourceibias.n436 gnd 0.009597f
C1630 commonsourceibias.n437 gnd 0.009461f
C1631 commonsourceibias.t8 gnd 0.176757f
C1632 commonsourceibias.n438 gnd 0.007653f
C1633 commonsourceibias.n439 gnd 0.009461f
C1634 commonsourceibias.t38 gnd 0.176757f
C1635 commonsourceibias.n440 gnd 0.009134f
C1636 commonsourceibias.n441 gnd 0.009461f
C1637 commonsourceibias.t26 gnd 0.176757f
C1638 commonsourceibias.n442 gnd 0.007641f
C1639 commonsourceibias.n443 gnd 0.009461f
C1640 commonsourceibias.t36 gnd 0.176757f
C1641 commonsourceibias.t56 gnd 0.176757f
C1642 commonsourceibias.n444 gnd 0.070526f
C1643 commonsourceibias.n445 gnd 0.009461f
C1644 commonsourceibias.t42 gnd 0.176757f
C1645 commonsourceibias.n446 gnd 0.070526f
C1646 commonsourceibias.n447 gnd 0.009461f
C1647 commonsourceibias.t52 gnd 0.176757f
C1648 commonsourceibias.n448 gnd 0.070526f
C1649 commonsourceibias.n449 gnd 0.009461f
C1650 commonsourceibias.t2 gnd 0.176757f
C1651 commonsourceibias.n450 gnd 0.010754f
C1652 commonsourceibias.n451 gnd 0.009461f
C1653 commonsourceibias.t40 gnd 0.176757f
C1654 commonsourceibias.n452 gnd 0.012717f
C1655 commonsourceibias.t22 gnd 0.196904f
C1656 commonsourceibias.t62 gnd 0.176757f
C1657 commonsourceibias.n453 gnd 0.078584f
C1658 commonsourceibias.n454 gnd 0.084191f
C1659 commonsourceibias.n455 gnd 0.04027f
C1660 commonsourceibias.n456 gnd 0.009461f
C1661 commonsourceibias.n457 gnd 0.00769f
C1662 commonsourceibias.n458 gnd 0.013037f
C1663 commonsourceibias.n459 gnd 0.070526f
C1664 commonsourceibias.n460 gnd 0.013093f
C1665 commonsourceibias.n461 gnd 0.009461f
C1666 commonsourceibias.n462 gnd 0.009461f
C1667 commonsourceibias.n463 gnd 0.009461f
C1668 commonsourceibias.n464 gnd 0.009597f
C1669 commonsourceibias.n465 gnd 0.070526f
C1670 commonsourceibias.n466 gnd 0.011661f
C1671 commonsourceibias.n467 gnd 0.0129f
C1672 commonsourceibias.n468 gnd 0.009461f
C1673 commonsourceibias.n469 gnd 0.009461f
C1674 commonsourceibias.n470 gnd 0.012816f
C1675 commonsourceibias.n471 gnd 0.007653f
C1676 commonsourceibias.n472 gnd 0.012975f
C1677 commonsourceibias.n473 gnd 0.009461f
C1678 commonsourceibias.n474 gnd 0.009461f
C1679 commonsourceibias.n475 gnd 0.013054f
C1680 commonsourceibias.n476 gnd 0.011256f
C1681 commonsourceibias.n477 gnd 0.009134f
C1682 commonsourceibias.n478 gnd 0.009461f
C1683 commonsourceibias.n479 gnd 0.009461f
C1684 commonsourceibias.n480 gnd 0.011572f
C1685 commonsourceibias.n481 gnd 0.012989f
C1686 commonsourceibias.n482 gnd 0.070526f
C1687 commonsourceibias.n483 gnd 0.012901f
C1688 commonsourceibias.n484 gnd 0.009461f
C1689 commonsourceibias.n485 gnd 0.009461f
C1690 commonsourceibias.n486 gnd 0.009461f
C1691 commonsourceibias.n487 gnd 0.012901f
C1692 commonsourceibias.n488 gnd 0.070526f
C1693 commonsourceibias.n489 gnd 0.012989f
C1694 commonsourceibias.t46 gnd 0.176757f
C1695 commonsourceibias.n490 gnd 0.070526f
C1696 commonsourceibias.n491 gnd 0.011572f
C1697 commonsourceibias.n492 gnd 0.009461f
C1698 commonsourceibias.n493 gnd 0.009461f
C1699 commonsourceibias.n494 gnd 0.009461f
C1700 commonsourceibias.n495 gnd 0.011256f
C1701 commonsourceibias.n496 gnd 0.013054f
C1702 commonsourceibias.n497 gnd 0.070526f
C1703 commonsourceibias.n498 gnd 0.012975f
C1704 commonsourceibias.n499 gnd 0.009461f
C1705 commonsourceibias.n500 gnd 0.009461f
C1706 commonsourceibias.n501 gnd 0.009461f
C1707 commonsourceibias.n502 gnd 0.012816f
C1708 commonsourceibias.n503 gnd 0.070526f
C1709 commonsourceibias.n504 gnd 0.0129f
C1710 commonsourceibias.t32 gnd 0.176757f
C1711 commonsourceibias.n505 gnd 0.070526f
C1712 commonsourceibias.n506 gnd 0.011661f
C1713 commonsourceibias.n507 gnd 0.009461f
C1714 commonsourceibias.n508 gnd 0.009461f
C1715 commonsourceibias.n509 gnd 0.009461f
C1716 commonsourceibias.n510 gnd 0.010754f
C1717 commonsourceibias.n511 gnd 0.013093f
C1718 commonsourceibias.n512 gnd 0.070526f
C1719 commonsourceibias.n513 gnd 0.013037f
C1720 commonsourceibias.n514 gnd 0.009461f
C1721 commonsourceibias.n515 gnd 0.009461f
C1722 commonsourceibias.n516 gnd 0.009461f
C1723 commonsourceibias.n517 gnd 0.012717f
C1724 commonsourceibias.n518 gnd 0.070526f
C1725 commonsourceibias.n519 gnd 0.012748f
C1726 commonsourceibias.t34 gnd 0.191163f
C1727 commonsourceibias.n520 gnd 0.085044f
C1728 commonsourceibias.n521 gnd 0.095092f
C1729 commonsourceibias.t61 gnd 0.020415f
C1730 commonsourceibias.t35 gnd 0.020415f
C1731 commonsourceibias.n522 gnd 0.180398f
C1732 commonsourceibias.n523 gnd 0.156264f
C1733 commonsourceibias.t33 gnd 0.020415f
C1734 commonsourceibias.t21 gnd 0.020415f
C1735 commonsourceibias.n524 gnd 0.180398f
C1736 commonsourceibias.n525 gnd 0.082864f
C1737 commonsourceibias.t39 gnd 0.020415f
C1738 commonsourceibias.t9 gnd 0.020415f
C1739 commonsourceibias.n526 gnd 0.180398f
C1740 commonsourceibias.n527 gnd 0.082864f
C1741 commonsourceibias.t27 gnd 0.020415f
C1742 commonsourceibias.t47 gnd 0.020415f
C1743 commonsourceibias.n528 gnd 0.180398f
C1744 commonsourceibias.n529 gnd 0.069229f
C1745 commonsourceibias.n530 gnd 0.083829f
C1746 commonsourceibias.n531 gnd 0.06839f
C1747 commonsourceibias.n532 gnd 0.009415f
C1748 commonsourceibias.n533 gnd 0.012901f
C1749 commonsourceibias.n534 gnd 0.070526f
C1750 commonsourceibias.n535 gnd 0.012989f
C1751 commonsourceibias.t73 gnd 0.176757f
C1752 commonsourceibias.n536 gnd 0.070526f
C1753 commonsourceibias.n537 gnd 0.011572f
C1754 commonsourceibias.n538 gnd 0.009461f
C1755 commonsourceibias.n539 gnd 0.009461f
C1756 commonsourceibias.n540 gnd 0.009461f
C1757 commonsourceibias.n541 gnd 0.011256f
C1758 commonsourceibias.n542 gnd 0.013054f
C1759 commonsourceibias.n543 gnd 0.070526f
C1760 commonsourceibias.n544 gnd 0.012975f
C1761 commonsourceibias.n545 gnd 0.009461f
C1762 commonsourceibias.n546 gnd 0.009461f
C1763 commonsourceibias.n547 gnd 0.009461f
C1764 commonsourceibias.n548 gnd 0.012816f
C1765 commonsourceibias.n549 gnd 0.070526f
C1766 commonsourceibias.n550 gnd 0.0129f
C1767 commonsourceibias.t95 gnd 0.176757f
C1768 commonsourceibias.n551 gnd 0.070526f
C1769 commonsourceibias.n552 gnd 0.011661f
C1770 commonsourceibias.n553 gnd 0.009461f
C1771 commonsourceibias.n554 gnd 0.009461f
C1772 commonsourceibias.n555 gnd 0.009461f
C1773 commonsourceibias.n556 gnd 0.010754f
C1774 commonsourceibias.n557 gnd 0.013093f
C1775 commonsourceibias.n558 gnd 0.070526f
C1776 commonsourceibias.n559 gnd 0.013037f
C1777 commonsourceibias.n560 gnd 0.009461f
C1778 commonsourceibias.n561 gnd 0.009461f
C1779 commonsourceibias.n562 gnd 0.009461f
C1780 commonsourceibias.n563 gnd 0.012717f
C1781 commonsourceibias.n564 gnd 0.070526f
C1782 commonsourceibias.n565 gnd 0.012748f
C1783 commonsourceibias.n566 gnd 0.085044f
C1784 commonsourceibias.n567 gnd 0.056182f
C1785 commonsourceibias.n568 gnd 0.012624f
C1786 commonsourceibias.t144 gnd 0.176757f
C1787 commonsourceibias.n569 gnd 0.00769f
C1788 commonsourceibias.n570 gnd 0.009461f
C1789 commonsourceibias.t66 gnd 0.176757f
C1790 commonsourceibias.n571 gnd 0.009597f
C1791 commonsourceibias.n572 gnd 0.009461f
C1792 commonsourceibias.t143 gnd 0.176757f
C1793 commonsourceibias.n573 gnd 0.007653f
C1794 commonsourceibias.n574 gnd 0.009461f
C1795 commonsourceibias.t65 gnd 0.176757f
C1796 commonsourceibias.n575 gnd 0.009134f
C1797 commonsourceibias.n576 gnd 0.009461f
C1798 commonsourceibias.t142 gnd 0.176757f
C1799 commonsourceibias.n577 gnd 0.007641f
C1800 commonsourceibias.n578 gnd 0.009461f
C1801 commonsourceibias.t72 gnd 0.176757f
C1802 commonsourceibias.t99 gnd 0.176757f
C1803 commonsourceibias.n579 gnd 0.070526f
C1804 commonsourceibias.n580 gnd 0.009461f
C1805 commonsourceibias.t80 gnd 0.176757f
C1806 commonsourceibias.n581 gnd 0.070526f
C1807 commonsourceibias.n582 gnd 0.009461f
C1808 commonsourceibias.t69 gnd 0.176757f
C1809 commonsourceibias.n583 gnd 0.070526f
C1810 commonsourceibias.n584 gnd 0.009461f
C1811 commonsourceibias.t98 gnd 0.176757f
C1812 commonsourceibias.n585 gnd 0.010754f
C1813 commonsourceibias.n586 gnd 0.009461f
C1814 commonsourceibias.t86 gnd 0.176757f
C1815 commonsourceibias.n587 gnd 0.012717f
C1816 commonsourceibias.t97 gnd 0.196904f
C1817 commonsourceibias.t68 gnd 0.176757f
C1818 commonsourceibias.n588 gnd 0.078584f
C1819 commonsourceibias.n589 gnd 0.084191f
C1820 commonsourceibias.n590 gnd 0.04027f
C1821 commonsourceibias.n591 gnd 0.009461f
C1822 commonsourceibias.n592 gnd 0.00769f
C1823 commonsourceibias.n593 gnd 0.013037f
C1824 commonsourceibias.n594 gnd 0.070526f
C1825 commonsourceibias.n595 gnd 0.013093f
C1826 commonsourceibias.n596 gnd 0.009461f
C1827 commonsourceibias.n597 gnd 0.009461f
C1828 commonsourceibias.n598 gnd 0.009461f
C1829 commonsourceibias.n599 gnd 0.009597f
C1830 commonsourceibias.n600 gnd 0.070526f
C1831 commonsourceibias.n601 gnd 0.011661f
C1832 commonsourceibias.n602 gnd 0.0129f
C1833 commonsourceibias.n603 gnd 0.009461f
C1834 commonsourceibias.n604 gnd 0.009461f
C1835 commonsourceibias.n605 gnd 0.012816f
C1836 commonsourceibias.n606 gnd 0.007653f
C1837 commonsourceibias.n607 gnd 0.012975f
C1838 commonsourceibias.n608 gnd 0.009461f
C1839 commonsourceibias.n609 gnd 0.009461f
C1840 commonsourceibias.n610 gnd 0.013054f
C1841 commonsourceibias.n611 gnd 0.011256f
C1842 commonsourceibias.n612 gnd 0.009134f
C1843 commonsourceibias.n613 gnd 0.009461f
C1844 commonsourceibias.n614 gnd 0.009461f
C1845 commonsourceibias.n615 gnd 0.011572f
C1846 commonsourceibias.n616 gnd 0.012989f
C1847 commonsourceibias.n617 gnd 0.070526f
C1848 commonsourceibias.n618 gnd 0.012901f
C1849 commonsourceibias.n619 gnd 0.009461f
C1850 commonsourceibias.n620 gnd 0.009461f
C1851 commonsourceibias.n621 gnd 0.009461f
C1852 commonsourceibias.n622 gnd 0.012901f
C1853 commonsourceibias.n623 gnd 0.070526f
C1854 commonsourceibias.n624 gnd 0.012989f
C1855 commonsourceibias.t100 gnd 0.176757f
C1856 commonsourceibias.n625 gnd 0.070526f
C1857 commonsourceibias.n626 gnd 0.011572f
C1858 commonsourceibias.n627 gnd 0.009461f
C1859 commonsourceibias.n628 gnd 0.009461f
C1860 commonsourceibias.n629 gnd 0.009461f
C1861 commonsourceibias.n630 gnd 0.011256f
C1862 commonsourceibias.n631 gnd 0.013054f
C1863 commonsourceibias.n632 gnd 0.070526f
C1864 commonsourceibias.n633 gnd 0.012975f
C1865 commonsourceibias.n634 gnd 0.009461f
C1866 commonsourceibias.n635 gnd 0.009461f
C1867 commonsourceibias.n636 gnd 0.009461f
C1868 commonsourceibias.n637 gnd 0.012816f
C1869 commonsourceibias.n638 gnd 0.070526f
C1870 commonsourceibias.n639 gnd 0.0129f
C1871 commonsourceibias.t154 gnd 0.176757f
C1872 commonsourceibias.n640 gnd 0.070526f
C1873 commonsourceibias.n641 gnd 0.011661f
C1874 commonsourceibias.n642 gnd 0.009461f
C1875 commonsourceibias.n643 gnd 0.009461f
C1876 commonsourceibias.n644 gnd 0.009461f
C1877 commonsourceibias.n645 gnd 0.010754f
C1878 commonsourceibias.n646 gnd 0.013093f
C1879 commonsourceibias.n647 gnd 0.070526f
C1880 commonsourceibias.n648 gnd 0.013037f
C1881 commonsourceibias.n649 gnd 0.009461f
C1882 commonsourceibias.n650 gnd 0.009461f
C1883 commonsourceibias.n651 gnd 0.009461f
C1884 commonsourceibias.n652 gnd 0.012717f
C1885 commonsourceibias.n653 gnd 0.070526f
C1886 commonsourceibias.n654 gnd 0.012748f
C1887 commonsourceibias.t151 gnd 0.191163f
C1888 commonsourceibias.n655 gnd 0.085044f
C1889 commonsourceibias.n656 gnd 0.030348f
C1890 commonsourceibias.n657 gnd 0.15151f
C1891 commonsourceibias.n658 gnd 0.012624f
C1892 commonsourceibias.t107 gnd 0.176757f
C1893 commonsourceibias.n659 gnd 0.00769f
C1894 commonsourceibias.n660 gnd 0.009461f
C1895 commonsourceibias.t122 gnd 0.176757f
C1896 commonsourceibias.n661 gnd 0.009597f
C1897 commonsourceibias.n662 gnd 0.009461f
C1898 commonsourceibias.t101 gnd 0.176757f
C1899 commonsourceibias.n663 gnd 0.007653f
C1900 commonsourceibias.n664 gnd 0.009461f
C1901 commonsourceibias.t115 gnd 0.176757f
C1902 commonsourceibias.n665 gnd 0.009134f
C1903 commonsourceibias.n666 gnd 0.009461f
C1904 commonsourceibias.t81 gnd 0.176757f
C1905 commonsourceibias.n667 gnd 0.007641f
C1906 commonsourceibias.n668 gnd 0.009461f
C1907 commonsourceibias.t70 gnd 0.176757f
C1908 commonsourceibias.t103 gnd 0.176757f
C1909 commonsourceibias.n669 gnd 0.070526f
C1910 commonsourceibias.n670 gnd 0.009461f
C1911 commonsourceibias.t132 gnd 0.176757f
C1912 commonsourceibias.n671 gnd 0.070526f
C1913 commonsourceibias.n672 gnd 0.009461f
C1914 commonsourceibias.t153 gnd 0.176757f
C1915 commonsourceibias.n673 gnd 0.070526f
C1916 commonsourceibias.n674 gnd 0.009461f
C1917 commonsourceibias.t87 gnd 0.176757f
C1918 commonsourceibias.n675 gnd 0.010754f
C1919 commonsourceibias.n676 gnd 0.009461f
C1920 commonsourceibias.t109 gnd 0.176757f
C1921 commonsourceibias.n677 gnd 0.012717f
C1922 commonsourceibias.t74 gnd 0.196904f
C1923 commonsourceibias.t145 gnd 0.176757f
C1924 commonsourceibias.n678 gnd 0.078584f
C1925 commonsourceibias.n679 gnd 0.084191f
C1926 commonsourceibias.n680 gnd 0.04027f
C1927 commonsourceibias.n681 gnd 0.009461f
C1928 commonsourceibias.n682 gnd 0.00769f
C1929 commonsourceibias.n683 gnd 0.013037f
C1930 commonsourceibias.n684 gnd 0.070526f
C1931 commonsourceibias.n685 gnd 0.013093f
C1932 commonsourceibias.n686 gnd 0.009461f
C1933 commonsourceibias.n687 gnd 0.009461f
C1934 commonsourceibias.n688 gnd 0.009461f
C1935 commonsourceibias.n689 gnd 0.009597f
C1936 commonsourceibias.n690 gnd 0.070526f
C1937 commonsourceibias.n691 gnd 0.011661f
C1938 commonsourceibias.n692 gnd 0.0129f
C1939 commonsourceibias.n693 gnd 0.009461f
C1940 commonsourceibias.n694 gnd 0.009461f
C1941 commonsourceibias.n695 gnd 0.012816f
C1942 commonsourceibias.n696 gnd 0.007653f
C1943 commonsourceibias.n697 gnd 0.012975f
C1944 commonsourceibias.n698 gnd 0.009461f
C1945 commonsourceibias.n699 gnd 0.009461f
C1946 commonsourceibias.n700 gnd 0.013054f
C1947 commonsourceibias.n701 gnd 0.011256f
C1948 commonsourceibias.n702 gnd 0.009134f
C1949 commonsourceibias.n703 gnd 0.009461f
C1950 commonsourceibias.n704 gnd 0.009461f
C1951 commonsourceibias.n705 gnd 0.011572f
C1952 commonsourceibias.n706 gnd 0.012989f
C1953 commonsourceibias.n707 gnd 0.070526f
C1954 commonsourceibias.n708 gnd 0.012901f
C1955 commonsourceibias.n709 gnd 0.009461f
C1956 commonsourceibias.n710 gnd 0.009461f
C1957 commonsourceibias.n711 gnd 0.009461f
C1958 commonsourceibias.n712 gnd 0.012901f
C1959 commonsourceibias.n713 gnd 0.070526f
C1960 commonsourceibias.n714 gnd 0.012989f
C1961 commonsourceibias.t110 gnd 0.176757f
C1962 commonsourceibias.n715 gnd 0.070526f
C1963 commonsourceibias.n716 gnd 0.011572f
C1964 commonsourceibias.n717 gnd 0.009461f
C1965 commonsourceibias.n718 gnd 0.009461f
C1966 commonsourceibias.n719 gnd 0.009461f
C1967 commonsourceibias.n720 gnd 0.011256f
C1968 commonsourceibias.n721 gnd 0.013054f
C1969 commonsourceibias.n722 gnd 0.070526f
C1970 commonsourceibias.n723 gnd 0.012975f
C1971 commonsourceibias.n724 gnd 0.009461f
C1972 commonsourceibias.n725 gnd 0.009461f
C1973 commonsourceibias.n726 gnd 0.009461f
C1974 commonsourceibias.n727 gnd 0.012816f
C1975 commonsourceibias.n728 gnd 0.070526f
C1976 commonsourceibias.n729 gnd 0.0129f
C1977 commonsourceibias.t135 gnd 0.176757f
C1978 commonsourceibias.n730 gnd 0.070526f
C1979 commonsourceibias.n731 gnd 0.011661f
C1980 commonsourceibias.n732 gnd 0.009461f
C1981 commonsourceibias.n733 gnd 0.009461f
C1982 commonsourceibias.n734 gnd 0.009461f
C1983 commonsourceibias.n735 gnd 0.010754f
C1984 commonsourceibias.n736 gnd 0.013093f
C1985 commonsourceibias.n737 gnd 0.070526f
C1986 commonsourceibias.n738 gnd 0.013037f
C1987 commonsourceibias.n739 gnd 0.009461f
C1988 commonsourceibias.n740 gnd 0.009461f
C1989 commonsourceibias.n741 gnd 0.009461f
C1990 commonsourceibias.n742 gnd 0.012717f
C1991 commonsourceibias.n743 gnd 0.070526f
C1992 commonsourceibias.n744 gnd 0.012748f
C1993 commonsourceibias.t82 gnd 0.191163f
C1994 commonsourceibias.n745 gnd 0.085044f
C1995 commonsourceibias.n746 gnd 0.030348f
C1996 commonsourceibias.n747 gnd 0.199656f
C1997 commonsourceibias.n748 gnd 5.01419f
C1998 vdd.t45 gnd 0.032405f
C1999 vdd.t25 gnd 0.032405f
C2000 vdd.n0 gnd 0.255579f
C2001 vdd.t4 gnd 0.032405f
C2002 vdd.t41 gnd 0.032405f
C2003 vdd.n1 gnd 0.255158f
C2004 vdd.n2 gnd 0.235304f
C2005 vdd.t22 gnd 0.032405f
C2006 vdd.t52 gnd 0.032405f
C2007 vdd.n3 gnd 0.255158f
C2008 vdd.n4 gnd 0.119002f
C2009 vdd.t50 gnd 0.032405f
C2010 vdd.t30 gnd 0.032405f
C2011 vdd.n5 gnd 0.255158f
C2012 vdd.n6 gnd 0.111661f
C2013 vdd.t56 gnd 0.032405f
C2014 vdd.t20 gnd 0.032405f
C2015 vdd.n7 gnd 0.255579f
C2016 vdd.t28 gnd 0.032405f
C2017 vdd.t48 gnd 0.032405f
C2018 vdd.n8 gnd 0.255158f
C2019 vdd.n9 gnd 0.235304f
C2020 vdd.t37 gnd 0.032405f
C2021 vdd.t8 gnd 0.032405f
C2022 vdd.n10 gnd 0.255158f
C2023 vdd.n11 gnd 0.119002f
C2024 vdd.t17 gnd 0.032405f
C2025 vdd.t35 gnd 0.032405f
C2026 vdd.n12 gnd 0.255158f
C2027 vdd.n13 gnd 0.111661f
C2028 vdd.n14 gnd 0.078943f
C2029 vdd.t156 gnd 0.018003f
C2030 vdd.t237 gnd 0.018003f
C2031 vdd.n15 gnd 0.165705f
C2032 vdd.t57 gnd 0.018003f
C2033 vdd.t58 gnd 0.018003f
C2034 vdd.n16 gnd 0.165221f
C2035 vdd.n17 gnd 0.287535f
C2036 vdd.t159 gnd 0.018003f
C2037 vdd.t238 gnd 0.018003f
C2038 vdd.n18 gnd 0.165221f
C2039 vdd.n19 gnd 0.118957f
C2040 vdd.t241 gnd 0.018003f
C2041 vdd.t59 gnd 0.018003f
C2042 vdd.n20 gnd 0.165705f
C2043 vdd.t157 gnd 0.018003f
C2044 vdd.t242 gnd 0.018003f
C2045 vdd.n21 gnd 0.165221f
C2046 vdd.n22 gnd 0.287535f
C2047 vdd.t239 gnd 0.018003f
C2048 vdd.t240 gnd 0.018003f
C2049 vdd.n23 gnd 0.165221f
C2050 vdd.n24 gnd 0.118957f
C2051 vdd.t243 gnd 0.018003f
C2052 vdd.t0 gnd 0.018003f
C2053 vdd.n25 gnd 0.165221f
C2054 vdd.t236 gnd 0.018003f
C2055 vdd.t158 gnd 0.018003f
C2056 vdd.n26 gnd 0.165221f
C2057 vdd.n27 gnd 18.1145f
C2058 vdd.n28 gnd 7.14758f
C2059 vdd.n29 gnd 0.00491f
C2060 vdd.n30 gnd 0.004556f
C2061 vdd.n31 gnd 0.00252f
C2062 vdd.n32 gnd 0.005787f
C2063 vdd.n33 gnd 0.002448f
C2064 vdd.n34 gnd 0.002592f
C2065 vdd.n35 gnd 0.004556f
C2066 vdd.n36 gnd 0.002448f
C2067 vdd.n37 gnd 0.005787f
C2068 vdd.n38 gnd 0.002592f
C2069 vdd.n39 gnd 0.004556f
C2070 vdd.n40 gnd 0.002448f
C2071 vdd.n41 gnd 0.00434f
C2072 vdd.n42 gnd 0.004353f
C2073 vdd.t113 gnd 0.012433f
C2074 vdd.n43 gnd 0.027663f
C2075 vdd.n44 gnd 0.143964f
C2076 vdd.n45 gnd 0.002448f
C2077 vdd.n46 gnd 0.002592f
C2078 vdd.n47 gnd 0.005787f
C2079 vdd.n48 gnd 0.005787f
C2080 vdd.n49 gnd 0.002592f
C2081 vdd.n50 gnd 0.002448f
C2082 vdd.n51 gnd 0.004556f
C2083 vdd.n52 gnd 0.004556f
C2084 vdd.n53 gnd 0.002448f
C2085 vdd.n54 gnd 0.002592f
C2086 vdd.n55 gnd 0.005787f
C2087 vdd.n56 gnd 0.005787f
C2088 vdd.n57 gnd 0.002592f
C2089 vdd.n58 gnd 0.002448f
C2090 vdd.n59 gnd 0.004556f
C2091 vdd.n60 gnd 0.004556f
C2092 vdd.n61 gnd 0.002448f
C2093 vdd.n62 gnd 0.002592f
C2094 vdd.n63 gnd 0.005787f
C2095 vdd.n64 gnd 0.005787f
C2096 vdd.n65 gnd 0.013682f
C2097 vdd.n66 gnd 0.00252f
C2098 vdd.n67 gnd 0.002448f
C2099 vdd.n68 gnd 0.011777f
C2100 vdd.n69 gnd 0.008222f
C2101 vdd.t93 gnd 0.028804f
C2102 vdd.t144 gnd 0.028804f
C2103 vdd.n70 gnd 0.197961f
C2104 vdd.n71 gnd 0.155666f
C2105 vdd.t78 gnd 0.028804f
C2106 vdd.t129 gnd 0.028804f
C2107 vdd.n72 gnd 0.197961f
C2108 vdd.n73 gnd 0.125622f
C2109 vdd.t83 gnd 0.028804f
C2110 vdd.t140 gnd 0.028804f
C2111 vdd.n74 gnd 0.197961f
C2112 vdd.n75 gnd 0.125622f
C2113 vdd.t105 gnd 0.028804f
C2114 vdd.t148 gnd 0.028804f
C2115 vdd.n76 gnd 0.197961f
C2116 vdd.n77 gnd 0.125622f
C2117 vdd.t116 gnd 0.028804f
C2118 vdd.t135 gnd 0.028804f
C2119 vdd.n78 gnd 0.197961f
C2120 vdd.n79 gnd 0.125622f
C2121 vdd.n80 gnd 0.00491f
C2122 vdd.n81 gnd 0.004556f
C2123 vdd.n82 gnd 0.00252f
C2124 vdd.n83 gnd 0.005787f
C2125 vdd.n84 gnd 0.002448f
C2126 vdd.n85 gnd 0.002592f
C2127 vdd.n86 gnd 0.004556f
C2128 vdd.n87 gnd 0.002448f
C2129 vdd.n88 gnd 0.005787f
C2130 vdd.n89 gnd 0.002592f
C2131 vdd.n90 gnd 0.004556f
C2132 vdd.n91 gnd 0.002448f
C2133 vdd.n92 gnd 0.00434f
C2134 vdd.n93 gnd 0.004353f
C2135 vdd.t97 gnd 0.012433f
C2136 vdd.n94 gnd 0.027663f
C2137 vdd.n95 gnd 0.143964f
C2138 vdd.n96 gnd 0.002448f
C2139 vdd.n97 gnd 0.002592f
C2140 vdd.n98 gnd 0.005787f
C2141 vdd.n99 gnd 0.005787f
C2142 vdd.n100 gnd 0.002592f
C2143 vdd.n101 gnd 0.002448f
C2144 vdd.n102 gnd 0.004556f
C2145 vdd.n103 gnd 0.004556f
C2146 vdd.n104 gnd 0.002448f
C2147 vdd.n105 gnd 0.002592f
C2148 vdd.n106 gnd 0.005787f
C2149 vdd.n107 gnd 0.005787f
C2150 vdd.n108 gnd 0.002592f
C2151 vdd.n109 gnd 0.002448f
C2152 vdd.n110 gnd 0.004556f
C2153 vdd.n111 gnd 0.004556f
C2154 vdd.n112 gnd 0.002448f
C2155 vdd.n113 gnd 0.002592f
C2156 vdd.n114 gnd 0.005787f
C2157 vdd.n115 gnd 0.005787f
C2158 vdd.n116 gnd 0.013682f
C2159 vdd.n117 gnd 0.00252f
C2160 vdd.n118 gnd 0.002448f
C2161 vdd.n119 gnd 0.011777f
C2162 vdd.n120 gnd 0.007964f
C2163 vdd.n121 gnd 0.093463f
C2164 vdd.n122 gnd 0.00491f
C2165 vdd.n123 gnd 0.004556f
C2166 vdd.n124 gnd 0.00252f
C2167 vdd.n125 gnd 0.005787f
C2168 vdd.n126 gnd 0.002448f
C2169 vdd.n127 gnd 0.002592f
C2170 vdd.n128 gnd 0.004556f
C2171 vdd.n129 gnd 0.002448f
C2172 vdd.n130 gnd 0.005787f
C2173 vdd.n131 gnd 0.002592f
C2174 vdd.n132 gnd 0.004556f
C2175 vdd.n133 gnd 0.002448f
C2176 vdd.n134 gnd 0.00434f
C2177 vdd.n135 gnd 0.004353f
C2178 vdd.t146 gnd 0.012433f
C2179 vdd.n136 gnd 0.027663f
C2180 vdd.n137 gnd 0.143964f
C2181 vdd.n138 gnd 0.002448f
C2182 vdd.n139 gnd 0.002592f
C2183 vdd.n140 gnd 0.005787f
C2184 vdd.n141 gnd 0.005787f
C2185 vdd.n142 gnd 0.002592f
C2186 vdd.n143 gnd 0.002448f
C2187 vdd.n144 gnd 0.004556f
C2188 vdd.n145 gnd 0.004556f
C2189 vdd.n146 gnd 0.002448f
C2190 vdd.n147 gnd 0.002592f
C2191 vdd.n148 gnd 0.005787f
C2192 vdd.n149 gnd 0.005787f
C2193 vdd.n150 gnd 0.002592f
C2194 vdd.n151 gnd 0.002448f
C2195 vdd.n152 gnd 0.004556f
C2196 vdd.n153 gnd 0.004556f
C2197 vdd.n154 gnd 0.002448f
C2198 vdd.n155 gnd 0.002592f
C2199 vdd.n156 gnd 0.005787f
C2200 vdd.n157 gnd 0.005787f
C2201 vdd.n158 gnd 0.013682f
C2202 vdd.n159 gnd 0.00252f
C2203 vdd.n160 gnd 0.002448f
C2204 vdd.n161 gnd 0.011777f
C2205 vdd.n162 gnd 0.008222f
C2206 vdd.t147 gnd 0.028804f
C2207 vdd.t75 gnd 0.028804f
C2208 vdd.n163 gnd 0.197961f
C2209 vdd.n164 gnd 0.155666f
C2210 vdd.t137 gnd 0.028804f
C2211 vdd.t143 gnd 0.028804f
C2212 vdd.n165 gnd 0.197961f
C2213 vdd.n166 gnd 0.125622f
C2214 vdd.t71 gnd 0.028804f
C2215 vdd.t111 gnd 0.028804f
C2216 vdd.n167 gnd 0.197961f
C2217 vdd.n168 gnd 0.125622f
C2218 vdd.t134 gnd 0.028804f
C2219 vdd.t151 gnd 0.028804f
C2220 vdd.n169 gnd 0.197961f
C2221 vdd.n170 gnd 0.125622f
C2222 vdd.t99 gnd 0.028804f
C2223 vdd.t133 gnd 0.028804f
C2224 vdd.n171 gnd 0.197961f
C2225 vdd.n172 gnd 0.125622f
C2226 vdd.n173 gnd 0.00491f
C2227 vdd.n174 gnd 0.004556f
C2228 vdd.n175 gnd 0.00252f
C2229 vdd.n176 gnd 0.005787f
C2230 vdd.n177 gnd 0.002448f
C2231 vdd.n178 gnd 0.002592f
C2232 vdd.n179 gnd 0.004556f
C2233 vdd.n180 gnd 0.002448f
C2234 vdd.n181 gnd 0.005787f
C2235 vdd.n182 gnd 0.002592f
C2236 vdd.n183 gnd 0.004556f
C2237 vdd.n184 gnd 0.002448f
C2238 vdd.n185 gnd 0.00434f
C2239 vdd.n186 gnd 0.004353f
C2240 vdd.t154 gnd 0.012433f
C2241 vdd.n187 gnd 0.027663f
C2242 vdd.n188 gnd 0.143964f
C2243 vdd.n189 gnd 0.002448f
C2244 vdd.n190 gnd 0.002592f
C2245 vdd.n191 gnd 0.005787f
C2246 vdd.n192 gnd 0.005787f
C2247 vdd.n193 gnd 0.002592f
C2248 vdd.n194 gnd 0.002448f
C2249 vdd.n195 gnd 0.004556f
C2250 vdd.n196 gnd 0.004556f
C2251 vdd.n197 gnd 0.002448f
C2252 vdd.n198 gnd 0.002592f
C2253 vdd.n199 gnd 0.005787f
C2254 vdd.n200 gnd 0.005787f
C2255 vdd.n201 gnd 0.002592f
C2256 vdd.n202 gnd 0.002448f
C2257 vdd.n203 gnd 0.004556f
C2258 vdd.n204 gnd 0.004556f
C2259 vdd.n205 gnd 0.002448f
C2260 vdd.n206 gnd 0.002592f
C2261 vdd.n207 gnd 0.005787f
C2262 vdd.n208 gnd 0.005787f
C2263 vdd.n209 gnd 0.013682f
C2264 vdd.n210 gnd 0.00252f
C2265 vdd.n211 gnd 0.002448f
C2266 vdd.n212 gnd 0.011777f
C2267 vdd.n213 gnd 0.007964f
C2268 vdd.n214 gnd 0.055601f
C2269 vdd.n215 gnd 0.200345f
C2270 vdd.n216 gnd 0.00491f
C2271 vdd.n217 gnd 0.004556f
C2272 vdd.n218 gnd 0.00252f
C2273 vdd.n219 gnd 0.005787f
C2274 vdd.n220 gnd 0.002448f
C2275 vdd.n221 gnd 0.002592f
C2276 vdd.n222 gnd 0.004556f
C2277 vdd.n223 gnd 0.002448f
C2278 vdd.n224 gnd 0.005787f
C2279 vdd.n225 gnd 0.002592f
C2280 vdd.n226 gnd 0.004556f
C2281 vdd.n227 gnd 0.002448f
C2282 vdd.n228 gnd 0.00434f
C2283 vdd.n229 gnd 0.004353f
C2284 vdd.t152 gnd 0.012433f
C2285 vdd.n230 gnd 0.027663f
C2286 vdd.n231 gnd 0.143964f
C2287 vdd.n232 gnd 0.002448f
C2288 vdd.n233 gnd 0.002592f
C2289 vdd.n234 gnd 0.005787f
C2290 vdd.n235 gnd 0.005787f
C2291 vdd.n236 gnd 0.002592f
C2292 vdd.n237 gnd 0.002448f
C2293 vdd.n238 gnd 0.004556f
C2294 vdd.n239 gnd 0.004556f
C2295 vdd.n240 gnd 0.002448f
C2296 vdd.n241 gnd 0.002592f
C2297 vdd.n242 gnd 0.005787f
C2298 vdd.n243 gnd 0.005787f
C2299 vdd.n244 gnd 0.002592f
C2300 vdd.n245 gnd 0.002448f
C2301 vdd.n246 gnd 0.004556f
C2302 vdd.n247 gnd 0.004556f
C2303 vdd.n248 gnd 0.002448f
C2304 vdd.n249 gnd 0.002592f
C2305 vdd.n250 gnd 0.005787f
C2306 vdd.n251 gnd 0.005787f
C2307 vdd.n252 gnd 0.013682f
C2308 vdd.n253 gnd 0.00252f
C2309 vdd.n254 gnd 0.002448f
C2310 vdd.n255 gnd 0.011777f
C2311 vdd.n256 gnd 0.008222f
C2312 vdd.t153 gnd 0.028804f
C2313 vdd.t91 gnd 0.028804f
C2314 vdd.n257 gnd 0.197961f
C2315 vdd.n258 gnd 0.155666f
C2316 vdd.t142 gnd 0.028804f
C2317 vdd.t150 gnd 0.028804f
C2318 vdd.n259 gnd 0.197961f
C2319 vdd.n260 gnd 0.125622f
C2320 vdd.t84 gnd 0.028804f
C2321 vdd.t124 gnd 0.028804f
C2322 vdd.n261 gnd 0.197961f
C2323 vdd.n262 gnd 0.125622f
C2324 vdd.t141 gnd 0.028804f
C2325 vdd.t65 gnd 0.028804f
C2326 vdd.n263 gnd 0.197961f
C2327 vdd.n264 gnd 0.125622f
C2328 vdd.t108 gnd 0.028804f
C2329 vdd.t139 gnd 0.028804f
C2330 vdd.n265 gnd 0.197961f
C2331 vdd.n266 gnd 0.125622f
C2332 vdd.n267 gnd 0.00491f
C2333 vdd.n268 gnd 0.004556f
C2334 vdd.n269 gnd 0.00252f
C2335 vdd.n270 gnd 0.005787f
C2336 vdd.n271 gnd 0.002448f
C2337 vdd.n272 gnd 0.002592f
C2338 vdd.n273 gnd 0.004556f
C2339 vdd.n274 gnd 0.002448f
C2340 vdd.n275 gnd 0.005787f
C2341 vdd.n276 gnd 0.002592f
C2342 vdd.n277 gnd 0.004556f
C2343 vdd.n278 gnd 0.002448f
C2344 vdd.n279 gnd 0.00434f
C2345 vdd.n280 gnd 0.004353f
C2346 vdd.t73 gnd 0.012433f
C2347 vdd.n281 gnd 0.027663f
C2348 vdd.n282 gnd 0.143964f
C2349 vdd.n283 gnd 0.002448f
C2350 vdd.n284 gnd 0.002592f
C2351 vdd.n285 gnd 0.005787f
C2352 vdd.n286 gnd 0.005787f
C2353 vdd.n287 gnd 0.002592f
C2354 vdd.n288 gnd 0.002448f
C2355 vdd.n289 gnd 0.004556f
C2356 vdd.n290 gnd 0.004556f
C2357 vdd.n291 gnd 0.002448f
C2358 vdd.n292 gnd 0.002592f
C2359 vdd.n293 gnd 0.005787f
C2360 vdd.n294 gnd 0.005787f
C2361 vdd.n295 gnd 0.002592f
C2362 vdd.n296 gnd 0.002448f
C2363 vdd.n297 gnd 0.004556f
C2364 vdd.n298 gnd 0.004556f
C2365 vdd.n299 gnd 0.002448f
C2366 vdd.n300 gnd 0.002592f
C2367 vdd.n301 gnd 0.005787f
C2368 vdd.n302 gnd 0.005787f
C2369 vdd.n303 gnd 0.013682f
C2370 vdd.n304 gnd 0.00252f
C2371 vdd.n305 gnd 0.002448f
C2372 vdd.n306 gnd 0.011777f
C2373 vdd.n307 gnd 0.007964f
C2374 vdd.n308 gnd 0.055601f
C2375 vdd.n309 gnd 0.220186f
C2376 vdd.n310 gnd 0.008916f
C2377 vdd.n311 gnd 0.008916f
C2378 vdd.n312 gnd 0.007201f
C2379 vdd.n313 gnd 0.007201f
C2380 vdd.n314 gnd 0.008947f
C2381 vdd.n315 gnd 0.008947f
C2382 vdd.t70 gnd 0.457154f
C2383 vdd.n316 gnd 0.008947f
C2384 vdd.n317 gnd 0.008947f
C2385 vdd.n318 gnd 0.008947f
C2386 vdd.t104 gnd 0.457154f
C2387 vdd.n319 gnd 0.008947f
C2388 vdd.n320 gnd 0.008947f
C2389 vdd.n321 gnd 0.008947f
C2390 vdd.n322 gnd 0.008947f
C2391 vdd.n323 gnd 0.007201f
C2392 vdd.n324 gnd 0.008947f
C2393 vdd.n325 gnd 0.736018f
C2394 vdd.n326 gnd 0.008947f
C2395 vdd.n327 gnd 0.008947f
C2396 vdd.n328 gnd 0.008947f
C2397 vdd.n329 gnd 0.626301f
C2398 vdd.n330 gnd 0.008947f
C2399 vdd.n331 gnd 0.008947f
C2400 vdd.n332 gnd 0.008947f
C2401 vdd.n333 gnd 0.008947f
C2402 vdd.n334 gnd 0.008947f
C2403 vdd.n335 gnd 0.007201f
C2404 vdd.n336 gnd 0.008947f
C2405 vdd.t132 gnd 0.457154f
C2406 vdd.n337 gnd 0.008947f
C2407 vdd.n338 gnd 0.008947f
C2408 vdd.n339 gnd 0.008947f
C2409 vdd.n340 gnd 0.914309f
C2410 vdd.n341 gnd 0.008947f
C2411 vdd.n342 gnd 0.008947f
C2412 vdd.n343 gnd 0.008947f
C2413 vdd.n344 gnd 0.008947f
C2414 vdd.n345 gnd 0.008947f
C2415 vdd.n346 gnd 0.007201f
C2416 vdd.n347 gnd 0.008947f
C2417 vdd.n348 gnd 0.008947f
C2418 vdd.n349 gnd 0.008947f
C2419 vdd.n350 gnd 0.021084f
C2420 vdd.n351 gnd 2.10291f
C2421 vdd.n352 gnd 0.021413f
C2422 vdd.n353 gnd 0.008947f
C2423 vdd.n354 gnd 0.008947f
C2424 vdd.n356 gnd 0.008947f
C2425 vdd.n357 gnd 0.008947f
C2426 vdd.n358 gnd 0.007201f
C2427 vdd.n359 gnd 0.007201f
C2428 vdd.n360 gnd 0.008947f
C2429 vdd.n361 gnd 0.008947f
C2430 vdd.n362 gnd 0.008947f
C2431 vdd.n363 gnd 0.008947f
C2432 vdd.n364 gnd 0.008947f
C2433 vdd.n365 gnd 0.008947f
C2434 vdd.n366 gnd 0.007201f
C2435 vdd.n368 gnd 0.008947f
C2436 vdd.n369 gnd 0.008947f
C2437 vdd.n370 gnd 0.008947f
C2438 vdd.n371 gnd 0.008947f
C2439 vdd.n372 gnd 0.008947f
C2440 vdd.n373 gnd 0.007201f
C2441 vdd.n375 gnd 0.008947f
C2442 vdd.n376 gnd 0.008947f
C2443 vdd.n377 gnd 0.008947f
C2444 vdd.n378 gnd 0.008947f
C2445 vdd.n379 gnd 0.008947f
C2446 vdd.n380 gnd 0.007201f
C2447 vdd.n382 gnd 0.008947f
C2448 vdd.n383 gnd 0.008947f
C2449 vdd.n384 gnd 0.008947f
C2450 vdd.n385 gnd 0.008947f
C2451 vdd.n386 gnd 0.006013f
C2452 vdd.t202 gnd 0.110068f
C2453 vdd.t201 gnd 0.117632f
C2454 vdd.t200 gnd 0.143747f
C2455 vdd.n387 gnd 0.184263f
C2456 vdd.n388 gnd 0.155535f
C2457 vdd.n390 gnd 0.008947f
C2458 vdd.n391 gnd 0.008947f
C2459 vdd.n392 gnd 0.007201f
C2460 vdd.n393 gnd 0.008947f
C2461 vdd.n395 gnd 0.008947f
C2462 vdd.n396 gnd 0.008947f
C2463 vdd.n397 gnd 0.008947f
C2464 vdd.n398 gnd 0.008947f
C2465 vdd.n399 gnd 0.007201f
C2466 vdd.n401 gnd 0.008947f
C2467 vdd.n402 gnd 0.008947f
C2468 vdd.n403 gnd 0.008947f
C2469 vdd.n404 gnd 0.008947f
C2470 vdd.n405 gnd 0.008947f
C2471 vdd.n406 gnd 0.007201f
C2472 vdd.n408 gnd 0.008947f
C2473 vdd.n409 gnd 0.008947f
C2474 vdd.n410 gnd 0.008947f
C2475 vdd.n411 gnd 0.008947f
C2476 vdd.n412 gnd 0.008947f
C2477 vdd.n413 gnd 0.007201f
C2478 vdd.n415 gnd 0.008947f
C2479 vdd.n416 gnd 0.008947f
C2480 vdd.n417 gnd 0.008947f
C2481 vdd.n418 gnd 0.008947f
C2482 vdd.n419 gnd 0.008947f
C2483 vdd.n420 gnd 0.007201f
C2484 vdd.n422 gnd 0.008947f
C2485 vdd.n423 gnd 0.008947f
C2486 vdd.n424 gnd 0.008947f
C2487 vdd.n425 gnd 0.008947f
C2488 vdd.n426 gnd 0.007129f
C2489 vdd.t185 gnd 0.110068f
C2490 vdd.t184 gnd 0.117632f
C2491 vdd.t182 gnd 0.143747f
C2492 vdd.n427 gnd 0.184263f
C2493 vdd.n428 gnd 0.155535f
C2494 vdd.n430 gnd 0.008947f
C2495 vdd.n431 gnd 0.008947f
C2496 vdd.n432 gnd 0.007201f
C2497 vdd.n433 gnd 0.008947f
C2498 vdd.n435 gnd 0.008947f
C2499 vdd.n436 gnd 0.008947f
C2500 vdd.n437 gnd 0.008947f
C2501 vdd.n438 gnd 0.008947f
C2502 vdd.n439 gnd 0.007201f
C2503 vdd.n441 gnd 0.008947f
C2504 vdd.n442 gnd 0.008947f
C2505 vdd.n443 gnd 0.008947f
C2506 vdd.n444 gnd 0.008947f
C2507 vdd.n445 gnd 0.008947f
C2508 vdd.n446 gnd 0.007201f
C2509 vdd.n448 gnd 0.008947f
C2510 vdd.n449 gnd 0.008947f
C2511 vdd.n450 gnd 0.008947f
C2512 vdd.n451 gnd 0.008947f
C2513 vdd.n452 gnd 0.008947f
C2514 vdd.n453 gnd 0.007201f
C2515 vdd.n455 gnd 0.008947f
C2516 vdd.n456 gnd 0.008947f
C2517 vdd.n457 gnd 0.008947f
C2518 vdd.n458 gnd 0.008947f
C2519 vdd.n459 gnd 0.008947f
C2520 vdd.n460 gnd 0.007201f
C2521 vdd.n462 gnd 0.008947f
C2522 vdd.n463 gnd 0.008947f
C2523 vdd.n464 gnd 0.008947f
C2524 vdd.n465 gnd 0.008947f
C2525 vdd.n466 gnd 0.008947f
C2526 vdd.n467 gnd 0.008947f
C2527 vdd.n468 gnd 0.007201f
C2528 vdd.n469 gnd 0.008947f
C2529 vdd.n470 gnd 0.008947f
C2530 vdd.n471 gnd 0.007201f
C2531 vdd.n472 gnd 0.008947f
C2532 vdd.n473 gnd 0.008947f
C2533 vdd.n474 gnd 0.007201f
C2534 vdd.n475 gnd 0.008947f
C2535 vdd.n476 gnd 0.007201f
C2536 vdd.n477 gnd 0.008947f
C2537 vdd.n478 gnd 0.007201f
C2538 vdd.n479 gnd 0.008947f
C2539 vdd.n480 gnd 0.008947f
C2540 vdd.t128 gnd 0.457154f
C2541 vdd.n481 gnd 0.489155f
C2542 vdd.n482 gnd 0.008947f
C2543 vdd.n483 gnd 0.007201f
C2544 vdd.n484 gnd 0.008947f
C2545 vdd.n485 gnd 0.007201f
C2546 vdd.n486 gnd 0.008947f
C2547 vdd.t77 gnd 0.457154f
C2548 vdd.n487 gnd 0.008947f
C2549 vdd.n488 gnd 0.007201f
C2550 vdd.n489 gnd 0.008947f
C2551 vdd.n490 gnd 0.007201f
C2552 vdd.n491 gnd 0.008947f
C2553 vdd.n492 gnd 0.717732f
C2554 vdd.n493 gnd 0.758876f
C2555 vdd.t74 gnd 0.457154f
C2556 vdd.n494 gnd 0.008947f
C2557 vdd.n495 gnd 0.007201f
C2558 vdd.n496 gnd 0.008947f
C2559 vdd.n497 gnd 0.007201f
C2560 vdd.n498 gnd 0.008947f
C2561 vdd.n499 gnd 0.5623f
C2562 vdd.n500 gnd 0.008947f
C2563 vdd.n501 gnd 0.007201f
C2564 vdd.n502 gnd 0.008947f
C2565 vdd.n503 gnd 0.007201f
C2566 vdd.n504 gnd 0.008947f
C2567 vdd.n505 gnd 0.914309f
C2568 vdd.t112 gnd 0.457154f
C2569 vdd.n506 gnd 0.008947f
C2570 vdd.n507 gnd 0.007201f
C2571 vdd.n508 gnd 0.008947f
C2572 vdd.n509 gnd 0.007201f
C2573 vdd.n510 gnd 0.008947f
C2574 vdd.n511 gnd 0.489155f
C2575 vdd.n512 gnd 0.008947f
C2576 vdd.n513 gnd 0.007201f
C2577 vdd.n514 gnd 0.021413f
C2578 vdd.n515 gnd 0.021413f
C2579 vdd.n516 gnd 11.0997f
C2580 vdd.t179 gnd 0.457154f
C2581 vdd.n517 gnd 0.021413f
C2582 vdd.n518 gnd 0.007694f
C2583 vdd.n519 gnd 0.007201f
C2584 vdd.n524 gnd 0.005726f
C2585 vdd.n525 gnd 0.007201f
C2586 vdd.n526 gnd 0.008947f
C2587 vdd.n527 gnd 0.008947f
C2588 vdd.n528 gnd 0.008947f
C2589 vdd.n529 gnd 0.008947f
C2590 vdd.n530 gnd 0.008947f
C2591 vdd.n531 gnd 0.007201f
C2592 vdd.n532 gnd 0.008947f
C2593 vdd.n533 gnd 0.008947f
C2594 vdd.n534 gnd 0.008947f
C2595 vdd.n535 gnd 0.008947f
C2596 vdd.n536 gnd 0.008947f
C2597 vdd.n537 gnd 0.007201f
C2598 vdd.n538 gnd 0.008947f
C2599 vdd.n539 gnd 0.008947f
C2600 vdd.n540 gnd 0.008947f
C2601 vdd.n541 gnd 0.008947f
C2602 vdd.n542 gnd 0.008947f
C2603 vdd.t214 gnd 0.110068f
C2604 vdd.t215 gnd 0.117632f
C2605 vdd.t213 gnd 0.143747f
C2606 vdd.n543 gnd 0.184263f
C2607 vdd.n544 gnd 0.154815f
C2608 vdd.n545 gnd 0.01469f
C2609 vdd.n546 gnd 0.008947f
C2610 vdd.n547 gnd 0.008947f
C2611 vdd.n548 gnd 0.008947f
C2612 vdd.n549 gnd 0.008947f
C2613 vdd.n550 gnd 0.008947f
C2614 vdd.n551 gnd 0.007201f
C2615 vdd.n552 gnd 0.008947f
C2616 vdd.n553 gnd 0.008947f
C2617 vdd.n554 gnd 0.008947f
C2618 vdd.n555 gnd 0.008947f
C2619 vdd.n556 gnd 0.008947f
C2620 vdd.n557 gnd 0.007201f
C2621 vdd.n558 gnd 0.008947f
C2622 vdd.n559 gnd 0.008947f
C2623 vdd.n560 gnd 0.008947f
C2624 vdd.n561 gnd 0.008947f
C2625 vdd.n562 gnd 0.008947f
C2626 vdd.n563 gnd 0.007201f
C2627 vdd.n564 gnd 0.008947f
C2628 vdd.n565 gnd 0.008947f
C2629 vdd.n566 gnd 0.008947f
C2630 vdd.n567 gnd 0.008947f
C2631 vdd.n568 gnd 0.008947f
C2632 vdd.n569 gnd 0.007201f
C2633 vdd.n570 gnd 0.008947f
C2634 vdd.n571 gnd 0.008947f
C2635 vdd.n572 gnd 0.008947f
C2636 vdd.n573 gnd 0.008947f
C2637 vdd.n574 gnd 0.008947f
C2638 vdd.n575 gnd 0.007201f
C2639 vdd.n576 gnd 0.008947f
C2640 vdd.n577 gnd 0.008947f
C2641 vdd.n578 gnd 0.008947f
C2642 vdd.n579 gnd 0.007129f
C2643 vdd.t204 gnd 0.110068f
C2644 vdd.t205 gnd 0.117632f
C2645 vdd.t203 gnd 0.143747f
C2646 vdd.n580 gnd 0.184263f
C2647 vdd.n581 gnd 0.154815f
C2648 vdd.n582 gnd 0.008947f
C2649 vdd.n583 gnd 0.007201f
C2650 vdd.n585 gnd 0.008947f
C2651 vdd.n587 gnd 0.008947f
C2652 vdd.n588 gnd 0.008947f
C2653 vdd.n589 gnd 0.007201f
C2654 vdd.n590 gnd 0.008947f
C2655 vdd.n591 gnd 0.008947f
C2656 vdd.n592 gnd 0.008947f
C2657 vdd.n593 gnd 0.008947f
C2658 vdd.n594 gnd 0.008947f
C2659 vdd.n595 gnd 0.007201f
C2660 vdd.n596 gnd 0.008947f
C2661 vdd.n597 gnd 0.008947f
C2662 vdd.n598 gnd 0.008947f
C2663 vdd.n599 gnd 0.008947f
C2664 vdd.n600 gnd 0.008947f
C2665 vdd.n601 gnd 0.007201f
C2666 vdd.n602 gnd 0.008947f
C2667 vdd.n603 gnd 0.008947f
C2668 vdd.n604 gnd 0.008947f
C2669 vdd.n605 gnd 0.005726f
C2670 vdd.n610 gnd 0.006084f
C2671 vdd.n611 gnd 0.006084f
C2672 vdd.n612 gnd 0.006084f
C2673 vdd.n613 gnd 10.797999f
C2674 vdd.n614 gnd 0.006084f
C2675 vdd.n615 gnd 0.006084f
C2676 vdd.n616 gnd 0.006084f
C2677 vdd.n618 gnd 0.006084f
C2678 vdd.n619 gnd 0.006084f
C2679 vdd.n621 gnd 0.006084f
C2680 vdd.n622 gnd 0.004429f
C2681 vdd.n624 gnd 0.006084f
C2682 vdd.t163 gnd 0.245843f
C2683 vdd.t162 gnd 0.251651f
C2684 vdd.t160 gnd 0.160496f
C2685 vdd.n625 gnd 0.086739f
C2686 vdd.n626 gnd 0.049201f
C2687 vdd.n627 gnd 0.008695f
C2688 vdd.n628 gnd 0.013814f
C2689 vdd.n630 gnd 0.006084f
C2690 vdd.n631 gnd 0.62173f
C2691 vdd.n632 gnd 0.013026f
C2692 vdd.n633 gnd 0.013026f
C2693 vdd.n634 gnd 0.006084f
C2694 vdd.n635 gnd 0.013814f
C2695 vdd.n636 gnd 0.006084f
C2696 vdd.n637 gnd 0.006084f
C2697 vdd.n638 gnd 0.006084f
C2698 vdd.n639 gnd 0.006084f
C2699 vdd.n640 gnd 0.006084f
C2700 vdd.n642 gnd 0.006084f
C2701 vdd.n643 gnd 0.006084f
C2702 vdd.n645 gnd 0.006084f
C2703 vdd.n646 gnd 0.006084f
C2704 vdd.n648 gnd 0.006084f
C2705 vdd.n649 gnd 0.006084f
C2706 vdd.n651 gnd 0.006084f
C2707 vdd.n652 gnd 0.006084f
C2708 vdd.n654 gnd 0.006084f
C2709 vdd.n655 gnd 0.006084f
C2710 vdd.n657 gnd 0.006084f
C2711 vdd.n658 gnd 0.004429f
C2712 vdd.n660 gnd 0.006084f
C2713 vdd.t177 gnd 0.245843f
C2714 vdd.t176 gnd 0.251651f
C2715 vdd.t175 gnd 0.160496f
C2716 vdd.n661 gnd 0.086739f
C2717 vdd.n662 gnd 0.049201f
C2718 vdd.n663 gnd 0.008695f
C2719 vdd.n664 gnd 0.006084f
C2720 vdd.n665 gnd 0.006084f
C2721 vdd.t161 gnd 0.310865f
C2722 vdd.n666 gnd 0.006084f
C2723 vdd.n667 gnd 0.006084f
C2724 vdd.n668 gnd 0.006084f
C2725 vdd.n669 gnd 0.006084f
C2726 vdd.n670 gnd 0.006084f
C2727 vdd.n671 gnd 0.62173f
C2728 vdd.n672 gnd 0.006084f
C2729 vdd.n673 gnd 0.006084f
C2730 vdd.n674 gnd 0.489155f
C2731 vdd.n675 gnd 0.006084f
C2732 vdd.n676 gnd 0.006084f
C2733 vdd.n677 gnd 0.006084f
C2734 vdd.n678 gnd 0.006084f
C2735 vdd.n679 gnd 0.62173f
C2736 vdd.n680 gnd 0.006084f
C2737 vdd.n681 gnd 0.006084f
C2738 vdd.n682 gnd 0.006084f
C2739 vdd.n683 gnd 0.006084f
C2740 vdd.n684 gnd 0.006084f
C2741 vdd.t15 gnd 0.310865f
C2742 vdd.n685 gnd 0.006084f
C2743 vdd.n686 gnd 0.006084f
C2744 vdd.n687 gnd 0.006084f
C2745 vdd.n688 gnd 0.006084f
C2746 vdd.n689 gnd 0.006084f
C2747 vdd.t32 gnd 0.310865f
C2748 vdd.n690 gnd 0.006084f
C2749 vdd.n691 gnd 0.006084f
C2750 vdd.n692 gnd 0.598872f
C2751 vdd.n693 gnd 0.006084f
C2752 vdd.n694 gnd 0.006084f
C2753 vdd.n695 gnd 0.006084f
C2754 vdd.t31 gnd 0.310865f
C2755 vdd.n696 gnd 0.006084f
C2756 vdd.n697 gnd 0.006084f
C2757 vdd.n698 gnd 0.461726f
C2758 vdd.n699 gnd 0.006084f
C2759 vdd.n700 gnd 0.006084f
C2760 vdd.n701 gnd 0.006084f
C2761 vdd.n702 gnd 0.434297f
C2762 vdd.n703 gnd 0.006084f
C2763 vdd.n704 gnd 0.006084f
C2764 vdd.n705 gnd 0.32458f
C2765 vdd.n706 gnd 0.006084f
C2766 vdd.n707 gnd 0.006084f
C2767 vdd.n708 gnd 0.006084f
C2768 vdd.n709 gnd 0.571443f
C2769 vdd.n710 gnd 0.006084f
C2770 vdd.n711 gnd 0.006084f
C2771 vdd.t38 gnd 0.310865f
C2772 vdd.n712 gnd 0.006084f
C2773 vdd.n713 gnd 0.006084f
C2774 vdd.n714 gnd 0.006084f
C2775 vdd.n715 gnd 0.62173f
C2776 vdd.n716 gnd 0.006084f
C2777 vdd.n717 gnd 0.006084f
C2778 vdd.t39 gnd 0.310865f
C2779 vdd.n718 gnd 0.006084f
C2780 vdd.n719 gnd 0.006084f
C2781 vdd.n720 gnd 0.006084f
C2782 vdd.t9 gnd 0.310865f
C2783 vdd.n721 gnd 0.006084f
C2784 vdd.n722 gnd 0.006084f
C2785 vdd.n723 gnd 0.006084f
C2786 vdd.t188 gnd 0.251651f
C2787 vdd.t186 gnd 0.160496f
C2788 vdd.t189 gnd 0.251651f
C2789 vdd.n724 gnd 0.141438f
C2790 vdd.n725 gnd 0.017624f
C2791 vdd.n726 gnd 0.006084f
C2792 vdd.t187 gnd 0.224006f
C2793 vdd.n727 gnd 0.006084f
C2794 vdd.n728 gnd 0.006084f
C2795 vdd.n729 gnd 0.534871f
C2796 vdd.n730 gnd 0.006084f
C2797 vdd.n731 gnd 0.006084f
C2798 vdd.n732 gnd 0.006084f
C2799 vdd.n733 gnd 0.361152f
C2800 vdd.n734 gnd 0.006084f
C2801 vdd.n735 gnd 0.006084f
C2802 vdd.t10 gnd 0.128003f
C2803 vdd.n736 gnd 0.397724f
C2804 vdd.n737 gnd 0.006084f
C2805 vdd.n738 gnd 0.006084f
C2806 vdd.n739 gnd 0.006084f
C2807 vdd.n740 gnd 0.498298f
C2808 vdd.n741 gnd 0.006084f
C2809 vdd.n742 gnd 0.006084f
C2810 vdd.t23 gnd 0.310865f
C2811 vdd.n743 gnd 0.006084f
C2812 vdd.n744 gnd 0.006084f
C2813 vdd.n745 gnd 0.006084f
C2814 vdd.t19 gnd 0.310865f
C2815 vdd.n746 gnd 0.006084f
C2816 vdd.n747 gnd 0.006084f
C2817 vdd.t42 gnd 0.310865f
C2818 vdd.n748 gnd 0.006084f
C2819 vdd.n749 gnd 0.006084f
C2820 vdd.n750 gnd 0.006084f
C2821 vdd.t1 gnd 0.210291f
C2822 vdd.n751 gnd 0.006084f
C2823 vdd.n752 gnd 0.006084f
C2824 vdd.n753 gnd 0.548585f
C2825 vdd.n754 gnd 0.006084f
C2826 vdd.n755 gnd 0.006084f
C2827 vdd.n756 gnd 0.006084f
C2828 vdd.t43 gnd 0.310865f
C2829 vdd.n757 gnd 0.006084f
C2830 vdd.n758 gnd 0.006084f
C2831 vdd.t55 gnd 0.29715f
C2832 vdd.n759 gnd 0.411439f
C2833 vdd.n760 gnd 0.006084f
C2834 vdd.n761 gnd 0.006084f
C2835 vdd.n762 gnd 0.006084f
C2836 vdd.t5 gnd 0.310865f
C2837 vdd.n763 gnd 0.006084f
C2838 vdd.n764 gnd 0.006084f
C2839 vdd.t47 gnd 0.310865f
C2840 vdd.n765 gnd 0.006084f
C2841 vdd.n766 gnd 0.006084f
C2842 vdd.n767 gnd 0.006084f
C2843 vdd.n768 gnd 0.62173f
C2844 vdd.n769 gnd 0.006084f
C2845 vdd.n770 gnd 0.006084f
C2846 vdd.t27 gnd 0.310865f
C2847 vdd.n771 gnd 0.006084f
C2848 vdd.n772 gnd 0.006084f
C2849 vdd.n773 gnd 0.006084f
C2850 vdd.n774 gnd 0.429725f
C2851 vdd.n775 gnd 0.006084f
C2852 vdd.n776 gnd 0.006084f
C2853 vdd.n777 gnd 0.006084f
C2854 vdd.n778 gnd 0.006084f
C2855 vdd.n779 gnd 0.006084f
C2856 vdd.t217 gnd 0.310865f
C2857 vdd.n780 gnd 0.006084f
C2858 vdd.n781 gnd 0.006084f
C2859 vdd.t7 gnd 0.310865f
C2860 vdd.n782 gnd 0.006084f
C2861 vdd.n783 gnd 0.013026f
C2862 vdd.n784 gnd 0.013026f
C2863 vdd.n785 gnd 0.704018f
C2864 vdd.n786 gnd 0.006084f
C2865 vdd.n787 gnd 0.006084f
C2866 vdd.t36 gnd 0.310865f
C2867 vdd.n788 gnd 0.013026f
C2868 vdd.n789 gnd 0.006084f
C2869 vdd.n790 gnd 0.006084f
C2870 vdd.t49 gnd 0.530299f
C2871 vdd.n808 gnd 0.013814f
C2872 vdd.n826 gnd 0.013026f
C2873 vdd.n827 gnd 0.006084f
C2874 vdd.n828 gnd 0.013026f
C2875 vdd.t235 gnd 0.245843f
C2876 vdd.t234 gnd 0.251651f
C2877 vdd.t233 gnd 0.160496f
C2878 vdd.n829 gnd 0.086739f
C2879 vdd.n830 gnd 0.049201f
C2880 vdd.n831 gnd 0.013814f
C2881 vdd.n832 gnd 0.006084f
C2882 vdd.n833 gnd 0.365723f
C2883 vdd.n834 gnd 0.013026f
C2884 vdd.n835 gnd 0.006084f
C2885 vdd.n836 gnd 0.013814f
C2886 vdd.n837 gnd 0.006084f
C2887 vdd.t212 gnd 0.245843f
C2888 vdd.t211 gnd 0.251651f
C2889 vdd.t209 gnd 0.160496f
C2890 vdd.n838 gnd 0.086739f
C2891 vdd.n839 gnd 0.049201f
C2892 vdd.n840 gnd 0.008695f
C2893 vdd.n841 gnd 0.006084f
C2894 vdd.n842 gnd 0.006084f
C2895 vdd.t210 gnd 0.310865f
C2896 vdd.n843 gnd 0.006084f
C2897 vdd.t51 gnd 0.310865f
C2898 vdd.n844 gnd 0.006084f
C2899 vdd.n845 gnd 0.006084f
C2900 vdd.n846 gnd 0.006084f
C2901 vdd.n847 gnd 0.006084f
C2902 vdd.n848 gnd 0.006084f
C2903 vdd.n849 gnd 0.62173f
C2904 vdd.n850 gnd 0.006084f
C2905 vdd.n851 gnd 0.006084f
C2906 vdd.t21 gnd 0.310865f
C2907 vdd.n852 gnd 0.006084f
C2908 vdd.n853 gnd 0.006084f
C2909 vdd.n854 gnd 0.006084f
C2910 vdd.n855 gnd 0.006084f
C2911 vdd.n856 gnd 0.448011f
C2912 vdd.n857 gnd 0.006084f
C2913 vdd.n858 gnd 0.006084f
C2914 vdd.n859 gnd 0.006084f
C2915 vdd.n860 gnd 0.006084f
C2916 vdd.n861 gnd 0.006084f
C2917 vdd.t2 gnd 0.310865f
C2918 vdd.n862 gnd 0.006084f
C2919 vdd.n863 gnd 0.006084f
C2920 vdd.t40 gnd 0.310865f
C2921 vdd.n864 gnd 0.006084f
C2922 vdd.n865 gnd 0.006084f
C2923 vdd.n866 gnd 0.006084f
C2924 vdd.t26 gnd 0.310865f
C2925 vdd.n867 gnd 0.006084f
C2926 vdd.n868 gnd 0.006084f
C2927 vdd.t3 gnd 0.310865f
C2928 vdd.n869 gnd 0.006084f
C2929 vdd.n870 gnd 0.006084f
C2930 vdd.n871 gnd 0.006084f
C2931 vdd.t24 gnd 0.29715f
C2932 vdd.n872 gnd 0.006084f
C2933 vdd.n873 gnd 0.006084f
C2934 vdd.n874 gnd 0.461726f
C2935 vdd.n875 gnd 0.006084f
C2936 vdd.n876 gnd 0.006084f
C2937 vdd.n877 gnd 0.006084f
C2938 vdd.t44 gnd 0.310865f
C2939 vdd.n878 gnd 0.006084f
C2940 vdd.n879 gnd 0.006084f
C2941 vdd.t12 gnd 0.210291f
C2942 vdd.n880 gnd 0.32458f
C2943 vdd.n881 gnd 0.006084f
C2944 vdd.n882 gnd 0.006084f
C2945 vdd.n883 gnd 0.006084f
C2946 vdd.n884 gnd 0.571443f
C2947 vdd.n885 gnd 0.006084f
C2948 vdd.n886 gnd 0.006084f
C2949 vdd.t53 gnd 0.310865f
C2950 vdd.n887 gnd 0.006084f
C2951 vdd.n888 gnd 0.006084f
C2952 vdd.n889 gnd 0.006084f
C2953 vdd.n890 gnd 0.62173f
C2954 vdd.n891 gnd 0.006084f
C2955 vdd.n892 gnd 0.006084f
C2956 vdd.t18 gnd 0.310865f
C2957 vdd.n893 gnd 0.006084f
C2958 vdd.n894 gnd 0.006084f
C2959 vdd.n895 gnd 0.006084f
C2960 vdd.t11 gnd 0.128003f
C2961 vdd.n896 gnd 0.006084f
C2962 vdd.n897 gnd 0.006084f
C2963 vdd.n898 gnd 0.006084f
C2964 vdd.t225 gnd 0.251651f
C2965 vdd.t223 gnd 0.160496f
C2966 vdd.t226 gnd 0.251651f
C2967 vdd.n899 gnd 0.141438f
C2968 vdd.n900 gnd 0.006084f
C2969 vdd.n901 gnd 0.006084f
C2970 vdd.t33 gnd 0.310865f
C2971 vdd.n902 gnd 0.006084f
C2972 vdd.n903 gnd 0.006084f
C2973 vdd.t224 gnd 0.224006f
C2974 vdd.n904 gnd 0.493727f
C2975 vdd.n905 gnd 0.006084f
C2976 vdd.n906 gnd 0.006084f
C2977 vdd.n907 gnd 0.006084f
C2978 vdd.n908 gnd 0.361152f
C2979 vdd.n909 gnd 0.006084f
C2980 vdd.n910 gnd 0.006084f
C2981 vdd.n911 gnd 0.397724f
C2982 vdd.n912 gnd 0.006084f
C2983 vdd.n913 gnd 0.006084f
C2984 vdd.n914 gnd 0.006084f
C2985 vdd.n915 gnd 0.498298f
C2986 vdd.n916 gnd 0.006084f
C2987 vdd.n917 gnd 0.006084f
C2988 vdd.t13 gnd 0.310865f
C2989 vdd.n918 gnd 0.006084f
C2990 vdd.n919 gnd 0.006084f
C2991 vdd.n920 gnd 0.006084f
C2992 vdd.n921 gnd 0.62173f
C2993 vdd.n922 gnd 0.006084f
C2994 vdd.n923 gnd 0.006084f
C2995 vdd.t14 gnd 0.310865f
C2996 vdd.n924 gnd 0.006084f
C2997 vdd.n925 gnd 0.006084f
C2998 vdd.n926 gnd 0.006084f
C2999 vdd.t54 gnd 0.310865f
C3000 vdd.n927 gnd 0.006084f
C3001 vdd.n928 gnd 0.006084f
C3002 vdd.n929 gnd 0.006084f
C3003 vdd.n930 gnd 0.006084f
C3004 vdd.n931 gnd 0.006084f
C3005 vdd.t46 gnd 0.310865f
C3006 vdd.n932 gnd 0.006084f
C3007 vdd.n933 gnd 0.006084f
C3008 vdd.n934 gnd 0.608015f
C3009 vdd.n935 gnd 0.006084f
C3010 vdd.n936 gnd 0.006084f
C3011 vdd.n937 gnd 0.006084f
C3012 vdd.t6 gnd 0.310865f
C3013 vdd.n938 gnd 0.006084f
C3014 vdd.n939 gnd 0.006084f
C3015 vdd.n940 gnd 0.470869f
C3016 vdd.n941 gnd 0.006084f
C3017 vdd.n942 gnd 0.006084f
C3018 vdd.n943 gnd 0.006084f
C3019 vdd.n944 gnd 0.62173f
C3020 vdd.n945 gnd 0.006084f
C3021 vdd.n946 gnd 0.006084f
C3022 vdd.n947 gnd 0.333723f
C3023 vdd.n948 gnd 0.006084f
C3024 vdd.n949 gnd 0.006084f
C3025 vdd.n950 gnd 0.006084f
C3026 vdd.n951 gnd 0.62173f
C3027 vdd.n952 gnd 0.006084f
C3028 vdd.n953 gnd 0.006084f
C3029 vdd.n954 gnd 0.006084f
C3030 vdd.n955 gnd 0.006084f
C3031 vdd.n956 gnd 0.006084f
C3032 vdd.t165 gnd 0.310865f
C3033 vdd.n957 gnd 0.006084f
C3034 vdd.n958 gnd 0.006084f
C3035 vdd.n959 gnd 0.006084f
C3036 vdd.n960 gnd 0.013026f
C3037 vdd.n961 gnd 0.013026f
C3038 vdd.n962 gnd 0.841164f
C3039 vdd.n963 gnd 0.006084f
C3040 vdd.n964 gnd 0.006084f
C3041 vdd.n965 gnd 0.44344f
C3042 vdd.n966 gnd 0.013026f
C3043 vdd.n967 gnd 0.006084f
C3044 vdd.n968 gnd 0.006084f
C3045 vdd.n969 gnd 11.0997f
C3046 vdd.n1003 gnd 0.013814f
C3047 vdd.n1004 gnd 0.006084f
C3048 vdd.n1005 gnd 0.006084f
C3049 vdd.n1006 gnd 0.005726f
C3050 vdd.n1009 gnd 0.021413f
C3051 vdd.n1010 gnd 0.005977f
C3052 vdd.n1011 gnd 0.007201f
C3053 vdd.n1013 gnd 0.008947f
C3054 vdd.n1014 gnd 0.008947f
C3055 vdd.n1015 gnd 0.007201f
C3056 vdd.n1017 gnd 0.008947f
C3057 vdd.n1018 gnd 0.008947f
C3058 vdd.n1019 gnd 0.008947f
C3059 vdd.n1020 gnd 0.008947f
C3060 vdd.n1021 gnd 0.008947f
C3061 vdd.n1022 gnd 0.007201f
C3062 vdd.n1024 gnd 0.008947f
C3063 vdd.n1025 gnd 0.008947f
C3064 vdd.n1026 gnd 0.008947f
C3065 vdd.n1027 gnd 0.008947f
C3066 vdd.n1028 gnd 0.008947f
C3067 vdd.n1029 gnd 0.007201f
C3068 vdd.n1031 gnd 0.008947f
C3069 vdd.n1032 gnd 0.008947f
C3070 vdd.n1033 gnd 0.008947f
C3071 vdd.n1034 gnd 0.008947f
C3072 vdd.n1035 gnd 0.006013f
C3073 vdd.t174 gnd 0.110068f
C3074 vdd.t173 gnd 0.117632f
C3075 vdd.t172 gnd 0.143747f
C3076 vdd.n1036 gnd 0.184263f
C3077 vdd.n1037 gnd 0.154815f
C3078 vdd.n1039 gnd 0.008947f
C3079 vdd.n1040 gnd 0.008947f
C3080 vdd.n1041 gnd 0.007201f
C3081 vdd.n1042 gnd 0.008947f
C3082 vdd.n1044 gnd 0.008947f
C3083 vdd.n1045 gnd 0.008947f
C3084 vdd.n1046 gnd 0.008947f
C3085 vdd.n1047 gnd 0.008947f
C3086 vdd.n1048 gnd 0.007201f
C3087 vdd.n1050 gnd 0.008947f
C3088 vdd.n1051 gnd 0.008947f
C3089 vdd.n1052 gnd 0.008947f
C3090 vdd.n1053 gnd 0.008947f
C3091 vdd.n1054 gnd 0.008947f
C3092 vdd.n1055 gnd 0.007201f
C3093 vdd.n1057 gnd 0.008947f
C3094 vdd.n1058 gnd 0.008947f
C3095 vdd.n1059 gnd 0.008947f
C3096 vdd.n1060 gnd 0.008947f
C3097 vdd.n1061 gnd 0.008947f
C3098 vdd.n1062 gnd 0.007201f
C3099 vdd.n1064 gnd 0.008947f
C3100 vdd.n1065 gnd 0.008947f
C3101 vdd.n1066 gnd 0.008947f
C3102 vdd.n1067 gnd 0.008947f
C3103 vdd.n1068 gnd 0.008947f
C3104 vdd.n1069 gnd 0.007201f
C3105 vdd.n1071 gnd 0.008947f
C3106 vdd.n1072 gnd 0.008947f
C3107 vdd.n1073 gnd 0.008947f
C3108 vdd.n1074 gnd 0.008947f
C3109 vdd.n1075 gnd 0.007129f
C3110 vdd.t171 gnd 0.110068f
C3111 vdd.t170 gnd 0.117632f
C3112 vdd.t168 gnd 0.143747f
C3113 vdd.n1076 gnd 0.184263f
C3114 vdd.n1077 gnd 0.154815f
C3115 vdd.n1079 gnd 0.008947f
C3116 vdd.n1080 gnd 0.008947f
C3117 vdd.n1081 gnd 0.007201f
C3118 vdd.n1082 gnd 0.008947f
C3119 vdd.n1084 gnd 0.008947f
C3120 vdd.n1085 gnd 0.008947f
C3121 vdd.n1086 gnd 0.008947f
C3122 vdd.n1087 gnd 0.008947f
C3123 vdd.n1088 gnd 0.007201f
C3124 vdd.n1090 gnd 0.008947f
C3125 vdd.n1091 gnd 0.008947f
C3126 vdd.n1092 gnd 0.008947f
C3127 vdd.n1093 gnd 0.008947f
C3128 vdd.n1094 gnd 0.008947f
C3129 vdd.n1095 gnd 0.007201f
C3130 vdd.n1097 gnd 0.008947f
C3131 vdd.n1098 gnd 0.008947f
C3132 vdd.n1099 gnd 0.008947f
C3133 vdd.n1100 gnd 0.008947f
C3134 vdd.n1101 gnd 0.008947f
C3135 vdd.n1102 gnd 0.007201f
C3136 vdd.n1104 gnd 0.008947f
C3137 vdd.n1105 gnd 0.008947f
C3138 vdd.n1106 gnd 0.005726f
C3139 vdd.n1107 gnd 0.007201f
C3140 vdd.n1108 gnd 0.013814f
C3141 vdd.n1109 gnd 0.013814f
C3142 vdd.n1110 gnd 0.006084f
C3143 vdd.n1111 gnd 0.006084f
C3144 vdd.n1112 gnd 0.006084f
C3145 vdd.n1113 gnd 0.006084f
C3146 vdd.n1114 gnd 0.006084f
C3147 vdd.n1115 gnd 0.006084f
C3148 vdd.n1116 gnd 0.006084f
C3149 vdd.n1117 gnd 0.006084f
C3150 vdd.n1118 gnd 0.006084f
C3151 vdd.n1119 gnd 0.006084f
C3152 vdd.n1120 gnd 0.006084f
C3153 vdd.n1121 gnd 0.006084f
C3154 vdd.n1122 gnd 0.006084f
C3155 vdd.n1123 gnd 0.006084f
C3156 vdd.n1124 gnd 0.006084f
C3157 vdd.n1125 gnd 0.006084f
C3158 vdd.n1126 gnd 0.006084f
C3159 vdd.n1127 gnd 0.006084f
C3160 vdd.n1128 gnd 0.006084f
C3161 vdd.n1129 gnd 0.006084f
C3162 vdd.n1130 gnd 0.006084f
C3163 vdd.n1131 gnd 0.006084f
C3164 vdd.n1132 gnd 0.006084f
C3165 vdd.n1133 gnd 0.006084f
C3166 vdd.n1134 gnd 0.006084f
C3167 vdd.n1135 gnd 0.006084f
C3168 vdd.n1136 gnd 0.006084f
C3169 vdd.n1137 gnd 0.006084f
C3170 vdd.n1138 gnd 0.006084f
C3171 vdd.n1139 gnd 0.006084f
C3172 vdd.n1140 gnd 0.006084f
C3173 vdd.n1141 gnd 0.006084f
C3174 vdd.n1142 gnd 0.006084f
C3175 vdd.t166 gnd 0.245843f
C3176 vdd.t167 gnd 0.251651f
C3177 vdd.t164 gnd 0.160496f
C3178 vdd.n1143 gnd 0.086739f
C3179 vdd.n1144 gnd 0.049201f
C3180 vdd.n1145 gnd 0.008695f
C3181 vdd.n1146 gnd 0.006084f
C3182 vdd.t207 gnd 0.245843f
C3183 vdd.t208 gnd 0.251651f
C3184 vdd.t206 gnd 0.160496f
C3185 vdd.n1147 gnd 0.086739f
C3186 vdd.n1148 gnd 0.049201f
C3187 vdd.n1149 gnd 0.006084f
C3188 vdd.n1150 gnd 0.006084f
C3189 vdd.n1151 gnd 0.006084f
C3190 vdd.n1152 gnd 0.006084f
C3191 vdd.n1153 gnd 0.006084f
C3192 vdd.n1154 gnd 0.006084f
C3193 vdd.n1155 gnd 0.006084f
C3194 vdd.n1156 gnd 0.006084f
C3195 vdd.n1157 gnd 0.006084f
C3196 vdd.n1158 gnd 0.006084f
C3197 vdd.n1159 gnd 0.006084f
C3198 vdd.n1160 gnd 0.006084f
C3199 vdd.n1161 gnd 0.006084f
C3200 vdd.n1162 gnd 0.006084f
C3201 vdd.n1163 gnd 0.006084f
C3202 vdd.n1164 gnd 0.006084f
C3203 vdd.n1165 gnd 0.006084f
C3204 vdd.n1166 gnd 0.006084f
C3205 vdd.n1167 gnd 0.006084f
C3206 vdd.n1168 gnd 0.006084f
C3207 vdd.n1169 gnd 0.006084f
C3208 vdd.n1170 gnd 0.006084f
C3209 vdd.n1171 gnd 0.006084f
C3210 vdd.n1172 gnd 0.006084f
C3211 vdd.n1173 gnd 0.006084f
C3212 vdd.n1174 gnd 0.006084f
C3213 vdd.n1175 gnd 0.004429f
C3214 vdd.n1176 gnd 0.008695f
C3215 vdd.n1177 gnd 0.004697f
C3216 vdd.n1178 gnd 0.006084f
C3217 vdd.n1179 gnd 0.006084f
C3218 vdd.n1180 gnd 0.006084f
C3219 vdd.n1181 gnd 0.013814f
C3220 vdd.n1182 gnd 0.013814f
C3221 vdd.n1183 gnd 0.013026f
C3222 vdd.n1184 gnd 0.013026f
C3223 vdd.n1185 gnd 0.006084f
C3224 vdd.n1186 gnd 0.006084f
C3225 vdd.n1187 gnd 0.006084f
C3226 vdd.n1188 gnd 0.006084f
C3227 vdd.n1189 gnd 0.006084f
C3228 vdd.n1190 gnd 0.006084f
C3229 vdd.n1191 gnd 0.006084f
C3230 vdd.n1192 gnd 0.006084f
C3231 vdd.n1193 gnd 0.006084f
C3232 vdd.n1194 gnd 0.006084f
C3233 vdd.n1195 gnd 0.006084f
C3234 vdd.n1196 gnd 0.006084f
C3235 vdd.n1197 gnd 0.006084f
C3236 vdd.n1198 gnd 0.006084f
C3237 vdd.n1199 gnd 0.006084f
C3238 vdd.n1200 gnd 0.006084f
C3239 vdd.n1201 gnd 0.006084f
C3240 vdd.n1202 gnd 0.006084f
C3241 vdd.n1203 gnd 0.006084f
C3242 vdd.n1204 gnd 0.006084f
C3243 vdd.n1205 gnd 0.006084f
C3244 vdd.n1206 gnd 0.006084f
C3245 vdd.n1207 gnd 0.006084f
C3246 vdd.n1208 gnd 0.006084f
C3247 vdd.n1209 gnd 0.006084f
C3248 vdd.n1210 gnd 0.006084f
C3249 vdd.n1211 gnd 0.006084f
C3250 vdd.n1212 gnd 0.006084f
C3251 vdd.n1213 gnd 0.006084f
C3252 vdd.n1214 gnd 0.006084f
C3253 vdd.n1215 gnd 0.006084f
C3254 vdd.n1216 gnd 0.006084f
C3255 vdd.n1217 gnd 0.006084f
C3256 vdd.n1218 gnd 0.006084f
C3257 vdd.n1219 gnd 0.006084f
C3258 vdd.n1220 gnd 0.006084f
C3259 vdd.n1221 gnd 0.006084f
C3260 vdd.n1222 gnd 0.006084f
C3261 vdd.n1223 gnd 0.006084f
C3262 vdd.n1224 gnd 0.006084f
C3263 vdd.n1225 gnd 0.006084f
C3264 vdd.n1226 gnd 0.006084f
C3265 vdd.n1227 gnd 0.370295f
C3266 vdd.n1228 gnd 0.006084f
C3267 vdd.n1229 gnd 0.006084f
C3268 vdd.n1230 gnd 0.006084f
C3269 vdd.n1231 gnd 0.006084f
C3270 vdd.n1232 gnd 0.006084f
C3271 vdd.n1233 gnd 0.006084f
C3272 vdd.n1234 gnd 0.006084f
C3273 vdd.n1235 gnd 0.006084f
C3274 vdd.n1236 gnd 0.006084f
C3275 vdd.n1237 gnd 0.006084f
C3276 vdd.n1238 gnd 0.006084f
C3277 vdd.n1239 gnd 0.006084f
C3278 vdd.n1240 gnd 0.006084f
C3279 vdd.n1241 gnd 0.006084f
C3280 vdd.n1242 gnd 0.006084f
C3281 vdd.n1243 gnd 0.006084f
C3282 vdd.n1244 gnd 0.006084f
C3283 vdd.n1245 gnd 0.006084f
C3284 vdd.n1246 gnd 0.006084f
C3285 vdd.n1247 gnd 0.006084f
C3286 vdd.n1248 gnd 0.006084f
C3287 vdd.n1249 gnd 0.006084f
C3288 vdd.n1250 gnd 0.006084f
C3289 vdd.n1251 gnd 0.006084f
C3290 vdd.n1252 gnd 0.006084f
C3291 vdd.n1253 gnd 0.5623f
C3292 vdd.n1254 gnd 0.006084f
C3293 vdd.n1255 gnd 0.006084f
C3294 vdd.n1256 gnd 0.006084f
C3295 vdd.n1257 gnd 0.006084f
C3296 vdd.n1258 gnd 0.006084f
C3297 vdd.n1259 gnd 0.006084f
C3298 vdd.n1260 gnd 0.006084f
C3299 vdd.n1261 gnd 0.006084f
C3300 vdd.n1262 gnd 0.006084f
C3301 vdd.n1263 gnd 0.006084f
C3302 vdd.n1264 gnd 0.006084f
C3303 vdd.n1265 gnd 0.196576f
C3304 vdd.n1266 gnd 0.006084f
C3305 vdd.n1267 gnd 0.006084f
C3306 vdd.n1268 gnd 0.006084f
C3307 vdd.n1269 gnd 0.006084f
C3308 vdd.n1270 gnd 0.006084f
C3309 vdd.n1271 gnd 0.006084f
C3310 vdd.n1272 gnd 0.006084f
C3311 vdd.n1273 gnd 0.006084f
C3312 vdd.n1274 gnd 0.006084f
C3313 vdd.n1275 gnd 0.006084f
C3314 vdd.n1276 gnd 0.006084f
C3315 vdd.n1277 gnd 0.006084f
C3316 vdd.n1278 gnd 0.006084f
C3317 vdd.n1279 gnd 0.006084f
C3318 vdd.n1280 gnd 0.006084f
C3319 vdd.n1281 gnd 0.006084f
C3320 vdd.n1282 gnd 0.006084f
C3321 vdd.n1283 gnd 0.006084f
C3322 vdd.n1284 gnd 0.006084f
C3323 vdd.n1285 gnd 0.006084f
C3324 vdd.n1286 gnd 0.006084f
C3325 vdd.n1287 gnd 0.006084f
C3326 vdd.n1288 gnd 0.006084f
C3327 vdd.n1289 gnd 0.006084f
C3328 vdd.n1290 gnd 0.006084f
C3329 vdd.n1291 gnd 0.006084f
C3330 vdd.n1292 gnd 0.006084f
C3331 vdd.n1293 gnd 0.006084f
C3332 vdd.n1294 gnd 0.006084f
C3333 vdd.n1295 gnd 0.006084f
C3334 vdd.n1296 gnd 0.006084f
C3335 vdd.n1297 gnd 0.006084f
C3336 vdd.n1298 gnd 0.006084f
C3337 vdd.n1299 gnd 0.006084f
C3338 vdd.n1300 gnd 0.006084f
C3339 vdd.n1301 gnd 0.006084f
C3340 vdd.n1302 gnd 0.006084f
C3341 vdd.n1303 gnd 0.006084f
C3342 vdd.n1304 gnd 0.006084f
C3343 vdd.n1305 gnd 0.006084f
C3344 vdd.n1306 gnd 0.006084f
C3345 vdd.n1307 gnd 0.006084f
C3346 vdd.n1308 gnd 0.013026f
C3347 vdd.n1309 gnd 0.013026f
C3348 vdd.n1310 gnd 0.013814f
C3349 vdd.n1311 gnd 0.006084f
C3350 vdd.n1312 gnd 0.006084f
C3351 vdd.n1313 gnd 0.004697f
C3352 vdd.n1314 gnd 0.006084f
C3353 vdd.n1315 gnd 0.006084f
C3354 vdd.n1316 gnd 0.004429f
C3355 vdd.n1317 gnd 0.006084f
C3356 vdd.n1318 gnd 0.006084f
C3357 vdd.n1319 gnd 0.006084f
C3358 vdd.n1320 gnd 0.006084f
C3359 vdd.n1321 gnd 0.006084f
C3360 vdd.n1322 gnd 0.006084f
C3361 vdd.n1323 gnd 0.006084f
C3362 vdd.n1324 gnd 0.006084f
C3363 vdd.n1325 gnd 0.006084f
C3364 vdd.n1326 gnd 0.006084f
C3365 vdd.n1327 gnd 0.006084f
C3366 vdd.n1328 gnd 0.006084f
C3367 vdd.n1329 gnd 0.006084f
C3368 vdd.n1330 gnd 0.006084f
C3369 vdd.n1331 gnd 0.006084f
C3370 vdd.n1332 gnd 0.006084f
C3371 vdd.n1333 gnd 0.006084f
C3372 vdd.n1334 gnd 0.006084f
C3373 vdd.n1335 gnd 0.006084f
C3374 vdd.n1336 gnd 0.006084f
C3375 vdd.n1337 gnd 0.006084f
C3376 vdd.n1338 gnd 0.006084f
C3377 vdd.n1339 gnd 0.006084f
C3378 vdd.n1340 gnd 0.006084f
C3379 vdd.n1341 gnd 0.006084f
C3380 vdd.n1342 gnd 0.006084f
C3381 vdd.n1343 gnd 0.040983f
C3382 vdd.n1345 gnd 0.021413f
C3383 vdd.n1346 gnd 0.007201f
C3384 vdd.n1348 gnd 0.008947f
C3385 vdd.n1349 gnd 0.007201f
C3386 vdd.n1350 gnd 0.008947f
C3387 vdd.n1352 gnd 0.008947f
C3388 vdd.n1353 gnd 0.008947f
C3389 vdd.n1355 gnd 0.008947f
C3390 vdd.n1356 gnd 0.005977f
C3391 vdd.t169 gnd 0.457154f
C3392 vdd.n1357 gnd 0.008947f
C3393 vdd.n1358 gnd 0.021413f
C3394 vdd.n1359 gnd 0.007201f
C3395 vdd.n1360 gnd 0.008947f
C3396 vdd.n1361 gnd 0.007201f
C3397 vdd.n1362 gnd 0.008947f
C3398 vdd.n1363 gnd 0.914309f
C3399 vdd.n1364 gnd 0.008947f
C3400 vdd.n1365 gnd 0.007201f
C3401 vdd.n1366 gnd 0.007201f
C3402 vdd.n1367 gnd 0.008947f
C3403 vdd.n1368 gnd 0.007201f
C3404 vdd.n1369 gnd 0.008947f
C3405 vdd.t89 gnd 0.457154f
C3406 vdd.n1370 gnd 0.008947f
C3407 vdd.n1371 gnd 0.007201f
C3408 vdd.n1372 gnd 0.008947f
C3409 vdd.n1373 gnd 0.007201f
C3410 vdd.n1374 gnd 0.008947f
C3411 vdd.t119 gnd 0.457154f
C3412 vdd.n1375 gnd 0.008947f
C3413 vdd.n1376 gnd 0.007201f
C3414 vdd.n1377 gnd 0.008947f
C3415 vdd.n1378 gnd 0.007201f
C3416 vdd.n1379 gnd 0.008947f
C3417 vdd.t121 gnd 0.457154f
C3418 vdd.n1380 gnd 0.717732f
C3419 vdd.n1381 gnd 0.008947f
C3420 vdd.n1382 gnd 0.007201f
C3421 vdd.n1383 gnd 0.008947f
C3422 vdd.n1384 gnd 0.007201f
C3423 vdd.n1385 gnd 0.008947f
C3424 vdd.n1386 gnd 0.644588f
C3425 vdd.n1387 gnd 0.008947f
C3426 vdd.n1388 gnd 0.007201f
C3427 vdd.n1389 gnd 0.008947f
C3428 vdd.n1390 gnd 0.007201f
C3429 vdd.n1391 gnd 0.008947f
C3430 vdd.n1392 gnd 0.489155f
C3431 vdd.t85 gnd 0.457154f
C3432 vdd.n1393 gnd 0.008947f
C3433 vdd.n1394 gnd 0.007201f
C3434 vdd.n1395 gnd 0.008916f
C3435 vdd.n1396 gnd 0.007201f
C3436 vdd.n1397 gnd 0.008947f
C3437 vdd.t62 gnd 0.457154f
C3438 vdd.n1398 gnd 0.008947f
C3439 vdd.n1399 gnd 0.007201f
C3440 vdd.n1400 gnd 0.008947f
C3441 vdd.n1401 gnd 0.007201f
C3442 vdd.n1402 gnd 0.008947f
C3443 vdd.t66 gnd 0.457154f
C3444 vdd.n1403 gnd 0.580586f
C3445 vdd.n1404 gnd 0.008947f
C3446 vdd.n1405 gnd 0.007201f
C3447 vdd.n1406 gnd 0.008947f
C3448 vdd.n1407 gnd 0.007201f
C3449 vdd.n1408 gnd 0.008947f
C3450 vdd.t102 gnd 0.457154f
C3451 vdd.n1409 gnd 0.008947f
C3452 vdd.n1410 gnd 0.007201f
C3453 vdd.n1411 gnd 0.008947f
C3454 vdd.n1412 gnd 0.007201f
C3455 vdd.n1413 gnd 0.008947f
C3456 vdd.n1414 gnd 0.626301f
C3457 vdd.n1415 gnd 0.758876f
C3458 vdd.t117 gnd 0.457154f
C3459 vdd.n1416 gnd 0.008947f
C3460 vdd.n1417 gnd 0.007201f
C3461 vdd.n1418 gnd 0.008947f
C3462 vdd.n1419 gnd 0.007201f
C3463 vdd.n1420 gnd 0.008947f
C3464 vdd.n1421 gnd 0.470869f
C3465 vdd.n1422 gnd 0.008947f
C3466 vdd.n1423 gnd 0.007201f
C3467 vdd.n1424 gnd 0.008947f
C3468 vdd.n1425 gnd 0.007201f
C3469 vdd.n1426 gnd 0.008947f
C3470 vdd.n1427 gnd 0.914309f
C3471 vdd.t94 gnd 0.457154f
C3472 vdd.n1428 gnd 0.008947f
C3473 vdd.n1429 gnd 0.007201f
C3474 vdd.n1430 gnd 0.008947f
C3475 vdd.n1431 gnd 0.007201f
C3476 vdd.n1432 gnd 0.008947f
C3477 vdd.t197 gnd 0.457154f
C3478 vdd.n1433 gnd 0.008947f
C3479 vdd.n1434 gnd 0.007201f
C3480 vdd.n1435 gnd 0.021413f
C3481 vdd.n1436 gnd 0.021413f
C3482 vdd.n1437 gnd 2.10291f
C3483 vdd.n1438 gnd 0.516584f
C3484 vdd.n1439 gnd 0.021413f
C3485 vdd.n1440 gnd 0.008947f
C3486 vdd.n1442 gnd 0.008947f
C3487 vdd.n1443 gnd 0.008947f
C3488 vdd.n1444 gnd 0.007201f
C3489 vdd.n1445 gnd 0.008947f
C3490 vdd.n1446 gnd 0.008947f
C3491 vdd.n1448 gnd 0.008947f
C3492 vdd.n1449 gnd 0.008947f
C3493 vdd.n1451 gnd 0.008947f
C3494 vdd.n1452 gnd 0.007201f
C3495 vdd.n1453 gnd 0.008947f
C3496 vdd.n1454 gnd 0.008947f
C3497 vdd.n1456 gnd 0.008947f
C3498 vdd.n1457 gnd 0.008947f
C3499 vdd.n1459 gnd 0.008947f
C3500 vdd.n1460 gnd 0.007201f
C3501 vdd.n1461 gnd 0.008947f
C3502 vdd.n1462 gnd 0.008947f
C3503 vdd.n1464 gnd 0.008947f
C3504 vdd.n1465 gnd 0.008947f
C3505 vdd.n1467 gnd 0.008947f
C3506 vdd.n1468 gnd 0.007201f
C3507 vdd.n1469 gnd 0.008947f
C3508 vdd.n1470 gnd 0.008947f
C3509 vdd.n1472 gnd 0.008947f
C3510 vdd.n1473 gnd 0.008947f
C3511 vdd.n1475 gnd 0.008947f
C3512 vdd.t231 gnd 0.110068f
C3513 vdd.t232 gnd 0.117632f
C3514 vdd.t230 gnd 0.143747f
C3515 vdd.n1476 gnd 0.184263f
C3516 vdd.n1477 gnd 0.155535f
C3517 vdd.n1478 gnd 0.01541f
C3518 vdd.n1479 gnd 0.008947f
C3519 vdd.n1480 gnd 0.008947f
C3520 vdd.n1482 gnd 0.008947f
C3521 vdd.n1483 gnd 0.008947f
C3522 vdd.n1485 gnd 0.008947f
C3523 vdd.n1486 gnd 0.007201f
C3524 vdd.n1487 gnd 0.008947f
C3525 vdd.n1488 gnd 0.008947f
C3526 vdd.n1490 gnd 0.008947f
C3527 vdd.n1491 gnd 0.008947f
C3528 vdd.n1493 gnd 0.008947f
C3529 vdd.n1494 gnd 0.007201f
C3530 vdd.n1495 gnd 0.008947f
C3531 vdd.n1496 gnd 0.008947f
C3532 vdd.n1498 gnd 0.008947f
C3533 vdd.n1499 gnd 0.008947f
C3534 vdd.n1501 gnd 0.008947f
C3535 vdd.n1502 gnd 0.007201f
C3536 vdd.n1503 gnd 0.008947f
C3537 vdd.n1504 gnd 0.008947f
C3538 vdd.n1506 gnd 0.008947f
C3539 vdd.n1507 gnd 0.008947f
C3540 vdd.n1509 gnd 0.008947f
C3541 vdd.n1510 gnd 0.007201f
C3542 vdd.n1511 gnd 0.008947f
C3543 vdd.n1512 gnd 0.008947f
C3544 vdd.n1514 gnd 0.008947f
C3545 vdd.n1515 gnd 0.008947f
C3546 vdd.n1517 gnd 0.008947f
C3547 vdd.n1518 gnd 0.007201f
C3548 vdd.n1519 gnd 0.008947f
C3549 vdd.n1520 gnd 0.008947f
C3550 vdd.n1522 gnd 0.008947f
C3551 vdd.n1523 gnd 0.007129f
C3552 vdd.n1525 gnd 0.007201f
C3553 vdd.n1526 gnd 0.008947f
C3554 vdd.n1527 gnd 0.008947f
C3555 vdd.n1528 gnd 0.008947f
C3556 vdd.n1529 gnd 0.008947f
C3557 vdd.n1531 gnd 0.008947f
C3558 vdd.n1532 gnd 0.008947f
C3559 vdd.n1533 gnd 0.007201f
C3560 vdd.n1534 gnd 0.008947f
C3561 vdd.n1536 gnd 0.008947f
C3562 vdd.n1537 gnd 0.008947f
C3563 vdd.n1539 gnd 0.008947f
C3564 vdd.n1540 gnd 0.008947f
C3565 vdd.n1541 gnd 0.007201f
C3566 vdd.n1542 gnd 0.008947f
C3567 vdd.n1544 gnd 0.008947f
C3568 vdd.n1545 gnd 0.008947f
C3569 vdd.n1547 gnd 0.008947f
C3570 vdd.n1548 gnd 0.008947f
C3571 vdd.n1549 gnd 0.007201f
C3572 vdd.n1550 gnd 0.008947f
C3573 vdd.n1552 gnd 0.008947f
C3574 vdd.n1553 gnd 0.008947f
C3575 vdd.n1555 gnd 0.008947f
C3576 vdd.n1556 gnd 0.008947f
C3577 vdd.n1557 gnd 0.007201f
C3578 vdd.n1558 gnd 0.008947f
C3579 vdd.n1560 gnd 0.008947f
C3580 vdd.n1561 gnd 0.008947f
C3581 vdd.n1563 gnd 0.008947f
C3582 vdd.n1564 gnd 0.00342f
C3583 vdd.t198 gnd 0.110068f
C3584 vdd.t199 gnd 0.117632f
C3585 vdd.t196 gnd 0.143747f
C3586 vdd.n1565 gnd 0.184263f
C3587 vdd.n1566 gnd 0.155535f
C3588 vdd.n1567 gnd 0.01181f
C3589 vdd.n1568 gnd 0.003781f
C3590 vdd.n1569 gnd 0.007201f
C3591 vdd.n1570 gnd 0.008947f
C3592 vdd.n1571 gnd 0.008947f
C3593 vdd.n1572 gnd 0.008947f
C3594 vdd.n1573 gnd 0.007201f
C3595 vdd.n1574 gnd 0.007201f
C3596 vdd.n1575 gnd 0.007201f
C3597 vdd.n1576 gnd 0.008947f
C3598 vdd.n1577 gnd 0.008947f
C3599 vdd.n1578 gnd 0.008947f
C3600 vdd.n1579 gnd 0.007201f
C3601 vdd.n1580 gnd 0.007201f
C3602 vdd.n1581 gnd 0.007201f
C3603 vdd.n1582 gnd 0.008947f
C3604 vdd.n1583 gnd 0.008947f
C3605 vdd.n1584 gnd 0.008947f
C3606 vdd.n1585 gnd 0.007201f
C3607 vdd.n1586 gnd 0.007201f
C3608 vdd.n1587 gnd 0.007201f
C3609 vdd.n1588 gnd 0.008947f
C3610 vdd.n1589 gnd 0.008947f
C3611 vdd.n1590 gnd 0.008947f
C3612 vdd.n1591 gnd 0.007201f
C3613 vdd.n1592 gnd 0.007201f
C3614 vdd.n1593 gnd 0.007201f
C3615 vdd.n1594 gnd 0.008947f
C3616 vdd.n1595 gnd 0.008947f
C3617 vdd.n1596 gnd 0.008947f
C3618 vdd.n1597 gnd 0.007201f
C3619 vdd.n1598 gnd 0.008947f
C3620 vdd.n1599 gnd 0.008947f
C3621 vdd.n1601 gnd 0.008947f
C3622 vdd.t221 gnd 0.110068f
C3623 vdd.t222 gnd 0.117632f
C3624 vdd.t220 gnd 0.143747f
C3625 vdd.n1602 gnd 0.184263f
C3626 vdd.n1603 gnd 0.155535f
C3627 vdd.n1604 gnd 0.01541f
C3628 vdd.n1605 gnd 0.004897f
C3629 vdd.n1606 gnd 0.008947f
C3630 vdd.n1607 gnd 0.008947f
C3631 vdd.n1608 gnd 0.008947f
C3632 vdd.n1609 gnd 0.007201f
C3633 vdd.n1610 gnd 0.007201f
C3634 vdd.n1611 gnd 0.007201f
C3635 vdd.n1612 gnd 0.008947f
C3636 vdd.n1613 gnd 0.008947f
C3637 vdd.n1614 gnd 0.008947f
C3638 vdd.n1615 gnd 0.007201f
C3639 vdd.n1616 gnd 0.007201f
C3640 vdd.n1617 gnd 0.007201f
C3641 vdd.n1618 gnd 0.008947f
C3642 vdd.n1619 gnd 0.008947f
C3643 vdd.n1620 gnd 0.008947f
C3644 vdd.n1621 gnd 0.007201f
C3645 vdd.n1622 gnd 0.007201f
C3646 vdd.n1623 gnd 0.007201f
C3647 vdd.n1624 gnd 0.008947f
C3648 vdd.n1625 gnd 0.008947f
C3649 vdd.n1626 gnd 0.008947f
C3650 vdd.n1627 gnd 0.007201f
C3651 vdd.n1628 gnd 0.007201f
C3652 vdd.n1629 gnd 0.007201f
C3653 vdd.n1630 gnd 0.008947f
C3654 vdd.n1631 gnd 0.008947f
C3655 vdd.n1632 gnd 0.008947f
C3656 vdd.n1633 gnd 0.007201f
C3657 vdd.n1634 gnd 0.007201f
C3658 vdd.n1635 gnd 0.006013f
C3659 vdd.n1636 gnd 0.008947f
C3660 vdd.n1637 gnd 0.008947f
C3661 vdd.n1638 gnd 0.008947f
C3662 vdd.n1639 gnd 0.006013f
C3663 vdd.n1640 gnd 0.007201f
C3664 vdd.n1641 gnd 0.007201f
C3665 vdd.n1642 gnd 0.008947f
C3666 vdd.n1643 gnd 0.008947f
C3667 vdd.n1644 gnd 0.008947f
C3668 vdd.n1645 gnd 0.007201f
C3669 vdd.n1646 gnd 0.007201f
C3670 vdd.n1647 gnd 0.007201f
C3671 vdd.n1648 gnd 0.008947f
C3672 vdd.n1649 gnd 0.008947f
C3673 vdd.n1650 gnd 0.008947f
C3674 vdd.n1651 gnd 0.007201f
C3675 vdd.n1652 gnd 0.007201f
C3676 vdd.n1653 gnd 0.007201f
C3677 vdd.n1654 gnd 0.008947f
C3678 vdd.n1655 gnd 0.008947f
C3679 vdd.n1656 gnd 0.008947f
C3680 vdd.n1657 gnd 0.007201f
C3681 vdd.n1658 gnd 0.007201f
C3682 vdd.n1659 gnd 0.007201f
C3683 vdd.n1660 gnd 0.008947f
C3684 vdd.n1661 gnd 0.008947f
C3685 vdd.n1662 gnd 0.008947f
C3686 vdd.n1663 gnd 0.007201f
C3687 vdd.n1664 gnd 0.007201f
C3688 vdd.n1665 gnd 0.005977f
C3689 vdd.n1666 gnd 0.021413f
C3690 vdd.n1667 gnd 0.021084f
C3691 vdd.n1668 gnd 0.005977f
C3692 vdd.n1669 gnd 0.021084f
C3693 vdd.n1670 gnd 1.28918f
C3694 vdd.n1671 gnd 0.021084f
C3695 vdd.n1672 gnd 0.005977f
C3696 vdd.n1673 gnd 0.021084f
C3697 vdd.n1674 gnd 0.008947f
C3698 vdd.n1675 gnd 0.008947f
C3699 vdd.n1676 gnd 0.007201f
C3700 vdd.n1677 gnd 0.008947f
C3701 vdd.n1678 gnd 0.854879f
C3702 vdd.n1679 gnd 0.008947f
C3703 vdd.n1680 gnd 0.007201f
C3704 vdd.n1681 gnd 0.008947f
C3705 vdd.n1682 gnd 0.008947f
C3706 vdd.n1683 gnd 0.008947f
C3707 vdd.n1684 gnd 0.007201f
C3708 vdd.n1685 gnd 0.008947f
C3709 vdd.n1686 gnd 0.900594f
C3710 vdd.n1687 gnd 0.008947f
C3711 vdd.n1688 gnd 0.007201f
C3712 vdd.n1689 gnd 0.008947f
C3713 vdd.n1690 gnd 0.008947f
C3714 vdd.n1691 gnd 0.008947f
C3715 vdd.n1692 gnd 0.007201f
C3716 vdd.n1693 gnd 0.008947f
C3717 vdd.t60 gnd 0.457154f
C3718 vdd.n1694 gnd 0.745162f
C3719 vdd.n1695 gnd 0.008947f
C3720 vdd.n1696 gnd 0.007201f
C3721 vdd.n1697 gnd 0.008947f
C3722 vdd.n1698 gnd 0.008947f
C3723 vdd.n1699 gnd 0.008947f
C3724 vdd.n1700 gnd 0.007201f
C3725 vdd.n1701 gnd 0.008947f
C3726 vdd.n1702 gnd 0.589729f
C3727 vdd.n1703 gnd 0.008947f
C3728 vdd.n1704 gnd 0.007201f
C3729 vdd.n1705 gnd 0.008947f
C3730 vdd.n1706 gnd 0.008947f
C3731 vdd.n1707 gnd 0.008947f
C3732 vdd.n1708 gnd 0.007201f
C3733 vdd.n1709 gnd 0.008947f
C3734 vdd.n1710 gnd 0.736018f
C3735 vdd.n1711 gnd 0.480012f
C3736 vdd.n1712 gnd 0.008947f
C3737 vdd.n1713 gnd 0.007201f
C3738 vdd.n1714 gnd 0.008947f
C3739 vdd.n1715 gnd 0.008947f
C3740 vdd.n1716 gnd 0.008947f
C3741 vdd.n1717 gnd 0.007201f
C3742 vdd.n1718 gnd 0.008947f
C3743 vdd.n1719 gnd 0.635445f
C3744 vdd.n1720 gnd 0.008947f
C3745 vdd.n1721 gnd 0.007201f
C3746 vdd.n1722 gnd 0.008947f
C3747 vdd.n1723 gnd 0.008947f
C3748 vdd.n1724 gnd 0.008947f
C3749 vdd.n1725 gnd 0.007201f
C3750 vdd.n1726 gnd 0.008947f
C3751 vdd.t87 gnd 0.457154f
C3752 vdd.n1727 gnd 0.758876f
C3753 vdd.n1728 gnd 0.008947f
C3754 vdd.n1729 gnd 0.007201f
C3755 vdd.n1730 gnd 0.00491f
C3756 vdd.n1731 gnd 0.004556f
C3757 vdd.n1732 gnd 0.00252f
C3758 vdd.n1733 gnd 0.005787f
C3759 vdd.n1734 gnd 0.002448f
C3760 vdd.n1735 gnd 0.002592f
C3761 vdd.n1736 gnd 0.004556f
C3762 vdd.n1737 gnd 0.002448f
C3763 vdd.n1738 gnd 0.005787f
C3764 vdd.n1739 gnd 0.002592f
C3765 vdd.n1740 gnd 0.004556f
C3766 vdd.n1741 gnd 0.002448f
C3767 vdd.n1742 gnd 0.00434f
C3768 vdd.n1743 gnd 0.004353f
C3769 vdd.t114 gnd 0.012433f
C3770 vdd.n1744 gnd 0.027663f
C3771 vdd.n1745 gnd 0.143964f
C3772 vdd.n1746 gnd 0.002448f
C3773 vdd.n1747 gnd 0.002592f
C3774 vdd.n1748 gnd 0.005787f
C3775 vdd.n1749 gnd 0.005787f
C3776 vdd.n1750 gnd 0.002592f
C3777 vdd.n1751 gnd 0.002448f
C3778 vdd.n1752 gnd 0.004556f
C3779 vdd.n1753 gnd 0.004556f
C3780 vdd.n1754 gnd 0.002448f
C3781 vdd.n1755 gnd 0.002592f
C3782 vdd.n1756 gnd 0.005787f
C3783 vdd.n1757 gnd 0.005787f
C3784 vdd.n1758 gnd 0.002592f
C3785 vdd.n1759 gnd 0.002448f
C3786 vdd.n1760 gnd 0.004556f
C3787 vdd.n1761 gnd 0.004556f
C3788 vdd.n1762 gnd 0.002448f
C3789 vdd.n1763 gnd 0.002592f
C3790 vdd.n1764 gnd 0.005787f
C3791 vdd.n1765 gnd 0.005787f
C3792 vdd.n1766 gnd 0.013682f
C3793 vdd.n1767 gnd 0.00252f
C3794 vdd.n1768 gnd 0.002448f
C3795 vdd.n1769 gnd 0.011777f
C3796 vdd.n1770 gnd 0.008222f
C3797 vdd.t145 gnd 0.028804f
C3798 vdd.t155 gnd 0.028804f
C3799 vdd.n1771 gnd 0.197961f
C3800 vdd.n1772 gnd 0.155666f
C3801 vdd.t130 gnd 0.028804f
C3802 vdd.t79 gnd 0.028804f
C3803 vdd.n1773 gnd 0.197961f
C3804 vdd.n1774 gnd 0.125622f
C3805 vdd.t123 gnd 0.028804f
C3806 vdd.t88 gnd 0.028804f
C3807 vdd.n1775 gnd 0.197961f
C3808 vdd.n1776 gnd 0.125622f
C3809 vdd.t149 gnd 0.028804f
C3810 vdd.t106 gnd 0.028804f
C3811 vdd.n1777 gnd 0.197961f
C3812 vdd.n1778 gnd 0.125622f
C3813 vdd.t136 gnd 0.028804f
C3814 vdd.t118 gnd 0.028804f
C3815 vdd.n1779 gnd 0.197961f
C3816 vdd.n1780 gnd 0.125622f
C3817 vdd.n1781 gnd 0.00491f
C3818 vdd.n1782 gnd 0.004556f
C3819 vdd.n1783 gnd 0.00252f
C3820 vdd.n1784 gnd 0.005787f
C3821 vdd.n1785 gnd 0.002448f
C3822 vdd.n1786 gnd 0.002592f
C3823 vdd.n1787 gnd 0.004556f
C3824 vdd.n1788 gnd 0.002448f
C3825 vdd.n1789 gnd 0.005787f
C3826 vdd.n1790 gnd 0.002592f
C3827 vdd.n1791 gnd 0.004556f
C3828 vdd.n1792 gnd 0.002448f
C3829 vdd.n1793 gnd 0.00434f
C3830 vdd.n1794 gnd 0.004353f
C3831 vdd.t96 gnd 0.012433f
C3832 vdd.n1795 gnd 0.027663f
C3833 vdd.n1796 gnd 0.143964f
C3834 vdd.n1797 gnd 0.002448f
C3835 vdd.n1798 gnd 0.002592f
C3836 vdd.n1799 gnd 0.005787f
C3837 vdd.n1800 gnd 0.005787f
C3838 vdd.n1801 gnd 0.002592f
C3839 vdd.n1802 gnd 0.002448f
C3840 vdd.n1803 gnd 0.004556f
C3841 vdd.n1804 gnd 0.004556f
C3842 vdd.n1805 gnd 0.002448f
C3843 vdd.n1806 gnd 0.002592f
C3844 vdd.n1807 gnd 0.005787f
C3845 vdd.n1808 gnd 0.005787f
C3846 vdd.n1809 gnd 0.002592f
C3847 vdd.n1810 gnd 0.002448f
C3848 vdd.n1811 gnd 0.004556f
C3849 vdd.n1812 gnd 0.004556f
C3850 vdd.n1813 gnd 0.002448f
C3851 vdd.n1814 gnd 0.002592f
C3852 vdd.n1815 gnd 0.005787f
C3853 vdd.n1816 gnd 0.005787f
C3854 vdd.n1817 gnd 0.013682f
C3855 vdd.n1818 gnd 0.00252f
C3856 vdd.n1819 gnd 0.002448f
C3857 vdd.n1820 gnd 0.011777f
C3858 vdd.n1821 gnd 0.007964f
C3859 vdd.n1822 gnd 0.093463f
C3860 vdd.n1823 gnd 0.00491f
C3861 vdd.n1824 gnd 0.004556f
C3862 vdd.n1825 gnd 0.00252f
C3863 vdd.n1826 gnd 0.005787f
C3864 vdd.n1827 gnd 0.002448f
C3865 vdd.n1828 gnd 0.002592f
C3866 vdd.n1829 gnd 0.004556f
C3867 vdd.n1830 gnd 0.002448f
C3868 vdd.n1831 gnd 0.005787f
C3869 vdd.n1832 gnd 0.002592f
C3870 vdd.n1833 gnd 0.004556f
C3871 vdd.n1834 gnd 0.002448f
C3872 vdd.n1835 gnd 0.00434f
C3873 vdd.n1836 gnd 0.004353f
C3874 vdd.t90 gnd 0.012433f
C3875 vdd.n1837 gnd 0.027663f
C3876 vdd.n1838 gnd 0.143964f
C3877 vdd.n1839 gnd 0.002448f
C3878 vdd.n1840 gnd 0.002592f
C3879 vdd.n1841 gnd 0.005787f
C3880 vdd.n1842 gnd 0.005787f
C3881 vdd.n1843 gnd 0.002592f
C3882 vdd.n1844 gnd 0.002448f
C3883 vdd.n1845 gnd 0.004556f
C3884 vdd.n1846 gnd 0.004556f
C3885 vdd.n1847 gnd 0.002448f
C3886 vdd.n1848 gnd 0.002592f
C3887 vdd.n1849 gnd 0.005787f
C3888 vdd.n1850 gnd 0.005787f
C3889 vdd.n1851 gnd 0.002592f
C3890 vdd.n1852 gnd 0.002448f
C3891 vdd.n1853 gnd 0.004556f
C3892 vdd.n1854 gnd 0.004556f
C3893 vdd.n1855 gnd 0.002448f
C3894 vdd.n1856 gnd 0.002592f
C3895 vdd.n1857 gnd 0.005787f
C3896 vdd.n1858 gnd 0.005787f
C3897 vdd.n1859 gnd 0.013682f
C3898 vdd.n1860 gnd 0.00252f
C3899 vdd.n1861 gnd 0.002448f
C3900 vdd.n1862 gnd 0.011777f
C3901 vdd.n1863 gnd 0.008222f
C3902 vdd.t122 gnd 0.028804f
C3903 vdd.t120 gnd 0.028804f
C3904 vdd.n1864 gnd 0.197961f
C3905 vdd.n1865 gnd 0.155666f
C3906 vdd.t86 gnd 0.028804f
C3907 vdd.t69 gnd 0.028804f
C3908 vdd.n1866 gnd 0.197961f
C3909 vdd.n1867 gnd 0.125622f
C3910 vdd.t63 gnd 0.028804f
C3911 vdd.t115 gnd 0.028804f
C3912 vdd.n1868 gnd 0.197961f
C3913 vdd.n1869 gnd 0.125622f
C3914 vdd.t103 gnd 0.028804f
C3915 vdd.t67 gnd 0.028804f
C3916 vdd.n1870 gnd 0.197961f
C3917 vdd.n1871 gnd 0.125622f
C3918 vdd.t61 gnd 0.028804f
C3919 vdd.t131 gnd 0.028804f
C3920 vdd.n1872 gnd 0.197961f
C3921 vdd.n1873 gnd 0.125622f
C3922 vdd.n1874 gnd 0.00491f
C3923 vdd.n1875 gnd 0.004556f
C3924 vdd.n1876 gnd 0.00252f
C3925 vdd.n1877 gnd 0.005787f
C3926 vdd.n1878 gnd 0.002448f
C3927 vdd.n1879 gnd 0.002592f
C3928 vdd.n1880 gnd 0.004556f
C3929 vdd.n1881 gnd 0.002448f
C3930 vdd.n1882 gnd 0.005787f
C3931 vdd.n1883 gnd 0.002592f
C3932 vdd.n1884 gnd 0.004556f
C3933 vdd.n1885 gnd 0.002448f
C3934 vdd.n1886 gnd 0.00434f
C3935 vdd.n1887 gnd 0.004353f
C3936 vdd.t95 gnd 0.012433f
C3937 vdd.n1888 gnd 0.027663f
C3938 vdd.n1889 gnd 0.143964f
C3939 vdd.n1890 gnd 0.002448f
C3940 vdd.n1891 gnd 0.002592f
C3941 vdd.n1892 gnd 0.005787f
C3942 vdd.n1893 gnd 0.005787f
C3943 vdd.n1894 gnd 0.002592f
C3944 vdd.n1895 gnd 0.002448f
C3945 vdd.n1896 gnd 0.004556f
C3946 vdd.n1897 gnd 0.004556f
C3947 vdd.n1898 gnd 0.002448f
C3948 vdd.n1899 gnd 0.002592f
C3949 vdd.n1900 gnd 0.005787f
C3950 vdd.n1901 gnd 0.005787f
C3951 vdd.n1902 gnd 0.002592f
C3952 vdd.n1903 gnd 0.002448f
C3953 vdd.n1904 gnd 0.004556f
C3954 vdd.n1905 gnd 0.004556f
C3955 vdd.n1906 gnd 0.002448f
C3956 vdd.n1907 gnd 0.002592f
C3957 vdd.n1908 gnd 0.005787f
C3958 vdd.n1909 gnd 0.005787f
C3959 vdd.n1910 gnd 0.013682f
C3960 vdd.n1911 gnd 0.00252f
C3961 vdd.n1912 gnd 0.002448f
C3962 vdd.n1913 gnd 0.011777f
C3963 vdd.n1914 gnd 0.007964f
C3964 vdd.n1915 gnd 0.055601f
C3965 vdd.n1916 gnd 0.200345f
C3966 vdd.n1917 gnd 0.00491f
C3967 vdd.n1918 gnd 0.004556f
C3968 vdd.n1919 gnd 0.00252f
C3969 vdd.n1920 gnd 0.005787f
C3970 vdd.n1921 gnd 0.002448f
C3971 vdd.n1922 gnd 0.002592f
C3972 vdd.n1923 gnd 0.004556f
C3973 vdd.n1924 gnd 0.002448f
C3974 vdd.n1925 gnd 0.005787f
C3975 vdd.n1926 gnd 0.002592f
C3976 vdd.n1927 gnd 0.004556f
C3977 vdd.n1928 gnd 0.002448f
C3978 vdd.n1929 gnd 0.00434f
C3979 vdd.n1930 gnd 0.004353f
C3980 vdd.t101 gnd 0.012433f
C3981 vdd.n1931 gnd 0.027663f
C3982 vdd.n1932 gnd 0.143964f
C3983 vdd.n1933 gnd 0.002448f
C3984 vdd.n1934 gnd 0.002592f
C3985 vdd.n1935 gnd 0.005787f
C3986 vdd.n1936 gnd 0.005787f
C3987 vdd.n1937 gnd 0.002592f
C3988 vdd.n1938 gnd 0.002448f
C3989 vdd.n1939 gnd 0.004556f
C3990 vdd.n1940 gnd 0.004556f
C3991 vdd.n1941 gnd 0.002448f
C3992 vdd.n1942 gnd 0.002592f
C3993 vdd.n1943 gnd 0.005787f
C3994 vdd.n1944 gnd 0.005787f
C3995 vdd.n1945 gnd 0.002592f
C3996 vdd.n1946 gnd 0.002448f
C3997 vdd.n1947 gnd 0.004556f
C3998 vdd.n1948 gnd 0.004556f
C3999 vdd.n1949 gnd 0.002448f
C4000 vdd.n1950 gnd 0.002592f
C4001 vdd.n1951 gnd 0.005787f
C4002 vdd.n1952 gnd 0.005787f
C4003 vdd.n1953 gnd 0.013682f
C4004 vdd.n1954 gnd 0.00252f
C4005 vdd.n1955 gnd 0.002448f
C4006 vdd.n1956 gnd 0.011777f
C4007 vdd.n1957 gnd 0.008222f
C4008 vdd.t127 gnd 0.028804f
C4009 vdd.t126 gnd 0.028804f
C4010 vdd.n1958 gnd 0.197961f
C4011 vdd.n1959 gnd 0.155666f
C4012 vdd.t100 gnd 0.028804f
C4013 vdd.t82 gnd 0.028804f
C4014 vdd.n1960 gnd 0.197961f
C4015 vdd.n1961 gnd 0.125622f
C4016 vdd.t80 gnd 0.028804f
C4017 vdd.t125 gnd 0.028804f
C4018 vdd.n1962 gnd 0.197961f
C4019 vdd.n1963 gnd 0.125622f
C4020 vdd.t109 gnd 0.028804f
C4021 vdd.t81 gnd 0.028804f
C4022 vdd.n1964 gnd 0.197961f
C4023 vdd.n1965 gnd 0.125622f
C4024 vdd.t76 gnd 0.028804f
C4025 vdd.t138 gnd 0.028804f
C4026 vdd.n1966 gnd 0.197961f
C4027 vdd.n1967 gnd 0.125622f
C4028 vdd.n1968 gnd 0.00491f
C4029 vdd.n1969 gnd 0.004556f
C4030 vdd.n1970 gnd 0.00252f
C4031 vdd.n1971 gnd 0.005787f
C4032 vdd.n1972 gnd 0.002448f
C4033 vdd.n1973 gnd 0.002592f
C4034 vdd.n1974 gnd 0.004556f
C4035 vdd.n1975 gnd 0.002448f
C4036 vdd.n1976 gnd 0.005787f
C4037 vdd.n1977 gnd 0.002592f
C4038 vdd.n1978 gnd 0.004556f
C4039 vdd.n1979 gnd 0.002448f
C4040 vdd.n1980 gnd 0.00434f
C4041 vdd.n1981 gnd 0.004353f
C4042 vdd.t107 gnd 0.012433f
C4043 vdd.n1982 gnd 0.027663f
C4044 vdd.n1983 gnd 0.143964f
C4045 vdd.n1984 gnd 0.002448f
C4046 vdd.n1985 gnd 0.002592f
C4047 vdd.n1986 gnd 0.005787f
C4048 vdd.n1987 gnd 0.005787f
C4049 vdd.n1988 gnd 0.002592f
C4050 vdd.n1989 gnd 0.002448f
C4051 vdd.n1990 gnd 0.004556f
C4052 vdd.n1991 gnd 0.004556f
C4053 vdd.n1992 gnd 0.002448f
C4054 vdd.n1993 gnd 0.002592f
C4055 vdd.n1994 gnd 0.005787f
C4056 vdd.n1995 gnd 0.005787f
C4057 vdd.n1996 gnd 0.002592f
C4058 vdd.n1997 gnd 0.002448f
C4059 vdd.n1998 gnd 0.004556f
C4060 vdd.n1999 gnd 0.004556f
C4061 vdd.n2000 gnd 0.002448f
C4062 vdd.n2001 gnd 0.002592f
C4063 vdd.n2002 gnd 0.005787f
C4064 vdd.n2003 gnd 0.005787f
C4065 vdd.n2004 gnd 0.013682f
C4066 vdd.n2005 gnd 0.00252f
C4067 vdd.n2006 gnd 0.002448f
C4068 vdd.n2007 gnd 0.011777f
C4069 vdd.n2008 gnd 0.007964f
C4070 vdd.n2009 gnd 0.055601f
C4071 vdd.n2010 gnd 0.220186f
C4072 vdd.n2011 gnd 2.30604f
C4073 vdd.n2012 gnd 0.532576f
C4074 vdd.n2013 gnd 0.008916f
C4075 vdd.n2014 gnd 0.008947f
C4076 vdd.n2015 gnd 0.007201f
C4077 vdd.n2016 gnd 0.008947f
C4078 vdd.n2017 gnd 0.726875f
C4079 vdd.n2018 gnd 0.008947f
C4080 vdd.n2019 gnd 0.007201f
C4081 vdd.n2020 gnd 0.008947f
C4082 vdd.n2021 gnd 0.008947f
C4083 vdd.n2022 gnd 0.008947f
C4084 vdd.n2023 gnd 0.007201f
C4085 vdd.n2024 gnd 0.008947f
C4086 vdd.n2025 gnd 0.758876f
C4087 vdd.t68 gnd 0.457154f
C4088 vdd.n2026 gnd 0.571443f
C4089 vdd.n2027 gnd 0.008947f
C4090 vdd.n2028 gnd 0.007201f
C4091 vdd.n2029 gnd 0.008947f
C4092 vdd.n2030 gnd 0.008947f
C4093 vdd.n2031 gnd 0.008947f
C4094 vdd.n2032 gnd 0.007201f
C4095 vdd.n2033 gnd 0.008947f
C4096 vdd.n2034 gnd 0.498298f
C4097 vdd.n2035 gnd 0.008947f
C4098 vdd.n2036 gnd 0.007201f
C4099 vdd.n2037 gnd 0.008947f
C4100 vdd.n2038 gnd 0.008947f
C4101 vdd.n2039 gnd 0.008947f
C4102 vdd.n2040 gnd 0.007201f
C4103 vdd.n2041 gnd 0.008947f
C4104 vdd.n2042 gnd 0.5623f
C4105 vdd.n2043 gnd 0.653731f
C4106 vdd.n2044 gnd 0.008947f
C4107 vdd.n2045 gnd 0.007201f
C4108 vdd.n2046 gnd 0.008947f
C4109 vdd.n2047 gnd 0.008947f
C4110 vdd.n2048 gnd 0.008947f
C4111 vdd.n2049 gnd 0.007201f
C4112 vdd.n2050 gnd 0.008947f
C4113 vdd.n2051 gnd 0.809163f
C4114 vdd.n2052 gnd 0.008947f
C4115 vdd.n2053 gnd 0.007201f
C4116 vdd.n2054 gnd 0.008947f
C4117 vdd.n2055 gnd 0.008947f
C4118 vdd.n2056 gnd 0.021084f
C4119 vdd.n2057 gnd 0.008947f
C4120 vdd.n2058 gnd 0.008947f
C4121 vdd.n2059 gnd 0.007201f
C4122 vdd.n2060 gnd 0.008947f
C4123 vdd.n2061 gnd 0.489155f
C4124 vdd.n2062 gnd 0.914309f
C4125 vdd.n2063 gnd 0.008947f
C4126 vdd.n2064 gnd 0.007201f
C4127 vdd.n2065 gnd 0.008947f
C4128 vdd.n2066 gnd 0.008947f
C4129 vdd.n2067 gnd 0.021084f
C4130 vdd.n2068 gnd 0.005977f
C4131 vdd.n2069 gnd 0.021084f
C4132 vdd.n2070 gnd 1.25717f
C4133 vdd.n2071 gnd 0.021084f
C4134 vdd.n2072 gnd 0.021413f
C4135 vdd.n2073 gnd 0.00342f
C4136 vdd.t192 gnd 0.110068f
C4137 vdd.t191 gnd 0.117632f
C4138 vdd.t190 gnd 0.143747f
C4139 vdd.n2074 gnd 0.184263f
C4140 vdd.n2075 gnd 0.154815f
C4141 vdd.n2076 gnd 0.01109f
C4142 vdd.n2077 gnd 0.003781f
C4143 vdd.n2078 gnd 0.007694f
C4144 vdd.n2079 gnd 0.949782f
C4145 vdd.n2081 gnd 0.007201f
C4146 vdd.n2082 gnd 0.007201f
C4147 vdd.n2083 gnd 0.008947f
C4148 vdd.n2085 gnd 0.008947f
C4149 vdd.n2086 gnd 0.008947f
C4150 vdd.n2087 gnd 0.007201f
C4151 vdd.n2088 gnd 0.007201f
C4152 vdd.n2089 gnd 0.007201f
C4153 vdd.n2090 gnd 0.008947f
C4154 vdd.n2092 gnd 0.008947f
C4155 vdd.n2093 gnd 0.008947f
C4156 vdd.n2094 gnd 0.007201f
C4157 vdd.n2095 gnd 0.007201f
C4158 vdd.n2096 gnd 0.007201f
C4159 vdd.n2097 gnd 0.008947f
C4160 vdd.n2099 gnd 0.008947f
C4161 vdd.n2100 gnd 0.008947f
C4162 vdd.n2101 gnd 0.007201f
C4163 vdd.n2102 gnd 0.007201f
C4164 vdd.n2103 gnd 0.007201f
C4165 vdd.n2104 gnd 0.008947f
C4166 vdd.n2106 gnd 0.008947f
C4167 vdd.n2107 gnd 0.008947f
C4168 vdd.n2108 gnd 0.007201f
C4169 vdd.n2109 gnd 0.008947f
C4170 vdd.n2110 gnd 0.008947f
C4171 vdd.n2111 gnd 0.008947f
C4172 vdd.n2112 gnd 0.01469f
C4173 vdd.n2113 gnd 0.004897f
C4174 vdd.n2114 gnd 0.007201f
C4175 vdd.n2115 gnd 0.008947f
C4176 vdd.n2117 gnd 0.008947f
C4177 vdd.n2118 gnd 0.008947f
C4178 vdd.n2119 gnd 0.007201f
C4179 vdd.n2120 gnd 0.007201f
C4180 vdd.n2121 gnd 0.007201f
C4181 vdd.n2122 gnd 0.008947f
C4182 vdd.n2124 gnd 0.008947f
C4183 vdd.n2125 gnd 0.008947f
C4184 vdd.n2126 gnd 0.007201f
C4185 vdd.n2127 gnd 0.007201f
C4186 vdd.n2128 gnd 0.007201f
C4187 vdd.n2129 gnd 0.008947f
C4188 vdd.n2131 gnd 0.008947f
C4189 vdd.n2132 gnd 0.008947f
C4190 vdd.n2133 gnd 0.007201f
C4191 vdd.n2134 gnd 0.007201f
C4192 vdd.n2135 gnd 0.007201f
C4193 vdd.n2136 gnd 0.008947f
C4194 vdd.n2138 gnd 0.008947f
C4195 vdd.n2139 gnd 0.008947f
C4196 vdd.n2140 gnd 0.007201f
C4197 vdd.n2141 gnd 0.007201f
C4198 vdd.n2142 gnd 0.007201f
C4199 vdd.n2143 gnd 0.008947f
C4200 vdd.n2145 gnd 0.008947f
C4201 vdd.n2146 gnd 0.008947f
C4202 vdd.n2147 gnd 0.007201f
C4203 vdd.n2148 gnd 0.008947f
C4204 vdd.n2149 gnd 0.008947f
C4205 vdd.n2150 gnd 0.008947f
C4206 vdd.n2151 gnd 0.01469f
C4207 vdd.n2152 gnd 0.006013f
C4208 vdd.n2153 gnd 0.007201f
C4209 vdd.n2154 gnd 0.008947f
C4210 vdd.n2156 gnd 0.008947f
C4211 vdd.n2157 gnd 0.008947f
C4212 vdd.n2158 gnd 0.007201f
C4213 vdd.n2159 gnd 0.007201f
C4214 vdd.n2160 gnd 0.007201f
C4215 vdd.n2161 gnd 0.008947f
C4216 vdd.n2163 gnd 0.008947f
C4217 vdd.n2164 gnd 0.008947f
C4218 vdd.n2165 gnd 0.007201f
C4219 vdd.n2166 gnd 0.007201f
C4220 vdd.n2167 gnd 0.007201f
C4221 vdd.n2168 gnd 0.008947f
C4222 vdd.n2170 gnd 0.008947f
C4223 vdd.n2171 gnd 0.008947f
C4224 vdd.n2172 gnd 0.007201f
C4225 vdd.n2173 gnd 0.007201f
C4226 vdd.n2174 gnd 0.007201f
C4227 vdd.n2175 gnd 0.008947f
C4228 vdd.n2177 gnd 0.008947f
C4229 vdd.n2178 gnd 0.007201f
C4230 vdd.n2179 gnd 0.007201f
C4231 vdd.n2180 gnd 0.008947f
C4232 vdd.n2182 gnd 0.008947f
C4233 vdd.n2183 gnd 0.008947f
C4234 vdd.n2184 gnd 0.007201f
C4235 vdd.n2185 gnd 0.007694f
C4236 vdd.n2186 gnd 0.949782f
C4237 vdd.n2187 gnd 0.040983f
C4238 vdd.n2188 gnd 0.006084f
C4239 vdd.n2189 gnd 0.006084f
C4240 vdd.n2190 gnd 0.006084f
C4241 vdd.n2191 gnd 0.006084f
C4242 vdd.n2192 gnd 0.006084f
C4243 vdd.n2193 gnd 0.006084f
C4244 vdd.n2194 gnd 0.006084f
C4245 vdd.n2195 gnd 0.006084f
C4246 vdd.n2196 gnd 0.006084f
C4247 vdd.n2197 gnd 0.006084f
C4248 vdd.n2198 gnd 0.006084f
C4249 vdd.n2199 gnd 0.006084f
C4250 vdd.n2200 gnd 0.006084f
C4251 vdd.n2201 gnd 0.006084f
C4252 vdd.n2202 gnd 0.006084f
C4253 vdd.n2203 gnd 0.006084f
C4254 vdd.n2204 gnd 0.006084f
C4255 vdd.n2205 gnd 0.006084f
C4256 vdd.n2206 gnd 0.006084f
C4257 vdd.n2207 gnd 0.006084f
C4258 vdd.n2208 gnd 0.006084f
C4259 vdd.n2209 gnd 0.006084f
C4260 vdd.n2210 gnd 0.006084f
C4261 vdd.n2211 gnd 0.006084f
C4262 vdd.n2212 gnd 0.006084f
C4263 vdd.n2213 gnd 0.006084f
C4264 vdd.n2214 gnd 0.006084f
C4265 vdd.n2215 gnd 0.006084f
C4266 vdd.n2216 gnd 0.006084f
C4267 vdd.n2217 gnd 0.006084f
C4268 vdd.n2218 gnd 10.797999f
C4269 vdd.n2220 gnd 0.013814f
C4270 vdd.n2221 gnd 0.013814f
C4271 vdd.n2222 gnd 0.013026f
C4272 vdd.n2223 gnd 0.006084f
C4273 vdd.n2224 gnd 0.006084f
C4274 vdd.n2225 gnd 0.62173f
C4275 vdd.n2226 gnd 0.006084f
C4276 vdd.n2227 gnd 0.006084f
C4277 vdd.n2228 gnd 0.006084f
C4278 vdd.n2229 gnd 0.006084f
C4279 vdd.n2230 gnd 0.006084f
C4280 vdd.n2231 gnd 0.489155f
C4281 vdd.n2232 gnd 0.006084f
C4282 vdd.n2233 gnd 0.006084f
C4283 vdd.n2234 gnd 0.006084f
C4284 vdd.n2235 gnd 0.006084f
C4285 vdd.n2236 gnd 0.006084f
C4286 vdd.n2237 gnd 0.62173f
C4287 vdd.n2238 gnd 0.006084f
C4288 vdd.n2239 gnd 0.006084f
C4289 vdd.n2240 gnd 0.006084f
C4290 vdd.n2241 gnd 0.006084f
C4291 vdd.n2242 gnd 0.006084f
C4292 vdd.n2243 gnd 0.62173f
C4293 vdd.n2244 gnd 0.006084f
C4294 vdd.n2245 gnd 0.006084f
C4295 vdd.n2246 gnd 0.006084f
C4296 vdd.n2247 gnd 0.006084f
C4297 vdd.n2248 gnd 0.006084f
C4298 vdd.n2249 gnd 0.598872f
C4299 vdd.n2250 gnd 0.006084f
C4300 vdd.n2251 gnd 0.006084f
C4301 vdd.n2252 gnd 0.006084f
C4302 vdd.n2253 gnd 0.006084f
C4303 vdd.n2254 gnd 0.006084f
C4304 vdd.n2255 gnd 0.461726f
C4305 vdd.n2256 gnd 0.006084f
C4306 vdd.n2257 gnd 0.006084f
C4307 vdd.n2258 gnd 0.006084f
C4308 vdd.n2259 gnd 0.006084f
C4309 vdd.n2260 gnd 0.006084f
C4310 vdd.n2261 gnd 0.32458f
C4311 vdd.n2262 gnd 0.006084f
C4312 vdd.n2263 gnd 0.006084f
C4313 vdd.n2264 gnd 0.006084f
C4314 vdd.n2265 gnd 0.006084f
C4315 vdd.n2266 gnd 0.006084f
C4316 vdd.n2267 gnd 0.434297f
C4317 vdd.n2268 gnd 0.006084f
C4318 vdd.n2269 gnd 0.006084f
C4319 vdd.n2270 gnd 0.006084f
C4320 vdd.n2271 gnd 0.006084f
C4321 vdd.n2272 gnd 0.006084f
C4322 vdd.n2273 gnd 0.571443f
C4323 vdd.n2274 gnd 0.006084f
C4324 vdd.n2275 gnd 0.006084f
C4325 vdd.n2276 gnd 0.006084f
C4326 vdd.n2277 gnd 0.006084f
C4327 vdd.n2278 gnd 0.006084f
C4328 vdd.n2279 gnd 0.62173f
C4329 vdd.n2280 gnd 0.006084f
C4330 vdd.n2281 gnd 0.006084f
C4331 vdd.n2282 gnd 0.006084f
C4332 vdd.n2283 gnd 0.006084f
C4333 vdd.n2284 gnd 0.006084f
C4334 vdd.n2285 gnd 0.534871f
C4335 vdd.n2286 gnd 0.006084f
C4336 vdd.n2287 gnd 0.006084f
C4337 vdd.n2288 gnd 0.004831f
C4338 vdd.n2289 gnd 0.017624f
C4339 vdd.n2290 gnd 0.004294f
C4340 vdd.n2291 gnd 0.006084f
C4341 vdd.n2292 gnd 0.397724f
C4342 vdd.n2293 gnd 0.006084f
C4343 vdd.n2294 gnd 0.006084f
C4344 vdd.n2295 gnd 0.006084f
C4345 vdd.n2296 gnd 0.006084f
C4346 vdd.n2297 gnd 0.006084f
C4347 vdd.n2298 gnd 0.361152f
C4348 vdd.n2299 gnd 0.006084f
C4349 vdd.n2300 gnd 0.006084f
C4350 vdd.n2301 gnd 0.006084f
C4351 vdd.n2302 gnd 0.006084f
C4352 vdd.n2303 gnd 0.006084f
C4353 vdd.n2304 gnd 0.498298f
C4354 vdd.n2305 gnd 0.006084f
C4355 vdd.n2306 gnd 0.006084f
C4356 vdd.n2307 gnd 0.006084f
C4357 vdd.n2308 gnd 0.006084f
C4358 vdd.n2309 gnd 0.006084f
C4359 vdd.n2310 gnd 0.548585f
C4360 vdd.n2311 gnd 0.006084f
C4361 vdd.n2312 gnd 0.006084f
C4362 vdd.n2313 gnd 0.006084f
C4363 vdd.n2314 gnd 0.006084f
C4364 vdd.n2315 gnd 0.006084f
C4365 vdd.n2316 gnd 0.411439f
C4366 vdd.n2317 gnd 0.006084f
C4367 vdd.n2318 gnd 0.006084f
C4368 vdd.n2319 gnd 0.006084f
C4369 vdd.n2320 gnd 0.006084f
C4370 vdd.n2321 gnd 0.006084f
C4371 vdd.n2322 gnd 0.196576f
C4372 vdd.n2323 gnd 0.006084f
C4373 vdd.n2324 gnd 0.006084f
C4374 vdd.n2325 gnd 0.006084f
C4375 vdd.n2326 gnd 0.006084f
C4376 vdd.n2327 gnd 0.006084f
C4377 vdd.n2328 gnd 0.196576f
C4378 vdd.n2329 gnd 0.006084f
C4379 vdd.n2330 gnd 0.006084f
C4380 vdd.n2331 gnd 0.006084f
C4381 vdd.n2332 gnd 0.006084f
C4382 vdd.n2333 gnd 0.006084f
C4383 vdd.n2334 gnd 0.62173f
C4384 vdd.n2335 gnd 0.006084f
C4385 vdd.n2336 gnd 0.006084f
C4386 vdd.n2337 gnd 0.006084f
C4387 vdd.n2338 gnd 0.006084f
C4388 vdd.n2339 gnd 0.006084f
C4389 vdd.n2340 gnd 0.006084f
C4390 vdd.n2341 gnd 0.006084f
C4391 vdd.n2342 gnd 0.429725f
C4392 vdd.n2343 gnd 0.006084f
C4393 vdd.n2344 gnd 0.006084f
C4394 vdd.n2345 gnd 0.006084f
C4395 vdd.n2346 gnd 0.006084f
C4396 vdd.n2347 gnd 0.006084f
C4397 vdd.n2348 gnd 0.006084f
C4398 vdd.n2349 gnd 0.388581f
C4399 vdd.n2350 gnd 0.006084f
C4400 vdd.n2351 gnd 0.006084f
C4401 vdd.n2352 gnd 0.006084f
C4402 vdd.n2353 gnd 0.013814f
C4403 vdd.n2354 gnd 0.013026f
C4404 vdd.n2355 gnd 0.006084f
C4405 vdd.n2356 gnd 0.006084f
C4406 vdd.n2357 gnd 0.004697f
C4407 vdd.n2358 gnd 0.006084f
C4408 vdd.n2359 gnd 0.006084f
C4409 vdd.n2360 gnd 0.004429f
C4410 vdd.n2361 gnd 0.006084f
C4411 vdd.n2362 gnd 0.006084f
C4412 vdd.n2363 gnd 0.006084f
C4413 vdd.n2364 gnd 0.006084f
C4414 vdd.n2365 gnd 0.006084f
C4415 vdd.n2366 gnd 0.006084f
C4416 vdd.n2367 gnd 0.006084f
C4417 vdd.n2368 gnd 0.006084f
C4418 vdd.n2369 gnd 0.006084f
C4419 vdd.n2370 gnd 0.006084f
C4420 vdd.n2371 gnd 0.006084f
C4421 vdd.n2372 gnd 0.006084f
C4422 vdd.n2373 gnd 0.006084f
C4423 vdd.n2374 gnd 0.006084f
C4424 vdd.n2375 gnd 0.006084f
C4425 vdd.n2376 gnd 0.006084f
C4426 vdd.n2377 gnd 0.006084f
C4427 vdd.n2378 gnd 0.006084f
C4428 vdd.n2379 gnd 0.006084f
C4429 vdd.n2380 gnd 0.006084f
C4430 vdd.n2381 gnd 0.006084f
C4431 vdd.n2382 gnd 0.006084f
C4432 vdd.n2383 gnd 0.006084f
C4433 vdd.n2384 gnd 0.006084f
C4434 vdd.n2385 gnd 0.006084f
C4435 vdd.n2386 gnd 0.006084f
C4436 vdd.n2387 gnd 0.006084f
C4437 vdd.n2388 gnd 0.006084f
C4438 vdd.n2389 gnd 0.006084f
C4439 vdd.n2390 gnd 0.006084f
C4440 vdd.n2391 gnd 0.006084f
C4441 vdd.n2392 gnd 0.006084f
C4442 vdd.n2393 gnd 0.006084f
C4443 vdd.n2394 gnd 0.006084f
C4444 vdd.n2395 gnd 0.006084f
C4445 vdd.n2396 gnd 0.006084f
C4446 vdd.n2397 gnd 0.006084f
C4447 vdd.n2398 gnd 0.006084f
C4448 vdd.n2399 gnd 0.006084f
C4449 vdd.n2400 gnd 0.006084f
C4450 vdd.n2401 gnd 0.006084f
C4451 vdd.n2402 gnd 0.006084f
C4452 vdd.n2403 gnd 0.006084f
C4453 vdd.n2404 gnd 0.006084f
C4454 vdd.n2405 gnd 0.006084f
C4455 vdd.n2406 gnd 0.006084f
C4456 vdd.n2407 gnd 0.006084f
C4457 vdd.n2408 gnd 0.006084f
C4458 vdd.n2409 gnd 0.006084f
C4459 vdd.n2410 gnd 0.006084f
C4460 vdd.n2411 gnd 0.006084f
C4461 vdd.n2412 gnd 0.006084f
C4462 vdd.n2413 gnd 0.006084f
C4463 vdd.n2414 gnd 0.006084f
C4464 vdd.n2415 gnd 0.006084f
C4465 vdd.n2416 gnd 0.006084f
C4466 vdd.n2417 gnd 0.006084f
C4467 vdd.n2418 gnd 0.006084f
C4468 vdd.n2419 gnd 0.006084f
C4469 vdd.n2420 gnd 0.006084f
C4470 vdd.n2421 gnd 0.013814f
C4471 vdd.n2422 gnd 0.013026f
C4472 vdd.n2423 gnd 0.013026f
C4473 vdd.n2424 gnd 0.704018f
C4474 vdd.n2425 gnd 0.013026f
C4475 vdd.n2426 gnd 0.013814f
C4476 vdd.n2427 gnd 0.013026f
C4477 vdd.n2428 gnd 0.006084f
C4478 vdd.n2429 gnd 0.006084f
C4479 vdd.n2430 gnd 0.006084f
C4480 vdd.n2431 gnd 0.004697f
C4481 vdd.n2432 gnd 0.008695f
C4482 vdd.n2433 gnd 0.004429f
C4483 vdd.n2434 gnd 0.006084f
C4484 vdd.n2435 gnd 0.006084f
C4485 vdd.n2436 gnd 0.006084f
C4486 vdd.n2437 gnd 0.006084f
C4487 vdd.n2438 gnd 0.006084f
C4488 vdd.n2439 gnd 0.006084f
C4489 vdd.n2440 gnd 0.006084f
C4490 vdd.n2441 gnd 0.006084f
C4491 vdd.n2442 gnd 0.006084f
C4492 vdd.n2443 gnd 0.006084f
C4493 vdd.n2444 gnd 0.006084f
C4494 vdd.n2445 gnd 0.006084f
C4495 vdd.n2446 gnd 0.006084f
C4496 vdd.n2447 gnd 0.006084f
C4497 vdd.n2448 gnd 0.006084f
C4498 vdd.n2449 gnd 0.006084f
C4499 vdd.n2450 gnd 0.006084f
C4500 vdd.n2451 gnd 0.006084f
C4501 vdd.n2452 gnd 0.006084f
C4502 vdd.n2453 gnd 0.006084f
C4503 vdd.n2454 gnd 0.006084f
C4504 vdd.n2455 gnd 0.006084f
C4505 vdd.n2456 gnd 0.006084f
C4506 vdd.n2457 gnd 0.006084f
C4507 vdd.n2458 gnd 0.006084f
C4508 vdd.n2459 gnd 0.006084f
C4509 vdd.n2460 gnd 0.006084f
C4510 vdd.n2461 gnd 0.006084f
C4511 vdd.n2462 gnd 0.006084f
C4512 vdd.n2463 gnd 0.006084f
C4513 vdd.n2464 gnd 0.006084f
C4514 vdd.n2465 gnd 0.006084f
C4515 vdd.n2466 gnd 0.006084f
C4516 vdd.n2467 gnd 0.006084f
C4517 vdd.n2468 gnd 0.006084f
C4518 vdd.n2469 gnd 0.006084f
C4519 vdd.n2470 gnd 0.006084f
C4520 vdd.n2471 gnd 0.006084f
C4521 vdd.n2472 gnd 0.006084f
C4522 vdd.n2473 gnd 0.006084f
C4523 vdd.n2474 gnd 0.006084f
C4524 vdd.n2475 gnd 0.006084f
C4525 vdd.n2476 gnd 0.006084f
C4526 vdd.n2477 gnd 0.006084f
C4527 vdd.n2478 gnd 0.006084f
C4528 vdd.n2479 gnd 0.006084f
C4529 vdd.n2480 gnd 0.006084f
C4530 vdd.n2481 gnd 0.006084f
C4531 vdd.n2482 gnd 0.006084f
C4532 vdd.n2483 gnd 0.006084f
C4533 vdd.n2484 gnd 0.006084f
C4534 vdd.n2485 gnd 0.006084f
C4535 vdd.n2486 gnd 0.006084f
C4536 vdd.n2487 gnd 0.006084f
C4537 vdd.n2488 gnd 0.006084f
C4538 vdd.n2489 gnd 0.006084f
C4539 vdd.n2490 gnd 0.006084f
C4540 vdd.n2491 gnd 0.006084f
C4541 vdd.n2492 gnd 0.006084f
C4542 vdd.n2493 gnd 0.006084f
C4543 vdd.n2494 gnd 0.013814f
C4544 vdd.n2495 gnd 0.013814f
C4545 vdd.n2496 gnd 0.758876f
C4546 vdd.t29 gnd 2.69721f
C4547 vdd.t16 gnd 2.69721f
C4548 vdd.n2530 gnd 0.013814f
C4549 vdd.t34 gnd 0.530299f
C4550 vdd.n2531 gnd 0.006084f
C4551 vdd.t218 gnd 0.245843f
C4552 vdd.t219 gnd 0.251651f
C4553 vdd.t216 gnd 0.160496f
C4554 vdd.n2532 gnd 0.086739f
C4555 vdd.n2533 gnd 0.049201f
C4556 vdd.n2534 gnd 0.006084f
C4557 vdd.t228 gnd 0.245843f
C4558 vdd.t229 gnd 0.251651f
C4559 vdd.t227 gnd 0.160496f
C4560 vdd.n2535 gnd 0.086739f
C4561 vdd.n2536 gnd 0.049201f
C4562 vdd.n2537 gnd 0.008695f
C4563 vdd.n2538 gnd 0.013814f
C4564 vdd.n2539 gnd 0.013814f
C4565 vdd.n2540 gnd 0.006084f
C4566 vdd.n2541 gnd 0.006084f
C4567 vdd.n2542 gnd 0.006084f
C4568 vdd.n2543 gnd 0.006084f
C4569 vdd.n2544 gnd 0.006084f
C4570 vdd.n2545 gnd 0.006084f
C4571 vdd.n2546 gnd 0.006084f
C4572 vdd.n2547 gnd 0.006084f
C4573 vdd.n2548 gnd 0.006084f
C4574 vdd.n2549 gnd 0.006084f
C4575 vdd.n2550 gnd 0.006084f
C4576 vdd.n2551 gnd 0.006084f
C4577 vdd.n2552 gnd 0.006084f
C4578 vdd.n2553 gnd 0.006084f
C4579 vdd.n2554 gnd 0.006084f
C4580 vdd.n2555 gnd 0.006084f
C4581 vdd.n2556 gnd 0.006084f
C4582 vdd.n2557 gnd 0.006084f
C4583 vdd.n2558 gnd 0.006084f
C4584 vdd.n2559 gnd 0.006084f
C4585 vdd.n2560 gnd 0.006084f
C4586 vdd.n2561 gnd 0.006084f
C4587 vdd.n2562 gnd 0.006084f
C4588 vdd.n2563 gnd 0.006084f
C4589 vdd.n2564 gnd 0.006084f
C4590 vdd.n2565 gnd 0.006084f
C4591 vdd.n2566 gnd 0.006084f
C4592 vdd.n2567 gnd 0.006084f
C4593 vdd.n2568 gnd 0.006084f
C4594 vdd.n2569 gnd 0.006084f
C4595 vdd.n2570 gnd 0.006084f
C4596 vdd.n2571 gnd 0.006084f
C4597 vdd.n2572 gnd 0.006084f
C4598 vdd.n2573 gnd 0.006084f
C4599 vdd.n2574 gnd 0.006084f
C4600 vdd.n2575 gnd 0.006084f
C4601 vdd.n2576 gnd 0.006084f
C4602 vdd.n2577 gnd 0.006084f
C4603 vdd.n2578 gnd 0.006084f
C4604 vdd.n2579 gnd 0.006084f
C4605 vdd.n2580 gnd 0.006084f
C4606 vdd.n2581 gnd 0.006084f
C4607 vdd.n2582 gnd 0.006084f
C4608 vdd.n2583 gnd 0.006084f
C4609 vdd.n2584 gnd 0.006084f
C4610 vdd.n2585 gnd 0.006084f
C4611 vdd.n2586 gnd 0.006084f
C4612 vdd.n2587 gnd 0.006084f
C4613 vdd.n2588 gnd 0.006084f
C4614 vdd.n2589 gnd 0.006084f
C4615 vdd.n2590 gnd 0.006084f
C4616 vdd.n2591 gnd 0.006084f
C4617 vdd.n2592 gnd 0.006084f
C4618 vdd.n2593 gnd 0.006084f
C4619 vdd.n2594 gnd 0.006084f
C4620 vdd.n2595 gnd 0.006084f
C4621 vdd.n2596 gnd 0.006084f
C4622 vdd.n2597 gnd 0.006084f
C4623 vdd.n2598 gnd 0.006084f
C4624 vdd.n2599 gnd 0.006084f
C4625 vdd.n2600 gnd 0.004429f
C4626 vdd.n2601 gnd 0.006084f
C4627 vdd.n2602 gnd 0.006084f
C4628 vdd.n2603 gnd 0.004697f
C4629 vdd.n2604 gnd 0.006084f
C4630 vdd.n2605 gnd 0.006084f
C4631 vdd.n2606 gnd 0.013814f
C4632 vdd.n2607 gnd 0.013026f
C4633 vdd.n2608 gnd 0.013026f
C4634 vdd.n2609 gnd 0.006084f
C4635 vdd.n2610 gnd 0.006084f
C4636 vdd.n2611 gnd 0.006084f
C4637 vdd.n2612 gnd 0.006084f
C4638 vdd.n2613 gnd 0.006084f
C4639 vdd.n2614 gnd 0.006084f
C4640 vdd.n2615 gnd 0.006084f
C4641 vdd.n2616 gnd 0.006084f
C4642 vdd.n2617 gnd 0.006084f
C4643 vdd.n2618 gnd 0.006084f
C4644 vdd.n2619 gnd 0.006084f
C4645 vdd.n2620 gnd 0.006084f
C4646 vdd.n2621 gnd 0.006084f
C4647 vdd.n2622 gnd 0.006084f
C4648 vdd.n2623 gnd 0.006084f
C4649 vdd.n2624 gnd 0.006084f
C4650 vdd.n2625 gnd 0.006084f
C4651 vdd.n2626 gnd 0.006084f
C4652 vdd.n2627 gnd 0.006084f
C4653 vdd.n2628 gnd 0.006084f
C4654 vdd.n2629 gnd 0.006084f
C4655 vdd.n2630 gnd 0.006084f
C4656 vdd.n2631 gnd 0.006084f
C4657 vdd.n2632 gnd 0.006084f
C4658 vdd.n2633 gnd 0.006084f
C4659 vdd.n2634 gnd 0.006084f
C4660 vdd.n2635 gnd 0.006084f
C4661 vdd.n2636 gnd 0.006084f
C4662 vdd.n2637 gnd 0.006084f
C4663 vdd.n2638 gnd 0.006084f
C4664 vdd.n2639 gnd 0.006084f
C4665 vdd.n2640 gnd 0.006084f
C4666 vdd.n2641 gnd 0.006084f
C4667 vdd.n2642 gnd 0.006084f
C4668 vdd.n2643 gnd 0.006084f
C4669 vdd.n2644 gnd 0.006084f
C4670 vdd.n2645 gnd 0.006084f
C4671 vdd.n2646 gnd 0.006084f
C4672 vdd.n2647 gnd 0.006084f
C4673 vdd.n2648 gnd 0.006084f
C4674 vdd.n2649 gnd 0.006084f
C4675 vdd.n2650 gnd 0.006084f
C4676 vdd.n2651 gnd 0.006084f
C4677 vdd.n2652 gnd 0.006084f
C4678 vdd.n2653 gnd 0.006084f
C4679 vdd.n2654 gnd 0.006084f
C4680 vdd.n2655 gnd 0.006084f
C4681 vdd.n2656 gnd 0.006084f
C4682 vdd.n2657 gnd 0.006084f
C4683 vdd.n2658 gnd 0.006084f
C4684 vdd.n2659 gnd 0.006084f
C4685 vdd.n2660 gnd 0.006084f
C4686 vdd.n2661 gnd 0.006084f
C4687 vdd.n2662 gnd 0.006084f
C4688 vdd.n2663 gnd 0.006084f
C4689 vdd.n2664 gnd 0.006084f
C4690 vdd.n2665 gnd 0.006084f
C4691 vdd.n2666 gnd 0.006084f
C4692 vdd.n2667 gnd 0.006084f
C4693 vdd.n2668 gnd 0.006084f
C4694 vdd.n2669 gnd 0.006084f
C4695 vdd.n2670 gnd 0.006084f
C4696 vdd.n2671 gnd 0.006084f
C4697 vdd.n2672 gnd 0.006084f
C4698 vdd.n2673 gnd 0.006084f
C4699 vdd.n2674 gnd 0.006084f
C4700 vdd.n2675 gnd 0.006084f
C4701 vdd.n2676 gnd 0.006084f
C4702 vdd.n2677 gnd 0.006084f
C4703 vdd.n2678 gnd 0.006084f
C4704 vdd.n2679 gnd 0.006084f
C4705 vdd.n2680 gnd 0.006084f
C4706 vdd.n2681 gnd 0.006084f
C4707 vdd.n2682 gnd 0.006084f
C4708 vdd.n2683 gnd 0.006084f
C4709 vdd.n2684 gnd 0.006084f
C4710 vdd.n2685 gnd 0.006084f
C4711 vdd.n2686 gnd 0.006084f
C4712 vdd.n2687 gnd 0.006084f
C4713 vdd.n2688 gnd 0.006084f
C4714 vdd.n2689 gnd 0.006084f
C4715 vdd.n2690 gnd 0.006084f
C4716 vdd.n2691 gnd 0.006084f
C4717 vdd.n2692 gnd 0.006084f
C4718 vdd.n2693 gnd 0.006084f
C4719 vdd.n2694 gnd 0.006084f
C4720 vdd.n2695 gnd 0.006084f
C4721 vdd.n2696 gnd 0.006084f
C4722 vdd.n2697 gnd 0.006084f
C4723 vdd.n2698 gnd 0.006084f
C4724 vdd.n2699 gnd 0.006084f
C4725 vdd.n2700 gnd 0.006084f
C4726 vdd.n2701 gnd 0.006084f
C4727 vdd.n2702 gnd 0.006084f
C4728 vdd.n2703 gnd 0.006084f
C4729 vdd.n2704 gnd 0.006084f
C4730 vdd.n2705 gnd 0.006084f
C4731 vdd.n2706 gnd 0.006084f
C4732 vdd.n2707 gnd 0.006084f
C4733 vdd.n2708 gnd 0.006084f
C4734 vdd.n2709 gnd 0.006084f
C4735 vdd.n2710 gnd 0.196576f
C4736 vdd.n2711 gnd 0.006084f
C4737 vdd.n2712 gnd 0.006084f
C4738 vdd.n2713 gnd 0.006084f
C4739 vdd.n2714 gnd 0.006084f
C4740 vdd.n2715 gnd 0.006084f
C4741 vdd.n2716 gnd 0.196576f
C4742 vdd.n2717 gnd 0.006084f
C4743 vdd.n2718 gnd 0.006084f
C4744 vdd.n2719 gnd 0.006084f
C4745 vdd.n2720 gnd 0.006084f
C4746 vdd.n2721 gnd 0.006084f
C4747 vdd.n2722 gnd 0.006084f
C4748 vdd.n2723 gnd 0.006084f
C4749 vdd.n2724 gnd 0.006084f
C4750 vdd.n2725 gnd 0.006084f
C4751 vdd.n2726 gnd 0.006084f
C4752 vdd.n2727 gnd 0.006084f
C4753 vdd.n2728 gnd 0.388581f
C4754 vdd.n2729 gnd 0.006084f
C4755 vdd.n2730 gnd 0.006084f
C4756 vdd.n2731 gnd 0.006084f
C4757 vdd.n2732 gnd 0.013026f
C4758 vdd.n2733 gnd 0.013026f
C4759 vdd.n2734 gnd 0.013814f
C4760 vdd.n2735 gnd 0.013814f
C4761 vdd.n2736 gnd 0.006084f
C4762 vdd.n2737 gnd 0.006084f
C4763 vdd.n2738 gnd 0.006084f
C4764 vdd.n2739 gnd 0.004697f
C4765 vdd.n2740 gnd 0.008695f
C4766 vdd.n2741 gnd 0.004429f
C4767 vdd.n2742 gnd 0.006084f
C4768 vdd.n2743 gnd 0.006084f
C4769 vdd.n2744 gnd 0.006084f
C4770 vdd.n2745 gnd 0.006084f
C4771 vdd.n2746 gnd 0.006084f
C4772 vdd.n2747 gnd 0.006084f
C4773 vdd.n2748 gnd 0.006084f
C4774 vdd.n2749 gnd 0.006084f
C4775 vdd.n2750 gnd 0.006084f
C4776 vdd.n2751 gnd 0.006084f
C4777 vdd.n2752 gnd 0.006084f
C4778 vdd.n2753 gnd 0.006084f
C4779 vdd.n2754 gnd 0.006084f
C4780 vdd.n2755 gnd 0.006084f
C4781 vdd.n2756 gnd 0.006084f
C4782 vdd.n2757 gnd 0.006084f
C4783 vdd.n2758 gnd 0.006084f
C4784 vdd.n2759 gnd 0.006084f
C4785 vdd.n2760 gnd 0.006084f
C4786 vdd.n2761 gnd 0.006084f
C4787 vdd.n2762 gnd 0.006084f
C4788 vdd.n2763 gnd 0.006084f
C4789 vdd.n2764 gnd 0.006084f
C4790 vdd.n2765 gnd 0.006084f
C4791 vdd.n2766 gnd 0.006084f
C4792 vdd.n2767 gnd 0.006084f
C4793 vdd.n2768 gnd 0.006084f
C4794 vdd.n2769 gnd 0.006084f
C4795 vdd.n2770 gnd 0.006084f
C4796 vdd.n2771 gnd 0.006084f
C4797 vdd.n2772 gnd 0.006084f
C4798 vdd.n2773 gnd 0.006084f
C4799 vdd.n2774 gnd 0.006084f
C4800 vdd.n2775 gnd 0.006084f
C4801 vdd.n2776 gnd 0.006084f
C4802 vdd.n2777 gnd 0.006084f
C4803 vdd.n2778 gnd 0.006084f
C4804 vdd.n2779 gnd 0.006084f
C4805 vdd.n2780 gnd 0.006084f
C4806 vdd.n2781 gnd 0.006084f
C4807 vdd.n2782 gnd 0.006084f
C4808 vdd.n2783 gnd 0.006084f
C4809 vdd.n2784 gnd 0.006084f
C4810 vdd.n2785 gnd 0.006084f
C4811 vdd.n2786 gnd 0.006084f
C4812 vdd.n2787 gnd 0.006084f
C4813 vdd.n2788 gnd 0.006084f
C4814 vdd.n2789 gnd 0.006084f
C4815 vdd.n2790 gnd 0.006084f
C4816 vdd.n2791 gnd 0.006084f
C4817 vdd.n2792 gnd 0.006084f
C4818 vdd.n2793 gnd 0.006084f
C4819 vdd.n2794 gnd 0.006084f
C4820 vdd.n2795 gnd 0.006084f
C4821 vdd.n2796 gnd 0.006084f
C4822 vdd.n2797 gnd 0.006084f
C4823 vdd.n2798 gnd 0.006084f
C4824 vdd.n2799 gnd 0.006084f
C4825 vdd.n2800 gnd 0.758876f
C4826 vdd.n2802 gnd 0.013814f
C4827 vdd.n2803 gnd 0.013814f
C4828 vdd.n2804 gnd 0.013026f
C4829 vdd.n2805 gnd 0.006084f
C4830 vdd.n2806 gnd 0.006084f
C4831 vdd.n2807 gnd 0.365723f
C4832 vdd.n2808 gnd 0.006084f
C4833 vdd.n2809 gnd 0.006084f
C4834 vdd.n2810 gnd 0.006084f
C4835 vdd.n2811 gnd 0.006084f
C4836 vdd.n2812 gnd 0.006084f
C4837 vdd.n2813 gnd 0.370295f
C4838 vdd.n2814 gnd 0.006084f
C4839 vdd.n2815 gnd 0.006084f
C4840 vdd.n2816 gnd 0.006084f
C4841 vdd.n2817 gnd 0.006084f
C4842 vdd.n2818 gnd 0.006084f
C4843 vdd.n2819 gnd 0.62173f
C4844 vdd.n2820 gnd 0.006084f
C4845 vdd.n2821 gnd 0.006084f
C4846 vdd.n2822 gnd 0.006084f
C4847 vdd.n2823 gnd 0.006084f
C4848 vdd.n2824 gnd 0.006084f
C4849 vdd.n2825 gnd 0.448011f
C4850 vdd.n2826 gnd 0.006084f
C4851 vdd.n2827 gnd 0.006084f
C4852 vdd.n2828 gnd 0.006084f
C4853 vdd.n2829 gnd 0.006084f
C4854 vdd.n2830 gnd 0.006084f
C4855 vdd.n2831 gnd 0.5623f
C4856 vdd.n2832 gnd 0.006084f
C4857 vdd.n2833 gnd 0.006084f
C4858 vdd.n2834 gnd 0.006084f
C4859 vdd.n2835 gnd 0.006084f
C4860 vdd.n2836 gnd 0.006084f
C4861 vdd.n2837 gnd 0.461726f
C4862 vdd.n2838 gnd 0.006084f
C4863 vdd.n2839 gnd 0.006084f
C4864 vdd.n2840 gnd 0.006084f
C4865 vdd.n2841 gnd 0.006084f
C4866 vdd.n2842 gnd 0.006084f
C4867 vdd.n2843 gnd 0.32458f
C4868 vdd.n2844 gnd 0.006084f
C4869 vdd.n2845 gnd 0.006084f
C4870 vdd.n2846 gnd 0.006084f
C4871 vdd.n2847 gnd 0.006084f
C4872 vdd.n2848 gnd 0.006084f
C4873 vdd.n2849 gnd 0.196576f
C4874 vdd.n2850 gnd 0.006084f
C4875 vdd.n2851 gnd 0.006084f
C4876 vdd.n2852 gnd 0.006084f
C4877 vdd.n2853 gnd 0.006084f
C4878 vdd.n2854 gnd 0.006084f
C4879 vdd.n2855 gnd 0.571443f
C4880 vdd.n2856 gnd 0.006084f
C4881 vdd.n2857 gnd 0.006084f
C4882 vdd.n2858 gnd 0.006084f
C4883 vdd.n2859 gnd 0.004294f
C4884 vdd.n2860 gnd 0.006084f
C4885 vdd.n2861 gnd 0.006084f
C4886 vdd.n2862 gnd 0.62173f
C4887 vdd.n2863 gnd 0.006084f
C4888 vdd.n2864 gnd 0.006084f
C4889 vdd.n2865 gnd 0.006084f
C4890 vdd.n2866 gnd 0.006084f
C4891 vdd.n2867 gnd 0.006084f
C4892 vdd.n2868 gnd 0.493727f
C4893 vdd.n2869 gnd 0.006084f
C4894 vdd.n2870 gnd 0.004831f
C4895 vdd.n2871 gnd 0.006084f
C4896 vdd.n2872 gnd 0.006084f
C4897 vdd.n2873 gnd 0.006084f
C4898 vdd.n2874 gnd 0.397724f
C4899 vdd.n2875 gnd 0.006084f
C4900 vdd.n2876 gnd 0.006084f
C4901 vdd.n2877 gnd 0.006084f
C4902 vdd.n2878 gnd 0.006084f
C4903 vdd.n2879 gnd 0.006084f
C4904 vdd.n2880 gnd 0.361152f
C4905 vdd.n2881 gnd 0.006084f
C4906 vdd.n2882 gnd 0.006084f
C4907 vdd.n2883 gnd 0.006084f
C4908 vdd.n2884 gnd 0.006084f
C4909 vdd.n2885 gnd 0.006084f
C4910 vdd.n2886 gnd 0.498298f
C4911 vdd.n2887 gnd 0.006084f
C4912 vdd.n2888 gnd 0.006084f
C4913 vdd.n2889 gnd 0.006084f
C4914 vdd.n2890 gnd 0.006084f
C4915 vdd.n2891 gnd 0.006084f
C4916 vdd.n2892 gnd 0.62173f
C4917 vdd.n2893 gnd 0.006084f
C4918 vdd.n2894 gnd 0.006084f
C4919 vdd.n2895 gnd 0.006084f
C4920 vdd.n2896 gnd 0.006084f
C4921 vdd.n2897 gnd 0.006084f
C4922 vdd.n2898 gnd 0.608015f
C4923 vdd.n2899 gnd 0.006084f
C4924 vdd.n2900 gnd 0.006084f
C4925 vdd.n2901 gnd 0.006084f
C4926 vdd.n2902 gnd 0.006084f
C4927 vdd.n2903 gnd 0.006084f
C4928 vdd.n2904 gnd 0.470869f
C4929 vdd.n2905 gnd 0.006084f
C4930 vdd.n2906 gnd 0.006084f
C4931 vdd.n2907 gnd 0.006084f
C4932 vdd.n2908 gnd 0.006084f
C4933 vdd.n2909 gnd 0.006084f
C4934 vdd.n2910 gnd 0.333723f
C4935 vdd.n2911 gnd 0.006084f
C4936 vdd.n2912 gnd 0.006084f
C4937 vdd.n2913 gnd 0.006084f
C4938 vdd.n2914 gnd 0.006084f
C4939 vdd.n2915 gnd 0.006084f
C4940 vdd.n2916 gnd 0.62173f
C4941 vdd.n2917 gnd 0.006084f
C4942 vdd.n2918 gnd 0.006084f
C4943 vdd.n2919 gnd 0.006084f
C4944 vdd.n2920 gnd 0.006084f
C4945 vdd.n2921 gnd 0.006084f
C4946 vdd.n2922 gnd 0.006084f
C4947 vdd.n2924 gnd 0.006084f
C4948 vdd.n2925 gnd 0.006084f
C4949 vdd.n2927 gnd 0.006084f
C4950 vdd.n2928 gnd 0.006084f
C4951 vdd.n2931 gnd 0.006084f
C4952 vdd.n2932 gnd 0.006084f
C4953 vdd.n2933 gnd 0.006084f
C4954 vdd.n2934 gnd 0.006084f
C4955 vdd.n2936 gnd 0.006084f
C4956 vdd.n2937 gnd 0.006084f
C4957 vdd.n2938 gnd 0.006084f
C4958 vdd.n2939 gnd 0.006084f
C4959 vdd.n2940 gnd 0.006084f
C4960 vdd.n2941 gnd 0.006084f
C4961 vdd.n2943 gnd 0.006084f
C4962 vdd.n2944 gnd 0.006084f
C4963 vdd.n2945 gnd 0.006084f
C4964 vdd.n2946 gnd 0.006084f
C4965 vdd.n2947 gnd 0.006084f
C4966 vdd.n2948 gnd 0.006084f
C4967 vdd.n2950 gnd 0.006084f
C4968 vdd.n2951 gnd 0.006084f
C4969 vdd.n2952 gnd 0.006084f
C4970 vdd.n2953 gnd 0.006084f
C4971 vdd.n2954 gnd 0.006084f
C4972 vdd.n2955 gnd 0.006084f
C4973 vdd.n2957 gnd 0.006084f
C4974 vdd.n2958 gnd 0.013814f
C4975 vdd.n2959 gnd 0.013814f
C4976 vdd.n2960 gnd 0.013026f
C4977 vdd.n2961 gnd 0.006084f
C4978 vdd.n2962 gnd 0.006084f
C4979 vdd.n2963 gnd 0.006084f
C4980 vdd.n2964 gnd 0.006084f
C4981 vdd.n2965 gnd 0.006084f
C4982 vdd.n2966 gnd 0.006084f
C4983 vdd.n2967 gnd 0.62173f
C4984 vdd.n2968 gnd 0.006084f
C4985 vdd.n2969 gnd 0.006084f
C4986 vdd.n2970 gnd 0.006084f
C4987 vdd.n2971 gnd 0.006084f
C4988 vdd.n2972 gnd 0.006084f
C4989 vdd.n2973 gnd 0.44344f
C4990 vdd.n2974 gnd 0.006084f
C4991 vdd.n2975 gnd 0.006084f
C4992 vdd.n2976 gnd 0.006084f
C4993 vdd.n2977 gnd 0.013814f
C4994 vdd.n2979 gnd 0.013814f
C4995 vdd.n2980 gnd 0.013026f
C4996 vdd.n2981 gnd 0.006084f
C4997 vdd.n2982 gnd 0.004697f
C4998 vdd.n2983 gnd 0.006084f
C4999 vdd.n2985 gnd 0.006084f
C5000 vdd.n2986 gnd 0.006084f
C5001 vdd.n2987 gnd 0.006084f
C5002 vdd.n2988 gnd 0.006084f
C5003 vdd.n2989 gnd 0.006084f
C5004 vdd.n2990 gnd 0.006084f
C5005 vdd.n2992 gnd 0.006084f
C5006 vdd.n2993 gnd 0.006084f
C5007 vdd.n2994 gnd 0.006084f
C5008 vdd.n2995 gnd 0.006084f
C5009 vdd.n2996 gnd 0.006084f
C5010 vdd.n2997 gnd 0.006084f
C5011 vdd.n2999 gnd 0.006084f
C5012 vdd.n3000 gnd 0.006084f
C5013 vdd.n3001 gnd 0.006084f
C5014 vdd.n3002 gnd 0.006084f
C5015 vdd.n3003 gnd 0.006084f
C5016 vdd.n3004 gnd 0.006084f
C5017 vdd.n3006 gnd 0.006084f
C5018 vdd.n3007 gnd 0.006084f
C5019 vdd.n3008 gnd 0.006084f
C5020 vdd.n3009 gnd 0.9532f
C5021 vdd.n3010 gnd 0.037566f
C5022 vdd.n3011 gnd 0.006084f
C5023 vdd.n3012 gnd 0.006084f
C5024 vdd.n3014 gnd 0.006084f
C5025 vdd.n3015 gnd 0.006084f
C5026 vdd.n3016 gnd 0.006084f
C5027 vdd.n3017 gnd 0.006084f
C5028 vdd.n3018 gnd 0.006084f
C5029 vdd.n3019 gnd 0.006084f
C5030 vdd.n3021 gnd 0.006084f
C5031 vdd.n3022 gnd 0.006084f
C5032 vdd.n3023 gnd 0.006084f
C5033 vdd.n3024 gnd 0.006084f
C5034 vdd.n3025 gnd 0.006084f
C5035 vdd.n3026 gnd 0.006084f
C5036 vdd.n3028 gnd 0.006084f
C5037 vdd.n3029 gnd 0.006084f
C5038 vdd.n3030 gnd 0.006084f
C5039 vdd.n3031 gnd 0.006084f
C5040 vdd.n3032 gnd 0.006084f
C5041 vdd.n3033 gnd 0.006084f
C5042 vdd.n3035 gnd 0.006084f
C5043 vdd.n3036 gnd 0.006084f
C5044 vdd.n3038 gnd 0.006084f
C5045 vdd.n3039 gnd 0.006084f
C5046 vdd.n3040 gnd 0.013814f
C5047 vdd.n3041 gnd 0.013026f
C5048 vdd.n3042 gnd 0.013026f
C5049 vdd.n3043 gnd 0.841164f
C5050 vdd.n3044 gnd 0.013026f
C5051 vdd.n3045 gnd 0.013814f
C5052 vdd.n3046 gnd 0.013026f
C5053 vdd.n3047 gnd 0.006084f
C5054 vdd.n3048 gnd 0.004697f
C5055 vdd.n3049 gnd 0.006084f
C5056 vdd.n3051 gnd 0.006084f
C5057 vdd.n3052 gnd 0.006084f
C5058 vdd.n3053 gnd 0.006084f
C5059 vdd.n3054 gnd 0.006084f
C5060 vdd.n3055 gnd 0.006084f
C5061 vdd.n3056 gnd 0.006084f
C5062 vdd.n3058 gnd 0.006084f
C5063 vdd.n3059 gnd 0.006084f
C5064 vdd.n3060 gnd 0.006084f
C5065 vdd.n3061 gnd 0.006084f
C5066 vdd.n3062 gnd 0.006084f
C5067 vdd.n3063 gnd 0.006084f
C5068 vdd.n3065 gnd 0.006084f
C5069 vdd.n3066 gnd 0.006084f
C5070 vdd.n3067 gnd 0.006084f
C5071 vdd.n3068 gnd 0.006084f
C5072 vdd.n3069 gnd 0.006084f
C5073 vdd.n3070 gnd 0.006084f
C5074 vdd.n3072 gnd 0.006084f
C5075 vdd.n3073 gnd 0.006084f
C5076 vdd.n3075 gnd 0.006084f
C5077 vdd.n3076 gnd 0.037566f
C5078 vdd.n3077 gnd 0.9532f
C5079 vdd.n3078 gnd 0.007694f
C5080 vdd.n3079 gnd 0.00342f
C5081 vdd.t180 gnd 0.110068f
C5082 vdd.t181 gnd 0.117632f
C5083 vdd.t178 gnd 0.143747f
C5084 vdd.n3080 gnd 0.184263f
C5085 vdd.n3081 gnd 0.154815f
C5086 vdd.n3082 gnd 0.01109f
C5087 vdd.n3083 gnd 0.008947f
C5088 vdd.n3084 gnd 0.003781f
C5089 vdd.n3085 gnd 0.007201f
C5090 vdd.n3086 gnd 0.008947f
C5091 vdd.n3087 gnd 0.008947f
C5092 vdd.n3088 gnd 0.007201f
C5093 vdd.n3089 gnd 0.007201f
C5094 vdd.n3090 gnd 0.008947f
C5095 vdd.n3092 gnd 0.008947f
C5096 vdd.n3093 gnd 0.007201f
C5097 vdd.n3094 gnd 0.007201f
C5098 vdd.n3095 gnd 0.007201f
C5099 vdd.n3096 gnd 0.008947f
C5100 vdd.n3098 gnd 0.008947f
C5101 vdd.n3100 gnd 0.008947f
C5102 vdd.n3101 gnd 0.007201f
C5103 vdd.n3102 gnd 0.007201f
C5104 vdd.n3103 gnd 0.007201f
C5105 vdd.n3104 gnd 0.008947f
C5106 vdd.n3106 gnd 0.008947f
C5107 vdd.n3108 gnd 0.008947f
C5108 vdd.n3109 gnd 0.007201f
C5109 vdd.n3110 gnd 0.007201f
C5110 vdd.n3111 gnd 0.007201f
C5111 vdd.n3112 gnd 0.008947f
C5112 vdd.n3114 gnd 0.008947f
C5113 vdd.n3115 gnd 0.008947f
C5114 vdd.n3116 gnd 0.007201f
C5115 vdd.n3117 gnd 0.007201f
C5116 vdd.n3118 gnd 0.008947f
C5117 vdd.n3119 gnd 0.008947f
C5118 vdd.n3121 gnd 0.008947f
C5119 vdd.n3122 gnd 0.007201f
C5120 vdd.n3123 gnd 0.008947f
C5121 vdd.n3124 gnd 0.008947f
C5122 vdd.n3125 gnd 0.008947f
C5123 vdd.n3126 gnd 0.01469f
C5124 vdd.n3127 gnd 0.004897f
C5125 vdd.n3128 gnd 0.008947f
C5126 vdd.n3130 gnd 0.008947f
C5127 vdd.n3132 gnd 0.008947f
C5128 vdd.n3133 gnd 0.007201f
C5129 vdd.n3134 gnd 0.007201f
C5130 vdd.n3135 gnd 0.007201f
C5131 vdd.n3136 gnd 0.008947f
C5132 vdd.n3138 gnd 0.008947f
C5133 vdd.n3140 gnd 0.008947f
C5134 vdd.n3141 gnd 0.007201f
C5135 vdd.n3142 gnd 0.007201f
C5136 vdd.n3143 gnd 0.007201f
C5137 vdd.n3144 gnd 0.008947f
C5138 vdd.n3146 gnd 0.008947f
C5139 vdd.n3148 gnd 0.008947f
C5140 vdd.n3149 gnd 0.007201f
C5141 vdd.n3150 gnd 0.007201f
C5142 vdd.n3151 gnd 0.007201f
C5143 vdd.n3152 gnd 0.008947f
C5144 vdd.n3154 gnd 0.008947f
C5145 vdd.n3156 gnd 0.008947f
C5146 vdd.n3157 gnd 0.007201f
C5147 vdd.n3158 gnd 0.007201f
C5148 vdd.n3159 gnd 0.007201f
C5149 vdd.n3160 gnd 0.008947f
C5150 vdd.n3162 gnd 0.008947f
C5151 vdd.n3164 gnd 0.008947f
C5152 vdd.n3165 gnd 0.007201f
C5153 vdd.n3166 gnd 0.007201f
C5154 vdd.n3167 gnd 0.006013f
C5155 vdd.n3168 gnd 0.008947f
C5156 vdd.n3170 gnd 0.008947f
C5157 vdd.n3172 gnd 0.008947f
C5158 vdd.n3173 gnd 0.006013f
C5159 vdd.n3174 gnd 0.007201f
C5160 vdd.n3175 gnd 0.007201f
C5161 vdd.n3176 gnd 0.008947f
C5162 vdd.n3178 gnd 0.008947f
C5163 vdd.n3180 gnd 0.008947f
C5164 vdd.n3181 gnd 0.007201f
C5165 vdd.n3182 gnd 0.007201f
C5166 vdd.n3183 gnd 0.007201f
C5167 vdd.n3184 gnd 0.008947f
C5168 vdd.n3186 gnd 0.008947f
C5169 vdd.n3188 gnd 0.008947f
C5170 vdd.n3189 gnd 0.007201f
C5171 vdd.n3190 gnd 0.007201f
C5172 vdd.n3191 gnd 0.007201f
C5173 vdd.n3192 gnd 0.008947f
C5174 vdd.n3194 gnd 0.008947f
C5175 vdd.n3195 gnd 0.008947f
C5176 vdd.n3196 gnd 0.007201f
C5177 vdd.n3197 gnd 0.007201f
C5178 vdd.n3198 gnd 0.008947f
C5179 vdd.n3199 gnd 0.008947f
C5180 vdd.n3200 gnd 0.007201f
C5181 vdd.n3201 gnd 0.007201f
C5182 vdd.n3202 gnd 0.008947f
C5183 vdd.n3203 gnd 0.008947f
C5184 vdd.n3205 gnd 0.008947f
C5185 vdd.n3206 gnd 0.007201f
C5186 vdd.n3207 gnd 0.005977f
C5187 vdd.n3208 gnd 0.021413f
C5188 vdd.n3209 gnd 0.021084f
C5189 vdd.n3210 gnd 0.005977f
C5190 vdd.n3211 gnd 0.021084f
C5191 vdd.n3212 gnd 1.25717f
C5192 vdd.n3213 gnd 0.021084f
C5193 vdd.n3214 gnd 0.005977f
C5194 vdd.n3215 gnd 0.021084f
C5195 vdd.n3216 gnd 0.008947f
C5196 vdd.n3217 gnd 0.008947f
C5197 vdd.n3218 gnd 0.007201f
C5198 vdd.n3219 gnd 0.008947f
C5199 vdd.n3220 gnd 0.914309f
C5200 vdd.n3221 gnd 0.008947f
C5201 vdd.n3222 gnd 0.007201f
C5202 vdd.n3223 gnd 0.008947f
C5203 vdd.n3224 gnd 0.008947f
C5204 vdd.n3225 gnd 0.008947f
C5205 vdd.n3226 gnd 0.007201f
C5206 vdd.n3227 gnd 0.008947f
C5207 vdd.n3228 gnd 0.809163f
C5208 vdd.n3229 gnd 0.008947f
C5209 vdd.n3230 gnd 0.007201f
C5210 vdd.n3231 gnd 0.008947f
C5211 vdd.n3232 gnd 0.008947f
C5212 vdd.n3233 gnd 0.008947f
C5213 vdd.n3234 gnd 0.007201f
C5214 vdd.n3235 gnd 0.008947f
C5215 vdd.t92 gnd 0.457154f
C5216 vdd.n3236 gnd 0.653731f
C5217 vdd.n3237 gnd 0.008947f
C5218 vdd.n3238 gnd 0.007201f
C5219 vdd.n3239 gnd 0.008947f
C5220 vdd.n3240 gnd 0.008947f
C5221 vdd.n3241 gnd 0.008947f
C5222 vdd.n3242 gnd 0.007201f
C5223 vdd.n3243 gnd 0.008947f
C5224 vdd.n3244 gnd 0.498298f
C5225 vdd.n3245 gnd 0.008947f
C5226 vdd.n3246 gnd 0.007201f
C5227 vdd.n3247 gnd 0.008947f
C5228 vdd.n3248 gnd 0.008947f
C5229 vdd.n3249 gnd 0.008947f
C5230 vdd.n3250 gnd 0.007201f
C5231 vdd.n3251 gnd 0.008947f
C5232 vdd.n3252 gnd 0.644588f
C5233 vdd.n3253 gnd 0.571443f
C5234 vdd.n3254 gnd 0.008947f
C5235 vdd.n3255 gnd 0.007201f
C5236 vdd.n3256 gnd 0.008947f
C5237 vdd.n3257 gnd 0.008947f
C5238 vdd.n3258 gnd 0.008947f
C5239 vdd.n3259 gnd 0.007201f
C5240 vdd.n3260 gnd 0.008947f
C5241 vdd.n3261 gnd 0.726875f
C5242 vdd.n3262 gnd 0.008947f
C5243 vdd.n3263 gnd 0.007201f
C5244 vdd.n3264 gnd 0.008947f
C5245 vdd.n3265 gnd 0.008947f
C5246 vdd.n3266 gnd 0.008947f
C5247 vdd.n3267 gnd 0.007201f
C5248 vdd.n3268 gnd 0.007201f
C5249 vdd.n3269 gnd 0.007201f
C5250 vdd.n3270 gnd 0.008947f
C5251 vdd.n3271 gnd 0.008947f
C5252 vdd.n3272 gnd 0.008947f
C5253 vdd.n3273 gnd 0.007201f
C5254 vdd.n3274 gnd 0.007201f
C5255 vdd.n3275 gnd 0.007201f
C5256 vdd.n3276 gnd 0.008947f
C5257 vdd.n3277 gnd 0.008947f
C5258 vdd.n3278 gnd 0.008947f
C5259 vdd.n3279 gnd 0.007201f
C5260 vdd.n3280 gnd 0.007201f
C5261 vdd.n3281 gnd 0.007201f
C5262 vdd.n3282 gnd 0.008947f
C5263 vdd.n3283 gnd 0.008947f
C5264 vdd.n3284 gnd 0.008947f
C5265 vdd.n3285 gnd 0.007201f
C5266 vdd.n3286 gnd 0.007201f
C5267 vdd.n3287 gnd 0.005977f
C5268 vdd.n3288 gnd 0.021084f
C5269 vdd.n3289 gnd 0.021413f
C5270 vdd.n3291 gnd 0.021413f
C5271 vdd.n3292 gnd 0.00342f
C5272 vdd.t195 gnd 0.110068f
C5273 vdd.t194 gnd 0.117632f
C5274 vdd.t193 gnd 0.143747f
C5275 vdd.n3293 gnd 0.184263f
C5276 vdd.n3294 gnd 0.155535f
C5277 vdd.n3295 gnd 0.01181f
C5278 vdd.n3296 gnd 0.003781f
C5279 vdd.n3297 gnd 0.007201f
C5280 vdd.n3298 gnd 0.008947f
C5281 vdd.n3300 gnd 0.008947f
C5282 vdd.n3301 gnd 0.008947f
C5283 vdd.n3302 gnd 0.007201f
C5284 vdd.n3303 gnd 0.007201f
C5285 vdd.n3304 gnd 0.007201f
C5286 vdd.n3305 gnd 0.008947f
C5287 vdd.n3307 gnd 0.008947f
C5288 vdd.n3308 gnd 0.008947f
C5289 vdd.n3309 gnd 0.007201f
C5290 vdd.n3310 gnd 0.007201f
C5291 vdd.n3311 gnd 0.007201f
C5292 vdd.n3312 gnd 0.008947f
C5293 vdd.n3314 gnd 0.008947f
C5294 vdd.n3315 gnd 0.008947f
C5295 vdd.n3316 gnd 0.007201f
C5296 vdd.n3317 gnd 0.007201f
C5297 vdd.n3318 gnd 0.007201f
C5298 vdd.n3319 gnd 0.008947f
C5299 vdd.n3321 gnd 0.008947f
C5300 vdd.n3322 gnd 0.008947f
C5301 vdd.n3323 gnd 0.007201f
C5302 vdd.n3324 gnd 0.007201f
C5303 vdd.n3325 gnd 0.007201f
C5304 vdd.n3326 gnd 0.008947f
C5305 vdd.n3328 gnd 0.008947f
C5306 vdd.n3329 gnd 0.008947f
C5307 vdd.n3330 gnd 0.007201f
C5308 vdd.n3331 gnd 0.008947f
C5309 vdd.n3332 gnd 0.008947f
C5310 vdd.n3333 gnd 0.008947f
C5311 vdd.n3334 gnd 0.01541f
C5312 vdd.n3335 gnd 0.004897f
C5313 vdd.n3336 gnd 0.007201f
C5314 vdd.n3337 gnd 0.008947f
C5315 vdd.n3339 gnd 0.008947f
C5316 vdd.n3340 gnd 0.008947f
C5317 vdd.n3341 gnd 0.007201f
C5318 vdd.n3342 gnd 0.007201f
C5319 vdd.n3343 gnd 0.007201f
C5320 vdd.n3344 gnd 0.008947f
C5321 vdd.n3346 gnd 0.008947f
C5322 vdd.n3347 gnd 0.008947f
C5323 vdd.n3348 gnd 0.007201f
C5324 vdd.n3349 gnd 0.007201f
C5325 vdd.n3350 gnd 0.007201f
C5326 vdd.n3351 gnd 0.008947f
C5327 vdd.n3353 gnd 0.008947f
C5328 vdd.n3354 gnd 0.008947f
C5329 vdd.n3355 gnd 0.007201f
C5330 vdd.n3356 gnd 0.007201f
C5331 vdd.n3357 gnd 0.007201f
C5332 vdd.n3358 gnd 0.008947f
C5333 vdd.n3360 gnd 0.008947f
C5334 vdd.n3361 gnd 0.008947f
C5335 vdd.n3362 gnd 0.007201f
C5336 vdd.n3363 gnd 0.007201f
C5337 vdd.n3364 gnd 0.007201f
C5338 vdd.n3365 gnd 0.008947f
C5339 vdd.n3367 gnd 0.008947f
C5340 vdd.n3368 gnd 0.008947f
C5341 vdd.n3369 gnd 0.007201f
C5342 vdd.n3370 gnd 0.008947f
C5343 vdd.n3371 gnd 0.008947f
C5344 vdd.n3372 gnd 0.008947f
C5345 vdd.n3373 gnd 0.01541f
C5346 vdd.n3374 gnd 0.006013f
C5347 vdd.n3375 gnd 0.007201f
C5348 vdd.n3376 gnd 0.008947f
C5349 vdd.n3378 gnd 0.008947f
C5350 vdd.n3379 gnd 0.008947f
C5351 vdd.n3380 gnd 0.007201f
C5352 vdd.n3381 gnd 0.007201f
C5353 vdd.n3382 gnd 0.007201f
C5354 vdd.n3383 gnd 0.008947f
C5355 vdd.n3385 gnd 0.008947f
C5356 vdd.n3386 gnd 0.008947f
C5357 vdd.n3387 gnd 0.007201f
C5358 vdd.n3388 gnd 0.007201f
C5359 vdd.n3389 gnd 0.007201f
C5360 vdd.n3390 gnd 0.008947f
C5361 vdd.n3392 gnd 0.008947f
C5362 vdd.n3393 gnd 0.008947f
C5363 vdd.n3394 gnd 0.007201f
C5364 vdd.n3395 gnd 0.007201f
C5365 vdd.n3396 gnd 0.007201f
C5366 vdd.n3397 gnd 0.008947f
C5367 vdd.n3399 gnd 0.008947f
C5368 vdd.n3400 gnd 0.008947f
C5369 vdd.n3402 gnd 0.008947f
C5370 vdd.n3403 gnd 0.007201f
C5371 vdd.n3404 gnd 0.007201f
C5372 vdd.n3405 gnd 0.005977f
C5373 vdd.n3406 gnd 0.021413f
C5374 vdd.n3407 gnd 0.021084f
C5375 vdd.n3408 gnd 0.005977f
C5376 vdd.n3409 gnd 0.021084f
C5377 vdd.n3410 gnd 1.28918f
C5378 vdd.n3411 gnd 0.516584f
C5379 vdd.t183 gnd 0.457154f
C5380 vdd.n3412 gnd 0.854879f
C5381 vdd.n3413 gnd 0.008947f
C5382 vdd.n3414 gnd 0.007201f
C5383 vdd.n3415 gnd 0.007201f
C5384 vdd.n3416 gnd 0.007201f
C5385 vdd.n3417 gnd 0.008947f
C5386 vdd.n3418 gnd 0.900594f
C5387 vdd.t72 gnd 0.457154f
C5388 vdd.n3419 gnd 0.470869f
C5389 vdd.n3420 gnd 0.745162f
C5390 vdd.n3421 gnd 0.008947f
C5391 vdd.n3422 gnd 0.007201f
C5392 vdd.n3423 gnd 0.007201f
C5393 vdd.n3424 gnd 0.007201f
C5394 vdd.n3425 gnd 0.008947f
C5395 vdd.n3426 gnd 0.589729f
C5396 vdd.t98 gnd 0.457154f
C5397 vdd.n3427 gnd 0.758876f
C5398 vdd.t64 gnd 0.457154f
C5399 vdd.n3428 gnd 0.480012f
C5400 vdd.n3429 gnd 0.008947f
C5401 vdd.n3430 gnd 0.007201f
C5402 vdd.n3431 gnd 0.007201f
C5403 vdd.n3432 gnd 0.007201f
C5404 vdd.n3433 gnd 0.008947f
C5405 vdd.n3434 gnd 0.635445f
C5406 vdd.n3435 gnd 0.580586f
C5407 vdd.t110 gnd 0.457154f
C5408 vdd.n3436 gnd 0.758876f
C5409 vdd.n3437 gnd 0.008947f
C5410 vdd.n3438 gnd 0.007201f
C5411 vdd.n3439 gnd 0.532576f
C5412 vdd.n3440 gnd 2.29632f
C5413 a_n2804_13878.t18 gnd 0.194556f
C5414 a_n2804_13878.t5 gnd 0.194556f
C5415 a_n2804_13878.t15 gnd 0.194556f
C5416 a_n2804_13878.n0 gnd 1.53358f
C5417 a_n2804_13878.t20 gnd 0.194556f
C5418 a_n2804_13878.t10 gnd 0.194556f
C5419 a_n2804_13878.n1 gnd 1.53196f
C5420 a_n2804_13878.n2 gnd 2.14061f
C5421 a_n2804_13878.t16 gnd 0.194556f
C5422 a_n2804_13878.t9 gnd 0.194556f
C5423 a_n2804_13878.n3 gnd 1.53196f
C5424 a_n2804_13878.n4 gnd 1.04414f
C5425 a_n2804_13878.t3 gnd 0.194556f
C5426 a_n2804_13878.t6 gnd 0.194556f
C5427 a_n2804_13878.n5 gnd 1.53196f
C5428 a_n2804_13878.n6 gnd 1.04414f
C5429 a_n2804_13878.t19 gnd 0.194556f
C5430 a_n2804_13878.t4 gnd 0.194556f
C5431 a_n2804_13878.n7 gnd 1.53196f
C5432 a_n2804_13878.n8 gnd 1.04414f
C5433 a_n2804_13878.t14 gnd 0.194556f
C5434 a_n2804_13878.t2 gnd 0.194556f
C5435 a_n2804_13878.n9 gnd 1.53196f
C5436 a_n2804_13878.n10 gnd 4.90178f
C5437 a_n2804_13878.t30 gnd 1.82172f
C5438 a_n2804_13878.t0 gnd 0.194556f
C5439 a_n2804_13878.t29 gnd 0.194556f
C5440 a_n2804_13878.n11 gnd 1.37045f
C5441 a_n2804_13878.n12 gnd 1.53128f
C5442 a_n2804_13878.t27 gnd 1.81809f
C5443 a_n2804_13878.n13 gnd 0.770559f
C5444 a_n2804_13878.t26 gnd 1.81809f
C5445 a_n2804_13878.n14 gnd 0.770559f
C5446 a_n2804_13878.t28 gnd 0.194556f
C5447 a_n2804_13878.t25 gnd 0.194556f
C5448 a_n2804_13878.n15 gnd 1.37045f
C5449 a_n2804_13878.n16 gnd 0.778022f
C5450 a_n2804_13878.t31 gnd 1.81809f
C5451 a_n2804_13878.n17 gnd 2.85814f
C5452 a_n2804_13878.n18 gnd 3.74876f
C5453 a_n2804_13878.t8 gnd 0.194556f
C5454 a_n2804_13878.t17 gnd 0.194556f
C5455 a_n2804_13878.n19 gnd 1.53195f
C5456 a_n2804_13878.n20 gnd 2.50239f
C5457 a_n2804_13878.t21 gnd 0.194556f
C5458 a_n2804_13878.t7 gnd 0.194556f
C5459 a_n2804_13878.n21 gnd 1.53196f
C5460 a_n2804_13878.n22 gnd 0.678771f
C5461 a_n2804_13878.t11 gnd 0.194556f
C5462 a_n2804_13878.t12 gnd 0.194556f
C5463 a_n2804_13878.n23 gnd 1.53196f
C5464 a_n2804_13878.n24 gnd 0.678771f
C5465 a_n2804_13878.t22 gnd 0.194556f
C5466 a_n2804_13878.t23 gnd 0.194556f
C5467 a_n2804_13878.n25 gnd 1.53196f
C5468 a_n2804_13878.n26 gnd 0.678771f
C5469 a_n2804_13878.t1 gnd 0.194556f
C5470 a_n2804_13878.t13 gnd 0.194556f
C5471 a_n2804_13878.n27 gnd 1.53196f
C5472 a_n2804_13878.n28 gnd 1.37704f
C5473 a_n2804_13878.n29 gnd 1.5345f
C5474 a_n2804_13878.t24 gnd 0.194556f
C5475 a_n2982_13878.n0 gnd 3.88594f
C5476 a_n2982_13878.n1 gnd 2.85743f
C5477 a_n2982_13878.n2 gnd 3.82475f
C5478 a_n2982_13878.n3 gnd 0.806598f
C5479 a_n2982_13878.n4 gnd 0.8066f
C5480 a_n2982_13878.n5 gnd 0.916876f
C5481 a_n2982_13878.n6 gnd 0.201555f
C5482 a_n2982_13878.n7 gnd 0.148449f
C5483 a_n2982_13878.n8 gnd 0.233314f
C5484 a_n2982_13878.n9 gnd 0.180209f
C5485 a_n2982_13878.n10 gnd 0.201555f
C5486 a_n2982_13878.n11 gnd 1.34265f
C5487 a_n2982_13878.n12 gnd 0.148449f
C5488 a_n2982_13878.n13 gnd 0.969982f
C5489 a_n2982_13878.n14 gnd 0.212423f
C5490 a_n2982_13878.n15 gnd 0.747657f
C5491 a_n2982_13878.n16 gnd 0.212423f
C5492 a_n2982_13878.n17 gnd 0.212423f
C5493 a_n2982_13878.n18 gnd 0.483791f
C5494 a_n2982_13878.n19 gnd 0.278519f
C5495 a_n2982_13878.n20 gnd 0.212423f
C5496 a_n2982_13878.n21 gnd 0.536897f
C5497 a_n2982_13878.n22 gnd 0.212423f
C5498 a_n2982_13878.n23 gnd 0.212423f
C5499 a_n2982_13878.n24 gnd 0.945129f
C5500 a_n2982_13878.n25 gnd 0.278519f
C5501 a_n2982_13878.n26 gnd 0.985614f
C5502 a_n2982_13878.n27 gnd 0.212423f
C5503 a_n2982_13878.n28 gnd 0.212423f
C5504 a_n2982_13878.n29 gnd 0.483791f
C5505 a_n2982_13878.n30 gnd 0.212423f
C5506 a_n2982_13878.n31 gnd 0.278519f
C5507 a_n2982_13878.n32 gnd 3.26746f
C5508 a_n2982_13878.n33 gnd 0.278518f
C5509 a_n2982_13878.n34 gnd 0.106212f
C5510 a_n2982_13878.n35 gnd 0.212423f
C5511 a_n2982_13878.n36 gnd 0.85592f
C5512 a_n2982_13878.n37 gnd 0.212423f
C5513 a_n2982_13878.n38 gnd 0.278519f
C5514 a_n2982_13878.n39 gnd 1.74886f
C5515 a_n2982_13878.n40 gnd 1.17841f
C5516 a_n2982_13878.n41 gnd 2.35355f
C5517 a_n2982_13878.n42 gnd 1.17841f
C5518 a_n2982_13878.n43 gnd 2.1518f
C5519 a_n2982_13878.n44 gnd 1.74886f
C5520 a_n2982_13878.n45 gnd 0.008523f
C5521 a_n2982_13878.n46 gnd 4.11e-19
C5522 a_n2982_13878.n48 gnd 0.008224f
C5523 a_n2982_13878.n49 gnd 0.011959f
C5524 a_n2982_13878.n50 gnd 0.004385f
C5525 a_n2982_13878.n51 gnd 0.008523f
C5526 a_n2982_13878.n52 gnd 4.11e-19
C5527 a_n2982_13878.n54 gnd 0.008224f
C5528 a_n2982_13878.n55 gnd 0.011959f
C5529 a_n2982_13878.n56 gnd 0.007912f
C5530 a_n2982_13878.n58 gnd 0.28176f
C5531 a_n2982_13878.n59 gnd 0.008523f
C5532 a_n2982_13878.n60 gnd 4.11e-19
C5533 a_n2982_13878.n62 gnd 0.008224f
C5534 a_n2982_13878.n63 gnd 0.011959f
C5535 a_n2982_13878.n64 gnd 0.007912f
C5536 a_n2982_13878.n66 gnd 0.28176f
C5537 a_n2982_13878.n67 gnd 0.008523f
C5538 a_n2982_13878.n68 gnd 4.11e-19
C5539 a_n2982_13878.n70 gnd 0.008224f
C5540 a_n2982_13878.n71 gnd 0.011959f
C5541 a_n2982_13878.n72 gnd 0.007912f
C5542 a_n2982_13878.n74 gnd 0.28176f
C5543 a_n2982_13878.n75 gnd 0.008224f
C5544 a_n2982_13878.n76 gnd 0.280611f
C5545 a_n2982_13878.n77 gnd 0.008224f
C5546 a_n2982_13878.n78 gnd 0.280611f
C5547 a_n2982_13878.n79 gnd 0.008224f
C5548 a_n2982_13878.n80 gnd 0.280611f
C5549 a_n2982_13878.n81 gnd 0.008224f
C5550 a_n2982_13878.n82 gnd 0.280611f
C5551 a_n2982_13878.n83 gnd 0.301308f
C5552 a_n2982_13878.t11 gnd 0.699618f
C5553 a_n2982_13878.t37 gnd 0.68535f
C5554 a_n2982_13878.t57 gnd 0.68535f
C5555 a_n2982_13878.t29 gnd 0.68535f
C5556 a_n2982_13878.n84 gnd 0.301188f
C5557 a_n2982_13878.t55 gnd 0.68535f
C5558 a_n2982_13878.t15 gnd 0.68535f
C5559 a_n2982_13878.t17 gnd 0.68535f
C5560 a_n2982_13878.n85 gnd 0.297497f
C5561 a_n2982_13878.t31 gnd 0.68535f
C5562 a_n2982_13878.t41 gnd 0.68535f
C5563 a_n2982_13878.t49 gnd 0.68535f
C5564 a_n2982_13878.t33 gnd 0.699618f
C5565 a_n2982_13878.t110 gnd 0.699618f
C5566 a_n2982_13878.t87 gnd 0.68535f
C5567 a_n2982_13878.t92 gnd 0.68535f
C5568 a_n2982_13878.t80 gnd 0.68535f
C5569 a_n2982_13878.n86 gnd 0.301188f
C5570 a_n2982_13878.t97 gnd 0.68535f
C5571 a_n2982_13878.t106 gnd 0.68535f
C5572 a_n2982_13878.t107 gnd 0.68535f
C5573 a_n2982_13878.n87 gnd 0.297497f
C5574 a_n2982_13878.t74 gnd 0.68535f
C5575 a_n2982_13878.t89 gnd 0.68535f
C5576 a_n2982_13878.t77 gnd 0.68535f
C5577 a_n2982_13878.n88 gnd 0.301308f
C5578 a_n2982_13878.t84 gnd 0.68535f
C5579 a_n2982_13878.t103 gnd 0.696376f
C5580 a_n2982_13878.t24 gnd 1.37961f
C5581 a_n2982_13878.t20 gnd 0.147339f
C5582 a_n2982_13878.t48 gnd 0.147339f
C5583 a_n2982_13878.n89 gnd 1.03786f
C5584 a_n2982_13878.t54 gnd 0.147339f
C5585 a_n2982_13878.t40 gnd 0.147339f
C5586 a_n2982_13878.n90 gnd 1.03786f
C5587 a_n2982_13878.t52 gnd 0.147339f
C5588 a_n2982_13878.t44 gnd 0.147339f
C5589 a_n2982_13878.n91 gnd 1.03786f
C5590 a_n2982_13878.t14 gnd 0.147339f
C5591 a_n2982_13878.t36 gnd 0.147339f
C5592 a_n2982_13878.n92 gnd 1.03786f
C5593 a_n2982_13878.t28 gnd 0.147339f
C5594 a_n2982_13878.t22 gnd 0.147339f
C5595 a_n2982_13878.n93 gnd 1.03786f
C5596 a_n2982_13878.t46 gnd 1.37686f
C5597 a_n2982_13878.t27 gnd 0.68535f
C5598 a_n2982_13878.n94 gnd 0.301308f
C5599 a_n2982_13878.t21 gnd 0.68535f
C5600 a_n2982_13878.t13 gnd 0.68535f
C5601 a_n2982_13878.n95 gnd 0.292258f
C5602 a_n2982_13878.t39 gnd 0.68535f
C5603 a_n2982_13878.n96 gnd 0.303898f
C5604 a_n2982_13878.t51 gnd 0.68535f
C5605 a_n2982_13878.t47 gnd 0.68535f
C5606 a_n2982_13878.n97 gnd 0.297169f
C5607 a_n2982_13878.t23 gnd 0.699618f
C5608 a_n2982_13878.t86 gnd 0.68535f
C5609 a_n2982_13878.n98 gnd 0.301308f
C5610 a_n2982_13878.t95 gnd 0.68535f
C5611 a_n2982_13878.t101 gnd 0.68535f
C5612 a_n2982_13878.n99 gnd 0.292258f
C5613 a_n2982_13878.t105 gnd 0.68535f
C5614 a_n2982_13878.n100 gnd 0.303898f
C5615 a_n2982_13878.t76 gnd 0.68535f
C5616 a_n2982_13878.t79 gnd 0.68535f
C5617 a_n2982_13878.n101 gnd 0.297169f
C5618 a_n2982_13878.t109 gnd 0.699618f
C5619 a_n2982_13878.t78 gnd 0.68535f
C5620 a_n2982_13878.n102 gnd 0.303453f
C5621 a_n2982_13878.t104 gnd 0.68535f
C5622 a_n2982_13878.n103 gnd 0.301188f
C5623 a_n2982_13878.n104 gnd 0.301323f
C5624 a_n2982_13878.t100 gnd 0.68535f
C5625 a_n2982_13878.n105 gnd 0.297497f
C5626 a_n2982_13878.t73 gnd 0.68535f
C5627 a_n2982_13878.n106 gnd 0.297752f
C5628 a_n2982_13878.n107 gnd 0.303454f
C5629 a_n2982_13878.t75 gnd 0.696376f
C5630 a_n2982_13878.t19 gnd 0.68535f
C5631 a_n2982_13878.n108 gnd 0.303453f
C5632 a_n2982_13878.t53 gnd 0.68535f
C5633 a_n2982_13878.n109 gnd 0.301188f
C5634 a_n2982_13878.n110 gnd 0.301323f
C5635 a_n2982_13878.t43 gnd 0.68535f
C5636 a_n2982_13878.n111 gnd 0.297497f
C5637 a_n2982_13878.t35 gnd 0.68535f
C5638 a_n2982_13878.n112 gnd 0.297752f
C5639 a_n2982_13878.n113 gnd 0.303454f
C5640 a_n2982_13878.t45 gnd 0.696376f
C5641 a_n2982_13878.n114 gnd 1.32692f
C5642 a_n2982_13878.t83 gnd 0.68535f
C5643 a_n2982_13878.n115 gnd 0.297497f
C5644 a_n2982_13878.t91 gnd 0.68535f
C5645 a_n2982_13878.n116 gnd 0.297497f
C5646 a_n2982_13878.t81 gnd 0.68535f
C5647 a_n2982_13878.n117 gnd 0.297497f
C5648 a_n2982_13878.t96 gnd 0.68535f
C5649 a_n2982_13878.n118 gnd 0.297497f
C5650 a_n2982_13878.t85 gnd 0.68535f
C5651 a_n2982_13878.n119 gnd 0.292094f
C5652 a_n2982_13878.t111 gnd 0.68535f
C5653 a_n2982_13878.n120 gnd 0.301323f
C5654 a_n2982_13878.t88 gnd 0.696834f
C5655 a_n2982_13878.t98 gnd 0.68535f
C5656 a_n2982_13878.n121 gnd 0.292094f
C5657 a_n2982_13878.t82 gnd 0.68535f
C5658 a_n2982_13878.n122 gnd 0.301323f
C5659 a_n2982_13878.t93 gnd 0.696834f
C5660 a_n2982_13878.t102 gnd 0.68535f
C5661 a_n2982_13878.n123 gnd 0.292094f
C5662 a_n2982_13878.t90 gnd 0.68535f
C5663 a_n2982_13878.n124 gnd 0.301323f
C5664 a_n2982_13878.t108 gnd 0.696834f
C5665 a_n2982_13878.t94 gnd 0.68535f
C5666 a_n2982_13878.n125 gnd 0.292094f
C5667 a_n2982_13878.t72 gnd 0.68535f
C5668 a_n2982_13878.n126 gnd 0.301323f
C5669 a_n2982_13878.t99 gnd 0.696834f
C5670 a_n2982_13878.n127 gnd 1.6691f
C5671 a_n2982_13878.n128 gnd 0.303454f
C5672 a_n2982_13878.n129 gnd 0.297752f
C5673 a_n2982_13878.n130 gnd 0.292258f
C5674 a_n2982_13878.n131 gnd 0.301323f
C5675 a_n2982_13878.n132 gnd 0.303898f
C5676 a_n2982_13878.n133 gnd 0.297169f
C5677 a_n2982_13878.n134 gnd 0.303453f
C5678 a_n2982_13878.t25 gnd 0.68535f
C5679 a_n2982_13878.n135 gnd 0.303454f
C5680 a_n2982_13878.t2 gnd 0.114597f
C5681 a_n2982_13878.t10 gnd 0.114597f
C5682 a_n2982_13878.n136 gnd 1.01487f
C5683 a_n2982_13878.t61 gnd 0.114597f
C5684 a_n2982_13878.t62 gnd 0.114597f
C5685 a_n2982_13878.n137 gnd 1.01262f
C5686 a_n2982_13878.t59 gnd 0.114597f
C5687 a_n2982_13878.t64 gnd 0.114597f
C5688 a_n2982_13878.n138 gnd 1.01262f
C5689 a_n2982_13878.t66 gnd 0.114597f
C5690 a_n2982_13878.t60 gnd 0.114597f
C5691 a_n2982_13878.n139 gnd 1.01487f
C5692 a_n2982_13878.t70 gnd 0.114597f
C5693 a_n2982_13878.t7 gnd 0.114597f
C5694 a_n2982_13878.n140 gnd 1.01262f
C5695 a_n2982_13878.t67 gnd 0.114597f
C5696 a_n2982_13878.t71 gnd 0.114597f
C5697 a_n2982_13878.n141 gnd 1.01262f
C5698 a_n2982_13878.t1 gnd 0.114597f
C5699 a_n2982_13878.t6 gnd 0.114597f
C5700 a_n2982_13878.n142 gnd 1.01262f
C5701 a_n2982_13878.t63 gnd 0.114597f
C5702 a_n2982_13878.t4 gnd 0.114597f
C5703 a_n2982_13878.n143 gnd 1.01262f
C5704 a_n2982_13878.t9 gnd 0.114597f
C5705 a_n2982_13878.t69 gnd 0.114597f
C5706 a_n2982_13878.n144 gnd 1.01262f
C5707 a_n2982_13878.t5 gnd 0.114597f
C5708 a_n2982_13878.t65 gnd 0.114597f
C5709 a_n2982_13878.n145 gnd 1.01487f
C5710 a_n2982_13878.t3 gnd 0.114597f
C5711 a_n2982_13878.t0 gnd 0.114597f
C5712 a_n2982_13878.n146 gnd 1.01262f
C5713 a_n2982_13878.t8 gnd 0.114597f
C5714 a_n2982_13878.t68 gnd 0.114597f
C5715 a_n2982_13878.n147 gnd 1.01262f
C5716 a_n2982_13878.n148 gnd 0.30128f
C5717 a_n2982_13878.n149 gnd 0.292258f
C5718 a_n2982_13878.n150 gnd 0.301323f
C5719 a_n2982_13878.n151 gnd 0.303898f
C5720 a_n2982_13878.n152 gnd 0.297169f
C5721 a_n2982_13878.n153 gnd 0.303453f
C5722 a_n2982_13878.n154 gnd 1.00893f
C5723 a_n2982_13878.t34 gnd 1.37961f
C5724 a_n2982_13878.t50 gnd 0.147339f
C5725 a_n2982_13878.t26 gnd 0.147339f
C5726 a_n2982_13878.n155 gnd 1.03786f
C5727 a_n2982_13878.t32 gnd 0.147339f
C5728 a_n2982_13878.t42 gnd 0.147339f
C5729 a_n2982_13878.n156 gnd 1.03786f
C5730 a_n2982_13878.t16 gnd 0.147339f
C5731 a_n2982_13878.t18 gnd 0.147339f
C5732 a_n2982_13878.n157 gnd 1.03786f
C5733 a_n2982_13878.t30 gnd 0.147339f
C5734 a_n2982_13878.t56 gnd 0.147339f
C5735 a_n2982_13878.n158 gnd 1.03786f
C5736 a_n2982_13878.t38 gnd 0.147339f
C5737 a_n2982_13878.t58 gnd 0.147339f
C5738 a_n2982_13878.n159 gnd 1.03786f
C5739 a_n2982_13878.t12 gnd 1.37686f
C5740 a_n8300_8799.t38 gnd 0.114398f
C5741 a_n8300_8799.t28 gnd 0.114398f
C5742 a_n8300_8799.t27 gnd 0.114398f
C5743 a_n8300_8799.n0 gnd 1.01311f
C5744 a_n8300_8799.t33 gnd 0.114398f
C5745 a_n8300_8799.t32 gnd 0.114398f
C5746 a_n8300_8799.n1 gnd 1.01086f
C5747 a_n8300_8799.n2 gnd 0.805199f
C5748 a_n8300_8799.t3 gnd 0.147083f
C5749 a_n8300_8799.t0 gnd 0.147083f
C5750 a_n8300_8799.n3 gnd 1.16006f
C5751 a_n8300_8799.t17 gnd 0.147083f
C5752 a_n8300_8799.t13 gnd 0.147083f
C5753 a_n8300_8799.n4 gnd 1.15815f
C5754 a_n8300_8799.n5 gnd 1.04104f
C5755 a_n8300_8799.t45 gnd 0.147083f
C5756 a_n8300_8799.t10 gnd 0.147083f
C5757 a_n8300_8799.n6 gnd 1.15815f
C5758 a_n8300_8799.n7 gnd 0.513147f
C5759 a_n8300_8799.t18 gnd 0.147083f
C5760 a_n8300_8799.t15 gnd 0.147083f
C5761 a_n8300_8799.n8 gnd 1.15815f
C5762 a_n8300_8799.n9 gnd 0.513147f
C5763 a_n8300_8799.t46 gnd 0.147083f
C5764 a_n8300_8799.t4 gnd 0.147083f
C5765 a_n8300_8799.n10 gnd 1.15815f
C5766 a_n8300_8799.n11 gnd 0.513147f
C5767 a_n8300_8799.t14 gnd 0.147083f
C5768 a_n8300_8799.t20 gnd 0.147083f
C5769 a_n8300_8799.n12 gnd 1.15815f
C5770 a_n8300_8799.n13 gnd 3.78853f
C5771 a_n8300_8799.t47 gnd 0.147083f
C5772 a_n8300_8799.t11 gnd 0.147083f
C5773 a_n8300_8799.n14 gnd 1.16007f
C5774 a_n8300_8799.t9 gnd 0.147083f
C5775 a_n8300_8799.t2 gnd 0.147083f
C5776 a_n8300_8799.n15 gnd 1.15815f
C5777 a_n8300_8799.n16 gnd 1.04104f
C5778 a_n8300_8799.t8 gnd 0.147083f
C5779 a_n8300_8799.t7 gnd 0.147083f
C5780 a_n8300_8799.n17 gnd 1.15815f
C5781 a_n8300_8799.n18 gnd 0.513147f
C5782 a_n8300_8799.t6 gnd 0.147083f
C5783 a_n8300_8799.t12 gnd 0.147083f
C5784 a_n8300_8799.n19 gnd 1.15815f
C5785 a_n8300_8799.n20 gnd 0.513147f
C5786 a_n8300_8799.t5 gnd 0.147083f
C5787 a_n8300_8799.t19 gnd 0.147083f
C5788 a_n8300_8799.n21 gnd 1.15815f
C5789 a_n8300_8799.n22 gnd 0.513147f
C5790 a_n8300_8799.t16 gnd 0.147083f
C5791 a_n8300_8799.t1 gnd 0.147083f
C5792 a_n8300_8799.n23 gnd 1.15815f
C5793 a_n8300_8799.n24 gnd 2.53268f
C5794 a_n8300_8799.n25 gnd 7.78082f
C5795 a_n8300_8799.n26 gnd 0.053014f
C5796 a_n8300_8799.t74 gnd 0.609875f
C5797 a_n8300_8799.n27 gnd 0.271892f
C5798 a_n8300_8799.t75 gnd 0.609875f
C5799 a_n8300_8799.n28 gnd 0.053014f
C5800 a_n8300_8799.t94 gnd 0.609875f
C5801 a_n8300_8799.n29 gnd 0.266989f
C5802 a_n8300_8799.n30 gnd 0.053014f
C5803 a_n8300_8799.t107 gnd 0.609875f
C5804 a_n8300_8799.n31 gnd 0.266989f
C5805 a_n8300_8799.t108 gnd 0.609875f
C5806 a_n8300_8799.n32 gnd 0.053014f
C5807 a_n8300_8799.t65 gnd 0.609875f
C5808 a_n8300_8799.n33 gnd 0.271892f
C5809 a_n8300_8799.t89 gnd 0.624209f
C5810 a_n8300_8799.t111 gnd 0.609875f
C5811 a_n8300_8799.n34 gnd 0.278164f
C5812 a_n8300_8799.n35 gnd 0.254229f
C5813 a_n8300_8799.n36 gnd 0.215257f
C5814 a_n8300_8799.n37 gnd 0.053014f
C5815 a_n8300_8799.n38 gnd 0.01203f
C5816 a_n8300_8799.t87 gnd 0.609875f
C5817 a_n8300_8799.n39 gnd 0.272382f
C5818 a_n8300_8799.n40 gnd 0.01203f
C5819 a_n8300_8799.n41 gnd 0.053014f
C5820 a_n8300_8799.n42 gnd 0.053014f
C5821 a_n8300_8799.n43 gnd 0.053014f
C5822 a_n8300_8799.n44 gnd 0.272219f
C5823 a_n8300_8799.n45 gnd 0.01203f
C5824 a_n8300_8799.t76 gnd 0.609875f
C5825 a_n8300_8799.n46 gnd 0.272219f
C5826 a_n8300_8799.n47 gnd 0.053014f
C5827 a_n8300_8799.n48 gnd 0.053014f
C5828 a_n8300_8799.n49 gnd 0.053014f
C5829 a_n8300_8799.n50 gnd 0.01203f
C5830 a_n8300_8799.t106 gnd 0.609875f
C5831 a_n8300_8799.n51 gnd 0.272382f
C5832 a_n8300_8799.n52 gnd 0.01203f
C5833 a_n8300_8799.n53 gnd 0.053014f
C5834 a_n8300_8799.n54 gnd 0.053014f
C5835 a_n8300_8799.n55 gnd 0.053014f
C5836 a_n8300_8799.n56 gnd 0.267316f
C5837 a_n8300_8799.n57 gnd 0.01203f
C5838 a_n8300_8799.t92 gnd 0.609875f
C5839 a_n8300_8799.n58 gnd 0.266335f
C5840 a_n8300_8799.n59 gnd 0.296767f
C5841 a_n8300_8799.n60 gnd 0.053014f
C5842 a_n8300_8799.t79 gnd 0.609875f
C5843 a_n8300_8799.n61 gnd 0.271892f
C5844 a_n8300_8799.t80 gnd 0.609875f
C5845 a_n8300_8799.n62 gnd 0.053014f
C5846 a_n8300_8799.t103 gnd 0.609875f
C5847 a_n8300_8799.n63 gnd 0.266989f
C5848 a_n8300_8799.n64 gnd 0.053014f
C5849 a_n8300_8799.t116 gnd 0.609875f
C5850 a_n8300_8799.n65 gnd 0.266989f
C5851 a_n8300_8799.t118 gnd 0.609875f
C5852 a_n8300_8799.n66 gnd 0.053014f
C5853 a_n8300_8799.t71 gnd 0.609875f
C5854 a_n8300_8799.n67 gnd 0.271892f
C5855 a_n8300_8799.t96 gnd 0.624209f
C5856 a_n8300_8799.t119 gnd 0.609875f
C5857 a_n8300_8799.n68 gnd 0.278164f
C5858 a_n8300_8799.n69 gnd 0.254229f
C5859 a_n8300_8799.n70 gnd 0.215257f
C5860 a_n8300_8799.n71 gnd 0.053014f
C5861 a_n8300_8799.n72 gnd 0.01203f
C5862 a_n8300_8799.t93 gnd 0.609875f
C5863 a_n8300_8799.n73 gnd 0.272382f
C5864 a_n8300_8799.n74 gnd 0.01203f
C5865 a_n8300_8799.n75 gnd 0.053014f
C5866 a_n8300_8799.n76 gnd 0.053014f
C5867 a_n8300_8799.n77 gnd 0.053014f
C5868 a_n8300_8799.n78 gnd 0.272219f
C5869 a_n8300_8799.n79 gnd 0.01203f
C5870 a_n8300_8799.t83 gnd 0.609875f
C5871 a_n8300_8799.n80 gnd 0.272219f
C5872 a_n8300_8799.n81 gnd 0.053014f
C5873 a_n8300_8799.n82 gnd 0.053014f
C5874 a_n8300_8799.n83 gnd 0.053014f
C5875 a_n8300_8799.n84 gnd 0.01203f
C5876 a_n8300_8799.t115 gnd 0.609875f
C5877 a_n8300_8799.n85 gnd 0.272382f
C5878 a_n8300_8799.n86 gnd 0.01203f
C5879 a_n8300_8799.n87 gnd 0.053014f
C5880 a_n8300_8799.n88 gnd 0.053014f
C5881 a_n8300_8799.n89 gnd 0.053014f
C5882 a_n8300_8799.n90 gnd 0.267316f
C5883 a_n8300_8799.n91 gnd 0.01203f
C5884 a_n8300_8799.t101 gnd 0.609875f
C5885 a_n8300_8799.n92 gnd 0.266335f
C5886 a_n8300_8799.n93 gnd 0.128065f
C5887 a_n8300_8799.n94 gnd 0.91559f
C5888 a_n8300_8799.n95 gnd 0.053014f
C5889 a_n8300_8799.t58 gnd 0.609875f
C5890 a_n8300_8799.n96 gnd 0.271892f
C5891 a_n8300_8799.t48 gnd 0.609875f
C5892 a_n8300_8799.n97 gnd 0.053014f
C5893 a_n8300_8799.t72 gnd 0.609875f
C5894 a_n8300_8799.n98 gnd 0.266989f
C5895 a_n8300_8799.n99 gnd 0.053014f
C5896 a_n8300_8799.t90 gnd 0.609875f
C5897 a_n8300_8799.n100 gnd 0.266989f
C5898 a_n8300_8799.t78 gnd 0.609875f
C5899 a_n8300_8799.n101 gnd 0.053014f
C5900 a_n8300_8799.t81 gnd 0.609875f
C5901 a_n8300_8799.n102 gnd 0.271892f
C5902 a_n8300_8799.t98 gnd 0.624209f
C5903 a_n8300_8799.t67 gnd 0.609875f
C5904 a_n8300_8799.n103 gnd 0.278164f
C5905 a_n8300_8799.n104 gnd 0.254229f
C5906 a_n8300_8799.n105 gnd 0.215257f
C5907 a_n8300_8799.n106 gnd 0.053014f
C5908 a_n8300_8799.n107 gnd 0.01203f
C5909 a_n8300_8799.t54 gnd 0.609875f
C5910 a_n8300_8799.n108 gnd 0.272382f
C5911 a_n8300_8799.n109 gnd 0.01203f
C5912 a_n8300_8799.n110 gnd 0.053014f
C5913 a_n8300_8799.n111 gnd 0.053014f
C5914 a_n8300_8799.n112 gnd 0.053014f
C5915 a_n8300_8799.n113 gnd 0.272219f
C5916 a_n8300_8799.n114 gnd 0.01203f
C5917 a_n8300_8799.t102 gnd 0.609875f
C5918 a_n8300_8799.n115 gnd 0.272219f
C5919 a_n8300_8799.n116 gnd 0.053014f
C5920 a_n8300_8799.n117 gnd 0.053014f
C5921 a_n8300_8799.n118 gnd 0.053014f
C5922 a_n8300_8799.n119 gnd 0.01203f
C5923 a_n8300_8799.t109 gnd 0.609875f
C5924 a_n8300_8799.n120 gnd 0.272382f
C5925 a_n8300_8799.n121 gnd 0.01203f
C5926 a_n8300_8799.n122 gnd 0.053014f
C5927 a_n8300_8799.n123 gnd 0.053014f
C5928 a_n8300_8799.n124 gnd 0.053014f
C5929 a_n8300_8799.n125 gnd 0.267316f
C5930 a_n8300_8799.n126 gnd 0.01203f
C5931 a_n8300_8799.t84 gnd 0.609875f
C5932 a_n8300_8799.n127 gnd 0.266335f
C5933 a_n8300_8799.n128 gnd 0.128065f
C5934 a_n8300_8799.n129 gnd 1.93713f
C5935 a_n8300_8799.n130 gnd 0.053014f
C5936 a_n8300_8799.t51 gnd 0.609875f
C5937 a_n8300_8799.t50 gnd 0.609875f
C5938 a_n8300_8799.n131 gnd 0.053014f
C5939 a_n8300_8799.t100 gnd 0.609875f
C5940 a_n8300_8799.n132 gnd 0.053014f
C5941 a_n8300_8799.t61 gnd 0.609875f
C5942 a_n8300_8799.n133 gnd 0.272382f
C5943 a_n8300_8799.n134 gnd 0.053014f
C5944 a_n8300_8799.t53 gnd 0.609875f
C5945 a_n8300_8799.t104 gnd 0.609875f
C5946 a_n8300_8799.n135 gnd 0.053014f
C5947 a_n8300_8799.t77 gnd 0.609875f
C5948 a_n8300_8799.n136 gnd 0.272219f
C5949 a_n8300_8799.n137 gnd 0.053014f
C5950 a_n8300_8799.t62 gnd 0.609875f
C5951 a_n8300_8799.t117 gnd 0.609875f
C5952 a_n8300_8799.n138 gnd 0.053014f
C5953 a_n8300_8799.t88 gnd 0.609875f
C5954 a_n8300_8799.n139 gnd 0.271892f
C5955 a_n8300_8799.t113 gnd 0.624209f
C5956 a_n8300_8799.t64 gnd 0.609875f
C5957 a_n8300_8799.n140 gnd 0.278164f
C5958 a_n8300_8799.n141 gnd 0.254229f
C5959 a_n8300_8799.n142 gnd 0.215257f
C5960 a_n8300_8799.n143 gnd 0.053014f
C5961 a_n8300_8799.n144 gnd 0.01203f
C5962 a_n8300_8799.n145 gnd 0.272382f
C5963 a_n8300_8799.n146 gnd 0.01203f
C5964 a_n8300_8799.n147 gnd 0.266989f
C5965 a_n8300_8799.n148 gnd 0.053014f
C5966 a_n8300_8799.n149 gnd 0.053014f
C5967 a_n8300_8799.n150 gnd 0.053014f
C5968 a_n8300_8799.n151 gnd 0.01203f
C5969 a_n8300_8799.n152 gnd 0.272219f
C5970 a_n8300_8799.n153 gnd 0.266989f
C5971 a_n8300_8799.n154 gnd 0.01203f
C5972 a_n8300_8799.n155 gnd 0.053014f
C5973 a_n8300_8799.n156 gnd 0.053014f
C5974 a_n8300_8799.n157 gnd 0.053014f
C5975 a_n8300_8799.n158 gnd 0.01203f
C5976 a_n8300_8799.n159 gnd 0.271892f
C5977 a_n8300_8799.n160 gnd 0.267316f
C5978 a_n8300_8799.n161 gnd 0.01203f
C5979 a_n8300_8799.n162 gnd 0.266335f
C5980 a_n8300_8799.n163 gnd 0.296767f
C5981 a_n8300_8799.n164 gnd 0.053014f
C5982 a_n8300_8799.t57 gnd 0.609875f
C5983 a_n8300_8799.t56 gnd 0.609875f
C5984 a_n8300_8799.n165 gnd 0.053014f
C5985 a_n8300_8799.t112 gnd 0.609875f
C5986 a_n8300_8799.n166 gnd 0.053014f
C5987 a_n8300_8799.t66 gnd 0.609875f
C5988 a_n8300_8799.n167 gnd 0.272382f
C5989 a_n8300_8799.n168 gnd 0.053014f
C5990 a_n8300_8799.t60 gnd 0.609875f
C5991 a_n8300_8799.t114 gnd 0.609875f
C5992 a_n8300_8799.n169 gnd 0.053014f
C5993 a_n8300_8799.t86 gnd 0.609875f
C5994 a_n8300_8799.n170 gnd 0.272219f
C5995 a_n8300_8799.n171 gnd 0.053014f
C5996 a_n8300_8799.t69 gnd 0.609875f
C5997 a_n8300_8799.t52 gnd 0.609875f
C5998 a_n8300_8799.n172 gnd 0.053014f
C5999 a_n8300_8799.t95 gnd 0.609875f
C6000 a_n8300_8799.n173 gnd 0.271892f
C6001 a_n8300_8799.t49 gnd 0.624209f
C6002 a_n8300_8799.t70 gnd 0.609875f
C6003 a_n8300_8799.n174 gnd 0.278164f
C6004 a_n8300_8799.n175 gnd 0.254229f
C6005 a_n8300_8799.n176 gnd 0.215257f
C6006 a_n8300_8799.n177 gnd 0.053014f
C6007 a_n8300_8799.n178 gnd 0.01203f
C6008 a_n8300_8799.n179 gnd 0.272382f
C6009 a_n8300_8799.n180 gnd 0.01203f
C6010 a_n8300_8799.n181 gnd 0.266989f
C6011 a_n8300_8799.n182 gnd 0.053014f
C6012 a_n8300_8799.n183 gnd 0.053014f
C6013 a_n8300_8799.n184 gnd 0.053014f
C6014 a_n8300_8799.n185 gnd 0.01203f
C6015 a_n8300_8799.n186 gnd 0.272219f
C6016 a_n8300_8799.n187 gnd 0.266989f
C6017 a_n8300_8799.n188 gnd 0.01203f
C6018 a_n8300_8799.n189 gnd 0.053014f
C6019 a_n8300_8799.n190 gnd 0.053014f
C6020 a_n8300_8799.n191 gnd 0.053014f
C6021 a_n8300_8799.n192 gnd 0.01203f
C6022 a_n8300_8799.n193 gnd 0.271892f
C6023 a_n8300_8799.n194 gnd 0.267316f
C6024 a_n8300_8799.n195 gnd 0.01203f
C6025 a_n8300_8799.n196 gnd 0.266335f
C6026 a_n8300_8799.n197 gnd 0.128065f
C6027 a_n8300_8799.n198 gnd 0.91559f
C6028 a_n8300_8799.n199 gnd 0.053014f
C6029 a_n8300_8799.t85 gnd 0.609875f
C6030 a_n8300_8799.t99 gnd 0.609875f
C6031 a_n8300_8799.n200 gnd 0.053014f
C6032 a_n8300_8799.t59 gnd 0.609875f
C6033 a_n8300_8799.n201 gnd 0.053014f
C6034 a_n8300_8799.t110 gnd 0.609875f
C6035 a_n8300_8799.n202 gnd 0.272382f
C6036 a_n8300_8799.n203 gnd 0.053014f
C6037 a_n8300_8799.t73 gnd 0.609875f
C6038 a_n8300_8799.t105 gnd 0.609875f
C6039 a_n8300_8799.n204 gnd 0.053014f
C6040 a_n8300_8799.t63 gnd 0.609875f
C6041 a_n8300_8799.n205 gnd 0.272219f
C6042 a_n8300_8799.n206 gnd 0.053014f
C6043 a_n8300_8799.t91 gnd 0.609875f
C6044 a_n8300_8799.t55 gnd 0.609875f
C6045 a_n8300_8799.n207 gnd 0.053014f
C6046 a_n8300_8799.t82 gnd 0.609875f
C6047 a_n8300_8799.n208 gnd 0.271892f
C6048 a_n8300_8799.t97 gnd 0.624209f
C6049 a_n8300_8799.t68 gnd 0.609875f
C6050 a_n8300_8799.n209 gnd 0.278164f
C6051 a_n8300_8799.n210 gnd 0.254229f
C6052 a_n8300_8799.n211 gnd 0.215257f
C6053 a_n8300_8799.n212 gnd 0.053014f
C6054 a_n8300_8799.n213 gnd 0.01203f
C6055 a_n8300_8799.n214 gnd 0.272382f
C6056 a_n8300_8799.n215 gnd 0.01203f
C6057 a_n8300_8799.n216 gnd 0.266989f
C6058 a_n8300_8799.n217 gnd 0.053014f
C6059 a_n8300_8799.n218 gnd 0.053014f
C6060 a_n8300_8799.n219 gnd 0.053014f
C6061 a_n8300_8799.n220 gnd 0.01203f
C6062 a_n8300_8799.n221 gnd 0.272219f
C6063 a_n8300_8799.n222 gnd 0.266989f
C6064 a_n8300_8799.n223 gnd 0.01203f
C6065 a_n8300_8799.n224 gnd 0.053014f
C6066 a_n8300_8799.n225 gnd 0.053014f
C6067 a_n8300_8799.n226 gnd 0.053014f
C6068 a_n8300_8799.n227 gnd 0.01203f
C6069 a_n8300_8799.n228 gnd 0.271892f
C6070 a_n8300_8799.n229 gnd 0.267316f
C6071 a_n8300_8799.n230 gnd 0.01203f
C6072 a_n8300_8799.n231 gnd 0.266335f
C6073 a_n8300_8799.n232 gnd 0.128065f
C6074 a_n8300_8799.n233 gnd 1.4042f
C6075 a_n8300_8799.n234 gnd 17.7114f
C6076 a_n8300_8799.n235 gnd 4.4634f
C6077 a_n8300_8799.t29 gnd 0.114398f
C6078 a_n8300_8799.t30 gnd 0.114398f
C6079 a_n8300_8799.n236 gnd 1.01311f
C6080 a_n8300_8799.t23 gnd 0.114398f
C6081 a_n8300_8799.t24 gnd 0.114398f
C6082 a_n8300_8799.n237 gnd 1.01086f
C6083 a_n8300_8799.n238 gnd 0.805197f
C6084 a_n8300_8799.t22 gnd 0.114398f
C6085 a_n8300_8799.t40 gnd 0.114398f
C6086 a_n8300_8799.n239 gnd 1.01086f
C6087 a_n8300_8799.n240 gnd 0.336223f
C6088 a_n8300_8799.n241 gnd 0.480018f
C6089 a_n8300_8799.t42 gnd 0.114398f
C6090 a_n8300_8799.t35 gnd 0.114398f
C6091 a_n8300_8799.n242 gnd 1.01086f
C6092 a_n8300_8799.n243 gnd 0.336223f
C6093 a_n8300_8799.t37 gnd 0.114398f
C6094 a_n8300_8799.t21 gnd 0.114398f
C6095 a_n8300_8799.n244 gnd 1.01086f
C6096 a_n8300_8799.n245 gnd 0.395393f
C6097 a_n8300_8799.t39 gnd 0.114398f
C6098 a_n8300_8799.t41 gnd 0.114398f
C6099 a_n8300_8799.n246 gnd 1.01086f
C6100 a_n8300_8799.n247 gnd 2.91093f
C6101 a_n8300_8799.t36 gnd 0.114398f
C6102 a_n8300_8799.t34 gnd 0.114398f
C6103 a_n8300_8799.n248 gnd 1.01311f
C6104 a_n8300_8799.t25 gnd 0.114398f
C6105 a_n8300_8799.t31 gnd 0.114398f
C6106 a_n8300_8799.n249 gnd 1.01086f
C6107 a_n8300_8799.n250 gnd 0.805199f
C6108 a_n8300_8799.t43 gnd 0.114398f
C6109 a_n8300_8799.t26 gnd 0.114398f
C6110 a_n8300_8799.n251 gnd 1.01086f
C6111 a_n8300_8799.n252 gnd 0.336224f
C6112 a_n8300_8799.n253 gnd 2.44997f
C6113 a_n8300_8799.n254 gnd 0.336226f
C6114 a_n8300_8799.n255 gnd 1.01086f
C6115 a_n8300_8799.t44 gnd 0.114398f
C6116 a_n2903_n3924.n0 gnd 2.10908f
C6117 a_n2903_n3924.n1 gnd 2.29654f
C6118 a_n2903_n3924.n2 gnd 1.52909f
C6119 a_n2903_n3924.n3 gnd 1.39023f
C6120 a_n2903_n3924.n4 gnd 1.91428f
C6121 a_n2903_n3924.n5 gnd 1.87222f
C6122 a_n2903_n3924.n6 gnd 1.87222f
C6123 a_n2903_n3924.n7 gnd 2.19334f
C6124 a_n2903_n3924.n8 gnd 1.00796f
C6125 a_n2903_n3924.n9 gnd 0.764541f
C6126 a_n2903_n3924.n10 gnd 1.34454f
C6127 a_n2903_n3924.n11 gnd 1.6947f
C6128 a_n2903_n3924.t5 gnd 0.102925f
C6129 a_n2903_n3924.t26 gnd 0.102925f
C6130 a_n2903_n3924.t3 gnd 0.102925f
C6131 a_n2903_n3924.n12 gnd 0.840609f
C6132 a_n2903_n3924.t15 gnd 1.3291f
C6133 a_n2903_n3924.t27 gnd 0.102925f
C6134 a_n2903_n3924.t8 gnd 0.102925f
C6135 a_n2903_n3924.n13 gnd 0.840609f
C6136 a_n2903_n3924.t4 gnd 0.102925f
C6137 a_n2903_n3924.t9 gnd 0.102925f
C6138 a_n2903_n3924.n14 gnd 0.840609f
C6139 a_n2903_n3924.t6 gnd 0.102925f
C6140 a_n2903_n3924.t18 gnd 0.102925f
C6141 a_n2903_n3924.n15 gnd 0.840609f
C6142 a_n2903_n3924.t1 gnd 1.06972f
C6143 a_n2903_n3924.t55 gnd 1.32974f
C6144 a_n2903_n3924.t19 gnd 1.3291f
C6145 a_n2903_n3924.t24 gnd 1.3291f
C6146 a_n2903_n3924.t21 gnd 1.3291f
C6147 a_n2903_n3924.t14 gnd 1.3291f
C6148 a_n2903_n3924.t53 gnd 1.3291f
C6149 a_n2903_n3924.t11 gnd 1.3291f
C6150 a_n2903_n3924.n16 gnd 0.965474f
C6151 a_n2903_n3924.t47 gnd 1.06972f
C6152 a_n2903_n3924.t46 gnd 0.102925f
C6153 a_n2903_n3924.t32 gnd 0.102925f
C6154 a_n2903_n3924.n17 gnd 0.840607f
C6155 a_n2903_n3924.t30 gnd 0.102925f
C6156 a_n2903_n3924.t29 gnd 0.102925f
C6157 a_n2903_n3924.n18 gnd 0.840607f
C6158 a_n2903_n3924.t45 gnd 0.102925f
C6159 a_n2903_n3924.t48 gnd 0.102925f
C6160 a_n2903_n3924.n19 gnd 0.840607f
C6161 a_n2903_n3924.t49 gnd 0.102925f
C6162 a_n2903_n3924.t43 gnd 0.102925f
C6163 a_n2903_n3924.n20 gnd 0.840607f
C6164 a_n2903_n3924.t39 gnd 0.102925f
C6165 a_n2903_n3924.t36 gnd 0.102925f
C6166 a_n2903_n3924.n21 gnd 0.840607f
C6167 a_n2903_n3924.t42 gnd 1.06972f
C6168 a_n2903_n3924.t2 gnd 1.06972f
C6169 a_n2903_n3924.t10 gnd 0.102925f
C6170 a_n2903_n3924.t16 gnd 0.102925f
C6171 a_n2903_n3924.n22 gnd 0.840607f
C6172 a_n2903_n3924.t17 gnd 0.102925f
C6173 a_n2903_n3924.t12 gnd 0.102925f
C6174 a_n2903_n3924.n23 gnd 0.840607f
C6175 a_n2903_n3924.t20 gnd 0.102925f
C6176 a_n2903_n3924.t25 gnd 0.102925f
C6177 a_n2903_n3924.n24 gnd 0.840607f
C6178 a_n2903_n3924.t54 gnd 0.102925f
C6179 a_n2903_n3924.t52 gnd 0.102925f
C6180 a_n2903_n3924.n25 gnd 0.840607f
C6181 a_n2903_n3924.t7 gnd 0.102925f
C6182 a_n2903_n3924.t23 gnd 0.102925f
C6183 a_n2903_n3924.n26 gnd 0.840607f
C6184 a_n2903_n3924.t13 gnd 1.06972f
C6185 a_n2903_n3924.n27 gnd 1.02539f
C6186 a_n2903_n3924.t37 gnd 1.06972f
C6187 a_n2903_n3924.t35 gnd 0.102925f
C6188 a_n2903_n3924.t33 gnd 0.102925f
C6189 a_n2903_n3924.n28 gnd 0.840609f
C6190 a_n2903_n3924.t31 gnd 0.102925f
C6191 a_n2903_n3924.t34 gnd 0.102925f
C6192 a_n2903_n3924.n29 gnd 0.840609f
C6193 a_n2903_n3924.t40 gnd 0.102925f
C6194 a_n2903_n3924.t41 gnd 0.102925f
C6195 a_n2903_n3924.n30 gnd 0.840609f
C6196 a_n2903_n3924.t38 gnd 0.102925f
C6197 a_n2903_n3924.t51 gnd 0.102925f
C6198 a_n2903_n3924.n31 gnd 0.840609f
C6199 a_n2903_n3924.t28 gnd 0.102925f
C6200 a_n2903_n3924.t44 gnd 0.102925f
C6201 a_n2903_n3924.n32 gnd 0.840609f
C6202 a_n2903_n3924.t50 gnd 1.06972f
C6203 a_n2903_n3924.t22 gnd 1.06972f
C6204 a_n2903_n3924.n33 gnd 0.84061f
C6205 a_n2903_n3924.t0 gnd 0.102925f
C6206 plus.n0 gnd 0.023894f
C6207 plus.t21 gnd 0.337957f
C6208 plus.n1 gnd 0.023894f
C6209 plus.t22 gnd 0.337957f
C6210 plus.t16 gnd 0.337957f
C6211 plus.n2 gnd 0.150131f
C6212 plus.n3 gnd 0.023894f
C6213 plus.t17 gnd 0.337957f
C6214 plus.t11 gnd 0.337957f
C6215 plus.n4 gnd 0.150131f
C6216 plus.n5 gnd 0.023894f
C6217 plus.t5 gnd 0.337957f
C6218 plus.t6 gnd 0.337957f
C6219 plus.n6 gnd 0.150131f
C6220 plus.n7 gnd 0.023894f
C6221 plus.t23 gnd 0.337957f
C6222 plus.t24 gnd 0.337957f
C6223 plus.n8 gnd 0.150131f
C6224 plus.n9 gnd 0.023894f
C6225 plus.t18 gnd 0.337957f
C6226 plus.t13 gnd 0.337957f
C6227 plus.n10 gnd 0.155021f
C6228 plus.t15 gnd 0.350224f
C6229 plus.n11 gnd 0.139136f
C6230 plus.n12 gnd 0.102865f
C6231 plus.n13 gnd 0.005422f
C6232 plus.n14 gnd 0.150131f
C6233 plus.n15 gnd 0.005422f
C6234 plus.n16 gnd 0.023894f
C6235 plus.n17 gnd 0.023894f
C6236 plus.n18 gnd 0.023894f
C6237 plus.n19 gnd 0.005422f
C6238 plus.n20 gnd 0.150131f
C6239 plus.n21 gnd 0.005422f
C6240 plus.n22 gnd 0.023894f
C6241 plus.n23 gnd 0.023894f
C6242 plus.n24 gnd 0.023894f
C6243 plus.n25 gnd 0.005422f
C6244 plus.n26 gnd 0.150131f
C6245 plus.n27 gnd 0.005422f
C6246 plus.n28 gnd 0.023894f
C6247 plus.n29 gnd 0.023894f
C6248 plus.n30 gnd 0.023894f
C6249 plus.n31 gnd 0.005422f
C6250 plus.n32 gnd 0.150131f
C6251 plus.n33 gnd 0.005422f
C6252 plus.n34 gnd 0.023894f
C6253 plus.n35 gnd 0.023894f
C6254 plus.n36 gnd 0.023894f
C6255 plus.n37 gnd 0.005422f
C6256 plus.n38 gnd 0.150131f
C6257 plus.n39 gnd 0.005422f
C6258 plus.n40 gnd 0.150352f
C6259 plus.n41 gnd 0.270561f
C6260 plus.n42 gnd 0.023894f
C6261 plus.n43 gnd 0.005422f
C6262 plus.t10 gnd 0.337957f
C6263 plus.n44 gnd 0.023894f
C6264 plus.n45 gnd 0.005422f
C6265 plus.t12 gnd 0.337957f
C6266 plus.n46 gnd 0.023894f
C6267 plus.n47 gnd 0.005422f
C6268 plus.t7 gnd 0.337957f
C6269 plus.n48 gnd 0.023894f
C6270 plus.n49 gnd 0.005422f
C6271 plus.t27 gnd 0.337957f
C6272 plus.n50 gnd 0.023894f
C6273 plus.n51 gnd 0.005422f
C6274 plus.t26 gnd 0.337957f
C6275 plus.t20 gnd 0.350224f
C6276 plus.t19 gnd 0.337957f
C6277 plus.n52 gnd 0.155021f
C6278 plus.n53 gnd 0.139136f
C6279 plus.n54 gnd 0.102865f
C6280 plus.n55 gnd 0.023894f
C6281 plus.n56 gnd 0.150131f
C6282 plus.n57 gnd 0.005422f
C6283 plus.t25 gnd 0.337957f
C6284 plus.n58 gnd 0.150131f
C6285 plus.n59 gnd 0.023894f
C6286 plus.n60 gnd 0.023894f
C6287 plus.n61 gnd 0.023894f
C6288 plus.n62 gnd 0.150131f
C6289 plus.n63 gnd 0.005422f
C6290 plus.t9 gnd 0.337957f
C6291 plus.n64 gnd 0.150131f
C6292 plus.n65 gnd 0.023894f
C6293 plus.n66 gnd 0.023894f
C6294 plus.n67 gnd 0.023894f
C6295 plus.n68 gnd 0.150131f
C6296 plus.n69 gnd 0.005422f
C6297 plus.t14 gnd 0.337957f
C6298 plus.n70 gnd 0.150131f
C6299 plus.n71 gnd 0.023894f
C6300 plus.n72 gnd 0.023894f
C6301 plus.n73 gnd 0.023894f
C6302 plus.n74 gnd 0.150131f
C6303 plus.n75 gnd 0.005422f
C6304 plus.t28 gnd 0.337957f
C6305 plus.n76 gnd 0.150131f
C6306 plus.n77 gnd 0.023894f
C6307 plus.n78 gnd 0.023894f
C6308 plus.n79 gnd 0.023894f
C6309 plus.n80 gnd 0.150131f
C6310 plus.n81 gnd 0.005422f
C6311 plus.t8 gnd 0.337957f
C6312 plus.n82 gnd 0.150352f
C6313 plus.n83 gnd 0.79089f
C6314 plus.n84 gnd 1.18323f
C6315 plus.t1 gnd 0.041248f
C6316 plus.t2 gnd 0.007366f
C6317 plus.t4 gnd 0.007366f
C6318 plus.n85 gnd 0.023889f
C6319 plus.n86 gnd 0.185449f
C6320 plus.t3 gnd 0.007366f
C6321 plus.t0 gnd 0.007366f
C6322 plus.n87 gnd 0.023889f
C6323 plus.n88 gnd 0.139202f
C6324 plus.n89 gnd 2.79427f
.ends

