* NGSPICE file created from opamp98.ext - technology: sky130A

.subckt opamp98 gnd CSoutput output vdd plus minus commonsourceibias outputibias diffpairibias
X0 gnd.t337 commonsourceibias.t80 CSoutput.t106 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X1 CSoutput.t150 a_n6972_8799.t40 vdd.t229 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X2 commonsourceibias.t47 commonsourceibias.t46 gnd.t336 gnd.t300 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X3 a_n2140_13878.t7 a_n2848_n452.t56 vdd.t107 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 a_n2140_13878.t23 a_n2848_n452.t18 a_n2848_n452.t19 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X5 vdd.t228 a_n6972_8799.t41 CSoutput.t24 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X6 vdd.t79 vdd.t77 vdd.t78 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X7 outputibias.t7 outputibias.t6 gnd.t138 gnd.t137 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X8 gnd.t134 gnd.t132 gnd.t133 gnd.t45 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X9 a_n6972_8799.t35 plus.t5 a_n3106_n452.t26 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X10 a_n3106_n452.t25 plus.t6 a_n6972_8799.t34 gnd.t168 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X11 gnd.t335 commonsourceibias.t81 CSoutput.t105 gnd.t293 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X12 CSoutput.t52 a_n6972_8799.t42 vdd.t227 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X13 CSoutput.t152 a_n2318_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X14 gnd.t330 commonsourceibias.t82 CSoutput.t101 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X15 gnd.t334 commonsourceibias.t44 commonsourceibias.t45 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X16 gnd.t333 commonsourceibias.t83 CSoutput.t104 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X17 a_n2318_8322.t27 a_n2848_n452.t57 a_n6972_8799.t16 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X18 gnd.t332 commonsourceibias.t84 CSoutput.t103 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 output.t15 CSoutput.t153 vdd.t88 gnd.t20 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X20 CSoutput.t39 a_n6972_8799.t43 vdd.t226 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X21 outputibias.t5 outputibias.t4 gnd.t158 gnd.t157 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X22 gnd.t331 commonsourceibias.t85 CSoutput.t102 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X23 vdd.t225 a_n6972_8799.t44 CSoutput.t0 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X24 a_n2848_n452.t46 minus.t5 a_n3106_n452.t41 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X25 gnd.t329 commonsourceibias.t42 commonsourceibias.t43 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X26 a_n6972_8799.t12 plus.t7 a_n3106_n452.t24 gnd.t145 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X27 a_n6972_8799.t30 a_n2848_n452.t58 a_n2318_8322.t26 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X28 a_n2848_n452.t45 minus.t6 a_n3106_n452.t40 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X29 plus.t4 gnd.t129 gnd.t131 gnd.t130 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X30 vdd.t224 a_n6972_8799.t45 CSoutput.t21 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X31 CSoutput.t10 a_n6972_8799.t46 vdd.t223 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X32 a_n6972_8799.t31 a_n2848_n452.t59 a_n2318_8322.t25 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X33 CSoutput.t100 commonsourceibias.t86 gnd.t328 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X34 gnd.t327 commonsourceibias.t40 commonsourceibias.t41 gnd.t289 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 vdd.t76 vdd.t74 vdd.t75 vdd.t5 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X36 CSoutput.t99 commonsourceibias.t87 gnd.t326 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 CSoutput.t45 a_n6972_8799.t47 vdd.t222 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X38 vdd.t93 CSoutput.t154 output.t14 gnd.t19 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X39 a_n3106_n452.t23 plus.t8 a_n6972_8799.t14 gnd.t161 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X40 CSoutput.t98 commonsourceibias.t88 gnd.t325 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X41 CSoutput.t115 commonsourceibias.t89 gnd.t324 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X42 a_n3106_n452.t49 diffpairibias.t16 gnd.t177 gnd.t176 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X43 CSoutput.t48 a_n6972_8799.t48 vdd.t221 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X44 a_n3106_n452.t39 minus.t7 a_n2848_n452.t44 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X45 vdd.t73 vdd.t71 vdd.t72 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X46 CSoutput.t114 commonsourceibias.t90 gnd.t323 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X47 CSoutput.t13 a_n6972_8799.t49 vdd.t220 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X48 gnd.t322 commonsourceibias.t56 commonsourceibias.t57 gnd.t252 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X49 outputibias.t3 outputibias.t2 gnd.t147 gnd.t146 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X50 output.t13 CSoutput.t155 vdd.t84 gnd.t18 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X51 a_n2140_13878.t22 a_n2848_n452.t22 a_n2848_n452.t23 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X52 CSoutput.t113 commonsourceibias.t91 gnd.t321 gnd.t300 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X53 commonsourceibias.t55 commonsourceibias.t54 gnd.t320 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X54 a_n2848_n452.t15 a_n2848_n452.t14 a_n2140_13878.t21 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X55 gnd.t128 gnd.t126 gnd.t127 gnd.t74 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X56 CSoutput.t156 a_n2318_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X57 CSoutput.t2 a_n6972_8799.t50 vdd.t219 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X58 vdd.t70 vdd.t68 vdd.t69 vdd.t51 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X59 a_n3106_n452.t22 plus.t9 a_n6972_8799.t23 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X60 vdd.t218 a_n6972_8799.t51 CSoutput.t15 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X61 diffpairibias.t15 diffpairibias.t14 gnd.t142 gnd.t141 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X62 a_n3106_n452.t21 plus.t10 a_n6972_8799.t4 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X63 a_n3106_n452.t38 minus.t8 a_n2848_n452.t43 gnd.t143 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X64 gnd.t125 gnd.t123 gnd.t124 gnd.t45 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X65 a_n6972_8799.t5 a_n2848_n452.t60 a_n2318_8322.t24 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X66 CSoutput.t143 a_n6972_8799.t52 vdd.t217 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X67 vdd.t216 a_n6972_8799.t53 CSoutput.t41 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X68 gnd.t319 commonsourceibias.t92 CSoutput.t112 gnd.t293 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X69 diffpairibias.t13 diffpairibias.t12 gnd.t339 gnd.t338 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X70 gnd.t318 commonsourceibias.t93 CSoutput.t111 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X71 CSoutput.t47 a_n6972_8799.t54 vdd.t215 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X72 output.t12 CSoutput.t157 vdd.t86 gnd.t17 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X73 commonsourceibias.t53 commonsourceibias.t52 gnd.t317 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X74 gnd.t316 commonsourceibias.t94 CSoutput.t110 gnd.t289 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X75 vdd.t214 a_n6972_8799.t55 CSoutput.t44 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X76 CSoutput.t149 a_n6972_8799.t56 vdd.t213 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X77 CSoutput.t144 a_n6972_8799.t57 vdd.t212 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X78 commonsourceibias.t51 commonsourceibias.t50 gnd.t315 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X79 gnd.t314 commonsourceibias.t95 CSoutput.t109 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 CSoutput.t11 a_n6972_8799.t58 vdd.t211 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 a_n3106_n452.t37 minus.t9 a_n2848_n452.t42 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X82 output.t11 CSoutput.t158 vdd.t81 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X83 a_n3106_n452.t20 plus.t11 a_n6972_8799.t20 gnd.t135 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X84 commonsourceibias.t49 commonsourceibias.t48 gnd.t313 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 a_n6972_8799.t36 plus.t12 a_n3106_n452.t19 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X86 gnd.t312 commonsourceibias.t96 CSoutput.t108 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X87 CSoutput.t107 commonsourceibias.t97 gnd.t311 gnd.t282 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 gnd.t310 commonsourceibias.t78 commonsourceibias.t79 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 a_n3106_n452.t35 diffpairibias.t17 gnd.t167 gnd.t166 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X90 CSoutput.t159 a_n2318_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X91 a_n2848_n452.t25 a_n2848_n452.t24 a_n2140_13878.t20 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X92 vdd.t210 a_n6972_8799.t59 CSoutput.t29 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X93 a_n3106_n452.t18 plus.t13 a_n6972_8799.t11 gnd.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X94 a_n6972_8799.t6 a_n2848_n452.t61 a_n2318_8322.t23 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X95 vdd.t209 a_n6972_8799.t60 CSoutput.t145 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X96 a_n2848_n452.t9 a_n2848_n452.t8 a_n2140_13878.t19 vdd.t3 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X97 gnd.t309 commonsourceibias.t76 commonsourceibias.t77 gnd.t274 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X98 commonsourceibias.t75 commonsourceibias.t74 gnd.t308 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X99 CSoutput.t141 commonsourceibias.t98 gnd.t307 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X100 vdd.t208 a_n6972_8799.t61 CSoutput.t142 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X101 CSoutput.t20 a_n6972_8799.t62 vdd.t207 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X102 CSoutput.t140 commonsourceibias.t99 gnd.t306 gnd.t269 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X103 a_n2848_n452.t47 minus.t10 a_n3106_n452.t42 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X104 vdd.t91 CSoutput.t160 output.t10 gnd.t15 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X105 vdd.t67 vdd.t65 vdd.t66 vdd.t55 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X106 vdd.t64 vdd.t62 vdd.t63 vdd.t17 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X107 CSoutput.t139 commonsourceibias.t100 gnd.t305 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 CSoutput.t14 a_n6972_8799.t63 vdd.t206 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X109 vdd.t61 vdd.t58 vdd.t60 vdd.t59 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X110 gnd.t304 commonsourceibias.t101 CSoutput.t138 gnd.t274 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X111 commonsourceibias.t73 commonsourceibias.t72 gnd.t303 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X112 CSoutput.t137 commonsourceibias.t102 gnd.t302 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X113 CSoutput.t136 commonsourceibias.t103 gnd.t301 gnd.t300 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X114 vdd.t98 a_n2848_n452.t62 a_n2318_8322.t11 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X115 a_n2848_n452.t13 a_n2848_n452.t12 a_n2140_13878.t18 vdd.t112 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X116 a_n2318_8322.t10 a_n2848_n452.t63 vdd.t100 vdd.t99 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X117 a_n3106_n452.t54 diffpairibias.t18 gnd.t353 gnd.t352 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X118 CSoutput.t36 a_n6972_8799.t64 vdd.t205 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X119 gnd.t299 commonsourceibias.t104 CSoutput.t135 gnd.t250 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X120 gnd.t122 gnd.t120 gnd.t121 gnd.t63 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X121 gnd.t119 gnd.t117 minus.t4 gnd.t118 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X122 commonsourceibias.t71 commonsourceibias.t70 gnd.t298 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X123 commonsourceibias.t69 commonsourceibias.t68 gnd.t297 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X124 vdd.t117 a_n2848_n452.t64 a_n2140_13878.t6 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X125 vdd.t57 vdd.t54 vdd.t56 vdd.t55 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X126 gnd.t296 commonsourceibias.t66 commonsourceibias.t67 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X127 gnd.t295 commonsourceibias.t105 CSoutput.t134 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X128 vdd.t203 a_n6972_8799.t65 CSoutput.t12 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X129 gnd.t294 commonsourceibias.t64 commonsourceibias.t65 gnd.t293 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X130 outputibias.t1 outputibias.t0 gnd.t349 gnd.t348 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X131 gnd.t116 gnd.t114 plus.t3 gnd.t115 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X132 a_n6972_8799.t13 plus.t14 a_n3106_n452.t17 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X133 a_n2848_n452.t52 minus.t11 a_n3106_n452.t47 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X134 vdd.t53 vdd.t50 vdd.t52 vdd.t51 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X135 a_n2318_8322.t9 a_n2848_n452.t65 vdd.t119 vdd.t118 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X136 commonsourceibias.t63 commonsourceibias.t62 gnd.t292 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X137 gnd.t291 commonsourceibias.t106 CSoutput.t133 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X138 gnd.t290 commonsourceibias.t107 CSoutput.t132 gnd.t289 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X139 a_n6972_8799.t26 a_n2848_n452.t66 a_n2318_8322.t22 vdd.t131 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X140 gnd.t288 commonsourceibias.t108 CSoutput.t131 gnd.t245 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X141 a_n6972_8799.t15 plus.t15 a_n3106_n452.t16 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X142 diffpairibias.t11 diffpairibias.t10 gnd.t153 gnd.t152 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X143 a_n2848_n452.t51 minus.t12 a_n3106_n452.t46 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X144 a_n2848_n452.t5 a_n2848_n452.t4 a_n2140_13878.t17 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X145 vdd.t201 a_n6972_8799.t66 CSoutput.t5 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X146 a_n6972_8799.t27 a_n2848_n452.t67 a_n2318_8322.t21 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X147 CSoutput.t28 a_n6972_8799.t67 vdd.t200 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X148 gnd.t287 commonsourceibias.t109 CSoutput.t130 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X149 output.t19 outputibias.t8 gnd.t160 gnd.t159 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X150 a_n2140_13878.t16 a_n2848_n452.t20 a_n2848_n452.t21 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X151 vdd.t49 vdd.t47 vdd.t48 vdd.t17 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X152 gnd.t286 commonsourceibias.t110 CSoutput.t129 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X153 CSoutput.t128 commonsourceibias.t111 gnd.t284 gnd.t282 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X154 commonsourceibias.t61 commonsourceibias.t60 gnd.t283 gnd.t282 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X155 a_n3106_n452.t45 minus.t13 a_n2848_n452.t50 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X156 CSoutput.t146 a_n6972_8799.t68 vdd.t199 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X157 gnd.t281 commonsourceibias.t112 CSoutput.t127 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X158 vdd.t125 a_n2848_n452.t68 a_n2318_8322.t8 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X159 CSoutput.t126 commonsourceibias.t113 gnd.t280 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X160 a_n2140_13878.t15 a_n2848_n452.t6 a_n2848_n452.t7 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X161 vdd.t198 a_n6972_8799.t69 CSoutput.t22 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X162 a_n2848_n452.t49 minus.t14 a_n3106_n452.t44 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X163 a_n3106_n452.t15 plus.t16 a_n6972_8799.t29 gnd.t149 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X164 a_n2848_n452.t33 a_n2848_n452.t32 a_n2140_13878.t14 vdd.t101 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X165 CSoutput.t125 commonsourceibias.t114 gnd.t279 gnd.t269 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X166 a_n3106_n452.t50 diffpairibias.t19 gnd.t343 gnd.t342 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X167 gnd.t113 gnd.t110 gnd.t112 gnd.t111 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X168 a_n3106_n452.t51 diffpairibias.t20 gnd.t345 gnd.t344 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X169 vdd.t89 CSoutput.t161 output.t9 gnd.t14 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X170 a_n6972_8799.t24 plus.t17 a_n3106_n452.t14 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X171 CSoutput.t124 commonsourceibias.t115 gnd.t278 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X172 CSoutput.t123 commonsourceibias.t116 gnd.t277 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X173 vdd.t197 a_n6972_8799.t70 CSoutput.t16 vdd.t159 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X174 gnd.t275 commonsourceibias.t117 CSoutput.t122 gnd.t274 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X175 gnd.t273 commonsourceibias.t118 CSoutput.t121 gnd.t252 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X176 CSoutput.t120 commonsourceibias.t119 gnd.t272 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X177 commonsourceibias.t59 commonsourceibias.t58 gnd.t270 gnd.t269 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X178 CSoutput.t119 commonsourceibias.t120 gnd.t268 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X179 gnd.t109 gnd.t107 gnd.t108 gnd.t38 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X180 a_n6972_8799.t2 plus.t18 a_n3106_n452.t13 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X181 gnd.t106 gnd.t103 gnd.t105 gnd.t104 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X182 gnd.t267 commonsourceibias.t121 CSoutput.t118 gnd.t250 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X183 CSoutput.t50 a_n6972_8799.t71 vdd.t196 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X184 minus.t3 gnd.t100 gnd.t102 gnd.t101 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X185 CSoutput.t51 a_n6972_8799.t72 vdd.t194 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X186 gnd.t99 gnd.t97 gnd.t98 gnd.t67 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X187 CSoutput.t117 commonsourceibias.t122 gnd.t266 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X188 diffpairibias.t9 diffpairibias.t8 gnd.t347 gnd.t346 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X189 a_n2140_13878.t5 a_n2848_n452.t69 vdd.t127 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X190 a_n2848_n452.t48 minus.t15 a_n3106_n452.t43 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X191 vdd.t130 a_n2848_n452.t70 a_n2140_13878.t4 vdd.t129 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X192 CSoutput.t31 a_n6972_8799.t73 vdd.t193 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X193 a_n3106_n452.t12 plus.t19 a_n6972_8799.t3 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X194 vdd.t191 a_n6972_8799.t74 CSoutput.t35 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X195 gnd.t265 commonsourceibias.t123 CSoutput.t116 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 CSoutput.t70 commonsourceibias.t124 gnd.t264 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X197 a_n2140_13878.t13 a_n2848_n452.t28 a_n2848_n452.t29 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X198 gnd.t263 commonsourceibias.t6 commonsourceibias.t7 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X199 gnd.t262 commonsourceibias.t125 CSoutput.t69 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X200 gnd.t261 commonsourceibias.t126 CSoutput.t68 gnd.t245 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X201 a_n3106_n452.t27 minus.t16 a_n2848_n452.t35 gnd.t144 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X202 gnd.t249 commonsourceibias.t127 CSoutput.t84 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X203 a_n2318_8322.t20 a_n2848_n452.t71 a_n6972_8799.t25 vdd.t80 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X204 vdd.t95 CSoutput.t162 output.t8 gnd.t13 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X205 CSoutput.t60 a_n6972_8799.t75 vdd.t189 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X206 diffpairibias.t7 diffpairibias.t6 gnd.t26 gnd.t25 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X207 CSoutput.t67 commonsourceibias.t128 gnd.t260 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X208 vdd.t188 a_n6972_8799.t76 CSoutput.t61 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X209 vdd.t121 a_n2848_n452.t72 a_n2318_8322.t7 vdd.t120 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X210 gnd.t259 commonsourceibias.t4 commonsourceibias.t5 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X211 vdd.t186 a_n6972_8799.t77 CSoutput.t42 vdd.t159 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X212 gnd.t96 gnd.t94 gnd.t95 gnd.t67 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X213 a_n3106_n452.t52 minus.t17 a_n2848_n452.t54 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X214 CSoutput.t66 commonsourceibias.t129 gnd.t258 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 a_n3106_n452.t11 plus.t20 a_n6972_8799.t9 gnd.t143 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X216 a_n3106_n452.t36 minus.t18 a_n2848_n452.t41 gnd.t168 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X217 gnd.t257 commonsourceibias.t130 CSoutput.t65 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X218 CSoutput.t64 commonsourceibias.t131 gnd.t256 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X219 a_n2140_13878.t3 a_n2848_n452.t73 vdd.t123 vdd.t122 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X220 vdd.t185 a_n6972_8799.t78 CSoutput.t53 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X221 CSoutput.t19 a_n6972_8799.t79 vdd.t184 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X222 CSoutput.t17 a_n6972_8799.t80 vdd.t183 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X223 gnd.t255 commonsourceibias.t2 commonsourceibias.t3 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X224 gnd.t93 gnd.t90 gnd.t92 gnd.t91 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X225 a_n3106_n452.t53 diffpairibias.t21 gnd.t351 gnd.t350 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X226 minus.t2 gnd.t87 gnd.t89 gnd.t88 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X227 CSoutput.t63 commonsourceibias.t132 gnd.t254 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X228 vdd.t235 a_n2848_n452.t74 a_n2318_8322.t6 vdd.t234 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X229 a_n2318_8322.t19 a_n2848_n452.t75 a_n6972_8799.t39 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X230 CSoutput.t163 a_n2318_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X231 CSoutput.t1 a_n6972_8799.t81 vdd.t182 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X232 a_n6972_8799.t8 plus.t21 a_n3106_n452.t10 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X233 vdd.t180 a_n6972_8799.t82 CSoutput.t4 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X234 vdd.t46 vdd.t44 vdd.t45 vdd.t25 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X235 a_n2848_n452.t36 minus.t19 a_n3106_n452.t28 gnd.t145 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X236 CSoutput.t83 commonsourceibias.t133 gnd.t247 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X237 CSoutput.t8 a_n6972_8799.t83 vdd.t179 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X238 a_n3106_n452.t2 minus.t20 a_n2848_n452.t34 gnd.t135 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X239 gnd.t253 commonsourceibias.t134 CSoutput.t62 gnd.t252 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X240 vdd.t178 a_n6972_8799.t84 CSoutput.t59 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X241 vdd.t177 a_n6972_8799.t85 CSoutput.t43 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X242 gnd.t251 commonsourceibias.t0 commonsourceibias.t1 gnd.t250 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X243 gnd.t246 commonsourceibias.t16 commonsourceibias.t17 gnd.t245 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X244 vdd.t94 CSoutput.t164 output.t7 gnd.t12 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X245 CSoutput.t82 commonsourceibias.t135 gnd.t244 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X246 output.t6 CSoutput.t165 vdd.t85 gnd.t11 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X247 CSoutput.t81 commonsourceibias.t136 gnd.t243 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X248 vdd.t43 vdd.t41 vdd.t42 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X249 gnd.t242 commonsourceibias.t137 CSoutput.t80 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X250 vdd.t40 vdd.t37 vdd.t39 vdd.t38 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X251 a_n3106_n452.t31 minus.t21 a_n2848_n452.t38 gnd.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X252 gnd.t86 gnd.t84 gnd.t85 gnd.t49 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X253 gnd.t83 gnd.t80 gnd.t82 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X254 a_n3106_n452.t48 minus.t22 a_n2848_n452.t53 gnd.t161 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X255 a_n2140_13878.t12 a_n2848_n452.t30 a_n2848_n452.t31 vdd.t113 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X256 CSoutput.t151 a_n6972_8799.t86 vdd.t176 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X257 gnd.t79 gnd.t77 gnd.t78 gnd.t49 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X258 CSoutput.t79 commonsourceibias.t138 gnd.t241 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X259 a_n2318_8322.t18 a_n2848_n452.t76 a_n6972_8799.t33 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X260 diffpairibias.t5 diffpairibias.t4 gnd.t171 gnd.t170 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X261 CSoutput.t166 a_n2318_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X262 commonsourceibias.t15 commonsourceibias.t14 gnd.t239 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X263 CSoutput.t56 a_n6972_8799.t87 vdd.t175 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X264 vdd.t173 a_n6972_8799.t88 CSoutput.t54 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X265 gnd.t238 commonsourceibias.t139 CSoutput.t78 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X266 CSoutput.t77 commonsourceibias.t140 gnd.t236 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X267 vdd.t172 a_n6972_8799.t89 CSoutput.t49 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X268 gnd.t76 gnd.t73 gnd.t75 gnd.t74 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X269 a_n2318_8322.t5 a_n2848_n452.t77 vdd.t231 vdd.t230 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X270 gnd.t235 commonsourceibias.t28 commonsourceibias.t29 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X271 gnd.t233 commonsourceibias.t141 CSoutput.t97 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X272 CSoutput.t37 a_n6972_8799.t90 vdd.t170 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 a_n3106_n452.t55 minus.t23 a_n2848_n452.t55 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X274 vdd.t36 vdd.t34 vdd.t35 vdd.t9 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X275 gnd.t72 gnd.t70 gnd.t71 gnd.t38 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X276 output.t18 outputibias.t9 gnd.t24 gnd.t23 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X277 CSoutput.t96 commonsourceibias.t142 gnd.t232 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 vdd.t233 a_n2848_n452.t78 a_n2140_13878.t2 vdd.t232 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X279 CSoutput.t25 a_n6972_8799.t91 vdd.t168 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X280 vdd.t33 vdd.t31 vdd.t32 vdd.t25 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X281 output.t5 CSoutput.t167 vdd.t87 gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X282 CSoutput.t58 a_n6972_8799.t92 vdd.t166 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X283 gnd.t69 gnd.t66 gnd.t68 gnd.t67 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X284 vdd.t83 CSoutput.t168 output.t4 gnd.t9 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X285 gnd.t230 commonsourceibias.t143 CSoutput.t95 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X286 gnd.t65 gnd.t62 gnd.t64 gnd.t63 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X287 CSoutput.t94 commonsourceibias.t144 gnd.t229 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X288 CSoutput.t93 commonsourceibias.t145 gnd.t228 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X289 gnd.t61 gnd.t59 plus.t2 gnd.t60 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X290 vdd.t165 a_n6972_8799.t93 CSoutput.t26 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X291 gnd.t226 commonsourceibias.t26 commonsourceibias.t27 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X292 vdd.t163 a_n6972_8799.t94 CSoutput.t34 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X293 output.t17 outputibias.t10 gnd.t140 gnd.t139 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X294 vdd.t30 vdd.t28 vdd.t29 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X295 a_n2318_8322.t17 a_n2848_n452.t79 a_n6972_8799.t38 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X296 CSoutput.t33 a_n6972_8799.t95 vdd.t162 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X297 a_n6972_8799.t19 a_n2848_n452.t80 a_n2318_8322.t16 vdd.t113 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X298 vdd.t160 a_n6972_8799.t96 CSoutput.t40 vdd.t159 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X299 a_n2140_13878.t1 a_n2848_n452.t81 vdd.t115 vdd.t114 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X300 output.t16 outputibias.t11 gnd.t341 gnd.t340 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X301 vdd.t82 CSoutput.t169 output.t3 gnd.t8 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X302 vdd.t158 a_n6972_8799.t97 CSoutput.t32 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X303 CSoutput.t27 a_n6972_8799.t98 vdd.t157 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X304 a_n3106_n452.t9 plus.t22 a_n6972_8799.t37 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X305 a_n2848_n452.t40 minus.t24 a_n3106_n452.t34 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X306 CSoutput.t92 commonsourceibias.t146 gnd.t224 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 gnd.t58 gnd.t55 gnd.t57 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X308 a_n6972_8799.t0 plus.t23 a_n3106_n452.t8 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X309 gnd.t54 gnd.t52 minus.t1 gnd.t53 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X310 vdd.t27 vdd.t24 vdd.t26 vdd.t25 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X311 a_n2318_8322.t15 a_n2848_n452.t82 a_n6972_8799.t21 vdd.t112 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X312 vdd.t23 vdd.t20 vdd.t22 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X313 a_n2848_n452.t0 minus.t25 a_n3106_n452.t0 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X314 output.t2 CSoutput.t170 vdd.t92 gnd.t7 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X315 a_n2140_13878.t11 a_n2848_n452.t26 a_n2848_n452.t27 vdd.t131 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X316 commonsourceibias.t25 commonsourceibias.t24 gnd.t222 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X317 gnd.t220 commonsourceibias.t147 CSoutput.t91 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X318 vdd.t155 a_n6972_8799.t99 CSoutput.t46 vdd.t140 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X319 gnd.t219 commonsourceibias.t12 commonsourceibias.t13 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X320 vdd.t19 vdd.t16 vdd.t18 vdd.t17 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X321 CSoutput.t76 commonsourceibias.t148 gnd.t218 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X322 gnd.t216 commonsourceibias.t149 CSoutput.t75 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X323 vdd.t15 vdd.t12 vdd.t14 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X324 a_n3106_n452.t29 minus.t26 a_n2848_n452.t37 gnd.t149 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X325 a_n3106_n452.t30 diffpairibias.t22 gnd.t151 gnd.t150 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X326 output.t1 CSoutput.t171 vdd.t90 gnd.t6 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X327 gnd.t214 commonsourceibias.t150 CSoutput.t74 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X328 vdd.t154 a_n6972_8799.t100 CSoutput.t9 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X329 gnd.t51 gnd.t48 gnd.t50 gnd.t49 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X330 gnd.t212 commonsourceibias.t151 CSoutput.t73 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X331 a_n2848_n452.t17 a_n2848_n452.t16 a_n2140_13878.t10 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X332 commonsourceibias.t11 commonsourceibias.t10 gnd.t210 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X333 a_n6972_8799.t22 a_n2848_n452.t83 a_n2318_8322.t14 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X334 gnd.t47 gnd.t44 gnd.t46 gnd.t45 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X335 a_n6972_8799.t32 plus.t24 a_n3106_n452.t7 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X336 gnd.t209 commonsourceibias.t152 CSoutput.t72 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X337 vdd.t153 a_n6972_8799.t101 CSoutput.t57 vdd.t140 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X338 CSoutput.t38 a_n6972_8799.t102 vdd.t152 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X339 vdd.t150 a_n6972_8799.t103 CSoutput.t7 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X340 diffpairibias.t3 diffpairibias.t2 gnd.t156 gnd.t155 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X341 vdd.t149 a_n6972_8799.t104 CSoutput.t18 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X342 CSoutput.t23 a_n6972_8799.t105 vdd.t147 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X343 a_n2318_8322.t13 a_n2848_n452.t84 a_n6972_8799.t7 vdd.t101 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X344 a_n2848_n452.t1 minus.t27 a_n3106_n452.t1 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X345 gnd.t43 gnd.t41 plus.t1 gnd.t42 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X346 commonsourceibias.t9 commonsourceibias.t8 gnd.t207 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X347 vdd.t145 a_n6972_8799.t106 CSoutput.t6 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X348 gnd.t205 commonsourceibias.t153 CSoutput.t71 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X349 diffpairibias.t1 diffpairibias.t0 gnd.t355 gnd.t354 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X350 CSoutput.t172 a_n2318_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X351 gnd.t40 gnd.t37 gnd.t39 gnd.t38 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X352 CSoutput.t90 commonsourceibias.t154 gnd.t203 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X353 vdd.t11 vdd.t8 vdd.t10 vdd.t9 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X354 vdd.t103 a_n2848_n452.t85 a_n2140_13878.t0 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X355 commonsourceibias.t23 commonsourceibias.t22 gnd.t201 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X356 gnd.t36 gnd.t33 gnd.t35 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X357 gnd.t200 commonsourceibias.t155 CSoutput.t89 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X358 vdd.t7 vdd.t4 vdd.t6 vdd.t5 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X359 CSoutput.t88 commonsourceibias.t156 gnd.t199 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X360 CSoutput.t87 commonsourceibias.t157 gnd.t197 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X361 plus.t0 gnd.t30 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X362 vdd.t143 a_n6972_8799.t107 CSoutput.t30 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X363 commonsourceibias.t21 commonsourceibias.t20 gnd.t195 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X364 vdd.t141 a_n6972_8799.t108 CSoutput.t3 vdd.t140 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X365 CSoutput.t86 commonsourceibias.t158 gnd.t193 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X366 CSoutput.t148 a_n6972_8799.t109 vdd.t139 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X367 gnd.t191 commonsourceibias.t18 commonsourceibias.t19 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X368 vdd.t96 CSoutput.t173 output.t0 gnd.t5 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X369 a_n6972_8799.t18 plus.t25 a_n3106_n452.t6 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X370 gnd.t29 gnd.t27 minus.t0 gnd.t28 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X371 a_n2848_n452.t39 minus.t28 a_n3106_n452.t33 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X372 CSoutput.t85 commonsourceibias.t159 gnd.t189 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X373 a_n6972_8799.t28 plus.t26 a_n3106_n452.t5 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X374 a_n2318_8322.t12 a_n2848_n452.t86 a_n6972_8799.t17 vdd.t3 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X375 gnd.t187 commonsourceibias.t38 commonsourceibias.t39 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X376 vdd.t137 a_n6972_8799.t110 CSoutput.t55 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X377 commonsourceibias.t37 commonsourceibias.t36 gnd.t185 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X378 gnd.t183 commonsourceibias.t34 commonsourceibias.t35 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X379 a_n2318_8322.t4 a_n2848_n452.t87 vdd.t111 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X380 a_n2140_13878.t9 a_n2848_n452.t2 a_n2848_n452.t3 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X381 vdd.t135 a_n6972_8799.t111 CSoutput.t147 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X382 commonsourceibias.t33 commonsourceibias.t32 gnd.t181 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X383 a_n3106_n452.t4 plus.t27 a_n6972_8799.t10 gnd.t144 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X384 a_n3106_n452.t32 diffpairibias.t23 gnd.t164 gnd.t163 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X385 gnd.t179 commonsourceibias.t30 commonsourceibias.t31 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X386 a_n2848_n452.t11 a_n2848_n452.t10 a_n2140_13878.t8 vdd.t80 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X387 a_n3106_n452.t3 plus.t28 a_n6972_8799.t1 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
R0 commonsourceibias.n281 commonsourceibias.t102 222.032
R1 commonsourceibias.n44 commonsourceibias.t54 222.032
R2 commonsourceibias.n166 commonsourceibias.t119 222.032
R3 commonsourceibias.n643 commonsourceibias.t108 222.032
R4 commonsourceibias.n413 commonsourceibias.t16 222.032
R5 commonsourceibias.n529 commonsourceibias.t126 222.032
R6 commonsourceibias.n364 commonsourceibias.t101 207.983
R7 commonsourceibias.n127 commonsourceibias.t76 207.983
R8 commonsourceibias.n249 commonsourceibias.t117 207.983
R9 commonsourceibias.n731 commonsourceibias.t124 207.983
R10 commonsourceibias.n501 commonsourceibias.t32 207.983
R11 commonsourceibias.n616 commonsourceibias.t140 207.983
R12 commonsourceibias.n280 commonsourceibias.t152 168.701
R13 commonsourceibias.n286 commonsourceibias.t157 168.701
R14 commonsourceibias.n292 commonsourceibias.t112 168.701
R15 commonsourceibias.n276 commonsourceibias.t97 168.701
R16 commonsourceibias.n300 commonsourceibias.t85 168.701
R17 commonsourceibias.n306 commonsourceibias.t122 168.701
R18 commonsourceibias.n271 commonsourceibias.t104 168.701
R19 commonsourceibias.n314 commonsourceibias.t91 168.701
R20 commonsourceibias.n320 commonsourceibias.t94 168.701
R21 commonsourceibias.n266 commonsourceibias.t113 168.701
R22 commonsourceibias.n328 commonsourceibias.t96 168.701
R23 commonsourceibias.n334 commonsourceibias.t100 168.701
R24 commonsourceibias.n261 commonsourceibias.t151 168.701
R25 commonsourceibias.n342 commonsourceibias.t129 168.701
R26 commonsourceibias.n348 commonsourceibias.t109 168.701
R27 commonsourceibias.n256 commonsourceibias.t159 168.701
R28 commonsourceibias.n356 commonsourceibias.t81 168.701
R29 commonsourceibias.n362 commonsourceibias.t120 168.701
R30 commonsourceibias.n125 commonsourceibias.t24 168.701
R31 commonsourceibias.n119 commonsourceibias.t64 168.701
R32 commonsourceibias.n19 commonsourceibias.t74 168.701
R33 commonsourceibias.n111 commonsourceibias.t4 168.701
R34 commonsourceibias.n105 commonsourceibias.t48 168.701
R35 commonsourceibias.n24 commonsourceibias.t44 168.701
R36 commonsourceibias.n97 commonsourceibias.t70 168.701
R37 commonsourceibias.n91 commonsourceibias.t78 168.701
R38 commonsourceibias.n29 commonsourceibias.t8 168.701
R39 commonsourceibias.n83 commonsourceibias.t40 168.701
R40 commonsourceibias.n77 commonsourceibias.t46 168.701
R41 commonsourceibias.n34 commonsourceibias.t0 168.701
R42 commonsourceibias.n69 commonsourceibias.t50 168.701
R43 commonsourceibias.n63 commonsourceibias.t26 168.701
R44 commonsourceibias.n39 commonsourceibias.t60 168.701
R45 commonsourceibias.n55 commonsourceibias.t34 168.701
R46 commonsourceibias.n49 commonsourceibias.t22 168.701
R47 commonsourceibias.n43 commonsourceibias.t12 168.701
R48 commonsourceibias.n247 commonsourceibias.t135 168.701
R49 commonsourceibias.n241 commonsourceibias.t92 168.701
R50 commonsourceibias.n5 commonsourceibias.t90 168.701
R51 commonsourceibias.n233 commonsourceibias.t127 168.701
R52 commonsourceibias.n227 commonsourceibias.t145 168.701
R53 commonsourceibias.n10 commonsourceibias.t83 168.701
R54 commonsourceibias.n219 commonsourceibias.t116 168.701
R55 commonsourceibias.n213 commonsourceibias.t110 168.701
R56 commonsourceibias.n150 commonsourceibias.t131 168.701
R57 commonsourceibias.n151 commonsourceibias.t107 168.701
R58 commonsourceibias.n153 commonsourceibias.t103 168.701
R59 commonsourceibias.n155 commonsourceibias.t121 168.701
R60 commonsourceibias.n191 commonsourceibias.t138 168.701
R61 commonsourceibias.n185 commonsourceibias.t95 168.701
R62 commonsourceibias.n161 commonsourceibias.t111 168.701
R63 commonsourceibias.n177 commonsourceibias.t130 168.701
R64 commonsourceibias.n171 commonsourceibias.t87 168.701
R65 commonsourceibias.n165 commonsourceibias.t84 168.701
R66 commonsourceibias.n642 commonsourceibias.t158 168.701
R67 commonsourceibias.n648 commonsourceibias.t150 168.701
R68 commonsourceibias.n654 commonsourceibias.t136 168.701
R69 commonsourceibias.n656 commonsourceibias.t118 168.701
R70 commonsourceibias.n663 commonsourceibias.t99 168.701
R71 commonsourceibias.n669 commonsourceibias.t143 168.701
R72 commonsourceibias.n671 commonsourceibias.t128 168.701
R73 commonsourceibias.n678 commonsourceibias.t106 168.701
R74 commonsourceibias.n684 commonsourceibias.t88 168.701
R75 commonsourceibias.n686 commonsourceibias.t137 168.701
R76 commonsourceibias.n693 commonsourceibias.t115 168.701
R77 commonsourceibias.n699 commonsourceibias.t123 168.701
R78 commonsourceibias.n701 commonsourceibias.t144 168.701
R79 commonsourceibias.n708 commonsourceibias.t147 168.701
R80 commonsourceibias.n714 commonsourceibias.t132 168.701
R81 commonsourceibias.n716 commonsourceibias.t93 168.701
R82 commonsourceibias.n723 commonsourceibias.t154 168.701
R83 commonsourceibias.n729 commonsourceibias.t141 168.701
R84 commonsourceibias.n412 commonsourceibias.t68 168.701
R85 commonsourceibias.n418 commonsourceibias.t66 168.701
R86 commonsourceibias.n424 commonsourceibias.t14 168.701
R87 commonsourceibias.n426 commonsourceibias.t56 168.701
R88 commonsourceibias.n433 commonsourceibias.t58 168.701
R89 commonsourceibias.n439 commonsourceibias.t18 168.701
R90 commonsourceibias.n441 commonsourceibias.t62 168.701
R91 commonsourceibias.n448 commonsourceibias.t28 168.701
R92 commonsourceibias.n454 commonsourceibias.t20 168.701
R93 commonsourceibias.n456 commonsourceibias.t2 168.701
R94 commonsourceibias.n463 commonsourceibias.t36 168.701
R95 commonsourceibias.n469 commonsourceibias.t42 168.701
R96 commonsourceibias.n471 commonsourceibias.t10 168.701
R97 commonsourceibias.n478 commonsourceibias.t38 168.701
R98 commonsourceibias.n484 commonsourceibias.t72 168.701
R99 commonsourceibias.n486 commonsourceibias.t30 168.701
R100 commonsourceibias.n493 commonsourceibias.t52 168.701
R101 commonsourceibias.n499 commonsourceibias.t6 168.701
R102 commonsourceibias.n614 commonsourceibias.t153 168.701
R103 commonsourceibias.n608 commonsourceibias.t86 168.701
R104 commonsourceibias.n601 commonsourceibias.t105 168.701
R105 commonsourceibias.n599 commonsourceibias.t146 168.701
R106 commonsourceibias.n593 commonsourceibias.t80 168.701
R107 commonsourceibias.n586 commonsourceibias.t156 168.701
R108 commonsourceibias.n584 commonsourceibias.t139 168.701
R109 commonsourceibias.n578 commonsourceibias.t133 168.701
R110 commonsourceibias.n571 commonsourceibias.t149 168.701
R111 commonsourceibias.n528 commonsourceibias.t89 168.701
R112 commonsourceibias.n534 commonsourceibias.t82 168.701
R113 commonsourceibias.n540 commonsourceibias.t148 168.701
R114 commonsourceibias.n542 commonsourceibias.t134 168.701
R115 commonsourceibias.n549 commonsourceibias.t114 168.701
R116 commonsourceibias.n555 commonsourceibias.t155 168.701
R117 commonsourceibias.n519 commonsourceibias.t142 168.701
R118 commonsourceibias.n517 commonsourceibias.t125 168.701
R119 commonsourceibias.n515 commonsourceibias.t98 168.701
R120 commonsourceibias.n363 commonsourceibias.n251 161.3
R121 commonsourceibias.n361 commonsourceibias.n360 161.3
R122 commonsourceibias.n359 commonsourceibias.n252 161.3
R123 commonsourceibias.n358 commonsourceibias.n357 161.3
R124 commonsourceibias.n355 commonsourceibias.n253 161.3
R125 commonsourceibias.n354 commonsourceibias.n353 161.3
R126 commonsourceibias.n352 commonsourceibias.n254 161.3
R127 commonsourceibias.n351 commonsourceibias.n350 161.3
R128 commonsourceibias.n349 commonsourceibias.n255 161.3
R129 commonsourceibias.n347 commonsourceibias.n346 161.3
R130 commonsourceibias.n345 commonsourceibias.n257 161.3
R131 commonsourceibias.n344 commonsourceibias.n343 161.3
R132 commonsourceibias.n341 commonsourceibias.n258 161.3
R133 commonsourceibias.n340 commonsourceibias.n339 161.3
R134 commonsourceibias.n338 commonsourceibias.n259 161.3
R135 commonsourceibias.n337 commonsourceibias.n336 161.3
R136 commonsourceibias.n335 commonsourceibias.n260 161.3
R137 commonsourceibias.n333 commonsourceibias.n332 161.3
R138 commonsourceibias.n331 commonsourceibias.n262 161.3
R139 commonsourceibias.n330 commonsourceibias.n329 161.3
R140 commonsourceibias.n327 commonsourceibias.n263 161.3
R141 commonsourceibias.n326 commonsourceibias.n325 161.3
R142 commonsourceibias.n324 commonsourceibias.n264 161.3
R143 commonsourceibias.n323 commonsourceibias.n322 161.3
R144 commonsourceibias.n321 commonsourceibias.n265 161.3
R145 commonsourceibias.n319 commonsourceibias.n318 161.3
R146 commonsourceibias.n317 commonsourceibias.n267 161.3
R147 commonsourceibias.n316 commonsourceibias.n315 161.3
R148 commonsourceibias.n313 commonsourceibias.n268 161.3
R149 commonsourceibias.n312 commonsourceibias.n311 161.3
R150 commonsourceibias.n310 commonsourceibias.n269 161.3
R151 commonsourceibias.n309 commonsourceibias.n308 161.3
R152 commonsourceibias.n307 commonsourceibias.n270 161.3
R153 commonsourceibias.n305 commonsourceibias.n304 161.3
R154 commonsourceibias.n303 commonsourceibias.n272 161.3
R155 commonsourceibias.n302 commonsourceibias.n301 161.3
R156 commonsourceibias.n299 commonsourceibias.n273 161.3
R157 commonsourceibias.n298 commonsourceibias.n297 161.3
R158 commonsourceibias.n296 commonsourceibias.n274 161.3
R159 commonsourceibias.n295 commonsourceibias.n294 161.3
R160 commonsourceibias.n293 commonsourceibias.n275 161.3
R161 commonsourceibias.n291 commonsourceibias.n290 161.3
R162 commonsourceibias.n289 commonsourceibias.n277 161.3
R163 commonsourceibias.n288 commonsourceibias.n287 161.3
R164 commonsourceibias.n285 commonsourceibias.n278 161.3
R165 commonsourceibias.n284 commonsourceibias.n283 161.3
R166 commonsourceibias.n282 commonsourceibias.n279 161.3
R167 commonsourceibias.n45 commonsourceibias.n42 161.3
R168 commonsourceibias.n47 commonsourceibias.n46 161.3
R169 commonsourceibias.n48 commonsourceibias.n41 161.3
R170 commonsourceibias.n51 commonsourceibias.n50 161.3
R171 commonsourceibias.n52 commonsourceibias.n40 161.3
R172 commonsourceibias.n54 commonsourceibias.n53 161.3
R173 commonsourceibias.n56 commonsourceibias.n38 161.3
R174 commonsourceibias.n58 commonsourceibias.n57 161.3
R175 commonsourceibias.n59 commonsourceibias.n37 161.3
R176 commonsourceibias.n61 commonsourceibias.n60 161.3
R177 commonsourceibias.n62 commonsourceibias.n36 161.3
R178 commonsourceibias.n65 commonsourceibias.n64 161.3
R179 commonsourceibias.n66 commonsourceibias.n35 161.3
R180 commonsourceibias.n68 commonsourceibias.n67 161.3
R181 commonsourceibias.n70 commonsourceibias.n33 161.3
R182 commonsourceibias.n72 commonsourceibias.n71 161.3
R183 commonsourceibias.n73 commonsourceibias.n32 161.3
R184 commonsourceibias.n75 commonsourceibias.n74 161.3
R185 commonsourceibias.n76 commonsourceibias.n31 161.3
R186 commonsourceibias.n79 commonsourceibias.n78 161.3
R187 commonsourceibias.n80 commonsourceibias.n30 161.3
R188 commonsourceibias.n82 commonsourceibias.n81 161.3
R189 commonsourceibias.n84 commonsourceibias.n28 161.3
R190 commonsourceibias.n86 commonsourceibias.n85 161.3
R191 commonsourceibias.n87 commonsourceibias.n27 161.3
R192 commonsourceibias.n89 commonsourceibias.n88 161.3
R193 commonsourceibias.n90 commonsourceibias.n26 161.3
R194 commonsourceibias.n93 commonsourceibias.n92 161.3
R195 commonsourceibias.n94 commonsourceibias.n25 161.3
R196 commonsourceibias.n96 commonsourceibias.n95 161.3
R197 commonsourceibias.n98 commonsourceibias.n23 161.3
R198 commonsourceibias.n100 commonsourceibias.n99 161.3
R199 commonsourceibias.n101 commonsourceibias.n22 161.3
R200 commonsourceibias.n103 commonsourceibias.n102 161.3
R201 commonsourceibias.n104 commonsourceibias.n21 161.3
R202 commonsourceibias.n107 commonsourceibias.n106 161.3
R203 commonsourceibias.n108 commonsourceibias.n20 161.3
R204 commonsourceibias.n110 commonsourceibias.n109 161.3
R205 commonsourceibias.n112 commonsourceibias.n18 161.3
R206 commonsourceibias.n114 commonsourceibias.n113 161.3
R207 commonsourceibias.n115 commonsourceibias.n17 161.3
R208 commonsourceibias.n117 commonsourceibias.n116 161.3
R209 commonsourceibias.n118 commonsourceibias.n16 161.3
R210 commonsourceibias.n121 commonsourceibias.n120 161.3
R211 commonsourceibias.n122 commonsourceibias.n15 161.3
R212 commonsourceibias.n124 commonsourceibias.n123 161.3
R213 commonsourceibias.n126 commonsourceibias.n14 161.3
R214 commonsourceibias.n167 commonsourceibias.n164 161.3
R215 commonsourceibias.n169 commonsourceibias.n168 161.3
R216 commonsourceibias.n170 commonsourceibias.n163 161.3
R217 commonsourceibias.n173 commonsourceibias.n172 161.3
R218 commonsourceibias.n174 commonsourceibias.n162 161.3
R219 commonsourceibias.n176 commonsourceibias.n175 161.3
R220 commonsourceibias.n178 commonsourceibias.n160 161.3
R221 commonsourceibias.n180 commonsourceibias.n179 161.3
R222 commonsourceibias.n181 commonsourceibias.n159 161.3
R223 commonsourceibias.n183 commonsourceibias.n182 161.3
R224 commonsourceibias.n184 commonsourceibias.n158 161.3
R225 commonsourceibias.n187 commonsourceibias.n186 161.3
R226 commonsourceibias.n188 commonsourceibias.n157 161.3
R227 commonsourceibias.n190 commonsourceibias.n189 161.3
R228 commonsourceibias.n192 commonsourceibias.n156 161.3
R229 commonsourceibias.n194 commonsourceibias.n193 161.3
R230 commonsourceibias.n196 commonsourceibias.n195 161.3
R231 commonsourceibias.n197 commonsourceibias.n154 161.3
R232 commonsourceibias.n199 commonsourceibias.n198 161.3
R233 commonsourceibias.n201 commonsourceibias.n200 161.3
R234 commonsourceibias.n202 commonsourceibias.n152 161.3
R235 commonsourceibias.n204 commonsourceibias.n203 161.3
R236 commonsourceibias.n206 commonsourceibias.n205 161.3
R237 commonsourceibias.n208 commonsourceibias.n207 161.3
R238 commonsourceibias.n209 commonsourceibias.n13 161.3
R239 commonsourceibias.n211 commonsourceibias.n210 161.3
R240 commonsourceibias.n212 commonsourceibias.n12 161.3
R241 commonsourceibias.n215 commonsourceibias.n214 161.3
R242 commonsourceibias.n216 commonsourceibias.n11 161.3
R243 commonsourceibias.n218 commonsourceibias.n217 161.3
R244 commonsourceibias.n220 commonsourceibias.n9 161.3
R245 commonsourceibias.n222 commonsourceibias.n221 161.3
R246 commonsourceibias.n223 commonsourceibias.n8 161.3
R247 commonsourceibias.n225 commonsourceibias.n224 161.3
R248 commonsourceibias.n226 commonsourceibias.n7 161.3
R249 commonsourceibias.n229 commonsourceibias.n228 161.3
R250 commonsourceibias.n230 commonsourceibias.n6 161.3
R251 commonsourceibias.n232 commonsourceibias.n231 161.3
R252 commonsourceibias.n234 commonsourceibias.n4 161.3
R253 commonsourceibias.n236 commonsourceibias.n235 161.3
R254 commonsourceibias.n237 commonsourceibias.n3 161.3
R255 commonsourceibias.n239 commonsourceibias.n238 161.3
R256 commonsourceibias.n240 commonsourceibias.n2 161.3
R257 commonsourceibias.n243 commonsourceibias.n242 161.3
R258 commonsourceibias.n244 commonsourceibias.n1 161.3
R259 commonsourceibias.n246 commonsourceibias.n245 161.3
R260 commonsourceibias.n248 commonsourceibias.n0 161.3
R261 commonsourceibias.n730 commonsourceibias.n618 161.3
R262 commonsourceibias.n728 commonsourceibias.n727 161.3
R263 commonsourceibias.n726 commonsourceibias.n619 161.3
R264 commonsourceibias.n725 commonsourceibias.n724 161.3
R265 commonsourceibias.n722 commonsourceibias.n620 161.3
R266 commonsourceibias.n721 commonsourceibias.n720 161.3
R267 commonsourceibias.n719 commonsourceibias.n621 161.3
R268 commonsourceibias.n718 commonsourceibias.n717 161.3
R269 commonsourceibias.n715 commonsourceibias.n622 161.3
R270 commonsourceibias.n713 commonsourceibias.n712 161.3
R271 commonsourceibias.n711 commonsourceibias.n623 161.3
R272 commonsourceibias.n710 commonsourceibias.n709 161.3
R273 commonsourceibias.n707 commonsourceibias.n624 161.3
R274 commonsourceibias.n706 commonsourceibias.n705 161.3
R275 commonsourceibias.n704 commonsourceibias.n625 161.3
R276 commonsourceibias.n703 commonsourceibias.n702 161.3
R277 commonsourceibias.n700 commonsourceibias.n626 161.3
R278 commonsourceibias.n698 commonsourceibias.n697 161.3
R279 commonsourceibias.n696 commonsourceibias.n627 161.3
R280 commonsourceibias.n695 commonsourceibias.n694 161.3
R281 commonsourceibias.n692 commonsourceibias.n628 161.3
R282 commonsourceibias.n691 commonsourceibias.n690 161.3
R283 commonsourceibias.n689 commonsourceibias.n629 161.3
R284 commonsourceibias.n688 commonsourceibias.n687 161.3
R285 commonsourceibias.n685 commonsourceibias.n630 161.3
R286 commonsourceibias.n683 commonsourceibias.n682 161.3
R287 commonsourceibias.n681 commonsourceibias.n631 161.3
R288 commonsourceibias.n680 commonsourceibias.n679 161.3
R289 commonsourceibias.n677 commonsourceibias.n632 161.3
R290 commonsourceibias.n676 commonsourceibias.n675 161.3
R291 commonsourceibias.n674 commonsourceibias.n633 161.3
R292 commonsourceibias.n673 commonsourceibias.n672 161.3
R293 commonsourceibias.n670 commonsourceibias.n634 161.3
R294 commonsourceibias.n668 commonsourceibias.n667 161.3
R295 commonsourceibias.n666 commonsourceibias.n635 161.3
R296 commonsourceibias.n665 commonsourceibias.n664 161.3
R297 commonsourceibias.n662 commonsourceibias.n636 161.3
R298 commonsourceibias.n661 commonsourceibias.n660 161.3
R299 commonsourceibias.n659 commonsourceibias.n637 161.3
R300 commonsourceibias.n658 commonsourceibias.n657 161.3
R301 commonsourceibias.n655 commonsourceibias.n638 161.3
R302 commonsourceibias.n653 commonsourceibias.n652 161.3
R303 commonsourceibias.n651 commonsourceibias.n639 161.3
R304 commonsourceibias.n650 commonsourceibias.n649 161.3
R305 commonsourceibias.n647 commonsourceibias.n640 161.3
R306 commonsourceibias.n646 commonsourceibias.n645 161.3
R307 commonsourceibias.n644 commonsourceibias.n641 161.3
R308 commonsourceibias.n500 commonsourceibias.n388 161.3
R309 commonsourceibias.n498 commonsourceibias.n497 161.3
R310 commonsourceibias.n496 commonsourceibias.n389 161.3
R311 commonsourceibias.n495 commonsourceibias.n494 161.3
R312 commonsourceibias.n492 commonsourceibias.n390 161.3
R313 commonsourceibias.n491 commonsourceibias.n490 161.3
R314 commonsourceibias.n489 commonsourceibias.n391 161.3
R315 commonsourceibias.n488 commonsourceibias.n487 161.3
R316 commonsourceibias.n485 commonsourceibias.n392 161.3
R317 commonsourceibias.n483 commonsourceibias.n482 161.3
R318 commonsourceibias.n481 commonsourceibias.n393 161.3
R319 commonsourceibias.n480 commonsourceibias.n479 161.3
R320 commonsourceibias.n477 commonsourceibias.n394 161.3
R321 commonsourceibias.n476 commonsourceibias.n475 161.3
R322 commonsourceibias.n474 commonsourceibias.n395 161.3
R323 commonsourceibias.n473 commonsourceibias.n472 161.3
R324 commonsourceibias.n470 commonsourceibias.n396 161.3
R325 commonsourceibias.n468 commonsourceibias.n467 161.3
R326 commonsourceibias.n466 commonsourceibias.n397 161.3
R327 commonsourceibias.n465 commonsourceibias.n464 161.3
R328 commonsourceibias.n462 commonsourceibias.n398 161.3
R329 commonsourceibias.n461 commonsourceibias.n460 161.3
R330 commonsourceibias.n459 commonsourceibias.n399 161.3
R331 commonsourceibias.n458 commonsourceibias.n457 161.3
R332 commonsourceibias.n455 commonsourceibias.n400 161.3
R333 commonsourceibias.n453 commonsourceibias.n452 161.3
R334 commonsourceibias.n451 commonsourceibias.n401 161.3
R335 commonsourceibias.n450 commonsourceibias.n449 161.3
R336 commonsourceibias.n447 commonsourceibias.n402 161.3
R337 commonsourceibias.n446 commonsourceibias.n445 161.3
R338 commonsourceibias.n444 commonsourceibias.n403 161.3
R339 commonsourceibias.n443 commonsourceibias.n442 161.3
R340 commonsourceibias.n440 commonsourceibias.n404 161.3
R341 commonsourceibias.n438 commonsourceibias.n437 161.3
R342 commonsourceibias.n436 commonsourceibias.n405 161.3
R343 commonsourceibias.n435 commonsourceibias.n434 161.3
R344 commonsourceibias.n432 commonsourceibias.n406 161.3
R345 commonsourceibias.n431 commonsourceibias.n430 161.3
R346 commonsourceibias.n429 commonsourceibias.n407 161.3
R347 commonsourceibias.n428 commonsourceibias.n427 161.3
R348 commonsourceibias.n425 commonsourceibias.n408 161.3
R349 commonsourceibias.n423 commonsourceibias.n422 161.3
R350 commonsourceibias.n421 commonsourceibias.n409 161.3
R351 commonsourceibias.n420 commonsourceibias.n419 161.3
R352 commonsourceibias.n417 commonsourceibias.n410 161.3
R353 commonsourceibias.n416 commonsourceibias.n415 161.3
R354 commonsourceibias.n414 commonsourceibias.n411 161.3
R355 commonsourceibias.n570 commonsourceibias.n569 161.3
R356 commonsourceibias.n568 commonsourceibias.n567 161.3
R357 commonsourceibias.n566 commonsourceibias.n516 161.3
R358 commonsourceibias.n565 commonsourceibias.n564 161.3
R359 commonsourceibias.n563 commonsourceibias.n562 161.3
R360 commonsourceibias.n561 commonsourceibias.n518 161.3
R361 commonsourceibias.n560 commonsourceibias.n559 161.3
R362 commonsourceibias.n558 commonsourceibias.n557 161.3
R363 commonsourceibias.n556 commonsourceibias.n520 161.3
R364 commonsourceibias.n554 commonsourceibias.n553 161.3
R365 commonsourceibias.n552 commonsourceibias.n521 161.3
R366 commonsourceibias.n551 commonsourceibias.n550 161.3
R367 commonsourceibias.n548 commonsourceibias.n522 161.3
R368 commonsourceibias.n547 commonsourceibias.n546 161.3
R369 commonsourceibias.n545 commonsourceibias.n523 161.3
R370 commonsourceibias.n544 commonsourceibias.n543 161.3
R371 commonsourceibias.n541 commonsourceibias.n524 161.3
R372 commonsourceibias.n539 commonsourceibias.n538 161.3
R373 commonsourceibias.n537 commonsourceibias.n525 161.3
R374 commonsourceibias.n536 commonsourceibias.n535 161.3
R375 commonsourceibias.n533 commonsourceibias.n526 161.3
R376 commonsourceibias.n532 commonsourceibias.n531 161.3
R377 commonsourceibias.n530 commonsourceibias.n527 161.3
R378 commonsourceibias.n615 commonsourceibias.n367 161.3
R379 commonsourceibias.n613 commonsourceibias.n612 161.3
R380 commonsourceibias.n611 commonsourceibias.n368 161.3
R381 commonsourceibias.n610 commonsourceibias.n609 161.3
R382 commonsourceibias.n607 commonsourceibias.n369 161.3
R383 commonsourceibias.n606 commonsourceibias.n605 161.3
R384 commonsourceibias.n604 commonsourceibias.n370 161.3
R385 commonsourceibias.n603 commonsourceibias.n602 161.3
R386 commonsourceibias.n600 commonsourceibias.n371 161.3
R387 commonsourceibias.n598 commonsourceibias.n597 161.3
R388 commonsourceibias.n596 commonsourceibias.n372 161.3
R389 commonsourceibias.n595 commonsourceibias.n594 161.3
R390 commonsourceibias.n592 commonsourceibias.n373 161.3
R391 commonsourceibias.n591 commonsourceibias.n590 161.3
R392 commonsourceibias.n589 commonsourceibias.n374 161.3
R393 commonsourceibias.n588 commonsourceibias.n587 161.3
R394 commonsourceibias.n585 commonsourceibias.n375 161.3
R395 commonsourceibias.n583 commonsourceibias.n582 161.3
R396 commonsourceibias.n581 commonsourceibias.n376 161.3
R397 commonsourceibias.n580 commonsourceibias.n579 161.3
R398 commonsourceibias.n577 commonsourceibias.n377 161.3
R399 commonsourceibias.n576 commonsourceibias.n575 161.3
R400 commonsourceibias.n574 commonsourceibias.n378 161.3
R401 commonsourceibias.n573 commonsourceibias.n572 161.3
R402 commonsourceibias.n141 commonsourceibias.n139 81.5057
R403 commonsourceibias.n381 commonsourceibias.n379 81.5057
R404 commonsourceibias.n141 commonsourceibias.n140 80.9324
R405 commonsourceibias.n143 commonsourceibias.n142 80.9324
R406 commonsourceibias.n145 commonsourceibias.n144 80.9324
R407 commonsourceibias.n147 commonsourceibias.n146 80.9324
R408 commonsourceibias.n138 commonsourceibias.n137 80.9324
R409 commonsourceibias.n136 commonsourceibias.n135 80.9324
R410 commonsourceibias.n134 commonsourceibias.n133 80.9324
R411 commonsourceibias.n132 commonsourceibias.n131 80.9324
R412 commonsourceibias.n130 commonsourceibias.n129 80.9324
R413 commonsourceibias.n504 commonsourceibias.n503 80.9324
R414 commonsourceibias.n506 commonsourceibias.n505 80.9324
R415 commonsourceibias.n508 commonsourceibias.n507 80.9324
R416 commonsourceibias.n510 commonsourceibias.n509 80.9324
R417 commonsourceibias.n512 commonsourceibias.n511 80.9324
R418 commonsourceibias.n387 commonsourceibias.n386 80.9324
R419 commonsourceibias.n385 commonsourceibias.n384 80.9324
R420 commonsourceibias.n383 commonsourceibias.n382 80.9324
R421 commonsourceibias.n381 commonsourceibias.n380 80.9324
R422 commonsourceibias.n365 commonsourceibias.n364 80.6037
R423 commonsourceibias.n128 commonsourceibias.n127 80.6037
R424 commonsourceibias.n250 commonsourceibias.n249 80.6037
R425 commonsourceibias.n732 commonsourceibias.n731 80.6037
R426 commonsourceibias.n502 commonsourceibias.n501 80.6037
R427 commonsourceibias.n617 commonsourceibias.n616 80.6037
R428 commonsourceibias.n322 commonsourceibias.n321 56.5617
R429 commonsourceibias.n336 commonsourceibias.n335 56.5617
R430 commonsourceibias.n85 commonsourceibias.n84 56.5617
R431 commonsourceibias.n71 commonsourceibias.n70 56.5617
R432 commonsourceibias.n207 commonsourceibias.n206 56.5617
R433 commonsourceibias.n193 commonsourceibias.n192 56.5617
R434 commonsourceibias.n687 commonsourceibias.n685 56.5617
R435 commonsourceibias.n702 commonsourceibias.n700 56.5617
R436 commonsourceibias.n457 commonsourceibias.n455 56.5617
R437 commonsourceibias.n472 commonsourceibias.n470 56.5617
R438 commonsourceibias.n572 commonsourceibias.n570 56.5617
R439 commonsourceibias.n294 commonsourceibias.n293 56.5617
R440 commonsourceibias.n308 commonsourceibias.n307 56.5617
R441 commonsourceibias.n350 commonsourceibias.n349 56.5617
R442 commonsourceibias.n113 commonsourceibias.n112 56.5617
R443 commonsourceibias.n99 commonsourceibias.n98 56.5617
R444 commonsourceibias.n57 commonsourceibias.n56 56.5617
R445 commonsourceibias.n235 commonsourceibias.n234 56.5617
R446 commonsourceibias.n221 commonsourceibias.n220 56.5617
R447 commonsourceibias.n179 commonsourceibias.n178 56.5617
R448 commonsourceibias.n657 commonsourceibias.n655 56.5617
R449 commonsourceibias.n672 commonsourceibias.n670 56.5617
R450 commonsourceibias.n717 commonsourceibias.n715 56.5617
R451 commonsourceibias.n427 commonsourceibias.n425 56.5617
R452 commonsourceibias.n442 commonsourceibias.n440 56.5617
R453 commonsourceibias.n487 commonsourceibias.n485 56.5617
R454 commonsourceibias.n602 commonsourceibias.n600 56.5617
R455 commonsourceibias.n587 commonsourceibias.n585 56.5617
R456 commonsourceibias.n543 commonsourceibias.n541 56.5617
R457 commonsourceibias.n557 commonsourceibias.n556 56.5617
R458 commonsourceibias.n285 commonsourceibias.n284 51.2335
R459 commonsourceibias.n357 commonsourceibias.n252 51.2335
R460 commonsourceibias.n120 commonsourceibias.n15 51.2335
R461 commonsourceibias.n48 commonsourceibias.n47 51.2335
R462 commonsourceibias.n242 commonsourceibias.n1 51.2335
R463 commonsourceibias.n170 commonsourceibias.n169 51.2335
R464 commonsourceibias.n647 commonsourceibias.n646 51.2335
R465 commonsourceibias.n724 commonsourceibias.n619 51.2335
R466 commonsourceibias.n417 commonsourceibias.n416 51.2335
R467 commonsourceibias.n494 commonsourceibias.n389 51.2335
R468 commonsourceibias.n609 commonsourceibias.n368 51.2335
R469 commonsourceibias.n533 commonsourceibias.n532 51.2335
R470 commonsourceibias.n364 commonsourceibias.n363 50.9056
R471 commonsourceibias.n127 commonsourceibias.n126 50.9056
R472 commonsourceibias.n249 commonsourceibias.n248 50.9056
R473 commonsourceibias.n731 commonsourceibias.n730 50.9056
R474 commonsourceibias.n501 commonsourceibias.n500 50.9056
R475 commonsourceibias.n616 commonsourceibias.n615 50.9056
R476 commonsourceibias.n299 commonsourceibias.n298 50.2647
R477 commonsourceibias.n343 commonsourceibias.n257 50.2647
R478 commonsourceibias.n106 commonsourceibias.n20 50.2647
R479 commonsourceibias.n62 commonsourceibias.n61 50.2647
R480 commonsourceibias.n228 commonsourceibias.n6 50.2647
R481 commonsourceibias.n184 commonsourceibias.n183 50.2647
R482 commonsourceibias.n662 commonsourceibias.n661 50.2647
R483 commonsourceibias.n709 commonsourceibias.n623 50.2647
R484 commonsourceibias.n432 commonsourceibias.n431 50.2647
R485 commonsourceibias.n479 commonsourceibias.n393 50.2647
R486 commonsourceibias.n594 commonsourceibias.n372 50.2647
R487 commonsourceibias.n548 commonsourceibias.n547 50.2647
R488 commonsourceibias.n281 commonsourceibias.n280 49.9027
R489 commonsourceibias.n44 commonsourceibias.n43 49.9027
R490 commonsourceibias.n166 commonsourceibias.n165 49.9027
R491 commonsourceibias.n643 commonsourceibias.n642 49.9027
R492 commonsourceibias.n413 commonsourceibias.n412 49.9027
R493 commonsourceibias.n529 commonsourceibias.n528 49.9027
R494 commonsourceibias.n313 commonsourceibias.n312 49.296
R495 commonsourceibias.n329 commonsourceibias.n262 49.296
R496 commonsourceibias.n92 commonsourceibias.n25 49.296
R497 commonsourceibias.n76 commonsourceibias.n75 49.296
R498 commonsourceibias.n214 commonsourceibias.n11 49.296
R499 commonsourceibias.n198 commonsourceibias.n197 49.296
R500 commonsourceibias.n677 commonsourceibias.n676 49.296
R501 commonsourceibias.n694 commonsourceibias.n627 49.296
R502 commonsourceibias.n447 commonsourceibias.n446 49.296
R503 commonsourceibias.n464 commonsourceibias.n397 49.296
R504 commonsourceibias.n579 commonsourceibias.n376 49.296
R505 commonsourceibias.n562 commonsourceibias.n561 49.296
R506 commonsourceibias.n315 commonsourceibias.n267 48.3272
R507 commonsourceibias.n327 commonsourceibias.n326 48.3272
R508 commonsourceibias.n90 commonsourceibias.n89 48.3272
R509 commonsourceibias.n78 commonsourceibias.n30 48.3272
R510 commonsourceibias.n212 commonsourceibias.n211 48.3272
R511 commonsourceibias.n202 commonsourceibias.n201 48.3272
R512 commonsourceibias.n679 commonsourceibias.n631 48.3272
R513 commonsourceibias.n692 commonsourceibias.n691 48.3272
R514 commonsourceibias.n449 commonsourceibias.n401 48.3272
R515 commonsourceibias.n462 commonsourceibias.n461 48.3272
R516 commonsourceibias.n577 commonsourceibias.n576 48.3272
R517 commonsourceibias.n566 commonsourceibias.n565 48.3272
R518 commonsourceibias.n301 commonsourceibias.n272 47.3584
R519 commonsourceibias.n341 commonsourceibias.n340 47.3584
R520 commonsourceibias.n104 commonsourceibias.n103 47.3584
R521 commonsourceibias.n64 commonsourceibias.n35 47.3584
R522 commonsourceibias.n226 commonsourceibias.n225 47.3584
R523 commonsourceibias.n186 commonsourceibias.n157 47.3584
R524 commonsourceibias.n664 commonsourceibias.n635 47.3584
R525 commonsourceibias.n707 commonsourceibias.n706 47.3584
R526 commonsourceibias.n434 commonsourceibias.n405 47.3584
R527 commonsourceibias.n477 commonsourceibias.n476 47.3584
R528 commonsourceibias.n592 commonsourceibias.n591 47.3584
R529 commonsourceibias.n550 commonsourceibias.n521 47.3584
R530 commonsourceibias.n287 commonsourceibias.n277 46.3896
R531 commonsourceibias.n355 commonsourceibias.n354 46.3896
R532 commonsourceibias.n118 commonsourceibias.n117 46.3896
R533 commonsourceibias.n50 commonsourceibias.n40 46.3896
R534 commonsourceibias.n240 commonsourceibias.n239 46.3896
R535 commonsourceibias.n172 commonsourceibias.n162 46.3896
R536 commonsourceibias.n649 commonsourceibias.n639 46.3896
R537 commonsourceibias.n722 commonsourceibias.n721 46.3896
R538 commonsourceibias.n419 commonsourceibias.n409 46.3896
R539 commonsourceibias.n492 commonsourceibias.n491 46.3896
R540 commonsourceibias.n607 commonsourceibias.n606 46.3896
R541 commonsourceibias.n535 commonsourceibias.n525 46.3896
R542 commonsourceibias.n282 commonsourceibias.n281 44.7059
R543 commonsourceibias.n644 commonsourceibias.n643 44.7059
R544 commonsourceibias.n414 commonsourceibias.n413 44.7059
R545 commonsourceibias.n530 commonsourceibias.n529 44.7059
R546 commonsourceibias.n45 commonsourceibias.n44 44.7059
R547 commonsourceibias.n167 commonsourceibias.n166 44.7059
R548 commonsourceibias.n291 commonsourceibias.n277 34.7644
R549 commonsourceibias.n354 commonsourceibias.n254 34.7644
R550 commonsourceibias.n117 commonsourceibias.n17 34.7644
R551 commonsourceibias.n54 commonsourceibias.n40 34.7644
R552 commonsourceibias.n239 commonsourceibias.n3 34.7644
R553 commonsourceibias.n176 commonsourceibias.n162 34.7644
R554 commonsourceibias.n653 commonsourceibias.n639 34.7644
R555 commonsourceibias.n721 commonsourceibias.n621 34.7644
R556 commonsourceibias.n423 commonsourceibias.n409 34.7644
R557 commonsourceibias.n491 commonsourceibias.n391 34.7644
R558 commonsourceibias.n606 commonsourceibias.n370 34.7644
R559 commonsourceibias.n539 commonsourceibias.n525 34.7644
R560 commonsourceibias.n305 commonsourceibias.n272 33.7956
R561 commonsourceibias.n340 commonsourceibias.n259 33.7956
R562 commonsourceibias.n103 commonsourceibias.n22 33.7956
R563 commonsourceibias.n68 commonsourceibias.n35 33.7956
R564 commonsourceibias.n225 commonsourceibias.n8 33.7956
R565 commonsourceibias.n190 commonsourceibias.n157 33.7956
R566 commonsourceibias.n668 commonsourceibias.n635 33.7956
R567 commonsourceibias.n706 commonsourceibias.n625 33.7956
R568 commonsourceibias.n438 commonsourceibias.n405 33.7956
R569 commonsourceibias.n476 commonsourceibias.n395 33.7956
R570 commonsourceibias.n591 commonsourceibias.n374 33.7956
R571 commonsourceibias.n554 commonsourceibias.n521 33.7956
R572 commonsourceibias.n319 commonsourceibias.n267 32.8269
R573 commonsourceibias.n326 commonsourceibias.n264 32.8269
R574 commonsourceibias.n89 commonsourceibias.n27 32.8269
R575 commonsourceibias.n82 commonsourceibias.n30 32.8269
R576 commonsourceibias.n211 commonsourceibias.n13 32.8269
R577 commonsourceibias.n203 commonsourceibias.n202 32.8269
R578 commonsourceibias.n683 commonsourceibias.n631 32.8269
R579 commonsourceibias.n691 commonsourceibias.n629 32.8269
R580 commonsourceibias.n453 commonsourceibias.n401 32.8269
R581 commonsourceibias.n461 commonsourceibias.n399 32.8269
R582 commonsourceibias.n576 commonsourceibias.n378 32.8269
R583 commonsourceibias.n567 commonsourceibias.n566 32.8269
R584 commonsourceibias.n312 commonsourceibias.n269 31.8581
R585 commonsourceibias.n333 commonsourceibias.n262 31.8581
R586 commonsourceibias.n96 commonsourceibias.n25 31.8581
R587 commonsourceibias.n75 commonsourceibias.n32 31.8581
R588 commonsourceibias.n218 commonsourceibias.n11 31.8581
R589 commonsourceibias.n197 commonsourceibias.n196 31.8581
R590 commonsourceibias.n676 commonsourceibias.n633 31.8581
R591 commonsourceibias.n698 commonsourceibias.n627 31.8581
R592 commonsourceibias.n446 commonsourceibias.n403 31.8581
R593 commonsourceibias.n468 commonsourceibias.n397 31.8581
R594 commonsourceibias.n583 commonsourceibias.n376 31.8581
R595 commonsourceibias.n561 commonsourceibias.n560 31.8581
R596 commonsourceibias.n298 commonsourceibias.n274 30.8893
R597 commonsourceibias.n347 commonsourceibias.n257 30.8893
R598 commonsourceibias.n110 commonsourceibias.n20 30.8893
R599 commonsourceibias.n61 commonsourceibias.n37 30.8893
R600 commonsourceibias.n232 commonsourceibias.n6 30.8893
R601 commonsourceibias.n183 commonsourceibias.n159 30.8893
R602 commonsourceibias.n661 commonsourceibias.n637 30.8893
R603 commonsourceibias.n713 commonsourceibias.n623 30.8893
R604 commonsourceibias.n431 commonsourceibias.n407 30.8893
R605 commonsourceibias.n483 commonsourceibias.n393 30.8893
R606 commonsourceibias.n598 commonsourceibias.n372 30.8893
R607 commonsourceibias.n547 commonsourceibias.n523 30.8893
R608 commonsourceibias.n284 commonsourceibias.n279 29.9206
R609 commonsourceibias.n361 commonsourceibias.n252 29.9206
R610 commonsourceibias.n124 commonsourceibias.n15 29.9206
R611 commonsourceibias.n47 commonsourceibias.n42 29.9206
R612 commonsourceibias.n246 commonsourceibias.n1 29.9206
R613 commonsourceibias.n169 commonsourceibias.n164 29.9206
R614 commonsourceibias.n646 commonsourceibias.n641 29.9206
R615 commonsourceibias.n728 commonsourceibias.n619 29.9206
R616 commonsourceibias.n416 commonsourceibias.n411 29.9206
R617 commonsourceibias.n498 commonsourceibias.n389 29.9206
R618 commonsourceibias.n613 commonsourceibias.n368 29.9206
R619 commonsourceibias.n532 commonsourceibias.n527 29.9206
R620 commonsourceibias.n363 commonsourceibias.n362 21.8872
R621 commonsourceibias.n126 commonsourceibias.n125 21.8872
R622 commonsourceibias.n248 commonsourceibias.n247 21.8872
R623 commonsourceibias.n730 commonsourceibias.n729 21.8872
R624 commonsourceibias.n500 commonsourceibias.n499 21.8872
R625 commonsourceibias.n615 commonsourceibias.n614 21.8872
R626 commonsourceibias.n294 commonsourceibias.n276 21.3954
R627 commonsourceibias.n349 commonsourceibias.n348 21.3954
R628 commonsourceibias.n112 commonsourceibias.n111 21.3954
R629 commonsourceibias.n57 commonsourceibias.n39 21.3954
R630 commonsourceibias.n234 commonsourceibias.n233 21.3954
R631 commonsourceibias.n179 commonsourceibias.n161 21.3954
R632 commonsourceibias.n657 commonsourceibias.n656 21.3954
R633 commonsourceibias.n715 commonsourceibias.n714 21.3954
R634 commonsourceibias.n427 commonsourceibias.n426 21.3954
R635 commonsourceibias.n485 commonsourceibias.n484 21.3954
R636 commonsourceibias.n600 commonsourceibias.n599 21.3954
R637 commonsourceibias.n543 commonsourceibias.n542 21.3954
R638 commonsourceibias.n308 commonsourceibias.n271 20.9036
R639 commonsourceibias.n335 commonsourceibias.n334 20.9036
R640 commonsourceibias.n98 commonsourceibias.n97 20.9036
R641 commonsourceibias.n71 commonsourceibias.n34 20.9036
R642 commonsourceibias.n220 commonsourceibias.n219 20.9036
R643 commonsourceibias.n193 commonsourceibias.n155 20.9036
R644 commonsourceibias.n672 commonsourceibias.n671 20.9036
R645 commonsourceibias.n700 commonsourceibias.n699 20.9036
R646 commonsourceibias.n442 commonsourceibias.n441 20.9036
R647 commonsourceibias.n470 commonsourceibias.n469 20.9036
R648 commonsourceibias.n585 commonsourceibias.n584 20.9036
R649 commonsourceibias.n557 commonsourceibias.n519 20.9036
R650 commonsourceibias.n321 commonsourceibias.n320 20.4117
R651 commonsourceibias.n322 commonsourceibias.n266 20.4117
R652 commonsourceibias.n85 commonsourceibias.n29 20.4117
R653 commonsourceibias.n84 commonsourceibias.n83 20.4117
R654 commonsourceibias.n207 commonsourceibias.n150 20.4117
R655 commonsourceibias.n206 commonsourceibias.n151 20.4117
R656 commonsourceibias.n685 commonsourceibias.n684 20.4117
R657 commonsourceibias.n687 commonsourceibias.n686 20.4117
R658 commonsourceibias.n455 commonsourceibias.n454 20.4117
R659 commonsourceibias.n457 commonsourceibias.n456 20.4117
R660 commonsourceibias.n572 commonsourceibias.n571 20.4117
R661 commonsourceibias.n570 commonsourceibias.n515 20.4117
R662 commonsourceibias.n307 commonsourceibias.n306 19.9199
R663 commonsourceibias.n336 commonsourceibias.n261 19.9199
R664 commonsourceibias.n99 commonsourceibias.n24 19.9199
R665 commonsourceibias.n70 commonsourceibias.n69 19.9199
R666 commonsourceibias.n221 commonsourceibias.n10 19.9199
R667 commonsourceibias.n192 commonsourceibias.n191 19.9199
R668 commonsourceibias.n670 commonsourceibias.n669 19.9199
R669 commonsourceibias.n702 commonsourceibias.n701 19.9199
R670 commonsourceibias.n440 commonsourceibias.n439 19.9199
R671 commonsourceibias.n472 commonsourceibias.n471 19.9199
R672 commonsourceibias.n587 commonsourceibias.n586 19.9199
R673 commonsourceibias.n556 commonsourceibias.n555 19.9199
R674 commonsourceibias.n293 commonsourceibias.n292 19.4281
R675 commonsourceibias.n350 commonsourceibias.n256 19.4281
R676 commonsourceibias.n113 commonsourceibias.n19 19.4281
R677 commonsourceibias.n56 commonsourceibias.n55 19.4281
R678 commonsourceibias.n235 commonsourceibias.n5 19.4281
R679 commonsourceibias.n178 commonsourceibias.n177 19.4281
R680 commonsourceibias.n655 commonsourceibias.n654 19.4281
R681 commonsourceibias.n717 commonsourceibias.n716 19.4281
R682 commonsourceibias.n425 commonsourceibias.n424 19.4281
R683 commonsourceibias.n487 commonsourceibias.n486 19.4281
R684 commonsourceibias.n602 commonsourceibias.n601 19.4281
R685 commonsourceibias.n541 commonsourceibias.n540 19.4281
R686 commonsourceibias.n286 commonsourceibias.n285 13.526
R687 commonsourceibias.n357 commonsourceibias.n356 13.526
R688 commonsourceibias.n120 commonsourceibias.n119 13.526
R689 commonsourceibias.n49 commonsourceibias.n48 13.526
R690 commonsourceibias.n242 commonsourceibias.n241 13.526
R691 commonsourceibias.n171 commonsourceibias.n170 13.526
R692 commonsourceibias.n648 commonsourceibias.n647 13.526
R693 commonsourceibias.n724 commonsourceibias.n723 13.526
R694 commonsourceibias.n418 commonsourceibias.n417 13.526
R695 commonsourceibias.n494 commonsourceibias.n493 13.526
R696 commonsourceibias.n609 commonsourceibias.n608 13.526
R697 commonsourceibias.n534 commonsourceibias.n533 13.526
R698 commonsourceibias.n130 commonsourceibias.n128 13.2322
R699 commonsourceibias.n504 commonsourceibias.n502 13.2322
R700 commonsourceibias.n300 commonsourceibias.n299 13.0342
R701 commonsourceibias.n343 commonsourceibias.n342 13.0342
R702 commonsourceibias.n106 commonsourceibias.n105 13.0342
R703 commonsourceibias.n63 commonsourceibias.n62 13.0342
R704 commonsourceibias.n228 commonsourceibias.n227 13.0342
R705 commonsourceibias.n185 commonsourceibias.n184 13.0342
R706 commonsourceibias.n663 commonsourceibias.n662 13.0342
R707 commonsourceibias.n709 commonsourceibias.n708 13.0342
R708 commonsourceibias.n433 commonsourceibias.n432 13.0342
R709 commonsourceibias.n479 commonsourceibias.n478 13.0342
R710 commonsourceibias.n594 commonsourceibias.n593 13.0342
R711 commonsourceibias.n549 commonsourceibias.n548 13.0342
R712 commonsourceibias.n314 commonsourceibias.n313 12.5423
R713 commonsourceibias.n329 commonsourceibias.n328 12.5423
R714 commonsourceibias.n92 commonsourceibias.n91 12.5423
R715 commonsourceibias.n77 commonsourceibias.n76 12.5423
R716 commonsourceibias.n214 commonsourceibias.n213 12.5423
R717 commonsourceibias.n198 commonsourceibias.n153 12.5423
R718 commonsourceibias.n678 commonsourceibias.n677 12.5423
R719 commonsourceibias.n694 commonsourceibias.n693 12.5423
R720 commonsourceibias.n448 commonsourceibias.n447 12.5423
R721 commonsourceibias.n464 commonsourceibias.n463 12.5423
R722 commonsourceibias.n579 commonsourceibias.n578 12.5423
R723 commonsourceibias.n562 commonsourceibias.n517 12.5423
R724 commonsourceibias.n315 commonsourceibias.n314 12.0505
R725 commonsourceibias.n328 commonsourceibias.n327 12.0505
R726 commonsourceibias.n91 commonsourceibias.n90 12.0505
R727 commonsourceibias.n78 commonsourceibias.n77 12.0505
R728 commonsourceibias.n213 commonsourceibias.n212 12.0505
R729 commonsourceibias.n201 commonsourceibias.n153 12.0505
R730 commonsourceibias.n679 commonsourceibias.n678 12.0505
R731 commonsourceibias.n693 commonsourceibias.n692 12.0505
R732 commonsourceibias.n449 commonsourceibias.n448 12.0505
R733 commonsourceibias.n463 commonsourceibias.n462 12.0505
R734 commonsourceibias.n578 commonsourceibias.n577 12.0505
R735 commonsourceibias.n565 commonsourceibias.n517 12.0505
R736 commonsourceibias.n734 commonsourceibias.n366 11.9876
R737 commonsourceibias.n301 commonsourceibias.n300 11.5587
R738 commonsourceibias.n342 commonsourceibias.n341 11.5587
R739 commonsourceibias.n105 commonsourceibias.n104 11.5587
R740 commonsourceibias.n64 commonsourceibias.n63 11.5587
R741 commonsourceibias.n227 commonsourceibias.n226 11.5587
R742 commonsourceibias.n186 commonsourceibias.n185 11.5587
R743 commonsourceibias.n664 commonsourceibias.n663 11.5587
R744 commonsourceibias.n708 commonsourceibias.n707 11.5587
R745 commonsourceibias.n434 commonsourceibias.n433 11.5587
R746 commonsourceibias.n478 commonsourceibias.n477 11.5587
R747 commonsourceibias.n593 commonsourceibias.n592 11.5587
R748 commonsourceibias.n550 commonsourceibias.n549 11.5587
R749 commonsourceibias.n287 commonsourceibias.n286 11.0668
R750 commonsourceibias.n356 commonsourceibias.n355 11.0668
R751 commonsourceibias.n119 commonsourceibias.n118 11.0668
R752 commonsourceibias.n50 commonsourceibias.n49 11.0668
R753 commonsourceibias.n241 commonsourceibias.n240 11.0668
R754 commonsourceibias.n172 commonsourceibias.n171 11.0668
R755 commonsourceibias.n649 commonsourceibias.n648 11.0668
R756 commonsourceibias.n723 commonsourceibias.n722 11.0668
R757 commonsourceibias.n419 commonsourceibias.n418 11.0668
R758 commonsourceibias.n493 commonsourceibias.n492 11.0668
R759 commonsourceibias.n608 commonsourceibias.n607 11.0668
R760 commonsourceibias.n535 commonsourceibias.n534 11.0668
R761 commonsourceibias.n734 commonsourceibias.n733 10.3347
R762 commonsourceibias.n149 commonsourceibias.n148 9.50363
R763 commonsourceibias.n514 commonsourceibias.n513 9.50363
R764 commonsourceibias.n366 commonsourceibias.n250 8.75852
R765 commonsourceibias.n733 commonsourceibias.n617 8.75852
R766 commonsourceibias.n292 commonsourceibias.n291 5.16479
R767 commonsourceibias.n256 commonsourceibias.n254 5.16479
R768 commonsourceibias.n19 commonsourceibias.n17 5.16479
R769 commonsourceibias.n55 commonsourceibias.n54 5.16479
R770 commonsourceibias.n5 commonsourceibias.n3 5.16479
R771 commonsourceibias.n177 commonsourceibias.n176 5.16479
R772 commonsourceibias.n654 commonsourceibias.n653 5.16479
R773 commonsourceibias.n716 commonsourceibias.n621 5.16479
R774 commonsourceibias.n424 commonsourceibias.n423 5.16479
R775 commonsourceibias.n486 commonsourceibias.n391 5.16479
R776 commonsourceibias.n601 commonsourceibias.n370 5.16479
R777 commonsourceibias.n540 commonsourceibias.n539 5.16479
R778 commonsourceibias.n366 commonsourceibias.n365 5.03125
R779 commonsourceibias.n733 commonsourceibias.n732 5.03125
R780 commonsourceibias.n306 commonsourceibias.n305 4.67295
R781 commonsourceibias.n261 commonsourceibias.n259 4.67295
R782 commonsourceibias.n24 commonsourceibias.n22 4.67295
R783 commonsourceibias.n69 commonsourceibias.n68 4.67295
R784 commonsourceibias.n10 commonsourceibias.n8 4.67295
R785 commonsourceibias.n191 commonsourceibias.n190 4.67295
R786 commonsourceibias.n669 commonsourceibias.n668 4.67295
R787 commonsourceibias.n701 commonsourceibias.n625 4.67295
R788 commonsourceibias.n439 commonsourceibias.n438 4.67295
R789 commonsourceibias.n471 commonsourceibias.n395 4.67295
R790 commonsourceibias.n586 commonsourceibias.n374 4.67295
R791 commonsourceibias.n555 commonsourceibias.n554 4.67295
R792 commonsourceibias commonsourceibias.n734 4.20978
R793 commonsourceibias.n320 commonsourceibias.n319 4.18111
R794 commonsourceibias.n266 commonsourceibias.n264 4.18111
R795 commonsourceibias.n29 commonsourceibias.n27 4.18111
R796 commonsourceibias.n83 commonsourceibias.n82 4.18111
R797 commonsourceibias.n150 commonsourceibias.n13 4.18111
R798 commonsourceibias.n203 commonsourceibias.n151 4.18111
R799 commonsourceibias.n684 commonsourceibias.n683 4.18111
R800 commonsourceibias.n686 commonsourceibias.n629 4.18111
R801 commonsourceibias.n454 commonsourceibias.n453 4.18111
R802 commonsourceibias.n456 commonsourceibias.n399 4.18111
R803 commonsourceibias.n571 commonsourceibias.n378 4.18111
R804 commonsourceibias.n567 commonsourceibias.n515 4.18111
R805 commonsourceibias.n271 commonsourceibias.n269 3.68928
R806 commonsourceibias.n334 commonsourceibias.n333 3.68928
R807 commonsourceibias.n97 commonsourceibias.n96 3.68928
R808 commonsourceibias.n34 commonsourceibias.n32 3.68928
R809 commonsourceibias.n219 commonsourceibias.n218 3.68928
R810 commonsourceibias.n196 commonsourceibias.n155 3.68928
R811 commonsourceibias.n671 commonsourceibias.n633 3.68928
R812 commonsourceibias.n699 commonsourceibias.n698 3.68928
R813 commonsourceibias.n441 commonsourceibias.n403 3.68928
R814 commonsourceibias.n469 commonsourceibias.n468 3.68928
R815 commonsourceibias.n584 commonsourceibias.n583 3.68928
R816 commonsourceibias.n560 commonsourceibias.n519 3.68928
R817 commonsourceibias.n276 commonsourceibias.n274 3.19744
R818 commonsourceibias.n348 commonsourceibias.n347 3.19744
R819 commonsourceibias.n111 commonsourceibias.n110 3.19744
R820 commonsourceibias.n39 commonsourceibias.n37 3.19744
R821 commonsourceibias.n233 commonsourceibias.n232 3.19744
R822 commonsourceibias.n161 commonsourceibias.n159 3.19744
R823 commonsourceibias.n656 commonsourceibias.n637 3.19744
R824 commonsourceibias.n714 commonsourceibias.n713 3.19744
R825 commonsourceibias.n426 commonsourceibias.n407 3.19744
R826 commonsourceibias.n484 commonsourceibias.n483 3.19744
R827 commonsourceibias.n599 commonsourceibias.n598 3.19744
R828 commonsourceibias.n542 commonsourceibias.n523 3.19744
R829 commonsourceibias.n139 commonsourceibias.t13 2.82907
R830 commonsourceibias.n139 commonsourceibias.t55 2.82907
R831 commonsourceibias.n140 commonsourceibias.t35 2.82907
R832 commonsourceibias.n140 commonsourceibias.t23 2.82907
R833 commonsourceibias.n142 commonsourceibias.t27 2.82907
R834 commonsourceibias.n142 commonsourceibias.t61 2.82907
R835 commonsourceibias.n144 commonsourceibias.t1 2.82907
R836 commonsourceibias.n144 commonsourceibias.t51 2.82907
R837 commonsourceibias.n146 commonsourceibias.t41 2.82907
R838 commonsourceibias.n146 commonsourceibias.t47 2.82907
R839 commonsourceibias.n137 commonsourceibias.t79 2.82907
R840 commonsourceibias.n137 commonsourceibias.t9 2.82907
R841 commonsourceibias.n135 commonsourceibias.t45 2.82907
R842 commonsourceibias.n135 commonsourceibias.t71 2.82907
R843 commonsourceibias.n133 commonsourceibias.t5 2.82907
R844 commonsourceibias.n133 commonsourceibias.t49 2.82907
R845 commonsourceibias.n131 commonsourceibias.t65 2.82907
R846 commonsourceibias.n131 commonsourceibias.t75 2.82907
R847 commonsourceibias.n129 commonsourceibias.t77 2.82907
R848 commonsourceibias.n129 commonsourceibias.t25 2.82907
R849 commonsourceibias.n503 commonsourceibias.t7 2.82907
R850 commonsourceibias.n503 commonsourceibias.t33 2.82907
R851 commonsourceibias.n505 commonsourceibias.t31 2.82907
R852 commonsourceibias.n505 commonsourceibias.t53 2.82907
R853 commonsourceibias.n507 commonsourceibias.t39 2.82907
R854 commonsourceibias.n507 commonsourceibias.t73 2.82907
R855 commonsourceibias.n509 commonsourceibias.t43 2.82907
R856 commonsourceibias.n509 commonsourceibias.t11 2.82907
R857 commonsourceibias.n511 commonsourceibias.t3 2.82907
R858 commonsourceibias.n511 commonsourceibias.t37 2.82907
R859 commonsourceibias.n386 commonsourceibias.t29 2.82907
R860 commonsourceibias.n386 commonsourceibias.t21 2.82907
R861 commonsourceibias.n384 commonsourceibias.t19 2.82907
R862 commonsourceibias.n384 commonsourceibias.t63 2.82907
R863 commonsourceibias.n382 commonsourceibias.t57 2.82907
R864 commonsourceibias.n382 commonsourceibias.t59 2.82907
R865 commonsourceibias.n380 commonsourceibias.t67 2.82907
R866 commonsourceibias.n380 commonsourceibias.t15 2.82907
R867 commonsourceibias.n379 commonsourceibias.t17 2.82907
R868 commonsourceibias.n379 commonsourceibias.t69 2.82907
R869 commonsourceibias.n280 commonsourceibias.n279 2.7056
R870 commonsourceibias.n362 commonsourceibias.n361 2.7056
R871 commonsourceibias.n125 commonsourceibias.n124 2.7056
R872 commonsourceibias.n43 commonsourceibias.n42 2.7056
R873 commonsourceibias.n247 commonsourceibias.n246 2.7056
R874 commonsourceibias.n165 commonsourceibias.n164 2.7056
R875 commonsourceibias.n642 commonsourceibias.n641 2.7056
R876 commonsourceibias.n729 commonsourceibias.n728 2.7056
R877 commonsourceibias.n412 commonsourceibias.n411 2.7056
R878 commonsourceibias.n499 commonsourceibias.n498 2.7056
R879 commonsourceibias.n614 commonsourceibias.n613 2.7056
R880 commonsourceibias.n528 commonsourceibias.n527 2.7056
R881 commonsourceibias.n132 commonsourceibias.n130 0.573776
R882 commonsourceibias.n134 commonsourceibias.n132 0.573776
R883 commonsourceibias.n136 commonsourceibias.n134 0.573776
R884 commonsourceibias.n138 commonsourceibias.n136 0.573776
R885 commonsourceibias.n147 commonsourceibias.n145 0.573776
R886 commonsourceibias.n145 commonsourceibias.n143 0.573776
R887 commonsourceibias.n143 commonsourceibias.n141 0.573776
R888 commonsourceibias.n383 commonsourceibias.n381 0.573776
R889 commonsourceibias.n385 commonsourceibias.n383 0.573776
R890 commonsourceibias.n387 commonsourceibias.n385 0.573776
R891 commonsourceibias.n512 commonsourceibias.n510 0.573776
R892 commonsourceibias.n510 commonsourceibias.n508 0.573776
R893 commonsourceibias.n508 commonsourceibias.n506 0.573776
R894 commonsourceibias.n506 commonsourceibias.n504 0.573776
R895 commonsourceibias.n148 commonsourceibias.n138 0.287138
R896 commonsourceibias.n148 commonsourceibias.n147 0.287138
R897 commonsourceibias.n513 commonsourceibias.n387 0.287138
R898 commonsourceibias.n513 commonsourceibias.n512 0.287138
R899 commonsourceibias.n365 commonsourceibias.n251 0.285035
R900 commonsourceibias.n128 commonsourceibias.n14 0.285035
R901 commonsourceibias.n250 commonsourceibias.n0 0.285035
R902 commonsourceibias.n732 commonsourceibias.n618 0.285035
R903 commonsourceibias.n502 commonsourceibias.n388 0.285035
R904 commonsourceibias.n617 commonsourceibias.n367 0.285035
R905 commonsourceibias.n360 commonsourceibias.n251 0.189894
R906 commonsourceibias.n360 commonsourceibias.n359 0.189894
R907 commonsourceibias.n359 commonsourceibias.n358 0.189894
R908 commonsourceibias.n358 commonsourceibias.n253 0.189894
R909 commonsourceibias.n353 commonsourceibias.n253 0.189894
R910 commonsourceibias.n353 commonsourceibias.n352 0.189894
R911 commonsourceibias.n352 commonsourceibias.n351 0.189894
R912 commonsourceibias.n351 commonsourceibias.n255 0.189894
R913 commonsourceibias.n346 commonsourceibias.n255 0.189894
R914 commonsourceibias.n346 commonsourceibias.n345 0.189894
R915 commonsourceibias.n345 commonsourceibias.n344 0.189894
R916 commonsourceibias.n344 commonsourceibias.n258 0.189894
R917 commonsourceibias.n339 commonsourceibias.n258 0.189894
R918 commonsourceibias.n339 commonsourceibias.n338 0.189894
R919 commonsourceibias.n338 commonsourceibias.n337 0.189894
R920 commonsourceibias.n337 commonsourceibias.n260 0.189894
R921 commonsourceibias.n332 commonsourceibias.n260 0.189894
R922 commonsourceibias.n332 commonsourceibias.n331 0.189894
R923 commonsourceibias.n331 commonsourceibias.n330 0.189894
R924 commonsourceibias.n330 commonsourceibias.n263 0.189894
R925 commonsourceibias.n325 commonsourceibias.n263 0.189894
R926 commonsourceibias.n325 commonsourceibias.n324 0.189894
R927 commonsourceibias.n324 commonsourceibias.n323 0.189894
R928 commonsourceibias.n323 commonsourceibias.n265 0.189894
R929 commonsourceibias.n318 commonsourceibias.n265 0.189894
R930 commonsourceibias.n318 commonsourceibias.n317 0.189894
R931 commonsourceibias.n317 commonsourceibias.n316 0.189894
R932 commonsourceibias.n316 commonsourceibias.n268 0.189894
R933 commonsourceibias.n311 commonsourceibias.n268 0.189894
R934 commonsourceibias.n311 commonsourceibias.n310 0.189894
R935 commonsourceibias.n310 commonsourceibias.n309 0.189894
R936 commonsourceibias.n309 commonsourceibias.n270 0.189894
R937 commonsourceibias.n304 commonsourceibias.n270 0.189894
R938 commonsourceibias.n304 commonsourceibias.n303 0.189894
R939 commonsourceibias.n303 commonsourceibias.n302 0.189894
R940 commonsourceibias.n302 commonsourceibias.n273 0.189894
R941 commonsourceibias.n297 commonsourceibias.n273 0.189894
R942 commonsourceibias.n297 commonsourceibias.n296 0.189894
R943 commonsourceibias.n296 commonsourceibias.n295 0.189894
R944 commonsourceibias.n295 commonsourceibias.n275 0.189894
R945 commonsourceibias.n290 commonsourceibias.n275 0.189894
R946 commonsourceibias.n290 commonsourceibias.n289 0.189894
R947 commonsourceibias.n289 commonsourceibias.n288 0.189894
R948 commonsourceibias.n288 commonsourceibias.n278 0.189894
R949 commonsourceibias.n283 commonsourceibias.n278 0.189894
R950 commonsourceibias.n283 commonsourceibias.n282 0.189894
R951 commonsourceibias.n123 commonsourceibias.n14 0.189894
R952 commonsourceibias.n123 commonsourceibias.n122 0.189894
R953 commonsourceibias.n122 commonsourceibias.n121 0.189894
R954 commonsourceibias.n121 commonsourceibias.n16 0.189894
R955 commonsourceibias.n116 commonsourceibias.n16 0.189894
R956 commonsourceibias.n116 commonsourceibias.n115 0.189894
R957 commonsourceibias.n115 commonsourceibias.n114 0.189894
R958 commonsourceibias.n114 commonsourceibias.n18 0.189894
R959 commonsourceibias.n109 commonsourceibias.n18 0.189894
R960 commonsourceibias.n109 commonsourceibias.n108 0.189894
R961 commonsourceibias.n108 commonsourceibias.n107 0.189894
R962 commonsourceibias.n107 commonsourceibias.n21 0.189894
R963 commonsourceibias.n102 commonsourceibias.n21 0.189894
R964 commonsourceibias.n102 commonsourceibias.n101 0.189894
R965 commonsourceibias.n101 commonsourceibias.n100 0.189894
R966 commonsourceibias.n100 commonsourceibias.n23 0.189894
R967 commonsourceibias.n95 commonsourceibias.n23 0.189894
R968 commonsourceibias.n95 commonsourceibias.n94 0.189894
R969 commonsourceibias.n94 commonsourceibias.n93 0.189894
R970 commonsourceibias.n93 commonsourceibias.n26 0.189894
R971 commonsourceibias.n88 commonsourceibias.n26 0.189894
R972 commonsourceibias.n88 commonsourceibias.n87 0.189894
R973 commonsourceibias.n87 commonsourceibias.n86 0.189894
R974 commonsourceibias.n86 commonsourceibias.n28 0.189894
R975 commonsourceibias.n81 commonsourceibias.n28 0.189894
R976 commonsourceibias.n81 commonsourceibias.n80 0.189894
R977 commonsourceibias.n80 commonsourceibias.n79 0.189894
R978 commonsourceibias.n79 commonsourceibias.n31 0.189894
R979 commonsourceibias.n74 commonsourceibias.n31 0.189894
R980 commonsourceibias.n74 commonsourceibias.n73 0.189894
R981 commonsourceibias.n73 commonsourceibias.n72 0.189894
R982 commonsourceibias.n72 commonsourceibias.n33 0.189894
R983 commonsourceibias.n67 commonsourceibias.n33 0.189894
R984 commonsourceibias.n67 commonsourceibias.n66 0.189894
R985 commonsourceibias.n66 commonsourceibias.n65 0.189894
R986 commonsourceibias.n65 commonsourceibias.n36 0.189894
R987 commonsourceibias.n60 commonsourceibias.n36 0.189894
R988 commonsourceibias.n60 commonsourceibias.n59 0.189894
R989 commonsourceibias.n59 commonsourceibias.n58 0.189894
R990 commonsourceibias.n58 commonsourceibias.n38 0.189894
R991 commonsourceibias.n53 commonsourceibias.n38 0.189894
R992 commonsourceibias.n53 commonsourceibias.n52 0.189894
R993 commonsourceibias.n52 commonsourceibias.n51 0.189894
R994 commonsourceibias.n51 commonsourceibias.n41 0.189894
R995 commonsourceibias.n46 commonsourceibias.n41 0.189894
R996 commonsourceibias.n46 commonsourceibias.n45 0.189894
R997 commonsourceibias.n205 commonsourceibias.n204 0.189894
R998 commonsourceibias.n204 commonsourceibias.n152 0.189894
R999 commonsourceibias.n200 commonsourceibias.n152 0.189894
R1000 commonsourceibias.n200 commonsourceibias.n199 0.189894
R1001 commonsourceibias.n199 commonsourceibias.n154 0.189894
R1002 commonsourceibias.n195 commonsourceibias.n154 0.189894
R1003 commonsourceibias.n195 commonsourceibias.n194 0.189894
R1004 commonsourceibias.n194 commonsourceibias.n156 0.189894
R1005 commonsourceibias.n189 commonsourceibias.n156 0.189894
R1006 commonsourceibias.n189 commonsourceibias.n188 0.189894
R1007 commonsourceibias.n188 commonsourceibias.n187 0.189894
R1008 commonsourceibias.n187 commonsourceibias.n158 0.189894
R1009 commonsourceibias.n182 commonsourceibias.n158 0.189894
R1010 commonsourceibias.n182 commonsourceibias.n181 0.189894
R1011 commonsourceibias.n181 commonsourceibias.n180 0.189894
R1012 commonsourceibias.n180 commonsourceibias.n160 0.189894
R1013 commonsourceibias.n175 commonsourceibias.n160 0.189894
R1014 commonsourceibias.n175 commonsourceibias.n174 0.189894
R1015 commonsourceibias.n174 commonsourceibias.n173 0.189894
R1016 commonsourceibias.n173 commonsourceibias.n163 0.189894
R1017 commonsourceibias.n168 commonsourceibias.n163 0.189894
R1018 commonsourceibias.n168 commonsourceibias.n167 0.189894
R1019 commonsourceibias.n245 commonsourceibias.n0 0.189894
R1020 commonsourceibias.n245 commonsourceibias.n244 0.189894
R1021 commonsourceibias.n244 commonsourceibias.n243 0.189894
R1022 commonsourceibias.n243 commonsourceibias.n2 0.189894
R1023 commonsourceibias.n238 commonsourceibias.n2 0.189894
R1024 commonsourceibias.n238 commonsourceibias.n237 0.189894
R1025 commonsourceibias.n237 commonsourceibias.n236 0.189894
R1026 commonsourceibias.n236 commonsourceibias.n4 0.189894
R1027 commonsourceibias.n231 commonsourceibias.n4 0.189894
R1028 commonsourceibias.n231 commonsourceibias.n230 0.189894
R1029 commonsourceibias.n230 commonsourceibias.n229 0.189894
R1030 commonsourceibias.n229 commonsourceibias.n7 0.189894
R1031 commonsourceibias.n224 commonsourceibias.n7 0.189894
R1032 commonsourceibias.n224 commonsourceibias.n223 0.189894
R1033 commonsourceibias.n223 commonsourceibias.n222 0.189894
R1034 commonsourceibias.n222 commonsourceibias.n9 0.189894
R1035 commonsourceibias.n217 commonsourceibias.n9 0.189894
R1036 commonsourceibias.n217 commonsourceibias.n216 0.189894
R1037 commonsourceibias.n216 commonsourceibias.n215 0.189894
R1038 commonsourceibias.n215 commonsourceibias.n12 0.189894
R1039 commonsourceibias.n210 commonsourceibias.n12 0.189894
R1040 commonsourceibias.n210 commonsourceibias.n209 0.189894
R1041 commonsourceibias.n209 commonsourceibias.n208 0.189894
R1042 commonsourceibias.n645 commonsourceibias.n644 0.189894
R1043 commonsourceibias.n645 commonsourceibias.n640 0.189894
R1044 commonsourceibias.n650 commonsourceibias.n640 0.189894
R1045 commonsourceibias.n651 commonsourceibias.n650 0.189894
R1046 commonsourceibias.n652 commonsourceibias.n651 0.189894
R1047 commonsourceibias.n652 commonsourceibias.n638 0.189894
R1048 commonsourceibias.n658 commonsourceibias.n638 0.189894
R1049 commonsourceibias.n659 commonsourceibias.n658 0.189894
R1050 commonsourceibias.n660 commonsourceibias.n659 0.189894
R1051 commonsourceibias.n660 commonsourceibias.n636 0.189894
R1052 commonsourceibias.n665 commonsourceibias.n636 0.189894
R1053 commonsourceibias.n666 commonsourceibias.n665 0.189894
R1054 commonsourceibias.n667 commonsourceibias.n666 0.189894
R1055 commonsourceibias.n667 commonsourceibias.n634 0.189894
R1056 commonsourceibias.n673 commonsourceibias.n634 0.189894
R1057 commonsourceibias.n674 commonsourceibias.n673 0.189894
R1058 commonsourceibias.n675 commonsourceibias.n674 0.189894
R1059 commonsourceibias.n675 commonsourceibias.n632 0.189894
R1060 commonsourceibias.n680 commonsourceibias.n632 0.189894
R1061 commonsourceibias.n681 commonsourceibias.n680 0.189894
R1062 commonsourceibias.n682 commonsourceibias.n681 0.189894
R1063 commonsourceibias.n682 commonsourceibias.n630 0.189894
R1064 commonsourceibias.n688 commonsourceibias.n630 0.189894
R1065 commonsourceibias.n689 commonsourceibias.n688 0.189894
R1066 commonsourceibias.n690 commonsourceibias.n689 0.189894
R1067 commonsourceibias.n690 commonsourceibias.n628 0.189894
R1068 commonsourceibias.n695 commonsourceibias.n628 0.189894
R1069 commonsourceibias.n696 commonsourceibias.n695 0.189894
R1070 commonsourceibias.n697 commonsourceibias.n696 0.189894
R1071 commonsourceibias.n697 commonsourceibias.n626 0.189894
R1072 commonsourceibias.n703 commonsourceibias.n626 0.189894
R1073 commonsourceibias.n704 commonsourceibias.n703 0.189894
R1074 commonsourceibias.n705 commonsourceibias.n704 0.189894
R1075 commonsourceibias.n705 commonsourceibias.n624 0.189894
R1076 commonsourceibias.n710 commonsourceibias.n624 0.189894
R1077 commonsourceibias.n711 commonsourceibias.n710 0.189894
R1078 commonsourceibias.n712 commonsourceibias.n711 0.189894
R1079 commonsourceibias.n712 commonsourceibias.n622 0.189894
R1080 commonsourceibias.n718 commonsourceibias.n622 0.189894
R1081 commonsourceibias.n719 commonsourceibias.n718 0.189894
R1082 commonsourceibias.n720 commonsourceibias.n719 0.189894
R1083 commonsourceibias.n720 commonsourceibias.n620 0.189894
R1084 commonsourceibias.n725 commonsourceibias.n620 0.189894
R1085 commonsourceibias.n726 commonsourceibias.n725 0.189894
R1086 commonsourceibias.n727 commonsourceibias.n726 0.189894
R1087 commonsourceibias.n727 commonsourceibias.n618 0.189894
R1088 commonsourceibias.n415 commonsourceibias.n414 0.189894
R1089 commonsourceibias.n415 commonsourceibias.n410 0.189894
R1090 commonsourceibias.n420 commonsourceibias.n410 0.189894
R1091 commonsourceibias.n421 commonsourceibias.n420 0.189894
R1092 commonsourceibias.n422 commonsourceibias.n421 0.189894
R1093 commonsourceibias.n422 commonsourceibias.n408 0.189894
R1094 commonsourceibias.n428 commonsourceibias.n408 0.189894
R1095 commonsourceibias.n429 commonsourceibias.n428 0.189894
R1096 commonsourceibias.n430 commonsourceibias.n429 0.189894
R1097 commonsourceibias.n430 commonsourceibias.n406 0.189894
R1098 commonsourceibias.n435 commonsourceibias.n406 0.189894
R1099 commonsourceibias.n436 commonsourceibias.n435 0.189894
R1100 commonsourceibias.n437 commonsourceibias.n436 0.189894
R1101 commonsourceibias.n437 commonsourceibias.n404 0.189894
R1102 commonsourceibias.n443 commonsourceibias.n404 0.189894
R1103 commonsourceibias.n444 commonsourceibias.n443 0.189894
R1104 commonsourceibias.n445 commonsourceibias.n444 0.189894
R1105 commonsourceibias.n445 commonsourceibias.n402 0.189894
R1106 commonsourceibias.n450 commonsourceibias.n402 0.189894
R1107 commonsourceibias.n451 commonsourceibias.n450 0.189894
R1108 commonsourceibias.n452 commonsourceibias.n451 0.189894
R1109 commonsourceibias.n452 commonsourceibias.n400 0.189894
R1110 commonsourceibias.n458 commonsourceibias.n400 0.189894
R1111 commonsourceibias.n459 commonsourceibias.n458 0.189894
R1112 commonsourceibias.n460 commonsourceibias.n459 0.189894
R1113 commonsourceibias.n460 commonsourceibias.n398 0.189894
R1114 commonsourceibias.n465 commonsourceibias.n398 0.189894
R1115 commonsourceibias.n466 commonsourceibias.n465 0.189894
R1116 commonsourceibias.n467 commonsourceibias.n466 0.189894
R1117 commonsourceibias.n467 commonsourceibias.n396 0.189894
R1118 commonsourceibias.n473 commonsourceibias.n396 0.189894
R1119 commonsourceibias.n474 commonsourceibias.n473 0.189894
R1120 commonsourceibias.n475 commonsourceibias.n474 0.189894
R1121 commonsourceibias.n475 commonsourceibias.n394 0.189894
R1122 commonsourceibias.n480 commonsourceibias.n394 0.189894
R1123 commonsourceibias.n481 commonsourceibias.n480 0.189894
R1124 commonsourceibias.n482 commonsourceibias.n481 0.189894
R1125 commonsourceibias.n482 commonsourceibias.n392 0.189894
R1126 commonsourceibias.n488 commonsourceibias.n392 0.189894
R1127 commonsourceibias.n489 commonsourceibias.n488 0.189894
R1128 commonsourceibias.n490 commonsourceibias.n489 0.189894
R1129 commonsourceibias.n490 commonsourceibias.n390 0.189894
R1130 commonsourceibias.n495 commonsourceibias.n390 0.189894
R1131 commonsourceibias.n496 commonsourceibias.n495 0.189894
R1132 commonsourceibias.n497 commonsourceibias.n496 0.189894
R1133 commonsourceibias.n497 commonsourceibias.n388 0.189894
R1134 commonsourceibias.n531 commonsourceibias.n530 0.189894
R1135 commonsourceibias.n531 commonsourceibias.n526 0.189894
R1136 commonsourceibias.n536 commonsourceibias.n526 0.189894
R1137 commonsourceibias.n537 commonsourceibias.n536 0.189894
R1138 commonsourceibias.n538 commonsourceibias.n537 0.189894
R1139 commonsourceibias.n538 commonsourceibias.n524 0.189894
R1140 commonsourceibias.n544 commonsourceibias.n524 0.189894
R1141 commonsourceibias.n545 commonsourceibias.n544 0.189894
R1142 commonsourceibias.n546 commonsourceibias.n545 0.189894
R1143 commonsourceibias.n546 commonsourceibias.n522 0.189894
R1144 commonsourceibias.n551 commonsourceibias.n522 0.189894
R1145 commonsourceibias.n552 commonsourceibias.n551 0.189894
R1146 commonsourceibias.n553 commonsourceibias.n552 0.189894
R1147 commonsourceibias.n553 commonsourceibias.n520 0.189894
R1148 commonsourceibias.n558 commonsourceibias.n520 0.189894
R1149 commonsourceibias.n559 commonsourceibias.n558 0.189894
R1150 commonsourceibias.n559 commonsourceibias.n518 0.189894
R1151 commonsourceibias.n563 commonsourceibias.n518 0.189894
R1152 commonsourceibias.n564 commonsourceibias.n563 0.189894
R1153 commonsourceibias.n564 commonsourceibias.n516 0.189894
R1154 commonsourceibias.n568 commonsourceibias.n516 0.189894
R1155 commonsourceibias.n569 commonsourceibias.n568 0.189894
R1156 commonsourceibias.n574 commonsourceibias.n573 0.189894
R1157 commonsourceibias.n575 commonsourceibias.n574 0.189894
R1158 commonsourceibias.n575 commonsourceibias.n377 0.189894
R1159 commonsourceibias.n580 commonsourceibias.n377 0.189894
R1160 commonsourceibias.n581 commonsourceibias.n580 0.189894
R1161 commonsourceibias.n582 commonsourceibias.n581 0.189894
R1162 commonsourceibias.n582 commonsourceibias.n375 0.189894
R1163 commonsourceibias.n588 commonsourceibias.n375 0.189894
R1164 commonsourceibias.n589 commonsourceibias.n588 0.189894
R1165 commonsourceibias.n590 commonsourceibias.n589 0.189894
R1166 commonsourceibias.n590 commonsourceibias.n373 0.189894
R1167 commonsourceibias.n595 commonsourceibias.n373 0.189894
R1168 commonsourceibias.n596 commonsourceibias.n595 0.189894
R1169 commonsourceibias.n597 commonsourceibias.n596 0.189894
R1170 commonsourceibias.n597 commonsourceibias.n371 0.189894
R1171 commonsourceibias.n603 commonsourceibias.n371 0.189894
R1172 commonsourceibias.n604 commonsourceibias.n603 0.189894
R1173 commonsourceibias.n605 commonsourceibias.n604 0.189894
R1174 commonsourceibias.n605 commonsourceibias.n369 0.189894
R1175 commonsourceibias.n610 commonsourceibias.n369 0.189894
R1176 commonsourceibias.n611 commonsourceibias.n610 0.189894
R1177 commonsourceibias.n612 commonsourceibias.n611 0.189894
R1178 commonsourceibias.n612 commonsourceibias.n367 0.189894
R1179 commonsourceibias.n205 commonsourceibias.n149 0.0762576
R1180 commonsourceibias.n208 commonsourceibias.n149 0.0762576
R1181 commonsourceibias.n569 commonsourceibias.n514 0.0762576
R1182 commonsourceibias.n573 commonsourceibias.n514 0.0762576
R1183 CSoutput.n19 CSoutput.t158 184.661
R1184 CSoutput.n78 CSoutput.n77 165.8
R1185 CSoutput.n76 CSoutput.n0 165.8
R1186 CSoutput.n75 CSoutput.n74 165.8
R1187 CSoutput.n73 CSoutput.n72 165.8
R1188 CSoutput.n71 CSoutput.n2 165.8
R1189 CSoutput.n69 CSoutput.n68 165.8
R1190 CSoutput.n67 CSoutput.n3 165.8
R1191 CSoutput.n66 CSoutput.n65 165.8
R1192 CSoutput.n63 CSoutput.n4 165.8
R1193 CSoutput.n61 CSoutput.n60 165.8
R1194 CSoutput.n59 CSoutput.n5 165.8
R1195 CSoutput.n58 CSoutput.n57 165.8
R1196 CSoutput.n55 CSoutput.n6 165.8
R1197 CSoutput.n54 CSoutput.n53 165.8
R1198 CSoutput.n52 CSoutput.n51 165.8
R1199 CSoutput.n50 CSoutput.n8 165.8
R1200 CSoutput.n48 CSoutput.n47 165.8
R1201 CSoutput.n46 CSoutput.n9 165.8
R1202 CSoutput.n45 CSoutput.n44 165.8
R1203 CSoutput.n42 CSoutput.n10 165.8
R1204 CSoutput.n41 CSoutput.n40 165.8
R1205 CSoutput.n39 CSoutput.n38 165.8
R1206 CSoutput.n37 CSoutput.n12 165.8
R1207 CSoutput.n35 CSoutput.n34 165.8
R1208 CSoutput.n33 CSoutput.n13 165.8
R1209 CSoutput.n32 CSoutput.n31 165.8
R1210 CSoutput.n29 CSoutput.n14 165.8
R1211 CSoutput.n28 CSoutput.n27 165.8
R1212 CSoutput.n26 CSoutput.n25 165.8
R1213 CSoutput.n24 CSoutput.n16 165.8
R1214 CSoutput.n22 CSoutput.n21 165.8
R1215 CSoutput.n20 CSoutput.n17 165.8
R1216 CSoutput.n77 CSoutput.t160 162.194
R1217 CSoutput.n18 CSoutput.t169 120.501
R1218 CSoutput.n23 CSoutput.t171 120.501
R1219 CSoutput.n15 CSoutput.t164 120.501
R1220 CSoutput.n30 CSoutput.t155 120.501
R1221 CSoutput.n36 CSoutput.t173 120.501
R1222 CSoutput.n11 CSoutput.t167 120.501
R1223 CSoutput.n43 CSoutput.t162 120.501
R1224 CSoutput.n49 CSoutput.t153 120.501
R1225 CSoutput.n7 CSoutput.t154 120.501
R1226 CSoutput.n56 CSoutput.t165 120.501
R1227 CSoutput.n62 CSoutput.t161 120.501
R1228 CSoutput.n64 CSoutput.t157 120.501
R1229 CSoutput.n70 CSoutput.t168 120.501
R1230 CSoutput.n1 CSoutput.t170 120.501
R1231 CSoutput.n290 CSoutput.n288 103.469
R1232 CSoutput.n278 CSoutput.n276 103.469
R1233 CSoutput.n267 CSoutput.n265 103.469
R1234 CSoutput.n104 CSoutput.n102 103.469
R1235 CSoutput.n92 CSoutput.n90 103.469
R1236 CSoutput.n81 CSoutput.n79 103.469
R1237 CSoutput.n296 CSoutput.n295 103.111
R1238 CSoutput.n294 CSoutput.n293 103.111
R1239 CSoutput.n292 CSoutput.n291 103.111
R1240 CSoutput.n290 CSoutput.n289 103.111
R1241 CSoutput.n286 CSoutput.n285 103.111
R1242 CSoutput.n284 CSoutput.n283 103.111
R1243 CSoutput.n282 CSoutput.n281 103.111
R1244 CSoutput.n280 CSoutput.n279 103.111
R1245 CSoutput.n278 CSoutput.n277 103.111
R1246 CSoutput.n275 CSoutput.n274 103.111
R1247 CSoutput.n273 CSoutput.n272 103.111
R1248 CSoutput.n271 CSoutput.n270 103.111
R1249 CSoutput.n269 CSoutput.n268 103.111
R1250 CSoutput.n267 CSoutput.n266 103.111
R1251 CSoutput.n104 CSoutput.n103 103.111
R1252 CSoutput.n106 CSoutput.n105 103.111
R1253 CSoutput.n108 CSoutput.n107 103.111
R1254 CSoutput.n110 CSoutput.n109 103.111
R1255 CSoutput.n112 CSoutput.n111 103.111
R1256 CSoutput.n92 CSoutput.n91 103.111
R1257 CSoutput.n94 CSoutput.n93 103.111
R1258 CSoutput.n96 CSoutput.n95 103.111
R1259 CSoutput.n98 CSoutput.n97 103.111
R1260 CSoutput.n100 CSoutput.n99 103.111
R1261 CSoutput.n81 CSoutput.n80 103.111
R1262 CSoutput.n83 CSoutput.n82 103.111
R1263 CSoutput.n85 CSoutput.n84 103.111
R1264 CSoutput.n87 CSoutput.n86 103.111
R1265 CSoutput.n89 CSoutput.n88 103.111
R1266 CSoutput.n298 CSoutput.n297 103.111
R1267 CSoutput.n322 CSoutput.n320 81.5057
R1268 CSoutput.n303 CSoutput.n301 81.5057
R1269 CSoutput.n362 CSoutput.n360 81.5057
R1270 CSoutput.n343 CSoutput.n341 81.5057
R1271 CSoutput.n338 CSoutput.n337 80.9324
R1272 CSoutput.n336 CSoutput.n335 80.9324
R1273 CSoutput.n334 CSoutput.n333 80.9324
R1274 CSoutput.n332 CSoutput.n331 80.9324
R1275 CSoutput.n330 CSoutput.n329 80.9324
R1276 CSoutput.n328 CSoutput.n327 80.9324
R1277 CSoutput.n326 CSoutput.n325 80.9324
R1278 CSoutput.n324 CSoutput.n323 80.9324
R1279 CSoutput.n322 CSoutput.n321 80.9324
R1280 CSoutput.n319 CSoutput.n318 80.9324
R1281 CSoutput.n317 CSoutput.n316 80.9324
R1282 CSoutput.n315 CSoutput.n314 80.9324
R1283 CSoutput.n313 CSoutput.n312 80.9324
R1284 CSoutput.n311 CSoutput.n310 80.9324
R1285 CSoutput.n309 CSoutput.n308 80.9324
R1286 CSoutput.n307 CSoutput.n306 80.9324
R1287 CSoutput.n305 CSoutput.n304 80.9324
R1288 CSoutput.n303 CSoutput.n302 80.9324
R1289 CSoutput.n362 CSoutput.n361 80.9324
R1290 CSoutput.n364 CSoutput.n363 80.9324
R1291 CSoutput.n366 CSoutput.n365 80.9324
R1292 CSoutput.n368 CSoutput.n367 80.9324
R1293 CSoutput.n370 CSoutput.n369 80.9324
R1294 CSoutput.n372 CSoutput.n371 80.9324
R1295 CSoutput.n374 CSoutput.n373 80.9324
R1296 CSoutput.n376 CSoutput.n375 80.9324
R1297 CSoutput.n378 CSoutput.n377 80.9324
R1298 CSoutput.n343 CSoutput.n342 80.9324
R1299 CSoutput.n345 CSoutput.n344 80.9324
R1300 CSoutput.n347 CSoutput.n346 80.9324
R1301 CSoutput.n349 CSoutput.n348 80.9324
R1302 CSoutput.n351 CSoutput.n350 80.9324
R1303 CSoutput.n353 CSoutput.n352 80.9324
R1304 CSoutput.n355 CSoutput.n354 80.9324
R1305 CSoutput.n357 CSoutput.n356 80.9324
R1306 CSoutput.n359 CSoutput.n358 80.9324
R1307 CSoutput.n25 CSoutput.n24 48.1486
R1308 CSoutput.n69 CSoutput.n3 48.1486
R1309 CSoutput.n38 CSoutput.n37 48.1486
R1310 CSoutput.n42 CSoutput.n41 48.1486
R1311 CSoutput.n51 CSoutput.n50 48.1486
R1312 CSoutput.n55 CSoutput.n54 48.1486
R1313 CSoutput.n22 CSoutput.n17 46.462
R1314 CSoutput.n72 CSoutput.n71 46.462
R1315 CSoutput.n20 CSoutput.n19 44.9055
R1316 CSoutput.n29 CSoutput.n28 43.7635
R1317 CSoutput.n65 CSoutput.n63 43.7635
R1318 CSoutput.n35 CSoutput.n13 41.7396
R1319 CSoutput.n57 CSoutput.n5 41.7396
R1320 CSoutput.n44 CSoutput.n9 37.0171
R1321 CSoutput.n48 CSoutput.n9 37.0171
R1322 CSoutput.n76 CSoutput.n75 34.9932
R1323 CSoutput.n31 CSoutput.n13 32.2947
R1324 CSoutput.n61 CSoutput.n5 32.2947
R1325 CSoutput.n30 CSoutput.n29 29.6014
R1326 CSoutput.n63 CSoutput.n62 29.6014
R1327 CSoutput.n19 CSoutput.n18 28.4085
R1328 CSoutput.n18 CSoutput.n17 25.1176
R1329 CSoutput.n72 CSoutput.n1 25.1176
R1330 CSoutput.n43 CSoutput.n42 22.0922
R1331 CSoutput.n50 CSoutput.n49 22.0922
R1332 CSoutput.n77 CSoutput.n76 21.8586
R1333 CSoutput.n37 CSoutput.n36 18.9681
R1334 CSoutput.n56 CSoutput.n55 18.9681
R1335 CSoutput.n25 CSoutput.n15 17.6292
R1336 CSoutput.n64 CSoutput.n3 17.6292
R1337 CSoutput.n24 CSoutput.n23 15.844
R1338 CSoutput.n70 CSoutput.n69 15.844
R1339 CSoutput.n38 CSoutput.n11 14.5051
R1340 CSoutput.n54 CSoutput.n7 14.5051
R1341 CSoutput.n381 CSoutput.n78 11.6139
R1342 CSoutput.n41 CSoutput.n11 11.3811
R1343 CSoutput.n51 CSoutput.n7 11.3811
R1344 CSoutput.n23 CSoutput.n22 10.0422
R1345 CSoutput.n71 CSoutput.n70 10.0422
R1346 CSoutput.n287 CSoutput.n275 9.25285
R1347 CSoutput.n101 CSoutput.n89 9.25285
R1348 CSoutput.n340 CSoutput.n300 9.05363
R1349 CSoutput.n339 CSoutput.n319 8.97993
R1350 CSoutput.n379 CSoutput.n359 8.97993
R1351 CSoutput.n28 CSoutput.n15 8.25698
R1352 CSoutput.n65 CSoutput.n64 8.25698
R1353 CSoutput.n340 CSoutput.n339 7.89345
R1354 CSoutput.n380 CSoutput.n379 7.89345
R1355 CSoutput.n300 CSoutput.n299 7.12641
R1356 CSoutput.n114 CSoutput.n113 7.12641
R1357 CSoutput.n36 CSoutput.n35 6.91809
R1358 CSoutput.n57 CSoutput.n56 6.91809
R1359 CSoutput.n381 CSoutput.n114 5.46119
R1360 CSoutput.n339 CSoutput.n338 5.25266
R1361 CSoutput.n379 CSoutput.n378 5.25266
R1362 CSoutput.n299 CSoutput.n298 5.1449
R1363 CSoutput.n287 CSoutput.n286 5.1449
R1364 CSoutput.n113 CSoutput.n112 5.1449
R1365 CSoutput.n101 CSoutput.n100 5.1449
R1366 CSoutput.n205 CSoutput.n158 4.5005
R1367 CSoutput.n174 CSoutput.n158 4.5005
R1368 CSoutput.n169 CSoutput.n153 4.5005
R1369 CSoutput.n169 CSoutput.n155 4.5005
R1370 CSoutput.n169 CSoutput.n152 4.5005
R1371 CSoutput.n169 CSoutput.n156 4.5005
R1372 CSoutput.n169 CSoutput.n151 4.5005
R1373 CSoutput.n169 CSoutput.t172 4.5005
R1374 CSoutput.n169 CSoutput.n150 4.5005
R1375 CSoutput.n169 CSoutput.n157 4.5005
R1376 CSoutput.n169 CSoutput.n158 4.5005
R1377 CSoutput.n167 CSoutput.n153 4.5005
R1378 CSoutput.n167 CSoutput.n155 4.5005
R1379 CSoutput.n167 CSoutput.n152 4.5005
R1380 CSoutput.n167 CSoutput.n156 4.5005
R1381 CSoutput.n167 CSoutput.n151 4.5005
R1382 CSoutput.n167 CSoutput.t172 4.5005
R1383 CSoutput.n167 CSoutput.n150 4.5005
R1384 CSoutput.n167 CSoutput.n157 4.5005
R1385 CSoutput.n167 CSoutput.n158 4.5005
R1386 CSoutput.n166 CSoutput.n153 4.5005
R1387 CSoutput.n166 CSoutput.n155 4.5005
R1388 CSoutput.n166 CSoutput.n152 4.5005
R1389 CSoutput.n166 CSoutput.n156 4.5005
R1390 CSoutput.n166 CSoutput.n151 4.5005
R1391 CSoutput.n166 CSoutput.t172 4.5005
R1392 CSoutput.n166 CSoutput.n150 4.5005
R1393 CSoutput.n166 CSoutput.n157 4.5005
R1394 CSoutput.n166 CSoutput.n158 4.5005
R1395 CSoutput.n251 CSoutput.n153 4.5005
R1396 CSoutput.n251 CSoutput.n155 4.5005
R1397 CSoutput.n251 CSoutput.n152 4.5005
R1398 CSoutput.n251 CSoutput.n156 4.5005
R1399 CSoutput.n251 CSoutput.n151 4.5005
R1400 CSoutput.n251 CSoutput.t172 4.5005
R1401 CSoutput.n251 CSoutput.n150 4.5005
R1402 CSoutput.n251 CSoutput.n157 4.5005
R1403 CSoutput.n251 CSoutput.n158 4.5005
R1404 CSoutput.n249 CSoutput.n153 4.5005
R1405 CSoutput.n249 CSoutput.n155 4.5005
R1406 CSoutput.n249 CSoutput.n152 4.5005
R1407 CSoutput.n249 CSoutput.n156 4.5005
R1408 CSoutput.n249 CSoutput.n151 4.5005
R1409 CSoutput.n249 CSoutput.t172 4.5005
R1410 CSoutput.n249 CSoutput.n150 4.5005
R1411 CSoutput.n249 CSoutput.n157 4.5005
R1412 CSoutput.n247 CSoutput.n153 4.5005
R1413 CSoutput.n247 CSoutput.n155 4.5005
R1414 CSoutput.n247 CSoutput.n152 4.5005
R1415 CSoutput.n247 CSoutput.n156 4.5005
R1416 CSoutput.n247 CSoutput.n151 4.5005
R1417 CSoutput.n247 CSoutput.t172 4.5005
R1418 CSoutput.n247 CSoutput.n150 4.5005
R1419 CSoutput.n247 CSoutput.n157 4.5005
R1420 CSoutput.n177 CSoutput.n153 4.5005
R1421 CSoutput.n177 CSoutput.n155 4.5005
R1422 CSoutput.n177 CSoutput.n152 4.5005
R1423 CSoutput.n177 CSoutput.n156 4.5005
R1424 CSoutput.n177 CSoutput.n151 4.5005
R1425 CSoutput.n177 CSoutput.t172 4.5005
R1426 CSoutput.n177 CSoutput.n150 4.5005
R1427 CSoutput.n177 CSoutput.n157 4.5005
R1428 CSoutput.n177 CSoutput.n158 4.5005
R1429 CSoutput.n176 CSoutput.n153 4.5005
R1430 CSoutput.n176 CSoutput.n155 4.5005
R1431 CSoutput.n176 CSoutput.n152 4.5005
R1432 CSoutput.n176 CSoutput.n156 4.5005
R1433 CSoutput.n176 CSoutput.n151 4.5005
R1434 CSoutput.n176 CSoutput.t172 4.5005
R1435 CSoutput.n176 CSoutput.n150 4.5005
R1436 CSoutput.n176 CSoutput.n157 4.5005
R1437 CSoutput.n176 CSoutput.n158 4.5005
R1438 CSoutput.n180 CSoutput.n153 4.5005
R1439 CSoutput.n180 CSoutput.n155 4.5005
R1440 CSoutput.n180 CSoutput.n152 4.5005
R1441 CSoutput.n180 CSoutput.n156 4.5005
R1442 CSoutput.n180 CSoutput.n151 4.5005
R1443 CSoutput.n180 CSoutput.t172 4.5005
R1444 CSoutput.n180 CSoutput.n150 4.5005
R1445 CSoutput.n180 CSoutput.n157 4.5005
R1446 CSoutput.n180 CSoutput.n158 4.5005
R1447 CSoutput.n179 CSoutput.n153 4.5005
R1448 CSoutput.n179 CSoutput.n155 4.5005
R1449 CSoutput.n179 CSoutput.n152 4.5005
R1450 CSoutput.n179 CSoutput.n156 4.5005
R1451 CSoutput.n179 CSoutput.n151 4.5005
R1452 CSoutput.n179 CSoutput.t172 4.5005
R1453 CSoutput.n179 CSoutput.n150 4.5005
R1454 CSoutput.n179 CSoutput.n157 4.5005
R1455 CSoutput.n179 CSoutput.n158 4.5005
R1456 CSoutput.n162 CSoutput.n153 4.5005
R1457 CSoutput.n162 CSoutput.n155 4.5005
R1458 CSoutput.n162 CSoutput.n152 4.5005
R1459 CSoutput.n162 CSoutput.n156 4.5005
R1460 CSoutput.n162 CSoutput.n151 4.5005
R1461 CSoutput.n162 CSoutput.t172 4.5005
R1462 CSoutput.n162 CSoutput.n150 4.5005
R1463 CSoutput.n162 CSoutput.n157 4.5005
R1464 CSoutput.n162 CSoutput.n158 4.5005
R1465 CSoutput.n254 CSoutput.n153 4.5005
R1466 CSoutput.n254 CSoutput.n155 4.5005
R1467 CSoutput.n254 CSoutput.n152 4.5005
R1468 CSoutput.n254 CSoutput.n156 4.5005
R1469 CSoutput.n254 CSoutput.n151 4.5005
R1470 CSoutput.n254 CSoutput.t172 4.5005
R1471 CSoutput.n254 CSoutput.n150 4.5005
R1472 CSoutput.n254 CSoutput.n157 4.5005
R1473 CSoutput.n254 CSoutput.n158 4.5005
R1474 CSoutput.n241 CSoutput.n212 4.5005
R1475 CSoutput.n241 CSoutput.n218 4.5005
R1476 CSoutput.n199 CSoutput.n188 4.5005
R1477 CSoutput.n199 CSoutput.n190 4.5005
R1478 CSoutput.n199 CSoutput.n187 4.5005
R1479 CSoutput.n199 CSoutput.n191 4.5005
R1480 CSoutput.n199 CSoutput.n186 4.5005
R1481 CSoutput.n199 CSoutput.t166 4.5005
R1482 CSoutput.n199 CSoutput.n185 4.5005
R1483 CSoutput.n199 CSoutput.n192 4.5005
R1484 CSoutput.n241 CSoutput.n199 4.5005
R1485 CSoutput.n220 CSoutput.n188 4.5005
R1486 CSoutput.n220 CSoutput.n190 4.5005
R1487 CSoutput.n220 CSoutput.n187 4.5005
R1488 CSoutput.n220 CSoutput.n191 4.5005
R1489 CSoutput.n220 CSoutput.n186 4.5005
R1490 CSoutput.n220 CSoutput.t166 4.5005
R1491 CSoutput.n220 CSoutput.n185 4.5005
R1492 CSoutput.n220 CSoutput.n192 4.5005
R1493 CSoutput.n241 CSoutput.n220 4.5005
R1494 CSoutput.n198 CSoutput.n188 4.5005
R1495 CSoutput.n198 CSoutput.n190 4.5005
R1496 CSoutput.n198 CSoutput.n187 4.5005
R1497 CSoutput.n198 CSoutput.n191 4.5005
R1498 CSoutput.n198 CSoutput.n186 4.5005
R1499 CSoutput.n198 CSoutput.t166 4.5005
R1500 CSoutput.n198 CSoutput.n185 4.5005
R1501 CSoutput.n198 CSoutput.n192 4.5005
R1502 CSoutput.n241 CSoutput.n198 4.5005
R1503 CSoutput.n222 CSoutput.n188 4.5005
R1504 CSoutput.n222 CSoutput.n190 4.5005
R1505 CSoutput.n222 CSoutput.n187 4.5005
R1506 CSoutput.n222 CSoutput.n191 4.5005
R1507 CSoutput.n222 CSoutput.n186 4.5005
R1508 CSoutput.n222 CSoutput.t166 4.5005
R1509 CSoutput.n222 CSoutput.n185 4.5005
R1510 CSoutput.n222 CSoutput.n192 4.5005
R1511 CSoutput.n241 CSoutput.n222 4.5005
R1512 CSoutput.n188 CSoutput.n183 4.5005
R1513 CSoutput.n190 CSoutput.n183 4.5005
R1514 CSoutput.n187 CSoutput.n183 4.5005
R1515 CSoutput.n191 CSoutput.n183 4.5005
R1516 CSoutput.n186 CSoutput.n183 4.5005
R1517 CSoutput.t166 CSoutput.n183 4.5005
R1518 CSoutput.n185 CSoutput.n183 4.5005
R1519 CSoutput.n192 CSoutput.n183 4.5005
R1520 CSoutput.n244 CSoutput.n188 4.5005
R1521 CSoutput.n244 CSoutput.n190 4.5005
R1522 CSoutput.n244 CSoutput.n187 4.5005
R1523 CSoutput.n244 CSoutput.n191 4.5005
R1524 CSoutput.n244 CSoutput.n186 4.5005
R1525 CSoutput.n244 CSoutput.t166 4.5005
R1526 CSoutput.n244 CSoutput.n185 4.5005
R1527 CSoutput.n244 CSoutput.n192 4.5005
R1528 CSoutput.n242 CSoutput.n188 4.5005
R1529 CSoutput.n242 CSoutput.n190 4.5005
R1530 CSoutput.n242 CSoutput.n187 4.5005
R1531 CSoutput.n242 CSoutput.n191 4.5005
R1532 CSoutput.n242 CSoutput.n186 4.5005
R1533 CSoutput.n242 CSoutput.t166 4.5005
R1534 CSoutput.n242 CSoutput.n185 4.5005
R1535 CSoutput.n242 CSoutput.n192 4.5005
R1536 CSoutput.n242 CSoutput.n241 4.5005
R1537 CSoutput.n224 CSoutput.n188 4.5005
R1538 CSoutput.n224 CSoutput.n190 4.5005
R1539 CSoutput.n224 CSoutput.n187 4.5005
R1540 CSoutput.n224 CSoutput.n191 4.5005
R1541 CSoutput.n224 CSoutput.n186 4.5005
R1542 CSoutput.n224 CSoutput.t166 4.5005
R1543 CSoutput.n224 CSoutput.n185 4.5005
R1544 CSoutput.n224 CSoutput.n192 4.5005
R1545 CSoutput.n241 CSoutput.n224 4.5005
R1546 CSoutput.n196 CSoutput.n188 4.5005
R1547 CSoutput.n196 CSoutput.n190 4.5005
R1548 CSoutput.n196 CSoutput.n187 4.5005
R1549 CSoutput.n196 CSoutput.n191 4.5005
R1550 CSoutput.n196 CSoutput.n186 4.5005
R1551 CSoutput.n196 CSoutput.t166 4.5005
R1552 CSoutput.n196 CSoutput.n185 4.5005
R1553 CSoutput.n196 CSoutput.n192 4.5005
R1554 CSoutput.n241 CSoutput.n196 4.5005
R1555 CSoutput.n226 CSoutput.n188 4.5005
R1556 CSoutput.n226 CSoutput.n190 4.5005
R1557 CSoutput.n226 CSoutput.n187 4.5005
R1558 CSoutput.n226 CSoutput.n191 4.5005
R1559 CSoutput.n226 CSoutput.n186 4.5005
R1560 CSoutput.n226 CSoutput.t166 4.5005
R1561 CSoutput.n226 CSoutput.n185 4.5005
R1562 CSoutput.n226 CSoutput.n192 4.5005
R1563 CSoutput.n241 CSoutput.n226 4.5005
R1564 CSoutput.n195 CSoutput.n188 4.5005
R1565 CSoutput.n195 CSoutput.n190 4.5005
R1566 CSoutput.n195 CSoutput.n187 4.5005
R1567 CSoutput.n195 CSoutput.n191 4.5005
R1568 CSoutput.n195 CSoutput.n186 4.5005
R1569 CSoutput.n195 CSoutput.t166 4.5005
R1570 CSoutput.n195 CSoutput.n185 4.5005
R1571 CSoutput.n195 CSoutput.n192 4.5005
R1572 CSoutput.n241 CSoutput.n195 4.5005
R1573 CSoutput.n240 CSoutput.n188 4.5005
R1574 CSoutput.n240 CSoutput.n190 4.5005
R1575 CSoutput.n240 CSoutput.n187 4.5005
R1576 CSoutput.n240 CSoutput.n191 4.5005
R1577 CSoutput.n240 CSoutput.n186 4.5005
R1578 CSoutput.n240 CSoutput.t166 4.5005
R1579 CSoutput.n240 CSoutput.n185 4.5005
R1580 CSoutput.n240 CSoutput.n192 4.5005
R1581 CSoutput.n241 CSoutput.n240 4.5005
R1582 CSoutput.n239 CSoutput.n124 4.5005
R1583 CSoutput.n140 CSoutput.n124 4.5005
R1584 CSoutput.n135 CSoutput.n119 4.5005
R1585 CSoutput.n135 CSoutput.n121 4.5005
R1586 CSoutput.n135 CSoutput.n118 4.5005
R1587 CSoutput.n135 CSoutput.n122 4.5005
R1588 CSoutput.n135 CSoutput.n117 4.5005
R1589 CSoutput.n135 CSoutput.t163 4.5005
R1590 CSoutput.n135 CSoutput.n116 4.5005
R1591 CSoutput.n135 CSoutput.n123 4.5005
R1592 CSoutput.n135 CSoutput.n124 4.5005
R1593 CSoutput.n133 CSoutput.n119 4.5005
R1594 CSoutput.n133 CSoutput.n121 4.5005
R1595 CSoutput.n133 CSoutput.n118 4.5005
R1596 CSoutput.n133 CSoutput.n122 4.5005
R1597 CSoutput.n133 CSoutput.n117 4.5005
R1598 CSoutput.n133 CSoutput.t163 4.5005
R1599 CSoutput.n133 CSoutput.n116 4.5005
R1600 CSoutput.n133 CSoutput.n123 4.5005
R1601 CSoutput.n133 CSoutput.n124 4.5005
R1602 CSoutput.n132 CSoutput.n119 4.5005
R1603 CSoutput.n132 CSoutput.n121 4.5005
R1604 CSoutput.n132 CSoutput.n118 4.5005
R1605 CSoutput.n132 CSoutput.n122 4.5005
R1606 CSoutput.n132 CSoutput.n117 4.5005
R1607 CSoutput.n132 CSoutput.t163 4.5005
R1608 CSoutput.n132 CSoutput.n116 4.5005
R1609 CSoutput.n132 CSoutput.n123 4.5005
R1610 CSoutput.n132 CSoutput.n124 4.5005
R1611 CSoutput.n261 CSoutput.n119 4.5005
R1612 CSoutput.n261 CSoutput.n121 4.5005
R1613 CSoutput.n261 CSoutput.n118 4.5005
R1614 CSoutput.n261 CSoutput.n122 4.5005
R1615 CSoutput.n261 CSoutput.n117 4.5005
R1616 CSoutput.n261 CSoutput.t163 4.5005
R1617 CSoutput.n261 CSoutput.n116 4.5005
R1618 CSoutput.n261 CSoutput.n123 4.5005
R1619 CSoutput.n261 CSoutput.n124 4.5005
R1620 CSoutput.n259 CSoutput.n119 4.5005
R1621 CSoutput.n259 CSoutput.n121 4.5005
R1622 CSoutput.n259 CSoutput.n118 4.5005
R1623 CSoutput.n259 CSoutput.n122 4.5005
R1624 CSoutput.n259 CSoutput.n117 4.5005
R1625 CSoutput.n259 CSoutput.t163 4.5005
R1626 CSoutput.n259 CSoutput.n116 4.5005
R1627 CSoutput.n259 CSoutput.n123 4.5005
R1628 CSoutput.n257 CSoutput.n119 4.5005
R1629 CSoutput.n257 CSoutput.n121 4.5005
R1630 CSoutput.n257 CSoutput.n118 4.5005
R1631 CSoutput.n257 CSoutput.n122 4.5005
R1632 CSoutput.n257 CSoutput.n117 4.5005
R1633 CSoutput.n257 CSoutput.t163 4.5005
R1634 CSoutput.n257 CSoutput.n116 4.5005
R1635 CSoutput.n257 CSoutput.n123 4.5005
R1636 CSoutput.n143 CSoutput.n119 4.5005
R1637 CSoutput.n143 CSoutput.n121 4.5005
R1638 CSoutput.n143 CSoutput.n118 4.5005
R1639 CSoutput.n143 CSoutput.n122 4.5005
R1640 CSoutput.n143 CSoutput.n117 4.5005
R1641 CSoutput.n143 CSoutput.t163 4.5005
R1642 CSoutput.n143 CSoutput.n116 4.5005
R1643 CSoutput.n143 CSoutput.n123 4.5005
R1644 CSoutput.n143 CSoutput.n124 4.5005
R1645 CSoutput.n142 CSoutput.n119 4.5005
R1646 CSoutput.n142 CSoutput.n121 4.5005
R1647 CSoutput.n142 CSoutput.n118 4.5005
R1648 CSoutput.n142 CSoutput.n122 4.5005
R1649 CSoutput.n142 CSoutput.n117 4.5005
R1650 CSoutput.n142 CSoutput.t163 4.5005
R1651 CSoutput.n142 CSoutput.n116 4.5005
R1652 CSoutput.n142 CSoutput.n123 4.5005
R1653 CSoutput.n142 CSoutput.n124 4.5005
R1654 CSoutput.n146 CSoutput.n119 4.5005
R1655 CSoutput.n146 CSoutput.n121 4.5005
R1656 CSoutput.n146 CSoutput.n118 4.5005
R1657 CSoutput.n146 CSoutput.n122 4.5005
R1658 CSoutput.n146 CSoutput.n117 4.5005
R1659 CSoutput.n146 CSoutput.t163 4.5005
R1660 CSoutput.n146 CSoutput.n116 4.5005
R1661 CSoutput.n146 CSoutput.n123 4.5005
R1662 CSoutput.n146 CSoutput.n124 4.5005
R1663 CSoutput.n145 CSoutput.n119 4.5005
R1664 CSoutput.n145 CSoutput.n121 4.5005
R1665 CSoutput.n145 CSoutput.n118 4.5005
R1666 CSoutput.n145 CSoutput.n122 4.5005
R1667 CSoutput.n145 CSoutput.n117 4.5005
R1668 CSoutput.n145 CSoutput.t163 4.5005
R1669 CSoutput.n145 CSoutput.n116 4.5005
R1670 CSoutput.n145 CSoutput.n123 4.5005
R1671 CSoutput.n145 CSoutput.n124 4.5005
R1672 CSoutput.n128 CSoutput.n119 4.5005
R1673 CSoutput.n128 CSoutput.n121 4.5005
R1674 CSoutput.n128 CSoutput.n118 4.5005
R1675 CSoutput.n128 CSoutput.n122 4.5005
R1676 CSoutput.n128 CSoutput.n117 4.5005
R1677 CSoutput.n128 CSoutput.t163 4.5005
R1678 CSoutput.n128 CSoutput.n116 4.5005
R1679 CSoutput.n128 CSoutput.n123 4.5005
R1680 CSoutput.n128 CSoutput.n124 4.5005
R1681 CSoutput.n264 CSoutput.n119 4.5005
R1682 CSoutput.n264 CSoutput.n121 4.5005
R1683 CSoutput.n264 CSoutput.n118 4.5005
R1684 CSoutput.n264 CSoutput.n122 4.5005
R1685 CSoutput.n264 CSoutput.n117 4.5005
R1686 CSoutput.n264 CSoutput.t163 4.5005
R1687 CSoutput.n264 CSoutput.n116 4.5005
R1688 CSoutput.n264 CSoutput.n123 4.5005
R1689 CSoutput.n264 CSoutput.n124 4.5005
R1690 CSoutput.n299 CSoutput.n287 4.10845
R1691 CSoutput.n113 CSoutput.n101 4.10845
R1692 CSoutput.n297 CSoutput.t32 4.06363
R1693 CSoutput.n297 CSoutput.t47 4.06363
R1694 CSoutput.n295 CSoutput.t0 4.06363
R1695 CSoutput.n295 CSoutput.t39 4.06363
R1696 CSoutput.n293 CSoutput.t59 4.06363
R1697 CSoutput.n293 CSoutput.t8 4.06363
R1698 CSoutput.n291 CSoutput.t53 4.06363
R1699 CSoutput.n291 CSoutput.t52 4.06363
R1700 CSoutput.n289 CSoutput.t7 4.06363
R1701 CSoutput.n289 CSoutput.t17 4.06363
R1702 CSoutput.n288 CSoutput.t16 4.06363
R1703 CSoutput.n288 CSoutput.t11 4.06363
R1704 CSoutput.n285 CSoutput.t6 4.06363
R1705 CSoutput.n285 CSoutput.t14 4.06363
R1706 CSoutput.n283 CSoutput.t15 4.06363
R1707 CSoutput.n283 CSoutput.t2 4.06363
R1708 CSoutput.n281 CSoutput.t26 4.06363
R1709 CSoutput.n281 CSoutput.t58 4.06363
R1710 CSoutput.n279 CSoutput.t49 4.06363
R1711 CSoutput.n279 CSoutput.t13 4.06363
R1712 CSoutput.n277 CSoutput.t147 4.06363
R1713 CSoutput.n277 CSoutput.t37 4.06363
R1714 CSoutput.n276 CSoutput.t42 4.06363
R1715 CSoutput.n276 CSoutput.t36 4.06363
R1716 CSoutput.n274 CSoutput.t41 4.06363
R1717 CSoutput.n274 CSoutput.t38 4.06363
R1718 CSoutput.n272 CSoutput.t61 4.06363
R1719 CSoutput.n272 CSoutput.t25 4.06363
R1720 CSoutput.n270 CSoutput.t54 4.06363
R1721 CSoutput.n270 CSoutput.t23 4.06363
R1722 CSoutput.n268 CSoutput.t29 4.06363
R1723 CSoutput.n268 CSoutput.t148 4.06363
R1724 CSoutput.n266 CSoutput.t4 4.06363
R1725 CSoutput.n266 CSoutput.t10 4.06363
R1726 CSoutput.n265 CSoutput.t40 4.06363
R1727 CSoutput.n265 CSoutput.t149 4.06363
R1728 CSoutput.n102 CSoutput.t9 4.06363
R1729 CSoutput.n102 CSoutput.t48 4.06363
R1730 CSoutput.n103 CSoutput.t145 4.06363
R1731 CSoutput.n103 CSoutput.t51 4.06363
R1732 CSoutput.n105 CSoutput.t43 4.06363
R1733 CSoutput.n105 CSoutput.t150 4.06363
R1734 CSoutput.n107 CSoutput.t142 4.06363
R1735 CSoutput.n107 CSoutput.t20 4.06363
R1736 CSoutput.n109 CSoutput.t22 4.06363
R1737 CSoutput.n109 CSoutput.t151 4.06363
R1738 CSoutput.n111 CSoutput.t46 4.06363
R1739 CSoutput.n111 CSoutput.t146 4.06363
R1740 CSoutput.n90 CSoutput.t55 4.06363
R1741 CSoutput.n90 CSoutput.t144 4.06363
R1742 CSoutput.n91 CSoutput.t12 4.06363
R1743 CSoutput.n91 CSoutput.t19 4.06363
R1744 CSoutput.n93 CSoutput.t34 4.06363
R1745 CSoutput.n93 CSoutput.t45 4.06363
R1746 CSoutput.n95 CSoutput.t5 4.06363
R1747 CSoutput.n95 CSoutput.t28 4.06363
R1748 CSoutput.n97 CSoutput.t35 4.06363
R1749 CSoutput.n97 CSoutput.t27 4.06363
R1750 CSoutput.n99 CSoutput.t3 4.06363
R1751 CSoutput.n99 CSoutput.t31 4.06363
R1752 CSoutput.n79 CSoutput.t44 4.06363
R1753 CSoutput.n79 CSoutput.t33 4.06363
R1754 CSoutput.n80 CSoutput.t21 4.06363
R1755 CSoutput.n80 CSoutput.t1 4.06363
R1756 CSoutput.n82 CSoutput.t30 4.06363
R1757 CSoutput.n82 CSoutput.t50 4.06363
R1758 CSoutput.n84 CSoutput.t18 4.06363
R1759 CSoutput.n84 CSoutput.t56 4.06363
R1760 CSoutput.n86 CSoutput.t24 4.06363
R1761 CSoutput.n86 CSoutput.t60 4.06363
R1762 CSoutput.n88 CSoutput.t57 4.06363
R1763 CSoutput.n88 CSoutput.t143 4.06363
R1764 CSoutput.n44 CSoutput.n43 3.79402
R1765 CSoutput.n49 CSoutput.n48 3.79402
R1766 CSoutput.n381 CSoutput.n380 3.57343
R1767 CSoutput.n380 CSoutput.n340 3.42304
R1768 CSoutput.n337 CSoutput.t72 2.82907
R1769 CSoutput.n337 CSoutput.t137 2.82907
R1770 CSoutput.n335 CSoutput.t127 2.82907
R1771 CSoutput.n335 CSoutput.t87 2.82907
R1772 CSoutput.n333 CSoutput.t102 2.82907
R1773 CSoutput.n333 CSoutput.t107 2.82907
R1774 CSoutput.n331 CSoutput.t135 2.82907
R1775 CSoutput.n331 CSoutput.t117 2.82907
R1776 CSoutput.n329 CSoutput.t110 2.82907
R1777 CSoutput.n329 CSoutput.t113 2.82907
R1778 CSoutput.n327 CSoutput.t108 2.82907
R1779 CSoutput.n327 CSoutput.t126 2.82907
R1780 CSoutput.n325 CSoutput.t73 2.82907
R1781 CSoutput.n325 CSoutput.t139 2.82907
R1782 CSoutput.n323 CSoutput.t130 2.82907
R1783 CSoutput.n323 CSoutput.t66 2.82907
R1784 CSoutput.n321 CSoutput.t105 2.82907
R1785 CSoutput.n321 CSoutput.t85 2.82907
R1786 CSoutput.n320 CSoutput.t138 2.82907
R1787 CSoutput.n320 CSoutput.t119 2.82907
R1788 CSoutput.n318 CSoutput.t103 2.82907
R1789 CSoutput.n318 CSoutput.t120 2.82907
R1790 CSoutput.n316 CSoutput.t65 2.82907
R1791 CSoutput.n316 CSoutput.t99 2.82907
R1792 CSoutput.n314 CSoutput.t109 2.82907
R1793 CSoutput.n314 CSoutput.t128 2.82907
R1794 CSoutput.n312 CSoutput.t118 2.82907
R1795 CSoutput.n312 CSoutput.t79 2.82907
R1796 CSoutput.n310 CSoutput.t132 2.82907
R1797 CSoutput.n310 CSoutput.t136 2.82907
R1798 CSoutput.n308 CSoutput.t129 2.82907
R1799 CSoutput.n308 CSoutput.t64 2.82907
R1800 CSoutput.n306 CSoutput.t104 2.82907
R1801 CSoutput.n306 CSoutput.t123 2.82907
R1802 CSoutput.n304 CSoutput.t84 2.82907
R1803 CSoutput.n304 CSoutput.t93 2.82907
R1804 CSoutput.n302 CSoutput.t112 2.82907
R1805 CSoutput.n302 CSoutput.t114 2.82907
R1806 CSoutput.n301 CSoutput.t122 2.82907
R1807 CSoutput.n301 CSoutput.t82 2.82907
R1808 CSoutput.n360 CSoutput.t97 2.82907
R1809 CSoutput.n360 CSoutput.t70 2.82907
R1810 CSoutput.n361 CSoutput.t111 2.82907
R1811 CSoutput.n361 CSoutput.t90 2.82907
R1812 CSoutput.n363 CSoutput.t91 2.82907
R1813 CSoutput.n363 CSoutput.t63 2.82907
R1814 CSoutput.n365 CSoutput.t116 2.82907
R1815 CSoutput.n365 CSoutput.t94 2.82907
R1816 CSoutput.n367 CSoutput.t80 2.82907
R1817 CSoutput.n367 CSoutput.t124 2.82907
R1818 CSoutput.n369 CSoutput.t133 2.82907
R1819 CSoutput.n369 CSoutput.t98 2.82907
R1820 CSoutput.n371 CSoutput.t95 2.82907
R1821 CSoutput.n371 CSoutput.t67 2.82907
R1822 CSoutput.n373 CSoutput.t121 2.82907
R1823 CSoutput.n373 CSoutput.t140 2.82907
R1824 CSoutput.n375 CSoutput.t74 2.82907
R1825 CSoutput.n375 CSoutput.t81 2.82907
R1826 CSoutput.n377 CSoutput.t131 2.82907
R1827 CSoutput.n377 CSoutput.t86 2.82907
R1828 CSoutput.n341 CSoutput.t71 2.82907
R1829 CSoutput.n341 CSoutput.t77 2.82907
R1830 CSoutput.n342 CSoutput.t134 2.82907
R1831 CSoutput.n342 CSoutput.t100 2.82907
R1832 CSoutput.n344 CSoutput.t106 2.82907
R1833 CSoutput.n344 CSoutput.t92 2.82907
R1834 CSoutput.n346 CSoutput.t78 2.82907
R1835 CSoutput.n346 CSoutput.t88 2.82907
R1836 CSoutput.n348 CSoutput.t75 2.82907
R1837 CSoutput.n348 CSoutput.t83 2.82907
R1838 CSoutput.n350 CSoutput.t69 2.82907
R1839 CSoutput.n350 CSoutput.t141 2.82907
R1840 CSoutput.n352 CSoutput.t89 2.82907
R1841 CSoutput.n352 CSoutput.t96 2.82907
R1842 CSoutput.n354 CSoutput.t62 2.82907
R1843 CSoutput.n354 CSoutput.t125 2.82907
R1844 CSoutput.n356 CSoutput.t101 2.82907
R1845 CSoutput.n356 CSoutput.t76 2.82907
R1846 CSoutput.n358 CSoutput.t68 2.82907
R1847 CSoutput.n358 CSoutput.t115 2.82907
R1848 CSoutput.n75 CSoutput.n1 2.45513
R1849 CSoutput.n300 CSoutput.n114 2.36742
R1850 CSoutput.n205 CSoutput.n203 2.251
R1851 CSoutput.n205 CSoutput.n202 2.251
R1852 CSoutput.n205 CSoutput.n201 2.251
R1853 CSoutput.n205 CSoutput.n200 2.251
R1854 CSoutput.n174 CSoutput.n173 2.251
R1855 CSoutput.n174 CSoutput.n172 2.251
R1856 CSoutput.n174 CSoutput.n171 2.251
R1857 CSoutput.n174 CSoutput.n170 2.251
R1858 CSoutput.n247 CSoutput.n246 2.251
R1859 CSoutput.n212 CSoutput.n210 2.251
R1860 CSoutput.n212 CSoutput.n209 2.251
R1861 CSoutput.n212 CSoutput.n208 2.251
R1862 CSoutput.n230 CSoutput.n212 2.251
R1863 CSoutput.n218 CSoutput.n217 2.251
R1864 CSoutput.n218 CSoutput.n216 2.251
R1865 CSoutput.n218 CSoutput.n215 2.251
R1866 CSoutput.n218 CSoutput.n214 2.251
R1867 CSoutput.n244 CSoutput.n184 2.251
R1868 CSoutput.n239 CSoutput.n237 2.251
R1869 CSoutput.n239 CSoutput.n236 2.251
R1870 CSoutput.n239 CSoutput.n235 2.251
R1871 CSoutput.n239 CSoutput.n234 2.251
R1872 CSoutput.n140 CSoutput.n139 2.251
R1873 CSoutput.n140 CSoutput.n138 2.251
R1874 CSoutput.n140 CSoutput.n137 2.251
R1875 CSoutput.n140 CSoutput.n136 2.251
R1876 CSoutput.n257 CSoutput.n256 2.251
R1877 CSoutput.n174 CSoutput.n154 2.2505
R1878 CSoutput.n169 CSoutput.n154 2.2505
R1879 CSoutput.n167 CSoutput.n154 2.2505
R1880 CSoutput.n166 CSoutput.n154 2.2505
R1881 CSoutput.n251 CSoutput.n154 2.2505
R1882 CSoutput.n249 CSoutput.n154 2.2505
R1883 CSoutput.n247 CSoutput.n154 2.2505
R1884 CSoutput.n177 CSoutput.n154 2.2505
R1885 CSoutput.n176 CSoutput.n154 2.2505
R1886 CSoutput.n180 CSoutput.n154 2.2505
R1887 CSoutput.n179 CSoutput.n154 2.2505
R1888 CSoutput.n162 CSoutput.n154 2.2505
R1889 CSoutput.n254 CSoutput.n154 2.2505
R1890 CSoutput.n254 CSoutput.n253 2.2505
R1891 CSoutput.n218 CSoutput.n189 2.2505
R1892 CSoutput.n199 CSoutput.n189 2.2505
R1893 CSoutput.n220 CSoutput.n189 2.2505
R1894 CSoutput.n198 CSoutput.n189 2.2505
R1895 CSoutput.n222 CSoutput.n189 2.2505
R1896 CSoutput.n189 CSoutput.n183 2.2505
R1897 CSoutput.n244 CSoutput.n189 2.2505
R1898 CSoutput.n242 CSoutput.n189 2.2505
R1899 CSoutput.n224 CSoutput.n189 2.2505
R1900 CSoutput.n196 CSoutput.n189 2.2505
R1901 CSoutput.n226 CSoutput.n189 2.2505
R1902 CSoutput.n195 CSoutput.n189 2.2505
R1903 CSoutput.n240 CSoutput.n189 2.2505
R1904 CSoutput.n240 CSoutput.n193 2.2505
R1905 CSoutput.n140 CSoutput.n120 2.2505
R1906 CSoutput.n135 CSoutput.n120 2.2505
R1907 CSoutput.n133 CSoutput.n120 2.2505
R1908 CSoutput.n132 CSoutput.n120 2.2505
R1909 CSoutput.n261 CSoutput.n120 2.2505
R1910 CSoutput.n259 CSoutput.n120 2.2505
R1911 CSoutput.n257 CSoutput.n120 2.2505
R1912 CSoutput.n143 CSoutput.n120 2.2505
R1913 CSoutput.n142 CSoutput.n120 2.2505
R1914 CSoutput.n146 CSoutput.n120 2.2505
R1915 CSoutput.n145 CSoutput.n120 2.2505
R1916 CSoutput.n128 CSoutput.n120 2.2505
R1917 CSoutput.n264 CSoutput.n120 2.2505
R1918 CSoutput.n264 CSoutput.n263 2.2505
R1919 CSoutput.n182 CSoutput.n175 2.25024
R1920 CSoutput.n182 CSoutput.n168 2.25024
R1921 CSoutput.n250 CSoutput.n182 2.25024
R1922 CSoutput.n182 CSoutput.n178 2.25024
R1923 CSoutput.n182 CSoutput.n181 2.25024
R1924 CSoutput.n182 CSoutput.n149 2.25024
R1925 CSoutput.n232 CSoutput.n229 2.25024
R1926 CSoutput.n232 CSoutput.n228 2.25024
R1927 CSoutput.n232 CSoutput.n227 2.25024
R1928 CSoutput.n232 CSoutput.n194 2.25024
R1929 CSoutput.n232 CSoutput.n231 2.25024
R1930 CSoutput.n233 CSoutput.n232 2.25024
R1931 CSoutput.n148 CSoutput.n141 2.25024
R1932 CSoutput.n148 CSoutput.n134 2.25024
R1933 CSoutput.n260 CSoutput.n148 2.25024
R1934 CSoutput.n148 CSoutput.n144 2.25024
R1935 CSoutput.n148 CSoutput.n147 2.25024
R1936 CSoutput.n148 CSoutput.n115 2.25024
R1937 CSoutput.n249 CSoutput.n159 1.50111
R1938 CSoutput.n197 CSoutput.n183 1.50111
R1939 CSoutput.n259 CSoutput.n125 1.50111
R1940 CSoutput.n205 CSoutput.n204 1.501
R1941 CSoutput.n212 CSoutput.n211 1.501
R1942 CSoutput.n239 CSoutput.n238 1.501
R1943 CSoutput.n253 CSoutput.n164 1.12536
R1944 CSoutput.n253 CSoutput.n165 1.12536
R1945 CSoutput.n253 CSoutput.n252 1.12536
R1946 CSoutput.n213 CSoutput.n193 1.12536
R1947 CSoutput.n219 CSoutput.n193 1.12536
R1948 CSoutput.n221 CSoutput.n193 1.12536
R1949 CSoutput.n263 CSoutput.n130 1.12536
R1950 CSoutput.n263 CSoutput.n131 1.12536
R1951 CSoutput.n263 CSoutput.n262 1.12536
R1952 CSoutput.n253 CSoutput.n160 1.12536
R1953 CSoutput.n253 CSoutput.n161 1.12536
R1954 CSoutput.n253 CSoutput.n163 1.12536
R1955 CSoutput.n243 CSoutput.n193 1.12536
R1956 CSoutput.n223 CSoutput.n193 1.12536
R1957 CSoutput.n225 CSoutput.n193 1.12536
R1958 CSoutput.n263 CSoutput.n126 1.12536
R1959 CSoutput.n263 CSoutput.n127 1.12536
R1960 CSoutput.n263 CSoutput.n129 1.12536
R1961 CSoutput.n31 CSoutput.n30 0.669944
R1962 CSoutput.n62 CSoutput.n61 0.669944
R1963 CSoutput.n324 CSoutput.n322 0.573776
R1964 CSoutput.n326 CSoutput.n324 0.573776
R1965 CSoutput.n328 CSoutput.n326 0.573776
R1966 CSoutput.n330 CSoutput.n328 0.573776
R1967 CSoutput.n332 CSoutput.n330 0.573776
R1968 CSoutput.n334 CSoutput.n332 0.573776
R1969 CSoutput.n336 CSoutput.n334 0.573776
R1970 CSoutput.n338 CSoutput.n336 0.573776
R1971 CSoutput.n305 CSoutput.n303 0.573776
R1972 CSoutput.n307 CSoutput.n305 0.573776
R1973 CSoutput.n309 CSoutput.n307 0.573776
R1974 CSoutput.n311 CSoutput.n309 0.573776
R1975 CSoutput.n313 CSoutput.n311 0.573776
R1976 CSoutput.n315 CSoutput.n313 0.573776
R1977 CSoutput.n317 CSoutput.n315 0.573776
R1978 CSoutput.n319 CSoutput.n317 0.573776
R1979 CSoutput.n378 CSoutput.n376 0.573776
R1980 CSoutput.n376 CSoutput.n374 0.573776
R1981 CSoutput.n374 CSoutput.n372 0.573776
R1982 CSoutput.n372 CSoutput.n370 0.573776
R1983 CSoutput.n370 CSoutput.n368 0.573776
R1984 CSoutput.n368 CSoutput.n366 0.573776
R1985 CSoutput.n366 CSoutput.n364 0.573776
R1986 CSoutput.n364 CSoutput.n362 0.573776
R1987 CSoutput.n359 CSoutput.n357 0.573776
R1988 CSoutput.n357 CSoutput.n355 0.573776
R1989 CSoutput.n355 CSoutput.n353 0.573776
R1990 CSoutput.n353 CSoutput.n351 0.573776
R1991 CSoutput.n351 CSoutput.n349 0.573776
R1992 CSoutput.n349 CSoutput.n347 0.573776
R1993 CSoutput.n347 CSoutput.n345 0.573776
R1994 CSoutput.n345 CSoutput.n343 0.573776
R1995 CSoutput.n381 CSoutput.n264 0.53442
R1996 CSoutput.n292 CSoutput.n290 0.358259
R1997 CSoutput.n294 CSoutput.n292 0.358259
R1998 CSoutput.n296 CSoutput.n294 0.358259
R1999 CSoutput.n298 CSoutput.n296 0.358259
R2000 CSoutput.n280 CSoutput.n278 0.358259
R2001 CSoutput.n282 CSoutput.n280 0.358259
R2002 CSoutput.n284 CSoutput.n282 0.358259
R2003 CSoutput.n286 CSoutput.n284 0.358259
R2004 CSoutput.n269 CSoutput.n267 0.358259
R2005 CSoutput.n271 CSoutput.n269 0.358259
R2006 CSoutput.n273 CSoutput.n271 0.358259
R2007 CSoutput.n275 CSoutput.n273 0.358259
R2008 CSoutput.n112 CSoutput.n110 0.358259
R2009 CSoutput.n110 CSoutput.n108 0.358259
R2010 CSoutput.n108 CSoutput.n106 0.358259
R2011 CSoutput.n106 CSoutput.n104 0.358259
R2012 CSoutput.n100 CSoutput.n98 0.358259
R2013 CSoutput.n98 CSoutput.n96 0.358259
R2014 CSoutput.n96 CSoutput.n94 0.358259
R2015 CSoutput.n94 CSoutput.n92 0.358259
R2016 CSoutput.n89 CSoutput.n87 0.358259
R2017 CSoutput.n87 CSoutput.n85 0.358259
R2018 CSoutput.n85 CSoutput.n83 0.358259
R2019 CSoutput.n83 CSoutput.n81 0.358259
R2020 CSoutput.n21 CSoutput.n20 0.169105
R2021 CSoutput.n21 CSoutput.n16 0.169105
R2022 CSoutput.n26 CSoutput.n16 0.169105
R2023 CSoutput.n27 CSoutput.n26 0.169105
R2024 CSoutput.n27 CSoutput.n14 0.169105
R2025 CSoutput.n32 CSoutput.n14 0.169105
R2026 CSoutput.n33 CSoutput.n32 0.169105
R2027 CSoutput.n34 CSoutput.n33 0.169105
R2028 CSoutput.n34 CSoutput.n12 0.169105
R2029 CSoutput.n39 CSoutput.n12 0.169105
R2030 CSoutput.n40 CSoutput.n39 0.169105
R2031 CSoutput.n40 CSoutput.n10 0.169105
R2032 CSoutput.n45 CSoutput.n10 0.169105
R2033 CSoutput.n46 CSoutput.n45 0.169105
R2034 CSoutput.n47 CSoutput.n46 0.169105
R2035 CSoutput.n47 CSoutput.n8 0.169105
R2036 CSoutput.n52 CSoutput.n8 0.169105
R2037 CSoutput.n53 CSoutput.n52 0.169105
R2038 CSoutput.n53 CSoutput.n6 0.169105
R2039 CSoutput.n58 CSoutput.n6 0.169105
R2040 CSoutput.n59 CSoutput.n58 0.169105
R2041 CSoutput.n60 CSoutput.n59 0.169105
R2042 CSoutput.n60 CSoutput.n4 0.169105
R2043 CSoutput.n66 CSoutput.n4 0.169105
R2044 CSoutput.n67 CSoutput.n66 0.169105
R2045 CSoutput.n68 CSoutput.n67 0.169105
R2046 CSoutput.n68 CSoutput.n2 0.169105
R2047 CSoutput.n73 CSoutput.n2 0.169105
R2048 CSoutput.n74 CSoutput.n73 0.169105
R2049 CSoutput.n74 CSoutput.n0 0.169105
R2050 CSoutput.n78 CSoutput.n0 0.169105
R2051 CSoutput.n207 CSoutput.n206 0.0910737
R2052 CSoutput.n258 CSoutput.n255 0.0723685
R2053 CSoutput.n212 CSoutput.n207 0.0522944
R2054 CSoutput.n255 CSoutput.n254 0.0499135
R2055 CSoutput.n206 CSoutput.n205 0.0499135
R2056 CSoutput.n240 CSoutput.n239 0.0464294
R2057 CSoutput.n248 CSoutput.n245 0.0391444
R2058 CSoutput.n207 CSoutput.t152 0.023435
R2059 CSoutput.n255 CSoutput.t156 0.02262
R2060 CSoutput.n206 CSoutput.t159 0.02262
R2061 CSoutput CSoutput.n381 0.0052
R2062 CSoutput.n177 CSoutput.n160 0.00365111
R2063 CSoutput.n180 CSoutput.n161 0.00365111
R2064 CSoutput.n163 CSoutput.n162 0.00365111
R2065 CSoutput.n205 CSoutput.n164 0.00365111
R2066 CSoutput.n169 CSoutput.n165 0.00365111
R2067 CSoutput.n252 CSoutput.n166 0.00365111
R2068 CSoutput.n243 CSoutput.n242 0.00365111
R2069 CSoutput.n223 CSoutput.n196 0.00365111
R2070 CSoutput.n225 CSoutput.n195 0.00365111
R2071 CSoutput.n213 CSoutput.n212 0.00365111
R2072 CSoutput.n219 CSoutput.n199 0.00365111
R2073 CSoutput.n221 CSoutput.n198 0.00365111
R2074 CSoutput.n143 CSoutput.n126 0.00365111
R2075 CSoutput.n146 CSoutput.n127 0.00365111
R2076 CSoutput.n129 CSoutput.n128 0.00365111
R2077 CSoutput.n239 CSoutput.n130 0.00365111
R2078 CSoutput.n135 CSoutput.n131 0.00365111
R2079 CSoutput.n262 CSoutput.n132 0.00365111
R2080 CSoutput.n174 CSoutput.n164 0.00340054
R2081 CSoutput.n167 CSoutput.n165 0.00340054
R2082 CSoutput.n252 CSoutput.n251 0.00340054
R2083 CSoutput.n247 CSoutput.n160 0.00340054
R2084 CSoutput.n176 CSoutput.n161 0.00340054
R2085 CSoutput.n179 CSoutput.n163 0.00340054
R2086 CSoutput.n218 CSoutput.n213 0.00340054
R2087 CSoutput.n220 CSoutput.n219 0.00340054
R2088 CSoutput.n222 CSoutput.n221 0.00340054
R2089 CSoutput.n244 CSoutput.n243 0.00340054
R2090 CSoutput.n224 CSoutput.n223 0.00340054
R2091 CSoutput.n226 CSoutput.n225 0.00340054
R2092 CSoutput.n140 CSoutput.n130 0.00340054
R2093 CSoutput.n133 CSoutput.n131 0.00340054
R2094 CSoutput.n262 CSoutput.n261 0.00340054
R2095 CSoutput.n257 CSoutput.n126 0.00340054
R2096 CSoutput.n142 CSoutput.n127 0.00340054
R2097 CSoutput.n145 CSoutput.n129 0.00340054
R2098 CSoutput.n175 CSoutput.n169 0.00252698
R2099 CSoutput.n168 CSoutput.n166 0.00252698
R2100 CSoutput.n250 CSoutput.n249 0.00252698
R2101 CSoutput.n178 CSoutput.n176 0.00252698
R2102 CSoutput.n181 CSoutput.n179 0.00252698
R2103 CSoutput.n254 CSoutput.n149 0.00252698
R2104 CSoutput.n175 CSoutput.n174 0.00252698
R2105 CSoutput.n168 CSoutput.n167 0.00252698
R2106 CSoutput.n251 CSoutput.n250 0.00252698
R2107 CSoutput.n178 CSoutput.n177 0.00252698
R2108 CSoutput.n181 CSoutput.n180 0.00252698
R2109 CSoutput.n162 CSoutput.n149 0.00252698
R2110 CSoutput.n229 CSoutput.n199 0.00252698
R2111 CSoutput.n228 CSoutput.n198 0.00252698
R2112 CSoutput.n227 CSoutput.n183 0.00252698
R2113 CSoutput.n224 CSoutput.n194 0.00252698
R2114 CSoutput.n231 CSoutput.n226 0.00252698
R2115 CSoutput.n240 CSoutput.n233 0.00252698
R2116 CSoutput.n229 CSoutput.n218 0.00252698
R2117 CSoutput.n228 CSoutput.n220 0.00252698
R2118 CSoutput.n227 CSoutput.n222 0.00252698
R2119 CSoutput.n242 CSoutput.n194 0.00252698
R2120 CSoutput.n231 CSoutput.n196 0.00252698
R2121 CSoutput.n233 CSoutput.n195 0.00252698
R2122 CSoutput.n141 CSoutput.n135 0.00252698
R2123 CSoutput.n134 CSoutput.n132 0.00252698
R2124 CSoutput.n260 CSoutput.n259 0.00252698
R2125 CSoutput.n144 CSoutput.n142 0.00252698
R2126 CSoutput.n147 CSoutput.n145 0.00252698
R2127 CSoutput.n264 CSoutput.n115 0.00252698
R2128 CSoutput.n141 CSoutput.n140 0.00252698
R2129 CSoutput.n134 CSoutput.n133 0.00252698
R2130 CSoutput.n261 CSoutput.n260 0.00252698
R2131 CSoutput.n144 CSoutput.n143 0.00252698
R2132 CSoutput.n147 CSoutput.n146 0.00252698
R2133 CSoutput.n128 CSoutput.n115 0.00252698
R2134 CSoutput.n249 CSoutput.n248 0.0020275
R2135 CSoutput.n248 CSoutput.n247 0.0020275
R2136 CSoutput.n245 CSoutput.n183 0.0020275
R2137 CSoutput.n245 CSoutput.n244 0.0020275
R2138 CSoutput.n259 CSoutput.n258 0.0020275
R2139 CSoutput.n258 CSoutput.n257 0.0020275
R2140 CSoutput.n159 CSoutput.n158 0.00166668
R2141 CSoutput.n241 CSoutput.n197 0.00166668
R2142 CSoutput.n125 CSoutput.n124 0.00166668
R2143 CSoutput.n263 CSoutput.n125 0.00133328
R2144 CSoutput.n197 CSoutput.n193 0.00133328
R2145 CSoutput.n253 CSoutput.n159 0.00133328
R2146 CSoutput.n256 CSoutput.n148 0.001
R2147 CSoutput.n234 CSoutput.n148 0.001
R2148 CSoutput.n136 CSoutput.n116 0.001
R2149 CSoutput.n235 CSoutput.n116 0.001
R2150 CSoutput.n137 CSoutput.n117 0.001
R2151 CSoutput.n236 CSoutput.n117 0.001
R2152 CSoutput.n138 CSoutput.n118 0.001
R2153 CSoutput.n237 CSoutput.n118 0.001
R2154 CSoutput.n139 CSoutput.n119 0.001
R2155 CSoutput.n238 CSoutput.n119 0.001
R2156 CSoutput.n232 CSoutput.n184 0.001
R2157 CSoutput.n232 CSoutput.n230 0.001
R2158 CSoutput.n214 CSoutput.n185 0.001
R2159 CSoutput.n208 CSoutput.n185 0.001
R2160 CSoutput.n215 CSoutput.n186 0.001
R2161 CSoutput.n209 CSoutput.n186 0.001
R2162 CSoutput.n216 CSoutput.n187 0.001
R2163 CSoutput.n210 CSoutput.n187 0.001
R2164 CSoutput.n217 CSoutput.n188 0.001
R2165 CSoutput.n211 CSoutput.n188 0.001
R2166 CSoutput.n246 CSoutput.n182 0.001
R2167 CSoutput.n200 CSoutput.n182 0.001
R2168 CSoutput.n170 CSoutput.n150 0.001
R2169 CSoutput.n201 CSoutput.n150 0.001
R2170 CSoutput.n171 CSoutput.n151 0.001
R2171 CSoutput.n202 CSoutput.n151 0.001
R2172 CSoutput.n172 CSoutput.n152 0.001
R2173 CSoutput.n203 CSoutput.n152 0.001
R2174 CSoutput.n173 CSoutput.n153 0.001
R2175 CSoutput.n204 CSoutput.n153 0.001
R2176 CSoutput.n204 CSoutput.n154 0.001
R2177 CSoutput.n203 CSoutput.n155 0.001
R2178 CSoutput.n202 CSoutput.n156 0.001
R2179 CSoutput.n201 CSoutput.t172 0.001
R2180 CSoutput.n200 CSoutput.n157 0.001
R2181 CSoutput.n173 CSoutput.n155 0.001
R2182 CSoutput.n172 CSoutput.n156 0.001
R2183 CSoutput.n171 CSoutput.t172 0.001
R2184 CSoutput.n170 CSoutput.n157 0.001
R2185 CSoutput.n246 CSoutput.n158 0.001
R2186 CSoutput.n211 CSoutput.n189 0.001
R2187 CSoutput.n210 CSoutput.n190 0.001
R2188 CSoutput.n209 CSoutput.n191 0.001
R2189 CSoutput.n208 CSoutput.t166 0.001
R2190 CSoutput.n230 CSoutput.n192 0.001
R2191 CSoutput.n217 CSoutput.n190 0.001
R2192 CSoutput.n216 CSoutput.n191 0.001
R2193 CSoutput.n215 CSoutput.t166 0.001
R2194 CSoutput.n214 CSoutput.n192 0.001
R2195 CSoutput.n241 CSoutput.n184 0.001
R2196 CSoutput.n238 CSoutput.n120 0.001
R2197 CSoutput.n237 CSoutput.n121 0.001
R2198 CSoutput.n236 CSoutput.n122 0.001
R2199 CSoutput.n235 CSoutput.t163 0.001
R2200 CSoutput.n234 CSoutput.n123 0.001
R2201 CSoutput.n139 CSoutput.n121 0.001
R2202 CSoutput.n138 CSoutput.n122 0.001
R2203 CSoutput.n137 CSoutput.t163 0.001
R2204 CSoutput.n136 CSoutput.n123 0.001
R2205 CSoutput.n256 CSoutput.n124 0.001
R2206 gnd.n2829 gnd.n2828 978.75
R2207 gnd.n4756 gnd.n4755 939.716
R2208 gnd.n5581 gnd.n1311 771.183
R2209 gnd.n6759 gnd.n6758 771.183
R2210 gnd.n5818 gnd.n1309 771.183
R2211 gnd.n6815 gnd.n632 771.183
R2212 gnd.n4663 gnd.n1989 766.379
R2213 gnd.n4666 gnd.n4665 766.379
R2214 gnd.n3968 gnd.n3871 766.379
R2215 gnd.n3964 gnd.n3869 766.379
R2216 gnd.n4754 gnd.n2011 756.769
R2217 gnd.n3363 gnd.n3362 756.769
R2218 gnd.n4061 gnd.n3778 756.769
R2219 gnd.n4059 gnd.n3781 756.769
R2220 gnd.n7417 gnd.n125 751.963
R2221 gnd.n7575 gnd.n7574 751.963
R2222 gnd.n6973 gnd.n517 751.963
R2223 gnd.n6621 gnd.n479 751.963
R2224 gnd.n5575 gnd.n1357 751.963
R2225 gnd.n5773 gnd.n5772 751.963
R2226 gnd.n4823 gnd.n4758 751.963
R2227 gnd.n5071 gnd.n1987 751.963
R2228 gnd.n7572 gnd.n127 732.745
R2229 gnd.n195 gnd.n123 732.745
R2230 gnd.n6976 gnd.n6975 732.745
R2231 gnd.n7048 gnd.n484 732.745
R2232 gnd.n5770 gnd.n1359 732.745
R2233 gnd.n5701 gnd.n1355 732.745
R2234 gnd.n4990 gnd.n4757 732.745
R2235 gnd.n5069 gnd.n4873 732.745
R2236 gnd.n3140 gnd.n2188 723.135
R2237 gnd.n2830 gnd.n2496 723.135
R2238 gnd.n7220 gnd.n343 723.135
R2239 gnd.n2064 gnd.n1798 723.135
R2240 gnd.n2188 gnd.n2187 585
R2241 gnd.n3142 gnd.n2188 585
R2242 gnd.n3145 gnd.n3144 585
R2243 gnd.n3144 gnd.n3143 585
R2244 gnd.n2185 gnd.n2184 585
R2245 gnd.n2184 gnd.n2183 585
R2246 gnd.n3150 gnd.n3149 585
R2247 gnd.n3151 gnd.n3150 585
R2248 gnd.n2182 gnd.n2181 585
R2249 gnd.n3152 gnd.n2182 585
R2250 gnd.n3155 gnd.n3154 585
R2251 gnd.n3154 gnd.n3153 585
R2252 gnd.n2179 gnd.n2178 585
R2253 gnd.n2178 gnd.n2177 585
R2254 gnd.n3160 gnd.n3159 585
R2255 gnd.n3161 gnd.n3160 585
R2256 gnd.n2176 gnd.n2175 585
R2257 gnd.n3162 gnd.n2176 585
R2258 gnd.n3165 gnd.n3164 585
R2259 gnd.n3164 gnd.n3163 585
R2260 gnd.n2173 gnd.n2172 585
R2261 gnd.n2172 gnd.n2171 585
R2262 gnd.n3170 gnd.n3169 585
R2263 gnd.n3171 gnd.n3170 585
R2264 gnd.n2170 gnd.n2169 585
R2265 gnd.n3172 gnd.n2170 585
R2266 gnd.n3175 gnd.n3174 585
R2267 gnd.n3174 gnd.n3173 585
R2268 gnd.n2167 gnd.n2166 585
R2269 gnd.n2166 gnd.n2165 585
R2270 gnd.n3180 gnd.n3179 585
R2271 gnd.n3181 gnd.n3180 585
R2272 gnd.n2164 gnd.n2163 585
R2273 gnd.n3182 gnd.n2164 585
R2274 gnd.n3185 gnd.n3184 585
R2275 gnd.n3184 gnd.n3183 585
R2276 gnd.n2161 gnd.n2160 585
R2277 gnd.n2160 gnd.n2159 585
R2278 gnd.n3190 gnd.n3189 585
R2279 gnd.n3191 gnd.n3190 585
R2280 gnd.n2158 gnd.n2157 585
R2281 gnd.n3192 gnd.n2158 585
R2282 gnd.n3195 gnd.n3194 585
R2283 gnd.n3194 gnd.n3193 585
R2284 gnd.n2155 gnd.n2154 585
R2285 gnd.n2154 gnd.n2153 585
R2286 gnd.n3200 gnd.n3199 585
R2287 gnd.n3201 gnd.n3200 585
R2288 gnd.n2152 gnd.n2151 585
R2289 gnd.n3202 gnd.n2152 585
R2290 gnd.n3205 gnd.n3204 585
R2291 gnd.n3204 gnd.n3203 585
R2292 gnd.n2149 gnd.n2148 585
R2293 gnd.n2148 gnd.n2147 585
R2294 gnd.n3210 gnd.n3209 585
R2295 gnd.n3211 gnd.n3210 585
R2296 gnd.n2146 gnd.n2145 585
R2297 gnd.n3212 gnd.n2146 585
R2298 gnd.n3215 gnd.n3214 585
R2299 gnd.n3214 gnd.n3213 585
R2300 gnd.n2143 gnd.n2142 585
R2301 gnd.n2142 gnd.n2141 585
R2302 gnd.n3220 gnd.n3219 585
R2303 gnd.n3221 gnd.n3220 585
R2304 gnd.n2140 gnd.n2139 585
R2305 gnd.n3222 gnd.n2140 585
R2306 gnd.n3225 gnd.n3224 585
R2307 gnd.n3224 gnd.n3223 585
R2308 gnd.n2137 gnd.n2136 585
R2309 gnd.n2136 gnd.n2135 585
R2310 gnd.n3230 gnd.n3229 585
R2311 gnd.n3231 gnd.n3230 585
R2312 gnd.n2134 gnd.n2133 585
R2313 gnd.n3232 gnd.n2134 585
R2314 gnd.n3235 gnd.n3234 585
R2315 gnd.n3234 gnd.n3233 585
R2316 gnd.n2131 gnd.n2130 585
R2317 gnd.n2130 gnd.n2129 585
R2318 gnd.n3240 gnd.n3239 585
R2319 gnd.n3241 gnd.n3240 585
R2320 gnd.n2128 gnd.n2127 585
R2321 gnd.n3242 gnd.n2128 585
R2322 gnd.n3245 gnd.n3244 585
R2323 gnd.n3244 gnd.n3243 585
R2324 gnd.n2125 gnd.n2124 585
R2325 gnd.n2124 gnd.n2123 585
R2326 gnd.n3250 gnd.n3249 585
R2327 gnd.n3251 gnd.n3250 585
R2328 gnd.n2122 gnd.n2121 585
R2329 gnd.n3252 gnd.n2122 585
R2330 gnd.n3255 gnd.n3254 585
R2331 gnd.n3254 gnd.n3253 585
R2332 gnd.n2119 gnd.n2118 585
R2333 gnd.n2118 gnd.n2117 585
R2334 gnd.n3260 gnd.n3259 585
R2335 gnd.n3261 gnd.n3260 585
R2336 gnd.n2116 gnd.n2115 585
R2337 gnd.n3262 gnd.n2116 585
R2338 gnd.n3265 gnd.n3264 585
R2339 gnd.n3264 gnd.n3263 585
R2340 gnd.n2113 gnd.n2112 585
R2341 gnd.n2112 gnd.n2111 585
R2342 gnd.n3270 gnd.n3269 585
R2343 gnd.n3271 gnd.n3270 585
R2344 gnd.n2110 gnd.n2109 585
R2345 gnd.n3272 gnd.n2110 585
R2346 gnd.n3275 gnd.n3274 585
R2347 gnd.n3274 gnd.n3273 585
R2348 gnd.n2107 gnd.n2106 585
R2349 gnd.n2106 gnd.n2105 585
R2350 gnd.n3280 gnd.n3279 585
R2351 gnd.n3281 gnd.n3280 585
R2352 gnd.n2104 gnd.n2103 585
R2353 gnd.n3282 gnd.n2104 585
R2354 gnd.n3285 gnd.n3284 585
R2355 gnd.n3284 gnd.n3283 585
R2356 gnd.n2101 gnd.n2100 585
R2357 gnd.n2100 gnd.n2099 585
R2358 gnd.n3290 gnd.n3289 585
R2359 gnd.n3291 gnd.n3290 585
R2360 gnd.n2098 gnd.n2097 585
R2361 gnd.n3292 gnd.n2098 585
R2362 gnd.n3295 gnd.n3294 585
R2363 gnd.n3294 gnd.n3293 585
R2364 gnd.n2095 gnd.n2094 585
R2365 gnd.n2094 gnd.n2093 585
R2366 gnd.n3300 gnd.n3299 585
R2367 gnd.n3301 gnd.n3300 585
R2368 gnd.n2092 gnd.n2091 585
R2369 gnd.n3302 gnd.n2092 585
R2370 gnd.n3305 gnd.n3304 585
R2371 gnd.n3304 gnd.n3303 585
R2372 gnd.n2089 gnd.n2088 585
R2373 gnd.n2088 gnd.n2087 585
R2374 gnd.n3310 gnd.n3309 585
R2375 gnd.n3311 gnd.n3310 585
R2376 gnd.n2086 gnd.n2085 585
R2377 gnd.n3312 gnd.n2086 585
R2378 gnd.n3315 gnd.n3314 585
R2379 gnd.n3314 gnd.n3313 585
R2380 gnd.n2083 gnd.n2082 585
R2381 gnd.n2082 gnd.n2081 585
R2382 gnd.n3320 gnd.n3319 585
R2383 gnd.n3321 gnd.n3320 585
R2384 gnd.n2080 gnd.n2079 585
R2385 gnd.n3322 gnd.n2080 585
R2386 gnd.n3325 gnd.n3324 585
R2387 gnd.n3324 gnd.n3323 585
R2388 gnd.n2077 gnd.n2076 585
R2389 gnd.n2076 gnd.n2075 585
R2390 gnd.n3330 gnd.n3329 585
R2391 gnd.n3331 gnd.n3330 585
R2392 gnd.n2074 gnd.n2073 585
R2393 gnd.n3332 gnd.n2074 585
R2394 gnd.n3335 gnd.n3334 585
R2395 gnd.n3334 gnd.n3333 585
R2396 gnd.n2071 gnd.n2070 585
R2397 gnd.n2070 gnd.n2069 585
R2398 gnd.n3340 gnd.n3339 585
R2399 gnd.n3341 gnd.n3340 585
R2400 gnd.n2068 gnd.n2067 585
R2401 gnd.n3342 gnd.n2068 585
R2402 gnd.n3345 gnd.n3344 585
R2403 gnd.n3344 gnd.n3343 585
R2404 gnd.n2065 gnd.n2063 585
R2405 gnd.n2063 gnd.n2062 585
R2406 gnd.n3353 gnd.n3352 585
R2407 gnd.n3354 gnd.n3353 585
R2408 gnd.n3140 gnd.n3139 585
R2409 gnd.n3141 gnd.n3140 585
R2410 gnd.n2191 gnd.n2190 585
R2411 gnd.n2190 gnd.n2189 585
R2412 gnd.n3135 gnd.n3134 585
R2413 gnd.n3134 gnd.n3133 585
R2414 gnd.n2194 gnd.n2193 585
R2415 gnd.n3132 gnd.n2194 585
R2416 gnd.n3130 gnd.n3129 585
R2417 gnd.n3131 gnd.n3130 585
R2418 gnd.n3128 gnd.n2196 585
R2419 gnd.n2196 gnd.n2195 585
R2420 gnd.n3127 gnd.n3126 585
R2421 gnd.n3126 gnd.n3125 585
R2422 gnd.n2201 gnd.n2200 585
R2423 gnd.n3124 gnd.n2201 585
R2424 gnd.n3122 gnd.n3121 585
R2425 gnd.n3123 gnd.n3122 585
R2426 gnd.n3120 gnd.n2203 585
R2427 gnd.n2203 gnd.n2202 585
R2428 gnd.n3119 gnd.n3118 585
R2429 gnd.n3118 gnd.n3117 585
R2430 gnd.n2209 gnd.n2208 585
R2431 gnd.n3116 gnd.n2209 585
R2432 gnd.n3114 gnd.n3113 585
R2433 gnd.n3115 gnd.n3114 585
R2434 gnd.n3112 gnd.n2211 585
R2435 gnd.n2211 gnd.n2210 585
R2436 gnd.n3111 gnd.n3110 585
R2437 gnd.n3110 gnd.n3109 585
R2438 gnd.n2217 gnd.n2216 585
R2439 gnd.n3108 gnd.n2217 585
R2440 gnd.n3106 gnd.n3105 585
R2441 gnd.n3107 gnd.n3106 585
R2442 gnd.n3104 gnd.n2219 585
R2443 gnd.n2219 gnd.n2218 585
R2444 gnd.n3103 gnd.n3102 585
R2445 gnd.n3102 gnd.n3101 585
R2446 gnd.n2225 gnd.n2224 585
R2447 gnd.n3100 gnd.n2225 585
R2448 gnd.n3098 gnd.n3097 585
R2449 gnd.n3099 gnd.n3098 585
R2450 gnd.n3096 gnd.n2227 585
R2451 gnd.n2227 gnd.n2226 585
R2452 gnd.n3095 gnd.n3094 585
R2453 gnd.n3094 gnd.n3093 585
R2454 gnd.n2233 gnd.n2232 585
R2455 gnd.n3092 gnd.n2233 585
R2456 gnd.n3090 gnd.n3089 585
R2457 gnd.n3091 gnd.n3090 585
R2458 gnd.n3088 gnd.n2235 585
R2459 gnd.n2235 gnd.n2234 585
R2460 gnd.n3087 gnd.n3086 585
R2461 gnd.n3086 gnd.n3085 585
R2462 gnd.n2241 gnd.n2240 585
R2463 gnd.n3084 gnd.n2241 585
R2464 gnd.n3082 gnd.n3081 585
R2465 gnd.n3083 gnd.n3082 585
R2466 gnd.n3080 gnd.n2243 585
R2467 gnd.n2243 gnd.n2242 585
R2468 gnd.n3079 gnd.n3078 585
R2469 gnd.n3078 gnd.n3077 585
R2470 gnd.n2249 gnd.n2248 585
R2471 gnd.n3076 gnd.n2249 585
R2472 gnd.n3074 gnd.n3073 585
R2473 gnd.n3075 gnd.n3074 585
R2474 gnd.n3072 gnd.n2251 585
R2475 gnd.n2251 gnd.n2250 585
R2476 gnd.n3071 gnd.n3070 585
R2477 gnd.n3070 gnd.n3069 585
R2478 gnd.n2257 gnd.n2256 585
R2479 gnd.n3068 gnd.n2257 585
R2480 gnd.n3066 gnd.n3065 585
R2481 gnd.n3067 gnd.n3066 585
R2482 gnd.n3064 gnd.n2259 585
R2483 gnd.n2259 gnd.n2258 585
R2484 gnd.n3063 gnd.n3062 585
R2485 gnd.n3062 gnd.n3061 585
R2486 gnd.n2265 gnd.n2264 585
R2487 gnd.n3060 gnd.n2265 585
R2488 gnd.n3058 gnd.n3057 585
R2489 gnd.n3059 gnd.n3058 585
R2490 gnd.n3056 gnd.n2267 585
R2491 gnd.n2267 gnd.n2266 585
R2492 gnd.n3055 gnd.n3054 585
R2493 gnd.n3054 gnd.n3053 585
R2494 gnd.n2273 gnd.n2272 585
R2495 gnd.n3052 gnd.n2273 585
R2496 gnd.n3050 gnd.n3049 585
R2497 gnd.n3051 gnd.n3050 585
R2498 gnd.n3048 gnd.n2275 585
R2499 gnd.n2275 gnd.n2274 585
R2500 gnd.n3047 gnd.n3046 585
R2501 gnd.n3046 gnd.n3045 585
R2502 gnd.n2281 gnd.n2280 585
R2503 gnd.n3044 gnd.n2281 585
R2504 gnd.n3042 gnd.n3041 585
R2505 gnd.n3043 gnd.n3042 585
R2506 gnd.n3040 gnd.n2283 585
R2507 gnd.n2283 gnd.n2282 585
R2508 gnd.n3039 gnd.n3038 585
R2509 gnd.n3038 gnd.n3037 585
R2510 gnd.n2289 gnd.n2288 585
R2511 gnd.n3036 gnd.n2289 585
R2512 gnd.n3034 gnd.n3033 585
R2513 gnd.n3035 gnd.n3034 585
R2514 gnd.n3032 gnd.n2291 585
R2515 gnd.n2291 gnd.n2290 585
R2516 gnd.n3031 gnd.n3030 585
R2517 gnd.n3030 gnd.n3029 585
R2518 gnd.n2297 gnd.n2296 585
R2519 gnd.n3028 gnd.n2297 585
R2520 gnd.n3026 gnd.n3025 585
R2521 gnd.n3027 gnd.n3026 585
R2522 gnd.n3024 gnd.n2299 585
R2523 gnd.n2299 gnd.n2298 585
R2524 gnd.n3023 gnd.n3022 585
R2525 gnd.n3022 gnd.n3021 585
R2526 gnd.n2305 gnd.n2304 585
R2527 gnd.n3020 gnd.n2305 585
R2528 gnd.n3018 gnd.n3017 585
R2529 gnd.n3019 gnd.n3018 585
R2530 gnd.n3016 gnd.n2307 585
R2531 gnd.n2307 gnd.n2306 585
R2532 gnd.n3015 gnd.n3014 585
R2533 gnd.n3014 gnd.n3013 585
R2534 gnd.n2313 gnd.n2312 585
R2535 gnd.n3012 gnd.n2313 585
R2536 gnd.n3010 gnd.n3009 585
R2537 gnd.n3011 gnd.n3010 585
R2538 gnd.n3008 gnd.n2315 585
R2539 gnd.n2315 gnd.n2314 585
R2540 gnd.n3007 gnd.n3006 585
R2541 gnd.n3006 gnd.n3005 585
R2542 gnd.n2321 gnd.n2320 585
R2543 gnd.n3004 gnd.n2321 585
R2544 gnd.n3002 gnd.n3001 585
R2545 gnd.n3003 gnd.n3002 585
R2546 gnd.n3000 gnd.n2323 585
R2547 gnd.n2323 gnd.n2322 585
R2548 gnd.n2999 gnd.n2998 585
R2549 gnd.n2998 gnd.n2997 585
R2550 gnd.n2329 gnd.n2328 585
R2551 gnd.n2996 gnd.n2329 585
R2552 gnd.n2994 gnd.n2993 585
R2553 gnd.n2995 gnd.n2994 585
R2554 gnd.n2992 gnd.n2331 585
R2555 gnd.n2331 gnd.n2330 585
R2556 gnd.n2991 gnd.n2990 585
R2557 gnd.n2990 gnd.n2989 585
R2558 gnd.n2337 gnd.n2336 585
R2559 gnd.n2988 gnd.n2337 585
R2560 gnd.n2986 gnd.n2985 585
R2561 gnd.n2987 gnd.n2986 585
R2562 gnd.n2984 gnd.n2339 585
R2563 gnd.n2339 gnd.n2338 585
R2564 gnd.n2983 gnd.n2982 585
R2565 gnd.n2982 gnd.n2981 585
R2566 gnd.n2345 gnd.n2344 585
R2567 gnd.n2980 gnd.n2345 585
R2568 gnd.n2978 gnd.n2977 585
R2569 gnd.n2979 gnd.n2978 585
R2570 gnd.n2976 gnd.n2347 585
R2571 gnd.n2347 gnd.n2346 585
R2572 gnd.n2975 gnd.n2974 585
R2573 gnd.n2974 gnd.n2973 585
R2574 gnd.n2353 gnd.n2352 585
R2575 gnd.n2972 gnd.n2353 585
R2576 gnd.n2970 gnd.n2969 585
R2577 gnd.n2971 gnd.n2970 585
R2578 gnd.n2968 gnd.n2355 585
R2579 gnd.n2355 gnd.n2354 585
R2580 gnd.n2967 gnd.n2966 585
R2581 gnd.n2966 gnd.n2965 585
R2582 gnd.n2361 gnd.n2360 585
R2583 gnd.n2964 gnd.n2361 585
R2584 gnd.n2962 gnd.n2961 585
R2585 gnd.n2963 gnd.n2962 585
R2586 gnd.n2960 gnd.n2363 585
R2587 gnd.n2363 gnd.n2362 585
R2588 gnd.n2959 gnd.n2958 585
R2589 gnd.n2958 gnd.n2957 585
R2590 gnd.n2369 gnd.n2368 585
R2591 gnd.n2956 gnd.n2369 585
R2592 gnd.n2954 gnd.n2953 585
R2593 gnd.n2955 gnd.n2954 585
R2594 gnd.n2952 gnd.n2371 585
R2595 gnd.n2371 gnd.n2370 585
R2596 gnd.n2951 gnd.n2950 585
R2597 gnd.n2950 gnd.n2949 585
R2598 gnd.n2377 gnd.n2376 585
R2599 gnd.n2948 gnd.n2377 585
R2600 gnd.n2946 gnd.n2945 585
R2601 gnd.n2947 gnd.n2946 585
R2602 gnd.n2944 gnd.n2379 585
R2603 gnd.n2379 gnd.n2378 585
R2604 gnd.n2943 gnd.n2942 585
R2605 gnd.n2942 gnd.n2941 585
R2606 gnd.n2385 gnd.n2384 585
R2607 gnd.n2940 gnd.n2385 585
R2608 gnd.n2938 gnd.n2937 585
R2609 gnd.n2939 gnd.n2938 585
R2610 gnd.n2936 gnd.n2387 585
R2611 gnd.n2387 gnd.n2386 585
R2612 gnd.n2935 gnd.n2934 585
R2613 gnd.n2934 gnd.n2933 585
R2614 gnd.n2393 gnd.n2392 585
R2615 gnd.n2932 gnd.n2393 585
R2616 gnd.n2930 gnd.n2929 585
R2617 gnd.n2931 gnd.n2930 585
R2618 gnd.n2928 gnd.n2395 585
R2619 gnd.n2395 gnd.n2394 585
R2620 gnd.n2927 gnd.n2926 585
R2621 gnd.n2926 gnd.n2925 585
R2622 gnd.n2401 gnd.n2400 585
R2623 gnd.n2924 gnd.n2401 585
R2624 gnd.n2922 gnd.n2921 585
R2625 gnd.n2923 gnd.n2922 585
R2626 gnd.n2920 gnd.n2403 585
R2627 gnd.n2403 gnd.n2402 585
R2628 gnd.n2919 gnd.n2918 585
R2629 gnd.n2918 gnd.n2917 585
R2630 gnd.n2409 gnd.n2408 585
R2631 gnd.n2916 gnd.n2409 585
R2632 gnd.n2914 gnd.n2913 585
R2633 gnd.n2915 gnd.n2914 585
R2634 gnd.n2912 gnd.n2411 585
R2635 gnd.n2411 gnd.n2410 585
R2636 gnd.n2911 gnd.n2910 585
R2637 gnd.n2910 gnd.n2909 585
R2638 gnd.n2417 gnd.n2416 585
R2639 gnd.n2908 gnd.n2417 585
R2640 gnd.n2906 gnd.n2905 585
R2641 gnd.n2907 gnd.n2906 585
R2642 gnd.n2904 gnd.n2419 585
R2643 gnd.n2419 gnd.n2418 585
R2644 gnd.n2903 gnd.n2902 585
R2645 gnd.n2902 gnd.n2901 585
R2646 gnd.n2425 gnd.n2424 585
R2647 gnd.n2900 gnd.n2425 585
R2648 gnd.n2898 gnd.n2897 585
R2649 gnd.n2899 gnd.n2898 585
R2650 gnd.n2896 gnd.n2427 585
R2651 gnd.n2427 gnd.n2426 585
R2652 gnd.n2895 gnd.n2894 585
R2653 gnd.n2894 gnd.n2893 585
R2654 gnd.n2433 gnd.n2432 585
R2655 gnd.n2892 gnd.n2433 585
R2656 gnd.n2890 gnd.n2889 585
R2657 gnd.n2891 gnd.n2890 585
R2658 gnd.n2888 gnd.n2435 585
R2659 gnd.n2435 gnd.n2434 585
R2660 gnd.n2887 gnd.n2886 585
R2661 gnd.n2886 gnd.n2885 585
R2662 gnd.n2441 gnd.n2440 585
R2663 gnd.n2884 gnd.n2441 585
R2664 gnd.n2882 gnd.n2881 585
R2665 gnd.n2883 gnd.n2882 585
R2666 gnd.n2880 gnd.n2443 585
R2667 gnd.n2443 gnd.n2442 585
R2668 gnd.n2879 gnd.n2878 585
R2669 gnd.n2878 gnd.n2877 585
R2670 gnd.n2449 gnd.n2448 585
R2671 gnd.n2876 gnd.n2449 585
R2672 gnd.n2874 gnd.n2873 585
R2673 gnd.n2875 gnd.n2874 585
R2674 gnd.n2872 gnd.n2451 585
R2675 gnd.n2451 gnd.n2450 585
R2676 gnd.n2871 gnd.n2870 585
R2677 gnd.n2870 gnd.n2869 585
R2678 gnd.n2457 gnd.n2456 585
R2679 gnd.n2868 gnd.n2457 585
R2680 gnd.n2866 gnd.n2865 585
R2681 gnd.n2867 gnd.n2866 585
R2682 gnd.n2864 gnd.n2459 585
R2683 gnd.n2459 gnd.n2458 585
R2684 gnd.n2863 gnd.n2862 585
R2685 gnd.n2862 gnd.n2861 585
R2686 gnd.n2465 gnd.n2464 585
R2687 gnd.n2860 gnd.n2465 585
R2688 gnd.n2858 gnd.n2857 585
R2689 gnd.n2859 gnd.n2858 585
R2690 gnd.n2856 gnd.n2467 585
R2691 gnd.n2467 gnd.n2466 585
R2692 gnd.n2855 gnd.n2854 585
R2693 gnd.n2854 gnd.n2853 585
R2694 gnd.n2473 gnd.n2472 585
R2695 gnd.n2852 gnd.n2473 585
R2696 gnd.n2850 gnd.n2849 585
R2697 gnd.n2851 gnd.n2850 585
R2698 gnd.n2848 gnd.n2475 585
R2699 gnd.n2475 gnd.n2474 585
R2700 gnd.n2847 gnd.n2846 585
R2701 gnd.n2846 gnd.n2845 585
R2702 gnd.n2481 gnd.n2480 585
R2703 gnd.n2844 gnd.n2481 585
R2704 gnd.n2842 gnd.n2841 585
R2705 gnd.n2843 gnd.n2842 585
R2706 gnd.n2840 gnd.n2483 585
R2707 gnd.n2483 gnd.n2482 585
R2708 gnd.n2839 gnd.n2838 585
R2709 gnd.n2838 gnd.n2837 585
R2710 gnd.n2489 gnd.n2488 585
R2711 gnd.n2836 gnd.n2489 585
R2712 gnd.n2834 gnd.n2833 585
R2713 gnd.n2835 gnd.n2834 585
R2714 gnd.n2832 gnd.n2491 585
R2715 gnd.n2491 gnd.n2490 585
R2716 gnd.n2831 gnd.n2830 585
R2717 gnd.n2830 gnd.n2829 585
R2718 gnd.n344 gnd.n342 585
R2719 gnd.n2656 gnd.n342 585
R2720 gnd.n2662 gnd.n2658 585
R2721 gnd.n2658 gnd.n2657 585
R2722 gnd.n2664 gnd.n2663 585
R2723 gnd.n2665 gnd.n2664 585
R2724 gnd.n2655 gnd.n2654 585
R2725 gnd.n2666 gnd.n2655 585
R2726 gnd.n2669 gnd.n2668 585
R2727 gnd.n2668 gnd.n2667 585
R2728 gnd.n2670 gnd.n2649 585
R2729 gnd.n2649 gnd.n2648 585
R2730 gnd.n2672 gnd.n2671 585
R2731 gnd.n2673 gnd.n2672 585
R2732 gnd.n2647 gnd.n2646 585
R2733 gnd.n2674 gnd.n2647 585
R2734 gnd.n2677 gnd.n2676 585
R2735 gnd.n2676 gnd.n2675 585
R2736 gnd.n2678 gnd.n2641 585
R2737 gnd.n2641 gnd.n2640 585
R2738 gnd.n2680 gnd.n2679 585
R2739 gnd.n2681 gnd.n2680 585
R2740 gnd.n2639 gnd.n2638 585
R2741 gnd.n2682 gnd.n2639 585
R2742 gnd.n2685 gnd.n2684 585
R2743 gnd.n2684 gnd.n2683 585
R2744 gnd.n2686 gnd.n2633 585
R2745 gnd.n2633 gnd.n2632 585
R2746 gnd.n2688 gnd.n2687 585
R2747 gnd.n2689 gnd.n2688 585
R2748 gnd.n2631 gnd.n2630 585
R2749 gnd.n2690 gnd.n2631 585
R2750 gnd.n2693 gnd.n2692 585
R2751 gnd.n2692 gnd.n2691 585
R2752 gnd.n2694 gnd.n2625 585
R2753 gnd.n2625 gnd.n2624 585
R2754 gnd.n2696 gnd.n2695 585
R2755 gnd.n2697 gnd.n2696 585
R2756 gnd.n2623 gnd.n2622 585
R2757 gnd.n2698 gnd.n2623 585
R2758 gnd.n2701 gnd.n2700 585
R2759 gnd.n2700 gnd.n2699 585
R2760 gnd.n2702 gnd.n2617 585
R2761 gnd.n2617 gnd.n2616 585
R2762 gnd.n2704 gnd.n2703 585
R2763 gnd.n2705 gnd.n2704 585
R2764 gnd.n2615 gnd.n2614 585
R2765 gnd.n2706 gnd.n2615 585
R2766 gnd.n2709 gnd.n2708 585
R2767 gnd.n2708 gnd.n2707 585
R2768 gnd.n2710 gnd.n2609 585
R2769 gnd.n2609 gnd.n2608 585
R2770 gnd.n2712 gnd.n2711 585
R2771 gnd.n2713 gnd.n2712 585
R2772 gnd.n2607 gnd.n2606 585
R2773 gnd.n2714 gnd.n2607 585
R2774 gnd.n2717 gnd.n2716 585
R2775 gnd.n2716 gnd.n2715 585
R2776 gnd.n2718 gnd.n2601 585
R2777 gnd.n2601 gnd.n2600 585
R2778 gnd.n2720 gnd.n2719 585
R2779 gnd.n2721 gnd.n2720 585
R2780 gnd.n2599 gnd.n2598 585
R2781 gnd.n2722 gnd.n2599 585
R2782 gnd.n2725 gnd.n2724 585
R2783 gnd.n2724 gnd.n2723 585
R2784 gnd.n2726 gnd.n2593 585
R2785 gnd.n2593 gnd.n2592 585
R2786 gnd.n2728 gnd.n2727 585
R2787 gnd.n2729 gnd.n2728 585
R2788 gnd.n2591 gnd.n2590 585
R2789 gnd.n2730 gnd.n2591 585
R2790 gnd.n2733 gnd.n2732 585
R2791 gnd.n2732 gnd.n2731 585
R2792 gnd.n2734 gnd.n2585 585
R2793 gnd.n2585 gnd.n2584 585
R2794 gnd.n2736 gnd.n2735 585
R2795 gnd.n2737 gnd.n2736 585
R2796 gnd.n2583 gnd.n2582 585
R2797 gnd.n2738 gnd.n2583 585
R2798 gnd.n2741 gnd.n2740 585
R2799 gnd.n2740 gnd.n2739 585
R2800 gnd.n2742 gnd.n2577 585
R2801 gnd.n2577 gnd.n2576 585
R2802 gnd.n2744 gnd.n2743 585
R2803 gnd.n2745 gnd.n2744 585
R2804 gnd.n2575 gnd.n2574 585
R2805 gnd.n2746 gnd.n2575 585
R2806 gnd.n2749 gnd.n2748 585
R2807 gnd.n2748 gnd.n2747 585
R2808 gnd.n2750 gnd.n2569 585
R2809 gnd.n2569 gnd.n2568 585
R2810 gnd.n2752 gnd.n2751 585
R2811 gnd.n2753 gnd.n2752 585
R2812 gnd.n2567 gnd.n2566 585
R2813 gnd.n2754 gnd.n2567 585
R2814 gnd.n2757 gnd.n2756 585
R2815 gnd.n2756 gnd.n2755 585
R2816 gnd.n2758 gnd.n2561 585
R2817 gnd.n2561 gnd.n2560 585
R2818 gnd.n2760 gnd.n2759 585
R2819 gnd.n2761 gnd.n2760 585
R2820 gnd.n2559 gnd.n2558 585
R2821 gnd.n2762 gnd.n2559 585
R2822 gnd.n2765 gnd.n2764 585
R2823 gnd.n2764 gnd.n2763 585
R2824 gnd.n2766 gnd.n2553 585
R2825 gnd.n2553 gnd.n2552 585
R2826 gnd.n2768 gnd.n2767 585
R2827 gnd.n2769 gnd.n2768 585
R2828 gnd.n2551 gnd.n2550 585
R2829 gnd.n2770 gnd.n2551 585
R2830 gnd.n2773 gnd.n2772 585
R2831 gnd.n2772 gnd.n2771 585
R2832 gnd.n2774 gnd.n2545 585
R2833 gnd.n2545 gnd.n2544 585
R2834 gnd.n2776 gnd.n2775 585
R2835 gnd.n2777 gnd.n2776 585
R2836 gnd.n2543 gnd.n2542 585
R2837 gnd.n2778 gnd.n2543 585
R2838 gnd.n2781 gnd.n2780 585
R2839 gnd.n2780 gnd.n2779 585
R2840 gnd.n2782 gnd.n2537 585
R2841 gnd.n2537 gnd.n2536 585
R2842 gnd.n2784 gnd.n2783 585
R2843 gnd.n2785 gnd.n2784 585
R2844 gnd.n2535 gnd.n2534 585
R2845 gnd.n2786 gnd.n2535 585
R2846 gnd.n2789 gnd.n2788 585
R2847 gnd.n2788 gnd.n2787 585
R2848 gnd.n2790 gnd.n2529 585
R2849 gnd.n2529 gnd.n2528 585
R2850 gnd.n2792 gnd.n2791 585
R2851 gnd.n2793 gnd.n2792 585
R2852 gnd.n2527 gnd.n2526 585
R2853 gnd.n2794 gnd.n2527 585
R2854 gnd.n2797 gnd.n2796 585
R2855 gnd.n2796 gnd.n2795 585
R2856 gnd.n2798 gnd.n2521 585
R2857 gnd.n2521 gnd.n2520 585
R2858 gnd.n2800 gnd.n2799 585
R2859 gnd.n2801 gnd.n2800 585
R2860 gnd.n2519 gnd.n2518 585
R2861 gnd.n2802 gnd.n2519 585
R2862 gnd.n2805 gnd.n2804 585
R2863 gnd.n2804 gnd.n2803 585
R2864 gnd.n2806 gnd.n2513 585
R2865 gnd.n2513 gnd.n2512 585
R2866 gnd.n2808 gnd.n2807 585
R2867 gnd.n2809 gnd.n2808 585
R2868 gnd.n2511 gnd.n2510 585
R2869 gnd.n2810 gnd.n2511 585
R2870 gnd.n2813 gnd.n2812 585
R2871 gnd.n2812 gnd.n2811 585
R2872 gnd.n2814 gnd.n2506 585
R2873 gnd.n2506 gnd.n2505 585
R2874 gnd.n2816 gnd.n2815 585
R2875 gnd.n2817 gnd.n2816 585
R2876 gnd.n2504 gnd.n2503 585
R2877 gnd.n2818 gnd.n2504 585
R2878 gnd.n2821 gnd.n2820 585
R2879 gnd.n2820 gnd.n2819 585
R2880 gnd.n2500 gnd.n2498 585
R2881 gnd.n2498 gnd.n2497 585
R2882 gnd.n2826 gnd.n2825 585
R2883 gnd.n2827 gnd.n2826 585
R2884 gnd.n2499 gnd.n2496 585
R2885 gnd.n2828 gnd.n2496 585
R2886 gnd.n5691 gnd.n1357 585
R2887 gnd.n5771 gnd.n1357 585
R2888 gnd.n5693 gnd.n5692 585
R2889 gnd.n5694 gnd.n5693 585
R2890 gnd.n1651 gnd.n1650 585
R2891 gnd.n5386 gnd.n1650 585
R2892 gnd.n5569 gnd.n5568 585
R2893 gnd.n5568 gnd.n5567 585
R2894 gnd.n1654 gnd.n1653 585
R2895 gnd.n5384 gnd.n1654 585
R2896 gnd.n5556 gnd.n5555 585
R2897 gnd.n5557 gnd.n5556 585
R2898 gnd.n1670 gnd.n1669 585
R2899 gnd.n5373 gnd.n1669 585
R2900 gnd.n5551 gnd.n5550 585
R2901 gnd.n5550 gnd.n5549 585
R2902 gnd.n1673 gnd.n1672 585
R2903 gnd.n5328 gnd.n1673 585
R2904 gnd.n5540 gnd.n5539 585
R2905 gnd.n5541 gnd.n5540 585
R2906 gnd.n1686 gnd.n1685 585
R2907 gnd.n5334 gnd.n1685 585
R2908 gnd.n5535 gnd.n5534 585
R2909 gnd.n5534 gnd.n5533 585
R2910 gnd.n1689 gnd.n1688 585
R2911 gnd.n5320 gnd.n1689 585
R2912 gnd.n5524 gnd.n5523 585
R2913 gnd.n5525 gnd.n5524 585
R2914 gnd.n1704 gnd.n1703 585
R2915 gnd.n5316 gnd.n1703 585
R2916 gnd.n5519 gnd.n5518 585
R2917 gnd.n5518 gnd.n5517 585
R2918 gnd.n1707 gnd.n1706 585
R2919 gnd.n5289 gnd.n1707 585
R2920 gnd.n5508 gnd.n5507 585
R2921 gnd.n5509 gnd.n5508 585
R2922 gnd.n1720 gnd.n1719 585
R2923 gnd.n5295 gnd.n1719 585
R2924 gnd.n5503 gnd.n5502 585
R2925 gnd.n5502 gnd.n5501 585
R2926 gnd.n1723 gnd.n1722 585
R2927 gnd.n5280 gnd.n1723 585
R2928 gnd.n5492 gnd.n5491 585
R2929 gnd.n5493 gnd.n5492 585
R2930 gnd.n1738 gnd.n1737 585
R2931 gnd.n5276 gnd.n1737 585
R2932 gnd.n5487 gnd.n5486 585
R2933 gnd.n5486 gnd.n5485 585
R2934 gnd.n1741 gnd.n1740 585
R2935 gnd.n5249 gnd.n1741 585
R2936 gnd.n5476 gnd.n5475 585
R2937 gnd.n5477 gnd.n5476 585
R2938 gnd.n1754 gnd.n1753 585
R2939 gnd.n5429 gnd.n1753 585
R2940 gnd.n5471 gnd.n5470 585
R2941 gnd.n5470 gnd.n5469 585
R2942 gnd.n1757 gnd.n1756 585
R2943 gnd.n5241 gnd.n1757 585
R2944 gnd.n5443 gnd.n5442 585
R2945 gnd.n5442 gnd.n5441 585
R2946 gnd.n5444 gnd.n1791 585
R2947 gnd.n5233 gnd.n1791 585
R2948 gnd.n5446 gnd.n5445 585
R2949 gnd.n5447 gnd.n5446 585
R2950 gnd.n1783 gnd.n1782 585
R2951 gnd.n1786 gnd.n1783 585
R2952 gnd.n5457 gnd.n5456 585
R2953 gnd.n5456 gnd.n5455 585
R2954 gnd.n5458 gnd.n1777 585
R2955 gnd.n1777 gnd.n1775 585
R2956 gnd.n5460 gnd.n5459 585
R2957 gnd.n5461 gnd.n5460 585
R2958 gnd.n1778 gnd.n1776 585
R2959 gnd.n5217 gnd.n1776 585
R2960 gnd.n1895 gnd.n1894 585
R2961 gnd.n1894 gnd.n1867 585
R2962 gnd.n1896 gnd.n1874 585
R2963 gnd.n5199 gnd.n1874 585
R2964 gnd.n5186 gnd.n5185 585
R2965 gnd.n5185 gnd.n5184 585
R2966 gnd.n5187 gnd.n1886 585
R2967 gnd.n1886 gnd.n1884 585
R2968 gnd.n5189 gnd.n5188 585
R2969 gnd.n5190 gnd.n5189 585
R2970 gnd.n1887 gnd.n1885 585
R2971 gnd.n5173 gnd.n1885 585
R2972 gnd.n5145 gnd.n5144 585
R2973 gnd.n5144 gnd.n1902 585
R2974 gnd.n5146 gnd.n1910 585
R2975 gnd.n5160 gnd.n1910 585
R2976 gnd.n5147 gnd.n1920 585
R2977 gnd.n1920 gnd.n1908 585
R2978 gnd.n5149 gnd.n5148 585
R2979 gnd.n5150 gnd.n5149 585
R2980 gnd.n1921 gnd.n1919 585
R2981 gnd.n1928 gnd.n1919 585
R2982 gnd.n5136 gnd.n5135 585
R2983 gnd.n5135 gnd.n5134 585
R2984 gnd.n1924 gnd.n1923 585
R2985 gnd.n1925 gnd.n1924 585
R2986 gnd.n5125 gnd.n5124 585
R2987 gnd.n5126 gnd.n5125 585
R2988 gnd.n1938 gnd.n1937 585
R2989 gnd.n1937 gnd.n1934 585
R2990 gnd.n5120 gnd.n5119 585
R2991 gnd.n5119 gnd.n5118 585
R2992 gnd.n1941 gnd.n1940 585
R2993 gnd.n1942 gnd.n1941 585
R2994 gnd.n5109 gnd.n5108 585
R2995 gnd.n5110 gnd.n5109 585
R2996 gnd.n1953 gnd.n1952 585
R2997 gnd.n1960 gnd.n1952 585
R2998 gnd.n5104 gnd.n5103 585
R2999 gnd.n5103 gnd.n5102 585
R3000 gnd.n1956 gnd.n1955 585
R3001 gnd.n1957 gnd.n1956 585
R3002 gnd.n5093 gnd.n5092 585
R3003 gnd.n5094 gnd.n5093 585
R3004 gnd.n1970 gnd.n1969 585
R3005 gnd.n1969 gnd.n1966 585
R3006 gnd.n5088 gnd.n5087 585
R3007 gnd.n5087 gnd.n5086 585
R3008 gnd.n1973 gnd.n1972 585
R3009 gnd.n1974 gnd.n1973 585
R3010 gnd.n5077 gnd.n5076 585
R3011 gnd.n5078 gnd.n5077 585
R3012 gnd.n1985 gnd.n1984 585
R3013 gnd.n4872 gnd.n1984 585
R3014 gnd.n5072 gnd.n5071 585
R3015 gnd.n5071 gnd.n5070 585
R3016 gnd.n4779 gnd.n1987 585
R3017 gnd.n4782 gnd.n4780 585
R3018 gnd.n4785 gnd.n4784 585
R3019 gnd.n4777 gnd.n4776 585
R3020 gnd.n4790 gnd.n4789 585
R3021 gnd.n4792 gnd.n4775 585
R3022 gnd.n4795 gnd.n4794 585
R3023 gnd.n4773 gnd.n4772 585
R3024 gnd.n4800 gnd.n4799 585
R3025 gnd.n4802 gnd.n4771 585
R3026 gnd.n4805 gnd.n4804 585
R3027 gnd.n4769 gnd.n4768 585
R3028 gnd.n4810 gnd.n4809 585
R3029 gnd.n4812 gnd.n4767 585
R3030 gnd.n4815 gnd.n4814 585
R3031 gnd.n4765 gnd.n4764 585
R3032 gnd.n4820 gnd.n4819 585
R3033 gnd.n4822 gnd.n4763 585
R3034 gnd.n4824 gnd.n4823 585
R3035 gnd.n4823 gnd.n4756 585
R3036 gnd.n5774 gnd.n5773 585
R3037 gnd.n5775 gnd.n1350 585
R3038 gnd.n5627 gnd.n1347 585
R3039 gnd.n5630 gnd.n5629 585
R3040 gnd.n5640 gnd.n5626 585
R3041 gnd.n5641 gnd.n5624 585
R3042 gnd.n5623 gnd.n5614 585
R3043 gnd.n5648 gnd.n5613 585
R3044 gnd.n5649 gnd.n5612 585
R3045 gnd.n5610 gnd.n5604 585
R3046 gnd.n5656 gnd.n5603 585
R3047 gnd.n5657 gnd.n5601 585
R3048 gnd.n5600 gnd.n5591 585
R3049 gnd.n5664 gnd.n5590 585
R3050 gnd.n5665 gnd.n5589 585
R3051 gnd.n5587 gnd.n5579 585
R3052 gnd.n5672 gnd.n5578 585
R3053 gnd.n5673 gnd.n5576 585
R3054 gnd.n5575 gnd.n5573 585
R3055 gnd.n5575 gnd.n1364 585
R3056 gnd.n5772 gnd.n1353 585
R3057 gnd.n5772 gnd.n5771 585
R3058 gnd.n5388 gnd.n1352 585
R3059 gnd.n5694 gnd.n1352 585
R3060 gnd.n5391 gnd.n5387 585
R3061 gnd.n5387 gnd.n5386 585
R3062 gnd.n5392 gnd.n1657 585
R3063 gnd.n5567 gnd.n1657 585
R3064 gnd.n5393 gnd.n5385 585
R3065 gnd.n5385 gnd.n5384 585
R3066 gnd.n1829 gnd.n1667 585
R3067 gnd.n5557 gnd.n1667 585
R3068 gnd.n5397 gnd.n1828 585
R3069 gnd.n5373 gnd.n1828 585
R3070 gnd.n5398 gnd.n1676 585
R3071 gnd.n5549 gnd.n1676 585
R3072 gnd.n5399 gnd.n1827 585
R3073 gnd.n5328 gnd.n1827 585
R3074 gnd.n1825 gnd.n1683 585
R3075 gnd.n5541 gnd.n1683 585
R3076 gnd.n5403 gnd.n1824 585
R3077 gnd.n5334 gnd.n1824 585
R3078 gnd.n5404 gnd.n1692 585
R3079 gnd.n5533 gnd.n1692 585
R3080 gnd.n5405 gnd.n1823 585
R3081 gnd.n5320 gnd.n1823 585
R3082 gnd.n1821 gnd.n1701 585
R3083 gnd.n5525 gnd.n1701 585
R3084 gnd.n5409 gnd.n1820 585
R3085 gnd.n5316 gnd.n1820 585
R3086 gnd.n5410 gnd.n1710 585
R3087 gnd.n5517 gnd.n1710 585
R3088 gnd.n5411 gnd.n1819 585
R3089 gnd.n5289 gnd.n1819 585
R3090 gnd.n1817 gnd.n1717 585
R3091 gnd.n5509 gnd.n1717 585
R3092 gnd.n5415 gnd.n1816 585
R3093 gnd.n5295 gnd.n1816 585
R3094 gnd.n5416 gnd.n1726 585
R3095 gnd.n5501 gnd.n1726 585
R3096 gnd.n5417 gnd.n1815 585
R3097 gnd.n5280 gnd.n1815 585
R3098 gnd.n1813 gnd.n1735 585
R3099 gnd.n5493 gnd.n1735 585
R3100 gnd.n5421 gnd.n1812 585
R3101 gnd.n5276 gnd.n1812 585
R3102 gnd.n5422 gnd.n1744 585
R3103 gnd.n5485 gnd.n1744 585
R3104 gnd.n5423 gnd.n1811 585
R3105 gnd.n5249 gnd.n1811 585
R3106 gnd.n1808 gnd.n1751 585
R3107 gnd.n5477 gnd.n1751 585
R3108 gnd.n5428 gnd.n5427 585
R3109 gnd.n5429 gnd.n5428 585
R3110 gnd.n1807 gnd.n1760 585
R3111 gnd.n5469 gnd.n1760 585
R3112 gnd.n5240 gnd.n5239 585
R3113 gnd.n5241 gnd.n5240 585
R3114 gnd.n1857 gnd.n1797 585
R3115 gnd.n5441 gnd.n1797 585
R3116 gnd.n5235 gnd.n5234 585
R3117 gnd.n5234 gnd.n5233 585
R3118 gnd.n1859 gnd.n1790 585
R3119 gnd.n5447 gnd.n1790 585
R3120 gnd.n5210 gnd.n5208 585
R3121 gnd.n5208 gnd.n1786 585
R3122 gnd.n5211 gnd.n1785 585
R3123 gnd.n5455 gnd.n1785 585
R3124 gnd.n5213 gnd.n5212 585
R3125 gnd.n5212 gnd.n1775 585
R3126 gnd.n5214 gnd.n1774 585
R3127 gnd.n5461 gnd.n1774 585
R3128 gnd.n5216 gnd.n5215 585
R3129 gnd.n5217 gnd.n5216 585
R3130 gnd.n1869 gnd.n1868 585
R3131 gnd.n1868 gnd.n1867 585
R3132 gnd.n5201 gnd.n5200 585
R3133 gnd.n5200 gnd.n5199 585
R3134 gnd.n1872 gnd.n1871 585
R3135 gnd.n5184 gnd.n1872 585
R3136 gnd.n5169 gnd.n5168 585
R3137 gnd.n5168 gnd.n1884 585
R3138 gnd.n5170 gnd.n1883 585
R3139 gnd.n5190 gnd.n1883 585
R3140 gnd.n5172 gnd.n5171 585
R3141 gnd.n5173 gnd.n5172 585
R3142 gnd.n1904 gnd.n1903 585
R3143 gnd.n1903 gnd.n1902 585
R3144 gnd.n5162 gnd.n5161 585
R3145 gnd.n5161 gnd.n5160 585
R3146 gnd.n1907 gnd.n1906 585
R3147 gnd.n1908 gnd.n1907 585
R3148 gnd.n4845 gnd.n1918 585
R3149 gnd.n5150 gnd.n1918 585
R3150 gnd.n4847 gnd.n4846 585
R3151 gnd.n4846 gnd.n1928 585
R3152 gnd.n4848 gnd.n1927 585
R3153 gnd.n5134 gnd.n1927 585
R3154 gnd.n4850 gnd.n4849 585
R3155 gnd.n4849 gnd.n1925 585
R3156 gnd.n4851 gnd.n1936 585
R3157 gnd.n5126 gnd.n1936 585
R3158 gnd.n4853 gnd.n4852 585
R3159 gnd.n4852 gnd.n1934 585
R3160 gnd.n4854 gnd.n1944 585
R3161 gnd.n5118 gnd.n1944 585
R3162 gnd.n4856 gnd.n4855 585
R3163 gnd.n4855 gnd.n1942 585
R3164 gnd.n4857 gnd.n1951 585
R3165 gnd.n5110 gnd.n1951 585
R3166 gnd.n4859 gnd.n4858 585
R3167 gnd.n4858 gnd.n1960 585
R3168 gnd.n4860 gnd.n1959 585
R3169 gnd.n5102 gnd.n1959 585
R3170 gnd.n4862 gnd.n4861 585
R3171 gnd.n4861 gnd.n1957 585
R3172 gnd.n4863 gnd.n1968 585
R3173 gnd.n5094 gnd.n1968 585
R3174 gnd.n4865 gnd.n4864 585
R3175 gnd.n4864 gnd.n1966 585
R3176 gnd.n4866 gnd.n1976 585
R3177 gnd.n5086 gnd.n1976 585
R3178 gnd.n4868 gnd.n4867 585
R3179 gnd.n4867 gnd.n1974 585
R3180 gnd.n4869 gnd.n1983 585
R3181 gnd.n5078 gnd.n1983 585
R3182 gnd.n4871 gnd.n4870 585
R3183 gnd.n4872 gnd.n4871 585
R3184 gnd.n4759 gnd.n4758 585
R3185 gnd.n5070 gnd.n4758 585
R3186 gnd.n7477 gnd.n125 585
R3187 gnd.n7573 gnd.n125 585
R3188 gnd.n7478 gnd.n7415 585
R3189 gnd.n7415 gnd.n122 585
R3190 gnd.n7479 gnd.n203 585
R3191 gnd.n7493 gnd.n203 585
R3192 gnd.n215 gnd.n213 585
R3193 gnd.n213 gnd.n202 585
R3194 gnd.n7484 gnd.n7483 585
R3195 gnd.n7485 gnd.n7484 585
R3196 gnd.n214 gnd.n212 585
R3197 gnd.n212 gnd.n209 585
R3198 gnd.n7411 gnd.n7410 585
R3199 gnd.n7410 gnd.n7409 585
R3200 gnd.n218 gnd.n217 585
R3201 gnd.n228 gnd.n218 585
R3202 gnd.n7400 gnd.n7399 585
R3203 gnd.n7401 gnd.n7400 585
R3204 gnd.n230 gnd.n229 585
R3205 gnd.n229 gnd.n225 585
R3206 gnd.n7395 gnd.n7394 585
R3207 gnd.n7394 gnd.n7393 585
R3208 gnd.n233 gnd.n232 585
R3209 gnd.n234 gnd.n233 585
R3210 gnd.n7384 gnd.n7383 585
R3211 gnd.n7385 gnd.n7384 585
R3212 gnd.n245 gnd.n244 585
R3213 gnd.n250 gnd.n244 585
R3214 gnd.n7379 gnd.n7378 585
R3215 gnd.n7378 gnd.n7377 585
R3216 gnd.n248 gnd.n247 585
R3217 gnd.n259 gnd.n248 585
R3218 gnd.n7368 gnd.n7367 585
R3219 gnd.n7369 gnd.n7368 585
R3220 gnd.n261 gnd.n260 585
R3221 gnd.n260 gnd.n256 585
R3222 gnd.n7363 gnd.n7362 585
R3223 gnd.n7362 gnd.n7361 585
R3224 gnd.n264 gnd.n263 585
R3225 gnd.n265 gnd.n264 585
R3226 gnd.n7352 gnd.n7351 585
R3227 gnd.n7353 gnd.n7352 585
R3228 gnd.n275 gnd.n274 585
R3229 gnd.n280 gnd.n274 585
R3230 gnd.n7347 gnd.n7346 585
R3231 gnd.n7346 gnd.n7345 585
R3232 gnd.n278 gnd.n277 585
R3233 gnd.n289 gnd.n278 585
R3234 gnd.n7336 gnd.n7335 585
R3235 gnd.n7337 gnd.n7336 585
R3236 gnd.n291 gnd.n290 585
R3237 gnd.n290 gnd.n286 585
R3238 gnd.n7331 gnd.n7330 585
R3239 gnd.n7330 gnd.n7329 585
R3240 gnd.n294 gnd.n293 585
R3241 gnd.n295 gnd.n294 585
R3242 gnd.n7307 gnd.n7306 585
R3243 gnd.n7306 gnd.n7305 585
R3244 gnd.n7308 gnd.n323 585
R3245 gnd.n7301 gnd.n323 585
R3246 gnd.n329 gnd.n321 585
R3247 gnd.n330 gnd.n329 585
R3248 gnd.n7312 gnd.n320 585
R3249 gnd.n7228 gnd.n320 585
R3250 gnd.n7313 gnd.n319 585
R3251 gnd.n336 gnd.n319 585
R3252 gnd.n7314 gnd.n318 585
R3253 gnd.n7222 gnd.n318 585
R3254 gnd.n315 gnd.n313 585
R3255 gnd.n7202 gnd.n313 585
R3256 gnd.n7319 gnd.n7318 585
R3257 gnd.n7320 gnd.n7319 585
R3258 gnd.n314 gnd.n312 585
R3259 gnd.n7211 gnd.n312 585
R3260 gnd.n7173 gnd.n7171 585
R3261 gnd.n7171 gnd.n349 585
R3262 gnd.n7174 gnd.n362 585
R3263 gnd.n7190 gnd.n362 585
R3264 gnd.n7175 gnd.n7170 585
R3265 gnd.n7170 gnd.n7169 585
R3266 gnd.n376 gnd.n374 585
R3267 gnd.n6930 gnd.n374 585
R3268 gnd.n7180 gnd.n7179 585
R3269 gnd.n7181 gnd.n7180 585
R3270 gnd.n375 gnd.n373 585
R3271 gnd.n7159 gnd.n373 585
R3272 gnd.n7124 gnd.n395 585
R3273 gnd.n7138 gnd.n395 585
R3274 gnd.n408 gnd.n406 585
R3275 gnd.n6938 gnd.n406 585
R3276 gnd.n7129 gnd.n7128 585
R3277 gnd.n7130 gnd.n7129 585
R3278 gnd.n407 gnd.n405 585
R3279 gnd.n6917 gnd.n405 585
R3280 gnd.n7121 gnd.n7120 585
R3281 gnd.n7120 gnd.n7119 585
R3282 gnd.n411 gnd.n410 585
R3283 gnd.n6898 gnd.n411 585
R3284 gnd.n7110 gnd.n7109 585
R3285 gnd.n7111 gnd.n7110 585
R3286 gnd.n424 gnd.n423 585
R3287 gnd.n6904 gnd.n423 585
R3288 gnd.n7105 gnd.n7104 585
R3289 gnd.n7104 gnd.n7103 585
R3290 gnd.n427 gnd.n426 585
R3291 gnd.n6890 gnd.n427 585
R3292 gnd.n7094 gnd.n7093 585
R3293 gnd.n7095 gnd.n7094 585
R3294 gnd.n442 gnd.n441 585
R3295 gnd.n6886 gnd.n441 585
R3296 gnd.n7089 gnd.n7088 585
R3297 gnd.n7088 gnd.n7087 585
R3298 gnd.n445 gnd.n444 585
R3299 gnd.n6859 gnd.n445 585
R3300 gnd.n7078 gnd.n7077 585
R3301 gnd.n7079 gnd.n7078 585
R3302 gnd.n458 gnd.n457 585
R3303 gnd.n6865 gnd.n457 585
R3304 gnd.n7073 gnd.n7072 585
R3305 gnd.n7072 gnd.n7071 585
R3306 gnd.n461 gnd.n460 585
R3307 gnd.n6850 gnd.n461 585
R3308 gnd.n7062 gnd.n7061 585
R3309 gnd.n7063 gnd.n7062 585
R3310 gnd.n476 gnd.n475 585
R3311 gnd.n6846 gnd.n475 585
R3312 gnd.n7057 gnd.n7056 585
R3313 gnd.n7056 gnd.n7055 585
R3314 gnd.n479 gnd.n478 585
R3315 gnd.n6974 gnd.n479 585
R3316 gnd.n6622 gnd.n6621 585
R3317 gnd.n6624 gnd.n6623 585
R3318 gnd.n6754 gnd.n6625 585
R3319 gnd.n6753 gnd.n6626 585
R3320 gnd.n6628 gnd.n6627 585
R3321 gnd.n6746 gnd.n6636 585
R3322 gnd.n6745 gnd.n6637 585
R3323 gnd.n6644 gnd.n6638 585
R3324 gnd.n6738 gnd.n6645 585
R3325 gnd.n6737 gnd.n6646 585
R3326 gnd.n6648 gnd.n6647 585
R3327 gnd.n6730 gnd.n6656 585
R3328 gnd.n6729 gnd.n6657 585
R3329 gnd.n6664 gnd.n6658 585
R3330 gnd.n6722 gnd.n6665 585
R3331 gnd.n6721 gnd.n6666 585
R3332 gnd.n6668 gnd.n6667 585
R3333 gnd.n6714 gnd.n6711 585
R3334 gnd.n6710 gnd.n517 585
R3335 gnd.n7046 gnd.n517 585
R3336 gnd.n7576 gnd.n7575 585
R3337 gnd.n7448 gnd.n120 585
R3338 gnd.n7450 gnd.n7449 585
R3339 gnd.n7446 gnd.n7445 585
R3340 gnd.n7454 gnd.n7444 585
R3341 gnd.n7455 gnd.n7442 585
R3342 gnd.n7456 gnd.n7441 585
R3343 gnd.n7439 gnd.n7437 585
R3344 gnd.n7460 gnd.n7436 585
R3345 gnd.n7461 gnd.n7434 585
R3346 gnd.n7462 gnd.n7433 585
R3347 gnd.n7431 gnd.n7429 585
R3348 gnd.n7466 gnd.n7428 585
R3349 gnd.n7467 gnd.n7426 585
R3350 gnd.n7468 gnd.n7425 585
R3351 gnd.n7423 gnd.n7421 585
R3352 gnd.n7472 gnd.n7420 585
R3353 gnd.n7473 gnd.n7418 585
R3354 gnd.n7474 gnd.n7417 585
R3355 gnd.n7417 gnd.n124 585
R3356 gnd.n7574 gnd.n116 585
R3357 gnd.n7574 gnd.n7573 585
R3358 gnd.n7580 gnd.n115 585
R3359 gnd.n122 gnd.n115 585
R3360 gnd.n7581 gnd.n114 585
R3361 gnd.n7493 gnd.n114 585
R3362 gnd.n7582 gnd.n113 585
R3363 gnd.n202 gnd.n113 585
R3364 gnd.n211 gnd.n111 585
R3365 gnd.n7485 gnd.n211 585
R3366 gnd.n7586 gnd.n110 585
R3367 gnd.n209 gnd.n110 585
R3368 gnd.n7587 gnd.n109 585
R3369 gnd.n7409 gnd.n109 585
R3370 gnd.n7588 gnd.n108 585
R3371 gnd.n228 gnd.n108 585
R3372 gnd.n227 gnd.n106 585
R3373 gnd.n7401 gnd.n227 585
R3374 gnd.n7592 gnd.n105 585
R3375 gnd.n225 gnd.n105 585
R3376 gnd.n7593 gnd.n104 585
R3377 gnd.n7393 gnd.n104 585
R3378 gnd.n7594 gnd.n103 585
R3379 gnd.n234 gnd.n103 585
R3380 gnd.n243 gnd.n101 585
R3381 gnd.n7385 gnd.n243 585
R3382 gnd.n7598 gnd.n100 585
R3383 gnd.n250 gnd.n100 585
R3384 gnd.n7599 gnd.n99 585
R3385 gnd.n7377 gnd.n99 585
R3386 gnd.n7600 gnd.n98 585
R3387 gnd.n259 gnd.n98 585
R3388 gnd.n258 gnd.n96 585
R3389 gnd.n7369 gnd.n258 585
R3390 gnd.n7604 gnd.n95 585
R3391 gnd.n256 gnd.n95 585
R3392 gnd.n7605 gnd.n94 585
R3393 gnd.n7361 gnd.n94 585
R3394 gnd.n7606 gnd.n93 585
R3395 gnd.n265 gnd.n93 585
R3396 gnd.n273 gnd.n91 585
R3397 gnd.n7353 gnd.n273 585
R3398 gnd.n7610 gnd.n90 585
R3399 gnd.n280 gnd.n90 585
R3400 gnd.n7611 gnd.n89 585
R3401 gnd.n7345 gnd.n89 585
R3402 gnd.n7612 gnd.n88 585
R3403 gnd.n289 gnd.n88 585
R3404 gnd.n288 gnd.n86 585
R3405 gnd.n7337 gnd.n288 585
R3406 gnd.n7616 gnd.n85 585
R3407 gnd.n286 gnd.n85 585
R3408 gnd.n7617 gnd.n84 585
R3409 gnd.n7329 gnd.n84 585
R3410 gnd.n7618 gnd.n83 585
R3411 gnd.n295 gnd.n83 585
R3412 gnd.n325 gnd.n81 585
R3413 gnd.n7305 gnd.n325 585
R3414 gnd.n7622 gnd.n80 585
R3415 gnd.n7301 gnd.n80 585
R3416 gnd.n7623 gnd.n79 585
R3417 gnd.n330 gnd.n79 585
R3418 gnd.n7624 gnd.n78 585
R3419 gnd.n7228 gnd.n78 585
R3420 gnd.n340 gnd.n76 585
R3421 gnd.n340 gnd.n336 585
R3422 gnd.n7204 gnd.n341 585
R3423 gnd.n7222 gnd.n341 585
R3424 gnd.n7205 gnd.n7203 585
R3425 gnd.n7203 gnd.n7202 585
R3426 gnd.n353 gnd.n310 585
R3427 gnd.n7320 gnd.n310 585
R3428 gnd.n7210 gnd.n7209 585
R3429 gnd.n7211 gnd.n7210 585
R3430 gnd.n352 gnd.n351 585
R3431 gnd.n351 gnd.n349 585
R3432 gnd.n382 gnd.n360 585
R3433 gnd.n7190 gnd.n360 585
R3434 gnd.n7168 gnd.n7167 585
R3435 gnd.n7169 gnd.n7168 585
R3436 gnd.n381 gnd.n380 585
R3437 gnd.n6930 gnd.n380 585
R3438 gnd.n7162 gnd.n371 585
R3439 gnd.n7181 gnd.n371 585
R3440 gnd.n7161 gnd.n7160 585
R3441 gnd.n7160 gnd.n7159 585
R3442 gnd.n385 gnd.n384 585
R3443 gnd.n7138 gnd.n385 585
R3444 gnd.n6942 gnd.n6939 585
R3445 gnd.n6939 gnd.n6938 585
R3446 gnd.n6943 gnd.n403 585
R3447 gnd.n7130 gnd.n403 585
R3448 gnd.n6944 gnd.n584 585
R3449 gnd.n6917 gnd.n584 585
R3450 gnd.n582 gnd.n414 585
R3451 gnd.n7119 gnd.n414 585
R3452 gnd.n6948 gnd.n581 585
R3453 gnd.n6898 gnd.n581 585
R3454 gnd.n6949 gnd.n421 585
R3455 gnd.n7111 gnd.n421 585
R3456 gnd.n6950 gnd.n580 585
R3457 gnd.n6904 gnd.n580 585
R3458 gnd.n578 gnd.n430 585
R3459 gnd.n7103 gnd.n430 585
R3460 gnd.n6954 gnd.n577 585
R3461 gnd.n6890 gnd.n577 585
R3462 gnd.n6955 gnd.n439 585
R3463 gnd.n7095 gnd.n439 585
R3464 gnd.n6956 gnd.n576 585
R3465 gnd.n6886 gnd.n576 585
R3466 gnd.n574 gnd.n448 585
R3467 gnd.n7087 gnd.n448 585
R3468 gnd.n6960 gnd.n573 585
R3469 gnd.n6859 gnd.n573 585
R3470 gnd.n6961 gnd.n455 585
R3471 gnd.n7079 gnd.n455 585
R3472 gnd.n6962 gnd.n572 585
R3473 gnd.n6865 gnd.n572 585
R3474 gnd.n570 gnd.n464 585
R3475 gnd.n7071 gnd.n464 585
R3476 gnd.n6966 gnd.n569 585
R3477 gnd.n6850 gnd.n569 585
R3478 gnd.n6967 gnd.n473 585
R3479 gnd.n7063 gnd.n473 585
R3480 gnd.n6968 gnd.n568 585
R3481 gnd.n6846 gnd.n568 585
R3482 gnd.n565 gnd.n482 585
R3483 gnd.n7055 gnd.n482 585
R3484 gnd.n6973 gnd.n6972 585
R3485 gnd.n6974 gnd.n6973 585
R3486 gnd.n4663 gnd.n4662 585
R3487 gnd.n4664 gnd.n4663 585
R3488 gnd.n3357 gnd.n3356 585
R3489 gnd.n3364 gnd.n3356 585
R3490 gnd.n4645 gnd.n4644 585
R3491 gnd.n4646 gnd.n4645 585
R3492 gnd.n3375 gnd.n3374 585
R3493 gnd.n3374 gnd.n3370 585
R3494 gnd.n4635 gnd.n4634 585
R3495 gnd.n4636 gnd.n4635 585
R3496 gnd.n3383 gnd.n3382 585
R3497 gnd.n3388 gnd.n3382 585
R3498 gnd.n4357 gnd.n3400 585
R3499 gnd.n3400 gnd.n3387 585
R3500 gnd.n4359 gnd.n4358 585
R3501 gnd.n4360 gnd.n4359 585
R3502 gnd.n3401 gnd.n3399 585
R3503 gnd.n3399 gnd.n3395 585
R3504 gnd.n4348 gnd.n4347 585
R3505 gnd.n4349 gnd.n4348 585
R3506 gnd.n3408 gnd.n3407 585
R3507 gnd.n3413 gnd.n3407 585
R3508 gnd.n4326 gnd.n3426 585
R3509 gnd.n3426 gnd.n3412 585
R3510 gnd.n4328 gnd.n4327 585
R3511 gnd.n4329 gnd.n4328 585
R3512 gnd.n3427 gnd.n3425 585
R3513 gnd.n3425 gnd.n3421 585
R3514 gnd.n4317 gnd.n4316 585
R3515 gnd.n4318 gnd.n4317 585
R3516 gnd.n3434 gnd.n3433 585
R3517 gnd.n3438 gnd.n3433 585
R3518 gnd.n4295 gnd.n3450 585
R3519 gnd.n3588 gnd.n3450 585
R3520 gnd.n4297 gnd.n4296 585
R3521 gnd.n4298 gnd.n4297 585
R3522 gnd.n3451 gnd.n3449 585
R3523 gnd.n3449 gnd.n3446 585
R3524 gnd.n4286 gnd.n4285 585
R3525 gnd.n4287 gnd.n4286 585
R3526 gnd.n3458 gnd.n3457 585
R3527 gnd.n3463 gnd.n3457 585
R3528 gnd.n4264 gnd.n3476 585
R3529 gnd.n3476 gnd.n3462 585
R3530 gnd.n4266 gnd.n4265 585
R3531 gnd.n4267 gnd.n4266 585
R3532 gnd.n3477 gnd.n3475 585
R3533 gnd.n3475 gnd.n3471 585
R3534 gnd.n4255 gnd.n4254 585
R3535 gnd.n4256 gnd.n4255 585
R3536 gnd.n3485 gnd.n3484 585
R3537 gnd.n3490 gnd.n3484 585
R3538 gnd.n4233 gnd.n3502 585
R3539 gnd.n3502 gnd.n3489 585
R3540 gnd.n4235 gnd.n4234 585
R3541 gnd.n4236 gnd.n4235 585
R3542 gnd.n3503 gnd.n3501 585
R3543 gnd.n3501 gnd.n3497 585
R3544 gnd.n4224 gnd.n4223 585
R3545 gnd.n4225 gnd.n4224 585
R3546 gnd.n3510 gnd.n3509 585
R3547 gnd.n3613 gnd.n3509 585
R3548 gnd.n4202 gnd.n3525 585
R3549 gnd.n3525 gnd.n3514 585
R3550 gnd.n4204 gnd.n4203 585
R3551 gnd.n4205 gnd.n4204 585
R3552 gnd.n3526 gnd.n3524 585
R3553 gnd.n4194 gnd.n3524 585
R3554 gnd.n3694 gnd.n3693 585
R3555 gnd.n3694 gnd.n3531 585
R3556 gnd.n4181 gnd.n4180 585
R3557 gnd.n4180 gnd.n4179 585
R3558 gnd.n4182 gnd.n3686 585
R3559 gnd.n4159 gnd.n3686 585
R3560 gnd.n4184 gnd.n4183 585
R3561 gnd.n4185 gnd.n4184 585
R3562 gnd.n3687 gnd.n3685 585
R3563 gnd.n4167 gnd.n3685 585
R3564 gnd.n4151 gnd.n4150 585
R3565 gnd.n4150 gnd.n3704 585
R3566 gnd.n4149 gnd.n3709 585
R3567 gnd.n4149 gnd.n4148 585
R3568 gnd.n4134 gnd.n3710 585
R3569 gnd.n3718 gnd.n3710 585
R3570 gnd.n4136 gnd.n4135 585
R3571 gnd.n4137 gnd.n4136 585
R3572 gnd.n3721 gnd.n3720 585
R3573 gnd.n3728 gnd.n3720 585
R3574 gnd.n4109 gnd.n4108 585
R3575 gnd.n4110 gnd.n4109 585
R3576 gnd.n3740 gnd.n3739 585
R3577 gnd.n3739 gnd.n3735 585
R3578 gnd.n4099 gnd.n4098 585
R3579 gnd.n4100 gnd.n4099 585
R3580 gnd.n3750 gnd.n3749 585
R3581 gnd.n3755 gnd.n3749 585
R3582 gnd.n4077 gnd.n3768 585
R3583 gnd.n3768 gnd.n3754 585
R3584 gnd.n4079 gnd.n4078 585
R3585 gnd.n4080 gnd.n4079 585
R3586 gnd.n3769 gnd.n3767 585
R3587 gnd.n3767 gnd.n3763 585
R3588 gnd.n4068 gnd.n4067 585
R3589 gnd.n4069 gnd.n4068 585
R3590 gnd.n3776 gnd.n3775 585
R3591 gnd.n3780 gnd.n3775 585
R3592 gnd.n4045 gnd.n3797 585
R3593 gnd.n3797 gnd.n3779 585
R3594 gnd.n4047 gnd.n4046 585
R3595 gnd.n4048 gnd.n4047 585
R3596 gnd.n3798 gnd.n3796 585
R3597 gnd.n3796 gnd.n3787 585
R3598 gnd.n4040 gnd.n4039 585
R3599 gnd.n4039 gnd.n4038 585
R3600 gnd.n3845 gnd.n3844 585
R3601 gnd.n3846 gnd.n3845 585
R3602 gnd.n3999 gnd.n3998 585
R3603 gnd.n4000 gnd.n3999 585
R3604 gnd.n3855 gnd.n3854 585
R3605 gnd.n3854 gnd.n3853 585
R3606 gnd.n3994 gnd.n3993 585
R3607 gnd.n3993 gnd.n3992 585
R3608 gnd.n3858 gnd.n3857 585
R3609 gnd.n3859 gnd.n3858 585
R3610 gnd.n3983 gnd.n3982 585
R3611 gnd.n3984 gnd.n3983 585
R3612 gnd.n3866 gnd.n3865 585
R3613 gnd.n3975 gnd.n3865 585
R3614 gnd.n3978 gnd.n3977 585
R3615 gnd.n3977 gnd.n3976 585
R3616 gnd.n3869 gnd.n3868 585
R3617 gnd.n3870 gnd.n3869 585
R3618 gnd.n3964 gnd.n3963 585
R3619 gnd.n3962 gnd.n3888 585
R3620 gnd.n3961 gnd.n3887 585
R3621 gnd.n3966 gnd.n3887 585
R3622 gnd.n3960 gnd.n3959 585
R3623 gnd.n3958 gnd.n3957 585
R3624 gnd.n3956 gnd.n3955 585
R3625 gnd.n3954 gnd.n3953 585
R3626 gnd.n3952 gnd.n3951 585
R3627 gnd.n3950 gnd.n3949 585
R3628 gnd.n3948 gnd.n3947 585
R3629 gnd.n3946 gnd.n3945 585
R3630 gnd.n3944 gnd.n3943 585
R3631 gnd.n3942 gnd.n3941 585
R3632 gnd.n3940 gnd.n3939 585
R3633 gnd.n3938 gnd.n3937 585
R3634 gnd.n3936 gnd.n3935 585
R3635 gnd.n3934 gnd.n3933 585
R3636 gnd.n3932 gnd.n3931 585
R3637 gnd.n3930 gnd.n3929 585
R3638 gnd.n3928 gnd.n3927 585
R3639 gnd.n3926 gnd.n3925 585
R3640 gnd.n3924 gnd.n3923 585
R3641 gnd.n3922 gnd.n3921 585
R3642 gnd.n3920 gnd.n3919 585
R3643 gnd.n3918 gnd.n3917 585
R3644 gnd.n3875 gnd.n3874 585
R3645 gnd.n3969 gnd.n3968 585
R3646 gnd.n4667 gnd.n4666 585
R3647 gnd.n4669 gnd.n4668 585
R3648 gnd.n4671 gnd.n4670 585
R3649 gnd.n4673 gnd.n4672 585
R3650 gnd.n4675 gnd.n4674 585
R3651 gnd.n4677 gnd.n4676 585
R3652 gnd.n4679 gnd.n4678 585
R3653 gnd.n4681 gnd.n4680 585
R3654 gnd.n4683 gnd.n4682 585
R3655 gnd.n4685 gnd.n4684 585
R3656 gnd.n4687 gnd.n4686 585
R3657 gnd.n4689 gnd.n4688 585
R3658 gnd.n4691 gnd.n4690 585
R3659 gnd.n4693 gnd.n4692 585
R3660 gnd.n4695 gnd.n4694 585
R3661 gnd.n4697 gnd.n4696 585
R3662 gnd.n4699 gnd.n4698 585
R3663 gnd.n4701 gnd.n4700 585
R3664 gnd.n4703 gnd.n4702 585
R3665 gnd.n4705 gnd.n4704 585
R3666 gnd.n4707 gnd.n4706 585
R3667 gnd.n4709 gnd.n4708 585
R3668 gnd.n4711 gnd.n4710 585
R3669 gnd.n4713 gnd.n4712 585
R3670 gnd.n4715 gnd.n4714 585
R3671 gnd.n4716 gnd.n2031 585
R3672 gnd.n4717 gnd.n1989 585
R3673 gnd.n4755 gnd.n1989 585
R3674 gnd.n4665 gnd.n2061 585
R3675 gnd.n4665 gnd.n4664 585
R3676 gnd.n3564 gnd.n2060 585
R3677 gnd.n3364 gnd.n2060 585
R3678 gnd.n3565 gnd.n3372 585
R3679 gnd.n4646 gnd.n3372 585
R3680 gnd.n3567 gnd.n3566 585
R3681 gnd.n3566 gnd.n3370 585
R3682 gnd.n3568 gnd.n3381 585
R3683 gnd.n4636 gnd.n3381 585
R3684 gnd.n3570 gnd.n3569 585
R3685 gnd.n3570 gnd.n3388 585
R3686 gnd.n3572 gnd.n3571 585
R3687 gnd.n3571 gnd.n3387 585
R3688 gnd.n3573 gnd.n3397 585
R3689 gnd.n4360 gnd.n3397 585
R3690 gnd.n3575 gnd.n3574 585
R3691 gnd.n3574 gnd.n3395 585
R3692 gnd.n3576 gnd.n3406 585
R3693 gnd.n4349 gnd.n3406 585
R3694 gnd.n3578 gnd.n3577 585
R3695 gnd.n3578 gnd.n3413 585
R3696 gnd.n3580 gnd.n3579 585
R3697 gnd.n3579 gnd.n3412 585
R3698 gnd.n3581 gnd.n3423 585
R3699 gnd.n4329 gnd.n3423 585
R3700 gnd.n3583 gnd.n3582 585
R3701 gnd.n3582 gnd.n3421 585
R3702 gnd.n3584 gnd.n3432 585
R3703 gnd.n4318 gnd.n3432 585
R3704 gnd.n3586 gnd.n3585 585
R3705 gnd.n3586 gnd.n3438 585
R3706 gnd.n3590 gnd.n3589 585
R3707 gnd.n3589 gnd.n3588 585
R3708 gnd.n3591 gnd.n3448 585
R3709 gnd.n4298 gnd.n3448 585
R3710 gnd.n3593 gnd.n3592 585
R3711 gnd.n3592 gnd.n3446 585
R3712 gnd.n3594 gnd.n3456 585
R3713 gnd.n4287 gnd.n3456 585
R3714 gnd.n3596 gnd.n3595 585
R3715 gnd.n3596 gnd.n3463 585
R3716 gnd.n3598 gnd.n3597 585
R3717 gnd.n3597 gnd.n3462 585
R3718 gnd.n3599 gnd.n3473 585
R3719 gnd.n4267 gnd.n3473 585
R3720 gnd.n3601 gnd.n3600 585
R3721 gnd.n3600 gnd.n3471 585
R3722 gnd.n3602 gnd.n3483 585
R3723 gnd.n4256 gnd.n3483 585
R3724 gnd.n3604 gnd.n3603 585
R3725 gnd.n3604 gnd.n3490 585
R3726 gnd.n3606 gnd.n3605 585
R3727 gnd.n3605 gnd.n3489 585
R3728 gnd.n3607 gnd.n3499 585
R3729 gnd.n4236 gnd.n3499 585
R3730 gnd.n3609 gnd.n3608 585
R3731 gnd.n3608 gnd.n3497 585
R3732 gnd.n3610 gnd.n3508 585
R3733 gnd.n4225 gnd.n3508 585
R3734 gnd.n3615 gnd.n3614 585
R3735 gnd.n3614 gnd.n3613 585
R3736 gnd.n3611 gnd.n3534 585
R3737 gnd.n3611 gnd.n3514 585
R3738 gnd.n4191 gnd.n3522 585
R3739 gnd.n4205 gnd.n3522 585
R3740 gnd.n4193 gnd.n4192 585
R3741 gnd.n4194 gnd.n4193 585
R3742 gnd.n3695 gnd.n3532 585
R3743 gnd.n3532 gnd.n3531 585
R3744 gnd.n3697 gnd.n3696 585
R3745 gnd.n4179 gnd.n3697 585
R3746 gnd.n3682 gnd.n3680 585
R3747 gnd.n4159 gnd.n3682 585
R3748 gnd.n4187 gnd.n4186 585
R3749 gnd.n4186 gnd.n4185 585
R3750 gnd.n3681 gnd.n3679 585
R3751 gnd.n4167 gnd.n3681 585
R3752 gnd.n4144 gnd.n3713 585
R3753 gnd.n3713 gnd.n3704 585
R3754 gnd.n4146 gnd.n4145 585
R3755 gnd.n4148 gnd.n4146 585
R3756 gnd.n3714 gnd.n3712 585
R3757 gnd.n3718 gnd.n3712 585
R3758 gnd.n4139 gnd.n4138 585
R3759 gnd.n4138 gnd.n4137 585
R3760 gnd.n3717 gnd.n3716 585
R3761 gnd.n3728 gnd.n3717 585
R3762 gnd.n4018 gnd.n3737 585
R3763 gnd.n4110 gnd.n3737 585
R3764 gnd.n4020 gnd.n4019 585
R3765 gnd.n4019 gnd.n3735 585
R3766 gnd.n4021 gnd.n3748 585
R3767 gnd.n4100 gnd.n3748 585
R3768 gnd.n4023 gnd.n4022 585
R3769 gnd.n4023 gnd.n3755 585
R3770 gnd.n4025 gnd.n4024 585
R3771 gnd.n4024 gnd.n3754 585
R3772 gnd.n4026 gnd.n3765 585
R3773 gnd.n4080 gnd.n3765 585
R3774 gnd.n4028 gnd.n4027 585
R3775 gnd.n4027 gnd.n3763 585
R3776 gnd.n4029 gnd.n3774 585
R3777 gnd.n4069 gnd.n3774 585
R3778 gnd.n4031 gnd.n4030 585
R3779 gnd.n4031 gnd.n3780 585
R3780 gnd.n4033 gnd.n4032 585
R3781 gnd.n4032 gnd.n3779 585
R3782 gnd.n4034 gnd.n3795 585
R3783 gnd.n4048 gnd.n3795 585
R3784 gnd.n4035 gnd.n3848 585
R3785 gnd.n3848 gnd.n3787 585
R3786 gnd.n4037 gnd.n4036 585
R3787 gnd.n4038 gnd.n4037 585
R3788 gnd.n3849 gnd.n3847 585
R3789 gnd.n3847 gnd.n3846 585
R3790 gnd.n4002 gnd.n4001 585
R3791 gnd.n4001 gnd.n4000 585
R3792 gnd.n3852 gnd.n3851 585
R3793 gnd.n3853 gnd.n3852 585
R3794 gnd.n3991 gnd.n3990 585
R3795 gnd.n3992 gnd.n3991 585
R3796 gnd.n3861 gnd.n3860 585
R3797 gnd.n3860 gnd.n3859 585
R3798 gnd.n3986 gnd.n3985 585
R3799 gnd.n3985 gnd.n3984 585
R3800 gnd.n3864 gnd.n3863 585
R3801 gnd.n3975 gnd.n3864 585
R3802 gnd.n3974 gnd.n3973 585
R3803 gnd.n3976 gnd.n3974 585
R3804 gnd.n3872 gnd.n3871 585
R3805 gnd.n3871 gnd.n3870 585
R3806 gnd.n4654 gnd.n2011 585
R3807 gnd.n2011 gnd.n1988 585
R3808 gnd.n4656 gnd.n4655 585
R3809 gnd.n4657 gnd.n4656 585
R3810 gnd.n3366 gnd.n3365 585
R3811 gnd.n3373 gnd.n3365 585
R3812 gnd.n4649 gnd.n4648 585
R3813 gnd.n4648 gnd.n4647 585
R3814 gnd.n3369 gnd.n3368 585
R3815 gnd.n4637 gnd.n3369 585
R3816 gnd.n4368 gnd.n3390 585
R3817 gnd.n3390 gnd.n3380 585
R3818 gnd.n4370 gnd.n4369 585
R3819 gnd.n4371 gnd.n4370 585
R3820 gnd.n3391 gnd.n3389 585
R3821 gnd.n3398 gnd.n3389 585
R3822 gnd.n4363 gnd.n4362 585
R3823 gnd.n4362 gnd.n4361 585
R3824 gnd.n3394 gnd.n3393 585
R3825 gnd.n4350 gnd.n3394 585
R3826 gnd.n4337 gnd.n3416 585
R3827 gnd.n3416 gnd.n3415 585
R3828 gnd.n4339 gnd.n4338 585
R3829 gnd.n4340 gnd.n4339 585
R3830 gnd.n3417 gnd.n3414 585
R3831 gnd.n3424 gnd.n3414 585
R3832 gnd.n4332 gnd.n4331 585
R3833 gnd.n4331 gnd.n4330 585
R3834 gnd.n3420 gnd.n3419 585
R3835 gnd.n4319 gnd.n3420 585
R3836 gnd.n4306 gnd.n3441 585
R3837 gnd.n3441 gnd.n3440 585
R3838 gnd.n4308 gnd.n4307 585
R3839 gnd.n4309 gnd.n4308 585
R3840 gnd.n3442 gnd.n3439 585
R3841 gnd.n3587 gnd.n3439 585
R3842 gnd.n4301 gnd.n4300 585
R3843 gnd.n4300 gnd.n4299 585
R3844 gnd.n3445 gnd.n3444 585
R3845 gnd.n4288 gnd.n3445 585
R3846 gnd.n4275 gnd.n3466 585
R3847 gnd.n3466 gnd.n3465 585
R3848 gnd.n4277 gnd.n4276 585
R3849 gnd.n4278 gnd.n4277 585
R3850 gnd.n3467 gnd.n3464 585
R3851 gnd.n3474 gnd.n3464 585
R3852 gnd.n4270 gnd.n4269 585
R3853 gnd.n4269 gnd.n4268 585
R3854 gnd.n3470 gnd.n3469 585
R3855 gnd.n4257 gnd.n3470 585
R3856 gnd.n4244 gnd.n3492 585
R3857 gnd.n3492 gnd.n3482 585
R3858 gnd.n4246 gnd.n4245 585
R3859 gnd.n4247 gnd.n4246 585
R3860 gnd.n3493 gnd.n3491 585
R3861 gnd.n3500 gnd.n3491 585
R3862 gnd.n4239 gnd.n4238 585
R3863 gnd.n4238 gnd.n4237 585
R3864 gnd.n3496 gnd.n3495 585
R3865 gnd.n4226 gnd.n3496 585
R3866 gnd.n4213 gnd.n3516 585
R3867 gnd.n3612 gnd.n3516 585
R3868 gnd.n4215 gnd.n4214 585
R3869 gnd.n4216 gnd.n4215 585
R3870 gnd.n3517 gnd.n3515 585
R3871 gnd.n3523 gnd.n3515 585
R3872 gnd.n4208 gnd.n4207 585
R3873 gnd.n4207 gnd.n4206 585
R3874 gnd.n3520 gnd.n3519 585
R3875 gnd.n4195 gnd.n3520 585
R3876 gnd.n4177 gnd.n4176 585
R3877 gnd.n4178 gnd.n4177 585
R3878 gnd.n3699 gnd.n3698 585
R3879 gnd.n4160 gnd.n3698 585
R3880 gnd.n4172 gnd.n4171 585
R3881 gnd.n4171 gnd.n3684 585
R3882 gnd.n4170 gnd.n3701 585
R3883 gnd.n4170 gnd.n3683 585
R3884 gnd.n4169 gnd.n3703 585
R3885 gnd.n4169 gnd.n4168 585
R3886 gnd.n4121 gnd.n3702 585
R3887 gnd.n4147 gnd.n3702 585
R3888 gnd.n4123 gnd.n4122 585
R3889 gnd.n4122 gnd.n3711 585
R3890 gnd.n4124 gnd.n3730 585
R3891 gnd.n3730 gnd.n3719 585
R3892 gnd.n4126 gnd.n4125 585
R3893 gnd.n4127 gnd.n4126 585
R3894 gnd.n3731 gnd.n3729 585
R3895 gnd.n3738 gnd.n3729 585
R3896 gnd.n4113 gnd.n4112 585
R3897 gnd.n4112 gnd.n4111 585
R3898 gnd.n3734 gnd.n3733 585
R3899 gnd.n4101 gnd.n3734 585
R3900 gnd.n4088 gnd.n3758 585
R3901 gnd.n3758 gnd.n3757 585
R3902 gnd.n4090 gnd.n4089 585
R3903 gnd.n4091 gnd.n4090 585
R3904 gnd.n3759 gnd.n3756 585
R3905 gnd.n3766 gnd.n3756 585
R3906 gnd.n4083 gnd.n4082 585
R3907 gnd.n4082 gnd.n4081 585
R3908 gnd.n3762 gnd.n3761 585
R3909 gnd.n4070 gnd.n3762 585
R3910 gnd.n4057 gnd.n3783 585
R3911 gnd.n3783 gnd.n3782 585
R3912 gnd.n4059 gnd.n4058 585
R3913 gnd.n4060 gnd.n4059 585
R3914 gnd.n4053 gnd.n3781 585
R3915 gnd.n4052 gnd.n4051 585
R3916 gnd.n3786 gnd.n3785 585
R3917 gnd.n4049 gnd.n3786 585
R3918 gnd.n3808 gnd.n3807 585
R3919 gnd.n3811 gnd.n3810 585
R3920 gnd.n3809 gnd.n3804 585
R3921 gnd.n3816 gnd.n3815 585
R3922 gnd.n3818 gnd.n3817 585
R3923 gnd.n3821 gnd.n3820 585
R3924 gnd.n3819 gnd.n3802 585
R3925 gnd.n3826 gnd.n3825 585
R3926 gnd.n3828 gnd.n3827 585
R3927 gnd.n3831 gnd.n3830 585
R3928 gnd.n3829 gnd.n3800 585
R3929 gnd.n3836 gnd.n3835 585
R3930 gnd.n3840 gnd.n3837 585
R3931 gnd.n3841 gnd.n3778 585
R3932 gnd.n3362 gnd.n2026 585
R3933 gnd.n4723 gnd.n4722 585
R3934 gnd.n4725 gnd.n4724 585
R3935 gnd.n4727 gnd.n4726 585
R3936 gnd.n4729 gnd.n4728 585
R3937 gnd.n4731 gnd.n4730 585
R3938 gnd.n4733 gnd.n4732 585
R3939 gnd.n4735 gnd.n4734 585
R3940 gnd.n4737 gnd.n4736 585
R3941 gnd.n4739 gnd.n4738 585
R3942 gnd.n4741 gnd.n4740 585
R3943 gnd.n4743 gnd.n4742 585
R3944 gnd.n4745 gnd.n4744 585
R3945 gnd.n4748 gnd.n4747 585
R3946 gnd.n4746 gnd.n2014 585
R3947 gnd.n4752 gnd.n2012 585
R3948 gnd.n4754 gnd.n4753 585
R3949 gnd.n4755 gnd.n4754 585
R3950 gnd.n3363 gnd.n3360 585
R3951 gnd.n3363 gnd.n1988 585
R3952 gnd.n4659 gnd.n4658 585
R3953 gnd.n4658 gnd.n4657 585
R3954 gnd.n3361 gnd.n3359 585
R3955 gnd.n3373 gnd.n3361 585
R3956 gnd.n4640 gnd.n3371 585
R3957 gnd.n4647 gnd.n3371 585
R3958 gnd.n4639 gnd.n4638 585
R3959 gnd.n4638 gnd.n4637 585
R3960 gnd.n3379 gnd.n3377 585
R3961 gnd.n3380 gnd.n3379 585
R3962 gnd.n4373 gnd.n4372 585
R3963 gnd.n4372 gnd.n4371 585
R3964 gnd.n3386 gnd.n3385 585
R3965 gnd.n3398 gnd.n3386 585
R3966 gnd.n4353 gnd.n3396 585
R3967 gnd.n4361 gnd.n3396 585
R3968 gnd.n4352 gnd.n4351 585
R3969 gnd.n4351 gnd.n4350 585
R3970 gnd.n3405 gnd.n3403 585
R3971 gnd.n3415 gnd.n3405 585
R3972 gnd.n4342 gnd.n4341 585
R3973 gnd.n4341 gnd.n4340 585
R3974 gnd.n3411 gnd.n3410 585
R3975 gnd.n3424 gnd.n3411 585
R3976 gnd.n4322 gnd.n3422 585
R3977 gnd.n4330 gnd.n3422 585
R3978 gnd.n4321 gnd.n4320 585
R3979 gnd.n4320 gnd.n4319 585
R3980 gnd.n3431 gnd.n3429 585
R3981 gnd.n3440 gnd.n3431 585
R3982 gnd.n4311 gnd.n4310 585
R3983 gnd.n4310 gnd.n4309 585
R3984 gnd.n3437 gnd.n3436 585
R3985 gnd.n3587 gnd.n3437 585
R3986 gnd.n4291 gnd.n3447 585
R3987 gnd.n4299 gnd.n3447 585
R3988 gnd.n4290 gnd.n4289 585
R3989 gnd.n4289 gnd.n4288 585
R3990 gnd.n3455 gnd.n3453 585
R3991 gnd.n3465 gnd.n3455 585
R3992 gnd.n4280 gnd.n4279 585
R3993 gnd.n4279 gnd.n4278 585
R3994 gnd.n3461 gnd.n3460 585
R3995 gnd.n3474 gnd.n3461 585
R3996 gnd.n4260 gnd.n3472 585
R3997 gnd.n4268 gnd.n3472 585
R3998 gnd.n4259 gnd.n4258 585
R3999 gnd.n4258 gnd.n4257 585
R4000 gnd.n3481 gnd.n3479 585
R4001 gnd.n3482 gnd.n3481 585
R4002 gnd.n4249 gnd.n4248 585
R4003 gnd.n4248 gnd.n4247 585
R4004 gnd.n3488 gnd.n3487 585
R4005 gnd.n3500 gnd.n3488 585
R4006 gnd.n4229 gnd.n3498 585
R4007 gnd.n4237 gnd.n3498 585
R4008 gnd.n4228 gnd.n4227 585
R4009 gnd.n4227 gnd.n4226 585
R4010 gnd.n3507 gnd.n3505 585
R4011 gnd.n3612 gnd.n3507 585
R4012 gnd.n4218 gnd.n4217 585
R4013 gnd.n4217 gnd.n4216 585
R4014 gnd.n3513 gnd.n3512 585
R4015 gnd.n3523 gnd.n3513 585
R4016 gnd.n4198 gnd.n3521 585
R4017 gnd.n4206 gnd.n3521 585
R4018 gnd.n4197 gnd.n4196 585
R4019 gnd.n4196 gnd.n4195 585
R4020 gnd.n3530 gnd.n3528 585
R4021 gnd.n4178 gnd.n3530 585
R4022 gnd.n4161 gnd.n4158 585
R4023 gnd.n4161 gnd.n4160 585
R4024 gnd.n4163 gnd.n4162 585
R4025 gnd.n4162 gnd.n3684 585
R4026 gnd.n4164 gnd.n3706 585
R4027 gnd.n3706 gnd.n3683 585
R4028 gnd.n4166 gnd.n4165 585
R4029 gnd.n4168 gnd.n4166 585
R4030 gnd.n3707 gnd.n3705 585
R4031 gnd.n4147 gnd.n3705 585
R4032 gnd.n4131 gnd.n4130 585
R4033 gnd.n4130 gnd.n3711 585
R4034 gnd.n4129 gnd.n3725 585
R4035 gnd.n4129 gnd.n3719 585
R4036 gnd.n4128 gnd.n3727 585
R4037 gnd.n4128 gnd.n4127 585
R4038 gnd.n4105 gnd.n3726 585
R4039 gnd.n3738 gnd.n3726 585
R4040 gnd.n4104 gnd.n3736 585
R4041 gnd.n4111 gnd.n3736 585
R4042 gnd.n4103 gnd.n4102 585
R4043 gnd.n4102 gnd.n4101 585
R4044 gnd.n3747 gnd.n3744 585
R4045 gnd.n3757 gnd.n3747 585
R4046 gnd.n4093 gnd.n4092 585
R4047 gnd.n4092 gnd.n4091 585
R4048 gnd.n3753 gnd.n3752 585
R4049 gnd.n3766 gnd.n3753 585
R4050 gnd.n4073 gnd.n3764 585
R4051 gnd.n4081 gnd.n3764 585
R4052 gnd.n4072 gnd.n4071 585
R4053 gnd.n4071 gnd.n4070 585
R4054 gnd.n3773 gnd.n3771 585
R4055 gnd.n3782 gnd.n3773 585
R4056 gnd.n4062 gnd.n4061 585
R4057 gnd.n4061 gnd.n4060 585
R4058 gnd.n5770 gnd.n5769 585
R4059 gnd.n5771 gnd.n5770 585
R4060 gnd.n1360 gnd.n1358 585
R4061 gnd.n5694 gnd.n1358 585
R4062 gnd.n5564 gnd.n1660 585
R4063 gnd.n5386 gnd.n1660 585
R4064 gnd.n5566 gnd.n5565 585
R4065 gnd.n5567 gnd.n5566 585
R4066 gnd.n1661 gnd.n1659 585
R4067 gnd.n5384 gnd.n1659 585
R4068 gnd.n5559 gnd.n5558 585
R4069 gnd.n5558 gnd.n5557 585
R4070 gnd.n1664 gnd.n1663 585
R4071 gnd.n5373 gnd.n1664 585
R4072 gnd.n5548 gnd.n5547 585
R4073 gnd.n5549 gnd.n5548 585
R4074 gnd.n1678 gnd.n1677 585
R4075 gnd.n5328 gnd.n1677 585
R4076 gnd.n5543 gnd.n5542 585
R4077 gnd.n5542 gnd.n5541 585
R4078 gnd.n1681 gnd.n1680 585
R4079 gnd.n5334 gnd.n1681 585
R4080 gnd.n5532 gnd.n5531 585
R4081 gnd.n5533 gnd.n5532 585
R4082 gnd.n1695 gnd.n1694 585
R4083 gnd.n5320 gnd.n1694 585
R4084 gnd.n5527 gnd.n5526 585
R4085 gnd.n5526 gnd.n5525 585
R4086 gnd.n1698 gnd.n1697 585
R4087 gnd.n5316 gnd.n1698 585
R4088 gnd.n5516 gnd.n5515 585
R4089 gnd.n5517 gnd.n5516 585
R4090 gnd.n1712 gnd.n1711 585
R4091 gnd.n5289 gnd.n1711 585
R4092 gnd.n5511 gnd.n5510 585
R4093 gnd.n5510 gnd.n5509 585
R4094 gnd.n1715 gnd.n1714 585
R4095 gnd.n5295 gnd.n1715 585
R4096 gnd.n5500 gnd.n5499 585
R4097 gnd.n5501 gnd.n5500 585
R4098 gnd.n1729 gnd.n1728 585
R4099 gnd.n5280 gnd.n1728 585
R4100 gnd.n5495 gnd.n5494 585
R4101 gnd.n5494 gnd.n5493 585
R4102 gnd.n1732 gnd.n1731 585
R4103 gnd.n5276 gnd.n1732 585
R4104 gnd.n5484 gnd.n5483 585
R4105 gnd.n5485 gnd.n5484 585
R4106 gnd.n1746 gnd.n1745 585
R4107 gnd.n5249 gnd.n1745 585
R4108 gnd.n5479 gnd.n5478 585
R4109 gnd.n5478 gnd.n5477 585
R4110 gnd.n1749 gnd.n1748 585
R4111 gnd.n5429 gnd.n1749 585
R4112 gnd.n5468 gnd.n5467 585
R4113 gnd.n5469 gnd.n5468 585
R4114 gnd.n1763 gnd.n1762 585
R4115 gnd.n5241 gnd.n1762 585
R4116 gnd.n5440 gnd.n5439 585
R4117 gnd.n5441 gnd.n5440 585
R4118 gnd.n5438 gnd.n1787 585
R4119 gnd.n5233 gnd.n1787 585
R4120 gnd.n5449 gnd.n5448 585
R4121 gnd.n5448 gnd.n5447 585
R4122 gnd.n5451 gnd.n5450 585
R4123 gnd.n5451 gnd.n1786 585
R4124 gnd.n5454 gnd.n5453 585
R4125 gnd.n5455 gnd.n5454 585
R4126 gnd.n5452 gnd.n1772 585
R4127 gnd.n1775 gnd.n1772 585
R4128 gnd.n5463 gnd.n5462 585
R4129 gnd.n5462 gnd.n5461 585
R4130 gnd.n5464 gnd.n1771 585
R4131 gnd.n5217 gnd.n1771 585
R4132 gnd.n1876 gnd.n1770 585
R4133 gnd.n1876 gnd.n1867 585
R4134 gnd.n5198 gnd.n5197 585
R4135 gnd.n5199 gnd.n5198 585
R4136 gnd.n5196 gnd.n1875 585
R4137 gnd.n5184 gnd.n1875 585
R4138 gnd.n1881 gnd.n1877 585
R4139 gnd.n1884 gnd.n1881 585
R4140 gnd.n5192 gnd.n5191 585
R4141 gnd.n5191 gnd.n5190 585
R4142 gnd.n1880 gnd.n1879 585
R4143 gnd.n5173 gnd.n1880 585
R4144 gnd.n5157 gnd.n1912 585
R4145 gnd.n1912 gnd.n1902 585
R4146 gnd.n5159 gnd.n5158 585
R4147 gnd.n5160 gnd.n5159 585
R4148 gnd.n1913 gnd.n1911 585
R4149 gnd.n1911 gnd.n1908 585
R4150 gnd.n5152 gnd.n5151 585
R4151 gnd.n5151 gnd.n5150 585
R4152 gnd.n1916 gnd.n1915 585
R4153 gnd.n1928 gnd.n1916 585
R4154 gnd.n5133 gnd.n5132 585
R4155 gnd.n5134 gnd.n5133 585
R4156 gnd.n1930 gnd.n1929 585
R4157 gnd.n1929 gnd.n1925 585
R4158 gnd.n5128 gnd.n5127 585
R4159 gnd.n5127 gnd.n5126 585
R4160 gnd.n1933 gnd.n1932 585
R4161 gnd.n1934 gnd.n1933 585
R4162 gnd.n5117 gnd.n5116 585
R4163 gnd.n5118 gnd.n5117 585
R4164 gnd.n1946 gnd.n1945 585
R4165 gnd.n1945 gnd.n1942 585
R4166 gnd.n5112 gnd.n5111 585
R4167 gnd.n5111 gnd.n5110 585
R4168 gnd.n1949 gnd.n1948 585
R4169 gnd.n1960 gnd.n1949 585
R4170 gnd.n5101 gnd.n5100 585
R4171 gnd.n5102 gnd.n5101 585
R4172 gnd.n1962 gnd.n1961 585
R4173 gnd.n1961 gnd.n1957 585
R4174 gnd.n5096 gnd.n5095 585
R4175 gnd.n5095 gnd.n5094 585
R4176 gnd.n1965 gnd.n1964 585
R4177 gnd.n1966 gnd.n1965 585
R4178 gnd.n5085 gnd.n5084 585
R4179 gnd.n5086 gnd.n5085 585
R4180 gnd.n1978 gnd.n1977 585
R4181 gnd.n1977 gnd.n1974 585
R4182 gnd.n5080 gnd.n5079 585
R4183 gnd.n5079 gnd.n5078 585
R4184 gnd.n1981 gnd.n1980 585
R4185 gnd.n4872 gnd.n1981 585
R4186 gnd.n5069 gnd.n5068 585
R4187 gnd.n5070 gnd.n5069 585
R4188 gnd.n5065 gnd.n4873 585
R4189 gnd.n5064 gnd.n5063 585
R4190 gnd.n5061 gnd.n4875 585
R4191 gnd.n5061 gnd.n4756 585
R4192 gnd.n5060 gnd.n5059 585
R4193 gnd.n5058 gnd.n5057 585
R4194 gnd.n5056 gnd.n4880 585
R4195 gnd.n5054 gnd.n5053 585
R4196 gnd.n5052 gnd.n4881 585
R4197 gnd.n5051 gnd.n5050 585
R4198 gnd.n5048 gnd.n4886 585
R4199 gnd.n5046 gnd.n5045 585
R4200 gnd.n5044 gnd.n4887 585
R4201 gnd.n5043 gnd.n5042 585
R4202 gnd.n5040 gnd.n4892 585
R4203 gnd.n5038 gnd.n5037 585
R4204 gnd.n5036 gnd.n4893 585
R4205 gnd.n5035 gnd.n5034 585
R4206 gnd.n5032 gnd.n4898 585
R4207 gnd.n5030 gnd.n5029 585
R4208 gnd.n5028 gnd.n4899 585
R4209 gnd.n5027 gnd.n5026 585
R4210 gnd.n5024 gnd.n4907 585
R4211 gnd.n5022 gnd.n5021 585
R4212 gnd.n5020 gnd.n4908 585
R4213 gnd.n5019 gnd.n5018 585
R4214 gnd.n5016 gnd.n4913 585
R4215 gnd.n5014 gnd.n5013 585
R4216 gnd.n5012 gnd.n4914 585
R4217 gnd.n5011 gnd.n5010 585
R4218 gnd.n5008 gnd.n4919 585
R4219 gnd.n5006 gnd.n5005 585
R4220 gnd.n5004 gnd.n4920 585
R4221 gnd.n5003 gnd.n5002 585
R4222 gnd.n5000 gnd.n4925 585
R4223 gnd.n4998 gnd.n4997 585
R4224 gnd.n4996 gnd.n4926 585
R4225 gnd.n4995 gnd.n4931 585
R4226 gnd.n4988 gnd.n4934 585
R4227 gnd.n4991 gnd.n4990 585
R4228 gnd.n5701 gnd.n5700 585
R4229 gnd.n5703 gnd.n1643 585
R4230 gnd.n5705 gnd.n5704 585
R4231 gnd.n5706 gnd.n1636 585
R4232 gnd.n5708 gnd.n5707 585
R4233 gnd.n5710 gnd.n1634 585
R4234 gnd.n5712 gnd.n5711 585
R4235 gnd.n5713 gnd.n1629 585
R4236 gnd.n5715 gnd.n5714 585
R4237 gnd.n5717 gnd.n1627 585
R4238 gnd.n5719 gnd.n5718 585
R4239 gnd.n5720 gnd.n1622 585
R4240 gnd.n5722 gnd.n5721 585
R4241 gnd.n5724 gnd.n1620 585
R4242 gnd.n5726 gnd.n5725 585
R4243 gnd.n5727 gnd.n1615 585
R4244 gnd.n5729 gnd.n5728 585
R4245 gnd.n5731 gnd.n1613 585
R4246 gnd.n5733 gnd.n5732 585
R4247 gnd.n5734 gnd.n1607 585
R4248 gnd.n5736 gnd.n5735 585
R4249 gnd.n5740 gnd.n1386 585
R4250 gnd.n5742 gnd.n5741 585
R4251 gnd.n5743 gnd.n1381 585
R4252 gnd.n5745 gnd.n5744 585
R4253 gnd.n5747 gnd.n1379 585
R4254 gnd.n5749 gnd.n5748 585
R4255 gnd.n5750 gnd.n1374 585
R4256 gnd.n5752 gnd.n5751 585
R4257 gnd.n5754 gnd.n1372 585
R4258 gnd.n5756 gnd.n5755 585
R4259 gnd.n5757 gnd.n1366 585
R4260 gnd.n5759 gnd.n5758 585
R4261 gnd.n5761 gnd.n1365 585
R4262 gnd.n5762 gnd.n1363 585
R4263 gnd.n5765 gnd.n5764 585
R4264 gnd.n5766 gnd.n1359 585
R4265 gnd.n1364 gnd.n1359 585
R4266 gnd.n5697 gnd.n1355 585
R4267 gnd.n5771 gnd.n1355 585
R4268 gnd.n5696 gnd.n5695 585
R4269 gnd.n5695 gnd.n5694 585
R4270 gnd.n1648 gnd.n1647 585
R4271 gnd.n5386 gnd.n1648 585
R4272 gnd.n5381 gnd.n1656 585
R4273 gnd.n5567 gnd.n1656 585
R4274 gnd.n5383 gnd.n5382 585
R4275 gnd.n5384 gnd.n5383 585
R4276 gnd.n1831 gnd.n1666 585
R4277 gnd.n5557 gnd.n1666 585
R4278 gnd.n5375 gnd.n5374 585
R4279 gnd.n5374 gnd.n5373 585
R4280 gnd.n1833 gnd.n1675 585
R4281 gnd.n5549 gnd.n1675 585
R4282 gnd.n5330 gnd.n5329 585
R4283 gnd.n5329 gnd.n5328 585
R4284 gnd.n5331 gnd.n1682 585
R4285 gnd.n5541 gnd.n1682 585
R4286 gnd.n5333 gnd.n5332 585
R4287 gnd.n5334 gnd.n5333 585
R4288 gnd.n1840 gnd.n1691 585
R4289 gnd.n5533 gnd.n1691 585
R4290 gnd.n5322 gnd.n5321 585
R4291 gnd.n5321 gnd.n5320 585
R4292 gnd.n5319 gnd.n1700 585
R4293 gnd.n5525 gnd.n1700 585
R4294 gnd.n5318 gnd.n5317 585
R4295 gnd.n5317 gnd.n5316 585
R4296 gnd.n1842 gnd.n1709 585
R4297 gnd.n5517 gnd.n1709 585
R4298 gnd.n5291 gnd.n5290 585
R4299 gnd.n5290 gnd.n5289 585
R4300 gnd.n5292 gnd.n1716 585
R4301 gnd.n5509 gnd.n1716 585
R4302 gnd.n5294 gnd.n5293 585
R4303 gnd.n5295 gnd.n5294 585
R4304 gnd.n1850 gnd.n1725 585
R4305 gnd.n5501 gnd.n1725 585
R4306 gnd.n5282 gnd.n5281 585
R4307 gnd.n5281 gnd.n5280 585
R4308 gnd.n5279 gnd.n1734 585
R4309 gnd.n5493 gnd.n1734 585
R4310 gnd.n5278 gnd.n5277 585
R4311 gnd.n5277 gnd.n5276 585
R4312 gnd.n1852 gnd.n1743 585
R4313 gnd.n5485 gnd.n1743 585
R4314 gnd.n5251 gnd.n5250 585
R4315 gnd.n5250 gnd.n5249 585
R4316 gnd.n5248 gnd.n1750 585
R4317 gnd.n5477 gnd.n1750 585
R4318 gnd.n5247 gnd.n1806 585
R4319 gnd.n5429 gnd.n1806 585
R4320 gnd.n1854 gnd.n1759 585
R4321 gnd.n5469 gnd.n1759 585
R4322 gnd.n5243 gnd.n5242 585
R4323 gnd.n5242 gnd.n5241 585
R4324 gnd.n1856 gnd.n1796 585
R4325 gnd.n5441 gnd.n1796 585
R4326 gnd.n5232 gnd.n5231 585
R4327 gnd.n5233 gnd.n5232 585
R4328 gnd.n1860 gnd.n1789 585
R4329 gnd.n5447 gnd.n1789 585
R4330 gnd.n5227 gnd.n5226 585
R4331 gnd.n5226 gnd.n1786 585
R4332 gnd.n5225 gnd.n1784 585
R4333 gnd.n5455 gnd.n1784 585
R4334 gnd.n5224 gnd.n5223 585
R4335 gnd.n5223 gnd.n1775 585
R4336 gnd.n1863 gnd.n1773 585
R4337 gnd.n5461 gnd.n1773 585
R4338 gnd.n5219 gnd.n5218 585
R4339 gnd.n5218 gnd.n5217 585
R4340 gnd.n1866 gnd.n1865 585
R4341 gnd.n1867 gnd.n1866 585
R4342 gnd.n5181 gnd.n1873 585
R4343 gnd.n5199 gnd.n1873 585
R4344 gnd.n5183 gnd.n5182 585
R4345 gnd.n5184 gnd.n5183 585
R4346 gnd.n1898 gnd.n1897 585
R4347 gnd.n1897 gnd.n1884 585
R4348 gnd.n5176 gnd.n1882 585
R4349 gnd.n5190 gnd.n1882 585
R4350 gnd.n5175 gnd.n5174 585
R4351 gnd.n5174 gnd.n5173 585
R4352 gnd.n1901 gnd.n1900 585
R4353 gnd.n1902 gnd.n1901 585
R4354 gnd.n4957 gnd.n1909 585
R4355 gnd.n5160 gnd.n1909 585
R4356 gnd.n4959 gnd.n4958 585
R4357 gnd.n4958 gnd.n1908 585
R4358 gnd.n4960 gnd.n1917 585
R4359 gnd.n5150 gnd.n1917 585
R4360 gnd.n4962 gnd.n4961 585
R4361 gnd.n4961 gnd.n1928 585
R4362 gnd.n4963 gnd.n1926 585
R4363 gnd.n5134 gnd.n1926 585
R4364 gnd.n4965 gnd.n4964 585
R4365 gnd.n4964 gnd.n1925 585
R4366 gnd.n4966 gnd.n1935 585
R4367 gnd.n5126 gnd.n1935 585
R4368 gnd.n4968 gnd.n4967 585
R4369 gnd.n4967 gnd.n1934 585
R4370 gnd.n4969 gnd.n1943 585
R4371 gnd.n5118 gnd.n1943 585
R4372 gnd.n4971 gnd.n4970 585
R4373 gnd.n4970 gnd.n1942 585
R4374 gnd.n4972 gnd.n1950 585
R4375 gnd.n5110 gnd.n1950 585
R4376 gnd.n4974 gnd.n4973 585
R4377 gnd.n4973 gnd.n1960 585
R4378 gnd.n4975 gnd.n1958 585
R4379 gnd.n5102 gnd.n1958 585
R4380 gnd.n4977 gnd.n4976 585
R4381 gnd.n4976 gnd.n1957 585
R4382 gnd.n4978 gnd.n1967 585
R4383 gnd.n5094 gnd.n1967 585
R4384 gnd.n4980 gnd.n4979 585
R4385 gnd.n4979 gnd.n1966 585
R4386 gnd.n4981 gnd.n1975 585
R4387 gnd.n5086 gnd.n1975 585
R4388 gnd.n4983 gnd.n4982 585
R4389 gnd.n4982 gnd.n1974 585
R4390 gnd.n4984 gnd.n1982 585
R4391 gnd.n5078 gnd.n1982 585
R4392 gnd.n4985 gnd.n4936 585
R4393 gnd.n4936 gnd.n4872 585
R4394 gnd.n4986 gnd.n4757 585
R4395 gnd.n5070 gnd.n4757 585
R4396 gnd.n7572 gnd.n7571 585
R4397 gnd.n7573 gnd.n7572 585
R4398 gnd.n128 gnd.n126 585
R4399 gnd.n126 gnd.n122 585
R4400 gnd.n7492 gnd.n7491 585
R4401 gnd.n7493 gnd.n7492 585
R4402 gnd.n205 gnd.n204 585
R4403 gnd.n204 gnd.n202 585
R4404 gnd.n7487 gnd.n7486 585
R4405 gnd.n7486 gnd.n7485 585
R4406 gnd.n208 gnd.n207 585
R4407 gnd.n209 gnd.n208 585
R4408 gnd.n7408 gnd.n7407 585
R4409 gnd.n7409 gnd.n7408 585
R4410 gnd.n221 gnd.n220 585
R4411 gnd.n228 gnd.n220 585
R4412 gnd.n7403 gnd.n7402 585
R4413 gnd.n7402 gnd.n7401 585
R4414 gnd.n224 gnd.n223 585
R4415 gnd.n225 gnd.n224 585
R4416 gnd.n7392 gnd.n7391 585
R4417 gnd.n7393 gnd.n7392 585
R4418 gnd.n238 gnd.n237 585
R4419 gnd.n237 gnd.n234 585
R4420 gnd.n7387 gnd.n7386 585
R4421 gnd.n7386 gnd.n7385 585
R4422 gnd.n241 gnd.n240 585
R4423 gnd.n250 gnd.n241 585
R4424 gnd.n7376 gnd.n7375 585
R4425 gnd.n7377 gnd.n7376 585
R4426 gnd.n252 gnd.n251 585
R4427 gnd.n259 gnd.n251 585
R4428 gnd.n7371 gnd.n7370 585
R4429 gnd.n7370 gnd.n7369 585
R4430 gnd.n255 gnd.n254 585
R4431 gnd.n256 gnd.n255 585
R4432 gnd.n7360 gnd.n7359 585
R4433 gnd.n7361 gnd.n7360 585
R4434 gnd.n268 gnd.n267 585
R4435 gnd.n267 gnd.n265 585
R4436 gnd.n7355 gnd.n7354 585
R4437 gnd.n7354 gnd.n7353 585
R4438 gnd.n271 gnd.n270 585
R4439 gnd.n280 gnd.n271 585
R4440 gnd.n7344 gnd.n7343 585
R4441 gnd.n7345 gnd.n7344 585
R4442 gnd.n282 gnd.n281 585
R4443 gnd.n289 gnd.n281 585
R4444 gnd.n7339 gnd.n7338 585
R4445 gnd.n7338 gnd.n7337 585
R4446 gnd.n285 gnd.n284 585
R4447 gnd.n286 gnd.n285 585
R4448 gnd.n7328 gnd.n7327 585
R4449 gnd.n7329 gnd.n7328 585
R4450 gnd.n298 gnd.n297 585
R4451 gnd.n297 gnd.n295 585
R4452 gnd.n7304 gnd.n7303 585
R4453 gnd.n7305 gnd.n7304 585
R4454 gnd.n7302 gnd.n328 585
R4455 gnd.n7302 gnd.n7301 585
R4456 gnd.n327 gnd.n326 585
R4457 gnd.n330 gnd.n326 585
R4458 gnd.n7227 gnd.n7226 585
R4459 gnd.n7228 gnd.n7227 585
R4460 gnd.n7225 gnd.n7224 585
R4461 gnd.n7224 gnd.n336 585
R4462 gnd.n7223 gnd.n338 585
R4463 gnd.n7223 gnd.n7222 585
R4464 gnd.n337 gnd.n307 585
R4465 gnd.n7202 gnd.n307 585
R4466 gnd.n7322 gnd.n7321 585
R4467 gnd.n7321 gnd.n7320 585
R4468 gnd.n7323 gnd.n306 585
R4469 gnd.n7211 gnd.n306 585
R4470 gnd.n364 gnd.n305 585
R4471 gnd.n364 gnd.n349 585
R4472 gnd.n7189 gnd.n7188 585
R4473 gnd.n7190 gnd.n7189 585
R4474 gnd.n7187 gnd.n363 585
R4475 gnd.n7169 gnd.n363 585
R4476 gnd.n369 gnd.n365 585
R4477 gnd.n6930 gnd.n369 585
R4478 gnd.n7183 gnd.n7182 585
R4479 gnd.n7182 gnd.n7181 585
R4480 gnd.n368 gnd.n367 585
R4481 gnd.n7159 gnd.n368 585
R4482 gnd.n7137 gnd.n7136 585
R4483 gnd.n7138 gnd.n7137 585
R4484 gnd.n397 gnd.n396 585
R4485 gnd.n6938 gnd.n396 585
R4486 gnd.n7132 gnd.n7131 585
R4487 gnd.n7131 gnd.n7130 585
R4488 gnd.n400 gnd.n399 585
R4489 gnd.n6917 gnd.n400 585
R4490 gnd.n7118 gnd.n7117 585
R4491 gnd.n7119 gnd.n7118 585
R4492 gnd.n416 gnd.n415 585
R4493 gnd.n6898 gnd.n415 585
R4494 gnd.n7113 gnd.n7112 585
R4495 gnd.n7112 gnd.n7111 585
R4496 gnd.n419 gnd.n418 585
R4497 gnd.n6904 gnd.n419 585
R4498 gnd.n7102 gnd.n7101 585
R4499 gnd.n7103 gnd.n7102 585
R4500 gnd.n433 gnd.n432 585
R4501 gnd.n6890 gnd.n432 585
R4502 gnd.n7097 gnd.n7096 585
R4503 gnd.n7096 gnd.n7095 585
R4504 gnd.n436 gnd.n435 585
R4505 gnd.n6886 gnd.n436 585
R4506 gnd.n7086 gnd.n7085 585
R4507 gnd.n7087 gnd.n7086 585
R4508 gnd.n450 gnd.n449 585
R4509 gnd.n6859 gnd.n449 585
R4510 gnd.n7081 gnd.n7080 585
R4511 gnd.n7080 gnd.n7079 585
R4512 gnd.n453 gnd.n452 585
R4513 gnd.n6865 gnd.n453 585
R4514 gnd.n7070 gnd.n7069 585
R4515 gnd.n7071 gnd.n7070 585
R4516 gnd.n467 gnd.n466 585
R4517 gnd.n6850 gnd.n466 585
R4518 gnd.n7065 gnd.n7064 585
R4519 gnd.n7064 gnd.n7063 585
R4520 gnd.n470 gnd.n469 585
R4521 gnd.n6846 gnd.n470 585
R4522 gnd.n7054 gnd.n7053 585
R4523 gnd.n7055 gnd.n7054 585
R4524 gnd.n485 gnd.n484 585
R4525 gnd.n6974 gnd.n484 585
R4526 gnd.n7049 gnd.n7048 585
R4527 gnd.n488 gnd.n487 585
R4528 gnd.n7045 gnd.n7044 585
R4529 gnd.n7046 gnd.n7045 585
R4530 gnd.n7043 gnd.n519 585
R4531 gnd.n7042 gnd.n7041 585
R4532 gnd.n7040 gnd.n7039 585
R4533 gnd.n7038 gnd.n7037 585
R4534 gnd.n7036 gnd.n7035 585
R4535 gnd.n7034 gnd.n7033 585
R4536 gnd.n7032 gnd.n7031 585
R4537 gnd.n7030 gnd.n7029 585
R4538 gnd.n7028 gnd.n7027 585
R4539 gnd.n7026 gnd.n7025 585
R4540 gnd.n7024 gnd.n7023 585
R4541 gnd.n7022 gnd.n7021 585
R4542 gnd.n7020 gnd.n7019 585
R4543 gnd.n7017 gnd.n7016 585
R4544 gnd.n7015 gnd.n7014 585
R4545 gnd.n7013 gnd.n7012 585
R4546 gnd.n7011 gnd.n7010 585
R4547 gnd.n7009 gnd.n7008 585
R4548 gnd.n7007 gnd.n7006 585
R4549 gnd.n7005 gnd.n7004 585
R4550 gnd.n7003 gnd.n7002 585
R4551 gnd.n7001 gnd.n7000 585
R4552 gnd.n6999 gnd.n6998 585
R4553 gnd.n6997 gnd.n6996 585
R4554 gnd.n6995 gnd.n6994 585
R4555 gnd.n6993 gnd.n6992 585
R4556 gnd.n6991 gnd.n6990 585
R4557 gnd.n6989 gnd.n6988 585
R4558 gnd.n6987 gnd.n6986 585
R4559 gnd.n6985 gnd.n6984 585
R4560 gnd.n6983 gnd.n6982 585
R4561 gnd.n6981 gnd.n557 585
R4562 gnd.n561 gnd.n558 585
R4563 gnd.n6977 gnd.n6976 585
R4564 gnd.n196 gnd.n195 585
R4565 gnd.n7501 gnd.n191 585
R4566 gnd.n7503 gnd.n7502 585
R4567 gnd.n7505 gnd.n189 585
R4568 gnd.n7507 gnd.n7506 585
R4569 gnd.n7508 gnd.n184 585
R4570 gnd.n7510 gnd.n7509 585
R4571 gnd.n7512 gnd.n182 585
R4572 gnd.n7514 gnd.n7513 585
R4573 gnd.n7515 gnd.n177 585
R4574 gnd.n7517 gnd.n7516 585
R4575 gnd.n7519 gnd.n175 585
R4576 gnd.n7521 gnd.n7520 585
R4577 gnd.n7522 gnd.n170 585
R4578 gnd.n7524 gnd.n7523 585
R4579 gnd.n7526 gnd.n168 585
R4580 gnd.n7528 gnd.n7527 585
R4581 gnd.n7529 gnd.n163 585
R4582 gnd.n7531 gnd.n7530 585
R4583 gnd.n7533 gnd.n161 585
R4584 gnd.n7535 gnd.n7534 585
R4585 gnd.n7539 gnd.n156 585
R4586 gnd.n7541 gnd.n7540 585
R4587 gnd.n7543 gnd.n154 585
R4588 gnd.n7545 gnd.n7544 585
R4589 gnd.n7546 gnd.n149 585
R4590 gnd.n7548 gnd.n7547 585
R4591 gnd.n7550 gnd.n147 585
R4592 gnd.n7552 gnd.n7551 585
R4593 gnd.n7553 gnd.n142 585
R4594 gnd.n7555 gnd.n7554 585
R4595 gnd.n7557 gnd.n140 585
R4596 gnd.n7559 gnd.n7558 585
R4597 gnd.n7560 gnd.n135 585
R4598 gnd.n7562 gnd.n7561 585
R4599 gnd.n7564 gnd.n133 585
R4600 gnd.n7566 gnd.n7565 585
R4601 gnd.n7567 gnd.n131 585
R4602 gnd.n7568 gnd.n127 585
R4603 gnd.n127 gnd.n124 585
R4604 gnd.n7497 gnd.n123 585
R4605 gnd.n7573 gnd.n123 585
R4606 gnd.n7496 gnd.n7495 585
R4607 gnd.n7495 gnd.n122 585
R4608 gnd.n7494 gnd.n200 585
R4609 gnd.n7494 gnd.n7493 585
R4610 gnd.n7261 gnd.n201 585
R4611 gnd.n202 gnd.n201 585
R4612 gnd.n7262 gnd.n210 585
R4613 gnd.n7485 gnd.n210 585
R4614 gnd.n7264 gnd.n7263 585
R4615 gnd.n7263 gnd.n209 585
R4616 gnd.n7265 gnd.n219 585
R4617 gnd.n7409 gnd.n219 585
R4618 gnd.n7267 gnd.n7266 585
R4619 gnd.n7266 gnd.n228 585
R4620 gnd.n7268 gnd.n226 585
R4621 gnd.n7401 gnd.n226 585
R4622 gnd.n7270 gnd.n7269 585
R4623 gnd.n7269 gnd.n225 585
R4624 gnd.n7271 gnd.n235 585
R4625 gnd.n7393 gnd.n235 585
R4626 gnd.n7273 gnd.n7272 585
R4627 gnd.n7272 gnd.n234 585
R4628 gnd.n7274 gnd.n242 585
R4629 gnd.n7385 gnd.n242 585
R4630 gnd.n7276 gnd.n7275 585
R4631 gnd.n7275 gnd.n250 585
R4632 gnd.n7277 gnd.n249 585
R4633 gnd.n7377 gnd.n249 585
R4634 gnd.n7279 gnd.n7278 585
R4635 gnd.n7278 gnd.n259 585
R4636 gnd.n7280 gnd.n257 585
R4637 gnd.n7369 gnd.n257 585
R4638 gnd.n7282 gnd.n7281 585
R4639 gnd.n7281 gnd.n256 585
R4640 gnd.n7283 gnd.n266 585
R4641 gnd.n7361 gnd.n266 585
R4642 gnd.n7285 gnd.n7284 585
R4643 gnd.n7284 gnd.n265 585
R4644 gnd.n7286 gnd.n272 585
R4645 gnd.n7353 gnd.n272 585
R4646 gnd.n7288 gnd.n7287 585
R4647 gnd.n7287 gnd.n280 585
R4648 gnd.n7289 gnd.n279 585
R4649 gnd.n7345 gnd.n279 585
R4650 gnd.n7291 gnd.n7290 585
R4651 gnd.n7290 gnd.n289 585
R4652 gnd.n7292 gnd.n287 585
R4653 gnd.n7337 gnd.n287 585
R4654 gnd.n7294 gnd.n7293 585
R4655 gnd.n7293 gnd.n286 585
R4656 gnd.n7295 gnd.n296 585
R4657 gnd.n7329 gnd.n296 585
R4658 gnd.n7297 gnd.n7296 585
R4659 gnd.n7296 gnd.n295 585
R4660 gnd.n7298 gnd.n324 585
R4661 gnd.n7305 gnd.n324 585
R4662 gnd.n7300 gnd.n7299 585
R4663 gnd.n7301 gnd.n7300 585
R4664 gnd.n332 gnd.n331 585
R4665 gnd.n331 gnd.n330 585
R4666 gnd.n7230 gnd.n7229 585
R4667 gnd.n7229 gnd.n7228 585
R4668 gnd.n335 gnd.n334 585
R4669 gnd.n336 gnd.n335 585
R4670 gnd.n7199 gnd.n339 585
R4671 gnd.n7222 gnd.n339 585
R4672 gnd.n7201 gnd.n7200 585
R4673 gnd.n7202 gnd.n7201 585
R4674 gnd.n355 gnd.n309 585
R4675 gnd.n7320 gnd.n309 585
R4676 gnd.n7194 gnd.n350 585
R4677 gnd.n7211 gnd.n350 585
R4678 gnd.n7193 gnd.n7192 585
R4679 gnd.n7192 gnd.n349 585
R4680 gnd.n7191 gnd.n357 585
R4681 gnd.n7191 gnd.n7190 585
R4682 gnd.n6929 gnd.n358 585
R4683 gnd.n7169 gnd.n358 585
R4684 gnd.n6932 gnd.n6931 585
R4685 gnd.n6931 gnd.n6930 585
R4686 gnd.n6933 gnd.n370 585
R4687 gnd.n7181 gnd.n370 585
R4688 gnd.n6934 gnd.n387 585
R4689 gnd.n7159 gnd.n387 585
R4690 gnd.n6935 gnd.n394 585
R4691 gnd.n7138 gnd.n394 585
R4692 gnd.n6937 gnd.n6936 585
R4693 gnd.n6938 gnd.n6937 585
R4694 gnd.n585 gnd.n402 585
R4695 gnd.n7130 gnd.n402 585
R4696 gnd.n6919 gnd.n6918 585
R4697 gnd.n6918 gnd.n6917 585
R4698 gnd.n587 gnd.n413 585
R4699 gnd.n7119 gnd.n413 585
R4700 gnd.n6900 gnd.n6899 585
R4701 gnd.n6899 gnd.n6898 585
R4702 gnd.n6901 gnd.n420 585
R4703 gnd.n7111 gnd.n420 585
R4704 gnd.n6903 gnd.n6902 585
R4705 gnd.n6904 gnd.n6903 585
R4706 gnd.n594 gnd.n429 585
R4707 gnd.n7103 gnd.n429 585
R4708 gnd.n6892 gnd.n6891 585
R4709 gnd.n6891 gnd.n6890 585
R4710 gnd.n6889 gnd.n438 585
R4711 gnd.n7095 gnd.n438 585
R4712 gnd.n6888 gnd.n6887 585
R4713 gnd.n6887 gnd.n6886 585
R4714 gnd.n596 gnd.n447 585
R4715 gnd.n7087 gnd.n447 585
R4716 gnd.n6861 gnd.n6860 585
R4717 gnd.n6860 gnd.n6859 585
R4718 gnd.n6862 gnd.n454 585
R4719 gnd.n7079 gnd.n454 585
R4720 gnd.n6864 gnd.n6863 585
R4721 gnd.n6865 gnd.n6864 585
R4722 gnd.n6841 gnd.n463 585
R4723 gnd.n7071 gnd.n463 585
R4724 gnd.n6852 gnd.n6851 585
R4725 gnd.n6851 gnd.n6850 585
R4726 gnd.n6849 gnd.n472 585
R4727 gnd.n7063 gnd.n472 585
R4728 gnd.n6848 gnd.n6847 585
R4729 gnd.n6847 gnd.n6846 585
R4730 gnd.n6843 gnd.n481 585
R4731 gnd.n7055 gnd.n481 585
R4732 gnd.n6975 gnd.n563 585
R4733 gnd.n6975 gnd.n6974 585
R4734 gnd.n675 gnd.n674 585
R4735 gnd.n675 gnd.n646 585
R4736 gnd.n6771 gnd.n6770 585
R4737 gnd.n6770 gnd.n6769 585
R4738 gnd.n6772 gnd.n672 585
R4739 gnd.n672 gnd.n655 585
R4740 gnd.n6774 gnd.n6773 585
R4741 gnd.n6775 gnd.n6774 585
R4742 gnd.n673 gnd.n671 585
R4743 gnd.n671 gnd.n670 585
R4744 gnd.n6573 gnd.n661 585
R4745 gnd.n6781 gnd.n661 585
R4746 gnd.n6575 gnd.n6574 585
R4747 gnd.n6576 gnd.n6575 585
R4748 gnd.n6572 gnd.n899 585
R4749 gnd.n899 gnd.n898 585
R4750 gnd.n6571 gnd.n6570 585
R4751 gnd.n6570 gnd.n6569 585
R4752 gnd.n901 gnd.n900 585
R4753 gnd.n901 gnd.n880 585
R4754 gnd.n6557 gnd.n908 585
R4755 gnd.n908 gnd.n879 585
R4756 gnd.n6559 gnd.n6558 585
R4757 gnd.n6560 gnd.n6559 585
R4758 gnd.n6556 gnd.n907 585
R4759 gnd.n907 gnd.n890 585
R4760 gnd.n6555 gnd.n6554 585
R4761 gnd.n6554 gnd.n888 585
R4762 gnd.n6553 gnd.n909 585
R4763 gnd.n6553 gnd.n6552 585
R4764 gnd.n6227 gnd.n910 585
R4765 gnd.n911 gnd.n910 585
R4766 gnd.n6228 gnd.n6226 585
R4767 gnd.n6226 gnd.n920 585
R4768 gnd.n6230 gnd.n6229 585
R4769 gnd.n6230 gnd.n919 585
R4770 gnd.n6231 gnd.n6225 585
R4771 gnd.n6372 gnd.n6231 585
R4772 gnd.n6376 gnd.n6375 585
R4773 gnd.n6375 gnd.n6374 585
R4774 gnd.n6377 gnd.n6223 585
R4775 gnd.n6223 gnd.n928 585
R4776 gnd.n6379 gnd.n6378 585
R4777 gnd.n6380 gnd.n6379 585
R4778 gnd.n6224 gnd.n6222 585
R4779 gnd.n6222 gnd.n939 585
R4780 gnd.n6349 gnd.n6239 585
R4781 gnd.n6239 gnd.n937 585
R4782 gnd.n6351 gnd.n6350 585
R4783 gnd.n6352 gnd.n6351 585
R4784 gnd.n6348 gnd.n6238 585
R4785 gnd.n6238 gnd.n947 585
R4786 gnd.n6347 gnd.n6346 585
R4787 gnd.n6346 gnd.n945 585
R4788 gnd.n6345 gnd.n6240 585
R4789 gnd.n6345 gnd.n6344 585
R4790 gnd.n6331 gnd.n6241 585
R4791 gnd.n6241 gnd.n955 585
R4792 gnd.n6332 gnd.n6249 585
R4793 gnd.n6249 gnd.n953 585
R4794 gnd.n6334 gnd.n6333 585
R4795 gnd.n6335 gnd.n6334 585
R4796 gnd.n6330 gnd.n6248 585
R4797 gnd.n6248 gnd.n6247 585
R4798 gnd.n6329 gnd.n6328 585
R4799 gnd.n6328 gnd.n961 585
R4800 gnd.n6327 gnd.n6250 585
R4801 gnd.n6327 gnd.n6326 585
R4802 gnd.n6312 gnd.n6251 585
R4803 gnd.n6251 gnd.n970 585
R4804 gnd.n6313 gnd.n6259 585
R4805 gnd.n6259 gnd.n968 585
R4806 gnd.n6315 gnd.n6314 585
R4807 gnd.n6316 gnd.n6315 585
R4808 gnd.n6311 gnd.n6258 585
R4809 gnd.n6258 gnd.n6256 585
R4810 gnd.n6310 gnd.n6309 585
R4811 gnd.n6309 gnd.n976 585
R4812 gnd.n6308 gnd.n6260 585
R4813 gnd.n6308 gnd.n6307 585
R4814 gnd.n6295 gnd.n6261 585
R4815 gnd.n6261 gnd.n984 585
R4816 gnd.n6297 gnd.n6296 585
R4817 gnd.n6298 gnd.n6297 585
R4818 gnd.n6294 gnd.n6268 585
R4819 gnd.n6268 gnd.n6267 585
R4820 gnd.n6293 gnd.n6292 585
R4821 gnd.n6292 gnd.n992 585
R4822 gnd.n6291 gnd.n6269 585
R4823 gnd.n6291 gnd.n990 585
R4824 gnd.n6290 gnd.n6273 585
R4825 gnd.n6290 gnd.n6289 585
R4826 gnd.n6272 gnd.n6270 585
R4827 gnd.n6270 gnd.n1000 585
R4828 gnd.n6271 gnd.n1038 585
R4829 gnd.n1038 gnd.n998 585
R4830 gnd.n6416 gnd.n1037 585
R4831 gnd.n6416 gnd.n6415 585
R4832 gnd.n6418 gnd.n6417 585
R4833 gnd.n6417 gnd.n1008 585
R4834 gnd.n6419 gnd.n1035 585
R4835 gnd.n1035 gnd.n1006 585
R4836 gnd.n6421 gnd.n6420 585
R4837 gnd.n6422 gnd.n6421 585
R4838 gnd.n1036 gnd.n1034 585
R4839 gnd.n1034 gnd.n1016 585
R4840 gnd.n1170 gnd.n1169 585
R4841 gnd.n1170 gnd.n1014 585
R4842 gnd.n1172 gnd.n1171 585
R4843 gnd.n1171 gnd.n1025 585
R4844 gnd.n1173 gnd.n1023 585
R4845 gnd.n6430 gnd.n1023 585
R4846 gnd.n1175 gnd.n1174 585
R4847 gnd.n1174 gnd.n1022 585
R4848 gnd.n1176 gnd.n1165 585
R4849 gnd.n1165 gnd.n1049 585
R4850 gnd.n1178 gnd.n1177 585
R4851 gnd.n1179 gnd.n1178 585
R4852 gnd.n1168 gnd.n1164 585
R4853 gnd.n1164 gnd.n1058 585
R4854 gnd.n1167 gnd.n1166 585
R4855 gnd.n1166 gnd.n1056 585
R4856 gnd.n1156 gnd.n1155 585
R4857 gnd.n6080 gnd.n1156 585
R4858 gnd.n6083 gnd.n6082 585
R4859 gnd.n6082 gnd.n6081 585
R4860 gnd.n6084 gnd.n1152 585
R4861 gnd.n1152 gnd.n1065 585
R4862 gnd.n6086 gnd.n6085 585
R4863 gnd.n6087 gnd.n6086 585
R4864 gnd.n1154 gnd.n1151 585
R4865 gnd.n1151 gnd.n1149 585
R4866 gnd.n1153 gnd.n1140 585
R4867 gnd.n6093 gnd.n1140 585
R4868 gnd.n6096 gnd.n1139 585
R4869 gnd.n6096 gnd.n6095 585
R4870 gnd.n6098 gnd.n6097 585
R4871 gnd.n6097 gnd.n1080 585
R4872 gnd.n6099 gnd.n1136 585
R4873 gnd.n1136 gnd.n1078 585
R4874 gnd.n6101 gnd.n6100 585
R4875 gnd.n6102 gnd.n6101 585
R4876 gnd.n1138 gnd.n1135 585
R4877 gnd.n1135 gnd.n1087 585
R4878 gnd.n1137 gnd.n1124 585
R4879 gnd.n6108 gnd.n1124 585
R4880 gnd.n6111 gnd.n1123 585
R4881 gnd.n6111 gnd.n6110 585
R4882 gnd.n6113 gnd.n6112 585
R4883 gnd.n6112 gnd.n1095 585
R4884 gnd.n6114 gnd.n1121 585
R4885 gnd.n1121 gnd.n1093 585
R4886 gnd.n6116 gnd.n6115 585
R4887 gnd.n6117 gnd.n6116 585
R4888 gnd.n1122 gnd.n1120 585
R4889 gnd.n1120 gnd.n1103 585
R4890 gnd.n5871 gnd.n5870 585
R4891 gnd.n5871 gnd.n1101 585
R4892 gnd.n5873 gnd.n5872 585
R4893 gnd.n5872 gnd.n1111 585
R4894 gnd.n5874 gnd.n1109 585
R4895 gnd.n6125 gnd.n1109 585
R4896 gnd.n5875 gnd.n5869 585
R4897 gnd.n5869 gnd.n1200 585
R4898 gnd.n5877 gnd.n5876 585
R4899 gnd.n5877 gnd.n1199 585
R4900 gnd.n5941 gnd.n5868 585
R4901 gnd.n5941 gnd.n5940 585
R4902 gnd.n5943 gnd.n5942 585
R4903 gnd.n5942 gnd.n1209 585
R4904 gnd.n5944 gnd.n5866 585
R4905 gnd.n5866 gnd.n1207 585
R4906 gnd.n5946 gnd.n5945 585
R4907 gnd.n5947 gnd.n5946 585
R4908 gnd.n5867 gnd.n5865 585
R4909 gnd.n5865 gnd.n1218 585
R4910 gnd.n5924 gnd.n5885 585
R4911 gnd.n5885 gnd.n1216 585
R4912 gnd.n5926 gnd.n5925 585
R4913 gnd.n5927 gnd.n5926 585
R4914 gnd.n5923 gnd.n5884 585
R4915 gnd.n5884 gnd.n1225 585
R4916 gnd.n5922 gnd.n5921 585
R4917 gnd.n5921 gnd.n5920 585
R4918 gnd.n5887 gnd.n5886 585
R4919 gnd.n5889 gnd.n5887 585
R4920 gnd.n5907 gnd.n5906 585
R4921 gnd.n5906 gnd.n1233 585
R4922 gnd.n5908 gnd.n5903 585
R4923 gnd.n5903 gnd.n1231 585
R4924 gnd.n5910 gnd.n5909 585
R4925 gnd.n5911 gnd.n5910 585
R4926 gnd.n5905 gnd.n5902 585
R4927 gnd.n5902 gnd.n1241 585
R4928 gnd.n5904 gnd.n1276 585
R4929 gnd.n1276 gnd.n1239 585
R4930 gnd.n5969 gnd.n1275 585
R4931 gnd.n5969 gnd.n5968 585
R4932 gnd.n5971 gnd.n5970 585
R4933 gnd.n5970 gnd.n1248 585
R4934 gnd.n5972 gnd.n1273 585
R4935 gnd.n5852 gnd.n1273 585
R4936 gnd.n5974 gnd.n5973 585
R4937 gnd.n5975 gnd.n5974 585
R4938 gnd.n1274 gnd.n1272 585
R4939 gnd.n1272 gnd.n1256 585
R4940 gnd.n1521 gnd.n1520 585
R4941 gnd.n1521 gnd.n1254 585
R4942 gnd.n1523 gnd.n1522 585
R4943 gnd.n1522 gnd.n1264 585
R4944 gnd.n1524 gnd.n1262 585
R4945 gnd.n5983 gnd.n1262 585
R4946 gnd.n1526 gnd.n1525 585
R4947 gnd.n1525 gnd.n1288 585
R4948 gnd.n1527 gnd.n1413 585
R4949 gnd.n1413 gnd.n1287 585
R4950 gnd.n1529 gnd.n1528 585
R4951 gnd.n1530 gnd.n1529 585
R4952 gnd.n1519 gnd.n1412 585
R4953 gnd.n1412 gnd.n1297 585
R4954 gnd.n1518 gnd.n1517 585
R4955 gnd.n1517 gnd.n1295 585
R4956 gnd.n1516 gnd.n1515 585
R4957 gnd.n1514 gnd.n1513 585
R4958 gnd.n1512 gnd.n1436 585
R4959 gnd.n1512 gnd.n1305 585
R4960 gnd.n1511 gnd.n1510 585
R4961 gnd.n1509 gnd.n1508 585
R4962 gnd.n1507 gnd.n1438 585
R4963 gnd.n1505 gnd.n1504 585
R4964 gnd.n1503 gnd.n1439 585
R4965 gnd.n1502 gnd.n1501 585
R4966 gnd.n1499 gnd.n1440 585
R4967 gnd.n1497 gnd.n1496 585
R4968 gnd.n1495 gnd.n1441 585
R4969 gnd.n1494 gnd.n1493 585
R4970 gnd.n1491 gnd.n1442 585
R4971 gnd.n1489 gnd.n1488 585
R4972 gnd.n1487 gnd.n1443 585
R4973 gnd.n1486 gnd.n1485 585
R4974 gnd.n1483 gnd.n1444 585
R4975 gnd.n1481 gnd.n1480 585
R4976 gnd.n1479 gnd.n1445 585
R4977 gnd.n1478 gnd.n1477 585
R4978 gnd.n1475 gnd.n1446 585
R4979 gnd.n1473 gnd.n1472 585
R4980 gnd.n1471 gnd.n1447 585
R4981 gnd.n1470 gnd.n1469 585
R4982 gnd.n1467 gnd.n1448 585
R4983 gnd.n1465 gnd.n1464 585
R4984 gnd.n1463 gnd.n1449 585
R4985 gnd.n1462 gnd.n1461 585
R4986 gnd.n1459 gnd.n1458 585
R4987 gnd.n1457 gnd.n1456 585
R4988 gnd.n1455 gnd.n1391 585
R4989 gnd.n1605 gnd.n1604 585
R4990 gnd.n1602 gnd.n1390 585
R4991 gnd.n1600 gnd.n1599 585
R4992 gnd.n1598 gnd.n1393 585
R4993 gnd.n1596 gnd.n1595 585
R4994 gnd.n1593 gnd.n1396 585
R4995 gnd.n1591 gnd.n1590 585
R4996 gnd.n1589 gnd.n1397 585
R4997 gnd.n1588 gnd.n1587 585
R4998 gnd.n1585 gnd.n1398 585
R4999 gnd.n1583 gnd.n1582 585
R5000 gnd.n1581 gnd.n1399 585
R5001 gnd.n1580 gnd.n1579 585
R5002 gnd.n1577 gnd.n1400 585
R5003 gnd.n1575 gnd.n1574 585
R5004 gnd.n1573 gnd.n1401 585
R5005 gnd.n1572 gnd.n1571 585
R5006 gnd.n1569 gnd.n1402 585
R5007 gnd.n1567 gnd.n1566 585
R5008 gnd.n1565 gnd.n1403 585
R5009 gnd.n1564 gnd.n1563 585
R5010 gnd.n1561 gnd.n1404 585
R5011 gnd.n1559 gnd.n1558 585
R5012 gnd.n1557 gnd.n1405 585
R5013 gnd.n1556 gnd.n1555 585
R5014 gnd.n1553 gnd.n1406 585
R5015 gnd.n1551 gnd.n1550 585
R5016 gnd.n1549 gnd.n1407 585
R5017 gnd.n1548 gnd.n1547 585
R5018 gnd.n1545 gnd.n1408 585
R5019 gnd.n1543 gnd.n1542 585
R5020 gnd.n1541 gnd.n1409 585
R5021 gnd.n1540 gnd.n1539 585
R5022 gnd.n866 gnd.n865 585
R5023 gnd.n863 gnd.n677 585
R5024 gnd.n862 gnd.n861 585
R5025 gnd.n860 gnd.n859 585
R5026 gnd.n858 gnd.n679 585
R5027 gnd.n856 gnd.n855 585
R5028 gnd.n854 gnd.n680 585
R5029 gnd.n853 gnd.n852 585
R5030 gnd.n850 gnd.n681 585
R5031 gnd.n848 gnd.n847 585
R5032 gnd.n846 gnd.n682 585
R5033 gnd.n845 gnd.n844 585
R5034 gnd.n842 gnd.n683 585
R5035 gnd.n840 gnd.n839 585
R5036 gnd.n838 gnd.n684 585
R5037 gnd.n837 gnd.n836 585
R5038 gnd.n834 gnd.n685 585
R5039 gnd.n832 gnd.n831 585
R5040 gnd.n830 gnd.n686 585
R5041 gnd.n829 gnd.n828 585
R5042 gnd.n826 gnd.n687 585
R5043 gnd.n824 gnd.n823 585
R5044 gnd.n822 gnd.n688 585
R5045 gnd.n821 gnd.n820 585
R5046 gnd.n818 gnd.n689 585
R5047 gnd.n816 gnd.n815 585
R5048 gnd.n814 gnd.n690 585
R5049 gnd.n813 gnd.n812 585
R5050 gnd.n810 gnd.n691 585
R5051 gnd.n808 gnd.n807 585
R5052 gnd.n803 gnd.n692 585
R5053 gnd.n802 gnd.n801 585
R5054 gnd.n799 gnd.n648 585
R5055 gnd.n796 gnd.n534 585
R5056 gnd.n795 gnd.n794 585
R5057 gnd.n793 gnd.n792 585
R5058 gnd.n791 gnd.n694 585
R5059 gnd.n789 gnd.n788 585
R5060 gnd.n784 gnd.n695 585
R5061 gnd.n783 gnd.n782 585
R5062 gnd.n780 gnd.n696 585
R5063 gnd.n778 gnd.n777 585
R5064 gnd.n776 gnd.n697 585
R5065 gnd.n775 gnd.n774 585
R5066 gnd.n772 gnd.n698 585
R5067 gnd.n770 gnd.n769 585
R5068 gnd.n768 gnd.n699 585
R5069 gnd.n767 gnd.n766 585
R5070 gnd.n764 gnd.n700 585
R5071 gnd.n762 gnd.n761 585
R5072 gnd.n760 gnd.n701 585
R5073 gnd.n759 gnd.n758 585
R5074 gnd.n756 gnd.n702 585
R5075 gnd.n754 gnd.n753 585
R5076 gnd.n752 gnd.n703 585
R5077 gnd.n751 gnd.n750 585
R5078 gnd.n748 gnd.n704 585
R5079 gnd.n746 gnd.n745 585
R5080 gnd.n744 gnd.n705 585
R5081 gnd.n743 gnd.n742 585
R5082 gnd.n740 gnd.n706 585
R5083 gnd.n738 gnd.n737 585
R5084 gnd.n736 gnd.n707 585
R5085 gnd.n735 gnd.n734 585
R5086 gnd.n732 gnd.n708 585
R5087 gnd.n730 gnd.n729 585
R5088 gnd.n867 gnd.n676 585
R5089 gnd.n676 gnd.n646 585
R5090 gnd.n869 gnd.n868 585
R5091 gnd.n6769 gnd.n869 585
R5092 gnd.n668 gnd.n667 585
R5093 gnd.n668 gnd.n655 585
R5094 gnd.n6777 gnd.n6776 585
R5095 gnd.n6776 gnd.n6775 585
R5096 gnd.n6778 gnd.n665 585
R5097 gnd.n670 gnd.n665 585
R5098 gnd.n6780 gnd.n6779 585
R5099 gnd.n6781 gnd.n6780 585
R5100 gnd.n666 gnd.n664 585
R5101 gnd.n6576 gnd.n664 585
R5102 gnd.n6565 gnd.n903 585
R5103 gnd.n903 gnd.n898 585
R5104 gnd.n6567 gnd.n6566 585
R5105 gnd.n6569 gnd.n6567 585
R5106 gnd.n6564 gnd.n902 585
R5107 gnd.n902 gnd.n880 585
R5108 gnd.n6563 gnd.n6562 585
R5109 gnd.n6562 gnd.n879 585
R5110 gnd.n6561 gnd.n904 585
R5111 gnd.n6561 gnd.n6560 585
R5112 gnd.n6361 gnd.n905 585
R5113 gnd.n905 gnd.n890 585
R5114 gnd.n6363 gnd.n6362 585
R5115 gnd.n6362 gnd.n888 585
R5116 gnd.n6364 gnd.n912 585
R5117 gnd.n6552 gnd.n912 585
R5118 gnd.n6366 gnd.n6365 585
R5119 gnd.n6366 gnd.n911 585
R5120 gnd.n6368 gnd.n6367 585
R5121 gnd.n6367 gnd.n920 585
R5122 gnd.n6369 gnd.n6233 585
R5123 gnd.n6233 gnd.n919 585
R5124 gnd.n6371 gnd.n6370 585
R5125 gnd.n6372 gnd.n6371 585
R5126 gnd.n6360 gnd.n6232 585
R5127 gnd.n6374 gnd.n6232 585
R5128 gnd.n6359 gnd.n6358 585
R5129 gnd.n6358 gnd.n928 585
R5130 gnd.n6357 gnd.n6221 585
R5131 gnd.n6380 gnd.n6221 585
R5132 gnd.n6356 gnd.n6355 585
R5133 gnd.n6355 gnd.n939 585
R5134 gnd.n6354 gnd.n6234 585
R5135 gnd.n6354 gnd.n937 585
R5136 gnd.n6353 gnd.n6236 585
R5137 gnd.n6353 gnd.n6352 585
R5138 gnd.n6340 gnd.n6235 585
R5139 gnd.n6235 gnd.n947 585
R5140 gnd.n6341 gnd.n6244 585
R5141 gnd.n6244 gnd.n945 585
R5142 gnd.n6343 gnd.n6342 585
R5143 gnd.n6344 gnd.n6343 585
R5144 gnd.n6339 gnd.n6243 585
R5145 gnd.n6243 gnd.n955 585
R5146 gnd.n6338 gnd.n6337 585
R5147 gnd.n6337 gnd.n953 585
R5148 gnd.n6336 gnd.n6245 585
R5149 gnd.n6336 gnd.n6335 585
R5150 gnd.n6321 gnd.n6246 585
R5151 gnd.n6247 gnd.n6246 585
R5152 gnd.n6322 gnd.n6253 585
R5153 gnd.n6253 gnd.n961 585
R5154 gnd.n6324 gnd.n6323 585
R5155 gnd.n6326 gnd.n6324 585
R5156 gnd.n6320 gnd.n6252 585
R5157 gnd.n6252 gnd.n970 585
R5158 gnd.n6319 gnd.n6318 585
R5159 gnd.n6318 gnd.n968 585
R5160 gnd.n6317 gnd.n6254 585
R5161 gnd.n6317 gnd.n6316 585
R5162 gnd.n6302 gnd.n6255 585
R5163 gnd.n6256 gnd.n6255 585
R5164 gnd.n6303 gnd.n6263 585
R5165 gnd.n6263 gnd.n976 585
R5166 gnd.n6305 gnd.n6304 585
R5167 gnd.n6307 gnd.n6305 585
R5168 gnd.n6301 gnd.n6262 585
R5169 gnd.n6262 gnd.n984 585
R5170 gnd.n6300 gnd.n6299 585
R5171 gnd.n6299 gnd.n6298 585
R5172 gnd.n6265 gnd.n6264 585
R5173 gnd.n6267 gnd.n6265 585
R5174 gnd.n6284 gnd.n6283 585
R5175 gnd.n6283 gnd.n992 585
R5176 gnd.n6285 gnd.n6275 585
R5177 gnd.n6275 gnd.n990 585
R5178 gnd.n6287 gnd.n6286 585
R5179 gnd.n6289 gnd.n6287 585
R5180 gnd.n6282 gnd.n6274 585
R5181 gnd.n6274 gnd.n1000 585
R5182 gnd.n6281 gnd.n6280 585
R5183 gnd.n6280 gnd.n998 585
R5184 gnd.n6279 gnd.n1039 585
R5185 gnd.n6415 gnd.n1039 585
R5186 gnd.n6278 gnd.n6277 585
R5187 gnd.n6277 gnd.n1008 585
R5188 gnd.n6276 gnd.n1031 585
R5189 gnd.n1031 gnd.n1006 585
R5190 gnd.n6423 gnd.n1032 585
R5191 gnd.n6423 gnd.n6422 585
R5192 gnd.n6424 gnd.n1030 585
R5193 gnd.n6424 gnd.n1016 585
R5194 gnd.n6426 gnd.n6425 585
R5195 gnd.n6425 gnd.n1014 585
R5196 gnd.n6427 gnd.n1028 585
R5197 gnd.n1028 gnd.n1025 585
R5198 gnd.n6429 gnd.n6428 585
R5199 gnd.n6430 gnd.n6429 585
R5200 gnd.n1029 gnd.n1027 585
R5201 gnd.n1027 gnd.n1022 585
R5202 gnd.n1162 gnd.n1161 585
R5203 gnd.n1162 gnd.n1049 585
R5204 gnd.n1180 gnd.n1160 585
R5205 gnd.n1180 gnd.n1179 585
R5206 gnd.n1182 gnd.n1181 585
R5207 gnd.n1181 gnd.n1058 585
R5208 gnd.n1183 gnd.n1158 585
R5209 gnd.n1158 gnd.n1056 585
R5210 gnd.n1185 gnd.n1184 585
R5211 gnd.n6080 gnd.n1185 585
R5212 gnd.n1159 gnd.n1157 585
R5213 gnd.n6081 gnd.n1157 585
R5214 gnd.n1148 gnd.n1147 585
R5215 gnd.n1148 gnd.n1065 585
R5216 gnd.n6089 gnd.n6088 585
R5217 gnd.n6088 gnd.n6087 585
R5218 gnd.n6090 gnd.n1143 585
R5219 gnd.n1149 gnd.n1143 585
R5220 gnd.n6092 gnd.n6091 585
R5221 gnd.n6093 gnd.n6092 585
R5222 gnd.n1146 gnd.n1141 585
R5223 gnd.n6095 gnd.n1141 585
R5224 gnd.n1145 gnd.n1144 585
R5225 gnd.n1144 gnd.n1080 585
R5226 gnd.n1133 gnd.n1132 585
R5227 gnd.n1133 gnd.n1078 585
R5228 gnd.n6104 gnd.n6103 585
R5229 gnd.n6103 gnd.n6102 585
R5230 gnd.n6105 gnd.n1127 585
R5231 gnd.n1127 gnd.n1087 585
R5232 gnd.n6107 gnd.n6106 585
R5233 gnd.n6108 gnd.n6107 585
R5234 gnd.n1131 gnd.n1125 585
R5235 gnd.n6110 gnd.n1125 585
R5236 gnd.n1130 gnd.n1129 585
R5237 gnd.n1129 gnd.n1095 585
R5238 gnd.n1128 gnd.n1117 585
R5239 gnd.n1117 gnd.n1093 585
R5240 gnd.n6118 gnd.n1118 585
R5241 gnd.n6118 gnd.n6117 585
R5242 gnd.n6119 gnd.n1116 585
R5243 gnd.n6119 gnd.n1103 585
R5244 gnd.n6121 gnd.n6120 585
R5245 gnd.n6120 gnd.n1101 585
R5246 gnd.n6122 gnd.n1114 585
R5247 gnd.n1114 gnd.n1111 585
R5248 gnd.n6124 gnd.n6123 585
R5249 gnd.n6125 gnd.n6124 585
R5250 gnd.n1115 gnd.n1113 585
R5251 gnd.n1200 gnd.n1113 585
R5252 gnd.n5936 gnd.n5879 585
R5253 gnd.n5879 gnd.n1199 585
R5254 gnd.n5938 gnd.n5937 585
R5255 gnd.n5940 gnd.n5938 585
R5256 gnd.n5935 gnd.n5878 585
R5257 gnd.n5878 gnd.n1209 585
R5258 gnd.n5934 gnd.n5933 585
R5259 gnd.n5933 gnd.n1207 585
R5260 gnd.n5932 gnd.n5864 585
R5261 gnd.n5947 gnd.n5864 585
R5262 gnd.n5931 gnd.n5930 585
R5263 gnd.n5930 gnd.n1218 585
R5264 gnd.n5929 gnd.n5880 585
R5265 gnd.n5929 gnd.n1216 585
R5266 gnd.n5928 gnd.n5882 585
R5267 gnd.n5928 gnd.n5927 585
R5268 gnd.n5917 gnd.n5881 585
R5269 gnd.n5881 gnd.n1225 585
R5270 gnd.n5919 gnd.n5918 585
R5271 gnd.n5920 gnd.n5919 585
R5272 gnd.n5916 gnd.n5890 585
R5273 gnd.n5890 gnd.n5889 585
R5274 gnd.n5915 gnd.n5914 585
R5275 gnd.n5914 gnd.n1233 585
R5276 gnd.n5913 gnd.n5891 585
R5277 gnd.n5913 gnd.n1231 585
R5278 gnd.n5912 gnd.n5900 585
R5279 gnd.n5912 gnd.n5911 585
R5280 gnd.n5899 gnd.n5892 585
R5281 gnd.n5892 gnd.n1241 585
R5282 gnd.n5898 gnd.n5897 585
R5283 gnd.n5897 gnd.n1239 585
R5284 gnd.n5896 gnd.n1277 585
R5285 gnd.n5968 gnd.n1277 585
R5286 gnd.n5895 gnd.n5894 585
R5287 gnd.n5894 gnd.n1248 585
R5288 gnd.n5893 gnd.n1270 585
R5289 gnd.n5852 gnd.n1270 585
R5290 gnd.n5976 gnd.n1271 585
R5291 gnd.n5976 gnd.n5975 585
R5292 gnd.n5977 gnd.n1269 585
R5293 gnd.n5977 gnd.n1256 585
R5294 gnd.n5979 gnd.n5978 585
R5295 gnd.n5978 gnd.n1254 585
R5296 gnd.n5980 gnd.n1267 585
R5297 gnd.n1267 gnd.n1264 585
R5298 gnd.n5982 gnd.n5981 585
R5299 gnd.n5983 gnd.n5982 585
R5300 gnd.n1268 gnd.n1266 585
R5301 gnd.n1288 gnd.n1266 585
R5302 gnd.n1533 gnd.n1532 585
R5303 gnd.n1532 gnd.n1287 585
R5304 gnd.n1534 gnd.n1531 585
R5305 gnd.n1531 gnd.n1530 585
R5306 gnd.n1536 gnd.n1535 585
R5307 gnd.n1536 gnd.n1297 585
R5308 gnd.n1537 gnd.n1410 585
R5309 gnd.n1537 gnd.n1295 585
R5310 gnd.n3351 gnd.n2064 585
R5311 gnd.n2064 gnd.n1788 585
R5312 gnd.n7220 gnd.n7219 585
R5313 gnd.n7221 gnd.n7220 585
R5314 gnd.n7216 gnd.n343 585
R5315 gnd.n343 gnd.n311 585
R5316 gnd.n7215 gnd.n7214 585
R5317 gnd.n7214 gnd.n308 585
R5318 gnd.n7213 gnd.n346 585
R5319 gnd.n7213 gnd.n7212 585
R5320 gnd.n7150 gnd.n348 585
R5321 gnd.n361 gnd.n348 585
R5322 gnd.n7152 gnd.n7151 585
R5323 gnd.n7152 gnd.n359 585
R5324 gnd.n7154 gnd.n7153 585
R5325 gnd.n7153 gnd.n379 585
R5326 gnd.n7155 gnd.n389 585
R5327 gnd.n389 gnd.n372 585
R5328 gnd.n7157 gnd.n7156 585
R5329 gnd.n7158 gnd.n7157 585
R5330 gnd.n390 gnd.n388 585
R5331 gnd.n388 gnd.n386 585
R5332 gnd.n7141 gnd.n7140 585
R5333 gnd.n7140 gnd.n7139 585
R5334 gnd.n393 gnd.n392 585
R5335 gnd.n404 gnd.n393 585
R5336 gnd.n6913 gnd.n589 585
R5337 gnd.n589 gnd.n401 585
R5338 gnd.n6915 gnd.n6914 585
R5339 gnd.n6916 gnd.n6915 585
R5340 gnd.n590 gnd.n588 585
R5341 gnd.n588 gnd.n412 585
R5342 gnd.n6908 gnd.n6907 585
R5343 gnd.n6907 gnd.n422 585
R5344 gnd.n6906 gnd.n592 585
R5345 gnd.n6906 gnd.n6905 585
R5346 gnd.n6877 gnd.n593 585
R5347 gnd.n593 gnd.n431 585
R5348 gnd.n6879 gnd.n6878 585
R5349 gnd.n6879 gnd.n428 585
R5350 gnd.n6881 gnd.n6880 585
R5351 gnd.n6880 gnd.n440 585
R5352 gnd.n6882 gnd.n599 585
R5353 gnd.n599 gnd.n437 585
R5354 gnd.n6884 gnd.n6883 585
R5355 gnd.n6885 gnd.n6884 585
R5356 gnd.n600 gnd.n598 585
R5357 gnd.n598 gnd.n446 585
R5358 gnd.n6869 gnd.n6868 585
R5359 gnd.n6868 gnd.n456 585
R5360 gnd.n6867 gnd.n602 585
R5361 gnd.n6867 gnd.n6866 585
R5362 gnd.n6840 gnd.n6839 585
R5363 gnd.n6840 gnd.n465 585
R5364 gnd.n604 gnd.n603 585
R5365 gnd.n603 gnd.n462 585
R5366 gnd.n6835 gnd.n6834 585
R5367 gnd.n6834 gnd.n474 585
R5368 gnd.n6833 gnd.n606 585
R5369 gnd.n6833 gnd.n471 585
R5370 gnd.n6832 gnd.n6831 585
R5371 gnd.n6832 gnd.n483 585
R5372 gnd.n608 gnd.n607 585
R5373 gnd.n607 gnd.n480 585
R5374 gnd.n6827 gnd.n6826 585
R5375 gnd.n6826 gnd.n564 585
R5376 gnd.n6825 gnd.n610 585
R5377 gnd.n6825 gnd.n518 585
R5378 gnd.n6824 gnd.n6823 585
R5379 gnd.n6824 gnd.n489 585
R5380 gnd.n612 gnd.n611 585
R5381 gnd.n6816 gnd.n611 585
R5382 gnd.n6819 gnd.n6818 585
R5383 gnd.n6818 gnd.n6817 585
R5384 gnd.n615 gnd.n614 585
R5385 gnd.n616 gnd.n615 585
R5386 gnd.n6805 gnd.n641 585
R5387 gnd.n641 gnd.n639 585
R5388 gnd.n6807 gnd.n6806 585
R5389 gnd.n6808 gnd.n6807 585
R5390 gnd.n642 gnd.n640 585
R5391 gnd.n6613 gnd.n640 585
R5392 gnd.n6800 gnd.n6799 585
R5393 gnd.n6799 gnd.n6798 585
R5394 gnd.n645 gnd.n644 585
R5395 gnd.n6768 gnd.n645 585
R5396 gnd.n6788 gnd.n6787 585
R5397 gnd.n6789 gnd.n6788 585
R5398 gnd.n657 gnd.n656 585
R5399 gnd.n669 gnd.n656 585
R5400 gnd.n6783 gnd.n6782 585
R5401 gnd.n6782 gnd.n6781 585
R5402 gnd.n660 gnd.n659 585
R5403 gnd.n6577 gnd.n660 585
R5404 gnd.n6597 gnd.n883 585
R5405 gnd.n6568 gnd.n883 585
R5406 gnd.n6599 gnd.n6598 585
R5407 gnd.n6600 gnd.n6599 585
R5408 gnd.n884 gnd.n882 585
R5409 gnd.n906 gnd.n882 585
R5410 gnd.n6592 gnd.n6591 585
R5411 gnd.n6591 gnd.n6590 585
R5412 gnd.n887 gnd.n886 585
R5413 gnd.n6551 gnd.n887 585
R5414 gnd.n6539 gnd.n923 585
R5415 gnd.n6523 gnd.n923 585
R5416 gnd.n6541 gnd.n6540 585
R5417 gnd.n6542 gnd.n6541 585
R5418 gnd.n924 gnd.n922 585
R5419 gnd.n6373 gnd.n922 585
R5420 gnd.n6534 gnd.n6533 585
R5421 gnd.n6533 gnd.n6532 585
R5422 gnd.n927 gnd.n926 585
R5423 gnd.n6381 gnd.n927 585
R5424 gnd.n6517 gnd.n6516 585
R5425 gnd.t4 gnd.n6517 585
R5426 gnd.n941 gnd.n940 585
R5427 gnd.n6237 gnd.n940 585
R5428 gnd.n6512 gnd.n6511 585
R5429 gnd.n6511 gnd.n6510 585
R5430 gnd.n944 gnd.n943 585
R5431 gnd.n6242 gnd.n944 585
R5432 gnd.n6501 gnd.n6500 585
R5433 gnd.n6502 gnd.n6501 585
R5434 gnd.n957 gnd.n956 585
R5435 gnd.n6335 gnd.n956 585
R5436 gnd.n6496 gnd.n6495 585
R5437 gnd.n6495 gnd.n6494 585
R5438 gnd.n960 gnd.n959 585
R5439 gnd.n6325 gnd.n960 585
R5440 gnd.n6485 gnd.n6484 585
R5441 gnd.n6486 gnd.n6485 585
R5442 gnd.n972 gnd.n971 585
R5443 gnd.n6257 gnd.n971 585
R5444 gnd.n6480 gnd.n6479 585
R5445 gnd.n6479 gnd.n6478 585
R5446 gnd.n975 gnd.n974 585
R5447 gnd.n6306 gnd.n975 585
R5448 gnd.n6469 gnd.n6468 585
R5449 gnd.n6470 gnd.n6469 585
R5450 gnd.n986 gnd.n985 585
R5451 gnd.n6266 gnd.n985 585
R5452 gnd.n6464 gnd.n6463 585
R5453 gnd.n6463 gnd.n6462 585
R5454 gnd.n989 gnd.n988 585
R5455 gnd.n6288 gnd.n989 585
R5456 gnd.n6453 gnd.n6452 585
R5457 gnd.n6454 gnd.n6453 585
R5458 gnd.n1002 gnd.n1001 585
R5459 gnd.n6414 gnd.n1001 585
R5460 gnd.n6448 gnd.n6447 585
R5461 gnd.n6447 gnd.n6446 585
R5462 gnd.n1005 gnd.n1004 585
R5463 gnd.n1033 gnd.n1005 585
R5464 gnd.n6437 gnd.n6436 585
R5465 gnd.n6438 gnd.n6437 585
R5466 gnd.n1018 gnd.n1017 585
R5467 gnd.n1044 gnd.n1017 585
R5468 gnd.n6432 gnd.n6431 585
R5469 gnd.n6431 gnd.n6430 585
R5470 gnd.n1021 gnd.n1020 585
R5471 gnd.n6192 gnd.n1021 585
R5472 gnd.n6180 gnd.n1060 585
R5473 gnd.n1163 gnd.n1060 585
R5474 gnd.n6182 gnd.n6181 585
R5475 gnd.n6183 gnd.n6182 585
R5476 gnd.n1061 gnd.n1059 585
R5477 gnd.n6079 gnd.n1059 585
R5478 gnd.n6175 gnd.n6174 585
R5479 gnd.n6174 gnd.n6173 585
R5480 gnd.n1064 gnd.n1063 585
R5481 gnd.n1150 gnd.n1064 585
R5482 gnd.n6164 gnd.n6163 585
R5483 gnd.n6165 gnd.n6164 585
R5484 gnd.n1074 gnd.n1073 585
R5485 gnd.n6094 gnd.n1073 585
R5486 gnd.n6159 gnd.n6158 585
R5487 gnd.n6158 gnd.n6157 585
R5488 gnd.n1077 gnd.n1076 585
R5489 gnd.n1134 gnd.n1077 585
R5490 gnd.n6148 gnd.n6147 585
R5491 gnd.n6149 gnd.n6148 585
R5492 gnd.n1089 gnd.n1088 585
R5493 gnd.n6109 gnd.n1088 585
R5494 gnd.n6143 gnd.n6142 585
R5495 gnd.n6142 gnd.n6141 585
R5496 gnd.n1092 gnd.n1091 585
R5497 gnd.n1119 gnd.n1092 585
R5498 gnd.n6132 gnd.n6131 585
R5499 gnd.n6133 gnd.n6132 585
R5500 gnd.n1105 gnd.n1104 585
R5501 gnd.n1194 gnd.n1104 585
R5502 gnd.n6127 gnd.n6126 585
R5503 gnd.n6126 gnd.n6125 585
R5504 gnd.n1108 gnd.n1107 585
R5505 gnd.n6049 gnd.n1108 585
R5506 gnd.n6037 gnd.n1211 585
R5507 gnd.n5939 gnd.n1211 585
R5508 gnd.n6039 gnd.n6038 585
R5509 gnd.n6040 gnd.n6039 585
R5510 gnd.n1212 gnd.n1210 585
R5511 gnd.n5948 gnd.n1210 585
R5512 gnd.n6032 gnd.n6031 585
R5513 gnd.n6031 gnd.t21 585
R5514 gnd.n1215 gnd.n1214 585
R5515 gnd.n5883 gnd.n1215 585
R5516 gnd.n6022 gnd.n6021 585
R5517 gnd.n6023 gnd.n6022 585
R5518 gnd.n1227 gnd.n1226 585
R5519 gnd.n5888 gnd.n1226 585
R5520 gnd.n6017 gnd.n6016 585
R5521 gnd.n6016 gnd.n6015 585
R5522 gnd.n1230 gnd.n1229 585
R5523 gnd.n5901 gnd.n1230 585
R5524 gnd.n6006 gnd.n6005 585
R5525 gnd.n6007 gnd.n6006 585
R5526 gnd.n1243 gnd.n1242 585
R5527 gnd.n5967 gnd.n1242 585
R5528 gnd.n6001 gnd.n6000 585
R5529 gnd.n6000 gnd.n5999 585
R5530 gnd.n1246 gnd.n1245 585
R5531 gnd.n5853 gnd.n1246 585
R5532 gnd.n5990 gnd.n5989 585
R5533 gnd.n5991 gnd.n5990 585
R5534 gnd.n1258 gnd.n1257 585
R5535 gnd.n1282 gnd.n1257 585
R5536 gnd.n5985 gnd.n5984 585
R5537 gnd.n5984 gnd.n5983 585
R5538 gnd.n1261 gnd.n1260 585
R5539 gnd.n5844 gnd.n1261 585
R5540 gnd.n5832 gnd.n1299 585
R5541 gnd.n1411 gnd.n1299 585
R5542 gnd.n5834 gnd.n5833 585
R5543 gnd.n5835 gnd.n5834 585
R5544 gnd.n1300 gnd.n1298 585
R5545 gnd.n5677 gnd.n1298 585
R5546 gnd.n5827 gnd.n5826 585
R5547 gnd.n5826 gnd.n5825 585
R5548 gnd.n1303 gnd.n1302 585
R5549 gnd.n1312 gnd.n1303 585
R5550 gnd.n5816 gnd.n5815 585
R5551 gnd.n5817 gnd.n5816 585
R5552 gnd.n1314 gnd.n1313 585
R5553 gnd.n1313 gnd.n1310 585
R5554 gnd.n5811 gnd.n5810 585
R5555 gnd.n5810 gnd.n5809 585
R5556 gnd.n1317 gnd.n1316 585
R5557 gnd.n1318 gnd.n1317 585
R5558 gnd.n5356 gnd.n5352 585
R5559 gnd.n5352 gnd.n5351 585
R5560 gnd.n5359 gnd.n5357 585
R5561 gnd.n5359 gnd.n5358 585
R5562 gnd.n5360 gnd.n5350 585
R5563 gnd.n5360 gnd.n1356 585
R5564 gnd.n5362 gnd.n5361 585
R5565 gnd.n5361 gnd.n1354 585
R5566 gnd.n5363 gnd.n5345 585
R5567 gnd.n5345 gnd.n1649 585
R5568 gnd.n5365 gnd.n5364 585
R5569 gnd.n5365 gnd.n1658 585
R5570 gnd.n5366 gnd.n5344 585
R5571 gnd.n5366 gnd.n1655 585
R5572 gnd.n5368 gnd.n5367 585
R5573 gnd.n5367 gnd.n1668 585
R5574 gnd.n5369 gnd.n1835 585
R5575 gnd.n1835 gnd.n1665 585
R5576 gnd.n5371 gnd.n5370 585
R5577 gnd.n5372 gnd.n5371 585
R5578 gnd.n1836 gnd.n1834 585
R5579 gnd.n1834 gnd.n1674 585
R5580 gnd.n5338 gnd.n5337 585
R5581 gnd.n5337 gnd.n1684 585
R5582 gnd.n5336 gnd.n1838 585
R5583 gnd.n5336 gnd.n5335 585
R5584 gnd.n5307 gnd.n1839 585
R5585 gnd.n1839 gnd.n1693 585
R5586 gnd.n5309 gnd.n5308 585
R5587 gnd.n5309 gnd.n1690 585
R5588 gnd.n5311 gnd.n5310 585
R5589 gnd.n5310 gnd.n1702 585
R5590 gnd.n5312 gnd.n1845 585
R5591 gnd.n1845 gnd.n1699 585
R5592 gnd.n5314 gnd.n5313 585
R5593 gnd.n5315 gnd.n5314 585
R5594 gnd.n1846 gnd.n1844 585
R5595 gnd.n1844 gnd.n1708 585
R5596 gnd.n5299 gnd.n5298 585
R5597 gnd.n5298 gnd.n1718 585
R5598 gnd.n5297 gnd.n1848 585
R5599 gnd.n5297 gnd.n5296 585
R5600 gnd.n5267 gnd.n1849 585
R5601 gnd.n1849 gnd.n1727 585
R5602 gnd.n5269 gnd.n5268 585
R5603 gnd.n5269 gnd.n1724 585
R5604 gnd.n5271 gnd.n5270 585
R5605 gnd.n5270 gnd.n1736 585
R5606 gnd.n5272 gnd.n5256 585
R5607 gnd.n5256 gnd.n1733 585
R5608 gnd.n5274 gnd.n5273 585
R5609 gnd.n5275 gnd.n5274 585
R5610 gnd.n5257 gnd.n5255 585
R5611 gnd.n5255 gnd.n1742 585
R5612 gnd.n5259 gnd.n1805 585
R5613 gnd.n1805 gnd.n1752 585
R5614 gnd.n5431 gnd.n1804 585
R5615 gnd.n5431 gnd.n5430 585
R5616 gnd.n5433 gnd.n5432 585
R5617 gnd.n5432 gnd.n1761 585
R5618 gnd.n5434 gnd.n1799 585
R5619 gnd.n1799 gnd.n1758 585
R5620 gnd.n5436 gnd.n5435 585
R5621 gnd.n5437 gnd.n5436 585
R5622 gnd.n1800 gnd.n1798 585
R5623 gnd.n1798 gnd.n1795 585
R5624 gnd.n6760 gnd.n6759 585
R5625 gnd.n6759 gnd.n639 585
R5626 gnd.n6761 gnd.n638 585
R5627 gnd.n6808 gnd.n638 585
R5628 gnd.n6762 gnd.n6614 585
R5629 gnd.n6614 gnd.n6613 585
R5630 gnd.n871 gnd.n647 585
R5631 gnd.n6798 gnd.n647 585
R5632 gnd.n6767 gnd.n6766 585
R5633 gnd.n6768 gnd.n6767 585
R5634 gnd.n870 gnd.n654 585
R5635 gnd.n6789 gnd.n654 585
R5636 gnd.n6609 gnd.n6608 585
R5637 gnd.n6608 gnd.n669 585
R5638 gnd.n6607 gnd.n662 585
R5639 gnd.n6781 gnd.n662 585
R5640 gnd.n6606 gnd.n874 585
R5641 gnd.n6577 gnd.n874 585
R5642 gnd.n878 gnd.n873 585
R5643 gnd.n6568 gnd.n878 585
R5644 gnd.n6602 gnd.n6601 585
R5645 gnd.n6601 gnd.n6600 585
R5646 gnd.n877 gnd.n876 585
R5647 gnd.n906 gnd.n877 585
R5648 gnd.n915 gnd.n889 585
R5649 gnd.n6590 gnd.n889 585
R5650 gnd.n6550 gnd.n6549 585
R5651 gnd.n6551 gnd.n6550 585
R5652 gnd.n914 gnd.n913 585
R5653 gnd.n6523 gnd.n913 585
R5654 gnd.n6544 gnd.n6543 585
R5655 gnd.n6543 gnd.n6542 585
R5656 gnd.n918 gnd.n917 585
R5657 gnd.n6373 gnd.n918 585
R5658 gnd.n6383 gnd.n929 585
R5659 gnd.n6532 gnd.n929 585
R5660 gnd.n6384 gnd.n6382 585
R5661 gnd.n6382 gnd.n6381 585
R5662 gnd.n6219 gnd.n938 585
R5663 gnd.t4 gnd.n938 585
R5664 gnd.n6388 gnd.n6218 585
R5665 gnd.n6237 gnd.n6218 585
R5666 gnd.n6389 gnd.n946 585
R5667 gnd.n6510 gnd.n946 585
R5668 gnd.n6390 gnd.n6217 585
R5669 gnd.n6242 gnd.n6217 585
R5670 gnd.n6215 gnd.n954 585
R5671 gnd.n6502 gnd.n954 585
R5672 gnd.n6394 gnd.n6214 585
R5673 gnd.n6335 gnd.n6214 585
R5674 gnd.n6395 gnd.n962 585
R5675 gnd.n6494 gnd.n962 585
R5676 gnd.n6396 gnd.n6213 585
R5677 gnd.n6325 gnd.n6213 585
R5678 gnd.n6211 gnd.n969 585
R5679 gnd.n6486 gnd.n969 585
R5680 gnd.n6400 gnd.n6210 585
R5681 gnd.n6257 gnd.n6210 585
R5682 gnd.n6401 gnd.n977 585
R5683 gnd.n6478 gnd.n977 585
R5684 gnd.n6402 gnd.n6209 585
R5685 gnd.n6306 gnd.n6209 585
R5686 gnd.n6207 gnd.n983 585
R5687 gnd.n6470 gnd.n983 585
R5688 gnd.n6406 gnd.n6206 585
R5689 gnd.n6266 gnd.n6206 585
R5690 gnd.n6407 gnd.n991 585
R5691 gnd.n6462 gnd.n991 585
R5692 gnd.n6408 gnd.n6205 585
R5693 gnd.n6288 gnd.n6205 585
R5694 gnd.n1041 gnd.n999 585
R5695 gnd.n6454 gnd.n999 585
R5696 gnd.n6413 gnd.n6412 585
R5697 gnd.n6414 gnd.n6413 585
R5698 gnd.n1040 gnd.n1007 585
R5699 gnd.n6446 gnd.n1007 585
R5700 gnd.n6201 gnd.n6200 585
R5701 gnd.n6200 gnd.n1033 585
R5702 gnd.n6199 gnd.n1015 585
R5703 gnd.n6438 gnd.n1015 585
R5704 gnd.n6198 gnd.n1045 585
R5705 gnd.n1045 gnd.n1044 585
R5706 gnd.n1043 gnd.n1024 585
R5707 gnd.n6430 gnd.n1024 585
R5708 gnd.n6194 gnd.n6193 585
R5709 gnd.n6193 gnd.n6192 585
R5710 gnd.n1048 gnd.n1047 585
R5711 gnd.n1163 gnd.n1048 585
R5712 gnd.n1187 gnd.n1057 585
R5713 gnd.n6183 gnd.n1057 585
R5714 gnd.n6078 gnd.n6077 585
R5715 gnd.n6079 gnd.n6078 585
R5716 gnd.n1186 gnd.n1066 585
R5717 gnd.n6173 gnd.n1066 585
R5718 gnd.n6072 gnd.n6071 585
R5719 gnd.n6071 gnd.n1150 585
R5720 gnd.n6070 gnd.n1072 585
R5721 gnd.n6165 gnd.n1072 585
R5722 gnd.n6069 gnd.n1142 585
R5723 gnd.n6094 gnd.n1142 585
R5724 gnd.n1189 gnd.n1079 585
R5725 gnd.n6157 gnd.n1079 585
R5726 gnd.n6065 gnd.n6064 585
R5727 gnd.n6064 gnd.n1134 585
R5728 gnd.n6063 gnd.n1086 585
R5729 gnd.n6149 gnd.n1086 585
R5730 gnd.n6062 gnd.n1126 585
R5731 gnd.n6109 gnd.n1126 585
R5732 gnd.n1191 gnd.n1094 585
R5733 gnd.n6141 gnd.n1094 585
R5734 gnd.n6058 gnd.n6057 585
R5735 gnd.n6057 gnd.n1119 585
R5736 gnd.n6056 gnd.n1102 585
R5737 gnd.n6133 gnd.n1102 585
R5738 gnd.n6055 gnd.n1195 585
R5739 gnd.n1195 gnd.n1194 585
R5740 gnd.n1193 gnd.n1110 585
R5741 gnd.n6125 gnd.n1110 585
R5742 gnd.n6051 gnd.n6050 585
R5743 gnd.n6050 gnd.n6049 585
R5744 gnd.n1198 gnd.n1197 585
R5745 gnd.n5939 gnd.n1198 585
R5746 gnd.n5950 gnd.n1208 585
R5747 gnd.n6040 gnd.n1208 585
R5748 gnd.n5953 gnd.n5949 585
R5749 gnd.n5949 gnd.n5948 585
R5750 gnd.n5954 gnd.n1217 585
R5751 gnd.t21 gnd.n1217 585
R5752 gnd.n5955 gnd.n5863 585
R5753 gnd.n5883 gnd.n5863 585
R5754 gnd.n5861 gnd.n1224 585
R5755 gnd.n6023 gnd.n1224 585
R5756 gnd.n5959 gnd.n5860 585
R5757 gnd.n5888 gnd.n5860 585
R5758 gnd.n5960 gnd.n1232 585
R5759 gnd.n6015 gnd.n1232 585
R5760 gnd.n5961 gnd.n5859 585
R5761 gnd.n5901 gnd.n5859 585
R5762 gnd.n1279 gnd.n1240 585
R5763 gnd.n6007 gnd.n1240 585
R5764 gnd.n5966 gnd.n5965 585
R5765 gnd.n5967 gnd.n5966 585
R5766 gnd.n1278 gnd.n1247 585
R5767 gnd.n5999 gnd.n1247 585
R5768 gnd.n5855 gnd.n5854 585
R5769 gnd.n5854 gnd.n5853 585
R5770 gnd.n5851 gnd.n1255 585
R5771 gnd.n5991 gnd.n1255 585
R5772 gnd.n5850 gnd.n1283 585
R5773 gnd.n1283 gnd.n1282 585
R5774 gnd.n1281 gnd.n1263 585
R5775 gnd.n5983 gnd.n1263 585
R5776 gnd.n5846 gnd.n5845 585
R5777 gnd.n5845 gnd.n5844 585
R5778 gnd.n1286 gnd.n1285 585
R5779 gnd.n1411 gnd.n1286 585
R5780 gnd.n5680 gnd.n1296 585
R5781 gnd.n5835 gnd.n1296 585
R5782 gnd.n5679 gnd.n5678 585
R5783 gnd.n5678 gnd.n5677 585
R5784 gnd.n5684 gnd.n1304 585
R5785 gnd.n5825 gnd.n1304 585
R5786 gnd.n5685 gnd.n5676 585
R5787 gnd.n5676 gnd.n1312 585
R5788 gnd.n5686 gnd.n1311 585
R5789 gnd.n5817 gnd.n1311 585
R5790 gnd.n5582 gnd.n5581 585
R5791 gnd.n5669 gnd.n5583 585
R5792 gnd.n5668 gnd.n5584 585
R5793 gnd.n5593 gnd.n5585 585
R5794 gnd.n5661 gnd.n5594 585
R5795 gnd.n5660 gnd.n5595 585
R5796 gnd.n5597 gnd.n5596 585
R5797 gnd.n5653 gnd.n5606 585
R5798 gnd.n5652 gnd.n5607 585
R5799 gnd.n5616 gnd.n5608 585
R5800 gnd.n5645 gnd.n5617 585
R5801 gnd.n5644 gnd.n5618 585
R5802 gnd.n5620 gnd.n5619 585
R5803 gnd.n5637 gnd.n5632 585
R5804 gnd.n5636 gnd.n5633 585
R5805 gnd.n1344 gnd.n1343 585
R5806 gnd.n5778 gnd.n1345 585
R5807 gnd.n5781 gnd.n5780 585
R5808 gnd.n5779 gnd.n1340 585
R5809 gnd.n5787 gnd.n5786 585
R5810 gnd.n5789 gnd.n5788 585
R5811 gnd.n5792 gnd.n5791 585
R5812 gnd.n5790 gnd.n1338 585
R5813 gnd.n5797 gnd.n5796 585
R5814 gnd.n5799 gnd.n5798 585
R5815 gnd.n5802 gnd.n5801 585
R5816 gnd.n1333 gnd.n1332 585
R5817 gnd.n5807 gnd.n5806 585
R5818 gnd.n1334 gnd.n1309 585
R5819 gnd.n5809 gnd.n1309 585
R5820 gnd.n6811 gnd.n632 585
R5821 gnd.n639 gnd.n632 585
R5822 gnd.n6810 gnd.n6809 585
R5823 gnd.n6809 gnd.n6808 585
R5824 gnd.n637 gnd.n636 585
R5825 gnd.n6613 gnd.n637 585
R5826 gnd.n6797 gnd.n6796 585
R5827 gnd.n6798 gnd.n6797 585
R5828 gnd.n650 gnd.n649 585
R5829 gnd.n6768 gnd.n649 585
R5830 gnd.n6791 gnd.n6790 585
R5831 gnd.n6790 gnd.n6789 585
R5832 gnd.n653 gnd.n652 585
R5833 gnd.n669 gnd.n653 585
R5834 gnd.n6579 gnd.n663 585
R5835 gnd.n6781 gnd.n663 585
R5836 gnd.n6582 gnd.n6578 585
R5837 gnd.n6578 gnd.n6577 585
R5838 gnd.n6583 gnd.n897 585
R5839 gnd.n6568 gnd.n897 585
R5840 gnd.n6584 gnd.n881 585
R5841 gnd.n6600 gnd.n881 585
R5842 gnd.n894 gnd.n892 585
R5843 gnd.n906 gnd.n892 585
R5844 gnd.n6589 gnd.n6588 585
R5845 gnd.n6590 gnd.n6589 585
R5846 gnd.n893 gnd.n891 585
R5847 gnd.n6551 gnd.n891 585
R5848 gnd.n6525 gnd.n6524 585
R5849 gnd.n6524 gnd.n6523 585
R5850 gnd.n6526 gnd.n921 585
R5851 gnd.n6542 gnd.n921 585
R5852 gnd.n933 gnd.n931 585
R5853 gnd.n6373 gnd.n931 585
R5854 gnd.n6531 gnd.n6530 585
R5855 gnd.n6532 gnd.n6531 585
R5856 gnd.n932 gnd.n930 585
R5857 gnd.n6381 gnd.n930 585
R5858 gnd.n6519 gnd.n6518 585
R5859 gnd.n6518 gnd.t4 585
R5860 gnd.n936 gnd.n935 585
R5861 gnd.n6237 gnd.n936 585
R5862 gnd.n6509 gnd.n6508 585
R5863 gnd.n6510 gnd.n6509 585
R5864 gnd.n949 gnd.n948 585
R5865 gnd.n6242 gnd.n948 585
R5866 gnd.n6504 gnd.n6503 585
R5867 gnd.n6503 gnd.n6502 585
R5868 gnd.n952 gnd.n951 585
R5869 gnd.n6335 gnd.n952 585
R5870 gnd.n6493 gnd.n6492 585
R5871 gnd.n6494 gnd.n6493 585
R5872 gnd.n964 gnd.n963 585
R5873 gnd.n6325 gnd.n963 585
R5874 gnd.n6488 gnd.n6487 585
R5875 gnd.n6487 gnd.n6486 585
R5876 gnd.n967 gnd.n966 585
R5877 gnd.n6257 gnd.n967 585
R5878 gnd.n6477 gnd.n6476 585
R5879 gnd.n6478 gnd.n6477 585
R5880 gnd.n979 gnd.n978 585
R5881 gnd.n6306 gnd.n978 585
R5882 gnd.n6472 gnd.n6471 585
R5883 gnd.n6471 gnd.n6470 585
R5884 gnd.n982 gnd.n981 585
R5885 gnd.n6266 gnd.n982 585
R5886 gnd.n6461 gnd.n6460 585
R5887 gnd.n6462 gnd.n6461 585
R5888 gnd.n994 gnd.n993 585
R5889 gnd.n6288 gnd.n993 585
R5890 gnd.n6456 gnd.n6455 585
R5891 gnd.n6455 gnd.n6454 585
R5892 gnd.n997 gnd.n996 585
R5893 gnd.n6414 gnd.n997 585
R5894 gnd.n6445 gnd.n6444 585
R5895 gnd.n6446 gnd.n6445 585
R5896 gnd.n1010 gnd.n1009 585
R5897 gnd.n1033 gnd.n1009 585
R5898 gnd.n6440 gnd.n6439 585
R5899 gnd.n6439 gnd.n6438 585
R5900 gnd.n1013 gnd.n1012 585
R5901 gnd.n1044 gnd.n1013 585
R5902 gnd.n1052 gnd.n1026 585
R5903 gnd.n6430 gnd.n1026 585
R5904 gnd.n6191 gnd.n6190 585
R5905 gnd.n6192 gnd.n6191 585
R5906 gnd.n1051 gnd.n1050 585
R5907 gnd.n1163 gnd.n1050 585
R5908 gnd.n6185 gnd.n6184 585
R5909 gnd.n6184 gnd.n6183 585
R5910 gnd.n1055 gnd.n1054 585
R5911 gnd.n6079 gnd.n1055 585
R5912 gnd.n6172 gnd.n6171 585
R5913 gnd.n6173 gnd.n6172 585
R5914 gnd.n1068 gnd.n1067 585
R5915 gnd.n1150 gnd.n1067 585
R5916 gnd.n6167 gnd.n6166 585
R5917 gnd.n6166 gnd.n6165 585
R5918 gnd.n1071 gnd.n1070 585
R5919 gnd.n6094 gnd.n1071 585
R5920 gnd.n6156 gnd.n6155 585
R5921 gnd.n6157 gnd.n6156 585
R5922 gnd.n1082 gnd.n1081 585
R5923 gnd.n1134 gnd.n1081 585
R5924 gnd.n6151 gnd.n6150 585
R5925 gnd.n6150 gnd.n6149 585
R5926 gnd.n1085 gnd.n1084 585
R5927 gnd.n6109 gnd.n1085 585
R5928 gnd.n6140 gnd.n6139 585
R5929 gnd.n6141 gnd.n6140 585
R5930 gnd.n1097 gnd.n1096 585
R5931 gnd.n1119 gnd.n1096 585
R5932 gnd.n6135 gnd.n6134 585
R5933 gnd.n6134 gnd.n6133 585
R5934 gnd.n1100 gnd.n1099 585
R5935 gnd.n1194 gnd.n1100 585
R5936 gnd.n1203 gnd.n1112 585
R5937 gnd.n6125 gnd.n1112 585
R5938 gnd.n6048 gnd.n6047 585
R5939 gnd.n6049 gnd.n6048 585
R5940 gnd.n1202 gnd.n1201 585
R5941 gnd.n5939 gnd.n1201 585
R5942 gnd.n6042 gnd.n6041 585
R5943 gnd.n6041 gnd.n6040 585
R5944 gnd.n1206 gnd.n1205 585
R5945 gnd.n5948 gnd.n1206 585
R5946 gnd.n6030 gnd.n6029 585
R5947 gnd.t21 gnd.n6030 585
R5948 gnd.n1220 gnd.n1219 585
R5949 gnd.n5883 gnd.n1219 585
R5950 gnd.n6025 gnd.n6024 585
R5951 gnd.n6024 gnd.n6023 585
R5952 gnd.n1223 gnd.n1222 585
R5953 gnd.n5888 gnd.n1223 585
R5954 gnd.n6014 gnd.n6013 585
R5955 gnd.n6015 gnd.n6014 585
R5956 gnd.n1235 gnd.n1234 585
R5957 gnd.n5901 gnd.n1234 585
R5958 gnd.n6009 gnd.n6008 585
R5959 gnd.n6008 gnd.n6007 585
R5960 gnd.n1238 gnd.n1237 585
R5961 gnd.n5967 gnd.n1238 585
R5962 gnd.n5998 gnd.n5997 585
R5963 gnd.n5999 gnd.n5998 585
R5964 gnd.n1250 gnd.n1249 585
R5965 gnd.n5853 gnd.n1249 585
R5966 gnd.n5993 gnd.n5992 585
R5967 gnd.n5992 gnd.n5991 585
R5968 gnd.n1253 gnd.n1252 585
R5969 gnd.n1282 gnd.n1253 585
R5970 gnd.n1291 gnd.n1265 585
R5971 gnd.n5983 gnd.n1265 585
R5972 gnd.n5843 gnd.n5842 585
R5973 gnd.n5844 gnd.n5843 585
R5974 gnd.n1290 gnd.n1289 585
R5975 gnd.n1411 gnd.n1289 585
R5976 gnd.n5837 gnd.n5836 585
R5977 gnd.n5836 gnd.n5835 585
R5978 gnd.n1294 gnd.n1293 585
R5979 gnd.n5677 gnd.n1294 585
R5980 gnd.n5824 gnd.n5823 585
R5981 gnd.n5825 gnd.n5824 585
R5982 gnd.n1307 gnd.n1306 585
R5983 gnd.n1312 gnd.n1306 585
R5984 gnd.n5819 gnd.n5818 585
R5985 gnd.n5818 gnd.n5817 585
R5986 gnd.n6815 gnd.n6814 585
R5987 gnd.n6817 gnd.n6815 585
R5988 gnd.n633 gnd.n631 585
R5989 gnd.n6694 gnd.n6693 585
R5990 gnd.n6695 gnd.n6692 585
R5991 gnd.n6687 gnd.n6686 585
R5992 gnd.n6699 gnd.n6685 585
R5993 gnd.n6700 gnd.n6684 585
R5994 gnd.n6701 gnd.n6683 585
R5995 gnd.n6681 gnd.n6680 585
R5996 gnd.n6705 gnd.n6679 585
R5997 gnd.n6706 gnd.n6678 585
R5998 gnd.n6707 gnd.n6677 585
R5999 gnd.n6674 gnd.n6673 585
R6000 gnd.n6717 gnd.n6672 585
R6001 gnd.n6718 gnd.n6671 585
R6002 gnd.n6670 gnd.n6662 585
R6003 gnd.n6725 gnd.n6661 585
R6004 gnd.n6726 gnd.n6660 585
R6005 gnd.n6654 gnd.n6653 585
R6006 gnd.n6733 gnd.n6652 585
R6007 gnd.n6734 gnd.n6651 585
R6008 gnd.n6650 gnd.n6642 585
R6009 gnd.n6741 gnd.n6641 585
R6010 gnd.n6742 gnd.n6640 585
R6011 gnd.n6634 gnd.n6633 585
R6012 gnd.n6749 gnd.n6632 585
R6013 gnd.n6750 gnd.n6631 585
R6014 gnd.n6630 gnd.n6616 585
R6015 gnd.n6758 gnd.n6757 585
R6016 gnd.n730 gnd.n675 506.916
R6017 gnd.n865 gnd.n676 506.916
R6018 gnd.n1539 gnd.n1537 506.916
R6019 gnd.n1517 gnd.n1516 506.916
R6020 gnd.n3142 gnd.n3141 414.56
R6021 gnd.n1394 gnd.t126 389.64
R6022 gnd.n804 gnd.t62 389.64
R6023 gnd.n1450 gnd.t73 389.64
R6024 gnd.n785 gnd.t120 389.64
R6025 gnd.n1336 gnd.t110 371.625
R6026 gnd.n118 gnd.t44 371.625
R6027 gnd.n6712 gnd.t84 371.625
R6028 gnd.n1348 gnd.t97 371.625
R6029 gnd.n537 gnd.t77 371.625
R6030 gnd.n559 gnd.t48 371.625
R6031 gnd.n197 gnd.t123 371.625
R6032 gnd.n7536 gnd.t132 371.625
R6033 gnd.n4900 gnd.t70 371.625
R6034 gnd.n4932 gnd.t37 371.625
R6035 gnd.n4761 gnd.t107 371.625
R6036 gnd.n1641 gnd.t66 371.625
R6037 gnd.n1388 gnd.t94 371.625
R6038 gnd.n6689 gnd.t90 371.625
R6039 gnd.n3838 gnd.t33 323.425
R6040 gnd.n2027 gnd.t80 323.425
R6041 gnd.n4625 gnd.n4599 289.615
R6042 gnd.n4593 gnd.n4567 289.615
R6043 gnd.n4561 gnd.n4535 289.615
R6044 gnd.n4530 gnd.n4504 289.615
R6045 gnd.n4498 gnd.n4472 289.615
R6046 gnd.n4466 gnd.n4440 289.615
R6047 gnd.n4434 gnd.n4408 289.615
R6048 gnd.n4403 gnd.n4377 289.615
R6049 gnd.n3912 gnd.t103 279.217
R6050 gnd.n2053 gnd.t55 279.217
R6051 gnd.n1420 gnd.t116 260.649
R6052 gnd.n720 gnd.t119 260.649
R6053 gnd.n1435 gnd.n1305 256.663
R6054 gnd.n1437 gnd.n1305 256.663
R6055 gnd.n1506 gnd.n1305 256.663
R6056 gnd.n1500 gnd.n1305 256.663
R6057 gnd.n1498 gnd.n1305 256.663
R6058 gnd.n1492 gnd.n1305 256.663
R6059 gnd.n1490 gnd.n1305 256.663
R6060 gnd.n1484 gnd.n1305 256.663
R6061 gnd.n1482 gnd.n1305 256.663
R6062 gnd.n1476 gnd.n1305 256.663
R6063 gnd.n1474 gnd.n1305 256.663
R6064 gnd.n1468 gnd.n1305 256.663
R6065 gnd.n1466 gnd.n1305 256.663
R6066 gnd.n1460 gnd.n1305 256.663
R6067 gnd.n1453 gnd.n1305 256.663
R6068 gnd.n1454 gnd.n1305 256.663
R6069 gnd.n1605 gnd.n1392 256.663
R6070 gnd.n1603 gnd.n1305 256.663
R6071 gnd.n1601 gnd.n1305 256.663
R6072 gnd.n1594 gnd.n1305 256.663
R6073 gnd.n1592 gnd.n1305 256.663
R6074 gnd.n1586 gnd.n1305 256.663
R6075 gnd.n1584 gnd.n1305 256.663
R6076 gnd.n1578 gnd.n1305 256.663
R6077 gnd.n1576 gnd.n1305 256.663
R6078 gnd.n1570 gnd.n1305 256.663
R6079 gnd.n1568 gnd.n1305 256.663
R6080 gnd.n1562 gnd.n1305 256.663
R6081 gnd.n1560 gnd.n1305 256.663
R6082 gnd.n1554 gnd.n1305 256.663
R6083 gnd.n1552 gnd.n1305 256.663
R6084 gnd.n1546 gnd.n1305 256.663
R6085 gnd.n1544 gnd.n1305 256.663
R6086 gnd.n1538 gnd.n1305 256.663
R6087 gnd.n864 gnd.n648 256.663
R6088 gnd.n678 gnd.n648 256.663
R6089 gnd.n857 gnd.n648 256.663
R6090 gnd.n851 gnd.n648 256.663
R6091 gnd.n849 gnd.n648 256.663
R6092 gnd.n843 gnd.n648 256.663
R6093 gnd.n841 gnd.n648 256.663
R6094 gnd.n835 gnd.n648 256.663
R6095 gnd.n833 gnd.n648 256.663
R6096 gnd.n827 gnd.n648 256.663
R6097 gnd.n825 gnd.n648 256.663
R6098 gnd.n819 gnd.n648 256.663
R6099 gnd.n817 gnd.n648 256.663
R6100 gnd.n811 gnd.n648 256.663
R6101 gnd.n809 gnd.n648 256.663
R6102 gnd.n800 gnd.n648 256.663
R6103 gnd.n798 gnd.n534 256.663
R6104 gnd.n797 gnd.n648 256.663
R6105 gnd.n693 gnd.n648 256.663
R6106 gnd.n790 gnd.n648 256.663
R6107 gnd.n781 gnd.n648 256.663
R6108 gnd.n779 gnd.n648 256.663
R6109 gnd.n773 gnd.n648 256.663
R6110 gnd.n771 gnd.n648 256.663
R6111 gnd.n765 gnd.n648 256.663
R6112 gnd.n763 gnd.n648 256.663
R6113 gnd.n757 gnd.n648 256.663
R6114 gnd.n755 gnd.n648 256.663
R6115 gnd.n749 gnd.n648 256.663
R6116 gnd.n747 gnd.n648 256.663
R6117 gnd.n741 gnd.n648 256.663
R6118 gnd.n739 gnd.n648 256.663
R6119 gnd.n733 gnd.n648 256.663
R6120 gnd.n731 gnd.n648 256.663
R6121 gnd.n4781 gnd.n4756 242.672
R6122 gnd.n4783 gnd.n4756 242.672
R6123 gnd.n4791 gnd.n4756 242.672
R6124 gnd.n4793 gnd.n4756 242.672
R6125 gnd.n4801 gnd.n4756 242.672
R6126 gnd.n4803 gnd.n4756 242.672
R6127 gnd.n4811 gnd.n4756 242.672
R6128 gnd.n4813 gnd.n4756 242.672
R6129 gnd.n4821 gnd.n4756 242.672
R6130 gnd.n1364 gnd.n1351 242.672
R6131 gnd.n5628 gnd.n1364 242.672
R6132 gnd.n5625 gnd.n1364 242.672
R6133 gnd.n5622 gnd.n1364 242.672
R6134 gnd.n5611 gnd.n1364 242.672
R6135 gnd.n5602 gnd.n1364 242.672
R6136 gnd.n5599 gnd.n1364 242.672
R6137 gnd.n5588 gnd.n1364 242.672
R6138 gnd.n5577 gnd.n1364 242.672
R6139 gnd.n7046 gnd.n508 242.672
R6140 gnd.n7046 gnd.n509 242.672
R6141 gnd.n7046 gnd.n510 242.672
R6142 gnd.n7046 gnd.n511 242.672
R6143 gnd.n7046 gnd.n512 242.672
R6144 gnd.n7046 gnd.n513 242.672
R6145 gnd.n7046 gnd.n514 242.672
R6146 gnd.n7046 gnd.n515 242.672
R6147 gnd.n7046 gnd.n516 242.672
R6148 gnd.n124 gnd.n121 242.672
R6149 gnd.n7447 gnd.n124 242.672
R6150 gnd.n7443 gnd.n124 242.672
R6151 gnd.n7440 gnd.n124 242.672
R6152 gnd.n7435 gnd.n124 242.672
R6153 gnd.n7432 gnd.n124 242.672
R6154 gnd.n7427 gnd.n124 242.672
R6155 gnd.n7424 gnd.n124 242.672
R6156 gnd.n7419 gnd.n124 242.672
R6157 gnd.n3966 gnd.n3965 242.672
R6158 gnd.n3966 gnd.n3876 242.672
R6159 gnd.n3966 gnd.n3877 242.672
R6160 gnd.n3966 gnd.n3878 242.672
R6161 gnd.n3966 gnd.n3879 242.672
R6162 gnd.n3966 gnd.n3880 242.672
R6163 gnd.n3966 gnd.n3881 242.672
R6164 gnd.n3966 gnd.n3882 242.672
R6165 gnd.n3966 gnd.n3883 242.672
R6166 gnd.n3966 gnd.n3884 242.672
R6167 gnd.n3966 gnd.n3885 242.672
R6168 gnd.n3966 gnd.n3886 242.672
R6169 gnd.n3967 gnd.n3966 242.672
R6170 gnd.n4755 gnd.n2002 242.672
R6171 gnd.n4755 gnd.n2001 242.672
R6172 gnd.n4755 gnd.n2000 242.672
R6173 gnd.n4755 gnd.n1999 242.672
R6174 gnd.n4755 gnd.n1998 242.672
R6175 gnd.n4755 gnd.n1997 242.672
R6176 gnd.n4755 gnd.n1996 242.672
R6177 gnd.n4755 gnd.n1995 242.672
R6178 gnd.n4755 gnd.n1994 242.672
R6179 gnd.n4755 gnd.n1993 242.672
R6180 gnd.n4755 gnd.n1992 242.672
R6181 gnd.n4755 gnd.n1991 242.672
R6182 gnd.n4755 gnd.n1990 242.672
R6183 gnd.n4050 gnd.n4049 242.672
R6184 gnd.n4049 gnd.n3788 242.672
R6185 gnd.n4049 gnd.n3789 242.672
R6186 gnd.n4049 gnd.n3790 242.672
R6187 gnd.n4049 gnd.n3791 242.672
R6188 gnd.n4049 gnd.n3792 242.672
R6189 gnd.n4049 gnd.n3793 242.672
R6190 gnd.n4049 gnd.n3794 242.672
R6191 gnd.n4755 gnd.n2003 242.672
R6192 gnd.n4755 gnd.n2004 242.672
R6193 gnd.n4755 gnd.n2005 242.672
R6194 gnd.n4755 gnd.n2006 242.672
R6195 gnd.n4755 gnd.n2007 242.672
R6196 gnd.n4755 gnd.n2008 242.672
R6197 gnd.n4755 gnd.n2009 242.672
R6198 gnd.n4755 gnd.n2010 242.672
R6199 gnd.n5062 gnd.n4756 242.672
R6200 gnd.n4876 gnd.n4756 242.672
R6201 gnd.n5055 gnd.n4756 242.672
R6202 gnd.n5049 gnd.n4756 242.672
R6203 gnd.n5047 gnd.n4756 242.672
R6204 gnd.n5041 gnd.n4756 242.672
R6205 gnd.n5039 gnd.n4756 242.672
R6206 gnd.n5033 gnd.n4756 242.672
R6207 gnd.n5031 gnd.n4756 242.672
R6208 gnd.n5025 gnd.n4756 242.672
R6209 gnd.n5023 gnd.n4756 242.672
R6210 gnd.n5017 gnd.n4756 242.672
R6211 gnd.n5015 gnd.n4756 242.672
R6212 gnd.n5009 gnd.n4756 242.672
R6213 gnd.n5007 gnd.n4756 242.672
R6214 gnd.n5001 gnd.n4756 242.672
R6215 gnd.n4999 gnd.n4756 242.672
R6216 gnd.n4930 gnd.n4756 242.672
R6217 gnd.n4989 gnd.n4756 242.672
R6218 gnd.n5702 gnd.n1364 242.672
R6219 gnd.n1644 gnd.n1364 242.672
R6220 gnd.n5709 gnd.n1364 242.672
R6221 gnd.n1635 gnd.n1364 242.672
R6222 gnd.n5716 gnd.n1364 242.672
R6223 gnd.n1628 gnd.n1364 242.672
R6224 gnd.n5723 gnd.n1364 242.672
R6225 gnd.n1621 gnd.n1364 242.672
R6226 gnd.n5730 gnd.n1364 242.672
R6227 gnd.n1614 gnd.n1364 242.672
R6228 gnd.n5737 gnd.n1364 242.672
R6229 gnd.n5738 gnd.n1606 242.672
R6230 gnd.n5739 gnd.n1364 242.672
R6231 gnd.n1387 gnd.n1364 242.672
R6232 gnd.n5746 gnd.n1364 242.672
R6233 gnd.n1380 gnd.n1364 242.672
R6234 gnd.n5753 gnd.n1364 242.672
R6235 gnd.n1373 gnd.n1364 242.672
R6236 gnd.n5760 gnd.n1364 242.672
R6237 gnd.n5763 gnd.n1364 242.672
R6238 gnd.n7047 gnd.n7046 242.672
R6239 gnd.n7046 gnd.n490 242.672
R6240 gnd.n7046 gnd.n491 242.672
R6241 gnd.n7046 gnd.n492 242.672
R6242 gnd.n7046 gnd.n493 242.672
R6243 gnd.n7046 gnd.n494 242.672
R6244 gnd.n7046 gnd.n495 242.672
R6245 gnd.n7046 gnd.n496 242.672
R6246 gnd.n7018 gnd.n535 242.672
R6247 gnd.n7046 gnd.n497 242.672
R6248 gnd.n7046 gnd.n498 242.672
R6249 gnd.n7046 gnd.n499 242.672
R6250 gnd.n7046 gnd.n500 242.672
R6251 gnd.n7046 gnd.n501 242.672
R6252 gnd.n7046 gnd.n502 242.672
R6253 gnd.n7046 gnd.n503 242.672
R6254 gnd.n7046 gnd.n504 242.672
R6255 gnd.n7046 gnd.n505 242.672
R6256 gnd.n7046 gnd.n506 242.672
R6257 gnd.n7046 gnd.n507 242.672
R6258 gnd.n194 gnd.n124 242.672
R6259 gnd.n7504 gnd.n124 242.672
R6260 gnd.n190 gnd.n124 242.672
R6261 gnd.n7511 gnd.n124 242.672
R6262 gnd.n183 gnd.n124 242.672
R6263 gnd.n7518 gnd.n124 242.672
R6264 gnd.n176 gnd.n124 242.672
R6265 gnd.n7525 gnd.n124 242.672
R6266 gnd.n169 gnd.n124 242.672
R6267 gnd.n7532 gnd.n124 242.672
R6268 gnd.n162 gnd.n124 242.672
R6269 gnd.n7542 gnd.n124 242.672
R6270 gnd.n155 gnd.n124 242.672
R6271 gnd.n7549 gnd.n124 242.672
R6272 gnd.n148 gnd.n124 242.672
R6273 gnd.n7556 gnd.n124 242.672
R6274 gnd.n141 gnd.n124 242.672
R6275 gnd.n7563 gnd.n124 242.672
R6276 gnd.n134 gnd.n124 242.672
R6277 gnd.n5809 gnd.n1319 242.672
R6278 gnd.n5809 gnd.n1320 242.672
R6279 gnd.n5809 gnd.n1321 242.672
R6280 gnd.n5809 gnd.n1322 242.672
R6281 gnd.n5809 gnd.n1323 242.672
R6282 gnd.n5809 gnd.n1324 242.672
R6283 gnd.n5809 gnd.n1325 242.672
R6284 gnd.n5809 gnd.n1326 242.672
R6285 gnd.n5809 gnd.n1327 242.672
R6286 gnd.n5809 gnd.n1328 242.672
R6287 gnd.n5809 gnd.n1329 242.672
R6288 gnd.n5809 gnd.n1330 242.672
R6289 gnd.n5809 gnd.n1331 242.672
R6290 gnd.n5809 gnd.n5808 242.672
R6291 gnd.n6817 gnd.n630 242.672
R6292 gnd.n6817 gnd.n629 242.672
R6293 gnd.n6817 gnd.n628 242.672
R6294 gnd.n6817 gnd.n627 242.672
R6295 gnd.n6817 gnd.n626 242.672
R6296 gnd.n6817 gnd.n625 242.672
R6297 gnd.n6817 gnd.n624 242.672
R6298 gnd.n6817 gnd.n623 242.672
R6299 gnd.n6817 gnd.n622 242.672
R6300 gnd.n6817 gnd.n621 242.672
R6301 gnd.n6817 gnd.n620 242.672
R6302 gnd.n6817 gnd.n619 242.672
R6303 gnd.n6817 gnd.n618 242.672
R6304 gnd.n6817 gnd.n617 242.672
R6305 gnd.n131 gnd.n127 240.244
R6306 gnd.n7565 gnd.n7564 240.244
R6307 gnd.n7562 gnd.n135 240.244
R6308 gnd.n7558 gnd.n7557 240.244
R6309 gnd.n7555 gnd.n142 240.244
R6310 gnd.n7551 gnd.n7550 240.244
R6311 gnd.n7548 gnd.n149 240.244
R6312 gnd.n7544 gnd.n7543 240.244
R6313 gnd.n7541 gnd.n156 240.244
R6314 gnd.n7534 gnd.n7533 240.244
R6315 gnd.n7531 gnd.n163 240.244
R6316 gnd.n7527 gnd.n7526 240.244
R6317 gnd.n7524 gnd.n170 240.244
R6318 gnd.n7520 gnd.n7519 240.244
R6319 gnd.n7517 gnd.n177 240.244
R6320 gnd.n7513 gnd.n7512 240.244
R6321 gnd.n7510 gnd.n184 240.244
R6322 gnd.n7506 gnd.n7505 240.244
R6323 gnd.n7503 gnd.n191 240.244
R6324 gnd.n6975 gnd.n481 240.244
R6325 gnd.n6847 gnd.n481 240.244
R6326 gnd.n6847 gnd.n472 240.244
R6327 gnd.n6851 gnd.n472 240.244
R6328 gnd.n6851 gnd.n463 240.244
R6329 gnd.n6864 gnd.n463 240.244
R6330 gnd.n6864 gnd.n454 240.244
R6331 gnd.n6860 gnd.n454 240.244
R6332 gnd.n6860 gnd.n447 240.244
R6333 gnd.n6887 gnd.n447 240.244
R6334 gnd.n6887 gnd.n438 240.244
R6335 gnd.n6891 gnd.n438 240.244
R6336 gnd.n6891 gnd.n429 240.244
R6337 gnd.n6903 gnd.n429 240.244
R6338 gnd.n6903 gnd.n420 240.244
R6339 gnd.n6899 gnd.n420 240.244
R6340 gnd.n6899 gnd.n413 240.244
R6341 gnd.n6918 gnd.n413 240.244
R6342 gnd.n6918 gnd.n402 240.244
R6343 gnd.n6937 gnd.n402 240.244
R6344 gnd.n6937 gnd.n394 240.244
R6345 gnd.n394 gnd.n387 240.244
R6346 gnd.n387 gnd.n370 240.244
R6347 gnd.n6931 gnd.n370 240.244
R6348 gnd.n6931 gnd.n358 240.244
R6349 gnd.n7191 gnd.n358 240.244
R6350 gnd.n7192 gnd.n7191 240.244
R6351 gnd.n7192 gnd.n350 240.244
R6352 gnd.n350 gnd.n309 240.244
R6353 gnd.n7201 gnd.n309 240.244
R6354 gnd.n7201 gnd.n339 240.244
R6355 gnd.n339 gnd.n335 240.244
R6356 gnd.n7229 gnd.n335 240.244
R6357 gnd.n7229 gnd.n331 240.244
R6358 gnd.n7300 gnd.n331 240.244
R6359 gnd.n7300 gnd.n324 240.244
R6360 gnd.n7296 gnd.n324 240.244
R6361 gnd.n7296 gnd.n296 240.244
R6362 gnd.n7293 gnd.n296 240.244
R6363 gnd.n7293 gnd.n287 240.244
R6364 gnd.n7290 gnd.n287 240.244
R6365 gnd.n7290 gnd.n279 240.244
R6366 gnd.n7287 gnd.n279 240.244
R6367 gnd.n7287 gnd.n272 240.244
R6368 gnd.n7284 gnd.n272 240.244
R6369 gnd.n7284 gnd.n266 240.244
R6370 gnd.n7281 gnd.n266 240.244
R6371 gnd.n7281 gnd.n257 240.244
R6372 gnd.n7278 gnd.n257 240.244
R6373 gnd.n7278 gnd.n249 240.244
R6374 gnd.n7275 gnd.n249 240.244
R6375 gnd.n7275 gnd.n242 240.244
R6376 gnd.n7272 gnd.n242 240.244
R6377 gnd.n7272 gnd.n235 240.244
R6378 gnd.n7269 gnd.n235 240.244
R6379 gnd.n7269 gnd.n226 240.244
R6380 gnd.n7266 gnd.n226 240.244
R6381 gnd.n7266 gnd.n219 240.244
R6382 gnd.n7263 gnd.n219 240.244
R6383 gnd.n7263 gnd.n210 240.244
R6384 gnd.n210 gnd.n201 240.244
R6385 gnd.n7494 gnd.n201 240.244
R6386 gnd.n7495 gnd.n7494 240.244
R6387 gnd.n7495 gnd.n123 240.244
R6388 gnd.n7045 gnd.n488 240.244
R6389 gnd.n7045 gnd.n519 240.244
R6390 gnd.n7041 gnd.n7040 240.244
R6391 gnd.n7037 gnd.n7036 240.244
R6392 gnd.n7033 gnd.n7032 240.244
R6393 gnd.n7029 gnd.n7028 240.244
R6394 gnd.n7025 gnd.n7024 240.244
R6395 gnd.n7021 gnd.n7020 240.244
R6396 gnd.n7016 gnd.n7015 240.244
R6397 gnd.n7012 gnd.n7011 240.244
R6398 gnd.n7008 gnd.n7007 240.244
R6399 gnd.n7004 gnd.n7003 240.244
R6400 gnd.n7000 gnd.n6999 240.244
R6401 gnd.n6996 gnd.n6995 240.244
R6402 gnd.n6992 gnd.n6991 240.244
R6403 gnd.n6988 gnd.n6987 240.244
R6404 gnd.n6984 gnd.n6983 240.244
R6405 gnd.n558 gnd.n557 240.244
R6406 gnd.n7054 gnd.n484 240.244
R6407 gnd.n7054 gnd.n470 240.244
R6408 gnd.n7064 gnd.n470 240.244
R6409 gnd.n7064 gnd.n466 240.244
R6410 gnd.n7070 gnd.n466 240.244
R6411 gnd.n7070 gnd.n453 240.244
R6412 gnd.n7080 gnd.n453 240.244
R6413 gnd.n7080 gnd.n449 240.244
R6414 gnd.n7086 gnd.n449 240.244
R6415 gnd.n7086 gnd.n436 240.244
R6416 gnd.n7096 gnd.n436 240.244
R6417 gnd.n7096 gnd.n432 240.244
R6418 gnd.n7102 gnd.n432 240.244
R6419 gnd.n7102 gnd.n419 240.244
R6420 gnd.n7112 gnd.n419 240.244
R6421 gnd.n7112 gnd.n415 240.244
R6422 gnd.n7118 gnd.n415 240.244
R6423 gnd.n7118 gnd.n400 240.244
R6424 gnd.n7131 gnd.n400 240.244
R6425 gnd.n7131 gnd.n396 240.244
R6426 gnd.n7137 gnd.n396 240.244
R6427 gnd.n7137 gnd.n368 240.244
R6428 gnd.n7182 gnd.n368 240.244
R6429 gnd.n7182 gnd.n369 240.244
R6430 gnd.n369 gnd.n363 240.244
R6431 gnd.n7189 gnd.n363 240.244
R6432 gnd.n7189 gnd.n364 240.244
R6433 gnd.n364 gnd.n306 240.244
R6434 gnd.n7321 gnd.n306 240.244
R6435 gnd.n7321 gnd.n307 240.244
R6436 gnd.n7223 gnd.n307 240.244
R6437 gnd.n7224 gnd.n7223 240.244
R6438 gnd.n7227 gnd.n7224 240.244
R6439 gnd.n7227 gnd.n326 240.244
R6440 gnd.n7302 gnd.n326 240.244
R6441 gnd.n7304 gnd.n7302 240.244
R6442 gnd.n7304 gnd.n297 240.244
R6443 gnd.n7328 gnd.n297 240.244
R6444 gnd.n7328 gnd.n285 240.244
R6445 gnd.n7338 gnd.n285 240.244
R6446 gnd.n7338 gnd.n281 240.244
R6447 gnd.n7344 gnd.n281 240.244
R6448 gnd.n7344 gnd.n271 240.244
R6449 gnd.n7354 gnd.n271 240.244
R6450 gnd.n7354 gnd.n267 240.244
R6451 gnd.n7360 gnd.n267 240.244
R6452 gnd.n7360 gnd.n255 240.244
R6453 gnd.n7370 gnd.n255 240.244
R6454 gnd.n7370 gnd.n251 240.244
R6455 gnd.n7376 gnd.n251 240.244
R6456 gnd.n7376 gnd.n241 240.244
R6457 gnd.n7386 gnd.n241 240.244
R6458 gnd.n7386 gnd.n237 240.244
R6459 gnd.n7392 gnd.n237 240.244
R6460 gnd.n7392 gnd.n224 240.244
R6461 gnd.n7402 gnd.n224 240.244
R6462 gnd.n7402 gnd.n220 240.244
R6463 gnd.n7408 gnd.n220 240.244
R6464 gnd.n7408 gnd.n208 240.244
R6465 gnd.n7486 gnd.n208 240.244
R6466 gnd.n7486 gnd.n204 240.244
R6467 gnd.n7492 gnd.n204 240.244
R6468 gnd.n7492 gnd.n126 240.244
R6469 gnd.n7572 gnd.n126 240.244
R6470 gnd.n5764 gnd.n1359 240.244
R6471 gnd.n5762 gnd.n5761 240.244
R6472 gnd.n5759 gnd.n1366 240.244
R6473 gnd.n5755 gnd.n5754 240.244
R6474 gnd.n5752 gnd.n1374 240.244
R6475 gnd.n5748 gnd.n5747 240.244
R6476 gnd.n5745 gnd.n1381 240.244
R6477 gnd.n5741 gnd.n5740 240.244
R6478 gnd.n5736 gnd.n1607 240.244
R6479 gnd.n5732 gnd.n5731 240.244
R6480 gnd.n5729 gnd.n1615 240.244
R6481 gnd.n5725 gnd.n5724 240.244
R6482 gnd.n5722 gnd.n1622 240.244
R6483 gnd.n5718 gnd.n5717 240.244
R6484 gnd.n5715 gnd.n1629 240.244
R6485 gnd.n5711 gnd.n5710 240.244
R6486 gnd.n5708 gnd.n1636 240.244
R6487 gnd.n5704 gnd.n5703 240.244
R6488 gnd.n4936 gnd.n4757 240.244
R6489 gnd.n4936 gnd.n1982 240.244
R6490 gnd.n4982 gnd.n1982 240.244
R6491 gnd.n4982 gnd.n1975 240.244
R6492 gnd.n4979 gnd.n1975 240.244
R6493 gnd.n4979 gnd.n1967 240.244
R6494 gnd.n4976 gnd.n1967 240.244
R6495 gnd.n4976 gnd.n1958 240.244
R6496 gnd.n4973 gnd.n1958 240.244
R6497 gnd.n4973 gnd.n1950 240.244
R6498 gnd.n4970 gnd.n1950 240.244
R6499 gnd.n4970 gnd.n1943 240.244
R6500 gnd.n4967 gnd.n1943 240.244
R6501 gnd.n4967 gnd.n1935 240.244
R6502 gnd.n4964 gnd.n1935 240.244
R6503 gnd.n4964 gnd.n1926 240.244
R6504 gnd.n4961 gnd.n1926 240.244
R6505 gnd.n4961 gnd.n1917 240.244
R6506 gnd.n4958 gnd.n1917 240.244
R6507 gnd.n4958 gnd.n1909 240.244
R6508 gnd.n1909 gnd.n1901 240.244
R6509 gnd.n5174 gnd.n1901 240.244
R6510 gnd.n5174 gnd.n1882 240.244
R6511 gnd.n1897 gnd.n1882 240.244
R6512 gnd.n5183 gnd.n1897 240.244
R6513 gnd.n5183 gnd.n1873 240.244
R6514 gnd.n1873 gnd.n1866 240.244
R6515 gnd.n5218 gnd.n1866 240.244
R6516 gnd.n5218 gnd.n1773 240.244
R6517 gnd.n5223 gnd.n1773 240.244
R6518 gnd.n5223 gnd.n1784 240.244
R6519 gnd.n5226 gnd.n1784 240.244
R6520 gnd.n5226 gnd.n1789 240.244
R6521 gnd.n5232 gnd.n1789 240.244
R6522 gnd.n5232 gnd.n1796 240.244
R6523 gnd.n5242 gnd.n1796 240.244
R6524 gnd.n5242 gnd.n1759 240.244
R6525 gnd.n1806 gnd.n1759 240.244
R6526 gnd.n1806 gnd.n1750 240.244
R6527 gnd.n5250 gnd.n1750 240.244
R6528 gnd.n5250 gnd.n1743 240.244
R6529 gnd.n5277 gnd.n1743 240.244
R6530 gnd.n5277 gnd.n1734 240.244
R6531 gnd.n5281 gnd.n1734 240.244
R6532 gnd.n5281 gnd.n1725 240.244
R6533 gnd.n5294 gnd.n1725 240.244
R6534 gnd.n5294 gnd.n1716 240.244
R6535 gnd.n5290 gnd.n1716 240.244
R6536 gnd.n5290 gnd.n1709 240.244
R6537 gnd.n5317 gnd.n1709 240.244
R6538 gnd.n5317 gnd.n1700 240.244
R6539 gnd.n5321 gnd.n1700 240.244
R6540 gnd.n5321 gnd.n1691 240.244
R6541 gnd.n5333 gnd.n1691 240.244
R6542 gnd.n5333 gnd.n1682 240.244
R6543 gnd.n5329 gnd.n1682 240.244
R6544 gnd.n5329 gnd.n1675 240.244
R6545 gnd.n5374 gnd.n1675 240.244
R6546 gnd.n5374 gnd.n1666 240.244
R6547 gnd.n5383 gnd.n1666 240.244
R6548 gnd.n5383 gnd.n1656 240.244
R6549 gnd.n1656 gnd.n1648 240.244
R6550 gnd.n5695 gnd.n1648 240.244
R6551 gnd.n5695 gnd.n1355 240.244
R6552 gnd.n5063 gnd.n5061 240.244
R6553 gnd.n5061 gnd.n5060 240.244
R6554 gnd.n5057 gnd.n5056 240.244
R6555 gnd.n5054 gnd.n4881 240.244
R6556 gnd.n5050 gnd.n5048 240.244
R6557 gnd.n5046 gnd.n4887 240.244
R6558 gnd.n5042 gnd.n5040 240.244
R6559 gnd.n5038 gnd.n4893 240.244
R6560 gnd.n5034 gnd.n5032 240.244
R6561 gnd.n5030 gnd.n4899 240.244
R6562 gnd.n5026 gnd.n5024 240.244
R6563 gnd.n5022 gnd.n4908 240.244
R6564 gnd.n5018 gnd.n5016 240.244
R6565 gnd.n5014 gnd.n4914 240.244
R6566 gnd.n5010 gnd.n5008 240.244
R6567 gnd.n5006 gnd.n4920 240.244
R6568 gnd.n5002 gnd.n5000 240.244
R6569 gnd.n4998 gnd.n4926 240.244
R6570 gnd.n4988 gnd.n4931 240.244
R6571 gnd.n5069 gnd.n1981 240.244
R6572 gnd.n5079 gnd.n1981 240.244
R6573 gnd.n5079 gnd.n1977 240.244
R6574 gnd.n5085 gnd.n1977 240.244
R6575 gnd.n5085 gnd.n1965 240.244
R6576 gnd.n5095 gnd.n1965 240.244
R6577 gnd.n5095 gnd.n1961 240.244
R6578 gnd.n5101 gnd.n1961 240.244
R6579 gnd.n5101 gnd.n1949 240.244
R6580 gnd.n5111 gnd.n1949 240.244
R6581 gnd.n5111 gnd.n1945 240.244
R6582 gnd.n5117 gnd.n1945 240.244
R6583 gnd.n5117 gnd.n1933 240.244
R6584 gnd.n5127 gnd.n1933 240.244
R6585 gnd.n5127 gnd.n1929 240.244
R6586 gnd.n5133 gnd.n1929 240.244
R6587 gnd.n5133 gnd.n1916 240.244
R6588 gnd.n5151 gnd.n1916 240.244
R6589 gnd.n5151 gnd.n1911 240.244
R6590 gnd.n5159 gnd.n1911 240.244
R6591 gnd.n5159 gnd.n1912 240.244
R6592 gnd.n1912 gnd.n1880 240.244
R6593 gnd.n5191 gnd.n1880 240.244
R6594 gnd.n5191 gnd.n1881 240.244
R6595 gnd.n1881 gnd.n1875 240.244
R6596 gnd.n5198 gnd.n1875 240.244
R6597 gnd.n5198 gnd.n1876 240.244
R6598 gnd.n1876 gnd.n1771 240.244
R6599 gnd.n5462 gnd.n1771 240.244
R6600 gnd.n5462 gnd.n1772 240.244
R6601 gnd.n5454 gnd.n1772 240.244
R6602 gnd.n5454 gnd.n5451 240.244
R6603 gnd.n5451 gnd.n5448 240.244
R6604 gnd.n5448 gnd.n1787 240.244
R6605 gnd.n5440 gnd.n1787 240.244
R6606 gnd.n5440 gnd.n1762 240.244
R6607 gnd.n5468 gnd.n1762 240.244
R6608 gnd.n5468 gnd.n1749 240.244
R6609 gnd.n5478 gnd.n1749 240.244
R6610 gnd.n5478 gnd.n1745 240.244
R6611 gnd.n5484 gnd.n1745 240.244
R6612 gnd.n5484 gnd.n1732 240.244
R6613 gnd.n5494 gnd.n1732 240.244
R6614 gnd.n5494 gnd.n1728 240.244
R6615 gnd.n5500 gnd.n1728 240.244
R6616 gnd.n5500 gnd.n1715 240.244
R6617 gnd.n5510 gnd.n1715 240.244
R6618 gnd.n5510 gnd.n1711 240.244
R6619 gnd.n5516 gnd.n1711 240.244
R6620 gnd.n5516 gnd.n1698 240.244
R6621 gnd.n5526 gnd.n1698 240.244
R6622 gnd.n5526 gnd.n1694 240.244
R6623 gnd.n5532 gnd.n1694 240.244
R6624 gnd.n5532 gnd.n1681 240.244
R6625 gnd.n5542 gnd.n1681 240.244
R6626 gnd.n5542 gnd.n1677 240.244
R6627 gnd.n5548 gnd.n1677 240.244
R6628 gnd.n5548 gnd.n1664 240.244
R6629 gnd.n5558 gnd.n1664 240.244
R6630 gnd.n5558 gnd.n1659 240.244
R6631 gnd.n5566 gnd.n1659 240.244
R6632 gnd.n5566 gnd.n1660 240.244
R6633 gnd.n1660 gnd.n1358 240.244
R6634 gnd.n5770 gnd.n1358 240.244
R6635 gnd.n4754 gnd.n2012 240.244
R6636 gnd.n4747 gnd.n4746 240.244
R6637 gnd.n4744 gnd.n4743 240.244
R6638 gnd.n4740 gnd.n4739 240.244
R6639 gnd.n4736 gnd.n4735 240.244
R6640 gnd.n4732 gnd.n4731 240.244
R6641 gnd.n4728 gnd.n4727 240.244
R6642 gnd.n4724 gnd.n4723 240.244
R6643 gnd.n4061 gnd.n3773 240.244
R6644 gnd.n4071 gnd.n3773 240.244
R6645 gnd.n4071 gnd.n3764 240.244
R6646 gnd.n3764 gnd.n3753 240.244
R6647 gnd.n4092 gnd.n3753 240.244
R6648 gnd.n4092 gnd.n3747 240.244
R6649 gnd.n4102 gnd.n3747 240.244
R6650 gnd.n4102 gnd.n3736 240.244
R6651 gnd.n3736 gnd.n3726 240.244
R6652 gnd.n4128 gnd.n3726 240.244
R6653 gnd.n4129 gnd.n4128 240.244
R6654 gnd.n4130 gnd.n4129 240.244
R6655 gnd.n4130 gnd.n3705 240.244
R6656 gnd.n4166 gnd.n3705 240.244
R6657 gnd.n4166 gnd.n3706 240.244
R6658 gnd.n4162 gnd.n3706 240.244
R6659 gnd.n4162 gnd.n4161 240.244
R6660 gnd.n4161 gnd.n3530 240.244
R6661 gnd.n4196 gnd.n3530 240.244
R6662 gnd.n4196 gnd.n3521 240.244
R6663 gnd.n3521 gnd.n3513 240.244
R6664 gnd.n4217 gnd.n3513 240.244
R6665 gnd.n4217 gnd.n3507 240.244
R6666 gnd.n4227 gnd.n3507 240.244
R6667 gnd.n4227 gnd.n3498 240.244
R6668 gnd.n3498 gnd.n3488 240.244
R6669 gnd.n4248 gnd.n3488 240.244
R6670 gnd.n4248 gnd.n3481 240.244
R6671 gnd.n4258 gnd.n3481 240.244
R6672 gnd.n4258 gnd.n3472 240.244
R6673 gnd.n3472 gnd.n3461 240.244
R6674 gnd.n4279 gnd.n3461 240.244
R6675 gnd.n4279 gnd.n3455 240.244
R6676 gnd.n4289 gnd.n3455 240.244
R6677 gnd.n4289 gnd.n3447 240.244
R6678 gnd.n3447 gnd.n3437 240.244
R6679 gnd.n4310 gnd.n3437 240.244
R6680 gnd.n4310 gnd.n3431 240.244
R6681 gnd.n4320 gnd.n3431 240.244
R6682 gnd.n4320 gnd.n3422 240.244
R6683 gnd.n3422 gnd.n3411 240.244
R6684 gnd.n4341 gnd.n3411 240.244
R6685 gnd.n4341 gnd.n3405 240.244
R6686 gnd.n4351 gnd.n3405 240.244
R6687 gnd.n4351 gnd.n3396 240.244
R6688 gnd.n3396 gnd.n3386 240.244
R6689 gnd.n4372 gnd.n3386 240.244
R6690 gnd.n4372 gnd.n3379 240.244
R6691 gnd.n4638 gnd.n3379 240.244
R6692 gnd.n4638 gnd.n3371 240.244
R6693 gnd.n3371 gnd.n3361 240.244
R6694 gnd.n4658 gnd.n3361 240.244
R6695 gnd.n4658 gnd.n3363 240.244
R6696 gnd.n4051 gnd.n3786 240.244
R6697 gnd.n3807 gnd.n3786 240.244
R6698 gnd.n3810 gnd.n3809 240.244
R6699 gnd.n3817 gnd.n3816 240.244
R6700 gnd.n3820 gnd.n3819 240.244
R6701 gnd.n3827 gnd.n3826 240.244
R6702 gnd.n3830 gnd.n3829 240.244
R6703 gnd.n3837 gnd.n3836 240.244
R6704 gnd.n4059 gnd.n3783 240.244
R6705 gnd.n3783 gnd.n3762 240.244
R6706 gnd.n4082 gnd.n3762 240.244
R6707 gnd.n4082 gnd.n3756 240.244
R6708 gnd.n4090 gnd.n3756 240.244
R6709 gnd.n4090 gnd.n3758 240.244
R6710 gnd.n3758 gnd.n3734 240.244
R6711 gnd.n4112 gnd.n3734 240.244
R6712 gnd.n4112 gnd.n3729 240.244
R6713 gnd.n4126 gnd.n3729 240.244
R6714 gnd.n4126 gnd.n3730 240.244
R6715 gnd.n4122 gnd.n3730 240.244
R6716 gnd.n4122 gnd.n3702 240.244
R6717 gnd.n4169 gnd.n3702 240.244
R6718 gnd.n4170 gnd.n4169 240.244
R6719 gnd.n4171 gnd.n4170 240.244
R6720 gnd.n4171 gnd.n3698 240.244
R6721 gnd.n4177 gnd.n3698 240.244
R6722 gnd.n4177 gnd.n3520 240.244
R6723 gnd.n4207 gnd.n3520 240.244
R6724 gnd.n4207 gnd.n3515 240.244
R6725 gnd.n4215 gnd.n3515 240.244
R6726 gnd.n4215 gnd.n3516 240.244
R6727 gnd.n3516 gnd.n3496 240.244
R6728 gnd.n4238 gnd.n3496 240.244
R6729 gnd.n4238 gnd.n3491 240.244
R6730 gnd.n4246 gnd.n3491 240.244
R6731 gnd.n4246 gnd.n3492 240.244
R6732 gnd.n3492 gnd.n3470 240.244
R6733 gnd.n4269 gnd.n3470 240.244
R6734 gnd.n4269 gnd.n3464 240.244
R6735 gnd.n4277 gnd.n3464 240.244
R6736 gnd.n4277 gnd.n3466 240.244
R6737 gnd.n3466 gnd.n3445 240.244
R6738 gnd.n4300 gnd.n3445 240.244
R6739 gnd.n4300 gnd.n3439 240.244
R6740 gnd.n4308 gnd.n3439 240.244
R6741 gnd.n4308 gnd.n3441 240.244
R6742 gnd.n3441 gnd.n3420 240.244
R6743 gnd.n4331 gnd.n3420 240.244
R6744 gnd.n4331 gnd.n3414 240.244
R6745 gnd.n4339 gnd.n3414 240.244
R6746 gnd.n4339 gnd.n3416 240.244
R6747 gnd.n3416 gnd.n3394 240.244
R6748 gnd.n4362 gnd.n3394 240.244
R6749 gnd.n4362 gnd.n3389 240.244
R6750 gnd.n4370 gnd.n3389 240.244
R6751 gnd.n4370 gnd.n3390 240.244
R6752 gnd.n3390 gnd.n3369 240.244
R6753 gnd.n4648 gnd.n3369 240.244
R6754 gnd.n4648 gnd.n3365 240.244
R6755 gnd.n4656 gnd.n3365 240.244
R6756 gnd.n4656 gnd.n2011 240.244
R6757 gnd.n2031 gnd.n1989 240.244
R6758 gnd.n4714 gnd.n4713 240.244
R6759 gnd.n4710 gnd.n4709 240.244
R6760 gnd.n4706 gnd.n4705 240.244
R6761 gnd.n4702 gnd.n4701 240.244
R6762 gnd.n4698 gnd.n4697 240.244
R6763 gnd.n4694 gnd.n4693 240.244
R6764 gnd.n4690 gnd.n4689 240.244
R6765 gnd.n4686 gnd.n4685 240.244
R6766 gnd.n4682 gnd.n4681 240.244
R6767 gnd.n4678 gnd.n4677 240.244
R6768 gnd.n4674 gnd.n4673 240.244
R6769 gnd.n4670 gnd.n4669 240.244
R6770 gnd.n3974 gnd.n3871 240.244
R6771 gnd.n3974 gnd.n3864 240.244
R6772 gnd.n3985 gnd.n3864 240.244
R6773 gnd.n3985 gnd.n3860 240.244
R6774 gnd.n3991 gnd.n3860 240.244
R6775 gnd.n3991 gnd.n3852 240.244
R6776 gnd.n4001 gnd.n3852 240.244
R6777 gnd.n4001 gnd.n3847 240.244
R6778 gnd.n4037 gnd.n3847 240.244
R6779 gnd.n4037 gnd.n3848 240.244
R6780 gnd.n3848 gnd.n3795 240.244
R6781 gnd.n4032 gnd.n3795 240.244
R6782 gnd.n4032 gnd.n4031 240.244
R6783 gnd.n4031 gnd.n3774 240.244
R6784 gnd.n4027 gnd.n3774 240.244
R6785 gnd.n4027 gnd.n3765 240.244
R6786 gnd.n4024 gnd.n3765 240.244
R6787 gnd.n4024 gnd.n4023 240.244
R6788 gnd.n4023 gnd.n3748 240.244
R6789 gnd.n4019 gnd.n3748 240.244
R6790 gnd.n4019 gnd.n3737 240.244
R6791 gnd.n3737 gnd.n3717 240.244
R6792 gnd.n4138 gnd.n3717 240.244
R6793 gnd.n4138 gnd.n3712 240.244
R6794 gnd.n4146 gnd.n3712 240.244
R6795 gnd.n4146 gnd.n3713 240.244
R6796 gnd.n3713 gnd.n3681 240.244
R6797 gnd.n4186 gnd.n3681 240.244
R6798 gnd.n4186 gnd.n3682 240.244
R6799 gnd.n3697 gnd.n3682 240.244
R6800 gnd.n3697 gnd.n3532 240.244
R6801 gnd.n4193 gnd.n3532 240.244
R6802 gnd.n4193 gnd.n3522 240.244
R6803 gnd.n3611 gnd.n3522 240.244
R6804 gnd.n3614 gnd.n3611 240.244
R6805 gnd.n3614 gnd.n3508 240.244
R6806 gnd.n3608 gnd.n3508 240.244
R6807 gnd.n3608 gnd.n3499 240.244
R6808 gnd.n3605 gnd.n3499 240.244
R6809 gnd.n3605 gnd.n3604 240.244
R6810 gnd.n3604 gnd.n3483 240.244
R6811 gnd.n3600 gnd.n3483 240.244
R6812 gnd.n3600 gnd.n3473 240.244
R6813 gnd.n3597 gnd.n3473 240.244
R6814 gnd.n3597 gnd.n3596 240.244
R6815 gnd.n3596 gnd.n3456 240.244
R6816 gnd.n3592 gnd.n3456 240.244
R6817 gnd.n3592 gnd.n3448 240.244
R6818 gnd.n3589 gnd.n3448 240.244
R6819 gnd.n3589 gnd.n3586 240.244
R6820 gnd.n3586 gnd.n3432 240.244
R6821 gnd.n3582 gnd.n3432 240.244
R6822 gnd.n3582 gnd.n3423 240.244
R6823 gnd.n3579 gnd.n3423 240.244
R6824 gnd.n3579 gnd.n3578 240.244
R6825 gnd.n3578 gnd.n3406 240.244
R6826 gnd.n3574 gnd.n3406 240.244
R6827 gnd.n3574 gnd.n3397 240.244
R6828 gnd.n3571 gnd.n3397 240.244
R6829 gnd.n3571 gnd.n3570 240.244
R6830 gnd.n3570 gnd.n3381 240.244
R6831 gnd.n3566 gnd.n3381 240.244
R6832 gnd.n3566 gnd.n3372 240.244
R6833 gnd.n3372 gnd.n2060 240.244
R6834 gnd.n4665 gnd.n2060 240.244
R6835 gnd.n3888 gnd.n3887 240.244
R6836 gnd.n3959 gnd.n3887 240.244
R6837 gnd.n3957 gnd.n3956 240.244
R6838 gnd.n3953 gnd.n3952 240.244
R6839 gnd.n3949 gnd.n3948 240.244
R6840 gnd.n3945 gnd.n3944 240.244
R6841 gnd.n3941 gnd.n3940 240.244
R6842 gnd.n3937 gnd.n3936 240.244
R6843 gnd.n3933 gnd.n3932 240.244
R6844 gnd.n3929 gnd.n3928 240.244
R6845 gnd.n3925 gnd.n3924 240.244
R6846 gnd.n3921 gnd.n3920 240.244
R6847 gnd.n3917 gnd.n3875 240.244
R6848 gnd.n3977 gnd.n3869 240.244
R6849 gnd.n3977 gnd.n3865 240.244
R6850 gnd.n3983 gnd.n3865 240.244
R6851 gnd.n3983 gnd.n3858 240.244
R6852 gnd.n3993 gnd.n3858 240.244
R6853 gnd.n3993 gnd.n3854 240.244
R6854 gnd.n3999 gnd.n3854 240.244
R6855 gnd.n3999 gnd.n3845 240.244
R6856 gnd.n4039 gnd.n3845 240.244
R6857 gnd.n4039 gnd.n3796 240.244
R6858 gnd.n4047 gnd.n3796 240.244
R6859 gnd.n4047 gnd.n3797 240.244
R6860 gnd.n3797 gnd.n3775 240.244
R6861 gnd.n4068 gnd.n3775 240.244
R6862 gnd.n4068 gnd.n3767 240.244
R6863 gnd.n4079 gnd.n3767 240.244
R6864 gnd.n4079 gnd.n3768 240.244
R6865 gnd.n3768 gnd.n3749 240.244
R6866 gnd.n4099 gnd.n3749 240.244
R6867 gnd.n4099 gnd.n3739 240.244
R6868 gnd.n4109 gnd.n3739 240.244
R6869 gnd.n4109 gnd.n3720 240.244
R6870 gnd.n4136 gnd.n3720 240.244
R6871 gnd.n4136 gnd.n3710 240.244
R6872 gnd.n4149 gnd.n3710 240.244
R6873 gnd.n4150 gnd.n4149 240.244
R6874 gnd.n4150 gnd.n3685 240.244
R6875 gnd.n4184 gnd.n3685 240.244
R6876 gnd.n4184 gnd.n3686 240.244
R6877 gnd.n4180 gnd.n3686 240.244
R6878 gnd.n4180 gnd.n3694 240.244
R6879 gnd.n3694 gnd.n3524 240.244
R6880 gnd.n4204 gnd.n3524 240.244
R6881 gnd.n4204 gnd.n3525 240.244
R6882 gnd.n3525 gnd.n3509 240.244
R6883 gnd.n4224 gnd.n3509 240.244
R6884 gnd.n4224 gnd.n3501 240.244
R6885 gnd.n4235 gnd.n3501 240.244
R6886 gnd.n4235 gnd.n3502 240.244
R6887 gnd.n3502 gnd.n3484 240.244
R6888 gnd.n4255 gnd.n3484 240.244
R6889 gnd.n4255 gnd.n3475 240.244
R6890 gnd.n4266 gnd.n3475 240.244
R6891 gnd.n4266 gnd.n3476 240.244
R6892 gnd.n3476 gnd.n3457 240.244
R6893 gnd.n4286 gnd.n3457 240.244
R6894 gnd.n4286 gnd.n3449 240.244
R6895 gnd.n4297 gnd.n3449 240.244
R6896 gnd.n4297 gnd.n3450 240.244
R6897 gnd.n3450 gnd.n3433 240.244
R6898 gnd.n4317 gnd.n3433 240.244
R6899 gnd.n4317 gnd.n3425 240.244
R6900 gnd.n4328 gnd.n3425 240.244
R6901 gnd.n4328 gnd.n3426 240.244
R6902 gnd.n3426 gnd.n3407 240.244
R6903 gnd.n4348 gnd.n3407 240.244
R6904 gnd.n4348 gnd.n3399 240.244
R6905 gnd.n4359 gnd.n3399 240.244
R6906 gnd.n4359 gnd.n3400 240.244
R6907 gnd.n3400 gnd.n3382 240.244
R6908 gnd.n4635 gnd.n3382 240.244
R6909 gnd.n4635 gnd.n3374 240.244
R6910 gnd.n4645 gnd.n3374 240.244
R6911 gnd.n4645 gnd.n3356 240.244
R6912 gnd.n4663 gnd.n3356 240.244
R6913 gnd.n7418 gnd.n7417 240.244
R6914 gnd.n7423 gnd.n7420 240.244
R6915 gnd.n7426 gnd.n7425 240.244
R6916 gnd.n7431 gnd.n7428 240.244
R6917 gnd.n7434 gnd.n7433 240.244
R6918 gnd.n7439 gnd.n7436 240.244
R6919 gnd.n7442 gnd.n7441 240.244
R6920 gnd.n7446 gnd.n7444 240.244
R6921 gnd.n7449 gnd.n7448 240.244
R6922 gnd.n6973 gnd.n482 240.244
R6923 gnd.n568 gnd.n482 240.244
R6924 gnd.n568 gnd.n473 240.244
R6925 gnd.n569 gnd.n473 240.244
R6926 gnd.n569 gnd.n464 240.244
R6927 gnd.n572 gnd.n464 240.244
R6928 gnd.n572 gnd.n455 240.244
R6929 gnd.n573 gnd.n455 240.244
R6930 gnd.n573 gnd.n448 240.244
R6931 gnd.n576 gnd.n448 240.244
R6932 gnd.n576 gnd.n439 240.244
R6933 gnd.n577 gnd.n439 240.244
R6934 gnd.n577 gnd.n430 240.244
R6935 gnd.n580 gnd.n430 240.244
R6936 gnd.n580 gnd.n421 240.244
R6937 gnd.n581 gnd.n421 240.244
R6938 gnd.n581 gnd.n414 240.244
R6939 gnd.n584 gnd.n414 240.244
R6940 gnd.n584 gnd.n403 240.244
R6941 gnd.n6939 gnd.n403 240.244
R6942 gnd.n6939 gnd.n385 240.244
R6943 gnd.n7160 gnd.n385 240.244
R6944 gnd.n7160 gnd.n371 240.244
R6945 gnd.n380 gnd.n371 240.244
R6946 gnd.n7168 gnd.n380 240.244
R6947 gnd.n7168 gnd.n360 240.244
R6948 gnd.n360 gnd.n351 240.244
R6949 gnd.n7210 gnd.n351 240.244
R6950 gnd.n7210 gnd.n310 240.244
R6951 gnd.n7203 gnd.n310 240.244
R6952 gnd.n7203 gnd.n341 240.244
R6953 gnd.n341 gnd.n340 240.244
R6954 gnd.n340 gnd.n78 240.244
R6955 gnd.n79 gnd.n78 240.244
R6956 gnd.n80 gnd.n79 240.244
R6957 gnd.n325 gnd.n80 240.244
R6958 gnd.n325 gnd.n83 240.244
R6959 gnd.n84 gnd.n83 240.244
R6960 gnd.n85 gnd.n84 240.244
R6961 gnd.n288 gnd.n85 240.244
R6962 gnd.n288 gnd.n88 240.244
R6963 gnd.n89 gnd.n88 240.244
R6964 gnd.n90 gnd.n89 240.244
R6965 gnd.n273 gnd.n90 240.244
R6966 gnd.n273 gnd.n93 240.244
R6967 gnd.n94 gnd.n93 240.244
R6968 gnd.n95 gnd.n94 240.244
R6969 gnd.n258 gnd.n95 240.244
R6970 gnd.n258 gnd.n98 240.244
R6971 gnd.n99 gnd.n98 240.244
R6972 gnd.n100 gnd.n99 240.244
R6973 gnd.n243 gnd.n100 240.244
R6974 gnd.n243 gnd.n103 240.244
R6975 gnd.n104 gnd.n103 240.244
R6976 gnd.n105 gnd.n104 240.244
R6977 gnd.n227 gnd.n105 240.244
R6978 gnd.n227 gnd.n108 240.244
R6979 gnd.n109 gnd.n108 240.244
R6980 gnd.n110 gnd.n109 240.244
R6981 gnd.n211 gnd.n110 240.244
R6982 gnd.n211 gnd.n113 240.244
R6983 gnd.n114 gnd.n113 240.244
R6984 gnd.n115 gnd.n114 240.244
R6985 gnd.n7574 gnd.n115 240.244
R6986 gnd.n6625 gnd.n6624 240.244
R6987 gnd.n6627 gnd.n6626 240.244
R6988 gnd.n6637 gnd.n6636 240.244
R6989 gnd.n6645 gnd.n6644 240.244
R6990 gnd.n6647 gnd.n6646 240.244
R6991 gnd.n6657 gnd.n6656 240.244
R6992 gnd.n6665 gnd.n6664 240.244
R6993 gnd.n6667 gnd.n6666 240.244
R6994 gnd.n6711 gnd.n517 240.244
R6995 gnd.n7056 gnd.n479 240.244
R6996 gnd.n7056 gnd.n475 240.244
R6997 gnd.n7062 gnd.n475 240.244
R6998 gnd.n7062 gnd.n461 240.244
R6999 gnd.n7072 gnd.n461 240.244
R7000 gnd.n7072 gnd.n457 240.244
R7001 gnd.n7078 gnd.n457 240.244
R7002 gnd.n7078 gnd.n445 240.244
R7003 gnd.n7088 gnd.n445 240.244
R7004 gnd.n7088 gnd.n441 240.244
R7005 gnd.n7094 gnd.n441 240.244
R7006 gnd.n7094 gnd.n427 240.244
R7007 gnd.n7104 gnd.n427 240.244
R7008 gnd.n7104 gnd.n423 240.244
R7009 gnd.n7110 gnd.n423 240.244
R7010 gnd.n7110 gnd.n411 240.244
R7011 gnd.n7120 gnd.n411 240.244
R7012 gnd.n7120 gnd.n405 240.244
R7013 gnd.n7129 gnd.n405 240.244
R7014 gnd.n7129 gnd.n406 240.244
R7015 gnd.n406 gnd.n395 240.244
R7016 gnd.n395 gnd.n373 240.244
R7017 gnd.n7180 gnd.n373 240.244
R7018 gnd.n7180 gnd.n374 240.244
R7019 gnd.n7170 gnd.n374 240.244
R7020 gnd.n7170 gnd.n362 240.244
R7021 gnd.n7171 gnd.n362 240.244
R7022 gnd.n7171 gnd.n312 240.244
R7023 gnd.n7319 gnd.n312 240.244
R7024 gnd.n7319 gnd.n313 240.244
R7025 gnd.n318 gnd.n313 240.244
R7026 gnd.n319 gnd.n318 240.244
R7027 gnd.n320 gnd.n319 240.244
R7028 gnd.n329 gnd.n320 240.244
R7029 gnd.n329 gnd.n323 240.244
R7030 gnd.n7306 gnd.n323 240.244
R7031 gnd.n7306 gnd.n294 240.244
R7032 gnd.n7330 gnd.n294 240.244
R7033 gnd.n7330 gnd.n290 240.244
R7034 gnd.n7336 gnd.n290 240.244
R7035 gnd.n7336 gnd.n278 240.244
R7036 gnd.n7346 gnd.n278 240.244
R7037 gnd.n7346 gnd.n274 240.244
R7038 gnd.n7352 gnd.n274 240.244
R7039 gnd.n7352 gnd.n264 240.244
R7040 gnd.n7362 gnd.n264 240.244
R7041 gnd.n7362 gnd.n260 240.244
R7042 gnd.n7368 gnd.n260 240.244
R7043 gnd.n7368 gnd.n248 240.244
R7044 gnd.n7378 gnd.n248 240.244
R7045 gnd.n7378 gnd.n244 240.244
R7046 gnd.n7384 gnd.n244 240.244
R7047 gnd.n7384 gnd.n233 240.244
R7048 gnd.n7394 gnd.n233 240.244
R7049 gnd.n7394 gnd.n229 240.244
R7050 gnd.n7400 gnd.n229 240.244
R7051 gnd.n7400 gnd.n218 240.244
R7052 gnd.n7410 gnd.n218 240.244
R7053 gnd.n7410 gnd.n212 240.244
R7054 gnd.n7484 gnd.n212 240.244
R7055 gnd.n7484 gnd.n213 240.244
R7056 gnd.n213 gnd.n203 240.244
R7057 gnd.n7415 gnd.n203 240.244
R7058 gnd.n7415 gnd.n125 240.244
R7059 gnd.n5576 gnd.n5575 240.244
R7060 gnd.n5587 gnd.n5578 240.244
R7061 gnd.n5590 gnd.n5589 240.244
R7062 gnd.n5601 gnd.n5600 240.244
R7063 gnd.n5610 gnd.n5603 240.244
R7064 gnd.n5613 gnd.n5612 240.244
R7065 gnd.n5624 gnd.n5623 240.244
R7066 gnd.n5629 gnd.n5626 240.244
R7067 gnd.n5627 gnd.n1350 240.244
R7068 gnd.n4871 gnd.n4758 240.244
R7069 gnd.n4871 gnd.n1983 240.244
R7070 gnd.n4867 gnd.n1983 240.244
R7071 gnd.n4867 gnd.n1976 240.244
R7072 gnd.n4864 gnd.n1976 240.244
R7073 gnd.n4864 gnd.n1968 240.244
R7074 gnd.n4861 gnd.n1968 240.244
R7075 gnd.n4861 gnd.n1959 240.244
R7076 gnd.n4858 gnd.n1959 240.244
R7077 gnd.n4858 gnd.n1951 240.244
R7078 gnd.n4855 gnd.n1951 240.244
R7079 gnd.n4855 gnd.n1944 240.244
R7080 gnd.n4852 gnd.n1944 240.244
R7081 gnd.n4852 gnd.n1936 240.244
R7082 gnd.n4849 gnd.n1936 240.244
R7083 gnd.n4849 gnd.n1927 240.244
R7084 gnd.n4846 gnd.n1927 240.244
R7085 gnd.n4846 gnd.n1918 240.244
R7086 gnd.n1918 gnd.n1907 240.244
R7087 gnd.n5161 gnd.n1907 240.244
R7088 gnd.n5161 gnd.n1903 240.244
R7089 gnd.n5172 gnd.n1903 240.244
R7090 gnd.n5172 gnd.n1883 240.244
R7091 gnd.n5168 gnd.n1883 240.244
R7092 gnd.n5168 gnd.n1872 240.244
R7093 gnd.n5200 gnd.n1872 240.244
R7094 gnd.n5200 gnd.n1868 240.244
R7095 gnd.n5216 gnd.n1868 240.244
R7096 gnd.n5216 gnd.n1774 240.244
R7097 gnd.n5212 gnd.n1774 240.244
R7098 gnd.n5212 gnd.n1785 240.244
R7099 gnd.n5208 gnd.n1785 240.244
R7100 gnd.n5208 gnd.n1790 240.244
R7101 gnd.n5234 gnd.n1790 240.244
R7102 gnd.n5234 gnd.n1797 240.244
R7103 gnd.n5240 gnd.n1797 240.244
R7104 gnd.n5240 gnd.n1760 240.244
R7105 gnd.n5428 gnd.n1760 240.244
R7106 gnd.n5428 gnd.n1751 240.244
R7107 gnd.n1811 gnd.n1751 240.244
R7108 gnd.n1811 gnd.n1744 240.244
R7109 gnd.n1812 gnd.n1744 240.244
R7110 gnd.n1812 gnd.n1735 240.244
R7111 gnd.n1815 gnd.n1735 240.244
R7112 gnd.n1815 gnd.n1726 240.244
R7113 gnd.n1816 gnd.n1726 240.244
R7114 gnd.n1816 gnd.n1717 240.244
R7115 gnd.n1819 gnd.n1717 240.244
R7116 gnd.n1819 gnd.n1710 240.244
R7117 gnd.n1820 gnd.n1710 240.244
R7118 gnd.n1820 gnd.n1701 240.244
R7119 gnd.n1823 gnd.n1701 240.244
R7120 gnd.n1823 gnd.n1692 240.244
R7121 gnd.n1824 gnd.n1692 240.244
R7122 gnd.n1824 gnd.n1683 240.244
R7123 gnd.n1827 gnd.n1683 240.244
R7124 gnd.n1827 gnd.n1676 240.244
R7125 gnd.n1828 gnd.n1676 240.244
R7126 gnd.n1828 gnd.n1667 240.244
R7127 gnd.n5385 gnd.n1667 240.244
R7128 gnd.n5385 gnd.n1657 240.244
R7129 gnd.n5387 gnd.n1657 240.244
R7130 gnd.n5387 gnd.n1352 240.244
R7131 gnd.n5772 gnd.n1352 240.244
R7132 gnd.n4784 gnd.n4782 240.244
R7133 gnd.n4790 gnd.n4776 240.244
R7134 gnd.n4794 gnd.n4792 240.244
R7135 gnd.n4800 gnd.n4772 240.244
R7136 gnd.n4804 gnd.n4802 240.244
R7137 gnd.n4810 gnd.n4768 240.244
R7138 gnd.n4814 gnd.n4812 240.244
R7139 gnd.n4820 gnd.n4764 240.244
R7140 gnd.n4823 gnd.n4822 240.244
R7141 gnd.n5071 gnd.n1984 240.244
R7142 gnd.n5077 gnd.n1984 240.244
R7143 gnd.n5077 gnd.n1973 240.244
R7144 gnd.n5087 gnd.n1973 240.244
R7145 gnd.n5087 gnd.n1969 240.244
R7146 gnd.n5093 gnd.n1969 240.244
R7147 gnd.n5093 gnd.n1956 240.244
R7148 gnd.n5103 gnd.n1956 240.244
R7149 gnd.n5103 gnd.n1952 240.244
R7150 gnd.n5109 gnd.n1952 240.244
R7151 gnd.n5109 gnd.n1941 240.244
R7152 gnd.n5119 gnd.n1941 240.244
R7153 gnd.n5119 gnd.n1937 240.244
R7154 gnd.n5125 gnd.n1937 240.244
R7155 gnd.n5125 gnd.n1924 240.244
R7156 gnd.n5135 gnd.n1924 240.244
R7157 gnd.n5135 gnd.n1919 240.244
R7158 gnd.n5149 gnd.n1919 240.244
R7159 gnd.n5149 gnd.n1920 240.244
R7160 gnd.n1920 gnd.n1910 240.244
R7161 gnd.n5144 gnd.n1910 240.244
R7162 gnd.n5144 gnd.n1885 240.244
R7163 gnd.n5189 gnd.n1885 240.244
R7164 gnd.n5189 gnd.n1886 240.244
R7165 gnd.n5185 gnd.n1886 240.244
R7166 gnd.n5185 gnd.n1874 240.244
R7167 gnd.n1894 gnd.n1874 240.244
R7168 gnd.n1894 gnd.n1776 240.244
R7169 gnd.n5460 gnd.n1776 240.244
R7170 gnd.n5460 gnd.n1777 240.244
R7171 gnd.n5456 gnd.n1777 240.244
R7172 gnd.n5456 gnd.n1783 240.244
R7173 gnd.n5446 gnd.n1783 240.244
R7174 gnd.n5446 gnd.n1791 240.244
R7175 gnd.n5442 gnd.n1791 240.244
R7176 gnd.n5442 gnd.n1757 240.244
R7177 gnd.n5470 gnd.n1757 240.244
R7178 gnd.n5470 gnd.n1753 240.244
R7179 gnd.n5476 gnd.n1753 240.244
R7180 gnd.n5476 gnd.n1741 240.244
R7181 gnd.n5486 gnd.n1741 240.244
R7182 gnd.n5486 gnd.n1737 240.244
R7183 gnd.n5492 gnd.n1737 240.244
R7184 gnd.n5492 gnd.n1723 240.244
R7185 gnd.n5502 gnd.n1723 240.244
R7186 gnd.n5502 gnd.n1719 240.244
R7187 gnd.n5508 gnd.n1719 240.244
R7188 gnd.n5508 gnd.n1707 240.244
R7189 gnd.n5518 gnd.n1707 240.244
R7190 gnd.n5518 gnd.n1703 240.244
R7191 gnd.n5524 gnd.n1703 240.244
R7192 gnd.n5524 gnd.n1689 240.244
R7193 gnd.n5534 gnd.n1689 240.244
R7194 gnd.n5534 gnd.n1685 240.244
R7195 gnd.n5540 gnd.n1685 240.244
R7196 gnd.n5540 gnd.n1673 240.244
R7197 gnd.n5550 gnd.n1673 240.244
R7198 gnd.n5550 gnd.n1669 240.244
R7199 gnd.n5556 gnd.n1669 240.244
R7200 gnd.n5556 gnd.n1654 240.244
R7201 gnd.n5568 gnd.n1654 240.244
R7202 gnd.n5568 gnd.n1650 240.244
R7203 gnd.n5693 gnd.n1650 240.244
R7204 gnd.n5693 gnd.n1357 240.244
R7205 gnd.n3140 gnd.n2190 240.244
R7206 gnd.n3134 gnd.n2190 240.244
R7207 gnd.n3134 gnd.n2194 240.244
R7208 gnd.n3130 gnd.n2194 240.244
R7209 gnd.n3130 gnd.n2196 240.244
R7210 gnd.n3126 gnd.n2196 240.244
R7211 gnd.n3126 gnd.n2201 240.244
R7212 gnd.n3122 gnd.n2201 240.244
R7213 gnd.n3122 gnd.n2203 240.244
R7214 gnd.n3118 gnd.n2203 240.244
R7215 gnd.n3118 gnd.n2209 240.244
R7216 gnd.n3114 gnd.n2209 240.244
R7217 gnd.n3114 gnd.n2211 240.244
R7218 gnd.n3110 gnd.n2211 240.244
R7219 gnd.n3110 gnd.n2217 240.244
R7220 gnd.n3106 gnd.n2217 240.244
R7221 gnd.n3106 gnd.n2219 240.244
R7222 gnd.n3102 gnd.n2219 240.244
R7223 gnd.n3102 gnd.n2225 240.244
R7224 gnd.n3098 gnd.n2225 240.244
R7225 gnd.n3098 gnd.n2227 240.244
R7226 gnd.n3094 gnd.n2227 240.244
R7227 gnd.n3094 gnd.n2233 240.244
R7228 gnd.n3090 gnd.n2233 240.244
R7229 gnd.n3090 gnd.n2235 240.244
R7230 gnd.n3086 gnd.n2235 240.244
R7231 gnd.n3086 gnd.n2241 240.244
R7232 gnd.n3082 gnd.n2241 240.244
R7233 gnd.n3082 gnd.n2243 240.244
R7234 gnd.n3078 gnd.n2243 240.244
R7235 gnd.n3078 gnd.n2249 240.244
R7236 gnd.n3074 gnd.n2249 240.244
R7237 gnd.n3074 gnd.n2251 240.244
R7238 gnd.n3070 gnd.n2251 240.244
R7239 gnd.n3070 gnd.n2257 240.244
R7240 gnd.n3066 gnd.n2257 240.244
R7241 gnd.n3066 gnd.n2259 240.244
R7242 gnd.n3062 gnd.n2259 240.244
R7243 gnd.n3062 gnd.n2265 240.244
R7244 gnd.n3058 gnd.n2265 240.244
R7245 gnd.n3058 gnd.n2267 240.244
R7246 gnd.n3054 gnd.n2267 240.244
R7247 gnd.n3054 gnd.n2273 240.244
R7248 gnd.n3050 gnd.n2273 240.244
R7249 gnd.n3050 gnd.n2275 240.244
R7250 gnd.n3046 gnd.n2275 240.244
R7251 gnd.n3046 gnd.n2281 240.244
R7252 gnd.n3042 gnd.n2281 240.244
R7253 gnd.n3042 gnd.n2283 240.244
R7254 gnd.n3038 gnd.n2283 240.244
R7255 gnd.n3038 gnd.n2289 240.244
R7256 gnd.n3034 gnd.n2289 240.244
R7257 gnd.n3034 gnd.n2291 240.244
R7258 gnd.n3030 gnd.n2291 240.244
R7259 gnd.n3030 gnd.n2297 240.244
R7260 gnd.n3026 gnd.n2297 240.244
R7261 gnd.n3026 gnd.n2299 240.244
R7262 gnd.n3022 gnd.n2299 240.244
R7263 gnd.n3022 gnd.n2305 240.244
R7264 gnd.n3018 gnd.n2305 240.244
R7265 gnd.n3018 gnd.n2307 240.244
R7266 gnd.n3014 gnd.n2307 240.244
R7267 gnd.n3014 gnd.n2313 240.244
R7268 gnd.n3010 gnd.n2313 240.244
R7269 gnd.n3010 gnd.n2315 240.244
R7270 gnd.n3006 gnd.n2315 240.244
R7271 gnd.n3006 gnd.n2321 240.244
R7272 gnd.n3002 gnd.n2321 240.244
R7273 gnd.n3002 gnd.n2323 240.244
R7274 gnd.n2998 gnd.n2323 240.244
R7275 gnd.n2998 gnd.n2329 240.244
R7276 gnd.n2994 gnd.n2329 240.244
R7277 gnd.n2994 gnd.n2331 240.244
R7278 gnd.n2990 gnd.n2331 240.244
R7279 gnd.n2990 gnd.n2337 240.244
R7280 gnd.n2986 gnd.n2337 240.244
R7281 gnd.n2986 gnd.n2339 240.244
R7282 gnd.n2982 gnd.n2339 240.244
R7283 gnd.n2982 gnd.n2345 240.244
R7284 gnd.n2978 gnd.n2345 240.244
R7285 gnd.n2978 gnd.n2347 240.244
R7286 gnd.n2974 gnd.n2347 240.244
R7287 gnd.n2974 gnd.n2353 240.244
R7288 gnd.n2970 gnd.n2353 240.244
R7289 gnd.n2970 gnd.n2355 240.244
R7290 gnd.n2966 gnd.n2355 240.244
R7291 gnd.n2966 gnd.n2361 240.244
R7292 gnd.n2962 gnd.n2361 240.244
R7293 gnd.n2962 gnd.n2363 240.244
R7294 gnd.n2958 gnd.n2363 240.244
R7295 gnd.n2958 gnd.n2369 240.244
R7296 gnd.n2954 gnd.n2369 240.244
R7297 gnd.n2954 gnd.n2371 240.244
R7298 gnd.n2950 gnd.n2371 240.244
R7299 gnd.n2950 gnd.n2377 240.244
R7300 gnd.n2946 gnd.n2377 240.244
R7301 gnd.n2946 gnd.n2379 240.244
R7302 gnd.n2942 gnd.n2379 240.244
R7303 gnd.n2942 gnd.n2385 240.244
R7304 gnd.n2938 gnd.n2385 240.244
R7305 gnd.n2938 gnd.n2387 240.244
R7306 gnd.n2934 gnd.n2387 240.244
R7307 gnd.n2934 gnd.n2393 240.244
R7308 gnd.n2930 gnd.n2393 240.244
R7309 gnd.n2930 gnd.n2395 240.244
R7310 gnd.n2926 gnd.n2395 240.244
R7311 gnd.n2926 gnd.n2401 240.244
R7312 gnd.n2922 gnd.n2401 240.244
R7313 gnd.n2922 gnd.n2403 240.244
R7314 gnd.n2918 gnd.n2403 240.244
R7315 gnd.n2918 gnd.n2409 240.244
R7316 gnd.n2914 gnd.n2409 240.244
R7317 gnd.n2914 gnd.n2411 240.244
R7318 gnd.n2910 gnd.n2411 240.244
R7319 gnd.n2910 gnd.n2417 240.244
R7320 gnd.n2906 gnd.n2417 240.244
R7321 gnd.n2906 gnd.n2419 240.244
R7322 gnd.n2902 gnd.n2419 240.244
R7323 gnd.n2902 gnd.n2425 240.244
R7324 gnd.n2898 gnd.n2425 240.244
R7325 gnd.n2898 gnd.n2427 240.244
R7326 gnd.n2894 gnd.n2427 240.244
R7327 gnd.n2894 gnd.n2433 240.244
R7328 gnd.n2890 gnd.n2433 240.244
R7329 gnd.n2890 gnd.n2435 240.244
R7330 gnd.n2886 gnd.n2435 240.244
R7331 gnd.n2886 gnd.n2441 240.244
R7332 gnd.n2882 gnd.n2441 240.244
R7333 gnd.n2882 gnd.n2443 240.244
R7334 gnd.n2878 gnd.n2443 240.244
R7335 gnd.n2878 gnd.n2449 240.244
R7336 gnd.n2874 gnd.n2449 240.244
R7337 gnd.n2874 gnd.n2451 240.244
R7338 gnd.n2870 gnd.n2451 240.244
R7339 gnd.n2870 gnd.n2457 240.244
R7340 gnd.n2866 gnd.n2457 240.244
R7341 gnd.n2866 gnd.n2459 240.244
R7342 gnd.n2862 gnd.n2459 240.244
R7343 gnd.n2862 gnd.n2465 240.244
R7344 gnd.n2858 gnd.n2465 240.244
R7345 gnd.n2858 gnd.n2467 240.244
R7346 gnd.n2854 gnd.n2467 240.244
R7347 gnd.n2854 gnd.n2473 240.244
R7348 gnd.n2850 gnd.n2473 240.244
R7349 gnd.n2850 gnd.n2475 240.244
R7350 gnd.n2846 gnd.n2475 240.244
R7351 gnd.n2846 gnd.n2481 240.244
R7352 gnd.n2842 gnd.n2481 240.244
R7353 gnd.n2842 gnd.n2483 240.244
R7354 gnd.n2838 gnd.n2483 240.244
R7355 gnd.n2838 gnd.n2489 240.244
R7356 gnd.n2834 gnd.n2489 240.244
R7357 gnd.n2834 gnd.n2491 240.244
R7358 gnd.n2830 gnd.n2491 240.244
R7359 gnd.n2826 gnd.n2496 240.244
R7360 gnd.n2826 gnd.n2498 240.244
R7361 gnd.n2820 gnd.n2498 240.244
R7362 gnd.n2820 gnd.n2504 240.244
R7363 gnd.n2816 gnd.n2504 240.244
R7364 gnd.n2816 gnd.n2506 240.244
R7365 gnd.n2812 gnd.n2506 240.244
R7366 gnd.n2812 gnd.n2511 240.244
R7367 gnd.n2808 gnd.n2511 240.244
R7368 gnd.n2808 gnd.n2513 240.244
R7369 gnd.n2804 gnd.n2513 240.244
R7370 gnd.n2804 gnd.n2519 240.244
R7371 gnd.n2800 gnd.n2519 240.244
R7372 gnd.n2800 gnd.n2521 240.244
R7373 gnd.n2796 gnd.n2521 240.244
R7374 gnd.n2796 gnd.n2527 240.244
R7375 gnd.n2792 gnd.n2527 240.244
R7376 gnd.n2792 gnd.n2529 240.244
R7377 gnd.n2788 gnd.n2529 240.244
R7378 gnd.n2788 gnd.n2535 240.244
R7379 gnd.n2784 gnd.n2535 240.244
R7380 gnd.n2784 gnd.n2537 240.244
R7381 gnd.n2780 gnd.n2537 240.244
R7382 gnd.n2780 gnd.n2543 240.244
R7383 gnd.n2776 gnd.n2543 240.244
R7384 gnd.n2776 gnd.n2545 240.244
R7385 gnd.n2772 gnd.n2545 240.244
R7386 gnd.n2772 gnd.n2551 240.244
R7387 gnd.n2768 gnd.n2551 240.244
R7388 gnd.n2768 gnd.n2553 240.244
R7389 gnd.n2764 gnd.n2553 240.244
R7390 gnd.n2764 gnd.n2559 240.244
R7391 gnd.n2760 gnd.n2559 240.244
R7392 gnd.n2760 gnd.n2561 240.244
R7393 gnd.n2756 gnd.n2561 240.244
R7394 gnd.n2756 gnd.n2567 240.244
R7395 gnd.n2752 gnd.n2567 240.244
R7396 gnd.n2752 gnd.n2569 240.244
R7397 gnd.n2748 gnd.n2569 240.244
R7398 gnd.n2748 gnd.n2575 240.244
R7399 gnd.n2744 gnd.n2575 240.244
R7400 gnd.n2744 gnd.n2577 240.244
R7401 gnd.n2740 gnd.n2577 240.244
R7402 gnd.n2740 gnd.n2583 240.244
R7403 gnd.n2736 gnd.n2583 240.244
R7404 gnd.n2736 gnd.n2585 240.244
R7405 gnd.n2732 gnd.n2585 240.244
R7406 gnd.n2732 gnd.n2591 240.244
R7407 gnd.n2728 gnd.n2591 240.244
R7408 gnd.n2728 gnd.n2593 240.244
R7409 gnd.n2724 gnd.n2593 240.244
R7410 gnd.n2724 gnd.n2599 240.244
R7411 gnd.n2720 gnd.n2599 240.244
R7412 gnd.n2720 gnd.n2601 240.244
R7413 gnd.n2716 gnd.n2601 240.244
R7414 gnd.n2716 gnd.n2607 240.244
R7415 gnd.n2712 gnd.n2607 240.244
R7416 gnd.n2712 gnd.n2609 240.244
R7417 gnd.n2708 gnd.n2609 240.244
R7418 gnd.n2708 gnd.n2615 240.244
R7419 gnd.n2704 gnd.n2615 240.244
R7420 gnd.n2704 gnd.n2617 240.244
R7421 gnd.n2700 gnd.n2617 240.244
R7422 gnd.n2700 gnd.n2623 240.244
R7423 gnd.n2696 gnd.n2623 240.244
R7424 gnd.n2696 gnd.n2625 240.244
R7425 gnd.n2692 gnd.n2625 240.244
R7426 gnd.n2692 gnd.n2631 240.244
R7427 gnd.n2688 gnd.n2631 240.244
R7428 gnd.n2688 gnd.n2633 240.244
R7429 gnd.n2684 gnd.n2633 240.244
R7430 gnd.n2684 gnd.n2639 240.244
R7431 gnd.n2680 gnd.n2639 240.244
R7432 gnd.n2680 gnd.n2641 240.244
R7433 gnd.n2676 gnd.n2641 240.244
R7434 gnd.n2676 gnd.n2647 240.244
R7435 gnd.n2672 gnd.n2647 240.244
R7436 gnd.n2672 gnd.n2649 240.244
R7437 gnd.n2668 gnd.n2649 240.244
R7438 gnd.n2668 gnd.n2655 240.244
R7439 gnd.n2664 gnd.n2655 240.244
R7440 gnd.n2664 gnd.n2658 240.244
R7441 gnd.n2658 gnd.n342 240.244
R7442 gnd.n7220 gnd.n342 240.244
R7443 gnd.n5436 gnd.n1798 240.244
R7444 gnd.n5436 gnd.n1799 240.244
R7445 gnd.n5432 gnd.n1799 240.244
R7446 gnd.n5432 gnd.n5431 240.244
R7447 gnd.n5431 gnd.n1805 240.244
R7448 gnd.n5255 gnd.n1805 240.244
R7449 gnd.n5274 gnd.n5255 240.244
R7450 gnd.n5274 gnd.n5256 240.244
R7451 gnd.n5270 gnd.n5256 240.244
R7452 gnd.n5270 gnd.n5269 240.244
R7453 gnd.n5269 gnd.n1849 240.244
R7454 gnd.n5297 gnd.n1849 240.244
R7455 gnd.n5298 gnd.n5297 240.244
R7456 gnd.n5298 gnd.n1844 240.244
R7457 gnd.n5314 gnd.n1844 240.244
R7458 gnd.n5314 gnd.n1845 240.244
R7459 gnd.n5310 gnd.n1845 240.244
R7460 gnd.n5310 gnd.n5309 240.244
R7461 gnd.n5309 gnd.n1839 240.244
R7462 gnd.n5336 gnd.n1839 240.244
R7463 gnd.n5337 gnd.n5336 240.244
R7464 gnd.n5337 gnd.n1834 240.244
R7465 gnd.n5371 gnd.n1834 240.244
R7466 gnd.n5371 gnd.n1835 240.244
R7467 gnd.n5367 gnd.n1835 240.244
R7468 gnd.n5367 gnd.n5366 240.244
R7469 gnd.n5366 gnd.n5365 240.244
R7470 gnd.n5365 gnd.n5345 240.244
R7471 gnd.n5361 gnd.n5345 240.244
R7472 gnd.n5361 gnd.n5360 240.244
R7473 gnd.n5360 gnd.n5359 240.244
R7474 gnd.n5359 gnd.n5352 240.244
R7475 gnd.n5352 gnd.n1317 240.244
R7476 gnd.n5810 gnd.n1317 240.244
R7477 gnd.n5810 gnd.n1313 240.244
R7478 gnd.n5816 gnd.n1313 240.244
R7479 gnd.n5816 gnd.n1303 240.244
R7480 gnd.n5826 gnd.n1303 240.244
R7481 gnd.n5826 gnd.n1298 240.244
R7482 gnd.n5834 gnd.n1298 240.244
R7483 gnd.n5834 gnd.n1299 240.244
R7484 gnd.n1299 gnd.n1261 240.244
R7485 gnd.n5984 gnd.n1261 240.244
R7486 gnd.n5984 gnd.n1257 240.244
R7487 gnd.n5990 gnd.n1257 240.244
R7488 gnd.n5990 gnd.n1246 240.244
R7489 gnd.n6000 gnd.n1246 240.244
R7490 gnd.n6000 gnd.n1242 240.244
R7491 gnd.n6006 gnd.n1242 240.244
R7492 gnd.n6006 gnd.n1230 240.244
R7493 gnd.n6016 gnd.n1230 240.244
R7494 gnd.n6016 gnd.n1226 240.244
R7495 gnd.n6022 gnd.n1226 240.244
R7496 gnd.n6022 gnd.n1215 240.244
R7497 gnd.n6031 gnd.n1215 240.244
R7498 gnd.n6031 gnd.n1210 240.244
R7499 gnd.n6039 gnd.n1210 240.244
R7500 gnd.n6039 gnd.n1211 240.244
R7501 gnd.n1211 gnd.n1108 240.244
R7502 gnd.n6126 gnd.n1108 240.244
R7503 gnd.n6126 gnd.n1104 240.244
R7504 gnd.n6132 gnd.n1104 240.244
R7505 gnd.n6132 gnd.n1092 240.244
R7506 gnd.n6142 gnd.n1092 240.244
R7507 gnd.n6142 gnd.n1088 240.244
R7508 gnd.n6148 gnd.n1088 240.244
R7509 gnd.n6148 gnd.n1077 240.244
R7510 gnd.n6158 gnd.n1077 240.244
R7511 gnd.n6158 gnd.n1073 240.244
R7512 gnd.n6164 gnd.n1073 240.244
R7513 gnd.n6164 gnd.n1064 240.244
R7514 gnd.n6174 gnd.n1064 240.244
R7515 gnd.n6174 gnd.n1059 240.244
R7516 gnd.n6182 gnd.n1059 240.244
R7517 gnd.n6182 gnd.n1060 240.244
R7518 gnd.n1060 gnd.n1021 240.244
R7519 gnd.n6431 gnd.n1021 240.244
R7520 gnd.n6431 gnd.n1017 240.244
R7521 gnd.n6437 gnd.n1017 240.244
R7522 gnd.n6437 gnd.n1005 240.244
R7523 gnd.n6447 gnd.n1005 240.244
R7524 gnd.n6447 gnd.n1001 240.244
R7525 gnd.n6453 gnd.n1001 240.244
R7526 gnd.n6453 gnd.n989 240.244
R7527 gnd.n6463 gnd.n989 240.244
R7528 gnd.n6463 gnd.n985 240.244
R7529 gnd.n6469 gnd.n985 240.244
R7530 gnd.n6469 gnd.n975 240.244
R7531 gnd.n6479 gnd.n975 240.244
R7532 gnd.n6479 gnd.n971 240.244
R7533 gnd.n6485 gnd.n971 240.244
R7534 gnd.n6485 gnd.n960 240.244
R7535 gnd.n6495 gnd.n960 240.244
R7536 gnd.n6495 gnd.n956 240.244
R7537 gnd.n6501 gnd.n956 240.244
R7538 gnd.n6501 gnd.n944 240.244
R7539 gnd.n6511 gnd.n944 240.244
R7540 gnd.n6511 gnd.n940 240.244
R7541 gnd.n6517 gnd.n940 240.244
R7542 gnd.n6517 gnd.n927 240.244
R7543 gnd.n6533 gnd.n927 240.244
R7544 gnd.n6533 gnd.n922 240.244
R7545 gnd.n6541 gnd.n922 240.244
R7546 gnd.n6541 gnd.n923 240.244
R7547 gnd.n923 gnd.n887 240.244
R7548 gnd.n6591 gnd.n887 240.244
R7549 gnd.n6591 gnd.n882 240.244
R7550 gnd.n6599 gnd.n882 240.244
R7551 gnd.n6599 gnd.n883 240.244
R7552 gnd.n883 gnd.n660 240.244
R7553 gnd.n6782 gnd.n660 240.244
R7554 gnd.n6782 gnd.n656 240.244
R7555 gnd.n6788 gnd.n656 240.244
R7556 gnd.n6788 gnd.n645 240.244
R7557 gnd.n6799 gnd.n645 240.244
R7558 gnd.n6799 gnd.n640 240.244
R7559 gnd.n6807 gnd.n640 240.244
R7560 gnd.n6807 gnd.n641 240.244
R7561 gnd.n641 gnd.n615 240.244
R7562 gnd.n6818 gnd.n615 240.244
R7563 gnd.n6818 gnd.n611 240.244
R7564 gnd.n6824 gnd.n611 240.244
R7565 gnd.n6825 gnd.n6824 240.244
R7566 gnd.n6826 gnd.n6825 240.244
R7567 gnd.n6826 gnd.n607 240.244
R7568 gnd.n6832 gnd.n607 240.244
R7569 gnd.n6833 gnd.n6832 240.244
R7570 gnd.n6834 gnd.n6833 240.244
R7571 gnd.n6834 gnd.n603 240.244
R7572 gnd.n6840 gnd.n603 240.244
R7573 gnd.n6867 gnd.n6840 240.244
R7574 gnd.n6868 gnd.n6867 240.244
R7575 gnd.n6868 gnd.n598 240.244
R7576 gnd.n6884 gnd.n598 240.244
R7577 gnd.n6884 gnd.n599 240.244
R7578 gnd.n6880 gnd.n599 240.244
R7579 gnd.n6880 gnd.n6879 240.244
R7580 gnd.n6879 gnd.n593 240.244
R7581 gnd.n6906 gnd.n593 240.244
R7582 gnd.n6907 gnd.n6906 240.244
R7583 gnd.n6907 gnd.n588 240.244
R7584 gnd.n6915 gnd.n588 240.244
R7585 gnd.n6915 gnd.n589 240.244
R7586 gnd.n589 gnd.n393 240.244
R7587 gnd.n7140 gnd.n393 240.244
R7588 gnd.n7140 gnd.n388 240.244
R7589 gnd.n7157 gnd.n388 240.244
R7590 gnd.n7157 gnd.n389 240.244
R7591 gnd.n7153 gnd.n389 240.244
R7592 gnd.n7153 gnd.n7152 240.244
R7593 gnd.n7152 gnd.n348 240.244
R7594 gnd.n7213 gnd.n348 240.244
R7595 gnd.n7214 gnd.n7213 240.244
R7596 gnd.n7214 gnd.n343 240.244
R7597 gnd.n3144 gnd.n2188 240.244
R7598 gnd.n3144 gnd.n2184 240.244
R7599 gnd.n3150 gnd.n2184 240.244
R7600 gnd.n3150 gnd.n2182 240.244
R7601 gnd.n3154 gnd.n2182 240.244
R7602 gnd.n3154 gnd.n2178 240.244
R7603 gnd.n3160 gnd.n2178 240.244
R7604 gnd.n3160 gnd.n2176 240.244
R7605 gnd.n3164 gnd.n2176 240.244
R7606 gnd.n3164 gnd.n2172 240.244
R7607 gnd.n3170 gnd.n2172 240.244
R7608 gnd.n3170 gnd.n2170 240.244
R7609 gnd.n3174 gnd.n2170 240.244
R7610 gnd.n3174 gnd.n2166 240.244
R7611 gnd.n3180 gnd.n2166 240.244
R7612 gnd.n3180 gnd.n2164 240.244
R7613 gnd.n3184 gnd.n2164 240.244
R7614 gnd.n3184 gnd.n2160 240.244
R7615 gnd.n3190 gnd.n2160 240.244
R7616 gnd.n3190 gnd.n2158 240.244
R7617 gnd.n3194 gnd.n2158 240.244
R7618 gnd.n3194 gnd.n2154 240.244
R7619 gnd.n3200 gnd.n2154 240.244
R7620 gnd.n3200 gnd.n2152 240.244
R7621 gnd.n3204 gnd.n2152 240.244
R7622 gnd.n3204 gnd.n2148 240.244
R7623 gnd.n3210 gnd.n2148 240.244
R7624 gnd.n3210 gnd.n2146 240.244
R7625 gnd.n3214 gnd.n2146 240.244
R7626 gnd.n3214 gnd.n2142 240.244
R7627 gnd.n3220 gnd.n2142 240.244
R7628 gnd.n3220 gnd.n2140 240.244
R7629 gnd.n3224 gnd.n2140 240.244
R7630 gnd.n3224 gnd.n2136 240.244
R7631 gnd.n3230 gnd.n2136 240.244
R7632 gnd.n3230 gnd.n2134 240.244
R7633 gnd.n3234 gnd.n2134 240.244
R7634 gnd.n3234 gnd.n2130 240.244
R7635 gnd.n3240 gnd.n2130 240.244
R7636 gnd.n3240 gnd.n2128 240.244
R7637 gnd.n3244 gnd.n2128 240.244
R7638 gnd.n3244 gnd.n2124 240.244
R7639 gnd.n3250 gnd.n2124 240.244
R7640 gnd.n3250 gnd.n2122 240.244
R7641 gnd.n3254 gnd.n2122 240.244
R7642 gnd.n3254 gnd.n2118 240.244
R7643 gnd.n3260 gnd.n2118 240.244
R7644 gnd.n3260 gnd.n2116 240.244
R7645 gnd.n3264 gnd.n2116 240.244
R7646 gnd.n3264 gnd.n2112 240.244
R7647 gnd.n3270 gnd.n2112 240.244
R7648 gnd.n3270 gnd.n2110 240.244
R7649 gnd.n3274 gnd.n2110 240.244
R7650 gnd.n3274 gnd.n2106 240.244
R7651 gnd.n3280 gnd.n2106 240.244
R7652 gnd.n3280 gnd.n2104 240.244
R7653 gnd.n3284 gnd.n2104 240.244
R7654 gnd.n3284 gnd.n2100 240.244
R7655 gnd.n3290 gnd.n2100 240.244
R7656 gnd.n3290 gnd.n2098 240.244
R7657 gnd.n3294 gnd.n2098 240.244
R7658 gnd.n3294 gnd.n2094 240.244
R7659 gnd.n3300 gnd.n2094 240.244
R7660 gnd.n3300 gnd.n2092 240.244
R7661 gnd.n3304 gnd.n2092 240.244
R7662 gnd.n3304 gnd.n2088 240.244
R7663 gnd.n3310 gnd.n2088 240.244
R7664 gnd.n3310 gnd.n2086 240.244
R7665 gnd.n3314 gnd.n2086 240.244
R7666 gnd.n3314 gnd.n2082 240.244
R7667 gnd.n3320 gnd.n2082 240.244
R7668 gnd.n3320 gnd.n2080 240.244
R7669 gnd.n3324 gnd.n2080 240.244
R7670 gnd.n3324 gnd.n2076 240.244
R7671 gnd.n3330 gnd.n2076 240.244
R7672 gnd.n3330 gnd.n2074 240.244
R7673 gnd.n3334 gnd.n2074 240.244
R7674 gnd.n3334 gnd.n2070 240.244
R7675 gnd.n3340 gnd.n2070 240.244
R7676 gnd.n3340 gnd.n2068 240.244
R7677 gnd.n3344 gnd.n2068 240.244
R7678 gnd.n3344 gnd.n2063 240.244
R7679 gnd.n3353 gnd.n2063 240.244
R7680 gnd.n3353 gnd.n2064 240.244
R7681 gnd.n5676 gnd.n1311 240.244
R7682 gnd.n5676 gnd.n1304 240.244
R7683 gnd.n5678 gnd.n1304 240.244
R7684 gnd.n5678 gnd.n1296 240.244
R7685 gnd.n1296 gnd.n1286 240.244
R7686 gnd.n5845 gnd.n1286 240.244
R7687 gnd.n5845 gnd.n1263 240.244
R7688 gnd.n1283 gnd.n1263 240.244
R7689 gnd.n1283 gnd.n1255 240.244
R7690 gnd.n5854 gnd.n1255 240.244
R7691 gnd.n5854 gnd.n1247 240.244
R7692 gnd.n5966 gnd.n1247 240.244
R7693 gnd.n5966 gnd.n1240 240.244
R7694 gnd.n5859 gnd.n1240 240.244
R7695 gnd.n5859 gnd.n1232 240.244
R7696 gnd.n5860 gnd.n1232 240.244
R7697 gnd.n5860 gnd.n1224 240.244
R7698 gnd.n5863 gnd.n1224 240.244
R7699 gnd.n5863 gnd.n1217 240.244
R7700 gnd.n5949 gnd.n1217 240.244
R7701 gnd.n5949 gnd.n1208 240.244
R7702 gnd.n1208 gnd.n1198 240.244
R7703 gnd.n6050 gnd.n1198 240.244
R7704 gnd.n6050 gnd.n1110 240.244
R7705 gnd.n1195 gnd.n1110 240.244
R7706 gnd.n1195 gnd.n1102 240.244
R7707 gnd.n6057 gnd.n1102 240.244
R7708 gnd.n6057 gnd.n1094 240.244
R7709 gnd.n1126 gnd.n1094 240.244
R7710 gnd.n1126 gnd.n1086 240.244
R7711 gnd.n6064 gnd.n1086 240.244
R7712 gnd.n6064 gnd.n1079 240.244
R7713 gnd.n1142 gnd.n1079 240.244
R7714 gnd.n1142 gnd.n1072 240.244
R7715 gnd.n6071 gnd.n1072 240.244
R7716 gnd.n6071 gnd.n1066 240.244
R7717 gnd.n6078 gnd.n1066 240.244
R7718 gnd.n6078 gnd.n1057 240.244
R7719 gnd.n1057 gnd.n1048 240.244
R7720 gnd.n6193 gnd.n1048 240.244
R7721 gnd.n6193 gnd.n1024 240.244
R7722 gnd.n1045 gnd.n1024 240.244
R7723 gnd.n1045 gnd.n1015 240.244
R7724 gnd.n6200 gnd.n1015 240.244
R7725 gnd.n6200 gnd.n1007 240.244
R7726 gnd.n6413 gnd.n1007 240.244
R7727 gnd.n6413 gnd.n999 240.244
R7728 gnd.n6205 gnd.n999 240.244
R7729 gnd.n6205 gnd.n991 240.244
R7730 gnd.n6206 gnd.n991 240.244
R7731 gnd.n6206 gnd.n983 240.244
R7732 gnd.n6209 gnd.n983 240.244
R7733 gnd.n6209 gnd.n977 240.244
R7734 gnd.n6210 gnd.n977 240.244
R7735 gnd.n6210 gnd.n969 240.244
R7736 gnd.n6213 gnd.n969 240.244
R7737 gnd.n6213 gnd.n962 240.244
R7738 gnd.n6214 gnd.n962 240.244
R7739 gnd.n6214 gnd.n954 240.244
R7740 gnd.n6217 gnd.n954 240.244
R7741 gnd.n6217 gnd.n946 240.244
R7742 gnd.n6218 gnd.n946 240.244
R7743 gnd.n6218 gnd.n938 240.244
R7744 gnd.n6382 gnd.n938 240.244
R7745 gnd.n6382 gnd.n929 240.244
R7746 gnd.n929 gnd.n918 240.244
R7747 gnd.n6543 gnd.n918 240.244
R7748 gnd.n6543 gnd.n913 240.244
R7749 gnd.n6550 gnd.n913 240.244
R7750 gnd.n6550 gnd.n889 240.244
R7751 gnd.n889 gnd.n877 240.244
R7752 gnd.n6601 gnd.n877 240.244
R7753 gnd.n6601 gnd.n878 240.244
R7754 gnd.n878 gnd.n874 240.244
R7755 gnd.n874 gnd.n662 240.244
R7756 gnd.n6608 gnd.n662 240.244
R7757 gnd.n6608 gnd.n654 240.244
R7758 gnd.n6767 gnd.n654 240.244
R7759 gnd.n6767 gnd.n647 240.244
R7760 gnd.n6614 gnd.n647 240.244
R7761 gnd.n6614 gnd.n638 240.244
R7762 gnd.n6759 gnd.n638 240.244
R7763 gnd.n5584 gnd.n5583 240.244
R7764 gnd.n5594 gnd.n5593 240.244
R7765 gnd.n5596 gnd.n5595 240.244
R7766 gnd.n5607 gnd.n5606 240.244
R7767 gnd.n5617 gnd.n5616 240.244
R7768 gnd.n5619 gnd.n5618 240.244
R7769 gnd.n5633 gnd.n5632 240.244
R7770 gnd.n1345 gnd.n1344 240.244
R7771 gnd.n5780 gnd.n5779 240.244
R7772 gnd.n5788 gnd.n5787 240.244
R7773 gnd.n5791 gnd.n5790 240.244
R7774 gnd.n5798 gnd.n5797 240.244
R7775 gnd.n5801 gnd.n1332 240.244
R7776 gnd.n5807 gnd.n1309 240.244
R7777 gnd.n5818 gnd.n1306 240.244
R7778 gnd.n5824 gnd.n1306 240.244
R7779 gnd.n5824 gnd.n1294 240.244
R7780 gnd.n5836 gnd.n1294 240.244
R7781 gnd.n5836 gnd.n1289 240.244
R7782 gnd.n5843 gnd.n1289 240.244
R7783 gnd.n5843 gnd.n1265 240.244
R7784 gnd.n1265 gnd.n1253 240.244
R7785 gnd.n5992 gnd.n1253 240.244
R7786 gnd.n5992 gnd.n1249 240.244
R7787 gnd.n5998 gnd.n1249 240.244
R7788 gnd.n5998 gnd.n1238 240.244
R7789 gnd.n6008 gnd.n1238 240.244
R7790 gnd.n6008 gnd.n1234 240.244
R7791 gnd.n6014 gnd.n1234 240.244
R7792 gnd.n6014 gnd.n1223 240.244
R7793 gnd.n6024 gnd.n1223 240.244
R7794 gnd.n6024 gnd.n1219 240.244
R7795 gnd.n6030 gnd.n1219 240.244
R7796 gnd.n6030 gnd.n1206 240.244
R7797 gnd.n6041 gnd.n1206 240.244
R7798 gnd.n6041 gnd.n1201 240.244
R7799 gnd.n6048 gnd.n1201 240.244
R7800 gnd.n6048 gnd.n1112 240.244
R7801 gnd.n1112 gnd.n1100 240.244
R7802 gnd.n6134 gnd.n1100 240.244
R7803 gnd.n6134 gnd.n1096 240.244
R7804 gnd.n6140 gnd.n1096 240.244
R7805 gnd.n6140 gnd.n1085 240.244
R7806 gnd.n6150 gnd.n1085 240.244
R7807 gnd.n6150 gnd.n1081 240.244
R7808 gnd.n6156 gnd.n1081 240.244
R7809 gnd.n6156 gnd.n1071 240.244
R7810 gnd.n6166 gnd.n1071 240.244
R7811 gnd.n6166 gnd.n1067 240.244
R7812 gnd.n6172 gnd.n1067 240.244
R7813 gnd.n6172 gnd.n1055 240.244
R7814 gnd.n6184 gnd.n1055 240.244
R7815 gnd.n6184 gnd.n1050 240.244
R7816 gnd.n6191 gnd.n1050 240.244
R7817 gnd.n6191 gnd.n1026 240.244
R7818 gnd.n1026 gnd.n1013 240.244
R7819 gnd.n6439 gnd.n1013 240.244
R7820 gnd.n6439 gnd.n1009 240.244
R7821 gnd.n6445 gnd.n1009 240.244
R7822 gnd.n6445 gnd.n997 240.244
R7823 gnd.n6455 gnd.n997 240.244
R7824 gnd.n6455 gnd.n993 240.244
R7825 gnd.n6461 gnd.n993 240.244
R7826 gnd.n6461 gnd.n982 240.244
R7827 gnd.n6471 gnd.n982 240.244
R7828 gnd.n6471 gnd.n978 240.244
R7829 gnd.n6477 gnd.n978 240.244
R7830 gnd.n6477 gnd.n967 240.244
R7831 gnd.n6487 gnd.n967 240.244
R7832 gnd.n6487 gnd.n963 240.244
R7833 gnd.n6493 gnd.n963 240.244
R7834 gnd.n6493 gnd.n952 240.244
R7835 gnd.n6503 gnd.n952 240.244
R7836 gnd.n6503 gnd.n948 240.244
R7837 gnd.n6509 gnd.n948 240.244
R7838 gnd.n6509 gnd.n936 240.244
R7839 gnd.n6518 gnd.n936 240.244
R7840 gnd.n6518 gnd.n930 240.244
R7841 gnd.n6531 gnd.n930 240.244
R7842 gnd.n6531 gnd.n931 240.244
R7843 gnd.n931 gnd.n921 240.244
R7844 gnd.n6524 gnd.n921 240.244
R7845 gnd.n6524 gnd.n891 240.244
R7846 gnd.n6589 gnd.n891 240.244
R7847 gnd.n6589 gnd.n892 240.244
R7848 gnd.n892 gnd.n881 240.244
R7849 gnd.n897 gnd.n881 240.244
R7850 gnd.n6578 gnd.n897 240.244
R7851 gnd.n6578 gnd.n663 240.244
R7852 gnd.n663 gnd.n653 240.244
R7853 gnd.n6790 gnd.n653 240.244
R7854 gnd.n6790 gnd.n649 240.244
R7855 gnd.n6797 gnd.n649 240.244
R7856 gnd.n6797 gnd.n637 240.244
R7857 gnd.n6809 gnd.n637 240.244
R7858 gnd.n6809 gnd.n632 240.244
R7859 gnd.n6631 gnd.n6630 240.244
R7860 gnd.n6633 gnd.n6632 240.244
R7861 gnd.n6641 gnd.n6640 240.244
R7862 gnd.n6651 gnd.n6650 240.244
R7863 gnd.n6653 gnd.n6652 240.244
R7864 gnd.n6661 gnd.n6660 240.244
R7865 gnd.n6671 gnd.n6670 240.244
R7866 gnd.n6673 gnd.n6672 240.244
R7867 gnd.n6678 gnd.n6677 240.244
R7868 gnd.n6680 gnd.n6679 240.244
R7869 gnd.n6684 gnd.n6683 240.244
R7870 gnd.n6686 gnd.n6685 240.244
R7871 gnd.n6693 gnd.n6692 240.244
R7872 gnd.n6815 gnd.n631 240.244
R7873 gnd.n1420 gnd.n1419 240.132
R7874 gnd.n720 gnd.n719 240.132
R7875 gnd.n3141 gnd.n2189 225.874
R7876 gnd.n3133 gnd.n2189 225.874
R7877 gnd.n3133 gnd.n3132 225.874
R7878 gnd.n3132 gnd.n3131 225.874
R7879 gnd.n3131 gnd.n2195 225.874
R7880 gnd.n3125 gnd.n2195 225.874
R7881 gnd.n3125 gnd.n3124 225.874
R7882 gnd.n3124 gnd.n3123 225.874
R7883 gnd.n3123 gnd.n2202 225.874
R7884 gnd.n3117 gnd.n2202 225.874
R7885 gnd.n3117 gnd.n3116 225.874
R7886 gnd.n3116 gnd.n3115 225.874
R7887 gnd.n3115 gnd.n2210 225.874
R7888 gnd.n3109 gnd.n2210 225.874
R7889 gnd.n3109 gnd.n3108 225.874
R7890 gnd.n3108 gnd.n3107 225.874
R7891 gnd.n3107 gnd.n2218 225.874
R7892 gnd.n3101 gnd.n2218 225.874
R7893 gnd.n3101 gnd.n3100 225.874
R7894 gnd.n3100 gnd.n3099 225.874
R7895 gnd.n3099 gnd.n2226 225.874
R7896 gnd.n3093 gnd.n2226 225.874
R7897 gnd.n3093 gnd.n3092 225.874
R7898 gnd.n3092 gnd.n3091 225.874
R7899 gnd.n3091 gnd.n2234 225.874
R7900 gnd.n3085 gnd.n2234 225.874
R7901 gnd.n3085 gnd.n3084 225.874
R7902 gnd.n3084 gnd.n3083 225.874
R7903 gnd.n3083 gnd.n2242 225.874
R7904 gnd.n3077 gnd.n2242 225.874
R7905 gnd.n3077 gnd.n3076 225.874
R7906 gnd.n3076 gnd.n3075 225.874
R7907 gnd.n3075 gnd.n2250 225.874
R7908 gnd.n3069 gnd.n2250 225.874
R7909 gnd.n3069 gnd.n3068 225.874
R7910 gnd.n3068 gnd.n3067 225.874
R7911 gnd.n3067 gnd.n2258 225.874
R7912 gnd.n3061 gnd.n2258 225.874
R7913 gnd.n3061 gnd.n3060 225.874
R7914 gnd.n3060 gnd.n3059 225.874
R7915 gnd.n3059 gnd.n2266 225.874
R7916 gnd.n3053 gnd.n2266 225.874
R7917 gnd.n3053 gnd.n3052 225.874
R7918 gnd.n3052 gnd.n3051 225.874
R7919 gnd.n3051 gnd.n2274 225.874
R7920 gnd.n3045 gnd.n2274 225.874
R7921 gnd.n3045 gnd.n3044 225.874
R7922 gnd.n3044 gnd.n3043 225.874
R7923 gnd.n3043 gnd.n2282 225.874
R7924 gnd.n3037 gnd.n2282 225.874
R7925 gnd.n3037 gnd.n3036 225.874
R7926 gnd.n3036 gnd.n3035 225.874
R7927 gnd.n3035 gnd.n2290 225.874
R7928 gnd.n3029 gnd.n2290 225.874
R7929 gnd.n3029 gnd.n3028 225.874
R7930 gnd.n3028 gnd.n3027 225.874
R7931 gnd.n3027 gnd.n2298 225.874
R7932 gnd.n3021 gnd.n2298 225.874
R7933 gnd.n3021 gnd.n3020 225.874
R7934 gnd.n3020 gnd.n3019 225.874
R7935 gnd.n3019 gnd.n2306 225.874
R7936 gnd.n3013 gnd.n2306 225.874
R7937 gnd.n3013 gnd.n3012 225.874
R7938 gnd.n3012 gnd.n3011 225.874
R7939 gnd.n3011 gnd.n2314 225.874
R7940 gnd.n3005 gnd.n2314 225.874
R7941 gnd.n3005 gnd.n3004 225.874
R7942 gnd.n3004 gnd.n3003 225.874
R7943 gnd.n3003 gnd.n2322 225.874
R7944 gnd.n2997 gnd.n2322 225.874
R7945 gnd.n2997 gnd.n2996 225.874
R7946 gnd.n2996 gnd.n2995 225.874
R7947 gnd.n2995 gnd.n2330 225.874
R7948 gnd.n2989 gnd.n2330 225.874
R7949 gnd.n2989 gnd.n2988 225.874
R7950 gnd.n2988 gnd.n2987 225.874
R7951 gnd.n2987 gnd.n2338 225.874
R7952 gnd.n2981 gnd.n2338 225.874
R7953 gnd.n2981 gnd.n2980 225.874
R7954 gnd.n2980 gnd.n2979 225.874
R7955 gnd.n2979 gnd.n2346 225.874
R7956 gnd.n2973 gnd.n2346 225.874
R7957 gnd.n2973 gnd.n2972 225.874
R7958 gnd.n2972 gnd.n2971 225.874
R7959 gnd.n2971 gnd.n2354 225.874
R7960 gnd.n2965 gnd.n2354 225.874
R7961 gnd.n2965 gnd.n2964 225.874
R7962 gnd.n2964 gnd.n2963 225.874
R7963 gnd.n2963 gnd.n2362 225.874
R7964 gnd.n2957 gnd.n2362 225.874
R7965 gnd.n2957 gnd.n2956 225.874
R7966 gnd.n2956 gnd.n2955 225.874
R7967 gnd.n2955 gnd.n2370 225.874
R7968 gnd.n2949 gnd.n2370 225.874
R7969 gnd.n2949 gnd.n2948 225.874
R7970 gnd.n2948 gnd.n2947 225.874
R7971 gnd.n2947 gnd.n2378 225.874
R7972 gnd.n2941 gnd.n2378 225.874
R7973 gnd.n2941 gnd.n2940 225.874
R7974 gnd.n2940 gnd.n2939 225.874
R7975 gnd.n2939 gnd.n2386 225.874
R7976 gnd.n2933 gnd.n2386 225.874
R7977 gnd.n2933 gnd.n2932 225.874
R7978 gnd.n2932 gnd.n2931 225.874
R7979 gnd.n2931 gnd.n2394 225.874
R7980 gnd.n2925 gnd.n2394 225.874
R7981 gnd.n2925 gnd.n2924 225.874
R7982 gnd.n2924 gnd.n2923 225.874
R7983 gnd.n2923 gnd.n2402 225.874
R7984 gnd.n2917 gnd.n2402 225.874
R7985 gnd.n2917 gnd.n2916 225.874
R7986 gnd.n2916 gnd.n2915 225.874
R7987 gnd.n2915 gnd.n2410 225.874
R7988 gnd.n2909 gnd.n2410 225.874
R7989 gnd.n2909 gnd.n2908 225.874
R7990 gnd.n2908 gnd.n2907 225.874
R7991 gnd.n2907 gnd.n2418 225.874
R7992 gnd.n2901 gnd.n2418 225.874
R7993 gnd.n2901 gnd.n2900 225.874
R7994 gnd.n2900 gnd.n2899 225.874
R7995 gnd.n2899 gnd.n2426 225.874
R7996 gnd.n2893 gnd.n2426 225.874
R7997 gnd.n2893 gnd.n2892 225.874
R7998 gnd.n2892 gnd.n2891 225.874
R7999 gnd.n2891 gnd.n2434 225.874
R8000 gnd.n2885 gnd.n2434 225.874
R8001 gnd.n2885 gnd.n2884 225.874
R8002 gnd.n2884 gnd.n2883 225.874
R8003 gnd.n2883 gnd.n2442 225.874
R8004 gnd.n2877 gnd.n2442 225.874
R8005 gnd.n2877 gnd.n2876 225.874
R8006 gnd.n2876 gnd.n2875 225.874
R8007 gnd.n2875 gnd.n2450 225.874
R8008 gnd.n2869 gnd.n2450 225.874
R8009 gnd.n2869 gnd.n2868 225.874
R8010 gnd.n2868 gnd.n2867 225.874
R8011 gnd.n2867 gnd.n2458 225.874
R8012 gnd.n2861 gnd.n2458 225.874
R8013 gnd.n2861 gnd.n2860 225.874
R8014 gnd.n2860 gnd.n2859 225.874
R8015 gnd.n2859 gnd.n2466 225.874
R8016 gnd.n2853 gnd.n2466 225.874
R8017 gnd.n2853 gnd.n2852 225.874
R8018 gnd.n2852 gnd.n2851 225.874
R8019 gnd.n2851 gnd.n2474 225.874
R8020 gnd.n2845 gnd.n2474 225.874
R8021 gnd.n2845 gnd.n2844 225.874
R8022 gnd.n2844 gnd.n2843 225.874
R8023 gnd.n2843 gnd.n2482 225.874
R8024 gnd.n2837 gnd.n2482 225.874
R8025 gnd.n2837 gnd.n2836 225.874
R8026 gnd.n2836 gnd.n2835 225.874
R8027 gnd.n2835 gnd.n2490 225.874
R8028 gnd.n2829 gnd.n2490 225.874
R8029 gnd.n3912 gnd.t106 224.174
R8030 gnd.n2053 gnd.t57 224.174
R8031 gnd.n535 gnd.n496 199.319
R8032 gnd.n535 gnd.n497 199.319
R8033 gnd.n5739 gnd.n5738 199.319
R8034 gnd.n5738 gnd.n5737 199.319
R8035 gnd.n1421 gnd.n1418 186.49
R8036 gnd.n721 gnd.n718 186.49
R8037 gnd.n4626 gnd.n4625 185
R8038 gnd.n4624 gnd.n4623 185
R8039 gnd.n4603 gnd.n4602 185
R8040 gnd.n4618 gnd.n4617 185
R8041 gnd.n4616 gnd.n4615 185
R8042 gnd.n4607 gnd.n4606 185
R8043 gnd.n4610 gnd.n4609 185
R8044 gnd.n4594 gnd.n4593 185
R8045 gnd.n4592 gnd.n4591 185
R8046 gnd.n4571 gnd.n4570 185
R8047 gnd.n4586 gnd.n4585 185
R8048 gnd.n4584 gnd.n4583 185
R8049 gnd.n4575 gnd.n4574 185
R8050 gnd.n4578 gnd.n4577 185
R8051 gnd.n4562 gnd.n4561 185
R8052 gnd.n4560 gnd.n4559 185
R8053 gnd.n4539 gnd.n4538 185
R8054 gnd.n4554 gnd.n4553 185
R8055 gnd.n4552 gnd.n4551 185
R8056 gnd.n4543 gnd.n4542 185
R8057 gnd.n4546 gnd.n4545 185
R8058 gnd.n4531 gnd.n4530 185
R8059 gnd.n4529 gnd.n4528 185
R8060 gnd.n4508 gnd.n4507 185
R8061 gnd.n4523 gnd.n4522 185
R8062 gnd.n4521 gnd.n4520 185
R8063 gnd.n4512 gnd.n4511 185
R8064 gnd.n4515 gnd.n4514 185
R8065 gnd.n4499 gnd.n4498 185
R8066 gnd.n4497 gnd.n4496 185
R8067 gnd.n4476 gnd.n4475 185
R8068 gnd.n4491 gnd.n4490 185
R8069 gnd.n4489 gnd.n4488 185
R8070 gnd.n4480 gnd.n4479 185
R8071 gnd.n4483 gnd.n4482 185
R8072 gnd.n4467 gnd.n4466 185
R8073 gnd.n4465 gnd.n4464 185
R8074 gnd.n4444 gnd.n4443 185
R8075 gnd.n4459 gnd.n4458 185
R8076 gnd.n4457 gnd.n4456 185
R8077 gnd.n4448 gnd.n4447 185
R8078 gnd.n4451 gnd.n4450 185
R8079 gnd.n4435 gnd.n4434 185
R8080 gnd.n4433 gnd.n4432 185
R8081 gnd.n4412 gnd.n4411 185
R8082 gnd.n4427 gnd.n4426 185
R8083 gnd.n4425 gnd.n4424 185
R8084 gnd.n4416 gnd.n4415 185
R8085 gnd.n4419 gnd.n4418 185
R8086 gnd.n4404 gnd.n4403 185
R8087 gnd.n4402 gnd.n4401 185
R8088 gnd.n4381 gnd.n4380 185
R8089 gnd.n4396 gnd.n4395 185
R8090 gnd.n4394 gnd.n4393 185
R8091 gnd.n4385 gnd.n4384 185
R8092 gnd.n4388 gnd.n4387 185
R8093 gnd.n3913 gnd.t105 178.987
R8094 gnd.n2054 gnd.t58 178.987
R8095 gnd.n1 gnd.t351 170.774
R8096 gnd.n7 gnd.t353 170.103
R8097 gnd.n6 gnd.t151 170.103
R8098 gnd.n5 gnd.t345 170.103
R8099 gnd.n4 gnd.t164 170.103
R8100 gnd.n3 gnd.t343 170.103
R8101 gnd.n2 gnd.t177 170.103
R8102 gnd.n1 gnd.t167 170.103
R8103 gnd.n734 gnd.n732 163.367
R8104 gnd.n738 gnd.n707 163.367
R8105 gnd.n742 gnd.n740 163.367
R8106 gnd.n746 gnd.n705 163.367
R8107 gnd.n750 gnd.n748 163.367
R8108 gnd.n754 gnd.n703 163.367
R8109 gnd.n758 gnd.n756 163.367
R8110 gnd.n762 gnd.n701 163.367
R8111 gnd.n766 gnd.n764 163.367
R8112 gnd.n770 gnd.n699 163.367
R8113 gnd.n774 gnd.n772 163.367
R8114 gnd.n778 gnd.n697 163.367
R8115 gnd.n782 gnd.n780 163.367
R8116 gnd.n789 gnd.n695 163.367
R8117 gnd.n792 gnd.n791 163.367
R8118 gnd.n796 gnd.n795 163.367
R8119 gnd.n801 gnd.n799 163.367
R8120 gnd.n808 gnd.n692 163.367
R8121 gnd.n812 gnd.n810 163.367
R8122 gnd.n816 gnd.n690 163.367
R8123 gnd.n820 gnd.n818 163.367
R8124 gnd.n824 gnd.n688 163.367
R8125 gnd.n828 gnd.n826 163.367
R8126 gnd.n832 gnd.n686 163.367
R8127 gnd.n836 gnd.n834 163.367
R8128 gnd.n840 gnd.n684 163.367
R8129 gnd.n844 gnd.n842 163.367
R8130 gnd.n848 gnd.n682 163.367
R8131 gnd.n852 gnd.n850 163.367
R8132 gnd.n856 gnd.n680 163.367
R8133 gnd.n859 gnd.n858 163.367
R8134 gnd.n863 gnd.n862 163.367
R8135 gnd.n1537 gnd.n1536 163.367
R8136 gnd.n1536 gnd.n1531 163.367
R8137 gnd.n1532 gnd.n1531 163.367
R8138 gnd.n1532 gnd.n1266 163.367
R8139 gnd.n5982 gnd.n1266 163.367
R8140 gnd.n5982 gnd.n1267 163.367
R8141 gnd.n5978 gnd.n1267 163.367
R8142 gnd.n5978 gnd.n5977 163.367
R8143 gnd.n5977 gnd.n5976 163.367
R8144 gnd.n5976 gnd.n1270 163.367
R8145 gnd.n5894 gnd.n1270 163.367
R8146 gnd.n5894 gnd.n1277 163.367
R8147 gnd.n5897 gnd.n1277 163.367
R8148 gnd.n5897 gnd.n5892 163.367
R8149 gnd.n5912 gnd.n5892 163.367
R8150 gnd.n5913 gnd.n5912 163.367
R8151 gnd.n5914 gnd.n5913 163.367
R8152 gnd.n5914 gnd.n5890 163.367
R8153 gnd.n5919 gnd.n5890 163.367
R8154 gnd.n5919 gnd.n5881 163.367
R8155 gnd.n5928 gnd.n5881 163.367
R8156 gnd.n5929 gnd.n5928 163.367
R8157 gnd.n5930 gnd.n5929 163.367
R8158 gnd.n5930 gnd.n5864 163.367
R8159 gnd.n5933 gnd.n5864 163.367
R8160 gnd.n5933 gnd.n5878 163.367
R8161 gnd.n5938 gnd.n5878 163.367
R8162 gnd.n5938 gnd.n5879 163.367
R8163 gnd.n5879 gnd.n1113 163.367
R8164 gnd.n6124 gnd.n1113 163.367
R8165 gnd.n6124 gnd.n1114 163.367
R8166 gnd.n6120 gnd.n1114 163.367
R8167 gnd.n6120 gnd.n6119 163.367
R8168 gnd.n6119 gnd.n6118 163.367
R8169 gnd.n6118 gnd.n1117 163.367
R8170 gnd.n1129 gnd.n1117 163.367
R8171 gnd.n1129 gnd.n1125 163.367
R8172 gnd.n6107 gnd.n1125 163.367
R8173 gnd.n6107 gnd.n1127 163.367
R8174 gnd.n6103 gnd.n1127 163.367
R8175 gnd.n6103 gnd.n1133 163.367
R8176 gnd.n1144 gnd.n1133 163.367
R8177 gnd.n1144 gnd.n1141 163.367
R8178 gnd.n6092 gnd.n1141 163.367
R8179 gnd.n6092 gnd.n1143 163.367
R8180 gnd.n6088 gnd.n1143 163.367
R8181 gnd.n6088 gnd.n1148 163.367
R8182 gnd.n1157 gnd.n1148 163.367
R8183 gnd.n1185 gnd.n1157 163.367
R8184 gnd.n1185 gnd.n1158 163.367
R8185 gnd.n1181 gnd.n1158 163.367
R8186 gnd.n1181 gnd.n1180 163.367
R8187 gnd.n1180 gnd.n1162 163.367
R8188 gnd.n1162 gnd.n1027 163.367
R8189 gnd.n6429 gnd.n1027 163.367
R8190 gnd.n6429 gnd.n1028 163.367
R8191 gnd.n6425 gnd.n1028 163.367
R8192 gnd.n6425 gnd.n6424 163.367
R8193 gnd.n6424 gnd.n6423 163.367
R8194 gnd.n6423 gnd.n1031 163.367
R8195 gnd.n6277 gnd.n1031 163.367
R8196 gnd.n6277 gnd.n1039 163.367
R8197 gnd.n6280 gnd.n1039 163.367
R8198 gnd.n6280 gnd.n6274 163.367
R8199 gnd.n6287 gnd.n6274 163.367
R8200 gnd.n6287 gnd.n6275 163.367
R8201 gnd.n6283 gnd.n6275 163.367
R8202 gnd.n6283 gnd.n6265 163.367
R8203 gnd.n6299 gnd.n6265 163.367
R8204 gnd.n6299 gnd.n6262 163.367
R8205 gnd.n6305 gnd.n6262 163.367
R8206 gnd.n6305 gnd.n6263 163.367
R8207 gnd.n6263 gnd.n6255 163.367
R8208 gnd.n6317 gnd.n6255 163.367
R8209 gnd.n6318 gnd.n6317 163.367
R8210 gnd.n6318 gnd.n6252 163.367
R8211 gnd.n6324 gnd.n6252 163.367
R8212 gnd.n6324 gnd.n6253 163.367
R8213 gnd.n6253 gnd.n6246 163.367
R8214 gnd.n6336 gnd.n6246 163.367
R8215 gnd.n6337 gnd.n6336 163.367
R8216 gnd.n6337 gnd.n6243 163.367
R8217 gnd.n6343 gnd.n6243 163.367
R8218 gnd.n6343 gnd.n6244 163.367
R8219 gnd.n6244 gnd.n6235 163.367
R8220 gnd.n6353 gnd.n6235 163.367
R8221 gnd.n6354 gnd.n6353 163.367
R8222 gnd.n6355 gnd.n6354 163.367
R8223 gnd.n6355 gnd.n6221 163.367
R8224 gnd.n6358 gnd.n6221 163.367
R8225 gnd.n6358 gnd.n6232 163.367
R8226 gnd.n6371 gnd.n6232 163.367
R8227 gnd.n6371 gnd.n6233 163.367
R8228 gnd.n6367 gnd.n6233 163.367
R8229 gnd.n6367 gnd.n6366 163.367
R8230 gnd.n6366 gnd.n912 163.367
R8231 gnd.n6362 gnd.n912 163.367
R8232 gnd.n6362 gnd.n905 163.367
R8233 gnd.n6561 gnd.n905 163.367
R8234 gnd.n6562 gnd.n6561 163.367
R8235 gnd.n6562 gnd.n902 163.367
R8236 gnd.n6567 gnd.n902 163.367
R8237 gnd.n6567 gnd.n903 163.367
R8238 gnd.n903 gnd.n664 163.367
R8239 gnd.n6780 gnd.n664 163.367
R8240 gnd.n6780 gnd.n665 163.367
R8241 gnd.n6776 gnd.n665 163.367
R8242 gnd.n6776 gnd.n668 163.367
R8243 gnd.n869 gnd.n668 163.367
R8244 gnd.n869 gnd.n676 163.367
R8245 gnd.n1513 gnd.n1512 163.367
R8246 gnd.n1512 gnd.n1511 163.367
R8247 gnd.n1508 gnd.n1507 163.367
R8248 gnd.n1505 gnd.n1439 163.367
R8249 gnd.n1501 gnd.n1499 163.367
R8250 gnd.n1497 gnd.n1441 163.367
R8251 gnd.n1493 gnd.n1491 163.367
R8252 gnd.n1489 gnd.n1443 163.367
R8253 gnd.n1485 gnd.n1483 163.367
R8254 gnd.n1481 gnd.n1445 163.367
R8255 gnd.n1477 gnd.n1475 163.367
R8256 gnd.n1473 gnd.n1447 163.367
R8257 gnd.n1469 gnd.n1467 163.367
R8258 gnd.n1465 gnd.n1449 163.367
R8259 gnd.n1461 gnd.n1459 163.367
R8260 gnd.n1456 gnd.n1455 163.367
R8261 gnd.n1604 gnd.n1602 163.367
R8262 gnd.n1600 gnd.n1393 163.367
R8263 gnd.n1595 gnd.n1593 163.367
R8264 gnd.n1591 gnd.n1397 163.367
R8265 gnd.n1587 gnd.n1585 163.367
R8266 gnd.n1583 gnd.n1399 163.367
R8267 gnd.n1579 gnd.n1577 163.367
R8268 gnd.n1575 gnd.n1401 163.367
R8269 gnd.n1571 gnd.n1569 163.367
R8270 gnd.n1567 gnd.n1403 163.367
R8271 gnd.n1563 gnd.n1561 163.367
R8272 gnd.n1559 gnd.n1405 163.367
R8273 gnd.n1555 gnd.n1553 163.367
R8274 gnd.n1551 gnd.n1407 163.367
R8275 gnd.n1547 gnd.n1545 163.367
R8276 gnd.n1543 gnd.n1409 163.367
R8277 gnd.n1517 gnd.n1412 163.367
R8278 gnd.n1529 gnd.n1412 163.367
R8279 gnd.n1529 gnd.n1413 163.367
R8280 gnd.n1525 gnd.n1413 163.367
R8281 gnd.n1525 gnd.n1262 163.367
R8282 gnd.n1522 gnd.n1262 163.367
R8283 gnd.n1522 gnd.n1521 163.367
R8284 gnd.n1521 gnd.n1272 163.367
R8285 gnd.n5974 gnd.n1272 163.367
R8286 gnd.n5974 gnd.n1273 163.367
R8287 gnd.n5970 gnd.n1273 163.367
R8288 gnd.n5970 gnd.n5969 163.367
R8289 gnd.n5969 gnd.n1276 163.367
R8290 gnd.n5902 gnd.n1276 163.367
R8291 gnd.n5910 gnd.n5902 163.367
R8292 gnd.n5910 gnd.n5903 163.367
R8293 gnd.n5906 gnd.n5903 163.367
R8294 gnd.n5906 gnd.n5887 163.367
R8295 gnd.n5921 gnd.n5887 163.367
R8296 gnd.n5921 gnd.n5884 163.367
R8297 gnd.n5926 gnd.n5884 163.367
R8298 gnd.n5926 gnd.n5885 163.367
R8299 gnd.n5885 gnd.n5865 163.367
R8300 gnd.n5946 gnd.n5865 163.367
R8301 gnd.n5946 gnd.n5866 163.367
R8302 gnd.n5942 gnd.n5866 163.367
R8303 gnd.n5942 gnd.n5941 163.367
R8304 gnd.n5941 gnd.n5877 163.367
R8305 gnd.n5877 gnd.n5869 163.367
R8306 gnd.n5869 gnd.n1109 163.367
R8307 gnd.n5872 gnd.n1109 163.367
R8308 gnd.n5872 gnd.n5871 163.367
R8309 gnd.n5871 gnd.n1120 163.367
R8310 gnd.n6116 gnd.n1120 163.367
R8311 gnd.n6116 gnd.n1121 163.367
R8312 gnd.n6112 gnd.n1121 163.367
R8313 gnd.n6112 gnd.n6111 163.367
R8314 gnd.n6111 gnd.n1124 163.367
R8315 gnd.n1135 gnd.n1124 163.367
R8316 gnd.n6101 gnd.n1135 163.367
R8317 gnd.n6101 gnd.n1136 163.367
R8318 gnd.n6097 gnd.n1136 163.367
R8319 gnd.n6097 gnd.n6096 163.367
R8320 gnd.n6096 gnd.n1140 163.367
R8321 gnd.n1151 gnd.n1140 163.367
R8322 gnd.n6086 gnd.n1151 163.367
R8323 gnd.n6086 gnd.n1152 163.367
R8324 gnd.n6082 gnd.n1152 163.367
R8325 gnd.n6082 gnd.n1156 163.367
R8326 gnd.n1166 gnd.n1156 163.367
R8327 gnd.n1166 gnd.n1164 163.367
R8328 gnd.n1178 gnd.n1164 163.367
R8329 gnd.n1178 gnd.n1165 163.367
R8330 gnd.n1174 gnd.n1165 163.367
R8331 gnd.n1174 gnd.n1023 163.367
R8332 gnd.n1171 gnd.n1023 163.367
R8333 gnd.n1171 gnd.n1170 163.367
R8334 gnd.n1170 gnd.n1034 163.367
R8335 gnd.n6421 gnd.n1034 163.367
R8336 gnd.n6421 gnd.n1035 163.367
R8337 gnd.n6417 gnd.n1035 163.367
R8338 gnd.n6417 gnd.n6416 163.367
R8339 gnd.n6416 gnd.n1038 163.367
R8340 gnd.n6270 gnd.n1038 163.367
R8341 gnd.n6290 gnd.n6270 163.367
R8342 gnd.n6291 gnd.n6290 163.367
R8343 gnd.n6292 gnd.n6291 163.367
R8344 gnd.n6292 gnd.n6268 163.367
R8345 gnd.n6297 gnd.n6268 163.367
R8346 gnd.n6297 gnd.n6261 163.367
R8347 gnd.n6308 gnd.n6261 163.367
R8348 gnd.n6309 gnd.n6308 163.367
R8349 gnd.n6309 gnd.n6258 163.367
R8350 gnd.n6315 gnd.n6258 163.367
R8351 gnd.n6315 gnd.n6259 163.367
R8352 gnd.n6259 gnd.n6251 163.367
R8353 gnd.n6327 gnd.n6251 163.367
R8354 gnd.n6328 gnd.n6327 163.367
R8355 gnd.n6328 gnd.n6248 163.367
R8356 gnd.n6334 gnd.n6248 163.367
R8357 gnd.n6334 gnd.n6249 163.367
R8358 gnd.n6249 gnd.n6241 163.367
R8359 gnd.n6345 gnd.n6241 163.367
R8360 gnd.n6346 gnd.n6345 163.367
R8361 gnd.n6346 gnd.n6238 163.367
R8362 gnd.n6351 gnd.n6238 163.367
R8363 gnd.n6351 gnd.n6239 163.367
R8364 gnd.n6239 gnd.n6222 163.367
R8365 gnd.n6379 gnd.n6222 163.367
R8366 gnd.n6379 gnd.n6223 163.367
R8367 gnd.n6375 gnd.n6223 163.367
R8368 gnd.n6375 gnd.n6231 163.367
R8369 gnd.n6231 gnd.n6230 163.367
R8370 gnd.n6230 gnd.n6226 163.367
R8371 gnd.n6226 gnd.n910 163.367
R8372 gnd.n6553 gnd.n910 163.367
R8373 gnd.n6554 gnd.n6553 163.367
R8374 gnd.n6554 gnd.n907 163.367
R8375 gnd.n6559 gnd.n907 163.367
R8376 gnd.n6559 gnd.n908 163.367
R8377 gnd.n908 gnd.n901 163.367
R8378 gnd.n6570 gnd.n901 163.367
R8379 gnd.n6570 gnd.n899 163.367
R8380 gnd.n6575 gnd.n899 163.367
R8381 gnd.n6575 gnd.n661 163.367
R8382 gnd.n671 gnd.n661 163.367
R8383 gnd.n6774 gnd.n671 163.367
R8384 gnd.n6774 gnd.n672 163.367
R8385 gnd.n6770 gnd.n672 163.367
R8386 gnd.n6770 gnd.n675 163.367
R8387 gnd.n727 gnd.n726 156.462
R8388 gnd.n4566 gnd.n4534 153.042
R8389 gnd.n4630 gnd.n4629 152.079
R8390 gnd.n4598 gnd.n4597 152.079
R8391 gnd.n4566 gnd.n4565 152.079
R8392 gnd.n1426 gnd.n1425 152
R8393 gnd.n1427 gnd.n1416 152
R8394 gnd.n1429 gnd.n1428 152
R8395 gnd.n1431 gnd.n1414 152
R8396 gnd.n1433 gnd.n1432 152
R8397 gnd.n725 gnd.n709 152
R8398 gnd.n717 gnd.n710 152
R8399 gnd.n716 gnd.n715 152
R8400 gnd.n714 gnd.n711 152
R8401 gnd.n712 gnd.t117 150.546
R8402 gnd.t24 gnd.n4608 147.661
R8403 gnd.t160 gnd.n4576 147.661
R8404 gnd.t140 gnd.n4544 147.661
R8405 gnd.t341 gnd.n4513 147.661
R8406 gnd.t138 gnd.n4481 147.661
R8407 gnd.t349 gnd.n4449 147.661
R8408 gnd.t147 gnd.n4417 147.661
R8409 gnd.t158 gnd.n4386 147.661
R8410 gnd.n798 gnd.n797 143.351
R8411 gnd.n1454 gnd.n1392 143.351
R8412 gnd.n1603 gnd.n1392 143.351
R8413 gnd.n1423 gnd.t41 130.484
R8414 gnd.n1432 gnd.t114 126.766
R8415 gnd.n1430 gnd.t30 126.766
R8416 gnd.n1416 gnd.t59 126.766
R8417 gnd.n1424 gnd.t129 126.766
R8418 gnd.n713 gnd.t100 126.766
R8419 gnd.n715 gnd.t27 126.766
R8420 gnd.n724 gnd.t87 126.766
R8421 gnd.n726 gnd.t52 126.766
R8422 gnd.n4625 gnd.n4624 104.615
R8423 gnd.n4624 gnd.n4602 104.615
R8424 gnd.n4617 gnd.n4602 104.615
R8425 gnd.n4617 gnd.n4616 104.615
R8426 gnd.n4616 gnd.n4606 104.615
R8427 gnd.n4609 gnd.n4606 104.615
R8428 gnd.n4593 gnd.n4592 104.615
R8429 gnd.n4592 gnd.n4570 104.615
R8430 gnd.n4585 gnd.n4570 104.615
R8431 gnd.n4585 gnd.n4584 104.615
R8432 gnd.n4584 gnd.n4574 104.615
R8433 gnd.n4577 gnd.n4574 104.615
R8434 gnd.n4561 gnd.n4560 104.615
R8435 gnd.n4560 gnd.n4538 104.615
R8436 gnd.n4553 gnd.n4538 104.615
R8437 gnd.n4553 gnd.n4552 104.615
R8438 gnd.n4552 gnd.n4542 104.615
R8439 gnd.n4545 gnd.n4542 104.615
R8440 gnd.n4530 gnd.n4529 104.615
R8441 gnd.n4529 gnd.n4507 104.615
R8442 gnd.n4522 gnd.n4507 104.615
R8443 gnd.n4522 gnd.n4521 104.615
R8444 gnd.n4521 gnd.n4511 104.615
R8445 gnd.n4514 gnd.n4511 104.615
R8446 gnd.n4498 gnd.n4497 104.615
R8447 gnd.n4497 gnd.n4475 104.615
R8448 gnd.n4490 gnd.n4475 104.615
R8449 gnd.n4490 gnd.n4489 104.615
R8450 gnd.n4489 gnd.n4479 104.615
R8451 gnd.n4482 gnd.n4479 104.615
R8452 gnd.n4466 gnd.n4465 104.615
R8453 gnd.n4465 gnd.n4443 104.615
R8454 gnd.n4458 gnd.n4443 104.615
R8455 gnd.n4458 gnd.n4457 104.615
R8456 gnd.n4457 gnd.n4447 104.615
R8457 gnd.n4450 gnd.n4447 104.615
R8458 gnd.n4434 gnd.n4433 104.615
R8459 gnd.n4433 gnd.n4411 104.615
R8460 gnd.n4426 gnd.n4411 104.615
R8461 gnd.n4426 gnd.n4425 104.615
R8462 gnd.n4425 gnd.n4415 104.615
R8463 gnd.n4418 gnd.n4415 104.615
R8464 gnd.n4403 gnd.n4402 104.615
R8465 gnd.n4402 gnd.n4380 104.615
R8466 gnd.n4395 gnd.n4380 104.615
R8467 gnd.n4395 gnd.n4394 104.615
R8468 gnd.n4394 gnd.n4384 104.615
R8469 gnd.n4387 gnd.n4384 104.615
R8470 gnd.n3838 gnd.t36 100.632
R8471 gnd.n2027 gnd.t82 100.632
R8472 gnd.n7565 gnd.n134 99.6594
R8473 gnd.n7563 gnd.n7562 99.6594
R8474 gnd.n7558 gnd.n141 99.6594
R8475 gnd.n7556 gnd.n7555 99.6594
R8476 gnd.n7551 gnd.n148 99.6594
R8477 gnd.n7549 gnd.n7548 99.6594
R8478 gnd.n7544 gnd.n155 99.6594
R8479 gnd.n7542 gnd.n7541 99.6594
R8480 gnd.n7534 gnd.n162 99.6594
R8481 gnd.n7532 gnd.n7531 99.6594
R8482 gnd.n7527 gnd.n169 99.6594
R8483 gnd.n7525 gnd.n7524 99.6594
R8484 gnd.n7520 gnd.n176 99.6594
R8485 gnd.n7518 gnd.n7517 99.6594
R8486 gnd.n7513 gnd.n183 99.6594
R8487 gnd.n7511 gnd.n7510 99.6594
R8488 gnd.n7506 gnd.n190 99.6594
R8489 gnd.n7504 gnd.n7503 99.6594
R8490 gnd.n195 gnd.n194 99.6594
R8491 gnd.n7048 gnd.n7047 99.6594
R8492 gnd.n519 gnd.n490 99.6594
R8493 gnd.n7040 gnd.n491 99.6594
R8494 gnd.n7036 gnd.n492 99.6594
R8495 gnd.n7032 gnd.n493 99.6594
R8496 gnd.n7028 gnd.n494 99.6594
R8497 gnd.n7024 gnd.n495 99.6594
R8498 gnd.n7020 gnd.n496 99.6594
R8499 gnd.n7015 gnd.n498 99.6594
R8500 gnd.n7011 gnd.n499 99.6594
R8501 gnd.n7007 gnd.n500 99.6594
R8502 gnd.n7003 gnd.n501 99.6594
R8503 gnd.n6999 gnd.n502 99.6594
R8504 gnd.n6995 gnd.n503 99.6594
R8505 gnd.n6991 gnd.n504 99.6594
R8506 gnd.n6987 gnd.n505 99.6594
R8507 gnd.n6983 gnd.n506 99.6594
R8508 gnd.n558 gnd.n507 99.6594
R8509 gnd.n5763 gnd.n5762 99.6594
R8510 gnd.n5760 gnd.n5759 99.6594
R8511 gnd.n5755 gnd.n1373 99.6594
R8512 gnd.n5753 gnd.n5752 99.6594
R8513 gnd.n5748 gnd.n1380 99.6594
R8514 gnd.n5746 gnd.n5745 99.6594
R8515 gnd.n5741 gnd.n1387 99.6594
R8516 gnd.n5737 gnd.n5736 99.6594
R8517 gnd.n5732 gnd.n1614 99.6594
R8518 gnd.n5730 gnd.n5729 99.6594
R8519 gnd.n5725 gnd.n1621 99.6594
R8520 gnd.n5723 gnd.n5722 99.6594
R8521 gnd.n5718 gnd.n1628 99.6594
R8522 gnd.n5716 gnd.n5715 99.6594
R8523 gnd.n5711 gnd.n1635 99.6594
R8524 gnd.n5709 gnd.n5708 99.6594
R8525 gnd.n5704 gnd.n1644 99.6594
R8526 gnd.n5702 gnd.n5701 99.6594
R8527 gnd.n5062 gnd.n4873 99.6594
R8528 gnd.n5060 gnd.n4876 99.6594
R8529 gnd.n5056 gnd.n5055 99.6594
R8530 gnd.n5049 gnd.n4881 99.6594
R8531 gnd.n5048 gnd.n5047 99.6594
R8532 gnd.n5041 gnd.n4887 99.6594
R8533 gnd.n5040 gnd.n5039 99.6594
R8534 gnd.n5033 gnd.n4893 99.6594
R8535 gnd.n5032 gnd.n5031 99.6594
R8536 gnd.n5025 gnd.n4899 99.6594
R8537 gnd.n5024 gnd.n5023 99.6594
R8538 gnd.n5017 gnd.n4908 99.6594
R8539 gnd.n5016 gnd.n5015 99.6594
R8540 gnd.n5009 gnd.n4914 99.6594
R8541 gnd.n5008 gnd.n5007 99.6594
R8542 gnd.n5001 gnd.n4920 99.6594
R8543 gnd.n5000 gnd.n4999 99.6594
R8544 gnd.n4930 gnd.n4926 99.6594
R8545 gnd.n4989 gnd.n4988 99.6594
R8546 gnd.n4746 gnd.n2010 99.6594
R8547 gnd.n4744 gnd.n2009 99.6594
R8548 gnd.n4740 gnd.n2008 99.6594
R8549 gnd.n4736 gnd.n2007 99.6594
R8550 gnd.n4732 gnd.n2006 99.6594
R8551 gnd.n4728 gnd.n2005 99.6594
R8552 gnd.n4724 gnd.n2004 99.6594
R8553 gnd.n3362 gnd.n2003 99.6594
R8554 gnd.n4050 gnd.n3781 99.6594
R8555 gnd.n3807 gnd.n3788 99.6594
R8556 gnd.n3809 gnd.n3789 99.6594
R8557 gnd.n3817 gnd.n3790 99.6594
R8558 gnd.n3819 gnd.n3791 99.6594
R8559 gnd.n3827 gnd.n3792 99.6594
R8560 gnd.n3829 gnd.n3793 99.6594
R8561 gnd.n3837 gnd.n3794 99.6594
R8562 gnd.n4714 gnd.n1990 99.6594
R8563 gnd.n4710 gnd.n1991 99.6594
R8564 gnd.n4706 gnd.n1992 99.6594
R8565 gnd.n4702 gnd.n1993 99.6594
R8566 gnd.n4698 gnd.n1994 99.6594
R8567 gnd.n4694 gnd.n1995 99.6594
R8568 gnd.n4690 gnd.n1996 99.6594
R8569 gnd.n4686 gnd.n1997 99.6594
R8570 gnd.n4682 gnd.n1998 99.6594
R8571 gnd.n4678 gnd.n1999 99.6594
R8572 gnd.n4674 gnd.n2000 99.6594
R8573 gnd.n4670 gnd.n2001 99.6594
R8574 gnd.n4666 gnd.n2002 99.6594
R8575 gnd.n3965 gnd.n3964 99.6594
R8576 gnd.n3959 gnd.n3876 99.6594
R8577 gnd.n3956 gnd.n3877 99.6594
R8578 gnd.n3952 gnd.n3878 99.6594
R8579 gnd.n3948 gnd.n3879 99.6594
R8580 gnd.n3944 gnd.n3880 99.6594
R8581 gnd.n3940 gnd.n3881 99.6594
R8582 gnd.n3936 gnd.n3882 99.6594
R8583 gnd.n3932 gnd.n3883 99.6594
R8584 gnd.n3928 gnd.n3884 99.6594
R8585 gnd.n3924 gnd.n3885 99.6594
R8586 gnd.n3920 gnd.n3886 99.6594
R8587 gnd.n3967 gnd.n3875 99.6594
R8588 gnd.n7420 gnd.n7419 99.6594
R8589 gnd.n7425 gnd.n7424 99.6594
R8590 gnd.n7428 gnd.n7427 99.6594
R8591 gnd.n7433 gnd.n7432 99.6594
R8592 gnd.n7436 gnd.n7435 99.6594
R8593 gnd.n7441 gnd.n7440 99.6594
R8594 gnd.n7444 gnd.n7443 99.6594
R8595 gnd.n7449 gnd.n7447 99.6594
R8596 gnd.n7575 gnd.n121 99.6594
R8597 gnd.n6621 gnd.n508 99.6594
R8598 gnd.n6625 gnd.n509 99.6594
R8599 gnd.n6627 gnd.n510 99.6594
R8600 gnd.n6637 gnd.n511 99.6594
R8601 gnd.n6645 gnd.n512 99.6594
R8602 gnd.n6647 gnd.n513 99.6594
R8603 gnd.n6657 gnd.n514 99.6594
R8604 gnd.n6665 gnd.n515 99.6594
R8605 gnd.n6667 gnd.n516 99.6594
R8606 gnd.n5578 gnd.n5577 99.6594
R8607 gnd.n5589 gnd.n5588 99.6594
R8608 gnd.n5600 gnd.n5599 99.6594
R8609 gnd.n5603 gnd.n5602 99.6594
R8610 gnd.n5612 gnd.n5611 99.6594
R8611 gnd.n5623 gnd.n5622 99.6594
R8612 gnd.n5626 gnd.n5625 99.6594
R8613 gnd.n5628 gnd.n5627 99.6594
R8614 gnd.n5773 gnd.n1351 99.6594
R8615 gnd.n4781 gnd.n1987 99.6594
R8616 gnd.n4784 gnd.n4783 99.6594
R8617 gnd.n4791 gnd.n4790 99.6594
R8618 gnd.n4794 gnd.n4793 99.6594
R8619 gnd.n4801 gnd.n4800 99.6594
R8620 gnd.n4804 gnd.n4803 99.6594
R8621 gnd.n4811 gnd.n4810 99.6594
R8622 gnd.n4814 gnd.n4813 99.6594
R8623 gnd.n4821 gnd.n4820 99.6594
R8624 gnd.n4782 gnd.n4781 99.6594
R8625 gnd.n4783 gnd.n4776 99.6594
R8626 gnd.n4792 gnd.n4791 99.6594
R8627 gnd.n4793 gnd.n4772 99.6594
R8628 gnd.n4802 gnd.n4801 99.6594
R8629 gnd.n4803 gnd.n4768 99.6594
R8630 gnd.n4812 gnd.n4811 99.6594
R8631 gnd.n4813 gnd.n4764 99.6594
R8632 gnd.n4822 gnd.n4821 99.6594
R8633 gnd.n1351 gnd.n1350 99.6594
R8634 gnd.n5629 gnd.n5628 99.6594
R8635 gnd.n5625 gnd.n5624 99.6594
R8636 gnd.n5622 gnd.n5613 99.6594
R8637 gnd.n5611 gnd.n5610 99.6594
R8638 gnd.n5602 gnd.n5601 99.6594
R8639 gnd.n5599 gnd.n5590 99.6594
R8640 gnd.n5588 gnd.n5587 99.6594
R8641 gnd.n5577 gnd.n5576 99.6594
R8642 gnd.n6624 gnd.n508 99.6594
R8643 gnd.n6626 gnd.n509 99.6594
R8644 gnd.n6636 gnd.n510 99.6594
R8645 gnd.n6644 gnd.n511 99.6594
R8646 gnd.n6646 gnd.n512 99.6594
R8647 gnd.n6656 gnd.n513 99.6594
R8648 gnd.n6664 gnd.n514 99.6594
R8649 gnd.n6666 gnd.n515 99.6594
R8650 gnd.n6711 gnd.n516 99.6594
R8651 gnd.n7448 gnd.n121 99.6594
R8652 gnd.n7447 gnd.n7446 99.6594
R8653 gnd.n7443 gnd.n7442 99.6594
R8654 gnd.n7440 gnd.n7439 99.6594
R8655 gnd.n7435 gnd.n7434 99.6594
R8656 gnd.n7432 gnd.n7431 99.6594
R8657 gnd.n7427 gnd.n7426 99.6594
R8658 gnd.n7424 gnd.n7423 99.6594
R8659 gnd.n7419 gnd.n7418 99.6594
R8660 gnd.n3965 gnd.n3888 99.6594
R8661 gnd.n3957 gnd.n3876 99.6594
R8662 gnd.n3953 gnd.n3877 99.6594
R8663 gnd.n3949 gnd.n3878 99.6594
R8664 gnd.n3945 gnd.n3879 99.6594
R8665 gnd.n3941 gnd.n3880 99.6594
R8666 gnd.n3937 gnd.n3881 99.6594
R8667 gnd.n3933 gnd.n3882 99.6594
R8668 gnd.n3929 gnd.n3883 99.6594
R8669 gnd.n3925 gnd.n3884 99.6594
R8670 gnd.n3921 gnd.n3885 99.6594
R8671 gnd.n3917 gnd.n3886 99.6594
R8672 gnd.n3968 gnd.n3967 99.6594
R8673 gnd.n4669 gnd.n2002 99.6594
R8674 gnd.n4673 gnd.n2001 99.6594
R8675 gnd.n4677 gnd.n2000 99.6594
R8676 gnd.n4681 gnd.n1999 99.6594
R8677 gnd.n4685 gnd.n1998 99.6594
R8678 gnd.n4689 gnd.n1997 99.6594
R8679 gnd.n4693 gnd.n1996 99.6594
R8680 gnd.n4697 gnd.n1995 99.6594
R8681 gnd.n4701 gnd.n1994 99.6594
R8682 gnd.n4705 gnd.n1993 99.6594
R8683 gnd.n4709 gnd.n1992 99.6594
R8684 gnd.n4713 gnd.n1991 99.6594
R8685 gnd.n2031 gnd.n1990 99.6594
R8686 gnd.n4051 gnd.n4050 99.6594
R8687 gnd.n3810 gnd.n3788 99.6594
R8688 gnd.n3816 gnd.n3789 99.6594
R8689 gnd.n3820 gnd.n3790 99.6594
R8690 gnd.n3826 gnd.n3791 99.6594
R8691 gnd.n3830 gnd.n3792 99.6594
R8692 gnd.n3836 gnd.n3793 99.6594
R8693 gnd.n3794 gnd.n3778 99.6594
R8694 gnd.n4723 gnd.n2003 99.6594
R8695 gnd.n4727 gnd.n2004 99.6594
R8696 gnd.n4731 gnd.n2005 99.6594
R8697 gnd.n4735 gnd.n2006 99.6594
R8698 gnd.n4739 gnd.n2007 99.6594
R8699 gnd.n4743 gnd.n2008 99.6594
R8700 gnd.n4747 gnd.n2009 99.6594
R8701 gnd.n2012 gnd.n2010 99.6594
R8702 gnd.n5063 gnd.n5062 99.6594
R8703 gnd.n5057 gnd.n4876 99.6594
R8704 gnd.n5055 gnd.n5054 99.6594
R8705 gnd.n5050 gnd.n5049 99.6594
R8706 gnd.n5047 gnd.n5046 99.6594
R8707 gnd.n5042 gnd.n5041 99.6594
R8708 gnd.n5039 gnd.n5038 99.6594
R8709 gnd.n5034 gnd.n5033 99.6594
R8710 gnd.n5031 gnd.n5030 99.6594
R8711 gnd.n5026 gnd.n5025 99.6594
R8712 gnd.n5023 gnd.n5022 99.6594
R8713 gnd.n5018 gnd.n5017 99.6594
R8714 gnd.n5015 gnd.n5014 99.6594
R8715 gnd.n5010 gnd.n5009 99.6594
R8716 gnd.n5007 gnd.n5006 99.6594
R8717 gnd.n5002 gnd.n5001 99.6594
R8718 gnd.n4999 gnd.n4998 99.6594
R8719 gnd.n4931 gnd.n4930 99.6594
R8720 gnd.n4990 gnd.n4989 99.6594
R8721 gnd.n5703 gnd.n5702 99.6594
R8722 gnd.n1644 gnd.n1636 99.6594
R8723 gnd.n5710 gnd.n5709 99.6594
R8724 gnd.n1635 gnd.n1629 99.6594
R8725 gnd.n5717 gnd.n5716 99.6594
R8726 gnd.n1628 gnd.n1622 99.6594
R8727 gnd.n5724 gnd.n5723 99.6594
R8728 gnd.n1621 gnd.n1615 99.6594
R8729 gnd.n5731 gnd.n5730 99.6594
R8730 gnd.n1614 gnd.n1607 99.6594
R8731 gnd.n5740 gnd.n5739 99.6594
R8732 gnd.n1387 gnd.n1381 99.6594
R8733 gnd.n5747 gnd.n5746 99.6594
R8734 gnd.n1380 gnd.n1374 99.6594
R8735 gnd.n5754 gnd.n5753 99.6594
R8736 gnd.n1373 gnd.n1366 99.6594
R8737 gnd.n5761 gnd.n5760 99.6594
R8738 gnd.n5764 gnd.n5763 99.6594
R8739 gnd.n7047 gnd.n488 99.6594
R8740 gnd.n7041 gnd.n490 99.6594
R8741 gnd.n7037 gnd.n491 99.6594
R8742 gnd.n7033 gnd.n492 99.6594
R8743 gnd.n7029 gnd.n493 99.6594
R8744 gnd.n7025 gnd.n494 99.6594
R8745 gnd.n7021 gnd.n495 99.6594
R8746 gnd.n7016 gnd.n497 99.6594
R8747 gnd.n7012 gnd.n498 99.6594
R8748 gnd.n7008 gnd.n499 99.6594
R8749 gnd.n7004 gnd.n500 99.6594
R8750 gnd.n7000 gnd.n501 99.6594
R8751 gnd.n6996 gnd.n502 99.6594
R8752 gnd.n6992 gnd.n503 99.6594
R8753 gnd.n6988 gnd.n504 99.6594
R8754 gnd.n6984 gnd.n505 99.6594
R8755 gnd.n557 gnd.n506 99.6594
R8756 gnd.n6976 gnd.n507 99.6594
R8757 gnd.n194 gnd.n191 99.6594
R8758 gnd.n7505 gnd.n7504 99.6594
R8759 gnd.n190 gnd.n184 99.6594
R8760 gnd.n7512 gnd.n7511 99.6594
R8761 gnd.n183 gnd.n177 99.6594
R8762 gnd.n7519 gnd.n7518 99.6594
R8763 gnd.n176 gnd.n170 99.6594
R8764 gnd.n7526 gnd.n7525 99.6594
R8765 gnd.n169 gnd.n163 99.6594
R8766 gnd.n7533 gnd.n7532 99.6594
R8767 gnd.n162 gnd.n156 99.6594
R8768 gnd.n7543 gnd.n7542 99.6594
R8769 gnd.n155 gnd.n149 99.6594
R8770 gnd.n7550 gnd.n7549 99.6594
R8771 gnd.n148 gnd.n142 99.6594
R8772 gnd.n7557 gnd.n7556 99.6594
R8773 gnd.n141 gnd.n135 99.6594
R8774 gnd.n7564 gnd.n7563 99.6594
R8775 gnd.n134 gnd.n131 99.6594
R8776 gnd.n5581 gnd.n1319 99.6594
R8777 gnd.n5584 gnd.n1320 99.6594
R8778 gnd.n5594 gnd.n1321 99.6594
R8779 gnd.n5596 gnd.n1322 99.6594
R8780 gnd.n5607 gnd.n1323 99.6594
R8781 gnd.n5617 gnd.n1324 99.6594
R8782 gnd.n5619 gnd.n1325 99.6594
R8783 gnd.n5633 gnd.n1326 99.6594
R8784 gnd.n1345 gnd.n1327 99.6594
R8785 gnd.n5779 gnd.n1328 99.6594
R8786 gnd.n5788 gnd.n1329 99.6594
R8787 gnd.n5790 gnd.n1330 99.6594
R8788 gnd.n5798 gnd.n1331 99.6594
R8789 gnd.n5808 gnd.n1332 99.6594
R8790 gnd.n5583 gnd.n1319 99.6594
R8791 gnd.n5593 gnd.n1320 99.6594
R8792 gnd.n5595 gnd.n1321 99.6594
R8793 gnd.n5606 gnd.n1322 99.6594
R8794 gnd.n5616 gnd.n1323 99.6594
R8795 gnd.n5618 gnd.n1324 99.6594
R8796 gnd.n5632 gnd.n1325 99.6594
R8797 gnd.n1344 gnd.n1326 99.6594
R8798 gnd.n5780 gnd.n1327 99.6594
R8799 gnd.n5787 gnd.n1328 99.6594
R8800 gnd.n5791 gnd.n1329 99.6594
R8801 gnd.n5797 gnd.n1330 99.6594
R8802 gnd.n5801 gnd.n1331 99.6594
R8803 gnd.n5808 gnd.n5807 99.6594
R8804 gnd.n6758 gnd.n617 99.6594
R8805 gnd.n6631 gnd.n618 99.6594
R8806 gnd.n6633 gnd.n619 99.6594
R8807 gnd.n6641 gnd.n620 99.6594
R8808 gnd.n6651 gnd.n621 99.6594
R8809 gnd.n6653 gnd.n622 99.6594
R8810 gnd.n6661 gnd.n623 99.6594
R8811 gnd.n6671 gnd.n624 99.6594
R8812 gnd.n6673 gnd.n625 99.6594
R8813 gnd.n6678 gnd.n626 99.6594
R8814 gnd.n6680 gnd.n627 99.6594
R8815 gnd.n6684 gnd.n628 99.6594
R8816 gnd.n6686 gnd.n629 99.6594
R8817 gnd.n6693 gnd.n630 99.6594
R8818 gnd.n631 gnd.n630 99.6594
R8819 gnd.n6692 gnd.n629 99.6594
R8820 gnd.n6685 gnd.n628 99.6594
R8821 gnd.n6683 gnd.n627 99.6594
R8822 gnd.n6679 gnd.n626 99.6594
R8823 gnd.n6677 gnd.n625 99.6594
R8824 gnd.n6672 gnd.n624 99.6594
R8825 gnd.n6670 gnd.n623 99.6594
R8826 gnd.n6660 gnd.n622 99.6594
R8827 gnd.n6652 gnd.n621 99.6594
R8828 gnd.n6650 gnd.n620 99.6594
R8829 gnd.n6640 gnd.n619 99.6594
R8830 gnd.n6632 gnd.n618 99.6594
R8831 gnd.n6630 gnd.n617 99.6594
R8832 gnd.n1336 gnd.t113 98.63
R8833 gnd.n118 gnd.t46 98.63
R8834 gnd.n6712 gnd.t86 98.63
R8835 gnd.n1348 gnd.t98 98.63
R8836 gnd.n537 gnd.t79 98.63
R8837 gnd.n559 gnd.t51 98.63
R8838 gnd.n197 gnd.t124 98.63
R8839 gnd.n7536 gnd.t133 98.63
R8840 gnd.n4900 gnd.t72 98.63
R8841 gnd.n4932 gnd.t40 98.63
R8842 gnd.n4761 gnd.t109 98.63
R8843 gnd.n1641 gnd.t68 98.63
R8844 gnd.n1388 gnd.t95 98.63
R8845 gnd.n6689 gnd.t92 98.63
R8846 gnd.n1394 gnd.t128 96.6984
R8847 gnd.n804 gnd.t64 96.6984
R8848 gnd.n1450 gnd.t76 96.6906
R8849 gnd.n785 gnd.t121 96.6906
R8850 gnd.n2828 gnd.n2827 89.3769
R8851 gnd.n2827 gnd.n2497 89.3769
R8852 gnd.n2819 gnd.n2497 89.3769
R8853 gnd.n2819 gnd.n2818 89.3769
R8854 gnd.n2818 gnd.n2817 89.3769
R8855 gnd.n2817 gnd.n2505 89.3769
R8856 gnd.n2811 gnd.n2505 89.3769
R8857 gnd.n2811 gnd.n2810 89.3769
R8858 gnd.n2810 gnd.n2809 89.3769
R8859 gnd.n2809 gnd.n2512 89.3769
R8860 gnd.n2803 gnd.n2512 89.3769
R8861 gnd.n2803 gnd.n2802 89.3769
R8862 gnd.n2802 gnd.n2801 89.3769
R8863 gnd.n2801 gnd.n2520 89.3769
R8864 gnd.n2795 gnd.n2520 89.3769
R8865 gnd.n2795 gnd.n2794 89.3769
R8866 gnd.n2794 gnd.n2793 89.3769
R8867 gnd.n2793 gnd.n2528 89.3769
R8868 gnd.n2787 gnd.n2528 89.3769
R8869 gnd.n2787 gnd.n2786 89.3769
R8870 gnd.n2786 gnd.n2785 89.3769
R8871 gnd.n2785 gnd.n2536 89.3769
R8872 gnd.n2779 gnd.n2536 89.3769
R8873 gnd.n2779 gnd.n2778 89.3769
R8874 gnd.n2778 gnd.n2777 89.3769
R8875 gnd.n2777 gnd.n2544 89.3769
R8876 gnd.n2771 gnd.n2544 89.3769
R8877 gnd.n2771 gnd.n2770 89.3769
R8878 gnd.n2770 gnd.n2769 89.3769
R8879 gnd.n2769 gnd.n2552 89.3769
R8880 gnd.n2763 gnd.n2552 89.3769
R8881 gnd.n2763 gnd.n2762 89.3769
R8882 gnd.n2762 gnd.n2761 89.3769
R8883 gnd.n2761 gnd.n2560 89.3769
R8884 gnd.n2755 gnd.n2560 89.3769
R8885 gnd.n2755 gnd.n2754 89.3769
R8886 gnd.n2754 gnd.n2753 89.3769
R8887 gnd.n2753 gnd.n2568 89.3769
R8888 gnd.n2747 gnd.n2568 89.3769
R8889 gnd.n2747 gnd.n2746 89.3769
R8890 gnd.n2746 gnd.n2745 89.3769
R8891 gnd.n2745 gnd.n2576 89.3769
R8892 gnd.n2739 gnd.n2576 89.3769
R8893 gnd.n2739 gnd.n2738 89.3769
R8894 gnd.n2738 gnd.n2737 89.3769
R8895 gnd.n2737 gnd.n2584 89.3769
R8896 gnd.n2731 gnd.n2584 89.3769
R8897 gnd.n2731 gnd.n2730 89.3769
R8898 gnd.n2730 gnd.n2729 89.3769
R8899 gnd.n2729 gnd.n2592 89.3769
R8900 gnd.n2723 gnd.n2592 89.3769
R8901 gnd.n2723 gnd.n2722 89.3769
R8902 gnd.n2722 gnd.n2721 89.3769
R8903 gnd.n2721 gnd.n2600 89.3769
R8904 gnd.n2715 gnd.n2600 89.3769
R8905 gnd.n2715 gnd.n2714 89.3769
R8906 gnd.n2714 gnd.n2713 89.3769
R8907 gnd.n2713 gnd.n2608 89.3769
R8908 gnd.n2707 gnd.n2608 89.3769
R8909 gnd.n2707 gnd.n2706 89.3769
R8910 gnd.n2706 gnd.n2705 89.3769
R8911 gnd.n2705 gnd.n2616 89.3769
R8912 gnd.n2699 gnd.n2616 89.3769
R8913 gnd.n2699 gnd.n2698 89.3769
R8914 gnd.n2698 gnd.n2697 89.3769
R8915 gnd.n2697 gnd.n2624 89.3769
R8916 gnd.n2691 gnd.n2624 89.3769
R8917 gnd.n2691 gnd.n2690 89.3769
R8918 gnd.n2690 gnd.n2689 89.3769
R8919 gnd.n2689 gnd.n2632 89.3769
R8920 gnd.n2683 gnd.n2632 89.3769
R8921 gnd.n2683 gnd.n2682 89.3769
R8922 gnd.n2682 gnd.n2681 89.3769
R8923 gnd.n2681 gnd.n2640 89.3769
R8924 gnd.n2675 gnd.n2640 89.3769
R8925 gnd.n2675 gnd.n2674 89.3769
R8926 gnd.n2674 gnd.n2673 89.3769
R8927 gnd.n2673 gnd.n2648 89.3769
R8928 gnd.n2667 gnd.n2648 89.3769
R8929 gnd.n2667 gnd.n2666 89.3769
R8930 gnd.n2666 gnd.n2665 89.3769
R8931 gnd.n2665 gnd.n2657 89.3769
R8932 gnd.n2657 gnd.n2656 89.3769
R8933 gnd.n1423 gnd.n1422 81.8399
R8934 gnd.n3839 gnd.t35 74.8376
R8935 gnd.n2028 gnd.t83 74.8376
R8936 gnd.n1395 gnd.t127 72.8438
R8937 gnd.n805 gnd.t65 72.8438
R8938 gnd.n1424 gnd.n1417 72.8411
R8939 gnd.n1430 gnd.n1415 72.8411
R8940 gnd.n724 gnd.n723 72.8411
R8941 gnd.n1337 gnd.t112 72.836
R8942 gnd.n1451 gnd.t75 72.836
R8943 gnd.n786 gnd.t122 72.836
R8944 gnd.n119 gnd.t47 72.836
R8945 gnd.n6713 gnd.t85 72.836
R8946 gnd.n1349 gnd.t99 72.836
R8947 gnd.n538 gnd.t78 72.836
R8948 gnd.n560 gnd.t50 72.836
R8949 gnd.n198 gnd.t125 72.836
R8950 gnd.n7537 gnd.t134 72.836
R8951 gnd.n4901 gnd.t71 72.836
R8952 gnd.n4933 gnd.t39 72.836
R8953 gnd.n4762 gnd.t108 72.836
R8954 gnd.n1642 gnd.t69 72.836
R8955 gnd.n1389 gnd.t96 72.836
R8956 gnd.n6690 gnd.t93 72.836
R8957 gnd.n732 gnd.n731 71.676
R8958 gnd.n733 gnd.n707 71.676
R8959 gnd.n740 gnd.n739 71.676
R8960 gnd.n741 gnd.n705 71.676
R8961 gnd.n748 gnd.n747 71.676
R8962 gnd.n749 gnd.n703 71.676
R8963 gnd.n756 gnd.n755 71.676
R8964 gnd.n757 gnd.n701 71.676
R8965 gnd.n764 gnd.n763 71.676
R8966 gnd.n765 gnd.n699 71.676
R8967 gnd.n772 gnd.n771 71.676
R8968 gnd.n773 gnd.n697 71.676
R8969 gnd.n780 gnd.n779 71.676
R8970 gnd.n781 gnd.n695 71.676
R8971 gnd.n791 gnd.n790 71.676
R8972 gnd.n795 gnd.n693 71.676
R8973 gnd.n799 gnd.n798 71.676
R8974 gnd.n800 gnd.n692 71.676
R8975 gnd.n810 gnd.n809 71.676
R8976 gnd.n811 gnd.n690 71.676
R8977 gnd.n818 gnd.n817 71.676
R8978 gnd.n819 gnd.n688 71.676
R8979 gnd.n826 gnd.n825 71.676
R8980 gnd.n827 gnd.n686 71.676
R8981 gnd.n834 gnd.n833 71.676
R8982 gnd.n835 gnd.n684 71.676
R8983 gnd.n842 gnd.n841 71.676
R8984 gnd.n843 gnd.n682 71.676
R8985 gnd.n850 gnd.n849 71.676
R8986 gnd.n851 gnd.n680 71.676
R8987 gnd.n858 gnd.n857 71.676
R8988 gnd.n862 gnd.n678 71.676
R8989 gnd.n865 gnd.n864 71.676
R8990 gnd.n1516 gnd.n1435 71.676
R8991 gnd.n1511 gnd.n1437 71.676
R8992 gnd.n1507 gnd.n1506 71.676
R8993 gnd.n1500 gnd.n1439 71.676
R8994 gnd.n1499 gnd.n1498 71.676
R8995 gnd.n1492 gnd.n1441 71.676
R8996 gnd.n1491 gnd.n1490 71.676
R8997 gnd.n1484 gnd.n1443 71.676
R8998 gnd.n1483 gnd.n1482 71.676
R8999 gnd.n1476 gnd.n1445 71.676
R9000 gnd.n1475 gnd.n1474 71.676
R9001 gnd.n1468 gnd.n1447 71.676
R9002 gnd.n1467 gnd.n1466 71.676
R9003 gnd.n1460 gnd.n1449 71.676
R9004 gnd.n1459 gnd.n1453 71.676
R9005 gnd.n1455 gnd.n1454 71.676
R9006 gnd.n1602 gnd.n1601 71.676
R9007 gnd.n1594 gnd.n1393 71.676
R9008 gnd.n1593 gnd.n1592 71.676
R9009 gnd.n1586 gnd.n1397 71.676
R9010 gnd.n1585 gnd.n1584 71.676
R9011 gnd.n1578 gnd.n1399 71.676
R9012 gnd.n1577 gnd.n1576 71.676
R9013 gnd.n1570 gnd.n1401 71.676
R9014 gnd.n1569 gnd.n1568 71.676
R9015 gnd.n1562 gnd.n1403 71.676
R9016 gnd.n1561 gnd.n1560 71.676
R9017 gnd.n1554 gnd.n1405 71.676
R9018 gnd.n1553 gnd.n1552 71.676
R9019 gnd.n1546 gnd.n1407 71.676
R9020 gnd.n1545 gnd.n1544 71.676
R9021 gnd.n1538 gnd.n1409 71.676
R9022 gnd.n1513 gnd.n1435 71.676
R9023 gnd.n1508 gnd.n1437 71.676
R9024 gnd.n1506 gnd.n1505 71.676
R9025 gnd.n1501 gnd.n1500 71.676
R9026 gnd.n1498 gnd.n1497 71.676
R9027 gnd.n1493 gnd.n1492 71.676
R9028 gnd.n1490 gnd.n1489 71.676
R9029 gnd.n1485 gnd.n1484 71.676
R9030 gnd.n1482 gnd.n1481 71.676
R9031 gnd.n1477 gnd.n1476 71.676
R9032 gnd.n1474 gnd.n1473 71.676
R9033 gnd.n1469 gnd.n1468 71.676
R9034 gnd.n1466 gnd.n1465 71.676
R9035 gnd.n1461 gnd.n1460 71.676
R9036 gnd.n1456 gnd.n1453 71.676
R9037 gnd.n1604 gnd.n1603 71.676
R9038 gnd.n1601 gnd.n1600 71.676
R9039 gnd.n1595 gnd.n1594 71.676
R9040 gnd.n1592 gnd.n1591 71.676
R9041 gnd.n1587 gnd.n1586 71.676
R9042 gnd.n1584 gnd.n1583 71.676
R9043 gnd.n1579 gnd.n1578 71.676
R9044 gnd.n1576 gnd.n1575 71.676
R9045 gnd.n1571 gnd.n1570 71.676
R9046 gnd.n1568 gnd.n1567 71.676
R9047 gnd.n1563 gnd.n1562 71.676
R9048 gnd.n1560 gnd.n1559 71.676
R9049 gnd.n1555 gnd.n1554 71.676
R9050 gnd.n1552 gnd.n1551 71.676
R9051 gnd.n1547 gnd.n1546 71.676
R9052 gnd.n1544 gnd.n1543 71.676
R9053 gnd.n1539 gnd.n1538 71.676
R9054 gnd.n864 gnd.n863 71.676
R9055 gnd.n859 gnd.n678 71.676
R9056 gnd.n857 gnd.n856 71.676
R9057 gnd.n852 gnd.n851 71.676
R9058 gnd.n849 gnd.n848 71.676
R9059 gnd.n844 gnd.n843 71.676
R9060 gnd.n841 gnd.n840 71.676
R9061 gnd.n836 gnd.n835 71.676
R9062 gnd.n833 gnd.n832 71.676
R9063 gnd.n828 gnd.n827 71.676
R9064 gnd.n825 gnd.n824 71.676
R9065 gnd.n820 gnd.n819 71.676
R9066 gnd.n817 gnd.n816 71.676
R9067 gnd.n812 gnd.n811 71.676
R9068 gnd.n809 gnd.n808 71.676
R9069 gnd.n801 gnd.n800 71.676
R9070 gnd.n797 gnd.n796 71.676
R9071 gnd.n792 gnd.n693 71.676
R9072 gnd.n790 gnd.n789 71.676
R9073 gnd.n782 gnd.n781 71.676
R9074 gnd.n779 gnd.n778 71.676
R9075 gnd.n774 gnd.n773 71.676
R9076 gnd.n771 gnd.n770 71.676
R9077 gnd.n766 gnd.n765 71.676
R9078 gnd.n763 gnd.n762 71.676
R9079 gnd.n758 gnd.n757 71.676
R9080 gnd.n755 gnd.n754 71.676
R9081 gnd.n750 gnd.n749 71.676
R9082 gnd.n747 gnd.n746 71.676
R9083 gnd.n742 gnd.n741 71.676
R9084 gnd.n739 gnd.n738 71.676
R9085 gnd.n734 gnd.n733 71.676
R9086 gnd.n731 gnd.n730 71.676
R9087 gnd.n8 gnd.t142 69.1507
R9088 gnd.n14 gnd.t355 68.4792
R9089 gnd.n13 gnd.t347 68.4792
R9090 gnd.n12 gnd.t153 68.4792
R9091 gnd.n11 gnd.t26 68.4792
R9092 gnd.n10 gnd.t156 68.4792
R9093 gnd.n9 gnd.t339 68.4792
R9094 gnd.n8 gnd.t171 68.4792
R9095 gnd.n3966 gnd.n3870 64.369
R9096 gnd.n1597 gnd.n1395 59.5399
R9097 gnd.n806 gnd.n805 59.5399
R9098 gnd.n1452 gnd.n1451 59.5399
R9099 gnd.n787 gnd.n786 59.5399
R9100 gnd.n1434 gnd.n1433 59.1804
R9101 gnd.n4755 gnd.n1988 57.3586
R9102 gnd.n3657 gnd.t181 56.607
R9103 gnd.n56 gnd.t309 56.607
R9104 gnd.n3618 gnd.t264 56.407
R9105 gnd.n3637 gnd.t236 56.407
R9106 gnd.n17 gnd.t304 56.407
R9107 gnd.n36 gnd.t275 56.407
R9108 gnd.n3674 gnd.t246 55.8337
R9109 gnd.n3635 gnd.t288 55.8337
R9110 gnd.n3654 gnd.t261 55.8337
R9111 gnd.n73 gnd.t320 55.8337
R9112 gnd.n34 gnd.t302 55.8337
R9113 gnd.n53 gnd.t272 55.8337
R9114 gnd.n1421 gnd.n1420 54.358
R9115 gnd.n721 gnd.n720 54.358
R9116 gnd.n2656 gnd.n236 53.6263
R9117 gnd.n3657 gnd.n3656 53.0052
R9118 gnd.n3659 gnd.n3658 53.0052
R9119 gnd.n3661 gnd.n3660 53.0052
R9120 gnd.n3663 gnd.n3662 53.0052
R9121 gnd.n3665 gnd.n3664 53.0052
R9122 gnd.n3667 gnd.n3666 53.0052
R9123 gnd.n3669 gnd.n3668 53.0052
R9124 gnd.n3671 gnd.n3670 53.0052
R9125 gnd.n3673 gnd.n3672 53.0052
R9126 gnd.n3618 gnd.n3617 53.0052
R9127 gnd.n3620 gnd.n3619 53.0052
R9128 gnd.n3622 gnd.n3621 53.0052
R9129 gnd.n3624 gnd.n3623 53.0052
R9130 gnd.n3626 gnd.n3625 53.0052
R9131 gnd.n3628 gnd.n3627 53.0052
R9132 gnd.n3630 gnd.n3629 53.0052
R9133 gnd.n3632 gnd.n3631 53.0052
R9134 gnd.n3634 gnd.n3633 53.0052
R9135 gnd.n3637 gnd.n3636 53.0052
R9136 gnd.n3639 gnd.n3638 53.0052
R9137 gnd.n3641 gnd.n3640 53.0052
R9138 gnd.n3643 gnd.n3642 53.0052
R9139 gnd.n3645 gnd.n3644 53.0052
R9140 gnd.n3647 gnd.n3646 53.0052
R9141 gnd.n3649 gnd.n3648 53.0052
R9142 gnd.n3651 gnd.n3650 53.0052
R9143 gnd.n3653 gnd.n3652 53.0052
R9144 gnd.n72 gnd.n71 53.0052
R9145 gnd.n70 gnd.n69 53.0052
R9146 gnd.n68 gnd.n67 53.0052
R9147 gnd.n66 gnd.n65 53.0052
R9148 gnd.n64 gnd.n63 53.0052
R9149 gnd.n62 gnd.n61 53.0052
R9150 gnd.n60 gnd.n59 53.0052
R9151 gnd.n58 gnd.n57 53.0052
R9152 gnd.n56 gnd.n55 53.0052
R9153 gnd.n33 gnd.n32 53.0052
R9154 gnd.n31 gnd.n30 53.0052
R9155 gnd.n29 gnd.n28 53.0052
R9156 gnd.n27 gnd.n26 53.0052
R9157 gnd.n25 gnd.n24 53.0052
R9158 gnd.n23 gnd.n22 53.0052
R9159 gnd.n21 gnd.n20 53.0052
R9160 gnd.n19 gnd.n18 53.0052
R9161 gnd.n17 gnd.n16 53.0052
R9162 gnd.n52 gnd.n51 53.0052
R9163 gnd.n50 gnd.n49 53.0052
R9164 gnd.n48 gnd.n47 53.0052
R9165 gnd.n46 gnd.n45 53.0052
R9166 gnd.n44 gnd.n43 53.0052
R9167 gnd.n42 gnd.n41 53.0052
R9168 gnd.n40 gnd.n39 53.0052
R9169 gnd.n38 gnd.n37 53.0052
R9170 gnd.n36 gnd.n35 53.0052
R9171 gnd.n712 gnd.n711 52.4801
R9172 gnd.n4609 gnd.t24 52.3082
R9173 gnd.n4577 gnd.t160 52.3082
R9174 gnd.n4545 gnd.t140 52.3082
R9175 gnd.n4514 gnd.t341 52.3082
R9176 gnd.n4482 gnd.t138 52.3082
R9177 gnd.n4450 gnd.t349 52.3082
R9178 gnd.n4418 gnd.t147 52.3082
R9179 gnd.n4387 gnd.t158 52.3082
R9180 gnd.n5070 gnd.n4756 51.6227
R9181 gnd.n7573 gnd.n124 51.6227
R9182 gnd.n4439 gnd.n4407 51.4173
R9183 gnd.n4503 gnd.n4502 50.455
R9184 gnd.n4471 gnd.n4470 50.455
R9185 gnd.n4439 gnd.n4438 50.455
R9186 gnd.n7018 gnd.n534 45.6325
R9187 gnd.n1606 gnd.n1605 45.6325
R9188 gnd.n3913 gnd.n3912 45.1884
R9189 gnd.n2054 gnd.n2053 45.1884
R9190 gnd.n728 gnd.n727 44.3322
R9191 gnd.n1424 gnd.n1423 44.3189
R9192 gnd.n5800 gnd.n1337 42.2793
R9193 gnd.n3914 gnd.n3913 42.2793
R9194 gnd.n2055 gnd.n2054 42.2793
R9195 gnd.n3840 gnd.n3839 42.2793
R9196 gnd.n4722 gnd.n2028 42.2793
R9197 gnd.n120 gnd.n119 42.2793
R9198 gnd.n6714 gnd.n6713 42.2793
R9199 gnd.n5775 gnd.n1349 42.2793
R9200 gnd.n561 gnd.n560 42.2793
R9201 gnd.n7501 gnd.n198 42.2793
R9202 gnd.n7538 gnd.n7537 42.2793
R9203 gnd.n4902 gnd.n4901 42.2793
R9204 gnd.n4934 gnd.n4933 42.2793
R9205 gnd.n4763 gnd.n4762 42.2793
R9206 gnd.n1643 gnd.n1642 42.2793
R9207 gnd.n6691 gnd.n6690 42.2793
R9208 gnd.n1422 gnd.n1421 41.6274
R9209 gnd.n722 gnd.n721 41.6274
R9210 gnd.n1431 gnd.n1430 40.8975
R9211 gnd.n725 gnd.n724 40.8975
R9212 gnd.n7018 gnd.n538 36.9518
R9213 gnd.n1606 gnd.n1389 36.9518
R9214 gnd.n1430 gnd.n1429 35.055
R9215 gnd.n1425 gnd.n1424 35.055
R9216 gnd.n714 gnd.n713 35.055
R9217 gnd.n724 gnd.n710 35.055
R9218 gnd.n867 gnd.n866 32.9371
R9219 gnd.n1540 gnd.n1410 32.9371
R9220 gnd.n3143 gnd.n3142 32.6173
R9221 gnd.n3143 gnd.n2183 32.6173
R9222 gnd.n3151 gnd.n2183 32.6173
R9223 gnd.n3152 gnd.n3151 32.6173
R9224 gnd.n3153 gnd.n3152 32.6173
R9225 gnd.n3153 gnd.n2177 32.6173
R9226 gnd.n3161 gnd.n2177 32.6173
R9227 gnd.n3162 gnd.n3161 32.6173
R9228 gnd.n3163 gnd.n3162 32.6173
R9229 gnd.n3163 gnd.n2171 32.6173
R9230 gnd.n3171 gnd.n2171 32.6173
R9231 gnd.n3172 gnd.n3171 32.6173
R9232 gnd.n3173 gnd.n3172 32.6173
R9233 gnd.n3173 gnd.n2165 32.6173
R9234 gnd.n3181 gnd.n2165 32.6173
R9235 gnd.n3182 gnd.n3181 32.6173
R9236 gnd.n3183 gnd.n3182 32.6173
R9237 gnd.n3183 gnd.n2159 32.6173
R9238 gnd.n3191 gnd.n2159 32.6173
R9239 gnd.n3192 gnd.n3191 32.6173
R9240 gnd.n3193 gnd.n3192 32.6173
R9241 gnd.n3193 gnd.n2153 32.6173
R9242 gnd.n3201 gnd.n2153 32.6173
R9243 gnd.n3202 gnd.n3201 32.6173
R9244 gnd.n3203 gnd.n3202 32.6173
R9245 gnd.n3203 gnd.n2147 32.6173
R9246 gnd.n3211 gnd.n2147 32.6173
R9247 gnd.n3212 gnd.n3211 32.6173
R9248 gnd.n3213 gnd.n3212 32.6173
R9249 gnd.n3213 gnd.n2141 32.6173
R9250 gnd.n3221 gnd.n2141 32.6173
R9251 gnd.n3222 gnd.n3221 32.6173
R9252 gnd.n3223 gnd.n3222 32.6173
R9253 gnd.n3223 gnd.n2135 32.6173
R9254 gnd.n3231 gnd.n2135 32.6173
R9255 gnd.n3232 gnd.n3231 32.6173
R9256 gnd.n3233 gnd.n3232 32.6173
R9257 gnd.n3233 gnd.n2129 32.6173
R9258 gnd.n3241 gnd.n2129 32.6173
R9259 gnd.n3242 gnd.n3241 32.6173
R9260 gnd.n3243 gnd.n3242 32.6173
R9261 gnd.n3243 gnd.n2123 32.6173
R9262 gnd.n3251 gnd.n2123 32.6173
R9263 gnd.n3252 gnd.n3251 32.6173
R9264 gnd.n3253 gnd.n3252 32.6173
R9265 gnd.n3253 gnd.n2117 32.6173
R9266 gnd.n3261 gnd.n2117 32.6173
R9267 gnd.n3262 gnd.n3261 32.6173
R9268 gnd.n3263 gnd.n3262 32.6173
R9269 gnd.n3263 gnd.n2111 32.6173
R9270 gnd.n3271 gnd.n2111 32.6173
R9271 gnd.n3272 gnd.n3271 32.6173
R9272 gnd.n3273 gnd.n3272 32.6173
R9273 gnd.n3273 gnd.n2105 32.6173
R9274 gnd.n3281 gnd.n2105 32.6173
R9275 gnd.n3282 gnd.n3281 32.6173
R9276 gnd.n3283 gnd.n3282 32.6173
R9277 gnd.n3283 gnd.n2099 32.6173
R9278 gnd.n3291 gnd.n2099 32.6173
R9279 gnd.n3292 gnd.n3291 32.6173
R9280 gnd.n3293 gnd.n3292 32.6173
R9281 gnd.n3293 gnd.n2093 32.6173
R9282 gnd.n3301 gnd.n2093 32.6173
R9283 gnd.n3302 gnd.n3301 32.6173
R9284 gnd.n3303 gnd.n3302 32.6173
R9285 gnd.n3303 gnd.n2087 32.6173
R9286 gnd.n3311 gnd.n2087 32.6173
R9287 gnd.n3312 gnd.n3311 32.6173
R9288 gnd.n3313 gnd.n3312 32.6173
R9289 gnd.n3313 gnd.n2081 32.6173
R9290 gnd.n3321 gnd.n2081 32.6173
R9291 gnd.n3322 gnd.n3321 32.6173
R9292 gnd.n3323 gnd.n3322 32.6173
R9293 gnd.n3323 gnd.n2075 32.6173
R9294 gnd.n3331 gnd.n2075 32.6173
R9295 gnd.n3332 gnd.n3331 32.6173
R9296 gnd.n3333 gnd.n3332 32.6173
R9297 gnd.n3333 gnd.n2069 32.6173
R9298 gnd.n3341 gnd.n2069 32.6173
R9299 gnd.n3342 gnd.n3341 32.6173
R9300 gnd.n3343 gnd.n3342 32.6173
R9301 gnd.n3343 gnd.n2062 32.6173
R9302 gnd.n3354 gnd.n2062 32.6173
R9303 gnd.n3976 gnd.n3870 31.8661
R9304 gnd.n3976 gnd.n3975 31.8661
R9305 gnd.n3984 gnd.n3859 31.8661
R9306 gnd.n3992 gnd.n3859 31.8661
R9307 gnd.n3992 gnd.n3853 31.8661
R9308 gnd.n4000 gnd.n3853 31.8661
R9309 gnd.n4000 gnd.n3846 31.8661
R9310 gnd.n4038 gnd.n3846 31.8661
R9311 gnd.n4048 gnd.n3779 31.8661
R9312 gnd.n5070 gnd.n4872 31.8661
R9313 gnd.n5078 gnd.n1974 31.8661
R9314 gnd.n5086 gnd.n1974 31.8661
R9315 gnd.n5086 gnd.n1966 31.8661
R9316 gnd.n5094 gnd.n1966 31.8661
R9317 gnd.n5102 gnd.n1957 31.8661
R9318 gnd.n5102 gnd.n1960 31.8661
R9319 gnd.n5110 gnd.n1942 31.8661
R9320 gnd.n5118 gnd.n1942 31.8661
R9321 gnd.n5126 gnd.n1934 31.8661
R9322 gnd.n5134 gnd.n1925 31.8661
R9323 gnd.n5134 gnd.n1928 31.8661
R9324 gnd.n5150 gnd.n1908 31.8661
R9325 gnd.n5160 gnd.n1908 31.8661
R9326 gnd.n5173 gnd.n1902 31.8661
R9327 gnd.n5190 gnd.n1884 31.8661
R9328 gnd.n5184 gnd.n1884 31.8661
R9329 gnd.n5199 gnd.n1867 31.8661
R9330 gnd.n5217 gnd.n1867 31.8661
R9331 gnd.n5461 gnd.n1775 31.8661
R9332 gnd.n5455 gnd.n1786 31.8661
R9333 gnd.n5358 gnd.n1356 31.8661
R9334 gnd.n5351 gnd.n1318 31.8661
R9335 gnd.n5809 gnd.n1318 31.8661
R9336 gnd.n5809 gnd.n1310 31.8661
R9337 gnd.n5817 gnd.n1310 31.8661
R9338 gnd.n5817 gnd.n1312 31.8661
R9339 gnd.n6808 gnd.n639 31.8661
R9340 gnd.n639 gnd.n616 31.8661
R9341 gnd.n6817 gnd.n616 31.8661
R9342 gnd.n6817 gnd.n6816 31.8661
R9343 gnd.n6816 gnd.n489 31.8661
R9344 gnd.n564 gnd.n518 31.8661
R9345 gnd.n7228 gnd.n336 31.8661
R9346 gnd.n7301 gnd.n330 31.8661
R9347 gnd.n7305 gnd.n295 31.8661
R9348 gnd.n7329 gnd.n295 31.8661
R9349 gnd.n7337 gnd.n286 31.8661
R9350 gnd.n7337 gnd.n289 31.8661
R9351 gnd.n7345 gnd.n280 31.8661
R9352 gnd.n7353 gnd.n265 31.8661
R9353 gnd.n7361 gnd.n265 31.8661
R9354 gnd.n7369 gnd.n256 31.8661
R9355 gnd.n7369 gnd.n259 31.8661
R9356 gnd.n7377 gnd.n250 31.8661
R9357 gnd.n7385 gnd.n234 31.8661
R9358 gnd.n7393 gnd.n234 31.8661
R9359 gnd.n7401 gnd.n225 31.8661
R9360 gnd.n7401 gnd.n228 31.8661
R9361 gnd.n7409 gnd.n209 31.8661
R9362 gnd.n7485 gnd.n209 31.8661
R9363 gnd.n7485 gnd.n202 31.8661
R9364 gnd.n7493 gnd.n202 31.8661
R9365 gnd.n7573 gnd.n122 31.8661
R9366 gnd.n5461 gnd.t234 31.5474
R9367 gnd.n7301 gnd.t300 31.5474
R9368 gnd.t269 gnd.n1902 30.9101
R9369 gnd.n280 gnd.t225 30.9101
R9370 gnd.t213 gnd.n1934 30.2728
R9371 gnd.n250 gnd.t196 30.2728
R9372 gnd.n4872 gnd.t38 28.3609
R9373 gnd.t45 gnd.n122 28.3609
R9374 gnd.n5351 gnd.n1364 27.4049
R9375 gnd.n7046 gnd.n489 27.4049
R9376 gnd.n1337 gnd.n1336 25.7944
R9377 gnd.n3839 gnd.n3838 25.7944
R9378 gnd.n2028 gnd.n2027 25.7944
R9379 gnd.n119 gnd.n118 25.7944
R9380 gnd.n6713 gnd.n6712 25.7944
R9381 gnd.n1349 gnd.n1348 25.7944
R9382 gnd.n538 gnd.n537 25.7944
R9383 gnd.n560 gnd.n559 25.7944
R9384 gnd.n198 gnd.n197 25.7944
R9385 gnd.n7537 gnd.n7536 25.7944
R9386 gnd.n4901 gnd.n4900 25.7944
R9387 gnd.n4933 gnd.n4932 25.7944
R9388 gnd.n4762 gnd.n4761 25.7944
R9389 gnd.n1642 gnd.n1641 25.7944
R9390 gnd.n1389 gnd.n1388 25.7944
R9391 gnd.n6690 gnd.n6689 25.7944
R9392 gnd.n4060 gnd.n3780 24.8557
R9393 gnd.n4070 gnd.n3763 24.8557
R9394 gnd.n3766 gnd.n3754 24.8557
R9395 gnd.n4091 gnd.n3755 24.8557
R9396 gnd.n4101 gnd.n3735 24.8557
R9397 gnd.n4111 gnd.n4110 24.8557
R9398 gnd.n3719 gnd.n3718 24.8557
R9399 gnd.n4148 gnd.n3711 24.8557
R9400 gnd.n4147 gnd.n3704 24.8557
R9401 gnd.n4185 gnd.n3683 24.8557
R9402 gnd.n4159 gnd.n3684 24.8557
R9403 gnd.n4178 gnd.n3531 24.8557
R9404 gnd.n4195 gnd.n4194 24.8557
R9405 gnd.n4206 gnd.n4205 24.8557
R9406 gnd.n3523 gnd.n3514 24.8557
R9407 gnd.n4226 gnd.n3497 24.8557
R9408 gnd.n3500 gnd.n3489 24.8557
R9409 gnd.n4247 gnd.n3490 24.8557
R9410 gnd.n4256 gnd.n3482 24.8557
R9411 gnd.n4257 gnd.n3471 24.8557
R9412 gnd.n3474 gnd.n3462 24.8557
R9413 gnd.n4278 gnd.n3463 24.8557
R9414 gnd.n4288 gnd.n3446 24.8557
R9415 gnd.n4299 gnd.n4298 24.8557
R9416 gnd.n3588 gnd.n3587 24.8557
R9417 gnd.n4309 gnd.n3438 24.8557
R9418 gnd.n4319 gnd.n3421 24.8557
R9419 gnd.n4330 gnd.n4329 24.8557
R9420 gnd.n4340 gnd.n3413 24.8557
R9421 gnd.n4350 gnd.n3395 24.8557
R9422 gnd.n4361 gnd.n4360 24.8557
R9423 gnd.n4371 gnd.n3388 24.8557
R9424 gnd.n4636 gnd.n3380 24.8557
R9425 gnd.n4637 gnd.n3370 24.8557
R9426 gnd.n1395 gnd.n1394 23.855
R9427 gnd.n805 gnd.n804 23.855
R9428 gnd.n1451 gnd.n1450 23.855
R9429 gnd.n786 gnd.n785 23.855
R9430 gnd.n4081 gnd.t157 23.2624
R9431 gnd.n5094 gnd.t245 23.2624
R9432 gnd.n5677 gnd.n1305 23.2624
R9433 gnd.n6798 gnd.n648 23.2624
R9434 gnd.n7409 gnd.t271 23.2624
R9435 gnd.n3782 gnd.t34 22.6251
R9436 gnd.n5126 gnd.t217 22.6251
R9437 gnd.n7377 gnd.t182 22.6251
R9438 gnd.n5173 gnd.t190 21.9878
R9439 gnd.n7345 gnd.t240 21.9878
R9440 gnd.n5983 gnd.n1264 21.6691
R9441 gnd.n5975 gnd.n1256 21.6691
R9442 gnd.n5911 gnd.n1241 21.6691
R9443 gnd.n5927 gnd.n1225 21.6691
R9444 gnd.n5947 gnd.n1218 21.6691
R9445 gnd.n6125 gnd.n1111 21.6691
R9446 gnd.n6110 gnd.n1095 21.6691
R9447 gnd.n6102 gnd.n1087 21.6691
R9448 gnd.n6095 gnd.n1080 21.6691
R9449 gnd.n6087 gnd.n1149 21.6691
R9450 gnd.n6081 gnd.n6080 21.6691
R9451 gnd.n6430 gnd.n1022 21.6691
R9452 gnd.n6430 gnd.n1025 21.6691
R9453 gnd.n6415 gnd.n1008 21.6691
R9454 gnd.n6289 gnd.n1000 21.6691
R9455 gnd.n6267 gnd.n992 21.6691
R9456 gnd.n6307 gnd.n984 21.6691
R9457 gnd.n6316 gnd.n6256 21.6691
R9458 gnd.n6335 gnd.n6247 21.6691
R9459 gnd.n6352 gnd.n937 21.6691
R9460 gnd.n6380 gnd.n928 21.6691
R9461 gnd.n6552 gnd.n911 21.6691
R9462 gnd.n6569 gnd.n880 21.6691
R9463 gnd.n6769 gnd.n655 21.6691
R9464 gnd.t340 gnd.n3787 21.3504
R9465 gnd.t194 gnd.n1775 21.3504
R9466 gnd.n1788 gnd.n1786 21.3504
R9467 gnd.n5233 gnd.t215 21.3504
R9468 gnd.n7202 gnd.t206 21.3504
R9469 gnd.n7221 gnd.n336 21.3504
R9470 gnd.t289 gnd.n330 21.3504
R9471 gnd.n1518 gnd.n1434 20.7615
R9472 gnd.n728 gnd.n674 20.7615
R9473 gnd.t9 gnd.n3412 20.7131
R9474 gnd.n5199 gnd.t231 20.7131
R9475 gnd.n7329 gnd.t250 20.7131
R9476 gnd.t31 gnd.n1297 20.3945
R9477 gnd.n1411 gnd.n1287 20.3945
R9478 gnd.n5991 gnd.n1254 20.3945
R9479 gnd.n5939 gnd.n1199 20.3945
R9480 gnd.n6133 gnd.n1101 20.3945
R9481 gnd.n1163 gnd.n1049 20.3945
R9482 gnd.n6438 gnd.n1014 20.3945
R9483 gnd.n6325 gnd.n961 20.3945
R9484 gnd.n6242 gnd.n955 20.3945
R9485 gnd.n4287 gnd.t11 20.0758
R9486 gnd.n5150 gnd.t252 20.0758
R9487 gnd.t354 gnd.t63 20.0758
R9488 gnd.n7361 gnd.t282 20.0758
R9489 gnd.n1418 gnd.t131 19.8005
R9490 gnd.n1418 gnd.t43 19.8005
R9491 gnd.n1419 gnd.t32 19.8005
R9492 gnd.n1419 gnd.t61 19.8005
R9493 gnd.n718 gnd.t89 19.8005
R9494 gnd.n718 gnd.t54 19.8005
R9495 gnd.n719 gnd.t102 19.8005
R9496 gnd.n719 gnd.t29 19.8005
R9497 gnd.n3355 gnd.n3354 19.5706
R9498 gnd.n1415 gnd.n1414 19.5087
R9499 gnd.n1428 gnd.n1415 19.5087
R9500 gnd.n1426 gnd.n1417 19.5087
R9501 gnd.n723 gnd.n717 19.5087
R9502 gnd.t13 gnd.n4236 19.4385
R9503 gnd.n5110 gnd.t192 19.4385
R9504 gnd.n5819 gnd.n1307 19.3944
R9505 gnd.n5823 gnd.n1307 19.3944
R9506 gnd.n5823 gnd.n1293 19.3944
R9507 gnd.n5837 gnd.n1293 19.3944
R9508 gnd.n5837 gnd.n1290 19.3944
R9509 gnd.n5842 gnd.n1290 19.3944
R9510 gnd.n5842 gnd.n1291 19.3944
R9511 gnd.n1291 gnd.n1252 19.3944
R9512 gnd.n5993 gnd.n1252 19.3944
R9513 gnd.n5993 gnd.n1250 19.3944
R9514 gnd.n5997 gnd.n1250 19.3944
R9515 gnd.n5997 gnd.n1237 19.3944
R9516 gnd.n6009 gnd.n1237 19.3944
R9517 gnd.n6009 gnd.n1235 19.3944
R9518 gnd.n6013 gnd.n1235 19.3944
R9519 gnd.n6013 gnd.n1222 19.3944
R9520 gnd.n6025 gnd.n1222 19.3944
R9521 gnd.n6025 gnd.n1220 19.3944
R9522 gnd.n6029 gnd.n1220 19.3944
R9523 gnd.n6029 gnd.n1205 19.3944
R9524 gnd.n6042 gnd.n1205 19.3944
R9525 gnd.n6042 gnd.n1202 19.3944
R9526 gnd.n6047 gnd.n1202 19.3944
R9527 gnd.n6047 gnd.n1203 19.3944
R9528 gnd.n1203 gnd.n1099 19.3944
R9529 gnd.n6135 gnd.n1099 19.3944
R9530 gnd.n6135 gnd.n1097 19.3944
R9531 gnd.n6139 gnd.n1097 19.3944
R9532 gnd.n6139 gnd.n1084 19.3944
R9533 gnd.n6151 gnd.n1084 19.3944
R9534 gnd.n6151 gnd.n1082 19.3944
R9535 gnd.n6155 gnd.n1082 19.3944
R9536 gnd.n6155 gnd.n1070 19.3944
R9537 gnd.n6167 gnd.n1070 19.3944
R9538 gnd.n6167 gnd.n1068 19.3944
R9539 gnd.n6171 gnd.n1068 19.3944
R9540 gnd.n6171 gnd.n1054 19.3944
R9541 gnd.n6185 gnd.n1054 19.3944
R9542 gnd.n6185 gnd.n1051 19.3944
R9543 gnd.n6190 gnd.n1051 19.3944
R9544 gnd.n6190 gnd.n1052 19.3944
R9545 gnd.n1052 gnd.n1012 19.3944
R9546 gnd.n6440 gnd.n1012 19.3944
R9547 gnd.n6440 gnd.n1010 19.3944
R9548 gnd.n6444 gnd.n1010 19.3944
R9549 gnd.n6444 gnd.n996 19.3944
R9550 gnd.n6456 gnd.n996 19.3944
R9551 gnd.n6456 gnd.n994 19.3944
R9552 gnd.n6460 gnd.n994 19.3944
R9553 gnd.n6460 gnd.n981 19.3944
R9554 gnd.n6472 gnd.n981 19.3944
R9555 gnd.n6472 gnd.n979 19.3944
R9556 gnd.n6476 gnd.n979 19.3944
R9557 gnd.n6476 gnd.n966 19.3944
R9558 gnd.n6488 gnd.n966 19.3944
R9559 gnd.n6488 gnd.n964 19.3944
R9560 gnd.n6492 gnd.n964 19.3944
R9561 gnd.n6492 gnd.n951 19.3944
R9562 gnd.n6504 gnd.n951 19.3944
R9563 gnd.n6504 gnd.n949 19.3944
R9564 gnd.n6508 gnd.n949 19.3944
R9565 gnd.n6508 gnd.n935 19.3944
R9566 gnd.n6519 gnd.n935 19.3944
R9567 gnd.n6519 gnd.n932 19.3944
R9568 gnd.n6530 gnd.n932 19.3944
R9569 gnd.n6530 gnd.n933 19.3944
R9570 gnd.n6526 gnd.n933 19.3944
R9571 gnd.n6526 gnd.n6525 19.3944
R9572 gnd.n6525 gnd.n893 19.3944
R9573 gnd.n6588 gnd.n893 19.3944
R9574 gnd.n6588 gnd.n894 19.3944
R9575 gnd.n6584 gnd.n894 19.3944
R9576 gnd.n6584 gnd.n6583 19.3944
R9577 gnd.n6583 gnd.n6582 19.3944
R9578 gnd.n6582 gnd.n6579 19.3944
R9579 gnd.n6579 gnd.n652 19.3944
R9580 gnd.n6791 gnd.n652 19.3944
R9581 gnd.n6791 gnd.n650 19.3944
R9582 gnd.n6796 gnd.n650 19.3944
R9583 gnd.n6796 gnd.n636 19.3944
R9584 gnd.n6810 gnd.n636 19.3944
R9585 gnd.n6811 gnd.n6810 19.3944
R9586 gnd.n5802 gnd.n1333 19.3944
R9587 gnd.n5806 gnd.n1333 19.3944
R9588 gnd.n5806 gnd.n1334 19.3944
R9589 gnd.n5669 gnd.n5582 19.3944
R9590 gnd.n5669 gnd.n5668 19.3944
R9591 gnd.n5668 gnd.n5585 19.3944
R9592 gnd.n5661 gnd.n5585 19.3944
R9593 gnd.n5661 gnd.n5660 19.3944
R9594 gnd.n5660 gnd.n5597 19.3944
R9595 gnd.n5653 gnd.n5597 19.3944
R9596 gnd.n5653 gnd.n5652 19.3944
R9597 gnd.n5652 gnd.n5608 19.3944
R9598 gnd.n5645 gnd.n5608 19.3944
R9599 gnd.n5645 gnd.n5644 19.3944
R9600 gnd.n5644 gnd.n5620 19.3944
R9601 gnd.n5637 gnd.n5620 19.3944
R9602 gnd.n5637 gnd.n5636 19.3944
R9603 gnd.n5636 gnd.n1343 19.3944
R9604 gnd.n5778 gnd.n1343 19.3944
R9605 gnd.n5781 gnd.n5778 19.3944
R9606 gnd.n5781 gnd.n1340 19.3944
R9607 gnd.n5786 gnd.n1340 19.3944
R9608 gnd.n5789 gnd.n5786 19.3944
R9609 gnd.n5792 gnd.n5789 19.3944
R9610 gnd.n5792 gnd.n1338 19.3944
R9611 gnd.n5796 gnd.n1338 19.3944
R9612 gnd.n5799 gnd.n5796 19.3944
R9613 gnd.n3963 gnd.n3962 19.3944
R9614 gnd.n3962 gnd.n3961 19.3944
R9615 gnd.n3961 gnd.n3960 19.3944
R9616 gnd.n3960 gnd.n3958 19.3944
R9617 gnd.n3958 gnd.n3955 19.3944
R9618 gnd.n3955 gnd.n3954 19.3944
R9619 gnd.n3954 gnd.n3951 19.3944
R9620 gnd.n3951 gnd.n3950 19.3944
R9621 gnd.n3950 gnd.n3947 19.3944
R9622 gnd.n3947 gnd.n3946 19.3944
R9623 gnd.n3946 gnd.n3943 19.3944
R9624 gnd.n3943 gnd.n3942 19.3944
R9625 gnd.n3942 gnd.n3939 19.3944
R9626 gnd.n3939 gnd.n3938 19.3944
R9627 gnd.n3938 gnd.n3935 19.3944
R9628 gnd.n3935 gnd.n3934 19.3944
R9629 gnd.n3934 gnd.n3931 19.3944
R9630 gnd.n3931 gnd.n3930 19.3944
R9631 gnd.n3930 gnd.n3927 19.3944
R9632 gnd.n3927 gnd.n3926 19.3944
R9633 gnd.n3926 gnd.n3923 19.3944
R9634 gnd.n3923 gnd.n3922 19.3944
R9635 gnd.n3919 gnd.n3918 19.3944
R9636 gnd.n3918 gnd.n3874 19.3944
R9637 gnd.n3969 gnd.n3874 19.3944
R9638 gnd.n4672 gnd.n4671 19.3944
R9639 gnd.n4671 gnd.n4668 19.3944
R9640 gnd.n4668 gnd.n4667 19.3944
R9641 gnd.n4717 gnd.n4716 19.3944
R9642 gnd.n4716 gnd.n4715 19.3944
R9643 gnd.n4715 gnd.n4712 19.3944
R9644 gnd.n4712 gnd.n4711 19.3944
R9645 gnd.n4711 gnd.n4708 19.3944
R9646 gnd.n4708 gnd.n4707 19.3944
R9647 gnd.n4707 gnd.n4704 19.3944
R9648 gnd.n4704 gnd.n4703 19.3944
R9649 gnd.n4703 gnd.n4700 19.3944
R9650 gnd.n4700 gnd.n4699 19.3944
R9651 gnd.n4699 gnd.n4696 19.3944
R9652 gnd.n4696 gnd.n4695 19.3944
R9653 gnd.n4695 gnd.n4692 19.3944
R9654 gnd.n4692 gnd.n4691 19.3944
R9655 gnd.n4691 gnd.n4688 19.3944
R9656 gnd.n4688 gnd.n4687 19.3944
R9657 gnd.n4687 gnd.n4684 19.3944
R9658 gnd.n4684 gnd.n4683 19.3944
R9659 gnd.n4683 gnd.n4680 19.3944
R9660 gnd.n4680 gnd.n4679 19.3944
R9661 gnd.n4679 gnd.n4676 19.3944
R9662 gnd.n4676 gnd.n4675 19.3944
R9663 gnd.n4062 gnd.n3771 19.3944
R9664 gnd.n4072 gnd.n3771 19.3944
R9665 gnd.n4073 gnd.n4072 19.3944
R9666 gnd.n4073 gnd.n3752 19.3944
R9667 gnd.n4093 gnd.n3752 19.3944
R9668 gnd.n4093 gnd.n3744 19.3944
R9669 gnd.n4103 gnd.n3744 19.3944
R9670 gnd.n4104 gnd.n4103 19.3944
R9671 gnd.n4105 gnd.n4104 19.3944
R9672 gnd.n4105 gnd.n3727 19.3944
R9673 gnd.n3727 gnd.n3725 19.3944
R9674 gnd.n4131 gnd.n3725 19.3944
R9675 gnd.n4131 gnd.n3707 19.3944
R9676 gnd.n4165 gnd.n3707 19.3944
R9677 gnd.n4165 gnd.n4164 19.3944
R9678 gnd.n4164 gnd.n4163 19.3944
R9679 gnd.n4163 gnd.n4158 19.3944
R9680 gnd.n4158 gnd.n3528 19.3944
R9681 gnd.n4197 gnd.n3528 19.3944
R9682 gnd.n4198 gnd.n4197 19.3944
R9683 gnd.n4198 gnd.n3512 19.3944
R9684 gnd.n4218 gnd.n3512 19.3944
R9685 gnd.n4218 gnd.n3505 19.3944
R9686 gnd.n4228 gnd.n3505 19.3944
R9687 gnd.n4229 gnd.n4228 19.3944
R9688 gnd.n4229 gnd.n3487 19.3944
R9689 gnd.n4249 gnd.n3487 19.3944
R9690 gnd.n4249 gnd.n3479 19.3944
R9691 gnd.n4259 gnd.n3479 19.3944
R9692 gnd.n4260 gnd.n4259 19.3944
R9693 gnd.n4260 gnd.n3460 19.3944
R9694 gnd.n4280 gnd.n3460 19.3944
R9695 gnd.n4280 gnd.n3453 19.3944
R9696 gnd.n4290 gnd.n3453 19.3944
R9697 gnd.n4291 gnd.n4290 19.3944
R9698 gnd.n4291 gnd.n3436 19.3944
R9699 gnd.n4311 gnd.n3436 19.3944
R9700 gnd.n4311 gnd.n3429 19.3944
R9701 gnd.n4321 gnd.n3429 19.3944
R9702 gnd.n4322 gnd.n4321 19.3944
R9703 gnd.n4322 gnd.n3410 19.3944
R9704 gnd.n4342 gnd.n3410 19.3944
R9705 gnd.n4342 gnd.n3403 19.3944
R9706 gnd.n4352 gnd.n3403 19.3944
R9707 gnd.n4353 gnd.n4352 19.3944
R9708 gnd.n4353 gnd.n3385 19.3944
R9709 gnd.n4373 gnd.n3385 19.3944
R9710 gnd.n4373 gnd.n3377 19.3944
R9711 gnd.n4639 gnd.n3377 19.3944
R9712 gnd.n4640 gnd.n4639 19.3944
R9713 gnd.n4640 gnd.n3359 19.3944
R9714 gnd.n4659 gnd.n3359 19.3944
R9715 gnd.n4659 gnd.n3360 19.3944
R9716 gnd.n4053 gnd.n4052 19.3944
R9717 gnd.n4052 gnd.n3785 19.3944
R9718 gnd.n3808 gnd.n3785 19.3944
R9719 gnd.n3811 gnd.n3808 19.3944
R9720 gnd.n3811 gnd.n3804 19.3944
R9721 gnd.n3815 gnd.n3804 19.3944
R9722 gnd.n3818 gnd.n3815 19.3944
R9723 gnd.n3821 gnd.n3818 19.3944
R9724 gnd.n3821 gnd.n3802 19.3944
R9725 gnd.n3825 gnd.n3802 19.3944
R9726 gnd.n3828 gnd.n3825 19.3944
R9727 gnd.n3831 gnd.n3828 19.3944
R9728 gnd.n3831 gnd.n3800 19.3944
R9729 gnd.n3835 gnd.n3800 19.3944
R9730 gnd.n4058 gnd.n4057 19.3944
R9731 gnd.n4057 gnd.n3761 19.3944
R9732 gnd.n4083 gnd.n3761 19.3944
R9733 gnd.n4083 gnd.n3759 19.3944
R9734 gnd.n4089 gnd.n3759 19.3944
R9735 gnd.n4089 gnd.n4088 19.3944
R9736 gnd.n4088 gnd.n3733 19.3944
R9737 gnd.n4113 gnd.n3733 19.3944
R9738 gnd.n4113 gnd.n3731 19.3944
R9739 gnd.n4125 gnd.n3731 19.3944
R9740 gnd.n4125 gnd.n4124 19.3944
R9741 gnd.n4124 gnd.n4123 19.3944
R9742 gnd.n4123 gnd.n4121 19.3944
R9743 gnd.n4121 gnd.n3703 19.3944
R9744 gnd.n3703 gnd.n3701 19.3944
R9745 gnd.n4172 gnd.n3701 19.3944
R9746 gnd.n4172 gnd.n3699 19.3944
R9747 gnd.n4176 gnd.n3699 19.3944
R9748 gnd.n4176 gnd.n3519 19.3944
R9749 gnd.n4208 gnd.n3519 19.3944
R9750 gnd.n4208 gnd.n3517 19.3944
R9751 gnd.n4214 gnd.n3517 19.3944
R9752 gnd.n4214 gnd.n4213 19.3944
R9753 gnd.n4213 gnd.n3495 19.3944
R9754 gnd.n4239 gnd.n3495 19.3944
R9755 gnd.n4239 gnd.n3493 19.3944
R9756 gnd.n4245 gnd.n3493 19.3944
R9757 gnd.n4245 gnd.n4244 19.3944
R9758 gnd.n4244 gnd.n3469 19.3944
R9759 gnd.n4270 gnd.n3469 19.3944
R9760 gnd.n4270 gnd.n3467 19.3944
R9761 gnd.n4276 gnd.n3467 19.3944
R9762 gnd.n4276 gnd.n4275 19.3944
R9763 gnd.n4275 gnd.n3444 19.3944
R9764 gnd.n4301 gnd.n3444 19.3944
R9765 gnd.n4301 gnd.n3442 19.3944
R9766 gnd.n4307 gnd.n3442 19.3944
R9767 gnd.n4307 gnd.n4306 19.3944
R9768 gnd.n4306 gnd.n3419 19.3944
R9769 gnd.n4332 gnd.n3419 19.3944
R9770 gnd.n4332 gnd.n3417 19.3944
R9771 gnd.n4338 gnd.n3417 19.3944
R9772 gnd.n4338 gnd.n4337 19.3944
R9773 gnd.n4337 gnd.n3393 19.3944
R9774 gnd.n4363 gnd.n3393 19.3944
R9775 gnd.n4363 gnd.n3391 19.3944
R9776 gnd.n4369 gnd.n3391 19.3944
R9777 gnd.n4369 gnd.n4368 19.3944
R9778 gnd.n4368 gnd.n3368 19.3944
R9779 gnd.n4649 gnd.n3368 19.3944
R9780 gnd.n4649 gnd.n3366 19.3944
R9781 gnd.n4655 gnd.n3366 19.3944
R9782 gnd.n4655 gnd.n4654 19.3944
R9783 gnd.n4753 gnd.n4752 19.3944
R9784 gnd.n4752 gnd.n2014 19.3944
R9785 gnd.n4748 gnd.n2014 19.3944
R9786 gnd.n4748 gnd.n4745 19.3944
R9787 gnd.n4745 gnd.n4742 19.3944
R9788 gnd.n4742 gnd.n4741 19.3944
R9789 gnd.n4741 gnd.n4738 19.3944
R9790 gnd.n4738 gnd.n4737 19.3944
R9791 gnd.n4737 gnd.n4734 19.3944
R9792 gnd.n4734 gnd.n4733 19.3944
R9793 gnd.n4733 gnd.n4730 19.3944
R9794 gnd.n4730 gnd.n4729 19.3944
R9795 gnd.n4729 gnd.n4726 19.3944
R9796 gnd.n4726 gnd.n4725 19.3944
R9797 gnd.n3973 gnd.n3872 19.3944
R9798 gnd.n3973 gnd.n3863 19.3944
R9799 gnd.n3986 gnd.n3863 19.3944
R9800 gnd.n3986 gnd.n3861 19.3944
R9801 gnd.n3990 gnd.n3861 19.3944
R9802 gnd.n3990 gnd.n3851 19.3944
R9803 gnd.n4002 gnd.n3851 19.3944
R9804 gnd.n4002 gnd.n3849 19.3944
R9805 gnd.n4036 gnd.n3849 19.3944
R9806 gnd.n4036 gnd.n4035 19.3944
R9807 gnd.n4035 gnd.n4034 19.3944
R9808 gnd.n4034 gnd.n4033 19.3944
R9809 gnd.n4033 gnd.n4030 19.3944
R9810 gnd.n4030 gnd.n4029 19.3944
R9811 gnd.n4029 gnd.n4028 19.3944
R9812 gnd.n4028 gnd.n4026 19.3944
R9813 gnd.n4026 gnd.n4025 19.3944
R9814 gnd.n4025 gnd.n4022 19.3944
R9815 gnd.n4022 gnd.n4021 19.3944
R9816 gnd.n4021 gnd.n4020 19.3944
R9817 gnd.n4020 gnd.n4018 19.3944
R9818 gnd.n4018 gnd.n3716 19.3944
R9819 gnd.n4139 gnd.n3716 19.3944
R9820 gnd.n4139 gnd.n3714 19.3944
R9821 gnd.n4145 gnd.n3714 19.3944
R9822 gnd.n4145 gnd.n4144 19.3944
R9823 gnd.n4144 gnd.n3679 19.3944
R9824 gnd.n4187 gnd.n3679 19.3944
R9825 gnd.n4187 gnd.n3680 19.3944
R9826 gnd.n3696 gnd.n3695 19.3944
R9827 gnd.n4192 gnd.n4191 19.3944
R9828 gnd.n3615 gnd.n3534 19.3944
R9829 gnd.n3610 gnd.n3609 19.3944
R9830 gnd.n3609 gnd.n3607 19.3944
R9831 gnd.n3607 gnd.n3606 19.3944
R9832 gnd.n3606 gnd.n3603 19.3944
R9833 gnd.n3603 gnd.n3602 19.3944
R9834 gnd.n3602 gnd.n3601 19.3944
R9835 gnd.n3601 gnd.n3599 19.3944
R9836 gnd.n3599 gnd.n3598 19.3944
R9837 gnd.n3598 gnd.n3595 19.3944
R9838 gnd.n3595 gnd.n3594 19.3944
R9839 gnd.n3594 gnd.n3593 19.3944
R9840 gnd.n3593 gnd.n3591 19.3944
R9841 gnd.n3591 gnd.n3590 19.3944
R9842 gnd.n3590 gnd.n3585 19.3944
R9843 gnd.n3585 gnd.n3584 19.3944
R9844 gnd.n3584 gnd.n3583 19.3944
R9845 gnd.n3583 gnd.n3581 19.3944
R9846 gnd.n3581 gnd.n3580 19.3944
R9847 gnd.n3580 gnd.n3577 19.3944
R9848 gnd.n3577 gnd.n3576 19.3944
R9849 gnd.n3576 gnd.n3575 19.3944
R9850 gnd.n3575 gnd.n3573 19.3944
R9851 gnd.n3573 gnd.n3572 19.3944
R9852 gnd.n3572 gnd.n3569 19.3944
R9853 gnd.n3569 gnd.n3568 19.3944
R9854 gnd.n3568 gnd.n3567 19.3944
R9855 gnd.n3567 gnd.n3565 19.3944
R9856 gnd.n3565 gnd.n3564 19.3944
R9857 gnd.n3564 gnd.n2061 19.3944
R9858 gnd.n3978 gnd.n3868 19.3944
R9859 gnd.n3978 gnd.n3866 19.3944
R9860 gnd.n3982 gnd.n3866 19.3944
R9861 gnd.n3982 gnd.n3857 19.3944
R9862 gnd.n3994 gnd.n3857 19.3944
R9863 gnd.n3994 gnd.n3855 19.3944
R9864 gnd.n3998 gnd.n3855 19.3944
R9865 gnd.n3998 gnd.n3844 19.3944
R9866 gnd.n4040 gnd.n3844 19.3944
R9867 gnd.n4040 gnd.n3798 19.3944
R9868 gnd.n4046 gnd.n3798 19.3944
R9869 gnd.n4046 gnd.n4045 19.3944
R9870 gnd.n4045 gnd.n3776 19.3944
R9871 gnd.n4067 gnd.n3776 19.3944
R9872 gnd.n4067 gnd.n3769 19.3944
R9873 gnd.n4078 gnd.n3769 19.3944
R9874 gnd.n4078 gnd.n4077 19.3944
R9875 gnd.n4077 gnd.n3750 19.3944
R9876 gnd.n4098 gnd.n3750 19.3944
R9877 gnd.n4098 gnd.n3740 19.3944
R9878 gnd.n4108 gnd.n3740 19.3944
R9879 gnd.n4108 gnd.n3721 19.3944
R9880 gnd.n4135 gnd.n3721 19.3944
R9881 gnd.n4135 gnd.n4134 19.3944
R9882 gnd.n4134 gnd.n3709 19.3944
R9883 gnd.n4151 gnd.n3709 19.3944
R9884 gnd.n4151 gnd.n3687 19.3944
R9885 gnd.n4183 gnd.n3687 19.3944
R9886 gnd.n4183 gnd.n4182 19.3944
R9887 gnd.n4182 gnd.n4181 19.3944
R9888 gnd.n4181 gnd.n3693 19.3944
R9889 gnd.n3693 gnd.n3526 19.3944
R9890 gnd.n4203 gnd.n3526 19.3944
R9891 gnd.n4203 gnd.n4202 19.3944
R9892 gnd.n4202 gnd.n3510 19.3944
R9893 gnd.n4223 gnd.n3510 19.3944
R9894 gnd.n4223 gnd.n3503 19.3944
R9895 gnd.n4234 gnd.n3503 19.3944
R9896 gnd.n4234 gnd.n4233 19.3944
R9897 gnd.n4233 gnd.n3485 19.3944
R9898 gnd.n4254 gnd.n3485 19.3944
R9899 gnd.n4254 gnd.n3477 19.3944
R9900 gnd.n4265 gnd.n3477 19.3944
R9901 gnd.n4265 gnd.n4264 19.3944
R9902 gnd.n4264 gnd.n3458 19.3944
R9903 gnd.n4285 gnd.n3458 19.3944
R9904 gnd.n4285 gnd.n3451 19.3944
R9905 gnd.n4296 gnd.n3451 19.3944
R9906 gnd.n4296 gnd.n4295 19.3944
R9907 gnd.n4295 gnd.n3434 19.3944
R9908 gnd.n4316 gnd.n3434 19.3944
R9909 gnd.n4316 gnd.n3427 19.3944
R9910 gnd.n4327 gnd.n3427 19.3944
R9911 gnd.n4327 gnd.n4326 19.3944
R9912 gnd.n4326 gnd.n3408 19.3944
R9913 gnd.n4347 gnd.n3408 19.3944
R9914 gnd.n4347 gnd.n3401 19.3944
R9915 gnd.n4358 gnd.n3401 19.3944
R9916 gnd.n4358 gnd.n4357 19.3944
R9917 gnd.n4357 gnd.n3383 19.3944
R9918 gnd.n4634 gnd.n3383 19.3944
R9919 gnd.n4634 gnd.n3375 19.3944
R9920 gnd.n4644 gnd.n3375 19.3944
R9921 gnd.n4644 gnd.n3357 19.3944
R9922 gnd.n4662 gnd.n3357 19.3944
R9923 gnd.n6972 gnd.n565 19.3944
R9924 gnd.n6968 gnd.n565 19.3944
R9925 gnd.n6968 gnd.n6967 19.3944
R9926 gnd.n6967 gnd.n6966 19.3944
R9927 gnd.n6966 gnd.n570 19.3944
R9928 gnd.n6962 gnd.n570 19.3944
R9929 gnd.n6962 gnd.n6961 19.3944
R9930 gnd.n6961 gnd.n6960 19.3944
R9931 gnd.n6960 gnd.n574 19.3944
R9932 gnd.n6956 gnd.n574 19.3944
R9933 gnd.n6956 gnd.n6955 19.3944
R9934 gnd.n6955 gnd.n6954 19.3944
R9935 gnd.n6954 gnd.n578 19.3944
R9936 gnd.n6950 gnd.n578 19.3944
R9937 gnd.n6950 gnd.n6949 19.3944
R9938 gnd.n6949 gnd.n6948 19.3944
R9939 gnd.n6948 gnd.n582 19.3944
R9940 gnd.n6944 gnd.n582 19.3944
R9941 gnd.n6944 gnd.n6943 19.3944
R9942 gnd.n6943 gnd.n6942 19.3944
R9943 gnd.n6942 gnd.n384 19.3944
R9944 gnd.n7161 gnd.n384 19.3944
R9945 gnd.n7162 gnd.n7161 19.3944
R9946 gnd.n7162 gnd.n381 19.3944
R9947 gnd.n7167 gnd.n381 19.3944
R9948 gnd.n7167 gnd.n382 19.3944
R9949 gnd.n382 gnd.n352 19.3944
R9950 gnd.n7209 gnd.n352 19.3944
R9951 gnd.n7209 gnd.n353 19.3944
R9952 gnd.n7205 gnd.n353 19.3944
R9953 gnd.n7205 gnd.n7204 19.3944
R9954 gnd.n7204 gnd.n76 19.3944
R9955 gnd.n7624 gnd.n76 19.3944
R9956 gnd.n7624 gnd.n7623 19.3944
R9957 gnd.n7623 gnd.n7622 19.3944
R9958 gnd.n7622 gnd.n81 19.3944
R9959 gnd.n7618 gnd.n81 19.3944
R9960 gnd.n7618 gnd.n7617 19.3944
R9961 gnd.n7617 gnd.n7616 19.3944
R9962 gnd.n7616 gnd.n86 19.3944
R9963 gnd.n7612 gnd.n86 19.3944
R9964 gnd.n7612 gnd.n7611 19.3944
R9965 gnd.n7611 gnd.n7610 19.3944
R9966 gnd.n7610 gnd.n91 19.3944
R9967 gnd.n7606 gnd.n91 19.3944
R9968 gnd.n7606 gnd.n7605 19.3944
R9969 gnd.n7605 gnd.n7604 19.3944
R9970 gnd.n7604 gnd.n96 19.3944
R9971 gnd.n7600 gnd.n96 19.3944
R9972 gnd.n7600 gnd.n7599 19.3944
R9973 gnd.n7599 gnd.n7598 19.3944
R9974 gnd.n7598 gnd.n101 19.3944
R9975 gnd.n7594 gnd.n101 19.3944
R9976 gnd.n7594 gnd.n7593 19.3944
R9977 gnd.n7593 gnd.n7592 19.3944
R9978 gnd.n7592 gnd.n106 19.3944
R9979 gnd.n7588 gnd.n106 19.3944
R9980 gnd.n7588 gnd.n7587 19.3944
R9981 gnd.n7587 gnd.n7586 19.3944
R9982 gnd.n7586 gnd.n111 19.3944
R9983 gnd.n7582 gnd.n111 19.3944
R9984 gnd.n7582 gnd.n7581 19.3944
R9985 gnd.n7581 gnd.n7580 19.3944
R9986 gnd.n7580 gnd.n116 19.3944
R9987 gnd.n7474 gnd.n7473 19.3944
R9988 gnd.n7473 gnd.n7472 19.3944
R9989 gnd.n7472 gnd.n7421 19.3944
R9990 gnd.n7468 gnd.n7421 19.3944
R9991 gnd.n7468 gnd.n7467 19.3944
R9992 gnd.n7467 gnd.n7466 19.3944
R9993 gnd.n7466 gnd.n7429 19.3944
R9994 gnd.n7462 gnd.n7429 19.3944
R9995 gnd.n7462 gnd.n7461 19.3944
R9996 gnd.n7461 gnd.n7460 19.3944
R9997 gnd.n7460 gnd.n7437 19.3944
R9998 gnd.n7456 gnd.n7437 19.3944
R9999 gnd.n7456 gnd.n7455 19.3944
R10000 gnd.n7455 gnd.n7454 19.3944
R10001 gnd.n7454 gnd.n7445 19.3944
R10002 gnd.n7450 gnd.n7445 19.3944
R10003 gnd.n6623 gnd.n6622 19.3944
R10004 gnd.n6754 gnd.n6623 19.3944
R10005 gnd.n6754 gnd.n6753 19.3944
R10006 gnd.n6753 gnd.n6628 19.3944
R10007 gnd.n6746 gnd.n6628 19.3944
R10008 gnd.n6746 gnd.n6745 19.3944
R10009 gnd.n6745 gnd.n6638 19.3944
R10010 gnd.n6738 gnd.n6638 19.3944
R10011 gnd.n6738 gnd.n6737 19.3944
R10012 gnd.n6737 gnd.n6648 19.3944
R10013 gnd.n6730 gnd.n6648 19.3944
R10014 gnd.n6730 gnd.n6729 19.3944
R10015 gnd.n6729 gnd.n6658 19.3944
R10016 gnd.n6722 gnd.n6658 19.3944
R10017 gnd.n6722 gnd.n6721 19.3944
R10018 gnd.n6721 gnd.n6668 19.3944
R10019 gnd.n7057 gnd.n478 19.3944
R10020 gnd.n7057 gnd.n476 19.3944
R10021 gnd.n7061 gnd.n476 19.3944
R10022 gnd.n7061 gnd.n460 19.3944
R10023 gnd.n7073 gnd.n460 19.3944
R10024 gnd.n7073 gnd.n458 19.3944
R10025 gnd.n7077 gnd.n458 19.3944
R10026 gnd.n7077 gnd.n444 19.3944
R10027 gnd.n7089 gnd.n444 19.3944
R10028 gnd.n7089 gnd.n442 19.3944
R10029 gnd.n7093 gnd.n442 19.3944
R10030 gnd.n7093 gnd.n426 19.3944
R10031 gnd.n7105 gnd.n426 19.3944
R10032 gnd.n7105 gnd.n424 19.3944
R10033 gnd.n7109 gnd.n424 19.3944
R10034 gnd.n7109 gnd.n410 19.3944
R10035 gnd.n7121 gnd.n410 19.3944
R10036 gnd.n7121 gnd.n407 19.3944
R10037 gnd.n7128 gnd.n407 19.3944
R10038 gnd.n7128 gnd.n408 19.3944
R10039 gnd.n7124 gnd.n408 19.3944
R10040 gnd.n7124 gnd.n375 19.3944
R10041 gnd.n7179 gnd.n375 19.3944
R10042 gnd.n7179 gnd.n376 19.3944
R10043 gnd.n7175 gnd.n376 19.3944
R10044 gnd.n7175 gnd.n7174 19.3944
R10045 gnd.n7174 gnd.n7173 19.3944
R10046 gnd.n7173 gnd.n314 19.3944
R10047 gnd.n7318 gnd.n314 19.3944
R10048 gnd.n7318 gnd.n315 19.3944
R10049 gnd.n7314 gnd.n315 19.3944
R10050 gnd.n7314 gnd.n7313 19.3944
R10051 gnd.n7313 gnd.n7312 19.3944
R10052 gnd.n7312 gnd.n321 19.3944
R10053 gnd.n7308 gnd.n321 19.3944
R10054 gnd.n7308 gnd.n7307 19.3944
R10055 gnd.n7307 gnd.n293 19.3944
R10056 gnd.n7331 gnd.n293 19.3944
R10057 gnd.n7331 gnd.n291 19.3944
R10058 gnd.n7335 gnd.n291 19.3944
R10059 gnd.n7335 gnd.n277 19.3944
R10060 gnd.n7347 gnd.n277 19.3944
R10061 gnd.n7347 gnd.n275 19.3944
R10062 gnd.n7351 gnd.n275 19.3944
R10063 gnd.n7351 gnd.n263 19.3944
R10064 gnd.n7363 gnd.n263 19.3944
R10065 gnd.n7363 gnd.n261 19.3944
R10066 gnd.n7367 gnd.n261 19.3944
R10067 gnd.n7367 gnd.n247 19.3944
R10068 gnd.n7379 gnd.n247 19.3944
R10069 gnd.n7379 gnd.n245 19.3944
R10070 gnd.n7383 gnd.n245 19.3944
R10071 gnd.n7383 gnd.n232 19.3944
R10072 gnd.n7395 gnd.n232 19.3944
R10073 gnd.n7395 gnd.n230 19.3944
R10074 gnd.n7399 gnd.n230 19.3944
R10075 gnd.n7399 gnd.n217 19.3944
R10076 gnd.n7411 gnd.n217 19.3944
R10077 gnd.n7411 gnd.n214 19.3944
R10078 gnd.n7483 gnd.n214 19.3944
R10079 gnd.n7483 gnd.n215 19.3944
R10080 gnd.n7479 gnd.n215 19.3944
R10081 gnd.n7479 gnd.n7478 19.3944
R10082 gnd.n7478 gnd.n7477 19.3944
R10083 gnd.n5673 gnd.n5573 19.3944
R10084 gnd.n5673 gnd.n5672 19.3944
R10085 gnd.n5672 gnd.n5579 19.3944
R10086 gnd.n5665 gnd.n5579 19.3944
R10087 gnd.n5665 gnd.n5664 19.3944
R10088 gnd.n5664 gnd.n5591 19.3944
R10089 gnd.n5657 gnd.n5591 19.3944
R10090 gnd.n5657 gnd.n5656 19.3944
R10091 gnd.n5656 gnd.n5604 19.3944
R10092 gnd.n5649 gnd.n5604 19.3944
R10093 gnd.n5649 gnd.n5648 19.3944
R10094 gnd.n5648 gnd.n5614 19.3944
R10095 gnd.n5641 gnd.n5614 19.3944
R10096 gnd.n5641 gnd.n5640 19.3944
R10097 gnd.n5640 gnd.n5630 19.3944
R10098 gnd.n5630 gnd.n1347 19.3944
R10099 gnd.n5435 gnd.n1800 19.3944
R10100 gnd.n5435 gnd.n5434 19.3944
R10101 gnd.n5434 gnd.n5433 19.3944
R10102 gnd.n5433 gnd.n1804 19.3944
R10103 gnd.n5259 gnd.n1804 19.3944
R10104 gnd.n5259 gnd.n5257 19.3944
R10105 gnd.n5273 gnd.n5257 19.3944
R10106 gnd.n5273 gnd.n5272 19.3944
R10107 gnd.n5272 gnd.n5271 19.3944
R10108 gnd.n5271 gnd.n5268 19.3944
R10109 gnd.n5268 gnd.n5267 19.3944
R10110 gnd.n5267 gnd.n1848 19.3944
R10111 gnd.n5299 gnd.n1848 19.3944
R10112 gnd.n5299 gnd.n1846 19.3944
R10113 gnd.n5313 gnd.n1846 19.3944
R10114 gnd.n5313 gnd.n5312 19.3944
R10115 gnd.n5312 gnd.n5311 19.3944
R10116 gnd.n5311 gnd.n5308 19.3944
R10117 gnd.n5308 gnd.n5307 19.3944
R10118 gnd.n5307 gnd.n1838 19.3944
R10119 gnd.n5338 gnd.n1838 19.3944
R10120 gnd.n5338 gnd.n1836 19.3944
R10121 gnd.n5370 gnd.n1836 19.3944
R10122 gnd.n5370 gnd.n5369 19.3944
R10123 gnd.n5369 gnd.n5368 19.3944
R10124 gnd.n5368 gnd.n5344 19.3944
R10125 gnd.n5364 gnd.n5344 19.3944
R10126 gnd.n5364 gnd.n5363 19.3944
R10127 gnd.n5363 gnd.n5362 19.3944
R10128 gnd.n5362 gnd.n5350 19.3944
R10129 gnd.n5357 gnd.n5350 19.3944
R10130 gnd.n5357 gnd.n5356 19.3944
R10131 gnd.n5356 gnd.n1316 19.3944
R10132 gnd.n5811 gnd.n1316 19.3944
R10133 gnd.n5811 gnd.n1314 19.3944
R10134 gnd.n5815 gnd.n1314 19.3944
R10135 gnd.n5815 gnd.n1302 19.3944
R10136 gnd.n5827 gnd.n1302 19.3944
R10137 gnd.n5827 gnd.n1300 19.3944
R10138 gnd.n5833 gnd.n1300 19.3944
R10139 gnd.n5833 gnd.n5832 19.3944
R10140 gnd.n5832 gnd.n1260 19.3944
R10141 gnd.n5985 gnd.n1260 19.3944
R10142 gnd.n5985 gnd.n1258 19.3944
R10143 gnd.n5989 gnd.n1258 19.3944
R10144 gnd.n5989 gnd.n1245 19.3944
R10145 gnd.n6001 gnd.n1245 19.3944
R10146 gnd.n6001 gnd.n1243 19.3944
R10147 gnd.n6005 gnd.n1243 19.3944
R10148 gnd.n6005 gnd.n1229 19.3944
R10149 gnd.n6017 gnd.n1229 19.3944
R10150 gnd.n6017 gnd.n1227 19.3944
R10151 gnd.n6021 gnd.n1227 19.3944
R10152 gnd.n6021 gnd.n1214 19.3944
R10153 gnd.n6032 gnd.n1214 19.3944
R10154 gnd.n6032 gnd.n1212 19.3944
R10155 gnd.n6038 gnd.n1212 19.3944
R10156 gnd.n6038 gnd.n6037 19.3944
R10157 gnd.n6037 gnd.n1107 19.3944
R10158 gnd.n6127 gnd.n1107 19.3944
R10159 gnd.n6127 gnd.n1105 19.3944
R10160 gnd.n6131 gnd.n1105 19.3944
R10161 gnd.n6131 gnd.n1091 19.3944
R10162 gnd.n6143 gnd.n1091 19.3944
R10163 gnd.n6143 gnd.n1089 19.3944
R10164 gnd.n6147 gnd.n1089 19.3944
R10165 gnd.n6147 gnd.n1076 19.3944
R10166 gnd.n6159 gnd.n1076 19.3944
R10167 gnd.n6159 gnd.n1074 19.3944
R10168 gnd.n6163 gnd.n1074 19.3944
R10169 gnd.n6163 gnd.n1063 19.3944
R10170 gnd.n6175 gnd.n1063 19.3944
R10171 gnd.n6175 gnd.n1061 19.3944
R10172 gnd.n6181 gnd.n1061 19.3944
R10173 gnd.n6181 gnd.n6180 19.3944
R10174 gnd.n6180 gnd.n1020 19.3944
R10175 gnd.n6432 gnd.n1020 19.3944
R10176 gnd.n6432 gnd.n1018 19.3944
R10177 gnd.n6436 gnd.n1018 19.3944
R10178 gnd.n6436 gnd.n1004 19.3944
R10179 gnd.n6448 gnd.n1004 19.3944
R10180 gnd.n6448 gnd.n1002 19.3944
R10181 gnd.n6452 gnd.n1002 19.3944
R10182 gnd.n6452 gnd.n988 19.3944
R10183 gnd.n6464 gnd.n988 19.3944
R10184 gnd.n6464 gnd.n986 19.3944
R10185 gnd.n6468 gnd.n986 19.3944
R10186 gnd.n6468 gnd.n974 19.3944
R10187 gnd.n6480 gnd.n974 19.3944
R10188 gnd.n6480 gnd.n972 19.3944
R10189 gnd.n6484 gnd.n972 19.3944
R10190 gnd.n6484 gnd.n959 19.3944
R10191 gnd.n6496 gnd.n959 19.3944
R10192 gnd.n6496 gnd.n957 19.3944
R10193 gnd.n6500 gnd.n957 19.3944
R10194 gnd.n6500 gnd.n943 19.3944
R10195 gnd.n6512 gnd.n943 19.3944
R10196 gnd.n6512 gnd.n941 19.3944
R10197 gnd.n6516 gnd.n941 19.3944
R10198 gnd.n6516 gnd.n926 19.3944
R10199 gnd.n6534 gnd.n926 19.3944
R10200 gnd.n6534 gnd.n924 19.3944
R10201 gnd.n6540 gnd.n924 19.3944
R10202 gnd.n6540 gnd.n6539 19.3944
R10203 gnd.n6539 gnd.n886 19.3944
R10204 gnd.n6592 gnd.n886 19.3944
R10205 gnd.n6592 gnd.n884 19.3944
R10206 gnd.n6598 gnd.n884 19.3944
R10207 gnd.n6598 gnd.n6597 19.3944
R10208 gnd.n6597 gnd.n659 19.3944
R10209 gnd.n6783 gnd.n659 19.3944
R10210 gnd.n6783 gnd.n657 19.3944
R10211 gnd.n6787 gnd.n657 19.3944
R10212 gnd.n6787 gnd.n644 19.3944
R10213 gnd.n6800 gnd.n644 19.3944
R10214 gnd.n6800 gnd.n642 19.3944
R10215 gnd.n6806 gnd.n642 19.3944
R10216 gnd.n6806 gnd.n6805 19.3944
R10217 gnd.n6805 gnd.n614 19.3944
R10218 gnd.n6819 gnd.n614 19.3944
R10219 gnd.n6819 gnd.n612 19.3944
R10220 gnd.n6823 gnd.n612 19.3944
R10221 gnd.n6823 gnd.n610 19.3944
R10222 gnd.n6827 gnd.n610 19.3944
R10223 gnd.n6827 gnd.n608 19.3944
R10224 gnd.n6831 gnd.n608 19.3944
R10225 gnd.n6831 gnd.n606 19.3944
R10226 gnd.n6835 gnd.n606 19.3944
R10227 gnd.n6835 gnd.n604 19.3944
R10228 gnd.n6839 gnd.n604 19.3944
R10229 gnd.n6839 gnd.n602 19.3944
R10230 gnd.n6869 gnd.n602 19.3944
R10231 gnd.n6869 gnd.n600 19.3944
R10232 gnd.n6883 gnd.n600 19.3944
R10233 gnd.n6883 gnd.n6882 19.3944
R10234 gnd.n6882 gnd.n6881 19.3944
R10235 gnd.n6881 gnd.n6878 19.3944
R10236 gnd.n6878 gnd.n6877 19.3944
R10237 gnd.n6877 gnd.n592 19.3944
R10238 gnd.n6908 gnd.n592 19.3944
R10239 gnd.n6908 gnd.n590 19.3944
R10240 gnd.n6914 gnd.n590 19.3944
R10241 gnd.n6914 gnd.n6913 19.3944
R10242 gnd.n6913 gnd.n392 19.3944
R10243 gnd.n7141 gnd.n392 19.3944
R10244 gnd.n7141 gnd.n390 19.3944
R10245 gnd.n7156 gnd.n390 19.3944
R10246 gnd.n7156 gnd.n7155 19.3944
R10247 gnd.n7155 gnd.n7154 19.3944
R10248 gnd.n7154 gnd.n7151 19.3944
R10249 gnd.n7151 gnd.n7150 19.3944
R10250 gnd.n7150 gnd.n346 19.3944
R10251 gnd.n7215 gnd.n346 19.3944
R10252 gnd.n7216 gnd.n7215 19.3944
R10253 gnd.n2825 gnd.n2499 19.3944
R10254 gnd.n2825 gnd.n2500 19.3944
R10255 gnd.n2821 gnd.n2500 19.3944
R10256 gnd.n2821 gnd.n2503 19.3944
R10257 gnd.n2815 gnd.n2503 19.3944
R10258 gnd.n2815 gnd.n2814 19.3944
R10259 gnd.n2814 gnd.n2813 19.3944
R10260 gnd.n2813 gnd.n2510 19.3944
R10261 gnd.n2807 gnd.n2510 19.3944
R10262 gnd.n2807 gnd.n2806 19.3944
R10263 gnd.n2806 gnd.n2805 19.3944
R10264 gnd.n2805 gnd.n2518 19.3944
R10265 gnd.n2799 gnd.n2518 19.3944
R10266 gnd.n2799 gnd.n2798 19.3944
R10267 gnd.n2798 gnd.n2797 19.3944
R10268 gnd.n2797 gnd.n2526 19.3944
R10269 gnd.n2791 gnd.n2526 19.3944
R10270 gnd.n2791 gnd.n2790 19.3944
R10271 gnd.n2790 gnd.n2789 19.3944
R10272 gnd.n2789 gnd.n2534 19.3944
R10273 gnd.n2783 gnd.n2534 19.3944
R10274 gnd.n2783 gnd.n2782 19.3944
R10275 gnd.n2782 gnd.n2781 19.3944
R10276 gnd.n2781 gnd.n2542 19.3944
R10277 gnd.n2775 gnd.n2542 19.3944
R10278 gnd.n2775 gnd.n2774 19.3944
R10279 gnd.n2774 gnd.n2773 19.3944
R10280 gnd.n2773 gnd.n2550 19.3944
R10281 gnd.n2767 gnd.n2550 19.3944
R10282 gnd.n2767 gnd.n2766 19.3944
R10283 gnd.n2766 gnd.n2765 19.3944
R10284 gnd.n2765 gnd.n2558 19.3944
R10285 gnd.n2759 gnd.n2558 19.3944
R10286 gnd.n2759 gnd.n2758 19.3944
R10287 gnd.n2758 gnd.n2757 19.3944
R10288 gnd.n2757 gnd.n2566 19.3944
R10289 gnd.n2751 gnd.n2566 19.3944
R10290 gnd.n2751 gnd.n2750 19.3944
R10291 gnd.n2750 gnd.n2749 19.3944
R10292 gnd.n2749 gnd.n2574 19.3944
R10293 gnd.n2743 gnd.n2574 19.3944
R10294 gnd.n2743 gnd.n2742 19.3944
R10295 gnd.n2742 gnd.n2741 19.3944
R10296 gnd.n2741 gnd.n2582 19.3944
R10297 gnd.n2735 gnd.n2582 19.3944
R10298 gnd.n2735 gnd.n2734 19.3944
R10299 gnd.n2734 gnd.n2733 19.3944
R10300 gnd.n2733 gnd.n2590 19.3944
R10301 gnd.n2727 gnd.n2590 19.3944
R10302 gnd.n2727 gnd.n2726 19.3944
R10303 gnd.n2726 gnd.n2725 19.3944
R10304 gnd.n2725 gnd.n2598 19.3944
R10305 gnd.n2719 gnd.n2598 19.3944
R10306 gnd.n2719 gnd.n2718 19.3944
R10307 gnd.n2718 gnd.n2717 19.3944
R10308 gnd.n2717 gnd.n2606 19.3944
R10309 gnd.n2711 gnd.n2606 19.3944
R10310 gnd.n2711 gnd.n2710 19.3944
R10311 gnd.n2710 gnd.n2709 19.3944
R10312 gnd.n2709 gnd.n2614 19.3944
R10313 gnd.n2703 gnd.n2614 19.3944
R10314 gnd.n2703 gnd.n2702 19.3944
R10315 gnd.n2702 gnd.n2701 19.3944
R10316 gnd.n2701 gnd.n2622 19.3944
R10317 gnd.n2695 gnd.n2622 19.3944
R10318 gnd.n2695 gnd.n2694 19.3944
R10319 gnd.n2694 gnd.n2693 19.3944
R10320 gnd.n2693 gnd.n2630 19.3944
R10321 gnd.n2687 gnd.n2630 19.3944
R10322 gnd.n2687 gnd.n2686 19.3944
R10323 gnd.n2686 gnd.n2685 19.3944
R10324 gnd.n2685 gnd.n2638 19.3944
R10325 gnd.n2679 gnd.n2638 19.3944
R10326 gnd.n2679 gnd.n2678 19.3944
R10327 gnd.n2678 gnd.n2677 19.3944
R10328 gnd.n2677 gnd.n2646 19.3944
R10329 gnd.n2671 gnd.n2646 19.3944
R10330 gnd.n2671 gnd.n2670 19.3944
R10331 gnd.n2670 gnd.n2669 19.3944
R10332 gnd.n2669 gnd.n2654 19.3944
R10333 gnd.n2663 gnd.n2654 19.3944
R10334 gnd.n2663 gnd.n2662 19.3944
R10335 gnd.n2662 gnd.n344 19.3944
R10336 gnd.n7219 gnd.n344 19.3944
R10337 gnd.n3139 gnd.n2191 19.3944
R10338 gnd.n3135 gnd.n2191 19.3944
R10339 gnd.n3135 gnd.n2193 19.3944
R10340 gnd.n3129 gnd.n2193 19.3944
R10341 gnd.n3129 gnd.n3128 19.3944
R10342 gnd.n3128 gnd.n3127 19.3944
R10343 gnd.n3127 gnd.n2200 19.3944
R10344 gnd.n3121 gnd.n2200 19.3944
R10345 gnd.n3121 gnd.n3120 19.3944
R10346 gnd.n3120 gnd.n3119 19.3944
R10347 gnd.n3119 gnd.n2208 19.3944
R10348 gnd.n3113 gnd.n2208 19.3944
R10349 gnd.n3113 gnd.n3112 19.3944
R10350 gnd.n3112 gnd.n3111 19.3944
R10351 gnd.n3111 gnd.n2216 19.3944
R10352 gnd.n3105 gnd.n2216 19.3944
R10353 gnd.n3105 gnd.n3104 19.3944
R10354 gnd.n3104 gnd.n3103 19.3944
R10355 gnd.n3103 gnd.n2224 19.3944
R10356 gnd.n3097 gnd.n2224 19.3944
R10357 gnd.n3097 gnd.n3096 19.3944
R10358 gnd.n3096 gnd.n3095 19.3944
R10359 gnd.n3095 gnd.n2232 19.3944
R10360 gnd.n3089 gnd.n2232 19.3944
R10361 gnd.n3089 gnd.n3088 19.3944
R10362 gnd.n3088 gnd.n3087 19.3944
R10363 gnd.n3087 gnd.n2240 19.3944
R10364 gnd.n3081 gnd.n2240 19.3944
R10365 gnd.n3081 gnd.n3080 19.3944
R10366 gnd.n3080 gnd.n3079 19.3944
R10367 gnd.n3079 gnd.n2248 19.3944
R10368 gnd.n3073 gnd.n2248 19.3944
R10369 gnd.n3073 gnd.n3072 19.3944
R10370 gnd.n3072 gnd.n3071 19.3944
R10371 gnd.n3071 gnd.n2256 19.3944
R10372 gnd.n3065 gnd.n2256 19.3944
R10373 gnd.n3065 gnd.n3064 19.3944
R10374 gnd.n3064 gnd.n3063 19.3944
R10375 gnd.n3063 gnd.n2264 19.3944
R10376 gnd.n3057 gnd.n2264 19.3944
R10377 gnd.n3057 gnd.n3056 19.3944
R10378 gnd.n3056 gnd.n3055 19.3944
R10379 gnd.n3055 gnd.n2272 19.3944
R10380 gnd.n3049 gnd.n2272 19.3944
R10381 gnd.n3049 gnd.n3048 19.3944
R10382 gnd.n3048 gnd.n3047 19.3944
R10383 gnd.n3047 gnd.n2280 19.3944
R10384 gnd.n3041 gnd.n2280 19.3944
R10385 gnd.n3041 gnd.n3040 19.3944
R10386 gnd.n3040 gnd.n3039 19.3944
R10387 gnd.n3039 gnd.n2288 19.3944
R10388 gnd.n3033 gnd.n2288 19.3944
R10389 gnd.n3033 gnd.n3032 19.3944
R10390 gnd.n3032 gnd.n3031 19.3944
R10391 gnd.n3031 gnd.n2296 19.3944
R10392 gnd.n3025 gnd.n2296 19.3944
R10393 gnd.n3025 gnd.n3024 19.3944
R10394 gnd.n3024 gnd.n3023 19.3944
R10395 gnd.n3023 gnd.n2304 19.3944
R10396 gnd.n3017 gnd.n2304 19.3944
R10397 gnd.n3017 gnd.n3016 19.3944
R10398 gnd.n3016 gnd.n3015 19.3944
R10399 gnd.n3015 gnd.n2312 19.3944
R10400 gnd.n3009 gnd.n2312 19.3944
R10401 gnd.n3009 gnd.n3008 19.3944
R10402 gnd.n3008 gnd.n3007 19.3944
R10403 gnd.n3007 gnd.n2320 19.3944
R10404 gnd.n3001 gnd.n2320 19.3944
R10405 gnd.n3001 gnd.n3000 19.3944
R10406 gnd.n3000 gnd.n2999 19.3944
R10407 gnd.n2999 gnd.n2328 19.3944
R10408 gnd.n2993 gnd.n2328 19.3944
R10409 gnd.n2993 gnd.n2992 19.3944
R10410 gnd.n2992 gnd.n2991 19.3944
R10411 gnd.n2991 gnd.n2336 19.3944
R10412 gnd.n2985 gnd.n2336 19.3944
R10413 gnd.n2985 gnd.n2984 19.3944
R10414 gnd.n2984 gnd.n2983 19.3944
R10415 gnd.n2983 gnd.n2344 19.3944
R10416 gnd.n2977 gnd.n2344 19.3944
R10417 gnd.n2977 gnd.n2976 19.3944
R10418 gnd.n2976 gnd.n2975 19.3944
R10419 gnd.n2975 gnd.n2352 19.3944
R10420 gnd.n2969 gnd.n2352 19.3944
R10421 gnd.n2969 gnd.n2968 19.3944
R10422 gnd.n2968 gnd.n2967 19.3944
R10423 gnd.n2967 gnd.n2360 19.3944
R10424 gnd.n2961 gnd.n2360 19.3944
R10425 gnd.n2961 gnd.n2960 19.3944
R10426 gnd.n2960 gnd.n2959 19.3944
R10427 gnd.n2959 gnd.n2368 19.3944
R10428 gnd.n2953 gnd.n2368 19.3944
R10429 gnd.n2953 gnd.n2952 19.3944
R10430 gnd.n2952 gnd.n2951 19.3944
R10431 gnd.n2951 gnd.n2376 19.3944
R10432 gnd.n2945 gnd.n2376 19.3944
R10433 gnd.n2945 gnd.n2944 19.3944
R10434 gnd.n2944 gnd.n2943 19.3944
R10435 gnd.n2943 gnd.n2384 19.3944
R10436 gnd.n2937 gnd.n2384 19.3944
R10437 gnd.n2937 gnd.n2936 19.3944
R10438 gnd.n2936 gnd.n2935 19.3944
R10439 gnd.n2935 gnd.n2392 19.3944
R10440 gnd.n2929 gnd.n2392 19.3944
R10441 gnd.n2929 gnd.n2928 19.3944
R10442 gnd.n2928 gnd.n2927 19.3944
R10443 gnd.n2927 gnd.n2400 19.3944
R10444 gnd.n2921 gnd.n2400 19.3944
R10445 gnd.n2921 gnd.n2920 19.3944
R10446 gnd.n2920 gnd.n2919 19.3944
R10447 gnd.n2919 gnd.n2408 19.3944
R10448 gnd.n2913 gnd.n2408 19.3944
R10449 gnd.n2913 gnd.n2912 19.3944
R10450 gnd.n2912 gnd.n2911 19.3944
R10451 gnd.n2911 gnd.n2416 19.3944
R10452 gnd.n2905 gnd.n2416 19.3944
R10453 gnd.n2905 gnd.n2904 19.3944
R10454 gnd.n2904 gnd.n2903 19.3944
R10455 gnd.n2903 gnd.n2424 19.3944
R10456 gnd.n2897 gnd.n2424 19.3944
R10457 gnd.n2897 gnd.n2896 19.3944
R10458 gnd.n2896 gnd.n2895 19.3944
R10459 gnd.n2895 gnd.n2432 19.3944
R10460 gnd.n2889 gnd.n2432 19.3944
R10461 gnd.n2889 gnd.n2888 19.3944
R10462 gnd.n2888 gnd.n2887 19.3944
R10463 gnd.n2887 gnd.n2440 19.3944
R10464 gnd.n2881 gnd.n2440 19.3944
R10465 gnd.n2881 gnd.n2880 19.3944
R10466 gnd.n2880 gnd.n2879 19.3944
R10467 gnd.n2879 gnd.n2448 19.3944
R10468 gnd.n2873 gnd.n2448 19.3944
R10469 gnd.n2873 gnd.n2872 19.3944
R10470 gnd.n2872 gnd.n2871 19.3944
R10471 gnd.n2871 gnd.n2456 19.3944
R10472 gnd.n2865 gnd.n2456 19.3944
R10473 gnd.n2865 gnd.n2864 19.3944
R10474 gnd.n2864 gnd.n2863 19.3944
R10475 gnd.n2863 gnd.n2464 19.3944
R10476 gnd.n2857 gnd.n2464 19.3944
R10477 gnd.n2857 gnd.n2856 19.3944
R10478 gnd.n2856 gnd.n2855 19.3944
R10479 gnd.n2855 gnd.n2472 19.3944
R10480 gnd.n2849 gnd.n2472 19.3944
R10481 gnd.n2849 gnd.n2848 19.3944
R10482 gnd.n2848 gnd.n2847 19.3944
R10483 gnd.n2847 gnd.n2480 19.3944
R10484 gnd.n2841 gnd.n2480 19.3944
R10485 gnd.n2841 gnd.n2840 19.3944
R10486 gnd.n2840 gnd.n2839 19.3944
R10487 gnd.n2839 gnd.n2488 19.3944
R10488 gnd.n2833 gnd.n2488 19.3944
R10489 gnd.n2833 gnd.n2832 19.3944
R10490 gnd.n2832 gnd.n2831 19.3944
R10491 gnd.n7049 gnd.n487 19.3944
R10492 gnd.n7044 gnd.n487 19.3944
R10493 gnd.n7044 gnd.n7043 19.3944
R10494 gnd.n7043 gnd.n7042 19.3944
R10495 gnd.n7042 gnd.n7039 19.3944
R10496 gnd.n7039 gnd.n7038 19.3944
R10497 gnd.n7038 gnd.n7035 19.3944
R10498 gnd.n7035 gnd.n7034 19.3944
R10499 gnd.n7034 gnd.n7031 19.3944
R10500 gnd.n7031 gnd.n7030 19.3944
R10501 gnd.n7030 gnd.n7027 19.3944
R10502 gnd.n7027 gnd.n7026 19.3944
R10503 gnd.n7026 gnd.n7023 19.3944
R10504 gnd.n7023 gnd.n7022 19.3944
R10505 gnd.n7022 gnd.n7019 19.3944
R10506 gnd.n7017 gnd.n7014 19.3944
R10507 gnd.n7014 gnd.n7013 19.3944
R10508 gnd.n7013 gnd.n7010 19.3944
R10509 gnd.n7010 gnd.n7009 19.3944
R10510 gnd.n7009 gnd.n7006 19.3944
R10511 gnd.n7006 gnd.n7005 19.3944
R10512 gnd.n7005 gnd.n7002 19.3944
R10513 gnd.n7002 gnd.n7001 19.3944
R10514 gnd.n7001 gnd.n6998 19.3944
R10515 gnd.n6998 gnd.n6997 19.3944
R10516 gnd.n6997 gnd.n6994 19.3944
R10517 gnd.n6994 gnd.n6993 19.3944
R10518 gnd.n6993 gnd.n6990 19.3944
R10519 gnd.n6990 gnd.n6989 19.3944
R10520 gnd.n6989 gnd.n6986 19.3944
R10521 gnd.n6986 gnd.n6985 19.3944
R10522 gnd.n6985 gnd.n6982 19.3944
R10523 gnd.n6982 gnd.n6981 19.3944
R10524 gnd.n6843 gnd.n563 19.3944
R10525 gnd.n6848 gnd.n6843 19.3944
R10526 gnd.n6849 gnd.n6848 19.3944
R10527 gnd.n6852 gnd.n6849 19.3944
R10528 gnd.n6852 gnd.n6841 19.3944
R10529 gnd.n6863 gnd.n6841 19.3944
R10530 gnd.n6863 gnd.n6862 19.3944
R10531 gnd.n6862 gnd.n6861 19.3944
R10532 gnd.n6861 gnd.n596 19.3944
R10533 gnd.n6888 gnd.n596 19.3944
R10534 gnd.n6889 gnd.n6888 19.3944
R10535 gnd.n6892 gnd.n6889 19.3944
R10536 gnd.n6892 gnd.n594 19.3944
R10537 gnd.n6902 gnd.n594 19.3944
R10538 gnd.n6902 gnd.n6901 19.3944
R10539 gnd.n6901 gnd.n6900 19.3944
R10540 gnd.n6900 gnd.n587 19.3944
R10541 gnd.n6919 gnd.n587 19.3944
R10542 gnd.n6919 gnd.n585 19.3944
R10543 gnd.n6936 gnd.n585 19.3944
R10544 gnd.n6936 gnd.n6935 19.3944
R10545 gnd.n6935 gnd.n6934 19.3944
R10546 gnd.n6934 gnd.n6933 19.3944
R10547 gnd.n6933 gnd.n6932 19.3944
R10548 gnd.n6932 gnd.n6929 19.3944
R10549 gnd.n6929 gnd.n357 19.3944
R10550 gnd.n7193 gnd.n357 19.3944
R10551 gnd.n7194 gnd.n7193 19.3944
R10552 gnd.n7194 gnd.n355 19.3944
R10553 gnd.n7200 gnd.n355 19.3944
R10554 gnd.n7200 gnd.n7199 19.3944
R10555 gnd.n7199 gnd.n334 19.3944
R10556 gnd.n7230 gnd.n334 19.3944
R10557 gnd.n7230 gnd.n332 19.3944
R10558 gnd.n7299 gnd.n332 19.3944
R10559 gnd.n7299 gnd.n7298 19.3944
R10560 gnd.n7298 gnd.n7297 19.3944
R10561 gnd.n7297 gnd.n7295 19.3944
R10562 gnd.n7295 gnd.n7294 19.3944
R10563 gnd.n7294 gnd.n7292 19.3944
R10564 gnd.n7292 gnd.n7291 19.3944
R10565 gnd.n7291 gnd.n7289 19.3944
R10566 gnd.n7289 gnd.n7288 19.3944
R10567 gnd.n7288 gnd.n7286 19.3944
R10568 gnd.n7286 gnd.n7285 19.3944
R10569 gnd.n7285 gnd.n7283 19.3944
R10570 gnd.n7283 gnd.n7282 19.3944
R10571 gnd.n7282 gnd.n7280 19.3944
R10572 gnd.n7280 gnd.n7279 19.3944
R10573 gnd.n7279 gnd.n7277 19.3944
R10574 gnd.n7277 gnd.n7276 19.3944
R10575 gnd.n7276 gnd.n7274 19.3944
R10576 gnd.n7274 gnd.n7273 19.3944
R10577 gnd.n7273 gnd.n7271 19.3944
R10578 gnd.n7271 gnd.n7270 19.3944
R10579 gnd.n7270 gnd.n7268 19.3944
R10580 gnd.n7268 gnd.n7267 19.3944
R10581 gnd.n7267 gnd.n7265 19.3944
R10582 gnd.n7265 gnd.n7264 19.3944
R10583 gnd.n7264 gnd.n7262 19.3944
R10584 gnd.n7262 gnd.n7261 19.3944
R10585 gnd.n7261 gnd.n200 19.3944
R10586 gnd.n7496 gnd.n200 19.3944
R10587 gnd.n7497 gnd.n7496 19.3944
R10588 gnd.n7535 gnd.n161 19.3944
R10589 gnd.n7530 gnd.n161 19.3944
R10590 gnd.n7530 gnd.n7529 19.3944
R10591 gnd.n7529 gnd.n7528 19.3944
R10592 gnd.n7528 gnd.n168 19.3944
R10593 gnd.n7523 gnd.n168 19.3944
R10594 gnd.n7523 gnd.n7522 19.3944
R10595 gnd.n7522 gnd.n7521 19.3944
R10596 gnd.n7521 gnd.n175 19.3944
R10597 gnd.n7516 gnd.n175 19.3944
R10598 gnd.n7516 gnd.n7515 19.3944
R10599 gnd.n7515 gnd.n7514 19.3944
R10600 gnd.n7514 gnd.n182 19.3944
R10601 gnd.n7509 gnd.n182 19.3944
R10602 gnd.n7509 gnd.n7508 19.3944
R10603 gnd.n7508 gnd.n7507 19.3944
R10604 gnd.n7507 gnd.n189 19.3944
R10605 gnd.n7502 gnd.n189 19.3944
R10606 gnd.n7568 gnd.n7567 19.3944
R10607 gnd.n7567 gnd.n7566 19.3944
R10608 gnd.n7566 gnd.n133 19.3944
R10609 gnd.n7561 gnd.n133 19.3944
R10610 gnd.n7561 gnd.n7560 19.3944
R10611 gnd.n7560 gnd.n7559 19.3944
R10612 gnd.n7559 gnd.n140 19.3944
R10613 gnd.n7554 gnd.n140 19.3944
R10614 gnd.n7554 gnd.n7553 19.3944
R10615 gnd.n7553 gnd.n7552 19.3944
R10616 gnd.n7552 gnd.n147 19.3944
R10617 gnd.n7547 gnd.n147 19.3944
R10618 gnd.n7547 gnd.n7546 19.3944
R10619 gnd.n7546 gnd.n7545 19.3944
R10620 gnd.n7545 gnd.n154 19.3944
R10621 gnd.n7540 gnd.n154 19.3944
R10622 gnd.n7540 gnd.n7539 19.3944
R10623 gnd.n7053 gnd.n485 19.3944
R10624 gnd.n7053 gnd.n469 19.3944
R10625 gnd.n7065 gnd.n469 19.3944
R10626 gnd.n7065 gnd.n467 19.3944
R10627 gnd.n7069 gnd.n467 19.3944
R10628 gnd.n7069 gnd.n452 19.3944
R10629 gnd.n7081 gnd.n452 19.3944
R10630 gnd.n7081 gnd.n450 19.3944
R10631 gnd.n7085 gnd.n450 19.3944
R10632 gnd.n7085 gnd.n435 19.3944
R10633 gnd.n7097 gnd.n435 19.3944
R10634 gnd.n7097 gnd.n433 19.3944
R10635 gnd.n7101 gnd.n433 19.3944
R10636 gnd.n7101 gnd.n418 19.3944
R10637 gnd.n7113 gnd.n418 19.3944
R10638 gnd.n7113 gnd.n416 19.3944
R10639 gnd.n7117 gnd.n416 19.3944
R10640 gnd.n7117 gnd.n399 19.3944
R10641 gnd.n7132 gnd.n399 19.3944
R10642 gnd.n7132 gnd.n397 19.3944
R10643 gnd.n7136 gnd.n397 19.3944
R10644 gnd.n7136 gnd.n367 19.3944
R10645 gnd.n7183 gnd.n367 19.3944
R10646 gnd.n7183 gnd.n365 19.3944
R10647 gnd.n7187 gnd.n365 19.3944
R10648 gnd.n7188 gnd.n7187 19.3944
R10649 gnd.n7188 gnd.n305 19.3944
R10650 gnd.n7323 gnd.n7322 19.3944
R10651 gnd.n338 gnd.n337 19.3944
R10652 gnd.n7226 gnd.n7225 19.3944
R10653 gnd.n328 gnd.n327 19.3944
R10654 gnd.n7303 gnd.n298 19.3944
R10655 gnd.n7327 gnd.n298 19.3944
R10656 gnd.n7327 gnd.n284 19.3944
R10657 gnd.n7339 gnd.n284 19.3944
R10658 gnd.n7339 gnd.n282 19.3944
R10659 gnd.n7343 gnd.n282 19.3944
R10660 gnd.n7343 gnd.n270 19.3944
R10661 gnd.n7355 gnd.n270 19.3944
R10662 gnd.n7355 gnd.n268 19.3944
R10663 gnd.n7359 gnd.n268 19.3944
R10664 gnd.n7359 gnd.n254 19.3944
R10665 gnd.n7371 gnd.n254 19.3944
R10666 gnd.n7371 gnd.n252 19.3944
R10667 gnd.n7375 gnd.n252 19.3944
R10668 gnd.n7375 gnd.n240 19.3944
R10669 gnd.n7387 gnd.n240 19.3944
R10670 gnd.n7387 gnd.n238 19.3944
R10671 gnd.n7391 gnd.n238 19.3944
R10672 gnd.n7391 gnd.n223 19.3944
R10673 gnd.n7403 gnd.n223 19.3944
R10674 gnd.n7403 gnd.n221 19.3944
R10675 gnd.n7407 gnd.n221 19.3944
R10676 gnd.n7407 gnd.n207 19.3944
R10677 gnd.n7487 gnd.n207 19.3944
R10678 gnd.n7487 gnd.n205 19.3944
R10679 gnd.n7491 gnd.n205 19.3944
R10680 gnd.n7491 gnd.n128 19.3944
R10681 gnd.n7571 gnd.n128 19.3944
R10682 gnd.n5065 gnd.n5064 19.3944
R10683 gnd.n5064 gnd.n4875 19.3944
R10684 gnd.n5059 gnd.n4875 19.3944
R10685 gnd.n5059 gnd.n5058 19.3944
R10686 gnd.n5058 gnd.n4880 19.3944
R10687 gnd.n5053 gnd.n4880 19.3944
R10688 gnd.n5053 gnd.n5052 19.3944
R10689 gnd.n5052 gnd.n5051 19.3944
R10690 gnd.n5051 gnd.n4886 19.3944
R10691 gnd.n5045 gnd.n4886 19.3944
R10692 gnd.n5045 gnd.n5044 19.3944
R10693 gnd.n5044 gnd.n5043 19.3944
R10694 gnd.n5043 gnd.n4892 19.3944
R10695 gnd.n5037 gnd.n4892 19.3944
R10696 gnd.n5037 gnd.n5036 19.3944
R10697 gnd.n5036 gnd.n5035 19.3944
R10698 gnd.n5035 gnd.n4898 19.3944
R10699 gnd.n5029 gnd.n5028 19.3944
R10700 gnd.n5028 gnd.n5027 19.3944
R10701 gnd.n5027 gnd.n4907 19.3944
R10702 gnd.n5021 gnd.n4907 19.3944
R10703 gnd.n5021 gnd.n5020 19.3944
R10704 gnd.n5020 gnd.n5019 19.3944
R10705 gnd.n5019 gnd.n4913 19.3944
R10706 gnd.n5013 gnd.n4913 19.3944
R10707 gnd.n5013 gnd.n5012 19.3944
R10708 gnd.n5012 gnd.n5011 19.3944
R10709 gnd.n5011 gnd.n4919 19.3944
R10710 gnd.n5005 gnd.n4919 19.3944
R10711 gnd.n5005 gnd.n5004 19.3944
R10712 gnd.n5004 gnd.n5003 19.3944
R10713 gnd.n5003 gnd.n4925 19.3944
R10714 gnd.n4997 gnd.n4925 19.3944
R10715 gnd.n4997 gnd.n4996 19.3944
R10716 gnd.n4996 gnd.n4995 19.3944
R10717 gnd.n5072 gnd.n1985 19.3944
R10718 gnd.n5076 gnd.n1985 19.3944
R10719 gnd.n5076 gnd.n1972 19.3944
R10720 gnd.n5088 gnd.n1972 19.3944
R10721 gnd.n5088 gnd.n1970 19.3944
R10722 gnd.n5092 gnd.n1970 19.3944
R10723 gnd.n5092 gnd.n1955 19.3944
R10724 gnd.n5104 gnd.n1955 19.3944
R10725 gnd.n5104 gnd.n1953 19.3944
R10726 gnd.n5108 gnd.n1953 19.3944
R10727 gnd.n5108 gnd.n1940 19.3944
R10728 gnd.n5120 gnd.n1940 19.3944
R10729 gnd.n5120 gnd.n1938 19.3944
R10730 gnd.n5124 gnd.n1938 19.3944
R10731 gnd.n5124 gnd.n1923 19.3944
R10732 gnd.n5136 gnd.n1923 19.3944
R10733 gnd.n5136 gnd.n1921 19.3944
R10734 gnd.n5148 gnd.n1921 19.3944
R10735 gnd.n5148 gnd.n5147 19.3944
R10736 gnd.n5147 gnd.n5146 19.3944
R10737 gnd.n5146 gnd.n5145 19.3944
R10738 gnd.n5145 gnd.n1887 19.3944
R10739 gnd.n5188 gnd.n1887 19.3944
R10740 gnd.n5188 gnd.n5187 19.3944
R10741 gnd.n5187 gnd.n5186 19.3944
R10742 gnd.n5186 gnd.n1896 19.3944
R10743 gnd.n1896 gnd.n1895 19.3944
R10744 gnd.n1895 gnd.n1778 19.3944
R10745 gnd.n5459 gnd.n1778 19.3944
R10746 gnd.n5459 gnd.n5458 19.3944
R10747 gnd.n5458 gnd.n5457 19.3944
R10748 gnd.n5457 gnd.n1782 19.3944
R10749 gnd.n5445 gnd.n1782 19.3944
R10750 gnd.n5445 gnd.n5444 19.3944
R10751 gnd.n5444 gnd.n5443 19.3944
R10752 gnd.n5443 gnd.n1756 19.3944
R10753 gnd.n5471 gnd.n1756 19.3944
R10754 gnd.n5471 gnd.n1754 19.3944
R10755 gnd.n5475 gnd.n1754 19.3944
R10756 gnd.n5475 gnd.n1740 19.3944
R10757 gnd.n5487 gnd.n1740 19.3944
R10758 gnd.n5487 gnd.n1738 19.3944
R10759 gnd.n5491 gnd.n1738 19.3944
R10760 gnd.n5491 gnd.n1722 19.3944
R10761 gnd.n5503 gnd.n1722 19.3944
R10762 gnd.n5503 gnd.n1720 19.3944
R10763 gnd.n5507 gnd.n1720 19.3944
R10764 gnd.n5507 gnd.n1706 19.3944
R10765 gnd.n5519 gnd.n1706 19.3944
R10766 gnd.n5519 gnd.n1704 19.3944
R10767 gnd.n5523 gnd.n1704 19.3944
R10768 gnd.n5523 gnd.n1688 19.3944
R10769 gnd.n5535 gnd.n1688 19.3944
R10770 gnd.n5535 gnd.n1686 19.3944
R10771 gnd.n5539 gnd.n1686 19.3944
R10772 gnd.n5539 gnd.n1672 19.3944
R10773 gnd.n5551 gnd.n1672 19.3944
R10774 gnd.n5551 gnd.n1670 19.3944
R10775 gnd.n5555 gnd.n1670 19.3944
R10776 gnd.n5555 gnd.n1653 19.3944
R10777 gnd.n5569 gnd.n1653 19.3944
R10778 gnd.n5569 gnd.n1651 19.3944
R10779 gnd.n5692 gnd.n1651 19.3944
R10780 gnd.n5692 gnd.n5691 19.3944
R10781 gnd.n4780 gnd.n4779 19.3944
R10782 gnd.n4785 gnd.n4780 19.3944
R10783 gnd.n4785 gnd.n4777 19.3944
R10784 gnd.n4789 gnd.n4777 19.3944
R10785 gnd.n4789 gnd.n4775 19.3944
R10786 gnd.n4795 gnd.n4775 19.3944
R10787 gnd.n4795 gnd.n4773 19.3944
R10788 gnd.n4799 gnd.n4773 19.3944
R10789 gnd.n4799 gnd.n4771 19.3944
R10790 gnd.n4805 gnd.n4771 19.3944
R10791 gnd.n4805 gnd.n4769 19.3944
R10792 gnd.n4809 gnd.n4769 19.3944
R10793 gnd.n4809 gnd.n4767 19.3944
R10794 gnd.n4815 gnd.n4767 19.3944
R10795 gnd.n4815 gnd.n4765 19.3944
R10796 gnd.n4819 gnd.n4765 19.3944
R10797 gnd.n4870 gnd.n4759 19.3944
R10798 gnd.n4870 gnd.n4869 19.3944
R10799 gnd.n4869 gnd.n4868 19.3944
R10800 gnd.n4868 gnd.n4866 19.3944
R10801 gnd.n4866 gnd.n4865 19.3944
R10802 gnd.n4865 gnd.n4863 19.3944
R10803 gnd.n4863 gnd.n4862 19.3944
R10804 gnd.n4862 gnd.n4860 19.3944
R10805 gnd.n4860 gnd.n4859 19.3944
R10806 gnd.n4859 gnd.n4857 19.3944
R10807 gnd.n4857 gnd.n4856 19.3944
R10808 gnd.n4856 gnd.n4854 19.3944
R10809 gnd.n4854 gnd.n4853 19.3944
R10810 gnd.n4853 gnd.n4851 19.3944
R10811 gnd.n4851 gnd.n4850 19.3944
R10812 gnd.n4850 gnd.n4848 19.3944
R10813 gnd.n4848 gnd.n4847 19.3944
R10814 gnd.n4847 gnd.n4845 19.3944
R10815 gnd.n4845 gnd.n1906 19.3944
R10816 gnd.n5162 gnd.n1906 19.3944
R10817 gnd.n5162 gnd.n1904 19.3944
R10818 gnd.n5171 gnd.n1904 19.3944
R10819 gnd.n5171 gnd.n5170 19.3944
R10820 gnd.n5170 gnd.n5169 19.3944
R10821 gnd.n5169 gnd.n1871 19.3944
R10822 gnd.n5201 gnd.n1871 19.3944
R10823 gnd.n5201 gnd.n1869 19.3944
R10824 gnd.n5215 gnd.n1869 19.3944
R10825 gnd.n5215 gnd.n5214 19.3944
R10826 gnd.n5214 gnd.n5213 19.3944
R10827 gnd.n5213 gnd.n5211 19.3944
R10828 gnd.n5211 gnd.n5210 19.3944
R10829 gnd.n5210 gnd.n1859 19.3944
R10830 gnd.n5235 gnd.n1859 19.3944
R10831 gnd.n5235 gnd.n1857 19.3944
R10832 gnd.n5239 gnd.n1857 19.3944
R10833 gnd.n5239 gnd.n1807 19.3944
R10834 gnd.n5427 gnd.n1807 19.3944
R10835 gnd.n5427 gnd.n1808 19.3944
R10836 gnd.n5423 gnd.n1808 19.3944
R10837 gnd.n5423 gnd.n5422 19.3944
R10838 gnd.n5422 gnd.n5421 19.3944
R10839 gnd.n5421 gnd.n1813 19.3944
R10840 gnd.n5417 gnd.n1813 19.3944
R10841 gnd.n5417 gnd.n5416 19.3944
R10842 gnd.n5416 gnd.n5415 19.3944
R10843 gnd.n5415 gnd.n1817 19.3944
R10844 gnd.n5411 gnd.n1817 19.3944
R10845 gnd.n5411 gnd.n5410 19.3944
R10846 gnd.n5410 gnd.n5409 19.3944
R10847 gnd.n5409 gnd.n1821 19.3944
R10848 gnd.n5405 gnd.n1821 19.3944
R10849 gnd.n5405 gnd.n5404 19.3944
R10850 gnd.n5404 gnd.n5403 19.3944
R10851 gnd.n5403 gnd.n1825 19.3944
R10852 gnd.n5399 gnd.n1825 19.3944
R10853 gnd.n5399 gnd.n5398 19.3944
R10854 gnd.n5398 gnd.n5397 19.3944
R10855 gnd.n5397 gnd.n1829 19.3944
R10856 gnd.n5393 gnd.n1829 19.3944
R10857 gnd.n5393 gnd.n5392 19.3944
R10858 gnd.n5392 gnd.n5391 19.3944
R10859 gnd.n5391 gnd.n5388 19.3944
R10860 gnd.n5388 gnd.n1353 19.3944
R10861 gnd.n4986 gnd.n4985 19.3944
R10862 gnd.n4985 gnd.n4984 19.3944
R10863 gnd.n4984 gnd.n4983 19.3944
R10864 gnd.n4983 gnd.n4981 19.3944
R10865 gnd.n4981 gnd.n4980 19.3944
R10866 gnd.n4980 gnd.n4978 19.3944
R10867 gnd.n4978 gnd.n4977 19.3944
R10868 gnd.n4977 gnd.n4975 19.3944
R10869 gnd.n4975 gnd.n4974 19.3944
R10870 gnd.n4974 gnd.n4972 19.3944
R10871 gnd.n4972 gnd.n4971 19.3944
R10872 gnd.n4971 gnd.n4969 19.3944
R10873 gnd.n4969 gnd.n4968 19.3944
R10874 gnd.n4968 gnd.n4966 19.3944
R10875 gnd.n4966 gnd.n4965 19.3944
R10876 gnd.n4965 gnd.n4963 19.3944
R10877 gnd.n4963 gnd.n4962 19.3944
R10878 gnd.n4962 gnd.n4960 19.3944
R10879 gnd.n4960 gnd.n4959 19.3944
R10880 gnd.n4959 gnd.n4957 19.3944
R10881 gnd.n4957 gnd.n1900 19.3944
R10882 gnd.n5175 gnd.n1900 19.3944
R10883 gnd.n5176 gnd.n5175 19.3944
R10884 gnd.n5176 gnd.n1898 19.3944
R10885 gnd.n5182 gnd.n1898 19.3944
R10886 gnd.n5182 gnd.n5181 19.3944
R10887 gnd.n5181 gnd.n1865 19.3944
R10888 gnd.n5219 gnd.n1865 19.3944
R10889 gnd.n5219 gnd.n1863 19.3944
R10890 gnd.n5224 gnd.n1863 19.3944
R10891 gnd.n5225 gnd.n5224 19.3944
R10892 gnd.n5227 gnd.n5225 19.3944
R10893 gnd.n5227 gnd.n1860 19.3944
R10894 gnd.n5231 gnd.n1860 19.3944
R10895 gnd.n5231 gnd.n1856 19.3944
R10896 gnd.n5243 gnd.n1856 19.3944
R10897 gnd.n5243 gnd.n1854 19.3944
R10898 gnd.n5247 gnd.n1854 19.3944
R10899 gnd.n5248 gnd.n5247 19.3944
R10900 gnd.n5251 gnd.n5248 19.3944
R10901 gnd.n5251 gnd.n1852 19.3944
R10902 gnd.n5278 gnd.n1852 19.3944
R10903 gnd.n5279 gnd.n5278 19.3944
R10904 gnd.n5282 gnd.n5279 19.3944
R10905 gnd.n5282 gnd.n1850 19.3944
R10906 gnd.n5293 gnd.n1850 19.3944
R10907 gnd.n5293 gnd.n5292 19.3944
R10908 gnd.n5292 gnd.n5291 19.3944
R10909 gnd.n5291 gnd.n1842 19.3944
R10910 gnd.n5318 gnd.n1842 19.3944
R10911 gnd.n5319 gnd.n5318 19.3944
R10912 gnd.n5322 gnd.n5319 19.3944
R10913 gnd.n5322 gnd.n1840 19.3944
R10914 gnd.n5332 gnd.n1840 19.3944
R10915 gnd.n5332 gnd.n5331 19.3944
R10916 gnd.n5331 gnd.n5330 19.3944
R10917 gnd.n5330 gnd.n1833 19.3944
R10918 gnd.n5375 gnd.n1833 19.3944
R10919 gnd.n5375 gnd.n1831 19.3944
R10920 gnd.n5382 gnd.n1831 19.3944
R10921 gnd.n5382 gnd.n5381 19.3944
R10922 gnd.n5381 gnd.n1647 19.3944
R10923 gnd.n5696 gnd.n1647 19.3944
R10924 gnd.n5697 gnd.n5696 19.3944
R10925 gnd.n5735 gnd.n5734 19.3944
R10926 gnd.n5734 gnd.n5733 19.3944
R10927 gnd.n5733 gnd.n1613 19.3944
R10928 gnd.n5728 gnd.n1613 19.3944
R10929 gnd.n5728 gnd.n5727 19.3944
R10930 gnd.n5727 gnd.n5726 19.3944
R10931 gnd.n5726 gnd.n1620 19.3944
R10932 gnd.n5721 gnd.n1620 19.3944
R10933 gnd.n5721 gnd.n5720 19.3944
R10934 gnd.n5720 gnd.n5719 19.3944
R10935 gnd.n5719 gnd.n1627 19.3944
R10936 gnd.n5714 gnd.n1627 19.3944
R10937 gnd.n5714 gnd.n5713 19.3944
R10938 gnd.n5713 gnd.n5712 19.3944
R10939 gnd.n5712 gnd.n1634 19.3944
R10940 gnd.n5707 gnd.n1634 19.3944
R10941 gnd.n5707 gnd.n5706 19.3944
R10942 gnd.n5706 gnd.n5705 19.3944
R10943 gnd.n5766 gnd.n5765 19.3944
R10944 gnd.n5765 gnd.n1363 19.3944
R10945 gnd.n1365 gnd.n1363 19.3944
R10946 gnd.n5758 gnd.n1365 19.3944
R10947 gnd.n5758 gnd.n5757 19.3944
R10948 gnd.n5757 gnd.n5756 19.3944
R10949 gnd.n5756 gnd.n1372 19.3944
R10950 gnd.n5751 gnd.n1372 19.3944
R10951 gnd.n5751 gnd.n5750 19.3944
R10952 gnd.n5750 gnd.n5749 19.3944
R10953 gnd.n5749 gnd.n1379 19.3944
R10954 gnd.n5744 gnd.n1379 19.3944
R10955 gnd.n5744 gnd.n5743 19.3944
R10956 gnd.n5743 gnd.n5742 19.3944
R10957 gnd.n5742 gnd.n1386 19.3944
R10958 gnd.n5068 gnd.n1980 19.3944
R10959 gnd.n5080 gnd.n1980 19.3944
R10960 gnd.n5080 gnd.n1978 19.3944
R10961 gnd.n5084 gnd.n1978 19.3944
R10962 gnd.n5084 gnd.n1964 19.3944
R10963 gnd.n5096 gnd.n1964 19.3944
R10964 gnd.n5096 gnd.n1962 19.3944
R10965 gnd.n5100 gnd.n1962 19.3944
R10966 gnd.n5100 gnd.n1948 19.3944
R10967 gnd.n5112 gnd.n1948 19.3944
R10968 gnd.n5112 gnd.n1946 19.3944
R10969 gnd.n5116 gnd.n1946 19.3944
R10970 gnd.n5116 gnd.n1932 19.3944
R10971 gnd.n5128 gnd.n1932 19.3944
R10972 gnd.n5128 gnd.n1930 19.3944
R10973 gnd.n5132 gnd.n1930 19.3944
R10974 gnd.n5132 gnd.n1915 19.3944
R10975 gnd.n5152 gnd.n1915 19.3944
R10976 gnd.n5152 gnd.n1913 19.3944
R10977 gnd.n5158 gnd.n1913 19.3944
R10978 gnd.n5158 gnd.n5157 19.3944
R10979 gnd.n5157 gnd.n1879 19.3944
R10980 gnd.n5192 gnd.n1879 19.3944
R10981 gnd.n5192 gnd.n1877 19.3944
R10982 gnd.n5196 gnd.n1877 19.3944
R10983 gnd.n5197 gnd.n5196 19.3944
R10984 gnd.n5197 gnd.n1770 19.3944
R10985 gnd.n5464 gnd.n5463 19.3944
R10986 gnd.n5453 gnd.n5452 19.3944
R10987 gnd.n5450 gnd.n5449 19.3944
R10988 gnd.n5439 gnd.n5438 19.3944
R10989 gnd.n5467 gnd.n1763 19.3944
R10990 gnd.n5467 gnd.n1748 19.3944
R10991 gnd.n5479 gnd.n1748 19.3944
R10992 gnd.n5479 gnd.n1746 19.3944
R10993 gnd.n5483 gnd.n1746 19.3944
R10994 gnd.n5483 gnd.n1731 19.3944
R10995 gnd.n5495 gnd.n1731 19.3944
R10996 gnd.n5495 gnd.n1729 19.3944
R10997 gnd.n5499 gnd.n1729 19.3944
R10998 gnd.n5499 gnd.n1714 19.3944
R10999 gnd.n5511 gnd.n1714 19.3944
R11000 gnd.n5511 gnd.n1712 19.3944
R11001 gnd.n5515 gnd.n1712 19.3944
R11002 gnd.n5515 gnd.n1697 19.3944
R11003 gnd.n5527 gnd.n1697 19.3944
R11004 gnd.n5527 gnd.n1695 19.3944
R11005 gnd.n5531 gnd.n1695 19.3944
R11006 gnd.n5531 gnd.n1680 19.3944
R11007 gnd.n5543 gnd.n1680 19.3944
R11008 gnd.n5543 gnd.n1678 19.3944
R11009 gnd.n5547 gnd.n1678 19.3944
R11010 gnd.n5547 gnd.n1663 19.3944
R11011 gnd.n5559 gnd.n1663 19.3944
R11012 gnd.n5559 gnd.n1661 19.3944
R11013 gnd.n5565 gnd.n1661 19.3944
R11014 gnd.n5565 gnd.n5564 19.3944
R11015 gnd.n5564 gnd.n1360 19.3944
R11016 gnd.n5769 gnd.n1360 19.3944
R11017 gnd.n3145 gnd.n2187 19.3944
R11018 gnd.n3145 gnd.n2185 19.3944
R11019 gnd.n3149 gnd.n2185 19.3944
R11020 gnd.n3149 gnd.n2181 19.3944
R11021 gnd.n3155 gnd.n2181 19.3944
R11022 gnd.n3155 gnd.n2179 19.3944
R11023 gnd.n3159 gnd.n2179 19.3944
R11024 gnd.n3159 gnd.n2175 19.3944
R11025 gnd.n3165 gnd.n2175 19.3944
R11026 gnd.n3165 gnd.n2173 19.3944
R11027 gnd.n3169 gnd.n2173 19.3944
R11028 gnd.n3169 gnd.n2169 19.3944
R11029 gnd.n3175 gnd.n2169 19.3944
R11030 gnd.n3175 gnd.n2167 19.3944
R11031 gnd.n3179 gnd.n2167 19.3944
R11032 gnd.n3179 gnd.n2163 19.3944
R11033 gnd.n3185 gnd.n2163 19.3944
R11034 gnd.n3185 gnd.n2161 19.3944
R11035 gnd.n3189 gnd.n2161 19.3944
R11036 gnd.n3189 gnd.n2157 19.3944
R11037 gnd.n3195 gnd.n2157 19.3944
R11038 gnd.n3195 gnd.n2155 19.3944
R11039 gnd.n3199 gnd.n2155 19.3944
R11040 gnd.n3199 gnd.n2151 19.3944
R11041 gnd.n3205 gnd.n2151 19.3944
R11042 gnd.n3205 gnd.n2149 19.3944
R11043 gnd.n3209 gnd.n2149 19.3944
R11044 gnd.n3209 gnd.n2145 19.3944
R11045 gnd.n3215 gnd.n2145 19.3944
R11046 gnd.n3215 gnd.n2143 19.3944
R11047 gnd.n3219 gnd.n2143 19.3944
R11048 gnd.n3219 gnd.n2139 19.3944
R11049 gnd.n3225 gnd.n2139 19.3944
R11050 gnd.n3225 gnd.n2137 19.3944
R11051 gnd.n3229 gnd.n2137 19.3944
R11052 gnd.n3229 gnd.n2133 19.3944
R11053 gnd.n3235 gnd.n2133 19.3944
R11054 gnd.n3235 gnd.n2131 19.3944
R11055 gnd.n3239 gnd.n2131 19.3944
R11056 gnd.n3239 gnd.n2127 19.3944
R11057 gnd.n3245 gnd.n2127 19.3944
R11058 gnd.n3245 gnd.n2125 19.3944
R11059 gnd.n3249 gnd.n2125 19.3944
R11060 gnd.n3249 gnd.n2121 19.3944
R11061 gnd.n3255 gnd.n2121 19.3944
R11062 gnd.n3255 gnd.n2119 19.3944
R11063 gnd.n3259 gnd.n2119 19.3944
R11064 gnd.n3259 gnd.n2115 19.3944
R11065 gnd.n3265 gnd.n2115 19.3944
R11066 gnd.n3265 gnd.n2113 19.3944
R11067 gnd.n3269 gnd.n2113 19.3944
R11068 gnd.n3269 gnd.n2109 19.3944
R11069 gnd.n3275 gnd.n2109 19.3944
R11070 gnd.n3275 gnd.n2107 19.3944
R11071 gnd.n3279 gnd.n2107 19.3944
R11072 gnd.n3279 gnd.n2103 19.3944
R11073 gnd.n3285 gnd.n2103 19.3944
R11074 gnd.n3285 gnd.n2101 19.3944
R11075 gnd.n3289 gnd.n2101 19.3944
R11076 gnd.n3289 gnd.n2097 19.3944
R11077 gnd.n3295 gnd.n2097 19.3944
R11078 gnd.n3295 gnd.n2095 19.3944
R11079 gnd.n3299 gnd.n2095 19.3944
R11080 gnd.n3299 gnd.n2091 19.3944
R11081 gnd.n3305 gnd.n2091 19.3944
R11082 gnd.n3305 gnd.n2089 19.3944
R11083 gnd.n3309 gnd.n2089 19.3944
R11084 gnd.n3309 gnd.n2085 19.3944
R11085 gnd.n3315 gnd.n2085 19.3944
R11086 gnd.n3315 gnd.n2083 19.3944
R11087 gnd.n3319 gnd.n2083 19.3944
R11088 gnd.n3319 gnd.n2079 19.3944
R11089 gnd.n3325 gnd.n2079 19.3944
R11090 gnd.n3325 gnd.n2077 19.3944
R11091 gnd.n3329 gnd.n2077 19.3944
R11092 gnd.n3329 gnd.n2073 19.3944
R11093 gnd.n3335 gnd.n2073 19.3944
R11094 gnd.n3335 gnd.n2071 19.3944
R11095 gnd.n3339 gnd.n2071 19.3944
R11096 gnd.n3339 gnd.n2067 19.3944
R11097 gnd.n3345 gnd.n2067 19.3944
R11098 gnd.n3345 gnd.n2065 19.3944
R11099 gnd.n3352 gnd.n2065 19.3944
R11100 gnd.n3352 gnd.n3351 19.3944
R11101 gnd.n5686 gnd.n5685 19.3944
R11102 gnd.n5685 gnd.n5684 19.3944
R11103 gnd.n5684 gnd.n5679 19.3944
R11104 gnd.n5680 gnd.n5679 19.3944
R11105 gnd.n5680 gnd.n1285 19.3944
R11106 gnd.n5846 gnd.n1285 19.3944
R11107 gnd.n5846 gnd.n1281 19.3944
R11108 gnd.n5850 gnd.n1281 19.3944
R11109 gnd.n5851 gnd.n5850 19.3944
R11110 gnd.n5855 gnd.n5851 19.3944
R11111 gnd.n5855 gnd.n1278 19.3944
R11112 gnd.n5965 gnd.n1278 19.3944
R11113 gnd.n5965 gnd.n1279 19.3944
R11114 gnd.n5961 gnd.n1279 19.3944
R11115 gnd.n5961 gnd.n5960 19.3944
R11116 gnd.n5960 gnd.n5959 19.3944
R11117 gnd.n5959 gnd.n5861 19.3944
R11118 gnd.n5955 gnd.n5861 19.3944
R11119 gnd.n5955 gnd.n5954 19.3944
R11120 gnd.n5954 gnd.n5953 19.3944
R11121 gnd.n5953 gnd.n5950 19.3944
R11122 gnd.n5950 gnd.n1197 19.3944
R11123 gnd.n6051 gnd.n1197 19.3944
R11124 gnd.n6051 gnd.n1193 19.3944
R11125 gnd.n6055 gnd.n1193 19.3944
R11126 gnd.n6056 gnd.n6055 19.3944
R11127 gnd.n6058 gnd.n6056 19.3944
R11128 gnd.n6058 gnd.n1191 19.3944
R11129 gnd.n6062 gnd.n1191 19.3944
R11130 gnd.n6063 gnd.n6062 19.3944
R11131 gnd.n6065 gnd.n6063 19.3944
R11132 gnd.n6065 gnd.n1189 19.3944
R11133 gnd.n6069 gnd.n1189 19.3944
R11134 gnd.n6070 gnd.n6069 19.3944
R11135 gnd.n6072 gnd.n6070 19.3944
R11136 gnd.n6072 gnd.n1186 19.3944
R11137 gnd.n6077 gnd.n1186 19.3944
R11138 gnd.n6077 gnd.n1187 19.3944
R11139 gnd.n1187 gnd.n1047 19.3944
R11140 gnd.n6194 gnd.n1047 19.3944
R11141 gnd.n6194 gnd.n1043 19.3944
R11142 gnd.n6198 gnd.n1043 19.3944
R11143 gnd.n6199 gnd.n6198 19.3944
R11144 gnd.n6201 gnd.n6199 19.3944
R11145 gnd.n6201 gnd.n1040 19.3944
R11146 gnd.n6412 gnd.n1040 19.3944
R11147 gnd.n6412 gnd.n1041 19.3944
R11148 gnd.n6408 gnd.n1041 19.3944
R11149 gnd.n6408 gnd.n6407 19.3944
R11150 gnd.n6407 gnd.n6406 19.3944
R11151 gnd.n6406 gnd.n6207 19.3944
R11152 gnd.n6402 gnd.n6207 19.3944
R11153 gnd.n6402 gnd.n6401 19.3944
R11154 gnd.n6401 gnd.n6400 19.3944
R11155 gnd.n6400 gnd.n6211 19.3944
R11156 gnd.n6396 gnd.n6211 19.3944
R11157 gnd.n6396 gnd.n6395 19.3944
R11158 gnd.n6395 gnd.n6394 19.3944
R11159 gnd.n6394 gnd.n6215 19.3944
R11160 gnd.n6390 gnd.n6215 19.3944
R11161 gnd.n6390 gnd.n6389 19.3944
R11162 gnd.n6389 gnd.n6388 19.3944
R11163 gnd.n6388 gnd.n6219 19.3944
R11164 gnd.n6384 gnd.n6219 19.3944
R11165 gnd.n6384 gnd.n6383 19.3944
R11166 gnd.n6383 gnd.n917 19.3944
R11167 gnd.n6544 gnd.n917 19.3944
R11168 gnd.n6544 gnd.n914 19.3944
R11169 gnd.n6549 gnd.n914 19.3944
R11170 gnd.n6549 gnd.n915 19.3944
R11171 gnd.n915 gnd.n876 19.3944
R11172 gnd.n6602 gnd.n876 19.3944
R11173 gnd.n6602 gnd.n873 19.3944
R11174 gnd.n6606 gnd.n873 19.3944
R11175 gnd.n6607 gnd.n6606 19.3944
R11176 gnd.n6609 gnd.n6607 19.3944
R11177 gnd.n6609 gnd.n870 19.3944
R11178 gnd.n6766 gnd.n870 19.3944
R11179 gnd.n6766 gnd.n871 19.3944
R11180 gnd.n6762 gnd.n871 19.3944
R11181 gnd.n6762 gnd.n6761 19.3944
R11182 gnd.n6761 gnd.n6760 19.3944
R11183 gnd.n6695 gnd.n6694 19.3944
R11184 gnd.n6694 gnd.n633 19.3944
R11185 gnd.n6814 gnd.n633 19.3944
R11186 gnd.n6757 gnd.n6616 19.3944
R11187 gnd.n6750 gnd.n6616 19.3944
R11188 gnd.n6750 gnd.n6749 19.3944
R11189 gnd.n6749 gnd.n6634 19.3944
R11190 gnd.n6742 gnd.n6634 19.3944
R11191 gnd.n6742 gnd.n6741 19.3944
R11192 gnd.n6741 gnd.n6642 19.3944
R11193 gnd.n6734 gnd.n6642 19.3944
R11194 gnd.n6734 gnd.n6733 19.3944
R11195 gnd.n6733 gnd.n6654 19.3944
R11196 gnd.n6726 gnd.n6654 19.3944
R11197 gnd.n6726 gnd.n6725 19.3944
R11198 gnd.n6725 gnd.n6662 19.3944
R11199 gnd.n6718 gnd.n6662 19.3944
R11200 gnd.n6718 gnd.n6717 19.3944
R11201 gnd.n6717 gnd.n6674 19.3944
R11202 gnd.n6707 gnd.n6674 19.3944
R11203 gnd.n6707 gnd.n6706 19.3944
R11204 gnd.n6706 gnd.n6705 19.3944
R11205 gnd.n6705 gnd.n6681 19.3944
R11206 gnd.n6701 gnd.n6681 19.3944
R11207 gnd.n6701 gnd.n6700 19.3944
R11208 gnd.n6700 gnd.n6699 19.3944
R11209 gnd.n6699 gnd.n6687 19.3944
R11210 gnd.n1200 gnd.t145 19.1199
R11211 gnd.n6141 gnd.n1093 19.1199
R11212 gnd.n6079 gnd.n1056 19.1199
R11213 gnd.n6446 gnd.n1006 19.1199
R11214 gnd.n6257 gnd.n968 19.1199
R11215 gnd.t148 gnd.n953 19.1199
R11216 gnd.n6798 gnd.n646 19.1199
R11217 gnd.n4179 gnd.t18 18.8012
R11218 gnd.n3612 gnd.t159 18.8012
R11219 gnd.n4049 gnd.n4048 18.4825
R11220 gnd.n6576 gnd.t101 18.4825
R11221 gnd.n7019 gnd.n7018 18.4247
R11222 gnd.n1606 gnd.n1386 18.4247
R11223 gnd.n7450 gnd.n120 18.2308
R11224 gnd.n6714 gnd.n6668 18.2308
R11225 gnd.n5775 gnd.n1347 18.2308
R11226 gnd.n4819 gnd.n4763 18.2308
R11227 gnd.t8 gnd.n3728 18.1639
R11228 gnd.n5852 gnd.t141 18.1639
R11229 gnd.t352 gnd.n879 18.1639
R11230 gnd.n6007 gnd.n1239 17.8452
R11231 gnd.n5883 gnd.n1216 17.8452
R11232 gnd.n1150 gnd.n1065 17.8452
R11233 gnd.n6454 gnd.n998 17.8452
R11234 gnd.n6381 gnd.n939 17.8452
R11235 gnd.n6551 gnd.n888 17.8452
R11236 gnd.n3757 gnd.t16 17.5266
R11237 gnd.n6149 gnd.t338 17.5266
R11238 gnd.n6306 gnd.t344 17.5266
R11239 gnd.n4657 gnd.n3355 17.2079
R11240 gnd.t143 gnd.n1248 17.2079
R11241 gnd.n6560 gnd.t173 17.2079
R11242 gnd.n7393 gnd.n236 17.2079
R11243 gnd.n4168 gnd.t12 16.8893
R11244 gnd.n5441 gnd.n1795 16.5706
R11245 gnd.n5469 gnd.n1758 16.5706
R11246 gnd.n5429 gnd.n1761 16.5706
R11247 gnd.n5249 gnd.n1752 16.5706
R11248 gnd.n5485 gnd.n1742 16.5706
R11249 gnd.n5276 gnd.n5275 16.5706
R11250 gnd.n5493 gnd.n1733 16.5706
R11251 gnd.n5501 gnd.n1724 16.5706
R11252 gnd.n5295 gnd.n1727 16.5706
R11253 gnd.n5289 gnd.n1718 16.5706
R11254 gnd.n5517 gnd.n1708 16.5706
R11255 gnd.n5316 gnd.n5315 16.5706
R11256 gnd.n5525 gnd.n1699 16.5706
R11257 gnd.n5533 gnd.n1690 16.5706
R11258 gnd.n5334 gnd.n1693 16.5706
R11259 gnd.n5328 gnd.n1684 16.5706
R11260 gnd.n5549 gnd.n1674 16.5706
R11261 gnd.n5373 gnd.n5372 16.5706
R11262 gnd.n5557 gnd.n1665 16.5706
R11263 gnd.n5384 gnd.n1668 16.5706
R11264 gnd.n5567 gnd.n1655 16.5706
R11265 gnd.n5386 gnd.n1658 16.5706
R11266 gnd.n5694 gnd.n1649 16.5706
R11267 gnd.n5771 gnd.n1354 16.5706
R11268 gnd.n6015 gnd.n1231 16.5706
R11269 gnd.n5920 gnd.n5888 16.5706
R11270 gnd.n6157 gnd.n1078 16.5706
R11271 gnd.n6094 gnd.n6093 16.5706
R11272 gnd.n6462 gnd.n990 16.5706
R11273 gnd.n6298 gnd.n6266 16.5706
R11274 gnd.n6374 gnd.n6373 16.5706
R11275 gnd.n6542 gnd.n920 16.5706
R11276 gnd.n6974 gnd.n480 16.5706
R11277 gnd.n7055 gnd.n483 16.5706
R11278 gnd.n6846 gnd.n471 16.5706
R11279 gnd.n7063 gnd.n474 16.5706
R11280 gnd.n6850 gnd.n462 16.5706
R11281 gnd.n7071 gnd.n465 16.5706
R11282 gnd.n6866 gnd.n6865 16.5706
R11283 gnd.n7079 gnd.n456 16.5706
R11284 gnd.n6859 gnd.n446 16.5706
R11285 gnd.n6886 gnd.n437 16.5706
R11286 gnd.n7095 gnd.n440 16.5706
R11287 gnd.n7103 gnd.n431 16.5706
R11288 gnd.n6905 gnd.n6904 16.5706
R11289 gnd.n7111 gnd.n422 16.5706
R11290 gnd.n6898 gnd.n412 16.5706
R11291 gnd.n6917 gnd.n401 16.5706
R11292 gnd.n7130 gnd.n404 16.5706
R11293 gnd.n7138 gnd.n386 16.5706
R11294 gnd.n7159 gnd.n7158 16.5706
R11295 gnd.n7181 gnd.n372 16.5706
R11296 gnd.n6930 gnd.n379 16.5706
R11297 gnd.n7190 gnd.n361 16.5706
R11298 gnd.n7212 gnd.n349 16.5706
R11299 gnd.n7320 gnd.n311 16.5706
R11300 gnd.n3984 gnd.t104 16.2519
R11301 gnd.n4216 gnd.t10 16.2519
R11302 gnd.n5437 gnd.t184 16.2519
R11303 gnd.n1312 gnd.t111 16.2519
R11304 gnd.n6808 gnd.t91 16.2519
R11305 gnd.t285 gnd.n308 16.2519
R11306 gnd.n5940 gnd.t161 15.9333
R11307 gnd.n6344 gnd.t162 15.9333
R11308 gnd.n4610 gnd.n4608 15.6674
R11309 gnd.n4578 gnd.n4576 15.6674
R11310 gnd.n4546 gnd.n4544 15.6674
R11311 gnd.n4515 gnd.n4513 15.6674
R11312 gnd.n4483 gnd.n4481 15.6674
R11313 gnd.n4451 gnd.n4449 15.6674
R11314 gnd.n4419 gnd.n4417 15.6674
R11315 gnd.n4388 gnd.n4386 15.6674
R11316 gnd.n3975 gnd.t104 15.6146
R11317 gnd.t56 gnd.n4646 15.6146
R11318 gnd.t81 gnd.n3364 15.6146
R11319 gnd.t186 gnd.n1736 15.6146
R11320 gnd.n5825 gnd.t111 15.6146
R11321 gnd.n6613 gnd.t91 15.6146
R11322 gnd.n7139 gnd.t227 15.6146
R11323 gnd.n5233 gnd.n1795 15.296
R11324 gnd.n5441 gnd.n5437 15.296
R11325 gnd.n5241 gnd.n1758 15.296
R11326 gnd.n5469 gnd.n1761 15.296
R11327 gnd.n5430 gnd.n5429 15.296
R11328 gnd.n5477 gnd.n1752 15.296
R11329 gnd.n5249 gnd.n1742 15.296
R11330 gnd.n5276 gnd.n1733 15.296
R11331 gnd.n5493 gnd.n1736 15.296
R11332 gnd.n5280 gnd.n1724 15.296
R11333 gnd.n5501 gnd.n1727 15.296
R11334 gnd.n5296 gnd.n5295 15.296
R11335 gnd.n5509 gnd.n1718 15.296
R11336 gnd.n5289 gnd.n1708 15.296
R11337 gnd.n5316 gnd.n1699 15.296
R11338 gnd.n5525 gnd.n1702 15.296
R11339 gnd.n5320 gnd.n1690 15.296
R11340 gnd.n5533 gnd.n1693 15.296
R11341 gnd.n5335 gnd.n5334 15.296
R11342 gnd.n5541 gnd.n1684 15.296
R11343 gnd.n5328 gnd.n1674 15.296
R11344 gnd.n5373 gnd.n1665 15.296
R11345 gnd.n5557 gnd.n1668 15.296
R11346 gnd.n5384 gnd.n1655 15.296
R11347 gnd.n5567 gnd.n1658 15.296
R11348 gnd.n5694 gnd.n1354 15.296
R11349 gnd.n5771 gnd.n1356 15.296
R11350 gnd.n6974 gnd.n564 15.296
R11351 gnd.n7055 gnd.n480 15.296
R11352 gnd.n7063 gnd.n471 15.296
R11353 gnd.n6850 gnd.n474 15.296
R11354 gnd.n7071 gnd.n462 15.296
R11355 gnd.n6865 gnd.n465 15.296
R11356 gnd.n6859 gnd.n456 15.296
R11357 gnd.n7087 gnd.n446 15.296
R11358 gnd.n6886 gnd.n6885 15.296
R11359 gnd.n7095 gnd.n437 15.296
R11360 gnd.n6890 gnd.n440 15.296
R11361 gnd.n7103 gnd.n428 15.296
R11362 gnd.n6904 gnd.n431 15.296
R11363 gnd.n6898 gnd.n422 15.296
R11364 gnd.n7119 gnd.n412 15.296
R11365 gnd.n6917 gnd.n6916 15.296
R11366 gnd.n7130 gnd.n401 15.296
R11367 gnd.n6938 gnd.n404 15.296
R11368 gnd.n7139 gnd.n7138 15.296
R11369 gnd.n7159 gnd.n386 15.296
R11370 gnd.n6930 gnd.n372 15.296
R11371 gnd.n7169 gnd.n379 15.296
R11372 gnd.n7190 gnd.n359 15.296
R11373 gnd.n361 gnd.n349 15.296
R11374 gnd.n7212 gnd.n7211 15.296
R11375 gnd.n7320 gnd.n308 15.296
R11376 gnd.n7202 gnd.n311 15.296
R11377 gnd.n713 gnd.n712 15.0827
R11378 gnd.n1422 gnd.n1417 15.0481
R11379 gnd.n723 gnd.n722 15.0481
R11380 gnd.n3440 gnd.t17 14.9773
R11381 gnd.t202 gnd.n1702 14.9773
R11382 gnd.t293 gnd.n428 14.9773
R11383 gnd.n6023 gnd.t168 14.6587
R11384 gnd.n6532 gnd.t175 14.6587
R11385 gnd.n3415 gnd.t137 14.34
R11386 gnd.n3398 gnd.t15 14.34
R11387 gnd.n5967 gnd.n1239 14.0214
R11388 gnd.t21 gnd.n1216 14.0214
R11389 gnd.n6109 gnd.n6108 14.0214
R11390 gnd.n6173 gnd.n1065 14.0214
R11391 gnd.n6414 gnd.n998 14.0214
R11392 gnd.n6478 gnd.n976 14.0214
R11393 gnd.t4 gnd.n939 14.0214
R11394 gnd.n6590 gnd.n888 14.0214
R11395 gnd.n6789 gnd.t28 14.0214
R11396 gnd.n4137 gnd.t139 13.7027
R11397 gnd.t166 gnd.n1233 13.7027
R11398 gnd.t346 gnd.n919 13.7027
R11399 gnd.n3841 gnd.n3840 13.5763
R11400 gnd.n4722 gnd.n2026 13.5763
R11401 gnd.n6981 gnd.n561 13.5763
R11402 gnd.n7502 gnd.n7501 13.5763
R11403 gnd.n4995 gnd.n4934 13.5763
R11404 gnd.n5705 gnd.n1643 13.5763
R11405 gnd.n4049 gnd.n3787 13.384
R11406 gnd.n1433 gnd.n1414 13.1884
R11407 gnd.n1428 gnd.n1427 13.1884
R11408 gnd.n1427 gnd.n1426 13.1884
R11409 gnd.n716 gnd.n711 13.1884
R11410 gnd.n717 gnd.n716 13.1884
R11411 gnd.n1429 gnd.n1416 13.146
R11412 gnd.n1425 gnd.n1416 13.146
R11413 gnd.n715 gnd.n714 13.146
R11414 gnd.n715 gnd.n710 13.146
R11415 gnd.n4611 gnd.n4607 12.8005
R11416 gnd.n4579 gnd.n4575 12.8005
R11417 gnd.n4547 gnd.n4543 12.8005
R11418 gnd.n4516 gnd.n4512 12.8005
R11419 gnd.n4484 gnd.n4480 12.8005
R11420 gnd.n4452 gnd.n4448 12.8005
R11421 gnd.n4420 gnd.n4416 12.8005
R11422 gnd.n4389 gnd.n4385 12.8005
R11423 gnd.n5835 gnd.n1295 12.7467
R11424 gnd.t60 gnd.t74 12.7467
R11425 gnd.n5853 gnd.n5852 12.7467
R11426 gnd.t0 gnd.n1231 12.7467
R11427 gnd.n6040 gnd.n1207 12.7467
R11428 gnd.n1119 gnd.n1093 12.7467
R11429 gnd.n6183 gnd.n1056 12.7467
R11430 gnd.t154 gnd.n1058 12.7467
R11431 gnd.n6422 gnd.t135 12.7467
R11432 gnd.n1033 gnd.n1006 12.7467
R11433 gnd.n6486 gnd.n968 12.7467
R11434 gnd.n6510 gnd.n947 12.7467
R11435 gnd.t1 gnd.n920 12.7467
R11436 gnd.n6600 gnd.n879 12.7467
R11437 gnd.t118 gnd.n898 12.7467
R11438 gnd.n1960 gnd.t192 12.4281
R11439 gnd.n5541 gnd.t204 12.4281
R11440 gnd.t170 gnd.n1207 12.4281
R11441 gnd.t150 gnd.n947 12.4281
R11442 gnd.n7087 gnd.t221 12.4281
R11443 gnd.t208 gnd.n225 12.4281
R11444 gnd.n3840 gnd.n3835 12.4126
R11445 gnd.n4725 gnd.n4722 12.4126
R11446 gnd.n6977 gnd.n561 12.4126
R11447 gnd.n7501 gnd.n196 12.4126
R11448 gnd.n4991 gnd.n4934 12.4126
R11449 gnd.n5700 gnd.n1643 12.4126
R11450 gnd.n1515 gnd.n1434 12.1761
R11451 gnd.n729 gnd.n728 12.1761
R11452 gnd.n4615 gnd.n4614 12.0247
R11453 gnd.n4583 gnd.n4582 12.0247
R11454 gnd.n4551 gnd.n4550 12.0247
R11455 gnd.n4520 gnd.n4519 12.0247
R11456 gnd.n4488 gnd.n4487 12.0247
R11457 gnd.n4456 gnd.n4455 12.0247
R11458 gnd.n4424 gnd.n4423 12.0247
R11459 gnd.n4393 gnd.n4392 12.0247
R11460 gnd.n1928 gnd.t252 11.7908
R11461 gnd.n5509 gnd.t223 11.7908
R11462 gnd.t67 gnd.n1649 11.7908
R11463 gnd.t49 gnd.n483 11.7908
R11464 gnd.n7119 gnd.t248 11.7908
R11465 gnd.t282 gnd.n256 11.7908
R11466 gnd.n5844 gnd.n1287 11.4721
R11467 gnd.n6049 gnd.n1199 11.4721
R11468 gnd.n1194 gnd.n1101 11.4721
R11469 gnd.n6192 gnd.n1049 11.4721
R11470 gnd.n1044 gnd.n1014 11.4721
R11471 gnd.n6494 gnd.n961 11.4721
R11472 gnd.n6502 gnd.n955 11.4721
R11473 gnd.n6577 gnd.n898 11.4721
R11474 gnd.n6775 gnd.n669 11.4721
R11475 gnd.n4618 gnd.n4605 11.249
R11476 gnd.n4586 gnd.n4573 11.249
R11477 gnd.n4554 gnd.n4541 11.249
R11478 gnd.n4523 gnd.n4510 11.249
R11479 gnd.n4491 gnd.n4478 11.249
R11480 gnd.n4459 gnd.n4446 11.249
R11481 gnd.n4427 gnd.n4414 11.249
R11482 gnd.n4396 gnd.n4383 11.249
R11483 gnd.n4127 gnd.t139 11.1535
R11484 gnd.n5184 gnd.t231 11.1535
R11485 gnd.n5477 gnd.t237 11.1535
R11486 gnd.n7169 gnd.t276 11.1535
R11487 gnd.t250 gnd.n286 11.1535
R11488 gnd.t115 gnd.n1295 10.8348
R11489 gnd.t3 gnd.n1103 10.8348
R11490 gnd.n6117 gnd.t3 10.8348
R11491 gnd.t22 gnd.n970 10.8348
R11492 gnd.n6326 gnd.t22 10.8348
R11493 gnd.n803 gnd.n802 10.6151
R11494 gnd.n807 gnd.n803 10.6151
R11495 gnd.n813 gnd.n691 10.6151
R11496 gnd.n814 gnd.n813 10.6151
R11497 gnd.n815 gnd.n814 10.6151
R11498 gnd.n815 gnd.n689 10.6151
R11499 gnd.n821 gnd.n689 10.6151
R11500 gnd.n822 gnd.n821 10.6151
R11501 gnd.n823 gnd.n822 10.6151
R11502 gnd.n823 gnd.n687 10.6151
R11503 gnd.n829 gnd.n687 10.6151
R11504 gnd.n830 gnd.n829 10.6151
R11505 gnd.n831 gnd.n830 10.6151
R11506 gnd.n831 gnd.n685 10.6151
R11507 gnd.n837 gnd.n685 10.6151
R11508 gnd.n838 gnd.n837 10.6151
R11509 gnd.n839 gnd.n838 10.6151
R11510 gnd.n839 gnd.n683 10.6151
R11511 gnd.n845 gnd.n683 10.6151
R11512 gnd.n846 gnd.n845 10.6151
R11513 gnd.n847 gnd.n846 10.6151
R11514 gnd.n847 gnd.n681 10.6151
R11515 gnd.n853 gnd.n681 10.6151
R11516 gnd.n854 gnd.n853 10.6151
R11517 gnd.n855 gnd.n854 10.6151
R11518 gnd.n855 gnd.n679 10.6151
R11519 gnd.n860 gnd.n679 10.6151
R11520 gnd.n861 gnd.n860 10.6151
R11521 gnd.n861 gnd.n677 10.6151
R11522 gnd.n866 gnd.n677 10.6151
R11523 gnd.n1535 gnd.n1410 10.6151
R11524 gnd.n1535 gnd.n1534 10.6151
R11525 gnd.n1534 gnd.n1533 10.6151
R11526 gnd.n1533 gnd.n1268 10.6151
R11527 gnd.n5981 gnd.n1268 10.6151
R11528 gnd.n5981 gnd.n5980 10.6151
R11529 gnd.n5980 gnd.n5979 10.6151
R11530 gnd.n5979 gnd.n1269 10.6151
R11531 gnd.n1271 gnd.n1269 10.6151
R11532 gnd.n5893 gnd.n1271 10.6151
R11533 gnd.n5895 gnd.n5893 10.6151
R11534 gnd.n5896 gnd.n5895 10.6151
R11535 gnd.n5898 gnd.n5896 10.6151
R11536 gnd.n5899 gnd.n5898 10.6151
R11537 gnd.n5900 gnd.n5899 10.6151
R11538 gnd.n5900 gnd.n5891 10.6151
R11539 gnd.n5915 gnd.n5891 10.6151
R11540 gnd.n5916 gnd.n5915 10.6151
R11541 gnd.n5918 gnd.n5916 10.6151
R11542 gnd.n5918 gnd.n5917 10.6151
R11543 gnd.n5917 gnd.n5882 10.6151
R11544 gnd.n5882 gnd.n5880 10.6151
R11545 gnd.n5931 gnd.n5880 10.6151
R11546 gnd.n5932 gnd.n5931 10.6151
R11547 gnd.n5934 gnd.n5932 10.6151
R11548 gnd.n5935 gnd.n5934 10.6151
R11549 gnd.n5937 gnd.n5935 10.6151
R11550 gnd.n5937 gnd.n5936 10.6151
R11551 gnd.n5936 gnd.n1115 10.6151
R11552 gnd.n6123 gnd.n1115 10.6151
R11553 gnd.n6123 gnd.n6122 10.6151
R11554 gnd.n6122 gnd.n6121 10.6151
R11555 gnd.n6121 gnd.n1116 10.6151
R11556 gnd.n1118 gnd.n1116 10.6151
R11557 gnd.n1128 gnd.n1118 10.6151
R11558 gnd.n1130 gnd.n1128 10.6151
R11559 gnd.n1131 gnd.n1130 10.6151
R11560 gnd.n6106 gnd.n1131 10.6151
R11561 gnd.n6106 gnd.n6105 10.6151
R11562 gnd.n6105 gnd.n6104 10.6151
R11563 gnd.n6104 gnd.n1132 10.6151
R11564 gnd.n1145 gnd.n1132 10.6151
R11565 gnd.n1146 gnd.n1145 10.6151
R11566 gnd.n6091 gnd.n1146 10.6151
R11567 gnd.n6091 gnd.n6090 10.6151
R11568 gnd.n6090 gnd.n6089 10.6151
R11569 gnd.n6089 gnd.n1147 10.6151
R11570 gnd.n1159 gnd.n1147 10.6151
R11571 gnd.n1184 gnd.n1159 10.6151
R11572 gnd.n1184 gnd.n1183 10.6151
R11573 gnd.n1183 gnd.n1182 10.6151
R11574 gnd.n1182 gnd.n1160 10.6151
R11575 gnd.n1161 gnd.n1160 10.6151
R11576 gnd.n1161 gnd.n1029 10.6151
R11577 gnd.n6428 gnd.n1029 10.6151
R11578 gnd.n6428 gnd.n6427 10.6151
R11579 gnd.n6427 gnd.n6426 10.6151
R11580 gnd.n6426 gnd.n1030 10.6151
R11581 gnd.n1032 gnd.n1030 10.6151
R11582 gnd.n6276 gnd.n1032 10.6151
R11583 gnd.n6278 gnd.n6276 10.6151
R11584 gnd.n6279 gnd.n6278 10.6151
R11585 gnd.n6281 gnd.n6279 10.6151
R11586 gnd.n6282 gnd.n6281 10.6151
R11587 gnd.n6286 gnd.n6282 10.6151
R11588 gnd.n6286 gnd.n6285 10.6151
R11589 gnd.n6285 gnd.n6284 10.6151
R11590 gnd.n6284 gnd.n6264 10.6151
R11591 gnd.n6300 gnd.n6264 10.6151
R11592 gnd.n6301 gnd.n6300 10.6151
R11593 gnd.n6304 gnd.n6301 10.6151
R11594 gnd.n6304 gnd.n6303 10.6151
R11595 gnd.n6303 gnd.n6302 10.6151
R11596 gnd.n6302 gnd.n6254 10.6151
R11597 gnd.n6319 gnd.n6254 10.6151
R11598 gnd.n6320 gnd.n6319 10.6151
R11599 gnd.n6323 gnd.n6320 10.6151
R11600 gnd.n6323 gnd.n6322 10.6151
R11601 gnd.n6322 gnd.n6321 10.6151
R11602 gnd.n6321 gnd.n6245 10.6151
R11603 gnd.n6338 gnd.n6245 10.6151
R11604 gnd.n6339 gnd.n6338 10.6151
R11605 gnd.n6342 gnd.n6339 10.6151
R11606 gnd.n6342 gnd.n6341 10.6151
R11607 gnd.n6341 gnd.n6340 10.6151
R11608 gnd.n6340 gnd.n6236 10.6151
R11609 gnd.n6236 gnd.n6234 10.6151
R11610 gnd.n6356 gnd.n6234 10.6151
R11611 gnd.n6357 gnd.n6356 10.6151
R11612 gnd.n6359 gnd.n6357 10.6151
R11613 gnd.n6360 gnd.n6359 10.6151
R11614 gnd.n6370 gnd.n6360 10.6151
R11615 gnd.n6370 gnd.n6369 10.6151
R11616 gnd.n6369 gnd.n6368 10.6151
R11617 gnd.n6368 gnd.n6365 10.6151
R11618 gnd.n6365 gnd.n6364 10.6151
R11619 gnd.n6364 gnd.n6363 10.6151
R11620 gnd.n6363 gnd.n6361 10.6151
R11621 gnd.n6361 gnd.n904 10.6151
R11622 gnd.n6563 gnd.n904 10.6151
R11623 gnd.n6564 gnd.n6563 10.6151
R11624 gnd.n6566 gnd.n6564 10.6151
R11625 gnd.n6566 gnd.n6565 10.6151
R11626 gnd.n6565 gnd.n666 10.6151
R11627 gnd.n6779 gnd.n666 10.6151
R11628 gnd.n6779 gnd.n6778 10.6151
R11629 gnd.n6778 gnd.n6777 10.6151
R11630 gnd.n6777 gnd.n667 10.6151
R11631 gnd.n868 gnd.n667 10.6151
R11632 gnd.n868 gnd.n867 10.6151
R11633 gnd.n1599 gnd.n1390 10.6151
R11634 gnd.n1599 gnd.n1598 10.6151
R11635 gnd.n1596 gnd.n1396 10.6151
R11636 gnd.n1590 gnd.n1396 10.6151
R11637 gnd.n1590 gnd.n1589 10.6151
R11638 gnd.n1589 gnd.n1588 10.6151
R11639 gnd.n1588 gnd.n1398 10.6151
R11640 gnd.n1582 gnd.n1398 10.6151
R11641 gnd.n1582 gnd.n1581 10.6151
R11642 gnd.n1581 gnd.n1580 10.6151
R11643 gnd.n1580 gnd.n1400 10.6151
R11644 gnd.n1574 gnd.n1400 10.6151
R11645 gnd.n1574 gnd.n1573 10.6151
R11646 gnd.n1573 gnd.n1572 10.6151
R11647 gnd.n1572 gnd.n1402 10.6151
R11648 gnd.n1566 gnd.n1402 10.6151
R11649 gnd.n1566 gnd.n1565 10.6151
R11650 gnd.n1565 gnd.n1564 10.6151
R11651 gnd.n1564 gnd.n1404 10.6151
R11652 gnd.n1558 gnd.n1404 10.6151
R11653 gnd.n1558 gnd.n1557 10.6151
R11654 gnd.n1557 gnd.n1556 10.6151
R11655 gnd.n1556 gnd.n1406 10.6151
R11656 gnd.n1550 gnd.n1406 10.6151
R11657 gnd.n1550 gnd.n1549 10.6151
R11658 gnd.n1549 gnd.n1548 10.6151
R11659 gnd.n1548 gnd.n1408 10.6151
R11660 gnd.n1542 gnd.n1408 10.6151
R11661 gnd.n1542 gnd.n1541 10.6151
R11662 gnd.n1541 gnd.n1540 10.6151
R11663 gnd.n1515 gnd.n1514 10.6151
R11664 gnd.n1514 gnd.n1436 10.6151
R11665 gnd.n1510 gnd.n1436 10.6151
R11666 gnd.n1510 gnd.n1509 10.6151
R11667 gnd.n1509 gnd.n1438 10.6151
R11668 gnd.n1504 gnd.n1438 10.6151
R11669 gnd.n1504 gnd.n1503 10.6151
R11670 gnd.n1503 gnd.n1502 10.6151
R11671 gnd.n1502 gnd.n1440 10.6151
R11672 gnd.n1496 gnd.n1440 10.6151
R11673 gnd.n1496 gnd.n1495 10.6151
R11674 gnd.n1495 gnd.n1494 10.6151
R11675 gnd.n1494 gnd.n1442 10.6151
R11676 gnd.n1488 gnd.n1442 10.6151
R11677 gnd.n1488 gnd.n1487 10.6151
R11678 gnd.n1487 gnd.n1486 10.6151
R11679 gnd.n1486 gnd.n1444 10.6151
R11680 gnd.n1480 gnd.n1444 10.6151
R11681 gnd.n1480 gnd.n1479 10.6151
R11682 gnd.n1479 gnd.n1478 10.6151
R11683 gnd.n1478 gnd.n1446 10.6151
R11684 gnd.n1472 gnd.n1446 10.6151
R11685 gnd.n1472 gnd.n1471 10.6151
R11686 gnd.n1471 gnd.n1470 10.6151
R11687 gnd.n1470 gnd.n1448 10.6151
R11688 gnd.n1464 gnd.n1448 10.6151
R11689 gnd.n1464 gnd.n1463 10.6151
R11690 gnd.n1463 gnd.n1462 10.6151
R11691 gnd.n1458 gnd.n1457 10.6151
R11692 gnd.n1457 gnd.n1391 10.6151
R11693 gnd.n729 gnd.n708 10.6151
R11694 gnd.n735 gnd.n708 10.6151
R11695 gnd.n736 gnd.n735 10.6151
R11696 gnd.n737 gnd.n736 10.6151
R11697 gnd.n737 gnd.n706 10.6151
R11698 gnd.n743 gnd.n706 10.6151
R11699 gnd.n744 gnd.n743 10.6151
R11700 gnd.n745 gnd.n744 10.6151
R11701 gnd.n745 gnd.n704 10.6151
R11702 gnd.n751 gnd.n704 10.6151
R11703 gnd.n752 gnd.n751 10.6151
R11704 gnd.n753 gnd.n752 10.6151
R11705 gnd.n753 gnd.n702 10.6151
R11706 gnd.n759 gnd.n702 10.6151
R11707 gnd.n760 gnd.n759 10.6151
R11708 gnd.n761 gnd.n760 10.6151
R11709 gnd.n761 gnd.n700 10.6151
R11710 gnd.n767 gnd.n700 10.6151
R11711 gnd.n768 gnd.n767 10.6151
R11712 gnd.n769 gnd.n768 10.6151
R11713 gnd.n769 gnd.n698 10.6151
R11714 gnd.n775 gnd.n698 10.6151
R11715 gnd.n776 gnd.n775 10.6151
R11716 gnd.n777 gnd.n776 10.6151
R11717 gnd.n777 gnd.n696 10.6151
R11718 gnd.n783 gnd.n696 10.6151
R11719 gnd.n784 gnd.n783 10.6151
R11720 gnd.n788 gnd.n784 10.6151
R11721 gnd.n793 gnd.n694 10.6151
R11722 gnd.n794 gnd.n793 10.6151
R11723 gnd.n1519 gnd.n1518 10.6151
R11724 gnd.n1528 gnd.n1519 10.6151
R11725 gnd.n1528 gnd.n1527 10.6151
R11726 gnd.n1527 gnd.n1526 10.6151
R11727 gnd.n1526 gnd.n1524 10.6151
R11728 gnd.n1524 gnd.n1523 10.6151
R11729 gnd.n1523 gnd.n1520 10.6151
R11730 gnd.n1520 gnd.n1274 10.6151
R11731 gnd.n5973 gnd.n1274 10.6151
R11732 gnd.n5973 gnd.n5972 10.6151
R11733 gnd.n5972 gnd.n5971 10.6151
R11734 gnd.n5971 gnd.n1275 10.6151
R11735 gnd.n5904 gnd.n1275 10.6151
R11736 gnd.n5905 gnd.n5904 10.6151
R11737 gnd.n5909 gnd.n5905 10.6151
R11738 gnd.n5909 gnd.n5908 10.6151
R11739 gnd.n5908 gnd.n5907 10.6151
R11740 gnd.n5907 gnd.n5886 10.6151
R11741 gnd.n5922 gnd.n5886 10.6151
R11742 gnd.n5923 gnd.n5922 10.6151
R11743 gnd.n5925 gnd.n5923 10.6151
R11744 gnd.n5925 gnd.n5924 10.6151
R11745 gnd.n5924 gnd.n5867 10.6151
R11746 gnd.n5945 gnd.n5867 10.6151
R11747 gnd.n5945 gnd.n5944 10.6151
R11748 gnd.n5944 gnd.n5943 10.6151
R11749 gnd.n5943 gnd.n5868 10.6151
R11750 gnd.n5876 gnd.n5868 10.6151
R11751 gnd.n5876 gnd.n5875 10.6151
R11752 gnd.n5875 gnd.n5874 10.6151
R11753 gnd.n5874 gnd.n5873 10.6151
R11754 gnd.n5873 gnd.n5870 10.6151
R11755 gnd.n5870 gnd.n1122 10.6151
R11756 gnd.n6115 gnd.n1122 10.6151
R11757 gnd.n6115 gnd.n6114 10.6151
R11758 gnd.n6114 gnd.n6113 10.6151
R11759 gnd.n6113 gnd.n1123 10.6151
R11760 gnd.n1137 gnd.n1123 10.6151
R11761 gnd.n1138 gnd.n1137 10.6151
R11762 gnd.n6100 gnd.n1138 10.6151
R11763 gnd.n6100 gnd.n6099 10.6151
R11764 gnd.n6099 gnd.n6098 10.6151
R11765 gnd.n6098 gnd.n1139 10.6151
R11766 gnd.n1153 gnd.n1139 10.6151
R11767 gnd.n1154 gnd.n1153 10.6151
R11768 gnd.n6085 gnd.n1154 10.6151
R11769 gnd.n6085 gnd.n6084 10.6151
R11770 gnd.n6084 gnd.n6083 10.6151
R11771 gnd.n6083 gnd.n1155 10.6151
R11772 gnd.n1167 gnd.n1155 10.6151
R11773 gnd.n1168 gnd.n1167 10.6151
R11774 gnd.n1177 gnd.n1168 10.6151
R11775 gnd.n1177 gnd.n1176 10.6151
R11776 gnd.n1176 gnd.n1175 10.6151
R11777 gnd.n1175 gnd.n1173 10.6151
R11778 gnd.n1173 gnd.n1172 10.6151
R11779 gnd.n1172 gnd.n1169 10.6151
R11780 gnd.n1169 gnd.n1036 10.6151
R11781 gnd.n6420 gnd.n1036 10.6151
R11782 gnd.n6420 gnd.n6419 10.6151
R11783 gnd.n6419 gnd.n6418 10.6151
R11784 gnd.n6418 gnd.n1037 10.6151
R11785 gnd.n6271 gnd.n1037 10.6151
R11786 gnd.n6272 gnd.n6271 10.6151
R11787 gnd.n6273 gnd.n6272 10.6151
R11788 gnd.n6273 gnd.n6269 10.6151
R11789 gnd.n6293 gnd.n6269 10.6151
R11790 gnd.n6294 gnd.n6293 10.6151
R11791 gnd.n6296 gnd.n6294 10.6151
R11792 gnd.n6296 gnd.n6295 10.6151
R11793 gnd.n6295 gnd.n6260 10.6151
R11794 gnd.n6310 gnd.n6260 10.6151
R11795 gnd.n6311 gnd.n6310 10.6151
R11796 gnd.n6314 gnd.n6311 10.6151
R11797 gnd.n6314 gnd.n6313 10.6151
R11798 gnd.n6313 gnd.n6312 10.6151
R11799 gnd.n6312 gnd.n6250 10.6151
R11800 gnd.n6329 gnd.n6250 10.6151
R11801 gnd.n6330 gnd.n6329 10.6151
R11802 gnd.n6333 gnd.n6330 10.6151
R11803 gnd.n6333 gnd.n6332 10.6151
R11804 gnd.n6332 gnd.n6331 10.6151
R11805 gnd.n6331 gnd.n6240 10.6151
R11806 gnd.n6347 gnd.n6240 10.6151
R11807 gnd.n6348 gnd.n6347 10.6151
R11808 gnd.n6350 gnd.n6348 10.6151
R11809 gnd.n6350 gnd.n6349 10.6151
R11810 gnd.n6349 gnd.n6224 10.6151
R11811 gnd.n6378 gnd.n6224 10.6151
R11812 gnd.n6378 gnd.n6377 10.6151
R11813 gnd.n6377 gnd.n6376 10.6151
R11814 gnd.n6376 gnd.n6225 10.6151
R11815 gnd.n6229 gnd.n6225 10.6151
R11816 gnd.n6229 gnd.n6228 10.6151
R11817 gnd.n6228 gnd.n6227 10.6151
R11818 gnd.n6227 gnd.n909 10.6151
R11819 gnd.n6555 gnd.n909 10.6151
R11820 gnd.n6556 gnd.n6555 10.6151
R11821 gnd.n6558 gnd.n6556 10.6151
R11822 gnd.n6558 gnd.n6557 10.6151
R11823 gnd.n6557 gnd.n900 10.6151
R11824 gnd.n6571 gnd.n900 10.6151
R11825 gnd.n6572 gnd.n6571 10.6151
R11826 gnd.n6574 gnd.n6572 10.6151
R11827 gnd.n6574 gnd.n6573 10.6151
R11828 gnd.n6573 gnd.n673 10.6151
R11829 gnd.n6773 gnd.n673 10.6151
R11830 gnd.n6773 gnd.n6772 10.6151
R11831 gnd.n6772 gnd.n6771 10.6151
R11832 gnd.n6771 gnd.n674 10.6151
R11833 gnd.n4038 gnd.t340 10.5161
R11834 gnd.n4349 gnd.t137 10.5161
R11835 gnd.t15 gnd.n3387 10.5161
R11836 gnd.n5455 gnd.t194 10.5161
R11837 gnd.n5447 gnd.n1788 10.5161
R11838 gnd.n5447 gnd.t215 10.5161
R11839 gnd.n7222 gnd.t206 10.5161
R11840 gnd.n7222 gnd.n7221 10.5161
R11841 gnd.n7228 gnd.t289 10.5161
R11842 gnd.n4619 gnd.n4603 10.4732
R11843 gnd.n4587 gnd.n4571 10.4732
R11844 gnd.n4555 gnd.n4539 10.4732
R11845 gnd.n4524 gnd.n4508 10.4732
R11846 gnd.n4492 gnd.n4476 10.4732
R11847 gnd.n4460 gnd.n4444 10.4732
R11848 gnd.n4428 gnd.n4412 10.4732
R11849 gnd.n4397 gnd.n4381 10.4732
R11850 gnd.n5844 gnd.n1288 10.1975
R11851 gnd.n1282 gnd.n1264 10.1975
R11852 gnd.n6049 gnd.n1200 10.1975
R11853 gnd.n6192 gnd.n1022 10.1975
R11854 gnd.n1044 gnd.n1025 10.1975
R11855 gnd.n6502 gnd.n953 10.1975
R11856 gnd.n6577 gnd.n6576 10.1975
R11857 gnd.n670 gnd.n669 10.1975
R11858 gnd.n4318 gnd.t17 9.87883
R11859 gnd.n5190 gnd.t190 9.87883
R11860 gnd.n5485 gnd.t198 9.87883
R11861 gnd.n7181 gnd.t211 9.87883
R11862 gnd.n289 gnd.t240 9.87883
R11863 gnd.n7627 gnd.n74 9.81789
R11864 gnd.n4623 gnd.n4622 9.69747
R11865 gnd.n4591 gnd.n4590 9.69747
R11866 gnd.n4559 gnd.n4558 9.69747
R11867 gnd.n4528 gnd.n4527 9.69747
R11868 gnd.n4496 gnd.n4495 9.69747
R11869 gnd.n4464 gnd.n4463 9.69747
R11870 gnd.n4432 gnd.n4431 9.69747
R11871 gnd.n4401 gnd.n4400 9.69747
R11872 gnd.n1134 gnd.t144 9.56018
R11873 gnd.n6470 gnd.t136 9.56018
R11874 gnd.n5689 gnd.n5573 9.45599
R11875 gnd.n6622 gnd.n6620 9.45599
R11876 gnd.n4629 gnd.n4628 9.45567
R11877 gnd.n4597 gnd.n4596 9.45567
R11878 gnd.n4565 gnd.n4564 9.45567
R11879 gnd.n4534 gnd.n4533 9.45567
R11880 gnd.n4502 gnd.n4501 9.45567
R11881 gnd.n4470 gnd.n4469 9.45567
R11882 gnd.n4438 gnd.n4437 9.45567
R11883 gnd.n4407 gnd.n4406 9.45567
R11884 gnd.n3676 gnd.n3675 9.39724
R11885 gnd.n4628 gnd.n4627 9.3005
R11886 gnd.n4601 gnd.n4600 9.3005
R11887 gnd.n4622 gnd.n4621 9.3005
R11888 gnd.n4620 gnd.n4619 9.3005
R11889 gnd.n4605 gnd.n4604 9.3005
R11890 gnd.n4614 gnd.n4613 9.3005
R11891 gnd.n4612 gnd.n4611 9.3005
R11892 gnd.n4596 gnd.n4595 9.3005
R11893 gnd.n4569 gnd.n4568 9.3005
R11894 gnd.n4590 gnd.n4589 9.3005
R11895 gnd.n4588 gnd.n4587 9.3005
R11896 gnd.n4573 gnd.n4572 9.3005
R11897 gnd.n4582 gnd.n4581 9.3005
R11898 gnd.n4580 gnd.n4579 9.3005
R11899 gnd.n4564 gnd.n4563 9.3005
R11900 gnd.n4537 gnd.n4536 9.3005
R11901 gnd.n4558 gnd.n4557 9.3005
R11902 gnd.n4556 gnd.n4555 9.3005
R11903 gnd.n4541 gnd.n4540 9.3005
R11904 gnd.n4550 gnd.n4549 9.3005
R11905 gnd.n4548 gnd.n4547 9.3005
R11906 gnd.n4533 gnd.n4532 9.3005
R11907 gnd.n4506 gnd.n4505 9.3005
R11908 gnd.n4527 gnd.n4526 9.3005
R11909 gnd.n4525 gnd.n4524 9.3005
R11910 gnd.n4510 gnd.n4509 9.3005
R11911 gnd.n4519 gnd.n4518 9.3005
R11912 gnd.n4517 gnd.n4516 9.3005
R11913 gnd.n4501 gnd.n4500 9.3005
R11914 gnd.n4474 gnd.n4473 9.3005
R11915 gnd.n4495 gnd.n4494 9.3005
R11916 gnd.n4493 gnd.n4492 9.3005
R11917 gnd.n4478 gnd.n4477 9.3005
R11918 gnd.n4487 gnd.n4486 9.3005
R11919 gnd.n4485 gnd.n4484 9.3005
R11920 gnd.n4469 gnd.n4468 9.3005
R11921 gnd.n4442 gnd.n4441 9.3005
R11922 gnd.n4463 gnd.n4462 9.3005
R11923 gnd.n4461 gnd.n4460 9.3005
R11924 gnd.n4446 gnd.n4445 9.3005
R11925 gnd.n4455 gnd.n4454 9.3005
R11926 gnd.n4453 gnd.n4452 9.3005
R11927 gnd.n4437 gnd.n4436 9.3005
R11928 gnd.n4410 gnd.n4409 9.3005
R11929 gnd.n4431 gnd.n4430 9.3005
R11930 gnd.n4429 gnd.n4428 9.3005
R11931 gnd.n4414 gnd.n4413 9.3005
R11932 gnd.n4423 gnd.n4422 9.3005
R11933 gnd.n4421 gnd.n4420 9.3005
R11934 gnd.n4406 gnd.n4405 9.3005
R11935 gnd.n4379 gnd.n4378 9.3005
R11936 gnd.n4400 gnd.n4399 9.3005
R11937 gnd.n4398 gnd.n4397 9.3005
R11938 gnd.n4383 gnd.n4382 9.3005
R11939 gnd.n4392 gnd.n4391 9.3005
R11940 gnd.n4390 gnd.n4389 9.3005
R11941 gnd.n4752 gnd.n4751 9.3005
R11942 gnd.n4750 gnd.n2014 9.3005
R11943 gnd.n4749 gnd.n4748 9.3005
R11944 gnd.n4745 gnd.n2015 9.3005
R11945 gnd.n4742 gnd.n2016 9.3005
R11946 gnd.n4741 gnd.n2017 9.3005
R11947 gnd.n4738 gnd.n2018 9.3005
R11948 gnd.n4737 gnd.n2019 9.3005
R11949 gnd.n4734 gnd.n2020 9.3005
R11950 gnd.n4733 gnd.n2021 9.3005
R11951 gnd.n4730 gnd.n2022 9.3005
R11952 gnd.n4729 gnd.n2023 9.3005
R11953 gnd.n4726 gnd.n2024 9.3005
R11954 gnd.n4725 gnd.n2025 9.3005
R11955 gnd.n4722 gnd.n4721 9.3005
R11956 gnd.n4720 gnd.n2026 9.3005
R11957 gnd.n4753 gnd.n2013 9.3005
R11958 gnd.n4057 gnd.n4056 9.3005
R11959 gnd.n3761 gnd.n3760 9.3005
R11960 gnd.n4084 gnd.n4083 9.3005
R11961 gnd.n4085 gnd.n3759 9.3005
R11962 gnd.n4089 gnd.n4086 9.3005
R11963 gnd.n4088 gnd.n4087 9.3005
R11964 gnd.n3733 gnd.n3732 9.3005
R11965 gnd.n4114 gnd.n4113 9.3005
R11966 gnd.n4115 gnd.n3731 9.3005
R11967 gnd.n4125 gnd.n4116 9.3005
R11968 gnd.n4124 gnd.n4117 9.3005
R11969 gnd.n4123 gnd.n4118 9.3005
R11970 gnd.n4121 gnd.n4120 9.3005
R11971 gnd.n4119 gnd.n3703 9.3005
R11972 gnd.n3701 gnd.n3700 9.3005
R11973 gnd.n4173 gnd.n4172 9.3005
R11974 gnd.n4174 gnd.n3699 9.3005
R11975 gnd.n4176 gnd.n4175 9.3005
R11976 gnd.n3519 gnd.n3518 9.3005
R11977 gnd.n4209 gnd.n4208 9.3005
R11978 gnd.n4210 gnd.n3517 9.3005
R11979 gnd.n4214 gnd.n4211 9.3005
R11980 gnd.n4213 gnd.n4212 9.3005
R11981 gnd.n3495 gnd.n3494 9.3005
R11982 gnd.n4240 gnd.n4239 9.3005
R11983 gnd.n4241 gnd.n3493 9.3005
R11984 gnd.n4245 gnd.n4242 9.3005
R11985 gnd.n4244 gnd.n4243 9.3005
R11986 gnd.n3469 gnd.n3468 9.3005
R11987 gnd.n4271 gnd.n4270 9.3005
R11988 gnd.n4272 gnd.n3467 9.3005
R11989 gnd.n4276 gnd.n4273 9.3005
R11990 gnd.n4275 gnd.n4274 9.3005
R11991 gnd.n3444 gnd.n3443 9.3005
R11992 gnd.n4302 gnd.n4301 9.3005
R11993 gnd.n4303 gnd.n3442 9.3005
R11994 gnd.n4307 gnd.n4304 9.3005
R11995 gnd.n4306 gnd.n4305 9.3005
R11996 gnd.n3419 gnd.n3418 9.3005
R11997 gnd.n4333 gnd.n4332 9.3005
R11998 gnd.n4334 gnd.n3417 9.3005
R11999 gnd.n4338 gnd.n4335 9.3005
R12000 gnd.n4337 gnd.n4336 9.3005
R12001 gnd.n3393 gnd.n3392 9.3005
R12002 gnd.n4364 gnd.n4363 9.3005
R12003 gnd.n4365 gnd.n3391 9.3005
R12004 gnd.n4369 gnd.n4366 9.3005
R12005 gnd.n4368 gnd.n4367 9.3005
R12006 gnd.n3368 gnd.n3367 9.3005
R12007 gnd.n4650 gnd.n4649 9.3005
R12008 gnd.n4651 gnd.n3366 9.3005
R12009 gnd.n4655 gnd.n4652 9.3005
R12010 gnd.n4654 gnd.n4653 9.3005
R12011 gnd.n4058 gnd.n4055 9.3005
R12012 gnd.n3840 gnd.n3799 9.3005
R12013 gnd.n3835 gnd.n3834 9.3005
R12014 gnd.n3833 gnd.n3800 9.3005
R12015 gnd.n3832 gnd.n3831 9.3005
R12016 gnd.n3828 gnd.n3801 9.3005
R12017 gnd.n3825 gnd.n3824 9.3005
R12018 gnd.n3823 gnd.n3802 9.3005
R12019 gnd.n3822 gnd.n3821 9.3005
R12020 gnd.n3818 gnd.n3803 9.3005
R12021 gnd.n3815 gnd.n3814 9.3005
R12022 gnd.n3813 gnd.n3804 9.3005
R12023 gnd.n3812 gnd.n3811 9.3005
R12024 gnd.n3808 gnd.n3806 9.3005
R12025 gnd.n3805 gnd.n3785 9.3005
R12026 gnd.n4052 gnd.n3784 9.3005
R12027 gnd.n4054 gnd.n4053 9.3005
R12028 gnd.n3842 gnd.n3841 9.3005
R12029 gnd.n4065 gnd.n3771 9.3005
R12030 gnd.n4072 gnd.n3772 9.3005
R12031 gnd.n4074 gnd.n4073 9.3005
R12032 gnd.n4075 gnd.n3752 9.3005
R12033 gnd.n4094 gnd.n4093 9.3005
R12034 gnd.n4096 gnd.n3744 9.3005
R12035 gnd.n4103 gnd.n3746 9.3005
R12036 gnd.n4104 gnd.n3741 9.3005
R12037 gnd.n4106 gnd.n4105 9.3005
R12038 gnd.n3742 gnd.n3727 9.3005
R12039 gnd.n3725 gnd.n3723 9.3005
R12040 gnd.n4132 gnd.n4131 9.3005
R12041 gnd.n3708 gnd.n3707 9.3005
R12042 gnd.n4165 gnd.n4153 9.3005
R12043 gnd.n4164 gnd.n4155 9.3005
R12044 gnd.n4163 gnd.n4156 9.3005
R12045 gnd.n4158 gnd.n4157 9.3005
R12046 gnd.n3691 gnd.n3528 9.3005
R12047 gnd.n4197 gnd.n3529 9.3005
R12048 gnd.n4199 gnd.n4198 9.3005
R12049 gnd.n4200 gnd.n3512 9.3005
R12050 gnd.n4219 gnd.n4218 9.3005
R12051 gnd.n4221 gnd.n3505 9.3005
R12052 gnd.n4228 gnd.n3506 9.3005
R12053 gnd.n4230 gnd.n4229 9.3005
R12054 gnd.n4231 gnd.n3487 9.3005
R12055 gnd.n4250 gnd.n4249 9.3005
R12056 gnd.n4252 gnd.n3479 9.3005
R12057 gnd.n4259 gnd.n3480 9.3005
R12058 gnd.n4261 gnd.n4260 9.3005
R12059 gnd.n4262 gnd.n3460 9.3005
R12060 gnd.n4281 gnd.n4280 9.3005
R12061 gnd.n4283 gnd.n3453 9.3005
R12062 gnd.n4290 gnd.n3454 9.3005
R12063 gnd.n4292 gnd.n4291 9.3005
R12064 gnd.n4293 gnd.n3436 9.3005
R12065 gnd.n4312 gnd.n4311 9.3005
R12066 gnd.n4314 gnd.n3429 9.3005
R12067 gnd.n4321 gnd.n3430 9.3005
R12068 gnd.n4323 gnd.n4322 9.3005
R12069 gnd.n4324 gnd.n3410 9.3005
R12070 gnd.n4343 gnd.n4342 9.3005
R12071 gnd.n4345 gnd.n3403 9.3005
R12072 gnd.n4352 gnd.n3404 9.3005
R12073 gnd.n4354 gnd.n4353 9.3005
R12074 gnd.n4355 gnd.n3385 9.3005
R12075 gnd.n4374 gnd.n4373 9.3005
R12076 gnd.n4376 gnd.n3377 9.3005
R12077 gnd.n4639 gnd.n3378 9.3005
R12078 gnd.n4641 gnd.n4640 9.3005
R12079 gnd.n4642 gnd.n3359 9.3005
R12080 gnd.n4660 gnd.n4659 9.3005
R12081 gnd.n3360 gnd.n2029 9.3005
R12082 gnd.n4063 gnd.n4062 9.3005
R12083 gnd.n4716 gnd.n2030 9.3005
R12084 gnd.n4715 gnd.n2032 9.3005
R12085 gnd.n4712 gnd.n2033 9.3005
R12086 gnd.n4711 gnd.n2034 9.3005
R12087 gnd.n4708 gnd.n2035 9.3005
R12088 gnd.n4707 gnd.n2036 9.3005
R12089 gnd.n4704 gnd.n2037 9.3005
R12090 gnd.n4703 gnd.n2038 9.3005
R12091 gnd.n4700 gnd.n2039 9.3005
R12092 gnd.n4699 gnd.n2040 9.3005
R12093 gnd.n4696 gnd.n2041 9.3005
R12094 gnd.n4695 gnd.n2042 9.3005
R12095 gnd.n4692 gnd.n2043 9.3005
R12096 gnd.n4691 gnd.n2044 9.3005
R12097 gnd.n4688 gnd.n2045 9.3005
R12098 gnd.n4687 gnd.n2046 9.3005
R12099 gnd.n4684 gnd.n2047 9.3005
R12100 gnd.n4683 gnd.n2048 9.3005
R12101 gnd.n4680 gnd.n2049 9.3005
R12102 gnd.n4679 gnd.n2050 9.3005
R12103 gnd.n4676 gnd.n2051 9.3005
R12104 gnd.n4675 gnd.n2052 9.3005
R12105 gnd.n4672 gnd.n2056 9.3005
R12106 gnd.n4671 gnd.n2057 9.3005
R12107 gnd.n4668 gnd.n2058 9.3005
R12108 gnd.n4667 gnd.n2059 9.3005
R12109 gnd.n4718 gnd.n4717 9.3005
R12110 gnd.n3609 gnd.n3535 9.3005
R12111 gnd.n3607 gnd.n3536 9.3005
R12112 gnd.n3606 gnd.n3537 9.3005
R12113 gnd.n3603 gnd.n3538 9.3005
R12114 gnd.n3602 gnd.n3539 9.3005
R12115 gnd.n3601 gnd.n3540 9.3005
R12116 gnd.n3599 gnd.n3541 9.3005
R12117 gnd.n3598 gnd.n3542 9.3005
R12118 gnd.n3595 gnd.n3543 9.3005
R12119 gnd.n3594 gnd.n3544 9.3005
R12120 gnd.n3593 gnd.n3545 9.3005
R12121 gnd.n3591 gnd.n3546 9.3005
R12122 gnd.n3590 gnd.n3547 9.3005
R12123 gnd.n3585 gnd.n3548 9.3005
R12124 gnd.n3584 gnd.n3549 9.3005
R12125 gnd.n3583 gnd.n3550 9.3005
R12126 gnd.n3581 gnd.n3551 9.3005
R12127 gnd.n3580 gnd.n3552 9.3005
R12128 gnd.n3577 gnd.n3553 9.3005
R12129 gnd.n3576 gnd.n3554 9.3005
R12130 gnd.n3575 gnd.n3555 9.3005
R12131 gnd.n3573 gnd.n3556 9.3005
R12132 gnd.n3572 gnd.n3557 9.3005
R12133 gnd.n3569 gnd.n3558 9.3005
R12134 gnd.n3568 gnd.n3559 9.3005
R12135 gnd.n3567 gnd.n3560 9.3005
R12136 gnd.n3565 gnd.n3561 9.3005
R12137 gnd.n3564 gnd.n3563 9.3005
R12138 gnd.n3562 gnd.n2061 9.3005
R12139 gnd.n3973 gnd.n3972 9.3005
R12140 gnd.n3863 gnd.n3862 9.3005
R12141 gnd.n3987 gnd.n3986 9.3005
R12142 gnd.n3988 gnd.n3861 9.3005
R12143 gnd.n3990 gnd.n3989 9.3005
R12144 gnd.n3851 gnd.n3850 9.3005
R12145 gnd.n4003 gnd.n4002 9.3005
R12146 gnd.n4004 gnd.n3849 9.3005
R12147 gnd.n4036 gnd.n4005 9.3005
R12148 gnd.n4035 gnd.n4006 9.3005
R12149 gnd.n4034 gnd.n4007 9.3005
R12150 gnd.n4033 gnd.n4008 9.3005
R12151 gnd.n4030 gnd.n4009 9.3005
R12152 gnd.n4029 gnd.n4010 9.3005
R12153 gnd.n4028 gnd.n4011 9.3005
R12154 gnd.n4026 gnd.n4012 9.3005
R12155 gnd.n4025 gnd.n4013 9.3005
R12156 gnd.n4022 gnd.n4014 9.3005
R12157 gnd.n4021 gnd.n4015 9.3005
R12158 gnd.n4020 gnd.n4016 9.3005
R12159 gnd.n4018 gnd.n4017 9.3005
R12160 gnd.n3716 gnd.n3715 9.3005
R12161 gnd.n4140 gnd.n4139 9.3005
R12162 gnd.n4141 gnd.n3714 9.3005
R12163 gnd.n4145 gnd.n4142 9.3005
R12164 gnd.n4144 gnd.n4143 9.3005
R12165 gnd.n3679 gnd.n3678 9.3005
R12166 gnd.n4188 gnd.n4187 9.3005
R12167 gnd.n3971 gnd.n3872 9.3005
R12168 gnd.n3874 gnd.n3873 9.3005
R12169 gnd.n3918 gnd.n3916 9.3005
R12170 gnd.n3919 gnd.n3915 9.3005
R12171 gnd.n3922 gnd.n3911 9.3005
R12172 gnd.n3923 gnd.n3910 9.3005
R12173 gnd.n3926 gnd.n3909 9.3005
R12174 gnd.n3927 gnd.n3908 9.3005
R12175 gnd.n3930 gnd.n3907 9.3005
R12176 gnd.n3931 gnd.n3906 9.3005
R12177 gnd.n3934 gnd.n3905 9.3005
R12178 gnd.n3935 gnd.n3904 9.3005
R12179 gnd.n3938 gnd.n3903 9.3005
R12180 gnd.n3939 gnd.n3902 9.3005
R12181 gnd.n3942 gnd.n3901 9.3005
R12182 gnd.n3943 gnd.n3900 9.3005
R12183 gnd.n3946 gnd.n3899 9.3005
R12184 gnd.n3947 gnd.n3898 9.3005
R12185 gnd.n3950 gnd.n3897 9.3005
R12186 gnd.n3951 gnd.n3896 9.3005
R12187 gnd.n3954 gnd.n3895 9.3005
R12188 gnd.n3955 gnd.n3894 9.3005
R12189 gnd.n3958 gnd.n3893 9.3005
R12190 gnd.n3960 gnd.n3892 9.3005
R12191 gnd.n3961 gnd.n3891 9.3005
R12192 gnd.n3962 gnd.n3890 9.3005
R12193 gnd.n3963 gnd.n3889 9.3005
R12194 gnd.n3970 gnd.n3969 9.3005
R12195 gnd.n3979 gnd.n3978 9.3005
R12196 gnd.n3980 gnd.n3866 9.3005
R12197 gnd.n3982 gnd.n3981 9.3005
R12198 gnd.n3857 gnd.n3856 9.3005
R12199 gnd.n3995 gnd.n3994 9.3005
R12200 gnd.n3996 gnd.n3855 9.3005
R12201 gnd.n3998 gnd.n3997 9.3005
R12202 gnd.n3844 gnd.n3843 9.3005
R12203 gnd.n4041 gnd.n4040 9.3005
R12204 gnd.n4042 gnd.n3798 9.3005
R12205 gnd.n4046 gnd.n4044 9.3005
R12206 gnd.n4045 gnd.n3777 9.3005
R12207 gnd.n4064 gnd.n3776 9.3005
R12208 gnd.n4067 gnd.n4066 9.3005
R12209 gnd.n3770 gnd.n3769 9.3005
R12210 gnd.n4078 gnd.n4076 9.3005
R12211 gnd.n4077 gnd.n3751 9.3005
R12212 gnd.n4095 gnd.n3750 9.3005
R12213 gnd.n4098 gnd.n4097 9.3005
R12214 gnd.n3745 gnd.n3740 9.3005
R12215 gnd.n4108 gnd.n4107 9.3005
R12216 gnd.n3743 gnd.n3721 9.3005
R12217 gnd.n4135 gnd.n3722 9.3005
R12218 gnd.n4134 gnd.n4133 9.3005
R12219 gnd.n3724 gnd.n3709 9.3005
R12220 gnd.n4152 gnd.n4151 9.3005
R12221 gnd.n4154 gnd.n3687 9.3005
R12222 gnd.n4183 gnd.n3688 9.3005
R12223 gnd.n4182 gnd.n3689 9.3005
R12224 gnd.n4181 gnd.n3690 9.3005
R12225 gnd.n3693 gnd.n3692 9.3005
R12226 gnd.n3527 gnd.n3526 9.3005
R12227 gnd.n4203 gnd.n4201 9.3005
R12228 gnd.n4202 gnd.n3511 9.3005
R12229 gnd.n4220 gnd.n3510 9.3005
R12230 gnd.n4223 gnd.n4222 9.3005
R12231 gnd.n3504 gnd.n3503 9.3005
R12232 gnd.n4234 gnd.n4232 9.3005
R12233 gnd.n4233 gnd.n3486 9.3005
R12234 gnd.n4251 gnd.n3485 9.3005
R12235 gnd.n4254 gnd.n4253 9.3005
R12236 gnd.n3478 gnd.n3477 9.3005
R12237 gnd.n4265 gnd.n4263 9.3005
R12238 gnd.n4264 gnd.n3459 9.3005
R12239 gnd.n4282 gnd.n3458 9.3005
R12240 gnd.n4285 gnd.n4284 9.3005
R12241 gnd.n3452 gnd.n3451 9.3005
R12242 gnd.n4296 gnd.n4294 9.3005
R12243 gnd.n4295 gnd.n3435 9.3005
R12244 gnd.n4313 gnd.n3434 9.3005
R12245 gnd.n4316 gnd.n4315 9.3005
R12246 gnd.n3428 gnd.n3427 9.3005
R12247 gnd.n4327 gnd.n4325 9.3005
R12248 gnd.n4326 gnd.n3409 9.3005
R12249 gnd.n4344 gnd.n3408 9.3005
R12250 gnd.n4347 gnd.n4346 9.3005
R12251 gnd.n3402 gnd.n3401 9.3005
R12252 gnd.n4358 gnd.n4356 9.3005
R12253 gnd.n4357 gnd.n3384 9.3005
R12254 gnd.n4375 gnd.n3383 9.3005
R12255 gnd.n4634 gnd.n4633 9.3005
R12256 gnd.n3376 gnd.n3375 9.3005
R12257 gnd.n4644 gnd.n4643 9.3005
R12258 gnd.n3358 gnd.n3357 9.3005
R12259 gnd.n4662 gnd.n4661 9.3005
R12260 gnd.n3868 gnd.n3867 9.3005
R12261 gnd.n3139 gnd.n3138 9.3005
R12262 gnd.n3137 gnd.n2191 9.3005
R12263 gnd.n3136 gnd.n3135 9.3005
R12264 gnd.n2193 gnd.n2192 9.3005
R12265 gnd.n3129 gnd.n2197 9.3005
R12266 gnd.n3128 gnd.n2198 9.3005
R12267 gnd.n3127 gnd.n2199 9.3005
R12268 gnd.n2204 gnd.n2200 9.3005
R12269 gnd.n3121 gnd.n2205 9.3005
R12270 gnd.n3120 gnd.n2206 9.3005
R12271 gnd.n3119 gnd.n2207 9.3005
R12272 gnd.n2212 gnd.n2208 9.3005
R12273 gnd.n3113 gnd.n2213 9.3005
R12274 gnd.n3112 gnd.n2214 9.3005
R12275 gnd.n3111 gnd.n2215 9.3005
R12276 gnd.n2220 gnd.n2216 9.3005
R12277 gnd.n3105 gnd.n2221 9.3005
R12278 gnd.n3104 gnd.n2222 9.3005
R12279 gnd.n3103 gnd.n2223 9.3005
R12280 gnd.n2228 gnd.n2224 9.3005
R12281 gnd.n3097 gnd.n2229 9.3005
R12282 gnd.n3096 gnd.n2230 9.3005
R12283 gnd.n3095 gnd.n2231 9.3005
R12284 gnd.n2236 gnd.n2232 9.3005
R12285 gnd.n3089 gnd.n2237 9.3005
R12286 gnd.n3088 gnd.n2238 9.3005
R12287 gnd.n3087 gnd.n2239 9.3005
R12288 gnd.n2244 gnd.n2240 9.3005
R12289 gnd.n3081 gnd.n2245 9.3005
R12290 gnd.n3080 gnd.n2246 9.3005
R12291 gnd.n3079 gnd.n2247 9.3005
R12292 gnd.n2252 gnd.n2248 9.3005
R12293 gnd.n3073 gnd.n2253 9.3005
R12294 gnd.n3072 gnd.n2254 9.3005
R12295 gnd.n3071 gnd.n2255 9.3005
R12296 gnd.n2260 gnd.n2256 9.3005
R12297 gnd.n3065 gnd.n2261 9.3005
R12298 gnd.n3064 gnd.n2262 9.3005
R12299 gnd.n3063 gnd.n2263 9.3005
R12300 gnd.n2268 gnd.n2264 9.3005
R12301 gnd.n3057 gnd.n2269 9.3005
R12302 gnd.n3056 gnd.n2270 9.3005
R12303 gnd.n3055 gnd.n2271 9.3005
R12304 gnd.n2276 gnd.n2272 9.3005
R12305 gnd.n3049 gnd.n2277 9.3005
R12306 gnd.n3048 gnd.n2278 9.3005
R12307 gnd.n3047 gnd.n2279 9.3005
R12308 gnd.n2284 gnd.n2280 9.3005
R12309 gnd.n3041 gnd.n2285 9.3005
R12310 gnd.n3040 gnd.n2286 9.3005
R12311 gnd.n3039 gnd.n2287 9.3005
R12312 gnd.n2292 gnd.n2288 9.3005
R12313 gnd.n3033 gnd.n2293 9.3005
R12314 gnd.n3032 gnd.n2294 9.3005
R12315 gnd.n3031 gnd.n2295 9.3005
R12316 gnd.n2300 gnd.n2296 9.3005
R12317 gnd.n3025 gnd.n2301 9.3005
R12318 gnd.n3024 gnd.n2302 9.3005
R12319 gnd.n3023 gnd.n2303 9.3005
R12320 gnd.n2308 gnd.n2304 9.3005
R12321 gnd.n3017 gnd.n2309 9.3005
R12322 gnd.n3016 gnd.n2310 9.3005
R12323 gnd.n3015 gnd.n2311 9.3005
R12324 gnd.n2316 gnd.n2312 9.3005
R12325 gnd.n3009 gnd.n2317 9.3005
R12326 gnd.n3008 gnd.n2318 9.3005
R12327 gnd.n3007 gnd.n2319 9.3005
R12328 gnd.n2324 gnd.n2320 9.3005
R12329 gnd.n3001 gnd.n2325 9.3005
R12330 gnd.n3000 gnd.n2326 9.3005
R12331 gnd.n2999 gnd.n2327 9.3005
R12332 gnd.n2332 gnd.n2328 9.3005
R12333 gnd.n2993 gnd.n2333 9.3005
R12334 gnd.n2992 gnd.n2334 9.3005
R12335 gnd.n2991 gnd.n2335 9.3005
R12336 gnd.n2340 gnd.n2336 9.3005
R12337 gnd.n2985 gnd.n2341 9.3005
R12338 gnd.n2984 gnd.n2342 9.3005
R12339 gnd.n2983 gnd.n2343 9.3005
R12340 gnd.n2348 gnd.n2344 9.3005
R12341 gnd.n2977 gnd.n2349 9.3005
R12342 gnd.n2976 gnd.n2350 9.3005
R12343 gnd.n2975 gnd.n2351 9.3005
R12344 gnd.n2356 gnd.n2352 9.3005
R12345 gnd.n2969 gnd.n2357 9.3005
R12346 gnd.n2968 gnd.n2358 9.3005
R12347 gnd.n2967 gnd.n2359 9.3005
R12348 gnd.n2364 gnd.n2360 9.3005
R12349 gnd.n2961 gnd.n2365 9.3005
R12350 gnd.n2960 gnd.n2366 9.3005
R12351 gnd.n2959 gnd.n2367 9.3005
R12352 gnd.n2372 gnd.n2368 9.3005
R12353 gnd.n2953 gnd.n2373 9.3005
R12354 gnd.n2952 gnd.n2374 9.3005
R12355 gnd.n2951 gnd.n2375 9.3005
R12356 gnd.n2380 gnd.n2376 9.3005
R12357 gnd.n2945 gnd.n2381 9.3005
R12358 gnd.n2944 gnd.n2382 9.3005
R12359 gnd.n2943 gnd.n2383 9.3005
R12360 gnd.n2388 gnd.n2384 9.3005
R12361 gnd.n2937 gnd.n2389 9.3005
R12362 gnd.n2936 gnd.n2390 9.3005
R12363 gnd.n2935 gnd.n2391 9.3005
R12364 gnd.n2396 gnd.n2392 9.3005
R12365 gnd.n2929 gnd.n2397 9.3005
R12366 gnd.n2928 gnd.n2398 9.3005
R12367 gnd.n2927 gnd.n2399 9.3005
R12368 gnd.n2404 gnd.n2400 9.3005
R12369 gnd.n2921 gnd.n2405 9.3005
R12370 gnd.n2920 gnd.n2406 9.3005
R12371 gnd.n2919 gnd.n2407 9.3005
R12372 gnd.n2412 gnd.n2408 9.3005
R12373 gnd.n2913 gnd.n2413 9.3005
R12374 gnd.n2912 gnd.n2414 9.3005
R12375 gnd.n2911 gnd.n2415 9.3005
R12376 gnd.n2420 gnd.n2416 9.3005
R12377 gnd.n2905 gnd.n2421 9.3005
R12378 gnd.n2904 gnd.n2422 9.3005
R12379 gnd.n2903 gnd.n2423 9.3005
R12380 gnd.n2428 gnd.n2424 9.3005
R12381 gnd.n2897 gnd.n2429 9.3005
R12382 gnd.n2896 gnd.n2430 9.3005
R12383 gnd.n2895 gnd.n2431 9.3005
R12384 gnd.n2436 gnd.n2432 9.3005
R12385 gnd.n2889 gnd.n2437 9.3005
R12386 gnd.n2888 gnd.n2438 9.3005
R12387 gnd.n2887 gnd.n2439 9.3005
R12388 gnd.n2444 gnd.n2440 9.3005
R12389 gnd.n2881 gnd.n2445 9.3005
R12390 gnd.n2880 gnd.n2446 9.3005
R12391 gnd.n2879 gnd.n2447 9.3005
R12392 gnd.n2452 gnd.n2448 9.3005
R12393 gnd.n2873 gnd.n2453 9.3005
R12394 gnd.n2872 gnd.n2454 9.3005
R12395 gnd.n2871 gnd.n2455 9.3005
R12396 gnd.n2460 gnd.n2456 9.3005
R12397 gnd.n2865 gnd.n2461 9.3005
R12398 gnd.n2864 gnd.n2462 9.3005
R12399 gnd.n2863 gnd.n2463 9.3005
R12400 gnd.n2468 gnd.n2464 9.3005
R12401 gnd.n2857 gnd.n2469 9.3005
R12402 gnd.n2856 gnd.n2470 9.3005
R12403 gnd.n2855 gnd.n2471 9.3005
R12404 gnd.n2476 gnd.n2472 9.3005
R12405 gnd.n2849 gnd.n2477 9.3005
R12406 gnd.n2848 gnd.n2478 9.3005
R12407 gnd.n2847 gnd.n2479 9.3005
R12408 gnd.n2484 gnd.n2480 9.3005
R12409 gnd.n2841 gnd.n2485 9.3005
R12410 gnd.n2840 gnd.n2486 9.3005
R12411 gnd.n2839 gnd.n2487 9.3005
R12412 gnd.n2492 gnd.n2488 9.3005
R12413 gnd.n2833 gnd.n2493 9.3005
R12414 gnd.n2832 gnd.n2494 9.3005
R12415 gnd.n2831 gnd.n2495 9.3005
R12416 gnd.n2825 gnd.n2824 9.3005
R12417 gnd.n2823 gnd.n2500 9.3005
R12418 gnd.n2822 gnd.n2821 9.3005
R12419 gnd.n2503 gnd.n2502 9.3005
R12420 gnd.n2815 gnd.n2507 9.3005
R12421 gnd.n2814 gnd.n2508 9.3005
R12422 gnd.n2813 gnd.n2509 9.3005
R12423 gnd.n2514 gnd.n2510 9.3005
R12424 gnd.n2807 gnd.n2515 9.3005
R12425 gnd.n2806 gnd.n2516 9.3005
R12426 gnd.n2805 gnd.n2517 9.3005
R12427 gnd.n2522 gnd.n2518 9.3005
R12428 gnd.n2799 gnd.n2523 9.3005
R12429 gnd.n2798 gnd.n2524 9.3005
R12430 gnd.n2797 gnd.n2525 9.3005
R12431 gnd.n2530 gnd.n2526 9.3005
R12432 gnd.n2791 gnd.n2531 9.3005
R12433 gnd.n2790 gnd.n2532 9.3005
R12434 gnd.n2789 gnd.n2533 9.3005
R12435 gnd.n2538 gnd.n2534 9.3005
R12436 gnd.n2783 gnd.n2539 9.3005
R12437 gnd.n2782 gnd.n2540 9.3005
R12438 gnd.n2781 gnd.n2541 9.3005
R12439 gnd.n2546 gnd.n2542 9.3005
R12440 gnd.n2775 gnd.n2547 9.3005
R12441 gnd.n2774 gnd.n2548 9.3005
R12442 gnd.n2773 gnd.n2549 9.3005
R12443 gnd.n2554 gnd.n2550 9.3005
R12444 gnd.n2767 gnd.n2555 9.3005
R12445 gnd.n2766 gnd.n2556 9.3005
R12446 gnd.n2765 gnd.n2557 9.3005
R12447 gnd.n2562 gnd.n2558 9.3005
R12448 gnd.n2759 gnd.n2563 9.3005
R12449 gnd.n2758 gnd.n2564 9.3005
R12450 gnd.n2757 gnd.n2565 9.3005
R12451 gnd.n2570 gnd.n2566 9.3005
R12452 gnd.n2751 gnd.n2571 9.3005
R12453 gnd.n2750 gnd.n2572 9.3005
R12454 gnd.n2749 gnd.n2573 9.3005
R12455 gnd.n2578 gnd.n2574 9.3005
R12456 gnd.n2743 gnd.n2579 9.3005
R12457 gnd.n2742 gnd.n2580 9.3005
R12458 gnd.n2741 gnd.n2581 9.3005
R12459 gnd.n2586 gnd.n2582 9.3005
R12460 gnd.n2735 gnd.n2587 9.3005
R12461 gnd.n2734 gnd.n2588 9.3005
R12462 gnd.n2733 gnd.n2589 9.3005
R12463 gnd.n2594 gnd.n2590 9.3005
R12464 gnd.n2727 gnd.n2595 9.3005
R12465 gnd.n2726 gnd.n2596 9.3005
R12466 gnd.n2725 gnd.n2597 9.3005
R12467 gnd.n2602 gnd.n2598 9.3005
R12468 gnd.n2719 gnd.n2603 9.3005
R12469 gnd.n2718 gnd.n2604 9.3005
R12470 gnd.n2717 gnd.n2605 9.3005
R12471 gnd.n2610 gnd.n2606 9.3005
R12472 gnd.n2711 gnd.n2611 9.3005
R12473 gnd.n2710 gnd.n2612 9.3005
R12474 gnd.n2709 gnd.n2613 9.3005
R12475 gnd.n2618 gnd.n2614 9.3005
R12476 gnd.n2703 gnd.n2619 9.3005
R12477 gnd.n2702 gnd.n2620 9.3005
R12478 gnd.n2701 gnd.n2621 9.3005
R12479 gnd.n2626 gnd.n2622 9.3005
R12480 gnd.n2695 gnd.n2627 9.3005
R12481 gnd.n2694 gnd.n2628 9.3005
R12482 gnd.n2693 gnd.n2629 9.3005
R12483 gnd.n2634 gnd.n2630 9.3005
R12484 gnd.n2687 gnd.n2635 9.3005
R12485 gnd.n2686 gnd.n2636 9.3005
R12486 gnd.n2685 gnd.n2637 9.3005
R12487 gnd.n2642 gnd.n2638 9.3005
R12488 gnd.n2679 gnd.n2643 9.3005
R12489 gnd.n2678 gnd.n2644 9.3005
R12490 gnd.n2677 gnd.n2645 9.3005
R12491 gnd.n2650 gnd.n2646 9.3005
R12492 gnd.n2671 gnd.n2651 9.3005
R12493 gnd.n2670 gnd.n2652 9.3005
R12494 gnd.n2669 gnd.n2653 9.3005
R12495 gnd.n2659 gnd.n2654 9.3005
R12496 gnd.n2663 gnd.n2660 9.3005
R12497 gnd.n2662 gnd.n2661 9.3005
R12498 gnd.n345 gnd.n344 9.3005
R12499 gnd.n7219 gnd.n7218 9.3005
R12500 gnd.n2501 gnd.n2499 9.3005
R12501 gnd.n7567 gnd.n130 9.3005
R12502 gnd.n7566 gnd.n132 9.3005
R12503 gnd.n136 gnd.n133 9.3005
R12504 gnd.n7561 gnd.n137 9.3005
R12505 gnd.n7560 gnd.n138 9.3005
R12506 gnd.n7559 gnd.n139 9.3005
R12507 gnd.n143 gnd.n140 9.3005
R12508 gnd.n7554 gnd.n144 9.3005
R12509 gnd.n7553 gnd.n145 9.3005
R12510 gnd.n7552 gnd.n146 9.3005
R12511 gnd.n150 gnd.n147 9.3005
R12512 gnd.n7547 gnd.n151 9.3005
R12513 gnd.n7546 gnd.n152 9.3005
R12514 gnd.n7545 gnd.n153 9.3005
R12515 gnd.n157 gnd.n154 9.3005
R12516 gnd.n7540 gnd.n158 9.3005
R12517 gnd.n7539 gnd.n159 9.3005
R12518 gnd.n7535 gnd.n160 9.3005
R12519 gnd.n164 gnd.n161 9.3005
R12520 gnd.n7530 gnd.n165 9.3005
R12521 gnd.n7529 gnd.n166 9.3005
R12522 gnd.n7528 gnd.n167 9.3005
R12523 gnd.n171 gnd.n168 9.3005
R12524 gnd.n7523 gnd.n172 9.3005
R12525 gnd.n7522 gnd.n173 9.3005
R12526 gnd.n7521 gnd.n174 9.3005
R12527 gnd.n178 gnd.n175 9.3005
R12528 gnd.n7516 gnd.n179 9.3005
R12529 gnd.n7515 gnd.n180 9.3005
R12530 gnd.n7514 gnd.n181 9.3005
R12531 gnd.n185 gnd.n182 9.3005
R12532 gnd.n7509 gnd.n186 9.3005
R12533 gnd.n7508 gnd.n187 9.3005
R12534 gnd.n7507 gnd.n188 9.3005
R12535 gnd.n192 gnd.n189 9.3005
R12536 gnd.n7502 gnd.n193 9.3005
R12537 gnd.n7501 gnd.n7500 9.3005
R12538 gnd.n7499 gnd.n196 9.3005
R12539 gnd.n7569 gnd.n7568 9.3005
R12540 gnd.n6844 gnd.n6843 9.3005
R12541 gnd.n6848 gnd.n6845 9.3005
R12542 gnd.n6849 gnd.n6842 9.3005
R12543 gnd.n6853 gnd.n6852 9.3005
R12544 gnd.n6854 gnd.n6841 9.3005
R12545 gnd.n6863 gnd.n6855 9.3005
R12546 gnd.n6862 gnd.n6856 9.3005
R12547 gnd.n6861 gnd.n6858 9.3005
R12548 gnd.n6857 gnd.n596 9.3005
R12549 gnd.n6888 gnd.n597 9.3005
R12550 gnd.n6889 gnd.n595 9.3005
R12551 gnd.n6893 gnd.n6892 9.3005
R12552 gnd.n6894 gnd.n594 9.3005
R12553 gnd.n6902 gnd.n6895 9.3005
R12554 gnd.n6901 gnd.n6896 9.3005
R12555 gnd.n6900 gnd.n6897 9.3005
R12556 gnd.n587 gnd.n586 9.3005
R12557 gnd.n6920 gnd.n6919 9.3005
R12558 gnd.n6921 gnd.n585 9.3005
R12559 gnd.n6936 gnd.n6922 9.3005
R12560 gnd.n6935 gnd.n6923 9.3005
R12561 gnd.n6934 gnd.n6924 9.3005
R12562 gnd.n6933 gnd.n6925 9.3005
R12563 gnd.n6932 gnd.n6926 9.3005
R12564 gnd.n6929 gnd.n6928 9.3005
R12565 gnd.n6927 gnd.n357 9.3005
R12566 gnd.n7193 gnd.n356 9.3005
R12567 gnd.n7195 gnd.n7194 9.3005
R12568 gnd.n7196 gnd.n355 9.3005
R12569 gnd.n7200 gnd.n7197 9.3005
R12570 gnd.n7199 gnd.n7198 9.3005
R12571 gnd.n334 gnd.n333 9.3005
R12572 gnd.n7231 gnd.n7230 9.3005
R12573 gnd.n7232 gnd.n332 9.3005
R12574 gnd.n7299 gnd.n7233 9.3005
R12575 gnd.n7298 gnd.n7234 9.3005
R12576 gnd.n7297 gnd.n7235 9.3005
R12577 gnd.n7295 gnd.n7236 9.3005
R12578 gnd.n7294 gnd.n7237 9.3005
R12579 gnd.n7292 gnd.n7238 9.3005
R12580 gnd.n7291 gnd.n7239 9.3005
R12581 gnd.n7289 gnd.n7240 9.3005
R12582 gnd.n7288 gnd.n7241 9.3005
R12583 gnd.n7286 gnd.n7242 9.3005
R12584 gnd.n7285 gnd.n7243 9.3005
R12585 gnd.n7283 gnd.n7244 9.3005
R12586 gnd.n7282 gnd.n7245 9.3005
R12587 gnd.n7280 gnd.n7246 9.3005
R12588 gnd.n7279 gnd.n7247 9.3005
R12589 gnd.n7277 gnd.n7248 9.3005
R12590 gnd.n7276 gnd.n7249 9.3005
R12591 gnd.n7274 gnd.n7250 9.3005
R12592 gnd.n7273 gnd.n7251 9.3005
R12593 gnd.n7271 gnd.n7252 9.3005
R12594 gnd.n7270 gnd.n7253 9.3005
R12595 gnd.n7268 gnd.n7254 9.3005
R12596 gnd.n7267 gnd.n7255 9.3005
R12597 gnd.n7265 gnd.n7256 9.3005
R12598 gnd.n7264 gnd.n7257 9.3005
R12599 gnd.n7262 gnd.n7258 9.3005
R12600 gnd.n7261 gnd.n7260 9.3005
R12601 gnd.n7259 gnd.n200 9.3005
R12602 gnd.n7496 gnd.n199 9.3005
R12603 gnd.n7498 gnd.n7497 9.3005
R12604 gnd.n563 gnd.n562 9.3005
R12605 gnd.n6981 gnd.n6980 9.3005
R12606 gnd.n6982 gnd.n556 9.3005
R12607 gnd.n6985 gnd.n555 9.3005
R12608 gnd.n6986 gnd.n554 9.3005
R12609 gnd.n6989 gnd.n553 9.3005
R12610 gnd.n6990 gnd.n552 9.3005
R12611 gnd.n6993 gnd.n551 9.3005
R12612 gnd.n6994 gnd.n550 9.3005
R12613 gnd.n6997 gnd.n549 9.3005
R12614 gnd.n6998 gnd.n548 9.3005
R12615 gnd.n7001 gnd.n547 9.3005
R12616 gnd.n7002 gnd.n546 9.3005
R12617 gnd.n7005 gnd.n545 9.3005
R12618 gnd.n7006 gnd.n544 9.3005
R12619 gnd.n7009 gnd.n543 9.3005
R12620 gnd.n7010 gnd.n542 9.3005
R12621 gnd.n7013 gnd.n541 9.3005
R12622 gnd.n7014 gnd.n540 9.3005
R12623 gnd.n7017 gnd.n539 9.3005
R12624 gnd.n7019 gnd.n533 9.3005
R12625 gnd.n7022 gnd.n532 9.3005
R12626 gnd.n7023 gnd.n531 9.3005
R12627 gnd.n7026 gnd.n530 9.3005
R12628 gnd.n7027 gnd.n529 9.3005
R12629 gnd.n7030 gnd.n528 9.3005
R12630 gnd.n7031 gnd.n527 9.3005
R12631 gnd.n7034 gnd.n526 9.3005
R12632 gnd.n7035 gnd.n525 9.3005
R12633 gnd.n7038 gnd.n524 9.3005
R12634 gnd.n7039 gnd.n523 9.3005
R12635 gnd.n7042 gnd.n522 9.3005
R12636 gnd.n7043 gnd.n521 9.3005
R12637 gnd.n7044 gnd.n520 9.3005
R12638 gnd.n487 gnd.n486 9.3005
R12639 gnd.n7050 gnd.n7049 9.3005
R12640 gnd.n6979 gnd.n561 9.3005
R12641 gnd.n6978 gnd.n6977 9.3005
R12642 gnd.n7053 gnd.n7052 9.3005
R12643 gnd.n469 gnd.n468 9.3005
R12644 gnd.n7066 gnd.n7065 9.3005
R12645 gnd.n7067 gnd.n467 9.3005
R12646 gnd.n7069 gnd.n7068 9.3005
R12647 gnd.n452 gnd.n451 9.3005
R12648 gnd.n7082 gnd.n7081 9.3005
R12649 gnd.n7083 gnd.n450 9.3005
R12650 gnd.n7085 gnd.n7084 9.3005
R12651 gnd.n435 gnd.n434 9.3005
R12652 gnd.n7098 gnd.n7097 9.3005
R12653 gnd.n7099 gnd.n433 9.3005
R12654 gnd.n7101 gnd.n7100 9.3005
R12655 gnd.n418 gnd.n417 9.3005
R12656 gnd.n7114 gnd.n7113 9.3005
R12657 gnd.n7115 gnd.n416 9.3005
R12658 gnd.n7117 gnd.n7116 9.3005
R12659 gnd.n399 gnd.n398 9.3005
R12660 gnd.n7133 gnd.n7132 9.3005
R12661 gnd.n7134 gnd.n397 9.3005
R12662 gnd.n7136 gnd.n7135 9.3005
R12663 gnd.n367 gnd.n366 9.3005
R12664 gnd.n7184 gnd.n7183 9.3005
R12665 gnd.n7185 gnd.n365 9.3005
R12666 gnd.n7187 gnd.n7186 9.3005
R12667 gnd.n7188 gnd.n299 9.3005
R12668 gnd.n7327 gnd.n7326 9.3005
R12669 gnd.n284 gnd.n283 9.3005
R12670 gnd.n7340 gnd.n7339 9.3005
R12671 gnd.n7341 gnd.n282 9.3005
R12672 gnd.n7343 gnd.n7342 9.3005
R12673 gnd.n270 gnd.n269 9.3005
R12674 gnd.n7356 gnd.n7355 9.3005
R12675 gnd.n7357 gnd.n268 9.3005
R12676 gnd.n7359 gnd.n7358 9.3005
R12677 gnd.n254 gnd.n253 9.3005
R12678 gnd.n7372 gnd.n7371 9.3005
R12679 gnd.n7373 gnd.n252 9.3005
R12680 gnd.n7375 gnd.n7374 9.3005
R12681 gnd.n240 gnd.n239 9.3005
R12682 gnd.n7388 gnd.n7387 9.3005
R12683 gnd.n7389 gnd.n238 9.3005
R12684 gnd.n7391 gnd.n7390 9.3005
R12685 gnd.n223 gnd.n222 9.3005
R12686 gnd.n7404 gnd.n7403 9.3005
R12687 gnd.n7405 gnd.n221 9.3005
R12688 gnd.n7407 gnd.n7406 9.3005
R12689 gnd.n207 gnd.n206 9.3005
R12690 gnd.n7488 gnd.n7487 9.3005
R12691 gnd.n7489 gnd.n205 9.3005
R12692 gnd.n7491 gnd.n7490 9.3005
R12693 gnd.n129 gnd.n128 9.3005
R12694 gnd.n7571 gnd.n7570 9.3005
R12695 gnd.n7051 gnd.n485 9.3005
R12696 gnd.n7325 gnd.n298 9.3005
R12697 gnd.n7148 gnd.n346 9.3005
R12698 gnd.n7215 gnd.n347 9.3005
R12699 gnd.n7217 gnd.n7216 9.3005
R12700 gnd.n5433 gnd.n1803 9.3005
R12701 gnd.n5258 gnd.n1804 9.3005
R12702 gnd.n5260 gnd.n5259 9.3005
R12703 gnd.n5261 gnd.n5257 9.3005
R12704 gnd.n5273 gnd.n5262 9.3005
R12705 gnd.n5272 gnd.n5263 9.3005
R12706 gnd.n5271 gnd.n5264 9.3005
R12707 gnd.n5268 gnd.n5265 9.3005
R12708 gnd.n5267 gnd.n5266 9.3005
R12709 gnd.n1848 gnd.n1847 9.3005
R12710 gnd.n5300 gnd.n5299 9.3005
R12711 gnd.n5301 gnd.n1846 9.3005
R12712 gnd.n5313 gnd.n5302 9.3005
R12713 gnd.n5312 gnd.n5303 9.3005
R12714 gnd.n5311 gnd.n5304 9.3005
R12715 gnd.n5308 gnd.n5305 9.3005
R12716 gnd.n5307 gnd.n5306 9.3005
R12717 gnd.n1838 gnd.n1837 9.3005
R12718 gnd.n5339 gnd.n5338 9.3005
R12719 gnd.n5340 gnd.n1836 9.3005
R12720 gnd.n5370 gnd.n5341 9.3005
R12721 gnd.n5369 gnd.n5342 9.3005
R12722 gnd.n5368 gnd.n5343 9.3005
R12723 gnd.n5346 gnd.n5344 9.3005
R12724 gnd.n5364 gnd.n5347 9.3005
R12725 gnd.n5363 gnd.n5348 9.3005
R12726 gnd.n5362 gnd.n5349 9.3005
R12727 gnd.n5353 gnd.n5350 9.3005
R12728 gnd.n5357 gnd.n5354 9.3005
R12729 gnd.n5356 gnd.n5355 9.3005
R12730 gnd.n1316 gnd.n1315 9.3005
R12731 gnd.n5812 gnd.n5811 9.3005
R12732 gnd.n5813 gnd.n1314 9.3005
R12733 gnd.n5815 gnd.n5814 9.3005
R12734 gnd.n1302 gnd.n1301 9.3005
R12735 gnd.n5828 gnd.n5827 9.3005
R12736 gnd.n5829 gnd.n1300 9.3005
R12737 gnd.n5833 gnd.n5830 9.3005
R12738 gnd.n5832 gnd.n5831 9.3005
R12739 gnd.n1260 gnd.n1259 9.3005
R12740 gnd.n5986 gnd.n5985 9.3005
R12741 gnd.n5987 gnd.n1258 9.3005
R12742 gnd.n5989 gnd.n5988 9.3005
R12743 gnd.n1245 gnd.n1244 9.3005
R12744 gnd.n6002 gnd.n6001 9.3005
R12745 gnd.n6003 gnd.n1243 9.3005
R12746 gnd.n6005 gnd.n6004 9.3005
R12747 gnd.n1229 gnd.n1228 9.3005
R12748 gnd.n6018 gnd.n6017 9.3005
R12749 gnd.n6019 gnd.n1227 9.3005
R12750 gnd.n6021 gnd.n6020 9.3005
R12751 gnd.n1214 gnd.n1213 9.3005
R12752 gnd.n6033 gnd.n6032 9.3005
R12753 gnd.n6034 gnd.n1212 9.3005
R12754 gnd.n6038 gnd.n6035 9.3005
R12755 gnd.n6037 gnd.n6036 9.3005
R12756 gnd.n1107 gnd.n1106 9.3005
R12757 gnd.n6128 gnd.n6127 9.3005
R12758 gnd.n6129 gnd.n1105 9.3005
R12759 gnd.n6131 gnd.n6130 9.3005
R12760 gnd.n1091 gnd.n1090 9.3005
R12761 gnd.n6144 gnd.n6143 9.3005
R12762 gnd.n6145 gnd.n1089 9.3005
R12763 gnd.n6147 gnd.n6146 9.3005
R12764 gnd.n1076 gnd.n1075 9.3005
R12765 gnd.n6160 gnd.n6159 9.3005
R12766 gnd.n6161 gnd.n1074 9.3005
R12767 gnd.n6163 gnd.n6162 9.3005
R12768 gnd.n1063 gnd.n1062 9.3005
R12769 gnd.n6176 gnd.n6175 9.3005
R12770 gnd.n6177 gnd.n1061 9.3005
R12771 gnd.n6181 gnd.n6178 9.3005
R12772 gnd.n6180 gnd.n6179 9.3005
R12773 gnd.n1020 gnd.n1019 9.3005
R12774 gnd.n6433 gnd.n6432 9.3005
R12775 gnd.n6434 gnd.n1018 9.3005
R12776 gnd.n6436 gnd.n6435 9.3005
R12777 gnd.n1004 gnd.n1003 9.3005
R12778 gnd.n6449 gnd.n6448 9.3005
R12779 gnd.n6450 gnd.n1002 9.3005
R12780 gnd.n6452 gnd.n6451 9.3005
R12781 gnd.n988 gnd.n987 9.3005
R12782 gnd.n6465 gnd.n6464 9.3005
R12783 gnd.n6466 gnd.n986 9.3005
R12784 gnd.n6468 gnd.n6467 9.3005
R12785 gnd.n974 gnd.n973 9.3005
R12786 gnd.n6481 gnd.n6480 9.3005
R12787 gnd.n6482 gnd.n972 9.3005
R12788 gnd.n6484 gnd.n6483 9.3005
R12789 gnd.n959 gnd.n958 9.3005
R12790 gnd.n6497 gnd.n6496 9.3005
R12791 gnd.n6498 gnd.n957 9.3005
R12792 gnd.n6500 gnd.n6499 9.3005
R12793 gnd.n943 gnd.n942 9.3005
R12794 gnd.n6513 gnd.n6512 9.3005
R12795 gnd.n6514 gnd.n941 9.3005
R12796 gnd.n6516 gnd.n6515 9.3005
R12797 gnd.n926 gnd.n925 9.3005
R12798 gnd.n6535 gnd.n6534 9.3005
R12799 gnd.n6536 gnd.n924 9.3005
R12800 gnd.n6540 gnd.n6537 9.3005
R12801 gnd.n6539 gnd.n6538 9.3005
R12802 gnd.n886 gnd.n885 9.3005
R12803 gnd.n6593 gnd.n6592 9.3005
R12804 gnd.n6594 gnd.n884 9.3005
R12805 gnd.n6598 gnd.n6595 9.3005
R12806 gnd.n6597 gnd.n6596 9.3005
R12807 gnd.n659 gnd.n658 9.3005
R12808 gnd.n6784 gnd.n6783 9.3005
R12809 gnd.n6785 gnd.n657 9.3005
R12810 gnd.n6787 gnd.n6786 9.3005
R12811 gnd.n644 gnd.n643 9.3005
R12812 gnd.n6801 gnd.n6800 9.3005
R12813 gnd.n6802 gnd.n642 9.3005
R12814 gnd.n6806 gnd.n6803 9.3005
R12815 gnd.n6805 gnd.n6804 9.3005
R12816 gnd.n614 gnd.n613 9.3005
R12817 gnd.n6820 gnd.n6819 9.3005
R12818 gnd.n6821 gnd.n612 9.3005
R12819 gnd.n6823 gnd.n6822 9.3005
R12820 gnd.n610 gnd.n609 9.3005
R12821 gnd.n6828 gnd.n6827 9.3005
R12822 gnd.n6829 gnd.n608 9.3005
R12823 gnd.n6831 gnd.n6830 9.3005
R12824 gnd.n606 gnd.n605 9.3005
R12825 gnd.n6836 gnd.n6835 9.3005
R12826 gnd.n6837 gnd.n604 9.3005
R12827 gnd.n6839 gnd.n6838 9.3005
R12828 gnd.n602 gnd.n601 9.3005
R12829 gnd.n6870 gnd.n6869 9.3005
R12830 gnd.n6871 gnd.n600 9.3005
R12831 gnd.n6883 gnd.n6872 9.3005
R12832 gnd.n6882 gnd.n6873 9.3005
R12833 gnd.n6881 gnd.n6874 9.3005
R12834 gnd.n6878 gnd.n6875 9.3005
R12835 gnd.n6877 gnd.n6876 9.3005
R12836 gnd.n592 gnd.n591 9.3005
R12837 gnd.n6909 gnd.n6908 9.3005
R12838 gnd.n6910 gnd.n590 9.3005
R12839 gnd.n6914 gnd.n6911 9.3005
R12840 gnd.n6913 gnd.n6912 9.3005
R12841 gnd.n392 gnd.n391 9.3005
R12842 gnd.n7142 gnd.n7141 9.3005
R12843 gnd.n7143 gnd.n390 9.3005
R12844 gnd.n7156 gnd.n7144 9.3005
R12845 gnd.n7155 gnd.n7145 9.3005
R12846 gnd.n7154 gnd.n7146 9.3005
R12847 gnd.n7151 gnd.n7147 9.3005
R12848 gnd.n7150 gnd.n7149 9.3005
R12849 gnd.n5210 gnd.n5209 9.3005
R12850 gnd.n4870 gnd.n4827 9.3005
R12851 gnd.n4869 gnd.n4828 9.3005
R12852 gnd.n4868 gnd.n4829 9.3005
R12853 gnd.n4866 gnd.n4830 9.3005
R12854 gnd.n4865 gnd.n4831 9.3005
R12855 gnd.n4863 gnd.n4832 9.3005
R12856 gnd.n4862 gnd.n4833 9.3005
R12857 gnd.n4860 gnd.n4834 9.3005
R12858 gnd.n4859 gnd.n4835 9.3005
R12859 gnd.n4857 gnd.n4836 9.3005
R12860 gnd.n4856 gnd.n4837 9.3005
R12861 gnd.n4854 gnd.n4838 9.3005
R12862 gnd.n4853 gnd.n4839 9.3005
R12863 gnd.n4851 gnd.n4840 9.3005
R12864 gnd.n4850 gnd.n4841 9.3005
R12865 gnd.n4848 gnd.n4842 9.3005
R12866 gnd.n4847 gnd.n4843 9.3005
R12867 gnd.n4845 gnd.n4844 9.3005
R12868 gnd.n1906 gnd.n1905 9.3005
R12869 gnd.n5163 gnd.n5162 9.3005
R12870 gnd.n5164 gnd.n1904 9.3005
R12871 gnd.n5171 gnd.n5165 9.3005
R12872 gnd.n5170 gnd.n5166 9.3005
R12873 gnd.n5169 gnd.n5167 9.3005
R12874 gnd.n1871 gnd.n1870 9.3005
R12875 gnd.n5202 gnd.n5201 9.3005
R12876 gnd.n5203 gnd.n1869 9.3005
R12877 gnd.n5215 gnd.n5204 9.3005
R12878 gnd.n5214 gnd.n5205 9.3005
R12879 gnd.n5213 gnd.n5206 9.3005
R12880 gnd.n5211 gnd.n5207 9.3005
R12881 gnd.n4826 gnd.n4759 9.3005
R12882 gnd.n4819 gnd.n4818 9.3005
R12883 gnd.n4817 gnd.n4765 9.3005
R12884 gnd.n4816 gnd.n4815 9.3005
R12885 gnd.n4767 gnd.n4766 9.3005
R12886 gnd.n4809 gnd.n4808 9.3005
R12887 gnd.n4807 gnd.n4769 9.3005
R12888 gnd.n4806 gnd.n4805 9.3005
R12889 gnd.n4771 gnd.n4770 9.3005
R12890 gnd.n4799 gnd.n4798 9.3005
R12891 gnd.n4797 gnd.n4773 9.3005
R12892 gnd.n4796 gnd.n4795 9.3005
R12893 gnd.n4775 gnd.n4774 9.3005
R12894 gnd.n4789 gnd.n4788 9.3005
R12895 gnd.n4787 gnd.n4777 9.3005
R12896 gnd.n4786 gnd.n4785 9.3005
R12897 gnd.n4780 gnd.n4778 9.3005
R12898 gnd.n4779 gnd.n1986 9.3005
R12899 gnd.n4763 gnd.n4760 9.3005
R12900 gnd.n4825 gnd.n4824 9.3005
R12901 gnd.n5074 gnd.n1985 9.3005
R12902 gnd.n5076 gnd.n5075 9.3005
R12903 gnd.n1972 gnd.n1971 9.3005
R12904 gnd.n5089 gnd.n5088 9.3005
R12905 gnd.n5090 gnd.n1970 9.3005
R12906 gnd.n5092 gnd.n5091 9.3005
R12907 gnd.n1955 gnd.n1954 9.3005
R12908 gnd.n5105 gnd.n5104 9.3005
R12909 gnd.n5106 gnd.n1953 9.3005
R12910 gnd.n5108 gnd.n5107 9.3005
R12911 gnd.n1940 gnd.n1939 9.3005
R12912 gnd.n5121 gnd.n5120 9.3005
R12913 gnd.n5122 gnd.n1938 9.3005
R12914 gnd.n5124 gnd.n5123 9.3005
R12915 gnd.n1923 gnd.n1922 9.3005
R12916 gnd.n5137 gnd.n5136 9.3005
R12917 gnd.n5138 gnd.n1921 9.3005
R12918 gnd.n5148 gnd.n5139 9.3005
R12919 gnd.n5147 gnd.n5140 9.3005
R12920 gnd.n5146 gnd.n5141 9.3005
R12921 gnd.n5145 gnd.n5143 9.3005
R12922 gnd.n5142 gnd.n1887 9.3005
R12923 gnd.n5188 gnd.n1888 9.3005
R12924 gnd.n5187 gnd.n1889 9.3005
R12925 gnd.n5186 gnd.n1890 9.3005
R12926 gnd.n1896 gnd.n1891 9.3005
R12927 gnd.n1895 gnd.n1893 9.3005
R12928 gnd.n1892 gnd.n1778 9.3005
R12929 gnd.n5459 gnd.n1779 9.3005
R12930 gnd.n5458 gnd.n1780 9.3005
R12931 gnd.n5457 gnd.n1781 9.3005
R12932 gnd.n1861 gnd.n1782 9.3005
R12933 gnd.n5445 gnd.n1792 9.3005
R12934 gnd.n5444 gnd.n1793 9.3005
R12935 gnd.n5443 gnd.n1794 9.3005
R12936 gnd.n1756 gnd.n1755 9.3005
R12937 gnd.n5472 gnd.n5471 9.3005
R12938 gnd.n5473 gnd.n1754 9.3005
R12939 gnd.n5475 gnd.n5474 9.3005
R12940 gnd.n1740 gnd.n1739 9.3005
R12941 gnd.n5488 gnd.n5487 9.3005
R12942 gnd.n5489 gnd.n1738 9.3005
R12943 gnd.n5491 gnd.n5490 9.3005
R12944 gnd.n1722 gnd.n1721 9.3005
R12945 gnd.n5504 gnd.n5503 9.3005
R12946 gnd.n5505 gnd.n1720 9.3005
R12947 gnd.n5507 gnd.n5506 9.3005
R12948 gnd.n1706 gnd.n1705 9.3005
R12949 gnd.n5520 gnd.n5519 9.3005
R12950 gnd.n5521 gnd.n1704 9.3005
R12951 gnd.n5523 gnd.n5522 9.3005
R12952 gnd.n1688 gnd.n1687 9.3005
R12953 gnd.n5536 gnd.n5535 9.3005
R12954 gnd.n5537 gnd.n1686 9.3005
R12955 gnd.n5539 gnd.n5538 9.3005
R12956 gnd.n1672 gnd.n1671 9.3005
R12957 gnd.n5552 gnd.n5551 9.3005
R12958 gnd.n5553 gnd.n1670 9.3005
R12959 gnd.n5555 gnd.n5554 9.3005
R12960 gnd.n1653 gnd.n1652 9.3005
R12961 gnd.n5570 gnd.n5569 9.3005
R12962 gnd.n5571 gnd.n1651 9.3005
R12963 gnd.n5692 gnd.n5572 9.3005
R12964 gnd.n5691 gnd.n5690 9.3005
R12965 gnd.n5073 gnd.n5072 9.3005
R12966 gnd.n1608 gnd.n1386 9.3005
R12967 gnd.n5742 gnd.n1385 9.3005
R12968 gnd.n5743 gnd.n1384 9.3005
R12969 gnd.n5744 gnd.n1383 9.3005
R12970 gnd.n1382 gnd.n1379 9.3005
R12971 gnd.n5749 gnd.n1378 9.3005
R12972 gnd.n5750 gnd.n1377 9.3005
R12973 gnd.n5751 gnd.n1376 9.3005
R12974 gnd.n1375 gnd.n1372 9.3005
R12975 gnd.n5756 gnd.n1371 9.3005
R12976 gnd.n5757 gnd.n1370 9.3005
R12977 gnd.n5758 gnd.n1369 9.3005
R12978 gnd.n1368 gnd.n1365 9.3005
R12979 gnd.n1367 gnd.n1363 9.3005
R12980 gnd.n5765 gnd.n1362 9.3005
R12981 gnd.n5767 gnd.n5766 9.3005
R12982 gnd.n5734 gnd.n1611 9.3005
R12983 gnd.n5733 gnd.n1612 9.3005
R12984 gnd.n1616 gnd.n1613 9.3005
R12985 gnd.n5728 gnd.n1617 9.3005
R12986 gnd.n5727 gnd.n1618 9.3005
R12987 gnd.n5726 gnd.n1619 9.3005
R12988 gnd.n1623 gnd.n1620 9.3005
R12989 gnd.n5721 gnd.n1624 9.3005
R12990 gnd.n5720 gnd.n1625 9.3005
R12991 gnd.n5719 gnd.n1626 9.3005
R12992 gnd.n1630 gnd.n1627 9.3005
R12993 gnd.n5714 gnd.n1631 9.3005
R12994 gnd.n5713 gnd.n1632 9.3005
R12995 gnd.n5712 gnd.n1633 9.3005
R12996 gnd.n1637 gnd.n1634 9.3005
R12997 gnd.n5707 gnd.n1638 9.3005
R12998 gnd.n5706 gnd.n1639 9.3005
R12999 gnd.n5705 gnd.n1640 9.3005
R13000 gnd.n1645 gnd.n1643 9.3005
R13001 gnd.n5700 gnd.n5699 9.3005
R13002 gnd.n5735 gnd.n1610 9.3005
R13003 gnd.n4985 gnd.n4935 9.3005
R13004 gnd.n4984 gnd.n4937 9.3005
R13005 gnd.n4983 gnd.n4938 9.3005
R13006 gnd.n4981 gnd.n4939 9.3005
R13007 gnd.n4980 gnd.n4940 9.3005
R13008 gnd.n4978 gnd.n4941 9.3005
R13009 gnd.n4977 gnd.n4942 9.3005
R13010 gnd.n4975 gnd.n4943 9.3005
R13011 gnd.n4974 gnd.n4944 9.3005
R13012 gnd.n4972 gnd.n4945 9.3005
R13013 gnd.n4971 gnd.n4946 9.3005
R13014 gnd.n4969 gnd.n4947 9.3005
R13015 gnd.n4968 gnd.n4948 9.3005
R13016 gnd.n4966 gnd.n4949 9.3005
R13017 gnd.n4965 gnd.n4950 9.3005
R13018 gnd.n4963 gnd.n4951 9.3005
R13019 gnd.n4962 gnd.n4952 9.3005
R13020 gnd.n4960 gnd.n4953 9.3005
R13021 gnd.n4959 gnd.n4954 9.3005
R13022 gnd.n4957 gnd.n4956 9.3005
R13023 gnd.n4955 gnd.n1900 9.3005
R13024 gnd.n5175 gnd.n1899 9.3005
R13025 gnd.n5177 gnd.n5176 9.3005
R13026 gnd.n5178 gnd.n1898 9.3005
R13027 gnd.n5182 gnd.n5179 9.3005
R13028 gnd.n5181 gnd.n5180 9.3005
R13029 gnd.n1865 gnd.n1864 9.3005
R13030 gnd.n5220 gnd.n5219 9.3005
R13031 gnd.n5221 gnd.n1863 9.3005
R13032 gnd.n5224 gnd.n5222 9.3005
R13033 gnd.n5225 gnd.n1862 9.3005
R13034 gnd.n5228 gnd.n5227 9.3005
R13035 gnd.n5229 gnd.n1860 9.3005
R13036 gnd.n5231 gnd.n5230 9.3005
R13037 gnd.n1856 gnd.n1855 9.3005
R13038 gnd.n5244 gnd.n5243 9.3005
R13039 gnd.n5245 gnd.n1854 9.3005
R13040 gnd.n5247 gnd.n5246 9.3005
R13041 gnd.n5248 gnd.n1853 9.3005
R13042 gnd.n5252 gnd.n5251 9.3005
R13043 gnd.n5253 gnd.n1852 9.3005
R13044 gnd.n5278 gnd.n5254 9.3005
R13045 gnd.n5279 gnd.n1851 9.3005
R13046 gnd.n5283 gnd.n5282 9.3005
R13047 gnd.n5284 gnd.n1850 9.3005
R13048 gnd.n5293 gnd.n5285 9.3005
R13049 gnd.n5292 gnd.n5286 9.3005
R13050 gnd.n5291 gnd.n5288 9.3005
R13051 gnd.n5287 gnd.n1842 9.3005
R13052 gnd.n5318 gnd.n1843 9.3005
R13053 gnd.n5319 gnd.n1841 9.3005
R13054 gnd.n5323 gnd.n5322 9.3005
R13055 gnd.n5324 gnd.n1840 9.3005
R13056 gnd.n5332 gnd.n5325 9.3005
R13057 gnd.n5331 gnd.n5326 9.3005
R13058 gnd.n5330 gnd.n5327 9.3005
R13059 gnd.n1833 gnd.n1832 9.3005
R13060 gnd.n5376 gnd.n5375 9.3005
R13061 gnd.n5377 gnd.n1831 9.3005
R13062 gnd.n5382 gnd.n5378 9.3005
R13063 gnd.n5381 gnd.n5380 9.3005
R13064 gnd.n5379 gnd.n1647 9.3005
R13065 gnd.n5696 gnd.n1646 9.3005
R13066 gnd.n5698 gnd.n5697 9.3005
R13067 gnd.n4987 gnd.n4986 9.3005
R13068 gnd.n4995 gnd.n4994 9.3005
R13069 gnd.n4996 gnd.n4929 9.3005
R13070 gnd.n4997 gnd.n4928 9.3005
R13071 gnd.n4927 gnd.n4925 9.3005
R13072 gnd.n5003 gnd.n4924 9.3005
R13073 gnd.n5004 gnd.n4923 9.3005
R13074 gnd.n5005 gnd.n4922 9.3005
R13075 gnd.n4921 gnd.n4919 9.3005
R13076 gnd.n5011 gnd.n4918 9.3005
R13077 gnd.n5012 gnd.n4917 9.3005
R13078 gnd.n5013 gnd.n4916 9.3005
R13079 gnd.n4915 gnd.n4913 9.3005
R13080 gnd.n5019 gnd.n4912 9.3005
R13081 gnd.n5020 gnd.n4911 9.3005
R13082 gnd.n5021 gnd.n4910 9.3005
R13083 gnd.n4909 gnd.n4907 9.3005
R13084 gnd.n5027 gnd.n4906 9.3005
R13085 gnd.n5028 gnd.n4905 9.3005
R13086 gnd.n5029 gnd.n4904 9.3005
R13087 gnd.n4903 gnd.n4898 9.3005
R13088 gnd.n5035 gnd.n4897 9.3005
R13089 gnd.n5036 gnd.n4896 9.3005
R13090 gnd.n5037 gnd.n4895 9.3005
R13091 gnd.n4894 gnd.n4892 9.3005
R13092 gnd.n5043 gnd.n4891 9.3005
R13093 gnd.n5044 gnd.n4890 9.3005
R13094 gnd.n5045 gnd.n4889 9.3005
R13095 gnd.n4888 gnd.n4886 9.3005
R13096 gnd.n5051 gnd.n4885 9.3005
R13097 gnd.n5052 gnd.n4884 9.3005
R13098 gnd.n5053 gnd.n4883 9.3005
R13099 gnd.n4882 gnd.n4880 9.3005
R13100 gnd.n5058 gnd.n4879 9.3005
R13101 gnd.n5059 gnd.n4878 9.3005
R13102 gnd.n4877 gnd.n4875 9.3005
R13103 gnd.n5064 gnd.n4874 9.3005
R13104 gnd.n5066 gnd.n5065 9.3005
R13105 gnd.n4993 gnd.n4934 9.3005
R13106 gnd.n4992 gnd.n4991 9.3005
R13107 gnd.n1980 gnd.n1979 9.3005
R13108 gnd.n5081 gnd.n5080 9.3005
R13109 gnd.n5082 gnd.n1978 9.3005
R13110 gnd.n5084 gnd.n5083 9.3005
R13111 gnd.n1964 gnd.n1963 9.3005
R13112 gnd.n5097 gnd.n5096 9.3005
R13113 gnd.n5098 gnd.n1962 9.3005
R13114 gnd.n5100 gnd.n5099 9.3005
R13115 gnd.n1948 gnd.n1947 9.3005
R13116 gnd.n5113 gnd.n5112 9.3005
R13117 gnd.n5114 gnd.n1946 9.3005
R13118 gnd.n5116 gnd.n5115 9.3005
R13119 gnd.n1932 gnd.n1931 9.3005
R13120 gnd.n5129 gnd.n5128 9.3005
R13121 gnd.n5130 gnd.n1930 9.3005
R13122 gnd.n5132 gnd.n5131 9.3005
R13123 gnd.n1915 gnd.n1914 9.3005
R13124 gnd.n5153 gnd.n5152 9.3005
R13125 gnd.n5154 gnd.n1913 9.3005
R13126 gnd.n5158 gnd.n5155 9.3005
R13127 gnd.n5157 gnd.n5156 9.3005
R13128 gnd.n1879 gnd.n1878 9.3005
R13129 gnd.n5193 gnd.n5192 9.3005
R13130 gnd.n5194 gnd.n1877 9.3005
R13131 gnd.n5196 gnd.n5195 9.3005
R13132 gnd.n5197 gnd.n1764 9.3005
R13133 gnd.n1748 gnd.n1747 9.3005
R13134 gnd.n5480 gnd.n5479 9.3005
R13135 gnd.n5481 gnd.n1746 9.3005
R13136 gnd.n5483 gnd.n5482 9.3005
R13137 gnd.n1731 gnd.n1730 9.3005
R13138 gnd.n5496 gnd.n5495 9.3005
R13139 gnd.n5497 gnd.n1729 9.3005
R13140 gnd.n5499 gnd.n5498 9.3005
R13141 gnd.n1714 gnd.n1713 9.3005
R13142 gnd.n5512 gnd.n5511 9.3005
R13143 gnd.n5513 gnd.n1712 9.3005
R13144 gnd.n5515 gnd.n5514 9.3005
R13145 gnd.n1697 gnd.n1696 9.3005
R13146 gnd.n5528 gnd.n5527 9.3005
R13147 gnd.n5529 gnd.n1695 9.3005
R13148 gnd.n5531 gnd.n5530 9.3005
R13149 gnd.n1680 gnd.n1679 9.3005
R13150 gnd.n5544 gnd.n5543 9.3005
R13151 gnd.n5545 gnd.n1678 9.3005
R13152 gnd.n5547 gnd.n5546 9.3005
R13153 gnd.n1663 gnd.n1662 9.3005
R13154 gnd.n5560 gnd.n5559 9.3005
R13155 gnd.n5561 gnd.n1661 9.3005
R13156 gnd.n5565 gnd.n5562 9.3005
R13157 gnd.n5564 gnd.n5563 9.3005
R13158 gnd.n1361 gnd.n1360 9.3005
R13159 gnd.n5769 gnd.n5768 9.3005
R13160 gnd.n5068 gnd.n5067 9.3005
R13161 gnd.n5467 gnd.n5466 9.3005
R13162 gnd.n5435 gnd.n1801 9.3005
R13163 gnd.n5434 gnd.n1802 9.3005
R13164 gnd.n3349 gnd.n1800 9.3005
R13165 gnd.n3352 gnd.n3348 9.3005
R13166 gnd.n3347 gnd.n2065 9.3005
R13167 gnd.n3346 gnd.n3345 9.3005
R13168 gnd.n2067 gnd.n2066 9.3005
R13169 gnd.n3339 gnd.n3338 9.3005
R13170 gnd.n3337 gnd.n2071 9.3005
R13171 gnd.n3336 gnd.n3335 9.3005
R13172 gnd.n2073 gnd.n2072 9.3005
R13173 gnd.n3329 gnd.n3328 9.3005
R13174 gnd.n3327 gnd.n2077 9.3005
R13175 gnd.n3326 gnd.n3325 9.3005
R13176 gnd.n2079 gnd.n2078 9.3005
R13177 gnd.n3319 gnd.n3318 9.3005
R13178 gnd.n3317 gnd.n2083 9.3005
R13179 gnd.n3316 gnd.n3315 9.3005
R13180 gnd.n2085 gnd.n2084 9.3005
R13181 gnd.n3309 gnd.n3308 9.3005
R13182 gnd.n3307 gnd.n2089 9.3005
R13183 gnd.n3306 gnd.n3305 9.3005
R13184 gnd.n2091 gnd.n2090 9.3005
R13185 gnd.n3299 gnd.n3298 9.3005
R13186 gnd.n3297 gnd.n2095 9.3005
R13187 gnd.n3296 gnd.n3295 9.3005
R13188 gnd.n2097 gnd.n2096 9.3005
R13189 gnd.n3289 gnd.n3288 9.3005
R13190 gnd.n3287 gnd.n2101 9.3005
R13191 gnd.n3286 gnd.n3285 9.3005
R13192 gnd.n2103 gnd.n2102 9.3005
R13193 gnd.n3279 gnd.n3278 9.3005
R13194 gnd.n3277 gnd.n2107 9.3005
R13195 gnd.n3276 gnd.n3275 9.3005
R13196 gnd.n2109 gnd.n2108 9.3005
R13197 gnd.n3269 gnd.n3268 9.3005
R13198 gnd.n3267 gnd.n2113 9.3005
R13199 gnd.n3266 gnd.n3265 9.3005
R13200 gnd.n2115 gnd.n2114 9.3005
R13201 gnd.n3259 gnd.n3258 9.3005
R13202 gnd.n3257 gnd.n2119 9.3005
R13203 gnd.n3256 gnd.n3255 9.3005
R13204 gnd.n2121 gnd.n2120 9.3005
R13205 gnd.n3249 gnd.n3248 9.3005
R13206 gnd.n3247 gnd.n2125 9.3005
R13207 gnd.n3246 gnd.n3245 9.3005
R13208 gnd.n2127 gnd.n2126 9.3005
R13209 gnd.n3239 gnd.n3238 9.3005
R13210 gnd.n3237 gnd.n2131 9.3005
R13211 gnd.n3236 gnd.n3235 9.3005
R13212 gnd.n2133 gnd.n2132 9.3005
R13213 gnd.n3229 gnd.n3228 9.3005
R13214 gnd.n3227 gnd.n2137 9.3005
R13215 gnd.n3226 gnd.n3225 9.3005
R13216 gnd.n2139 gnd.n2138 9.3005
R13217 gnd.n3219 gnd.n3218 9.3005
R13218 gnd.n3217 gnd.n2143 9.3005
R13219 gnd.n3216 gnd.n3215 9.3005
R13220 gnd.n2145 gnd.n2144 9.3005
R13221 gnd.n3209 gnd.n3208 9.3005
R13222 gnd.n3207 gnd.n2149 9.3005
R13223 gnd.n3206 gnd.n3205 9.3005
R13224 gnd.n2151 gnd.n2150 9.3005
R13225 gnd.n3199 gnd.n3198 9.3005
R13226 gnd.n3197 gnd.n2155 9.3005
R13227 gnd.n3196 gnd.n3195 9.3005
R13228 gnd.n2157 gnd.n2156 9.3005
R13229 gnd.n3189 gnd.n3188 9.3005
R13230 gnd.n3187 gnd.n2161 9.3005
R13231 gnd.n3186 gnd.n3185 9.3005
R13232 gnd.n2163 gnd.n2162 9.3005
R13233 gnd.n3179 gnd.n3178 9.3005
R13234 gnd.n3177 gnd.n2167 9.3005
R13235 gnd.n3176 gnd.n3175 9.3005
R13236 gnd.n2169 gnd.n2168 9.3005
R13237 gnd.n3169 gnd.n3168 9.3005
R13238 gnd.n3167 gnd.n2173 9.3005
R13239 gnd.n3166 gnd.n3165 9.3005
R13240 gnd.n2175 gnd.n2174 9.3005
R13241 gnd.n3159 gnd.n3158 9.3005
R13242 gnd.n3157 gnd.n2179 9.3005
R13243 gnd.n3156 gnd.n3155 9.3005
R13244 gnd.n2181 gnd.n2180 9.3005
R13245 gnd.n3149 gnd.n3148 9.3005
R13246 gnd.n3147 gnd.n2185 9.3005
R13247 gnd.n3146 gnd.n3145 9.3005
R13248 gnd.n2187 gnd.n2186 9.3005
R13249 gnd.n3351 gnd.n3350 9.3005
R13250 gnd.n6618 gnd.n6616 9.3005
R13251 gnd.n6751 gnd.n6750 9.3005
R13252 gnd.n6749 gnd.n6748 9.3005
R13253 gnd.n6635 gnd.n6634 9.3005
R13254 gnd.n6743 gnd.n6742 9.3005
R13255 gnd.n6741 gnd.n6740 9.3005
R13256 gnd.n6643 gnd.n6642 9.3005
R13257 gnd.n6735 gnd.n6734 9.3005
R13258 gnd.n6733 gnd.n6732 9.3005
R13259 gnd.n6655 gnd.n6654 9.3005
R13260 gnd.n6727 gnd.n6726 9.3005
R13261 gnd.n6725 gnd.n6724 9.3005
R13262 gnd.n6663 gnd.n6662 9.3005
R13263 gnd.n6719 gnd.n6718 9.3005
R13264 gnd.n6717 gnd.n6716 9.3005
R13265 gnd.n6675 gnd.n6674 9.3005
R13266 gnd.n6708 gnd.n6707 9.3005
R13267 gnd.n6706 gnd.n6676 9.3005
R13268 gnd.n6757 gnd.n6756 9.3005
R13269 gnd.n6669 gnd.n6668 9.3005
R13270 gnd.n6721 gnd.n6720 9.3005
R13271 gnd.n6723 gnd.n6722 9.3005
R13272 gnd.n6659 gnd.n6658 9.3005
R13273 gnd.n6729 gnd.n6728 9.3005
R13274 gnd.n6731 gnd.n6730 9.3005
R13275 gnd.n6649 gnd.n6648 9.3005
R13276 gnd.n6737 gnd.n6736 9.3005
R13277 gnd.n6739 gnd.n6738 9.3005
R13278 gnd.n6639 gnd.n6638 9.3005
R13279 gnd.n6745 gnd.n6744 9.3005
R13280 gnd.n6747 gnd.n6746 9.3005
R13281 gnd.n6629 gnd.n6628 9.3005
R13282 gnd.n6753 gnd.n6752 9.3005
R13283 gnd.n6755 gnd.n6754 9.3005
R13284 gnd.n6623 gnd.n6617 9.3005
R13285 gnd.n6715 gnd.n6714 9.3005
R13286 gnd.n6710 gnd.n6709 9.3005
R13287 gnd.n6705 gnd.n6704 9.3005
R13288 gnd.n6703 gnd.n6681 9.3005
R13289 gnd.n6702 gnd.n6701 9.3005
R13290 gnd.n6700 gnd.n6682 9.3005
R13291 gnd.n6699 gnd.n6698 9.3005
R13292 gnd.n6697 gnd.n6687 9.3005
R13293 gnd.n6696 gnd.n6695 9.3005
R13294 gnd.n6694 gnd.n6688 9.3005
R13295 gnd.n634 gnd.n633 9.3005
R13296 gnd.n6814 gnd.n6813 9.3005
R13297 gnd.n5821 gnd.n1307 9.3005
R13298 gnd.n5823 gnd.n5822 9.3005
R13299 gnd.n1293 gnd.n1292 9.3005
R13300 gnd.n5838 gnd.n5837 9.3005
R13301 gnd.n5839 gnd.n1290 9.3005
R13302 gnd.n5842 gnd.n5841 9.3005
R13303 gnd.n5840 gnd.n1291 9.3005
R13304 gnd.n1252 gnd.n1251 9.3005
R13305 gnd.n5994 gnd.n5993 9.3005
R13306 gnd.n5995 gnd.n1250 9.3005
R13307 gnd.n5997 gnd.n5996 9.3005
R13308 gnd.n1237 gnd.n1236 9.3005
R13309 gnd.n6010 gnd.n6009 9.3005
R13310 gnd.n6011 gnd.n1235 9.3005
R13311 gnd.n6013 gnd.n6012 9.3005
R13312 gnd.n1222 gnd.n1221 9.3005
R13313 gnd.n6026 gnd.n6025 9.3005
R13314 gnd.n6027 gnd.n1220 9.3005
R13315 gnd.n6029 gnd.n6028 9.3005
R13316 gnd.n1205 gnd.n1204 9.3005
R13317 gnd.n6043 gnd.n6042 9.3005
R13318 gnd.n6044 gnd.n1202 9.3005
R13319 gnd.n6047 gnd.n6046 9.3005
R13320 gnd.n6045 gnd.n1203 9.3005
R13321 gnd.n1099 gnd.n1098 9.3005
R13322 gnd.n6136 gnd.n6135 9.3005
R13323 gnd.n6137 gnd.n1097 9.3005
R13324 gnd.n6139 gnd.n6138 9.3005
R13325 gnd.n1084 gnd.n1083 9.3005
R13326 gnd.n6152 gnd.n6151 9.3005
R13327 gnd.n6153 gnd.n1082 9.3005
R13328 gnd.n6155 gnd.n6154 9.3005
R13329 gnd.n1070 gnd.n1069 9.3005
R13330 gnd.n6168 gnd.n6167 9.3005
R13331 gnd.n6169 gnd.n1068 9.3005
R13332 gnd.n6171 gnd.n6170 9.3005
R13333 gnd.n1054 gnd.n1053 9.3005
R13334 gnd.n6186 gnd.n6185 9.3005
R13335 gnd.n6187 gnd.n1051 9.3005
R13336 gnd.n6190 gnd.n6189 9.3005
R13337 gnd.n6188 gnd.n1052 9.3005
R13338 gnd.n1012 gnd.n1011 9.3005
R13339 gnd.n6441 gnd.n6440 9.3005
R13340 gnd.n6442 gnd.n1010 9.3005
R13341 gnd.n6444 gnd.n6443 9.3005
R13342 gnd.n996 gnd.n995 9.3005
R13343 gnd.n6457 gnd.n6456 9.3005
R13344 gnd.n6458 gnd.n994 9.3005
R13345 gnd.n6460 gnd.n6459 9.3005
R13346 gnd.n981 gnd.n980 9.3005
R13347 gnd.n6473 gnd.n6472 9.3005
R13348 gnd.n6474 gnd.n979 9.3005
R13349 gnd.n6476 gnd.n6475 9.3005
R13350 gnd.n966 gnd.n965 9.3005
R13351 gnd.n6489 gnd.n6488 9.3005
R13352 gnd.n6490 gnd.n964 9.3005
R13353 gnd.n6492 gnd.n6491 9.3005
R13354 gnd.n951 gnd.n950 9.3005
R13355 gnd.n6505 gnd.n6504 9.3005
R13356 gnd.n6506 gnd.n949 9.3005
R13357 gnd.n6508 gnd.n6507 9.3005
R13358 gnd.n935 gnd.n934 9.3005
R13359 gnd.n6520 gnd.n6519 9.3005
R13360 gnd.n6521 gnd.n932 9.3005
R13361 gnd.n6530 gnd.n6529 9.3005
R13362 gnd.n6528 gnd.n933 9.3005
R13363 gnd.n6527 gnd.n6526 9.3005
R13364 gnd.n6525 gnd.n6522 9.3005
R13365 gnd.n895 gnd.n893 9.3005
R13366 gnd.n6588 gnd.n6587 9.3005
R13367 gnd.n6586 gnd.n894 9.3005
R13368 gnd.n6585 gnd.n6584 9.3005
R13369 gnd.n6583 gnd.n896 9.3005
R13370 gnd.n6582 gnd.n6581 9.3005
R13371 gnd.n6580 gnd.n6579 9.3005
R13372 gnd.n652 gnd.n651 9.3005
R13373 gnd.n6792 gnd.n6791 9.3005
R13374 gnd.n6793 gnd.n650 9.3005
R13375 gnd.n6796 gnd.n6795 9.3005
R13376 gnd.n6794 gnd.n636 9.3005
R13377 gnd.n6810 gnd.n635 9.3005
R13378 gnd.n6812 gnd.n6811 9.3005
R13379 gnd.n5820 gnd.n5819 9.3005
R13380 gnd.n5806 gnd.n5805 9.3005
R13381 gnd.n5804 gnd.n1333 9.3005
R13382 gnd.n5803 gnd.n5802 9.3005
R13383 gnd.n5799 gnd.n1335 9.3005
R13384 gnd.n5796 gnd.n5795 9.3005
R13385 gnd.n5794 gnd.n1338 9.3005
R13386 gnd.n5793 gnd.n5792 9.3005
R13387 gnd.n5789 gnd.n1339 9.3005
R13388 gnd.n5786 gnd.n5785 9.3005
R13389 gnd.n1334 gnd.n1308 9.3005
R13390 gnd.n1859 gnd.n1858 9.3005
R13391 gnd.n5236 gnd.n5235 9.3005
R13392 gnd.n5237 gnd.n1857 9.3005
R13393 gnd.n5239 gnd.n5238 9.3005
R13394 gnd.n1809 gnd.n1807 9.3005
R13395 gnd.n5427 gnd.n5426 9.3005
R13396 gnd.n5425 gnd.n1808 9.3005
R13397 gnd.n5424 gnd.n5423 9.3005
R13398 gnd.n5422 gnd.n1810 9.3005
R13399 gnd.n5421 gnd.n5420 9.3005
R13400 gnd.n5419 gnd.n1813 9.3005
R13401 gnd.n5418 gnd.n5417 9.3005
R13402 gnd.n5416 gnd.n1814 9.3005
R13403 gnd.n5415 gnd.n5414 9.3005
R13404 gnd.n5413 gnd.n1817 9.3005
R13405 gnd.n5412 gnd.n5411 9.3005
R13406 gnd.n5410 gnd.n1818 9.3005
R13407 gnd.n5409 gnd.n5408 9.3005
R13408 gnd.n5407 gnd.n1821 9.3005
R13409 gnd.n5406 gnd.n5405 9.3005
R13410 gnd.n5404 gnd.n1822 9.3005
R13411 gnd.n5403 gnd.n5402 9.3005
R13412 gnd.n5401 gnd.n1825 9.3005
R13413 gnd.n5400 gnd.n5399 9.3005
R13414 gnd.n5398 gnd.n1826 9.3005
R13415 gnd.n5397 gnd.n5396 9.3005
R13416 gnd.n5395 gnd.n1829 9.3005
R13417 gnd.n5394 gnd.n5393 9.3005
R13418 gnd.n5392 gnd.n1830 9.3005
R13419 gnd.n5391 gnd.n5390 9.3005
R13420 gnd.n5389 gnd.n5388 9.3005
R13421 gnd.n1353 gnd.n1341 9.3005
R13422 gnd.n5783 gnd.n1340 9.3005
R13423 gnd.n5782 gnd.n5781 9.3005
R13424 gnd.n5778 gnd.n5777 9.3005
R13425 gnd.n1346 gnd.n1343 9.3005
R13426 gnd.n5636 gnd.n5635 9.3005
R13427 gnd.n5638 gnd.n5637 9.3005
R13428 gnd.n5621 gnd.n5620 9.3005
R13429 gnd.n5644 gnd.n5643 9.3005
R13430 gnd.n5646 gnd.n5645 9.3005
R13431 gnd.n5609 gnd.n5608 9.3005
R13432 gnd.n5652 gnd.n5651 9.3005
R13433 gnd.n5654 gnd.n5653 9.3005
R13434 gnd.n5598 gnd.n5597 9.3005
R13435 gnd.n5660 gnd.n5659 9.3005
R13436 gnd.n5662 gnd.n5661 9.3005
R13437 gnd.n5586 gnd.n5585 9.3005
R13438 gnd.n5668 gnd.n5667 9.3005
R13439 gnd.n5670 gnd.n5669 9.3005
R13440 gnd.n5582 gnd.n5574 9.3005
R13441 gnd.n5674 gnd.n5673 9.3005
R13442 gnd.n5672 gnd.n5671 9.3005
R13443 gnd.n5580 gnd.n5579 9.3005
R13444 gnd.n5666 gnd.n5665 9.3005
R13445 gnd.n5664 gnd.n5663 9.3005
R13446 gnd.n5592 gnd.n5591 9.3005
R13447 gnd.n5658 gnd.n5657 9.3005
R13448 gnd.n5656 gnd.n5655 9.3005
R13449 gnd.n5605 gnd.n5604 9.3005
R13450 gnd.n5650 gnd.n5649 9.3005
R13451 gnd.n5648 gnd.n5647 9.3005
R13452 gnd.n5615 gnd.n5614 9.3005
R13453 gnd.n5642 gnd.n5641 9.3005
R13454 gnd.n5640 gnd.n5639 9.3005
R13455 gnd.n5631 gnd.n5630 9.3005
R13456 gnd.n5634 gnd.n1347 9.3005
R13457 gnd.n5776 gnd.n5775 9.3005
R13458 gnd.n5774 gnd.n1342 9.3005
R13459 gnd.n5685 gnd.n5675 9.3005
R13460 gnd.n5684 gnd.n5683 9.3005
R13461 gnd.n5682 gnd.n5679 9.3005
R13462 gnd.n5681 gnd.n5680 9.3005
R13463 gnd.n1285 gnd.n1284 9.3005
R13464 gnd.n5847 gnd.n5846 9.3005
R13465 gnd.n5848 gnd.n1281 9.3005
R13466 gnd.n5850 gnd.n5849 9.3005
R13467 gnd.n5851 gnd.n1280 9.3005
R13468 gnd.n5856 gnd.n5855 9.3005
R13469 gnd.n5857 gnd.n1278 9.3005
R13470 gnd.n5965 gnd.n5964 9.3005
R13471 gnd.n5963 gnd.n1279 9.3005
R13472 gnd.n5962 gnd.n5961 9.3005
R13473 gnd.n5960 gnd.n5858 9.3005
R13474 gnd.n5959 gnd.n5958 9.3005
R13475 gnd.n5957 gnd.n5861 9.3005
R13476 gnd.n5956 gnd.n5955 9.3005
R13477 gnd.n5954 gnd.n5862 9.3005
R13478 gnd.n5953 gnd.n5952 9.3005
R13479 gnd.n5951 gnd.n5950 9.3005
R13480 gnd.n1197 gnd.n1196 9.3005
R13481 gnd.n6052 gnd.n6051 9.3005
R13482 gnd.n6053 gnd.n1193 9.3005
R13483 gnd.n6055 gnd.n6054 9.3005
R13484 gnd.n6056 gnd.n1192 9.3005
R13485 gnd.n6059 gnd.n6058 9.3005
R13486 gnd.n6060 gnd.n1191 9.3005
R13487 gnd.n6062 gnd.n6061 9.3005
R13488 gnd.n6063 gnd.n1190 9.3005
R13489 gnd.n6066 gnd.n6065 9.3005
R13490 gnd.n6067 gnd.n1189 9.3005
R13491 gnd.n6069 gnd.n6068 9.3005
R13492 gnd.n6070 gnd.n1188 9.3005
R13493 gnd.n6073 gnd.n6072 9.3005
R13494 gnd.n6074 gnd.n1186 9.3005
R13495 gnd.n6077 gnd.n6076 9.3005
R13496 gnd.n6075 gnd.n1187 9.3005
R13497 gnd.n1047 gnd.n1046 9.3005
R13498 gnd.n6195 gnd.n6194 9.3005
R13499 gnd.n6196 gnd.n1043 9.3005
R13500 gnd.n6198 gnd.n6197 9.3005
R13501 gnd.n6199 gnd.n1042 9.3005
R13502 gnd.n6202 gnd.n6201 9.3005
R13503 gnd.n6203 gnd.n1040 9.3005
R13504 gnd.n6412 gnd.n6411 9.3005
R13505 gnd.n6410 gnd.n1041 9.3005
R13506 gnd.n6409 gnd.n6408 9.3005
R13507 gnd.n6407 gnd.n6204 9.3005
R13508 gnd.n6406 gnd.n6405 9.3005
R13509 gnd.n6404 gnd.n6207 9.3005
R13510 gnd.n6403 gnd.n6402 9.3005
R13511 gnd.n6401 gnd.n6208 9.3005
R13512 gnd.n6400 gnd.n6399 9.3005
R13513 gnd.n6398 gnd.n6211 9.3005
R13514 gnd.n6397 gnd.n6396 9.3005
R13515 gnd.n6395 gnd.n6212 9.3005
R13516 gnd.n6394 gnd.n6393 9.3005
R13517 gnd.n6392 gnd.n6215 9.3005
R13518 gnd.n6391 gnd.n6390 9.3005
R13519 gnd.n6389 gnd.n6216 9.3005
R13520 gnd.n6388 gnd.n6387 9.3005
R13521 gnd.n6386 gnd.n6219 9.3005
R13522 gnd.n6385 gnd.n6384 9.3005
R13523 gnd.n6383 gnd.n6220 9.3005
R13524 gnd.n917 gnd.n916 9.3005
R13525 gnd.n6545 gnd.n6544 9.3005
R13526 gnd.n6546 gnd.n914 9.3005
R13527 gnd.n6549 gnd.n6548 9.3005
R13528 gnd.n6547 gnd.n915 9.3005
R13529 gnd.n876 gnd.n875 9.3005
R13530 gnd.n6603 gnd.n6602 9.3005
R13531 gnd.n6604 gnd.n873 9.3005
R13532 gnd.n6606 gnd.n6605 9.3005
R13533 gnd.n6607 gnd.n872 9.3005
R13534 gnd.n6610 gnd.n6609 9.3005
R13535 gnd.n6611 gnd.n870 9.3005
R13536 gnd.n6766 gnd.n6765 9.3005
R13537 gnd.n6764 gnd.n871 9.3005
R13538 gnd.n6763 gnd.n6762 9.3005
R13539 gnd.n6761 gnd.n6612 9.3005
R13540 gnd.n6760 gnd.n6615 9.3005
R13541 gnd.n5687 gnd.n5686 9.3005
R13542 gnd.n7058 gnd.n7057 9.3005
R13543 gnd.n7059 gnd.n476 9.3005
R13544 gnd.n7061 gnd.n7060 9.3005
R13545 gnd.n460 gnd.n459 9.3005
R13546 gnd.n7074 gnd.n7073 9.3005
R13547 gnd.n7075 gnd.n458 9.3005
R13548 gnd.n7077 gnd.n7076 9.3005
R13549 gnd.n444 gnd.n443 9.3005
R13550 gnd.n7090 gnd.n7089 9.3005
R13551 gnd.n7091 gnd.n442 9.3005
R13552 gnd.n7093 gnd.n7092 9.3005
R13553 gnd.n426 gnd.n425 9.3005
R13554 gnd.n7106 gnd.n7105 9.3005
R13555 gnd.n7107 gnd.n424 9.3005
R13556 gnd.n7109 gnd.n7108 9.3005
R13557 gnd.n410 gnd.n409 9.3005
R13558 gnd.n7122 gnd.n7121 9.3005
R13559 gnd.n7123 gnd.n407 9.3005
R13560 gnd.n7128 gnd.n7127 9.3005
R13561 gnd.n7126 gnd.n408 9.3005
R13562 gnd.n7125 gnd.n7124 9.3005
R13563 gnd.n377 gnd.n375 9.3005
R13564 gnd.n7179 gnd.n7178 9.3005
R13565 gnd.n7177 gnd.n376 9.3005
R13566 gnd.n7176 gnd.n7175 9.3005
R13567 gnd.n7174 gnd.n378 9.3005
R13568 gnd.n7173 gnd.n7172 9.3005
R13569 gnd.n316 gnd.n314 9.3005
R13570 gnd.n7318 gnd.n7317 9.3005
R13571 gnd.n7316 gnd.n315 9.3005
R13572 gnd.n7315 gnd.n7314 9.3005
R13573 gnd.n7313 gnd.n317 9.3005
R13574 gnd.n7312 gnd.n7311 9.3005
R13575 gnd.n7310 gnd.n321 9.3005
R13576 gnd.n7309 gnd.n7308 9.3005
R13577 gnd.n7307 gnd.n322 9.3005
R13578 gnd.n293 gnd.n292 9.3005
R13579 gnd.n7332 gnd.n7331 9.3005
R13580 gnd.n7333 gnd.n291 9.3005
R13581 gnd.n7335 gnd.n7334 9.3005
R13582 gnd.n277 gnd.n276 9.3005
R13583 gnd.n7348 gnd.n7347 9.3005
R13584 gnd.n7349 gnd.n275 9.3005
R13585 gnd.n7351 gnd.n7350 9.3005
R13586 gnd.n263 gnd.n262 9.3005
R13587 gnd.n7364 gnd.n7363 9.3005
R13588 gnd.n7365 gnd.n261 9.3005
R13589 gnd.n7367 gnd.n7366 9.3005
R13590 gnd.n247 gnd.n246 9.3005
R13591 gnd.n7380 gnd.n7379 9.3005
R13592 gnd.n7381 gnd.n245 9.3005
R13593 gnd.n7383 gnd.n7382 9.3005
R13594 gnd.n232 gnd.n231 9.3005
R13595 gnd.n7396 gnd.n7395 9.3005
R13596 gnd.n7397 gnd.n230 9.3005
R13597 gnd.n7399 gnd.n7398 9.3005
R13598 gnd.n217 gnd.n216 9.3005
R13599 gnd.n7412 gnd.n7411 9.3005
R13600 gnd.n7413 gnd.n214 9.3005
R13601 gnd.n7483 gnd.n7482 9.3005
R13602 gnd.n7481 gnd.n215 9.3005
R13603 gnd.n7480 gnd.n7479 9.3005
R13604 gnd.n7478 gnd.n7414 9.3005
R13605 gnd.n7477 gnd.n7476 9.3005
R13606 gnd.n478 gnd.n477 9.3005
R13607 gnd.n7473 gnd.n7416 9.3005
R13608 gnd.n7472 gnd.n7471 9.3005
R13609 gnd.n7470 gnd.n7421 9.3005
R13610 gnd.n7469 gnd.n7468 9.3005
R13611 gnd.n7467 gnd.n7422 9.3005
R13612 gnd.n7466 gnd.n7465 9.3005
R13613 gnd.n7464 gnd.n7429 9.3005
R13614 gnd.n7463 gnd.n7462 9.3005
R13615 gnd.n7461 gnd.n7430 9.3005
R13616 gnd.n7460 gnd.n7459 9.3005
R13617 gnd.n7458 gnd.n7437 9.3005
R13618 gnd.n7457 gnd.n7456 9.3005
R13619 gnd.n7455 gnd.n7438 9.3005
R13620 gnd.n7454 gnd.n7453 9.3005
R13621 gnd.n7452 gnd.n7445 9.3005
R13622 gnd.n7451 gnd.n7450 9.3005
R13623 gnd.n120 gnd.n117 9.3005
R13624 gnd.n7577 gnd.n7576 9.3005
R13625 gnd.n7475 gnd.n7474 9.3005
R13626 gnd.n6970 gnd.n565 9.3005
R13627 gnd.n6969 gnd.n6968 9.3005
R13628 gnd.n6967 gnd.n567 9.3005
R13629 gnd.n6966 gnd.n6965 9.3005
R13630 gnd.n6964 gnd.n570 9.3005
R13631 gnd.n6963 gnd.n6962 9.3005
R13632 gnd.n6961 gnd.n571 9.3005
R13633 gnd.n6960 gnd.n6959 9.3005
R13634 gnd.n6958 gnd.n574 9.3005
R13635 gnd.n6957 gnd.n6956 9.3005
R13636 gnd.n6955 gnd.n575 9.3005
R13637 gnd.n6954 gnd.n6953 9.3005
R13638 gnd.n6952 gnd.n578 9.3005
R13639 gnd.n6951 gnd.n6950 9.3005
R13640 gnd.n6949 gnd.n579 9.3005
R13641 gnd.n6948 gnd.n6947 9.3005
R13642 gnd.n6946 gnd.n582 9.3005
R13643 gnd.n6945 gnd.n6944 9.3005
R13644 gnd.n6943 gnd.n583 9.3005
R13645 gnd.n6942 gnd.n6941 9.3005
R13646 gnd.n6940 gnd.n384 9.3005
R13647 gnd.n7161 gnd.n383 9.3005
R13648 gnd.n7163 gnd.n7162 9.3005
R13649 gnd.n7164 gnd.n381 9.3005
R13650 gnd.n7167 gnd.n7166 9.3005
R13651 gnd.n7165 gnd.n382 9.3005
R13652 gnd.n354 gnd.n352 9.3005
R13653 gnd.n7209 gnd.n7208 9.3005
R13654 gnd.n7207 gnd.n353 9.3005
R13655 gnd.n7206 gnd.n7205 9.3005
R13656 gnd.n7204 gnd.n75 9.3005
R13657 gnd.n7626 gnd.n76 9.3005
R13658 gnd.n7625 gnd.n7624 9.3005
R13659 gnd.n7623 gnd.n77 9.3005
R13660 gnd.n7622 gnd.n7621 9.3005
R13661 gnd.n7620 gnd.n81 9.3005
R13662 gnd.n7619 gnd.n7618 9.3005
R13663 gnd.n7617 gnd.n82 9.3005
R13664 gnd.n7616 gnd.n7615 9.3005
R13665 gnd.n7614 gnd.n86 9.3005
R13666 gnd.n7613 gnd.n7612 9.3005
R13667 gnd.n7611 gnd.n87 9.3005
R13668 gnd.n7610 gnd.n7609 9.3005
R13669 gnd.n7608 gnd.n91 9.3005
R13670 gnd.n7607 gnd.n7606 9.3005
R13671 gnd.n7605 gnd.n92 9.3005
R13672 gnd.n7604 gnd.n7603 9.3005
R13673 gnd.n7602 gnd.n96 9.3005
R13674 gnd.n7601 gnd.n7600 9.3005
R13675 gnd.n7599 gnd.n97 9.3005
R13676 gnd.n7598 gnd.n7597 9.3005
R13677 gnd.n7596 gnd.n101 9.3005
R13678 gnd.n7595 gnd.n7594 9.3005
R13679 gnd.n7593 gnd.n102 9.3005
R13680 gnd.n7592 gnd.n7591 9.3005
R13681 gnd.n7590 gnd.n106 9.3005
R13682 gnd.n7589 gnd.n7588 9.3005
R13683 gnd.n7587 gnd.n107 9.3005
R13684 gnd.n7586 gnd.n7585 9.3005
R13685 gnd.n7584 gnd.n111 9.3005
R13686 gnd.n7583 gnd.n7582 9.3005
R13687 gnd.n7581 gnd.n112 9.3005
R13688 gnd.n7580 gnd.n7579 9.3005
R13689 gnd.n7578 gnd.n116 9.3005
R13690 gnd.n6972 gnd.n6971 9.3005
R13691 gnd.t19 gnd.n4267 9.24152
R13692 gnd.n4647 gnd.t56 9.24152
R13693 gnd.n3373 gnd.t81 9.24152
R13694 gnd.t217 gnd.n1925 9.24152
R13695 gnd.n5517 gnd.t178 9.24152
R13696 gnd.n7111 gnd.t188 9.24152
R13697 gnd.n259 gnd.t182 9.24152
R13698 gnd.t348 gnd.t19 8.92286
R13699 gnd.n5835 gnd.n1297 8.92286
R13700 gnd.n6040 gnd.n1209 8.92286
R13701 gnd.n6117 gnd.n1119 8.92286
R13702 gnd.n6183 gnd.n1058 8.92286
R13703 gnd.n6422 gnd.n1033 8.92286
R13704 gnd.n6486 gnd.n970 8.92286
R13705 gnd.n6510 gnd.n945 8.92286
R13706 gnd.n6600 gnd.n880 8.92286
R13707 gnd.n6769 gnd.n6768 8.92286
R13708 gnd.n4626 gnd.n4601 8.92171
R13709 gnd.n4594 gnd.n4569 8.92171
R13710 gnd.n4562 gnd.n4537 8.92171
R13711 gnd.n4531 gnd.n4506 8.92171
R13712 gnd.n4499 gnd.n4474 8.92171
R13713 gnd.n4467 gnd.n4442 8.92171
R13714 gnd.n4435 gnd.n4410 8.92171
R13715 gnd.n4404 gnd.n4379 8.92171
R13716 gnd.n727 gnd.n709 8.72777
R13717 gnd.n3613 gnd.t10 8.60421
R13718 gnd.t245 gnd.n1957 8.60421
R13719 gnd.n5549 gnd.t180 8.60421
R13720 gnd.n5825 gnd.n1305 8.60421
R13721 gnd.n1179 gnd.t155 8.60421
R13722 gnd.t163 gnd.n1016 8.60421
R13723 gnd.n7079 gnd.t274 8.60421
R13724 gnd.n228 gnd.t271 8.60421
R13725 gnd.n3655 gnd.n3635 8.43467
R13726 gnd.n54 gnd.n34 8.43467
R13727 gnd.n5209 gnd.n0 8.41456
R13728 gnd.n7627 gnd.n7626 8.41456
R13729 gnd.n5677 gnd.t115 8.28555
R13730 gnd.n4627 gnd.n4599 8.14595
R13731 gnd.n4595 gnd.n4567 8.14595
R13732 gnd.n4563 gnd.n4535 8.14595
R13733 gnd.n4532 gnd.n4504 8.14595
R13734 gnd.n4500 gnd.n4472 8.14595
R13735 gnd.n4468 gnd.n4440 8.14595
R13736 gnd.n4436 gnd.n4408 8.14595
R13737 gnd.n4405 gnd.n4377 8.14595
R13738 gnd.n4632 gnd.n4631 7.97301
R13739 gnd.t12 gnd.n4167 7.9669
R13740 gnd.n5889 gnd.t166 7.9669
R13741 gnd.n6372 gnd.t346 7.9669
R13742 gnd.n7576 gnd.n120 7.75808
R13743 gnd.n6714 gnd.n6710 7.75808
R13744 gnd.n5775 gnd.n5774 7.75808
R13745 gnd.n4824 gnd.n4763 7.75808
R13746 gnd.n4664 gnd.n3355 7.64824
R13747 gnd.n1282 gnd.t130 7.64824
R13748 gnd.n5968 gnd.n5967 7.64824
R13749 gnd.t21 gnd.n1218 7.64824
R13750 gnd.n6093 gnd.t165 7.64824
R13751 gnd.n6165 gnd.t165 7.64824
R13752 gnd.n6288 gnd.t172 7.64824
R13753 gnd.t172 gnd.n990 7.64824
R13754 gnd.t4 gnd.n937 7.64824
R13755 gnd.n6590 gnd.n890 7.64824
R13756 gnd.n6568 gnd.t118 7.64824
R13757 gnd.n4100 gnd.t16 7.32958
R13758 gnd.t350 gnd.t60 7.32958
R13759 gnd.n1432 gnd.n1431 7.30353
R13760 gnd.n726 gnd.n725 7.30353
R13761 gnd.n4060 gnd.n3779 7.01093
R13762 gnd.n3782 gnd.n3780 7.01093
R13763 gnd.n4070 gnd.n4069 7.01093
R13764 gnd.n4081 gnd.n3763 7.01093
R13765 gnd.n4080 gnd.n3766 7.01093
R13766 gnd.n4091 gnd.n3754 7.01093
R13767 gnd.n3757 gnd.n3755 7.01093
R13768 gnd.n4101 gnd.n4100 7.01093
R13769 gnd.n4111 gnd.n3735 7.01093
R13770 gnd.n4110 gnd.n3738 7.01093
R13771 gnd.n4127 gnd.n3728 7.01093
R13772 gnd.n4137 gnd.n3719 7.01093
R13773 gnd.n4148 gnd.n4147 7.01093
R13774 gnd.n4168 gnd.n3704 7.01093
R13775 gnd.n4167 gnd.n3683 7.01093
R13776 gnd.n4185 gnd.n3684 7.01093
R13777 gnd.n4179 gnd.n4178 7.01093
R13778 gnd.n4195 gnd.n3531 7.01093
R13779 gnd.n4205 gnd.n3523 7.01093
R13780 gnd.n4216 gnd.n3514 7.01093
R13781 gnd.n3613 gnd.n3612 7.01093
R13782 gnd.n4226 gnd.n4225 7.01093
R13783 gnd.n4237 gnd.n3497 7.01093
R13784 gnd.n4236 gnd.n3500 7.01093
R13785 gnd.n4247 gnd.n3489 7.01093
R13786 gnd.n4257 gnd.n4256 7.01093
R13787 gnd.n4268 gnd.n3471 7.01093
R13788 gnd.n4267 gnd.n3474 7.01093
R13789 gnd.n4278 gnd.n3462 7.01093
R13790 gnd.n3465 gnd.n3463 7.01093
R13791 gnd.n4288 gnd.n4287 7.01093
R13792 gnd.n4299 gnd.n3446 7.01093
R13793 gnd.n3440 gnd.n3438 7.01093
R13794 gnd.n4319 gnd.n4318 7.01093
R13795 gnd.n4330 gnd.n3421 7.01093
R13796 gnd.n4329 gnd.n3424 7.01093
R13797 gnd.n4340 gnd.n3412 7.01093
R13798 gnd.n3415 gnd.n3413 7.01093
R13799 gnd.n4361 gnd.n3395 7.01093
R13800 gnd.n4360 gnd.n3398 7.01093
R13801 gnd.n4371 gnd.n3387 7.01093
R13802 gnd.n3388 gnd.n3380 7.01093
R13803 gnd.n4637 gnd.n4636 7.01093
R13804 gnd.n4647 gnd.n3370 7.01093
R13805 gnd.n4646 gnd.n3373 7.01093
R13806 gnd.n4657 gnd.n3364 7.01093
R13807 gnd.n4664 gnd.n1988 7.01093
R13808 gnd.n6173 gnd.t169 7.01093
R13809 gnd.t174 gnd.n6414 7.01093
R13810 gnd.n6768 gnd.t88 7.01093
R13811 gnd.n3738 gnd.t8 6.69227
R13812 gnd.n4268 gnd.t348 6.69227
R13813 gnd.n4350 gnd.t7 6.69227
R13814 gnd.n5372 gnd.t180 6.69227
R13815 gnd.n5948 gnd.t170 6.69227
R13816 gnd.n6237 gnd.t150 6.69227
R13817 gnd.n6866 gnd.t274 6.69227
R13818 gnd.n807 gnd.n806 6.5566
R13819 gnd.n1598 gnd.n1597 6.5566
R13820 gnd.n1458 gnd.n1452 6.5566
R13821 gnd.n787 gnd.n694 6.5566
R13822 gnd.n5911 gnd.n5901 6.37362
R13823 gnd.n6023 gnd.n1225 6.37362
R13824 gnd.n6102 gnd.n1134 6.37362
R13825 gnd.n6470 gnd.n984 6.37362
R13826 gnd.n6532 gnd.n928 6.37362
R13827 gnd.n6523 gnd.n911 6.37362
R13828 gnd.n6775 gnd.t28 6.37362
R13829 gnd.n5802 gnd.n5800 6.20656
R13830 gnd.n7538 gnd.n7535 6.20656
R13831 gnd.n5029 gnd.n4902 6.20656
R13832 gnd.n6695 gnd.n6691 6.20656
R13833 gnd.t146 gnd.n4159 6.05496
R13834 gnd.n4160 gnd.t18 6.05496
R13835 gnd.n4225 gnd.t159 6.05496
R13836 gnd.n3587 gnd.t14 6.05496
R13837 gnd.n5315 gnd.t178 6.05496
R13838 gnd.n6905 gnd.t188 6.05496
R13839 gnd.n4629 gnd.n4599 5.81868
R13840 gnd.n4597 gnd.n4567 5.81868
R13841 gnd.n4565 gnd.n4535 5.81868
R13842 gnd.n4534 gnd.n4504 5.81868
R13843 gnd.n4502 gnd.n4472 5.81868
R13844 gnd.n4470 gnd.n4440 5.81868
R13845 gnd.n4438 gnd.n4408 5.81868
R13846 gnd.n4407 gnd.n4377 5.81868
R13847 gnd.n5975 gnd.t42 5.73631
R13848 gnd.t161 gnd.n1209 5.73631
R13849 gnd.t144 gnd.n1078 5.73631
R13850 gnd.n6298 gnd.t136 5.73631
R13851 gnd.t162 gnd.n945 5.73631
R13852 gnd.t88 gnd.n646 5.73631
R13853 gnd.n802 gnd.n534 5.62001
R13854 gnd.n1605 gnd.n1390 5.62001
R13855 gnd.n1605 gnd.n1391 5.62001
R13856 gnd.n794 gnd.n534 5.62001
R13857 gnd.n3919 gnd.n3914 5.4308
R13858 gnd.n4672 gnd.n2055 5.4308
R13859 gnd.n4237 gnd.t13 5.41765
R13860 gnd.t20 gnd.n3482 5.41765
R13861 gnd.n4309 gnd.t23 5.41765
R13862 gnd.n5430 gnd.t237 5.41765
R13863 gnd.n5275 gnd.t198 5.41765
R13864 gnd.n1194 gnd.t176 5.41765
R13865 gnd.n6494 gnd.t152 5.41765
R13866 gnd.n7158 gnd.t211 5.41765
R13867 gnd.t276 gnd.n359 5.41765
R13868 gnd.n6015 gnd.n1233 5.09899
R13869 gnd.n5889 gnd.n5888 5.09899
R13870 gnd.t2 gnd.n6109 5.09899
R13871 gnd.n6157 gnd.n1080 5.09899
R13872 gnd.n6095 gnd.n6094 5.09899
R13873 gnd.n6462 gnd.n992 5.09899
R13874 gnd.n6267 gnd.n6266 5.09899
R13875 gnd.n6478 gnd.t149 5.09899
R13876 gnd.n6373 gnd.n6372 5.09899
R13877 gnd.n6542 gnd.n919 5.09899
R13878 gnd.n4627 gnd.n4626 5.04292
R13879 gnd.n4595 gnd.n4594 5.04292
R13880 gnd.n4563 gnd.n4562 5.04292
R13881 gnd.n4532 gnd.n4531 5.04292
R13882 gnd.n4500 gnd.n4499 5.04292
R13883 gnd.n4468 gnd.n4467 5.04292
R13884 gnd.n4436 gnd.n4435 5.04292
R13885 gnd.n4405 gnd.n4404 5.04292
R13886 gnd.n3675 gnd.n3674 4.82753
R13887 gnd.n74 gnd.n73 4.82753
R13888 gnd.n4206 gnd.t5 4.78034
R13889 gnd.n3465 gnd.t11 4.78034
R13890 gnd.n5296 gnd.t223 4.78034
R13891 gnd.t176 gnd.n1111 4.78034
R13892 gnd.n6247 gnd.t152 4.78034
R13893 gnd.t53 gnd.n648 4.78034
R13894 gnd.n6916 gnd.t248 4.78034
R13895 gnd.n3680 gnd.n3677 4.74817
R13896 gnd.n4192 gnd.n3533 4.74817
R13897 gnd.n4190 gnd.n3534 4.74817
R13898 gnd.n3616 gnd.n3610 4.74817
R13899 gnd.n3696 gnd.n3677 4.74817
R13900 gnd.n3695 gnd.n3533 4.74817
R13901 gnd.n4191 gnd.n4190 4.74817
R13902 gnd.n3616 gnd.n3615 4.74817
R13903 gnd.n7324 gnd.n7323 4.74817
R13904 gnd.n337 gnd.n304 4.74817
R13905 gnd.n7225 gnd.n303 4.74817
R13906 gnd.n327 gnd.n302 4.74817
R13907 gnd.n7303 gnd.n301 4.74817
R13908 gnd.n7324 gnd.n305 4.74817
R13909 gnd.n7322 gnd.n304 4.74817
R13910 gnd.n338 gnd.n303 4.74817
R13911 gnd.n7226 gnd.n302 4.74817
R13912 gnd.n328 gnd.n301 4.74817
R13913 gnd.n5465 gnd.n5464 4.74817
R13914 gnd.n5452 gnd.n1769 4.74817
R13915 gnd.n5450 gnd.n1768 4.74817
R13916 gnd.n5438 gnd.n1767 4.74817
R13917 gnd.n1766 gnd.n1763 4.74817
R13918 gnd.n5465 gnd.n1770 4.74817
R13919 gnd.n5463 gnd.n1769 4.74817
R13920 gnd.n5453 gnd.n1768 4.74817
R13921 gnd.n5449 gnd.n1767 4.74817
R13922 gnd.n5439 gnd.n1766 4.74817
R13923 gnd.n3655 gnd.n3654 4.7074
R13924 gnd.n54 gnd.n53 4.7074
R13925 gnd.n3675 gnd.n3655 4.65959
R13926 gnd.n74 gnd.n54 4.65959
R13927 gnd.n7018 gnd.n536 4.6132
R13928 gnd.n1609 gnd.n1606 4.6132
R13929 gnd.n5358 gnd.n1364 4.46168
R13930 gnd.n5968 gnd.t143 4.46168
R13931 gnd.t173 gnd.n890 4.46168
R13932 gnd.n7046 gnd.n518 4.46168
R13933 gnd.n722 gnd.n709 4.46111
R13934 gnd.n4612 gnd.n4608 4.38594
R13935 gnd.n4580 gnd.n4576 4.38594
R13936 gnd.n4548 gnd.n4544 4.38594
R13937 gnd.n4517 gnd.n4513 4.38594
R13938 gnd.n4485 gnd.n4481 4.38594
R13939 gnd.n4453 gnd.n4449 4.38594
R13940 gnd.n4421 gnd.n4417 4.38594
R13941 gnd.n4390 gnd.n4386 4.38594
R13942 gnd.n4623 gnd.n4601 4.26717
R13943 gnd.n4591 gnd.n4569 4.26717
R13944 gnd.n4559 gnd.n4537 4.26717
R13945 gnd.n4528 gnd.n4506 4.26717
R13946 gnd.n4496 gnd.n4474 4.26717
R13947 gnd.n4464 gnd.n4442 4.26717
R13948 gnd.n4432 gnd.n4410 4.26717
R13949 gnd.n4401 gnd.n4379 4.26717
R13950 gnd.t6 gnd.n3711 4.14303
R13951 gnd.n3424 gnd.t9 4.14303
R13952 gnd.n5335 gnd.t204 4.14303
R13953 gnd.n1149 gnd.t342 4.14303
R13954 gnd.n6289 gnd.t25 4.14303
R13955 gnd.n6885 gnd.t221 4.14303
R13956 gnd.n4631 gnd.n4630 4.08274
R13957 gnd.n806 gnd.n691 4.05904
R13958 gnd.n1597 gnd.n1596 4.05904
R13959 gnd.n1462 gnd.n1452 4.05904
R13960 gnd.n788 gnd.n787 4.05904
R13961 gnd.n15 gnd.n7 3.99943
R13962 gnd.t130 gnd.n1254 3.82437
R13963 gnd.n6007 gnd.n1241 3.82437
R13964 gnd.n5927 gnd.n5883 3.82437
R13965 gnd.n6149 gnd.n1087 3.82437
R13966 gnd.n6087 gnd.n1150 3.82437
R13967 gnd.n6454 gnd.n1000 3.82437
R13968 gnd.n6307 gnd.n6306 3.82437
R13969 gnd.n6381 gnd.n6380 3.82437
R13970 gnd.n6552 gnd.n6551 3.82437
R13971 gnd.n6613 gnd.t53 3.82437
R13972 gnd.n4631 gnd.n4503 3.70378
R13973 gnd.n4189 gnd.n3676 3.65935
R13974 gnd.n15 gnd.n14 3.60163
R13975 gnd.n5078 gnd.t38 3.50571
R13976 gnd.n5386 gnd.t67 3.50571
R13977 gnd.n6846 gnd.t49 3.50571
R13978 gnd.n7493 gnd.t45 3.50571
R13979 gnd.n4622 gnd.n4603 3.49141
R13980 gnd.n4590 gnd.n4571 3.49141
R13981 gnd.n4558 gnd.n4539 3.49141
R13982 gnd.n4527 gnd.n4508 3.49141
R13983 gnd.n4495 gnd.n4476 3.49141
R13984 gnd.n4463 gnd.n4444 3.49141
R13985 gnd.n4431 gnd.n4412 3.49141
R13986 gnd.n4400 gnd.n4381 3.49141
R13987 gnd.n5853 gnd.t42 3.18706
R13988 gnd.n6781 gnd.t101 3.18706
R13989 gnd.n3718 gnd.t6 2.8684
R13990 gnd.n3656 gnd.t317 2.82907
R13991 gnd.n3656 gnd.t263 2.82907
R13992 gnd.n3658 gnd.t303 2.82907
R13993 gnd.n3658 gnd.t179 2.82907
R13994 gnd.n3660 gnd.t210 2.82907
R13995 gnd.n3660 gnd.t187 2.82907
R13996 gnd.n3662 gnd.t185 2.82907
R13997 gnd.n3662 gnd.t329 2.82907
R13998 gnd.n3664 gnd.t195 2.82907
R13999 gnd.n3664 gnd.t255 2.82907
R14000 gnd.n3666 gnd.t292 2.82907
R14001 gnd.n3666 gnd.t235 2.82907
R14002 gnd.n3668 gnd.t270 2.82907
R14003 gnd.n3668 gnd.t191 2.82907
R14004 gnd.n3670 gnd.t239 2.82907
R14005 gnd.n3670 gnd.t322 2.82907
R14006 gnd.n3672 gnd.t297 2.82907
R14007 gnd.n3672 gnd.t296 2.82907
R14008 gnd.n3617 gnd.t203 2.82907
R14009 gnd.n3617 gnd.t233 2.82907
R14010 gnd.n3619 gnd.t254 2.82907
R14011 gnd.n3619 gnd.t318 2.82907
R14012 gnd.n3621 gnd.t229 2.82907
R14013 gnd.n3621 gnd.t220 2.82907
R14014 gnd.n3623 gnd.t278 2.82907
R14015 gnd.n3623 gnd.t265 2.82907
R14016 gnd.n3625 gnd.t325 2.82907
R14017 gnd.n3625 gnd.t242 2.82907
R14018 gnd.n3627 gnd.t260 2.82907
R14019 gnd.n3627 gnd.t291 2.82907
R14020 gnd.n3629 gnd.t306 2.82907
R14021 gnd.n3629 gnd.t230 2.82907
R14022 gnd.n3631 gnd.t243 2.82907
R14023 gnd.n3631 gnd.t273 2.82907
R14024 gnd.n3633 gnd.t193 2.82907
R14025 gnd.n3633 gnd.t214 2.82907
R14026 gnd.n3636 gnd.t328 2.82907
R14027 gnd.n3636 gnd.t205 2.82907
R14028 gnd.n3638 gnd.t224 2.82907
R14029 gnd.n3638 gnd.t295 2.82907
R14030 gnd.n3640 gnd.t199 2.82907
R14031 gnd.n3640 gnd.t337 2.82907
R14032 gnd.n3642 gnd.t247 2.82907
R14033 gnd.n3642 gnd.t238 2.82907
R14034 gnd.n3644 gnd.t307 2.82907
R14035 gnd.n3644 gnd.t216 2.82907
R14036 gnd.n3646 gnd.t232 2.82907
R14037 gnd.n3646 gnd.t262 2.82907
R14038 gnd.n3648 gnd.t279 2.82907
R14039 gnd.n3648 gnd.t200 2.82907
R14040 gnd.n3650 gnd.t218 2.82907
R14041 gnd.n3650 gnd.t253 2.82907
R14042 gnd.n3652 gnd.t324 2.82907
R14043 gnd.n3652 gnd.t330 2.82907
R14044 gnd.n71 gnd.t201 2.82907
R14045 gnd.n71 gnd.t219 2.82907
R14046 gnd.n69 gnd.t283 2.82907
R14047 gnd.n69 gnd.t183 2.82907
R14048 gnd.n67 gnd.t315 2.82907
R14049 gnd.n67 gnd.t226 2.82907
R14050 gnd.n65 gnd.t336 2.82907
R14051 gnd.n65 gnd.t251 2.82907
R14052 gnd.n63 gnd.t207 2.82907
R14053 gnd.n63 gnd.t327 2.82907
R14054 gnd.n61 gnd.t298 2.82907
R14055 gnd.n61 gnd.t310 2.82907
R14056 gnd.n59 gnd.t313 2.82907
R14057 gnd.n59 gnd.t334 2.82907
R14058 gnd.n57 gnd.t308 2.82907
R14059 gnd.n57 gnd.t259 2.82907
R14060 gnd.n55 gnd.t222 2.82907
R14061 gnd.n55 gnd.t294 2.82907
R14062 gnd.n32 gnd.t197 2.82907
R14063 gnd.n32 gnd.t209 2.82907
R14064 gnd.n30 gnd.t311 2.82907
R14065 gnd.n30 gnd.t281 2.82907
R14066 gnd.n28 gnd.t266 2.82907
R14067 gnd.n28 gnd.t331 2.82907
R14068 gnd.n26 gnd.t321 2.82907
R14069 gnd.n26 gnd.t299 2.82907
R14070 gnd.n24 gnd.t280 2.82907
R14071 gnd.n24 gnd.t316 2.82907
R14072 gnd.n22 gnd.t305 2.82907
R14073 gnd.n22 gnd.t312 2.82907
R14074 gnd.n20 gnd.t258 2.82907
R14075 gnd.n20 gnd.t212 2.82907
R14076 gnd.n18 gnd.t189 2.82907
R14077 gnd.n18 gnd.t287 2.82907
R14078 gnd.n16 gnd.t268 2.82907
R14079 gnd.n16 gnd.t335 2.82907
R14080 gnd.n51 gnd.t326 2.82907
R14081 gnd.n51 gnd.t332 2.82907
R14082 gnd.n49 gnd.t284 2.82907
R14083 gnd.n49 gnd.t257 2.82907
R14084 gnd.n47 gnd.t241 2.82907
R14085 gnd.n47 gnd.t314 2.82907
R14086 gnd.n45 gnd.t301 2.82907
R14087 gnd.n45 gnd.t267 2.82907
R14088 gnd.n43 gnd.t256 2.82907
R14089 gnd.n43 gnd.t290 2.82907
R14090 gnd.n41 gnd.t277 2.82907
R14091 gnd.n41 gnd.t286 2.82907
R14092 gnd.n39 gnd.t228 2.82907
R14093 gnd.n39 gnd.t333 2.82907
R14094 gnd.n37 gnd.t323 2.82907
R14095 gnd.n37 gnd.t249 2.82907
R14096 gnd.n35 gnd.t244 2.82907
R14097 gnd.n35 gnd.t319 2.82907
R14098 gnd.n4619 gnd.n4618 2.71565
R14099 gnd.n4587 gnd.n4586 2.71565
R14100 gnd.n4555 gnd.n4554 2.71565
R14101 gnd.n4524 gnd.n4523 2.71565
R14102 gnd.n4492 gnd.n4491 2.71565
R14103 gnd.n4460 gnd.n4459 2.71565
R14104 gnd.n4428 gnd.n4427 2.71565
R14105 gnd.n4397 gnd.n4396 2.71565
R14106 gnd.n5999 gnd.n1248 2.54975
R14107 gnd.n5901 gnd.t0 2.54975
R14108 gnd.n5948 gnd.n5947 2.54975
R14109 gnd.n6125 gnd.t145 2.54975
R14110 gnd.n6141 gnd.n1095 2.54975
R14111 gnd.n6110 gnd.t2 2.54975
R14112 gnd.n6080 gnd.n6079 2.54975
R14113 gnd.n6446 gnd.n1008 2.54975
R14114 gnd.n6256 gnd.t149 2.54975
R14115 gnd.n6316 gnd.n6257 2.54975
R14116 gnd.n6335 gnd.t148 2.54975
R14117 gnd.n6352 gnd.n6237 2.54975
R14118 gnd.n6523 gnd.t1 2.54975
R14119 gnd.n6560 gnd.n906 2.54975
R14120 gnd.n4189 gnd.n3677 2.27742
R14121 gnd.n4189 gnd.n3533 2.27742
R14122 gnd.n4190 gnd.n4189 2.27742
R14123 gnd.n4189 gnd.n3616 2.27742
R14124 gnd.n7325 gnd.n7324 2.27742
R14125 gnd.n7325 gnd.n304 2.27742
R14126 gnd.n7325 gnd.n303 2.27742
R14127 gnd.n7325 gnd.n302 2.27742
R14128 gnd.n7325 gnd.n301 2.27742
R14129 gnd.n5466 gnd.n5465 2.27742
R14130 gnd.n5466 gnd.n1769 2.27742
R14131 gnd.n5466 gnd.n1768 2.27742
R14132 gnd.n5466 gnd.n1767 2.27742
R14133 gnd.n5466 gnd.n1766 2.27742
R14134 gnd.n4069 gnd.t34 2.23109
R14135 gnd.n4194 gnd.t5 2.23109
R14136 gnd.n6165 gnd.t342 2.23109
R14137 gnd.t25 gnd.n6288 2.23109
R14138 gnd.n236 gnd.t208 2.23109
R14139 gnd.n4615 gnd.n4605 1.93989
R14140 gnd.n4583 gnd.n4573 1.93989
R14141 gnd.n4551 gnd.n4541 1.93989
R14142 gnd.n4520 gnd.n4510 1.93989
R14143 gnd.n4488 gnd.n4478 1.93989
R14144 gnd.n4456 gnd.n4446 1.93989
R14145 gnd.n4424 gnd.n4414 1.93989
R14146 gnd.n4393 gnd.n4383 1.93989
R14147 gnd.t157 gnd.n4080 1.59378
R14148 gnd.n3490 gnd.t20 1.59378
R14149 gnd.n3588 gnd.t23 1.59378
R14150 gnd.n5118 gnd.t213 1.59378
R14151 gnd.n5320 gnd.t202 1.59378
R14152 gnd.n6890 gnd.t293 1.59378
R14153 gnd.n7385 gnd.t196 1.59378
R14154 gnd.n1530 gnd.t31 1.27512
R14155 gnd.n1530 gnd.n1411 1.27512
R14156 gnd.n5991 gnd.n1256 1.27512
R14157 gnd.n5940 gnd.n5939 1.27512
R14158 gnd.n6133 gnd.n1103 1.27512
R14159 gnd.n1179 gnd.n1163 1.27512
R14160 gnd.n6438 gnd.n1016 1.27512
R14161 gnd.n6326 gnd.n6325 1.27512
R14162 gnd.n6344 gnd.n6242 1.27512
R14163 gnd.n6569 gnd.n6568 1.27512
R14164 gnd.n6789 gnd.n655 1.27512
R14165 gnd.n3922 gnd.n3914 1.16414
R14166 gnd.n4675 gnd.n2055 1.16414
R14167 gnd.n4614 gnd.n4607 1.16414
R14168 gnd.n4582 gnd.n4575 1.16414
R14169 gnd.n4550 gnd.n4543 1.16414
R14170 gnd.n4519 gnd.n4512 1.16414
R14171 gnd.n4487 gnd.n4480 1.16414
R14172 gnd.n4455 gnd.n4448 1.16414
R14173 gnd.n4423 gnd.n4416 1.16414
R14174 gnd.n4392 gnd.n4385 1.16414
R14175 gnd.n7018 gnd.n7017 0.970197
R14176 gnd.n5735 gnd.n1606 0.970197
R14177 gnd.n4598 gnd.n4566 0.962709
R14178 gnd.n4630 gnd.n4598 0.962709
R14179 gnd.n4471 gnd.n4439 0.962709
R14180 gnd.n4503 gnd.n4471 0.962709
R14181 gnd.n4160 gnd.t146 0.956468
R14182 gnd.n4298 gnd.t14 0.956468
R14183 gnd.n5160 gnd.t269 0.956468
R14184 gnd.n5280 gnd.t186 0.956468
R14185 gnd.n1288 gnd.t350 0.956468
R14186 gnd.n5999 gnd.t141 0.956468
R14187 gnd.n906 gnd.t352 0.956468
R14188 gnd.n670 gnd.t354 0.956468
R14189 gnd.n6938 gnd.t227 0.956468
R14190 gnd.n7353 gnd.t225 0.956468
R14191 gnd.n3667 gnd.n3665 0.773756
R14192 gnd.n66 gnd.n64 0.773756
R14193 gnd.n3674 gnd.n3673 0.773756
R14194 gnd.n3673 gnd.n3671 0.773756
R14195 gnd.n3671 gnd.n3669 0.773756
R14196 gnd.n3669 gnd.n3667 0.773756
R14197 gnd.n3665 gnd.n3663 0.773756
R14198 gnd.n3663 gnd.n3661 0.773756
R14199 gnd.n3661 gnd.n3659 0.773756
R14200 gnd.n3659 gnd.n3657 0.773756
R14201 gnd.n58 gnd.n56 0.773756
R14202 gnd.n60 gnd.n58 0.773756
R14203 gnd.n62 gnd.n60 0.773756
R14204 gnd.n64 gnd.n62 0.773756
R14205 gnd.n68 gnd.n66 0.773756
R14206 gnd.n70 gnd.n68 0.773756
R14207 gnd.n72 gnd.n70 0.773756
R14208 gnd.n73 gnd.n72 0.773756
R14209 gnd.n2 gnd.n1 0.672012
R14210 gnd.n3 gnd.n2 0.672012
R14211 gnd.n4 gnd.n3 0.672012
R14212 gnd.n5 gnd.n4 0.672012
R14213 gnd.n6 gnd.n5 0.672012
R14214 gnd.n7 gnd.n6 0.672012
R14215 gnd.n9 gnd.n8 0.672012
R14216 gnd.n10 gnd.n9 0.672012
R14217 gnd.n11 gnd.n10 0.672012
R14218 gnd.n12 gnd.n11 0.672012
R14219 gnd.n13 gnd.n12 0.672012
R14220 gnd.n14 gnd.n13 0.672012
R14221 gnd.n5983 gnd.t74 0.637812
R14222 gnd.n5920 gnd.t168 0.637812
R14223 gnd.n6081 gnd.t169 0.637812
R14224 gnd.n6415 gnd.t174 0.637812
R14225 gnd.n6374 gnd.t175 0.637812
R14226 gnd.n6781 gnd.t63 0.637812
R14227 gnd.n7628 gnd.n7627 0.63688
R14228 gnd gnd.n0 0.634843
R14229 gnd.n3635 gnd.n3634 0.573776
R14230 gnd.n3634 gnd.n3632 0.573776
R14231 gnd.n3632 gnd.n3630 0.573776
R14232 gnd.n3630 gnd.n3628 0.573776
R14233 gnd.n3628 gnd.n3626 0.573776
R14234 gnd.n3626 gnd.n3624 0.573776
R14235 gnd.n3624 gnd.n3622 0.573776
R14236 gnd.n3622 gnd.n3620 0.573776
R14237 gnd.n3620 gnd.n3618 0.573776
R14238 gnd.n3654 gnd.n3653 0.573776
R14239 gnd.n3653 gnd.n3651 0.573776
R14240 gnd.n3651 gnd.n3649 0.573776
R14241 gnd.n3649 gnd.n3647 0.573776
R14242 gnd.n3647 gnd.n3645 0.573776
R14243 gnd.n3645 gnd.n3643 0.573776
R14244 gnd.n3643 gnd.n3641 0.573776
R14245 gnd.n3641 gnd.n3639 0.573776
R14246 gnd.n3639 gnd.n3637 0.573776
R14247 gnd.n19 gnd.n17 0.573776
R14248 gnd.n21 gnd.n19 0.573776
R14249 gnd.n23 gnd.n21 0.573776
R14250 gnd.n25 gnd.n23 0.573776
R14251 gnd.n27 gnd.n25 0.573776
R14252 gnd.n29 gnd.n27 0.573776
R14253 gnd.n31 gnd.n29 0.573776
R14254 gnd.n33 gnd.n31 0.573776
R14255 gnd.n34 gnd.n33 0.573776
R14256 gnd.n38 gnd.n36 0.573776
R14257 gnd.n40 gnd.n38 0.573776
R14258 gnd.n42 gnd.n40 0.573776
R14259 gnd.n44 gnd.n42 0.573776
R14260 gnd.n46 gnd.n44 0.573776
R14261 gnd.n48 gnd.n46 0.573776
R14262 gnd.n50 gnd.n48 0.573776
R14263 gnd.n52 gnd.n50 0.573776
R14264 gnd.n53 gnd.n52 0.573776
R14265 gnd.n7325 gnd.n300 0.5435
R14266 gnd.n5466 gnd.n1765 0.5435
R14267 gnd.n5688 gnd.n5687 0.523366
R14268 gnd.n6619 gnd.n6615 0.523366
R14269 gnd.n6813 gnd.n6812 0.489829
R14270 gnd.n5820 gnd.n1308 0.489829
R14271 gnd.n3562 gnd.n2059 0.486781
R14272 gnd.n3971 gnd.n3970 0.48678
R14273 gnd.n4653 gnd.n2013 0.480683
R14274 gnd.n4055 gnd.n4054 0.480683
R14275 gnd.n4826 gnd.n4825 0.477634
R14276 gnd.n5073 gnd.n1986 0.477634
R14277 gnd.n7476 gnd.n7475 0.477634
R14278 gnd.n7578 gnd.n7577 0.477634
R14279 gnd.n7570 gnd.n7569 0.465439
R14280 gnd.n7499 gnd.n7498 0.465439
R14281 gnd.n6978 gnd.n562 0.465439
R14282 gnd.n7051 gnd.n7050 0.465439
R14283 gnd.n5768 gnd.n5767 0.465439
R14284 gnd.n5699 gnd.n5698 0.465439
R14285 gnd.n4992 gnd.n4987 0.465439
R14286 gnd.n5067 gnd.n5066 0.465439
R14287 gnd.n3138 gnd.n2186 0.459342
R14288 gnd.n2501 gnd.n2495 0.459342
R14289 gnd.n7218 gnd.n7217 0.459342
R14290 gnd.n3350 gnd.n3349 0.459342
R14291 gnd.n5800 gnd.n5799 0.388379
R14292 gnd.n4611 gnd.n4610 0.388379
R14293 gnd.n4579 gnd.n4578 0.388379
R14294 gnd.n4547 gnd.n4546 0.388379
R14295 gnd.n4516 gnd.n4515 0.388379
R14296 gnd.n4484 gnd.n4483 0.388379
R14297 gnd.n4452 gnd.n4451 0.388379
R14298 gnd.n4420 gnd.n4419 0.388379
R14299 gnd.n4389 gnd.n4388 0.388379
R14300 gnd.n7539 gnd.n7538 0.388379
R14301 gnd.n4902 gnd.n4898 0.388379
R14302 gnd.n6691 gnd.n6687 0.388379
R14303 gnd.n5690 gnd.n5689 0.377553
R14304 gnd.n6620 gnd.n477 0.377553
R14305 gnd.n7628 gnd.n15 0.374463
R14306 gnd.t7 gnd.n4349 0.319156
R14307 gnd.n5217 gnd.t234 0.319156
R14308 gnd.n5241 gnd.t184 0.319156
R14309 gnd.n6108 gnd.t338 0.319156
R14310 gnd.t155 gnd.t154 0.319156
R14311 gnd.t135 gnd.t163 0.319156
R14312 gnd.t344 gnd.n976 0.319156
R14313 gnd.n7211 gnd.t285 0.319156
R14314 gnd.n7305 gnd.t300 0.319156
R14315 gnd.n3889 gnd.n3867 0.311721
R14316 gnd gnd.n7628 0.295112
R14317 gnd.n4720 gnd.n4719 0.268793
R14318 gnd.n5784 gnd.n1341 0.247451
R14319 gnd.n6971 gnd.n566 0.247451
R14320 gnd.n4719 gnd.n4718 0.241354
R14321 gnd.n536 gnd.n533 0.229039
R14322 gnd.n539 gnd.n536 0.229039
R14323 gnd.n1609 gnd.n1608 0.229039
R14324 gnd.n1610 gnd.n1609 0.229039
R14325 gnd.n3676 gnd.n0 0.210825
R14326 gnd.n4043 gnd.n3842 0.206293
R14327 gnd.n4628 gnd.n4600 0.155672
R14328 gnd.n4621 gnd.n4600 0.155672
R14329 gnd.n4621 gnd.n4620 0.155672
R14330 gnd.n4620 gnd.n4604 0.155672
R14331 gnd.n4613 gnd.n4604 0.155672
R14332 gnd.n4613 gnd.n4612 0.155672
R14333 gnd.n4596 gnd.n4568 0.155672
R14334 gnd.n4589 gnd.n4568 0.155672
R14335 gnd.n4589 gnd.n4588 0.155672
R14336 gnd.n4588 gnd.n4572 0.155672
R14337 gnd.n4581 gnd.n4572 0.155672
R14338 gnd.n4581 gnd.n4580 0.155672
R14339 gnd.n4564 gnd.n4536 0.155672
R14340 gnd.n4557 gnd.n4536 0.155672
R14341 gnd.n4557 gnd.n4556 0.155672
R14342 gnd.n4556 gnd.n4540 0.155672
R14343 gnd.n4549 gnd.n4540 0.155672
R14344 gnd.n4549 gnd.n4548 0.155672
R14345 gnd.n4533 gnd.n4505 0.155672
R14346 gnd.n4526 gnd.n4505 0.155672
R14347 gnd.n4526 gnd.n4525 0.155672
R14348 gnd.n4525 gnd.n4509 0.155672
R14349 gnd.n4518 gnd.n4509 0.155672
R14350 gnd.n4518 gnd.n4517 0.155672
R14351 gnd.n4501 gnd.n4473 0.155672
R14352 gnd.n4494 gnd.n4473 0.155672
R14353 gnd.n4494 gnd.n4493 0.155672
R14354 gnd.n4493 gnd.n4477 0.155672
R14355 gnd.n4486 gnd.n4477 0.155672
R14356 gnd.n4486 gnd.n4485 0.155672
R14357 gnd.n4469 gnd.n4441 0.155672
R14358 gnd.n4462 gnd.n4441 0.155672
R14359 gnd.n4462 gnd.n4461 0.155672
R14360 gnd.n4461 gnd.n4445 0.155672
R14361 gnd.n4454 gnd.n4445 0.155672
R14362 gnd.n4454 gnd.n4453 0.155672
R14363 gnd.n4437 gnd.n4409 0.155672
R14364 gnd.n4430 gnd.n4409 0.155672
R14365 gnd.n4430 gnd.n4429 0.155672
R14366 gnd.n4429 gnd.n4413 0.155672
R14367 gnd.n4422 gnd.n4413 0.155672
R14368 gnd.n4422 gnd.n4421 0.155672
R14369 gnd.n4406 gnd.n4378 0.155672
R14370 gnd.n4399 gnd.n4378 0.155672
R14371 gnd.n4399 gnd.n4398 0.155672
R14372 gnd.n4398 gnd.n4382 0.155672
R14373 gnd.n4391 gnd.n4382 0.155672
R14374 gnd.n4391 gnd.n4390 0.155672
R14375 gnd.n4751 gnd.n2013 0.152939
R14376 gnd.n4751 gnd.n4750 0.152939
R14377 gnd.n4750 gnd.n4749 0.152939
R14378 gnd.n4749 gnd.n2015 0.152939
R14379 gnd.n2016 gnd.n2015 0.152939
R14380 gnd.n2017 gnd.n2016 0.152939
R14381 gnd.n2018 gnd.n2017 0.152939
R14382 gnd.n2019 gnd.n2018 0.152939
R14383 gnd.n2020 gnd.n2019 0.152939
R14384 gnd.n2021 gnd.n2020 0.152939
R14385 gnd.n2022 gnd.n2021 0.152939
R14386 gnd.n2023 gnd.n2022 0.152939
R14387 gnd.n2024 gnd.n2023 0.152939
R14388 gnd.n2025 gnd.n2024 0.152939
R14389 gnd.n4721 gnd.n2025 0.152939
R14390 gnd.n4721 gnd.n4720 0.152939
R14391 gnd.n4056 gnd.n4055 0.152939
R14392 gnd.n4056 gnd.n3760 0.152939
R14393 gnd.n4084 gnd.n3760 0.152939
R14394 gnd.n4085 gnd.n4084 0.152939
R14395 gnd.n4086 gnd.n4085 0.152939
R14396 gnd.n4087 gnd.n4086 0.152939
R14397 gnd.n4087 gnd.n3732 0.152939
R14398 gnd.n4114 gnd.n3732 0.152939
R14399 gnd.n4115 gnd.n4114 0.152939
R14400 gnd.n4116 gnd.n4115 0.152939
R14401 gnd.n4117 gnd.n4116 0.152939
R14402 gnd.n4118 gnd.n4117 0.152939
R14403 gnd.n4120 gnd.n4118 0.152939
R14404 gnd.n4120 gnd.n4119 0.152939
R14405 gnd.n4119 gnd.n3700 0.152939
R14406 gnd.n4173 gnd.n3700 0.152939
R14407 gnd.n4174 gnd.n4173 0.152939
R14408 gnd.n4175 gnd.n4174 0.152939
R14409 gnd.n4175 gnd.n3518 0.152939
R14410 gnd.n4209 gnd.n3518 0.152939
R14411 gnd.n4210 gnd.n4209 0.152939
R14412 gnd.n4211 gnd.n4210 0.152939
R14413 gnd.n4212 gnd.n4211 0.152939
R14414 gnd.n4212 gnd.n3494 0.152939
R14415 gnd.n4240 gnd.n3494 0.152939
R14416 gnd.n4241 gnd.n4240 0.152939
R14417 gnd.n4242 gnd.n4241 0.152939
R14418 gnd.n4243 gnd.n4242 0.152939
R14419 gnd.n4243 gnd.n3468 0.152939
R14420 gnd.n4271 gnd.n3468 0.152939
R14421 gnd.n4272 gnd.n4271 0.152939
R14422 gnd.n4273 gnd.n4272 0.152939
R14423 gnd.n4274 gnd.n4273 0.152939
R14424 gnd.n4274 gnd.n3443 0.152939
R14425 gnd.n4302 gnd.n3443 0.152939
R14426 gnd.n4303 gnd.n4302 0.152939
R14427 gnd.n4304 gnd.n4303 0.152939
R14428 gnd.n4305 gnd.n4304 0.152939
R14429 gnd.n4305 gnd.n3418 0.152939
R14430 gnd.n4333 gnd.n3418 0.152939
R14431 gnd.n4334 gnd.n4333 0.152939
R14432 gnd.n4335 gnd.n4334 0.152939
R14433 gnd.n4336 gnd.n4335 0.152939
R14434 gnd.n4336 gnd.n3392 0.152939
R14435 gnd.n4364 gnd.n3392 0.152939
R14436 gnd.n4365 gnd.n4364 0.152939
R14437 gnd.n4366 gnd.n4365 0.152939
R14438 gnd.n4367 gnd.n4366 0.152939
R14439 gnd.n4367 gnd.n3367 0.152939
R14440 gnd.n4650 gnd.n3367 0.152939
R14441 gnd.n4651 gnd.n4650 0.152939
R14442 gnd.n4652 gnd.n4651 0.152939
R14443 gnd.n4653 gnd.n4652 0.152939
R14444 gnd.n4054 gnd.n3784 0.152939
R14445 gnd.n3805 gnd.n3784 0.152939
R14446 gnd.n3806 gnd.n3805 0.152939
R14447 gnd.n3812 gnd.n3806 0.152939
R14448 gnd.n3813 gnd.n3812 0.152939
R14449 gnd.n3814 gnd.n3813 0.152939
R14450 gnd.n3814 gnd.n3803 0.152939
R14451 gnd.n3822 gnd.n3803 0.152939
R14452 gnd.n3823 gnd.n3822 0.152939
R14453 gnd.n3824 gnd.n3823 0.152939
R14454 gnd.n3824 gnd.n3801 0.152939
R14455 gnd.n3832 gnd.n3801 0.152939
R14456 gnd.n3833 gnd.n3832 0.152939
R14457 gnd.n3834 gnd.n3833 0.152939
R14458 gnd.n3834 gnd.n3799 0.152939
R14459 gnd.n3842 gnd.n3799 0.152939
R14460 gnd.n4718 gnd.n2030 0.152939
R14461 gnd.n2032 gnd.n2030 0.152939
R14462 gnd.n2033 gnd.n2032 0.152939
R14463 gnd.n2034 gnd.n2033 0.152939
R14464 gnd.n2035 gnd.n2034 0.152939
R14465 gnd.n2036 gnd.n2035 0.152939
R14466 gnd.n2037 gnd.n2036 0.152939
R14467 gnd.n2038 gnd.n2037 0.152939
R14468 gnd.n2039 gnd.n2038 0.152939
R14469 gnd.n2040 gnd.n2039 0.152939
R14470 gnd.n2041 gnd.n2040 0.152939
R14471 gnd.n2042 gnd.n2041 0.152939
R14472 gnd.n2043 gnd.n2042 0.152939
R14473 gnd.n2044 gnd.n2043 0.152939
R14474 gnd.n2045 gnd.n2044 0.152939
R14475 gnd.n2046 gnd.n2045 0.152939
R14476 gnd.n2047 gnd.n2046 0.152939
R14477 gnd.n2048 gnd.n2047 0.152939
R14478 gnd.n2049 gnd.n2048 0.152939
R14479 gnd.n2050 gnd.n2049 0.152939
R14480 gnd.n2051 gnd.n2050 0.152939
R14481 gnd.n2052 gnd.n2051 0.152939
R14482 gnd.n2056 gnd.n2052 0.152939
R14483 gnd.n2057 gnd.n2056 0.152939
R14484 gnd.n2058 gnd.n2057 0.152939
R14485 gnd.n2059 gnd.n2058 0.152939
R14486 gnd.n3536 gnd.n3535 0.152939
R14487 gnd.n3537 gnd.n3536 0.152939
R14488 gnd.n3538 gnd.n3537 0.152939
R14489 gnd.n3539 gnd.n3538 0.152939
R14490 gnd.n3540 gnd.n3539 0.152939
R14491 gnd.n3541 gnd.n3540 0.152939
R14492 gnd.n3542 gnd.n3541 0.152939
R14493 gnd.n3543 gnd.n3542 0.152939
R14494 gnd.n3544 gnd.n3543 0.152939
R14495 gnd.n3545 gnd.n3544 0.152939
R14496 gnd.n3546 gnd.n3545 0.152939
R14497 gnd.n3547 gnd.n3546 0.152939
R14498 gnd.n3548 gnd.n3547 0.152939
R14499 gnd.n3549 gnd.n3548 0.152939
R14500 gnd.n3550 gnd.n3549 0.152939
R14501 gnd.n3551 gnd.n3550 0.152939
R14502 gnd.n3552 gnd.n3551 0.152939
R14503 gnd.n3553 gnd.n3552 0.152939
R14504 gnd.n3554 gnd.n3553 0.152939
R14505 gnd.n3555 gnd.n3554 0.152939
R14506 gnd.n3556 gnd.n3555 0.152939
R14507 gnd.n3557 gnd.n3556 0.152939
R14508 gnd.n3558 gnd.n3557 0.152939
R14509 gnd.n3559 gnd.n3558 0.152939
R14510 gnd.n3560 gnd.n3559 0.152939
R14511 gnd.n3561 gnd.n3560 0.152939
R14512 gnd.n3563 gnd.n3561 0.152939
R14513 gnd.n3563 gnd.n3562 0.152939
R14514 gnd.n3972 gnd.n3971 0.152939
R14515 gnd.n3972 gnd.n3862 0.152939
R14516 gnd.n3987 gnd.n3862 0.152939
R14517 gnd.n3988 gnd.n3987 0.152939
R14518 gnd.n3989 gnd.n3988 0.152939
R14519 gnd.n3989 gnd.n3850 0.152939
R14520 gnd.n4003 gnd.n3850 0.152939
R14521 gnd.n4004 gnd.n4003 0.152939
R14522 gnd.n4005 gnd.n4004 0.152939
R14523 gnd.n4006 gnd.n4005 0.152939
R14524 gnd.n4007 gnd.n4006 0.152939
R14525 gnd.n4008 gnd.n4007 0.152939
R14526 gnd.n4009 gnd.n4008 0.152939
R14527 gnd.n4010 gnd.n4009 0.152939
R14528 gnd.n4011 gnd.n4010 0.152939
R14529 gnd.n4012 gnd.n4011 0.152939
R14530 gnd.n4013 gnd.n4012 0.152939
R14531 gnd.n4014 gnd.n4013 0.152939
R14532 gnd.n4015 gnd.n4014 0.152939
R14533 gnd.n4016 gnd.n4015 0.152939
R14534 gnd.n4017 gnd.n4016 0.152939
R14535 gnd.n4017 gnd.n3715 0.152939
R14536 gnd.n4140 gnd.n3715 0.152939
R14537 gnd.n4141 gnd.n4140 0.152939
R14538 gnd.n4142 gnd.n4141 0.152939
R14539 gnd.n4143 gnd.n4142 0.152939
R14540 gnd.n4143 gnd.n3678 0.152939
R14541 gnd.n4188 gnd.n3678 0.152939
R14542 gnd.n3890 gnd.n3889 0.152939
R14543 gnd.n3891 gnd.n3890 0.152939
R14544 gnd.n3892 gnd.n3891 0.152939
R14545 gnd.n3893 gnd.n3892 0.152939
R14546 gnd.n3894 gnd.n3893 0.152939
R14547 gnd.n3895 gnd.n3894 0.152939
R14548 gnd.n3896 gnd.n3895 0.152939
R14549 gnd.n3897 gnd.n3896 0.152939
R14550 gnd.n3898 gnd.n3897 0.152939
R14551 gnd.n3899 gnd.n3898 0.152939
R14552 gnd.n3900 gnd.n3899 0.152939
R14553 gnd.n3901 gnd.n3900 0.152939
R14554 gnd.n3902 gnd.n3901 0.152939
R14555 gnd.n3903 gnd.n3902 0.152939
R14556 gnd.n3904 gnd.n3903 0.152939
R14557 gnd.n3905 gnd.n3904 0.152939
R14558 gnd.n3906 gnd.n3905 0.152939
R14559 gnd.n3907 gnd.n3906 0.152939
R14560 gnd.n3908 gnd.n3907 0.152939
R14561 gnd.n3909 gnd.n3908 0.152939
R14562 gnd.n3910 gnd.n3909 0.152939
R14563 gnd.n3911 gnd.n3910 0.152939
R14564 gnd.n3915 gnd.n3911 0.152939
R14565 gnd.n3916 gnd.n3915 0.152939
R14566 gnd.n3916 gnd.n3873 0.152939
R14567 gnd.n3970 gnd.n3873 0.152939
R14568 gnd.n3138 gnd.n3137 0.152939
R14569 gnd.n3137 gnd.n3136 0.152939
R14570 gnd.n3136 gnd.n2192 0.152939
R14571 gnd.n2197 gnd.n2192 0.152939
R14572 gnd.n2198 gnd.n2197 0.152939
R14573 gnd.n2199 gnd.n2198 0.152939
R14574 gnd.n2204 gnd.n2199 0.152939
R14575 gnd.n2205 gnd.n2204 0.152939
R14576 gnd.n2206 gnd.n2205 0.152939
R14577 gnd.n2207 gnd.n2206 0.152939
R14578 gnd.n2212 gnd.n2207 0.152939
R14579 gnd.n2213 gnd.n2212 0.152939
R14580 gnd.n2214 gnd.n2213 0.152939
R14581 gnd.n2215 gnd.n2214 0.152939
R14582 gnd.n2220 gnd.n2215 0.152939
R14583 gnd.n2221 gnd.n2220 0.152939
R14584 gnd.n2222 gnd.n2221 0.152939
R14585 gnd.n2223 gnd.n2222 0.152939
R14586 gnd.n2228 gnd.n2223 0.152939
R14587 gnd.n2229 gnd.n2228 0.152939
R14588 gnd.n2230 gnd.n2229 0.152939
R14589 gnd.n2231 gnd.n2230 0.152939
R14590 gnd.n2236 gnd.n2231 0.152939
R14591 gnd.n2237 gnd.n2236 0.152939
R14592 gnd.n2238 gnd.n2237 0.152939
R14593 gnd.n2239 gnd.n2238 0.152939
R14594 gnd.n2244 gnd.n2239 0.152939
R14595 gnd.n2245 gnd.n2244 0.152939
R14596 gnd.n2246 gnd.n2245 0.152939
R14597 gnd.n2247 gnd.n2246 0.152939
R14598 gnd.n2252 gnd.n2247 0.152939
R14599 gnd.n2253 gnd.n2252 0.152939
R14600 gnd.n2254 gnd.n2253 0.152939
R14601 gnd.n2255 gnd.n2254 0.152939
R14602 gnd.n2260 gnd.n2255 0.152939
R14603 gnd.n2261 gnd.n2260 0.152939
R14604 gnd.n2262 gnd.n2261 0.152939
R14605 gnd.n2263 gnd.n2262 0.152939
R14606 gnd.n2268 gnd.n2263 0.152939
R14607 gnd.n2269 gnd.n2268 0.152939
R14608 gnd.n2270 gnd.n2269 0.152939
R14609 gnd.n2271 gnd.n2270 0.152939
R14610 gnd.n2276 gnd.n2271 0.152939
R14611 gnd.n2277 gnd.n2276 0.152939
R14612 gnd.n2278 gnd.n2277 0.152939
R14613 gnd.n2279 gnd.n2278 0.152939
R14614 gnd.n2284 gnd.n2279 0.152939
R14615 gnd.n2285 gnd.n2284 0.152939
R14616 gnd.n2286 gnd.n2285 0.152939
R14617 gnd.n2287 gnd.n2286 0.152939
R14618 gnd.n2292 gnd.n2287 0.152939
R14619 gnd.n2293 gnd.n2292 0.152939
R14620 gnd.n2294 gnd.n2293 0.152939
R14621 gnd.n2295 gnd.n2294 0.152939
R14622 gnd.n2300 gnd.n2295 0.152939
R14623 gnd.n2301 gnd.n2300 0.152939
R14624 gnd.n2302 gnd.n2301 0.152939
R14625 gnd.n2303 gnd.n2302 0.152939
R14626 gnd.n2308 gnd.n2303 0.152939
R14627 gnd.n2309 gnd.n2308 0.152939
R14628 gnd.n2310 gnd.n2309 0.152939
R14629 gnd.n2311 gnd.n2310 0.152939
R14630 gnd.n2316 gnd.n2311 0.152939
R14631 gnd.n2317 gnd.n2316 0.152939
R14632 gnd.n2318 gnd.n2317 0.152939
R14633 gnd.n2319 gnd.n2318 0.152939
R14634 gnd.n2324 gnd.n2319 0.152939
R14635 gnd.n2325 gnd.n2324 0.152939
R14636 gnd.n2326 gnd.n2325 0.152939
R14637 gnd.n2327 gnd.n2326 0.152939
R14638 gnd.n2332 gnd.n2327 0.152939
R14639 gnd.n2333 gnd.n2332 0.152939
R14640 gnd.n2334 gnd.n2333 0.152939
R14641 gnd.n2335 gnd.n2334 0.152939
R14642 gnd.n2340 gnd.n2335 0.152939
R14643 gnd.n2341 gnd.n2340 0.152939
R14644 gnd.n2342 gnd.n2341 0.152939
R14645 gnd.n2343 gnd.n2342 0.152939
R14646 gnd.n2348 gnd.n2343 0.152939
R14647 gnd.n2349 gnd.n2348 0.152939
R14648 gnd.n2350 gnd.n2349 0.152939
R14649 gnd.n2351 gnd.n2350 0.152939
R14650 gnd.n2356 gnd.n2351 0.152939
R14651 gnd.n2357 gnd.n2356 0.152939
R14652 gnd.n2358 gnd.n2357 0.152939
R14653 gnd.n2359 gnd.n2358 0.152939
R14654 gnd.n2364 gnd.n2359 0.152939
R14655 gnd.n2365 gnd.n2364 0.152939
R14656 gnd.n2366 gnd.n2365 0.152939
R14657 gnd.n2367 gnd.n2366 0.152939
R14658 gnd.n2372 gnd.n2367 0.152939
R14659 gnd.n2373 gnd.n2372 0.152939
R14660 gnd.n2374 gnd.n2373 0.152939
R14661 gnd.n2375 gnd.n2374 0.152939
R14662 gnd.n2380 gnd.n2375 0.152939
R14663 gnd.n2381 gnd.n2380 0.152939
R14664 gnd.n2382 gnd.n2381 0.152939
R14665 gnd.n2383 gnd.n2382 0.152939
R14666 gnd.n2388 gnd.n2383 0.152939
R14667 gnd.n2389 gnd.n2388 0.152939
R14668 gnd.n2390 gnd.n2389 0.152939
R14669 gnd.n2391 gnd.n2390 0.152939
R14670 gnd.n2396 gnd.n2391 0.152939
R14671 gnd.n2397 gnd.n2396 0.152939
R14672 gnd.n2398 gnd.n2397 0.152939
R14673 gnd.n2399 gnd.n2398 0.152939
R14674 gnd.n2404 gnd.n2399 0.152939
R14675 gnd.n2405 gnd.n2404 0.152939
R14676 gnd.n2406 gnd.n2405 0.152939
R14677 gnd.n2407 gnd.n2406 0.152939
R14678 gnd.n2412 gnd.n2407 0.152939
R14679 gnd.n2413 gnd.n2412 0.152939
R14680 gnd.n2414 gnd.n2413 0.152939
R14681 gnd.n2415 gnd.n2414 0.152939
R14682 gnd.n2420 gnd.n2415 0.152939
R14683 gnd.n2421 gnd.n2420 0.152939
R14684 gnd.n2422 gnd.n2421 0.152939
R14685 gnd.n2423 gnd.n2422 0.152939
R14686 gnd.n2428 gnd.n2423 0.152939
R14687 gnd.n2429 gnd.n2428 0.152939
R14688 gnd.n2430 gnd.n2429 0.152939
R14689 gnd.n2431 gnd.n2430 0.152939
R14690 gnd.n2436 gnd.n2431 0.152939
R14691 gnd.n2437 gnd.n2436 0.152939
R14692 gnd.n2438 gnd.n2437 0.152939
R14693 gnd.n2439 gnd.n2438 0.152939
R14694 gnd.n2444 gnd.n2439 0.152939
R14695 gnd.n2445 gnd.n2444 0.152939
R14696 gnd.n2446 gnd.n2445 0.152939
R14697 gnd.n2447 gnd.n2446 0.152939
R14698 gnd.n2452 gnd.n2447 0.152939
R14699 gnd.n2453 gnd.n2452 0.152939
R14700 gnd.n2454 gnd.n2453 0.152939
R14701 gnd.n2455 gnd.n2454 0.152939
R14702 gnd.n2460 gnd.n2455 0.152939
R14703 gnd.n2461 gnd.n2460 0.152939
R14704 gnd.n2462 gnd.n2461 0.152939
R14705 gnd.n2463 gnd.n2462 0.152939
R14706 gnd.n2468 gnd.n2463 0.152939
R14707 gnd.n2469 gnd.n2468 0.152939
R14708 gnd.n2470 gnd.n2469 0.152939
R14709 gnd.n2471 gnd.n2470 0.152939
R14710 gnd.n2476 gnd.n2471 0.152939
R14711 gnd.n2477 gnd.n2476 0.152939
R14712 gnd.n2478 gnd.n2477 0.152939
R14713 gnd.n2479 gnd.n2478 0.152939
R14714 gnd.n2484 gnd.n2479 0.152939
R14715 gnd.n2485 gnd.n2484 0.152939
R14716 gnd.n2486 gnd.n2485 0.152939
R14717 gnd.n2487 gnd.n2486 0.152939
R14718 gnd.n2492 gnd.n2487 0.152939
R14719 gnd.n2493 gnd.n2492 0.152939
R14720 gnd.n2494 gnd.n2493 0.152939
R14721 gnd.n2495 gnd.n2494 0.152939
R14722 gnd.n2824 gnd.n2501 0.152939
R14723 gnd.n2824 gnd.n2823 0.152939
R14724 gnd.n2823 gnd.n2822 0.152939
R14725 gnd.n2822 gnd.n2502 0.152939
R14726 gnd.n2507 gnd.n2502 0.152939
R14727 gnd.n2508 gnd.n2507 0.152939
R14728 gnd.n2509 gnd.n2508 0.152939
R14729 gnd.n2514 gnd.n2509 0.152939
R14730 gnd.n2515 gnd.n2514 0.152939
R14731 gnd.n2516 gnd.n2515 0.152939
R14732 gnd.n2517 gnd.n2516 0.152939
R14733 gnd.n2522 gnd.n2517 0.152939
R14734 gnd.n2523 gnd.n2522 0.152939
R14735 gnd.n2524 gnd.n2523 0.152939
R14736 gnd.n2525 gnd.n2524 0.152939
R14737 gnd.n2530 gnd.n2525 0.152939
R14738 gnd.n2531 gnd.n2530 0.152939
R14739 gnd.n2532 gnd.n2531 0.152939
R14740 gnd.n2533 gnd.n2532 0.152939
R14741 gnd.n2538 gnd.n2533 0.152939
R14742 gnd.n2539 gnd.n2538 0.152939
R14743 gnd.n2540 gnd.n2539 0.152939
R14744 gnd.n2541 gnd.n2540 0.152939
R14745 gnd.n2546 gnd.n2541 0.152939
R14746 gnd.n2547 gnd.n2546 0.152939
R14747 gnd.n2548 gnd.n2547 0.152939
R14748 gnd.n2549 gnd.n2548 0.152939
R14749 gnd.n2554 gnd.n2549 0.152939
R14750 gnd.n2555 gnd.n2554 0.152939
R14751 gnd.n2556 gnd.n2555 0.152939
R14752 gnd.n2557 gnd.n2556 0.152939
R14753 gnd.n2562 gnd.n2557 0.152939
R14754 gnd.n2563 gnd.n2562 0.152939
R14755 gnd.n2564 gnd.n2563 0.152939
R14756 gnd.n2565 gnd.n2564 0.152939
R14757 gnd.n2570 gnd.n2565 0.152939
R14758 gnd.n2571 gnd.n2570 0.152939
R14759 gnd.n2572 gnd.n2571 0.152939
R14760 gnd.n2573 gnd.n2572 0.152939
R14761 gnd.n2578 gnd.n2573 0.152939
R14762 gnd.n2579 gnd.n2578 0.152939
R14763 gnd.n2580 gnd.n2579 0.152939
R14764 gnd.n2581 gnd.n2580 0.152939
R14765 gnd.n2586 gnd.n2581 0.152939
R14766 gnd.n2587 gnd.n2586 0.152939
R14767 gnd.n2588 gnd.n2587 0.152939
R14768 gnd.n2589 gnd.n2588 0.152939
R14769 gnd.n2594 gnd.n2589 0.152939
R14770 gnd.n2595 gnd.n2594 0.152939
R14771 gnd.n2596 gnd.n2595 0.152939
R14772 gnd.n2597 gnd.n2596 0.152939
R14773 gnd.n2602 gnd.n2597 0.152939
R14774 gnd.n2603 gnd.n2602 0.152939
R14775 gnd.n2604 gnd.n2603 0.152939
R14776 gnd.n2605 gnd.n2604 0.152939
R14777 gnd.n2610 gnd.n2605 0.152939
R14778 gnd.n2611 gnd.n2610 0.152939
R14779 gnd.n2612 gnd.n2611 0.152939
R14780 gnd.n2613 gnd.n2612 0.152939
R14781 gnd.n2618 gnd.n2613 0.152939
R14782 gnd.n2619 gnd.n2618 0.152939
R14783 gnd.n2620 gnd.n2619 0.152939
R14784 gnd.n2621 gnd.n2620 0.152939
R14785 gnd.n2626 gnd.n2621 0.152939
R14786 gnd.n2627 gnd.n2626 0.152939
R14787 gnd.n2628 gnd.n2627 0.152939
R14788 gnd.n2629 gnd.n2628 0.152939
R14789 gnd.n2634 gnd.n2629 0.152939
R14790 gnd.n2635 gnd.n2634 0.152939
R14791 gnd.n2636 gnd.n2635 0.152939
R14792 gnd.n2637 gnd.n2636 0.152939
R14793 gnd.n2642 gnd.n2637 0.152939
R14794 gnd.n2643 gnd.n2642 0.152939
R14795 gnd.n2644 gnd.n2643 0.152939
R14796 gnd.n2645 gnd.n2644 0.152939
R14797 gnd.n2650 gnd.n2645 0.152939
R14798 gnd.n2651 gnd.n2650 0.152939
R14799 gnd.n2652 gnd.n2651 0.152939
R14800 gnd.n2653 gnd.n2652 0.152939
R14801 gnd.n2659 gnd.n2653 0.152939
R14802 gnd.n2660 gnd.n2659 0.152939
R14803 gnd.n2661 gnd.n2660 0.152939
R14804 gnd.n2661 gnd.n345 0.152939
R14805 gnd.n7218 gnd.n345 0.152939
R14806 gnd.n7326 gnd.n7325 0.152939
R14807 gnd.n7326 gnd.n283 0.152939
R14808 gnd.n7340 gnd.n283 0.152939
R14809 gnd.n7341 gnd.n7340 0.152939
R14810 gnd.n7342 gnd.n7341 0.152939
R14811 gnd.n7342 gnd.n269 0.152939
R14812 gnd.n7356 gnd.n269 0.152939
R14813 gnd.n7357 gnd.n7356 0.152939
R14814 gnd.n7358 gnd.n7357 0.152939
R14815 gnd.n7358 gnd.n253 0.152939
R14816 gnd.n7372 gnd.n253 0.152939
R14817 gnd.n7373 gnd.n7372 0.152939
R14818 gnd.n7374 gnd.n7373 0.152939
R14819 gnd.n7374 gnd.n239 0.152939
R14820 gnd.n7388 gnd.n239 0.152939
R14821 gnd.n7389 gnd.n7388 0.152939
R14822 gnd.n7390 gnd.n7389 0.152939
R14823 gnd.n7390 gnd.n222 0.152939
R14824 gnd.n7404 gnd.n222 0.152939
R14825 gnd.n7405 gnd.n7404 0.152939
R14826 gnd.n7406 gnd.n7405 0.152939
R14827 gnd.n7406 gnd.n206 0.152939
R14828 gnd.n7488 gnd.n206 0.152939
R14829 gnd.n7489 gnd.n7488 0.152939
R14830 gnd.n7490 gnd.n7489 0.152939
R14831 gnd.n7490 gnd.n129 0.152939
R14832 gnd.n7570 gnd.n129 0.152939
R14833 gnd.n7569 gnd.n130 0.152939
R14834 gnd.n132 gnd.n130 0.152939
R14835 gnd.n136 gnd.n132 0.152939
R14836 gnd.n137 gnd.n136 0.152939
R14837 gnd.n138 gnd.n137 0.152939
R14838 gnd.n139 gnd.n138 0.152939
R14839 gnd.n143 gnd.n139 0.152939
R14840 gnd.n144 gnd.n143 0.152939
R14841 gnd.n145 gnd.n144 0.152939
R14842 gnd.n146 gnd.n145 0.152939
R14843 gnd.n150 gnd.n146 0.152939
R14844 gnd.n151 gnd.n150 0.152939
R14845 gnd.n152 gnd.n151 0.152939
R14846 gnd.n153 gnd.n152 0.152939
R14847 gnd.n157 gnd.n153 0.152939
R14848 gnd.n158 gnd.n157 0.152939
R14849 gnd.n159 gnd.n158 0.152939
R14850 gnd.n160 gnd.n159 0.152939
R14851 gnd.n164 gnd.n160 0.152939
R14852 gnd.n165 gnd.n164 0.152939
R14853 gnd.n166 gnd.n165 0.152939
R14854 gnd.n167 gnd.n166 0.152939
R14855 gnd.n171 gnd.n167 0.152939
R14856 gnd.n172 gnd.n171 0.152939
R14857 gnd.n173 gnd.n172 0.152939
R14858 gnd.n174 gnd.n173 0.152939
R14859 gnd.n178 gnd.n174 0.152939
R14860 gnd.n179 gnd.n178 0.152939
R14861 gnd.n180 gnd.n179 0.152939
R14862 gnd.n181 gnd.n180 0.152939
R14863 gnd.n185 gnd.n181 0.152939
R14864 gnd.n186 gnd.n185 0.152939
R14865 gnd.n187 gnd.n186 0.152939
R14866 gnd.n188 gnd.n187 0.152939
R14867 gnd.n192 gnd.n188 0.152939
R14868 gnd.n193 gnd.n192 0.152939
R14869 gnd.n7500 gnd.n193 0.152939
R14870 gnd.n7500 gnd.n7499 0.152939
R14871 gnd.n6844 gnd.n562 0.152939
R14872 gnd.n6845 gnd.n6844 0.152939
R14873 gnd.n6845 gnd.n6842 0.152939
R14874 gnd.n6853 gnd.n6842 0.152939
R14875 gnd.n6854 gnd.n6853 0.152939
R14876 gnd.n6855 gnd.n6854 0.152939
R14877 gnd.n6856 gnd.n6855 0.152939
R14878 gnd.n6858 gnd.n6856 0.152939
R14879 gnd.n6858 gnd.n6857 0.152939
R14880 gnd.n6857 gnd.n597 0.152939
R14881 gnd.n597 gnd.n595 0.152939
R14882 gnd.n6893 gnd.n595 0.152939
R14883 gnd.n6894 gnd.n6893 0.152939
R14884 gnd.n6895 gnd.n6894 0.152939
R14885 gnd.n6896 gnd.n6895 0.152939
R14886 gnd.n6897 gnd.n6896 0.152939
R14887 gnd.n6897 gnd.n586 0.152939
R14888 gnd.n6920 gnd.n586 0.152939
R14889 gnd.n6921 gnd.n6920 0.152939
R14890 gnd.n6922 gnd.n6921 0.152939
R14891 gnd.n6923 gnd.n6922 0.152939
R14892 gnd.n6924 gnd.n6923 0.152939
R14893 gnd.n6925 gnd.n6924 0.152939
R14894 gnd.n6926 gnd.n6925 0.152939
R14895 gnd.n6928 gnd.n6926 0.152939
R14896 gnd.n6928 gnd.n6927 0.152939
R14897 gnd.n6927 gnd.n356 0.152939
R14898 gnd.n7195 gnd.n356 0.152939
R14899 gnd.n7196 gnd.n7195 0.152939
R14900 gnd.n7197 gnd.n7196 0.152939
R14901 gnd.n7198 gnd.n7197 0.152939
R14902 gnd.n7198 gnd.n333 0.152939
R14903 gnd.n7231 gnd.n333 0.152939
R14904 gnd.n7232 gnd.n7231 0.152939
R14905 gnd.n7233 gnd.n7232 0.152939
R14906 gnd.n7234 gnd.n7233 0.152939
R14907 gnd.n7235 gnd.n7234 0.152939
R14908 gnd.n7236 gnd.n7235 0.152939
R14909 gnd.n7237 gnd.n7236 0.152939
R14910 gnd.n7238 gnd.n7237 0.152939
R14911 gnd.n7239 gnd.n7238 0.152939
R14912 gnd.n7240 gnd.n7239 0.152939
R14913 gnd.n7241 gnd.n7240 0.152939
R14914 gnd.n7242 gnd.n7241 0.152939
R14915 gnd.n7243 gnd.n7242 0.152939
R14916 gnd.n7244 gnd.n7243 0.152939
R14917 gnd.n7245 gnd.n7244 0.152939
R14918 gnd.n7246 gnd.n7245 0.152939
R14919 gnd.n7247 gnd.n7246 0.152939
R14920 gnd.n7248 gnd.n7247 0.152939
R14921 gnd.n7249 gnd.n7248 0.152939
R14922 gnd.n7250 gnd.n7249 0.152939
R14923 gnd.n7251 gnd.n7250 0.152939
R14924 gnd.n7252 gnd.n7251 0.152939
R14925 gnd.n7253 gnd.n7252 0.152939
R14926 gnd.n7254 gnd.n7253 0.152939
R14927 gnd.n7255 gnd.n7254 0.152939
R14928 gnd.n7256 gnd.n7255 0.152939
R14929 gnd.n7257 gnd.n7256 0.152939
R14930 gnd.n7258 gnd.n7257 0.152939
R14931 gnd.n7260 gnd.n7258 0.152939
R14932 gnd.n7260 gnd.n7259 0.152939
R14933 gnd.n7259 gnd.n199 0.152939
R14934 gnd.n7498 gnd.n199 0.152939
R14935 gnd.n7050 gnd.n486 0.152939
R14936 gnd.n520 gnd.n486 0.152939
R14937 gnd.n521 gnd.n520 0.152939
R14938 gnd.n522 gnd.n521 0.152939
R14939 gnd.n523 gnd.n522 0.152939
R14940 gnd.n524 gnd.n523 0.152939
R14941 gnd.n525 gnd.n524 0.152939
R14942 gnd.n526 gnd.n525 0.152939
R14943 gnd.n527 gnd.n526 0.152939
R14944 gnd.n528 gnd.n527 0.152939
R14945 gnd.n529 gnd.n528 0.152939
R14946 gnd.n530 gnd.n529 0.152939
R14947 gnd.n531 gnd.n530 0.152939
R14948 gnd.n532 gnd.n531 0.152939
R14949 gnd.n533 gnd.n532 0.152939
R14950 gnd.n540 gnd.n539 0.152939
R14951 gnd.n541 gnd.n540 0.152939
R14952 gnd.n542 gnd.n541 0.152939
R14953 gnd.n543 gnd.n542 0.152939
R14954 gnd.n544 gnd.n543 0.152939
R14955 gnd.n545 gnd.n544 0.152939
R14956 gnd.n546 gnd.n545 0.152939
R14957 gnd.n547 gnd.n546 0.152939
R14958 gnd.n548 gnd.n547 0.152939
R14959 gnd.n549 gnd.n548 0.152939
R14960 gnd.n550 gnd.n549 0.152939
R14961 gnd.n551 gnd.n550 0.152939
R14962 gnd.n552 gnd.n551 0.152939
R14963 gnd.n553 gnd.n552 0.152939
R14964 gnd.n554 gnd.n553 0.152939
R14965 gnd.n555 gnd.n554 0.152939
R14966 gnd.n556 gnd.n555 0.152939
R14967 gnd.n6980 gnd.n556 0.152939
R14968 gnd.n6980 gnd.n6979 0.152939
R14969 gnd.n6979 gnd.n6978 0.152939
R14970 gnd.n7052 gnd.n7051 0.152939
R14971 gnd.n7052 gnd.n468 0.152939
R14972 gnd.n7066 gnd.n468 0.152939
R14973 gnd.n7067 gnd.n7066 0.152939
R14974 gnd.n7068 gnd.n7067 0.152939
R14975 gnd.n7068 gnd.n451 0.152939
R14976 gnd.n7082 gnd.n451 0.152939
R14977 gnd.n7083 gnd.n7082 0.152939
R14978 gnd.n7084 gnd.n7083 0.152939
R14979 gnd.n7084 gnd.n434 0.152939
R14980 gnd.n7098 gnd.n434 0.152939
R14981 gnd.n7099 gnd.n7098 0.152939
R14982 gnd.n7100 gnd.n7099 0.152939
R14983 gnd.n7100 gnd.n417 0.152939
R14984 gnd.n7114 gnd.n417 0.152939
R14985 gnd.n7115 gnd.n7114 0.152939
R14986 gnd.n7116 gnd.n7115 0.152939
R14987 gnd.n7116 gnd.n398 0.152939
R14988 gnd.n7133 gnd.n398 0.152939
R14989 gnd.n7134 gnd.n7133 0.152939
R14990 gnd.n7135 gnd.n7134 0.152939
R14991 gnd.n7135 gnd.n366 0.152939
R14992 gnd.n7184 gnd.n366 0.152939
R14993 gnd.n7185 gnd.n7184 0.152939
R14994 gnd.n7186 gnd.n7185 0.152939
R14995 gnd.n7186 gnd.n299 0.152939
R14996 gnd.n7325 gnd.n299 0.152939
R14997 gnd.n7149 gnd.n7148 0.152939
R14998 gnd.n7148 gnd.n347 0.152939
R14999 gnd.n1803 gnd.n1802 0.152939
R15000 gnd.n5258 gnd.n1803 0.152939
R15001 gnd.n5260 gnd.n5258 0.152939
R15002 gnd.n5261 gnd.n5260 0.152939
R15003 gnd.n5262 gnd.n5261 0.152939
R15004 gnd.n5263 gnd.n5262 0.152939
R15005 gnd.n5264 gnd.n5263 0.152939
R15006 gnd.n5265 gnd.n5264 0.152939
R15007 gnd.n5266 gnd.n5265 0.152939
R15008 gnd.n5266 gnd.n1847 0.152939
R15009 gnd.n5300 gnd.n1847 0.152939
R15010 gnd.n5301 gnd.n5300 0.152939
R15011 gnd.n5302 gnd.n5301 0.152939
R15012 gnd.n5303 gnd.n5302 0.152939
R15013 gnd.n5304 gnd.n5303 0.152939
R15014 gnd.n5305 gnd.n5304 0.152939
R15015 gnd.n5306 gnd.n5305 0.152939
R15016 gnd.n5306 gnd.n1837 0.152939
R15017 gnd.n5339 gnd.n1837 0.152939
R15018 gnd.n5340 gnd.n5339 0.152939
R15019 gnd.n5341 gnd.n5340 0.152939
R15020 gnd.n5342 gnd.n5341 0.152939
R15021 gnd.n5343 gnd.n5342 0.152939
R15022 gnd.n5346 gnd.n5343 0.152939
R15023 gnd.n5347 gnd.n5346 0.152939
R15024 gnd.n5348 gnd.n5347 0.152939
R15025 gnd.n5349 gnd.n5348 0.152939
R15026 gnd.n5353 gnd.n5349 0.152939
R15027 gnd.n5354 gnd.n5353 0.152939
R15028 gnd.n5355 gnd.n5354 0.152939
R15029 gnd.n5355 gnd.n1315 0.152939
R15030 gnd.n5812 gnd.n1315 0.152939
R15031 gnd.n5813 gnd.n5812 0.152939
R15032 gnd.n5814 gnd.n5813 0.152939
R15033 gnd.n5814 gnd.n1301 0.152939
R15034 gnd.n5828 gnd.n1301 0.152939
R15035 gnd.n5829 gnd.n5828 0.152939
R15036 gnd.n5830 gnd.n5829 0.152939
R15037 gnd.n5831 gnd.n5830 0.152939
R15038 gnd.n5831 gnd.n1259 0.152939
R15039 gnd.n5986 gnd.n1259 0.152939
R15040 gnd.n5987 gnd.n5986 0.152939
R15041 gnd.n5988 gnd.n5987 0.152939
R15042 gnd.n5988 gnd.n1244 0.152939
R15043 gnd.n6002 gnd.n1244 0.152939
R15044 gnd.n6003 gnd.n6002 0.152939
R15045 gnd.n6004 gnd.n6003 0.152939
R15046 gnd.n6004 gnd.n1228 0.152939
R15047 gnd.n6018 gnd.n1228 0.152939
R15048 gnd.n6019 gnd.n6018 0.152939
R15049 gnd.n6020 gnd.n6019 0.152939
R15050 gnd.n6020 gnd.n1213 0.152939
R15051 gnd.n6033 gnd.n1213 0.152939
R15052 gnd.n6034 gnd.n6033 0.152939
R15053 gnd.n6035 gnd.n6034 0.152939
R15054 gnd.n6036 gnd.n6035 0.152939
R15055 gnd.n6036 gnd.n1106 0.152939
R15056 gnd.n6128 gnd.n1106 0.152939
R15057 gnd.n6129 gnd.n6128 0.152939
R15058 gnd.n6130 gnd.n6129 0.152939
R15059 gnd.n6130 gnd.n1090 0.152939
R15060 gnd.n6144 gnd.n1090 0.152939
R15061 gnd.n6145 gnd.n6144 0.152939
R15062 gnd.n6146 gnd.n6145 0.152939
R15063 gnd.n6146 gnd.n1075 0.152939
R15064 gnd.n6160 gnd.n1075 0.152939
R15065 gnd.n6161 gnd.n6160 0.152939
R15066 gnd.n6162 gnd.n6161 0.152939
R15067 gnd.n6162 gnd.n1062 0.152939
R15068 gnd.n6176 gnd.n1062 0.152939
R15069 gnd.n6177 gnd.n6176 0.152939
R15070 gnd.n6178 gnd.n6177 0.152939
R15071 gnd.n6179 gnd.n6178 0.152939
R15072 gnd.n6179 gnd.n1019 0.152939
R15073 gnd.n6433 gnd.n1019 0.152939
R15074 gnd.n6434 gnd.n6433 0.152939
R15075 gnd.n6435 gnd.n6434 0.152939
R15076 gnd.n6435 gnd.n1003 0.152939
R15077 gnd.n6449 gnd.n1003 0.152939
R15078 gnd.n6450 gnd.n6449 0.152939
R15079 gnd.n6451 gnd.n6450 0.152939
R15080 gnd.n6451 gnd.n987 0.152939
R15081 gnd.n6465 gnd.n987 0.152939
R15082 gnd.n6466 gnd.n6465 0.152939
R15083 gnd.n6467 gnd.n6466 0.152939
R15084 gnd.n6467 gnd.n973 0.152939
R15085 gnd.n6481 gnd.n973 0.152939
R15086 gnd.n6482 gnd.n6481 0.152939
R15087 gnd.n6483 gnd.n6482 0.152939
R15088 gnd.n6483 gnd.n958 0.152939
R15089 gnd.n6497 gnd.n958 0.152939
R15090 gnd.n6498 gnd.n6497 0.152939
R15091 gnd.n6499 gnd.n6498 0.152939
R15092 gnd.n6499 gnd.n942 0.152939
R15093 gnd.n6513 gnd.n942 0.152939
R15094 gnd.n6514 gnd.n6513 0.152939
R15095 gnd.n6515 gnd.n6514 0.152939
R15096 gnd.n6515 gnd.n925 0.152939
R15097 gnd.n6535 gnd.n925 0.152939
R15098 gnd.n6536 gnd.n6535 0.152939
R15099 gnd.n6537 gnd.n6536 0.152939
R15100 gnd.n6538 gnd.n6537 0.152939
R15101 gnd.n6538 gnd.n885 0.152939
R15102 gnd.n6593 gnd.n885 0.152939
R15103 gnd.n6594 gnd.n6593 0.152939
R15104 gnd.n6595 gnd.n6594 0.152939
R15105 gnd.n6596 gnd.n6595 0.152939
R15106 gnd.n6596 gnd.n658 0.152939
R15107 gnd.n6784 gnd.n658 0.152939
R15108 gnd.n6785 gnd.n6784 0.152939
R15109 gnd.n6786 gnd.n6785 0.152939
R15110 gnd.n6786 gnd.n643 0.152939
R15111 gnd.n6801 gnd.n643 0.152939
R15112 gnd.n6802 gnd.n6801 0.152939
R15113 gnd.n6803 gnd.n6802 0.152939
R15114 gnd.n6804 gnd.n6803 0.152939
R15115 gnd.n6804 gnd.n613 0.152939
R15116 gnd.n6820 gnd.n613 0.152939
R15117 gnd.n6821 gnd.n6820 0.152939
R15118 gnd.n6822 gnd.n6821 0.152939
R15119 gnd.n6822 gnd.n609 0.152939
R15120 gnd.n6828 gnd.n609 0.152939
R15121 gnd.n6829 gnd.n6828 0.152939
R15122 gnd.n6830 gnd.n6829 0.152939
R15123 gnd.n6830 gnd.n605 0.152939
R15124 gnd.n6836 gnd.n605 0.152939
R15125 gnd.n6837 gnd.n6836 0.152939
R15126 gnd.n6838 gnd.n6837 0.152939
R15127 gnd.n6838 gnd.n601 0.152939
R15128 gnd.n6870 gnd.n601 0.152939
R15129 gnd.n6871 gnd.n6870 0.152939
R15130 gnd.n6872 gnd.n6871 0.152939
R15131 gnd.n6873 gnd.n6872 0.152939
R15132 gnd.n6874 gnd.n6873 0.152939
R15133 gnd.n6875 gnd.n6874 0.152939
R15134 gnd.n6876 gnd.n6875 0.152939
R15135 gnd.n6876 gnd.n591 0.152939
R15136 gnd.n6909 gnd.n591 0.152939
R15137 gnd.n6910 gnd.n6909 0.152939
R15138 gnd.n6911 gnd.n6910 0.152939
R15139 gnd.n6912 gnd.n6911 0.152939
R15140 gnd.n6912 gnd.n391 0.152939
R15141 gnd.n7142 gnd.n391 0.152939
R15142 gnd.n7143 gnd.n7142 0.152939
R15143 gnd.n7144 gnd.n7143 0.152939
R15144 gnd.n7145 gnd.n7144 0.152939
R15145 gnd.n7146 gnd.n7145 0.152939
R15146 gnd.n7147 gnd.n7146 0.152939
R15147 gnd.n7149 gnd.n7147 0.152939
R15148 gnd.n4827 gnd.n4826 0.152939
R15149 gnd.n4828 gnd.n4827 0.152939
R15150 gnd.n4829 gnd.n4828 0.152939
R15151 gnd.n4830 gnd.n4829 0.152939
R15152 gnd.n4831 gnd.n4830 0.152939
R15153 gnd.n4832 gnd.n4831 0.152939
R15154 gnd.n4833 gnd.n4832 0.152939
R15155 gnd.n4834 gnd.n4833 0.152939
R15156 gnd.n4835 gnd.n4834 0.152939
R15157 gnd.n4836 gnd.n4835 0.152939
R15158 gnd.n4837 gnd.n4836 0.152939
R15159 gnd.n4838 gnd.n4837 0.152939
R15160 gnd.n4839 gnd.n4838 0.152939
R15161 gnd.n4840 gnd.n4839 0.152939
R15162 gnd.n4841 gnd.n4840 0.152939
R15163 gnd.n4842 gnd.n4841 0.152939
R15164 gnd.n4843 gnd.n4842 0.152939
R15165 gnd.n4844 gnd.n4843 0.152939
R15166 gnd.n4844 gnd.n1905 0.152939
R15167 gnd.n5163 gnd.n1905 0.152939
R15168 gnd.n5164 gnd.n5163 0.152939
R15169 gnd.n5165 gnd.n5164 0.152939
R15170 gnd.n5166 gnd.n5165 0.152939
R15171 gnd.n5167 gnd.n5166 0.152939
R15172 gnd.n5167 gnd.n1870 0.152939
R15173 gnd.n5202 gnd.n1870 0.152939
R15174 gnd.n5203 gnd.n5202 0.152939
R15175 gnd.n5204 gnd.n5203 0.152939
R15176 gnd.n5205 gnd.n5204 0.152939
R15177 gnd.n5206 gnd.n5205 0.152939
R15178 gnd.n5207 gnd.n5206 0.152939
R15179 gnd.n4778 gnd.n1986 0.152939
R15180 gnd.n4786 gnd.n4778 0.152939
R15181 gnd.n4787 gnd.n4786 0.152939
R15182 gnd.n4788 gnd.n4787 0.152939
R15183 gnd.n4788 gnd.n4774 0.152939
R15184 gnd.n4796 gnd.n4774 0.152939
R15185 gnd.n4797 gnd.n4796 0.152939
R15186 gnd.n4798 gnd.n4797 0.152939
R15187 gnd.n4798 gnd.n4770 0.152939
R15188 gnd.n4806 gnd.n4770 0.152939
R15189 gnd.n4807 gnd.n4806 0.152939
R15190 gnd.n4808 gnd.n4807 0.152939
R15191 gnd.n4808 gnd.n4766 0.152939
R15192 gnd.n4816 gnd.n4766 0.152939
R15193 gnd.n4817 gnd.n4816 0.152939
R15194 gnd.n4818 gnd.n4817 0.152939
R15195 gnd.n4818 gnd.n4760 0.152939
R15196 gnd.n4825 gnd.n4760 0.152939
R15197 gnd.n5074 gnd.n5073 0.152939
R15198 gnd.n5075 gnd.n5074 0.152939
R15199 gnd.n5075 gnd.n1971 0.152939
R15200 gnd.n5089 gnd.n1971 0.152939
R15201 gnd.n5090 gnd.n5089 0.152939
R15202 gnd.n5091 gnd.n5090 0.152939
R15203 gnd.n5091 gnd.n1954 0.152939
R15204 gnd.n5105 gnd.n1954 0.152939
R15205 gnd.n5106 gnd.n5105 0.152939
R15206 gnd.n5107 gnd.n5106 0.152939
R15207 gnd.n5107 gnd.n1939 0.152939
R15208 gnd.n5121 gnd.n1939 0.152939
R15209 gnd.n5122 gnd.n5121 0.152939
R15210 gnd.n5123 gnd.n5122 0.152939
R15211 gnd.n5123 gnd.n1922 0.152939
R15212 gnd.n5137 gnd.n1922 0.152939
R15213 gnd.n5138 gnd.n5137 0.152939
R15214 gnd.n5139 gnd.n5138 0.152939
R15215 gnd.n5140 gnd.n5139 0.152939
R15216 gnd.n5141 gnd.n5140 0.152939
R15217 gnd.n5143 gnd.n5141 0.152939
R15218 gnd.n5143 gnd.n5142 0.152939
R15219 gnd.n5142 gnd.n1888 0.152939
R15220 gnd.n1889 gnd.n1888 0.152939
R15221 gnd.n1890 gnd.n1889 0.152939
R15222 gnd.n1891 gnd.n1890 0.152939
R15223 gnd.n1893 gnd.n1891 0.152939
R15224 gnd.n1893 gnd.n1892 0.152939
R15225 gnd.n1892 gnd.n1779 0.152939
R15226 gnd.n1780 gnd.n1779 0.152939
R15227 gnd.n1781 gnd.n1780 0.152939
R15228 gnd.n1861 gnd.n1781 0.152939
R15229 gnd.n1861 gnd.n1792 0.152939
R15230 gnd.n1793 gnd.n1792 0.152939
R15231 gnd.n1794 gnd.n1793 0.152939
R15232 gnd.n1794 gnd.n1755 0.152939
R15233 gnd.n5472 gnd.n1755 0.152939
R15234 gnd.n5473 gnd.n5472 0.152939
R15235 gnd.n5474 gnd.n5473 0.152939
R15236 gnd.n5474 gnd.n1739 0.152939
R15237 gnd.n5488 gnd.n1739 0.152939
R15238 gnd.n5489 gnd.n5488 0.152939
R15239 gnd.n5490 gnd.n5489 0.152939
R15240 gnd.n5490 gnd.n1721 0.152939
R15241 gnd.n5504 gnd.n1721 0.152939
R15242 gnd.n5505 gnd.n5504 0.152939
R15243 gnd.n5506 gnd.n5505 0.152939
R15244 gnd.n5506 gnd.n1705 0.152939
R15245 gnd.n5520 gnd.n1705 0.152939
R15246 gnd.n5521 gnd.n5520 0.152939
R15247 gnd.n5522 gnd.n5521 0.152939
R15248 gnd.n5522 gnd.n1687 0.152939
R15249 gnd.n5536 gnd.n1687 0.152939
R15250 gnd.n5537 gnd.n5536 0.152939
R15251 gnd.n5538 gnd.n5537 0.152939
R15252 gnd.n5538 gnd.n1671 0.152939
R15253 gnd.n5552 gnd.n1671 0.152939
R15254 gnd.n5553 gnd.n5552 0.152939
R15255 gnd.n5554 gnd.n5553 0.152939
R15256 gnd.n5554 gnd.n1652 0.152939
R15257 gnd.n5570 gnd.n1652 0.152939
R15258 gnd.n5571 gnd.n5570 0.152939
R15259 gnd.n5572 gnd.n5571 0.152939
R15260 gnd.n5690 gnd.n5572 0.152939
R15261 gnd.n5466 gnd.n1747 0.152939
R15262 gnd.n5480 gnd.n1747 0.152939
R15263 gnd.n5481 gnd.n5480 0.152939
R15264 gnd.n5482 gnd.n5481 0.152939
R15265 gnd.n5482 gnd.n1730 0.152939
R15266 gnd.n5496 gnd.n1730 0.152939
R15267 gnd.n5497 gnd.n5496 0.152939
R15268 gnd.n5498 gnd.n5497 0.152939
R15269 gnd.n5498 gnd.n1713 0.152939
R15270 gnd.n5512 gnd.n1713 0.152939
R15271 gnd.n5513 gnd.n5512 0.152939
R15272 gnd.n5514 gnd.n5513 0.152939
R15273 gnd.n5514 gnd.n1696 0.152939
R15274 gnd.n5528 gnd.n1696 0.152939
R15275 gnd.n5529 gnd.n5528 0.152939
R15276 gnd.n5530 gnd.n5529 0.152939
R15277 gnd.n5530 gnd.n1679 0.152939
R15278 gnd.n5544 gnd.n1679 0.152939
R15279 gnd.n5545 gnd.n5544 0.152939
R15280 gnd.n5546 gnd.n5545 0.152939
R15281 gnd.n5546 gnd.n1662 0.152939
R15282 gnd.n5560 gnd.n1662 0.152939
R15283 gnd.n5561 gnd.n5560 0.152939
R15284 gnd.n5562 gnd.n5561 0.152939
R15285 gnd.n5563 gnd.n5562 0.152939
R15286 gnd.n5563 gnd.n1361 0.152939
R15287 gnd.n5768 gnd.n1361 0.152939
R15288 gnd.n5767 gnd.n1362 0.152939
R15289 gnd.n1367 gnd.n1362 0.152939
R15290 gnd.n1368 gnd.n1367 0.152939
R15291 gnd.n1369 gnd.n1368 0.152939
R15292 gnd.n1370 gnd.n1369 0.152939
R15293 gnd.n1371 gnd.n1370 0.152939
R15294 gnd.n1375 gnd.n1371 0.152939
R15295 gnd.n1376 gnd.n1375 0.152939
R15296 gnd.n1377 gnd.n1376 0.152939
R15297 gnd.n1378 gnd.n1377 0.152939
R15298 gnd.n1382 gnd.n1378 0.152939
R15299 gnd.n1383 gnd.n1382 0.152939
R15300 gnd.n1384 gnd.n1383 0.152939
R15301 gnd.n1385 gnd.n1384 0.152939
R15302 gnd.n1608 gnd.n1385 0.152939
R15303 gnd.n1611 gnd.n1610 0.152939
R15304 gnd.n1612 gnd.n1611 0.152939
R15305 gnd.n1616 gnd.n1612 0.152939
R15306 gnd.n1617 gnd.n1616 0.152939
R15307 gnd.n1618 gnd.n1617 0.152939
R15308 gnd.n1619 gnd.n1618 0.152939
R15309 gnd.n1623 gnd.n1619 0.152939
R15310 gnd.n1624 gnd.n1623 0.152939
R15311 gnd.n1625 gnd.n1624 0.152939
R15312 gnd.n1626 gnd.n1625 0.152939
R15313 gnd.n1630 gnd.n1626 0.152939
R15314 gnd.n1631 gnd.n1630 0.152939
R15315 gnd.n1632 gnd.n1631 0.152939
R15316 gnd.n1633 gnd.n1632 0.152939
R15317 gnd.n1637 gnd.n1633 0.152939
R15318 gnd.n1638 gnd.n1637 0.152939
R15319 gnd.n1639 gnd.n1638 0.152939
R15320 gnd.n1640 gnd.n1639 0.152939
R15321 gnd.n1645 gnd.n1640 0.152939
R15322 gnd.n5699 gnd.n1645 0.152939
R15323 gnd.n4987 gnd.n4935 0.152939
R15324 gnd.n4937 gnd.n4935 0.152939
R15325 gnd.n4938 gnd.n4937 0.152939
R15326 gnd.n4939 gnd.n4938 0.152939
R15327 gnd.n4940 gnd.n4939 0.152939
R15328 gnd.n4941 gnd.n4940 0.152939
R15329 gnd.n4942 gnd.n4941 0.152939
R15330 gnd.n4943 gnd.n4942 0.152939
R15331 gnd.n4944 gnd.n4943 0.152939
R15332 gnd.n4945 gnd.n4944 0.152939
R15333 gnd.n4946 gnd.n4945 0.152939
R15334 gnd.n4947 gnd.n4946 0.152939
R15335 gnd.n4948 gnd.n4947 0.152939
R15336 gnd.n4949 gnd.n4948 0.152939
R15337 gnd.n4950 gnd.n4949 0.152939
R15338 gnd.n4951 gnd.n4950 0.152939
R15339 gnd.n4952 gnd.n4951 0.152939
R15340 gnd.n4953 gnd.n4952 0.152939
R15341 gnd.n4954 gnd.n4953 0.152939
R15342 gnd.n4956 gnd.n4954 0.152939
R15343 gnd.n4956 gnd.n4955 0.152939
R15344 gnd.n4955 gnd.n1899 0.152939
R15345 gnd.n5177 gnd.n1899 0.152939
R15346 gnd.n5178 gnd.n5177 0.152939
R15347 gnd.n5179 gnd.n5178 0.152939
R15348 gnd.n5180 gnd.n5179 0.152939
R15349 gnd.n5180 gnd.n1864 0.152939
R15350 gnd.n5220 gnd.n1864 0.152939
R15351 gnd.n5221 gnd.n5220 0.152939
R15352 gnd.n5222 gnd.n5221 0.152939
R15353 gnd.n5222 gnd.n1862 0.152939
R15354 gnd.n5228 gnd.n1862 0.152939
R15355 gnd.n5229 gnd.n5228 0.152939
R15356 gnd.n5230 gnd.n5229 0.152939
R15357 gnd.n5230 gnd.n1855 0.152939
R15358 gnd.n5244 gnd.n1855 0.152939
R15359 gnd.n5245 gnd.n5244 0.152939
R15360 gnd.n5246 gnd.n5245 0.152939
R15361 gnd.n5246 gnd.n1853 0.152939
R15362 gnd.n5252 gnd.n1853 0.152939
R15363 gnd.n5253 gnd.n5252 0.152939
R15364 gnd.n5254 gnd.n5253 0.152939
R15365 gnd.n5254 gnd.n1851 0.152939
R15366 gnd.n5283 gnd.n1851 0.152939
R15367 gnd.n5284 gnd.n5283 0.152939
R15368 gnd.n5285 gnd.n5284 0.152939
R15369 gnd.n5286 gnd.n5285 0.152939
R15370 gnd.n5288 gnd.n5286 0.152939
R15371 gnd.n5288 gnd.n5287 0.152939
R15372 gnd.n5287 gnd.n1843 0.152939
R15373 gnd.n1843 gnd.n1841 0.152939
R15374 gnd.n5323 gnd.n1841 0.152939
R15375 gnd.n5324 gnd.n5323 0.152939
R15376 gnd.n5325 gnd.n5324 0.152939
R15377 gnd.n5326 gnd.n5325 0.152939
R15378 gnd.n5327 gnd.n5326 0.152939
R15379 gnd.n5327 gnd.n1832 0.152939
R15380 gnd.n5376 gnd.n1832 0.152939
R15381 gnd.n5377 gnd.n5376 0.152939
R15382 gnd.n5378 gnd.n5377 0.152939
R15383 gnd.n5380 gnd.n5378 0.152939
R15384 gnd.n5380 gnd.n5379 0.152939
R15385 gnd.n5379 gnd.n1646 0.152939
R15386 gnd.n5698 gnd.n1646 0.152939
R15387 gnd.n5066 gnd.n4874 0.152939
R15388 gnd.n4877 gnd.n4874 0.152939
R15389 gnd.n4878 gnd.n4877 0.152939
R15390 gnd.n4879 gnd.n4878 0.152939
R15391 gnd.n4882 gnd.n4879 0.152939
R15392 gnd.n4883 gnd.n4882 0.152939
R15393 gnd.n4884 gnd.n4883 0.152939
R15394 gnd.n4885 gnd.n4884 0.152939
R15395 gnd.n4888 gnd.n4885 0.152939
R15396 gnd.n4889 gnd.n4888 0.152939
R15397 gnd.n4890 gnd.n4889 0.152939
R15398 gnd.n4891 gnd.n4890 0.152939
R15399 gnd.n4894 gnd.n4891 0.152939
R15400 gnd.n4895 gnd.n4894 0.152939
R15401 gnd.n4896 gnd.n4895 0.152939
R15402 gnd.n4897 gnd.n4896 0.152939
R15403 gnd.n4903 gnd.n4897 0.152939
R15404 gnd.n4904 gnd.n4903 0.152939
R15405 gnd.n4905 gnd.n4904 0.152939
R15406 gnd.n4906 gnd.n4905 0.152939
R15407 gnd.n4909 gnd.n4906 0.152939
R15408 gnd.n4910 gnd.n4909 0.152939
R15409 gnd.n4911 gnd.n4910 0.152939
R15410 gnd.n4912 gnd.n4911 0.152939
R15411 gnd.n4915 gnd.n4912 0.152939
R15412 gnd.n4916 gnd.n4915 0.152939
R15413 gnd.n4917 gnd.n4916 0.152939
R15414 gnd.n4918 gnd.n4917 0.152939
R15415 gnd.n4921 gnd.n4918 0.152939
R15416 gnd.n4922 gnd.n4921 0.152939
R15417 gnd.n4923 gnd.n4922 0.152939
R15418 gnd.n4924 gnd.n4923 0.152939
R15419 gnd.n4927 gnd.n4924 0.152939
R15420 gnd.n4928 gnd.n4927 0.152939
R15421 gnd.n4929 gnd.n4928 0.152939
R15422 gnd.n4994 gnd.n4929 0.152939
R15423 gnd.n4994 gnd.n4993 0.152939
R15424 gnd.n4993 gnd.n4992 0.152939
R15425 gnd.n5067 gnd.n1979 0.152939
R15426 gnd.n5081 gnd.n1979 0.152939
R15427 gnd.n5082 gnd.n5081 0.152939
R15428 gnd.n5083 gnd.n5082 0.152939
R15429 gnd.n5083 gnd.n1963 0.152939
R15430 gnd.n5097 gnd.n1963 0.152939
R15431 gnd.n5098 gnd.n5097 0.152939
R15432 gnd.n5099 gnd.n5098 0.152939
R15433 gnd.n5099 gnd.n1947 0.152939
R15434 gnd.n5113 gnd.n1947 0.152939
R15435 gnd.n5114 gnd.n5113 0.152939
R15436 gnd.n5115 gnd.n5114 0.152939
R15437 gnd.n5115 gnd.n1931 0.152939
R15438 gnd.n5129 gnd.n1931 0.152939
R15439 gnd.n5130 gnd.n5129 0.152939
R15440 gnd.n5131 gnd.n5130 0.152939
R15441 gnd.n5131 gnd.n1914 0.152939
R15442 gnd.n5153 gnd.n1914 0.152939
R15443 gnd.n5154 gnd.n5153 0.152939
R15444 gnd.n5155 gnd.n5154 0.152939
R15445 gnd.n5156 gnd.n5155 0.152939
R15446 gnd.n5156 gnd.n1878 0.152939
R15447 gnd.n5193 gnd.n1878 0.152939
R15448 gnd.n5194 gnd.n5193 0.152939
R15449 gnd.n5195 gnd.n5194 0.152939
R15450 gnd.n5195 gnd.n1764 0.152939
R15451 gnd.n5466 gnd.n1764 0.152939
R15452 gnd.n1802 gnd.n1801 0.152939
R15453 gnd.n3146 gnd.n2186 0.152939
R15454 gnd.n3147 gnd.n3146 0.152939
R15455 gnd.n3148 gnd.n3147 0.152939
R15456 gnd.n3148 gnd.n2180 0.152939
R15457 gnd.n3156 gnd.n2180 0.152939
R15458 gnd.n3157 gnd.n3156 0.152939
R15459 gnd.n3158 gnd.n3157 0.152939
R15460 gnd.n3158 gnd.n2174 0.152939
R15461 gnd.n3166 gnd.n2174 0.152939
R15462 gnd.n3167 gnd.n3166 0.152939
R15463 gnd.n3168 gnd.n3167 0.152939
R15464 gnd.n3168 gnd.n2168 0.152939
R15465 gnd.n3176 gnd.n2168 0.152939
R15466 gnd.n3177 gnd.n3176 0.152939
R15467 gnd.n3178 gnd.n3177 0.152939
R15468 gnd.n3178 gnd.n2162 0.152939
R15469 gnd.n3186 gnd.n2162 0.152939
R15470 gnd.n3187 gnd.n3186 0.152939
R15471 gnd.n3188 gnd.n3187 0.152939
R15472 gnd.n3188 gnd.n2156 0.152939
R15473 gnd.n3196 gnd.n2156 0.152939
R15474 gnd.n3197 gnd.n3196 0.152939
R15475 gnd.n3198 gnd.n3197 0.152939
R15476 gnd.n3198 gnd.n2150 0.152939
R15477 gnd.n3206 gnd.n2150 0.152939
R15478 gnd.n3207 gnd.n3206 0.152939
R15479 gnd.n3208 gnd.n3207 0.152939
R15480 gnd.n3208 gnd.n2144 0.152939
R15481 gnd.n3216 gnd.n2144 0.152939
R15482 gnd.n3217 gnd.n3216 0.152939
R15483 gnd.n3218 gnd.n3217 0.152939
R15484 gnd.n3218 gnd.n2138 0.152939
R15485 gnd.n3226 gnd.n2138 0.152939
R15486 gnd.n3227 gnd.n3226 0.152939
R15487 gnd.n3228 gnd.n3227 0.152939
R15488 gnd.n3228 gnd.n2132 0.152939
R15489 gnd.n3236 gnd.n2132 0.152939
R15490 gnd.n3237 gnd.n3236 0.152939
R15491 gnd.n3238 gnd.n3237 0.152939
R15492 gnd.n3238 gnd.n2126 0.152939
R15493 gnd.n3246 gnd.n2126 0.152939
R15494 gnd.n3247 gnd.n3246 0.152939
R15495 gnd.n3248 gnd.n3247 0.152939
R15496 gnd.n3248 gnd.n2120 0.152939
R15497 gnd.n3256 gnd.n2120 0.152939
R15498 gnd.n3257 gnd.n3256 0.152939
R15499 gnd.n3258 gnd.n3257 0.152939
R15500 gnd.n3258 gnd.n2114 0.152939
R15501 gnd.n3266 gnd.n2114 0.152939
R15502 gnd.n3267 gnd.n3266 0.152939
R15503 gnd.n3268 gnd.n3267 0.152939
R15504 gnd.n3268 gnd.n2108 0.152939
R15505 gnd.n3276 gnd.n2108 0.152939
R15506 gnd.n3277 gnd.n3276 0.152939
R15507 gnd.n3278 gnd.n3277 0.152939
R15508 gnd.n3278 gnd.n2102 0.152939
R15509 gnd.n3286 gnd.n2102 0.152939
R15510 gnd.n3287 gnd.n3286 0.152939
R15511 gnd.n3288 gnd.n3287 0.152939
R15512 gnd.n3288 gnd.n2096 0.152939
R15513 gnd.n3296 gnd.n2096 0.152939
R15514 gnd.n3297 gnd.n3296 0.152939
R15515 gnd.n3298 gnd.n3297 0.152939
R15516 gnd.n3298 gnd.n2090 0.152939
R15517 gnd.n3306 gnd.n2090 0.152939
R15518 gnd.n3307 gnd.n3306 0.152939
R15519 gnd.n3308 gnd.n3307 0.152939
R15520 gnd.n3308 gnd.n2084 0.152939
R15521 gnd.n3316 gnd.n2084 0.152939
R15522 gnd.n3317 gnd.n3316 0.152939
R15523 gnd.n3318 gnd.n3317 0.152939
R15524 gnd.n3318 gnd.n2078 0.152939
R15525 gnd.n3326 gnd.n2078 0.152939
R15526 gnd.n3327 gnd.n3326 0.152939
R15527 gnd.n3328 gnd.n3327 0.152939
R15528 gnd.n3328 gnd.n2072 0.152939
R15529 gnd.n3336 gnd.n2072 0.152939
R15530 gnd.n3337 gnd.n3336 0.152939
R15531 gnd.n3338 gnd.n3337 0.152939
R15532 gnd.n3338 gnd.n2066 0.152939
R15533 gnd.n3346 gnd.n2066 0.152939
R15534 gnd.n3347 gnd.n3346 0.152939
R15535 gnd.n3348 gnd.n3347 0.152939
R15536 gnd.n3350 gnd.n3348 0.152939
R15537 gnd.n6704 gnd.n6703 0.152939
R15538 gnd.n6703 gnd.n6702 0.152939
R15539 gnd.n6702 gnd.n6682 0.152939
R15540 gnd.n6698 gnd.n6682 0.152939
R15541 gnd.n6698 gnd.n6697 0.152939
R15542 gnd.n6697 gnd.n6696 0.152939
R15543 gnd.n6696 gnd.n6688 0.152939
R15544 gnd.n6688 gnd.n634 0.152939
R15545 gnd.n6813 gnd.n634 0.152939
R15546 gnd.n5821 gnd.n5820 0.152939
R15547 gnd.n5822 gnd.n5821 0.152939
R15548 gnd.n5822 gnd.n1292 0.152939
R15549 gnd.n5838 gnd.n1292 0.152939
R15550 gnd.n5839 gnd.n5838 0.152939
R15551 gnd.n5841 gnd.n5839 0.152939
R15552 gnd.n5841 gnd.n5840 0.152939
R15553 gnd.n5840 gnd.n1251 0.152939
R15554 gnd.n5994 gnd.n1251 0.152939
R15555 gnd.n5995 gnd.n5994 0.152939
R15556 gnd.n5996 gnd.n5995 0.152939
R15557 gnd.n5996 gnd.n1236 0.152939
R15558 gnd.n6010 gnd.n1236 0.152939
R15559 gnd.n6011 gnd.n6010 0.152939
R15560 gnd.n6012 gnd.n6011 0.152939
R15561 gnd.n6012 gnd.n1221 0.152939
R15562 gnd.n6026 gnd.n1221 0.152939
R15563 gnd.n6027 gnd.n6026 0.152939
R15564 gnd.n6028 gnd.n6027 0.152939
R15565 gnd.n6028 gnd.n1204 0.152939
R15566 gnd.n6043 gnd.n1204 0.152939
R15567 gnd.n6044 gnd.n6043 0.152939
R15568 gnd.n6046 gnd.n6044 0.152939
R15569 gnd.n6046 gnd.n6045 0.152939
R15570 gnd.n6045 gnd.n1098 0.152939
R15571 gnd.n6136 gnd.n1098 0.152939
R15572 gnd.n6137 gnd.n6136 0.152939
R15573 gnd.n6138 gnd.n6137 0.152939
R15574 gnd.n6138 gnd.n1083 0.152939
R15575 gnd.n6152 gnd.n1083 0.152939
R15576 gnd.n6153 gnd.n6152 0.152939
R15577 gnd.n6154 gnd.n6153 0.152939
R15578 gnd.n6154 gnd.n1069 0.152939
R15579 gnd.n6168 gnd.n1069 0.152939
R15580 gnd.n6169 gnd.n6168 0.152939
R15581 gnd.n6170 gnd.n6169 0.152939
R15582 gnd.n6170 gnd.n1053 0.152939
R15583 gnd.n6186 gnd.n1053 0.152939
R15584 gnd.n6187 gnd.n6186 0.152939
R15585 gnd.n6189 gnd.n6187 0.152939
R15586 gnd.n6189 gnd.n6188 0.152939
R15587 gnd.n6188 gnd.n1011 0.152939
R15588 gnd.n6441 gnd.n1011 0.152939
R15589 gnd.n6442 gnd.n6441 0.152939
R15590 gnd.n6443 gnd.n6442 0.152939
R15591 gnd.n6443 gnd.n995 0.152939
R15592 gnd.n6457 gnd.n995 0.152939
R15593 gnd.n6458 gnd.n6457 0.152939
R15594 gnd.n6459 gnd.n6458 0.152939
R15595 gnd.n6459 gnd.n980 0.152939
R15596 gnd.n6473 gnd.n980 0.152939
R15597 gnd.n6474 gnd.n6473 0.152939
R15598 gnd.n6475 gnd.n6474 0.152939
R15599 gnd.n6475 gnd.n965 0.152939
R15600 gnd.n6489 gnd.n965 0.152939
R15601 gnd.n6490 gnd.n6489 0.152939
R15602 gnd.n6491 gnd.n6490 0.152939
R15603 gnd.n6491 gnd.n950 0.152939
R15604 gnd.n6505 gnd.n950 0.152939
R15605 gnd.n6506 gnd.n6505 0.152939
R15606 gnd.n6507 gnd.n6506 0.152939
R15607 gnd.n6507 gnd.n934 0.152939
R15608 gnd.n6520 gnd.n934 0.152939
R15609 gnd.n6521 gnd.n6520 0.152939
R15610 gnd.n6529 gnd.n6521 0.152939
R15611 gnd.n6529 gnd.n6528 0.152939
R15612 gnd.n6528 gnd.n6527 0.152939
R15613 gnd.n6527 gnd.n6522 0.152939
R15614 gnd.n6522 gnd.n895 0.152939
R15615 gnd.n6587 gnd.n895 0.152939
R15616 gnd.n6587 gnd.n6586 0.152939
R15617 gnd.n6586 gnd.n6585 0.152939
R15618 gnd.n6585 gnd.n896 0.152939
R15619 gnd.n6581 gnd.n896 0.152939
R15620 gnd.n6581 gnd.n6580 0.152939
R15621 gnd.n6580 gnd.n651 0.152939
R15622 gnd.n6792 gnd.n651 0.152939
R15623 gnd.n6793 gnd.n6792 0.152939
R15624 gnd.n6795 gnd.n6793 0.152939
R15625 gnd.n6795 gnd.n6794 0.152939
R15626 gnd.n6794 gnd.n635 0.152939
R15627 gnd.n6812 gnd.n635 0.152939
R15628 gnd.n5785 gnd.n1339 0.152939
R15629 gnd.n5793 gnd.n1339 0.152939
R15630 gnd.n5794 gnd.n5793 0.152939
R15631 gnd.n5795 gnd.n5794 0.152939
R15632 gnd.n5795 gnd.n1335 0.152939
R15633 gnd.n5803 gnd.n1335 0.152939
R15634 gnd.n5804 gnd.n5803 0.152939
R15635 gnd.n5805 gnd.n5804 0.152939
R15636 gnd.n5805 gnd.n1308 0.152939
R15637 gnd.n5236 gnd.n1858 0.152939
R15638 gnd.n5237 gnd.n5236 0.152939
R15639 gnd.n5238 gnd.n5237 0.152939
R15640 gnd.n5238 gnd.n1809 0.152939
R15641 gnd.n5426 gnd.n1809 0.152939
R15642 gnd.n5426 gnd.n5425 0.152939
R15643 gnd.n5425 gnd.n5424 0.152939
R15644 gnd.n5424 gnd.n1810 0.152939
R15645 gnd.n5420 gnd.n1810 0.152939
R15646 gnd.n5420 gnd.n5419 0.152939
R15647 gnd.n5419 gnd.n5418 0.152939
R15648 gnd.n5418 gnd.n1814 0.152939
R15649 gnd.n5414 gnd.n1814 0.152939
R15650 gnd.n5414 gnd.n5413 0.152939
R15651 gnd.n5413 gnd.n5412 0.152939
R15652 gnd.n5412 gnd.n1818 0.152939
R15653 gnd.n5408 gnd.n1818 0.152939
R15654 gnd.n5408 gnd.n5407 0.152939
R15655 gnd.n5407 gnd.n5406 0.152939
R15656 gnd.n5406 gnd.n1822 0.152939
R15657 gnd.n5402 gnd.n1822 0.152939
R15658 gnd.n5402 gnd.n5401 0.152939
R15659 gnd.n5401 gnd.n5400 0.152939
R15660 gnd.n5400 gnd.n1826 0.152939
R15661 gnd.n5396 gnd.n1826 0.152939
R15662 gnd.n5396 gnd.n5395 0.152939
R15663 gnd.n5395 gnd.n5394 0.152939
R15664 gnd.n5394 gnd.n1830 0.152939
R15665 gnd.n5390 gnd.n1830 0.152939
R15666 gnd.n5390 gnd.n5389 0.152939
R15667 gnd.n5389 gnd.n1341 0.152939
R15668 gnd.n5687 gnd.n5675 0.152939
R15669 gnd.n5683 gnd.n5675 0.152939
R15670 gnd.n5683 gnd.n5682 0.152939
R15671 gnd.n5682 gnd.n5681 0.152939
R15672 gnd.n5681 gnd.n1284 0.152939
R15673 gnd.n5847 gnd.n1284 0.152939
R15674 gnd.n5848 gnd.n5847 0.152939
R15675 gnd.n5849 gnd.n5848 0.152939
R15676 gnd.n5849 gnd.n1280 0.152939
R15677 gnd.n5856 gnd.n1280 0.152939
R15678 gnd.n5857 gnd.n5856 0.152939
R15679 gnd.n5964 gnd.n5857 0.152939
R15680 gnd.n5964 gnd.n5963 0.152939
R15681 gnd.n5963 gnd.n5962 0.152939
R15682 gnd.n5962 gnd.n5858 0.152939
R15683 gnd.n5958 gnd.n5858 0.152939
R15684 gnd.n5958 gnd.n5957 0.152939
R15685 gnd.n5957 gnd.n5956 0.152939
R15686 gnd.n5956 gnd.n5862 0.152939
R15687 gnd.n5952 gnd.n5862 0.152939
R15688 gnd.n5952 gnd.n5951 0.152939
R15689 gnd.n5951 gnd.n1196 0.152939
R15690 gnd.n6052 gnd.n1196 0.152939
R15691 gnd.n6053 gnd.n6052 0.152939
R15692 gnd.n6054 gnd.n6053 0.152939
R15693 gnd.n6054 gnd.n1192 0.152939
R15694 gnd.n6059 gnd.n1192 0.152939
R15695 gnd.n6060 gnd.n6059 0.152939
R15696 gnd.n6061 gnd.n6060 0.152939
R15697 gnd.n6061 gnd.n1190 0.152939
R15698 gnd.n6066 gnd.n1190 0.152939
R15699 gnd.n6067 gnd.n6066 0.152939
R15700 gnd.n6068 gnd.n6067 0.152939
R15701 gnd.n6068 gnd.n1188 0.152939
R15702 gnd.n6073 gnd.n1188 0.152939
R15703 gnd.n6074 gnd.n6073 0.152939
R15704 gnd.n6076 gnd.n6074 0.152939
R15705 gnd.n6076 gnd.n6075 0.152939
R15706 gnd.n6075 gnd.n1046 0.152939
R15707 gnd.n6195 gnd.n1046 0.152939
R15708 gnd.n6196 gnd.n6195 0.152939
R15709 gnd.n6197 gnd.n6196 0.152939
R15710 gnd.n6197 gnd.n1042 0.152939
R15711 gnd.n6202 gnd.n1042 0.152939
R15712 gnd.n6203 gnd.n6202 0.152939
R15713 gnd.n6411 gnd.n6203 0.152939
R15714 gnd.n6411 gnd.n6410 0.152939
R15715 gnd.n6410 gnd.n6409 0.152939
R15716 gnd.n6409 gnd.n6204 0.152939
R15717 gnd.n6405 gnd.n6204 0.152939
R15718 gnd.n6405 gnd.n6404 0.152939
R15719 gnd.n6404 gnd.n6403 0.152939
R15720 gnd.n6403 gnd.n6208 0.152939
R15721 gnd.n6399 gnd.n6208 0.152939
R15722 gnd.n6399 gnd.n6398 0.152939
R15723 gnd.n6398 gnd.n6397 0.152939
R15724 gnd.n6397 gnd.n6212 0.152939
R15725 gnd.n6393 gnd.n6212 0.152939
R15726 gnd.n6393 gnd.n6392 0.152939
R15727 gnd.n6392 gnd.n6391 0.152939
R15728 gnd.n6391 gnd.n6216 0.152939
R15729 gnd.n6387 gnd.n6216 0.152939
R15730 gnd.n6387 gnd.n6386 0.152939
R15731 gnd.n6386 gnd.n6385 0.152939
R15732 gnd.n6385 gnd.n6220 0.152939
R15733 gnd.n6220 gnd.n916 0.152939
R15734 gnd.n6545 gnd.n916 0.152939
R15735 gnd.n6546 gnd.n6545 0.152939
R15736 gnd.n6548 gnd.n6546 0.152939
R15737 gnd.n6548 gnd.n6547 0.152939
R15738 gnd.n6547 gnd.n875 0.152939
R15739 gnd.n6603 gnd.n875 0.152939
R15740 gnd.n6604 gnd.n6603 0.152939
R15741 gnd.n6605 gnd.n6604 0.152939
R15742 gnd.n6605 gnd.n872 0.152939
R15743 gnd.n6610 gnd.n872 0.152939
R15744 gnd.n6611 gnd.n6610 0.152939
R15745 gnd.n6765 gnd.n6611 0.152939
R15746 gnd.n6765 gnd.n6764 0.152939
R15747 gnd.n6764 gnd.n6763 0.152939
R15748 gnd.n6763 gnd.n6612 0.152939
R15749 gnd.n6615 gnd.n6612 0.152939
R15750 gnd.n7058 gnd.n477 0.152939
R15751 gnd.n7059 gnd.n7058 0.152939
R15752 gnd.n7060 gnd.n7059 0.152939
R15753 gnd.n7060 gnd.n459 0.152939
R15754 gnd.n7074 gnd.n459 0.152939
R15755 gnd.n7075 gnd.n7074 0.152939
R15756 gnd.n7076 gnd.n7075 0.152939
R15757 gnd.n7076 gnd.n443 0.152939
R15758 gnd.n7090 gnd.n443 0.152939
R15759 gnd.n7091 gnd.n7090 0.152939
R15760 gnd.n7092 gnd.n7091 0.152939
R15761 gnd.n7092 gnd.n425 0.152939
R15762 gnd.n7106 gnd.n425 0.152939
R15763 gnd.n7107 gnd.n7106 0.152939
R15764 gnd.n7108 gnd.n7107 0.152939
R15765 gnd.n7108 gnd.n409 0.152939
R15766 gnd.n7122 gnd.n409 0.152939
R15767 gnd.n7123 gnd.n7122 0.152939
R15768 gnd.n7127 gnd.n7123 0.152939
R15769 gnd.n7127 gnd.n7126 0.152939
R15770 gnd.n7126 gnd.n7125 0.152939
R15771 gnd.n7125 gnd.n377 0.152939
R15772 gnd.n7178 gnd.n377 0.152939
R15773 gnd.n7178 gnd.n7177 0.152939
R15774 gnd.n7177 gnd.n7176 0.152939
R15775 gnd.n7176 gnd.n378 0.152939
R15776 gnd.n7172 gnd.n378 0.152939
R15777 gnd.n7172 gnd.n316 0.152939
R15778 gnd.n7317 gnd.n316 0.152939
R15779 gnd.n7317 gnd.n7316 0.152939
R15780 gnd.n7316 gnd.n7315 0.152939
R15781 gnd.n7315 gnd.n317 0.152939
R15782 gnd.n7311 gnd.n317 0.152939
R15783 gnd.n7311 gnd.n7310 0.152939
R15784 gnd.n7310 gnd.n7309 0.152939
R15785 gnd.n7309 gnd.n322 0.152939
R15786 gnd.n322 gnd.n292 0.152939
R15787 gnd.n7332 gnd.n292 0.152939
R15788 gnd.n7333 gnd.n7332 0.152939
R15789 gnd.n7334 gnd.n7333 0.152939
R15790 gnd.n7334 gnd.n276 0.152939
R15791 gnd.n7348 gnd.n276 0.152939
R15792 gnd.n7349 gnd.n7348 0.152939
R15793 gnd.n7350 gnd.n7349 0.152939
R15794 gnd.n7350 gnd.n262 0.152939
R15795 gnd.n7364 gnd.n262 0.152939
R15796 gnd.n7365 gnd.n7364 0.152939
R15797 gnd.n7366 gnd.n7365 0.152939
R15798 gnd.n7366 gnd.n246 0.152939
R15799 gnd.n7380 gnd.n246 0.152939
R15800 gnd.n7381 gnd.n7380 0.152939
R15801 gnd.n7382 gnd.n7381 0.152939
R15802 gnd.n7382 gnd.n231 0.152939
R15803 gnd.n7396 gnd.n231 0.152939
R15804 gnd.n7397 gnd.n7396 0.152939
R15805 gnd.n7398 gnd.n7397 0.152939
R15806 gnd.n7398 gnd.n216 0.152939
R15807 gnd.n7412 gnd.n216 0.152939
R15808 gnd.n7413 gnd.n7412 0.152939
R15809 gnd.n7482 gnd.n7413 0.152939
R15810 gnd.n7482 gnd.n7481 0.152939
R15811 gnd.n7481 gnd.n7480 0.152939
R15812 gnd.n7480 gnd.n7414 0.152939
R15813 gnd.n7476 gnd.n7414 0.152939
R15814 gnd.n7475 gnd.n7416 0.152939
R15815 gnd.n7471 gnd.n7416 0.152939
R15816 gnd.n7471 gnd.n7470 0.152939
R15817 gnd.n7470 gnd.n7469 0.152939
R15818 gnd.n7469 gnd.n7422 0.152939
R15819 gnd.n7465 gnd.n7422 0.152939
R15820 gnd.n7465 gnd.n7464 0.152939
R15821 gnd.n7464 gnd.n7463 0.152939
R15822 gnd.n7463 gnd.n7430 0.152939
R15823 gnd.n7459 gnd.n7430 0.152939
R15824 gnd.n7459 gnd.n7458 0.152939
R15825 gnd.n7458 gnd.n7457 0.152939
R15826 gnd.n7457 gnd.n7438 0.152939
R15827 gnd.n7453 gnd.n7438 0.152939
R15828 gnd.n7453 gnd.n7452 0.152939
R15829 gnd.n7452 gnd.n7451 0.152939
R15830 gnd.n7451 gnd.n117 0.152939
R15831 gnd.n7577 gnd.n117 0.152939
R15832 gnd.n6971 gnd.n6970 0.152939
R15833 gnd.n6970 gnd.n6969 0.152939
R15834 gnd.n6969 gnd.n567 0.152939
R15835 gnd.n6965 gnd.n567 0.152939
R15836 gnd.n6965 gnd.n6964 0.152939
R15837 gnd.n6964 gnd.n6963 0.152939
R15838 gnd.n6963 gnd.n571 0.152939
R15839 gnd.n6959 gnd.n571 0.152939
R15840 gnd.n6959 gnd.n6958 0.152939
R15841 gnd.n6958 gnd.n6957 0.152939
R15842 gnd.n6957 gnd.n575 0.152939
R15843 gnd.n6953 gnd.n575 0.152939
R15844 gnd.n6953 gnd.n6952 0.152939
R15845 gnd.n6952 gnd.n6951 0.152939
R15846 gnd.n6951 gnd.n579 0.152939
R15847 gnd.n6947 gnd.n579 0.152939
R15848 gnd.n6947 gnd.n6946 0.152939
R15849 gnd.n6946 gnd.n6945 0.152939
R15850 gnd.n6945 gnd.n583 0.152939
R15851 gnd.n6941 gnd.n583 0.152939
R15852 gnd.n6941 gnd.n6940 0.152939
R15853 gnd.n6940 gnd.n383 0.152939
R15854 gnd.n7163 gnd.n383 0.152939
R15855 gnd.n7164 gnd.n7163 0.152939
R15856 gnd.n7166 gnd.n7164 0.152939
R15857 gnd.n7166 gnd.n7165 0.152939
R15858 gnd.n7165 gnd.n354 0.152939
R15859 gnd.n7208 gnd.n354 0.152939
R15860 gnd.n7208 gnd.n7207 0.152939
R15861 gnd.n7207 gnd.n7206 0.152939
R15862 gnd.n7206 gnd.n75 0.152939
R15863 gnd.n7626 gnd.n75 0.152939
R15864 gnd.n7626 gnd.n7625 0.152939
R15865 gnd.n7625 gnd.n77 0.152939
R15866 gnd.n7621 gnd.n77 0.152939
R15867 gnd.n7621 gnd.n7620 0.152939
R15868 gnd.n7620 gnd.n7619 0.152939
R15869 gnd.n7619 gnd.n82 0.152939
R15870 gnd.n7615 gnd.n82 0.152939
R15871 gnd.n7615 gnd.n7614 0.152939
R15872 gnd.n7614 gnd.n7613 0.152939
R15873 gnd.n7613 gnd.n87 0.152939
R15874 gnd.n7609 gnd.n87 0.152939
R15875 gnd.n7609 gnd.n7608 0.152939
R15876 gnd.n7608 gnd.n7607 0.152939
R15877 gnd.n7607 gnd.n92 0.152939
R15878 gnd.n7603 gnd.n92 0.152939
R15879 gnd.n7603 gnd.n7602 0.152939
R15880 gnd.n7602 gnd.n7601 0.152939
R15881 gnd.n7601 gnd.n97 0.152939
R15882 gnd.n7597 gnd.n97 0.152939
R15883 gnd.n7597 gnd.n7596 0.152939
R15884 gnd.n7596 gnd.n7595 0.152939
R15885 gnd.n7595 gnd.n102 0.152939
R15886 gnd.n7591 gnd.n102 0.152939
R15887 gnd.n7591 gnd.n7590 0.152939
R15888 gnd.n7590 gnd.n7589 0.152939
R15889 gnd.n7589 gnd.n107 0.152939
R15890 gnd.n7585 gnd.n107 0.152939
R15891 gnd.n7585 gnd.n7584 0.152939
R15892 gnd.n7584 gnd.n7583 0.152939
R15893 gnd.n7583 gnd.n112 0.152939
R15894 gnd.n7579 gnd.n112 0.152939
R15895 gnd.n7579 gnd.n7578 0.152939
R15896 gnd.n6704 gnd.n566 0.151415
R15897 gnd.n5785 gnd.n5784 0.151415
R15898 gnd.n5209 gnd.n5207 0.145814
R15899 gnd.n5209 gnd.n1858 0.145814
R15900 gnd.n347 gnd.n300 0.130073
R15901 gnd.n1801 gnd.n1765 0.130073
R15902 gnd.n4189 gnd.n3535 0.0767195
R15903 gnd.n4189 gnd.n4188 0.0767195
R15904 gnd.n5689 gnd.n5688 0.063
R15905 gnd.n6620 gnd.n6619 0.063
R15906 gnd.n4719 gnd.n2029 0.0477147
R15907 gnd.n3979 gnd.n3867 0.0442063
R15908 gnd.n3980 gnd.n3979 0.0442063
R15909 gnd.n3981 gnd.n3980 0.0442063
R15910 gnd.n3981 gnd.n3856 0.0442063
R15911 gnd.n3995 gnd.n3856 0.0442063
R15912 gnd.n3996 gnd.n3995 0.0442063
R15913 gnd.n3997 gnd.n3996 0.0442063
R15914 gnd.n3997 gnd.n3843 0.0442063
R15915 gnd.n4041 gnd.n3843 0.0442063
R15916 gnd.n4042 gnd.n4041 0.0442063
R15917 gnd.n4044 gnd.n3777 0.0344674
R15918 gnd.n6708 gnd.n6676 0.0344674
R15919 gnd.n5783 gnd.n5782 0.0344674
R15920 gnd.n4064 gnd.n4063 0.0269946
R15921 gnd.n4066 gnd.n4065 0.0269946
R15922 gnd.n3772 gnd.n3770 0.0269946
R15923 gnd.n4076 gnd.n4074 0.0269946
R15924 gnd.n4075 gnd.n3751 0.0269946
R15925 gnd.n4095 gnd.n4094 0.0269946
R15926 gnd.n4097 gnd.n4096 0.0269946
R15927 gnd.n3746 gnd.n3745 0.0269946
R15928 gnd.n4107 gnd.n3741 0.0269946
R15929 gnd.n4106 gnd.n3743 0.0269946
R15930 gnd.n3742 gnd.n3722 0.0269946
R15931 gnd.n4133 gnd.n3723 0.0269946
R15932 gnd.n4132 gnd.n3724 0.0269946
R15933 gnd.n4152 gnd.n3708 0.0269946
R15934 gnd.n4154 gnd.n4153 0.0269946
R15935 gnd.n4155 gnd.n3688 0.0269946
R15936 gnd.n4156 gnd.n3689 0.0269946
R15937 gnd.n4157 gnd.n3690 0.0269946
R15938 gnd.n3692 gnd.n3691 0.0269946
R15939 gnd.n3529 gnd.n3527 0.0269946
R15940 gnd.n4201 gnd.n4199 0.0269946
R15941 gnd.n4200 gnd.n3511 0.0269946
R15942 gnd.n4220 gnd.n4219 0.0269946
R15943 gnd.n4222 gnd.n4221 0.0269946
R15944 gnd.n3506 gnd.n3504 0.0269946
R15945 gnd.n4232 gnd.n4230 0.0269946
R15946 gnd.n4231 gnd.n3486 0.0269946
R15947 gnd.n4251 gnd.n4250 0.0269946
R15948 gnd.n4253 gnd.n4252 0.0269946
R15949 gnd.n3480 gnd.n3478 0.0269946
R15950 gnd.n4263 gnd.n4261 0.0269946
R15951 gnd.n4262 gnd.n3459 0.0269946
R15952 gnd.n4282 gnd.n4281 0.0269946
R15953 gnd.n4284 gnd.n4283 0.0269946
R15954 gnd.n3454 gnd.n3452 0.0269946
R15955 gnd.n4294 gnd.n4292 0.0269946
R15956 gnd.n4293 gnd.n3435 0.0269946
R15957 gnd.n4313 gnd.n4312 0.0269946
R15958 gnd.n4315 gnd.n4314 0.0269946
R15959 gnd.n3430 gnd.n3428 0.0269946
R15960 gnd.n4325 gnd.n4323 0.0269946
R15961 gnd.n4324 gnd.n3409 0.0269946
R15962 gnd.n4344 gnd.n4343 0.0269946
R15963 gnd.n4346 gnd.n4345 0.0269946
R15964 gnd.n3404 gnd.n3402 0.0269946
R15965 gnd.n4356 gnd.n4354 0.0269946
R15966 gnd.n4355 gnd.n3384 0.0269946
R15967 gnd.n4375 gnd.n4374 0.0269946
R15968 gnd.n3378 gnd.n3376 0.0269946
R15969 gnd.n4643 gnd.n4641 0.0269946
R15970 gnd.n4642 gnd.n3358 0.0269946
R15971 gnd.n4661 gnd.n4660 0.0269946
R15972 gnd.n6619 gnd.n6617 0.0246168
R15973 gnd.n5688 gnd.n5674 0.0246168
R15974 gnd.n7217 gnd.n300 0.0233659
R15975 gnd.n3349 gnd.n1765 0.0233659
R15976 gnd.n4044 gnd.n4043 0.0202011
R15977 gnd.n6756 gnd.n6617 0.0174837
R15978 gnd.n6756 gnd.n6755 0.0174837
R15979 gnd.n6755 gnd.n6618 0.0174837
R15980 gnd.n6752 gnd.n6618 0.0174837
R15981 gnd.n6752 gnd.n6751 0.0174837
R15982 gnd.n6751 gnd.n6629 0.0174837
R15983 gnd.n6748 gnd.n6629 0.0174837
R15984 gnd.n6748 gnd.n6747 0.0174837
R15985 gnd.n6747 gnd.n6635 0.0174837
R15986 gnd.n6744 gnd.n6635 0.0174837
R15987 gnd.n6744 gnd.n6743 0.0174837
R15988 gnd.n6743 gnd.n6639 0.0174837
R15989 gnd.n6740 gnd.n6639 0.0174837
R15990 gnd.n6740 gnd.n6739 0.0174837
R15991 gnd.n6739 gnd.n6643 0.0174837
R15992 gnd.n6736 gnd.n6643 0.0174837
R15993 gnd.n6736 gnd.n6735 0.0174837
R15994 gnd.n6735 gnd.n6649 0.0174837
R15995 gnd.n6732 gnd.n6649 0.0174837
R15996 gnd.n6732 gnd.n6731 0.0174837
R15997 gnd.n6731 gnd.n6655 0.0174837
R15998 gnd.n6728 gnd.n6655 0.0174837
R15999 gnd.n6728 gnd.n6727 0.0174837
R16000 gnd.n6727 gnd.n6659 0.0174837
R16001 gnd.n6724 gnd.n6659 0.0174837
R16002 gnd.n6724 gnd.n6723 0.0174837
R16003 gnd.n6723 gnd.n6663 0.0174837
R16004 gnd.n6720 gnd.n6663 0.0174837
R16005 gnd.n6720 gnd.n6719 0.0174837
R16006 gnd.n6719 gnd.n6669 0.0174837
R16007 gnd.n6716 gnd.n6669 0.0174837
R16008 gnd.n6716 gnd.n6715 0.0174837
R16009 gnd.n6715 gnd.n6675 0.0174837
R16010 gnd.n6709 gnd.n6675 0.0174837
R16011 gnd.n6709 gnd.n6708 0.0174837
R16012 gnd.n5674 gnd.n5574 0.0174837
R16013 gnd.n5671 gnd.n5574 0.0174837
R16014 gnd.n5671 gnd.n5670 0.0174837
R16015 gnd.n5670 gnd.n5580 0.0174837
R16016 gnd.n5667 gnd.n5580 0.0174837
R16017 gnd.n5667 gnd.n5666 0.0174837
R16018 gnd.n5666 gnd.n5586 0.0174837
R16019 gnd.n5663 gnd.n5586 0.0174837
R16020 gnd.n5663 gnd.n5662 0.0174837
R16021 gnd.n5662 gnd.n5592 0.0174837
R16022 gnd.n5659 gnd.n5592 0.0174837
R16023 gnd.n5659 gnd.n5658 0.0174837
R16024 gnd.n5658 gnd.n5598 0.0174837
R16025 gnd.n5655 gnd.n5598 0.0174837
R16026 gnd.n5655 gnd.n5654 0.0174837
R16027 gnd.n5654 gnd.n5605 0.0174837
R16028 gnd.n5651 gnd.n5605 0.0174837
R16029 gnd.n5651 gnd.n5650 0.0174837
R16030 gnd.n5650 gnd.n5609 0.0174837
R16031 gnd.n5647 gnd.n5609 0.0174837
R16032 gnd.n5647 gnd.n5646 0.0174837
R16033 gnd.n5646 gnd.n5615 0.0174837
R16034 gnd.n5643 gnd.n5615 0.0174837
R16035 gnd.n5643 gnd.n5642 0.0174837
R16036 gnd.n5642 gnd.n5621 0.0174837
R16037 gnd.n5639 gnd.n5621 0.0174837
R16038 gnd.n5639 gnd.n5638 0.0174837
R16039 gnd.n5638 gnd.n5631 0.0174837
R16040 gnd.n5635 gnd.n5631 0.0174837
R16041 gnd.n5635 gnd.n5634 0.0174837
R16042 gnd.n5634 gnd.n1346 0.0174837
R16043 gnd.n5776 gnd.n1346 0.0174837
R16044 gnd.n5777 gnd.n5776 0.0174837
R16045 gnd.n5777 gnd.n1342 0.0174837
R16046 gnd.n5782 gnd.n1342 0.0174837
R16047 gnd.n4043 gnd.n4042 0.0148637
R16048 gnd.n4632 gnd.n4376 0.0144266
R16049 gnd.n4633 gnd.n4632 0.0130679
R16050 gnd.n4063 gnd.n3777 0.00797283
R16051 gnd.n4065 gnd.n4064 0.00797283
R16052 gnd.n4066 gnd.n3772 0.00797283
R16053 gnd.n4074 gnd.n3770 0.00797283
R16054 gnd.n4076 gnd.n4075 0.00797283
R16055 gnd.n4094 gnd.n3751 0.00797283
R16056 gnd.n4096 gnd.n4095 0.00797283
R16057 gnd.n4097 gnd.n3746 0.00797283
R16058 gnd.n3745 gnd.n3741 0.00797283
R16059 gnd.n4107 gnd.n4106 0.00797283
R16060 gnd.n3743 gnd.n3742 0.00797283
R16061 gnd.n3723 gnd.n3722 0.00797283
R16062 gnd.n4133 gnd.n4132 0.00797283
R16063 gnd.n3724 gnd.n3708 0.00797283
R16064 gnd.n4153 gnd.n4152 0.00797283
R16065 gnd.n4155 gnd.n4154 0.00797283
R16066 gnd.n4156 gnd.n3688 0.00797283
R16067 gnd.n4157 gnd.n3689 0.00797283
R16068 gnd.n3691 gnd.n3690 0.00797283
R16069 gnd.n3692 gnd.n3529 0.00797283
R16070 gnd.n4199 gnd.n3527 0.00797283
R16071 gnd.n4201 gnd.n4200 0.00797283
R16072 gnd.n4219 gnd.n3511 0.00797283
R16073 gnd.n4221 gnd.n4220 0.00797283
R16074 gnd.n4222 gnd.n3506 0.00797283
R16075 gnd.n4230 gnd.n3504 0.00797283
R16076 gnd.n4232 gnd.n4231 0.00797283
R16077 gnd.n4250 gnd.n3486 0.00797283
R16078 gnd.n4252 gnd.n4251 0.00797283
R16079 gnd.n4253 gnd.n3480 0.00797283
R16080 gnd.n4261 gnd.n3478 0.00797283
R16081 gnd.n4263 gnd.n4262 0.00797283
R16082 gnd.n4281 gnd.n3459 0.00797283
R16083 gnd.n4283 gnd.n4282 0.00797283
R16084 gnd.n4284 gnd.n3454 0.00797283
R16085 gnd.n4292 gnd.n3452 0.00797283
R16086 gnd.n4294 gnd.n4293 0.00797283
R16087 gnd.n4312 gnd.n3435 0.00797283
R16088 gnd.n4314 gnd.n4313 0.00797283
R16089 gnd.n4315 gnd.n3430 0.00797283
R16090 gnd.n4323 gnd.n3428 0.00797283
R16091 gnd.n4325 gnd.n4324 0.00797283
R16092 gnd.n4343 gnd.n3409 0.00797283
R16093 gnd.n4345 gnd.n4344 0.00797283
R16094 gnd.n4346 gnd.n3404 0.00797283
R16095 gnd.n4354 gnd.n3402 0.00797283
R16096 gnd.n4356 gnd.n4355 0.00797283
R16097 gnd.n4374 gnd.n3384 0.00797283
R16098 gnd.n4376 gnd.n4375 0.00797283
R16099 gnd.n4633 gnd.n3378 0.00797283
R16100 gnd.n4641 gnd.n3376 0.00797283
R16101 gnd.n4643 gnd.n4642 0.00797283
R16102 gnd.n4660 gnd.n3358 0.00797283
R16103 gnd.n4661 gnd.n2029 0.00797283
R16104 gnd.n333 gnd.n317 0.00433921
R16105 gnd.n5228 gnd.n1861 0.00433921
R16106 gnd.n6676 gnd.n566 0.000839674
R16107 gnd.n5784 gnd.n5783 0.000839674
R16108 a_n6972_8799.n140 a_n6972_8799.t54 490.524
R16109 a_n6972_8799.n151 a_n6972_8799.t63 490.524
R16110 a_n6972_8799.n163 a_n6972_8799.t102 490.524
R16111 a_n6972_8799.n106 a_n6972_8799.t99 490.524
R16112 a_n6972_8799.n117 a_n6972_8799.t108 490.524
R16113 a_n6972_8799.n129 a_n6972_8799.t101 490.524
R16114 a_n6972_8799.n31 a_n6972_8799.t70 484.3
R16115 a_n6972_8799.n146 a_n6972_8799.t58 464.166
R16116 a_n6972_8799.n145 a_n6972_8799.t103 464.166
R16117 a_n6972_8799.n136 a_n6972_8799.t80 464.166
R16118 a_n6972_8799.n144 a_n6972_8799.t78 464.166
R16119 a_n6972_8799.n143 a_n6972_8799.t42 464.166
R16120 a_n6972_8799.n137 a_n6972_8799.t84 464.166
R16121 a_n6972_8799.n142 a_n6972_8799.t83 464.166
R16122 a_n6972_8799.n141 a_n6972_8799.t44 464.166
R16123 a_n6972_8799.n138 a_n6972_8799.t43 464.166
R16124 a_n6972_8799.n139 a_n6972_8799.t97 464.166
R16125 a_n6972_8799.n40 a_n6972_8799.t77 484.3
R16126 a_n6972_8799.n157 a_n6972_8799.t64 464.166
R16127 a_n6972_8799.n156 a_n6972_8799.t111 464.166
R16128 a_n6972_8799.n147 a_n6972_8799.t90 464.166
R16129 a_n6972_8799.n155 a_n6972_8799.t89 464.166
R16130 a_n6972_8799.n154 a_n6972_8799.t49 464.166
R16131 a_n6972_8799.n148 a_n6972_8799.t93 464.166
R16132 a_n6972_8799.n153 a_n6972_8799.t92 464.166
R16133 a_n6972_8799.n152 a_n6972_8799.t51 464.166
R16134 a_n6972_8799.n149 a_n6972_8799.t50 464.166
R16135 a_n6972_8799.n150 a_n6972_8799.t106 464.166
R16136 a_n6972_8799.n49 a_n6972_8799.t96 484.3
R16137 a_n6972_8799.n169 a_n6972_8799.t56 464.166
R16138 a_n6972_8799.n168 a_n6972_8799.t82 464.166
R16139 a_n6972_8799.n159 a_n6972_8799.t46 464.166
R16140 a_n6972_8799.n167 a_n6972_8799.t59 464.166
R16141 a_n6972_8799.n166 a_n6972_8799.t109 464.166
R16142 a_n6972_8799.n160 a_n6972_8799.t88 464.166
R16143 a_n6972_8799.n165 a_n6972_8799.t105 464.166
R16144 a_n6972_8799.n164 a_n6972_8799.t76 464.166
R16145 a_n6972_8799.n161 a_n6972_8799.t91 464.166
R16146 a_n6972_8799.n162 a_n6972_8799.t53 464.166
R16147 a_n6972_8799.n105 a_n6972_8799.t68 464.166
R16148 a_n6972_8799.n104 a_n6972_8799.t69 464.166
R16149 a_n6972_8799.n107 a_n6972_8799.t86 464.166
R16150 a_n6972_8799.n103 a_n6972_8799.t61 464.166
R16151 a_n6972_8799.n108 a_n6972_8799.t62 464.166
R16152 a_n6972_8799.n109 a_n6972_8799.t85 464.166
R16153 a_n6972_8799.n102 a_n6972_8799.t40 464.166
R16154 a_n6972_8799.n110 a_n6972_8799.t60 464.166
R16155 a_n6972_8799.n101 a_n6972_8799.t72 464.166
R16156 a_n6972_8799.n111 a_n6972_8799.t100 464.166
R16157 a_n6972_8799.n116 a_n6972_8799.t73 464.166
R16158 a_n6972_8799.n115 a_n6972_8799.t74 464.166
R16159 a_n6972_8799.n118 a_n6972_8799.t98 464.166
R16160 a_n6972_8799.n114 a_n6972_8799.t66 464.166
R16161 a_n6972_8799.n119 a_n6972_8799.t67 464.166
R16162 a_n6972_8799.n120 a_n6972_8799.t94 464.166
R16163 a_n6972_8799.n113 a_n6972_8799.t47 464.166
R16164 a_n6972_8799.n121 a_n6972_8799.t65 464.166
R16165 a_n6972_8799.n112 a_n6972_8799.t79 464.166
R16166 a_n6972_8799.n122 a_n6972_8799.t110 464.166
R16167 a_n6972_8799.n128 a_n6972_8799.t52 464.166
R16168 a_n6972_8799.n127 a_n6972_8799.t41 464.166
R16169 a_n6972_8799.n130 a_n6972_8799.t75 464.166
R16170 a_n6972_8799.n126 a_n6972_8799.t104 464.166
R16171 a_n6972_8799.n131 a_n6972_8799.t87 464.166
R16172 a_n6972_8799.n132 a_n6972_8799.t107 464.166
R16173 a_n6972_8799.n125 a_n6972_8799.t71 464.166
R16174 a_n6972_8799.n133 a_n6972_8799.t45 464.166
R16175 a_n6972_8799.n124 a_n6972_8799.t81 464.166
R16176 a_n6972_8799.n134 a_n6972_8799.t55 464.166
R16177 a_n6972_8799.n39 a_n6972_8799.n38 75.3623
R16178 a_n6972_8799.n37 a_n6972_8799.n24 70.3058
R16179 a_n6972_8799.n24 a_n6972_8799.n36 70.1674
R16180 a_n6972_8799.n36 a_n6972_8799.n137 20.9683
R16181 a_n6972_8799.n35 a_n6972_8799.n25 75.0448
R16182 a_n6972_8799.n143 a_n6972_8799.n35 11.2134
R16183 a_n6972_8799.n34 a_n6972_8799.n25 80.4688
R16184 a_n6972_8799.n27 a_n6972_8799.n33 74.73
R16185 a_n6972_8799.n32 a_n6972_8799.n27 70.1674
R16186 a_n6972_8799.n146 a_n6972_8799.n32 20.9683
R16187 a_n6972_8799.n26 a_n6972_8799.n31 70.5844
R16188 a_n6972_8799.n48 a_n6972_8799.n47 75.3623
R16189 a_n6972_8799.n46 a_n6972_8799.n20 70.3058
R16190 a_n6972_8799.n20 a_n6972_8799.n45 70.1674
R16191 a_n6972_8799.n45 a_n6972_8799.n148 20.9683
R16192 a_n6972_8799.n44 a_n6972_8799.n21 75.0448
R16193 a_n6972_8799.n154 a_n6972_8799.n44 11.2134
R16194 a_n6972_8799.n43 a_n6972_8799.n21 80.4688
R16195 a_n6972_8799.n23 a_n6972_8799.n42 74.73
R16196 a_n6972_8799.n41 a_n6972_8799.n23 70.1674
R16197 a_n6972_8799.n157 a_n6972_8799.n41 20.9683
R16198 a_n6972_8799.n22 a_n6972_8799.n40 70.5844
R16199 a_n6972_8799.n57 a_n6972_8799.n56 75.3623
R16200 a_n6972_8799.n55 a_n6972_8799.n16 70.3058
R16201 a_n6972_8799.n16 a_n6972_8799.n54 70.1674
R16202 a_n6972_8799.n54 a_n6972_8799.n160 20.9683
R16203 a_n6972_8799.n53 a_n6972_8799.n17 75.0448
R16204 a_n6972_8799.n166 a_n6972_8799.n53 11.2134
R16205 a_n6972_8799.n52 a_n6972_8799.n17 80.4688
R16206 a_n6972_8799.n19 a_n6972_8799.n51 74.73
R16207 a_n6972_8799.n50 a_n6972_8799.n19 70.1674
R16208 a_n6972_8799.n169 a_n6972_8799.n50 20.9683
R16209 a_n6972_8799.n18 a_n6972_8799.n49 70.5844
R16210 a_n6972_8799.n12 a_n6972_8799.n66 70.5844
R16211 a_n6972_8799.n65 a_n6972_8799.n13 70.1674
R16212 a_n6972_8799.n65 a_n6972_8799.n101 20.9683
R16213 a_n6972_8799.n13 a_n6972_8799.n64 74.73
R16214 a_n6972_8799.n110 a_n6972_8799.n64 11.843
R16215 a_n6972_8799.n63 a_n6972_8799.n14 80.4688
R16216 a_n6972_8799.n63 a_n6972_8799.n102 0.365327
R16217 a_n6972_8799.n14 a_n6972_8799.n62 75.0448
R16218 a_n6972_8799.n61 a_n6972_8799.n15 70.1674
R16219 a_n6972_8799.n61 a_n6972_8799.n103 20.9683
R16220 a_n6972_8799.n15 a_n6972_8799.n60 70.3058
R16221 a_n6972_8799.n107 a_n6972_8799.n60 20.6913
R16222 a_n6972_8799.n59 a_n6972_8799.n58 75.3623
R16223 a_n6972_8799.n8 a_n6972_8799.n75 70.5844
R16224 a_n6972_8799.n74 a_n6972_8799.n9 70.1674
R16225 a_n6972_8799.n74 a_n6972_8799.n112 20.9683
R16226 a_n6972_8799.n9 a_n6972_8799.n73 74.73
R16227 a_n6972_8799.n121 a_n6972_8799.n73 11.843
R16228 a_n6972_8799.n72 a_n6972_8799.n10 80.4688
R16229 a_n6972_8799.n72 a_n6972_8799.n113 0.365327
R16230 a_n6972_8799.n10 a_n6972_8799.n71 75.0448
R16231 a_n6972_8799.n70 a_n6972_8799.n11 70.1674
R16232 a_n6972_8799.n70 a_n6972_8799.n114 20.9683
R16233 a_n6972_8799.n11 a_n6972_8799.n69 70.3058
R16234 a_n6972_8799.n118 a_n6972_8799.n69 20.6913
R16235 a_n6972_8799.n68 a_n6972_8799.n67 75.3623
R16236 a_n6972_8799.n4 a_n6972_8799.n84 70.5844
R16237 a_n6972_8799.n83 a_n6972_8799.n5 70.1674
R16238 a_n6972_8799.n83 a_n6972_8799.n124 20.9683
R16239 a_n6972_8799.n5 a_n6972_8799.n82 74.73
R16240 a_n6972_8799.n133 a_n6972_8799.n82 11.843
R16241 a_n6972_8799.n81 a_n6972_8799.n6 80.4688
R16242 a_n6972_8799.n81 a_n6972_8799.n125 0.365327
R16243 a_n6972_8799.n6 a_n6972_8799.n80 75.0448
R16244 a_n6972_8799.n79 a_n6972_8799.n7 70.1674
R16245 a_n6972_8799.n79 a_n6972_8799.n126 20.9683
R16246 a_n6972_8799.n7 a_n6972_8799.n78 70.3058
R16247 a_n6972_8799.n130 a_n6972_8799.n78 20.6913
R16248 a_n6972_8799.n77 a_n6972_8799.n76 75.3623
R16249 a_n6972_8799.n28 a_n6972_8799.n85 98.9633
R16250 a_n6972_8799.n30 a_n6972_8799.n174 98.9631
R16251 a_n6972_8799.n30 a_n6972_8799.n175 98.6055
R16252 a_n6972_8799.n30 a_n6972_8799.n176 98.6055
R16253 a_n6972_8799.n29 a_n6972_8799.n88 98.6055
R16254 a_n6972_8799.n29 a_n6972_8799.n87 98.6055
R16255 a_n6972_8799.n28 a_n6972_8799.n86 98.6055
R16256 a_n6972_8799.n178 a_n6972_8799.n177 98.6054
R16257 a_n6972_8799.n1 a_n6972_8799.n89 81.4626
R16258 a_n6972_8799.n3 a_n6972_8799.n95 81.4626
R16259 a_n6972_8799.n0 a_n6972_8799.n92 81.4626
R16260 a_n6972_8799.n2 a_n6972_8799.n98 80.9324
R16261 a_n6972_8799.n2 a_n6972_8799.n99 80.9324
R16262 a_n6972_8799.n1 a_n6972_8799.n100 80.9324
R16263 a_n6972_8799.n1 a_n6972_8799.n91 80.9324
R16264 a_n6972_8799.n1 a_n6972_8799.n90 80.9324
R16265 a_n6972_8799.n3 a_n6972_8799.n96 80.9324
R16266 a_n6972_8799.n0 a_n6972_8799.n97 80.9324
R16267 a_n6972_8799.n0 a_n6972_8799.n94 80.9324
R16268 a_n6972_8799.n0 a_n6972_8799.n93 80.9324
R16269 a_n6972_8799.n32 a_n6972_8799.n145 20.9683
R16270 a_n6972_8799.n144 a_n6972_8799.n143 48.2005
R16271 a_n6972_8799.n142 a_n6972_8799.n36 20.9683
R16272 a_n6972_8799.n139 a_n6972_8799.n138 48.2005
R16273 a_n6972_8799.n41 a_n6972_8799.n156 20.9683
R16274 a_n6972_8799.n155 a_n6972_8799.n154 48.2005
R16275 a_n6972_8799.n153 a_n6972_8799.n45 20.9683
R16276 a_n6972_8799.n150 a_n6972_8799.n149 48.2005
R16277 a_n6972_8799.n50 a_n6972_8799.n168 20.9683
R16278 a_n6972_8799.n167 a_n6972_8799.n166 48.2005
R16279 a_n6972_8799.n165 a_n6972_8799.n54 20.9683
R16280 a_n6972_8799.n162 a_n6972_8799.n161 48.2005
R16281 a_n6972_8799.n105 a_n6972_8799.n104 48.2005
R16282 a_n6972_8799.n108 a_n6972_8799.n61 20.9683
R16283 a_n6972_8799.n109 a_n6972_8799.n102 48.2005
R16284 a_n6972_8799.n111 a_n6972_8799.n65 20.9683
R16285 a_n6972_8799.n116 a_n6972_8799.n115 48.2005
R16286 a_n6972_8799.n119 a_n6972_8799.n70 20.9683
R16287 a_n6972_8799.n120 a_n6972_8799.n113 48.2005
R16288 a_n6972_8799.n122 a_n6972_8799.n74 20.9683
R16289 a_n6972_8799.n128 a_n6972_8799.n127 48.2005
R16290 a_n6972_8799.n131 a_n6972_8799.n79 20.9683
R16291 a_n6972_8799.n132 a_n6972_8799.n125 48.2005
R16292 a_n6972_8799.n134 a_n6972_8799.n83 20.9683
R16293 a_n6972_8799.n34 a_n6972_8799.n136 47.835
R16294 a_n6972_8799.n37 a_n6972_8799.n141 20.6913
R16295 a_n6972_8799.n43 a_n6972_8799.n147 47.835
R16296 a_n6972_8799.n46 a_n6972_8799.n152 20.6913
R16297 a_n6972_8799.n52 a_n6972_8799.n159 47.835
R16298 a_n6972_8799.n55 a_n6972_8799.n164 20.6913
R16299 a_n6972_8799.n103 a_n6972_8799.n60 21.4216
R16300 a_n6972_8799.n114 a_n6972_8799.n69 21.4216
R16301 a_n6972_8799.n126 a_n6972_8799.n78 21.4216
R16302 a_n6972_8799.t48 a_n6972_8799.n66 484.3
R16303 a_n6972_8799.t57 a_n6972_8799.n75 484.3
R16304 a_n6972_8799.t95 a_n6972_8799.n84 484.3
R16305 a_n6972_8799.n59 a_n6972_8799.n106 45.0871
R16306 a_n6972_8799.n68 a_n6972_8799.n117 45.0871
R16307 a_n6972_8799.n77 a_n6972_8799.n129 45.0871
R16308 a_n6972_8799.n39 a_n6972_8799.n140 45.0871
R16309 a_n6972_8799.n48 a_n6972_8799.n151 45.0871
R16310 a_n6972_8799.n57 a_n6972_8799.n163 45.0871
R16311 a_n6972_8799.n2 a_n6972_8799.n0 34.3237
R16312 a_n6972_8799.n177 a_n6972_8799.n173 32.2674
R16313 a_n6972_8799.n33 a_n6972_8799.n136 11.843
R16314 a_n6972_8799.n141 a_n6972_8799.n38 36.139
R16315 a_n6972_8799.n42 a_n6972_8799.n147 11.843
R16316 a_n6972_8799.n152 a_n6972_8799.n47 36.139
R16317 a_n6972_8799.n51 a_n6972_8799.n159 11.843
R16318 a_n6972_8799.n164 a_n6972_8799.n56 36.139
R16319 a_n6972_8799.n107 a_n6972_8799.n58 36.139
R16320 a_n6972_8799.n101 a_n6972_8799.n64 34.4824
R16321 a_n6972_8799.n118 a_n6972_8799.n67 36.139
R16322 a_n6972_8799.n112 a_n6972_8799.n73 34.4824
R16323 a_n6972_8799.n130 a_n6972_8799.n76 36.139
R16324 a_n6972_8799.n124 a_n6972_8799.n82 34.4824
R16325 a_n6972_8799.n35 a_n6972_8799.n137 35.3134
R16326 a_n6972_8799.n44 a_n6972_8799.n148 35.3134
R16327 a_n6972_8799.n53 a_n6972_8799.n160 35.3134
R16328 a_n6972_8799.n62 a_n6972_8799.n108 35.3134
R16329 a_n6972_8799.n109 a_n6972_8799.n62 11.2134
R16330 a_n6972_8799.n71 a_n6972_8799.n119 35.3134
R16331 a_n6972_8799.n120 a_n6972_8799.n71 11.2134
R16332 a_n6972_8799.n80 a_n6972_8799.n131 35.3134
R16333 a_n6972_8799.n132 a_n6972_8799.n80 11.2134
R16334 a_n6972_8799.n145 a_n6972_8799.n33 34.4824
R16335 a_n6972_8799.n38 a_n6972_8799.n138 10.5784
R16336 a_n6972_8799.n156 a_n6972_8799.n42 34.4824
R16337 a_n6972_8799.n47 a_n6972_8799.n149 10.5784
R16338 a_n6972_8799.n168 a_n6972_8799.n51 34.4824
R16339 a_n6972_8799.n56 a_n6972_8799.n161 10.5784
R16340 a_n6972_8799.n58 a_n6972_8799.n104 10.5784
R16341 a_n6972_8799.n67 a_n6972_8799.n115 10.5784
R16342 a_n6972_8799.n76 a_n6972_8799.n127 10.5784
R16343 a_n6972_8799.n173 a_n6972_8799.n29 18.3287
R16344 a_n6972_8799.n140 a_n6972_8799.n139 14.1472
R16345 a_n6972_8799.n151 a_n6972_8799.n150 14.1472
R16346 a_n6972_8799.n163 a_n6972_8799.n162 14.1472
R16347 a_n6972_8799.n106 a_n6972_8799.n105 14.1472
R16348 a_n6972_8799.n117 a_n6972_8799.n116 14.1472
R16349 a_n6972_8799.n129 a_n6972_8799.n128 14.1472
R16350 a_n6972_8799.n172 a_n6972_8799.n1 12.3339
R16351 a_n6972_8799.n173 a_n6972_8799.n172 11.4887
R16352 a_n6972_8799.n158 a_n6972_8799.n26 9.01755
R16353 a_n6972_8799.n123 a_n6972_8799.n12 9.01755
R16354 a_n6972_8799.n171 a_n6972_8799.n135 7.04375
R16355 a_n6972_8799.n171 a_n6972_8799.n170 6.54711
R16356 a_n6972_8799.n158 a_n6972_8799.n22 4.90959
R16357 a_n6972_8799.n170 a_n6972_8799.n18 4.90959
R16358 a_n6972_8799.n123 a_n6972_8799.n8 4.90959
R16359 a_n6972_8799.n135 a_n6972_8799.n4 4.90959
R16360 a_n6972_8799.n170 a_n6972_8799.n158 4.10845
R16361 a_n6972_8799.n135 a_n6972_8799.n123 4.10845
R16362 a_n6972_8799.n174 a_n6972_8799.t39 3.61217
R16363 a_n6972_8799.n174 a_n6972_8799.t31 3.61217
R16364 a_n6972_8799.n175 a_n6972_8799.t16 3.61217
R16365 a_n6972_8799.n175 a_n6972_8799.t26 3.61217
R16366 a_n6972_8799.n176 a_n6972_8799.t38 3.61217
R16367 a_n6972_8799.n176 a_n6972_8799.t19 3.61217
R16368 a_n6972_8799.n88 a_n6972_8799.t7 3.61217
R16369 a_n6972_8799.n88 a_n6972_8799.t30 3.61217
R16370 a_n6972_8799.n87 a_n6972_8799.t33 3.61217
R16371 a_n6972_8799.n87 a_n6972_8799.t22 3.61217
R16372 a_n6972_8799.n86 a_n6972_8799.t25 3.61217
R16373 a_n6972_8799.n86 a_n6972_8799.t6 3.61217
R16374 a_n6972_8799.n85 a_n6972_8799.t17 3.61217
R16375 a_n6972_8799.n85 a_n6972_8799.t27 3.61217
R16376 a_n6972_8799.n178 a_n6972_8799.t21 3.61217
R16377 a_n6972_8799.t5 a_n6972_8799.n178 3.61217
R16378 a_n6972_8799.n172 a_n6972_8799.n171 3.4105
R16379 a_n6972_8799.n98 a_n6972_8799.t1 2.82907
R16380 a_n6972_8799.n98 a_n6972_8799.t32 2.82907
R16381 a_n6972_8799.n99 a_n6972_8799.t4 2.82907
R16382 a_n6972_8799.n99 a_n6972_8799.t28 2.82907
R16383 a_n6972_8799.n100 a_n6972_8799.t11 2.82907
R16384 a_n6972_8799.n100 a_n6972_8799.t15 2.82907
R16385 a_n6972_8799.n91 a_n6972_8799.t29 2.82907
R16386 a_n6972_8799.n91 a_n6972_8799.t24 2.82907
R16387 a_n6972_8799.n90 a_n6972_8799.t37 2.82907
R16388 a_n6972_8799.n90 a_n6972_8799.t8 2.82907
R16389 a_n6972_8799.n89 a_n6972_8799.t20 2.82907
R16390 a_n6972_8799.n89 a_n6972_8799.t35 2.82907
R16391 a_n6972_8799.n95 a_n6972_8799.t23 2.82907
R16392 a_n6972_8799.n95 a_n6972_8799.t13 2.82907
R16393 a_n6972_8799.n96 a_n6972_8799.t10 2.82907
R16394 a_n6972_8799.n96 a_n6972_8799.t18 2.82907
R16395 a_n6972_8799.n97 a_n6972_8799.t3 2.82907
R16396 a_n6972_8799.n97 a_n6972_8799.t2 2.82907
R16397 a_n6972_8799.n94 a_n6972_8799.t14 2.82907
R16398 a_n6972_8799.n94 a_n6972_8799.t12 2.82907
R16399 a_n6972_8799.n93 a_n6972_8799.t34 2.82907
R16400 a_n6972_8799.n93 a_n6972_8799.t36 2.82907
R16401 a_n6972_8799.n92 a_n6972_8799.t9 2.82907
R16402 a_n6972_8799.n92 a_n6972_8799.t0 2.82907
R16403 a_n6972_8799.n31 a_n6972_8799.n146 22.3251
R16404 a_n6972_8799.n40 a_n6972_8799.n157 22.3251
R16405 a_n6972_8799.n49 a_n6972_8799.n169 22.3251
R16406 a_n6972_8799.n66 a_n6972_8799.n111 22.3251
R16407 a_n6972_8799.n75 a_n6972_8799.n122 22.3251
R16408 a_n6972_8799.n84 a_n6972_8799.n134 22.3251
R16409 a_n6972_8799.n34 a_n6972_8799.n144 0.365327
R16410 a_n6972_8799.n142 a_n6972_8799.n37 21.4216
R16411 a_n6972_8799.n43 a_n6972_8799.n155 0.365327
R16412 a_n6972_8799.n153 a_n6972_8799.n46 21.4216
R16413 a_n6972_8799.n52 a_n6972_8799.n167 0.365327
R16414 a_n6972_8799.n165 a_n6972_8799.n55 21.4216
R16415 a_n6972_8799.n110 a_n6972_8799.n63 47.835
R16416 a_n6972_8799.n121 a_n6972_8799.n72 47.835
R16417 a_n6972_8799.n133 a_n6972_8799.n81 47.835
R16418 a_n6972_8799.n1 a_n6972_8799.n2 2.12119
R16419 a_n6972_8799.n0 a_n6972_8799.n3 1.59102
R16420 a_n6972_8799.n27 a_n6972_8799.n25 0.758076
R16421 a_n6972_8799.n25 a_n6972_8799.n24 0.758076
R16422 a_n6972_8799.n39 a_n6972_8799.n24 0.758076
R16423 a_n6972_8799.n23 a_n6972_8799.n21 0.758076
R16424 a_n6972_8799.n21 a_n6972_8799.n20 0.758076
R16425 a_n6972_8799.n48 a_n6972_8799.n20 0.758076
R16426 a_n6972_8799.n19 a_n6972_8799.n17 0.758076
R16427 a_n6972_8799.n17 a_n6972_8799.n16 0.758076
R16428 a_n6972_8799.n57 a_n6972_8799.n16 0.758076
R16429 a_n6972_8799.n15 a_n6972_8799.n14 0.758076
R16430 a_n6972_8799.n14 a_n6972_8799.n13 0.758076
R16431 a_n6972_8799.n13 a_n6972_8799.n12 0.758076
R16432 a_n6972_8799.n11 a_n6972_8799.n10 0.758076
R16433 a_n6972_8799.n10 a_n6972_8799.n9 0.758076
R16434 a_n6972_8799.n9 a_n6972_8799.n8 0.758076
R16435 a_n6972_8799.n7 a_n6972_8799.n6 0.758076
R16436 a_n6972_8799.n6 a_n6972_8799.n5 0.758076
R16437 a_n6972_8799.n5 a_n6972_8799.n4 0.758076
R16438 a_n6972_8799.n177 a_n6972_8799.n30 0.716017
R16439 a_n6972_8799.n29 a_n6972_8799.n28 0.716017
R16440 a_n6972_8799.n77 a_n6972_8799.n7 0.568682
R16441 a_n6972_8799.n68 a_n6972_8799.n11 0.568682
R16442 a_n6972_8799.n59 a_n6972_8799.n15 0.568682
R16443 a_n6972_8799.n19 a_n6972_8799.n18 0.568682
R16444 a_n6972_8799.n23 a_n6972_8799.n22 0.568682
R16445 a_n6972_8799.n27 a_n6972_8799.n26 0.568682
R16446 vdd.n303 vdd.n267 756.745
R16447 vdd.n252 vdd.n216 756.745
R16448 vdd.n209 vdd.n173 756.745
R16449 vdd.n158 vdd.n122 756.745
R16450 vdd.n116 vdd.n80 756.745
R16451 vdd.n65 vdd.n29 756.745
R16452 vdd.n1860 vdd.n1824 756.745
R16453 vdd.n1911 vdd.n1875 756.745
R16454 vdd.n1766 vdd.n1730 756.745
R16455 vdd.n1817 vdd.n1781 756.745
R16456 vdd.n1673 vdd.n1637 756.745
R16457 vdd.n1724 vdd.n1688 756.745
R16458 vdd.n1081 vdd.t8 640.208
R16459 vdd.n809 vdd.t50 640.208
R16460 vdd.n1101 vdd.t34 640.208
R16461 vdd.n800 vdd.t68 640.208
R16462 vdd.n700 vdd.t37 640.208
R16463 vdd.n2416 vdd.t65 640.208
R16464 vdd.n661 vdd.t74 640.208
R16465 vdd.n2413 vdd.t54 640.208
R16466 vdd.n625 vdd.t4 640.208
R16467 vdd.n871 vdd.t58 640.208
R16468 vdd.n1472 vdd.t24 592.009
R16469 vdd.n1509 vdd.t31 592.009
R16470 vdd.n1383 vdd.t44 592.009
R16471 vdd.n1981 vdd.t16 592.009
R16472 vdd.n1018 vdd.t47 592.009
R16473 vdd.n978 vdd.t62 592.009
R16474 vdd.n3113 vdd.t20 592.009
R16475 vdd.n427 vdd.t71 592.009
R16476 vdd.n387 vdd.t77 592.009
R16477 vdd.n580 vdd.t28 592.009
R16478 vdd.n543 vdd.t41 592.009
R16479 vdd.n2900 vdd.t12 592.009
R16480 vdd.n304 vdd.n303 585
R16481 vdd.n302 vdd.n269 585
R16482 vdd.n301 vdd.n300 585
R16483 vdd.n272 vdd.n270 585
R16484 vdd.n295 vdd.n294 585
R16485 vdd.n293 vdd.n292 585
R16486 vdd.n276 vdd.n275 585
R16487 vdd.n287 vdd.n286 585
R16488 vdd.n285 vdd.n284 585
R16489 vdd.n280 vdd.n279 585
R16490 vdd.n253 vdd.n252 585
R16491 vdd.n251 vdd.n218 585
R16492 vdd.n250 vdd.n249 585
R16493 vdd.n221 vdd.n219 585
R16494 vdd.n244 vdd.n243 585
R16495 vdd.n242 vdd.n241 585
R16496 vdd.n225 vdd.n224 585
R16497 vdd.n236 vdd.n235 585
R16498 vdd.n234 vdd.n233 585
R16499 vdd.n229 vdd.n228 585
R16500 vdd.n210 vdd.n209 585
R16501 vdd.n208 vdd.n175 585
R16502 vdd.n207 vdd.n206 585
R16503 vdd.n178 vdd.n176 585
R16504 vdd.n201 vdd.n200 585
R16505 vdd.n199 vdd.n198 585
R16506 vdd.n182 vdd.n181 585
R16507 vdd.n193 vdd.n192 585
R16508 vdd.n191 vdd.n190 585
R16509 vdd.n186 vdd.n185 585
R16510 vdd.n159 vdd.n158 585
R16511 vdd.n157 vdd.n124 585
R16512 vdd.n156 vdd.n155 585
R16513 vdd.n127 vdd.n125 585
R16514 vdd.n150 vdd.n149 585
R16515 vdd.n148 vdd.n147 585
R16516 vdd.n131 vdd.n130 585
R16517 vdd.n142 vdd.n141 585
R16518 vdd.n140 vdd.n139 585
R16519 vdd.n135 vdd.n134 585
R16520 vdd.n117 vdd.n116 585
R16521 vdd.n115 vdd.n82 585
R16522 vdd.n114 vdd.n113 585
R16523 vdd.n85 vdd.n83 585
R16524 vdd.n108 vdd.n107 585
R16525 vdd.n106 vdd.n105 585
R16526 vdd.n89 vdd.n88 585
R16527 vdd.n100 vdd.n99 585
R16528 vdd.n98 vdd.n97 585
R16529 vdd.n93 vdd.n92 585
R16530 vdd.n66 vdd.n65 585
R16531 vdd.n64 vdd.n31 585
R16532 vdd.n63 vdd.n62 585
R16533 vdd.n34 vdd.n32 585
R16534 vdd.n57 vdd.n56 585
R16535 vdd.n55 vdd.n54 585
R16536 vdd.n38 vdd.n37 585
R16537 vdd.n49 vdd.n48 585
R16538 vdd.n47 vdd.n46 585
R16539 vdd.n42 vdd.n41 585
R16540 vdd.n1861 vdd.n1860 585
R16541 vdd.n1859 vdd.n1826 585
R16542 vdd.n1858 vdd.n1857 585
R16543 vdd.n1829 vdd.n1827 585
R16544 vdd.n1852 vdd.n1851 585
R16545 vdd.n1850 vdd.n1849 585
R16546 vdd.n1833 vdd.n1832 585
R16547 vdd.n1844 vdd.n1843 585
R16548 vdd.n1842 vdd.n1841 585
R16549 vdd.n1837 vdd.n1836 585
R16550 vdd.n1912 vdd.n1911 585
R16551 vdd.n1910 vdd.n1877 585
R16552 vdd.n1909 vdd.n1908 585
R16553 vdd.n1880 vdd.n1878 585
R16554 vdd.n1903 vdd.n1902 585
R16555 vdd.n1901 vdd.n1900 585
R16556 vdd.n1884 vdd.n1883 585
R16557 vdd.n1895 vdd.n1894 585
R16558 vdd.n1893 vdd.n1892 585
R16559 vdd.n1888 vdd.n1887 585
R16560 vdd.n1767 vdd.n1766 585
R16561 vdd.n1765 vdd.n1732 585
R16562 vdd.n1764 vdd.n1763 585
R16563 vdd.n1735 vdd.n1733 585
R16564 vdd.n1758 vdd.n1757 585
R16565 vdd.n1756 vdd.n1755 585
R16566 vdd.n1739 vdd.n1738 585
R16567 vdd.n1750 vdd.n1749 585
R16568 vdd.n1748 vdd.n1747 585
R16569 vdd.n1743 vdd.n1742 585
R16570 vdd.n1818 vdd.n1817 585
R16571 vdd.n1816 vdd.n1783 585
R16572 vdd.n1815 vdd.n1814 585
R16573 vdd.n1786 vdd.n1784 585
R16574 vdd.n1809 vdd.n1808 585
R16575 vdd.n1807 vdd.n1806 585
R16576 vdd.n1790 vdd.n1789 585
R16577 vdd.n1801 vdd.n1800 585
R16578 vdd.n1799 vdd.n1798 585
R16579 vdd.n1794 vdd.n1793 585
R16580 vdd.n1674 vdd.n1673 585
R16581 vdd.n1672 vdd.n1639 585
R16582 vdd.n1671 vdd.n1670 585
R16583 vdd.n1642 vdd.n1640 585
R16584 vdd.n1665 vdd.n1664 585
R16585 vdd.n1663 vdd.n1662 585
R16586 vdd.n1646 vdd.n1645 585
R16587 vdd.n1657 vdd.n1656 585
R16588 vdd.n1655 vdd.n1654 585
R16589 vdd.n1650 vdd.n1649 585
R16590 vdd.n1725 vdd.n1724 585
R16591 vdd.n1723 vdd.n1690 585
R16592 vdd.n1722 vdd.n1721 585
R16593 vdd.n1693 vdd.n1691 585
R16594 vdd.n1716 vdd.n1715 585
R16595 vdd.n1714 vdd.n1713 585
R16596 vdd.n1697 vdd.n1696 585
R16597 vdd.n1708 vdd.n1707 585
R16598 vdd.n1706 vdd.n1705 585
R16599 vdd.n1701 vdd.n1700 585
R16600 vdd.n3229 vdd.n352 488.781
R16601 vdd.n3111 vdd.n350 488.781
R16602 vdd.n3033 vdd.n515 488.781
R16603 vdd.n3031 vdd.n517 488.781
R16604 vdd.n1976 vdd.n1265 488.781
R16605 vdd.n1979 vdd.n1978 488.781
R16606 vdd.n1578 vdd.n1343 488.781
R16607 vdd.n1576 vdd.n1346 488.781
R16608 vdd.n281 vdd.t215 329.043
R16609 vdd.n230 vdd.t197 329.043
R16610 vdd.n187 vdd.t206 329.043
R16611 vdd.n136 vdd.t186 329.043
R16612 vdd.n94 vdd.t152 329.043
R16613 vdd.n43 vdd.t160 329.043
R16614 vdd.n1838 vdd.t221 329.043
R16615 vdd.n1889 vdd.t155 329.043
R16616 vdd.n1744 vdd.t212 329.043
R16617 vdd.n1795 vdd.t141 329.043
R16618 vdd.n1651 vdd.t162 329.043
R16619 vdd.n1702 vdd.t153 329.043
R16620 vdd.n1472 vdd.t27 319.788
R16621 vdd.n1509 vdd.t33 319.788
R16622 vdd.n1383 vdd.t46 319.788
R16623 vdd.n1981 vdd.t18 319.788
R16624 vdd.n1018 vdd.t48 319.788
R16625 vdd.n978 vdd.t63 319.788
R16626 vdd.n3113 vdd.t22 319.788
R16627 vdd.n427 vdd.t72 319.788
R16628 vdd.n387 vdd.t78 319.788
R16629 vdd.n580 vdd.t30 319.788
R16630 vdd.n543 vdd.t43 319.788
R16631 vdd.n2900 vdd.t15 319.788
R16632 vdd.n1473 vdd.t26 303.69
R16633 vdd.n1510 vdd.t32 303.69
R16634 vdd.n1384 vdd.t45 303.69
R16635 vdd.n1982 vdd.t19 303.69
R16636 vdd.n1019 vdd.t49 303.69
R16637 vdd.n979 vdd.t64 303.69
R16638 vdd.n3114 vdd.t23 303.69
R16639 vdd.n428 vdd.t73 303.69
R16640 vdd.n388 vdd.t79 303.69
R16641 vdd.n581 vdd.t29 303.69
R16642 vdd.n544 vdd.t42 303.69
R16643 vdd.n2901 vdd.t14 303.69
R16644 vdd.n2648 vdd.n755 291.221
R16645 vdd.n2862 vdd.n635 291.221
R16646 vdd.n2799 vdd.n632 291.221
R16647 vdd.n2580 vdd.n2579 291.221
R16648 vdd.n2376 vdd.n797 291.221
R16649 vdd.n2307 vdd.n2306 291.221
R16650 vdd.n1137 vdd.n1136 291.221
R16651 vdd.n2127 vdd.n903 291.221
R16652 vdd.n2778 vdd.n633 291.221
R16653 vdd.n2865 vdd.n2864 291.221
R16654 vdd.n2484 vdd.n2410 291.221
R16655 vdd.n2652 vdd.n759 291.221
R16656 vdd.n2304 vdd.n807 291.221
R16657 vdd.n805 vdd.n779 291.221
R16658 vdd.n1215 vdd.n944 291.221
R16659 vdd.n2131 vdd.n908 291.221
R16660 vdd.n2780 vdd.n633 185
R16661 vdd.n2863 vdd.n633 185
R16662 vdd.n2782 vdd.n2781 185
R16663 vdd.n2781 vdd.n631 185
R16664 vdd.n2783 vdd.n667 185
R16665 vdd.n2793 vdd.n667 185
R16666 vdd.n2784 vdd.n676 185
R16667 vdd.n676 vdd.n674 185
R16668 vdd.n2786 vdd.n2785 185
R16669 vdd.n2787 vdd.n2786 185
R16670 vdd.n2739 vdd.n675 185
R16671 vdd.n675 vdd.n671 185
R16672 vdd.n2738 vdd.n2737 185
R16673 vdd.n2737 vdd.n2736 185
R16674 vdd.n678 vdd.n677 185
R16675 vdd.n679 vdd.n678 185
R16676 vdd.n2729 vdd.n2728 185
R16677 vdd.n2730 vdd.n2729 185
R16678 vdd.n2727 vdd.n688 185
R16679 vdd.n688 vdd.n685 185
R16680 vdd.n2726 vdd.n2725 185
R16681 vdd.n2725 vdd.n2724 185
R16682 vdd.n690 vdd.n689 185
R16683 vdd.n698 vdd.n690 185
R16684 vdd.n2717 vdd.n2716 185
R16685 vdd.n2718 vdd.n2717 185
R16686 vdd.n2714 vdd.n699 185
R16687 vdd.n706 vdd.n699 185
R16688 vdd.n2713 vdd.n2712 185
R16689 vdd.n2712 vdd.n2711 185
R16690 vdd.n702 vdd.n701 185
R16691 vdd.n703 vdd.n702 185
R16692 vdd.n2704 vdd.n2703 185
R16693 vdd.n2705 vdd.n2704 185
R16694 vdd.n2702 vdd.n713 185
R16695 vdd.n713 vdd.n710 185
R16696 vdd.n2701 vdd.n2700 185
R16697 vdd.n2700 vdd.n2699 185
R16698 vdd.n715 vdd.n714 185
R16699 vdd.n723 vdd.n715 185
R16700 vdd.n2692 vdd.n2691 185
R16701 vdd.n2693 vdd.n2692 185
R16702 vdd.n2690 vdd.n724 185
R16703 vdd.n729 vdd.n724 185
R16704 vdd.n2689 vdd.n2688 185
R16705 vdd.n2688 vdd.n2687 185
R16706 vdd.n726 vdd.n725 185
R16707 vdd.n2559 vdd.n726 185
R16708 vdd.n2680 vdd.n2679 185
R16709 vdd.n2681 vdd.n2680 185
R16710 vdd.n2678 vdd.n736 185
R16711 vdd.n736 vdd.n733 185
R16712 vdd.n2677 vdd.n2676 185
R16713 vdd.n2676 vdd.n2675 185
R16714 vdd.n738 vdd.n737 185
R16715 vdd.n739 vdd.n738 185
R16716 vdd.n2668 vdd.n2667 185
R16717 vdd.n2669 vdd.n2668 185
R16718 vdd.n2666 vdd.n748 185
R16719 vdd.n748 vdd.n745 185
R16720 vdd.n2665 vdd.n2664 185
R16721 vdd.n2664 vdd.n2663 185
R16722 vdd.n750 vdd.n749 185
R16723 vdd.n2574 vdd.n750 185
R16724 vdd.n2656 vdd.n2655 185
R16725 vdd.n2657 vdd.n2656 185
R16726 vdd.n2654 vdd.n759 185
R16727 vdd.n759 vdd.n756 185
R16728 vdd.n2653 vdd.n2652 185
R16729 vdd.n761 vdd.n760 185
R16730 vdd.n2420 vdd.n2419 185
R16731 vdd.n2422 vdd.n2421 185
R16732 vdd.n2424 vdd.n2423 185
R16733 vdd.n2426 vdd.n2425 185
R16734 vdd.n2428 vdd.n2427 185
R16735 vdd.n2430 vdd.n2429 185
R16736 vdd.n2432 vdd.n2431 185
R16737 vdd.n2434 vdd.n2433 185
R16738 vdd.n2436 vdd.n2435 185
R16739 vdd.n2438 vdd.n2437 185
R16740 vdd.n2440 vdd.n2439 185
R16741 vdd.n2442 vdd.n2441 185
R16742 vdd.n2444 vdd.n2443 185
R16743 vdd.n2446 vdd.n2445 185
R16744 vdd.n2448 vdd.n2447 185
R16745 vdd.n2450 vdd.n2449 185
R16746 vdd.n2452 vdd.n2451 185
R16747 vdd.n2454 vdd.n2453 185
R16748 vdd.n2456 vdd.n2455 185
R16749 vdd.n2458 vdd.n2457 185
R16750 vdd.n2460 vdd.n2459 185
R16751 vdd.n2462 vdd.n2461 185
R16752 vdd.n2464 vdd.n2463 185
R16753 vdd.n2466 vdd.n2465 185
R16754 vdd.n2468 vdd.n2467 185
R16755 vdd.n2470 vdd.n2469 185
R16756 vdd.n2472 vdd.n2471 185
R16757 vdd.n2474 vdd.n2473 185
R16758 vdd.n2476 vdd.n2475 185
R16759 vdd.n2478 vdd.n2477 185
R16760 vdd.n2480 vdd.n2479 185
R16761 vdd.n2482 vdd.n2481 185
R16762 vdd.n2483 vdd.n2410 185
R16763 vdd.n2650 vdd.n2410 185
R16764 vdd.n2866 vdd.n2865 185
R16765 vdd.n2867 vdd.n624 185
R16766 vdd.n2869 vdd.n2868 185
R16767 vdd.n2871 vdd.n622 185
R16768 vdd.n2873 vdd.n2872 185
R16769 vdd.n2874 vdd.n621 185
R16770 vdd.n2876 vdd.n2875 185
R16771 vdd.n2878 vdd.n619 185
R16772 vdd.n2880 vdd.n2879 185
R16773 vdd.n2881 vdd.n618 185
R16774 vdd.n2883 vdd.n2882 185
R16775 vdd.n2885 vdd.n616 185
R16776 vdd.n2887 vdd.n2886 185
R16777 vdd.n2888 vdd.n615 185
R16778 vdd.n2890 vdd.n2889 185
R16779 vdd.n2892 vdd.n614 185
R16780 vdd.n2893 vdd.n611 185
R16781 vdd.n2896 vdd.n2895 185
R16782 vdd.n612 vdd.n610 185
R16783 vdd.n2752 vdd.n2751 185
R16784 vdd.n2754 vdd.n2753 185
R16785 vdd.n2756 vdd.n2748 185
R16786 vdd.n2758 vdd.n2757 185
R16787 vdd.n2759 vdd.n2747 185
R16788 vdd.n2761 vdd.n2760 185
R16789 vdd.n2763 vdd.n2745 185
R16790 vdd.n2765 vdd.n2764 185
R16791 vdd.n2766 vdd.n2744 185
R16792 vdd.n2768 vdd.n2767 185
R16793 vdd.n2770 vdd.n2742 185
R16794 vdd.n2772 vdd.n2771 185
R16795 vdd.n2773 vdd.n2741 185
R16796 vdd.n2775 vdd.n2774 185
R16797 vdd.n2777 vdd.n2740 185
R16798 vdd.n2779 vdd.n2778 185
R16799 vdd.n2778 vdd.n613 185
R16800 vdd.n2864 vdd.n628 185
R16801 vdd.n2864 vdd.n2863 185
R16802 vdd.n2487 vdd.n630 185
R16803 vdd.n631 vdd.n630 185
R16804 vdd.n2488 vdd.n666 185
R16805 vdd.n2793 vdd.n666 185
R16806 vdd.n2490 vdd.n2489 185
R16807 vdd.n2489 vdd.n674 185
R16808 vdd.n2491 vdd.n673 185
R16809 vdd.n2787 vdd.n673 185
R16810 vdd.n2493 vdd.n2492 185
R16811 vdd.n2492 vdd.n671 185
R16812 vdd.n2494 vdd.n681 185
R16813 vdd.n2736 vdd.n681 185
R16814 vdd.n2496 vdd.n2495 185
R16815 vdd.n2495 vdd.n679 185
R16816 vdd.n2497 vdd.n687 185
R16817 vdd.n2730 vdd.n687 185
R16818 vdd.n2499 vdd.n2498 185
R16819 vdd.n2498 vdd.n685 185
R16820 vdd.n2500 vdd.n692 185
R16821 vdd.n2724 vdd.n692 185
R16822 vdd.n2502 vdd.n2501 185
R16823 vdd.n2501 vdd.n698 185
R16824 vdd.n2503 vdd.n697 185
R16825 vdd.n2718 vdd.n697 185
R16826 vdd.n2505 vdd.n2504 185
R16827 vdd.n2504 vdd.n706 185
R16828 vdd.n2506 vdd.n705 185
R16829 vdd.n2711 vdd.n705 185
R16830 vdd.n2508 vdd.n2507 185
R16831 vdd.n2507 vdd.n703 185
R16832 vdd.n2509 vdd.n712 185
R16833 vdd.n2705 vdd.n712 185
R16834 vdd.n2511 vdd.n2510 185
R16835 vdd.n2510 vdd.n710 185
R16836 vdd.n2512 vdd.n717 185
R16837 vdd.n2699 vdd.n717 185
R16838 vdd.n2514 vdd.n2513 185
R16839 vdd.n2513 vdd.n723 185
R16840 vdd.n2515 vdd.n722 185
R16841 vdd.n2693 vdd.n722 185
R16842 vdd.n2517 vdd.n2516 185
R16843 vdd.n2516 vdd.n729 185
R16844 vdd.n2518 vdd.n728 185
R16845 vdd.n2687 vdd.n728 185
R16846 vdd.n2561 vdd.n2560 185
R16847 vdd.n2560 vdd.n2559 185
R16848 vdd.n2562 vdd.n735 185
R16849 vdd.n2681 vdd.n735 185
R16850 vdd.n2564 vdd.n2563 185
R16851 vdd.n2563 vdd.n733 185
R16852 vdd.n2565 vdd.n741 185
R16853 vdd.n2675 vdd.n741 185
R16854 vdd.n2567 vdd.n2566 185
R16855 vdd.n2566 vdd.n739 185
R16856 vdd.n2568 vdd.n747 185
R16857 vdd.n2669 vdd.n747 185
R16858 vdd.n2570 vdd.n2569 185
R16859 vdd.n2569 vdd.n745 185
R16860 vdd.n2571 vdd.n752 185
R16861 vdd.n2663 vdd.n752 185
R16862 vdd.n2573 vdd.n2572 185
R16863 vdd.n2574 vdd.n2573 185
R16864 vdd.n2486 vdd.n758 185
R16865 vdd.n2657 vdd.n758 185
R16866 vdd.n2485 vdd.n2484 185
R16867 vdd.n2484 vdd.n756 185
R16868 vdd.n1976 vdd.n1975 185
R16869 vdd.n1977 vdd.n1976 185
R16870 vdd.n1266 vdd.n1264 185
R16871 vdd.n1968 vdd.n1264 185
R16872 vdd.n1971 vdd.n1970 185
R16873 vdd.n1970 vdd.n1969 185
R16874 vdd.n1269 vdd.n1268 185
R16875 vdd.n1270 vdd.n1269 185
R16876 vdd.n1957 vdd.n1956 185
R16877 vdd.n1958 vdd.n1957 185
R16878 vdd.n1278 vdd.n1277 185
R16879 vdd.n1949 vdd.n1277 185
R16880 vdd.n1952 vdd.n1951 185
R16881 vdd.n1951 vdd.n1950 185
R16882 vdd.n1281 vdd.n1280 185
R16883 vdd.n1287 vdd.n1281 185
R16884 vdd.n1940 vdd.n1939 185
R16885 vdd.n1941 vdd.n1940 185
R16886 vdd.n1289 vdd.n1288 185
R16887 vdd.n1932 vdd.n1288 185
R16888 vdd.n1935 vdd.n1934 185
R16889 vdd.n1934 vdd.n1933 185
R16890 vdd.n1292 vdd.n1291 185
R16891 vdd.n1293 vdd.n1292 185
R16892 vdd.n1923 vdd.n1922 185
R16893 vdd.n1924 vdd.n1923 185
R16894 vdd.n1301 vdd.n1300 185
R16895 vdd.n1300 vdd.n1299 185
R16896 vdd.n1636 vdd.n1635 185
R16897 vdd.n1635 vdd.n1634 185
R16898 vdd.n1304 vdd.n1303 185
R16899 vdd.n1310 vdd.n1304 185
R16900 vdd.n1625 vdd.n1624 185
R16901 vdd.n1626 vdd.n1625 185
R16902 vdd.n1312 vdd.n1311 185
R16903 vdd.n1617 vdd.n1311 185
R16904 vdd.n1620 vdd.n1619 185
R16905 vdd.n1619 vdd.n1618 185
R16906 vdd.n1315 vdd.n1314 185
R16907 vdd.n1322 vdd.n1315 185
R16908 vdd.n1608 vdd.n1607 185
R16909 vdd.n1609 vdd.n1608 185
R16910 vdd.n1324 vdd.n1323 185
R16911 vdd.n1323 vdd.n1321 185
R16912 vdd.n1603 vdd.n1602 185
R16913 vdd.n1602 vdd.n1601 185
R16914 vdd.n1327 vdd.n1326 185
R16915 vdd.n1328 vdd.n1327 185
R16916 vdd.n1592 vdd.n1591 185
R16917 vdd.n1593 vdd.n1592 185
R16918 vdd.n1336 vdd.n1335 185
R16919 vdd.n1335 vdd.n1334 185
R16920 vdd.n1587 vdd.n1586 185
R16921 vdd.n1586 vdd.n1585 185
R16922 vdd.n1339 vdd.n1338 185
R16923 vdd.n1345 vdd.n1339 185
R16924 vdd.n1576 vdd.n1575 185
R16925 vdd.n1577 vdd.n1576 185
R16926 vdd.n1572 vdd.n1346 185
R16927 vdd.n1571 vdd.n1349 185
R16928 vdd.n1570 vdd.n1350 185
R16929 vdd.n1350 vdd.n1344 185
R16930 vdd.n1353 vdd.n1351 185
R16931 vdd.n1566 vdd.n1355 185
R16932 vdd.n1565 vdd.n1356 185
R16933 vdd.n1564 vdd.n1358 185
R16934 vdd.n1361 vdd.n1359 185
R16935 vdd.n1560 vdd.n1363 185
R16936 vdd.n1559 vdd.n1364 185
R16937 vdd.n1558 vdd.n1366 185
R16938 vdd.n1369 vdd.n1367 185
R16939 vdd.n1554 vdd.n1371 185
R16940 vdd.n1553 vdd.n1372 185
R16941 vdd.n1552 vdd.n1374 185
R16942 vdd.n1377 vdd.n1375 185
R16943 vdd.n1548 vdd.n1379 185
R16944 vdd.n1547 vdd.n1380 185
R16945 vdd.n1546 vdd.n1382 185
R16946 vdd.n1387 vdd.n1385 185
R16947 vdd.n1542 vdd.n1389 185
R16948 vdd.n1541 vdd.n1390 185
R16949 vdd.n1540 vdd.n1392 185
R16950 vdd.n1395 vdd.n1393 185
R16951 vdd.n1536 vdd.n1397 185
R16952 vdd.n1535 vdd.n1398 185
R16953 vdd.n1534 vdd.n1400 185
R16954 vdd.n1403 vdd.n1401 185
R16955 vdd.n1530 vdd.n1405 185
R16956 vdd.n1529 vdd.n1406 185
R16957 vdd.n1528 vdd.n1408 185
R16958 vdd.n1411 vdd.n1409 185
R16959 vdd.n1524 vdd.n1413 185
R16960 vdd.n1523 vdd.n1414 185
R16961 vdd.n1522 vdd.n1416 185
R16962 vdd.n1419 vdd.n1417 185
R16963 vdd.n1518 vdd.n1421 185
R16964 vdd.n1517 vdd.n1422 185
R16965 vdd.n1516 vdd.n1424 185
R16966 vdd.n1427 vdd.n1425 185
R16967 vdd.n1512 vdd.n1429 185
R16968 vdd.n1511 vdd.n1508 185
R16969 vdd.n1506 vdd.n1430 185
R16970 vdd.n1505 vdd.n1504 185
R16971 vdd.n1435 vdd.n1432 185
R16972 vdd.n1500 vdd.n1436 185
R16973 vdd.n1499 vdd.n1438 185
R16974 vdd.n1498 vdd.n1439 185
R16975 vdd.n1443 vdd.n1440 185
R16976 vdd.n1494 vdd.n1444 185
R16977 vdd.n1493 vdd.n1446 185
R16978 vdd.n1492 vdd.n1447 185
R16979 vdd.n1451 vdd.n1448 185
R16980 vdd.n1488 vdd.n1452 185
R16981 vdd.n1487 vdd.n1454 185
R16982 vdd.n1486 vdd.n1455 185
R16983 vdd.n1459 vdd.n1456 185
R16984 vdd.n1482 vdd.n1460 185
R16985 vdd.n1481 vdd.n1462 185
R16986 vdd.n1480 vdd.n1463 185
R16987 vdd.n1467 vdd.n1464 185
R16988 vdd.n1476 vdd.n1468 185
R16989 vdd.n1475 vdd.n1470 185
R16990 vdd.n1471 vdd.n1343 185
R16991 vdd.n1344 vdd.n1343 185
R16992 vdd.n1980 vdd.n1979 185
R16993 vdd.n1984 vdd.n1260 185
R16994 vdd.n1259 vdd.n1253 185
R16995 vdd.n1257 vdd.n1256 185
R16996 vdd.n1255 vdd.n1049 185
R16997 vdd.n1988 vdd.n1046 185
R16998 vdd.n1990 vdd.n1989 185
R16999 vdd.n1992 vdd.n1044 185
R17000 vdd.n1994 vdd.n1993 185
R17001 vdd.n1995 vdd.n1039 185
R17002 vdd.n1997 vdd.n1996 185
R17003 vdd.n1999 vdd.n1037 185
R17004 vdd.n2001 vdd.n2000 185
R17005 vdd.n2002 vdd.n1032 185
R17006 vdd.n2004 vdd.n2003 185
R17007 vdd.n2006 vdd.n1030 185
R17008 vdd.n2008 vdd.n2007 185
R17009 vdd.n2009 vdd.n1026 185
R17010 vdd.n2011 vdd.n2010 185
R17011 vdd.n2013 vdd.n1023 185
R17012 vdd.n2015 vdd.n2014 185
R17013 vdd.n1024 vdd.n1017 185
R17014 vdd.n2019 vdd.n1021 185
R17015 vdd.n2020 vdd.n1013 185
R17016 vdd.n2022 vdd.n2021 185
R17017 vdd.n2024 vdd.n1011 185
R17018 vdd.n2026 vdd.n2025 185
R17019 vdd.n2027 vdd.n1006 185
R17020 vdd.n2029 vdd.n2028 185
R17021 vdd.n2031 vdd.n1004 185
R17022 vdd.n2033 vdd.n2032 185
R17023 vdd.n2034 vdd.n999 185
R17024 vdd.n2036 vdd.n2035 185
R17025 vdd.n2038 vdd.n997 185
R17026 vdd.n2040 vdd.n2039 185
R17027 vdd.n2041 vdd.n992 185
R17028 vdd.n2043 vdd.n2042 185
R17029 vdd.n2045 vdd.n990 185
R17030 vdd.n2047 vdd.n2046 185
R17031 vdd.n2048 vdd.n986 185
R17032 vdd.n2050 vdd.n2049 185
R17033 vdd.n2052 vdd.n983 185
R17034 vdd.n2054 vdd.n2053 185
R17035 vdd.n984 vdd.n977 185
R17036 vdd.n2058 vdd.n981 185
R17037 vdd.n2059 vdd.n973 185
R17038 vdd.n2061 vdd.n2060 185
R17039 vdd.n2063 vdd.n971 185
R17040 vdd.n2065 vdd.n2064 185
R17041 vdd.n2066 vdd.n966 185
R17042 vdd.n2068 vdd.n2067 185
R17043 vdd.n2070 vdd.n964 185
R17044 vdd.n2072 vdd.n2071 185
R17045 vdd.n2073 vdd.n959 185
R17046 vdd.n2075 vdd.n2074 185
R17047 vdd.n2077 vdd.n957 185
R17048 vdd.n2079 vdd.n2078 185
R17049 vdd.n2080 vdd.n955 185
R17050 vdd.n2082 vdd.n2081 185
R17051 vdd.n2085 vdd.n2084 185
R17052 vdd.n2087 vdd.n2086 185
R17053 vdd.n2089 vdd.n953 185
R17054 vdd.n2091 vdd.n2090 185
R17055 vdd.n1265 vdd.n952 185
R17056 vdd.n1978 vdd.n1263 185
R17057 vdd.n1978 vdd.n1977 185
R17058 vdd.n1273 vdd.n1262 185
R17059 vdd.n1968 vdd.n1262 185
R17060 vdd.n1967 vdd.n1966 185
R17061 vdd.n1969 vdd.n1967 185
R17062 vdd.n1272 vdd.n1271 185
R17063 vdd.n1271 vdd.n1270 185
R17064 vdd.n1960 vdd.n1959 185
R17065 vdd.n1959 vdd.n1958 185
R17066 vdd.n1276 vdd.n1275 185
R17067 vdd.n1949 vdd.n1276 185
R17068 vdd.n1948 vdd.n1947 185
R17069 vdd.n1950 vdd.n1948 185
R17070 vdd.n1283 vdd.n1282 185
R17071 vdd.n1287 vdd.n1282 185
R17072 vdd.n1943 vdd.n1942 185
R17073 vdd.n1942 vdd.n1941 185
R17074 vdd.n1286 vdd.n1285 185
R17075 vdd.n1932 vdd.n1286 185
R17076 vdd.n1931 vdd.n1930 185
R17077 vdd.n1933 vdd.n1931 185
R17078 vdd.n1295 vdd.n1294 185
R17079 vdd.n1294 vdd.n1293 185
R17080 vdd.n1926 vdd.n1925 185
R17081 vdd.n1925 vdd.n1924 185
R17082 vdd.n1298 vdd.n1297 185
R17083 vdd.n1299 vdd.n1298 185
R17084 vdd.n1633 vdd.n1632 185
R17085 vdd.n1634 vdd.n1633 185
R17086 vdd.n1306 vdd.n1305 185
R17087 vdd.n1310 vdd.n1305 185
R17088 vdd.n1628 vdd.n1627 185
R17089 vdd.n1627 vdd.n1626 185
R17090 vdd.n1309 vdd.n1308 185
R17091 vdd.n1617 vdd.n1309 185
R17092 vdd.n1616 vdd.n1615 185
R17093 vdd.n1618 vdd.n1616 185
R17094 vdd.n1317 vdd.n1316 185
R17095 vdd.n1322 vdd.n1316 185
R17096 vdd.n1611 vdd.n1610 185
R17097 vdd.n1610 vdd.n1609 185
R17098 vdd.n1320 vdd.n1319 185
R17099 vdd.n1321 vdd.n1320 185
R17100 vdd.n1600 vdd.n1599 185
R17101 vdd.n1601 vdd.n1600 185
R17102 vdd.n1330 vdd.n1329 185
R17103 vdd.n1329 vdd.n1328 185
R17104 vdd.n1595 vdd.n1594 185
R17105 vdd.n1594 vdd.n1593 185
R17106 vdd.n1333 vdd.n1332 185
R17107 vdd.n1334 vdd.n1333 185
R17108 vdd.n1584 vdd.n1583 185
R17109 vdd.n1585 vdd.n1584 185
R17110 vdd.n1341 vdd.n1340 185
R17111 vdd.n1345 vdd.n1340 185
R17112 vdd.n1579 vdd.n1578 185
R17113 vdd.n1578 vdd.n1577 185
R17114 vdd.n799 vdd.n797 185
R17115 vdd.n2305 vdd.n797 185
R17116 vdd.n2227 vdd.n817 185
R17117 vdd.n817 vdd.n804 185
R17118 vdd.n2229 vdd.n2228 185
R17119 vdd.n2230 vdd.n2229 185
R17120 vdd.n2226 vdd.n816 185
R17121 vdd.n1166 vdd.n816 185
R17122 vdd.n2225 vdd.n2224 185
R17123 vdd.n2224 vdd.n2223 185
R17124 vdd.n819 vdd.n818 185
R17125 vdd.n820 vdd.n819 185
R17126 vdd.n2214 vdd.n2213 185
R17127 vdd.n2215 vdd.n2214 185
R17128 vdd.n2212 vdd.n830 185
R17129 vdd.n830 vdd.n827 185
R17130 vdd.n2211 vdd.n2210 185
R17131 vdd.n2210 vdd.n2209 185
R17132 vdd.n832 vdd.n831 185
R17133 vdd.n833 vdd.n832 185
R17134 vdd.n2202 vdd.n2201 185
R17135 vdd.n2203 vdd.n2202 185
R17136 vdd.n2200 vdd.n841 185
R17137 vdd.n846 vdd.n841 185
R17138 vdd.n2199 vdd.n2198 185
R17139 vdd.n2198 vdd.n2197 185
R17140 vdd.n843 vdd.n842 185
R17141 vdd.n852 vdd.n843 185
R17142 vdd.n2190 vdd.n2189 185
R17143 vdd.n2191 vdd.n2190 185
R17144 vdd.n2188 vdd.n853 185
R17145 vdd.n1187 vdd.n853 185
R17146 vdd.n2187 vdd.n2186 185
R17147 vdd.n2186 vdd.n2185 185
R17148 vdd.n855 vdd.n854 185
R17149 vdd.n856 vdd.n855 185
R17150 vdd.n2178 vdd.n2177 185
R17151 vdd.n2179 vdd.n2178 185
R17152 vdd.n2176 vdd.n865 185
R17153 vdd.n865 vdd.n862 185
R17154 vdd.n2175 vdd.n2174 185
R17155 vdd.n2174 vdd.n2173 185
R17156 vdd.n867 vdd.n866 185
R17157 vdd.n876 vdd.n867 185
R17158 vdd.n2165 vdd.n2164 185
R17159 vdd.n2166 vdd.n2165 185
R17160 vdd.n2163 vdd.n877 185
R17161 vdd.n883 vdd.n877 185
R17162 vdd.n2162 vdd.n2161 185
R17163 vdd.n2161 vdd.n2160 185
R17164 vdd.n879 vdd.n878 185
R17165 vdd.n880 vdd.n879 185
R17166 vdd.n2153 vdd.n2152 185
R17167 vdd.n2154 vdd.n2153 185
R17168 vdd.n2151 vdd.n890 185
R17169 vdd.n890 vdd.n887 185
R17170 vdd.n2150 vdd.n2149 185
R17171 vdd.n2149 vdd.n2148 185
R17172 vdd.n892 vdd.n891 185
R17173 vdd.n893 vdd.n892 185
R17174 vdd.n2141 vdd.n2140 185
R17175 vdd.n2142 vdd.n2141 185
R17176 vdd.n2139 vdd.n901 185
R17177 vdd.n907 vdd.n901 185
R17178 vdd.n2138 vdd.n2137 185
R17179 vdd.n2137 vdd.n2136 185
R17180 vdd.n903 vdd.n902 185
R17181 vdd.n904 vdd.n903 185
R17182 vdd.n2127 vdd.n2126 185
R17183 vdd.n2125 vdd.n946 185
R17184 vdd.n2124 vdd.n945 185
R17185 vdd.n2129 vdd.n945 185
R17186 vdd.n2123 vdd.n2122 185
R17187 vdd.n2121 vdd.n2120 185
R17188 vdd.n2119 vdd.n2118 185
R17189 vdd.n2117 vdd.n2116 185
R17190 vdd.n2115 vdd.n2114 185
R17191 vdd.n2113 vdd.n2112 185
R17192 vdd.n2111 vdd.n2110 185
R17193 vdd.n2109 vdd.n2108 185
R17194 vdd.n2107 vdd.n2106 185
R17195 vdd.n2105 vdd.n2104 185
R17196 vdd.n2103 vdd.n2102 185
R17197 vdd.n2101 vdd.n2100 185
R17198 vdd.n2099 vdd.n2098 185
R17199 vdd.n2097 vdd.n2096 185
R17200 vdd.n2095 vdd.n2094 185
R17201 vdd.n1103 vdd.n947 185
R17202 vdd.n1105 vdd.n1104 185
R17203 vdd.n1107 vdd.n1106 185
R17204 vdd.n1109 vdd.n1108 185
R17205 vdd.n1111 vdd.n1110 185
R17206 vdd.n1113 vdd.n1112 185
R17207 vdd.n1115 vdd.n1114 185
R17208 vdd.n1117 vdd.n1116 185
R17209 vdd.n1119 vdd.n1118 185
R17210 vdd.n1121 vdd.n1120 185
R17211 vdd.n1123 vdd.n1122 185
R17212 vdd.n1125 vdd.n1124 185
R17213 vdd.n1127 vdd.n1126 185
R17214 vdd.n1129 vdd.n1128 185
R17215 vdd.n1132 vdd.n1131 185
R17216 vdd.n1134 vdd.n1133 185
R17217 vdd.n1136 vdd.n1135 185
R17218 vdd.n2308 vdd.n2307 185
R17219 vdd.n2310 vdd.n2309 185
R17220 vdd.n2312 vdd.n2311 185
R17221 vdd.n2315 vdd.n2314 185
R17222 vdd.n2317 vdd.n2316 185
R17223 vdd.n2319 vdd.n2318 185
R17224 vdd.n2321 vdd.n2320 185
R17225 vdd.n2323 vdd.n2322 185
R17226 vdd.n2325 vdd.n2324 185
R17227 vdd.n2327 vdd.n2326 185
R17228 vdd.n2329 vdd.n2328 185
R17229 vdd.n2331 vdd.n2330 185
R17230 vdd.n2333 vdd.n2332 185
R17231 vdd.n2335 vdd.n2334 185
R17232 vdd.n2337 vdd.n2336 185
R17233 vdd.n2339 vdd.n2338 185
R17234 vdd.n2341 vdd.n2340 185
R17235 vdd.n2343 vdd.n2342 185
R17236 vdd.n2345 vdd.n2344 185
R17237 vdd.n2347 vdd.n2346 185
R17238 vdd.n2349 vdd.n2348 185
R17239 vdd.n2351 vdd.n2350 185
R17240 vdd.n2353 vdd.n2352 185
R17241 vdd.n2355 vdd.n2354 185
R17242 vdd.n2357 vdd.n2356 185
R17243 vdd.n2359 vdd.n2358 185
R17244 vdd.n2361 vdd.n2360 185
R17245 vdd.n2363 vdd.n2362 185
R17246 vdd.n2365 vdd.n2364 185
R17247 vdd.n2367 vdd.n2366 185
R17248 vdd.n2369 vdd.n2368 185
R17249 vdd.n2371 vdd.n2370 185
R17250 vdd.n2373 vdd.n2372 185
R17251 vdd.n2374 vdd.n798 185
R17252 vdd.n2376 vdd.n2375 185
R17253 vdd.n2377 vdd.n2376 185
R17254 vdd.n2306 vdd.n802 185
R17255 vdd.n2306 vdd.n2305 185
R17256 vdd.n1164 vdd.n803 185
R17257 vdd.n804 vdd.n803 185
R17258 vdd.n1165 vdd.n814 185
R17259 vdd.n2230 vdd.n814 185
R17260 vdd.n1168 vdd.n1167 185
R17261 vdd.n1167 vdd.n1166 185
R17262 vdd.n1169 vdd.n821 185
R17263 vdd.n2223 vdd.n821 185
R17264 vdd.n1171 vdd.n1170 185
R17265 vdd.n1170 vdd.n820 185
R17266 vdd.n1172 vdd.n828 185
R17267 vdd.n2215 vdd.n828 185
R17268 vdd.n1174 vdd.n1173 185
R17269 vdd.n1173 vdd.n827 185
R17270 vdd.n1175 vdd.n834 185
R17271 vdd.n2209 vdd.n834 185
R17272 vdd.n1177 vdd.n1176 185
R17273 vdd.n1176 vdd.n833 185
R17274 vdd.n1178 vdd.n839 185
R17275 vdd.n2203 vdd.n839 185
R17276 vdd.n1180 vdd.n1179 185
R17277 vdd.n1179 vdd.n846 185
R17278 vdd.n1181 vdd.n844 185
R17279 vdd.n2197 vdd.n844 185
R17280 vdd.n1183 vdd.n1182 185
R17281 vdd.n1182 vdd.n852 185
R17282 vdd.n1184 vdd.n850 185
R17283 vdd.n2191 vdd.n850 185
R17284 vdd.n1186 vdd.n1185 185
R17285 vdd.n1187 vdd.n1186 185
R17286 vdd.n1163 vdd.n857 185
R17287 vdd.n2185 vdd.n857 185
R17288 vdd.n1162 vdd.n1161 185
R17289 vdd.n1161 vdd.n856 185
R17290 vdd.n1160 vdd.n863 185
R17291 vdd.n2179 vdd.n863 185
R17292 vdd.n1159 vdd.n1158 185
R17293 vdd.n1158 vdd.n862 185
R17294 vdd.n1157 vdd.n868 185
R17295 vdd.n2173 vdd.n868 185
R17296 vdd.n1156 vdd.n1155 185
R17297 vdd.n1155 vdd.n876 185
R17298 vdd.n1154 vdd.n874 185
R17299 vdd.n2166 vdd.n874 185
R17300 vdd.n1153 vdd.n1152 185
R17301 vdd.n1152 vdd.n883 185
R17302 vdd.n1151 vdd.n881 185
R17303 vdd.n2160 vdd.n881 185
R17304 vdd.n1150 vdd.n1149 185
R17305 vdd.n1149 vdd.n880 185
R17306 vdd.n1148 vdd.n888 185
R17307 vdd.n2154 vdd.n888 185
R17308 vdd.n1147 vdd.n1146 185
R17309 vdd.n1146 vdd.n887 185
R17310 vdd.n1145 vdd.n894 185
R17311 vdd.n2148 vdd.n894 185
R17312 vdd.n1144 vdd.n1143 185
R17313 vdd.n1143 vdd.n893 185
R17314 vdd.n1142 vdd.n899 185
R17315 vdd.n2142 vdd.n899 185
R17316 vdd.n1141 vdd.n1140 185
R17317 vdd.n1140 vdd.n907 185
R17318 vdd.n1139 vdd.n905 185
R17319 vdd.n2136 vdd.n905 185
R17320 vdd.n1138 vdd.n1137 185
R17321 vdd.n1137 vdd.n904 185
R17322 vdd.n3229 vdd.n3228 185
R17323 vdd.n3230 vdd.n3229 185
R17324 vdd.n347 vdd.n346 185
R17325 vdd.n3231 vdd.n347 185
R17326 vdd.n3234 vdd.n3233 185
R17327 vdd.n3233 vdd.n3232 185
R17328 vdd.n3235 vdd.n341 185
R17329 vdd.n341 vdd.n340 185
R17330 vdd.n3237 vdd.n3236 185
R17331 vdd.n3238 vdd.n3237 185
R17332 vdd.n336 vdd.n335 185
R17333 vdd.n3239 vdd.n336 185
R17334 vdd.n3242 vdd.n3241 185
R17335 vdd.n3241 vdd.n3240 185
R17336 vdd.n3243 vdd.n330 185
R17337 vdd.n330 vdd.n329 185
R17338 vdd.n3245 vdd.n3244 185
R17339 vdd.n3246 vdd.n3245 185
R17340 vdd.n324 vdd.n323 185
R17341 vdd.n3247 vdd.n324 185
R17342 vdd.n3250 vdd.n3249 185
R17343 vdd.n3249 vdd.n3248 185
R17344 vdd.n3251 vdd.n319 185
R17345 vdd.n325 vdd.n319 185
R17346 vdd.n3253 vdd.n3252 185
R17347 vdd.n3254 vdd.n3253 185
R17348 vdd.n315 vdd.n313 185
R17349 vdd.n3255 vdd.n315 185
R17350 vdd.n3258 vdd.n3257 185
R17351 vdd.n3257 vdd.n3256 185
R17352 vdd.n314 vdd.n312 185
R17353 vdd.n481 vdd.n314 185
R17354 vdd.n3080 vdd.n3079 185
R17355 vdd.n3081 vdd.n3080 185
R17356 vdd.n483 vdd.n482 185
R17357 vdd.n3072 vdd.n482 185
R17358 vdd.n3075 vdd.n3074 185
R17359 vdd.n3074 vdd.n3073 185
R17360 vdd.n486 vdd.n485 185
R17361 vdd.n493 vdd.n486 185
R17362 vdd.n3063 vdd.n3062 185
R17363 vdd.n3064 vdd.n3063 185
R17364 vdd.n495 vdd.n494 185
R17365 vdd.n494 vdd.n492 185
R17366 vdd.n3058 vdd.n3057 185
R17367 vdd.n3057 vdd.n3056 185
R17368 vdd.n498 vdd.n497 185
R17369 vdd.n499 vdd.n498 185
R17370 vdd.n3047 vdd.n3046 185
R17371 vdd.n3048 vdd.n3047 185
R17372 vdd.n507 vdd.n506 185
R17373 vdd.n506 vdd.n505 185
R17374 vdd.n3042 vdd.n3041 185
R17375 vdd.n3041 vdd.n3040 185
R17376 vdd.n510 vdd.n509 185
R17377 vdd.n511 vdd.n510 185
R17378 vdd.n3031 vdd.n3030 185
R17379 vdd.n3032 vdd.n3031 185
R17380 vdd.n3027 vdd.n517 185
R17381 vdd.n3026 vdd.n3025 185
R17382 vdd.n3023 vdd.n519 185
R17383 vdd.n3023 vdd.n516 185
R17384 vdd.n3022 vdd.n3021 185
R17385 vdd.n3020 vdd.n3019 185
R17386 vdd.n3018 vdd.n3017 185
R17387 vdd.n3016 vdd.n3015 185
R17388 vdd.n3014 vdd.n525 185
R17389 vdd.n3012 vdd.n3011 185
R17390 vdd.n3010 vdd.n526 185
R17391 vdd.n3009 vdd.n3008 185
R17392 vdd.n3006 vdd.n531 185
R17393 vdd.n3004 vdd.n3003 185
R17394 vdd.n3002 vdd.n532 185
R17395 vdd.n3001 vdd.n3000 185
R17396 vdd.n2998 vdd.n537 185
R17397 vdd.n2996 vdd.n2995 185
R17398 vdd.n2994 vdd.n538 185
R17399 vdd.n2993 vdd.n2992 185
R17400 vdd.n2990 vdd.n545 185
R17401 vdd.n2988 vdd.n2987 185
R17402 vdd.n2986 vdd.n546 185
R17403 vdd.n2985 vdd.n2984 185
R17404 vdd.n2982 vdd.n551 185
R17405 vdd.n2980 vdd.n2979 185
R17406 vdd.n2978 vdd.n552 185
R17407 vdd.n2977 vdd.n2976 185
R17408 vdd.n2974 vdd.n557 185
R17409 vdd.n2972 vdd.n2971 185
R17410 vdd.n2970 vdd.n558 185
R17411 vdd.n2969 vdd.n2968 185
R17412 vdd.n2966 vdd.n563 185
R17413 vdd.n2964 vdd.n2963 185
R17414 vdd.n2962 vdd.n564 185
R17415 vdd.n2961 vdd.n2960 185
R17416 vdd.n2958 vdd.n569 185
R17417 vdd.n2956 vdd.n2955 185
R17418 vdd.n2954 vdd.n570 185
R17419 vdd.n2953 vdd.n2952 185
R17420 vdd.n2950 vdd.n575 185
R17421 vdd.n2948 vdd.n2947 185
R17422 vdd.n2946 vdd.n576 185
R17423 vdd.n585 vdd.n579 185
R17424 vdd.n2942 vdd.n2941 185
R17425 vdd.n2939 vdd.n583 185
R17426 vdd.n2938 vdd.n2937 185
R17427 vdd.n2936 vdd.n2935 185
R17428 vdd.n2934 vdd.n589 185
R17429 vdd.n2932 vdd.n2931 185
R17430 vdd.n2930 vdd.n590 185
R17431 vdd.n2929 vdd.n2928 185
R17432 vdd.n2926 vdd.n595 185
R17433 vdd.n2924 vdd.n2923 185
R17434 vdd.n2922 vdd.n596 185
R17435 vdd.n2921 vdd.n2920 185
R17436 vdd.n2918 vdd.n601 185
R17437 vdd.n2916 vdd.n2915 185
R17438 vdd.n2914 vdd.n602 185
R17439 vdd.n2913 vdd.n2912 185
R17440 vdd.n2910 vdd.n2909 185
R17441 vdd.n2908 vdd.n2907 185
R17442 vdd.n2906 vdd.n2905 185
R17443 vdd.n2904 vdd.n2903 185
R17444 vdd.n2899 vdd.n515 185
R17445 vdd.n516 vdd.n515 185
R17446 vdd.n3112 vdd.n3111 185
R17447 vdd.n3116 vdd.n462 185
R17448 vdd.n3118 vdd.n3117 185
R17449 vdd.n3120 vdd.n460 185
R17450 vdd.n3122 vdd.n3121 185
R17451 vdd.n3123 vdd.n455 185
R17452 vdd.n3125 vdd.n3124 185
R17453 vdd.n3127 vdd.n453 185
R17454 vdd.n3129 vdd.n3128 185
R17455 vdd.n3130 vdd.n448 185
R17456 vdd.n3132 vdd.n3131 185
R17457 vdd.n3134 vdd.n446 185
R17458 vdd.n3136 vdd.n3135 185
R17459 vdd.n3137 vdd.n441 185
R17460 vdd.n3139 vdd.n3138 185
R17461 vdd.n3141 vdd.n439 185
R17462 vdd.n3143 vdd.n3142 185
R17463 vdd.n3144 vdd.n435 185
R17464 vdd.n3146 vdd.n3145 185
R17465 vdd.n3148 vdd.n432 185
R17466 vdd.n3150 vdd.n3149 185
R17467 vdd.n433 vdd.n426 185
R17468 vdd.n3154 vdd.n430 185
R17469 vdd.n3155 vdd.n422 185
R17470 vdd.n3157 vdd.n3156 185
R17471 vdd.n3159 vdd.n420 185
R17472 vdd.n3161 vdd.n3160 185
R17473 vdd.n3162 vdd.n415 185
R17474 vdd.n3164 vdd.n3163 185
R17475 vdd.n3166 vdd.n413 185
R17476 vdd.n3168 vdd.n3167 185
R17477 vdd.n3169 vdd.n408 185
R17478 vdd.n3171 vdd.n3170 185
R17479 vdd.n3173 vdd.n406 185
R17480 vdd.n3175 vdd.n3174 185
R17481 vdd.n3176 vdd.n401 185
R17482 vdd.n3178 vdd.n3177 185
R17483 vdd.n3180 vdd.n399 185
R17484 vdd.n3182 vdd.n3181 185
R17485 vdd.n3183 vdd.n395 185
R17486 vdd.n3185 vdd.n3184 185
R17487 vdd.n3187 vdd.n392 185
R17488 vdd.n3189 vdd.n3188 185
R17489 vdd.n393 vdd.n386 185
R17490 vdd.n3193 vdd.n390 185
R17491 vdd.n3194 vdd.n382 185
R17492 vdd.n3196 vdd.n3195 185
R17493 vdd.n3198 vdd.n380 185
R17494 vdd.n3200 vdd.n3199 185
R17495 vdd.n3201 vdd.n375 185
R17496 vdd.n3203 vdd.n3202 185
R17497 vdd.n3205 vdd.n373 185
R17498 vdd.n3207 vdd.n3206 185
R17499 vdd.n3208 vdd.n368 185
R17500 vdd.n3210 vdd.n3209 185
R17501 vdd.n3212 vdd.n366 185
R17502 vdd.n3214 vdd.n3213 185
R17503 vdd.n3215 vdd.n360 185
R17504 vdd.n3217 vdd.n3216 185
R17505 vdd.n3219 vdd.n359 185
R17506 vdd.n3220 vdd.n358 185
R17507 vdd.n3223 vdd.n3222 185
R17508 vdd.n3224 vdd.n356 185
R17509 vdd.n3225 vdd.n352 185
R17510 vdd.n3107 vdd.n350 185
R17511 vdd.n3230 vdd.n350 185
R17512 vdd.n3106 vdd.n349 185
R17513 vdd.n3231 vdd.n349 185
R17514 vdd.n3105 vdd.n348 185
R17515 vdd.n3232 vdd.n348 185
R17516 vdd.n468 vdd.n467 185
R17517 vdd.n467 vdd.n340 185
R17518 vdd.n3101 vdd.n339 185
R17519 vdd.n3238 vdd.n339 185
R17520 vdd.n3100 vdd.n338 185
R17521 vdd.n3239 vdd.n338 185
R17522 vdd.n3099 vdd.n337 185
R17523 vdd.n3240 vdd.n337 185
R17524 vdd.n471 vdd.n470 185
R17525 vdd.n470 vdd.n329 185
R17526 vdd.n3095 vdd.n328 185
R17527 vdd.n3246 vdd.n328 185
R17528 vdd.n3094 vdd.n327 185
R17529 vdd.n3247 vdd.n327 185
R17530 vdd.n3093 vdd.n326 185
R17531 vdd.n3248 vdd.n326 185
R17532 vdd.n474 vdd.n473 185
R17533 vdd.n473 vdd.n325 185
R17534 vdd.n3089 vdd.n318 185
R17535 vdd.n3254 vdd.n318 185
R17536 vdd.n3088 vdd.n317 185
R17537 vdd.n3255 vdd.n317 185
R17538 vdd.n3087 vdd.n316 185
R17539 vdd.n3256 vdd.n316 185
R17540 vdd.n480 vdd.n476 185
R17541 vdd.n481 vdd.n480 185
R17542 vdd.n3083 vdd.n3082 185
R17543 vdd.n3082 vdd.n3081 185
R17544 vdd.n479 vdd.n478 185
R17545 vdd.n3072 vdd.n479 185
R17546 vdd.n3071 vdd.n3070 185
R17547 vdd.n3073 vdd.n3071 185
R17548 vdd.n488 vdd.n487 185
R17549 vdd.n493 vdd.n487 185
R17550 vdd.n3066 vdd.n3065 185
R17551 vdd.n3065 vdd.n3064 185
R17552 vdd.n491 vdd.n490 185
R17553 vdd.n492 vdd.n491 185
R17554 vdd.n3055 vdd.n3054 185
R17555 vdd.n3056 vdd.n3055 185
R17556 vdd.n501 vdd.n500 185
R17557 vdd.n500 vdd.n499 185
R17558 vdd.n3050 vdd.n3049 185
R17559 vdd.n3049 vdd.n3048 185
R17560 vdd.n504 vdd.n503 185
R17561 vdd.n505 vdd.n504 185
R17562 vdd.n3039 vdd.n3038 185
R17563 vdd.n3040 vdd.n3039 185
R17564 vdd.n513 vdd.n512 185
R17565 vdd.n512 vdd.n511 185
R17566 vdd.n3034 vdd.n3033 185
R17567 vdd.n3033 vdd.n3032 185
R17568 vdd.n2648 vdd.n2647 185
R17569 vdd.n2646 vdd.n2412 185
R17570 vdd.n2645 vdd.n2411 185
R17571 vdd.n2650 vdd.n2411 185
R17572 vdd.n2644 vdd.n2643 185
R17573 vdd.n2642 vdd.n2641 185
R17574 vdd.n2640 vdd.n2639 185
R17575 vdd.n2638 vdd.n2637 185
R17576 vdd.n2636 vdd.n2635 185
R17577 vdd.n2634 vdd.n2633 185
R17578 vdd.n2632 vdd.n2631 185
R17579 vdd.n2630 vdd.n2629 185
R17580 vdd.n2628 vdd.n2627 185
R17581 vdd.n2626 vdd.n2625 185
R17582 vdd.n2624 vdd.n2623 185
R17583 vdd.n2622 vdd.n2621 185
R17584 vdd.n2620 vdd.n2619 185
R17585 vdd.n2618 vdd.n2617 185
R17586 vdd.n2616 vdd.n2615 185
R17587 vdd.n2614 vdd.n2613 185
R17588 vdd.n2612 vdd.n2611 185
R17589 vdd.n2610 vdd.n2609 185
R17590 vdd.n2608 vdd.n2607 185
R17591 vdd.n2606 vdd.n2605 185
R17592 vdd.n2604 vdd.n2603 185
R17593 vdd.n2602 vdd.n2601 185
R17594 vdd.n2600 vdd.n2599 185
R17595 vdd.n2598 vdd.n2597 185
R17596 vdd.n2596 vdd.n2595 185
R17597 vdd.n2594 vdd.n2593 185
R17598 vdd.n2592 vdd.n2591 185
R17599 vdd.n2590 vdd.n2589 185
R17600 vdd.n2588 vdd.n2587 185
R17601 vdd.n2585 vdd.n2584 185
R17602 vdd.n2583 vdd.n2582 185
R17603 vdd.n2581 vdd.n2580 185
R17604 vdd.n2800 vdd.n2799 185
R17605 vdd.n2801 vdd.n660 185
R17606 vdd.n2803 vdd.n2802 185
R17607 vdd.n2805 vdd.n658 185
R17608 vdd.n2807 vdd.n2806 185
R17609 vdd.n2808 vdd.n657 185
R17610 vdd.n2810 vdd.n2809 185
R17611 vdd.n2812 vdd.n655 185
R17612 vdd.n2814 vdd.n2813 185
R17613 vdd.n2815 vdd.n654 185
R17614 vdd.n2817 vdd.n2816 185
R17615 vdd.n2819 vdd.n652 185
R17616 vdd.n2821 vdd.n2820 185
R17617 vdd.n2822 vdd.n651 185
R17618 vdd.n2824 vdd.n2823 185
R17619 vdd.n2826 vdd.n649 185
R17620 vdd.n2828 vdd.n2827 185
R17621 vdd.n2830 vdd.n648 185
R17622 vdd.n2832 vdd.n2831 185
R17623 vdd.n2834 vdd.n646 185
R17624 vdd.n2836 vdd.n2835 185
R17625 vdd.n2837 vdd.n645 185
R17626 vdd.n2839 vdd.n2838 185
R17627 vdd.n2841 vdd.n643 185
R17628 vdd.n2843 vdd.n2842 185
R17629 vdd.n2844 vdd.n642 185
R17630 vdd.n2846 vdd.n2845 185
R17631 vdd.n2848 vdd.n640 185
R17632 vdd.n2850 vdd.n2849 185
R17633 vdd.n2851 vdd.n639 185
R17634 vdd.n2853 vdd.n2852 185
R17635 vdd.n2855 vdd.n638 185
R17636 vdd.n2856 vdd.n637 185
R17637 vdd.n2859 vdd.n2858 185
R17638 vdd.n2860 vdd.n635 185
R17639 vdd.n635 vdd.n613 185
R17640 vdd.n2797 vdd.n632 185
R17641 vdd.n2863 vdd.n632 185
R17642 vdd.n2796 vdd.n2795 185
R17643 vdd.n2795 vdd.n631 185
R17644 vdd.n2794 vdd.n664 185
R17645 vdd.n2794 vdd.n2793 185
R17646 vdd.n2528 vdd.n665 185
R17647 vdd.n674 vdd.n665 185
R17648 vdd.n2529 vdd.n672 185
R17649 vdd.n2787 vdd.n672 185
R17650 vdd.n2531 vdd.n2530 185
R17651 vdd.n2530 vdd.n671 185
R17652 vdd.n2532 vdd.n680 185
R17653 vdd.n2736 vdd.n680 185
R17654 vdd.n2534 vdd.n2533 185
R17655 vdd.n2533 vdd.n679 185
R17656 vdd.n2535 vdd.n686 185
R17657 vdd.n2730 vdd.n686 185
R17658 vdd.n2537 vdd.n2536 185
R17659 vdd.n2536 vdd.n685 185
R17660 vdd.n2538 vdd.n691 185
R17661 vdd.n2724 vdd.n691 185
R17662 vdd.n2540 vdd.n2539 185
R17663 vdd.n2539 vdd.n698 185
R17664 vdd.n2541 vdd.n696 185
R17665 vdd.n2718 vdd.n696 185
R17666 vdd.n2543 vdd.n2542 185
R17667 vdd.n2542 vdd.n706 185
R17668 vdd.n2544 vdd.n704 185
R17669 vdd.n2711 vdd.n704 185
R17670 vdd.n2546 vdd.n2545 185
R17671 vdd.n2545 vdd.n703 185
R17672 vdd.n2547 vdd.n711 185
R17673 vdd.n2705 vdd.n711 185
R17674 vdd.n2549 vdd.n2548 185
R17675 vdd.n2548 vdd.n710 185
R17676 vdd.n2550 vdd.n716 185
R17677 vdd.n2699 vdd.n716 185
R17678 vdd.n2552 vdd.n2551 185
R17679 vdd.n2551 vdd.n723 185
R17680 vdd.n2553 vdd.n721 185
R17681 vdd.n2693 vdd.n721 185
R17682 vdd.n2555 vdd.n2554 185
R17683 vdd.n2554 vdd.n729 185
R17684 vdd.n2556 vdd.n727 185
R17685 vdd.n2687 vdd.n727 185
R17686 vdd.n2558 vdd.n2557 185
R17687 vdd.n2559 vdd.n2558 185
R17688 vdd.n2527 vdd.n734 185
R17689 vdd.n2681 vdd.n734 185
R17690 vdd.n2526 vdd.n2525 185
R17691 vdd.n2525 vdd.n733 185
R17692 vdd.n2524 vdd.n740 185
R17693 vdd.n2675 vdd.n740 185
R17694 vdd.n2523 vdd.n2522 185
R17695 vdd.n2522 vdd.n739 185
R17696 vdd.n2521 vdd.n746 185
R17697 vdd.n2669 vdd.n746 185
R17698 vdd.n2520 vdd.n2519 185
R17699 vdd.n2519 vdd.n745 185
R17700 vdd.n2415 vdd.n751 185
R17701 vdd.n2663 vdd.n751 185
R17702 vdd.n2576 vdd.n2575 185
R17703 vdd.n2575 vdd.n2574 185
R17704 vdd.n2577 vdd.n757 185
R17705 vdd.n2657 vdd.n757 185
R17706 vdd.n2579 vdd.n2578 185
R17707 vdd.n2579 vdd.n756 185
R17708 vdd.n755 vdd.n754 185
R17709 vdd.n756 vdd.n755 185
R17710 vdd.n2659 vdd.n2658 185
R17711 vdd.n2658 vdd.n2657 185
R17712 vdd.n2660 vdd.n753 185
R17713 vdd.n2574 vdd.n753 185
R17714 vdd.n2662 vdd.n2661 185
R17715 vdd.n2663 vdd.n2662 185
R17716 vdd.n744 vdd.n743 185
R17717 vdd.n745 vdd.n744 185
R17718 vdd.n2671 vdd.n2670 185
R17719 vdd.n2670 vdd.n2669 185
R17720 vdd.n2672 vdd.n742 185
R17721 vdd.n742 vdd.n739 185
R17722 vdd.n2674 vdd.n2673 185
R17723 vdd.n2675 vdd.n2674 185
R17724 vdd.n732 vdd.n731 185
R17725 vdd.n733 vdd.n732 185
R17726 vdd.n2683 vdd.n2682 185
R17727 vdd.n2682 vdd.n2681 185
R17728 vdd.n2684 vdd.n730 185
R17729 vdd.n2559 vdd.n730 185
R17730 vdd.n2686 vdd.n2685 185
R17731 vdd.n2687 vdd.n2686 185
R17732 vdd.n720 vdd.n719 185
R17733 vdd.n729 vdd.n720 185
R17734 vdd.n2695 vdd.n2694 185
R17735 vdd.n2694 vdd.n2693 185
R17736 vdd.n2696 vdd.n718 185
R17737 vdd.n723 vdd.n718 185
R17738 vdd.n2698 vdd.n2697 185
R17739 vdd.n2699 vdd.n2698 185
R17740 vdd.n709 vdd.n708 185
R17741 vdd.n710 vdd.n709 185
R17742 vdd.n2707 vdd.n2706 185
R17743 vdd.n2706 vdd.n2705 185
R17744 vdd.n2708 vdd.n707 185
R17745 vdd.n707 vdd.n703 185
R17746 vdd.n2710 vdd.n2709 185
R17747 vdd.n2711 vdd.n2710 185
R17748 vdd.n695 vdd.n694 185
R17749 vdd.n706 vdd.n695 185
R17750 vdd.n2720 vdd.n2719 185
R17751 vdd.n2719 vdd.n2718 185
R17752 vdd.n2721 vdd.n693 185
R17753 vdd.n698 vdd.n693 185
R17754 vdd.n2723 vdd.n2722 185
R17755 vdd.n2724 vdd.n2723 185
R17756 vdd.n684 vdd.n683 185
R17757 vdd.n685 vdd.n684 185
R17758 vdd.n2732 vdd.n2731 185
R17759 vdd.n2731 vdd.n2730 185
R17760 vdd.n2733 vdd.n682 185
R17761 vdd.n682 vdd.n679 185
R17762 vdd.n2735 vdd.n2734 185
R17763 vdd.n2736 vdd.n2735 185
R17764 vdd.n670 vdd.n669 185
R17765 vdd.n671 vdd.n670 185
R17766 vdd.n2789 vdd.n2788 185
R17767 vdd.n2788 vdd.n2787 185
R17768 vdd.n2790 vdd.n668 185
R17769 vdd.n674 vdd.n668 185
R17770 vdd.n2792 vdd.n2791 185
R17771 vdd.n2793 vdd.n2792 185
R17772 vdd.n636 vdd.n634 185
R17773 vdd.n634 vdd.n631 185
R17774 vdd.n2862 vdd.n2861 185
R17775 vdd.n2863 vdd.n2862 185
R17776 vdd.n2304 vdd.n2303 185
R17777 vdd.n2305 vdd.n2304 185
R17778 vdd.n808 vdd.n806 185
R17779 vdd.n806 vdd.n804 185
R17780 vdd.n2219 vdd.n815 185
R17781 vdd.n2230 vdd.n815 185
R17782 vdd.n2220 vdd.n824 185
R17783 vdd.n1166 vdd.n824 185
R17784 vdd.n2222 vdd.n2221 185
R17785 vdd.n2223 vdd.n2222 185
R17786 vdd.n2218 vdd.n823 185
R17787 vdd.n823 vdd.n820 185
R17788 vdd.n2217 vdd.n2216 185
R17789 vdd.n2216 vdd.n2215 185
R17790 vdd.n826 vdd.n825 185
R17791 vdd.n827 vdd.n826 185
R17792 vdd.n2208 vdd.n2207 185
R17793 vdd.n2209 vdd.n2208 185
R17794 vdd.n2206 vdd.n836 185
R17795 vdd.n836 vdd.n833 185
R17796 vdd.n2205 vdd.n2204 185
R17797 vdd.n2204 vdd.n2203 185
R17798 vdd.n838 vdd.n837 185
R17799 vdd.n846 vdd.n838 185
R17800 vdd.n2196 vdd.n2195 185
R17801 vdd.n2197 vdd.n2196 185
R17802 vdd.n2194 vdd.n847 185
R17803 vdd.n852 vdd.n847 185
R17804 vdd.n2193 vdd.n2192 185
R17805 vdd.n2192 vdd.n2191 185
R17806 vdd.n849 vdd.n848 185
R17807 vdd.n1187 vdd.n849 185
R17808 vdd.n2184 vdd.n2183 185
R17809 vdd.n2185 vdd.n2184 185
R17810 vdd.n2182 vdd.n859 185
R17811 vdd.n859 vdd.n856 185
R17812 vdd.n2181 vdd.n2180 185
R17813 vdd.n2180 vdd.n2179 185
R17814 vdd.n861 vdd.n860 185
R17815 vdd.n862 vdd.n861 185
R17816 vdd.n2172 vdd.n2171 185
R17817 vdd.n2173 vdd.n2172 185
R17818 vdd.n2169 vdd.n870 185
R17819 vdd.n876 vdd.n870 185
R17820 vdd.n2168 vdd.n2167 185
R17821 vdd.n2167 vdd.n2166 185
R17822 vdd.n873 vdd.n872 185
R17823 vdd.n883 vdd.n873 185
R17824 vdd.n2159 vdd.n2158 185
R17825 vdd.n2160 vdd.n2159 185
R17826 vdd.n2157 vdd.n884 185
R17827 vdd.n884 vdd.n880 185
R17828 vdd.n2156 vdd.n2155 185
R17829 vdd.n2155 vdd.n2154 185
R17830 vdd.n886 vdd.n885 185
R17831 vdd.n887 vdd.n886 185
R17832 vdd.n2147 vdd.n2146 185
R17833 vdd.n2148 vdd.n2147 185
R17834 vdd.n2145 vdd.n896 185
R17835 vdd.n896 vdd.n893 185
R17836 vdd.n2144 vdd.n2143 185
R17837 vdd.n2143 vdd.n2142 185
R17838 vdd.n898 vdd.n897 185
R17839 vdd.n907 vdd.n898 185
R17840 vdd.n2135 vdd.n2134 185
R17841 vdd.n2136 vdd.n2135 185
R17842 vdd.n2133 vdd.n908 185
R17843 vdd.n908 vdd.n904 185
R17844 vdd.n2235 vdd.n779 185
R17845 vdd.n2377 vdd.n779 185
R17846 vdd.n2237 vdd.n2236 185
R17847 vdd.n2239 vdd.n2238 185
R17848 vdd.n2241 vdd.n2240 185
R17849 vdd.n2243 vdd.n2242 185
R17850 vdd.n2245 vdd.n2244 185
R17851 vdd.n2247 vdd.n2246 185
R17852 vdd.n2249 vdd.n2248 185
R17853 vdd.n2251 vdd.n2250 185
R17854 vdd.n2253 vdd.n2252 185
R17855 vdd.n2255 vdd.n2254 185
R17856 vdd.n2257 vdd.n2256 185
R17857 vdd.n2259 vdd.n2258 185
R17858 vdd.n2261 vdd.n2260 185
R17859 vdd.n2263 vdd.n2262 185
R17860 vdd.n2265 vdd.n2264 185
R17861 vdd.n2267 vdd.n2266 185
R17862 vdd.n2269 vdd.n2268 185
R17863 vdd.n2271 vdd.n2270 185
R17864 vdd.n2273 vdd.n2272 185
R17865 vdd.n2275 vdd.n2274 185
R17866 vdd.n2277 vdd.n2276 185
R17867 vdd.n2279 vdd.n2278 185
R17868 vdd.n2281 vdd.n2280 185
R17869 vdd.n2283 vdd.n2282 185
R17870 vdd.n2285 vdd.n2284 185
R17871 vdd.n2287 vdd.n2286 185
R17872 vdd.n2289 vdd.n2288 185
R17873 vdd.n2291 vdd.n2290 185
R17874 vdd.n2293 vdd.n2292 185
R17875 vdd.n2295 vdd.n2294 185
R17876 vdd.n2297 vdd.n2296 185
R17877 vdd.n2299 vdd.n2298 185
R17878 vdd.n2301 vdd.n2300 185
R17879 vdd.n2302 vdd.n807 185
R17880 vdd.n2234 vdd.n805 185
R17881 vdd.n2305 vdd.n805 185
R17882 vdd.n2233 vdd.n2232 185
R17883 vdd.n2232 vdd.n804 185
R17884 vdd.n2231 vdd.n812 185
R17885 vdd.n2231 vdd.n2230 185
R17886 vdd.n1084 vdd.n813 185
R17887 vdd.n1166 vdd.n813 185
R17888 vdd.n1085 vdd.n822 185
R17889 vdd.n2223 vdd.n822 185
R17890 vdd.n1087 vdd.n1086 185
R17891 vdd.n1086 vdd.n820 185
R17892 vdd.n1088 vdd.n829 185
R17893 vdd.n2215 vdd.n829 185
R17894 vdd.n1090 vdd.n1089 185
R17895 vdd.n1089 vdd.n827 185
R17896 vdd.n1091 vdd.n835 185
R17897 vdd.n2209 vdd.n835 185
R17898 vdd.n1093 vdd.n1092 185
R17899 vdd.n1092 vdd.n833 185
R17900 vdd.n1094 vdd.n840 185
R17901 vdd.n2203 vdd.n840 185
R17902 vdd.n1096 vdd.n1095 185
R17903 vdd.n1095 vdd.n846 185
R17904 vdd.n1097 vdd.n845 185
R17905 vdd.n2197 vdd.n845 185
R17906 vdd.n1099 vdd.n1098 185
R17907 vdd.n1098 vdd.n852 185
R17908 vdd.n1100 vdd.n851 185
R17909 vdd.n2191 vdd.n851 185
R17910 vdd.n1189 vdd.n1188 185
R17911 vdd.n1188 vdd.n1187 185
R17912 vdd.n1190 vdd.n858 185
R17913 vdd.n2185 vdd.n858 185
R17914 vdd.n1192 vdd.n1191 185
R17915 vdd.n1191 vdd.n856 185
R17916 vdd.n1193 vdd.n864 185
R17917 vdd.n2179 vdd.n864 185
R17918 vdd.n1195 vdd.n1194 185
R17919 vdd.n1194 vdd.n862 185
R17920 vdd.n1196 vdd.n869 185
R17921 vdd.n2173 vdd.n869 185
R17922 vdd.n1198 vdd.n1197 185
R17923 vdd.n1197 vdd.n876 185
R17924 vdd.n1199 vdd.n875 185
R17925 vdd.n2166 vdd.n875 185
R17926 vdd.n1201 vdd.n1200 185
R17927 vdd.n1200 vdd.n883 185
R17928 vdd.n1202 vdd.n882 185
R17929 vdd.n2160 vdd.n882 185
R17930 vdd.n1204 vdd.n1203 185
R17931 vdd.n1203 vdd.n880 185
R17932 vdd.n1205 vdd.n889 185
R17933 vdd.n2154 vdd.n889 185
R17934 vdd.n1207 vdd.n1206 185
R17935 vdd.n1206 vdd.n887 185
R17936 vdd.n1208 vdd.n895 185
R17937 vdd.n2148 vdd.n895 185
R17938 vdd.n1210 vdd.n1209 185
R17939 vdd.n1209 vdd.n893 185
R17940 vdd.n1211 vdd.n900 185
R17941 vdd.n2142 vdd.n900 185
R17942 vdd.n1213 vdd.n1212 185
R17943 vdd.n1212 vdd.n907 185
R17944 vdd.n1214 vdd.n906 185
R17945 vdd.n2136 vdd.n906 185
R17946 vdd.n1216 vdd.n1215 185
R17947 vdd.n1215 vdd.n904 185
R17948 vdd.n2132 vdd.n2131 185
R17949 vdd.n910 vdd.n909 185
R17950 vdd.n1051 vdd.n1050 185
R17951 vdd.n1053 vdd.n1052 185
R17952 vdd.n1055 vdd.n1054 185
R17953 vdd.n1057 vdd.n1056 185
R17954 vdd.n1059 vdd.n1058 185
R17955 vdd.n1061 vdd.n1060 185
R17956 vdd.n1063 vdd.n1062 185
R17957 vdd.n1065 vdd.n1064 185
R17958 vdd.n1067 vdd.n1066 185
R17959 vdd.n1069 vdd.n1068 185
R17960 vdd.n1071 vdd.n1070 185
R17961 vdd.n1073 vdd.n1072 185
R17962 vdd.n1075 vdd.n1074 185
R17963 vdd.n1077 vdd.n1076 185
R17964 vdd.n1079 vdd.n1078 185
R17965 vdd.n1250 vdd.n1080 185
R17966 vdd.n1249 vdd.n1248 185
R17967 vdd.n1247 vdd.n1246 185
R17968 vdd.n1245 vdd.n1244 185
R17969 vdd.n1243 vdd.n1242 185
R17970 vdd.n1241 vdd.n1240 185
R17971 vdd.n1239 vdd.n1238 185
R17972 vdd.n1237 vdd.n1236 185
R17973 vdd.n1235 vdd.n1234 185
R17974 vdd.n1233 vdd.n1232 185
R17975 vdd.n1231 vdd.n1230 185
R17976 vdd.n1229 vdd.n1228 185
R17977 vdd.n1227 vdd.n1226 185
R17978 vdd.n1225 vdd.n1224 185
R17979 vdd.n1223 vdd.n1222 185
R17980 vdd.n1221 vdd.n1220 185
R17981 vdd.n1219 vdd.n1218 185
R17982 vdd.n1217 vdd.n944 185
R17983 vdd.n2129 vdd.n944 185
R17984 vdd.n2129 vdd.n911 179.345
R17985 vdd.n613 vdd.n516 179.345
R17986 vdd.n303 vdd.n302 171.744
R17987 vdd.n302 vdd.n301 171.744
R17988 vdd.n301 vdd.n270 171.744
R17989 vdd.n294 vdd.n270 171.744
R17990 vdd.n294 vdd.n293 171.744
R17991 vdd.n293 vdd.n275 171.744
R17992 vdd.n286 vdd.n275 171.744
R17993 vdd.n286 vdd.n285 171.744
R17994 vdd.n285 vdd.n279 171.744
R17995 vdd.n252 vdd.n251 171.744
R17996 vdd.n251 vdd.n250 171.744
R17997 vdd.n250 vdd.n219 171.744
R17998 vdd.n243 vdd.n219 171.744
R17999 vdd.n243 vdd.n242 171.744
R18000 vdd.n242 vdd.n224 171.744
R18001 vdd.n235 vdd.n224 171.744
R18002 vdd.n235 vdd.n234 171.744
R18003 vdd.n234 vdd.n228 171.744
R18004 vdd.n209 vdd.n208 171.744
R18005 vdd.n208 vdd.n207 171.744
R18006 vdd.n207 vdd.n176 171.744
R18007 vdd.n200 vdd.n176 171.744
R18008 vdd.n200 vdd.n199 171.744
R18009 vdd.n199 vdd.n181 171.744
R18010 vdd.n192 vdd.n181 171.744
R18011 vdd.n192 vdd.n191 171.744
R18012 vdd.n191 vdd.n185 171.744
R18013 vdd.n158 vdd.n157 171.744
R18014 vdd.n157 vdd.n156 171.744
R18015 vdd.n156 vdd.n125 171.744
R18016 vdd.n149 vdd.n125 171.744
R18017 vdd.n149 vdd.n148 171.744
R18018 vdd.n148 vdd.n130 171.744
R18019 vdd.n141 vdd.n130 171.744
R18020 vdd.n141 vdd.n140 171.744
R18021 vdd.n140 vdd.n134 171.744
R18022 vdd.n116 vdd.n115 171.744
R18023 vdd.n115 vdd.n114 171.744
R18024 vdd.n114 vdd.n83 171.744
R18025 vdd.n107 vdd.n83 171.744
R18026 vdd.n107 vdd.n106 171.744
R18027 vdd.n106 vdd.n88 171.744
R18028 vdd.n99 vdd.n88 171.744
R18029 vdd.n99 vdd.n98 171.744
R18030 vdd.n98 vdd.n92 171.744
R18031 vdd.n65 vdd.n64 171.744
R18032 vdd.n64 vdd.n63 171.744
R18033 vdd.n63 vdd.n32 171.744
R18034 vdd.n56 vdd.n32 171.744
R18035 vdd.n56 vdd.n55 171.744
R18036 vdd.n55 vdd.n37 171.744
R18037 vdd.n48 vdd.n37 171.744
R18038 vdd.n48 vdd.n47 171.744
R18039 vdd.n47 vdd.n41 171.744
R18040 vdd.n1860 vdd.n1859 171.744
R18041 vdd.n1859 vdd.n1858 171.744
R18042 vdd.n1858 vdd.n1827 171.744
R18043 vdd.n1851 vdd.n1827 171.744
R18044 vdd.n1851 vdd.n1850 171.744
R18045 vdd.n1850 vdd.n1832 171.744
R18046 vdd.n1843 vdd.n1832 171.744
R18047 vdd.n1843 vdd.n1842 171.744
R18048 vdd.n1842 vdd.n1836 171.744
R18049 vdd.n1911 vdd.n1910 171.744
R18050 vdd.n1910 vdd.n1909 171.744
R18051 vdd.n1909 vdd.n1878 171.744
R18052 vdd.n1902 vdd.n1878 171.744
R18053 vdd.n1902 vdd.n1901 171.744
R18054 vdd.n1901 vdd.n1883 171.744
R18055 vdd.n1894 vdd.n1883 171.744
R18056 vdd.n1894 vdd.n1893 171.744
R18057 vdd.n1893 vdd.n1887 171.744
R18058 vdd.n1766 vdd.n1765 171.744
R18059 vdd.n1765 vdd.n1764 171.744
R18060 vdd.n1764 vdd.n1733 171.744
R18061 vdd.n1757 vdd.n1733 171.744
R18062 vdd.n1757 vdd.n1756 171.744
R18063 vdd.n1756 vdd.n1738 171.744
R18064 vdd.n1749 vdd.n1738 171.744
R18065 vdd.n1749 vdd.n1748 171.744
R18066 vdd.n1748 vdd.n1742 171.744
R18067 vdd.n1817 vdd.n1816 171.744
R18068 vdd.n1816 vdd.n1815 171.744
R18069 vdd.n1815 vdd.n1784 171.744
R18070 vdd.n1808 vdd.n1784 171.744
R18071 vdd.n1808 vdd.n1807 171.744
R18072 vdd.n1807 vdd.n1789 171.744
R18073 vdd.n1800 vdd.n1789 171.744
R18074 vdd.n1800 vdd.n1799 171.744
R18075 vdd.n1799 vdd.n1793 171.744
R18076 vdd.n1673 vdd.n1672 171.744
R18077 vdd.n1672 vdd.n1671 171.744
R18078 vdd.n1671 vdd.n1640 171.744
R18079 vdd.n1664 vdd.n1640 171.744
R18080 vdd.n1664 vdd.n1663 171.744
R18081 vdd.n1663 vdd.n1645 171.744
R18082 vdd.n1656 vdd.n1645 171.744
R18083 vdd.n1656 vdd.n1655 171.744
R18084 vdd.n1655 vdd.n1649 171.744
R18085 vdd.n1724 vdd.n1723 171.744
R18086 vdd.n1723 vdd.n1722 171.744
R18087 vdd.n1722 vdd.n1691 171.744
R18088 vdd.n1715 vdd.n1691 171.744
R18089 vdd.n1715 vdd.n1714 171.744
R18090 vdd.n1714 vdd.n1696 171.744
R18091 vdd.n1707 vdd.n1696 171.744
R18092 vdd.n1707 vdd.n1706 171.744
R18093 vdd.n1706 vdd.n1700 171.744
R18094 vdd.n3222 vdd.n356 146.341
R18095 vdd.n3220 vdd.n3219 146.341
R18096 vdd.n3217 vdd.n360 146.341
R18097 vdd.n3213 vdd.n3212 146.341
R18098 vdd.n3210 vdd.n368 146.341
R18099 vdd.n3206 vdd.n3205 146.341
R18100 vdd.n3203 vdd.n375 146.341
R18101 vdd.n3199 vdd.n3198 146.341
R18102 vdd.n3196 vdd.n382 146.341
R18103 vdd.n393 vdd.n390 146.341
R18104 vdd.n3188 vdd.n3187 146.341
R18105 vdd.n3185 vdd.n395 146.341
R18106 vdd.n3181 vdd.n3180 146.341
R18107 vdd.n3178 vdd.n401 146.341
R18108 vdd.n3174 vdd.n3173 146.341
R18109 vdd.n3171 vdd.n408 146.341
R18110 vdd.n3167 vdd.n3166 146.341
R18111 vdd.n3164 vdd.n415 146.341
R18112 vdd.n3160 vdd.n3159 146.341
R18113 vdd.n3157 vdd.n422 146.341
R18114 vdd.n433 vdd.n430 146.341
R18115 vdd.n3149 vdd.n3148 146.341
R18116 vdd.n3146 vdd.n435 146.341
R18117 vdd.n3142 vdd.n3141 146.341
R18118 vdd.n3139 vdd.n441 146.341
R18119 vdd.n3135 vdd.n3134 146.341
R18120 vdd.n3132 vdd.n448 146.341
R18121 vdd.n3128 vdd.n3127 146.341
R18122 vdd.n3125 vdd.n455 146.341
R18123 vdd.n3121 vdd.n3120 146.341
R18124 vdd.n3118 vdd.n462 146.341
R18125 vdd.n3033 vdd.n512 146.341
R18126 vdd.n3039 vdd.n512 146.341
R18127 vdd.n3039 vdd.n504 146.341
R18128 vdd.n3049 vdd.n504 146.341
R18129 vdd.n3049 vdd.n500 146.341
R18130 vdd.n3055 vdd.n500 146.341
R18131 vdd.n3055 vdd.n491 146.341
R18132 vdd.n3065 vdd.n491 146.341
R18133 vdd.n3065 vdd.n487 146.341
R18134 vdd.n3071 vdd.n487 146.341
R18135 vdd.n3071 vdd.n479 146.341
R18136 vdd.n3082 vdd.n479 146.341
R18137 vdd.n3082 vdd.n480 146.341
R18138 vdd.n480 vdd.n316 146.341
R18139 vdd.n317 vdd.n316 146.341
R18140 vdd.n318 vdd.n317 146.341
R18141 vdd.n473 vdd.n318 146.341
R18142 vdd.n473 vdd.n326 146.341
R18143 vdd.n327 vdd.n326 146.341
R18144 vdd.n328 vdd.n327 146.341
R18145 vdd.n470 vdd.n328 146.341
R18146 vdd.n470 vdd.n337 146.341
R18147 vdd.n338 vdd.n337 146.341
R18148 vdd.n339 vdd.n338 146.341
R18149 vdd.n467 vdd.n339 146.341
R18150 vdd.n467 vdd.n348 146.341
R18151 vdd.n349 vdd.n348 146.341
R18152 vdd.n350 vdd.n349 146.341
R18153 vdd.n3025 vdd.n3023 146.341
R18154 vdd.n3023 vdd.n3022 146.341
R18155 vdd.n3019 vdd.n3018 146.341
R18156 vdd.n3015 vdd.n3014 146.341
R18157 vdd.n3012 vdd.n526 146.341
R18158 vdd.n3008 vdd.n3006 146.341
R18159 vdd.n3004 vdd.n532 146.341
R18160 vdd.n3000 vdd.n2998 146.341
R18161 vdd.n2996 vdd.n538 146.341
R18162 vdd.n2992 vdd.n2990 146.341
R18163 vdd.n2988 vdd.n546 146.341
R18164 vdd.n2984 vdd.n2982 146.341
R18165 vdd.n2980 vdd.n552 146.341
R18166 vdd.n2976 vdd.n2974 146.341
R18167 vdd.n2972 vdd.n558 146.341
R18168 vdd.n2968 vdd.n2966 146.341
R18169 vdd.n2964 vdd.n564 146.341
R18170 vdd.n2960 vdd.n2958 146.341
R18171 vdd.n2956 vdd.n570 146.341
R18172 vdd.n2952 vdd.n2950 146.341
R18173 vdd.n2948 vdd.n576 146.341
R18174 vdd.n2941 vdd.n585 146.341
R18175 vdd.n2939 vdd.n2938 146.341
R18176 vdd.n2935 vdd.n2934 146.341
R18177 vdd.n2932 vdd.n590 146.341
R18178 vdd.n2928 vdd.n2926 146.341
R18179 vdd.n2924 vdd.n596 146.341
R18180 vdd.n2920 vdd.n2918 146.341
R18181 vdd.n2916 vdd.n602 146.341
R18182 vdd.n2912 vdd.n2910 146.341
R18183 vdd.n2907 vdd.n2906 146.341
R18184 vdd.n2903 vdd.n515 146.341
R18185 vdd.n3031 vdd.n510 146.341
R18186 vdd.n3041 vdd.n510 146.341
R18187 vdd.n3041 vdd.n506 146.341
R18188 vdd.n3047 vdd.n506 146.341
R18189 vdd.n3047 vdd.n498 146.341
R18190 vdd.n3057 vdd.n498 146.341
R18191 vdd.n3057 vdd.n494 146.341
R18192 vdd.n3063 vdd.n494 146.341
R18193 vdd.n3063 vdd.n486 146.341
R18194 vdd.n3074 vdd.n486 146.341
R18195 vdd.n3074 vdd.n482 146.341
R18196 vdd.n3080 vdd.n482 146.341
R18197 vdd.n3080 vdd.n314 146.341
R18198 vdd.n3257 vdd.n314 146.341
R18199 vdd.n3257 vdd.n315 146.341
R18200 vdd.n3253 vdd.n315 146.341
R18201 vdd.n3253 vdd.n319 146.341
R18202 vdd.n3249 vdd.n319 146.341
R18203 vdd.n3249 vdd.n324 146.341
R18204 vdd.n3245 vdd.n324 146.341
R18205 vdd.n3245 vdd.n330 146.341
R18206 vdd.n3241 vdd.n330 146.341
R18207 vdd.n3241 vdd.n336 146.341
R18208 vdd.n3237 vdd.n336 146.341
R18209 vdd.n3237 vdd.n341 146.341
R18210 vdd.n3233 vdd.n341 146.341
R18211 vdd.n3233 vdd.n347 146.341
R18212 vdd.n3229 vdd.n347 146.341
R18213 vdd.n2090 vdd.n2089 146.341
R18214 vdd.n2087 vdd.n2084 146.341
R18215 vdd.n2082 vdd.n955 146.341
R18216 vdd.n2078 vdd.n2077 146.341
R18217 vdd.n2075 vdd.n959 146.341
R18218 vdd.n2071 vdd.n2070 146.341
R18219 vdd.n2068 vdd.n966 146.341
R18220 vdd.n2064 vdd.n2063 146.341
R18221 vdd.n2061 vdd.n973 146.341
R18222 vdd.n984 vdd.n981 146.341
R18223 vdd.n2053 vdd.n2052 146.341
R18224 vdd.n2050 vdd.n986 146.341
R18225 vdd.n2046 vdd.n2045 146.341
R18226 vdd.n2043 vdd.n992 146.341
R18227 vdd.n2039 vdd.n2038 146.341
R18228 vdd.n2036 vdd.n999 146.341
R18229 vdd.n2032 vdd.n2031 146.341
R18230 vdd.n2029 vdd.n1006 146.341
R18231 vdd.n2025 vdd.n2024 146.341
R18232 vdd.n2022 vdd.n1013 146.341
R18233 vdd.n1024 vdd.n1021 146.341
R18234 vdd.n2014 vdd.n2013 146.341
R18235 vdd.n2011 vdd.n1026 146.341
R18236 vdd.n2007 vdd.n2006 146.341
R18237 vdd.n2004 vdd.n1032 146.341
R18238 vdd.n2000 vdd.n1999 146.341
R18239 vdd.n1997 vdd.n1039 146.341
R18240 vdd.n1993 vdd.n1992 146.341
R18241 vdd.n1990 vdd.n1046 146.341
R18242 vdd.n1257 vdd.n1255 146.341
R18243 vdd.n1260 vdd.n1259 146.341
R18244 vdd.n1578 vdd.n1340 146.341
R18245 vdd.n1584 vdd.n1340 146.341
R18246 vdd.n1584 vdd.n1333 146.341
R18247 vdd.n1594 vdd.n1333 146.341
R18248 vdd.n1594 vdd.n1329 146.341
R18249 vdd.n1600 vdd.n1329 146.341
R18250 vdd.n1600 vdd.n1320 146.341
R18251 vdd.n1610 vdd.n1320 146.341
R18252 vdd.n1610 vdd.n1316 146.341
R18253 vdd.n1616 vdd.n1316 146.341
R18254 vdd.n1616 vdd.n1309 146.341
R18255 vdd.n1627 vdd.n1309 146.341
R18256 vdd.n1627 vdd.n1305 146.341
R18257 vdd.n1633 vdd.n1305 146.341
R18258 vdd.n1633 vdd.n1298 146.341
R18259 vdd.n1925 vdd.n1298 146.341
R18260 vdd.n1925 vdd.n1294 146.341
R18261 vdd.n1931 vdd.n1294 146.341
R18262 vdd.n1931 vdd.n1286 146.341
R18263 vdd.n1942 vdd.n1286 146.341
R18264 vdd.n1942 vdd.n1282 146.341
R18265 vdd.n1948 vdd.n1282 146.341
R18266 vdd.n1948 vdd.n1276 146.341
R18267 vdd.n1959 vdd.n1276 146.341
R18268 vdd.n1959 vdd.n1271 146.341
R18269 vdd.n1967 vdd.n1271 146.341
R18270 vdd.n1967 vdd.n1262 146.341
R18271 vdd.n1978 vdd.n1262 146.341
R18272 vdd.n1350 vdd.n1349 146.341
R18273 vdd.n1353 vdd.n1350 146.341
R18274 vdd.n1356 vdd.n1355 146.341
R18275 vdd.n1361 vdd.n1358 146.341
R18276 vdd.n1364 vdd.n1363 146.341
R18277 vdd.n1369 vdd.n1366 146.341
R18278 vdd.n1372 vdd.n1371 146.341
R18279 vdd.n1377 vdd.n1374 146.341
R18280 vdd.n1380 vdd.n1379 146.341
R18281 vdd.n1387 vdd.n1382 146.341
R18282 vdd.n1390 vdd.n1389 146.341
R18283 vdd.n1395 vdd.n1392 146.341
R18284 vdd.n1398 vdd.n1397 146.341
R18285 vdd.n1403 vdd.n1400 146.341
R18286 vdd.n1406 vdd.n1405 146.341
R18287 vdd.n1411 vdd.n1408 146.341
R18288 vdd.n1414 vdd.n1413 146.341
R18289 vdd.n1419 vdd.n1416 146.341
R18290 vdd.n1422 vdd.n1421 146.341
R18291 vdd.n1427 vdd.n1424 146.341
R18292 vdd.n1508 vdd.n1429 146.341
R18293 vdd.n1506 vdd.n1505 146.341
R18294 vdd.n1436 vdd.n1435 146.341
R18295 vdd.n1439 vdd.n1438 146.341
R18296 vdd.n1444 vdd.n1443 146.341
R18297 vdd.n1447 vdd.n1446 146.341
R18298 vdd.n1452 vdd.n1451 146.341
R18299 vdd.n1455 vdd.n1454 146.341
R18300 vdd.n1460 vdd.n1459 146.341
R18301 vdd.n1463 vdd.n1462 146.341
R18302 vdd.n1468 vdd.n1467 146.341
R18303 vdd.n1470 vdd.n1343 146.341
R18304 vdd.n1576 vdd.n1339 146.341
R18305 vdd.n1586 vdd.n1339 146.341
R18306 vdd.n1586 vdd.n1335 146.341
R18307 vdd.n1592 vdd.n1335 146.341
R18308 vdd.n1592 vdd.n1327 146.341
R18309 vdd.n1602 vdd.n1327 146.341
R18310 vdd.n1602 vdd.n1323 146.341
R18311 vdd.n1608 vdd.n1323 146.341
R18312 vdd.n1608 vdd.n1315 146.341
R18313 vdd.n1619 vdd.n1315 146.341
R18314 vdd.n1619 vdd.n1311 146.341
R18315 vdd.n1625 vdd.n1311 146.341
R18316 vdd.n1625 vdd.n1304 146.341
R18317 vdd.n1635 vdd.n1304 146.341
R18318 vdd.n1635 vdd.n1300 146.341
R18319 vdd.n1923 vdd.n1300 146.341
R18320 vdd.n1923 vdd.n1292 146.341
R18321 vdd.n1934 vdd.n1292 146.341
R18322 vdd.n1934 vdd.n1288 146.341
R18323 vdd.n1940 vdd.n1288 146.341
R18324 vdd.n1940 vdd.n1281 146.341
R18325 vdd.n1951 vdd.n1281 146.341
R18326 vdd.n1951 vdd.n1277 146.341
R18327 vdd.n1957 vdd.n1277 146.341
R18328 vdd.n1957 vdd.n1269 146.341
R18329 vdd.n1970 vdd.n1269 146.341
R18330 vdd.n1970 vdd.n1264 146.341
R18331 vdd.n1976 vdd.n1264 146.341
R18332 vdd.n1081 vdd.t11 127.284
R18333 vdd.n809 vdd.t52 127.284
R18334 vdd.n1101 vdd.t36 127.284
R18335 vdd.n800 vdd.t69 127.284
R18336 vdd.n700 vdd.t39 127.284
R18337 vdd.n700 vdd.t40 127.284
R18338 vdd.n2416 vdd.t67 127.284
R18339 vdd.n661 vdd.t75 127.284
R18340 vdd.n2413 vdd.t57 127.284
R18341 vdd.n625 vdd.t6 127.284
R18342 vdd.n871 vdd.t60 127.284
R18343 vdd.n871 vdd.t61 127.284
R18344 vdd.n22 vdd.n20 117.314
R18345 vdd.n17 vdd.n15 117.314
R18346 vdd.n27 vdd.n26 116.927
R18347 vdd.n24 vdd.n23 116.927
R18348 vdd.n22 vdd.n21 116.927
R18349 vdd.n17 vdd.n16 116.927
R18350 vdd.n19 vdd.n18 116.927
R18351 vdd.n27 vdd.n25 116.927
R18352 vdd.n1082 vdd.t10 111.188
R18353 vdd.n810 vdd.t53 111.188
R18354 vdd.n1102 vdd.t35 111.188
R18355 vdd.n801 vdd.t70 111.188
R18356 vdd.n2417 vdd.t66 111.188
R18357 vdd.n662 vdd.t76 111.188
R18358 vdd.n2414 vdd.t56 111.188
R18359 vdd.n626 vdd.t7 111.188
R18360 vdd.n2658 vdd.n755 99.5127
R18361 vdd.n2658 vdd.n753 99.5127
R18362 vdd.n2662 vdd.n753 99.5127
R18363 vdd.n2662 vdd.n744 99.5127
R18364 vdd.n2670 vdd.n744 99.5127
R18365 vdd.n2670 vdd.n742 99.5127
R18366 vdd.n2674 vdd.n742 99.5127
R18367 vdd.n2674 vdd.n732 99.5127
R18368 vdd.n2682 vdd.n732 99.5127
R18369 vdd.n2682 vdd.n730 99.5127
R18370 vdd.n2686 vdd.n730 99.5127
R18371 vdd.n2686 vdd.n720 99.5127
R18372 vdd.n2694 vdd.n720 99.5127
R18373 vdd.n2694 vdd.n718 99.5127
R18374 vdd.n2698 vdd.n718 99.5127
R18375 vdd.n2698 vdd.n709 99.5127
R18376 vdd.n2706 vdd.n709 99.5127
R18377 vdd.n2706 vdd.n707 99.5127
R18378 vdd.n2710 vdd.n707 99.5127
R18379 vdd.n2710 vdd.n695 99.5127
R18380 vdd.n2719 vdd.n695 99.5127
R18381 vdd.n2719 vdd.n693 99.5127
R18382 vdd.n2723 vdd.n693 99.5127
R18383 vdd.n2723 vdd.n684 99.5127
R18384 vdd.n2731 vdd.n684 99.5127
R18385 vdd.n2731 vdd.n682 99.5127
R18386 vdd.n2735 vdd.n682 99.5127
R18387 vdd.n2735 vdd.n670 99.5127
R18388 vdd.n2788 vdd.n670 99.5127
R18389 vdd.n2788 vdd.n668 99.5127
R18390 vdd.n2792 vdd.n668 99.5127
R18391 vdd.n2792 vdd.n634 99.5127
R18392 vdd.n2862 vdd.n634 99.5127
R18393 vdd.n2858 vdd.n635 99.5127
R18394 vdd.n2856 vdd.n2855 99.5127
R18395 vdd.n2853 vdd.n639 99.5127
R18396 vdd.n2849 vdd.n2848 99.5127
R18397 vdd.n2846 vdd.n642 99.5127
R18398 vdd.n2842 vdd.n2841 99.5127
R18399 vdd.n2839 vdd.n645 99.5127
R18400 vdd.n2835 vdd.n2834 99.5127
R18401 vdd.n2832 vdd.n648 99.5127
R18402 vdd.n2827 vdd.n2826 99.5127
R18403 vdd.n2824 vdd.n651 99.5127
R18404 vdd.n2820 vdd.n2819 99.5127
R18405 vdd.n2817 vdd.n654 99.5127
R18406 vdd.n2813 vdd.n2812 99.5127
R18407 vdd.n2810 vdd.n657 99.5127
R18408 vdd.n2806 vdd.n2805 99.5127
R18409 vdd.n2803 vdd.n660 99.5127
R18410 vdd.n2579 vdd.n757 99.5127
R18411 vdd.n2575 vdd.n757 99.5127
R18412 vdd.n2575 vdd.n751 99.5127
R18413 vdd.n2519 vdd.n751 99.5127
R18414 vdd.n2519 vdd.n746 99.5127
R18415 vdd.n2522 vdd.n746 99.5127
R18416 vdd.n2522 vdd.n740 99.5127
R18417 vdd.n2525 vdd.n740 99.5127
R18418 vdd.n2525 vdd.n734 99.5127
R18419 vdd.n2558 vdd.n734 99.5127
R18420 vdd.n2558 vdd.n727 99.5127
R18421 vdd.n2554 vdd.n727 99.5127
R18422 vdd.n2554 vdd.n721 99.5127
R18423 vdd.n2551 vdd.n721 99.5127
R18424 vdd.n2551 vdd.n716 99.5127
R18425 vdd.n2548 vdd.n716 99.5127
R18426 vdd.n2548 vdd.n711 99.5127
R18427 vdd.n2545 vdd.n711 99.5127
R18428 vdd.n2545 vdd.n704 99.5127
R18429 vdd.n2542 vdd.n704 99.5127
R18430 vdd.n2542 vdd.n696 99.5127
R18431 vdd.n2539 vdd.n696 99.5127
R18432 vdd.n2539 vdd.n691 99.5127
R18433 vdd.n2536 vdd.n691 99.5127
R18434 vdd.n2536 vdd.n686 99.5127
R18435 vdd.n2533 vdd.n686 99.5127
R18436 vdd.n2533 vdd.n680 99.5127
R18437 vdd.n2530 vdd.n680 99.5127
R18438 vdd.n2530 vdd.n672 99.5127
R18439 vdd.n672 vdd.n665 99.5127
R18440 vdd.n2794 vdd.n665 99.5127
R18441 vdd.n2795 vdd.n2794 99.5127
R18442 vdd.n2795 vdd.n632 99.5127
R18443 vdd.n2412 vdd.n2411 99.5127
R18444 vdd.n2643 vdd.n2411 99.5127
R18445 vdd.n2641 vdd.n2640 99.5127
R18446 vdd.n2637 vdd.n2636 99.5127
R18447 vdd.n2633 vdd.n2632 99.5127
R18448 vdd.n2629 vdd.n2628 99.5127
R18449 vdd.n2625 vdd.n2624 99.5127
R18450 vdd.n2621 vdd.n2620 99.5127
R18451 vdd.n2617 vdd.n2616 99.5127
R18452 vdd.n2613 vdd.n2612 99.5127
R18453 vdd.n2609 vdd.n2608 99.5127
R18454 vdd.n2605 vdd.n2604 99.5127
R18455 vdd.n2601 vdd.n2600 99.5127
R18456 vdd.n2597 vdd.n2596 99.5127
R18457 vdd.n2593 vdd.n2592 99.5127
R18458 vdd.n2589 vdd.n2588 99.5127
R18459 vdd.n2584 vdd.n2583 99.5127
R18460 vdd.n2376 vdd.n798 99.5127
R18461 vdd.n2372 vdd.n2371 99.5127
R18462 vdd.n2368 vdd.n2367 99.5127
R18463 vdd.n2364 vdd.n2363 99.5127
R18464 vdd.n2360 vdd.n2359 99.5127
R18465 vdd.n2356 vdd.n2355 99.5127
R18466 vdd.n2352 vdd.n2351 99.5127
R18467 vdd.n2348 vdd.n2347 99.5127
R18468 vdd.n2344 vdd.n2343 99.5127
R18469 vdd.n2340 vdd.n2339 99.5127
R18470 vdd.n2336 vdd.n2335 99.5127
R18471 vdd.n2332 vdd.n2331 99.5127
R18472 vdd.n2328 vdd.n2327 99.5127
R18473 vdd.n2324 vdd.n2323 99.5127
R18474 vdd.n2320 vdd.n2319 99.5127
R18475 vdd.n2316 vdd.n2315 99.5127
R18476 vdd.n2311 vdd.n2310 99.5127
R18477 vdd.n1137 vdd.n905 99.5127
R18478 vdd.n1140 vdd.n905 99.5127
R18479 vdd.n1140 vdd.n899 99.5127
R18480 vdd.n1143 vdd.n899 99.5127
R18481 vdd.n1143 vdd.n894 99.5127
R18482 vdd.n1146 vdd.n894 99.5127
R18483 vdd.n1146 vdd.n888 99.5127
R18484 vdd.n1149 vdd.n888 99.5127
R18485 vdd.n1149 vdd.n881 99.5127
R18486 vdd.n1152 vdd.n881 99.5127
R18487 vdd.n1152 vdd.n874 99.5127
R18488 vdd.n1155 vdd.n874 99.5127
R18489 vdd.n1155 vdd.n868 99.5127
R18490 vdd.n1158 vdd.n868 99.5127
R18491 vdd.n1158 vdd.n863 99.5127
R18492 vdd.n1161 vdd.n863 99.5127
R18493 vdd.n1161 vdd.n857 99.5127
R18494 vdd.n1186 vdd.n857 99.5127
R18495 vdd.n1186 vdd.n850 99.5127
R18496 vdd.n1182 vdd.n850 99.5127
R18497 vdd.n1182 vdd.n844 99.5127
R18498 vdd.n1179 vdd.n844 99.5127
R18499 vdd.n1179 vdd.n839 99.5127
R18500 vdd.n1176 vdd.n839 99.5127
R18501 vdd.n1176 vdd.n834 99.5127
R18502 vdd.n1173 vdd.n834 99.5127
R18503 vdd.n1173 vdd.n828 99.5127
R18504 vdd.n1170 vdd.n828 99.5127
R18505 vdd.n1170 vdd.n821 99.5127
R18506 vdd.n1167 vdd.n821 99.5127
R18507 vdd.n1167 vdd.n814 99.5127
R18508 vdd.n814 vdd.n803 99.5127
R18509 vdd.n2306 vdd.n803 99.5127
R18510 vdd.n946 vdd.n945 99.5127
R18511 vdd.n2122 vdd.n945 99.5127
R18512 vdd.n2120 vdd.n2119 99.5127
R18513 vdd.n2116 vdd.n2115 99.5127
R18514 vdd.n2112 vdd.n2111 99.5127
R18515 vdd.n2108 vdd.n2107 99.5127
R18516 vdd.n2104 vdd.n2103 99.5127
R18517 vdd.n2100 vdd.n2099 99.5127
R18518 vdd.n2096 vdd.n2095 99.5127
R18519 vdd.n1104 vdd.n1103 99.5127
R18520 vdd.n1108 vdd.n1107 99.5127
R18521 vdd.n1112 vdd.n1111 99.5127
R18522 vdd.n1116 vdd.n1115 99.5127
R18523 vdd.n1120 vdd.n1119 99.5127
R18524 vdd.n1124 vdd.n1123 99.5127
R18525 vdd.n1128 vdd.n1127 99.5127
R18526 vdd.n1133 vdd.n1132 99.5127
R18527 vdd.n2137 vdd.n903 99.5127
R18528 vdd.n2137 vdd.n901 99.5127
R18529 vdd.n2141 vdd.n901 99.5127
R18530 vdd.n2141 vdd.n892 99.5127
R18531 vdd.n2149 vdd.n892 99.5127
R18532 vdd.n2149 vdd.n890 99.5127
R18533 vdd.n2153 vdd.n890 99.5127
R18534 vdd.n2153 vdd.n879 99.5127
R18535 vdd.n2161 vdd.n879 99.5127
R18536 vdd.n2161 vdd.n877 99.5127
R18537 vdd.n2165 vdd.n877 99.5127
R18538 vdd.n2165 vdd.n867 99.5127
R18539 vdd.n2174 vdd.n867 99.5127
R18540 vdd.n2174 vdd.n865 99.5127
R18541 vdd.n2178 vdd.n865 99.5127
R18542 vdd.n2178 vdd.n855 99.5127
R18543 vdd.n2186 vdd.n855 99.5127
R18544 vdd.n2186 vdd.n853 99.5127
R18545 vdd.n2190 vdd.n853 99.5127
R18546 vdd.n2190 vdd.n843 99.5127
R18547 vdd.n2198 vdd.n843 99.5127
R18548 vdd.n2198 vdd.n841 99.5127
R18549 vdd.n2202 vdd.n841 99.5127
R18550 vdd.n2202 vdd.n832 99.5127
R18551 vdd.n2210 vdd.n832 99.5127
R18552 vdd.n2210 vdd.n830 99.5127
R18553 vdd.n2214 vdd.n830 99.5127
R18554 vdd.n2214 vdd.n819 99.5127
R18555 vdd.n2224 vdd.n819 99.5127
R18556 vdd.n2224 vdd.n816 99.5127
R18557 vdd.n2229 vdd.n816 99.5127
R18558 vdd.n2229 vdd.n817 99.5127
R18559 vdd.n817 vdd.n797 99.5127
R18560 vdd.n2778 vdd.n2777 99.5127
R18561 vdd.n2775 vdd.n2741 99.5127
R18562 vdd.n2771 vdd.n2770 99.5127
R18563 vdd.n2768 vdd.n2744 99.5127
R18564 vdd.n2764 vdd.n2763 99.5127
R18565 vdd.n2761 vdd.n2747 99.5127
R18566 vdd.n2757 vdd.n2756 99.5127
R18567 vdd.n2754 vdd.n2751 99.5127
R18568 vdd.n2895 vdd.n612 99.5127
R18569 vdd.n2893 vdd.n2892 99.5127
R18570 vdd.n2890 vdd.n615 99.5127
R18571 vdd.n2886 vdd.n2885 99.5127
R18572 vdd.n2883 vdd.n618 99.5127
R18573 vdd.n2879 vdd.n2878 99.5127
R18574 vdd.n2876 vdd.n621 99.5127
R18575 vdd.n2872 vdd.n2871 99.5127
R18576 vdd.n2869 vdd.n624 99.5127
R18577 vdd.n2484 vdd.n758 99.5127
R18578 vdd.n2573 vdd.n758 99.5127
R18579 vdd.n2573 vdd.n752 99.5127
R18580 vdd.n2569 vdd.n752 99.5127
R18581 vdd.n2569 vdd.n747 99.5127
R18582 vdd.n2566 vdd.n747 99.5127
R18583 vdd.n2566 vdd.n741 99.5127
R18584 vdd.n2563 vdd.n741 99.5127
R18585 vdd.n2563 vdd.n735 99.5127
R18586 vdd.n2560 vdd.n735 99.5127
R18587 vdd.n2560 vdd.n728 99.5127
R18588 vdd.n2516 vdd.n728 99.5127
R18589 vdd.n2516 vdd.n722 99.5127
R18590 vdd.n2513 vdd.n722 99.5127
R18591 vdd.n2513 vdd.n717 99.5127
R18592 vdd.n2510 vdd.n717 99.5127
R18593 vdd.n2510 vdd.n712 99.5127
R18594 vdd.n2507 vdd.n712 99.5127
R18595 vdd.n2507 vdd.n705 99.5127
R18596 vdd.n2504 vdd.n705 99.5127
R18597 vdd.n2504 vdd.n697 99.5127
R18598 vdd.n2501 vdd.n697 99.5127
R18599 vdd.n2501 vdd.n692 99.5127
R18600 vdd.n2498 vdd.n692 99.5127
R18601 vdd.n2498 vdd.n687 99.5127
R18602 vdd.n2495 vdd.n687 99.5127
R18603 vdd.n2495 vdd.n681 99.5127
R18604 vdd.n2492 vdd.n681 99.5127
R18605 vdd.n2492 vdd.n673 99.5127
R18606 vdd.n2489 vdd.n673 99.5127
R18607 vdd.n2489 vdd.n666 99.5127
R18608 vdd.n666 vdd.n630 99.5127
R18609 vdd.n2864 vdd.n630 99.5127
R18610 vdd.n2419 vdd.n761 99.5127
R18611 vdd.n2423 vdd.n2422 99.5127
R18612 vdd.n2427 vdd.n2426 99.5127
R18613 vdd.n2431 vdd.n2430 99.5127
R18614 vdd.n2435 vdd.n2434 99.5127
R18615 vdd.n2439 vdd.n2438 99.5127
R18616 vdd.n2443 vdd.n2442 99.5127
R18617 vdd.n2447 vdd.n2446 99.5127
R18618 vdd.n2451 vdd.n2450 99.5127
R18619 vdd.n2455 vdd.n2454 99.5127
R18620 vdd.n2459 vdd.n2458 99.5127
R18621 vdd.n2463 vdd.n2462 99.5127
R18622 vdd.n2467 vdd.n2466 99.5127
R18623 vdd.n2471 vdd.n2470 99.5127
R18624 vdd.n2475 vdd.n2474 99.5127
R18625 vdd.n2479 vdd.n2478 99.5127
R18626 vdd.n2481 vdd.n2410 99.5127
R18627 vdd.n2656 vdd.n759 99.5127
R18628 vdd.n2656 vdd.n750 99.5127
R18629 vdd.n2664 vdd.n750 99.5127
R18630 vdd.n2664 vdd.n748 99.5127
R18631 vdd.n2668 vdd.n748 99.5127
R18632 vdd.n2668 vdd.n738 99.5127
R18633 vdd.n2676 vdd.n738 99.5127
R18634 vdd.n2676 vdd.n736 99.5127
R18635 vdd.n2680 vdd.n736 99.5127
R18636 vdd.n2680 vdd.n726 99.5127
R18637 vdd.n2688 vdd.n726 99.5127
R18638 vdd.n2688 vdd.n724 99.5127
R18639 vdd.n2692 vdd.n724 99.5127
R18640 vdd.n2692 vdd.n715 99.5127
R18641 vdd.n2700 vdd.n715 99.5127
R18642 vdd.n2700 vdd.n713 99.5127
R18643 vdd.n2704 vdd.n713 99.5127
R18644 vdd.n2704 vdd.n702 99.5127
R18645 vdd.n2712 vdd.n702 99.5127
R18646 vdd.n2712 vdd.n699 99.5127
R18647 vdd.n2717 vdd.n699 99.5127
R18648 vdd.n2717 vdd.n690 99.5127
R18649 vdd.n2725 vdd.n690 99.5127
R18650 vdd.n2725 vdd.n688 99.5127
R18651 vdd.n2729 vdd.n688 99.5127
R18652 vdd.n2729 vdd.n678 99.5127
R18653 vdd.n2737 vdd.n678 99.5127
R18654 vdd.n2737 vdd.n675 99.5127
R18655 vdd.n2786 vdd.n675 99.5127
R18656 vdd.n2786 vdd.n676 99.5127
R18657 vdd.n676 vdd.n667 99.5127
R18658 vdd.n2781 vdd.n667 99.5127
R18659 vdd.n2781 vdd.n633 99.5127
R18660 vdd.n2300 vdd.n2299 99.5127
R18661 vdd.n2296 vdd.n2295 99.5127
R18662 vdd.n2292 vdd.n2291 99.5127
R18663 vdd.n2288 vdd.n2287 99.5127
R18664 vdd.n2284 vdd.n2283 99.5127
R18665 vdd.n2280 vdd.n2279 99.5127
R18666 vdd.n2276 vdd.n2275 99.5127
R18667 vdd.n2272 vdd.n2271 99.5127
R18668 vdd.n2268 vdd.n2267 99.5127
R18669 vdd.n2264 vdd.n2263 99.5127
R18670 vdd.n2260 vdd.n2259 99.5127
R18671 vdd.n2256 vdd.n2255 99.5127
R18672 vdd.n2252 vdd.n2251 99.5127
R18673 vdd.n2248 vdd.n2247 99.5127
R18674 vdd.n2244 vdd.n2243 99.5127
R18675 vdd.n2240 vdd.n2239 99.5127
R18676 vdd.n2236 vdd.n779 99.5127
R18677 vdd.n1215 vdd.n906 99.5127
R18678 vdd.n1212 vdd.n906 99.5127
R18679 vdd.n1212 vdd.n900 99.5127
R18680 vdd.n1209 vdd.n900 99.5127
R18681 vdd.n1209 vdd.n895 99.5127
R18682 vdd.n1206 vdd.n895 99.5127
R18683 vdd.n1206 vdd.n889 99.5127
R18684 vdd.n1203 vdd.n889 99.5127
R18685 vdd.n1203 vdd.n882 99.5127
R18686 vdd.n1200 vdd.n882 99.5127
R18687 vdd.n1200 vdd.n875 99.5127
R18688 vdd.n1197 vdd.n875 99.5127
R18689 vdd.n1197 vdd.n869 99.5127
R18690 vdd.n1194 vdd.n869 99.5127
R18691 vdd.n1194 vdd.n864 99.5127
R18692 vdd.n1191 vdd.n864 99.5127
R18693 vdd.n1191 vdd.n858 99.5127
R18694 vdd.n1188 vdd.n858 99.5127
R18695 vdd.n1188 vdd.n851 99.5127
R18696 vdd.n1098 vdd.n851 99.5127
R18697 vdd.n1098 vdd.n845 99.5127
R18698 vdd.n1095 vdd.n845 99.5127
R18699 vdd.n1095 vdd.n840 99.5127
R18700 vdd.n1092 vdd.n840 99.5127
R18701 vdd.n1092 vdd.n835 99.5127
R18702 vdd.n1089 vdd.n835 99.5127
R18703 vdd.n1089 vdd.n829 99.5127
R18704 vdd.n1086 vdd.n829 99.5127
R18705 vdd.n1086 vdd.n822 99.5127
R18706 vdd.n822 vdd.n813 99.5127
R18707 vdd.n2231 vdd.n813 99.5127
R18708 vdd.n2232 vdd.n2231 99.5127
R18709 vdd.n2232 vdd.n805 99.5127
R18710 vdd.n1050 vdd.n910 99.5127
R18711 vdd.n1054 vdd.n1053 99.5127
R18712 vdd.n1058 vdd.n1057 99.5127
R18713 vdd.n1062 vdd.n1061 99.5127
R18714 vdd.n1066 vdd.n1065 99.5127
R18715 vdd.n1070 vdd.n1069 99.5127
R18716 vdd.n1074 vdd.n1073 99.5127
R18717 vdd.n1078 vdd.n1077 99.5127
R18718 vdd.n1248 vdd.n1080 99.5127
R18719 vdd.n1246 vdd.n1245 99.5127
R18720 vdd.n1242 vdd.n1241 99.5127
R18721 vdd.n1238 vdd.n1237 99.5127
R18722 vdd.n1234 vdd.n1233 99.5127
R18723 vdd.n1230 vdd.n1229 99.5127
R18724 vdd.n1226 vdd.n1225 99.5127
R18725 vdd.n1222 vdd.n1221 99.5127
R18726 vdd.n1218 vdd.n944 99.5127
R18727 vdd.n2135 vdd.n908 99.5127
R18728 vdd.n2135 vdd.n898 99.5127
R18729 vdd.n2143 vdd.n898 99.5127
R18730 vdd.n2143 vdd.n896 99.5127
R18731 vdd.n2147 vdd.n896 99.5127
R18732 vdd.n2147 vdd.n886 99.5127
R18733 vdd.n2155 vdd.n886 99.5127
R18734 vdd.n2155 vdd.n884 99.5127
R18735 vdd.n2159 vdd.n884 99.5127
R18736 vdd.n2159 vdd.n873 99.5127
R18737 vdd.n2167 vdd.n873 99.5127
R18738 vdd.n2167 vdd.n870 99.5127
R18739 vdd.n2172 vdd.n870 99.5127
R18740 vdd.n2172 vdd.n861 99.5127
R18741 vdd.n2180 vdd.n861 99.5127
R18742 vdd.n2180 vdd.n859 99.5127
R18743 vdd.n2184 vdd.n859 99.5127
R18744 vdd.n2184 vdd.n849 99.5127
R18745 vdd.n2192 vdd.n849 99.5127
R18746 vdd.n2192 vdd.n847 99.5127
R18747 vdd.n2196 vdd.n847 99.5127
R18748 vdd.n2196 vdd.n838 99.5127
R18749 vdd.n2204 vdd.n838 99.5127
R18750 vdd.n2204 vdd.n836 99.5127
R18751 vdd.n2208 vdd.n836 99.5127
R18752 vdd.n2208 vdd.n826 99.5127
R18753 vdd.n2216 vdd.n826 99.5127
R18754 vdd.n2216 vdd.n823 99.5127
R18755 vdd.n2222 vdd.n823 99.5127
R18756 vdd.n2222 vdd.n824 99.5127
R18757 vdd.n824 vdd.n815 99.5127
R18758 vdd.n815 vdd.n806 99.5127
R18759 vdd.n2304 vdd.n806 99.5127
R18760 vdd.n9 vdd.n7 98.9633
R18761 vdd.n2 vdd.n0 98.9633
R18762 vdd.n9 vdd.n8 98.6055
R18763 vdd.n11 vdd.n10 98.6055
R18764 vdd.n13 vdd.n12 98.6055
R18765 vdd.n6 vdd.n5 98.6055
R18766 vdd.n4 vdd.n3 98.6055
R18767 vdd.n2 vdd.n1 98.6055
R18768 vdd.t215 vdd.n279 85.8723
R18769 vdd.t197 vdd.n228 85.8723
R18770 vdd.t206 vdd.n185 85.8723
R18771 vdd.t186 vdd.n134 85.8723
R18772 vdd.t152 vdd.n92 85.8723
R18773 vdd.t160 vdd.n41 85.8723
R18774 vdd.t221 vdd.n1836 85.8723
R18775 vdd.t155 vdd.n1887 85.8723
R18776 vdd.t212 vdd.n1742 85.8723
R18777 vdd.t141 vdd.n1793 85.8723
R18778 vdd.t162 vdd.n1649 85.8723
R18779 vdd.t153 vdd.n1700 85.8723
R18780 vdd.n2715 vdd.n700 78.546
R18781 vdd.n2170 vdd.n871 78.546
R18782 vdd.n266 vdd.n265 75.1835
R18783 vdd.n264 vdd.n263 75.1835
R18784 vdd.n262 vdd.n261 75.1835
R18785 vdd.n260 vdd.n259 75.1835
R18786 vdd.n258 vdd.n257 75.1835
R18787 vdd.n172 vdd.n171 75.1835
R18788 vdd.n170 vdd.n169 75.1835
R18789 vdd.n168 vdd.n167 75.1835
R18790 vdd.n166 vdd.n165 75.1835
R18791 vdd.n164 vdd.n163 75.1835
R18792 vdd.n79 vdd.n78 75.1835
R18793 vdd.n77 vdd.n76 75.1835
R18794 vdd.n75 vdd.n74 75.1835
R18795 vdd.n73 vdd.n72 75.1835
R18796 vdd.n71 vdd.n70 75.1835
R18797 vdd.n1866 vdd.n1865 75.1835
R18798 vdd.n1868 vdd.n1867 75.1835
R18799 vdd.n1870 vdd.n1869 75.1835
R18800 vdd.n1872 vdd.n1871 75.1835
R18801 vdd.n1874 vdd.n1873 75.1835
R18802 vdd.n1772 vdd.n1771 75.1835
R18803 vdd.n1774 vdd.n1773 75.1835
R18804 vdd.n1776 vdd.n1775 75.1835
R18805 vdd.n1778 vdd.n1777 75.1835
R18806 vdd.n1780 vdd.n1779 75.1835
R18807 vdd.n1679 vdd.n1678 75.1835
R18808 vdd.n1681 vdd.n1680 75.1835
R18809 vdd.n1683 vdd.n1682 75.1835
R18810 vdd.n1685 vdd.n1684 75.1835
R18811 vdd.n1687 vdd.n1686 75.1835
R18812 vdd.n2651 vdd.n2650 72.8958
R18813 vdd.n2650 vdd.n2394 72.8958
R18814 vdd.n2650 vdd.n2395 72.8958
R18815 vdd.n2650 vdd.n2396 72.8958
R18816 vdd.n2650 vdd.n2397 72.8958
R18817 vdd.n2650 vdd.n2398 72.8958
R18818 vdd.n2650 vdd.n2399 72.8958
R18819 vdd.n2650 vdd.n2400 72.8958
R18820 vdd.n2650 vdd.n2401 72.8958
R18821 vdd.n2650 vdd.n2402 72.8958
R18822 vdd.n2650 vdd.n2403 72.8958
R18823 vdd.n2650 vdd.n2404 72.8958
R18824 vdd.n2650 vdd.n2405 72.8958
R18825 vdd.n2650 vdd.n2406 72.8958
R18826 vdd.n2650 vdd.n2407 72.8958
R18827 vdd.n2650 vdd.n2408 72.8958
R18828 vdd.n2650 vdd.n2409 72.8958
R18829 vdd.n629 vdd.n613 72.8958
R18830 vdd.n2870 vdd.n613 72.8958
R18831 vdd.n623 vdd.n613 72.8958
R18832 vdd.n2877 vdd.n613 72.8958
R18833 vdd.n620 vdd.n613 72.8958
R18834 vdd.n2884 vdd.n613 72.8958
R18835 vdd.n617 vdd.n613 72.8958
R18836 vdd.n2891 vdd.n613 72.8958
R18837 vdd.n2894 vdd.n613 72.8958
R18838 vdd.n2750 vdd.n613 72.8958
R18839 vdd.n2755 vdd.n613 72.8958
R18840 vdd.n2749 vdd.n613 72.8958
R18841 vdd.n2762 vdd.n613 72.8958
R18842 vdd.n2746 vdd.n613 72.8958
R18843 vdd.n2769 vdd.n613 72.8958
R18844 vdd.n2743 vdd.n613 72.8958
R18845 vdd.n2776 vdd.n613 72.8958
R18846 vdd.n2129 vdd.n2128 72.8958
R18847 vdd.n2129 vdd.n912 72.8958
R18848 vdd.n2129 vdd.n913 72.8958
R18849 vdd.n2129 vdd.n914 72.8958
R18850 vdd.n2129 vdd.n915 72.8958
R18851 vdd.n2129 vdd.n916 72.8958
R18852 vdd.n2129 vdd.n917 72.8958
R18853 vdd.n2129 vdd.n918 72.8958
R18854 vdd.n2129 vdd.n919 72.8958
R18855 vdd.n2129 vdd.n920 72.8958
R18856 vdd.n2129 vdd.n921 72.8958
R18857 vdd.n2129 vdd.n922 72.8958
R18858 vdd.n2129 vdd.n923 72.8958
R18859 vdd.n2129 vdd.n924 72.8958
R18860 vdd.n2129 vdd.n925 72.8958
R18861 vdd.n2129 vdd.n926 72.8958
R18862 vdd.n2129 vdd.n927 72.8958
R18863 vdd.n2377 vdd.n780 72.8958
R18864 vdd.n2377 vdd.n781 72.8958
R18865 vdd.n2377 vdd.n782 72.8958
R18866 vdd.n2377 vdd.n783 72.8958
R18867 vdd.n2377 vdd.n784 72.8958
R18868 vdd.n2377 vdd.n785 72.8958
R18869 vdd.n2377 vdd.n786 72.8958
R18870 vdd.n2377 vdd.n787 72.8958
R18871 vdd.n2377 vdd.n788 72.8958
R18872 vdd.n2377 vdd.n789 72.8958
R18873 vdd.n2377 vdd.n790 72.8958
R18874 vdd.n2377 vdd.n791 72.8958
R18875 vdd.n2377 vdd.n792 72.8958
R18876 vdd.n2377 vdd.n793 72.8958
R18877 vdd.n2377 vdd.n794 72.8958
R18878 vdd.n2377 vdd.n795 72.8958
R18879 vdd.n2377 vdd.n796 72.8958
R18880 vdd.n2650 vdd.n2649 72.8958
R18881 vdd.n2650 vdd.n2378 72.8958
R18882 vdd.n2650 vdd.n2379 72.8958
R18883 vdd.n2650 vdd.n2380 72.8958
R18884 vdd.n2650 vdd.n2381 72.8958
R18885 vdd.n2650 vdd.n2382 72.8958
R18886 vdd.n2650 vdd.n2383 72.8958
R18887 vdd.n2650 vdd.n2384 72.8958
R18888 vdd.n2650 vdd.n2385 72.8958
R18889 vdd.n2650 vdd.n2386 72.8958
R18890 vdd.n2650 vdd.n2387 72.8958
R18891 vdd.n2650 vdd.n2388 72.8958
R18892 vdd.n2650 vdd.n2389 72.8958
R18893 vdd.n2650 vdd.n2390 72.8958
R18894 vdd.n2650 vdd.n2391 72.8958
R18895 vdd.n2650 vdd.n2392 72.8958
R18896 vdd.n2650 vdd.n2393 72.8958
R18897 vdd.n2798 vdd.n613 72.8958
R18898 vdd.n2804 vdd.n613 72.8958
R18899 vdd.n659 vdd.n613 72.8958
R18900 vdd.n2811 vdd.n613 72.8958
R18901 vdd.n656 vdd.n613 72.8958
R18902 vdd.n2818 vdd.n613 72.8958
R18903 vdd.n653 vdd.n613 72.8958
R18904 vdd.n2825 vdd.n613 72.8958
R18905 vdd.n650 vdd.n613 72.8958
R18906 vdd.n2833 vdd.n613 72.8958
R18907 vdd.n647 vdd.n613 72.8958
R18908 vdd.n2840 vdd.n613 72.8958
R18909 vdd.n644 vdd.n613 72.8958
R18910 vdd.n2847 vdd.n613 72.8958
R18911 vdd.n641 vdd.n613 72.8958
R18912 vdd.n2854 vdd.n613 72.8958
R18913 vdd.n2857 vdd.n613 72.8958
R18914 vdd.n2377 vdd.n778 72.8958
R18915 vdd.n2377 vdd.n777 72.8958
R18916 vdd.n2377 vdd.n776 72.8958
R18917 vdd.n2377 vdd.n775 72.8958
R18918 vdd.n2377 vdd.n774 72.8958
R18919 vdd.n2377 vdd.n773 72.8958
R18920 vdd.n2377 vdd.n772 72.8958
R18921 vdd.n2377 vdd.n771 72.8958
R18922 vdd.n2377 vdd.n770 72.8958
R18923 vdd.n2377 vdd.n769 72.8958
R18924 vdd.n2377 vdd.n768 72.8958
R18925 vdd.n2377 vdd.n767 72.8958
R18926 vdd.n2377 vdd.n766 72.8958
R18927 vdd.n2377 vdd.n765 72.8958
R18928 vdd.n2377 vdd.n764 72.8958
R18929 vdd.n2377 vdd.n763 72.8958
R18930 vdd.n2377 vdd.n762 72.8958
R18931 vdd.n2130 vdd.n2129 72.8958
R18932 vdd.n2129 vdd.n928 72.8958
R18933 vdd.n2129 vdd.n929 72.8958
R18934 vdd.n2129 vdd.n930 72.8958
R18935 vdd.n2129 vdd.n931 72.8958
R18936 vdd.n2129 vdd.n932 72.8958
R18937 vdd.n2129 vdd.n933 72.8958
R18938 vdd.n2129 vdd.n934 72.8958
R18939 vdd.n2129 vdd.n935 72.8958
R18940 vdd.n2129 vdd.n936 72.8958
R18941 vdd.n2129 vdd.n937 72.8958
R18942 vdd.n2129 vdd.n938 72.8958
R18943 vdd.n2129 vdd.n939 72.8958
R18944 vdd.n2129 vdd.n940 72.8958
R18945 vdd.n2129 vdd.n941 72.8958
R18946 vdd.n2129 vdd.n942 72.8958
R18947 vdd.n2129 vdd.n943 72.8958
R18948 vdd.n1348 vdd.n1344 66.2847
R18949 vdd.n1354 vdd.n1344 66.2847
R18950 vdd.n1357 vdd.n1344 66.2847
R18951 vdd.n1362 vdd.n1344 66.2847
R18952 vdd.n1365 vdd.n1344 66.2847
R18953 vdd.n1370 vdd.n1344 66.2847
R18954 vdd.n1373 vdd.n1344 66.2847
R18955 vdd.n1378 vdd.n1344 66.2847
R18956 vdd.n1381 vdd.n1344 66.2847
R18957 vdd.n1388 vdd.n1344 66.2847
R18958 vdd.n1391 vdd.n1344 66.2847
R18959 vdd.n1396 vdd.n1344 66.2847
R18960 vdd.n1399 vdd.n1344 66.2847
R18961 vdd.n1404 vdd.n1344 66.2847
R18962 vdd.n1407 vdd.n1344 66.2847
R18963 vdd.n1412 vdd.n1344 66.2847
R18964 vdd.n1415 vdd.n1344 66.2847
R18965 vdd.n1420 vdd.n1344 66.2847
R18966 vdd.n1423 vdd.n1344 66.2847
R18967 vdd.n1428 vdd.n1344 66.2847
R18968 vdd.n1507 vdd.n1344 66.2847
R18969 vdd.n1431 vdd.n1344 66.2847
R18970 vdd.n1437 vdd.n1344 66.2847
R18971 vdd.n1442 vdd.n1344 66.2847
R18972 vdd.n1445 vdd.n1344 66.2847
R18973 vdd.n1450 vdd.n1344 66.2847
R18974 vdd.n1453 vdd.n1344 66.2847
R18975 vdd.n1458 vdd.n1344 66.2847
R18976 vdd.n1461 vdd.n1344 66.2847
R18977 vdd.n1466 vdd.n1344 66.2847
R18978 vdd.n1469 vdd.n1344 66.2847
R18979 vdd.n1261 vdd.n911 66.2847
R18980 vdd.n1258 vdd.n911 66.2847
R18981 vdd.n1254 vdd.n911 66.2847
R18982 vdd.n1991 vdd.n911 66.2847
R18983 vdd.n1045 vdd.n911 66.2847
R18984 vdd.n1998 vdd.n911 66.2847
R18985 vdd.n1038 vdd.n911 66.2847
R18986 vdd.n2005 vdd.n911 66.2847
R18987 vdd.n1031 vdd.n911 66.2847
R18988 vdd.n2012 vdd.n911 66.2847
R18989 vdd.n1025 vdd.n911 66.2847
R18990 vdd.n1020 vdd.n911 66.2847
R18991 vdd.n2023 vdd.n911 66.2847
R18992 vdd.n1012 vdd.n911 66.2847
R18993 vdd.n2030 vdd.n911 66.2847
R18994 vdd.n1005 vdd.n911 66.2847
R18995 vdd.n2037 vdd.n911 66.2847
R18996 vdd.n998 vdd.n911 66.2847
R18997 vdd.n2044 vdd.n911 66.2847
R18998 vdd.n991 vdd.n911 66.2847
R18999 vdd.n2051 vdd.n911 66.2847
R19000 vdd.n985 vdd.n911 66.2847
R19001 vdd.n980 vdd.n911 66.2847
R19002 vdd.n2062 vdd.n911 66.2847
R19003 vdd.n972 vdd.n911 66.2847
R19004 vdd.n2069 vdd.n911 66.2847
R19005 vdd.n965 vdd.n911 66.2847
R19006 vdd.n2076 vdd.n911 66.2847
R19007 vdd.n958 vdd.n911 66.2847
R19008 vdd.n2083 vdd.n911 66.2847
R19009 vdd.n2088 vdd.n911 66.2847
R19010 vdd.n954 vdd.n911 66.2847
R19011 vdd.n3024 vdd.n516 66.2847
R19012 vdd.n520 vdd.n516 66.2847
R19013 vdd.n523 vdd.n516 66.2847
R19014 vdd.n3013 vdd.n516 66.2847
R19015 vdd.n3007 vdd.n516 66.2847
R19016 vdd.n3005 vdd.n516 66.2847
R19017 vdd.n2999 vdd.n516 66.2847
R19018 vdd.n2997 vdd.n516 66.2847
R19019 vdd.n2991 vdd.n516 66.2847
R19020 vdd.n2989 vdd.n516 66.2847
R19021 vdd.n2983 vdd.n516 66.2847
R19022 vdd.n2981 vdd.n516 66.2847
R19023 vdd.n2975 vdd.n516 66.2847
R19024 vdd.n2973 vdd.n516 66.2847
R19025 vdd.n2967 vdd.n516 66.2847
R19026 vdd.n2965 vdd.n516 66.2847
R19027 vdd.n2959 vdd.n516 66.2847
R19028 vdd.n2957 vdd.n516 66.2847
R19029 vdd.n2951 vdd.n516 66.2847
R19030 vdd.n2949 vdd.n516 66.2847
R19031 vdd.n584 vdd.n516 66.2847
R19032 vdd.n2940 vdd.n516 66.2847
R19033 vdd.n586 vdd.n516 66.2847
R19034 vdd.n2933 vdd.n516 66.2847
R19035 vdd.n2927 vdd.n516 66.2847
R19036 vdd.n2925 vdd.n516 66.2847
R19037 vdd.n2919 vdd.n516 66.2847
R19038 vdd.n2917 vdd.n516 66.2847
R19039 vdd.n2911 vdd.n516 66.2847
R19040 vdd.n607 vdd.n516 66.2847
R19041 vdd.n609 vdd.n516 66.2847
R19042 vdd.n3110 vdd.n351 66.2847
R19043 vdd.n3119 vdd.n351 66.2847
R19044 vdd.n461 vdd.n351 66.2847
R19045 vdd.n3126 vdd.n351 66.2847
R19046 vdd.n454 vdd.n351 66.2847
R19047 vdd.n3133 vdd.n351 66.2847
R19048 vdd.n447 vdd.n351 66.2847
R19049 vdd.n3140 vdd.n351 66.2847
R19050 vdd.n440 vdd.n351 66.2847
R19051 vdd.n3147 vdd.n351 66.2847
R19052 vdd.n434 vdd.n351 66.2847
R19053 vdd.n429 vdd.n351 66.2847
R19054 vdd.n3158 vdd.n351 66.2847
R19055 vdd.n421 vdd.n351 66.2847
R19056 vdd.n3165 vdd.n351 66.2847
R19057 vdd.n414 vdd.n351 66.2847
R19058 vdd.n3172 vdd.n351 66.2847
R19059 vdd.n407 vdd.n351 66.2847
R19060 vdd.n3179 vdd.n351 66.2847
R19061 vdd.n400 vdd.n351 66.2847
R19062 vdd.n3186 vdd.n351 66.2847
R19063 vdd.n394 vdd.n351 66.2847
R19064 vdd.n389 vdd.n351 66.2847
R19065 vdd.n3197 vdd.n351 66.2847
R19066 vdd.n381 vdd.n351 66.2847
R19067 vdd.n3204 vdd.n351 66.2847
R19068 vdd.n374 vdd.n351 66.2847
R19069 vdd.n3211 vdd.n351 66.2847
R19070 vdd.n367 vdd.n351 66.2847
R19071 vdd.n3218 vdd.n351 66.2847
R19072 vdd.n3221 vdd.n351 66.2847
R19073 vdd.n355 vdd.n351 66.2847
R19074 vdd.n356 vdd.n355 52.4337
R19075 vdd.n3221 vdd.n3220 52.4337
R19076 vdd.n3218 vdd.n3217 52.4337
R19077 vdd.n3213 vdd.n367 52.4337
R19078 vdd.n3211 vdd.n3210 52.4337
R19079 vdd.n3206 vdd.n374 52.4337
R19080 vdd.n3204 vdd.n3203 52.4337
R19081 vdd.n3199 vdd.n381 52.4337
R19082 vdd.n3197 vdd.n3196 52.4337
R19083 vdd.n390 vdd.n389 52.4337
R19084 vdd.n3188 vdd.n394 52.4337
R19085 vdd.n3186 vdd.n3185 52.4337
R19086 vdd.n3181 vdd.n400 52.4337
R19087 vdd.n3179 vdd.n3178 52.4337
R19088 vdd.n3174 vdd.n407 52.4337
R19089 vdd.n3172 vdd.n3171 52.4337
R19090 vdd.n3167 vdd.n414 52.4337
R19091 vdd.n3165 vdd.n3164 52.4337
R19092 vdd.n3160 vdd.n421 52.4337
R19093 vdd.n3158 vdd.n3157 52.4337
R19094 vdd.n430 vdd.n429 52.4337
R19095 vdd.n3149 vdd.n434 52.4337
R19096 vdd.n3147 vdd.n3146 52.4337
R19097 vdd.n3142 vdd.n440 52.4337
R19098 vdd.n3140 vdd.n3139 52.4337
R19099 vdd.n3135 vdd.n447 52.4337
R19100 vdd.n3133 vdd.n3132 52.4337
R19101 vdd.n3128 vdd.n454 52.4337
R19102 vdd.n3126 vdd.n3125 52.4337
R19103 vdd.n3121 vdd.n461 52.4337
R19104 vdd.n3119 vdd.n3118 52.4337
R19105 vdd.n3111 vdd.n3110 52.4337
R19106 vdd.n3024 vdd.n517 52.4337
R19107 vdd.n3022 vdd.n520 52.4337
R19108 vdd.n3018 vdd.n523 52.4337
R19109 vdd.n3014 vdd.n3013 52.4337
R19110 vdd.n3007 vdd.n526 52.4337
R19111 vdd.n3006 vdd.n3005 52.4337
R19112 vdd.n2999 vdd.n532 52.4337
R19113 vdd.n2998 vdd.n2997 52.4337
R19114 vdd.n2991 vdd.n538 52.4337
R19115 vdd.n2990 vdd.n2989 52.4337
R19116 vdd.n2983 vdd.n546 52.4337
R19117 vdd.n2982 vdd.n2981 52.4337
R19118 vdd.n2975 vdd.n552 52.4337
R19119 vdd.n2974 vdd.n2973 52.4337
R19120 vdd.n2967 vdd.n558 52.4337
R19121 vdd.n2966 vdd.n2965 52.4337
R19122 vdd.n2959 vdd.n564 52.4337
R19123 vdd.n2958 vdd.n2957 52.4337
R19124 vdd.n2951 vdd.n570 52.4337
R19125 vdd.n2950 vdd.n2949 52.4337
R19126 vdd.n584 vdd.n576 52.4337
R19127 vdd.n2941 vdd.n2940 52.4337
R19128 vdd.n2938 vdd.n586 52.4337
R19129 vdd.n2934 vdd.n2933 52.4337
R19130 vdd.n2927 vdd.n590 52.4337
R19131 vdd.n2926 vdd.n2925 52.4337
R19132 vdd.n2919 vdd.n596 52.4337
R19133 vdd.n2918 vdd.n2917 52.4337
R19134 vdd.n2911 vdd.n602 52.4337
R19135 vdd.n2910 vdd.n607 52.4337
R19136 vdd.n2906 vdd.n609 52.4337
R19137 vdd.n2090 vdd.n954 52.4337
R19138 vdd.n2088 vdd.n2087 52.4337
R19139 vdd.n2083 vdd.n2082 52.4337
R19140 vdd.n2078 vdd.n958 52.4337
R19141 vdd.n2076 vdd.n2075 52.4337
R19142 vdd.n2071 vdd.n965 52.4337
R19143 vdd.n2069 vdd.n2068 52.4337
R19144 vdd.n2064 vdd.n972 52.4337
R19145 vdd.n2062 vdd.n2061 52.4337
R19146 vdd.n981 vdd.n980 52.4337
R19147 vdd.n2053 vdd.n985 52.4337
R19148 vdd.n2051 vdd.n2050 52.4337
R19149 vdd.n2046 vdd.n991 52.4337
R19150 vdd.n2044 vdd.n2043 52.4337
R19151 vdd.n2039 vdd.n998 52.4337
R19152 vdd.n2037 vdd.n2036 52.4337
R19153 vdd.n2032 vdd.n1005 52.4337
R19154 vdd.n2030 vdd.n2029 52.4337
R19155 vdd.n2025 vdd.n1012 52.4337
R19156 vdd.n2023 vdd.n2022 52.4337
R19157 vdd.n1021 vdd.n1020 52.4337
R19158 vdd.n2014 vdd.n1025 52.4337
R19159 vdd.n2012 vdd.n2011 52.4337
R19160 vdd.n2007 vdd.n1031 52.4337
R19161 vdd.n2005 vdd.n2004 52.4337
R19162 vdd.n2000 vdd.n1038 52.4337
R19163 vdd.n1998 vdd.n1997 52.4337
R19164 vdd.n1993 vdd.n1045 52.4337
R19165 vdd.n1991 vdd.n1990 52.4337
R19166 vdd.n1255 vdd.n1254 52.4337
R19167 vdd.n1259 vdd.n1258 52.4337
R19168 vdd.n1979 vdd.n1261 52.4337
R19169 vdd.n1348 vdd.n1346 52.4337
R19170 vdd.n1354 vdd.n1353 52.4337
R19171 vdd.n1357 vdd.n1356 52.4337
R19172 vdd.n1362 vdd.n1361 52.4337
R19173 vdd.n1365 vdd.n1364 52.4337
R19174 vdd.n1370 vdd.n1369 52.4337
R19175 vdd.n1373 vdd.n1372 52.4337
R19176 vdd.n1378 vdd.n1377 52.4337
R19177 vdd.n1381 vdd.n1380 52.4337
R19178 vdd.n1388 vdd.n1387 52.4337
R19179 vdd.n1391 vdd.n1390 52.4337
R19180 vdd.n1396 vdd.n1395 52.4337
R19181 vdd.n1399 vdd.n1398 52.4337
R19182 vdd.n1404 vdd.n1403 52.4337
R19183 vdd.n1407 vdd.n1406 52.4337
R19184 vdd.n1412 vdd.n1411 52.4337
R19185 vdd.n1415 vdd.n1414 52.4337
R19186 vdd.n1420 vdd.n1419 52.4337
R19187 vdd.n1423 vdd.n1422 52.4337
R19188 vdd.n1428 vdd.n1427 52.4337
R19189 vdd.n1508 vdd.n1507 52.4337
R19190 vdd.n1505 vdd.n1431 52.4337
R19191 vdd.n1437 vdd.n1436 52.4337
R19192 vdd.n1442 vdd.n1439 52.4337
R19193 vdd.n1445 vdd.n1444 52.4337
R19194 vdd.n1450 vdd.n1447 52.4337
R19195 vdd.n1453 vdd.n1452 52.4337
R19196 vdd.n1458 vdd.n1455 52.4337
R19197 vdd.n1461 vdd.n1460 52.4337
R19198 vdd.n1466 vdd.n1463 52.4337
R19199 vdd.n1469 vdd.n1468 52.4337
R19200 vdd.n1349 vdd.n1348 52.4337
R19201 vdd.n1355 vdd.n1354 52.4337
R19202 vdd.n1358 vdd.n1357 52.4337
R19203 vdd.n1363 vdd.n1362 52.4337
R19204 vdd.n1366 vdd.n1365 52.4337
R19205 vdd.n1371 vdd.n1370 52.4337
R19206 vdd.n1374 vdd.n1373 52.4337
R19207 vdd.n1379 vdd.n1378 52.4337
R19208 vdd.n1382 vdd.n1381 52.4337
R19209 vdd.n1389 vdd.n1388 52.4337
R19210 vdd.n1392 vdd.n1391 52.4337
R19211 vdd.n1397 vdd.n1396 52.4337
R19212 vdd.n1400 vdd.n1399 52.4337
R19213 vdd.n1405 vdd.n1404 52.4337
R19214 vdd.n1408 vdd.n1407 52.4337
R19215 vdd.n1413 vdd.n1412 52.4337
R19216 vdd.n1416 vdd.n1415 52.4337
R19217 vdd.n1421 vdd.n1420 52.4337
R19218 vdd.n1424 vdd.n1423 52.4337
R19219 vdd.n1429 vdd.n1428 52.4337
R19220 vdd.n1507 vdd.n1506 52.4337
R19221 vdd.n1435 vdd.n1431 52.4337
R19222 vdd.n1438 vdd.n1437 52.4337
R19223 vdd.n1443 vdd.n1442 52.4337
R19224 vdd.n1446 vdd.n1445 52.4337
R19225 vdd.n1451 vdd.n1450 52.4337
R19226 vdd.n1454 vdd.n1453 52.4337
R19227 vdd.n1459 vdd.n1458 52.4337
R19228 vdd.n1462 vdd.n1461 52.4337
R19229 vdd.n1467 vdd.n1466 52.4337
R19230 vdd.n1470 vdd.n1469 52.4337
R19231 vdd.n1261 vdd.n1260 52.4337
R19232 vdd.n1258 vdd.n1257 52.4337
R19233 vdd.n1254 vdd.n1046 52.4337
R19234 vdd.n1992 vdd.n1991 52.4337
R19235 vdd.n1045 vdd.n1039 52.4337
R19236 vdd.n1999 vdd.n1998 52.4337
R19237 vdd.n1038 vdd.n1032 52.4337
R19238 vdd.n2006 vdd.n2005 52.4337
R19239 vdd.n1031 vdd.n1026 52.4337
R19240 vdd.n2013 vdd.n2012 52.4337
R19241 vdd.n1025 vdd.n1024 52.4337
R19242 vdd.n1020 vdd.n1013 52.4337
R19243 vdd.n2024 vdd.n2023 52.4337
R19244 vdd.n1012 vdd.n1006 52.4337
R19245 vdd.n2031 vdd.n2030 52.4337
R19246 vdd.n1005 vdd.n999 52.4337
R19247 vdd.n2038 vdd.n2037 52.4337
R19248 vdd.n998 vdd.n992 52.4337
R19249 vdd.n2045 vdd.n2044 52.4337
R19250 vdd.n991 vdd.n986 52.4337
R19251 vdd.n2052 vdd.n2051 52.4337
R19252 vdd.n985 vdd.n984 52.4337
R19253 vdd.n980 vdd.n973 52.4337
R19254 vdd.n2063 vdd.n2062 52.4337
R19255 vdd.n972 vdd.n966 52.4337
R19256 vdd.n2070 vdd.n2069 52.4337
R19257 vdd.n965 vdd.n959 52.4337
R19258 vdd.n2077 vdd.n2076 52.4337
R19259 vdd.n958 vdd.n955 52.4337
R19260 vdd.n2084 vdd.n2083 52.4337
R19261 vdd.n2089 vdd.n2088 52.4337
R19262 vdd.n1265 vdd.n954 52.4337
R19263 vdd.n3025 vdd.n3024 52.4337
R19264 vdd.n3019 vdd.n520 52.4337
R19265 vdd.n3015 vdd.n523 52.4337
R19266 vdd.n3013 vdd.n3012 52.4337
R19267 vdd.n3008 vdd.n3007 52.4337
R19268 vdd.n3005 vdd.n3004 52.4337
R19269 vdd.n3000 vdd.n2999 52.4337
R19270 vdd.n2997 vdd.n2996 52.4337
R19271 vdd.n2992 vdd.n2991 52.4337
R19272 vdd.n2989 vdd.n2988 52.4337
R19273 vdd.n2984 vdd.n2983 52.4337
R19274 vdd.n2981 vdd.n2980 52.4337
R19275 vdd.n2976 vdd.n2975 52.4337
R19276 vdd.n2973 vdd.n2972 52.4337
R19277 vdd.n2968 vdd.n2967 52.4337
R19278 vdd.n2965 vdd.n2964 52.4337
R19279 vdd.n2960 vdd.n2959 52.4337
R19280 vdd.n2957 vdd.n2956 52.4337
R19281 vdd.n2952 vdd.n2951 52.4337
R19282 vdd.n2949 vdd.n2948 52.4337
R19283 vdd.n585 vdd.n584 52.4337
R19284 vdd.n2940 vdd.n2939 52.4337
R19285 vdd.n2935 vdd.n586 52.4337
R19286 vdd.n2933 vdd.n2932 52.4337
R19287 vdd.n2928 vdd.n2927 52.4337
R19288 vdd.n2925 vdd.n2924 52.4337
R19289 vdd.n2920 vdd.n2919 52.4337
R19290 vdd.n2917 vdd.n2916 52.4337
R19291 vdd.n2912 vdd.n2911 52.4337
R19292 vdd.n2907 vdd.n607 52.4337
R19293 vdd.n2903 vdd.n609 52.4337
R19294 vdd.n3110 vdd.n462 52.4337
R19295 vdd.n3120 vdd.n3119 52.4337
R19296 vdd.n461 vdd.n455 52.4337
R19297 vdd.n3127 vdd.n3126 52.4337
R19298 vdd.n454 vdd.n448 52.4337
R19299 vdd.n3134 vdd.n3133 52.4337
R19300 vdd.n447 vdd.n441 52.4337
R19301 vdd.n3141 vdd.n3140 52.4337
R19302 vdd.n440 vdd.n435 52.4337
R19303 vdd.n3148 vdd.n3147 52.4337
R19304 vdd.n434 vdd.n433 52.4337
R19305 vdd.n429 vdd.n422 52.4337
R19306 vdd.n3159 vdd.n3158 52.4337
R19307 vdd.n421 vdd.n415 52.4337
R19308 vdd.n3166 vdd.n3165 52.4337
R19309 vdd.n414 vdd.n408 52.4337
R19310 vdd.n3173 vdd.n3172 52.4337
R19311 vdd.n407 vdd.n401 52.4337
R19312 vdd.n3180 vdd.n3179 52.4337
R19313 vdd.n400 vdd.n395 52.4337
R19314 vdd.n3187 vdd.n3186 52.4337
R19315 vdd.n394 vdd.n393 52.4337
R19316 vdd.n389 vdd.n382 52.4337
R19317 vdd.n3198 vdd.n3197 52.4337
R19318 vdd.n381 vdd.n375 52.4337
R19319 vdd.n3205 vdd.n3204 52.4337
R19320 vdd.n374 vdd.n368 52.4337
R19321 vdd.n3212 vdd.n3211 52.4337
R19322 vdd.n367 vdd.n360 52.4337
R19323 vdd.n3219 vdd.n3218 52.4337
R19324 vdd.n3222 vdd.n3221 52.4337
R19325 vdd.n355 vdd.n352 52.4337
R19326 vdd.t114 vdd.t120 51.4683
R19327 vdd.n258 vdd.n256 42.0461
R19328 vdd.n164 vdd.n162 42.0461
R19329 vdd.n71 vdd.n69 42.0461
R19330 vdd.n1866 vdd.n1864 42.0461
R19331 vdd.n1772 vdd.n1770 42.0461
R19332 vdd.n1679 vdd.n1677 42.0461
R19333 vdd.n308 vdd.n307 41.6884
R19334 vdd.n214 vdd.n213 41.6884
R19335 vdd.n121 vdd.n120 41.6884
R19336 vdd.n1916 vdd.n1915 41.6884
R19337 vdd.n1822 vdd.n1821 41.6884
R19338 vdd.n1729 vdd.n1728 41.6884
R19339 vdd.n1474 vdd.n1473 41.1157
R19340 vdd.n1511 vdd.n1510 41.1157
R19341 vdd.n1385 vdd.n1384 41.1157
R19342 vdd.n3115 vdd.n3114 41.1157
R19343 vdd.n3154 vdd.n428 41.1157
R19344 vdd.n3193 vdd.n388 41.1157
R19345 vdd.n2857 vdd.n2856 39.2114
R19346 vdd.n2854 vdd.n2853 39.2114
R19347 vdd.n2849 vdd.n641 39.2114
R19348 vdd.n2847 vdd.n2846 39.2114
R19349 vdd.n2842 vdd.n644 39.2114
R19350 vdd.n2840 vdd.n2839 39.2114
R19351 vdd.n2835 vdd.n647 39.2114
R19352 vdd.n2833 vdd.n2832 39.2114
R19353 vdd.n2827 vdd.n650 39.2114
R19354 vdd.n2825 vdd.n2824 39.2114
R19355 vdd.n2820 vdd.n653 39.2114
R19356 vdd.n2818 vdd.n2817 39.2114
R19357 vdd.n2813 vdd.n656 39.2114
R19358 vdd.n2811 vdd.n2810 39.2114
R19359 vdd.n2806 vdd.n659 39.2114
R19360 vdd.n2804 vdd.n2803 39.2114
R19361 vdd.n2799 vdd.n2798 39.2114
R19362 vdd.n2649 vdd.n2648 39.2114
R19363 vdd.n2643 vdd.n2378 39.2114
R19364 vdd.n2640 vdd.n2379 39.2114
R19365 vdd.n2636 vdd.n2380 39.2114
R19366 vdd.n2632 vdd.n2381 39.2114
R19367 vdd.n2628 vdd.n2382 39.2114
R19368 vdd.n2624 vdd.n2383 39.2114
R19369 vdd.n2620 vdd.n2384 39.2114
R19370 vdd.n2616 vdd.n2385 39.2114
R19371 vdd.n2612 vdd.n2386 39.2114
R19372 vdd.n2608 vdd.n2387 39.2114
R19373 vdd.n2604 vdd.n2388 39.2114
R19374 vdd.n2600 vdd.n2389 39.2114
R19375 vdd.n2596 vdd.n2390 39.2114
R19376 vdd.n2592 vdd.n2391 39.2114
R19377 vdd.n2588 vdd.n2392 39.2114
R19378 vdd.n2583 vdd.n2393 39.2114
R19379 vdd.n2372 vdd.n796 39.2114
R19380 vdd.n2368 vdd.n795 39.2114
R19381 vdd.n2364 vdd.n794 39.2114
R19382 vdd.n2360 vdd.n793 39.2114
R19383 vdd.n2356 vdd.n792 39.2114
R19384 vdd.n2352 vdd.n791 39.2114
R19385 vdd.n2348 vdd.n790 39.2114
R19386 vdd.n2344 vdd.n789 39.2114
R19387 vdd.n2340 vdd.n788 39.2114
R19388 vdd.n2336 vdd.n787 39.2114
R19389 vdd.n2332 vdd.n786 39.2114
R19390 vdd.n2328 vdd.n785 39.2114
R19391 vdd.n2324 vdd.n784 39.2114
R19392 vdd.n2320 vdd.n783 39.2114
R19393 vdd.n2316 vdd.n782 39.2114
R19394 vdd.n2311 vdd.n781 39.2114
R19395 vdd.n2307 vdd.n780 39.2114
R19396 vdd.n2128 vdd.n2127 39.2114
R19397 vdd.n2122 vdd.n912 39.2114
R19398 vdd.n2119 vdd.n913 39.2114
R19399 vdd.n2115 vdd.n914 39.2114
R19400 vdd.n2111 vdd.n915 39.2114
R19401 vdd.n2107 vdd.n916 39.2114
R19402 vdd.n2103 vdd.n917 39.2114
R19403 vdd.n2099 vdd.n918 39.2114
R19404 vdd.n2095 vdd.n919 39.2114
R19405 vdd.n1104 vdd.n920 39.2114
R19406 vdd.n1108 vdd.n921 39.2114
R19407 vdd.n1112 vdd.n922 39.2114
R19408 vdd.n1116 vdd.n923 39.2114
R19409 vdd.n1120 vdd.n924 39.2114
R19410 vdd.n1124 vdd.n925 39.2114
R19411 vdd.n1128 vdd.n926 39.2114
R19412 vdd.n1133 vdd.n927 39.2114
R19413 vdd.n2776 vdd.n2775 39.2114
R19414 vdd.n2771 vdd.n2743 39.2114
R19415 vdd.n2769 vdd.n2768 39.2114
R19416 vdd.n2764 vdd.n2746 39.2114
R19417 vdd.n2762 vdd.n2761 39.2114
R19418 vdd.n2757 vdd.n2749 39.2114
R19419 vdd.n2755 vdd.n2754 39.2114
R19420 vdd.n2750 vdd.n612 39.2114
R19421 vdd.n2894 vdd.n2893 39.2114
R19422 vdd.n2891 vdd.n2890 39.2114
R19423 vdd.n2886 vdd.n617 39.2114
R19424 vdd.n2884 vdd.n2883 39.2114
R19425 vdd.n2879 vdd.n620 39.2114
R19426 vdd.n2877 vdd.n2876 39.2114
R19427 vdd.n2872 vdd.n623 39.2114
R19428 vdd.n2870 vdd.n2869 39.2114
R19429 vdd.n2865 vdd.n629 39.2114
R19430 vdd.n2652 vdd.n2651 39.2114
R19431 vdd.n2419 vdd.n2394 39.2114
R19432 vdd.n2423 vdd.n2395 39.2114
R19433 vdd.n2427 vdd.n2396 39.2114
R19434 vdd.n2431 vdd.n2397 39.2114
R19435 vdd.n2435 vdd.n2398 39.2114
R19436 vdd.n2439 vdd.n2399 39.2114
R19437 vdd.n2443 vdd.n2400 39.2114
R19438 vdd.n2447 vdd.n2401 39.2114
R19439 vdd.n2451 vdd.n2402 39.2114
R19440 vdd.n2455 vdd.n2403 39.2114
R19441 vdd.n2459 vdd.n2404 39.2114
R19442 vdd.n2463 vdd.n2405 39.2114
R19443 vdd.n2467 vdd.n2406 39.2114
R19444 vdd.n2471 vdd.n2407 39.2114
R19445 vdd.n2475 vdd.n2408 39.2114
R19446 vdd.n2479 vdd.n2409 39.2114
R19447 vdd.n2651 vdd.n761 39.2114
R19448 vdd.n2422 vdd.n2394 39.2114
R19449 vdd.n2426 vdd.n2395 39.2114
R19450 vdd.n2430 vdd.n2396 39.2114
R19451 vdd.n2434 vdd.n2397 39.2114
R19452 vdd.n2438 vdd.n2398 39.2114
R19453 vdd.n2442 vdd.n2399 39.2114
R19454 vdd.n2446 vdd.n2400 39.2114
R19455 vdd.n2450 vdd.n2401 39.2114
R19456 vdd.n2454 vdd.n2402 39.2114
R19457 vdd.n2458 vdd.n2403 39.2114
R19458 vdd.n2462 vdd.n2404 39.2114
R19459 vdd.n2466 vdd.n2405 39.2114
R19460 vdd.n2470 vdd.n2406 39.2114
R19461 vdd.n2474 vdd.n2407 39.2114
R19462 vdd.n2478 vdd.n2408 39.2114
R19463 vdd.n2481 vdd.n2409 39.2114
R19464 vdd.n629 vdd.n624 39.2114
R19465 vdd.n2871 vdd.n2870 39.2114
R19466 vdd.n623 vdd.n621 39.2114
R19467 vdd.n2878 vdd.n2877 39.2114
R19468 vdd.n620 vdd.n618 39.2114
R19469 vdd.n2885 vdd.n2884 39.2114
R19470 vdd.n617 vdd.n615 39.2114
R19471 vdd.n2892 vdd.n2891 39.2114
R19472 vdd.n2895 vdd.n2894 39.2114
R19473 vdd.n2751 vdd.n2750 39.2114
R19474 vdd.n2756 vdd.n2755 39.2114
R19475 vdd.n2749 vdd.n2747 39.2114
R19476 vdd.n2763 vdd.n2762 39.2114
R19477 vdd.n2746 vdd.n2744 39.2114
R19478 vdd.n2770 vdd.n2769 39.2114
R19479 vdd.n2743 vdd.n2741 39.2114
R19480 vdd.n2777 vdd.n2776 39.2114
R19481 vdd.n2128 vdd.n946 39.2114
R19482 vdd.n2120 vdd.n912 39.2114
R19483 vdd.n2116 vdd.n913 39.2114
R19484 vdd.n2112 vdd.n914 39.2114
R19485 vdd.n2108 vdd.n915 39.2114
R19486 vdd.n2104 vdd.n916 39.2114
R19487 vdd.n2100 vdd.n917 39.2114
R19488 vdd.n2096 vdd.n918 39.2114
R19489 vdd.n1103 vdd.n919 39.2114
R19490 vdd.n1107 vdd.n920 39.2114
R19491 vdd.n1111 vdd.n921 39.2114
R19492 vdd.n1115 vdd.n922 39.2114
R19493 vdd.n1119 vdd.n923 39.2114
R19494 vdd.n1123 vdd.n924 39.2114
R19495 vdd.n1127 vdd.n925 39.2114
R19496 vdd.n1132 vdd.n926 39.2114
R19497 vdd.n1136 vdd.n927 39.2114
R19498 vdd.n2310 vdd.n780 39.2114
R19499 vdd.n2315 vdd.n781 39.2114
R19500 vdd.n2319 vdd.n782 39.2114
R19501 vdd.n2323 vdd.n783 39.2114
R19502 vdd.n2327 vdd.n784 39.2114
R19503 vdd.n2331 vdd.n785 39.2114
R19504 vdd.n2335 vdd.n786 39.2114
R19505 vdd.n2339 vdd.n787 39.2114
R19506 vdd.n2343 vdd.n788 39.2114
R19507 vdd.n2347 vdd.n789 39.2114
R19508 vdd.n2351 vdd.n790 39.2114
R19509 vdd.n2355 vdd.n791 39.2114
R19510 vdd.n2359 vdd.n792 39.2114
R19511 vdd.n2363 vdd.n793 39.2114
R19512 vdd.n2367 vdd.n794 39.2114
R19513 vdd.n2371 vdd.n795 39.2114
R19514 vdd.n798 vdd.n796 39.2114
R19515 vdd.n2649 vdd.n2412 39.2114
R19516 vdd.n2641 vdd.n2378 39.2114
R19517 vdd.n2637 vdd.n2379 39.2114
R19518 vdd.n2633 vdd.n2380 39.2114
R19519 vdd.n2629 vdd.n2381 39.2114
R19520 vdd.n2625 vdd.n2382 39.2114
R19521 vdd.n2621 vdd.n2383 39.2114
R19522 vdd.n2617 vdd.n2384 39.2114
R19523 vdd.n2613 vdd.n2385 39.2114
R19524 vdd.n2609 vdd.n2386 39.2114
R19525 vdd.n2605 vdd.n2387 39.2114
R19526 vdd.n2601 vdd.n2388 39.2114
R19527 vdd.n2597 vdd.n2389 39.2114
R19528 vdd.n2593 vdd.n2390 39.2114
R19529 vdd.n2589 vdd.n2391 39.2114
R19530 vdd.n2584 vdd.n2392 39.2114
R19531 vdd.n2580 vdd.n2393 39.2114
R19532 vdd.n2798 vdd.n660 39.2114
R19533 vdd.n2805 vdd.n2804 39.2114
R19534 vdd.n659 vdd.n657 39.2114
R19535 vdd.n2812 vdd.n2811 39.2114
R19536 vdd.n656 vdd.n654 39.2114
R19537 vdd.n2819 vdd.n2818 39.2114
R19538 vdd.n653 vdd.n651 39.2114
R19539 vdd.n2826 vdd.n2825 39.2114
R19540 vdd.n650 vdd.n648 39.2114
R19541 vdd.n2834 vdd.n2833 39.2114
R19542 vdd.n647 vdd.n645 39.2114
R19543 vdd.n2841 vdd.n2840 39.2114
R19544 vdd.n644 vdd.n642 39.2114
R19545 vdd.n2848 vdd.n2847 39.2114
R19546 vdd.n641 vdd.n639 39.2114
R19547 vdd.n2855 vdd.n2854 39.2114
R19548 vdd.n2858 vdd.n2857 39.2114
R19549 vdd.n807 vdd.n762 39.2114
R19550 vdd.n2299 vdd.n763 39.2114
R19551 vdd.n2295 vdd.n764 39.2114
R19552 vdd.n2291 vdd.n765 39.2114
R19553 vdd.n2287 vdd.n766 39.2114
R19554 vdd.n2283 vdd.n767 39.2114
R19555 vdd.n2279 vdd.n768 39.2114
R19556 vdd.n2275 vdd.n769 39.2114
R19557 vdd.n2271 vdd.n770 39.2114
R19558 vdd.n2267 vdd.n771 39.2114
R19559 vdd.n2263 vdd.n772 39.2114
R19560 vdd.n2259 vdd.n773 39.2114
R19561 vdd.n2255 vdd.n774 39.2114
R19562 vdd.n2251 vdd.n775 39.2114
R19563 vdd.n2247 vdd.n776 39.2114
R19564 vdd.n2243 vdd.n777 39.2114
R19565 vdd.n2239 vdd.n778 39.2114
R19566 vdd.n2131 vdd.n2130 39.2114
R19567 vdd.n1050 vdd.n928 39.2114
R19568 vdd.n1054 vdd.n929 39.2114
R19569 vdd.n1058 vdd.n930 39.2114
R19570 vdd.n1062 vdd.n931 39.2114
R19571 vdd.n1066 vdd.n932 39.2114
R19572 vdd.n1070 vdd.n933 39.2114
R19573 vdd.n1074 vdd.n934 39.2114
R19574 vdd.n1078 vdd.n935 39.2114
R19575 vdd.n1248 vdd.n936 39.2114
R19576 vdd.n1245 vdd.n937 39.2114
R19577 vdd.n1241 vdd.n938 39.2114
R19578 vdd.n1237 vdd.n939 39.2114
R19579 vdd.n1233 vdd.n940 39.2114
R19580 vdd.n1229 vdd.n941 39.2114
R19581 vdd.n1225 vdd.n942 39.2114
R19582 vdd.n1221 vdd.n943 39.2114
R19583 vdd.n2236 vdd.n778 39.2114
R19584 vdd.n2240 vdd.n777 39.2114
R19585 vdd.n2244 vdd.n776 39.2114
R19586 vdd.n2248 vdd.n775 39.2114
R19587 vdd.n2252 vdd.n774 39.2114
R19588 vdd.n2256 vdd.n773 39.2114
R19589 vdd.n2260 vdd.n772 39.2114
R19590 vdd.n2264 vdd.n771 39.2114
R19591 vdd.n2268 vdd.n770 39.2114
R19592 vdd.n2272 vdd.n769 39.2114
R19593 vdd.n2276 vdd.n768 39.2114
R19594 vdd.n2280 vdd.n767 39.2114
R19595 vdd.n2284 vdd.n766 39.2114
R19596 vdd.n2288 vdd.n765 39.2114
R19597 vdd.n2292 vdd.n764 39.2114
R19598 vdd.n2296 vdd.n763 39.2114
R19599 vdd.n2300 vdd.n762 39.2114
R19600 vdd.n2130 vdd.n910 39.2114
R19601 vdd.n1053 vdd.n928 39.2114
R19602 vdd.n1057 vdd.n929 39.2114
R19603 vdd.n1061 vdd.n930 39.2114
R19604 vdd.n1065 vdd.n931 39.2114
R19605 vdd.n1069 vdd.n932 39.2114
R19606 vdd.n1073 vdd.n933 39.2114
R19607 vdd.n1077 vdd.n934 39.2114
R19608 vdd.n1080 vdd.n935 39.2114
R19609 vdd.n1246 vdd.n936 39.2114
R19610 vdd.n1242 vdd.n937 39.2114
R19611 vdd.n1238 vdd.n938 39.2114
R19612 vdd.n1234 vdd.n939 39.2114
R19613 vdd.n1230 vdd.n940 39.2114
R19614 vdd.n1226 vdd.n941 39.2114
R19615 vdd.n1222 vdd.n942 39.2114
R19616 vdd.n1218 vdd.n943 39.2114
R19617 vdd.n1983 vdd.n1982 37.2369
R19618 vdd.n2019 vdd.n1019 37.2369
R19619 vdd.n2058 vdd.n979 37.2369
R19620 vdd.n2946 vdd.n581 37.2369
R19621 vdd.n545 vdd.n544 37.2369
R19622 vdd.n2902 vdd.n2901 37.2369
R19623 vdd.n2126 vdd.n902 31.0639
R19624 vdd.n2375 vdd.n799 31.0639
R19625 vdd.n2308 vdd.n802 31.0639
R19626 vdd.n1138 vdd.n1135 31.0639
R19627 vdd.n2581 vdd.n2578 31.0639
R19628 vdd.n2800 vdd.n2797 31.0639
R19629 vdd.n2647 vdd.n754 31.0639
R19630 vdd.n2861 vdd.n2860 31.0639
R19631 vdd.n2780 vdd.n2779 31.0639
R19632 vdd.n2866 vdd.n628 31.0639
R19633 vdd.n2485 vdd.n2483 31.0639
R19634 vdd.n2654 vdd.n2653 31.0639
R19635 vdd.n2133 vdd.n2132 31.0639
R19636 vdd.n2303 vdd.n2302 31.0639
R19637 vdd.n2235 vdd.n2234 31.0639
R19638 vdd.n1217 vdd.n1216 31.0639
R19639 vdd.n1083 vdd.n1082 30.449
R19640 vdd.n811 vdd.n810 30.449
R19641 vdd.n1130 vdd.n1102 30.449
R19642 vdd.n2313 vdd.n801 30.449
R19643 vdd.n2418 vdd.n2417 30.449
R19644 vdd.n663 vdd.n662 30.449
R19645 vdd.n2586 vdd.n2414 30.449
R19646 vdd.n627 vdd.n626 30.449
R19647 vdd.n1577 vdd.n1344 20.633
R19648 vdd.n1977 vdd.n911 20.633
R19649 vdd.n3032 vdd.n516 20.633
R19650 vdd.n3230 vdd.n351 20.633
R19651 vdd.n1579 vdd.n1341 19.3944
R19652 vdd.n1583 vdd.n1341 19.3944
R19653 vdd.n1583 vdd.n1332 19.3944
R19654 vdd.n1595 vdd.n1332 19.3944
R19655 vdd.n1595 vdd.n1330 19.3944
R19656 vdd.n1599 vdd.n1330 19.3944
R19657 vdd.n1599 vdd.n1319 19.3944
R19658 vdd.n1611 vdd.n1319 19.3944
R19659 vdd.n1611 vdd.n1317 19.3944
R19660 vdd.n1615 vdd.n1317 19.3944
R19661 vdd.n1615 vdd.n1308 19.3944
R19662 vdd.n1628 vdd.n1308 19.3944
R19663 vdd.n1628 vdd.n1306 19.3944
R19664 vdd.n1632 vdd.n1306 19.3944
R19665 vdd.n1632 vdd.n1297 19.3944
R19666 vdd.n1926 vdd.n1297 19.3944
R19667 vdd.n1926 vdd.n1295 19.3944
R19668 vdd.n1930 vdd.n1295 19.3944
R19669 vdd.n1930 vdd.n1285 19.3944
R19670 vdd.n1943 vdd.n1285 19.3944
R19671 vdd.n1943 vdd.n1283 19.3944
R19672 vdd.n1947 vdd.n1283 19.3944
R19673 vdd.n1947 vdd.n1275 19.3944
R19674 vdd.n1960 vdd.n1275 19.3944
R19675 vdd.n1960 vdd.n1272 19.3944
R19676 vdd.n1966 vdd.n1272 19.3944
R19677 vdd.n1966 vdd.n1273 19.3944
R19678 vdd.n1273 vdd.n1263 19.3944
R19679 vdd.n1504 vdd.n1430 19.3944
R19680 vdd.n1504 vdd.n1432 19.3944
R19681 vdd.n1500 vdd.n1432 19.3944
R19682 vdd.n1500 vdd.n1499 19.3944
R19683 vdd.n1499 vdd.n1498 19.3944
R19684 vdd.n1498 vdd.n1440 19.3944
R19685 vdd.n1494 vdd.n1440 19.3944
R19686 vdd.n1494 vdd.n1493 19.3944
R19687 vdd.n1493 vdd.n1492 19.3944
R19688 vdd.n1492 vdd.n1448 19.3944
R19689 vdd.n1488 vdd.n1448 19.3944
R19690 vdd.n1488 vdd.n1487 19.3944
R19691 vdd.n1487 vdd.n1486 19.3944
R19692 vdd.n1486 vdd.n1456 19.3944
R19693 vdd.n1482 vdd.n1456 19.3944
R19694 vdd.n1482 vdd.n1481 19.3944
R19695 vdd.n1481 vdd.n1480 19.3944
R19696 vdd.n1480 vdd.n1464 19.3944
R19697 vdd.n1476 vdd.n1464 19.3944
R19698 vdd.n1476 vdd.n1475 19.3944
R19699 vdd.n1542 vdd.n1541 19.3944
R19700 vdd.n1541 vdd.n1540 19.3944
R19701 vdd.n1540 vdd.n1393 19.3944
R19702 vdd.n1536 vdd.n1393 19.3944
R19703 vdd.n1536 vdd.n1535 19.3944
R19704 vdd.n1535 vdd.n1534 19.3944
R19705 vdd.n1534 vdd.n1401 19.3944
R19706 vdd.n1530 vdd.n1401 19.3944
R19707 vdd.n1530 vdd.n1529 19.3944
R19708 vdd.n1529 vdd.n1528 19.3944
R19709 vdd.n1528 vdd.n1409 19.3944
R19710 vdd.n1524 vdd.n1409 19.3944
R19711 vdd.n1524 vdd.n1523 19.3944
R19712 vdd.n1523 vdd.n1522 19.3944
R19713 vdd.n1522 vdd.n1417 19.3944
R19714 vdd.n1518 vdd.n1417 19.3944
R19715 vdd.n1518 vdd.n1517 19.3944
R19716 vdd.n1517 vdd.n1516 19.3944
R19717 vdd.n1516 vdd.n1425 19.3944
R19718 vdd.n1512 vdd.n1425 19.3944
R19719 vdd.n1572 vdd.n1571 19.3944
R19720 vdd.n1571 vdd.n1570 19.3944
R19721 vdd.n1570 vdd.n1351 19.3944
R19722 vdd.n1566 vdd.n1351 19.3944
R19723 vdd.n1566 vdd.n1565 19.3944
R19724 vdd.n1565 vdd.n1564 19.3944
R19725 vdd.n1564 vdd.n1359 19.3944
R19726 vdd.n1560 vdd.n1359 19.3944
R19727 vdd.n1560 vdd.n1559 19.3944
R19728 vdd.n1559 vdd.n1558 19.3944
R19729 vdd.n1558 vdd.n1367 19.3944
R19730 vdd.n1554 vdd.n1367 19.3944
R19731 vdd.n1554 vdd.n1553 19.3944
R19732 vdd.n1553 vdd.n1552 19.3944
R19733 vdd.n1552 vdd.n1375 19.3944
R19734 vdd.n1548 vdd.n1375 19.3944
R19735 vdd.n1548 vdd.n1547 19.3944
R19736 vdd.n1547 vdd.n1546 19.3944
R19737 vdd.n2015 vdd.n1017 19.3944
R19738 vdd.n2015 vdd.n1023 19.3944
R19739 vdd.n2010 vdd.n1023 19.3944
R19740 vdd.n2010 vdd.n2009 19.3944
R19741 vdd.n2009 vdd.n2008 19.3944
R19742 vdd.n2008 vdd.n1030 19.3944
R19743 vdd.n2003 vdd.n1030 19.3944
R19744 vdd.n2003 vdd.n2002 19.3944
R19745 vdd.n2002 vdd.n2001 19.3944
R19746 vdd.n2001 vdd.n1037 19.3944
R19747 vdd.n1996 vdd.n1037 19.3944
R19748 vdd.n1996 vdd.n1995 19.3944
R19749 vdd.n1995 vdd.n1994 19.3944
R19750 vdd.n1994 vdd.n1044 19.3944
R19751 vdd.n1989 vdd.n1044 19.3944
R19752 vdd.n1989 vdd.n1988 19.3944
R19753 vdd.n1256 vdd.n1049 19.3944
R19754 vdd.n1984 vdd.n1253 19.3944
R19755 vdd.n2054 vdd.n977 19.3944
R19756 vdd.n2054 vdd.n983 19.3944
R19757 vdd.n2049 vdd.n983 19.3944
R19758 vdd.n2049 vdd.n2048 19.3944
R19759 vdd.n2048 vdd.n2047 19.3944
R19760 vdd.n2047 vdd.n990 19.3944
R19761 vdd.n2042 vdd.n990 19.3944
R19762 vdd.n2042 vdd.n2041 19.3944
R19763 vdd.n2041 vdd.n2040 19.3944
R19764 vdd.n2040 vdd.n997 19.3944
R19765 vdd.n2035 vdd.n997 19.3944
R19766 vdd.n2035 vdd.n2034 19.3944
R19767 vdd.n2034 vdd.n2033 19.3944
R19768 vdd.n2033 vdd.n1004 19.3944
R19769 vdd.n2028 vdd.n1004 19.3944
R19770 vdd.n2028 vdd.n2027 19.3944
R19771 vdd.n2027 vdd.n2026 19.3944
R19772 vdd.n2026 vdd.n1011 19.3944
R19773 vdd.n2021 vdd.n1011 19.3944
R19774 vdd.n2021 vdd.n2020 19.3944
R19775 vdd.n2091 vdd.n952 19.3944
R19776 vdd.n2091 vdd.n953 19.3944
R19777 vdd.n2086 vdd.n2085 19.3944
R19778 vdd.n2081 vdd.n2080 19.3944
R19779 vdd.n2080 vdd.n2079 19.3944
R19780 vdd.n2079 vdd.n957 19.3944
R19781 vdd.n2074 vdd.n957 19.3944
R19782 vdd.n2074 vdd.n2073 19.3944
R19783 vdd.n2073 vdd.n2072 19.3944
R19784 vdd.n2072 vdd.n964 19.3944
R19785 vdd.n2067 vdd.n964 19.3944
R19786 vdd.n2067 vdd.n2066 19.3944
R19787 vdd.n2066 vdd.n2065 19.3944
R19788 vdd.n2065 vdd.n971 19.3944
R19789 vdd.n2060 vdd.n971 19.3944
R19790 vdd.n2060 vdd.n2059 19.3944
R19791 vdd.n1575 vdd.n1338 19.3944
R19792 vdd.n1587 vdd.n1338 19.3944
R19793 vdd.n1587 vdd.n1336 19.3944
R19794 vdd.n1591 vdd.n1336 19.3944
R19795 vdd.n1591 vdd.n1326 19.3944
R19796 vdd.n1603 vdd.n1326 19.3944
R19797 vdd.n1603 vdd.n1324 19.3944
R19798 vdd.n1607 vdd.n1324 19.3944
R19799 vdd.n1607 vdd.n1314 19.3944
R19800 vdd.n1620 vdd.n1314 19.3944
R19801 vdd.n1620 vdd.n1312 19.3944
R19802 vdd.n1624 vdd.n1312 19.3944
R19803 vdd.n1624 vdd.n1303 19.3944
R19804 vdd.n1636 vdd.n1303 19.3944
R19805 vdd.n1636 vdd.n1301 19.3944
R19806 vdd.n1922 vdd.n1301 19.3944
R19807 vdd.n1922 vdd.n1291 19.3944
R19808 vdd.n1935 vdd.n1291 19.3944
R19809 vdd.n1935 vdd.n1289 19.3944
R19810 vdd.n1939 vdd.n1289 19.3944
R19811 vdd.n1939 vdd.n1280 19.3944
R19812 vdd.n1952 vdd.n1280 19.3944
R19813 vdd.n1952 vdd.n1278 19.3944
R19814 vdd.n1956 vdd.n1278 19.3944
R19815 vdd.n1956 vdd.n1268 19.3944
R19816 vdd.n1971 vdd.n1268 19.3944
R19817 vdd.n1971 vdd.n1266 19.3944
R19818 vdd.n1975 vdd.n1266 19.3944
R19819 vdd.n3034 vdd.n513 19.3944
R19820 vdd.n3038 vdd.n513 19.3944
R19821 vdd.n3038 vdd.n503 19.3944
R19822 vdd.n3050 vdd.n503 19.3944
R19823 vdd.n3050 vdd.n501 19.3944
R19824 vdd.n3054 vdd.n501 19.3944
R19825 vdd.n3054 vdd.n490 19.3944
R19826 vdd.n3066 vdd.n490 19.3944
R19827 vdd.n3066 vdd.n488 19.3944
R19828 vdd.n3070 vdd.n488 19.3944
R19829 vdd.n3070 vdd.n478 19.3944
R19830 vdd.n3083 vdd.n478 19.3944
R19831 vdd.n3083 vdd.n476 19.3944
R19832 vdd.n3087 vdd.n476 19.3944
R19833 vdd.n3088 vdd.n3087 19.3944
R19834 vdd.n3089 vdd.n3088 19.3944
R19835 vdd.n3089 vdd.n474 19.3944
R19836 vdd.n3093 vdd.n474 19.3944
R19837 vdd.n3094 vdd.n3093 19.3944
R19838 vdd.n3095 vdd.n3094 19.3944
R19839 vdd.n3095 vdd.n471 19.3944
R19840 vdd.n3099 vdd.n471 19.3944
R19841 vdd.n3100 vdd.n3099 19.3944
R19842 vdd.n3101 vdd.n3100 19.3944
R19843 vdd.n3101 vdd.n468 19.3944
R19844 vdd.n3105 vdd.n468 19.3944
R19845 vdd.n3106 vdd.n3105 19.3944
R19846 vdd.n3107 vdd.n3106 19.3944
R19847 vdd.n3150 vdd.n426 19.3944
R19848 vdd.n3150 vdd.n432 19.3944
R19849 vdd.n3145 vdd.n432 19.3944
R19850 vdd.n3145 vdd.n3144 19.3944
R19851 vdd.n3144 vdd.n3143 19.3944
R19852 vdd.n3143 vdd.n439 19.3944
R19853 vdd.n3138 vdd.n439 19.3944
R19854 vdd.n3138 vdd.n3137 19.3944
R19855 vdd.n3137 vdd.n3136 19.3944
R19856 vdd.n3136 vdd.n446 19.3944
R19857 vdd.n3131 vdd.n446 19.3944
R19858 vdd.n3131 vdd.n3130 19.3944
R19859 vdd.n3130 vdd.n3129 19.3944
R19860 vdd.n3129 vdd.n453 19.3944
R19861 vdd.n3124 vdd.n453 19.3944
R19862 vdd.n3124 vdd.n3123 19.3944
R19863 vdd.n3123 vdd.n3122 19.3944
R19864 vdd.n3122 vdd.n460 19.3944
R19865 vdd.n3117 vdd.n460 19.3944
R19866 vdd.n3117 vdd.n3116 19.3944
R19867 vdd.n3189 vdd.n386 19.3944
R19868 vdd.n3189 vdd.n392 19.3944
R19869 vdd.n3184 vdd.n392 19.3944
R19870 vdd.n3184 vdd.n3183 19.3944
R19871 vdd.n3183 vdd.n3182 19.3944
R19872 vdd.n3182 vdd.n399 19.3944
R19873 vdd.n3177 vdd.n399 19.3944
R19874 vdd.n3177 vdd.n3176 19.3944
R19875 vdd.n3176 vdd.n3175 19.3944
R19876 vdd.n3175 vdd.n406 19.3944
R19877 vdd.n3170 vdd.n406 19.3944
R19878 vdd.n3170 vdd.n3169 19.3944
R19879 vdd.n3169 vdd.n3168 19.3944
R19880 vdd.n3168 vdd.n413 19.3944
R19881 vdd.n3163 vdd.n413 19.3944
R19882 vdd.n3163 vdd.n3162 19.3944
R19883 vdd.n3162 vdd.n3161 19.3944
R19884 vdd.n3161 vdd.n420 19.3944
R19885 vdd.n3156 vdd.n420 19.3944
R19886 vdd.n3156 vdd.n3155 19.3944
R19887 vdd.n3225 vdd.n3224 19.3944
R19888 vdd.n3224 vdd.n3223 19.3944
R19889 vdd.n3223 vdd.n358 19.3944
R19890 vdd.n359 vdd.n358 19.3944
R19891 vdd.n3216 vdd.n359 19.3944
R19892 vdd.n3216 vdd.n3215 19.3944
R19893 vdd.n3215 vdd.n3214 19.3944
R19894 vdd.n3214 vdd.n366 19.3944
R19895 vdd.n3209 vdd.n366 19.3944
R19896 vdd.n3209 vdd.n3208 19.3944
R19897 vdd.n3208 vdd.n3207 19.3944
R19898 vdd.n3207 vdd.n373 19.3944
R19899 vdd.n3202 vdd.n373 19.3944
R19900 vdd.n3202 vdd.n3201 19.3944
R19901 vdd.n3201 vdd.n3200 19.3944
R19902 vdd.n3200 vdd.n380 19.3944
R19903 vdd.n3195 vdd.n380 19.3944
R19904 vdd.n3195 vdd.n3194 19.3944
R19905 vdd.n3030 vdd.n509 19.3944
R19906 vdd.n3042 vdd.n509 19.3944
R19907 vdd.n3042 vdd.n507 19.3944
R19908 vdd.n3046 vdd.n507 19.3944
R19909 vdd.n3046 vdd.n497 19.3944
R19910 vdd.n3058 vdd.n497 19.3944
R19911 vdd.n3058 vdd.n495 19.3944
R19912 vdd.n3062 vdd.n495 19.3944
R19913 vdd.n3062 vdd.n485 19.3944
R19914 vdd.n3075 vdd.n485 19.3944
R19915 vdd.n3075 vdd.n483 19.3944
R19916 vdd.n3079 vdd.n483 19.3944
R19917 vdd.n3079 vdd.n312 19.3944
R19918 vdd.n3258 vdd.n312 19.3944
R19919 vdd.n3258 vdd.n313 19.3944
R19920 vdd.n3252 vdd.n313 19.3944
R19921 vdd.n3252 vdd.n3251 19.3944
R19922 vdd.n3251 vdd.n3250 19.3944
R19923 vdd.n3250 vdd.n323 19.3944
R19924 vdd.n3244 vdd.n323 19.3944
R19925 vdd.n3244 vdd.n3243 19.3944
R19926 vdd.n3243 vdd.n3242 19.3944
R19927 vdd.n3242 vdd.n335 19.3944
R19928 vdd.n3236 vdd.n335 19.3944
R19929 vdd.n3236 vdd.n3235 19.3944
R19930 vdd.n3235 vdd.n3234 19.3944
R19931 vdd.n3234 vdd.n346 19.3944
R19932 vdd.n3228 vdd.n346 19.3944
R19933 vdd.n2987 vdd.n2986 19.3944
R19934 vdd.n2986 vdd.n2985 19.3944
R19935 vdd.n2985 vdd.n551 19.3944
R19936 vdd.n2979 vdd.n551 19.3944
R19937 vdd.n2979 vdd.n2978 19.3944
R19938 vdd.n2978 vdd.n2977 19.3944
R19939 vdd.n2977 vdd.n557 19.3944
R19940 vdd.n2971 vdd.n557 19.3944
R19941 vdd.n2971 vdd.n2970 19.3944
R19942 vdd.n2970 vdd.n2969 19.3944
R19943 vdd.n2969 vdd.n563 19.3944
R19944 vdd.n2963 vdd.n563 19.3944
R19945 vdd.n2963 vdd.n2962 19.3944
R19946 vdd.n2962 vdd.n2961 19.3944
R19947 vdd.n2961 vdd.n569 19.3944
R19948 vdd.n2955 vdd.n569 19.3944
R19949 vdd.n2955 vdd.n2954 19.3944
R19950 vdd.n2954 vdd.n2953 19.3944
R19951 vdd.n2953 vdd.n575 19.3944
R19952 vdd.n2947 vdd.n575 19.3944
R19953 vdd.n3027 vdd.n3026 19.3944
R19954 vdd.n3026 vdd.n519 19.3944
R19955 vdd.n3021 vdd.n3020 19.3944
R19956 vdd.n3017 vdd.n3016 19.3944
R19957 vdd.n3016 vdd.n525 19.3944
R19958 vdd.n3011 vdd.n525 19.3944
R19959 vdd.n3011 vdd.n3010 19.3944
R19960 vdd.n3010 vdd.n3009 19.3944
R19961 vdd.n3009 vdd.n531 19.3944
R19962 vdd.n3003 vdd.n531 19.3944
R19963 vdd.n3003 vdd.n3002 19.3944
R19964 vdd.n3002 vdd.n3001 19.3944
R19965 vdd.n3001 vdd.n537 19.3944
R19966 vdd.n2995 vdd.n537 19.3944
R19967 vdd.n2995 vdd.n2994 19.3944
R19968 vdd.n2994 vdd.n2993 19.3944
R19969 vdd.n2942 vdd.n579 19.3944
R19970 vdd.n2942 vdd.n583 19.3944
R19971 vdd.n2937 vdd.n583 19.3944
R19972 vdd.n2937 vdd.n2936 19.3944
R19973 vdd.n2936 vdd.n589 19.3944
R19974 vdd.n2931 vdd.n589 19.3944
R19975 vdd.n2931 vdd.n2930 19.3944
R19976 vdd.n2930 vdd.n2929 19.3944
R19977 vdd.n2929 vdd.n595 19.3944
R19978 vdd.n2923 vdd.n595 19.3944
R19979 vdd.n2923 vdd.n2922 19.3944
R19980 vdd.n2922 vdd.n2921 19.3944
R19981 vdd.n2921 vdd.n601 19.3944
R19982 vdd.n2915 vdd.n601 19.3944
R19983 vdd.n2915 vdd.n2914 19.3944
R19984 vdd.n2914 vdd.n2913 19.3944
R19985 vdd.n2909 vdd.n2908 19.3944
R19986 vdd.n2905 vdd.n2904 19.3944
R19987 vdd.n1511 vdd.n1430 19.0066
R19988 vdd.n2019 vdd.n1017 19.0066
R19989 vdd.n3154 vdd.n426 19.0066
R19990 vdd.n2946 vdd.n579 19.0066
R19991 vdd.n1082 vdd.n1081 16.0975
R19992 vdd.n810 vdd.n809 16.0975
R19993 vdd.n1473 vdd.n1472 16.0975
R19994 vdd.n1510 vdd.n1509 16.0975
R19995 vdd.n1384 vdd.n1383 16.0975
R19996 vdd.n1982 vdd.n1981 16.0975
R19997 vdd.n1019 vdd.n1018 16.0975
R19998 vdd.n979 vdd.n978 16.0975
R19999 vdd.n1102 vdd.n1101 16.0975
R20000 vdd.n801 vdd.n800 16.0975
R20001 vdd.n2417 vdd.n2416 16.0975
R20002 vdd.n3114 vdd.n3113 16.0975
R20003 vdd.n428 vdd.n427 16.0975
R20004 vdd.n388 vdd.n387 16.0975
R20005 vdd.n581 vdd.n580 16.0975
R20006 vdd.n544 vdd.n543 16.0975
R20007 vdd.n662 vdd.n661 16.0975
R20008 vdd.n2414 vdd.n2413 16.0975
R20009 vdd.n2901 vdd.n2900 16.0975
R20010 vdd.n626 vdd.n625 16.0975
R20011 vdd.t120 vdd.n2377 15.4182
R20012 vdd.n2650 vdd.t114 15.4182
R20013 vdd.n28 vdd.n27 14.8572
R20014 vdd.n2129 vdd.n904 14.0578
R20015 vdd.n2863 vdd.n613 14.0578
R20016 vdd.n304 vdd.n269 13.1884
R20017 vdd.n253 vdd.n218 13.1884
R20018 vdd.n210 vdd.n175 13.1884
R20019 vdd.n159 vdd.n124 13.1884
R20020 vdd.n117 vdd.n82 13.1884
R20021 vdd.n66 vdd.n31 13.1884
R20022 vdd.n1861 vdd.n1826 13.1884
R20023 vdd.n1912 vdd.n1877 13.1884
R20024 vdd.n1767 vdd.n1732 13.1884
R20025 vdd.n1818 vdd.n1783 13.1884
R20026 vdd.n1674 vdd.n1639 13.1884
R20027 vdd.n1725 vdd.n1690 13.1884
R20028 vdd.n1542 vdd.n1385 12.9944
R20029 vdd.n1546 vdd.n1385 12.9944
R20030 vdd.n2058 vdd.n977 12.9944
R20031 vdd.n2059 vdd.n2058 12.9944
R20032 vdd.n3193 vdd.n386 12.9944
R20033 vdd.n3194 vdd.n3193 12.9944
R20034 vdd.n2987 vdd.n545 12.9944
R20035 vdd.n2993 vdd.n545 12.9944
R20036 vdd.n305 vdd.n267 12.8005
R20037 vdd.n300 vdd.n271 12.8005
R20038 vdd.n254 vdd.n216 12.8005
R20039 vdd.n249 vdd.n220 12.8005
R20040 vdd.n211 vdd.n173 12.8005
R20041 vdd.n206 vdd.n177 12.8005
R20042 vdd.n160 vdd.n122 12.8005
R20043 vdd.n155 vdd.n126 12.8005
R20044 vdd.n118 vdd.n80 12.8005
R20045 vdd.n113 vdd.n84 12.8005
R20046 vdd.n67 vdd.n29 12.8005
R20047 vdd.n62 vdd.n33 12.8005
R20048 vdd.n1862 vdd.n1824 12.8005
R20049 vdd.n1857 vdd.n1828 12.8005
R20050 vdd.n1913 vdd.n1875 12.8005
R20051 vdd.n1908 vdd.n1879 12.8005
R20052 vdd.n1768 vdd.n1730 12.8005
R20053 vdd.n1763 vdd.n1734 12.8005
R20054 vdd.n1819 vdd.n1781 12.8005
R20055 vdd.n1814 vdd.n1785 12.8005
R20056 vdd.n1675 vdd.n1637 12.8005
R20057 vdd.n1670 vdd.n1641 12.8005
R20058 vdd.n1726 vdd.n1688 12.8005
R20059 vdd.n1721 vdd.n1692 12.8005
R20060 vdd.n299 vdd.n272 12.0247
R20061 vdd.n248 vdd.n221 12.0247
R20062 vdd.n205 vdd.n178 12.0247
R20063 vdd.n154 vdd.n127 12.0247
R20064 vdd.n112 vdd.n85 12.0247
R20065 vdd.n61 vdd.n34 12.0247
R20066 vdd.n1856 vdd.n1829 12.0247
R20067 vdd.n1907 vdd.n1880 12.0247
R20068 vdd.n1762 vdd.n1735 12.0247
R20069 vdd.n1813 vdd.n1786 12.0247
R20070 vdd.n1669 vdd.n1642 12.0247
R20071 vdd.n1720 vdd.n1693 12.0247
R20072 vdd.n1577 vdd.n1345 11.337
R20073 vdd.n1585 vdd.n1334 11.337
R20074 vdd.n1593 vdd.n1334 11.337
R20075 vdd.n1601 vdd.n1328 11.337
R20076 vdd.n1609 vdd.n1321 11.337
R20077 vdd.n1618 vdd.n1617 11.337
R20078 vdd.n1626 vdd.n1310 11.337
R20079 vdd.n1924 vdd.n1299 11.337
R20080 vdd.n1933 vdd.n1293 11.337
R20081 vdd.n1941 vdd.n1287 11.337
R20082 vdd.n1950 vdd.n1949 11.337
R20083 vdd.n1958 vdd.n1270 11.337
R20084 vdd.n1969 vdd.n1270 11.337
R20085 vdd.n1969 vdd.n1968 11.337
R20086 vdd.n3040 vdd.n511 11.337
R20087 vdd.n3040 vdd.n505 11.337
R20088 vdd.n3048 vdd.n505 11.337
R20089 vdd.n3056 vdd.n499 11.337
R20090 vdd.n3064 vdd.n492 11.337
R20091 vdd.n3073 vdd.n3072 11.337
R20092 vdd.n3081 vdd.n481 11.337
R20093 vdd.n3255 vdd.n3254 11.337
R20094 vdd.n3248 vdd.n325 11.337
R20095 vdd.n3246 vdd.n329 11.337
R20096 vdd.n3240 vdd.n3239 11.337
R20097 vdd.n3238 vdd.n340 11.337
R20098 vdd.n3232 vdd.n340 11.337
R20099 vdd.n3231 vdd.n3230 11.337
R20100 vdd.n296 vdd.n295 11.249
R20101 vdd.n245 vdd.n244 11.249
R20102 vdd.n202 vdd.n201 11.249
R20103 vdd.n151 vdd.n150 11.249
R20104 vdd.n109 vdd.n108 11.249
R20105 vdd.n58 vdd.n57 11.249
R20106 vdd.n1853 vdd.n1852 11.249
R20107 vdd.n1904 vdd.n1903 11.249
R20108 vdd.n1759 vdd.n1758 11.249
R20109 vdd.n1810 vdd.n1809 11.249
R20110 vdd.n1666 vdd.n1665 11.249
R20111 vdd.n1717 vdd.n1716 11.249
R20112 vdd.n1593 vdd.t140 10.9969
R20113 vdd.t151 vdd.n3238 10.9969
R20114 vdd.n1322 vdd.t156 10.7702
R20115 vdd.t187 vdd.n3247 10.7702
R20116 vdd.n281 vdd.n280 10.7238
R20117 vdd.n230 vdd.n229 10.7238
R20118 vdd.n187 vdd.n186 10.7238
R20119 vdd.n136 vdd.n135 10.7238
R20120 vdd.n94 vdd.n93 10.7238
R20121 vdd.n43 vdd.n42 10.7238
R20122 vdd.n1838 vdd.n1837 10.7238
R20123 vdd.n1889 vdd.n1888 10.7238
R20124 vdd.n1744 vdd.n1743 10.7238
R20125 vdd.n1795 vdd.n1794 10.7238
R20126 vdd.n1651 vdd.n1650 10.7238
R20127 vdd.n1702 vdd.n1701 10.7238
R20128 vdd.n2305 vdd.t99 10.6568
R20129 vdd.t129 vdd.n756 10.6568
R20130 vdd.n2138 vdd.n902 10.6151
R20131 vdd.n2139 vdd.n2138 10.6151
R20132 vdd.n2140 vdd.n2139 10.6151
R20133 vdd.n2140 vdd.n891 10.6151
R20134 vdd.n2150 vdd.n891 10.6151
R20135 vdd.n2151 vdd.n2150 10.6151
R20136 vdd.n2152 vdd.n2151 10.6151
R20137 vdd.n2152 vdd.n878 10.6151
R20138 vdd.n2162 vdd.n878 10.6151
R20139 vdd.n2163 vdd.n2162 10.6151
R20140 vdd.n2164 vdd.n2163 10.6151
R20141 vdd.n2164 vdd.n866 10.6151
R20142 vdd.n2175 vdd.n866 10.6151
R20143 vdd.n2176 vdd.n2175 10.6151
R20144 vdd.n2177 vdd.n2176 10.6151
R20145 vdd.n2177 vdd.n854 10.6151
R20146 vdd.n2187 vdd.n854 10.6151
R20147 vdd.n2188 vdd.n2187 10.6151
R20148 vdd.n2189 vdd.n2188 10.6151
R20149 vdd.n2189 vdd.n842 10.6151
R20150 vdd.n2199 vdd.n842 10.6151
R20151 vdd.n2200 vdd.n2199 10.6151
R20152 vdd.n2201 vdd.n2200 10.6151
R20153 vdd.n2201 vdd.n831 10.6151
R20154 vdd.n2211 vdd.n831 10.6151
R20155 vdd.n2212 vdd.n2211 10.6151
R20156 vdd.n2213 vdd.n2212 10.6151
R20157 vdd.n2213 vdd.n818 10.6151
R20158 vdd.n2225 vdd.n818 10.6151
R20159 vdd.n2226 vdd.n2225 10.6151
R20160 vdd.n2228 vdd.n2226 10.6151
R20161 vdd.n2228 vdd.n2227 10.6151
R20162 vdd.n2227 vdd.n799 10.6151
R20163 vdd.n2375 vdd.n2374 10.6151
R20164 vdd.n2374 vdd.n2373 10.6151
R20165 vdd.n2373 vdd.n2370 10.6151
R20166 vdd.n2370 vdd.n2369 10.6151
R20167 vdd.n2369 vdd.n2366 10.6151
R20168 vdd.n2366 vdd.n2365 10.6151
R20169 vdd.n2365 vdd.n2362 10.6151
R20170 vdd.n2362 vdd.n2361 10.6151
R20171 vdd.n2361 vdd.n2358 10.6151
R20172 vdd.n2358 vdd.n2357 10.6151
R20173 vdd.n2357 vdd.n2354 10.6151
R20174 vdd.n2354 vdd.n2353 10.6151
R20175 vdd.n2353 vdd.n2350 10.6151
R20176 vdd.n2350 vdd.n2349 10.6151
R20177 vdd.n2349 vdd.n2346 10.6151
R20178 vdd.n2346 vdd.n2345 10.6151
R20179 vdd.n2345 vdd.n2342 10.6151
R20180 vdd.n2342 vdd.n2341 10.6151
R20181 vdd.n2341 vdd.n2338 10.6151
R20182 vdd.n2338 vdd.n2337 10.6151
R20183 vdd.n2337 vdd.n2334 10.6151
R20184 vdd.n2334 vdd.n2333 10.6151
R20185 vdd.n2333 vdd.n2330 10.6151
R20186 vdd.n2330 vdd.n2329 10.6151
R20187 vdd.n2329 vdd.n2326 10.6151
R20188 vdd.n2326 vdd.n2325 10.6151
R20189 vdd.n2325 vdd.n2322 10.6151
R20190 vdd.n2322 vdd.n2321 10.6151
R20191 vdd.n2321 vdd.n2318 10.6151
R20192 vdd.n2318 vdd.n2317 10.6151
R20193 vdd.n2317 vdd.n2314 10.6151
R20194 vdd.n2312 vdd.n2309 10.6151
R20195 vdd.n2309 vdd.n2308 10.6151
R20196 vdd.n1139 vdd.n1138 10.6151
R20197 vdd.n1141 vdd.n1139 10.6151
R20198 vdd.n1142 vdd.n1141 10.6151
R20199 vdd.n1144 vdd.n1142 10.6151
R20200 vdd.n1145 vdd.n1144 10.6151
R20201 vdd.n1147 vdd.n1145 10.6151
R20202 vdd.n1148 vdd.n1147 10.6151
R20203 vdd.n1150 vdd.n1148 10.6151
R20204 vdd.n1151 vdd.n1150 10.6151
R20205 vdd.n1153 vdd.n1151 10.6151
R20206 vdd.n1154 vdd.n1153 10.6151
R20207 vdd.n1156 vdd.n1154 10.6151
R20208 vdd.n1157 vdd.n1156 10.6151
R20209 vdd.n1159 vdd.n1157 10.6151
R20210 vdd.n1160 vdd.n1159 10.6151
R20211 vdd.n1162 vdd.n1160 10.6151
R20212 vdd.n1163 vdd.n1162 10.6151
R20213 vdd.n1185 vdd.n1163 10.6151
R20214 vdd.n1185 vdd.n1184 10.6151
R20215 vdd.n1184 vdd.n1183 10.6151
R20216 vdd.n1183 vdd.n1181 10.6151
R20217 vdd.n1181 vdd.n1180 10.6151
R20218 vdd.n1180 vdd.n1178 10.6151
R20219 vdd.n1178 vdd.n1177 10.6151
R20220 vdd.n1177 vdd.n1175 10.6151
R20221 vdd.n1175 vdd.n1174 10.6151
R20222 vdd.n1174 vdd.n1172 10.6151
R20223 vdd.n1172 vdd.n1171 10.6151
R20224 vdd.n1171 vdd.n1169 10.6151
R20225 vdd.n1169 vdd.n1168 10.6151
R20226 vdd.n1168 vdd.n1165 10.6151
R20227 vdd.n1165 vdd.n1164 10.6151
R20228 vdd.n1164 vdd.n802 10.6151
R20229 vdd.n2126 vdd.n2125 10.6151
R20230 vdd.n2125 vdd.n2124 10.6151
R20231 vdd.n2124 vdd.n2123 10.6151
R20232 vdd.n2123 vdd.n2121 10.6151
R20233 vdd.n2121 vdd.n2118 10.6151
R20234 vdd.n2118 vdd.n2117 10.6151
R20235 vdd.n2117 vdd.n2114 10.6151
R20236 vdd.n2114 vdd.n2113 10.6151
R20237 vdd.n2113 vdd.n2110 10.6151
R20238 vdd.n2110 vdd.n2109 10.6151
R20239 vdd.n2109 vdd.n2106 10.6151
R20240 vdd.n2106 vdd.n2105 10.6151
R20241 vdd.n2105 vdd.n2102 10.6151
R20242 vdd.n2102 vdd.n2101 10.6151
R20243 vdd.n2101 vdd.n2098 10.6151
R20244 vdd.n2098 vdd.n2097 10.6151
R20245 vdd.n2097 vdd.n2094 10.6151
R20246 vdd.n2094 vdd.n947 10.6151
R20247 vdd.n1105 vdd.n947 10.6151
R20248 vdd.n1106 vdd.n1105 10.6151
R20249 vdd.n1109 vdd.n1106 10.6151
R20250 vdd.n1110 vdd.n1109 10.6151
R20251 vdd.n1113 vdd.n1110 10.6151
R20252 vdd.n1114 vdd.n1113 10.6151
R20253 vdd.n1117 vdd.n1114 10.6151
R20254 vdd.n1118 vdd.n1117 10.6151
R20255 vdd.n1121 vdd.n1118 10.6151
R20256 vdd.n1122 vdd.n1121 10.6151
R20257 vdd.n1125 vdd.n1122 10.6151
R20258 vdd.n1126 vdd.n1125 10.6151
R20259 vdd.n1129 vdd.n1126 10.6151
R20260 vdd.n1134 vdd.n1131 10.6151
R20261 vdd.n1135 vdd.n1134 10.6151
R20262 vdd.n2578 vdd.n2577 10.6151
R20263 vdd.n2577 vdd.n2576 10.6151
R20264 vdd.n2576 vdd.n2415 10.6151
R20265 vdd.n2520 vdd.n2415 10.6151
R20266 vdd.n2521 vdd.n2520 10.6151
R20267 vdd.n2523 vdd.n2521 10.6151
R20268 vdd.n2524 vdd.n2523 10.6151
R20269 vdd.n2526 vdd.n2524 10.6151
R20270 vdd.n2527 vdd.n2526 10.6151
R20271 vdd.n2557 vdd.n2527 10.6151
R20272 vdd.n2557 vdd.n2556 10.6151
R20273 vdd.n2556 vdd.n2555 10.6151
R20274 vdd.n2555 vdd.n2553 10.6151
R20275 vdd.n2553 vdd.n2552 10.6151
R20276 vdd.n2552 vdd.n2550 10.6151
R20277 vdd.n2550 vdd.n2549 10.6151
R20278 vdd.n2549 vdd.n2547 10.6151
R20279 vdd.n2547 vdd.n2546 10.6151
R20280 vdd.n2546 vdd.n2544 10.6151
R20281 vdd.n2544 vdd.n2543 10.6151
R20282 vdd.n2543 vdd.n2541 10.6151
R20283 vdd.n2541 vdd.n2540 10.6151
R20284 vdd.n2540 vdd.n2538 10.6151
R20285 vdd.n2538 vdd.n2537 10.6151
R20286 vdd.n2537 vdd.n2535 10.6151
R20287 vdd.n2535 vdd.n2534 10.6151
R20288 vdd.n2534 vdd.n2532 10.6151
R20289 vdd.n2532 vdd.n2531 10.6151
R20290 vdd.n2531 vdd.n2529 10.6151
R20291 vdd.n2529 vdd.n2528 10.6151
R20292 vdd.n2528 vdd.n664 10.6151
R20293 vdd.n2796 vdd.n664 10.6151
R20294 vdd.n2797 vdd.n2796 10.6151
R20295 vdd.n2647 vdd.n2646 10.6151
R20296 vdd.n2646 vdd.n2645 10.6151
R20297 vdd.n2645 vdd.n2644 10.6151
R20298 vdd.n2644 vdd.n2642 10.6151
R20299 vdd.n2642 vdd.n2639 10.6151
R20300 vdd.n2639 vdd.n2638 10.6151
R20301 vdd.n2638 vdd.n2635 10.6151
R20302 vdd.n2635 vdd.n2634 10.6151
R20303 vdd.n2634 vdd.n2631 10.6151
R20304 vdd.n2631 vdd.n2630 10.6151
R20305 vdd.n2630 vdd.n2627 10.6151
R20306 vdd.n2627 vdd.n2626 10.6151
R20307 vdd.n2626 vdd.n2623 10.6151
R20308 vdd.n2623 vdd.n2622 10.6151
R20309 vdd.n2622 vdd.n2619 10.6151
R20310 vdd.n2619 vdd.n2618 10.6151
R20311 vdd.n2618 vdd.n2615 10.6151
R20312 vdd.n2615 vdd.n2614 10.6151
R20313 vdd.n2614 vdd.n2611 10.6151
R20314 vdd.n2611 vdd.n2610 10.6151
R20315 vdd.n2610 vdd.n2607 10.6151
R20316 vdd.n2607 vdd.n2606 10.6151
R20317 vdd.n2606 vdd.n2603 10.6151
R20318 vdd.n2603 vdd.n2602 10.6151
R20319 vdd.n2602 vdd.n2599 10.6151
R20320 vdd.n2599 vdd.n2598 10.6151
R20321 vdd.n2598 vdd.n2595 10.6151
R20322 vdd.n2595 vdd.n2594 10.6151
R20323 vdd.n2594 vdd.n2591 10.6151
R20324 vdd.n2591 vdd.n2590 10.6151
R20325 vdd.n2590 vdd.n2587 10.6151
R20326 vdd.n2585 vdd.n2582 10.6151
R20327 vdd.n2582 vdd.n2581 10.6151
R20328 vdd.n2659 vdd.n754 10.6151
R20329 vdd.n2660 vdd.n2659 10.6151
R20330 vdd.n2661 vdd.n2660 10.6151
R20331 vdd.n2661 vdd.n743 10.6151
R20332 vdd.n2671 vdd.n743 10.6151
R20333 vdd.n2672 vdd.n2671 10.6151
R20334 vdd.n2673 vdd.n2672 10.6151
R20335 vdd.n2673 vdd.n731 10.6151
R20336 vdd.n2683 vdd.n731 10.6151
R20337 vdd.n2684 vdd.n2683 10.6151
R20338 vdd.n2685 vdd.n2684 10.6151
R20339 vdd.n2685 vdd.n719 10.6151
R20340 vdd.n2695 vdd.n719 10.6151
R20341 vdd.n2696 vdd.n2695 10.6151
R20342 vdd.n2697 vdd.n2696 10.6151
R20343 vdd.n2697 vdd.n708 10.6151
R20344 vdd.n2707 vdd.n708 10.6151
R20345 vdd.n2708 vdd.n2707 10.6151
R20346 vdd.n2709 vdd.n2708 10.6151
R20347 vdd.n2709 vdd.n694 10.6151
R20348 vdd.n2720 vdd.n694 10.6151
R20349 vdd.n2721 vdd.n2720 10.6151
R20350 vdd.n2722 vdd.n2721 10.6151
R20351 vdd.n2722 vdd.n683 10.6151
R20352 vdd.n2732 vdd.n683 10.6151
R20353 vdd.n2733 vdd.n2732 10.6151
R20354 vdd.n2734 vdd.n2733 10.6151
R20355 vdd.n2734 vdd.n669 10.6151
R20356 vdd.n2789 vdd.n669 10.6151
R20357 vdd.n2790 vdd.n2789 10.6151
R20358 vdd.n2791 vdd.n2790 10.6151
R20359 vdd.n2791 vdd.n636 10.6151
R20360 vdd.n2861 vdd.n636 10.6151
R20361 vdd.n2860 vdd.n2859 10.6151
R20362 vdd.n2859 vdd.n637 10.6151
R20363 vdd.n638 vdd.n637 10.6151
R20364 vdd.n2852 vdd.n638 10.6151
R20365 vdd.n2852 vdd.n2851 10.6151
R20366 vdd.n2851 vdd.n2850 10.6151
R20367 vdd.n2850 vdd.n640 10.6151
R20368 vdd.n2845 vdd.n640 10.6151
R20369 vdd.n2845 vdd.n2844 10.6151
R20370 vdd.n2844 vdd.n2843 10.6151
R20371 vdd.n2843 vdd.n643 10.6151
R20372 vdd.n2838 vdd.n643 10.6151
R20373 vdd.n2838 vdd.n2837 10.6151
R20374 vdd.n2837 vdd.n2836 10.6151
R20375 vdd.n2836 vdd.n646 10.6151
R20376 vdd.n2831 vdd.n646 10.6151
R20377 vdd.n2831 vdd.n2830 10.6151
R20378 vdd.n2830 vdd.n2828 10.6151
R20379 vdd.n2828 vdd.n649 10.6151
R20380 vdd.n2823 vdd.n649 10.6151
R20381 vdd.n2823 vdd.n2822 10.6151
R20382 vdd.n2822 vdd.n2821 10.6151
R20383 vdd.n2821 vdd.n652 10.6151
R20384 vdd.n2816 vdd.n652 10.6151
R20385 vdd.n2816 vdd.n2815 10.6151
R20386 vdd.n2815 vdd.n2814 10.6151
R20387 vdd.n2814 vdd.n655 10.6151
R20388 vdd.n2809 vdd.n655 10.6151
R20389 vdd.n2809 vdd.n2808 10.6151
R20390 vdd.n2808 vdd.n2807 10.6151
R20391 vdd.n2807 vdd.n658 10.6151
R20392 vdd.n2802 vdd.n2801 10.6151
R20393 vdd.n2801 vdd.n2800 10.6151
R20394 vdd.n2779 vdd.n2740 10.6151
R20395 vdd.n2774 vdd.n2740 10.6151
R20396 vdd.n2774 vdd.n2773 10.6151
R20397 vdd.n2773 vdd.n2772 10.6151
R20398 vdd.n2772 vdd.n2742 10.6151
R20399 vdd.n2767 vdd.n2742 10.6151
R20400 vdd.n2767 vdd.n2766 10.6151
R20401 vdd.n2766 vdd.n2765 10.6151
R20402 vdd.n2765 vdd.n2745 10.6151
R20403 vdd.n2760 vdd.n2745 10.6151
R20404 vdd.n2760 vdd.n2759 10.6151
R20405 vdd.n2759 vdd.n2758 10.6151
R20406 vdd.n2758 vdd.n2748 10.6151
R20407 vdd.n2753 vdd.n2748 10.6151
R20408 vdd.n2753 vdd.n2752 10.6151
R20409 vdd.n2752 vdd.n610 10.6151
R20410 vdd.n2896 vdd.n610 10.6151
R20411 vdd.n2896 vdd.n611 10.6151
R20412 vdd.n614 vdd.n611 10.6151
R20413 vdd.n2889 vdd.n614 10.6151
R20414 vdd.n2889 vdd.n2888 10.6151
R20415 vdd.n2888 vdd.n2887 10.6151
R20416 vdd.n2887 vdd.n616 10.6151
R20417 vdd.n2882 vdd.n616 10.6151
R20418 vdd.n2882 vdd.n2881 10.6151
R20419 vdd.n2881 vdd.n2880 10.6151
R20420 vdd.n2880 vdd.n619 10.6151
R20421 vdd.n2875 vdd.n619 10.6151
R20422 vdd.n2875 vdd.n2874 10.6151
R20423 vdd.n2874 vdd.n2873 10.6151
R20424 vdd.n2873 vdd.n622 10.6151
R20425 vdd.n2868 vdd.n2867 10.6151
R20426 vdd.n2867 vdd.n2866 10.6151
R20427 vdd.n2486 vdd.n2485 10.6151
R20428 vdd.n2572 vdd.n2486 10.6151
R20429 vdd.n2572 vdd.n2571 10.6151
R20430 vdd.n2571 vdd.n2570 10.6151
R20431 vdd.n2570 vdd.n2568 10.6151
R20432 vdd.n2568 vdd.n2567 10.6151
R20433 vdd.n2567 vdd.n2565 10.6151
R20434 vdd.n2565 vdd.n2564 10.6151
R20435 vdd.n2564 vdd.n2562 10.6151
R20436 vdd.n2562 vdd.n2561 10.6151
R20437 vdd.n2561 vdd.n2518 10.6151
R20438 vdd.n2518 vdd.n2517 10.6151
R20439 vdd.n2517 vdd.n2515 10.6151
R20440 vdd.n2515 vdd.n2514 10.6151
R20441 vdd.n2514 vdd.n2512 10.6151
R20442 vdd.n2512 vdd.n2511 10.6151
R20443 vdd.n2511 vdd.n2509 10.6151
R20444 vdd.n2509 vdd.n2508 10.6151
R20445 vdd.n2508 vdd.n2506 10.6151
R20446 vdd.n2506 vdd.n2505 10.6151
R20447 vdd.n2505 vdd.n2503 10.6151
R20448 vdd.n2503 vdd.n2502 10.6151
R20449 vdd.n2502 vdd.n2500 10.6151
R20450 vdd.n2500 vdd.n2499 10.6151
R20451 vdd.n2499 vdd.n2497 10.6151
R20452 vdd.n2497 vdd.n2496 10.6151
R20453 vdd.n2496 vdd.n2494 10.6151
R20454 vdd.n2494 vdd.n2493 10.6151
R20455 vdd.n2493 vdd.n2491 10.6151
R20456 vdd.n2491 vdd.n2490 10.6151
R20457 vdd.n2490 vdd.n2488 10.6151
R20458 vdd.n2488 vdd.n2487 10.6151
R20459 vdd.n2487 vdd.n628 10.6151
R20460 vdd.n2653 vdd.n760 10.6151
R20461 vdd.n2420 vdd.n760 10.6151
R20462 vdd.n2421 vdd.n2420 10.6151
R20463 vdd.n2424 vdd.n2421 10.6151
R20464 vdd.n2425 vdd.n2424 10.6151
R20465 vdd.n2428 vdd.n2425 10.6151
R20466 vdd.n2429 vdd.n2428 10.6151
R20467 vdd.n2432 vdd.n2429 10.6151
R20468 vdd.n2433 vdd.n2432 10.6151
R20469 vdd.n2436 vdd.n2433 10.6151
R20470 vdd.n2437 vdd.n2436 10.6151
R20471 vdd.n2440 vdd.n2437 10.6151
R20472 vdd.n2441 vdd.n2440 10.6151
R20473 vdd.n2444 vdd.n2441 10.6151
R20474 vdd.n2445 vdd.n2444 10.6151
R20475 vdd.n2448 vdd.n2445 10.6151
R20476 vdd.n2449 vdd.n2448 10.6151
R20477 vdd.n2452 vdd.n2449 10.6151
R20478 vdd.n2453 vdd.n2452 10.6151
R20479 vdd.n2456 vdd.n2453 10.6151
R20480 vdd.n2457 vdd.n2456 10.6151
R20481 vdd.n2460 vdd.n2457 10.6151
R20482 vdd.n2461 vdd.n2460 10.6151
R20483 vdd.n2464 vdd.n2461 10.6151
R20484 vdd.n2465 vdd.n2464 10.6151
R20485 vdd.n2468 vdd.n2465 10.6151
R20486 vdd.n2469 vdd.n2468 10.6151
R20487 vdd.n2472 vdd.n2469 10.6151
R20488 vdd.n2473 vdd.n2472 10.6151
R20489 vdd.n2476 vdd.n2473 10.6151
R20490 vdd.n2477 vdd.n2476 10.6151
R20491 vdd.n2482 vdd.n2480 10.6151
R20492 vdd.n2483 vdd.n2482 10.6151
R20493 vdd.n2655 vdd.n2654 10.6151
R20494 vdd.n2655 vdd.n749 10.6151
R20495 vdd.n2665 vdd.n749 10.6151
R20496 vdd.n2666 vdd.n2665 10.6151
R20497 vdd.n2667 vdd.n2666 10.6151
R20498 vdd.n2667 vdd.n737 10.6151
R20499 vdd.n2677 vdd.n737 10.6151
R20500 vdd.n2678 vdd.n2677 10.6151
R20501 vdd.n2679 vdd.n2678 10.6151
R20502 vdd.n2679 vdd.n725 10.6151
R20503 vdd.n2689 vdd.n725 10.6151
R20504 vdd.n2690 vdd.n2689 10.6151
R20505 vdd.n2691 vdd.n2690 10.6151
R20506 vdd.n2691 vdd.n714 10.6151
R20507 vdd.n2701 vdd.n714 10.6151
R20508 vdd.n2702 vdd.n2701 10.6151
R20509 vdd.n2703 vdd.n2702 10.6151
R20510 vdd.n2703 vdd.n701 10.6151
R20511 vdd.n2713 vdd.n701 10.6151
R20512 vdd.n2714 vdd.n2713 10.6151
R20513 vdd.n2716 vdd.n689 10.6151
R20514 vdd.n2726 vdd.n689 10.6151
R20515 vdd.n2727 vdd.n2726 10.6151
R20516 vdd.n2728 vdd.n2727 10.6151
R20517 vdd.n2728 vdd.n677 10.6151
R20518 vdd.n2738 vdd.n677 10.6151
R20519 vdd.n2739 vdd.n2738 10.6151
R20520 vdd.n2785 vdd.n2739 10.6151
R20521 vdd.n2785 vdd.n2784 10.6151
R20522 vdd.n2784 vdd.n2783 10.6151
R20523 vdd.n2783 vdd.n2782 10.6151
R20524 vdd.n2782 vdd.n2780 10.6151
R20525 vdd.n2134 vdd.n2133 10.6151
R20526 vdd.n2134 vdd.n897 10.6151
R20527 vdd.n2144 vdd.n897 10.6151
R20528 vdd.n2145 vdd.n2144 10.6151
R20529 vdd.n2146 vdd.n2145 10.6151
R20530 vdd.n2146 vdd.n885 10.6151
R20531 vdd.n2156 vdd.n885 10.6151
R20532 vdd.n2157 vdd.n2156 10.6151
R20533 vdd.n2158 vdd.n2157 10.6151
R20534 vdd.n2158 vdd.n872 10.6151
R20535 vdd.n2168 vdd.n872 10.6151
R20536 vdd.n2169 vdd.n2168 10.6151
R20537 vdd.n2171 vdd.n860 10.6151
R20538 vdd.n2181 vdd.n860 10.6151
R20539 vdd.n2182 vdd.n2181 10.6151
R20540 vdd.n2183 vdd.n2182 10.6151
R20541 vdd.n2183 vdd.n848 10.6151
R20542 vdd.n2193 vdd.n848 10.6151
R20543 vdd.n2194 vdd.n2193 10.6151
R20544 vdd.n2195 vdd.n2194 10.6151
R20545 vdd.n2195 vdd.n837 10.6151
R20546 vdd.n2205 vdd.n837 10.6151
R20547 vdd.n2206 vdd.n2205 10.6151
R20548 vdd.n2207 vdd.n2206 10.6151
R20549 vdd.n2207 vdd.n825 10.6151
R20550 vdd.n2217 vdd.n825 10.6151
R20551 vdd.n2218 vdd.n2217 10.6151
R20552 vdd.n2221 vdd.n2218 10.6151
R20553 vdd.n2221 vdd.n2220 10.6151
R20554 vdd.n2220 vdd.n2219 10.6151
R20555 vdd.n2219 vdd.n808 10.6151
R20556 vdd.n2303 vdd.n808 10.6151
R20557 vdd.n2302 vdd.n2301 10.6151
R20558 vdd.n2301 vdd.n2298 10.6151
R20559 vdd.n2298 vdd.n2297 10.6151
R20560 vdd.n2297 vdd.n2294 10.6151
R20561 vdd.n2294 vdd.n2293 10.6151
R20562 vdd.n2293 vdd.n2290 10.6151
R20563 vdd.n2290 vdd.n2289 10.6151
R20564 vdd.n2289 vdd.n2286 10.6151
R20565 vdd.n2286 vdd.n2285 10.6151
R20566 vdd.n2285 vdd.n2282 10.6151
R20567 vdd.n2282 vdd.n2281 10.6151
R20568 vdd.n2281 vdd.n2278 10.6151
R20569 vdd.n2278 vdd.n2277 10.6151
R20570 vdd.n2277 vdd.n2274 10.6151
R20571 vdd.n2274 vdd.n2273 10.6151
R20572 vdd.n2273 vdd.n2270 10.6151
R20573 vdd.n2270 vdd.n2269 10.6151
R20574 vdd.n2269 vdd.n2266 10.6151
R20575 vdd.n2266 vdd.n2265 10.6151
R20576 vdd.n2265 vdd.n2262 10.6151
R20577 vdd.n2262 vdd.n2261 10.6151
R20578 vdd.n2261 vdd.n2258 10.6151
R20579 vdd.n2258 vdd.n2257 10.6151
R20580 vdd.n2257 vdd.n2254 10.6151
R20581 vdd.n2254 vdd.n2253 10.6151
R20582 vdd.n2253 vdd.n2250 10.6151
R20583 vdd.n2250 vdd.n2249 10.6151
R20584 vdd.n2249 vdd.n2246 10.6151
R20585 vdd.n2246 vdd.n2245 10.6151
R20586 vdd.n2245 vdd.n2242 10.6151
R20587 vdd.n2242 vdd.n2241 10.6151
R20588 vdd.n2238 vdd.n2237 10.6151
R20589 vdd.n2237 vdd.n2235 10.6151
R20590 vdd.n1216 vdd.n1214 10.6151
R20591 vdd.n1214 vdd.n1213 10.6151
R20592 vdd.n1213 vdd.n1211 10.6151
R20593 vdd.n1211 vdd.n1210 10.6151
R20594 vdd.n1210 vdd.n1208 10.6151
R20595 vdd.n1208 vdd.n1207 10.6151
R20596 vdd.n1207 vdd.n1205 10.6151
R20597 vdd.n1205 vdd.n1204 10.6151
R20598 vdd.n1204 vdd.n1202 10.6151
R20599 vdd.n1202 vdd.n1201 10.6151
R20600 vdd.n1201 vdd.n1199 10.6151
R20601 vdd.n1199 vdd.n1198 10.6151
R20602 vdd.n1198 vdd.n1196 10.6151
R20603 vdd.n1196 vdd.n1195 10.6151
R20604 vdd.n1195 vdd.n1193 10.6151
R20605 vdd.n1193 vdd.n1192 10.6151
R20606 vdd.n1192 vdd.n1190 10.6151
R20607 vdd.n1190 vdd.n1189 10.6151
R20608 vdd.n1189 vdd.n1100 10.6151
R20609 vdd.n1100 vdd.n1099 10.6151
R20610 vdd.n1099 vdd.n1097 10.6151
R20611 vdd.n1097 vdd.n1096 10.6151
R20612 vdd.n1096 vdd.n1094 10.6151
R20613 vdd.n1094 vdd.n1093 10.6151
R20614 vdd.n1093 vdd.n1091 10.6151
R20615 vdd.n1091 vdd.n1090 10.6151
R20616 vdd.n1090 vdd.n1088 10.6151
R20617 vdd.n1088 vdd.n1087 10.6151
R20618 vdd.n1087 vdd.n1085 10.6151
R20619 vdd.n1085 vdd.n1084 10.6151
R20620 vdd.n1084 vdd.n812 10.6151
R20621 vdd.n2233 vdd.n812 10.6151
R20622 vdd.n2234 vdd.n2233 10.6151
R20623 vdd.n2132 vdd.n909 10.6151
R20624 vdd.n1051 vdd.n909 10.6151
R20625 vdd.n1052 vdd.n1051 10.6151
R20626 vdd.n1055 vdd.n1052 10.6151
R20627 vdd.n1056 vdd.n1055 10.6151
R20628 vdd.n1059 vdd.n1056 10.6151
R20629 vdd.n1060 vdd.n1059 10.6151
R20630 vdd.n1063 vdd.n1060 10.6151
R20631 vdd.n1064 vdd.n1063 10.6151
R20632 vdd.n1067 vdd.n1064 10.6151
R20633 vdd.n1068 vdd.n1067 10.6151
R20634 vdd.n1071 vdd.n1068 10.6151
R20635 vdd.n1072 vdd.n1071 10.6151
R20636 vdd.n1075 vdd.n1072 10.6151
R20637 vdd.n1076 vdd.n1075 10.6151
R20638 vdd.n1079 vdd.n1076 10.6151
R20639 vdd.n1250 vdd.n1079 10.6151
R20640 vdd.n1250 vdd.n1249 10.6151
R20641 vdd.n1249 vdd.n1247 10.6151
R20642 vdd.n1247 vdd.n1244 10.6151
R20643 vdd.n1244 vdd.n1243 10.6151
R20644 vdd.n1243 vdd.n1240 10.6151
R20645 vdd.n1240 vdd.n1239 10.6151
R20646 vdd.n1239 vdd.n1236 10.6151
R20647 vdd.n1236 vdd.n1235 10.6151
R20648 vdd.n1235 vdd.n1232 10.6151
R20649 vdd.n1232 vdd.n1231 10.6151
R20650 vdd.n1231 vdd.n1228 10.6151
R20651 vdd.n1228 vdd.n1227 10.6151
R20652 vdd.n1227 vdd.n1224 10.6151
R20653 vdd.n1224 vdd.n1223 10.6151
R20654 vdd.n1220 vdd.n1219 10.6151
R20655 vdd.n1219 vdd.n1217 10.6151
R20656 vdd.n1634 vdd.t142 10.5435
R20657 vdd.n1977 vdd.t17 10.5435
R20658 vdd.n3032 vdd.t13 10.5435
R20659 vdd.n3256 vdd.t138 10.5435
R20660 vdd.n292 vdd.n274 10.4732
R20661 vdd.n241 vdd.n223 10.4732
R20662 vdd.n198 vdd.n180 10.4732
R20663 vdd.n147 vdd.n129 10.4732
R20664 vdd.n105 vdd.n87 10.4732
R20665 vdd.n54 vdd.n36 10.4732
R20666 vdd.n1849 vdd.n1831 10.4732
R20667 vdd.n1900 vdd.n1882 10.4732
R20668 vdd.n1755 vdd.n1737 10.4732
R20669 vdd.n1806 vdd.n1788 10.4732
R20670 vdd.n1662 vdd.n1644 10.4732
R20671 vdd.n1713 vdd.n1695 10.4732
R20672 vdd.n1932 vdd.t181 10.3167
R20673 vdd.t134 vdd.n493 10.3167
R20674 vdd.n1585 vdd.t25 9.86327
R20675 vdd.n3232 vdd.t21 9.86327
R20676 vdd.n2094 vdd.n2093 9.78206
R20677 vdd.n2830 vdd.n2829 9.78206
R20678 vdd.n2897 vdd.n2896 9.78206
R20679 vdd.n1986 vdd.n1250 9.78206
R20680 vdd.n291 vdd.n276 9.69747
R20681 vdd.n240 vdd.n225 9.69747
R20682 vdd.n197 vdd.n182 9.69747
R20683 vdd.n146 vdd.n131 9.69747
R20684 vdd.n104 vdd.n89 9.69747
R20685 vdd.n53 vdd.n38 9.69747
R20686 vdd.n1848 vdd.n1833 9.69747
R20687 vdd.n1899 vdd.n1884 9.69747
R20688 vdd.n1754 vdd.n1739 9.69747
R20689 vdd.n1805 vdd.n1790 9.69747
R20690 vdd.n1661 vdd.n1646 9.69747
R20691 vdd.n1712 vdd.n1697 9.69747
R20692 vdd.n307 vdd.n306 9.45567
R20693 vdd.n256 vdd.n255 9.45567
R20694 vdd.n213 vdd.n212 9.45567
R20695 vdd.n162 vdd.n161 9.45567
R20696 vdd.n120 vdd.n119 9.45567
R20697 vdd.n69 vdd.n68 9.45567
R20698 vdd.n1864 vdd.n1863 9.45567
R20699 vdd.n1915 vdd.n1914 9.45567
R20700 vdd.n1770 vdd.n1769 9.45567
R20701 vdd.n1821 vdd.n1820 9.45567
R20702 vdd.n1677 vdd.n1676 9.45567
R20703 vdd.n1728 vdd.n1727 9.45567
R20704 vdd.n2056 vdd.n977 9.3005
R20705 vdd.n2055 vdd.n2054 9.3005
R20706 vdd.n983 vdd.n982 9.3005
R20707 vdd.n2049 vdd.n987 9.3005
R20708 vdd.n2048 vdd.n988 9.3005
R20709 vdd.n2047 vdd.n989 9.3005
R20710 vdd.n993 vdd.n990 9.3005
R20711 vdd.n2042 vdd.n994 9.3005
R20712 vdd.n2041 vdd.n995 9.3005
R20713 vdd.n2040 vdd.n996 9.3005
R20714 vdd.n1000 vdd.n997 9.3005
R20715 vdd.n2035 vdd.n1001 9.3005
R20716 vdd.n2034 vdd.n1002 9.3005
R20717 vdd.n2033 vdd.n1003 9.3005
R20718 vdd.n1007 vdd.n1004 9.3005
R20719 vdd.n2028 vdd.n1008 9.3005
R20720 vdd.n2027 vdd.n1009 9.3005
R20721 vdd.n2026 vdd.n1010 9.3005
R20722 vdd.n1014 vdd.n1011 9.3005
R20723 vdd.n2021 vdd.n1015 9.3005
R20724 vdd.n2020 vdd.n1016 9.3005
R20725 vdd.n2019 vdd.n2018 9.3005
R20726 vdd.n2017 vdd.n1017 9.3005
R20727 vdd.n2016 vdd.n2015 9.3005
R20728 vdd.n1023 vdd.n1022 9.3005
R20729 vdd.n2010 vdd.n1027 9.3005
R20730 vdd.n2009 vdd.n1028 9.3005
R20731 vdd.n2008 vdd.n1029 9.3005
R20732 vdd.n1033 vdd.n1030 9.3005
R20733 vdd.n2003 vdd.n1034 9.3005
R20734 vdd.n2002 vdd.n1035 9.3005
R20735 vdd.n2001 vdd.n1036 9.3005
R20736 vdd.n1040 vdd.n1037 9.3005
R20737 vdd.n1996 vdd.n1041 9.3005
R20738 vdd.n1995 vdd.n1042 9.3005
R20739 vdd.n1994 vdd.n1043 9.3005
R20740 vdd.n1047 vdd.n1044 9.3005
R20741 vdd.n1989 vdd.n1048 9.3005
R20742 vdd.n2058 vdd.n2057 9.3005
R20743 vdd.n2080 vdd.n948 9.3005
R20744 vdd.n2079 vdd.n956 9.3005
R20745 vdd.n960 vdd.n957 9.3005
R20746 vdd.n2074 vdd.n961 9.3005
R20747 vdd.n2073 vdd.n962 9.3005
R20748 vdd.n2072 vdd.n963 9.3005
R20749 vdd.n967 vdd.n964 9.3005
R20750 vdd.n2067 vdd.n968 9.3005
R20751 vdd.n2066 vdd.n969 9.3005
R20752 vdd.n2065 vdd.n970 9.3005
R20753 vdd.n974 vdd.n971 9.3005
R20754 vdd.n2060 vdd.n975 9.3005
R20755 vdd.n2059 vdd.n976 9.3005
R20756 vdd.n2092 vdd.n2091 9.3005
R20757 vdd.n952 vdd.n951 9.3005
R20758 vdd.n1920 vdd.n1301 9.3005
R20759 vdd.n1922 vdd.n1921 9.3005
R20760 vdd.n1291 vdd.n1290 9.3005
R20761 vdd.n1936 vdd.n1935 9.3005
R20762 vdd.n1937 vdd.n1289 9.3005
R20763 vdd.n1939 vdd.n1938 9.3005
R20764 vdd.n1280 vdd.n1279 9.3005
R20765 vdd.n1953 vdd.n1952 9.3005
R20766 vdd.n1954 vdd.n1278 9.3005
R20767 vdd.n1956 vdd.n1955 9.3005
R20768 vdd.n1268 vdd.n1267 9.3005
R20769 vdd.n1972 vdd.n1971 9.3005
R20770 vdd.n1973 vdd.n1266 9.3005
R20771 vdd.n1975 vdd.n1974 9.3005
R20772 vdd.n283 vdd.n282 9.3005
R20773 vdd.n278 vdd.n277 9.3005
R20774 vdd.n289 vdd.n288 9.3005
R20775 vdd.n291 vdd.n290 9.3005
R20776 vdd.n274 vdd.n273 9.3005
R20777 vdd.n297 vdd.n296 9.3005
R20778 vdd.n299 vdd.n298 9.3005
R20779 vdd.n271 vdd.n268 9.3005
R20780 vdd.n306 vdd.n305 9.3005
R20781 vdd.n232 vdd.n231 9.3005
R20782 vdd.n227 vdd.n226 9.3005
R20783 vdd.n238 vdd.n237 9.3005
R20784 vdd.n240 vdd.n239 9.3005
R20785 vdd.n223 vdd.n222 9.3005
R20786 vdd.n246 vdd.n245 9.3005
R20787 vdd.n248 vdd.n247 9.3005
R20788 vdd.n220 vdd.n217 9.3005
R20789 vdd.n255 vdd.n254 9.3005
R20790 vdd.n189 vdd.n188 9.3005
R20791 vdd.n184 vdd.n183 9.3005
R20792 vdd.n195 vdd.n194 9.3005
R20793 vdd.n197 vdd.n196 9.3005
R20794 vdd.n180 vdd.n179 9.3005
R20795 vdd.n203 vdd.n202 9.3005
R20796 vdd.n205 vdd.n204 9.3005
R20797 vdd.n177 vdd.n174 9.3005
R20798 vdd.n212 vdd.n211 9.3005
R20799 vdd.n138 vdd.n137 9.3005
R20800 vdd.n133 vdd.n132 9.3005
R20801 vdd.n144 vdd.n143 9.3005
R20802 vdd.n146 vdd.n145 9.3005
R20803 vdd.n129 vdd.n128 9.3005
R20804 vdd.n152 vdd.n151 9.3005
R20805 vdd.n154 vdd.n153 9.3005
R20806 vdd.n126 vdd.n123 9.3005
R20807 vdd.n161 vdd.n160 9.3005
R20808 vdd.n96 vdd.n95 9.3005
R20809 vdd.n91 vdd.n90 9.3005
R20810 vdd.n102 vdd.n101 9.3005
R20811 vdd.n104 vdd.n103 9.3005
R20812 vdd.n87 vdd.n86 9.3005
R20813 vdd.n110 vdd.n109 9.3005
R20814 vdd.n112 vdd.n111 9.3005
R20815 vdd.n84 vdd.n81 9.3005
R20816 vdd.n119 vdd.n118 9.3005
R20817 vdd.n45 vdd.n44 9.3005
R20818 vdd.n40 vdd.n39 9.3005
R20819 vdd.n51 vdd.n50 9.3005
R20820 vdd.n53 vdd.n52 9.3005
R20821 vdd.n36 vdd.n35 9.3005
R20822 vdd.n59 vdd.n58 9.3005
R20823 vdd.n61 vdd.n60 9.3005
R20824 vdd.n33 vdd.n30 9.3005
R20825 vdd.n68 vdd.n67 9.3005
R20826 vdd.n2946 vdd.n2945 9.3005
R20827 vdd.n2947 vdd.n578 9.3005
R20828 vdd.n577 vdd.n575 9.3005
R20829 vdd.n2953 vdd.n574 9.3005
R20830 vdd.n2954 vdd.n573 9.3005
R20831 vdd.n2955 vdd.n572 9.3005
R20832 vdd.n571 vdd.n569 9.3005
R20833 vdd.n2961 vdd.n568 9.3005
R20834 vdd.n2962 vdd.n567 9.3005
R20835 vdd.n2963 vdd.n566 9.3005
R20836 vdd.n565 vdd.n563 9.3005
R20837 vdd.n2969 vdd.n562 9.3005
R20838 vdd.n2970 vdd.n561 9.3005
R20839 vdd.n2971 vdd.n560 9.3005
R20840 vdd.n559 vdd.n557 9.3005
R20841 vdd.n2977 vdd.n556 9.3005
R20842 vdd.n2978 vdd.n555 9.3005
R20843 vdd.n2979 vdd.n554 9.3005
R20844 vdd.n553 vdd.n551 9.3005
R20845 vdd.n2985 vdd.n550 9.3005
R20846 vdd.n2986 vdd.n549 9.3005
R20847 vdd.n2987 vdd.n548 9.3005
R20848 vdd.n547 vdd.n545 9.3005
R20849 vdd.n2993 vdd.n542 9.3005
R20850 vdd.n2994 vdd.n541 9.3005
R20851 vdd.n2995 vdd.n540 9.3005
R20852 vdd.n539 vdd.n537 9.3005
R20853 vdd.n3001 vdd.n536 9.3005
R20854 vdd.n3002 vdd.n535 9.3005
R20855 vdd.n3003 vdd.n534 9.3005
R20856 vdd.n533 vdd.n531 9.3005
R20857 vdd.n3009 vdd.n530 9.3005
R20858 vdd.n3010 vdd.n529 9.3005
R20859 vdd.n3011 vdd.n528 9.3005
R20860 vdd.n527 vdd.n525 9.3005
R20861 vdd.n3016 vdd.n524 9.3005
R20862 vdd.n3026 vdd.n518 9.3005
R20863 vdd.n3028 vdd.n3027 9.3005
R20864 vdd.n509 vdd.n508 9.3005
R20865 vdd.n3043 vdd.n3042 9.3005
R20866 vdd.n3044 vdd.n507 9.3005
R20867 vdd.n3046 vdd.n3045 9.3005
R20868 vdd.n497 vdd.n496 9.3005
R20869 vdd.n3059 vdd.n3058 9.3005
R20870 vdd.n3060 vdd.n495 9.3005
R20871 vdd.n3062 vdd.n3061 9.3005
R20872 vdd.n485 vdd.n484 9.3005
R20873 vdd.n3076 vdd.n3075 9.3005
R20874 vdd.n3077 vdd.n483 9.3005
R20875 vdd.n3079 vdd.n3078 9.3005
R20876 vdd.n312 vdd.n310 9.3005
R20877 vdd.n3030 vdd.n3029 9.3005
R20878 vdd.n3259 vdd.n3258 9.3005
R20879 vdd.n313 vdd.n311 9.3005
R20880 vdd.n3252 vdd.n320 9.3005
R20881 vdd.n3251 vdd.n321 9.3005
R20882 vdd.n3250 vdd.n322 9.3005
R20883 vdd.n331 vdd.n323 9.3005
R20884 vdd.n3244 vdd.n332 9.3005
R20885 vdd.n3243 vdd.n333 9.3005
R20886 vdd.n3242 vdd.n334 9.3005
R20887 vdd.n342 vdd.n335 9.3005
R20888 vdd.n3236 vdd.n343 9.3005
R20889 vdd.n3235 vdd.n344 9.3005
R20890 vdd.n3234 vdd.n345 9.3005
R20891 vdd.n353 vdd.n346 9.3005
R20892 vdd.n3228 vdd.n3227 9.3005
R20893 vdd.n3224 vdd.n354 9.3005
R20894 vdd.n3223 vdd.n357 9.3005
R20895 vdd.n361 vdd.n358 9.3005
R20896 vdd.n362 vdd.n359 9.3005
R20897 vdd.n3216 vdd.n363 9.3005
R20898 vdd.n3215 vdd.n364 9.3005
R20899 vdd.n3214 vdd.n365 9.3005
R20900 vdd.n369 vdd.n366 9.3005
R20901 vdd.n3209 vdd.n370 9.3005
R20902 vdd.n3208 vdd.n371 9.3005
R20903 vdd.n3207 vdd.n372 9.3005
R20904 vdd.n376 vdd.n373 9.3005
R20905 vdd.n3202 vdd.n377 9.3005
R20906 vdd.n3201 vdd.n378 9.3005
R20907 vdd.n3200 vdd.n379 9.3005
R20908 vdd.n383 vdd.n380 9.3005
R20909 vdd.n3195 vdd.n384 9.3005
R20910 vdd.n3194 vdd.n385 9.3005
R20911 vdd.n3193 vdd.n3192 9.3005
R20912 vdd.n3191 vdd.n386 9.3005
R20913 vdd.n3190 vdd.n3189 9.3005
R20914 vdd.n392 vdd.n391 9.3005
R20915 vdd.n3184 vdd.n396 9.3005
R20916 vdd.n3183 vdd.n397 9.3005
R20917 vdd.n3182 vdd.n398 9.3005
R20918 vdd.n402 vdd.n399 9.3005
R20919 vdd.n3177 vdd.n403 9.3005
R20920 vdd.n3176 vdd.n404 9.3005
R20921 vdd.n3175 vdd.n405 9.3005
R20922 vdd.n409 vdd.n406 9.3005
R20923 vdd.n3170 vdd.n410 9.3005
R20924 vdd.n3169 vdd.n411 9.3005
R20925 vdd.n3168 vdd.n412 9.3005
R20926 vdd.n416 vdd.n413 9.3005
R20927 vdd.n3163 vdd.n417 9.3005
R20928 vdd.n3162 vdd.n418 9.3005
R20929 vdd.n3161 vdd.n419 9.3005
R20930 vdd.n423 vdd.n420 9.3005
R20931 vdd.n3156 vdd.n424 9.3005
R20932 vdd.n3155 vdd.n425 9.3005
R20933 vdd.n3154 vdd.n3153 9.3005
R20934 vdd.n3152 vdd.n426 9.3005
R20935 vdd.n3151 vdd.n3150 9.3005
R20936 vdd.n432 vdd.n431 9.3005
R20937 vdd.n3145 vdd.n436 9.3005
R20938 vdd.n3144 vdd.n437 9.3005
R20939 vdd.n3143 vdd.n438 9.3005
R20940 vdd.n442 vdd.n439 9.3005
R20941 vdd.n3138 vdd.n443 9.3005
R20942 vdd.n3137 vdd.n444 9.3005
R20943 vdd.n3136 vdd.n445 9.3005
R20944 vdd.n449 vdd.n446 9.3005
R20945 vdd.n3131 vdd.n450 9.3005
R20946 vdd.n3130 vdd.n451 9.3005
R20947 vdd.n3129 vdd.n452 9.3005
R20948 vdd.n456 vdd.n453 9.3005
R20949 vdd.n3124 vdd.n457 9.3005
R20950 vdd.n3123 vdd.n458 9.3005
R20951 vdd.n3122 vdd.n459 9.3005
R20952 vdd.n463 vdd.n460 9.3005
R20953 vdd.n3117 vdd.n464 9.3005
R20954 vdd.n3116 vdd.n465 9.3005
R20955 vdd.n3112 vdd.n3109 9.3005
R20956 vdd.n3226 vdd.n3225 9.3005
R20957 vdd.n3036 vdd.n513 9.3005
R20958 vdd.n3038 vdd.n3037 9.3005
R20959 vdd.n503 vdd.n502 9.3005
R20960 vdd.n3051 vdd.n3050 9.3005
R20961 vdd.n3052 vdd.n501 9.3005
R20962 vdd.n3054 vdd.n3053 9.3005
R20963 vdd.n490 vdd.n489 9.3005
R20964 vdd.n3067 vdd.n3066 9.3005
R20965 vdd.n3068 vdd.n488 9.3005
R20966 vdd.n3070 vdd.n3069 9.3005
R20967 vdd.n478 vdd.n477 9.3005
R20968 vdd.n3084 vdd.n3083 9.3005
R20969 vdd.n3085 vdd.n476 9.3005
R20970 vdd.n3087 vdd.n3086 9.3005
R20971 vdd.n3088 vdd.n475 9.3005
R20972 vdd.n3090 vdd.n3089 9.3005
R20973 vdd.n3091 vdd.n474 9.3005
R20974 vdd.n3093 vdd.n3092 9.3005
R20975 vdd.n3094 vdd.n472 9.3005
R20976 vdd.n3096 vdd.n3095 9.3005
R20977 vdd.n3097 vdd.n471 9.3005
R20978 vdd.n3099 vdd.n3098 9.3005
R20979 vdd.n3100 vdd.n469 9.3005
R20980 vdd.n3102 vdd.n3101 9.3005
R20981 vdd.n3103 vdd.n468 9.3005
R20982 vdd.n3105 vdd.n3104 9.3005
R20983 vdd.n3106 vdd.n466 9.3005
R20984 vdd.n3108 vdd.n3107 9.3005
R20985 vdd.n3035 vdd.n3034 9.3005
R20986 vdd.n2899 vdd.n514 9.3005
R20987 vdd.n2904 vdd.n2898 9.3005
R20988 vdd.n2914 vdd.n605 9.3005
R20989 vdd.n2915 vdd.n604 9.3005
R20990 vdd.n603 vdd.n601 9.3005
R20991 vdd.n2921 vdd.n600 9.3005
R20992 vdd.n2922 vdd.n599 9.3005
R20993 vdd.n2923 vdd.n598 9.3005
R20994 vdd.n597 vdd.n595 9.3005
R20995 vdd.n2929 vdd.n594 9.3005
R20996 vdd.n2930 vdd.n593 9.3005
R20997 vdd.n2931 vdd.n592 9.3005
R20998 vdd.n591 vdd.n589 9.3005
R20999 vdd.n2936 vdd.n588 9.3005
R21000 vdd.n2937 vdd.n587 9.3005
R21001 vdd.n583 vdd.n582 9.3005
R21002 vdd.n2943 vdd.n2942 9.3005
R21003 vdd.n2944 vdd.n579 9.3005
R21004 vdd.n1985 vdd.n1984 9.3005
R21005 vdd.n1980 vdd.n1252 9.3005
R21006 vdd.n1581 vdd.n1341 9.3005
R21007 vdd.n1583 vdd.n1582 9.3005
R21008 vdd.n1332 vdd.n1331 9.3005
R21009 vdd.n1596 vdd.n1595 9.3005
R21010 vdd.n1597 vdd.n1330 9.3005
R21011 vdd.n1599 vdd.n1598 9.3005
R21012 vdd.n1319 vdd.n1318 9.3005
R21013 vdd.n1612 vdd.n1611 9.3005
R21014 vdd.n1613 vdd.n1317 9.3005
R21015 vdd.n1615 vdd.n1614 9.3005
R21016 vdd.n1308 vdd.n1307 9.3005
R21017 vdd.n1629 vdd.n1628 9.3005
R21018 vdd.n1630 vdd.n1306 9.3005
R21019 vdd.n1632 vdd.n1631 9.3005
R21020 vdd.n1297 vdd.n1296 9.3005
R21021 vdd.n1927 vdd.n1926 9.3005
R21022 vdd.n1928 vdd.n1295 9.3005
R21023 vdd.n1930 vdd.n1929 9.3005
R21024 vdd.n1285 vdd.n1284 9.3005
R21025 vdd.n1944 vdd.n1943 9.3005
R21026 vdd.n1945 vdd.n1283 9.3005
R21027 vdd.n1947 vdd.n1946 9.3005
R21028 vdd.n1275 vdd.n1274 9.3005
R21029 vdd.n1961 vdd.n1960 9.3005
R21030 vdd.n1962 vdd.n1272 9.3005
R21031 vdd.n1966 vdd.n1965 9.3005
R21032 vdd.n1964 vdd.n1273 9.3005
R21033 vdd.n1963 vdd.n1263 9.3005
R21034 vdd.n1580 vdd.n1579 9.3005
R21035 vdd.n1475 vdd.n1465 9.3005
R21036 vdd.n1477 vdd.n1476 9.3005
R21037 vdd.n1478 vdd.n1464 9.3005
R21038 vdd.n1480 vdd.n1479 9.3005
R21039 vdd.n1481 vdd.n1457 9.3005
R21040 vdd.n1483 vdd.n1482 9.3005
R21041 vdd.n1484 vdd.n1456 9.3005
R21042 vdd.n1486 vdd.n1485 9.3005
R21043 vdd.n1487 vdd.n1449 9.3005
R21044 vdd.n1489 vdd.n1488 9.3005
R21045 vdd.n1490 vdd.n1448 9.3005
R21046 vdd.n1492 vdd.n1491 9.3005
R21047 vdd.n1493 vdd.n1441 9.3005
R21048 vdd.n1495 vdd.n1494 9.3005
R21049 vdd.n1496 vdd.n1440 9.3005
R21050 vdd.n1498 vdd.n1497 9.3005
R21051 vdd.n1499 vdd.n1434 9.3005
R21052 vdd.n1501 vdd.n1500 9.3005
R21053 vdd.n1502 vdd.n1432 9.3005
R21054 vdd.n1504 vdd.n1503 9.3005
R21055 vdd.n1433 vdd.n1430 9.3005
R21056 vdd.n1511 vdd.n1426 9.3005
R21057 vdd.n1513 vdd.n1512 9.3005
R21058 vdd.n1514 vdd.n1425 9.3005
R21059 vdd.n1516 vdd.n1515 9.3005
R21060 vdd.n1517 vdd.n1418 9.3005
R21061 vdd.n1519 vdd.n1518 9.3005
R21062 vdd.n1520 vdd.n1417 9.3005
R21063 vdd.n1522 vdd.n1521 9.3005
R21064 vdd.n1523 vdd.n1410 9.3005
R21065 vdd.n1525 vdd.n1524 9.3005
R21066 vdd.n1526 vdd.n1409 9.3005
R21067 vdd.n1528 vdd.n1527 9.3005
R21068 vdd.n1529 vdd.n1402 9.3005
R21069 vdd.n1531 vdd.n1530 9.3005
R21070 vdd.n1532 vdd.n1401 9.3005
R21071 vdd.n1534 vdd.n1533 9.3005
R21072 vdd.n1535 vdd.n1394 9.3005
R21073 vdd.n1537 vdd.n1536 9.3005
R21074 vdd.n1538 vdd.n1393 9.3005
R21075 vdd.n1540 vdd.n1539 9.3005
R21076 vdd.n1541 vdd.n1386 9.3005
R21077 vdd.n1543 vdd.n1542 9.3005
R21078 vdd.n1544 vdd.n1385 9.3005
R21079 vdd.n1546 vdd.n1545 9.3005
R21080 vdd.n1547 vdd.n1376 9.3005
R21081 vdd.n1549 vdd.n1548 9.3005
R21082 vdd.n1550 vdd.n1375 9.3005
R21083 vdd.n1552 vdd.n1551 9.3005
R21084 vdd.n1553 vdd.n1368 9.3005
R21085 vdd.n1555 vdd.n1554 9.3005
R21086 vdd.n1556 vdd.n1367 9.3005
R21087 vdd.n1558 vdd.n1557 9.3005
R21088 vdd.n1559 vdd.n1360 9.3005
R21089 vdd.n1561 vdd.n1560 9.3005
R21090 vdd.n1562 vdd.n1359 9.3005
R21091 vdd.n1564 vdd.n1563 9.3005
R21092 vdd.n1565 vdd.n1352 9.3005
R21093 vdd.n1567 vdd.n1566 9.3005
R21094 vdd.n1568 vdd.n1351 9.3005
R21095 vdd.n1570 vdd.n1569 9.3005
R21096 vdd.n1571 vdd.n1347 9.3005
R21097 vdd.n1573 vdd.n1572 9.3005
R21098 vdd.n1471 vdd.n1342 9.3005
R21099 vdd.n1338 vdd.n1337 9.3005
R21100 vdd.n1588 vdd.n1587 9.3005
R21101 vdd.n1589 vdd.n1336 9.3005
R21102 vdd.n1591 vdd.n1590 9.3005
R21103 vdd.n1326 vdd.n1325 9.3005
R21104 vdd.n1604 vdd.n1603 9.3005
R21105 vdd.n1605 vdd.n1324 9.3005
R21106 vdd.n1607 vdd.n1606 9.3005
R21107 vdd.n1314 vdd.n1313 9.3005
R21108 vdd.n1621 vdd.n1620 9.3005
R21109 vdd.n1622 vdd.n1312 9.3005
R21110 vdd.n1624 vdd.n1623 9.3005
R21111 vdd.n1303 vdd.n1302 9.3005
R21112 vdd.n1575 vdd.n1574 9.3005
R21113 vdd.n1919 vdd.n1636 9.3005
R21114 vdd.n1840 vdd.n1839 9.3005
R21115 vdd.n1835 vdd.n1834 9.3005
R21116 vdd.n1846 vdd.n1845 9.3005
R21117 vdd.n1848 vdd.n1847 9.3005
R21118 vdd.n1831 vdd.n1830 9.3005
R21119 vdd.n1854 vdd.n1853 9.3005
R21120 vdd.n1856 vdd.n1855 9.3005
R21121 vdd.n1828 vdd.n1825 9.3005
R21122 vdd.n1863 vdd.n1862 9.3005
R21123 vdd.n1891 vdd.n1890 9.3005
R21124 vdd.n1886 vdd.n1885 9.3005
R21125 vdd.n1897 vdd.n1896 9.3005
R21126 vdd.n1899 vdd.n1898 9.3005
R21127 vdd.n1882 vdd.n1881 9.3005
R21128 vdd.n1905 vdd.n1904 9.3005
R21129 vdd.n1907 vdd.n1906 9.3005
R21130 vdd.n1879 vdd.n1876 9.3005
R21131 vdd.n1914 vdd.n1913 9.3005
R21132 vdd.n1746 vdd.n1745 9.3005
R21133 vdd.n1741 vdd.n1740 9.3005
R21134 vdd.n1752 vdd.n1751 9.3005
R21135 vdd.n1754 vdd.n1753 9.3005
R21136 vdd.n1737 vdd.n1736 9.3005
R21137 vdd.n1760 vdd.n1759 9.3005
R21138 vdd.n1762 vdd.n1761 9.3005
R21139 vdd.n1734 vdd.n1731 9.3005
R21140 vdd.n1769 vdd.n1768 9.3005
R21141 vdd.n1797 vdd.n1796 9.3005
R21142 vdd.n1792 vdd.n1791 9.3005
R21143 vdd.n1803 vdd.n1802 9.3005
R21144 vdd.n1805 vdd.n1804 9.3005
R21145 vdd.n1788 vdd.n1787 9.3005
R21146 vdd.n1811 vdd.n1810 9.3005
R21147 vdd.n1813 vdd.n1812 9.3005
R21148 vdd.n1785 vdd.n1782 9.3005
R21149 vdd.n1820 vdd.n1819 9.3005
R21150 vdd.n1653 vdd.n1652 9.3005
R21151 vdd.n1648 vdd.n1647 9.3005
R21152 vdd.n1659 vdd.n1658 9.3005
R21153 vdd.n1661 vdd.n1660 9.3005
R21154 vdd.n1644 vdd.n1643 9.3005
R21155 vdd.n1667 vdd.n1666 9.3005
R21156 vdd.n1669 vdd.n1668 9.3005
R21157 vdd.n1641 vdd.n1638 9.3005
R21158 vdd.n1676 vdd.n1675 9.3005
R21159 vdd.n1704 vdd.n1703 9.3005
R21160 vdd.n1699 vdd.n1698 9.3005
R21161 vdd.n1710 vdd.n1709 9.3005
R21162 vdd.n1712 vdd.n1711 9.3005
R21163 vdd.n1695 vdd.n1694 9.3005
R21164 vdd.n1718 vdd.n1717 9.3005
R21165 vdd.n1720 vdd.n1719 9.3005
R21166 vdd.n1692 vdd.n1689 9.3005
R21167 vdd.n1727 vdd.n1726 9.3005
R21168 vdd.n288 vdd.n287 8.92171
R21169 vdd.n237 vdd.n236 8.92171
R21170 vdd.n194 vdd.n193 8.92171
R21171 vdd.n143 vdd.n142 8.92171
R21172 vdd.n101 vdd.n100 8.92171
R21173 vdd.n50 vdd.n49 8.92171
R21174 vdd.n1845 vdd.n1844 8.92171
R21175 vdd.n1896 vdd.n1895 8.92171
R21176 vdd.n1751 vdd.n1750 8.92171
R21177 vdd.n1802 vdd.n1801 8.92171
R21178 vdd.n1658 vdd.n1657 8.92171
R21179 vdd.n1709 vdd.n1708 8.92171
R21180 vdd.n215 vdd.n121 8.81535
R21181 vdd.n1823 vdd.n1729 8.81535
R21182 vdd.n1958 vdd.t161 8.72962
R21183 vdd.n3048 vdd.t159 8.72962
R21184 vdd.t202 vdd.n1932 8.50289
R21185 vdd.n493 vdd.t169 8.50289
R21186 vdd.n28 vdd.n14 8.42249
R21187 vdd.n1634 vdd.t174 8.27616
R21188 vdd.n3256 vdd.t164 8.27616
R21189 vdd.n3260 vdd.n3259 8.16225
R21190 vdd.n1919 vdd.n1918 8.16225
R21191 vdd.n284 vdd.n278 8.14595
R21192 vdd.n233 vdd.n227 8.14595
R21193 vdd.n190 vdd.n184 8.14595
R21194 vdd.n139 vdd.n133 8.14595
R21195 vdd.n97 vdd.n91 8.14595
R21196 vdd.n46 vdd.n40 8.14595
R21197 vdd.n1841 vdd.n1835 8.14595
R21198 vdd.n1892 vdd.n1886 8.14595
R21199 vdd.n1747 vdd.n1741 8.14595
R21200 vdd.n1798 vdd.n1792 8.14595
R21201 vdd.n1654 vdd.n1648 8.14595
R21202 vdd.n1705 vdd.n1699 8.14595
R21203 vdd.t190 vdd.n1322 8.04943
R21204 vdd.n3247 vdd.t167 8.04943
R21205 vdd.n2136 vdd.n904 7.70933
R21206 vdd.n2136 vdd.n907 7.70933
R21207 vdd.n2142 vdd.n893 7.70933
R21208 vdd.n2148 vdd.n893 7.70933
R21209 vdd.n2148 vdd.n887 7.70933
R21210 vdd.n2154 vdd.n887 7.70933
R21211 vdd.n2160 vdd.n880 7.70933
R21212 vdd.n2160 vdd.n883 7.70933
R21213 vdd.n2166 vdd.n876 7.70933
R21214 vdd.n2173 vdd.n862 7.70933
R21215 vdd.n2179 vdd.n862 7.70933
R21216 vdd.n2185 vdd.n856 7.70933
R21217 vdd.n2191 vdd.n852 7.70933
R21218 vdd.n2197 vdd.n846 7.70933
R21219 vdd.n2209 vdd.n833 7.70933
R21220 vdd.n2215 vdd.n827 7.70933
R21221 vdd.n2215 vdd.n820 7.70933
R21222 vdd.n2223 vdd.n820 7.70933
R21223 vdd.n2305 vdd.n804 7.70933
R21224 vdd.n2657 vdd.n756 7.70933
R21225 vdd.n2669 vdd.n745 7.70933
R21226 vdd.n2669 vdd.n739 7.70933
R21227 vdd.n2675 vdd.n739 7.70933
R21228 vdd.n2681 vdd.n733 7.70933
R21229 vdd.n2687 vdd.n729 7.70933
R21230 vdd.n2693 vdd.n723 7.70933
R21231 vdd.n2705 vdd.n710 7.70933
R21232 vdd.n2711 vdd.n703 7.70933
R21233 vdd.n2711 vdd.n706 7.70933
R21234 vdd.n2718 vdd.n698 7.70933
R21235 vdd.n2724 vdd.n685 7.70933
R21236 vdd.n2730 vdd.n685 7.70933
R21237 vdd.n2736 vdd.n679 7.70933
R21238 vdd.n2736 vdd.n671 7.70933
R21239 vdd.n2787 vdd.n671 7.70933
R21240 vdd.n2787 vdd.n674 7.70933
R21241 vdd.n2793 vdd.n631 7.70933
R21242 vdd.n2863 vdd.n631 7.70933
R21243 vdd.n2716 vdd.n2715 7.49318
R21244 vdd.n2170 vdd.n2169 7.49318
R21245 vdd.n283 vdd.n280 7.3702
R21246 vdd.n232 vdd.n229 7.3702
R21247 vdd.n189 vdd.n186 7.3702
R21248 vdd.n138 vdd.n135 7.3702
R21249 vdd.n96 vdd.n93 7.3702
R21250 vdd.n45 vdd.n42 7.3702
R21251 vdd.n1840 vdd.n1837 7.3702
R21252 vdd.n1891 vdd.n1888 7.3702
R21253 vdd.n1746 vdd.n1743 7.3702
R21254 vdd.n1797 vdd.n1794 7.3702
R21255 vdd.n1653 vdd.n1650 7.3702
R21256 vdd.n1704 vdd.n1701 7.3702
R21257 vdd.n2154 vdd.t112 7.36923
R21258 vdd.t132 vdd.n679 7.36923
R21259 vdd.n2230 vdd.t97 7.25587
R21260 vdd.n2574 vdd.t126 7.25587
R21261 vdd.n1601 vdd.t192 7.1425
R21262 vdd.n3240 vdd.t144 7.1425
R21263 vdd.n1512 vdd.n1511 6.98232
R21264 vdd.n2020 vdd.n2019 6.98232
R21265 vdd.n3155 vdd.n3154 6.98232
R21266 vdd.n2947 vdd.n2946 6.98232
R21267 vdd.n1617 vdd.t148 6.91577
R21268 vdd.n325 vdd.t146 6.91577
R21269 vdd.n1924 vdd.t195 6.68904
R21270 vdd.n3081 vdd.t171 6.68904
R21271 vdd.n1287 vdd.t136 6.46231
R21272 vdd.t204 vdd.n492 6.46231
R21273 vdd.n3260 vdd.n309 6.27748
R21274 vdd.n1918 vdd.n1917 6.27748
R21275 vdd.t110 vdd.n833 5.89549
R21276 vdd.n2681 vdd.t116 5.89549
R21277 vdd.n284 vdd.n283 5.81868
R21278 vdd.n233 vdd.n232 5.81868
R21279 vdd.n190 vdd.n189 5.81868
R21280 vdd.n139 vdd.n138 5.81868
R21281 vdd.n97 vdd.n96 5.81868
R21282 vdd.n46 vdd.n45 5.81868
R21283 vdd.n1841 vdd.n1840 5.81868
R21284 vdd.n1892 vdd.n1891 5.81868
R21285 vdd.n1747 vdd.n1746 5.81868
R21286 vdd.n1798 vdd.n1797 5.81868
R21287 vdd.n1654 vdd.n1653 5.81868
R21288 vdd.n1705 vdd.n1704 5.81868
R21289 vdd.n2313 vdd.n2312 5.77611
R21290 vdd.n1131 vdd.n1130 5.77611
R21291 vdd.n2586 vdd.n2585 5.77611
R21292 vdd.n2802 vdd.n663 5.77611
R21293 vdd.n2868 vdd.n627 5.77611
R21294 vdd.n2480 vdd.n2418 5.77611
R21295 vdd.n2238 vdd.n811 5.77611
R21296 vdd.n1220 vdd.n1083 5.77611
R21297 vdd.n1474 vdd.n1471 5.62474
R21298 vdd.n1983 vdd.n1980 5.62474
R21299 vdd.n3115 vdd.n3112 5.62474
R21300 vdd.n2902 vdd.n2899 5.62474
R21301 vdd.t113 vdd.n856 5.55539
R21302 vdd.n2185 vdd.t108 5.55539
R21303 vdd.t1 vdd.n710 5.55539
R21304 vdd.n2705 vdd.t104 5.55539
R21305 vdd.n876 vdd.t59 5.44203
R21306 vdd.n2718 vdd.t38 5.44203
R21307 vdd.n2142 vdd.t9 5.32866
R21308 vdd.n1166 vdd.t51 5.32866
R21309 vdd.n2663 vdd.t55 5.32866
R21310 vdd.n674 vdd.t5 5.32866
R21311 vdd.n287 vdd.n278 5.04292
R21312 vdd.n236 vdd.n227 5.04292
R21313 vdd.n193 vdd.n184 5.04292
R21314 vdd.n142 vdd.n133 5.04292
R21315 vdd.n100 vdd.n91 5.04292
R21316 vdd.n49 vdd.n40 5.04292
R21317 vdd.n1844 vdd.n1835 5.04292
R21318 vdd.n1895 vdd.n1886 5.04292
R21319 vdd.n1750 vdd.n1741 5.04292
R21320 vdd.n1801 vdd.n1792 5.04292
R21321 vdd.n1657 vdd.n1648 5.04292
R21322 vdd.n1708 vdd.n1699 5.04292
R21323 vdd.n2191 vdd.t118 4.98857
R21324 vdd.n723 vdd.t232 4.98857
R21325 vdd.n1950 vdd.t136 4.8752
R21326 vdd.t131 vdd.t234 4.8752
R21327 vdd.t128 vdd.t124 4.8752
R21328 vdd.t122 vdd.t3 4.8752
R21329 vdd.t106 vdd.t80 4.8752
R21330 vdd.n3056 vdd.t204 4.8752
R21331 vdd.n2314 vdd.n2313 4.83952
R21332 vdd.n1130 vdd.n1129 4.83952
R21333 vdd.n2587 vdd.n2586 4.83952
R21334 vdd.n663 vdd.n658 4.83952
R21335 vdd.n627 vdd.n622 4.83952
R21336 vdd.n2477 vdd.n2418 4.83952
R21337 vdd.n2241 vdd.n811 4.83952
R21338 vdd.n1223 vdd.n1083 4.83952
R21339 vdd.n1988 vdd.n1987 4.74817
R21340 vdd.n1256 vdd.n1251 4.74817
R21341 vdd.n953 vdd.n950 4.74817
R21342 vdd.n2081 vdd.n949 4.74817
R21343 vdd.n2086 vdd.n950 4.74817
R21344 vdd.n2085 vdd.n949 4.74817
R21345 vdd.n521 vdd.n519 4.74817
R21346 vdd.n3017 vdd.n522 4.74817
R21347 vdd.n3020 vdd.n522 4.74817
R21348 vdd.n3021 vdd.n521 4.74817
R21349 vdd.n2909 vdd.n606 4.74817
R21350 vdd.n2905 vdd.n608 4.74817
R21351 vdd.n2908 vdd.n608 4.74817
R21352 vdd.n2913 vdd.n606 4.74817
R21353 vdd.n1987 vdd.n1049 4.74817
R21354 vdd.n1253 vdd.n1251 4.74817
R21355 vdd.n309 vdd.n308 4.7074
R21356 vdd.n215 vdd.n214 4.7074
R21357 vdd.n1917 vdd.n1916 4.7074
R21358 vdd.n1823 vdd.n1822 4.7074
R21359 vdd.t195 vdd.n1293 4.64847
R21360 vdd.n2166 vdd.t0 4.64847
R21361 vdd.n846 vdd.t133 4.64847
R21362 vdd.n2687 vdd.t109 4.64847
R21363 vdd.n698 vdd.t101 4.64847
R21364 vdd.n3072 vdd.t171 4.64847
R21365 vdd.n1626 vdd.t148 4.42174
R21366 vdd.n3254 vdd.t146 4.42174
R21367 vdd.n288 vdd.n276 4.26717
R21368 vdd.n237 vdd.n225 4.26717
R21369 vdd.n194 vdd.n182 4.26717
R21370 vdd.n143 vdd.n131 4.26717
R21371 vdd.n101 vdd.n89 4.26717
R21372 vdd.n50 vdd.n38 4.26717
R21373 vdd.n1845 vdd.n1833 4.26717
R21374 vdd.n1896 vdd.n1884 4.26717
R21375 vdd.n1751 vdd.n1739 4.26717
R21376 vdd.n1802 vdd.n1790 4.26717
R21377 vdd.n1658 vdd.n1646 4.26717
R21378 vdd.n1709 vdd.n1697 4.26717
R21379 vdd.t192 vdd.n1321 4.19501
R21380 vdd.t144 vdd.n329 4.19501
R21381 vdd.n309 vdd.n215 4.10845
R21382 vdd.n1917 vdd.n1823 4.10845
R21383 vdd.n265 vdd.t226 4.06363
R21384 vdd.n265 vdd.t158 4.06363
R21385 vdd.n263 vdd.t179 4.06363
R21386 vdd.n263 vdd.t225 4.06363
R21387 vdd.n261 vdd.t227 4.06363
R21388 vdd.n261 vdd.t178 4.06363
R21389 vdd.n259 vdd.t183 4.06363
R21390 vdd.n259 vdd.t185 4.06363
R21391 vdd.n257 vdd.t211 4.06363
R21392 vdd.n257 vdd.t150 4.06363
R21393 vdd.n171 vdd.t219 4.06363
R21394 vdd.n171 vdd.t145 4.06363
R21395 vdd.n169 vdd.t166 4.06363
R21396 vdd.n169 vdd.t218 4.06363
R21397 vdd.n167 vdd.t220 4.06363
R21398 vdd.n167 vdd.t165 4.06363
R21399 vdd.n165 vdd.t170 4.06363
R21400 vdd.n165 vdd.t172 4.06363
R21401 vdd.n163 vdd.t205 4.06363
R21402 vdd.n163 vdd.t135 4.06363
R21403 vdd.n78 vdd.t168 4.06363
R21404 vdd.n78 vdd.t216 4.06363
R21405 vdd.n76 vdd.t147 4.06363
R21406 vdd.n76 vdd.t188 4.06363
R21407 vdd.n74 vdd.t139 4.06363
R21408 vdd.n74 vdd.t173 4.06363
R21409 vdd.n72 vdd.t223 4.06363
R21410 vdd.n72 vdd.t210 4.06363
R21411 vdd.n70 vdd.t213 4.06363
R21412 vdd.n70 vdd.t180 4.06363
R21413 vdd.n1865 vdd.t194 4.06363
R21414 vdd.n1865 vdd.t154 4.06363
R21415 vdd.n1867 vdd.t229 4.06363
R21416 vdd.n1867 vdd.t209 4.06363
R21417 vdd.n1869 vdd.t207 4.06363
R21418 vdd.n1869 vdd.t177 4.06363
R21419 vdd.n1871 vdd.t176 4.06363
R21420 vdd.n1871 vdd.t208 4.06363
R21421 vdd.n1873 vdd.t199 4.06363
R21422 vdd.n1873 vdd.t198 4.06363
R21423 vdd.n1771 vdd.t184 4.06363
R21424 vdd.n1771 vdd.t137 4.06363
R21425 vdd.n1773 vdd.t222 4.06363
R21426 vdd.n1773 vdd.t203 4.06363
R21427 vdd.n1775 vdd.t200 4.06363
R21428 vdd.n1775 vdd.t163 4.06363
R21429 vdd.n1777 vdd.t157 4.06363
R21430 vdd.n1777 vdd.t201 4.06363
R21431 vdd.n1779 vdd.t193 4.06363
R21432 vdd.n1779 vdd.t191 4.06363
R21433 vdd.n1678 vdd.t182 4.06363
R21434 vdd.n1678 vdd.t214 4.06363
R21435 vdd.n1680 vdd.t196 4.06363
R21436 vdd.n1680 vdd.t224 4.06363
R21437 vdd.n1682 vdd.t175 4.06363
R21438 vdd.n1682 vdd.t143 4.06363
R21439 vdd.n1684 vdd.t189 4.06363
R21440 vdd.n1684 vdd.t149 4.06363
R21441 vdd.n1686 vdd.t217 4.06363
R21442 vdd.n1686 vdd.t228 4.06363
R21443 vdd.n26 vdd.t88 3.9605
R21444 vdd.n26 vdd.t93 3.9605
R21445 vdd.n23 vdd.t84 3.9605
R21446 vdd.n23 vdd.t96 3.9605
R21447 vdd.n21 vdd.t90 3.9605
R21448 vdd.n21 vdd.t94 3.9605
R21449 vdd.n20 vdd.t81 3.9605
R21450 vdd.n20 vdd.t82 3.9605
R21451 vdd.n15 vdd.t92 3.9605
R21452 vdd.n15 vdd.t91 3.9605
R21453 vdd.n16 vdd.t86 3.9605
R21454 vdd.n16 vdd.t83 3.9605
R21455 vdd.n18 vdd.t85 3.9605
R21456 vdd.n18 vdd.t89 3.9605
R21457 vdd.n25 vdd.t87 3.9605
R21458 vdd.n25 vdd.t95 3.9605
R21459 vdd.n2223 vdd.t230 3.85492
R21460 vdd.n1166 vdd.t230 3.85492
R21461 vdd.n2663 vdd.t102 3.85492
R21462 vdd.t102 vdd.n745 3.85492
R21463 vdd.n7 vdd.t107 3.61217
R21464 vdd.n7 vdd.t233 3.61217
R21465 vdd.n8 vdd.t123 3.61217
R21466 vdd.n8 vdd.t117 3.61217
R21467 vdd.n10 vdd.t127 3.61217
R21468 vdd.n10 vdd.t103 3.61217
R21469 vdd.n12 vdd.t115 3.61217
R21470 vdd.n12 vdd.t130 3.61217
R21471 vdd.n5 vdd.t100 3.61217
R21472 vdd.n5 vdd.t121 3.61217
R21473 vdd.n3 vdd.t231 3.61217
R21474 vdd.n3 vdd.t98 3.61217
R21475 vdd.n1 vdd.t111 3.61217
R21476 vdd.n1 vdd.t125 3.61217
R21477 vdd.n0 vdd.t119 3.61217
R21478 vdd.n0 vdd.t235 3.61217
R21479 vdd.n292 vdd.n291 3.49141
R21480 vdd.n241 vdd.n240 3.49141
R21481 vdd.n198 vdd.n197 3.49141
R21482 vdd.n147 vdd.n146 3.49141
R21483 vdd.n105 vdd.n104 3.49141
R21484 vdd.n54 vdd.n53 3.49141
R21485 vdd.n1849 vdd.n1848 3.49141
R21486 vdd.n1900 vdd.n1899 3.49141
R21487 vdd.n1755 vdd.n1754 3.49141
R21488 vdd.n1806 vdd.n1805 3.49141
R21489 vdd.n1662 vdd.n1661 3.49141
R21490 vdd.n1713 vdd.n1712 3.49141
R21491 vdd.n2377 vdd.t99 3.40145
R21492 vdd.n2650 vdd.t129 3.40145
R21493 vdd.n1609 vdd.t190 3.28809
R21494 vdd.t167 vdd.n3246 3.28809
R21495 vdd.n2715 vdd.n2714 3.12245
R21496 vdd.n2171 vdd.n2170 3.12245
R21497 vdd.n1310 vdd.t174 3.06136
R21498 vdd.n883 vdd.t0 3.06136
R21499 vdd.n2203 vdd.t133 3.06136
R21500 vdd.n2559 vdd.t109 3.06136
R21501 vdd.n2724 vdd.t101 3.06136
R21502 vdd.t164 vdd.n3255 3.06136
R21503 vdd.n1933 vdd.t202 2.83463
R21504 vdd.n3073 vdd.t169 2.83463
R21505 vdd.n1187 vdd.t118 2.72126
R21506 vdd.n2699 vdd.t232 2.72126
R21507 vdd.n295 vdd.n274 2.71565
R21508 vdd.n244 vdd.n223 2.71565
R21509 vdd.n201 vdd.n180 2.71565
R21510 vdd.n150 vdd.n129 2.71565
R21511 vdd.n108 vdd.n87 2.71565
R21512 vdd.n57 vdd.n36 2.71565
R21513 vdd.n1852 vdd.n1831 2.71565
R21514 vdd.n1903 vdd.n1882 2.71565
R21515 vdd.n1758 vdd.n1737 2.71565
R21516 vdd.n1809 vdd.n1788 2.71565
R21517 vdd.n1665 vdd.n1644 2.71565
R21518 vdd.n1716 vdd.n1695 2.71565
R21519 vdd.n1949 vdd.t161 2.6079
R21520 vdd.t159 vdd.n499 2.6079
R21521 vdd.t124 vdd.n827 2.49453
R21522 vdd.n2675 vdd.t122 2.49453
R21523 vdd.n282 vdd.n281 2.4129
R21524 vdd.n231 vdd.n230 2.4129
R21525 vdd.n188 vdd.n187 2.4129
R21526 vdd.n137 vdd.n136 2.4129
R21527 vdd.n95 vdd.n94 2.4129
R21528 vdd.n44 vdd.n43 2.4129
R21529 vdd.n1839 vdd.n1838 2.4129
R21530 vdd.n1890 vdd.n1889 2.4129
R21531 vdd.n1745 vdd.n1744 2.4129
R21532 vdd.n1796 vdd.n1795 2.4129
R21533 vdd.n1652 vdd.n1651 2.4129
R21534 vdd.n1703 vdd.n1702 2.4129
R21535 vdd.n907 vdd.t9 2.38117
R21536 vdd.n2230 vdd.t51 2.38117
R21537 vdd.n2574 vdd.t55 2.38117
R21538 vdd.n2793 vdd.t5 2.38117
R21539 vdd.n2093 vdd.n950 2.27742
R21540 vdd.n2093 vdd.n949 2.27742
R21541 vdd.n2829 vdd.n522 2.27742
R21542 vdd.n2829 vdd.n521 2.27742
R21543 vdd.n2897 vdd.n608 2.27742
R21544 vdd.n2897 vdd.n606 2.27742
R21545 vdd.n1987 vdd.n1986 2.27742
R21546 vdd.n1986 vdd.n1251 2.27742
R21547 vdd.n2179 vdd.t113 2.15444
R21548 vdd.n1187 vdd.t108 2.15444
R21549 vdd.n2699 vdd.t1 2.15444
R21550 vdd.t104 vdd.n703 2.15444
R21551 vdd.n296 vdd.n272 1.93989
R21552 vdd.n245 vdd.n221 1.93989
R21553 vdd.n202 vdd.n178 1.93989
R21554 vdd.n151 vdd.n127 1.93989
R21555 vdd.n109 vdd.n85 1.93989
R21556 vdd.n58 vdd.n34 1.93989
R21557 vdd.n1853 vdd.n1829 1.93989
R21558 vdd.n1904 vdd.n1880 1.93989
R21559 vdd.n1759 vdd.n1735 1.93989
R21560 vdd.n1810 vdd.n1786 1.93989
R21561 vdd.n1666 vdd.n1642 1.93989
R21562 vdd.n1717 vdd.n1693 1.93989
R21563 vdd.n2203 vdd.t110 1.81434
R21564 vdd.n2559 vdd.t116 1.81434
R21565 vdd.n2197 vdd.t234 1.58761
R21566 vdd.n729 vdd.t106 1.58761
R21567 vdd.n1345 vdd.t25 1.47425
R21568 vdd.t21 vdd.n3231 1.47425
R21569 vdd.n2173 vdd.t105 1.24752
R21570 vdd.n852 vdd.t131 1.24752
R21571 vdd.n2693 vdd.t80 1.24752
R21572 vdd.n706 vdd.t2 1.24752
R21573 vdd.n307 vdd.n267 1.16414
R21574 vdd.n300 vdd.n299 1.16414
R21575 vdd.n256 vdd.n216 1.16414
R21576 vdd.n249 vdd.n248 1.16414
R21577 vdd.n213 vdd.n173 1.16414
R21578 vdd.n206 vdd.n205 1.16414
R21579 vdd.n162 vdd.n122 1.16414
R21580 vdd.n155 vdd.n154 1.16414
R21581 vdd.n120 vdd.n80 1.16414
R21582 vdd.n113 vdd.n112 1.16414
R21583 vdd.n69 vdd.n29 1.16414
R21584 vdd.n62 vdd.n61 1.16414
R21585 vdd.n1864 vdd.n1824 1.16414
R21586 vdd.n1857 vdd.n1856 1.16414
R21587 vdd.n1915 vdd.n1875 1.16414
R21588 vdd.n1908 vdd.n1907 1.16414
R21589 vdd.n1770 vdd.n1730 1.16414
R21590 vdd.n1763 vdd.n1762 1.16414
R21591 vdd.n1821 vdd.n1781 1.16414
R21592 vdd.n1814 vdd.n1813 1.16414
R21593 vdd.n1677 vdd.n1637 1.16414
R21594 vdd.n1670 vdd.n1669 1.16414
R21595 vdd.n1728 vdd.n1688 1.16414
R21596 vdd.n1721 vdd.n1720 1.16414
R21597 vdd.n1941 vdd.t181 1.02079
R21598 vdd.t59 vdd.t105 1.02079
R21599 vdd.t2 vdd.t38 1.02079
R21600 vdd.n3064 vdd.t134 1.02079
R21601 vdd.n1475 vdd.n1474 0.970197
R21602 vdd.n1984 vdd.n1983 0.970197
R21603 vdd.n3116 vdd.n3115 0.970197
R21604 vdd.n2904 vdd.n2902 0.970197
R21605 vdd.n1918 vdd.n28 0.90431
R21606 vdd vdd.n3260 0.896477
R21607 vdd.t142 vdd.n1299 0.794056
R21608 vdd.n1968 vdd.t17 0.794056
R21609 vdd.t13 vdd.n511 0.794056
R21610 vdd.n481 vdd.t138 0.794056
R21611 vdd.n1618 vdd.t156 0.567326
R21612 vdd.n3248 vdd.t187 0.567326
R21613 vdd.n1974 vdd.n951 0.509646
R21614 vdd.n3029 vdd.n3028 0.509646
R21615 vdd.n3227 vdd.n3226 0.509646
R21616 vdd.n3109 vdd.n3108 0.509646
R21617 vdd.n3035 vdd.n514 0.509646
R21618 vdd.n1963 vdd.n1252 0.509646
R21619 vdd.n1580 vdd.n1342 0.509646
R21620 vdd.n1574 vdd.n1573 0.509646
R21621 vdd.n4 vdd.n2 0.459552
R21622 vdd.n11 vdd.n9 0.459552
R21623 vdd.t97 vdd.n804 0.453961
R21624 vdd.n2657 vdd.t126 0.453961
R21625 vdd.n305 vdd.n304 0.388379
R21626 vdd.n271 vdd.n269 0.388379
R21627 vdd.n254 vdd.n253 0.388379
R21628 vdd.n220 vdd.n218 0.388379
R21629 vdd.n211 vdd.n210 0.388379
R21630 vdd.n177 vdd.n175 0.388379
R21631 vdd.n160 vdd.n159 0.388379
R21632 vdd.n126 vdd.n124 0.388379
R21633 vdd.n118 vdd.n117 0.388379
R21634 vdd.n84 vdd.n82 0.388379
R21635 vdd.n67 vdd.n66 0.388379
R21636 vdd.n33 vdd.n31 0.388379
R21637 vdd.n1862 vdd.n1861 0.388379
R21638 vdd.n1828 vdd.n1826 0.388379
R21639 vdd.n1913 vdd.n1912 0.388379
R21640 vdd.n1879 vdd.n1877 0.388379
R21641 vdd.n1768 vdd.n1767 0.388379
R21642 vdd.n1734 vdd.n1732 0.388379
R21643 vdd.n1819 vdd.n1818 0.388379
R21644 vdd.n1785 vdd.n1783 0.388379
R21645 vdd.n1675 vdd.n1674 0.388379
R21646 vdd.n1641 vdd.n1639 0.388379
R21647 vdd.n1726 vdd.n1725 0.388379
R21648 vdd.n1692 vdd.n1690 0.388379
R21649 vdd.n19 vdd.n17 0.387128
R21650 vdd.n24 vdd.n22 0.387128
R21651 vdd.n6 vdd.n4 0.358259
R21652 vdd.n13 vdd.n11 0.358259
R21653 vdd.n260 vdd.n258 0.358259
R21654 vdd.n262 vdd.n260 0.358259
R21655 vdd.n264 vdd.n262 0.358259
R21656 vdd.n266 vdd.n264 0.358259
R21657 vdd.n308 vdd.n266 0.358259
R21658 vdd.n166 vdd.n164 0.358259
R21659 vdd.n168 vdd.n166 0.358259
R21660 vdd.n170 vdd.n168 0.358259
R21661 vdd.n172 vdd.n170 0.358259
R21662 vdd.n214 vdd.n172 0.358259
R21663 vdd.n73 vdd.n71 0.358259
R21664 vdd.n75 vdd.n73 0.358259
R21665 vdd.n77 vdd.n75 0.358259
R21666 vdd.n79 vdd.n77 0.358259
R21667 vdd.n121 vdd.n79 0.358259
R21668 vdd.n1916 vdd.n1874 0.358259
R21669 vdd.n1874 vdd.n1872 0.358259
R21670 vdd.n1872 vdd.n1870 0.358259
R21671 vdd.n1870 vdd.n1868 0.358259
R21672 vdd.n1868 vdd.n1866 0.358259
R21673 vdd.n1822 vdd.n1780 0.358259
R21674 vdd.n1780 vdd.n1778 0.358259
R21675 vdd.n1778 vdd.n1776 0.358259
R21676 vdd.n1776 vdd.n1774 0.358259
R21677 vdd.n1774 vdd.n1772 0.358259
R21678 vdd.n1729 vdd.n1687 0.358259
R21679 vdd.n1687 vdd.n1685 0.358259
R21680 vdd.n1685 vdd.n1683 0.358259
R21681 vdd.n1683 vdd.n1681 0.358259
R21682 vdd.n1681 vdd.n1679 0.358259
R21683 vdd.t140 vdd.n1328 0.340595
R21684 vdd.t112 vdd.n880 0.340595
R21685 vdd.n2209 vdd.t128 0.340595
R21686 vdd.t3 vdd.n733 0.340595
R21687 vdd.n2730 vdd.t132 0.340595
R21688 vdd.n3239 vdd.t151 0.340595
R21689 vdd.n14 vdd.n6 0.334552
R21690 vdd.n14 vdd.n13 0.334552
R21691 vdd.n27 vdd.n19 0.21707
R21692 vdd.n27 vdd.n24 0.21707
R21693 vdd.n306 vdd.n268 0.155672
R21694 vdd.n298 vdd.n268 0.155672
R21695 vdd.n298 vdd.n297 0.155672
R21696 vdd.n297 vdd.n273 0.155672
R21697 vdd.n290 vdd.n273 0.155672
R21698 vdd.n290 vdd.n289 0.155672
R21699 vdd.n289 vdd.n277 0.155672
R21700 vdd.n282 vdd.n277 0.155672
R21701 vdd.n255 vdd.n217 0.155672
R21702 vdd.n247 vdd.n217 0.155672
R21703 vdd.n247 vdd.n246 0.155672
R21704 vdd.n246 vdd.n222 0.155672
R21705 vdd.n239 vdd.n222 0.155672
R21706 vdd.n239 vdd.n238 0.155672
R21707 vdd.n238 vdd.n226 0.155672
R21708 vdd.n231 vdd.n226 0.155672
R21709 vdd.n212 vdd.n174 0.155672
R21710 vdd.n204 vdd.n174 0.155672
R21711 vdd.n204 vdd.n203 0.155672
R21712 vdd.n203 vdd.n179 0.155672
R21713 vdd.n196 vdd.n179 0.155672
R21714 vdd.n196 vdd.n195 0.155672
R21715 vdd.n195 vdd.n183 0.155672
R21716 vdd.n188 vdd.n183 0.155672
R21717 vdd.n161 vdd.n123 0.155672
R21718 vdd.n153 vdd.n123 0.155672
R21719 vdd.n153 vdd.n152 0.155672
R21720 vdd.n152 vdd.n128 0.155672
R21721 vdd.n145 vdd.n128 0.155672
R21722 vdd.n145 vdd.n144 0.155672
R21723 vdd.n144 vdd.n132 0.155672
R21724 vdd.n137 vdd.n132 0.155672
R21725 vdd.n119 vdd.n81 0.155672
R21726 vdd.n111 vdd.n81 0.155672
R21727 vdd.n111 vdd.n110 0.155672
R21728 vdd.n110 vdd.n86 0.155672
R21729 vdd.n103 vdd.n86 0.155672
R21730 vdd.n103 vdd.n102 0.155672
R21731 vdd.n102 vdd.n90 0.155672
R21732 vdd.n95 vdd.n90 0.155672
R21733 vdd.n68 vdd.n30 0.155672
R21734 vdd.n60 vdd.n30 0.155672
R21735 vdd.n60 vdd.n59 0.155672
R21736 vdd.n59 vdd.n35 0.155672
R21737 vdd.n52 vdd.n35 0.155672
R21738 vdd.n52 vdd.n51 0.155672
R21739 vdd.n51 vdd.n39 0.155672
R21740 vdd.n44 vdd.n39 0.155672
R21741 vdd.n1863 vdd.n1825 0.155672
R21742 vdd.n1855 vdd.n1825 0.155672
R21743 vdd.n1855 vdd.n1854 0.155672
R21744 vdd.n1854 vdd.n1830 0.155672
R21745 vdd.n1847 vdd.n1830 0.155672
R21746 vdd.n1847 vdd.n1846 0.155672
R21747 vdd.n1846 vdd.n1834 0.155672
R21748 vdd.n1839 vdd.n1834 0.155672
R21749 vdd.n1914 vdd.n1876 0.155672
R21750 vdd.n1906 vdd.n1876 0.155672
R21751 vdd.n1906 vdd.n1905 0.155672
R21752 vdd.n1905 vdd.n1881 0.155672
R21753 vdd.n1898 vdd.n1881 0.155672
R21754 vdd.n1898 vdd.n1897 0.155672
R21755 vdd.n1897 vdd.n1885 0.155672
R21756 vdd.n1890 vdd.n1885 0.155672
R21757 vdd.n1769 vdd.n1731 0.155672
R21758 vdd.n1761 vdd.n1731 0.155672
R21759 vdd.n1761 vdd.n1760 0.155672
R21760 vdd.n1760 vdd.n1736 0.155672
R21761 vdd.n1753 vdd.n1736 0.155672
R21762 vdd.n1753 vdd.n1752 0.155672
R21763 vdd.n1752 vdd.n1740 0.155672
R21764 vdd.n1745 vdd.n1740 0.155672
R21765 vdd.n1820 vdd.n1782 0.155672
R21766 vdd.n1812 vdd.n1782 0.155672
R21767 vdd.n1812 vdd.n1811 0.155672
R21768 vdd.n1811 vdd.n1787 0.155672
R21769 vdd.n1804 vdd.n1787 0.155672
R21770 vdd.n1804 vdd.n1803 0.155672
R21771 vdd.n1803 vdd.n1791 0.155672
R21772 vdd.n1796 vdd.n1791 0.155672
R21773 vdd.n1676 vdd.n1638 0.155672
R21774 vdd.n1668 vdd.n1638 0.155672
R21775 vdd.n1668 vdd.n1667 0.155672
R21776 vdd.n1667 vdd.n1643 0.155672
R21777 vdd.n1660 vdd.n1643 0.155672
R21778 vdd.n1660 vdd.n1659 0.155672
R21779 vdd.n1659 vdd.n1647 0.155672
R21780 vdd.n1652 vdd.n1647 0.155672
R21781 vdd.n1727 vdd.n1689 0.155672
R21782 vdd.n1719 vdd.n1689 0.155672
R21783 vdd.n1719 vdd.n1718 0.155672
R21784 vdd.n1718 vdd.n1694 0.155672
R21785 vdd.n1711 vdd.n1694 0.155672
R21786 vdd.n1711 vdd.n1710 0.155672
R21787 vdd.n1710 vdd.n1698 0.155672
R21788 vdd.n1703 vdd.n1698 0.155672
R21789 vdd.n956 vdd.n948 0.152939
R21790 vdd.n960 vdd.n956 0.152939
R21791 vdd.n961 vdd.n960 0.152939
R21792 vdd.n962 vdd.n961 0.152939
R21793 vdd.n963 vdd.n962 0.152939
R21794 vdd.n967 vdd.n963 0.152939
R21795 vdd.n968 vdd.n967 0.152939
R21796 vdd.n969 vdd.n968 0.152939
R21797 vdd.n970 vdd.n969 0.152939
R21798 vdd.n974 vdd.n970 0.152939
R21799 vdd.n975 vdd.n974 0.152939
R21800 vdd.n976 vdd.n975 0.152939
R21801 vdd.n2057 vdd.n976 0.152939
R21802 vdd.n2057 vdd.n2056 0.152939
R21803 vdd.n2056 vdd.n2055 0.152939
R21804 vdd.n2055 vdd.n982 0.152939
R21805 vdd.n987 vdd.n982 0.152939
R21806 vdd.n988 vdd.n987 0.152939
R21807 vdd.n989 vdd.n988 0.152939
R21808 vdd.n993 vdd.n989 0.152939
R21809 vdd.n994 vdd.n993 0.152939
R21810 vdd.n995 vdd.n994 0.152939
R21811 vdd.n996 vdd.n995 0.152939
R21812 vdd.n1000 vdd.n996 0.152939
R21813 vdd.n1001 vdd.n1000 0.152939
R21814 vdd.n1002 vdd.n1001 0.152939
R21815 vdd.n1003 vdd.n1002 0.152939
R21816 vdd.n1007 vdd.n1003 0.152939
R21817 vdd.n1008 vdd.n1007 0.152939
R21818 vdd.n1009 vdd.n1008 0.152939
R21819 vdd.n1010 vdd.n1009 0.152939
R21820 vdd.n1014 vdd.n1010 0.152939
R21821 vdd.n1015 vdd.n1014 0.152939
R21822 vdd.n1016 vdd.n1015 0.152939
R21823 vdd.n2018 vdd.n1016 0.152939
R21824 vdd.n2018 vdd.n2017 0.152939
R21825 vdd.n2017 vdd.n2016 0.152939
R21826 vdd.n2016 vdd.n1022 0.152939
R21827 vdd.n1027 vdd.n1022 0.152939
R21828 vdd.n1028 vdd.n1027 0.152939
R21829 vdd.n1029 vdd.n1028 0.152939
R21830 vdd.n1033 vdd.n1029 0.152939
R21831 vdd.n1034 vdd.n1033 0.152939
R21832 vdd.n1035 vdd.n1034 0.152939
R21833 vdd.n1036 vdd.n1035 0.152939
R21834 vdd.n1040 vdd.n1036 0.152939
R21835 vdd.n1041 vdd.n1040 0.152939
R21836 vdd.n1042 vdd.n1041 0.152939
R21837 vdd.n1043 vdd.n1042 0.152939
R21838 vdd.n1047 vdd.n1043 0.152939
R21839 vdd.n1048 vdd.n1047 0.152939
R21840 vdd.n2092 vdd.n951 0.152939
R21841 vdd.n1921 vdd.n1920 0.152939
R21842 vdd.n1921 vdd.n1290 0.152939
R21843 vdd.n1936 vdd.n1290 0.152939
R21844 vdd.n1937 vdd.n1936 0.152939
R21845 vdd.n1938 vdd.n1937 0.152939
R21846 vdd.n1938 vdd.n1279 0.152939
R21847 vdd.n1953 vdd.n1279 0.152939
R21848 vdd.n1954 vdd.n1953 0.152939
R21849 vdd.n1955 vdd.n1954 0.152939
R21850 vdd.n1955 vdd.n1267 0.152939
R21851 vdd.n1972 vdd.n1267 0.152939
R21852 vdd.n1973 vdd.n1972 0.152939
R21853 vdd.n1974 vdd.n1973 0.152939
R21854 vdd.n527 vdd.n524 0.152939
R21855 vdd.n528 vdd.n527 0.152939
R21856 vdd.n529 vdd.n528 0.152939
R21857 vdd.n530 vdd.n529 0.152939
R21858 vdd.n533 vdd.n530 0.152939
R21859 vdd.n534 vdd.n533 0.152939
R21860 vdd.n535 vdd.n534 0.152939
R21861 vdd.n536 vdd.n535 0.152939
R21862 vdd.n539 vdd.n536 0.152939
R21863 vdd.n540 vdd.n539 0.152939
R21864 vdd.n541 vdd.n540 0.152939
R21865 vdd.n542 vdd.n541 0.152939
R21866 vdd.n547 vdd.n542 0.152939
R21867 vdd.n548 vdd.n547 0.152939
R21868 vdd.n549 vdd.n548 0.152939
R21869 vdd.n550 vdd.n549 0.152939
R21870 vdd.n553 vdd.n550 0.152939
R21871 vdd.n554 vdd.n553 0.152939
R21872 vdd.n555 vdd.n554 0.152939
R21873 vdd.n556 vdd.n555 0.152939
R21874 vdd.n559 vdd.n556 0.152939
R21875 vdd.n560 vdd.n559 0.152939
R21876 vdd.n561 vdd.n560 0.152939
R21877 vdd.n562 vdd.n561 0.152939
R21878 vdd.n565 vdd.n562 0.152939
R21879 vdd.n566 vdd.n565 0.152939
R21880 vdd.n567 vdd.n566 0.152939
R21881 vdd.n568 vdd.n567 0.152939
R21882 vdd.n571 vdd.n568 0.152939
R21883 vdd.n572 vdd.n571 0.152939
R21884 vdd.n573 vdd.n572 0.152939
R21885 vdd.n574 vdd.n573 0.152939
R21886 vdd.n577 vdd.n574 0.152939
R21887 vdd.n578 vdd.n577 0.152939
R21888 vdd.n2945 vdd.n578 0.152939
R21889 vdd.n2945 vdd.n2944 0.152939
R21890 vdd.n2944 vdd.n2943 0.152939
R21891 vdd.n2943 vdd.n582 0.152939
R21892 vdd.n587 vdd.n582 0.152939
R21893 vdd.n588 vdd.n587 0.152939
R21894 vdd.n591 vdd.n588 0.152939
R21895 vdd.n592 vdd.n591 0.152939
R21896 vdd.n593 vdd.n592 0.152939
R21897 vdd.n594 vdd.n593 0.152939
R21898 vdd.n597 vdd.n594 0.152939
R21899 vdd.n598 vdd.n597 0.152939
R21900 vdd.n599 vdd.n598 0.152939
R21901 vdd.n600 vdd.n599 0.152939
R21902 vdd.n603 vdd.n600 0.152939
R21903 vdd.n604 vdd.n603 0.152939
R21904 vdd.n605 vdd.n604 0.152939
R21905 vdd.n3028 vdd.n518 0.152939
R21906 vdd.n3029 vdd.n508 0.152939
R21907 vdd.n3043 vdd.n508 0.152939
R21908 vdd.n3044 vdd.n3043 0.152939
R21909 vdd.n3045 vdd.n3044 0.152939
R21910 vdd.n3045 vdd.n496 0.152939
R21911 vdd.n3059 vdd.n496 0.152939
R21912 vdd.n3060 vdd.n3059 0.152939
R21913 vdd.n3061 vdd.n3060 0.152939
R21914 vdd.n3061 vdd.n484 0.152939
R21915 vdd.n3076 vdd.n484 0.152939
R21916 vdd.n3077 vdd.n3076 0.152939
R21917 vdd.n3078 vdd.n3077 0.152939
R21918 vdd.n3078 vdd.n310 0.152939
R21919 vdd.n320 vdd.n311 0.152939
R21920 vdd.n321 vdd.n320 0.152939
R21921 vdd.n322 vdd.n321 0.152939
R21922 vdd.n331 vdd.n322 0.152939
R21923 vdd.n332 vdd.n331 0.152939
R21924 vdd.n333 vdd.n332 0.152939
R21925 vdd.n334 vdd.n333 0.152939
R21926 vdd.n342 vdd.n334 0.152939
R21927 vdd.n343 vdd.n342 0.152939
R21928 vdd.n344 vdd.n343 0.152939
R21929 vdd.n345 vdd.n344 0.152939
R21930 vdd.n353 vdd.n345 0.152939
R21931 vdd.n3227 vdd.n353 0.152939
R21932 vdd.n3226 vdd.n354 0.152939
R21933 vdd.n357 vdd.n354 0.152939
R21934 vdd.n361 vdd.n357 0.152939
R21935 vdd.n362 vdd.n361 0.152939
R21936 vdd.n363 vdd.n362 0.152939
R21937 vdd.n364 vdd.n363 0.152939
R21938 vdd.n365 vdd.n364 0.152939
R21939 vdd.n369 vdd.n365 0.152939
R21940 vdd.n370 vdd.n369 0.152939
R21941 vdd.n371 vdd.n370 0.152939
R21942 vdd.n372 vdd.n371 0.152939
R21943 vdd.n376 vdd.n372 0.152939
R21944 vdd.n377 vdd.n376 0.152939
R21945 vdd.n378 vdd.n377 0.152939
R21946 vdd.n379 vdd.n378 0.152939
R21947 vdd.n383 vdd.n379 0.152939
R21948 vdd.n384 vdd.n383 0.152939
R21949 vdd.n385 vdd.n384 0.152939
R21950 vdd.n3192 vdd.n385 0.152939
R21951 vdd.n3192 vdd.n3191 0.152939
R21952 vdd.n3191 vdd.n3190 0.152939
R21953 vdd.n3190 vdd.n391 0.152939
R21954 vdd.n396 vdd.n391 0.152939
R21955 vdd.n397 vdd.n396 0.152939
R21956 vdd.n398 vdd.n397 0.152939
R21957 vdd.n402 vdd.n398 0.152939
R21958 vdd.n403 vdd.n402 0.152939
R21959 vdd.n404 vdd.n403 0.152939
R21960 vdd.n405 vdd.n404 0.152939
R21961 vdd.n409 vdd.n405 0.152939
R21962 vdd.n410 vdd.n409 0.152939
R21963 vdd.n411 vdd.n410 0.152939
R21964 vdd.n412 vdd.n411 0.152939
R21965 vdd.n416 vdd.n412 0.152939
R21966 vdd.n417 vdd.n416 0.152939
R21967 vdd.n418 vdd.n417 0.152939
R21968 vdd.n419 vdd.n418 0.152939
R21969 vdd.n423 vdd.n419 0.152939
R21970 vdd.n424 vdd.n423 0.152939
R21971 vdd.n425 vdd.n424 0.152939
R21972 vdd.n3153 vdd.n425 0.152939
R21973 vdd.n3153 vdd.n3152 0.152939
R21974 vdd.n3152 vdd.n3151 0.152939
R21975 vdd.n3151 vdd.n431 0.152939
R21976 vdd.n436 vdd.n431 0.152939
R21977 vdd.n437 vdd.n436 0.152939
R21978 vdd.n438 vdd.n437 0.152939
R21979 vdd.n442 vdd.n438 0.152939
R21980 vdd.n443 vdd.n442 0.152939
R21981 vdd.n444 vdd.n443 0.152939
R21982 vdd.n445 vdd.n444 0.152939
R21983 vdd.n449 vdd.n445 0.152939
R21984 vdd.n450 vdd.n449 0.152939
R21985 vdd.n451 vdd.n450 0.152939
R21986 vdd.n452 vdd.n451 0.152939
R21987 vdd.n456 vdd.n452 0.152939
R21988 vdd.n457 vdd.n456 0.152939
R21989 vdd.n458 vdd.n457 0.152939
R21990 vdd.n459 vdd.n458 0.152939
R21991 vdd.n463 vdd.n459 0.152939
R21992 vdd.n464 vdd.n463 0.152939
R21993 vdd.n465 vdd.n464 0.152939
R21994 vdd.n3109 vdd.n465 0.152939
R21995 vdd.n3036 vdd.n3035 0.152939
R21996 vdd.n3037 vdd.n3036 0.152939
R21997 vdd.n3037 vdd.n502 0.152939
R21998 vdd.n3051 vdd.n502 0.152939
R21999 vdd.n3052 vdd.n3051 0.152939
R22000 vdd.n3053 vdd.n3052 0.152939
R22001 vdd.n3053 vdd.n489 0.152939
R22002 vdd.n3067 vdd.n489 0.152939
R22003 vdd.n3068 vdd.n3067 0.152939
R22004 vdd.n3069 vdd.n3068 0.152939
R22005 vdd.n3069 vdd.n477 0.152939
R22006 vdd.n3084 vdd.n477 0.152939
R22007 vdd.n3085 vdd.n3084 0.152939
R22008 vdd.n3086 vdd.n3085 0.152939
R22009 vdd.n3086 vdd.n475 0.152939
R22010 vdd.n3090 vdd.n475 0.152939
R22011 vdd.n3091 vdd.n3090 0.152939
R22012 vdd.n3092 vdd.n3091 0.152939
R22013 vdd.n3092 vdd.n472 0.152939
R22014 vdd.n3096 vdd.n472 0.152939
R22015 vdd.n3097 vdd.n3096 0.152939
R22016 vdd.n3098 vdd.n3097 0.152939
R22017 vdd.n3098 vdd.n469 0.152939
R22018 vdd.n3102 vdd.n469 0.152939
R22019 vdd.n3103 vdd.n3102 0.152939
R22020 vdd.n3104 vdd.n3103 0.152939
R22021 vdd.n3104 vdd.n466 0.152939
R22022 vdd.n3108 vdd.n466 0.152939
R22023 vdd.n2898 vdd.n514 0.152939
R22024 vdd.n1985 vdd.n1252 0.152939
R22025 vdd.n1581 vdd.n1580 0.152939
R22026 vdd.n1582 vdd.n1581 0.152939
R22027 vdd.n1582 vdd.n1331 0.152939
R22028 vdd.n1596 vdd.n1331 0.152939
R22029 vdd.n1597 vdd.n1596 0.152939
R22030 vdd.n1598 vdd.n1597 0.152939
R22031 vdd.n1598 vdd.n1318 0.152939
R22032 vdd.n1612 vdd.n1318 0.152939
R22033 vdd.n1613 vdd.n1612 0.152939
R22034 vdd.n1614 vdd.n1613 0.152939
R22035 vdd.n1614 vdd.n1307 0.152939
R22036 vdd.n1629 vdd.n1307 0.152939
R22037 vdd.n1630 vdd.n1629 0.152939
R22038 vdd.n1631 vdd.n1630 0.152939
R22039 vdd.n1631 vdd.n1296 0.152939
R22040 vdd.n1927 vdd.n1296 0.152939
R22041 vdd.n1928 vdd.n1927 0.152939
R22042 vdd.n1929 vdd.n1928 0.152939
R22043 vdd.n1929 vdd.n1284 0.152939
R22044 vdd.n1944 vdd.n1284 0.152939
R22045 vdd.n1945 vdd.n1944 0.152939
R22046 vdd.n1946 vdd.n1945 0.152939
R22047 vdd.n1946 vdd.n1274 0.152939
R22048 vdd.n1961 vdd.n1274 0.152939
R22049 vdd.n1962 vdd.n1961 0.152939
R22050 vdd.n1965 vdd.n1962 0.152939
R22051 vdd.n1965 vdd.n1964 0.152939
R22052 vdd.n1964 vdd.n1963 0.152939
R22053 vdd.n1573 vdd.n1347 0.152939
R22054 vdd.n1569 vdd.n1347 0.152939
R22055 vdd.n1569 vdd.n1568 0.152939
R22056 vdd.n1568 vdd.n1567 0.152939
R22057 vdd.n1567 vdd.n1352 0.152939
R22058 vdd.n1563 vdd.n1352 0.152939
R22059 vdd.n1563 vdd.n1562 0.152939
R22060 vdd.n1562 vdd.n1561 0.152939
R22061 vdd.n1561 vdd.n1360 0.152939
R22062 vdd.n1557 vdd.n1360 0.152939
R22063 vdd.n1557 vdd.n1556 0.152939
R22064 vdd.n1556 vdd.n1555 0.152939
R22065 vdd.n1555 vdd.n1368 0.152939
R22066 vdd.n1551 vdd.n1368 0.152939
R22067 vdd.n1551 vdd.n1550 0.152939
R22068 vdd.n1550 vdd.n1549 0.152939
R22069 vdd.n1549 vdd.n1376 0.152939
R22070 vdd.n1545 vdd.n1376 0.152939
R22071 vdd.n1545 vdd.n1544 0.152939
R22072 vdd.n1544 vdd.n1543 0.152939
R22073 vdd.n1543 vdd.n1386 0.152939
R22074 vdd.n1539 vdd.n1386 0.152939
R22075 vdd.n1539 vdd.n1538 0.152939
R22076 vdd.n1538 vdd.n1537 0.152939
R22077 vdd.n1537 vdd.n1394 0.152939
R22078 vdd.n1533 vdd.n1394 0.152939
R22079 vdd.n1533 vdd.n1532 0.152939
R22080 vdd.n1532 vdd.n1531 0.152939
R22081 vdd.n1531 vdd.n1402 0.152939
R22082 vdd.n1527 vdd.n1402 0.152939
R22083 vdd.n1527 vdd.n1526 0.152939
R22084 vdd.n1526 vdd.n1525 0.152939
R22085 vdd.n1525 vdd.n1410 0.152939
R22086 vdd.n1521 vdd.n1410 0.152939
R22087 vdd.n1521 vdd.n1520 0.152939
R22088 vdd.n1520 vdd.n1519 0.152939
R22089 vdd.n1519 vdd.n1418 0.152939
R22090 vdd.n1515 vdd.n1418 0.152939
R22091 vdd.n1515 vdd.n1514 0.152939
R22092 vdd.n1514 vdd.n1513 0.152939
R22093 vdd.n1513 vdd.n1426 0.152939
R22094 vdd.n1433 vdd.n1426 0.152939
R22095 vdd.n1503 vdd.n1433 0.152939
R22096 vdd.n1503 vdd.n1502 0.152939
R22097 vdd.n1502 vdd.n1501 0.152939
R22098 vdd.n1501 vdd.n1434 0.152939
R22099 vdd.n1497 vdd.n1434 0.152939
R22100 vdd.n1497 vdd.n1496 0.152939
R22101 vdd.n1496 vdd.n1495 0.152939
R22102 vdd.n1495 vdd.n1441 0.152939
R22103 vdd.n1491 vdd.n1441 0.152939
R22104 vdd.n1491 vdd.n1490 0.152939
R22105 vdd.n1490 vdd.n1489 0.152939
R22106 vdd.n1489 vdd.n1449 0.152939
R22107 vdd.n1485 vdd.n1449 0.152939
R22108 vdd.n1485 vdd.n1484 0.152939
R22109 vdd.n1484 vdd.n1483 0.152939
R22110 vdd.n1483 vdd.n1457 0.152939
R22111 vdd.n1479 vdd.n1457 0.152939
R22112 vdd.n1479 vdd.n1478 0.152939
R22113 vdd.n1478 vdd.n1477 0.152939
R22114 vdd.n1477 vdd.n1465 0.152939
R22115 vdd.n1465 vdd.n1342 0.152939
R22116 vdd.n1574 vdd.n1337 0.152939
R22117 vdd.n1588 vdd.n1337 0.152939
R22118 vdd.n1589 vdd.n1588 0.152939
R22119 vdd.n1590 vdd.n1589 0.152939
R22120 vdd.n1590 vdd.n1325 0.152939
R22121 vdd.n1604 vdd.n1325 0.152939
R22122 vdd.n1605 vdd.n1604 0.152939
R22123 vdd.n1606 vdd.n1605 0.152939
R22124 vdd.n1606 vdd.n1313 0.152939
R22125 vdd.n1621 vdd.n1313 0.152939
R22126 vdd.n1622 vdd.n1621 0.152939
R22127 vdd.n1623 vdd.n1622 0.152939
R22128 vdd.n1623 vdd.n1302 0.152939
R22129 vdd.n1920 vdd.n1919 0.145814
R22130 vdd.n3259 vdd.n310 0.145814
R22131 vdd.n3259 vdd.n311 0.145814
R22132 vdd.n1919 vdd.n1302 0.145814
R22133 vdd.n2093 vdd.n2092 0.110256
R22134 vdd.n2829 vdd.n518 0.110256
R22135 vdd.n2898 vdd.n2897 0.110256
R22136 vdd.n1986 vdd.n1985 0.110256
R22137 vdd.n2093 vdd.n948 0.0431829
R22138 vdd.n1986 vdd.n1048 0.0431829
R22139 vdd.n2829 vdd.n524 0.0431829
R22140 vdd.n2897 vdd.n605 0.0431829
R22141 vdd vdd.n28 0.00833333
R22142 a_n2848_n452.n55 a_n2848_n452.t86 533.335
R22143 a_n2848_n452.n112 a_n2848_n452.t67 512.366
R22144 a_n2848_n452.n78 a_n2848_n452.t71 512.366
R22145 a_n2848_n452.n111 a_n2848_n452.t61 512.366
R22146 a_n2848_n452.n110 a_n2848_n452.t76 512.366
R22147 a_n2848_n452.n79 a_n2848_n452.t83 512.366
R22148 a_n2848_n452.n109 a_n2848_n452.t84 512.366
R22149 a_n2848_n452.n61 a_n2848_n452.t12 533.335
R22150 a_n2848_n452.n118 a_n2848_n452.t28 512.366
R22151 a_n2848_n452.n64 a_n2848_n452.t16 512.366
R22152 a_n2848_n452.n116 a_n2848_n452.t30 512.366
R22153 a_n2848_n452.n115 a_n2848_n452.t24 512.366
R22154 a_n2848_n452.n77 a_n2848_n452.t26 512.366
R22155 a_n2848_n452.n113 a_n2848_n452.t4 512.366
R22156 a_n2848_n452.n38 a_n2848_n452.t8 533.335
R22157 a_n2848_n452.n90 a_n2848_n452.t18 512.366
R22158 a_n2848_n452.n91 a_n2848_n452.t10 512.366
R22159 a_n2848_n452.n92 a_n2848_n452.t20 512.366
R22160 a_n2848_n452.n93 a_n2848_n452.t14 512.366
R22161 a_n2848_n452.n83 a_n2848_n452.t22 512.366
R22162 a_n2848_n452.n94 a_n2848_n452.t32 512.366
R22163 a_n2848_n452.n31 a_n2848_n452.t82 533.335
R22164 a_n2848_n452.n85 a_n2848_n452.t60 512.366
R22165 a_n2848_n452.n86 a_n2848_n452.t79 512.366
R22166 a_n2848_n452.n87 a_n2848_n452.t80 512.366
R22167 a_n2848_n452.n88 a_n2848_n452.t57 512.366
R22168 a_n2848_n452.n84 a_n2848_n452.t66 512.366
R22169 a_n2848_n452.n89 a_n2848_n452.t75 512.366
R22170 a_n2848_n452.n106 a_n2848_n452.t73 512.366
R22171 a_n2848_n452.n96 a_n2848_n452.t64 512.366
R22172 a_n2848_n452.n107 a_n2848_n452.t56 512.366
R22173 a_n2848_n452.n104 a_n2848_n452.t81 512.366
R22174 a_n2848_n452.n97 a_n2848_n452.t70 512.366
R22175 a_n2848_n452.n105 a_n2848_n452.t69 512.366
R22176 a_n2848_n452.n102 a_n2848_n452.t77 512.366
R22177 a_n2848_n452.n98 a_n2848_n452.t62 512.366
R22178 a_n2848_n452.n103 a_n2848_n452.t63 512.366
R22179 a_n2848_n452.n100 a_n2848_n452.t65 512.366
R22180 a_n2848_n452.n99 a_n2848_n452.t74 512.366
R22181 a_n2848_n452.n101 a_n2848_n452.t87 512.366
R22182 a_n2848_n452.n60 a_n2848_n452.n8 70.1674
R22183 a_n2848_n452.n54 a_n2848_n452.n11 70.1674
R22184 a_n2848_n452.n21 a_n2848_n452.n44 70.1674
R22185 a_n2848_n452.n24 a_n2848_n452.n37 70.1674
R22186 a_n2848_n452.n89 a_n2848_n452.n37 20.9683
R22187 a_n2848_n452.n36 a_n2848_n452.n25 72.3034
R22188 a_n2848_n452.n36 a_n2848_n452.n84 16.6962
R22189 a_n2848_n452.n25 a_n2848_n452.n35 77.6622
R22190 a_n2848_n452.n88 a_n2848_n452.n35 5.97853
R22191 a_n2848_n452.n34 a_n2848_n452.n26 77.6622
R22192 a_n2848_n452.n26 a_n2848_n452.n33 72.3034
R22193 a_n2848_n452.n85 a_n2848_n452.n31 20.9683
R22194 a_n2848_n452.n32 a_n2848_n452.n31 70.1674
R22195 a_n2848_n452.n94 a_n2848_n452.n44 20.9683
R22196 a_n2848_n452.n43 a_n2848_n452.n22 72.3034
R22197 a_n2848_n452.n43 a_n2848_n452.n83 16.6962
R22198 a_n2848_n452.n22 a_n2848_n452.n42 77.6622
R22199 a_n2848_n452.n93 a_n2848_n452.n42 5.97853
R22200 a_n2848_n452.n41 a_n2848_n452.n23 77.6622
R22201 a_n2848_n452.n23 a_n2848_n452.n40 72.3034
R22202 a_n2848_n452.n90 a_n2848_n452.n38 20.9683
R22203 a_n2848_n452.n39 a_n2848_n452.n38 70.1674
R22204 a_n2848_n452.n12 a_n2848_n452.n52 70.1674
R22205 a_n2848_n452.n14 a_n2848_n452.n50 70.1674
R22206 a_n2848_n452.n16 a_n2848_n452.n48 70.1674
R22207 a_n2848_n452.n19 a_n2848_n452.n46 70.1674
R22208 a_n2848_n452.n101 a_n2848_n452.n46 20.9683
R22209 a_n2848_n452.n45 a_n2848_n452.n20 75.0448
R22210 a_n2848_n452.n45 a_n2848_n452.n99 11.2134
R22211 a_n2848_n452.n20 a_n2848_n452.n100 161.3
R22212 a_n2848_n452.n103 a_n2848_n452.n48 20.9683
R22213 a_n2848_n452.n47 a_n2848_n452.n17 75.0448
R22214 a_n2848_n452.n47 a_n2848_n452.n98 11.2134
R22215 a_n2848_n452.n17 a_n2848_n452.n102 161.3
R22216 a_n2848_n452.n105 a_n2848_n452.n50 20.9683
R22217 a_n2848_n452.n49 a_n2848_n452.n15 75.0448
R22218 a_n2848_n452.n49 a_n2848_n452.n97 11.2134
R22219 a_n2848_n452.n15 a_n2848_n452.n104 161.3
R22220 a_n2848_n452.n107 a_n2848_n452.n52 20.9683
R22221 a_n2848_n452.n51 a_n2848_n452.n13 75.0448
R22222 a_n2848_n452.n51 a_n2848_n452.n96 11.2134
R22223 a_n2848_n452.n13 a_n2848_n452.n106 161.3
R22224 a_n2848_n452.n113 a_n2848_n452.n54 20.9683
R22225 a_n2848_n452.n11 a_n2848_n452.n53 72.3034
R22226 a_n2848_n452.n53 a_n2848_n452.n77 16.6962
R22227 a_n2848_n452.n114 a_n2848_n452.n6 161.3
R22228 a_n2848_n452.n109 a_n2848_n452.n60 20.9683
R22229 a_n2848_n452.n9 a_n2848_n452.n59 72.3034
R22230 a_n2848_n452.n59 a_n2848_n452.n79 16.6962
R22231 a_n2848_n452.n58 a_n2848_n452.n9 77.6622
R22232 a_n2848_n452.n110 a_n2848_n452.n58 5.97853
R22233 a_n2848_n452.n57 a_n2848_n452.n7 77.6622
R22234 a_n2848_n452.n7 a_n2848_n452.n56 72.3034
R22235 a_n2848_n452.n112 a_n2848_n452.n55 20.9683
R22236 a_n2848_n452.n10 a_n2848_n452.n55 70.1674
R22237 a_n2848_n452.n115 a_n2848_n452.n63 20.9683
R22238 a_n2848_n452.n63 a_n2848_n452.n6 70.1674
R22239 a_n2848_n452.n6 a_n2848_n452.n117 161.3
R22240 a_n2848_n452.n6 a_n2848_n452.n62 72.3034
R22241 a_n2848_n452.n118 a_n2848_n452.n61 20.9683
R22242 a_n2848_n452.n5 a_n2848_n452.n61 70.1674
R22243 a_n2848_n452.n3 a_n2848_n452.n74 81.4626
R22244 a_n2848_n452.n4 a_n2848_n452.n68 81.4626
R22245 a_n2848_n452.n0 a_n2848_n452.n65 81.4626
R22246 a_n2848_n452.n3 a_n2848_n452.n75 80.9324
R22247 a_n2848_n452.n2 a_n2848_n452.n76 80.9324
R22248 a_n2848_n452.n2 a_n2848_n452.n73 80.9324
R22249 a_n2848_n452.n2 a_n2848_n452.n72 80.9324
R22250 a_n2848_n452.n1 a_n2848_n452.n71 80.9324
R22251 a_n2848_n452.n4 a_n2848_n452.n69 80.9324
R22252 a_n2848_n452.n0 a_n2848_n452.n70 80.9324
R22253 a_n2848_n452.n0 a_n2848_n452.n67 80.9324
R22254 a_n2848_n452.n0 a_n2848_n452.n66 80.9324
R22255 a_n2848_n452.n27 a_n2848_n452.t9 74.6477
R22256 a_n2848_n452.t3 a_n2848_n452.n30 74.6477
R22257 a_n2848_n452.n29 a_n2848_n452.t13 74.2899
R22258 a_n2848_n452.n28 a_n2848_n452.t7 74.2897
R22259 a_n2848_n452.n30 a_n2848_n452.n122 70.6783
R22260 a_n2848_n452.n30 a_n2848_n452.n121 70.6783
R22261 a_n2848_n452.n29 a_n2848_n452.n120 70.6783
R22262 a_n2848_n452.n28 a_n2848_n452.n82 70.6783
R22263 a_n2848_n452.n27 a_n2848_n452.n81 70.6783
R22264 a_n2848_n452.n27 a_n2848_n452.n80 70.6783
R22265 a_n2848_n452.n111 a_n2848_n452.n110 48.2005
R22266 a_n2848_n452.n60 a_n2848_n452.t58 533.335
R22267 a_n2848_n452.n116 a_n2848_n452.n63 20.9683
R22268 a_n2848_n452.n54 a_n2848_n452.t2 533.335
R22269 a_n2848_n452.n93 a_n2848_n452.n92 48.2005
R22270 a_n2848_n452.t6 a_n2848_n452.n44 533.335
R22271 a_n2848_n452.n88 a_n2848_n452.n87 48.2005
R22272 a_n2848_n452.t59 a_n2848_n452.n37 533.335
R22273 a_n2848_n452.n106 a_n2848_n452.n96 48.2005
R22274 a_n2848_n452.t78 a_n2848_n452.n52 533.335
R22275 a_n2848_n452.n104 a_n2848_n452.n97 48.2005
R22276 a_n2848_n452.t85 a_n2848_n452.n50 533.335
R22277 a_n2848_n452.n102 a_n2848_n452.n98 48.2005
R22278 a_n2848_n452.t72 a_n2848_n452.n48 533.335
R22279 a_n2848_n452.n100 a_n2848_n452.n99 48.2005
R22280 a_n2848_n452.t68 a_n2848_n452.n46 533.335
R22281 a_n2848_n452.n56 a_n2848_n452.n78 16.6962
R22282 a_n2848_n452.n109 a_n2848_n452.n59 27.6507
R22283 a_n2848_n452.n62 a_n2848_n452.n64 16.6962
R22284 a_n2848_n452.n113 a_n2848_n452.n53 27.6507
R22285 a_n2848_n452.n91 a_n2848_n452.n40 16.6962
R22286 a_n2848_n452.n94 a_n2848_n452.n43 27.6507
R22287 a_n2848_n452.n86 a_n2848_n452.n33 16.6962
R22288 a_n2848_n452.n89 a_n2848_n452.n36 27.6507
R22289 a_n2848_n452.n57 a_n2848_n452.n78 41.7634
R22290 a_n2848_n452.n117 a_n2848_n452.n64 35.7853
R22291 a_n2848_n452.n114 a_n2848_n452.n77 35.7853
R22292 a_n2848_n452.n91 a_n2848_n452.n41 41.7634
R22293 a_n2848_n452.n86 a_n2848_n452.n34 41.7634
R22294 a_n2848_n452.n1 a_n2848_n452.n0 33.585
R22295 a_n2848_n452.n107 a_n2848_n452.n51 35.3134
R22296 a_n2848_n452.n105 a_n2848_n452.n49 35.3134
R22297 a_n2848_n452.n103 a_n2848_n452.n47 35.3134
R22298 a_n2848_n452.n101 a_n2848_n452.n45 35.3134
R22299 a_n2848_n452.n6 a_n2848_n452.n2 23.891
R22300 a_n2848_n452.n32 a_n2848_n452.n18 12.705
R22301 a_n2848_n452.n8 a_n2848_n452.n108 12.5005
R22302 a_n2848_n452.n57 a_n2848_n452.n111 5.97853
R22303 a_n2848_n452.n58 a_n2848_n452.n79 41.7634
R22304 a_n2848_n452.n117 a_n2848_n452.n116 12.4157
R22305 a_n2848_n452.n115 a_n2848_n452.n114 12.4157
R22306 a_n2848_n452.n92 a_n2848_n452.n41 5.97853
R22307 a_n2848_n452.n83 a_n2848_n452.n42 41.7634
R22308 a_n2848_n452.n87 a_n2848_n452.n34 5.97853
R22309 a_n2848_n452.n84 a_n2848_n452.n35 41.7634
R22310 a_n2848_n452.n119 a_n2848_n452.n5 11.1956
R22311 a_n2848_n452.n112 a_n2848_n452.n56 27.6507
R22312 a_n2848_n452.n118 a_n2848_n452.n62 27.6507
R22313 a_n2848_n452.n40 a_n2848_n452.n90 27.6507
R22314 a_n2848_n452.n33 a_n2848_n452.n85 27.6507
R22315 a_n2848_n452.n95 a_n2848_n452.n28 9.85898
R22316 a_n2848_n452.n20 a_n2848_n452.n18 8.73345
R22317 a_n2848_n452.n108 a_n2848_n452.n12 8.73345
R22318 a_n2848_n452.n95 a_n2848_n452.n21 7.36035
R22319 a_n2848_n452.n29 a_n2848_n452.n119 6.01559
R22320 a_n2848_n452.n108 a_n2848_n452.n95 5.3452
R22321 a_n2848_n452.n39 a_n2848_n452.n24 4.01186
R22322 a_n2848_n452.n11 a_n2848_n452.n10 4.01186
R22323 a_n2848_n452.n122 a_n2848_n452.t27 3.61217
R22324 a_n2848_n452.n122 a_n2848_n452.t5 3.61217
R22325 a_n2848_n452.n121 a_n2848_n452.t31 3.61217
R22326 a_n2848_n452.n121 a_n2848_n452.t25 3.61217
R22327 a_n2848_n452.n120 a_n2848_n452.t29 3.61217
R22328 a_n2848_n452.n120 a_n2848_n452.t17 3.61217
R22329 a_n2848_n452.n82 a_n2848_n452.t23 3.61217
R22330 a_n2848_n452.n82 a_n2848_n452.t33 3.61217
R22331 a_n2848_n452.n81 a_n2848_n452.t21 3.61217
R22332 a_n2848_n452.n81 a_n2848_n452.t15 3.61217
R22333 a_n2848_n452.n80 a_n2848_n452.t19 3.61217
R22334 a_n2848_n452.n80 a_n2848_n452.t11 3.61217
R22335 a_n2848_n452.n74 a_n2848_n452.t55 2.82907
R22336 a_n2848_n452.n74 a_n2848_n452.t39 2.82907
R22337 a_n2848_n452.n75 a_n2848_n452.t35 2.82907
R22338 a_n2848_n452.n75 a_n2848_n452.t48 2.82907
R22339 a_n2848_n452.n76 a_n2848_n452.t44 2.82907
R22340 a_n2848_n452.n76 a_n2848_n452.t45 2.82907
R22341 a_n2848_n452.n73 a_n2848_n452.t53 2.82907
R22342 a_n2848_n452.n73 a_n2848_n452.t36 2.82907
R22343 a_n2848_n452.n72 a_n2848_n452.t41 2.82907
R22344 a_n2848_n452.n72 a_n2848_n452.t0 2.82907
R22345 a_n2848_n452.n71 a_n2848_n452.t43 2.82907
R22346 a_n2848_n452.n71 a_n2848_n452.t51 2.82907
R22347 a_n2848_n452.n68 a_n2848_n452.t50 2.82907
R22348 a_n2848_n452.n68 a_n2848_n452.t47 2.82907
R22349 a_n2848_n452.n69 a_n2848_n452.t54 2.82907
R22350 a_n2848_n452.n69 a_n2848_n452.t52 2.82907
R22351 a_n2848_n452.n70 a_n2848_n452.t38 2.82907
R22352 a_n2848_n452.n70 a_n2848_n452.t40 2.82907
R22353 a_n2848_n452.n67 a_n2848_n452.t37 2.82907
R22354 a_n2848_n452.n67 a_n2848_n452.t1 2.82907
R22355 a_n2848_n452.n66 a_n2848_n452.t42 2.82907
R22356 a_n2848_n452.n66 a_n2848_n452.t46 2.82907
R22357 a_n2848_n452.n65 a_n2848_n452.t34 2.82907
R22358 a_n2848_n452.n65 a_n2848_n452.t49 2.82907
R22359 a_n2848_n452.n0 a_n2848_n452.n4 1.59102
R22360 a_n2848_n452.n119 a_n2848_n452.n18 1.30542
R22361 a_n2848_n452.n6 a_n2848_n452.n11 1.09898
R22362 a_n2848_n452.n30 a_n2848_n452.n29 1.07378
R22363 a_n2848_n452.n28 a_n2848_n452.n27 1.07378
R22364 a_n2848_n452.n2 a_n2848_n452.n3 1.06084
R22365 a_n2848_n452.n2 a_n2848_n452.n1 1.06084
R22366 a_n2848_n452.n15 a_n2848_n452.n16 1.04595
R22367 a_n2848_n452.n6 a_n2848_n452.n5 0.94747
R22368 a_n2848_n452.n26 a_n2848_n452.n25 0.758076
R22369 a_n2848_n452.n25 a_n2848_n452.n24 0.758076
R22370 a_n2848_n452.n23 a_n2848_n452.n22 0.758076
R22371 a_n2848_n452.n22 a_n2848_n452.n21 0.758076
R22372 a_n2848_n452.n20 a_n2848_n452.n19 0.758076
R22373 a_n2848_n452.n17 a_n2848_n452.n16 0.758076
R22374 a_n2848_n452.n15 a_n2848_n452.n14 0.758076
R22375 a_n2848_n452.n13 a_n2848_n452.n12 0.758076
R22376 a_n2848_n452.n9 a_n2848_n452.n7 0.758076
R22377 a_n2848_n452.n9 a_n2848_n452.n8 0.758076
R22378 a_n2848_n452.n17 a_n2848_n452.n19 0.67853
R22379 a_n2848_n452.n13 a_n2848_n452.n14 0.67853
R22380 a_n2848_n452.n7 a_n2848_n452.n10 0.568682
R22381 a_n2848_n452.n39 a_n2848_n452.n23 0.568682
R22382 a_n2848_n452.n32 a_n2848_n452.n26 0.568682
R22383 a_n2140_13878.n2 a_n2140_13878.n0 98.9633
R22384 a_n2140_13878.n5 a_n2140_13878.n3 98.7517
R22385 a_n2140_13878.n2 a_n2140_13878.n1 98.6055
R22386 a_n2140_13878.n9 a_n2140_13878.n8 98.6055
R22387 a_n2140_13878.n7 a_n2140_13878.n6 98.6055
R22388 a_n2140_13878.n5 a_n2140_13878.n4 98.6055
R22389 a_n2140_13878.n21 a_n2140_13878.n20 98.6054
R22390 a_n2140_13878.n19 a_n2140_13878.n18 98.6054
R22391 a_n2140_13878.n11 a_n2140_13878.t1 74.6477
R22392 a_n2140_13878.n16 a_n2140_13878.t2 74.2899
R22393 a_n2140_13878.n13 a_n2140_13878.t3 74.2899
R22394 a_n2140_13878.n12 a_n2140_13878.t0 74.2899
R22395 a_n2140_13878.n15 a_n2140_13878.n14 70.6783
R22396 a_n2140_13878.n11 a_n2140_13878.n10 70.6783
R22397 a_n2140_13878.n17 a_n2140_13878.n9 14.2849
R22398 a_n2140_13878.n19 a_n2140_13878.n17 11.9339
R22399 a_n2140_13878.n17 a_n2140_13878.n16 6.95632
R22400 a_n2140_13878.n18 a_n2140_13878.t14 3.61217
R22401 a_n2140_13878.n18 a_n2140_13878.t15 3.61217
R22402 a_n2140_13878.n1 a_n2140_13878.t8 3.61217
R22403 a_n2140_13878.n1 a_n2140_13878.t16 3.61217
R22404 a_n2140_13878.n0 a_n2140_13878.t19 3.61217
R22405 a_n2140_13878.n0 a_n2140_13878.t23 3.61217
R22406 a_n2140_13878.n14 a_n2140_13878.t6 3.61217
R22407 a_n2140_13878.n14 a_n2140_13878.t7 3.61217
R22408 a_n2140_13878.n10 a_n2140_13878.t4 3.61217
R22409 a_n2140_13878.n10 a_n2140_13878.t5 3.61217
R22410 a_n2140_13878.n8 a_n2140_13878.t17 3.61217
R22411 a_n2140_13878.n8 a_n2140_13878.t9 3.61217
R22412 a_n2140_13878.n6 a_n2140_13878.t20 3.61217
R22413 a_n2140_13878.n6 a_n2140_13878.t11 3.61217
R22414 a_n2140_13878.n4 a_n2140_13878.t10 3.61217
R22415 a_n2140_13878.n4 a_n2140_13878.t12 3.61217
R22416 a_n2140_13878.n3 a_n2140_13878.t18 3.61217
R22417 a_n2140_13878.n3 a_n2140_13878.t13 3.61217
R22418 a_n2140_13878.n21 a_n2140_13878.t21 3.61217
R22419 a_n2140_13878.t22 a_n2140_13878.n21 3.61217
R22420 a_n2140_13878.n12 a_n2140_13878.n11 0.358259
R22421 a_n2140_13878.n15 a_n2140_13878.n13 0.358259
R22422 a_n2140_13878.n16 a_n2140_13878.n15 0.358259
R22423 a_n2140_13878.n20 a_n2140_13878.n2 0.358259
R22424 a_n2140_13878.n20 a_n2140_13878.n19 0.358259
R22425 a_n2140_13878.n7 a_n2140_13878.n5 0.146627
R22426 a_n2140_13878.n9 a_n2140_13878.n7 0.146627
R22427 a_n2140_13878.n13 a_n2140_13878.n12 0.101793
R22428 outputibias.n27 outputibias.n1 289.615
R22429 outputibias.n58 outputibias.n32 289.615
R22430 outputibias.n90 outputibias.n64 289.615
R22431 outputibias.n122 outputibias.n96 289.615
R22432 outputibias.n28 outputibias.n27 185
R22433 outputibias.n26 outputibias.n25 185
R22434 outputibias.n5 outputibias.n4 185
R22435 outputibias.n20 outputibias.n19 185
R22436 outputibias.n18 outputibias.n17 185
R22437 outputibias.n9 outputibias.n8 185
R22438 outputibias.n12 outputibias.n11 185
R22439 outputibias.n59 outputibias.n58 185
R22440 outputibias.n57 outputibias.n56 185
R22441 outputibias.n36 outputibias.n35 185
R22442 outputibias.n51 outputibias.n50 185
R22443 outputibias.n49 outputibias.n48 185
R22444 outputibias.n40 outputibias.n39 185
R22445 outputibias.n43 outputibias.n42 185
R22446 outputibias.n91 outputibias.n90 185
R22447 outputibias.n89 outputibias.n88 185
R22448 outputibias.n68 outputibias.n67 185
R22449 outputibias.n83 outputibias.n82 185
R22450 outputibias.n81 outputibias.n80 185
R22451 outputibias.n72 outputibias.n71 185
R22452 outputibias.n75 outputibias.n74 185
R22453 outputibias.n123 outputibias.n122 185
R22454 outputibias.n121 outputibias.n120 185
R22455 outputibias.n100 outputibias.n99 185
R22456 outputibias.n115 outputibias.n114 185
R22457 outputibias.n113 outputibias.n112 185
R22458 outputibias.n104 outputibias.n103 185
R22459 outputibias.n107 outputibias.n106 185
R22460 outputibias.n0 outputibias.t9 178.945
R22461 outputibias.n133 outputibias.t10 177.018
R22462 outputibias.n132 outputibias.t11 177.018
R22463 outputibias.n0 outputibias.t8 177.018
R22464 outputibias.t7 outputibias.n10 147.661
R22465 outputibias.t1 outputibias.n41 147.661
R22466 outputibias.t3 outputibias.n73 147.661
R22467 outputibias.t5 outputibias.n105 147.661
R22468 outputibias.n128 outputibias.t6 132.363
R22469 outputibias.n128 outputibias.t0 130.436
R22470 outputibias.n129 outputibias.t2 130.436
R22471 outputibias.n130 outputibias.t4 130.436
R22472 outputibias.n27 outputibias.n26 104.615
R22473 outputibias.n26 outputibias.n4 104.615
R22474 outputibias.n19 outputibias.n4 104.615
R22475 outputibias.n19 outputibias.n18 104.615
R22476 outputibias.n18 outputibias.n8 104.615
R22477 outputibias.n11 outputibias.n8 104.615
R22478 outputibias.n58 outputibias.n57 104.615
R22479 outputibias.n57 outputibias.n35 104.615
R22480 outputibias.n50 outputibias.n35 104.615
R22481 outputibias.n50 outputibias.n49 104.615
R22482 outputibias.n49 outputibias.n39 104.615
R22483 outputibias.n42 outputibias.n39 104.615
R22484 outputibias.n90 outputibias.n89 104.615
R22485 outputibias.n89 outputibias.n67 104.615
R22486 outputibias.n82 outputibias.n67 104.615
R22487 outputibias.n82 outputibias.n81 104.615
R22488 outputibias.n81 outputibias.n71 104.615
R22489 outputibias.n74 outputibias.n71 104.615
R22490 outputibias.n122 outputibias.n121 104.615
R22491 outputibias.n121 outputibias.n99 104.615
R22492 outputibias.n114 outputibias.n99 104.615
R22493 outputibias.n114 outputibias.n113 104.615
R22494 outputibias.n113 outputibias.n103 104.615
R22495 outputibias.n106 outputibias.n103 104.615
R22496 outputibias.n63 outputibias.n31 95.6354
R22497 outputibias.n63 outputibias.n62 94.6732
R22498 outputibias.n95 outputibias.n94 94.6732
R22499 outputibias.n127 outputibias.n126 94.6732
R22500 outputibias.n11 outputibias.t7 52.3082
R22501 outputibias.n42 outputibias.t1 52.3082
R22502 outputibias.n74 outputibias.t3 52.3082
R22503 outputibias.n106 outputibias.t5 52.3082
R22504 outputibias.n12 outputibias.n10 15.6674
R22505 outputibias.n43 outputibias.n41 15.6674
R22506 outputibias.n75 outputibias.n73 15.6674
R22507 outputibias.n107 outputibias.n105 15.6674
R22508 outputibias.n13 outputibias.n9 12.8005
R22509 outputibias.n44 outputibias.n40 12.8005
R22510 outputibias.n76 outputibias.n72 12.8005
R22511 outputibias.n108 outputibias.n104 12.8005
R22512 outputibias.n17 outputibias.n16 12.0247
R22513 outputibias.n48 outputibias.n47 12.0247
R22514 outputibias.n80 outputibias.n79 12.0247
R22515 outputibias.n112 outputibias.n111 12.0247
R22516 outputibias.n20 outputibias.n7 11.249
R22517 outputibias.n51 outputibias.n38 11.249
R22518 outputibias.n83 outputibias.n70 11.249
R22519 outputibias.n115 outputibias.n102 11.249
R22520 outputibias.n21 outputibias.n5 10.4732
R22521 outputibias.n52 outputibias.n36 10.4732
R22522 outputibias.n84 outputibias.n68 10.4732
R22523 outputibias.n116 outputibias.n100 10.4732
R22524 outputibias.n25 outputibias.n24 9.69747
R22525 outputibias.n56 outputibias.n55 9.69747
R22526 outputibias.n88 outputibias.n87 9.69747
R22527 outputibias.n120 outputibias.n119 9.69747
R22528 outputibias.n31 outputibias.n30 9.45567
R22529 outputibias.n62 outputibias.n61 9.45567
R22530 outputibias.n94 outputibias.n93 9.45567
R22531 outputibias.n126 outputibias.n125 9.45567
R22532 outputibias.n30 outputibias.n29 9.3005
R22533 outputibias.n3 outputibias.n2 9.3005
R22534 outputibias.n24 outputibias.n23 9.3005
R22535 outputibias.n22 outputibias.n21 9.3005
R22536 outputibias.n7 outputibias.n6 9.3005
R22537 outputibias.n16 outputibias.n15 9.3005
R22538 outputibias.n14 outputibias.n13 9.3005
R22539 outputibias.n61 outputibias.n60 9.3005
R22540 outputibias.n34 outputibias.n33 9.3005
R22541 outputibias.n55 outputibias.n54 9.3005
R22542 outputibias.n53 outputibias.n52 9.3005
R22543 outputibias.n38 outputibias.n37 9.3005
R22544 outputibias.n47 outputibias.n46 9.3005
R22545 outputibias.n45 outputibias.n44 9.3005
R22546 outputibias.n93 outputibias.n92 9.3005
R22547 outputibias.n66 outputibias.n65 9.3005
R22548 outputibias.n87 outputibias.n86 9.3005
R22549 outputibias.n85 outputibias.n84 9.3005
R22550 outputibias.n70 outputibias.n69 9.3005
R22551 outputibias.n79 outputibias.n78 9.3005
R22552 outputibias.n77 outputibias.n76 9.3005
R22553 outputibias.n125 outputibias.n124 9.3005
R22554 outputibias.n98 outputibias.n97 9.3005
R22555 outputibias.n119 outputibias.n118 9.3005
R22556 outputibias.n117 outputibias.n116 9.3005
R22557 outputibias.n102 outputibias.n101 9.3005
R22558 outputibias.n111 outputibias.n110 9.3005
R22559 outputibias.n109 outputibias.n108 9.3005
R22560 outputibias.n28 outputibias.n3 8.92171
R22561 outputibias.n59 outputibias.n34 8.92171
R22562 outputibias.n91 outputibias.n66 8.92171
R22563 outputibias.n123 outputibias.n98 8.92171
R22564 outputibias.n29 outputibias.n1 8.14595
R22565 outputibias.n60 outputibias.n32 8.14595
R22566 outputibias.n92 outputibias.n64 8.14595
R22567 outputibias.n124 outputibias.n96 8.14595
R22568 outputibias.n31 outputibias.n1 5.81868
R22569 outputibias.n62 outputibias.n32 5.81868
R22570 outputibias.n94 outputibias.n64 5.81868
R22571 outputibias.n126 outputibias.n96 5.81868
R22572 outputibias.n131 outputibias.n130 5.20947
R22573 outputibias.n29 outputibias.n28 5.04292
R22574 outputibias.n60 outputibias.n59 5.04292
R22575 outputibias.n92 outputibias.n91 5.04292
R22576 outputibias.n124 outputibias.n123 5.04292
R22577 outputibias.n131 outputibias.n127 4.42209
R22578 outputibias.n14 outputibias.n10 4.38594
R22579 outputibias.n45 outputibias.n41 4.38594
R22580 outputibias.n77 outputibias.n73 4.38594
R22581 outputibias.n109 outputibias.n105 4.38594
R22582 outputibias.n132 outputibias.n131 4.28454
R22583 outputibias.n25 outputibias.n3 4.26717
R22584 outputibias.n56 outputibias.n34 4.26717
R22585 outputibias.n88 outputibias.n66 4.26717
R22586 outputibias.n120 outputibias.n98 4.26717
R22587 outputibias.n24 outputibias.n5 3.49141
R22588 outputibias.n55 outputibias.n36 3.49141
R22589 outputibias.n87 outputibias.n68 3.49141
R22590 outputibias.n119 outputibias.n100 3.49141
R22591 outputibias.n21 outputibias.n20 2.71565
R22592 outputibias.n52 outputibias.n51 2.71565
R22593 outputibias.n84 outputibias.n83 2.71565
R22594 outputibias.n116 outputibias.n115 2.71565
R22595 outputibias.n17 outputibias.n7 1.93989
R22596 outputibias.n48 outputibias.n38 1.93989
R22597 outputibias.n80 outputibias.n70 1.93989
R22598 outputibias.n112 outputibias.n102 1.93989
R22599 outputibias.n130 outputibias.n129 1.9266
R22600 outputibias.n129 outputibias.n128 1.9266
R22601 outputibias.n133 outputibias.n132 1.92658
R22602 outputibias.n134 outputibias.n133 1.29913
R22603 outputibias.n16 outputibias.n9 1.16414
R22604 outputibias.n47 outputibias.n40 1.16414
R22605 outputibias.n79 outputibias.n72 1.16414
R22606 outputibias.n111 outputibias.n104 1.16414
R22607 outputibias.n127 outputibias.n95 0.962709
R22608 outputibias.n95 outputibias.n63 0.962709
R22609 outputibias.n13 outputibias.n12 0.388379
R22610 outputibias.n44 outputibias.n43 0.388379
R22611 outputibias.n76 outputibias.n75 0.388379
R22612 outputibias.n108 outputibias.n107 0.388379
R22613 outputibias.n134 outputibias.n0 0.337251
R22614 outputibias outputibias.n134 0.302375
R22615 outputibias.n30 outputibias.n2 0.155672
R22616 outputibias.n23 outputibias.n2 0.155672
R22617 outputibias.n23 outputibias.n22 0.155672
R22618 outputibias.n22 outputibias.n6 0.155672
R22619 outputibias.n15 outputibias.n6 0.155672
R22620 outputibias.n15 outputibias.n14 0.155672
R22621 outputibias.n61 outputibias.n33 0.155672
R22622 outputibias.n54 outputibias.n33 0.155672
R22623 outputibias.n54 outputibias.n53 0.155672
R22624 outputibias.n53 outputibias.n37 0.155672
R22625 outputibias.n46 outputibias.n37 0.155672
R22626 outputibias.n46 outputibias.n45 0.155672
R22627 outputibias.n93 outputibias.n65 0.155672
R22628 outputibias.n86 outputibias.n65 0.155672
R22629 outputibias.n86 outputibias.n85 0.155672
R22630 outputibias.n85 outputibias.n69 0.155672
R22631 outputibias.n78 outputibias.n69 0.155672
R22632 outputibias.n78 outputibias.n77 0.155672
R22633 outputibias.n125 outputibias.n97 0.155672
R22634 outputibias.n118 outputibias.n97 0.155672
R22635 outputibias.n118 outputibias.n117 0.155672
R22636 outputibias.n117 outputibias.n101 0.155672
R22637 outputibias.n110 outputibias.n101 0.155672
R22638 outputibias.n110 outputibias.n109 0.155672
R22639 plus.n76 plus.t11 250.337
R22640 plus.n15 plus.t14 250.337
R22641 plus.n124 plus.t1 243.97
R22642 plus.n120 plus.t24 231.093
R22643 plus.n59 plus.t20 231.093
R22644 plus.n124 plus.n123 223.454
R22645 plus.n126 plus.n125 223.454
R22646 plus.n77 plus.t5 187.445
R22647 plus.n74 plus.t22 187.445
R22648 plus.n72 plus.t21 187.445
R22649 plus.n89 plus.t16 187.445
R22650 plus.n95 plus.t17 187.445
R22651 plus.n68 plus.t13 187.445
R22652 plus.n66 plus.t15 187.445
R22653 plus.n107 plus.t10 187.445
R22654 plus.n113 plus.t26 187.445
R22655 plus.n62 plus.t28 187.445
R22656 plus.n1 plus.t23 187.445
R22657 plus.n52 plus.t6 187.445
R22658 plus.n46 plus.t12 187.445
R22659 plus.n5 plus.t8 187.445
R22660 plus.n7 plus.t7 187.445
R22661 plus.n34 plus.t19 187.445
R22662 plus.n28 plus.t18 187.445
R22663 plus.n11 plus.t27 187.445
R22664 plus.n13 plus.t25 187.445
R22665 plus.n16 plus.t9 187.445
R22666 plus.n121 plus.n120 161.3
R22667 plus.n119 plus.n61 161.3
R22668 plus.n118 plus.n117 161.3
R22669 plus.n116 plus.n115 161.3
R22670 plus.n114 plus.n63 161.3
R22671 plus.n112 plus.n111 161.3
R22672 plus.n110 plus.n64 161.3
R22673 plus.n109 plus.n108 161.3
R22674 plus.n106 plus.n65 161.3
R22675 plus.n105 plus.n104 161.3
R22676 plus.n103 plus.n102 161.3
R22677 plus.n101 plus.n67 161.3
R22678 plus.n100 plus.n99 161.3
R22679 plus.n98 plus.n97 161.3
R22680 plus.n96 plus.n69 161.3
R22681 plus.n94 plus.n93 161.3
R22682 plus.n92 plus.n70 161.3
R22683 plus.n91 plus.n90 161.3
R22684 plus.n88 plus.n71 161.3
R22685 plus.n87 plus.n86 161.3
R22686 plus.n85 plus.n84 161.3
R22687 plus.n83 plus.n73 161.3
R22688 plus.n82 plus.n81 161.3
R22689 plus.n80 plus.n79 161.3
R22690 plus.n78 plus.n75 161.3
R22691 plus.n17 plus.n14 161.3
R22692 plus.n19 plus.n18 161.3
R22693 plus.n21 plus.n20 161.3
R22694 plus.n22 plus.n12 161.3
R22695 plus.n24 plus.n23 161.3
R22696 plus.n26 plus.n25 161.3
R22697 plus.n27 plus.n10 161.3
R22698 plus.n30 plus.n29 161.3
R22699 plus.n31 plus.n9 161.3
R22700 plus.n33 plus.n32 161.3
R22701 plus.n35 plus.n8 161.3
R22702 plus.n37 plus.n36 161.3
R22703 plus.n39 plus.n38 161.3
R22704 plus.n40 plus.n6 161.3
R22705 plus.n42 plus.n41 161.3
R22706 plus.n44 plus.n43 161.3
R22707 plus.n45 plus.n4 161.3
R22708 plus.n48 plus.n47 161.3
R22709 plus.n49 plus.n3 161.3
R22710 plus.n51 plus.n50 161.3
R22711 plus.n53 plus.n2 161.3
R22712 plus.n55 plus.n54 161.3
R22713 plus.n57 plus.n56 161.3
R22714 plus.n58 plus.n0 161.3
R22715 plus.n60 plus.n59 161.3
R22716 plus.n88 plus.n87 56.5617
R22717 plus.n97 plus.n96 56.5617
R22718 plus.n106 plus.n105 56.5617
R22719 plus.n45 plus.n44 56.5617
R22720 plus.n36 plus.n35 56.5617
R22721 plus.n27 plus.n26 56.5617
R22722 plus.n79 plus.n78 56.5617
R22723 plus.n115 plus.n114 56.5617
R22724 plus.n54 plus.n53 56.5617
R22725 plus.n18 plus.n17 56.5617
R22726 plus.n119 plus.n118 50.2647
R22727 plus.n58 plus.n57 50.2647
R22728 plus.n84 plus.n83 46.3896
R22729 plus.n108 plus.n64 46.3896
R22730 plus.n47 plus.n3 46.3896
R22731 plus.n23 plus.n22 46.3896
R22732 plus.n76 plus.n75 43.1929
R22733 plus.n15 plus.n14 43.1929
R22734 plus.n94 plus.n70 42.5146
R22735 plus.n101 plus.n100 42.5146
R22736 plus.n40 plus.n39 42.5146
R22737 plus.n33 plus.n9 42.5146
R22738 plus.n77 plus.n76 40.6041
R22739 plus.n16 plus.n15 40.6041
R22740 plus.n90 plus.n70 38.6395
R22741 plus.n102 plus.n101 38.6395
R22742 plus.n41 plus.n40 38.6395
R22743 plus.n29 plus.n9 38.6395
R22744 plus.n122 plus.n121 35.2031
R22745 plus.n83 plus.n82 34.7644
R22746 plus.n112 plus.n64 34.7644
R22747 plus.n51 plus.n3 34.7644
R22748 plus.n22 plus.n21 34.7644
R22749 plus.n79 plus.n74 21.8872
R22750 plus.n114 plus.n113 21.8872
R22751 plus.n53 plus.n52 21.8872
R22752 plus.n18 plus.n13 21.8872
R22753 plus.n89 plus.n88 19.9199
R22754 plus.n105 plus.n66 19.9199
R22755 plus.n44 plus.n5 19.9199
R22756 plus.n28 plus.n27 19.9199
R22757 plus.n123 plus.t2 19.8005
R22758 plus.n123 plus.t4 19.8005
R22759 plus.n125 plus.t3 19.8005
R22760 plus.n125 plus.t0 19.8005
R22761 plus.n96 plus.n95 17.9525
R22762 plus.n97 plus.n68 17.9525
R22763 plus.n36 plus.n7 17.9525
R22764 plus.n35 plus.n34 17.9525
R22765 plus.n87 plus.n72 15.9852
R22766 plus.n107 plus.n106 15.9852
R22767 plus.n46 plus.n45 15.9852
R22768 plus.n26 plus.n11 15.9852
R22769 plus plus.n127 15.0684
R22770 plus.n78 plus.n77 14.0178
R22771 plus.n115 plus.n62 14.0178
R22772 plus.n54 plus.n1 14.0178
R22773 plus.n17 plus.n16 14.0178
R22774 plus.n122 plus.n60 11.9342
R22775 plus.n118 plus.n62 10.575
R22776 plus.n57 plus.n1 10.575
R22777 plus.n120 plus.n119 9.49444
R22778 plus.n59 plus.n58 9.49444
R22779 plus.n84 plus.n72 8.60764
R22780 plus.n108 plus.n107 8.60764
R22781 plus.n47 plus.n46 8.60764
R22782 plus.n23 plus.n11 8.60764
R22783 plus.n95 plus.n94 6.6403
R22784 plus.n100 plus.n68 6.6403
R22785 plus.n39 plus.n7 6.6403
R22786 plus.n34 plus.n33 6.6403
R22787 plus.n127 plus.n126 5.40567
R22788 plus.n90 plus.n89 4.67295
R22789 plus.n102 plus.n66 4.67295
R22790 plus.n41 plus.n5 4.67295
R22791 plus.n29 plus.n28 4.67295
R22792 plus.n82 plus.n74 2.7056
R22793 plus.n113 plus.n112 2.7056
R22794 plus.n52 plus.n51 2.7056
R22795 plus.n21 plus.n13 2.7056
R22796 plus.n127 plus.n122 1.188
R22797 plus.n126 plus.n124 0.716017
R22798 plus.n80 plus.n75 0.189894
R22799 plus.n81 plus.n80 0.189894
R22800 plus.n81 plus.n73 0.189894
R22801 plus.n85 plus.n73 0.189894
R22802 plus.n86 plus.n85 0.189894
R22803 plus.n86 plus.n71 0.189894
R22804 plus.n91 plus.n71 0.189894
R22805 plus.n92 plus.n91 0.189894
R22806 plus.n93 plus.n92 0.189894
R22807 plus.n93 plus.n69 0.189894
R22808 plus.n98 plus.n69 0.189894
R22809 plus.n99 plus.n98 0.189894
R22810 plus.n99 plus.n67 0.189894
R22811 plus.n103 plus.n67 0.189894
R22812 plus.n104 plus.n103 0.189894
R22813 plus.n104 plus.n65 0.189894
R22814 plus.n109 plus.n65 0.189894
R22815 plus.n110 plus.n109 0.189894
R22816 plus.n111 plus.n110 0.189894
R22817 plus.n111 plus.n63 0.189894
R22818 plus.n116 plus.n63 0.189894
R22819 plus.n117 plus.n116 0.189894
R22820 plus.n117 plus.n61 0.189894
R22821 plus.n121 plus.n61 0.189894
R22822 plus.n60 plus.n0 0.189894
R22823 plus.n56 plus.n0 0.189894
R22824 plus.n56 plus.n55 0.189894
R22825 plus.n55 plus.n2 0.189894
R22826 plus.n50 plus.n2 0.189894
R22827 plus.n50 plus.n49 0.189894
R22828 plus.n49 plus.n48 0.189894
R22829 plus.n48 plus.n4 0.189894
R22830 plus.n43 plus.n4 0.189894
R22831 plus.n43 plus.n42 0.189894
R22832 plus.n42 plus.n6 0.189894
R22833 plus.n38 plus.n6 0.189894
R22834 plus.n38 plus.n37 0.189894
R22835 plus.n37 plus.n8 0.189894
R22836 plus.n32 plus.n8 0.189894
R22837 plus.n32 plus.n31 0.189894
R22838 plus.n31 plus.n30 0.189894
R22839 plus.n30 plus.n10 0.189894
R22840 plus.n25 plus.n10 0.189894
R22841 plus.n25 plus.n24 0.189894
R22842 plus.n24 plus.n12 0.189894
R22843 plus.n20 plus.n12 0.189894
R22844 plus.n20 plus.n19 0.189894
R22845 plus.n19 plus.n14 0.189894
R22846 a_n3106_n452.n1 a_n3106_n452.t54 214.321
R22847 a_n3106_n452.n14 a_n3106_n452.t30 214.321
R22848 a_n3106_n452.n15 a_n3106_n452.t51 214.321
R22849 a_n3106_n452.n16 a_n3106_n452.t32 214.321
R22850 a_n3106_n452.n17 a_n3106_n452.t50 214.321
R22851 a_n3106_n452.n18 a_n3106_n452.t49 214.321
R22852 a_n3106_n452.n19 a_n3106_n452.t35 214.321
R22853 a_n3106_n452.n20 a_n3106_n452.t53 214.321
R22854 a_n3106_n452.n0 a_n3106_n452.t20 55.8337
R22855 a_n3106_n452.n2 a_n3106_n452.t33 55.8337
R22856 a_n3106_n452.n13 a_n3106_n452.t38 55.8337
R22857 a_n3106_n452.n47 a_n3106_n452.t7 55.8335
R22858 a_n3106_n452.n45 a_n3106_n452.t42 55.8335
R22859 a_n3106_n452.n34 a_n3106_n452.t2 55.8335
R22860 a_n3106_n452.n33 a_n3106_n452.t17 55.8335
R22861 a_n3106_n452.n22 a_n3106_n452.t11 55.8335
R22862 a_n3106_n452.n49 a_n3106_n452.n48 53.0052
R22863 a_n3106_n452.n51 a_n3106_n452.n50 53.0052
R22864 a_n3106_n452.n53 a_n3106_n452.n52 53.0052
R22865 a_n3106_n452.n55 a_n3106_n452.n54 53.0052
R22866 a_n3106_n452.n4 a_n3106_n452.n3 53.0052
R22867 a_n3106_n452.n6 a_n3106_n452.n5 53.0052
R22868 a_n3106_n452.n8 a_n3106_n452.n7 53.0052
R22869 a_n3106_n452.n10 a_n3106_n452.n9 53.0052
R22870 a_n3106_n452.n12 a_n3106_n452.n11 53.0052
R22871 a_n3106_n452.n44 a_n3106_n452.n43 53.0051
R22872 a_n3106_n452.n42 a_n3106_n452.n41 53.0051
R22873 a_n3106_n452.n40 a_n3106_n452.n39 53.0051
R22874 a_n3106_n452.n38 a_n3106_n452.n37 53.0051
R22875 a_n3106_n452.n36 a_n3106_n452.n35 53.0051
R22876 a_n3106_n452.n32 a_n3106_n452.n31 53.0051
R22877 a_n3106_n452.n30 a_n3106_n452.n29 53.0051
R22878 a_n3106_n452.n28 a_n3106_n452.n27 53.0051
R22879 a_n3106_n452.n26 a_n3106_n452.n25 53.0051
R22880 a_n3106_n452.n24 a_n3106_n452.n23 53.0051
R22881 a_n3106_n452.n57 a_n3106_n452.n56 53.0051
R22882 a_n3106_n452.n21 a_n3106_n452.n13 12.2417
R22883 a_n3106_n452.n47 a_n3106_n452.n46 12.2417
R22884 a_n3106_n452.n22 a_n3106_n452.n21 5.16214
R22885 a_n3106_n452.n46 a_n3106_n452.n45 5.16214
R22886 a_n3106_n452.n48 a_n3106_n452.t5 2.82907
R22887 a_n3106_n452.n48 a_n3106_n452.t3 2.82907
R22888 a_n3106_n452.n50 a_n3106_n452.t16 2.82907
R22889 a_n3106_n452.n50 a_n3106_n452.t21 2.82907
R22890 a_n3106_n452.n52 a_n3106_n452.t14 2.82907
R22891 a_n3106_n452.n52 a_n3106_n452.t18 2.82907
R22892 a_n3106_n452.n54 a_n3106_n452.t10 2.82907
R22893 a_n3106_n452.n54 a_n3106_n452.t15 2.82907
R22894 a_n3106_n452.n3 a_n3106_n452.t43 2.82907
R22895 a_n3106_n452.n3 a_n3106_n452.t55 2.82907
R22896 a_n3106_n452.n5 a_n3106_n452.t40 2.82907
R22897 a_n3106_n452.n5 a_n3106_n452.t27 2.82907
R22898 a_n3106_n452.n7 a_n3106_n452.t28 2.82907
R22899 a_n3106_n452.n7 a_n3106_n452.t39 2.82907
R22900 a_n3106_n452.n9 a_n3106_n452.t0 2.82907
R22901 a_n3106_n452.n9 a_n3106_n452.t48 2.82907
R22902 a_n3106_n452.n11 a_n3106_n452.t46 2.82907
R22903 a_n3106_n452.n11 a_n3106_n452.t36 2.82907
R22904 a_n3106_n452.n43 a_n3106_n452.t47 2.82907
R22905 a_n3106_n452.n43 a_n3106_n452.t45 2.82907
R22906 a_n3106_n452.n41 a_n3106_n452.t34 2.82907
R22907 a_n3106_n452.n41 a_n3106_n452.t52 2.82907
R22908 a_n3106_n452.n39 a_n3106_n452.t1 2.82907
R22909 a_n3106_n452.n39 a_n3106_n452.t31 2.82907
R22910 a_n3106_n452.n37 a_n3106_n452.t41 2.82907
R22911 a_n3106_n452.n37 a_n3106_n452.t29 2.82907
R22912 a_n3106_n452.n35 a_n3106_n452.t44 2.82907
R22913 a_n3106_n452.n35 a_n3106_n452.t37 2.82907
R22914 a_n3106_n452.n31 a_n3106_n452.t6 2.82907
R22915 a_n3106_n452.n31 a_n3106_n452.t22 2.82907
R22916 a_n3106_n452.n29 a_n3106_n452.t13 2.82907
R22917 a_n3106_n452.n29 a_n3106_n452.t4 2.82907
R22918 a_n3106_n452.n27 a_n3106_n452.t24 2.82907
R22919 a_n3106_n452.n27 a_n3106_n452.t12 2.82907
R22920 a_n3106_n452.n25 a_n3106_n452.t19 2.82907
R22921 a_n3106_n452.n25 a_n3106_n452.t23 2.82907
R22922 a_n3106_n452.n23 a_n3106_n452.t8 2.82907
R22923 a_n3106_n452.n23 a_n3106_n452.t25 2.82907
R22924 a_n3106_n452.t26 a_n3106_n452.n57 2.82907
R22925 a_n3106_n452.n57 a_n3106_n452.t9 2.82907
R22926 a_n3106_n452.n46 a_n3106_n452.n1 2.54197
R22927 a_n3106_n452.n21 a_n3106_n452.n20 2.0129
R22928 a_n3106_n452.n20 a_n3106_n452.n19 0.672012
R22929 a_n3106_n452.n19 a_n3106_n452.n18 0.672012
R22930 a_n3106_n452.n18 a_n3106_n452.n17 0.672012
R22931 a_n3106_n452.n17 a_n3106_n452.n16 0.672012
R22932 a_n3106_n452.n16 a_n3106_n452.n15 0.672012
R22933 a_n3106_n452.n15 a_n3106_n452.n14 0.672012
R22934 a_n3106_n452.n14 a_n3106_n452.n1 0.672012
R22935 a_n3106_n452.n24 a_n3106_n452.n22 0.530672
R22936 a_n3106_n452.n26 a_n3106_n452.n24 0.530672
R22937 a_n3106_n452.n28 a_n3106_n452.n26 0.530672
R22938 a_n3106_n452.n30 a_n3106_n452.n28 0.530672
R22939 a_n3106_n452.n32 a_n3106_n452.n30 0.530672
R22940 a_n3106_n452.n33 a_n3106_n452.n32 0.530672
R22941 a_n3106_n452.n36 a_n3106_n452.n34 0.530672
R22942 a_n3106_n452.n38 a_n3106_n452.n36 0.530672
R22943 a_n3106_n452.n40 a_n3106_n452.n38 0.530672
R22944 a_n3106_n452.n42 a_n3106_n452.n40 0.530672
R22945 a_n3106_n452.n44 a_n3106_n452.n42 0.530672
R22946 a_n3106_n452.n45 a_n3106_n452.n44 0.530672
R22947 a_n3106_n452.n13 a_n3106_n452.n12 0.530672
R22948 a_n3106_n452.n12 a_n3106_n452.n10 0.530672
R22949 a_n3106_n452.n10 a_n3106_n452.n8 0.530672
R22950 a_n3106_n452.n8 a_n3106_n452.n6 0.530672
R22951 a_n3106_n452.n6 a_n3106_n452.n4 0.530672
R22952 a_n3106_n452.n4 a_n3106_n452.n2 0.530672
R22953 a_n3106_n452.n56 a_n3106_n452.n0 0.530672
R22954 a_n3106_n452.n56 a_n3106_n452.n55 0.530672
R22955 a_n3106_n452.n55 a_n3106_n452.n53 0.530672
R22956 a_n3106_n452.n53 a_n3106_n452.n51 0.530672
R22957 a_n3106_n452.n51 a_n3106_n452.n49 0.530672
R22958 a_n3106_n452.n49 a_n3106_n452.n47 0.530672
R22959 a_n3106_n452.n34 a_n3106_n452.n33 0.235414
R22960 a_n3106_n452.n2 a_n3106_n452.n0 0.235414
R22961 a_n2318_8322.n9 a_n2318_8322.t7 74.6477
R22962 a_n2318_8322.t26 a_n2318_8322.n22 74.6477
R22963 a_n2318_8322.n1 a_n2318_8322.t25 74.6474
R22964 a_n2318_8322.n16 a_n2318_8322.t12 74.2899
R22965 a_n2318_8322.n6 a_n2318_8322.t15 74.2899
R22966 a_n2318_8322.n10 a_n2318_8322.t5 74.2899
R22967 a_n2318_8322.n11 a_n2318_8322.t8 74.2899
R22968 a_n2318_8322.n14 a_n2318_8322.t9 74.2899
R22969 a_n2318_8322.n22 a_n2318_8322.n21 70.6783
R22970 a_n2318_8322.n20 a_n2318_8322.n19 70.6783
R22971 a_n2318_8322.n18 a_n2318_8322.n17 70.6783
R22972 a_n2318_8322.n1 a_n2318_8322.n0 70.6783
R22973 a_n2318_8322.n3 a_n2318_8322.n2 70.6783
R22974 a_n2318_8322.n5 a_n2318_8322.n4 70.6783
R22975 a_n2318_8322.n9 a_n2318_8322.n8 70.6783
R22976 a_n2318_8322.n13 a_n2318_8322.n12 70.6783
R22977 a_n2318_8322.n16 a_n2318_8322.n15 23.4712
R22978 a_n2318_8322.n7 a_n2318_8322.t3 10.0266
R22979 a_n2318_8322.n15 a_n2318_8322.n14 6.95632
R22980 a_n2318_8322.n7 a_n2318_8322.n6 6.19447
R22981 a_n2318_8322.n15 a_n2318_8322.n7 5.3452
R22982 a_n2318_8322.n21 a_n2318_8322.t14 3.61217
R22983 a_n2318_8322.n21 a_n2318_8322.t13 3.61217
R22984 a_n2318_8322.n19 a_n2318_8322.t23 3.61217
R22985 a_n2318_8322.n19 a_n2318_8322.t18 3.61217
R22986 a_n2318_8322.n17 a_n2318_8322.t21 3.61217
R22987 a_n2318_8322.n17 a_n2318_8322.t20 3.61217
R22988 a_n2318_8322.n0 a_n2318_8322.t22 3.61217
R22989 a_n2318_8322.n0 a_n2318_8322.t19 3.61217
R22990 a_n2318_8322.n2 a_n2318_8322.t16 3.61217
R22991 a_n2318_8322.n2 a_n2318_8322.t27 3.61217
R22992 a_n2318_8322.n4 a_n2318_8322.t24 3.61217
R22993 a_n2318_8322.n4 a_n2318_8322.t17 3.61217
R22994 a_n2318_8322.n8 a_n2318_8322.t11 3.61217
R22995 a_n2318_8322.n8 a_n2318_8322.t10 3.61217
R22996 a_n2318_8322.n12 a_n2318_8322.t6 3.61217
R22997 a_n2318_8322.n12 a_n2318_8322.t4 3.61217
R22998 a_n2318_8322.n6 a_n2318_8322.n5 0.358259
R22999 a_n2318_8322.n5 a_n2318_8322.n3 0.358259
R23000 a_n2318_8322.n3 a_n2318_8322.n1 0.358259
R23001 a_n2318_8322.n14 a_n2318_8322.n13 0.358259
R23002 a_n2318_8322.n13 a_n2318_8322.n11 0.358259
R23003 a_n2318_8322.n10 a_n2318_8322.n9 0.358259
R23004 a_n2318_8322.n18 a_n2318_8322.n16 0.358259
R23005 a_n2318_8322.n20 a_n2318_8322.n18 0.358259
R23006 a_n2318_8322.n22 a_n2318_8322.n20 0.358259
R23007 a_n2318_8322.n11 a_n2318_8322.n10 0.101793
R23008 a_n2318_8322.t2 a_n2318_8322.t1 0.0788333
R23009 a_n2318_8322.t0 a_n2318_8322.t2 0.0631667
R23010 a_n2318_8322.t3 a_n2318_8322.t0 0.0471944
R23011 a_n2318_8322.t3 a_n2318_8322.t1 0.0453889
R23012 output.n41 output.n15 289.615
R23013 output.n72 output.n46 289.615
R23014 output.n104 output.n78 289.615
R23015 output.n136 output.n110 289.615
R23016 output.n77 output.n45 197.26
R23017 output.n77 output.n76 196.298
R23018 output.n109 output.n108 196.298
R23019 output.n141 output.n140 196.298
R23020 output.n42 output.n41 185
R23021 output.n40 output.n39 185
R23022 output.n19 output.n18 185
R23023 output.n34 output.n33 185
R23024 output.n32 output.n31 185
R23025 output.n23 output.n22 185
R23026 output.n26 output.n25 185
R23027 output.n73 output.n72 185
R23028 output.n71 output.n70 185
R23029 output.n50 output.n49 185
R23030 output.n65 output.n64 185
R23031 output.n63 output.n62 185
R23032 output.n54 output.n53 185
R23033 output.n57 output.n56 185
R23034 output.n105 output.n104 185
R23035 output.n103 output.n102 185
R23036 output.n82 output.n81 185
R23037 output.n97 output.n96 185
R23038 output.n95 output.n94 185
R23039 output.n86 output.n85 185
R23040 output.n89 output.n88 185
R23041 output.n137 output.n136 185
R23042 output.n135 output.n134 185
R23043 output.n114 output.n113 185
R23044 output.n129 output.n128 185
R23045 output.n127 output.n126 185
R23046 output.n118 output.n117 185
R23047 output.n121 output.n120 185
R23048 output.t18 output.n24 147.661
R23049 output.t19 output.n55 147.661
R23050 output.t17 output.n87 147.661
R23051 output.t16 output.n119 147.661
R23052 output.n41 output.n40 104.615
R23053 output.n40 output.n18 104.615
R23054 output.n33 output.n18 104.615
R23055 output.n33 output.n32 104.615
R23056 output.n32 output.n22 104.615
R23057 output.n25 output.n22 104.615
R23058 output.n72 output.n71 104.615
R23059 output.n71 output.n49 104.615
R23060 output.n64 output.n49 104.615
R23061 output.n64 output.n63 104.615
R23062 output.n63 output.n53 104.615
R23063 output.n56 output.n53 104.615
R23064 output.n104 output.n103 104.615
R23065 output.n103 output.n81 104.615
R23066 output.n96 output.n81 104.615
R23067 output.n96 output.n95 104.615
R23068 output.n95 output.n85 104.615
R23069 output.n88 output.n85 104.615
R23070 output.n136 output.n135 104.615
R23071 output.n135 output.n113 104.615
R23072 output.n128 output.n113 104.615
R23073 output.n128 output.n127 104.615
R23074 output.n127 output.n117 104.615
R23075 output.n120 output.n117 104.615
R23076 output.n1 output.t10 77.056
R23077 output.n14 output.t11 76.6694
R23078 output.n1 output.n0 72.7095
R23079 output.n3 output.n2 72.7095
R23080 output.n5 output.n4 72.7095
R23081 output.n7 output.n6 72.7095
R23082 output.n9 output.n8 72.7095
R23083 output.n11 output.n10 72.7095
R23084 output.n13 output.n12 72.7095
R23085 output.n25 output.t18 52.3082
R23086 output.n56 output.t19 52.3082
R23087 output.n88 output.t17 52.3082
R23088 output.n120 output.t16 52.3082
R23089 output.n26 output.n24 15.6674
R23090 output.n57 output.n55 15.6674
R23091 output.n89 output.n87 15.6674
R23092 output.n121 output.n119 15.6674
R23093 output.n27 output.n23 12.8005
R23094 output.n58 output.n54 12.8005
R23095 output.n90 output.n86 12.8005
R23096 output.n122 output.n118 12.8005
R23097 output.n31 output.n30 12.0247
R23098 output.n62 output.n61 12.0247
R23099 output.n94 output.n93 12.0247
R23100 output.n126 output.n125 12.0247
R23101 output.n34 output.n21 11.249
R23102 output.n65 output.n52 11.249
R23103 output.n97 output.n84 11.249
R23104 output.n129 output.n116 11.249
R23105 output.n35 output.n19 10.4732
R23106 output.n66 output.n50 10.4732
R23107 output.n98 output.n82 10.4732
R23108 output.n130 output.n114 10.4732
R23109 output.n39 output.n38 9.69747
R23110 output.n70 output.n69 9.69747
R23111 output.n102 output.n101 9.69747
R23112 output.n134 output.n133 9.69747
R23113 output.n45 output.n44 9.45567
R23114 output.n76 output.n75 9.45567
R23115 output.n108 output.n107 9.45567
R23116 output.n140 output.n139 9.45567
R23117 output.n44 output.n43 9.3005
R23118 output.n17 output.n16 9.3005
R23119 output.n38 output.n37 9.3005
R23120 output.n36 output.n35 9.3005
R23121 output.n21 output.n20 9.3005
R23122 output.n30 output.n29 9.3005
R23123 output.n28 output.n27 9.3005
R23124 output.n75 output.n74 9.3005
R23125 output.n48 output.n47 9.3005
R23126 output.n69 output.n68 9.3005
R23127 output.n67 output.n66 9.3005
R23128 output.n52 output.n51 9.3005
R23129 output.n61 output.n60 9.3005
R23130 output.n59 output.n58 9.3005
R23131 output.n107 output.n106 9.3005
R23132 output.n80 output.n79 9.3005
R23133 output.n101 output.n100 9.3005
R23134 output.n99 output.n98 9.3005
R23135 output.n84 output.n83 9.3005
R23136 output.n93 output.n92 9.3005
R23137 output.n91 output.n90 9.3005
R23138 output.n139 output.n138 9.3005
R23139 output.n112 output.n111 9.3005
R23140 output.n133 output.n132 9.3005
R23141 output.n131 output.n130 9.3005
R23142 output.n116 output.n115 9.3005
R23143 output.n125 output.n124 9.3005
R23144 output.n123 output.n122 9.3005
R23145 output.n42 output.n17 8.92171
R23146 output.n73 output.n48 8.92171
R23147 output.n105 output.n80 8.92171
R23148 output.n137 output.n112 8.92171
R23149 output output.n141 8.15037
R23150 output.n43 output.n15 8.14595
R23151 output.n74 output.n46 8.14595
R23152 output.n106 output.n78 8.14595
R23153 output.n138 output.n110 8.14595
R23154 output.n45 output.n15 5.81868
R23155 output.n76 output.n46 5.81868
R23156 output.n108 output.n78 5.81868
R23157 output.n140 output.n110 5.81868
R23158 output.n43 output.n42 5.04292
R23159 output.n74 output.n73 5.04292
R23160 output.n106 output.n105 5.04292
R23161 output.n138 output.n137 5.04292
R23162 output.n28 output.n24 4.38594
R23163 output.n59 output.n55 4.38594
R23164 output.n91 output.n87 4.38594
R23165 output.n123 output.n119 4.38594
R23166 output.n39 output.n17 4.26717
R23167 output.n70 output.n48 4.26717
R23168 output.n102 output.n80 4.26717
R23169 output.n134 output.n112 4.26717
R23170 output.n0 output.t4 3.9605
R23171 output.n0 output.t2 3.9605
R23172 output.n2 output.t9 3.9605
R23173 output.n2 output.t12 3.9605
R23174 output.n4 output.t14 3.9605
R23175 output.n4 output.t6 3.9605
R23176 output.n6 output.t8 3.9605
R23177 output.n6 output.t15 3.9605
R23178 output.n8 output.t0 3.9605
R23179 output.n8 output.t5 3.9605
R23180 output.n10 output.t7 3.9605
R23181 output.n10 output.t13 3.9605
R23182 output.n12 output.t3 3.9605
R23183 output.n12 output.t1 3.9605
R23184 output.n38 output.n19 3.49141
R23185 output.n69 output.n50 3.49141
R23186 output.n101 output.n82 3.49141
R23187 output.n133 output.n114 3.49141
R23188 output.n35 output.n34 2.71565
R23189 output.n66 output.n65 2.71565
R23190 output.n98 output.n97 2.71565
R23191 output.n130 output.n129 2.71565
R23192 output.n31 output.n21 1.93989
R23193 output.n62 output.n52 1.93989
R23194 output.n94 output.n84 1.93989
R23195 output.n126 output.n116 1.93989
R23196 output.n30 output.n23 1.16414
R23197 output.n61 output.n54 1.16414
R23198 output.n93 output.n86 1.16414
R23199 output.n125 output.n118 1.16414
R23200 output.n141 output.n109 0.962709
R23201 output.n109 output.n77 0.962709
R23202 output.n27 output.n26 0.388379
R23203 output.n58 output.n57 0.388379
R23204 output.n90 output.n89 0.388379
R23205 output.n122 output.n121 0.388379
R23206 output.n14 output.n13 0.387128
R23207 output.n13 output.n11 0.387128
R23208 output.n11 output.n9 0.387128
R23209 output.n9 output.n7 0.387128
R23210 output.n7 output.n5 0.387128
R23211 output.n5 output.n3 0.387128
R23212 output.n3 output.n1 0.387128
R23213 output.n44 output.n16 0.155672
R23214 output.n37 output.n16 0.155672
R23215 output.n37 output.n36 0.155672
R23216 output.n36 output.n20 0.155672
R23217 output.n29 output.n20 0.155672
R23218 output.n29 output.n28 0.155672
R23219 output.n75 output.n47 0.155672
R23220 output.n68 output.n47 0.155672
R23221 output.n68 output.n67 0.155672
R23222 output.n67 output.n51 0.155672
R23223 output.n60 output.n51 0.155672
R23224 output.n60 output.n59 0.155672
R23225 output.n107 output.n79 0.155672
R23226 output.n100 output.n79 0.155672
R23227 output.n100 output.n99 0.155672
R23228 output.n99 output.n83 0.155672
R23229 output.n92 output.n83 0.155672
R23230 output.n92 output.n91 0.155672
R23231 output.n139 output.n111 0.155672
R23232 output.n132 output.n111 0.155672
R23233 output.n132 output.n131 0.155672
R23234 output.n131 output.n115 0.155672
R23235 output.n124 output.n115 0.155672
R23236 output.n124 output.n123 0.155672
R23237 output output.n14 0.126227
R23238 minus.n76 minus.t28 250.337
R23239 minus.n15 minus.t20 250.337
R23240 minus.n126 minus.t1 243.255
R23241 minus.n120 minus.t8 231.093
R23242 minus.n59 minus.t10 231.093
R23243 minus.n125 minus.n123 224.169
R23244 minus.n125 minus.n124 223.454
R23245 minus.n62 minus.t12 187.445
R23246 minus.n113 minus.t18 187.445
R23247 minus.n107 minus.t25 187.445
R23248 minus.n66 minus.t22 187.445
R23249 minus.n68 minus.t19 187.445
R23250 minus.n95 minus.t7 187.445
R23251 minus.n89 minus.t6 187.445
R23252 minus.n72 minus.t16 187.445
R23253 minus.n74 minus.t15 187.445
R23254 minus.n77 minus.t23 187.445
R23255 minus.n16 minus.t14 187.445
R23256 minus.n13 minus.t9 187.445
R23257 minus.n11 minus.t5 187.445
R23258 minus.n28 minus.t26 187.445
R23259 minus.n34 minus.t27 187.445
R23260 minus.n7 minus.t21 187.445
R23261 minus.n5 minus.t24 187.445
R23262 minus.n46 minus.t17 187.445
R23263 minus.n52 minus.t11 187.445
R23264 minus.n1 minus.t13 187.445
R23265 minus.n78 minus.n75 161.3
R23266 minus.n80 minus.n79 161.3
R23267 minus.n82 minus.n81 161.3
R23268 minus.n83 minus.n73 161.3
R23269 minus.n85 minus.n84 161.3
R23270 minus.n87 minus.n86 161.3
R23271 minus.n88 minus.n71 161.3
R23272 minus.n91 minus.n90 161.3
R23273 minus.n92 minus.n70 161.3
R23274 minus.n94 minus.n93 161.3
R23275 minus.n96 minus.n69 161.3
R23276 minus.n98 minus.n97 161.3
R23277 minus.n100 minus.n99 161.3
R23278 minus.n101 minus.n67 161.3
R23279 minus.n103 minus.n102 161.3
R23280 minus.n105 minus.n104 161.3
R23281 minus.n106 minus.n65 161.3
R23282 minus.n109 minus.n108 161.3
R23283 minus.n110 minus.n64 161.3
R23284 minus.n112 minus.n111 161.3
R23285 minus.n114 minus.n63 161.3
R23286 minus.n116 minus.n115 161.3
R23287 minus.n118 minus.n117 161.3
R23288 minus.n119 minus.n61 161.3
R23289 minus.n121 minus.n120 161.3
R23290 minus.n60 minus.n59 161.3
R23291 minus.n58 minus.n0 161.3
R23292 minus.n57 minus.n56 161.3
R23293 minus.n55 minus.n54 161.3
R23294 minus.n53 minus.n2 161.3
R23295 minus.n51 minus.n50 161.3
R23296 minus.n49 minus.n3 161.3
R23297 minus.n48 minus.n47 161.3
R23298 minus.n45 minus.n4 161.3
R23299 minus.n44 minus.n43 161.3
R23300 minus.n42 minus.n41 161.3
R23301 minus.n40 minus.n6 161.3
R23302 minus.n39 minus.n38 161.3
R23303 minus.n37 minus.n36 161.3
R23304 minus.n35 minus.n8 161.3
R23305 minus.n33 minus.n32 161.3
R23306 minus.n31 minus.n9 161.3
R23307 minus.n30 minus.n29 161.3
R23308 minus.n27 minus.n10 161.3
R23309 minus.n26 minus.n25 161.3
R23310 minus.n24 minus.n23 161.3
R23311 minus.n22 minus.n12 161.3
R23312 minus.n21 minus.n20 161.3
R23313 minus.n19 minus.n18 161.3
R23314 minus.n17 minus.n14 161.3
R23315 minus.n106 minus.n105 56.5617
R23316 minus.n97 minus.n96 56.5617
R23317 minus.n88 minus.n87 56.5617
R23318 minus.n27 minus.n26 56.5617
R23319 minus.n36 minus.n35 56.5617
R23320 minus.n45 minus.n44 56.5617
R23321 minus.n115 minus.n114 56.5617
R23322 minus.n79 minus.n78 56.5617
R23323 minus.n18 minus.n17 56.5617
R23324 minus.n54 minus.n53 56.5617
R23325 minus.n119 minus.n118 50.2647
R23326 minus.n58 minus.n57 50.2647
R23327 minus.n108 minus.n64 46.3896
R23328 minus.n84 minus.n83 46.3896
R23329 minus.n23 minus.n22 46.3896
R23330 minus.n47 minus.n3 46.3896
R23331 minus.n76 minus.n75 43.1929
R23332 minus.n15 minus.n14 43.1929
R23333 minus.n101 minus.n100 42.5146
R23334 minus.n94 minus.n70 42.5146
R23335 minus.n33 minus.n9 42.5146
R23336 minus.n40 minus.n39 42.5146
R23337 minus.n77 minus.n76 40.6041
R23338 minus.n16 minus.n15 40.6041
R23339 minus.n102 minus.n101 38.6395
R23340 minus.n90 minus.n70 38.6395
R23341 minus.n29 minus.n9 38.6395
R23342 minus.n41 minus.n40 38.6395
R23343 minus.n122 minus.n121 35.4191
R23344 minus.n112 minus.n64 34.7644
R23345 minus.n83 minus.n82 34.7644
R23346 minus.n22 minus.n21 34.7644
R23347 minus.n51 minus.n3 34.7644
R23348 minus.n114 minus.n113 21.8872
R23349 minus.n79 minus.n74 21.8872
R23350 minus.n18 minus.n13 21.8872
R23351 minus.n53 minus.n52 21.8872
R23352 minus.n105 minus.n66 19.9199
R23353 minus.n89 minus.n88 19.9199
R23354 minus.n28 minus.n27 19.9199
R23355 minus.n44 minus.n5 19.9199
R23356 minus.n124 minus.t0 19.8005
R23357 minus.n124 minus.t2 19.8005
R23358 minus.n123 minus.t4 19.8005
R23359 minus.n123 minus.t3 19.8005
R23360 minus.n97 minus.n68 17.9525
R23361 minus.n96 minus.n95 17.9525
R23362 minus.n35 minus.n34 17.9525
R23363 minus.n36 minus.n7 17.9525
R23364 minus.n107 minus.n106 15.9852
R23365 minus.n87 minus.n72 15.9852
R23366 minus.n26 minus.n11 15.9852
R23367 minus.n46 minus.n45 15.9852
R23368 minus.n115 minus.n62 14.0178
R23369 minus.n78 minus.n77 14.0178
R23370 minus.n17 minus.n16 14.0178
R23371 minus.n54 minus.n1 14.0178
R23372 minus.n122 minus.n60 12.1501
R23373 minus minus.n127 11.5812
R23374 minus.n118 minus.n62 10.575
R23375 minus.n57 minus.n1 10.575
R23376 minus.n120 minus.n119 9.49444
R23377 minus.n59 minus.n58 9.49444
R23378 minus.n108 minus.n107 8.60764
R23379 minus.n84 minus.n72 8.60764
R23380 minus.n23 minus.n11 8.60764
R23381 minus.n47 minus.n46 8.60764
R23382 minus.n100 minus.n68 6.6403
R23383 minus.n95 minus.n94 6.6403
R23384 minus.n34 minus.n33 6.6403
R23385 minus.n39 minus.n7 6.6403
R23386 minus.n127 minus.n126 4.80222
R23387 minus.n102 minus.n66 4.67295
R23388 minus.n90 minus.n89 4.67295
R23389 minus.n29 minus.n28 4.67295
R23390 minus.n41 minus.n5 4.67295
R23391 minus.n113 minus.n112 2.7056
R23392 minus.n82 minus.n74 2.7056
R23393 minus.n21 minus.n13 2.7056
R23394 minus.n52 minus.n51 2.7056
R23395 minus.n127 minus.n122 0.972091
R23396 minus.n126 minus.n125 0.716017
R23397 minus.n121 minus.n61 0.189894
R23398 minus.n117 minus.n61 0.189894
R23399 minus.n117 minus.n116 0.189894
R23400 minus.n116 minus.n63 0.189894
R23401 minus.n111 minus.n63 0.189894
R23402 minus.n111 minus.n110 0.189894
R23403 minus.n110 minus.n109 0.189894
R23404 minus.n109 minus.n65 0.189894
R23405 minus.n104 minus.n65 0.189894
R23406 minus.n104 minus.n103 0.189894
R23407 minus.n103 minus.n67 0.189894
R23408 minus.n99 minus.n67 0.189894
R23409 minus.n99 minus.n98 0.189894
R23410 minus.n98 minus.n69 0.189894
R23411 minus.n93 minus.n69 0.189894
R23412 minus.n93 minus.n92 0.189894
R23413 minus.n92 minus.n91 0.189894
R23414 minus.n91 minus.n71 0.189894
R23415 minus.n86 minus.n71 0.189894
R23416 minus.n86 minus.n85 0.189894
R23417 minus.n85 minus.n73 0.189894
R23418 minus.n81 minus.n73 0.189894
R23419 minus.n81 minus.n80 0.189894
R23420 minus.n80 minus.n75 0.189894
R23421 minus.n19 minus.n14 0.189894
R23422 minus.n20 minus.n19 0.189894
R23423 minus.n20 minus.n12 0.189894
R23424 minus.n24 minus.n12 0.189894
R23425 minus.n25 minus.n24 0.189894
R23426 minus.n25 minus.n10 0.189894
R23427 minus.n30 minus.n10 0.189894
R23428 minus.n31 minus.n30 0.189894
R23429 minus.n32 minus.n31 0.189894
R23430 minus.n32 minus.n8 0.189894
R23431 minus.n37 minus.n8 0.189894
R23432 minus.n38 minus.n37 0.189894
R23433 minus.n38 minus.n6 0.189894
R23434 minus.n42 minus.n6 0.189894
R23435 minus.n43 minus.n42 0.189894
R23436 minus.n43 minus.n4 0.189894
R23437 minus.n48 minus.n4 0.189894
R23438 minus.n49 minus.n48 0.189894
R23439 minus.n50 minus.n49 0.189894
R23440 minus.n50 minus.n2 0.189894
R23441 minus.n55 minus.n2 0.189894
R23442 minus.n56 minus.n55 0.189894
R23443 minus.n56 minus.n0 0.189894
R23444 minus.n60 minus.n0 0.189894
R23445 diffpairibias.n0 diffpairibias.t18 436.822
R23446 diffpairibias.n21 diffpairibias.t19 435.479
R23447 diffpairibias.n20 diffpairibias.t16 435.479
R23448 diffpairibias.n19 diffpairibias.t17 435.479
R23449 diffpairibias.n18 diffpairibias.t21 435.479
R23450 diffpairibias.n0 diffpairibias.t22 435.479
R23451 diffpairibias.n1 diffpairibias.t20 435.479
R23452 diffpairibias.n2 diffpairibias.t23 435.479
R23453 diffpairibias.n10 diffpairibias.t0 377.536
R23454 diffpairibias.n10 diffpairibias.t8 376.193
R23455 diffpairibias.n11 diffpairibias.t10 376.193
R23456 diffpairibias.n12 diffpairibias.t6 376.193
R23457 diffpairibias.n13 diffpairibias.t2 376.193
R23458 diffpairibias.n14 diffpairibias.t12 376.193
R23459 diffpairibias.n15 diffpairibias.t4 376.193
R23460 diffpairibias.n16 diffpairibias.t14 376.193
R23461 diffpairibias.n3 diffpairibias.t1 113.368
R23462 diffpairibias.n3 diffpairibias.t9 112.698
R23463 diffpairibias.n4 diffpairibias.t11 112.698
R23464 diffpairibias.n5 diffpairibias.t7 112.698
R23465 diffpairibias.n6 diffpairibias.t3 112.698
R23466 diffpairibias.n7 diffpairibias.t13 112.698
R23467 diffpairibias.n8 diffpairibias.t5 112.698
R23468 diffpairibias.n9 diffpairibias.t15 112.698
R23469 diffpairibias.n17 diffpairibias.n16 4.77242
R23470 diffpairibias.n17 diffpairibias.n9 4.30807
R23471 diffpairibias.n18 diffpairibias.n17 4.13945
R23472 diffpairibias.n16 diffpairibias.n15 1.34352
R23473 diffpairibias.n15 diffpairibias.n14 1.34352
R23474 diffpairibias.n14 diffpairibias.n13 1.34352
R23475 diffpairibias.n13 diffpairibias.n12 1.34352
R23476 diffpairibias.n12 diffpairibias.n11 1.34352
R23477 diffpairibias.n11 diffpairibias.n10 1.34352
R23478 diffpairibias.n2 diffpairibias.n1 1.34352
R23479 diffpairibias.n1 diffpairibias.n0 1.34352
R23480 diffpairibias.n19 diffpairibias.n18 1.34352
R23481 diffpairibias.n20 diffpairibias.n19 1.34352
R23482 diffpairibias.n21 diffpairibias.n20 1.34352
R23483 diffpairibias.n22 diffpairibias.n21 0.862419
R23484 diffpairibias diffpairibias.n22 0.684875
R23485 diffpairibias.n9 diffpairibias.n8 0.672012
R23486 diffpairibias.n8 diffpairibias.n7 0.672012
R23487 diffpairibias.n7 diffpairibias.n6 0.672012
R23488 diffpairibias.n6 diffpairibias.n5 0.672012
R23489 diffpairibias.n5 diffpairibias.n4 0.672012
R23490 diffpairibias.n4 diffpairibias.n3 0.672012
R23491 diffpairibias.n22 diffpairibias.n2 0.190907
C0 commonsourceibias output 0.006808f
C1 minus diffpairibias 5.39e-19
C2 CSoutput minus 2.80108f
C3 vdd plus 0.083679f
C4 plus diffpairibias 4.4e-19
C5 commonsourceibias outputibias 0.003832f
C6 vdd commonsourceibias 0.004218f
C7 CSoutput plus 0.9147f
C8 commonsourceibias diffpairibias 0.052851f
C9 CSoutput commonsourceibias 44.9728f
C10 minus plus 10.4342f
C11 minus commonsourceibias 0.515369f
C12 plus commonsourceibias 0.498793f
C13 output outputibias 2.34152f
C14 vdd output 7.23429f
C15 CSoutput output 6.13571f
C16 CSoutput outputibias 0.032386f
C17 vdd CSoutput 92.2856f
C18 diffpairibias gnd 48.95304f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.180656p
C22 plus gnd 39.338802f
C23 minus gnd 31.268171f
C24 CSoutput gnd 0.114548p
C25 vdd gnd 0.412024p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 minus.n0 gnd 0.030662f
C74 minus.t13 gnd 0.515581f
C75 minus.n1 gnd 0.208524f
C76 minus.n2 gnd 0.030662f
C77 minus.t11 gnd 0.515581f
C78 minus.n3 gnd 0.026202f
C79 minus.n4 gnd 0.030662f
C80 minus.t17 gnd 0.515581f
C81 minus.t24 gnd 0.515581f
C82 minus.n5 gnd 0.208524f
C83 minus.n6 gnd 0.030662f
C84 minus.t21 gnd 0.515581f
C85 minus.n7 gnd 0.208524f
C86 minus.n8 gnd 0.030662f
C87 minus.t27 gnd 0.515581f
C88 minus.n9 gnd 0.024922f
C89 minus.n10 gnd 0.030662f
C90 minus.t26 gnd 0.515581f
C91 minus.t5 gnd 0.515581f
C92 minus.n11 gnd 0.208524f
C93 minus.n12 gnd 0.030662f
C94 minus.t9 gnd 0.515581f
C95 minus.n13 gnd 0.208524f
C96 minus.n14 gnd 0.130127f
C97 minus.t14 gnd 0.515581f
C98 minus.t20 gnd 0.576771f
C99 minus.n15 gnd 0.243785f
C100 minus.n16 gnd 0.238799f
C101 minus.n17 gnd 0.039289f
C102 minus.n18 gnd 0.034698f
C103 minus.n19 gnd 0.030662f
C104 minus.n20 gnd 0.030662f
C105 minus.n21 gnd 0.036642f
C106 minus.n22 gnd 0.026202f
C107 minus.n23 gnd 0.039934f
C108 minus.n24 gnd 0.030662f
C109 minus.n25 gnd 0.030662f
C110 minus.n26 gnd 0.038141f
C111 minus.n27 gnd 0.035846f
C112 minus.n28 gnd 0.208524f
C113 minus.n29 gnd 0.038409f
C114 minus.n30 gnd 0.030662f
C115 minus.n31 gnd 0.030662f
C116 minus.n32 gnd 0.030662f
C117 minus.n33 gnd 0.039446f
C118 minus.n34 gnd 0.208524f
C119 minus.n35 gnd 0.036993f
C120 minus.n36 gnd 0.036993f
C121 minus.n37 gnd 0.030662f
C122 minus.n38 gnd 0.030662f
C123 minus.n39 gnd 0.039446f
C124 minus.n40 gnd 0.024922f
C125 minus.n41 gnd 0.038409f
C126 minus.n42 gnd 0.030662f
C127 minus.n43 gnd 0.030662f
C128 minus.n44 gnd 0.035846f
C129 minus.n45 gnd 0.038141f
C130 minus.n46 gnd 0.208524f
C131 minus.n47 gnd 0.039934f
C132 minus.n48 gnd 0.030662f
C133 minus.n49 gnd 0.030662f
C134 minus.n50 gnd 0.030662f
C135 minus.n51 gnd 0.036642f
C136 minus.n52 gnd 0.208524f
C137 minus.n53 gnd 0.034698f
C138 minus.n54 gnd 0.039289f
C139 minus.n55 gnd 0.030662f
C140 minus.n56 gnd 0.030662f
C141 minus.n57 gnd 0.04f
C142 minus.n58 gnd 0.011144f
C143 minus.t10 gnd 0.557601f
C144 minus.n59 gnd 0.241436f
C145 minus.n60 gnd 0.359197f
C146 minus.n61 gnd 0.030662f
C147 minus.t8 gnd 0.557601f
C148 minus.t12 gnd 0.515581f
C149 minus.n62 gnd 0.208524f
C150 minus.n63 gnd 0.030662f
C151 minus.t18 gnd 0.515581f
C152 minus.n64 gnd 0.026202f
C153 minus.n65 gnd 0.030662f
C154 minus.t25 gnd 0.515581f
C155 minus.t22 gnd 0.515581f
C156 minus.n66 gnd 0.208524f
C157 minus.n67 gnd 0.030662f
C158 minus.t19 gnd 0.515581f
C159 minus.n68 gnd 0.208524f
C160 minus.n69 gnd 0.030662f
C161 minus.t7 gnd 0.515581f
C162 minus.n70 gnd 0.024922f
C163 minus.n71 gnd 0.030662f
C164 minus.t6 gnd 0.515581f
C165 minus.t16 gnd 0.515581f
C166 minus.n72 gnd 0.208524f
C167 minus.n73 gnd 0.030662f
C168 minus.t15 gnd 0.515581f
C169 minus.n74 gnd 0.208524f
C170 minus.n75 gnd 0.130127f
C171 minus.t23 gnd 0.515581f
C172 minus.t28 gnd 0.576771f
C173 minus.n76 gnd 0.243785f
C174 minus.n77 gnd 0.238799f
C175 minus.n78 gnd 0.039289f
C176 minus.n79 gnd 0.034698f
C177 minus.n80 gnd 0.030662f
C178 minus.n81 gnd 0.030662f
C179 minus.n82 gnd 0.036642f
C180 minus.n83 gnd 0.026202f
C181 minus.n84 gnd 0.039934f
C182 minus.n85 gnd 0.030662f
C183 minus.n86 gnd 0.030662f
C184 minus.n87 gnd 0.038141f
C185 minus.n88 gnd 0.035846f
C186 minus.n89 gnd 0.208524f
C187 minus.n90 gnd 0.038409f
C188 minus.n91 gnd 0.030662f
C189 minus.n92 gnd 0.030662f
C190 minus.n93 gnd 0.030662f
C191 minus.n94 gnd 0.039446f
C192 minus.n95 gnd 0.208524f
C193 minus.n96 gnd 0.036993f
C194 minus.n97 gnd 0.036993f
C195 minus.n98 gnd 0.030662f
C196 minus.n99 gnd 0.030662f
C197 minus.n100 gnd 0.039446f
C198 minus.n101 gnd 0.024922f
C199 minus.n102 gnd 0.038409f
C200 minus.n103 gnd 0.030662f
C201 minus.n104 gnd 0.030662f
C202 minus.n105 gnd 0.035846f
C203 minus.n106 gnd 0.038141f
C204 minus.n107 gnd 0.208524f
C205 minus.n108 gnd 0.039934f
C206 minus.n109 gnd 0.030662f
C207 minus.n110 gnd 0.030662f
C208 minus.n111 gnd 0.030662f
C209 minus.n112 gnd 0.036642f
C210 minus.n113 gnd 0.208524f
C211 minus.n114 gnd 0.034698f
C212 minus.n115 gnd 0.039289f
C213 minus.n116 gnd 0.030662f
C214 minus.n117 gnd 0.030662f
C215 minus.n118 gnd 0.04f
C216 minus.n119 gnd 0.011144f
C217 minus.n120 gnd 0.241436f
C218 minus.n121 gnd 1.11855f
C219 minus.n122 gnd 1.64306f
C220 minus.t4 gnd 0.009452f
C221 minus.t3 gnd 0.009452f
C222 minus.n123 gnd 0.031081f
C223 minus.t0 gnd 0.009452f
C224 minus.t2 gnd 0.009452f
C225 minus.n124 gnd 0.030655f
C226 minus.n125 gnd 0.26163f
C227 minus.t1 gnd 0.05261f
C228 minus.n126 gnd 0.142769f
C229 minus.n127 gnd 1.95331f
C230 output.t10 gnd 0.464308f
C231 output.t4 gnd 0.044422f
C232 output.t2 gnd 0.044422f
C233 output.n0 gnd 0.364624f
C234 output.n1 gnd 0.614102f
C235 output.t9 gnd 0.044422f
C236 output.t12 gnd 0.044422f
C237 output.n2 gnd 0.364624f
C238 output.n3 gnd 0.350265f
C239 output.t14 gnd 0.044422f
C240 output.t6 gnd 0.044422f
C241 output.n4 gnd 0.364624f
C242 output.n5 gnd 0.350265f
C243 output.t8 gnd 0.044422f
C244 output.t15 gnd 0.044422f
C245 output.n6 gnd 0.364624f
C246 output.n7 gnd 0.350265f
C247 output.t0 gnd 0.044422f
C248 output.t5 gnd 0.044422f
C249 output.n8 gnd 0.364624f
C250 output.n9 gnd 0.350265f
C251 output.t7 gnd 0.044422f
C252 output.t13 gnd 0.044422f
C253 output.n10 gnd 0.364624f
C254 output.n11 gnd 0.350265f
C255 output.t3 gnd 0.044422f
C256 output.t1 gnd 0.044422f
C257 output.n12 gnd 0.364624f
C258 output.n13 gnd 0.350265f
C259 output.t11 gnd 0.462979f
C260 output.n14 gnd 0.28994f
C261 output.n15 gnd 0.015803f
C262 output.n16 gnd 0.011243f
C263 output.n17 gnd 0.006041f
C264 output.n18 gnd 0.01428f
C265 output.n19 gnd 0.006397f
C266 output.n20 gnd 0.011243f
C267 output.n21 gnd 0.006041f
C268 output.n22 gnd 0.01428f
C269 output.n23 gnd 0.006397f
C270 output.n24 gnd 0.048111f
C271 output.t18 gnd 0.023274f
C272 output.n25 gnd 0.01071f
C273 output.n26 gnd 0.008435f
C274 output.n27 gnd 0.006041f
C275 output.n28 gnd 0.267512f
C276 output.n29 gnd 0.011243f
C277 output.n30 gnd 0.006041f
C278 output.n31 gnd 0.006397f
C279 output.n32 gnd 0.01428f
C280 output.n33 gnd 0.01428f
C281 output.n34 gnd 0.006397f
C282 output.n35 gnd 0.006041f
C283 output.n36 gnd 0.011243f
C284 output.n37 gnd 0.011243f
C285 output.n38 gnd 0.006041f
C286 output.n39 gnd 0.006397f
C287 output.n40 gnd 0.01428f
C288 output.n41 gnd 0.030913f
C289 output.n42 gnd 0.006397f
C290 output.n43 gnd 0.006041f
C291 output.n44 gnd 0.025987f
C292 output.n45 gnd 0.097665f
C293 output.n46 gnd 0.015803f
C294 output.n47 gnd 0.011243f
C295 output.n48 gnd 0.006041f
C296 output.n49 gnd 0.01428f
C297 output.n50 gnd 0.006397f
C298 output.n51 gnd 0.011243f
C299 output.n52 gnd 0.006041f
C300 output.n53 gnd 0.01428f
C301 output.n54 gnd 0.006397f
C302 output.n55 gnd 0.048111f
C303 output.t19 gnd 0.023274f
C304 output.n56 gnd 0.01071f
C305 output.n57 gnd 0.008435f
C306 output.n58 gnd 0.006041f
C307 output.n59 gnd 0.267512f
C308 output.n60 gnd 0.011243f
C309 output.n61 gnd 0.006041f
C310 output.n62 gnd 0.006397f
C311 output.n63 gnd 0.01428f
C312 output.n64 gnd 0.01428f
C313 output.n65 gnd 0.006397f
C314 output.n66 gnd 0.006041f
C315 output.n67 gnd 0.011243f
C316 output.n68 gnd 0.011243f
C317 output.n69 gnd 0.006041f
C318 output.n70 gnd 0.006397f
C319 output.n71 gnd 0.01428f
C320 output.n72 gnd 0.030913f
C321 output.n73 gnd 0.006397f
C322 output.n74 gnd 0.006041f
C323 output.n75 gnd 0.025987f
C324 output.n76 gnd 0.09306f
C325 output.n77 gnd 1.65264f
C326 output.n78 gnd 0.015803f
C327 output.n79 gnd 0.011243f
C328 output.n80 gnd 0.006041f
C329 output.n81 gnd 0.01428f
C330 output.n82 gnd 0.006397f
C331 output.n83 gnd 0.011243f
C332 output.n84 gnd 0.006041f
C333 output.n85 gnd 0.01428f
C334 output.n86 gnd 0.006397f
C335 output.n87 gnd 0.048111f
C336 output.t17 gnd 0.023274f
C337 output.n88 gnd 0.01071f
C338 output.n89 gnd 0.008435f
C339 output.n90 gnd 0.006041f
C340 output.n91 gnd 0.267512f
C341 output.n92 gnd 0.011243f
C342 output.n93 gnd 0.006041f
C343 output.n94 gnd 0.006397f
C344 output.n95 gnd 0.01428f
C345 output.n96 gnd 0.01428f
C346 output.n97 gnd 0.006397f
C347 output.n98 gnd 0.006041f
C348 output.n99 gnd 0.011243f
C349 output.n100 gnd 0.011243f
C350 output.n101 gnd 0.006041f
C351 output.n102 gnd 0.006397f
C352 output.n103 gnd 0.01428f
C353 output.n104 gnd 0.030913f
C354 output.n105 gnd 0.006397f
C355 output.n106 gnd 0.006041f
C356 output.n107 gnd 0.025987f
C357 output.n108 gnd 0.09306f
C358 output.n109 gnd 0.713089f
C359 output.n110 gnd 0.015803f
C360 output.n111 gnd 0.011243f
C361 output.n112 gnd 0.006041f
C362 output.n113 gnd 0.01428f
C363 output.n114 gnd 0.006397f
C364 output.n115 gnd 0.011243f
C365 output.n116 gnd 0.006041f
C366 output.n117 gnd 0.01428f
C367 output.n118 gnd 0.006397f
C368 output.n119 gnd 0.048111f
C369 output.t16 gnd 0.023274f
C370 output.n120 gnd 0.01071f
C371 output.n121 gnd 0.008435f
C372 output.n122 gnd 0.006041f
C373 output.n123 gnd 0.267512f
C374 output.n124 gnd 0.011243f
C375 output.n125 gnd 0.006041f
C376 output.n126 gnd 0.006397f
C377 output.n127 gnd 0.01428f
C378 output.n128 gnd 0.01428f
C379 output.n129 gnd 0.006397f
C380 output.n130 gnd 0.006041f
C381 output.n131 gnd 0.011243f
C382 output.n132 gnd 0.011243f
C383 output.n133 gnd 0.006041f
C384 output.n134 gnd 0.006397f
C385 output.n135 gnd 0.01428f
C386 output.n136 gnd 0.030913f
C387 output.n137 gnd 0.006397f
C388 output.n138 gnd 0.006041f
C389 output.n139 gnd 0.025987f
C390 output.n140 gnd 0.09306f
C391 output.n141 gnd 1.67353f
C392 a_n2318_8322.t1 gnd 39.602997f
C393 a_n2318_8322.t3 gnd 29.1868f
C394 a_n2318_8322.t2 gnd 19.7318f
C395 a_n2318_8322.t0 gnd 39.602997f
C396 a_n2318_8322.t25 gnd 0.896865f
C397 a_n2318_8322.t22 gnd 0.095784f
C398 a_n2318_8322.t19 gnd 0.095784f
C399 a_n2318_8322.n0 gnd 0.674698f
C400 a_n2318_8322.n1 gnd 0.753878f
C401 a_n2318_8322.t16 gnd 0.095784f
C402 a_n2318_8322.t27 gnd 0.095784f
C403 a_n2318_8322.n2 gnd 0.674698f
C404 a_n2318_8322.n3 gnd 0.383035f
C405 a_n2318_8322.t24 gnd 0.095784f
C406 a_n2318_8322.t17 gnd 0.095784f
C407 a_n2318_8322.n4 gnd 0.674698f
C408 a_n2318_8322.n5 gnd 0.383035f
C409 a_n2318_8322.t15 gnd 0.895081f
C410 a_n2318_8322.n6 gnd 0.881139f
C411 a_n2318_8322.n7 gnd 3.71089f
C412 a_n2318_8322.t7 gnd 0.896867f
C413 a_n2318_8322.t11 gnd 0.095784f
C414 a_n2318_8322.t10 gnd 0.095784f
C415 a_n2318_8322.n8 gnd 0.674698f
C416 a_n2318_8322.n9 gnd 0.753876f
C417 a_n2318_8322.t5 gnd 0.895081f
C418 a_n2318_8322.n10 gnd 0.379361f
C419 a_n2318_8322.t8 gnd 0.895081f
C420 a_n2318_8322.n11 gnd 0.379361f
C421 a_n2318_8322.t6 gnd 0.095784f
C422 a_n2318_8322.t4 gnd 0.095784f
C423 a_n2318_8322.n12 gnd 0.674698f
C424 a_n2318_8322.n13 gnd 0.383035f
C425 a_n2318_8322.t9 gnd 0.895081f
C426 a_n2318_8322.n14 gnd 1.07426f
C427 a_n2318_8322.n15 gnd 1.82616f
C428 a_n2318_8322.t12 gnd 0.895081f
C429 a_n2318_8322.n16 gnd 1.55131f
C430 a_n2318_8322.t21 gnd 0.095784f
C431 a_n2318_8322.t20 gnd 0.095784f
C432 a_n2318_8322.n17 gnd 0.674698f
C433 a_n2318_8322.n18 gnd 0.383035f
C434 a_n2318_8322.t23 gnd 0.095784f
C435 a_n2318_8322.t18 gnd 0.095784f
C436 a_n2318_8322.n19 gnd 0.674698f
C437 a_n2318_8322.n20 gnd 0.383035f
C438 a_n2318_8322.t14 gnd 0.095784f
C439 a_n2318_8322.t13 gnd 0.095784f
C440 a_n2318_8322.n21 gnd 0.674698f
C441 a_n2318_8322.n22 gnd 0.753876f
C442 a_n2318_8322.t26 gnd 0.896867f
C443 a_n3106_n452.t9 gnd 0.10001f
C444 a_n3106_n452.t20 gnd 1.03942f
C445 a_n3106_n452.n0 gnd 0.392946f
C446 a_n3106_n452.t54 gnd 1.29145f
C447 a_n3106_n452.n1 gnd 1.22854f
C448 a_n3106_n452.t33 gnd 1.03942f
C449 a_n3106_n452.n2 gnd 0.392946f
C450 a_n3106_n452.t43 gnd 0.10001f
C451 a_n3106_n452.t55 gnd 0.10001f
C452 a_n3106_n452.n3 gnd 0.816794f
C453 a_n3106_n452.n4 gnd 0.411618f
C454 a_n3106_n452.t40 gnd 0.10001f
C455 a_n3106_n452.t27 gnd 0.10001f
C456 a_n3106_n452.n5 gnd 0.816794f
C457 a_n3106_n452.n6 gnd 0.411618f
C458 a_n3106_n452.t28 gnd 0.10001f
C459 a_n3106_n452.t39 gnd 0.10001f
C460 a_n3106_n452.n7 gnd 0.816794f
C461 a_n3106_n452.n8 gnd 0.411618f
C462 a_n3106_n452.t0 gnd 0.10001f
C463 a_n3106_n452.t48 gnd 0.10001f
C464 a_n3106_n452.n9 gnd 0.816794f
C465 a_n3106_n452.n10 gnd 0.411618f
C466 a_n3106_n452.t46 gnd 0.10001f
C467 a_n3106_n452.t36 gnd 0.10001f
C468 a_n3106_n452.n11 gnd 0.816794f
C469 a_n3106_n452.n12 gnd 0.411618f
C470 a_n3106_n452.t38 gnd 1.03942f
C471 a_n3106_n452.n13 gnd 0.972974f
C472 a_n3106_n452.t30 gnd 1.29145f
C473 a_n3106_n452.n14 gnd 0.909591f
C474 a_n3106_n452.t51 gnd 1.29145f
C475 a_n3106_n452.n15 gnd 0.909591f
C476 a_n3106_n452.t32 gnd 1.29145f
C477 a_n3106_n452.n16 gnd 0.909591f
C478 a_n3106_n452.t50 gnd 1.29145f
C479 a_n3106_n452.n17 gnd 0.909591f
C480 a_n3106_n452.t49 gnd 1.29145f
C481 a_n3106_n452.n18 gnd 0.909591f
C482 a_n3106_n452.t35 gnd 1.29145f
C483 a_n3106_n452.n19 gnd 0.909591f
C484 a_n3106_n452.t53 gnd 1.29145f
C485 a_n3106_n452.n20 gnd 0.789472f
C486 a_n3106_n452.n21 gnd 0.948419f
C487 a_n3106_n452.t11 gnd 1.03941f
C488 a_n3106_n452.n22 gnd 0.645631f
C489 a_n3106_n452.t8 gnd 0.10001f
C490 a_n3106_n452.t25 gnd 0.10001f
C491 a_n3106_n452.n23 gnd 0.816793f
C492 a_n3106_n452.n24 gnd 0.41162f
C493 a_n3106_n452.t19 gnd 0.10001f
C494 a_n3106_n452.t23 gnd 0.10001f
C495 a_n3106_n452.n25 gnd 0.816793f
C496 a_n3106_n452.n26 gnd 0.41162f
C497 a_n3106_n452.t24 gnd 0.10001f
C498 a_n3106_n452.t12 gnd 0.10001f
C499 a_n3106_n452.n27 gnd 0.816793f
C500 a_n3106_n452.n28 gnd 0.41162f
C501 a_n3106_n452.t13 gnd 0.10001f
C502 a_n3106_n452.t4 gnd 0.10001f
C503 a_n3106_n452.n29 gnd 0.816793f
C504 a_n3106_n452.n30 gnd 0.41162f
C505 a_n3106_n452.t6 gnd 0.10001f
C506 a_n3106_n452.t22 gnd 0.10001f
C507 a_n3106_n452.n31 gnd 0.816793f
C508 a_n3106_n452.n32 gnd 0.41162f
C509 a_n3106_n452.t17 gnd 1.03941f
C510 a_n3106_n452.n33 gnd 0.39295f
C511 a_n3106_n452.t2 gnd 1.03941f
C512 a_n3106_n452.n34 gnd 0.39295f
C513 a_n3106_n452.t44 gnd 0.10001f
C514 a_n3106_n452.t37 gnd 0.10001f
C515 a_n3106_n452.n35 gnd 0.816793f
C516 a_n3106_n452.n36 gnd 0.41162f
C517 a_n3106_n452.t41 gnd 0.10001f
C518 a_n3106_n452.t29 gnd 0.10001f
C519 a_n3106_n452.n37 gnd 0.816793f
C520 a_n3106_n452.n38 gnd 0.41162f
C521 a_n3106_n452.t1 gnd 0.10001f
C522 a_n3106_n452.t31 gnd 0.10001f
C523 a_n3106_n452.n39 gnd 0.816793f
C524 a_n3106_n452.n40 gnd 0.41162f
C525 a_n3106_n452.t34 gnd 0.10001f
C526 a_n3106_n452.t52 gnd 0.10001f
C527 a_n3106_n452.n41 gnd 0.816793f
C528 a_n3106_n452.n42 gnd 0.41162f
C529 a_n3106_n452.t47 gnd 0.10001f
C530 a_n3106_n452.t45 gnd 0.10001f
C531 a_n3106_n452.n43 gnd 0.816793f
C532 a_n3106_n452.n44 gnd 0.41162f
C533 a_n3106_n452.t42 gnd 1.03941f
C534 a_n3106_n452.n45 gnd 0.645631f
C535 a_n3106_n452.n46 gnd 1.05146f
C536 a_n3106_n452.t7 gnd 1.03941f
C537 a_n3106_n452.n47 gnd 0.972978f
C538 a_n3106_n452.t5 gnd 0.10001f
C539 a_n3106_n452.t3 gnd 0.10001f
C540 a_n3106_n452.n48 gnd 0.816794f
C541 a_n3106_n452.n49 gnd 0.411618f
C542 a_n3106_n452.t16 gnd 0.10001f
C543 a_n3106_n452.t21 gnd 0.10001f
C544 a_n3106_n452.n50 gnd 0.816794f
C545 a_n3106_n452.n51 gnd 0.411618f
C546 a_n3106_n452.t14 gnd 0.10001f
C547 a_n3106_n452.t18 gnd 0.10001f
C548 a_n3106_n452.n52 gnd 0.816794f
C549 a_n3106_n452.n53 gnd 0.411618f
C550 a_n3106_n452.t10 gnd 0.10001f
C551 a_n3106_n452.t15 gnd 0.10001f
C552 a_n3106_n452.n54 gnd 0.816794f
C553 a_n3106_n452.n55 gnd 0.411618f
C554 a_n3106_n452.n56 gnd 0.411617f
C555 a_n3106_n452.n57 gnd 0.816796f
C556 a_n3106_n452.t26 gnd 0.10001f
C557 plus.n0 gnd 0.022838f
C558 plus.t20 gnd 0.415311f
C559 plus.t23 gnd 0.384014f
C560 plus.n1 gnd 0.155312f
C561 plus.n2 gnd 0.022838f
C562 plus.t6 gnd 0.384014f
C563 plus.n3 gnd 0.019515f
C564 plus.n4 gnd 0.022838f
C565 plus.t12 gnd 0.384014f
C566 plus.t8 gnd 0.384014f
C567 plus.n5 gnd 0.155312f
C568 plus.n6 gnd 0.022838f
C569 plus.t7 gnd 0.384014f
C570 plus.n7 gnd 0.155312f
C571 plus.n8 gnd 0.022838f
C572 plus.t19 gnd 0.384014f
C573 plus.n9 gnd 0.018562f
C574 plus.n10 gnd 0.022838f
C575 plus.t18 gnd 0.384014f
C576 plus.t27 gnd 0.384014f
C577 plus.n11 gnd 0.155312f
C578 plus.n12 gnd 0.022838f
C579 plus.t25 gnd 0.384014f
C580 plus.n13 gnd 0.155312f
C581 plus.n14 gnd 0.096921f
C582 plus.t9 gnd 0.384014f
C583 plus.t14 gnd 0.429589f
C584 plus.n15 gnd 0.181575f
C585 plus.n16 gnd 0.177861f
C586 plus.n17 gnd 0.029263f
C587 plus.n18 gnd 0.025844f
C588 plus.n19 gnd 0.022838f
C589 plus.n20 gnd 0.022838f
C590 plus.n21 gnd 0.027291f
C591 plus.n22 gnd 0.019515f
C592 plus.n23 gnd 0.029743f
C593 plus.n24 gnd 0.022838f
C594 plus.n25 gnd 0.022838f
C595 plus.n26 gnd 0.028408f
C596 plus.n27 gnd 0.026698f
C597 plus.n28 gnd 0.155312f
C598 plus.n29 gnd 0.028608f
C599 plus.n30 gnd 0.022838f
C600 plus.n31 gnd 0.022838f
C601 plus.n32 gnd 0.022838f
C602 plus.n33 gnd 0.02938f
C603 plus.n34 gnd 0.155312f
C604 plus.n35 gnd 0.027553f
C605 plus.n36 gnd 0.027553f
C606 plus.n37 gnd 0.022838f
C607 plus.n38 gnd 0.022838f
C608 plus.n39 gnd 0.02938f
C609 plus.n40 gnd 0.018562f
C610 plus.n41 gnd 0.028608f
C611 plus.n42 gnd 0.022838f
C612 plus.n43 gnd 0.022838f
C613 plus.n44 gnd 0.026698f
C614 plus.n45 gnd 0.028408f
C615 plus.n46 gnd 0.155312f
C616 plus.n47 gnd 0.029743f
C617 plus.n48 gnd 0.022838f
C618 plus.n49 gnd 0.022838f
C619 plus.n50 gnd 0.022838f
C620 plus.n51 gnd 0.027291f
C621 plus.n52 gnd 0.155312f
C622 plus.n53 gnd 0.025844f
C623 plus.n54 gnd 0.029263f
C624 plus.n55 gnd 0.022838f
C625 plus.n56 gnd 0.022838f
C626 plus.n57 gnd 0.029793f
C627 plus.n58 gnd 0.0083f
C628 plus.n59 gnd 0.179825f
C629 plus.n60 gnd 0.261661f
C630 plus.n61 gnd 0.022838f
C631 plus.t28 gnd 0.384014f
C632 plus.n62 gnd 0.155312f
C633 plus.n63 gnd 0.022838f
C634 plus.t26 gnd 0.384014f
C635 plus.n64 gnd 0.019515f
C636 plus.n65 gnd 0.022838f
C637 plus.t10 gnd 0.384014f
C638 plus.t15 gnd 0.384014f
C639 plus.n66 gnd 0.155312f
C640 plus.n67 gnd 0.022838f
C641 plus.t13 gnd 0.384014f
C642 plus.n68 gnd 0.155312f
C643 plus.n69 gnd 0.022838f
C644 plus.t17 gnd 0.384014f
C645 plus.n70 gnd 0.018562f
C646 plus.n71 gnd 0.022838f
C647 plus.t16 gnd 0.384014f
C648 plus.t21 gnd 0.384014f
C649 plus.n72 gnd 0.155312f
C650 plus.n73 gnd 0.022838f
C651 plus.t22 gnd 0.384014f
C652 plus.n74 gnd 0.155312f
C653 plus.n75 gnd 0.096921f
C654 plus.t5 gnd 0.384014f
C655 plus.t11 gnd 0.429589f
C656 plus.n76 gnd 0.181575f
C657 plus.n77 gnd 0.177861f
C658 plus.n78 gnd 0.029263f
C659 plus.n79 gnd 0.025844f
C660 plus.n80 gnd 0.022838f
C661 plus.n81 gnd 0.022838f
C662 plus.n82 gnd 0.027291f
C663 plus.n83 gnd 0.019515f
C664 plus.n84 gnd 0.029743f
C665 plus.n85 gnd 0.022838f
C666 plus.n86 gnd 0.022838f
C667 plus.n87 gnd 0.028408f
C668 plus.n88 gnd 0.026698f
C669 plus.n89 gnd 0.155312f
C670 plus.n90 gnd 0.028608f
C671 plus.n91 gnd 0.022838f
C672 plus.n92 gnd 0.022838f
C673 plus.n93 gnd 0.022838f
C674 plus.n94 gnd 0.02938f
C675 plus.n95 gnd 0.155312f
C676 plus.n96 gnd 0.027553f
C677 plus.n97 gnd 0.027553f
C678 plus.n98 gnd 0.022838f
C679 plus.n99 gnd 0.022838f
C680 plus.n100 gnd 0.02938f
C681 plus.n101 gnd 0.018562f
C682 plus.n102 gnd 0.028608f
C683 plus.n103 gnd 0.022838f
C684 plus.n104 gnd 0.022838f
C685 plus.n105 gnd 0.026698f
C686 plus.n106 gnd 0.028408f
C687 plus.n107 gnd 0.155312f
C688 plus.n108 gnd 0.029743f
C689 plus.n109 gnd 0.022838f
C690 plus.n110 gnd 0.022838f
C691 plus.n111 gnd 0.022838f
C692 plus.n112 gnd 0.027291f
C693 plus.n113 gnd 0.155312f
C694 plus.n114 gnd 0.025844f
C695 plus.n115 gnd 0.029263f
C696 plus.n116 gnd 0.022838f
C697 plus.n117 gnd 0.022838f
C698 plus.n118 gnd 0.029793f
C699 plus.n119 gnd 0.0083f
C700 plus.t24 gnd 0.415311f
C701 plus.n120 gnd 0.179825f
C702 plus.n121 gnd 0.823978f
C703 plus.n122 gnd 1.21471f
C704 plus.t1 gnd 0.039425f
C705 plus.t2 gnd 0.00704f
C706 plus.t4 gnd 0.00704f
C707 plus.n123 gnd 0.022833f
C708 plus.n124 gnd 0.177252f
C709 plus.t3 gnd 0.00704f
C710 plus.t0 gnd 0.00704f
C711 plus.n125 gnd 0.022833f
C712 plus.n126 gnd 0.133049f
C713 plus.n127 gnd 3.03081f
C714 outputibias.t8 gnd 0.11477f
C715 outputibias.t9 gnd 0.115567f
C716 outputibias.n0 gnd 0.130108f
C717 outputibias.n1 gnd 0.001372f
C718 outputibias.n2 gnd 9.76e-19
C719 outputibias.n3 gnd 5.24e-19
C720 outputibias.n4 gnd 0.001239f
C721 outputibias.n5 gnd 5.55e-19
C722 outputibias.n6 gnd 9.76e-19
C723 outputibias.n7 gnd 5.24e-19
C724 outputibias.n8 gnd 0.001239f
C725 outputibias.n9 gnd 5.55e-19
C726 outputibias.n10 gnd 0.004176f
C727 outputibias.t7 gnd 0.00202f
C728 outputibias.n11 gnd 9.3e-19
C729 outputibias.n12 gnd 7.32e-19
C730 outputibias.n13 gnd 5.24e-19
C731 outputibias.n14 gnd 0.02322f
C732 outputibias.n15 gnd 9.76e-19
C733 outputibias.n16 gnd 5.24e-19
C734 outputibias.n17 gnd 5.55e-19
C735 outputibias.n18 gnd 0.001239f
C736 outputibias.n19 gnd 0.001239f
C737 outputibias.n20 gnd 5.55e-19
C738 outputibias.n21 gnd 5.24e-19
C739 outputibias.n22 gnd 9.76e-19
C740 outputibias.n23 gnd 9.76e-19
C741 outputibias.n24 gnd 5.24e-19
C742 outputibias.n25 gnd 5.55e-19
C743 outputibias.n26 gnd 0.001239f
C744 outputibias.n27 gnd 0.002683f
C745 outputibias.n28 gnd 5.55e-19
C746 outputibias.n29 gnd 5.24e-19
C747 outputibias.n30 gnd 0.002256f
C748 outputibias.n31 gnd 0.005781f
C749 outputibias.n32 gnd 0.001372f
C750 outputibias.n33 gnd 9.76e-19
C751 outputibias.n34 gnd 5.24e-19
C752 outputibias.n35 gnd 0.001239f
C753 outputibias.n36 gnd 5.55e-19
C754 outputibias.n37 gnd 9.76e-19
C755 outputibias.n38 gnd 5.24e-19
C756 outputibias.n39 gnd 0.001239f
C757 outputibias.n40 gnd 5.55e-19
C758 outputibias.n41 gnd 0.004176f
C759 outputibias.t1 gnd 0.00202f
C760 outputibias.n42 gnd 9.3e-19
C761 outputibias.n43 gnd 7.32e-19
C762 outputibias.n44 gnd 5.24e-19
C763 outputibias.n45 gnd 0.02322f
C764 outputibias.n46 gnd 9.76e-19
C765 outputibias.n47 gnd 5.24e-19
C766 outputibias.n48 gnd 5.55e-19
C767 outputibias.n49 gnd 0.001239f
C768 outputibias.n50 gnd 0.001239f
C769 outputibias.n51 gnd 5.55e-19
C770 outputibias.n52 gnd 5.24e-19
C771 outputibias.n53 gnd 9.76e-19
C772 outputibias.n54 gnd 9.76e-19
C773 outputibias.n55 gnd 5.24e-19
C774 outputibias.n56 gnd 5.55e-19
C775 outputibias.n57 gnd 0.001239f
C776 outputibias.n58 gnd 0.002683f
C777 outputibias.n59 gnd 5.55e-19
C778 outputibias.n60 gnd 5.24e-19
C779 outputibias.n61 gnd 0.002256f
C780 outputibias.n62 gnd 0.005197f
C781 outputibias.n63 gnd 0.121892f
C782 outputibias.n64 gnd 0.001372f
C783 outputibias.n65 gnd 9.76e-19
C784 outputibias.n66 gnd 5.24e-19
C785 outputibias.n67 gnd 0.001239f
C786 outputibias.n68 gnd 5.55e-19
C787 outputibias.n69 gnd 9.76e-19
C788 outputibias.n70 gnd 5.24e-19
C789 outputibias.n71 gnd 0.001239f
C790 outputibias.n72 gnd 5.55e-19
C791 outputibias.n73 gnd 0.004176f
C792 outputibias.t3 gnd 0.00202f
C793 outputibias.n74 gnd 9.3e-19
C794 outputibias.n75 gnd 7.32e-19
C795 outputibias.n76 gnd 5.24e-19
C796 outputibias.n77 gnd 0.02322f
C797 outputibias.n78 gnd 9.76e-19
C798 outputibias.n79 gnd 5.24e-19
C799 outputibias.n80 gnd 5.55e-19
C800 outputibias.n81 gnd 0.001239f
C801 outputibias.n82 gnd 0.001239f
C802 outputibias.n83 gnd 5.55e-19
C803 outputibias.n84 gnd 5.24e-19
C804 outputibias.n85 gnd 9.76e-19
C805 outputibias.n86 gnd 9.76e-19
C806 outputibias.n87 gnd 5.24e-19
C807 outputibias.n88 gnd 5.55e-19
C808 outputibias.n89 gnd 0.001239f
C809 outputibias.n90 gnd 0.002683f
C810 outputibias.n91 gnd 5.55e-19
C811 outputibias.n92 gnd 5.24e-19
C812 outputibias.n93 gnd 0.002256f
C813 outputibias.n94 gnd 0.005197f
C814 outputibias.n95 gnd 0.064513f
C815 outputibias.n96 gnd 0.001372f
C816 outputibias.n97 gnd 9.76e-19
C817 outputibias.n98 gnd 5.24e-19
C818 outputibias.n99 gnd 0.001239f
C819 outputibias.n100 gnd 5.55e-19
C820 outputibias.n101 gnd 9.76e-19
C821 outputibias.n102 gnd 5.24e-19
C822 outputibias.n103 gnd 0.001239f
C823 outputibias.n104 gnd 5.55e-19
C824 outputibias.n105 gnd 0.004176f
C825 outputibias.t5 gnd 0.00202f
C826 outputibias.n106 gnd 9.3e-19
C827 outputibias.n107 gnd 7.32e-19
C828 outputibias.n108 gnd 5.24e-19
C829 outputibias.n109 gnd 0.02322f
C830 outputibias.n110 gnd 9.76e-19
C831 outputibias.n111 gnd 5.24e-19
C832 outputibias.n112 gnd 5.55e-19
C833 outputibias.n113 gnd 0.001239f
C834 outputibias.n114 gnd 0.001239f
C835 outputibias.n115 gnd 5.55e-19
C836 outputibias.n116 gnd 5.24e-19
C837 outputibias.n117 gnd 9.76e-19
C838 outputibias.n118 gnd 9.76e-19
C839 outputibias.n119 gnd 5.24e-19
C840 outputibias.n120 gnd 5.55e-19
C841 outputibias.n121 gnd 0.001239f
C842 outputibias.n122 gnd 0.002683f
C843 outputibias.n123 gnd 5.55e-19
C844 outputibias.n124 gnd 5.24e-19
C845 outputibias.n125 gnd 0.002256f
C846 outputibias.n126 gnd 0.005197f
C847 outputibias.n127 gnd 0.084814f
C848 outputibias.t4 gnd 0.108319f
C849 outputibias.t2 gnd 0.108319f
C850 outputibias.t0 gnd 0.108319f
C851 outputibias.t6 gnd 0.109238f
C852 outputibias.n128 gnd 0.134674f
C853 outputibias.n129 gnd 0.07244f
C854 outputibias.n130 gnd 0.079818f
C855 outputibias.n131 gnd 0.164901f
C856 outputibias.t11 gnd 0.11477f
C857 outputibias.n132 gnd 0.067481f
C858 outputibias.t10 gnd 0.11477f
C859 outputibias.n133 gnd 0.065115f
C860 outputibias.n134 gnd 0.029159f
C861 a_n2140_13878.t21 gnd 0.186868f
C862 a_n2140_13878.t19 gnd 0.186868f
C863 a_n2140_13878.t23 gnd 0.186868f
C864 a_n2140_13878.n0 gnd 1.47386f
C865 a_n2140_13878.t8 gnd 0.186868f
C866 a_n2140_13878.t16 gnd 0.186868f
C867 a_n2140_13878.n1 gnd 1.47143f
C868 a_n2140_13878.n2 gnd 1.32263f
C869 a_n2140_13878.t18 gnd 0.186868f
C870 a_n2140_13878.t13 gnd 0.186868f
C871 a_n2140_13878.n3 gnd 1.47299f
C872 a_n2140_13878.t10 gnd 0.186868f
C873 a_n2140_13878.t12 gnd 0.186868f
C874 a_n2140_13878.n4 gnd 1.47143f
C875 a_n2140_13878.n5 gnd 2.05603f
C876 a_n2140_13878.t20 gnd 0.186868f
C877 a_n2140_13878.t11 gnd 0.186868f
C878 a_n2140_13878.n6 gnd 1.47143f
C879 a_n2140_13878.n7 gnd 1.00289f
C880 a_n2140_13878.t17 gnd 0.186868f
C881 a_n2140_13878.t9 gnd 0.186868f
C882 a_n2140_13878.n8 gnd 1.47143f
C883 a_n2140_13878.n9 gnd 4.06212f
C884 a_n2140_13878.t1 gnd 1.74974f
C885 a_n2140_13878.t4 gnd 0.186868f
C886 a_n2140_13878.t5 gnd 0.186868f
C887 a_n2140_13878.n10 gnd 1.3163f
C888 a_n2140_13878.n11 gnd 1.47077f
C889 a_n2140_13878.t0 gnd 1.74626f
C890 a_n2140_13878.n12 gnd 0.740113f
C891 a_n2140_13878.t3 gnd 1.74626f
C892 a_n2140_13878.n13 gnd 0.740113f
C893 a_n2140_13878.t6 gnd 0.186868f
C894 a_n2140_13878.t7 gnd 0.186868f
C895 a_n2140_13878.n14 gnd 1.3163f
C896 a_n2140_13878.n15 gnd 0.74728f
C897 a_n2140_13878.t2 gnd 1.74626f
C898 a_n2140_13878.n16 gnd 2.09583f
C899 a_n2140_13878.n17 gnd 2.85974f
C900 a_n2140_13878.t14 gnd 0.186868f
C901 a_n2140_13878.t15 gnd 0.186868f
C902 a_n2140_13878.n18 gnd 1.47142f
C903 a_n2140_13878.n19 gnd 2.01665f
C904 a_n2140_13878.n20 gnd 0.651948f
C905 a_n2140_13878.n21 gnd 1.47143f
C906 a_n2140_13878.t22 gnd 0.186868f
C907 a_n2848_n452.n0 gnd 4.35918f
C908 a_n2848_n452.n1 gnd 3.11675f
C909 a_n2848_n452.n2 gnd 3.98565f
C910 a_n2848_n452.n3 gnd 0.903102f
C911 a_n2848_n452.n4 gnd 0.903104f
C912 a_n2848_n452.n5 gnd 0.661444f
C913 a_n2848_n452.n6 gnd 2.95991f
C914 a_n2848_n452.n7 gnd 0.213645f
C915 a_n2848_n452.n8 gnd 0.739044f
C916 a_n2848_n452.n9 gnd 0.213645f
C917 a_n2848_n452.n10 gnd 0.439089f
C918 a_n2848_n452.n11 gnd 0.545911f
C919 a_n2848_n452.n12 gnd 0.66142f
C920 a_n2848_n452.n13 gnd 0.202714f
C921 a_n2848_n452.n14 gnd 0.149302f
C922 a_n2848_n452.n15 gnd 0.234656f
C923 a_n2848_n452.n16 gnd 0.181245f
C924 a_n2848_n452.n17 gnd 0.202714f
C925 a_n2848_n452.n18 gnd 1.10633f
C926 a_n2848_n452.n19 gnd 0.149302f
C927 a_n2848_n452.n20 gnd 0.714831f
C928 a_n2848_n452.n21 gnd 0.506946f
C929 a_n2848_n452.n22 gnd 0.213645f
C930 a_n2848_n452.n23 gnd 0.213645f
C931 a_n2848_n452.n24 gnd 0.439089f
C932 a_n2848_n452.n25 gnd 0.213645f
C933 a_n2848_n452.n26 gnd 0.213645f
C934 a_n2848_n452.n27 gnd 1.75891f
C935 a_n2848_n452.n28 gnd 2.057f
C936 a_n2848_n452.n29 gnd 1.87737f
C937 a_n2848_n452.n30 gnd 1.75891f
C938 a_n2848_n452.n31 gnd 0.282224f
C939 a_n2848_n452.n32 gnd 0.751876f
C940 a_n2848_n452.n33 gnd 0.004802f
C941 a_n2848_n452.n34 gnd 0.010385f
C942 a_n2848_n452.n35 gnd 0.010385f
C943 a_n2848_n452.n36 gnd 0.004802f
C944 a_n2848_n452.n37 gnd 0.282224f
C945 a_n2848_n452.n38 gnd 0.282224f
C946 a_n2848_n452.n39 gnd 0.439089f
C947 a_n2848_n452.n40 gnd 0.004802f
C948 a_n2848_n452.n41 gnd 0.010385f
C949 a_n2848_n452.n42 gnd 0.010385f
C950 a_n2848_n452.n43 gnd 0.004802f
C951 a_n2848_n452.n44 gnd 0.282224f
C952 a_n2848_n452.n45 gnd 0.008272f
C953 a_n2848_n452.n46 gnd 0.282224f
C954 a_n2848_n452.n47 gnd 0.008272f
C955 a_n2848_n452.n48 gnd 0.282224f
C956 a_n2848_n452.n49 gnd 0.008272f
C957 a_n2848_n452.n50 gnd 0.282224f
C958 a_n2848_n452.n51 gnd 0.008272f
C959 a_n2848_n452.n52 gnd 0.282224f
C960 a_n2848_n452.n53 gnd 0.004802f
C961 a_n2848_n452.n54 gnd 0.282224f
C962 a_n2848_n452.n55 gnd 0.282224f
C963 a_n2848_n452.n56 gnd 0.004802f
C964 a_n2848_n452.n57 gnd 0.010385f
C965 a_n2848_n452.n58 gnd 0.010385f
C966 a_n2848_n452.n59 gnd 0.004802f
C967 a_n2848_n452.n60 gnd 0.282224f
C968 a_n2848_n452.n61 gnd 0.282224f
C969 a_n2848_n452.n62 gnd 0.004802f
C970 a_n2848_n452.t12 gnd 0.70084f
C971 a_n2848_n452.t28 gnd 0.689291f
C972 a_n2848_n452.t16 gnd 0.689291f
C973 a_n2848_n452.n64 gnd 0.299372f
C974 a_n2848_n452.t30 gnd 0.689291f
C975 a_n2848_n452.t24 gnd 0.689291f
C976 a_n2848_n452.t34 gnd 0.115256f
C977 a_n2848_n452.t49 gnd 0.115256f
C978 a_n2848_n452.n65 gnd 1.02144f
C979 a_n2848_n452.t42 gnd 0.115256f
C980 a_n2848_n452.t46 gnd 0.115256f
C981 a_n2848_n452.n66 gnd 1.01844f
C982 a_n2848_n452.t37 gnd 0.115256f
C983 a_n2848_n452.t1 gnd 0.115256f
C984 a_n2848_n452.n67 gnd 1.01844f
C985 a_n2848_n452.t50 gnd 0.115256f
C986 a_n2848_n452.t47 gnd 0.115256f
C987 a_n2848_n452.n68 gnd 1.02144f
C988 a_n2848_n452.t54 gnd 0.115256f
C989 a_n2848_n452.t52 gnd 0.115256f
C990 a_n2848_n452.n69 gnd 1.01844f
C991 a_n2848_n452.t38 gnd 0.115256f
C992 a_n2848_n452.t40 gnd 0.115256f
C993 a_n2848_n452.n70 gnd 1.01844f
C994 a_n2848_n452.t43 gnd 0.115256f
C995 a_n2848_n452.t51 gnd 0.115256f
C996 a_n2848_n452.n71 gnd 1.01844f
C997 a_n2848_n452.t41 gnd 0.115256f
C998 a_n2848_n452.t0 gnd 0.115256f
C999 a_n2848_n452.n72 gnd 1.01844f
C1000 a_n2848_n452.t53 gnd 0.115256f
C1001 a_n2848_n452.t36 gnd 0.115256f
C1002 a_n2848_n452.n73 gnd 1.01844f
C1003 a_n2848_n452.t55 gnd 0.115256f
C1004 a_n2848_n452.t39 gnd 0.115256f
C1005 a_n2848_n452.n74 gnd 1.02145f
C1006 a_n2848_n452.t35 gnd 0.115256f
C1007 a_n2848_n452.t48 gnd 0.115256f
C1008 a_n2848_n452.n75 gnd 1.01844f
C1009 a_n2848_n452.t44 gnd 0.115256f
C1010 a_n2848_n452.t45 gnd 0.115256f
C1011 a_n2848_n452.n76 gnd 1.01844f
C1012 a_n2848_n452.t26 gnd 0.689291f
C1013 a_n2848_n452.n77 gnd 0.299372f
C1014 a_n2848_n452.t4 gnd 0.689291f
C1015 a_n2848_n452.t2 gnd 0.70084f
C1016 a_n2848_n452.t86 gnd 0.70084f
C1017 a_n2848_n452.t67 gnd 0.689291f
C1018 a_n2848_n452.t71 gnd 0.689291f
C1019 a_n2848_n452.n78 gnd 0.301107f
C1020 a_n2848_n452.t61 gnd 0.689291f
C1021 a_n2848_n452.t76 gnd 0.689291f
C1022 a_n2848_n452.t83 gnd 0.689291f
C1023 a_n2848_n452.n79 gnd 0.301107f
C1024 a_n2848_n452.t84 gnd 0.689291f
C1025 a_n2848_n452.t58 gnd 0.70084f
C1026 a_n2848_n452.t9 gnd 1.38754f
C1027 a_n2848_n452.t19 gnd 0.148186f
C1028 a_n2848_n452.t11 gnd 0.148186f
C1029 a_n2848_n452.n80 gnd 1.04382f
C1030 a_n2848_n452.t21 gnd 0.148186f
C1031 a_n2848_n452.t15 gnd 0.148186f
C1032 a_n2848_n452.n81 gnd 1.04382f
C1033 a_n2848_n452.t23 gnd 0.148186f
C1034 a_n2848_n452.t33 gnd 0.148186f
C1035 a_n2848_n452.n82 gnd 1.04382f
C1036 a_n2848_n452.t7 gnd 1.38477f
C1037 a_n2848_n452.t22 gnd 0.689291f
C1038 a_n2848_n452.n83 gnd 0.301107f
C1039 a_n2848_n452.t20 gnd 0.689291f
C1040 a_n2848_n452.t8 gnd 0.70084f
C1041 a_n2848_n452.t18 gnd 0.689291f
C1042 a_n2848_n452.t66 gnd 0.689291f
C1043 a_n2848_n452.n84 gnd 0.301107f
C1044 a_n2848_n452.t80 gnd 0.689291f
C1045 a_n2848_n452.t82 gnd 0.70084f
C1046 a_n2848_n452.t60 gnd 0.689291f
C1047 a_n2848_n452.n85 gnd 0.303562f
C1048 a_n2848_n452.t79 gnd 0.689291f
C1049 a_n2848_n452.n86 gnd 0.301107f
C1050 a_n2848_n452.n87 gnd 0.296573f
C1051 a_n2848_n452.t57 gnd 0.689291f
C1052 a_n2848_n452.n88 gnd 0.296573f
C1053 a_n2848_n452.t75 gnd 0.689291f
C1054 a_n2848_n452.n89 gnd 0.303562f
C1055 a_n2848_n452.t59 gnd 0.70084f
C1056 a_n2848_n452.n90 gnd 0.303562f
C1057 a_n2848_n452.t10 gnd 0.689291f
C1058 a_n2848_n452.n91 gnd 0.301107f
C1059 a_n2848_n452.n92 gnd 0.296573f
C1060 a_n2848_n452.t14 gnd 0.689291f
C1061 a_n2848_n452.n93 gnd 0.296573f
C1062 a_n2848_n452.t32 gnd 0.689291f
C1063 a_n2848_n452.n94 gnd 0.303562f
C1064 a_n2848_n452.t6 gnd 0.70084f
C1065 a_n2848_n452.n95 gnd 1.18578f
C1066 a_n2848_n452.t64 gnd 0.689291f
C1067 a_n2848_n452.n96 gnd 0.299207f
C1068 a_n2848_n452.t70 gnd 0.689291f
C1069 a_n2848_n452.n97 gnd 0.299207f
C1070 a_n2848_n452.t62 gnd 0.689291f
C1071 a_n2848_n452.n98 gnd 0.299207f
C1072 a_n2848_n452.t74 gnd 0.689291f
C1073 a_n2848_n452.n99 gnd 0.299207f
C1074 a_n2848_n452.t65 gnd 0.689291f
C1075 a_n2848_n452.n100 gnd 0.293774f
C1076 a_n2848_n452.t87 gnd 0.689291f
C1077 a_n2848_n452.n101 gnd 0.303056f
C1078 a_n2848_n452.t68 gnd 0.70084f
C1079 a_n2848_n452.t77 gnd 0.689291f
C1080 a_n2848_n452.n102 gnd 0.293774f
C1081 a_n2848_n452.t63 gnd 0.689291f
C1082 a_n2848_n452.n103 gnd 0.303056f
C1083 a_n2848_n452.t72 gnd 0.70084f
C1084 a_n2848_n452.t81 gnd 0.689291f
C1085 a_n2848_n452.n104 gnd 0.293774f
C1086 a_n2848_n452.t69 gnd 0.689291f
C1087 a_n2848_n452.n105 gnd 0.303056f
C1088 a_n2848_n452.t85 gnd 0.70084f
C1089 a_n2848_n452.t73 gnd 0.689291f
C1090 a_n2848_n452.n106 gnd 0.293774f
C1091 a_n2848_n452.t56 gnd 0.689291f
C1092 a_n2848_n452.n107 gnd 0.303056f
C1093 a_n2848_n452.t78 gnd 0.70084f
C1094 a_n2848_n452.n108 gnd 1.4348f
C1095 a_n2848_n452.n109 gnd 0.303562f
C1096 a_n2848_n452.n110 gnd 0.296573f
C1097 a_n2848_n452.n111 gnd 0.296573f
C1098 a_n2848_n452.n112 gnd 0.303562f
C1099 a_n2848_n452.n113 gnd 0.303562f
C1100 a_n2848_n452.n114 gnd 0.01212f
C1101 a_n2848_n452.n115 gnd 0.296573f
C1102 a_n2848_n452.n116 gnd 0.296573f
C1103 a_n2848_n452.n117 gnd 0.01212f
C1104 a_n2848_n452.n118 gnd 0.303562f
C1105 a_n2848_n452.n119 gnd 0.850479f
C1106 a_n2848_n452.t13 gnd 1.38478f
C1107 a_n2848_n452.t29 gnd 0.148186f
C1108 a_n2848_n452.t17 gnd 0.148186f
C1109 a_n2848_n452.n120 gnd 1.04382f
C1110 a_n2848_n452.t31 gnd 0.148186f
C1111 a_n2848_n452.t25 gnd 0.148186f
C1112 a_n2848_n452.n121 gnd 1.04382f
C1113 a_n2848_n452.t27 gnd 0.148186f
C1114 a_n2848_n452.t5 gnd 0.148186f
C1115 a_n2848_n452.n122 gnd 1.04382f
C1116 a_n2848_n452.t3 gnd 1.38754f
C1117 vdd.t119 gnd 0.034504f
C1118 vdd.t235 gnd 0.034504f
C1119 vdd.n0 gnd 0.272138f
C1120 vdd.t111 gnd 0.034504f
C1121 vdd.t125 gnd 0.034504f
C1122 vdd.n1 gnd 0.271688f
C1123 vdd.n2 gnd 0.250549f
C1124 vdd.t231 gnd 0.034504f
C1125 vdd.t98 gnd 0.034504f
C1126 vdd.n3 gnd 0.271688f
C1127 vdd.n4 gnd 0.126712f
C1128 vdd.t100 gnd 0.034504f
C1129 vdd.t121 gnd 0.034504f
C1130 vdd.n5 gnd 0.271688f
C1131 vdd.n6 gnd 0.118896f
C1132 vdd.t107 gnd 0.034504f
C1133 vdd.t233 gnd 0.034504f
C1134 vdd.n7 gnd 0.272138f
C1135 vdd.t123 gnd 0.034504f
C1136 vdd.t117 gnd 0.034504f
C1137 vdd.n8 gnd 0.271688f
C1138 vdd.n9 gnd 0.250549f
C1139 vdd.t127 gnd 0.034504f
C1140 vdd.t103 gnd 0.034504f
C1141 vdd.n10 gnd 0.271688f
C1142 vdd.n11 gnd 0.126712f
C1143 vdd.t115 gnd 0.034504f
C1144 vdd.t130 gnd 0.034504f
C1145 vdd.n12 gnd 0.271688f
C1146 vdd.n13 gnd 0.118896f
C1147 vdd.n14 gnd 0.084057f
C1148 vdd.t92 gnd 0.019169f
C1149 vdd.t91 gnd 0.019169f
C1150 vdd.n15 gnd 0.176441f
C1151 vdd.t86 gnd 0.019169f
C1152 vdd.t83 gnd 0.019169f
C1153 vdd.n16 gnd 0.175925f
C1154 vdd.n17 gnd 0.306164f
C1155 vdd.t85 gnd 0.019169f
C1156 vdd.t89 gnd 0.019169f
C1157 vdd.n18 gnd 0.175925f
C1158 vdd.n19 gnd 0.126664f
C1159 vdd.t81 gnd 0.019169f
C1160 vdd.t82 gnd 0.019169f
C1161 vdd.n20 gnd 0.176441f
C1162 vdd.t90 gnd 0.019169f
C1163 vdd.t94 gnd 0.019169f
C1164 vdd.n21 gnd 0.175925f
C1165 vdd.n22 gnd 0.306164f
C1166 vdd.t84 gnd 0.019169f
C1167 vdd.t96 gnd 0.019169f
C1168 vdd.n23 gnd 0.175925f
C1169 vdd.n24 gnd 0.126664f
C1170 vdd.t87 gnd 0.019169f
C1171 vdd.t95 gnd 0.019169f
C1172 vdd.n25 gnd 0.175925f
C1173 vdd.t88 gnd 0.019169f
C1174 vdd.t93 gnd 0.019169f
C1175 vdd.n26 gnd 0.175925f
C1176 vdd.n27 gnd 20.4786f
C1177 vdd.n28 gnd 7.7028f
C1178 vdd.n29 gnd 0.005228f
C1179 vdd.n30 gnd 0.004851f
C1180 vdd.n31 gnd 0.002684f
C1181 vdd.n32 gnd 0.006162f
C1182 vdd.n33 gnd 0.002607f
C1183 vdd.n34 gnd 0.00276f
C1184 vdd.n35 gnd 0.004851f
C1185 vdd.n36 gnd 0.002607f
C1186 vdd.n37 gnd 0.006162f
C1187 vdd.n38 gnd 0.00276f
C1188 vdd.n39 gnd 0.004851f
C1189 vdd.n40 gnd 0.002607f
C1190 vdd.n41 gnd 0.004621f
C1191 vdd.n42 gnd 0.004635f
C1192 vdd.t160 gnd 0.013238f
C1193 vdd.n43 gnd 0.029455f
C1194 vdd.n44 gnd 0.153291f
C1195 vdd.n45 gnd 0.002607f
C1196 vdd.n46 gnd 0.00276f
C1197 vdd.n47 gnd 0.006162f
C1198 vdd.n48 gnd 0.006162f
C1199 vdd.n49 gnd 0.00276f
C1200 vdd.n50 gnd 0.002607f
C1201 vdd.n51 gnd 0.004851f
C1202 vdd.n52 gnd 0.004851f
C1203 vdd.n53 gnd 0.002607f
C1204 vdd.n54 gnd 0.00276f
C1205 vdd.n55 gnd 0.006162f
C1206 vdd.n56 gnd 0.006162f
C1207 vdd.n57 gnd 0.00276f
C1208 vdd.n58 gnd 0.002607f
C1209 vdd.n59 gnd 0.004851f
C1210 vdd.n60 gnd 0.004851f
C1211 vdd.n61 gnd 0.002607f
C1212 vdd.n62 gnd 0.00276f
C1213 vdd.n63 gnd 0.006162f
C1214 vdd.n64 gnd 0.006162f
C1215 vdd.n65 gnd 0.014568f
C1216 vdd.n66 gnd 0.002684f
C1217 vdd.n67 gnd 0.002607f
C1218 vdd.n68 gnd 0.012539f
C1219 vdd.n69 gnd 0.008754f
C1220 vdd.t213 gnd 0.03067f
C1221 vdd.t180 gnd 0.03067f
C1222 vdd.n70 gnd 0.210786f
C1223 vdd.n71 gnd 0.165751f
C1224 vdd.t223 gnd 0.03067f
C1225 vdd.t210 gnd 0.03067f
C1226 vdd.n72 gnd 0.210786f
C1227 vdd.n73 gnd 0.13376f
C1228 vdd.t139 gnd 0.03067f
C1229 vdd.t173 gnd 0.03067f
C1230 vdd.n74 gnd 0.210786f
C1231 vdd.n75 gnd 0.13376f
C1232 vdd.t147 gnd 0.03067f
C1233 vdd.t188 gnd 0.03067f
C1234 vdd.n76 gnd 0.210786f
C1235 vdd.n77 gnd 0.13376f
C1236 vdd.t168 gnd 0.03067f
C1237 vdd.t216 gnd 0.03067f
C1238 vdd.n78 gnd 0.210786f
C1239 vdd.n79 gnd 0.13376f
C1240 vdd.n80 gnd 0.005228f
C1241 vdd.n81 gnd 0.004851f
C1242 vdd.n82 gnd 0.002684f
C1243 vdd.n83 gnd 0.006162f
C1244 vdd.n84 gnd 0.002607f
C1245 vdd.n85 gnd 0.00276f
C1246 vdd.n86 gnd 0.004851f
C1247 vdd.n87 gnd 0.002607f
C1248 vdd.n88 gnd 0.006162f
C1249 vdd.n89 gnd 0.00276f
C1250 vdd.n90 gnd 0.004851f
C1251 vdd.n91 gnd 0.002607f
C1252 vdd.n92 gnd 0.004621f
C1253 vdd.n93 gnd 0.004635f
C1254 vdd.t152 gnd 0.013238f
C1255 vdd.n94 gnd 0.029455f
C1256 vdd.n95 gnd 0.153291f
C1257 vdd.n96 gnd 0.002607f
C1258 vdd.n97 gnd 0.00276f
C1259 vdd.n98 gnd 0.006162f
C1260 vdd.n99 gnd 0.006162f
C1261 vdd.n100 gnd 0.00276f
C1262 vdd.n101 gnd 0.002607f
C1263 vdd.n102 gnd 0.004851f
C1264 vdd.n103 gnd 0.004851f
C1265 vdd.n104 gnd 0.002607f
C1266 vdd.n105 gnd 0.00276f
C1267 vdd.n106 gnd 0.006162f
C1268 vdd.n107 gnd 0.006162f
C1269 vdd.n108 gnd 0.00276f
C1270 vdd.n109 gnd 0.002607f
C1271 vdd.n110 gnd 0.004851f
C1272 vdd.n111 gnd 0.004851f
C1273 vdd.n112 gnd 0.002607f
C1274 vdd.n113 gnd 0.00276f
C1275 vdd.n114 gnd 0.006162f
C1276 vdd.n115 gnd 0.006162f
C1277 vdd.n116 gnd 0.014568f
C1278 vdd.n117 gnd 0.002684f
C1279 vdd.n118 gnd 0.002607f
C1280 vdd.n119 gnd 0.012539f
C1281 vdd.n120 gnd 0.00848f
C1282 vdd.n121 gnd 0.099518f
C1283 vdd.n122 gnd 0.005228f
C1284 vdd.n123 gnd 0.004851f
C1285 vdd.n124 gnd 0.002684f
C1286 vdd.n125 gnd 0.006162f
C1287 vdd.n126 gnd 0.002607f
C1288 vdd.n127 gnd 0.00276f
C1289 vdd.n128 gnd 0.004851f
C1290 vdd.n129 gnd 0.002607f
C1291 vdd.n130 gnd 0.006162f
C1292 vdd.n131 gnd 0.00276f
C1293 vdd.n132 gnd 0.004851f
C1294 vdd.n133 gnd 0.002607f
C1295 vdd.n134 gnd 0.004621f
C1296 vdd.n135 gnd 0.004635f
C1297 vdd.t186 gnd 0.013238f
C1298 vdd.n136 gnd 0.029455f
C1299 vdd.n137 gnd 0.153291f
C1300 vdd.n138 gnd 0.002607f
C1301 vdd.n139 gnd 0.00276f
C1302 vdd.n140 gnd 0.006162f
C1303 vdd.n141 gnd 0.006162f
C1304 vdd.n142 gnd 0.00276f
C1305 vdd.n143 gnd 0.002607f
C1306 vdd.n144 gnd 0.004851f
C1307 vdd.n145 gnd 0.004851f
C1308 vdd.n146 gnd 0.002607f
C1309 vdd.n147 gnd 0.00276f
C1310 vdd.n148 gnd 0.006162f
C1311 vdd.n149 gnd 0.006162f
C1312 vdd.n150 gnd 0.00276f
C1313 vdd.n151 gnd 0.002607f
C1314 vdd.n152 gnd 0.004851f
C1315 vdd.n153 gnd 0.004851f
C1316 vdd.n154 gnd 0.002607f
C1317 vdd.n155 gnd 0.00276f
C1318 vdd.n156 gnd 0.006162f
C1319 vdd.n157 gnd 0.006162f
C1320 vdd.n158 gnd 0.014568f
C1321 vdd.n159 gnd 0.002684f
C1322 vdd.n160 gnd 0.002607f
C1323 vdd.n161 gnd 0.012539f
C1324 vdd.n162 gnd 0.008754f
C1325 vdd.t205 gnd 0.03067f
C1326 vdd.t135 gnd 0.03067f
C1327 vdd.n163 gnd 0.210786f
C1328 vdd.n164 gnd 0.165751f
C1329 vdd.t170 gnd 0.03067f
C1330 vdd.t172 gnd 0.03067f
C1331 vdd.n165 gnd 0.210786f
C1332 vdd.n166 gnd 0.13376f
C1333 vdd.t220 gnd 0.03067f
C1334 vdd.t165 gnd 0.03067f
C1335 vdd.n167 gnd 0.210786f
C1336 vdd.n168 gnd 0.13376f
C1337 vdd.t166 gnd 0.03067f
C1338 vdd.t218 gnd 0.03067f
C1339 vdd.n169 gnd 0.210786f
C1340 vdd.n170 gnd 0.13376f
C1341 vdd.t219 gnd 0.03067f
C1342 vdd.t145 gnd 0.03067f
C1343 vdd.n171 gnd 0.210786f
C1344 vdd.n172 gnd 0.13376f
C1345 vdd.n173 gnd 0.005228f
C1346 vdd.n174 gnd 0.004851f
C1347 vdd.n175 gnd 0.002684f
C1348 vdd.n176 gnd 0.006162f
C1349 vdd.n177 gnd 0.002607f
C1350 vdd.n178 gnd 0.00276f
C1351 vdd.n179 gnd 0.004851f
C1352 vdd.n180 gnd 0.002607f
C1353 vdd.n181 gnd 0.006162f
C1354 vdd.n182 gnd 0.00276f
C1355 vdd.n183 gnd 0.004851f
C1356 vdd.n184 gnd 0.002607f
C1357 vdd.n185 gnd 0.004621f
C1358 vdd.n186 gnd 0.004635f
C1359 vdd.t206 gnd 0.013238f
C1360 vdd.n187 gnd 0.029455f
C1361 vdd.n188 gnd 0.153291f
C1362 vdd.n189 gnd 0.002607f
C1363 vdd.n190 gnd 0.00276f
C1364 vdd.n191 gnd 0.006162f
C1365 vdd.n192 gnd 0.006162f
C1366 vdd.n193 gnd 0.00276f
C1367 vdd.n194 gnd 0.002607f
C1368 vdd.n195 gnd 0.004851f
C1369 vdd.n196 gnd 0.004851f
C1370 vdd.n197 gnd 0.002607f
C1371 vdd.n198 gnd 0.00276f
C1372 vdd.n199 gnd 0.006162f
C1373 vdd.n200 gnd 0.006162f
C1374 vdd.n201 gnd 0.00276f
C1375 vdd.n202 gnd 0.002607f
C1376 vdd.n203 gnd 0.004851f
C1377 vdd.n204 gnd 0.004851f
C1378 vdd.n205 gnd 0.002607f
C1379 vdd.n206 gnd 0.00276f
C1380 vdd.n207 gnd 0.006162f
C1381 vdd.n208 gnd 0.006162f
C1382 vdd.n209 gnd 0.014568f
C1383 vdd.n210 gnd 0.002684f
C1384 vdd.n211 gnd 0.002607f
C1385 vdd.n212 gnd 0.012539f
C1386 vdd.n213 gnd 0.00848f
C1387 vdd.n214 gnd 0.059203f
C1388 vdd.n215 gnd 0.213325f
C1389 vdd.n216 gnd 0.005228f
C1390 vdd.n217 gnd 0.004851f
C1391 vdd.n218 gnd 0.002684f
C1392 vdd.n219 gnd 0.006162f
C1393 vdd.n220 gnd 0.002607f
C1394 vdd.n221 gnd 0.00276f
C1395 vdd.n222 gnd 0.004851f
C1396 vdd.n223 gnd 0.002607f
C1397 vdd.n224 gnd 0.006162f
C1398 vdd.n225 gnd 0.00276f
C1399 vdd.n226 gnd 0.004851f
C1400 vdd.n227 gnd 0.002607f
C1401 vdd.n228 gnd 0.004621f
C1402 vdd.n229 gnd 0.004635f
C1403 vdd.t197 gnd 0.013238f
C1404 vdd.n230 gnd 0.029455f
C1405 vdd.n231 gnd 0.153291f
C1406 vdd.n232 gnd 0.002607f
C1407 vdd.n233 gnd 0.00276f
C1408 vdd.n234 gnd 0.006162f
C1409 vdd.n235 gnd 0.006162f
C1410 vdd.n236 gnd 0.00276f
C1411 vdd.n237 gnd 0.002607f
C1412 vdd.n238 gnd 0.004851f
C1413 vdd.n239 gnd 0.004851f
C1414 vdd.n240 gnd 0.002607f
C1415 vdd.n241 gnd 0.00276f
C1416 vdd.n242 gnd 0.006162f
C1417 vdd.n243 gnd 0.006162f
C1418 vdd.n244 gnd 0.00276f
C1419 vdd.n245 gnd 0.002607f
C1420 vdd.n246 gnd 0.004851f
C1421 vdd.n247 gnd 0.004851f
C1422 vdd.n248 gnd 0.002607f
C1423 vdd.n249 gnd 0.00276f
C1424 vdd.n250 gnd 0.006162f
C1425 vdd.n251 gnd 0.006162f
C1426 vdd.n252 gnd 0.014568f
C1427 vdd.n253 gnd 0.002684f
C1428 vdd.n254 gnd 0.002607f
C1429 vdd.n255 gnd 0.012539f
C1430 vdd.n256 gnd 0.008754f
C1431 vdd.t211 gnd 0.03067f
C1432 vdd.t150 gnd 0.03067f
C1433 vdd.n257 gnd 0.210786f
C1434 vdd.n258 gnd 0.165751f
C1435 vdd.t183 gnd 0.03067f
C1436 vdd.t185 gnd 0.03067f
C1437 vdd.n259 gnd 0.210786f
C1438 vdd.n260 gnd 0.13376f
C1439 vdd.t227 gnd 0.03067f
C1440 vdd.t178 gnd 0.03067f
C1441 vdd.n261 gnd 0.210786f
C1442 vdd.n262 gnd 0.13376f
C1443 vdd.t179 gnd 0.03067f
C1444 vdd.t225 gnd 0.03067f
C1445 vdd.n263 gnd 0.210786f
C1446 vdd.n264 gnd 0.13376f
C1447 vdd.t226 gnd 0.03067f
C1448 vdd.t158 gnd 0.03067f
C1449 vdd.n265 gnd 0.210786f
C1450 vdd.n266 gnd 0.13376f
C1451 vdd.n267 gnd 0.005228f
C1452 vdd.n268 gnd 0.004851f
C1453 vdd.n269 gnd 0.002684f
C1454 vdd.n270 gnd 0.006162f
C1455 vdd.n271 gnd 0.002607f
C1456 vdd.n272 gnd 0.00276f
C1457 vdd.n273 gnd 0.004851f
C1458 vdd.n274 gnd 0.002607f
C1459 vdd.n275 gnd 0.006162f
C1460 vdd.n276 gnd 0.00276f
C1461 vdd.n277 gnd 0.004851f
C1462 vdd.n278 gnd 0.002607f
C1463 vdd.n279 gnd 0.004621f
C1464 vdd.n280 gnd 0.004635f
C1465 vdd.t215 gnd 0.013238f
C1466 vdd.n281 gnd 0.029455f
C1467 vdd.n282 gnd 0.153291f
C1468 vdd.n283 gnd 0.002607f
C1469 vdd.n284 gnd 0.00276f
C1470 vdd.n285 gnd 0.006162f
C1471 vdd.n286 gnd 0.006162f
C1472 vdd.n287 gnd 0.00276f
C1473 vdd.n288 gnd 0.002607f
C1474 vdd.n289 gnd 0.004851f
C1475 vdd.n290 gnd 0.004851f
C1476 vdd.n291 gnd 0.002607f
C1477 vdd.n292 gnd 0.00276f
C1478 vdd.n293 gnd 0.006162f
C1479 vdd.n294 gnd 0.006162f
C1480 vdd.n295 gnd 0.00276f
C1481 vdd.n296 gnd 0.002607f
C1482 vdd.n297 gnd 0.004851f
C1483 vdd.n298 gnd 0.004851f
C1484 vdd.n299 gnd 0.002607f
C1485 vdd.n300 gnd 0.00276f
C1486 vdd.n301 gnd 0.006162f
C1487 vdd.n302 gnd 0.006162f
C1488 vdd.n303 gnd 0.014568f
C1489 vdd.n304 gnd 0.002684f
C1490 vdd.n305 gnd 0.002607f
C1491 vdd.n306 gnd 0.012539f
C1492 vdd.n307 gnd 0.00848f
C1493 vdd.n308 gnd 0.059203f
C1494 vdd.n309 gnd 0.234451f
C1495 vdd.n310 gnd 0.009494f
C1496 vdd.n311 gnd 0.009494f
C1497 vdd.n312 gnd 0.007668f
C1498 vdd.n313 gnd 0.007668f
C1499 vdd.n314 gnd 0.009526f
C1500 vdd.n315 gnd 0.009526f
C1501 vdd.t138 gnd 0.486772f
C1502 vdd.n316 gnd 0.009526f
C1503 vdd.n317 gnd 0.009526f
C1504 vdd.n318 gnd 0.009526f
C1505 vdd.t146 gnd 0.486772f
C1506 vdd.n319 gnd 0.009526f
C1507 vdd.n320 gnd 0.009526f
C1508 vdd.n321 gnd 0.009526f
C1509 vdd.n322 gnd 0.009526f
C1510 vdd.n323 gnd 0.007668f
C1511 vdd.n324 gnd 0.009526f
C1512 vdd.n325 gnd 0.783703f
C1513 vdd.n326 gnd 0.009526f
C1514 vdd.n327 gnd 0.009526f
C1515 vdd.n328 gnd 0.009526f
C1516 vdd.n329 gnd 0.666878f
C1517 vdd.n330 gnd 0.009526f
C1518 vdd.n331 gnd 0.009526f
C1519 vdd.n332 gnd 0.009526f
C1520 vdd.n333 gnd 0.009526f
C1521 vdd.n334 gnd 0.009526f
C1522 vdd.n335 gnd 0.007668f
C1523 vdd.n336 gnd 0.009526f
C1524 vdd.t144 gnd 0.486772f
C1525 vdd.n337 gnd 0.009526f
C1526 vdd.n338 gnd 0.009526f
C1527 vdd.n339 gnd 0.009526f
C1528 vdd.n340 gnd 0.973544f
C1529 vdd.n341 gnd 0.009526f
C1530 vdd.n342 gnd 0.009526f
C1531 vdd.n343 gnd 0.009526f
C1532 vdd.n344 gnd 0.009526f
C1533 vdd.n345 gnd 0.009526f
C1534 vdd.n346 gnd 0.007668f
C1535 vdd.n347 gnd 0.009526f
C1536 vdd.n348 gnd 0.009526f
C1537 vdd.n349 gnd 0.009526f
C1538 vdd.n350 gnd 0.02245f
C1539 vdd.n351 gnd 2.23915f
C1540 vdd.n352 gnd 0.0228f
C1541 vdd.n353 gnd 0.009526f
C1542 vdd.n354 gnd 0.009526f
C1543 vdd.n356 gnd 0.009526f
C1544 vdd.n357 gnd 0.009526f
C1545 vdd.n358 gnd 0.007668f
C1546 vdd.n359 gnd 0.007668f
C1547 vdd.n360 gnd 0.009526f
C1548 vdd.n361 gnd 0.009526f
C1549 vdd.n362 gnd 0.009526f
C1550 vdd.n363 gnd 0.009526f
C1551 vdd.n364 gnd 0.009526f
C1552 vdd.n365 gnd 0.009526f
C1553 vdd.n366 gnd 0.007668f
C1554 vdd.n368 gnd 0.009526f
C1555 vdd.n369 gnd 0.009526f
C1556 vdd.n370 gnd 0.009526f
C1557 vdd.n371 gnd 0.009526f
C1558 vdd.n372 gnd 0.009526f
C1559 vdd.n373 gnd 0.007668f
C1560 vdd.n375 gnd 0.009526f
C1561 vdd.n376 gnd 0.009526f
C1562 vdd.n377 gnd 0.009526f
C1563 vdd.n378 gnd 0.009526f
C1564 vdd.n379 gnd 0.009526f
C1565 vdd.n380 gnd 0.007668f
C1566 vdd.n382 gnd 0.009526f
C1567 vdd.n383 gnd 0.009526f
C1568 vdd.n384 gnd 0.009526f
C1569 vdd.n385 gnd 0.009526f
C1570 vdd.n386 gnd 0.006402f
C1571 vdd.t79 gnd 0.117199f
C1572 vdd.t78 gnd 0.125253f
C1573 vdd.t77 gnd 0.15306f
C1574 vdd.n387 gnd 0.196201f
C1575 vdd.n388 gnd 0.165611f
C1576 vdd.n390 gnd 0.009526f
C1577 vdd.n391 gnd 0.009526f
C1578 vdd.n392 gnd 0.007668f
C1579 vdd.n393 gnd 0.009526f
C1580 vdd.n395 gnd 0.009526f
C1581 vdd.n396 gnd 0.009526f
C1582 vdd.n397 gnd 0.009526f
C1583 vdd.n398 gnd 0.009526f
C1584 vdd.n399 gnd 0.007668f
C1585 vdd.n401 gnd 0.009526f
C1586 vdd.n402 gnd 0.009526f
C1587 vdd.n403 gnd 0.009526f
C1588 vdd.n404 gnd 0.009526f
C1589 vdd.n405 gnd 0.009526f
C1590 vdd.n406 gnd 0.007668f
C1591 vdd.n408 gnd 0.009526f
C1592 vdd.n409 gnd 0.009526f
C1593 vdd.n410 gnd 0.009526f
C1594 vdd.n411 gnd 0.009526f
C1595 vdd.n412 gnd 0.009526f
C1596 vdd.n413 gnd 0.007668f
C1597 vdd.n415 gnd 0.009526f
C1598 vdd.n416 gnd 0.009526f
C1599 vdd.n417 gnd 0.009526f
C1600 vdd.n418 gnd 0.009526f
C1601 vdd.n419 gnd 0.009526f
C1602 vdd.n420 gnd 0.007668f
C1603 vdd.n422 gnd 0.009526f
C1604 vdd.n423 gnd 0.009526f
C1605 vdd.n424 gnd 0.009526f
C1606 vdd.n425 gnd 0.009526f
C1607 vdd.n426 gnd 0.007591f
C1608 vdd.t73 gnd 0.117199f
C1609 vdd.t72 gnd 0.125253f
C1610 vdd.t71 gnd 0.15306f
C1611 vdd.n427 gnd 0.196201f
C1612 vdd.n428 gnd 0.165611f
C1613 vdd.n430 gnd 0.009526f
C1614 vdd.n431 gnd 0.009526f
C1615 vdd.n432 gnd 0.007668f
C1616 vdd.n433 gnd 0.009526f
C1617 vdd.n435 gnd 0.009526f
C1618 vdd.n436 gnd 0.009526f
C1619 vdd.n437 gnd 0.009526f
C1620 vdd.n438 gnd 0.009526f
C1621 vdd.n439 gnd 0.007668f
C1622 vdd.n441 gnd 0.009526f
C1623 vdd.n442 gnd 0.009526f
C1624 vdd.n443 gnd 0.009526f
C1625 vdd.n444 gnd 0.009526f
C1626 vdd.n445 gnd 0.009526f
C1627 vdd.n446 gnd 0.007668f
C1628 vdd.n448 gnd 0.009526f
C1629 vdd.n449 gnd 0.009526f
C1630 vdd.n450 gnd 0.009526f
C1631 vdd.n451 gnd 0.009526f
C1632 vdd.n452 gnd 0.009526f
C1633 vdd.n453 gnd 0.007668f
C1634 vdd.n455 gnd 0.009526f
C1635 vdd.n456 gnd 0.009526f
C1636 vdd.n457 gnd 0.009526f
C1637 vdd.n458 gnd 0.009526f
C1638 vdd.n459 gnd 0.009526f
C1639 vdd.n460 gnd 0.007668f
C1640 vdd.n462 gnd 0.009526f
C1641 vdd.n463 gnd 0.009526f
C1642 vdd.n464 gnd 0.009526f
C1643 vdd.n465 gnd 0.009526f
C1644 vdd.n466 gnd 0.009526f
C1645 vdd.n467 gnd 0.009526f
C1646 vdd.n468 gnd 0.007668f
C1647 vdd.n469 gnd 0.009526f
C1648 vdd.n470 gnd 0.009526f
C1649 vdd.n471 gnd 0.007668f
C1650 vdd.n472 gnd 0.009526f
C1651 vdd.n473 gnd 0.009526f
C1652 vdd.n474 gnd 0.007668f
C1653 vdd.n475 gnd 0.009526f
C1654 vdd.n476 gnd 0.007668f
C1655 vdd.n477 gnd 0.009526f
C1656 vdd.n478 gnd 0.007668f
C1657 vdd.n479 gnd 0.009526f
C1658 vdd.n480 gnd 0.009526f
C1659 vdd.t171 gnd 0.486772f
C1660 vdd.n481 gnd 0.520846f
C1661 vdd.n482 gnd 0.009526f
C1662 vdd.n483 gnd 0.007668f
C1663 vdd.n484 gnd 0.009526f
C1664 vdd.n485 gnd 0.007668f
C1665 vdd.n486 gnd 0.009526f
C1666 vdd.t169 gnd 0.486772f
C1667 vdd.n487 gnd 0.009526f
C1668 vdd.n488 gnd 0.007668f
C1669 vdd.n489 gnd 0.009526f
C1670 vdd.n490 gnd 0.007668f
C1671 vdd.n491 gnd 0.009526f
C1672 vdd.n492 gnd 0.764232f
C1673 vdd.n493 gnd 0.808041f
C1674 vdd.t134 gnd 0.486772f
C1675 vdd.n494 gnd 0.009526f
C1676 vdd.n495 gnd 0.007668f
C1677 vdd.n496 gnd 0.009526f
C1678 vdd.n497 gnd 0.007668f
C1679 vdd.n498 gnd 0.009526f
C1680 vdd.n499 gnd 0.598729f
C1681 vdd.n500 gnd 0.009526f
C1682 vdd.n501 gnd 0.007668f
C1683 vdd.n502 gnd 0.009526f
C1684 vdd.n503 gnd 0.007668f
C1685 vdd.n504 gnd 0.009526f
C1686 vdd.n505 gnd 0.973544f
C1687 vdd.t159 gnd 0.486772f
C1688 vdd.n506 gnd 0.009526f
C1689 vdd.n507 gnd 0.007668f
C1690 vdd.n508 gnd 0.009526f
C1691 vdd.n509 gnd 0.007668f
C1692 vdd.n510 gnd 0.009526f
C1693 vdd.n511 gnd 0.520846f
C1694 vdd.n512 gnd 0.009526f
C1695 vdd.n513 gnd 0.007668f
C1696 vdd.n514 gnd 0.0228f
C1697 vdd.n515 gnd 0.0228f
C1698 vdd.n516 gnd 8.58666f
C1699 vdd.t13 gnd 0.486772f
C1700 vdd.n517 gnd 0.0228f
C1701 vdd.n518 gnd 0.008193f
C1702 vdd.n519 gnd 0.007668f
C1703 vdd.n524 gnd 0.006097f
C1704 vdd.n525 gnd 0.007668f
C1705 vdd.n526 gnd 0.009526f
C1706 vdd.n527 gnd 0.009526f
C1707 vdd.n528 gnd 0.009526f
C1708 vdd.n529 gnd 0.009526f
C1709 vdd.n530 gnd 0.009526f
C1710 vdd.n531 gnd 0.007668f
C1711 vdd.n532 gnd 0.009526f
C1712 vdd.n533 gnd 0.009526f
C1713 vdd.n534 gnd 0.009526f
C1714 vdd.n535 gnd 0.009526f
C1715 vdd.n536 gnd 0.009526f
C1716 vdd.n537 gnd 0.007668f
C1717 vdd.n538 gnd 0.009526f
C1718 vdd.n539 gnd 0.009526f
C1719 vdd.n540 gnd 0.009526f
C1720 vdd.n541 gnd 0.009526f
C1721 vdd.n542 gnd 0.009526f
C1722 vdd.t42 gnd 0.117199f
C1723 vdd.t43 gnd 0.125253f
C1724 vdd.t41 gnd 0.15306f
C1725 vdd.n543 gnd 0.196201f
C1726 vdd.n544 gnd 0.164844f
C1727 vdd.n545 gnd 0.015642f
C1728 vdd.n546 gnd 0.009526f
C1729 vdd.n547 gnd 0.009526f
C1730 vdd.n548 gnd 0.009526f
C1731 vdd.n549 gnd 0.009526f
C1732 vdd.n550 gnd 0.009526f
C1733 vdd.n551 gnd 0.007668f
C1734 vdd.n552 gnd 0.009526f
C1735 vdd.n553 gnd 0.009526f
C1736 vdd.n554 gnd 0.009526f
C1737 vdd.n555 gnd 0.009526f
C1738 vdd.n556 gnd 0.009526f
C1739 vdd.n557 gnd 0.007668f
C1740 vdd.n558 gnd 0.009526f
C1741 vdd.n559 gnd 0.009526f
C1742 vdd.n560 gnd 0.009526f
C1743 vdd.n561 gnd 0.009526f
C1744 vdd.n562 gnd 0.009526f
C1745 vdd.n563 gnd 0.007668f
C1746 vdd.n564 gnd 0.009526f
C1747 vdd.n565 gnd 0.009526f
C1748 vdd.n566 gnd 0.009526f
C1749 vdd.n567 gnd 0.009526f
C1750 vdd.n568 gnd 0.009526f
C1751 vdd.n569 gnd 0.007668f
C1752 vdd.n570 gnd 0.009526f
C1753 vdd.n571 gnd 0.009526f
C1754 vdd.n572 gnd 0.009526f
C1755 vdd.n573 gnd 0.009526f
C1756 vdd.n574 gnd 0.009526f
C1757 vdd.n575 gnd 0.007668f
C1758 vdd.n576 gnd 0.009526f
C1759 vdd.n577 gnd 0.009526f
C1760 vdd.n578 gnd 0.009526f
C1761 vdd.n579 gnd 0.007591f
C1762 vdd.t29 gnd 0.117199f
C1763 vdd.t30 gnd 0.125253f
C1764 vdd.t28 gnd 0.15306f
C1765 vdd.n580 gnd 0.196201f
C1766 vdd.n581 gnd 0.164844f
C1767 vdd.n582 gnd 0.009526f
C1768 vdd.n583 gnd 0.007668f
C1769 vdd.n585 gnd 0.009526f
C1770 vdd.n587 gnd 0.009526f
C1771 vdd.n588 gnd 0.009526f
C1772 vdd.n589 gnd 0.007668f
C1773 vdd.n590 gnd 0.009526f
C1774 vdd.n591 gnd 0.009526f
C1775 vdd.n592 gnd 0.009526f
C1776 vdd.n593 gnd 0.009526f
C1777 vdd.n594 gnd 0.009526f
C1778 vdd.n595 gnd 0.007668f
C1779 vdd.n596 gnd 0.009526f
C1780 vdd.n597 gnd 0.009526f
C1781 vdd.n598 gnd 0.009526f
C1782 vdd.n599 gnd 0.009526f
C1783 vdd.n600 gnd 0.009526f
C1784 vdd.n601 gnd 0.007668f
C1785 vdd.n602 gnd 0.009526f
C1786 vdd.n603 gnd 0.009526f
C1787 vdd.n604 gnd 0.009526f
C1788 vdd.n605 gnd 0.006097f
C1789 vdd.n610 gnd 0.006478f
C1790 vdd.n611 gnd 0.006478f
C1791 vdd.n612 gnd 0.006478f
C1792 vdd.n613 gnd 8.304331f
C1793 vdd.n614 gnd 0.006478f
C1794 vdd.n615 gnd 0.006478f
C1795 vdd.n616 gnd 0.006478f
C1796 vdd.n618 gnd 0.006478f
C1797 vdd.n619 gnd 0.006478f
C1798 vdd.n621 gnd 0.006478f
C1799 vdd.n622 gnd 0.004716f
C1800 vdd.n624 gnd 0.006478f
C1801 vdd.t7 gnd 0.261771f
C1802 vdd.t6 gnd 0.267955f
C1803 vdd.t4 gnd 0.170894f
C1804 vdd.n625 gnd 0.092359f
C1805 vdd.n626 gnd 0.052389f
C1806 vdd.n627 gnd 0.009258f
C1807 vdd.n628 gnd 0.014994f
C1808 vdd.n630 gnd 0.006478f
C1809 vdd.n631 gnd 0.66201f
C1810 vdd.n632 gnd 0.01419f
C1811 vdd.n633 gnd 0.01419f
C1812 vdd.n634 gnd 0.006478f
C1813 vdd.n635 gnd 0.015151f
C1814 vdd.n636 gnd 0.006478f
C1815 vdd.n637 gnd 0.006478f
C1816 vdd.n638 gnd 0.006478f
C1817 vdd.n639 gnd 0.006478f
C1818 vdd.n640 gnd 0.006478f
C1819 vdd.n642 gnd 0.006478f
C1820 vdd.n643 gnd 0.006478f
C1821 vdd.n645 gnd 0.006478f
C1822 vdd.n646 gnd 0.006478f
C1823 vdd.n648 gnd 0.006478f
C1824 vdd.n649 gnd 0.006478f
C1825 vdd.n651 gnd 0.006478f
C1826 vdd.n652 gnd 0.006478f
C1827 vdd.n654 gnd 0.006478f
C1828 vdd.n655 gnd 0.006478f
C1829 vdd.n657 gnd 0.006478f
C1830 vdd.n658 gnd 0.004716f
C1831 vdd.n660 gnd 0.006478f
C1832 vdd.t76 gnd 0.261771f
C1833 vdd.t75 gnd 0.267955f
C1834 vdd.t74 gnd 0.170894f
C1835 vdd.n661 gnd 0.092359f
C1836 vdd.n662 gnd 0.052389f
C1837 vdd.n663 gnd 0.009258f
C1838 vdd.n664 gnd 0.006478f
C1839 vdd.n665 gnd 0.006478f
C1840 vdd.t5 gnd 0.331005f
C1841 vdd.n666 gnd 0.006478f
C1842 vdd.n667 gnd 0.006478f
C1843 vdd.n668 gnd 0.006478f
C1844 vdd.n669 gnd 0.006478f
C1845 vdd.n670 gnd 0.006478f
C1846 vdd.n671 gnd 0.66201f
C1847 vdd.n672 gnd 0.006478f
C1848 vdd.n673 gnd 0.006478f
C1849 vdd.n674 gnd 0.559788f
C1850 vdd.n675 gnd 0.006478f
C1851 vdd.n676 gnd 0.006478f
C1852 vdd.n677 gnd 0.006478f
C1853 vdd.n678 gnd 0.006478f
C1854 vdd.n679 gnd 0.647407f
C1855 vdd.n680 gnd 0.006478f
C1856 vdd.n681 gnd 0.006478f
C1857 vdd.n682 gnd 0.006478f
C1858 vdd.n683 gnd 0.006478f
C1859 vdd.n684 gnd 0.006478f
C1860 vdd.n685 gnd 0.66201f
C1861 vdd.n686 gnd 0.006478f
C1862 vdd.n687 gnd 0.006478f
C1863 vdd.t132 gnd 0.331005f
C1864 vdd.n688 gnd 0.006478f
C1865 vdd.n689 gnd 0.006478f
C1866 vdd.n690 gnd 0.006478f
C1867 vdd.t101 gnd 0.331005f
C1868 vdd.n691 gnd 0.006478f
C1869 vdd.n692 gnd 0.006478f
C1870 vdd.n693 gnd 0.006478f
C1871 vdd.n694 gnd 0.006478f
C1872 vdd.n695 gnd 0.006478f
C1873 vdd.t38 gnd 0.27746f
C1874 vdd.n696 gnd 0.006478f
C1875 vdd.n697 gnd 0.006478f
C1876 vdd.n698 gnd 0.530581f
C1877 vdd.n699 gnd 0.006478f
C1878 vdd.t39 gnd 0.267955f
C1879 vdd.t37 gnd 0.170894f
C1880 vdd.t40 gnd 0.267955f
C1881 vdd.n700 gnd 0.150602f
C1882 vdd.n701 gnd 0.006478f
C1883 vdd.n702 gnd 0.006478f
C1884 vdd.n703 gnd 0.423492f
C1885 vdd.n704 gnd 0.006478f
C1886 vdd.n705 gnd 0.006478f
C1887 vdd.t2 gnd 0.097354f
C1888 vdd.n706 gnd 0.38455f
C1889 vdd.n707 gnd 0.006478f
C1890 vdd.n708 gnd 0.006478f
C1891 vdd.n709 gnd 0.006478f
C1892 vdd.n710 gnd 0.569523f
C1893 vdd.n711 gnd 0.006478f
C1894 vdd.n712 gnd 0.006478f
C1895 vdd.t104 gnd 0.331005f
C1896 vdd.n713 gnd 0.006478f
C1897 vdd.n714 gnd 0.006478f
C1898 vdd.n715 gnd 0.006478f
C1899 vdd.t232 gnd 0.331005f
C1900 vdd.n716 gnd 0.006478f
C1901 vdd.n717 gnd 0.006478f
C1902 vdd.t1 gnd 0.331005f
C1903 vdd.n718 gnd 0.006478f
C1904 vdd.n719 gnd 0.006478f
C1905 vdd.n720 gnd 0.006478f
C1906 vdd.t80 gnd 0.262857f
C1907 vdd.n721 gnd 0.006478f
C1908 vdd.n722 gnd 0.006478f
C1909 vdd.n723 gnd 0.545185f
C1910 vdd.n724 gnd 0.006478f
C1911 vdd.n725 gnd 0.006478f
C1912 vdd.n726 gnd 0.006478f
C1913 vdd.t109 gnd 0.331005f
C1914 vdd.n727 gnd 0.006478f
C1915 vdd.n728 gnd 0.006478f
C1916 vdd.t106 gnd 0.27746f
C1917 vdd.n729 gnd 0.399153f
C1918 vdd.n730 gnd 0.006478f
C1919 vdd.n731 gnd 0.006478f
C1920 vdd.n732 gnd 0.006478f
C1921 vdd.n733 gnd 0.345608f
C1922 vdd.n734 gnd 0.006478f
C1923 vdd.n735 gnd 0.006478f
C1924 vdd.t116 gnd 0.331005f
C1925 vdd.n736 gnd 0.006478f
C1926 vdd.n737 gnd 0.006478f
C1927 vdd.n738 gnd 0.006478f
C1928 vdd.n739 gnd 0.66201f
C1929 vdd.n740 gnd 0.006478f
C1930 vdd.n741 gnd 0.006478f
C1931 vdd.t3 gnd 0.223915f
C1932 vdd.t122 gnd 0.316402f
C1933 vdd.n742 gnd 0.006478f
C1934 vdd.n743 gnd 0.006478f
C1935 vdd.n744 gnd 0.006478f
C1936 vdd.n745 gnd 0.496507f
C1937 vdd.n746 gnd 0.006478f
C1938 vdd.n747 gnd 0.006478f
C1939 vdd.n748 gnd 0.006478f
C1940 vdd.n749 gnd 0.006478f
C1941 vdd.n750 gnd 0.006478f
C1942 vdd.t55 gnd 0.331005f
C1943 vdd.n751 gnd 0.006478f
C1944 vdd.n752 gnd 0.006478f
C1945 vdd.t102 gnd 0.331005f
C1946 vdd.n753 gnd 0.006478f
C1947 vdd.n754 gnd 0.01419f
C1948 vdd.n755 gnd 0.01419f
C1949 vdd.n756 gnd 0.78857f
C1950 vdd.n757 gnd 0.006478f
C1951 vdd.n758 gnd 0.006478f
C1952 vdd.t126 gnd 0.331005f
C1953 vdd.n759 gnd 0.01419f
C1954 vdd.n760 gnd 0.006478f
C1955 vdd.n761 gnd 0.006478f
C1956 vdd.t99 gnd 0.603597f
C1957 vdd.n779 gnd 0.015151f
C1958 vdd.n797 gnd 0.01419f
C1959 vdd.n798 gnd 0.006478f
C1960 vdd.n799 gnd 0.01419f
C1961 vdd.t70 gnd 0.261771f
C1962 vdd.t69 gnd 0.267955f
C1963 vdd.t68 gnd 0.170894f
C1964 vdd.n800 gnd 0.092359f
C1965 vdd.n801 gnd 0.052389f
C1966 vdd.n802 gnd 0.014994f
C1967 vdd.n803 gnd 0.006478f
C1968 vdd.n804 gnd 0.350476f
C1969 vdd.n805 gnd 0.01419f
C1970 vdd.n806 gnd 0.006478f
C1971 vdd.n807 gnd 0.015151f
C1972 vdd.n808 gnd 0.006478f
C1973 vdd.t53 gnd 0.261771f
C1974 vdd.t52 gnd 0.267955f
C1975 vdd.t50 gnd 0.170894f
C1976 vdd.n809 gnd 0.092359f
C1977 vdd.n810 gnd 0.052389f
C1978 vdd.n811 gnd 0.009258f
C1979 vdd.n812 gnd 0.006478f
C1980 vdd.n813 gnd 0.006478f
C1981 vdd.t51 gnd 0.331005f
C1982 vdd.n814 gnd 0.006478f
C1983 vdd.t97 gnd 0.331005f
C1984 vdd.n815 gnd 0.006478f
C1985 vdd.n816 gnd 0.006478f
C1986 vdd.n817 gnd 0.006478f
C1987 vdd.n818 gnd 0.006478f
C1988 vdd.n819 gnd 0.006478f
C1989 vdd.n820 gnd 0.66201f
C1990 vdd.n821 gnd 0.006478f
C1991 vdd.n822 gnd 0.006478f
C1992 vdd.t230 gnd 0.331005f
C1993 vdd.n823 gnd 0.006478f
C1994 vdd.n824 gnd 0.006478f
C1995 vdd.n825 gnd 0.006478f
C1996 vdd.n826 gnd 0.006478f
C1997 vdd.n827 gnd 0.438095f
C1998 vdd.n828 gnd 0.006478f
C1999 vdd.n829 gnd 0.006478f
C2000 vdd.n830 gnd 0.006478f
C2001 vdd.n831 gnd 0.006478f
C2002 vdd.n832 gnd 0.006478f
C2003 vdd.n833 gnd 0.584126f
C2004 vdd.n834 gnd 0.006478f
C2005 vdd.n835 gnd 0.006478f
C2006 vdd.t124 gnd 0.316402f
C2007 vdd.t128 gnd 0.223915f
C2008 vdd.n836 gnd 0.006478f
C2009 vdd.n837 gnd 0.006478f
C2010 vdd.n838 gnd 0.006478f
C2011 vdd.t133 gnd 0.331005f
C2012 vdd.n839 gnd 0.006478f
C2013 vdd.n840 gnd 0.006478f
C2014 vdd.t110 gnd 0.331005f
C2015 vdd.n841 gnd 0.006478f
C2016 vdd.n842 gnd 0.006478f
C2017 vdd.n843 gnd 0.006478f
C2018 vdd.t234 gnd 0.27746f
C2019 vdd.n844 gnd 0.006478f
C2020 vdd.n845 gnd 0.006478f
C2021 vdd.n846 gnd 0.530581f
C2022 vdd.n847 gnd 0.006478f
C2023 vdd.n848 gnd 0.006478f
C2024 vdd.n849 gnd 0.006478f
C2025 vdd.t118 gnd 0.331005f
C2026 vdd.n850 gnd 0.006478f
C2027 vdd.n851 gnd 0.006478f
C2028 vdd.t131 gnd 0.262857f
C2029 vdd.n852 gnd 0.38455f
C2030 vdd.n853 gnd 0.006478f
C2031 vdd.n854 gnd 0.006478f
C2032 vdd.n855 gnd 0.006478f
C2033 vdd.n856 gnd 0.569523f
C2034 vdd.n857 gnd 0.006478f
C2035 vdd.n858 gnd 0.006478f
C2036 vdd.t108 gnd 0.331005f
C2037 vdd.n859 gnd 0.006478f
C2038 vdd.n860 gnd 0.006478f
C2039 vdd.n861 gnd 0.006478f
C2040 vdd.n862 gnd 0.66201f
C2041 vdd.n863 gnd 0.006478f
C2042 vdd.n864 gnd 0.006478f
C2043 vdd.t113 gnd 0.331005f
C2044 vdd.n865 gnd 0.006478f
C2045 vdd.n866 gnd 0.006478f
C2046 vdd.n867 gnd 0.006478f
C2047 vdd.t105 gnd 0.097354f
C2048 vdd.n868 gnd 0.006478f
C2049 vdd.n869 gnd 0.006478f
C2050 vdd.n870 gnd 0.006478f
C2051 vdd.t60 gnd 0.267955f
C2052 vdd.t58 gnd 0.170894f
C2053 vdd.t61 gnd 0.267955f
C2054 vdd.n871 gnd 0.150602f
C2055 vdd.n872 gnd 0.006478f
C2056 vdd.n873 gnd 0.006478f
C2057 vdd.t0 gnd 0.331005f
C2058 vdd.n874 gnd 0.006478f
C2059 vdd.n875 gnd 0.006478f
C2060 vdd.t59 gnd 0.27746f
C2061 vdd.n876 gnd 0.564655f
C2062 vdd.n877 gnd 0.006478f
C2063 vdd.n878 gnd 0.006478f
C2064 vdd.n879 gnd 0.006478f
C2065 vdd.n880 gnd 0.345608f
C2066 vdd.n881 gnd 0.006478f
C2067 vdd.n882 gnd 0.006478f
C2068 vdd.n883 gnd 0.462433f
C2069 vdd.n884 gnd 0.006478f
C2070 vdd.n885 gnd 0.006478f
C2071 vdd.n886 gnd 0.006478f
C2072 vdd.n887 gnd 0.66201f
C2073 vdd.n888 gnd 0.006478f
C2074 vdd.n889 gnd 0.006478f
C2075 vdd.t112 gnd 0.331005f
C2076 vdd.n890 gnd 0.006478f
C2077 vdd.n891 gnd 0.006478f
C2078 vdd.n892 gnd 0.006478f
C2079 vdd.n893 gnd 0.66201f
C2080 vdd.n894 gnd 0.006478f
C2081 vdd.n895 gnd 0.006478f
C2082 vdd.n896 gnd 0.006478f
C2083 vdd.n897 gnd 0.006478f
C2084 vdd.n898 gnd 0.006478f
C2085 vdd.t9 gnd 0.331005f
C2086 vdd.n899 gnd 0.006478f
C2087 vdd.n900 gnd 0.006478f
C2088 vdd.n901 gnd 0.006478f
C2089 vdd.n902 gnd 0.01419f
C2090 vdd.n903 gnd 0.01419f
C2091 vdd.n904 gnd 0.934602f
C2092 vdd.n905 gnd 0.006478f
C2093 vdd.n906 gnd 0.006478f
C2094 vdd.n907 gnd 0.433227f
C2095 vdd.n908 gnd 0.01419f
C2096 vdd.n909 gnd 0.006478f
C2097 vdd.n910 gnd 0.006478f
C2098 vdd.n911 gnd 8.58666f
C2099 vdd.n944 gnd 0.015151f
C2100 vdd.n945 gnd 0.006478f
C2101 vdd.n946 gnd 0.006478f
C2102 vdd.n947 gnd 0.006478f
C2103 vdd.n948 gnd 0.006097f
C2104 vdd.n951 gnd 0.0228f
C2105 vdd.n952 gnd 0.006364f
C2106 vdd.n953 gnd 0.007668f
C2107 vdd.n955 gnd 0.009526f
C2108 vdd.n956 gnd 0.009526f
C2109 vdd.n957 gnd 0.007668f
C2110 vdd.n959 gnd 0.009526f
C2111 vdd.n960 gnd 0.009526f
C2112 vdd.n961 gnd 0.009526f
C2113 vdd.n962 gnd 0.009526f
C2114 vdd.n963 gnd 0.009526f
C2115 vdd.n964 gnd 0.007668f
C2116 vdd.n966 gnd 0.009526f
C2117 vdd.n967 gnd 0.009526f
C2118 vdd.n968 gnd 0.009526f
C2119 vdd.n969 gnd 0.009526f
C2120 vdd.n970 gnd 0.009526f
C2121 vdd.n971 gnd 0.007668f
C2122 vdd.n973 gnd 0.009526f
C2123 vdd.n974 gnd 0.009526f
C2124 vdd.n975 gnd 0.009526f
C2125 vdd.n976 gnd 0.009526f
C2126 vdd.n977 gnd 0.006402f
C2127 vdd.t64 gnd 0.117199f
C2128 vdd.t63 gnd 0.125253f
C2129 vdd.t62 gnd 0.15306f
C2130 vdd.n978 gnd 0.196201f
C2131 vdd.n979 gnd 0.164844f
C2132 vdd.n981 gnd 0.009526f
C2133 vdd.n982 gnd 0.009526f
C2134 vdd.n983 gnd 0.007668f
C2135 vdd.n984 gnd 0.009526f
C2136 vdd.n986 gnd 0.009526f
C2137 vdd.n987 gnd 0.009526f
C2138 vdd.n988 gnd 0.009526f
C2139 vdd.n989 gnd 0.009526f
C2140 vdd.n990 gnd 0.007668f
C2141 vdd.n992 gnd 0.009526f
C2142 vdd.n993 gnd 0.009526f
C2143 vdd.n994 gnd 0.009526f
C2144 vdd.n995 gnd 0.009526f
C2145 vdd.n996 gnd 0.009526f
C2146 vdd.n997 gnd 0.007668f
C2147 vdd.n999 gnd 0.009526f
C2148 vdd.n1000 gnd 0.009526f
C2149 vdd.n1001 gnd 0.009526f
C2150 vdd.n1002 gnd 0.009526f
C2151 vdd.n1003 gnd 0.009526f
C2152 vdd.n1004 gnd 0.007668f
C2153 vdd.n1006 gnd 0.009526f
C2154 vdd.n1007 gnd 0.009526f
C2155 vdd.n1008 gnd 0.009526f
C2156 vdd.n1009 gnd 0.009526f
C2157 vdd.n1010 gnd 0.009526f
C2158 vdd.n1011 gnd 0.007668f
C2159 vdd.n1013 gnd 0.009526f
C2160 vdd.n1014 gnd 0.009526f
C2161 vdd.n1015 gnd 0.009526f
C2162 vdd.n1016 gnd 0.009526f
C2163 vdd.n1017 gnd 0.007591f
C2164 vdd.t49 gnd 0.117199f
C2165 vdd.t48 gnd 0.125253f
C2166 vdd.t47 gnd 0.15306f
C2167 vdd.n1018 gnd 0.196201f
C2168 vdd.n1019 gnd 0.164844f
C2169 vdd.n1021 gnd 0.009526f
C2170 vdd.n1022 gnd 0.009526f
C2171 vdd.n1023 gnd 0.007668f
C2172 vdd.n1024 gnd 0.009526f
C2173 vdd.n1026 gnd 0.009526f
C2174 vdd.n1027 gnd 0.009526f
C2175 vdd.n1028 gnd 0.009526f
C2176 vdd.n1029 gnd 0.009526f
C2177 vdd.n1030 gnd 0.007668f
C2178 vdd.n1032 gnd 0.009526f
C2179 vdd.n1033 gnd 0.009526f
C2180 vdd.n1034 gnd 0.009526f
C2181 vdd.n1035 gnd 0.009526f
C2182 vdd.n1036 gnd 0.009526f
C2183 vdd.n1037 gnd 0.007668f
C2184 vdd.n1039 gnd 0.009526f
C2185 vdd.n1040 gnd 0.009526f
C2186 vdd.n1041 gnd 0.009526f
C2187 vdd.n1042 gnd 0.009526f
C2188 vdd.n1043 gnd 0.009526f
C2189 vdd.n1044 gnd 0.007668f
C2190 vdd.n1046 gnd 0.009526f
C2191 vdd.n1047 gnd 0.009526f
C2192 vdd.n1048 gnd 0.006097f
C2193 vdd.n1049 gnd 0.007668f
C2194 vdd.n1050 gnd 0.006478f
C2195 vdd.n1051 gnd 0.006478f
C2196 vdd.n1052 gnd 0.006478f
C2197 vdd.n1053 gnd 0.006478f
C2198 vdd.n1054 gnd 0.006478f
C2199 vdd.n1055 gnd 0.006478f
C2200 vdd.n1056 gnd 0.006478f
C2201 vdd.n1057 gnd 0.006478f
C2202 vdd.n1058 gnd 0.006478f
C2203 vdd.n1059 gnd 0.006478f
C2204 vdd.n1060 gnd 0.006478f
C2205 vdd.n1061 gnd 0.006478f
C2206 vdd.n1062 gnd 0.006478f
C2207 vdd.n1063 gnd 0.006478f
C2208 vdd.n1064 gnd 0.006478f
C2209 vdd.n1065 gnd 0.006478f
C2210 vdd.n1066 gnd 0.006478f
C2211 vdd.n1067 gnd 0.006478f
C2212 vdd.n1068 gnd 0.006478f
C2213 vdd.n1069 gnd 0.006478f
C2214 vdd.n1070 gnd 0.006478f
C2215 vdd.n1071 gnd 0.006478f
C2216 vdd.n1072 gnd 0.006478f
C2217 vdd.n1073 gnd 0.006478f
C2218 vdd.n1074 gnd 0.006478f
C2219 vdd.n1075 gnd 0.006478f
C2220 vdd.n1076 gnd 0.006478f
C2221 vdd.n1077 gnd 0.006478f
C2222 vdd.n1078 gnd 0.006478f
C2223 vdd.n1079 gnd 0.006478f
C2224 vdd.n1080 gnd 0.006478f
C2225 vdd.t10 gnd 0.261771f
C2226 vdd.t11 gnd 0.267955f
C2227 vdd.t8 gnd 0.170894f
C2228 vdd.n1081 gnd 0.092359f
C2229 vdd.n1082 gnd 0.052389f
C2230 vdd.n1083 gnd 0.009258f
C2231 vdd.n1084 gnd 0.006478f
C2232 vdd.n1085 gnd 0.006478f
C2233 vdd.n1086 gnd 0.006478f
C2234 vdd.n1087 gnd 0.006478f
C2235 vdd.n1088 gnd 0.006478f
C2236 vdd.n1089 gnd 0.006478f
C2237 vdd.n1090 gnd 0.006478f
C2238 vdd.n1091 gnd 0.006478f
C2239 vdd.n1092 gnd 0.006478f
C2240 vdd.n1093 gnd 0.006478f
C2241 vdd.n1094 gnd 0.006478f
C2242 vdd.n1095 gnd 0.006478f
C2243 vdd.n1096 gnd 0.006478f
C2244 vdd.n1097 gnd 0.006478f
C2245 vdd.n1098 gnd 0.006478f
C2246 vdd.n1099 gnd 0.006478f
C2247 vdd.n1100 gnd 0.006478f
C2248 vdd.t35 gnd 0.261771f
C2249 vdd.t36 gnd 0.267955f
C2250 vdd.t34 gnd 0.170894f
C2251 vdd.n1101 gnd 0.092359f
C2252 vdd.n1102 gnd 0.052389f
C2253 vdd.n1103 gnd 0.006478f
C2254 vdd.n1104 gnd 0.006478f
C2255 vdd.n1105 gnd 0.006478f
C2256 vdd.n1106 gnd 0.006478f
C2257 vdd.n1107 gnd 0.006478f
C2258 vdd.n1108 gnd 0.006478f
C2259 vdd.n1109 gnd 0.006478f
C2260 vdd.n1110 gnd 0.006478f
C2261 vdd.n1111 gnd 0.006478f
C2262 vdd.n1112 gnd 0.006478f
C2263 vdd.n1113 gnd 0.006478f
C2264 vdd.n1114 gnd 0.006478f
C2265 vdd.n1115 gnd 0.006478f
C2266 vdd.n1116 gnd 0.006478f
C2267 vdd.n1117 gnd 0.006478f
C2268 vdd.n1118 gnd 0.006478f
C2269 vdd.n1119 gnd 0.006478f
C2270 vdd.n1120 gnd 0.006478f
C2271 vdd.n1121 gnd 0.006478f
C2272 vdd.n1122 gnd 0.006478f
C2273 vdd.n1123 gnd 0.006478f
C2274 vdd.n1124 gnd 0.006478f
C2275 vdd.n1125 gnd 0.006478f
C2276 vdd.n1126 gnd 0.006478f
C2277 vdd.n1127 gnd 0.006478f
C2278 vdd.n1128 gnd 0.006478f
C2279 vdd.n1129 gnd 0.004716f
C2280 vdd.n1130 gnd 0.009258f
C2281 vdd.n1131 gnd 0.005001f
C2282 vdd.n1132 gnd 0.006478f
C2283 vdd.n1133 gnd 0.006478f
C2284 vdd.n1134 gnd 0.006478f
C2285 vdd.n1135 gnd 0.015151f
C2286 vdd.n1136 gnd 0.015151f
C2287 vdd.n1137 gnd 0.01419f
C2288 vdd.n1138 gnd 0.01419f
C2289 vdd.n1139 gnd 0.006478f
C2290 vdd.n1140 gnd 0.006478f
C2291 vdd.n1141 gnd 0.006478f
C2292 vdd.n1142 gnd 0.006478f
C2293 vdd.n1143 gnd 0.006478f
C2294 vdd.n1144 gnd 0.006478f
C2295 vdd.n1145 gnd 0.006478f
C2296 vdd.n1146 gnd 0.006478f
C2297 vdd.n1147 gnd 0.006478f
C2298 vdd.n1148 gnd 0.006478f
C2299 vdd.n1149 gnd 0.006478f
C2300 vdd.n1150 gnd 0.006478f
C2301 vdd.n1151 gnd 0.006478f
C2302 vdd.n1152 gnd 0.006478f
C2303 vdd.n1153 gnd 0.006478f
C2304 vdd.n1154 gnd 0.006478f
C2305 vdd.n1155 gnd 0.006478f
C2306 vdd.n1156 gnd 0.006478f
C2307 vdd.n1157 gnd 0.006478f
C2308 vdd.n1158 gnd 0.006478f
C2309 vdd.n1159 gnd 0.006478f
C2310 vdd.n1160 gnd 0.006478f
C2311 vdd.n1161 gnd 0.006478f
C2312 vdd.n1162 gnd 0.006478f
C2313 vdd.n1163 gnd 0.006478f
C2314 vdd.n1164 gnd 0.006478f
C2315 vdd.n1165 gnd 0.006478f
C2316 vdd.n1166 gnd 0.394285f
C2317 vdd.n1167 gnd 0.006478f
C2318 vdd.n1168 gnd 0.006478f
C2319 vdd.n1169 gnd 0.006478f
C2320 vdd.n1170 gnd 0.006478f
C2321 vdd.n1171 gnd 0.006478f
C2322 vdd.n1172 gnd 0.006478f
C2323 vdd.n1173 gnd 0.006478f
C2324 vdd.n1174 gnd 0.006478f
C2325 vdd.n1175 gnd 0.006478f
C2326 vdd.n1176 gnd 0.006478f
C2327 vdd.n1177 gnd 0.006478f
C2328 vdd.n1178 gnd 0.006478f
C2329 vdd.n1179 gnd 0.006478f
C2330 vdd.n1180 gnd 0.006478f
C2331 vdd.n1181 gnd 0.006478f
C2332 vdd.n1182 gnd 0.006478f
C2333 vdd.n1183 gnd 0.006478f
C2334 vdd.n1184 gnd 0.006478f
C2335 vdd.n1185 gnd 0.006478f
C2336 vdd.n1186 gnd 0.006478f
C2337 vdd.n1187 gnd 0.209312f
C2338 vdd.n1188 gnd 0.006478f
C2339 vdd.n1189 gnd 0.006478f
C2340 vdd.n1190 gnd 0.006478f
C2341 vdd.n1191 gnd 0.006478f
C2342 vdd.n1192 gnd 0.006478f
C2343 vdd.n1193 gnd 0.006478f
C2344 vdd.n1194 gnd 0.006478f
C2345 vdd.n1195 gnd 0.006478f
C2346 vdd.n1196 gnd 0.006478f
C2347 vdd.n1197 gnd 0.006478f
C2348 vdd.n1198 gnd 0.006478f
C2349 vdd.n1199 gnd 0.006478f
C2350 vdd.n1200 gnd 0.006478f
C2351 vdd.n1201 gnd 0.006478f
C2352 vdd.n1202 gnd 0.006478f
C2353 vdd.n1203 gnd 0.006478f
C2354 vdd.n1204 gnd 0.006478f
C2355 vdd.n1205 gnd 0.006478f
C2356 vdd.n1206 gnd 0.006478f
C2357 vdd.n1207 gnd 0.006478f
C2358 vdd.n1208 gnd 0.006478f
C2359 vdd.n1209 gnd 0.006478f
C2360 vdd.n1210 gnd 0.006478f
C2361 vdd.n1211 gnd 0.006478f
C2362 vdd.n1212 gnd 0.006478f
C2363 vdd.n1213 gnd 0.006478f
C2364 vdd.n1214 gnd 0.006478f
C2365 vdd.n1215 gnd 0.01419f
C2366 vdd.n1216 gnd 0.01419f
C2367 vdd.n1217 gnd 0.015151f
C2368 vdd.n1218 gnd 0.006478f
C2369 vdd.n1219 gnd 0.006478f
C2370 vdd.n1220 gnd 0.005001f
C2371 vdd.n1221 gnd 0.006478f
C2372 vdd.n1222 gnd 0.006478f
C2373 vdd.n1223 gnd 0.004716f
C2374 vdd.n1224 gnd 0.006478f
C2375 vdd.n1225 gnd 0.006478f
C2376 vdd.n1226 gnd 0.006478f
C2377 vdd.n1227 gnd 0.006478f
C2378 vdd.n1228 gnd 0.006478f
C2379 vdd.n1229 gnd 0.006478f
C2380 vdd.n1230 gnd 0.006478f
C2381 vdd.n1231 gnd 0.006478f
C2382 vdd.n1232 gnd 0.006478f
C2383 vdd.n1233 gnd 0.006478f
C2384 vdd.n1234 gnd 0.006478f
C2385 vdd.n1235 gnd 0.006478f
C2386 vdd.n1236 gnd 0.006478f
C2387 vdd.n1237 gnd 0.006478f
C2388 vdd.n1238 gnd 0.006478f
C2389 vdd.n1239 gnd 0.006478f
C2390 vdd.n1240 gnd 0.006478f
C2391 vdd.n1241 gnd 0.006478f
C2392 vdd.n1242 gnd 0.006478f
C2393 vdd.n1243 gnd 0.006478f
C2394 vdd.n1244 gnd 0.006478f
C2395 vdd.n1245 gnd 0.006478f
C2396 vdd.n1246 gnd 0.006478f
C2397 vdd.n1247 gnd 0.006478f
C2398 vdd.n1248 gnd 0.006478f
C2399 vdd.n1249 gnd 0.006478f
C2400 vdd.n1250 gnd 0.025963f
C2401 vdd.n1252 gnd 0.0228f
C2402 vdd.n1253 gnd 0.007668f
C2403 vdd.n1255 gnd 0.009526f
C2404 vdd.n1256 gnd 0.007668f
C2405 vdd.n1257 gnd 0.009526f
C2406 vdd.n1259 gnd 0.009526f
C2407 vdd.n1260 gnd 0.009526f
C2408 vdd.n1262 gnd 0.009526f
C2409 vdd.n1263 gnd 0.006364f
C2410 vdd.t17 gnd 0.486772f
C2411 vdd.n1264 gnd 0.009526f
C2412 vdd.n1265 gnd 0.0228f
C2413 vdd.n1266 gnd 0.007668f
C2414 vdd.n1267 gnd 0.009526f
C2415 vdd.n1268 gnd 0.007668f
C2416 vdd.n1269 gnd 0.009526f
C2417 vdd.n1270 gnd 0.973544f
C2418 vdd.n1271 gnd 0.009526f
C2419 vdd.n1272 gnd 0.007668f
C2420 vdd.n1273 gnd 0.007668f
C2421 vdd.n1274 gnd 0.009526f
C2422 vdd.n1275 gnd 0.007668f
C2423 vdd.n1276 gnd 0.009526f
C2424 vdd.t161 gnd 0.486772f
C2425 vdd.n1277 gnd 0.009526f
C2426 vdd.n1278 gnd 0.007668f
C2427 vdd.n1279 gnd 0.009526f
C2428 vdd.n1280 gnd 0.007668f
C2429 vdd.n1281 gnd 0.009526f
C2430 vdd.t136 gnd 0.486772f
C2431 vdd.n1282 gnd 0.009526f
C2432 vdd.n1283 gnd 0.007668f
C2433 vdd.n1284 gnd 0.009526f
C2434 vdd.n1285 gnd 0.007668f
C2435 vdd.n1286 gnd 0.009526f
C2436 vdd.t181 gnd 0.486772f
C2437 vdd.n1287 gnd 0.764232f
C2438 vdd.n1288 gnd 0.009526f
C2439 vdd.n1289 gnd 0.007668f
C2440 vdd.n1290 gnd 0.009526f
C2441 vdd.n1291 gnd 0.007668f
C2442 vdd.n1292 gnd 0.009526f
C2443 vdd.n1293 gnd 0.686348f
C2444 vdd.n1294 gnd 0.009526f
C2445 vdd.n1295 gnd 0.007668f
C2446 vdd.n1296 gnd 0.009526f
C2447 vdd.n1297 gnd 0.007668f
C2448 vdd.n1298 gnd 0.009526f
C2449 vdd.n1299 gnd 0.520846f
C2450 vdd.t195 gnd 0.486772f
C2451 vdd.n1300 gnd 0.009526f
C2452 vdd.n1301 gnd 0.007668f
C2453 vdd.n1302 gnd 0.009494f
C2454 vdd.n1303 gnd 0.007668f
C2455 vdd.n1304 gnd 0.009526f
C2456 vdd.t174 gnd 0.486772f
C2457 vdd.n1305 gnd 0.009526f
C2458 vdd.n1306 gnd 0.007668f
C2459 vdd.n1307 gnd 0.009526f
C2460 vdd.n1308 gnd 0.007668f
C2461 vdd.n1309 gnd 0.009526f
C2462 vdd.t148 gnd 0.486772f
C2463 vdd.n1310 gnd 0.6182f
C2464 vdd.n1311 gnd 0.009526f
C2465 vdd.n1312 gnd 0.007668f
C2466 vdd.n1313 gnd 0.009526f
C2467 vdd.n1314 gnd 0.007668f
C2468 vdd.n1315 gnd 0.009526f
C2469 vdd.t156 gnd 0.486772f
C2470 vdd.n1316 gnd 0.009526f
C2471 vdd.n1317 gnd 0.007668f
C2472 vdd.n1318 gnd 0.009526f
C2473 vdd.n1319 gnd 0.007668f
C2474 vdd.n1320 gnd 0.009526f
C2475 vdd.n1321 gnd 0.666878f
C2476 vdd.n1322 gnd 0.808041f
C2477 vdd.t190 gnd 0.486772f
C2478 vdd.n1323 gnd 0.009526f
C2479 vdd.n1324 gnd 0.007668f
C2480 vdd.n1325 gnd 0.009526f
C2481 vdd.n1326 gnd 0.007668f
C2482 vdd.n1327 gnd 0.009526f
C2483 vdd.n1328 gnd 0.501375f
C2484 vdd.n1329 gnd 0.009526f
C2485 vdd.n1330 gnd 0.007668f
C2486 vdd.n1331 gnd 0.009526f
C2487 vdd.n1332 gnd 0.007668f
C2488 vdd.n1333 gnd 0.009526f
C2489 vdd.n1334 gnd 0.973544f
C2490 vdd.t140 gnd 0.486772f
C2491 vdd.n1335 gnd 0.009526f
C2492 vdd.n1336 gnd 0.007668f
C2493 vdd.n1337 gnd 0.009526f
C2494 vdd.n1338 gnd 0.007668f
C2495 vdd.n1339 gnd 0.009526f
C2496 vdd.t25 gnd 0.486772f
C2497 vdd.n1340 gnd 0.009526f
C2498 vdd.n1341 gnd 0.007668f
C2499 vdd.n1342 gnd 0.0228f
C2500 vdd.n1343 gnd 0.0228f
C2501 vdd.n1344 gnd 2.23915f
C2502 vdd.n1345 gnd 0.550052f
C2503 vdd.n1346 gnd 0.0228f
C2504 vdd.n1347 gnd 0.009526f
C2505 vdd.n1349 gnd 0.009526f
C2506 vdd.n1350 gnd 0.009526f
C2507 vdd.n1351 gnd 0.007668f
C2508 vdd.n1352 gnd 0.009526f
C2509 vdd.n1353 gnd 0.009526f
C2510 vdd.n1355 gnd 0.009526f
C2511 vdd.n1356 gnd 0.009526f
C2512 vdd.n1358 gnd 0.009526f
C2513 vdd.n1359 gnd 0.007668f
C2514 vdd.n1360 gnd 0.009526f
C2515 vdd.n1361 gnd 0.009526f
C2516 vdd.n1363 gnd 0.009526f
C2517 vdd.n1364 gnd 0.009526f
C2518 vdd.n1366 gnd 0.009526f
C2519 vdd.n1367 gnd 0.007668f
C2520 vdd.n1368 gnd 0.009526f
C2521 vdd.n1369 gnd 0.009526f
C2522 vdd.n1371 gnd 0.009526f
C2523 vdd.n1372 gnd 0.009526f
C2524 vdd.n1374 gnd 0.009526f
C2525 vdd.n1375 gnd 0.007668f
C2526 vdd.n1376 gnd 0.009526f
C2527 vdd.n1377 gnd 0.009526f
C2528 vdd.n1379 gnd 0.009526f
C2529 vdd.n1380 gnd 0.009526f
C2530 vdd.n1382 gnd 0.009526f
C2531 vdd.t45 gnd 0.117199f
C2532 vdd.t46 gnd 0.125253f
C2533 vdd.t44 gnd 0.15306f
C2534 vdd.n1383 gnd 0.196201f
C2535 vdd.n1384 gnd 0.165611f
C2536 vdd.n1385 gnd 0.016409f
C2537 vdd.n1386 gnd 0.009526f
C2538 vdd.n1387 gnd 0.009526f
C2539 vdd.n1389 gnd 0.009526f
C2540 vdd.n1390 gnd 0.009526f
C2541 vdd.n1392 gnd 0.009526f
C2542 vdd.n1393 gnd 0.007668f
C2543 vdd.n1394 gnd 0.009526f
C2544 vdd.n1395 gnd 0.009526f
C2545 vdd.n1397 gnd 0.009526f
C2546 vdd.n1398 gnd 0.009526f
C2547 vdd.n1400 gnd 0.009526f
C2548 vdd.n1401 gnd 0.007668f
C2549 vdd.n1402 gnd 0.009526f
C2550 vdd.n1403 gnd 0.009526f
C2551 vdd.n1405 gnd 0.009526f
C2552 vdd.n1406 gnd 0.009526f
C2553 vdd.n1408 gnd 0.009526f
C2554 vdd.n1409 gnd 0.007668f
C2555 vdd.n1410 gnd 0.009526f
C2556 vdd.n1411 gnd 0.009526f
C2557 vdd.n1413 gnd 0.009526f
C2558 vdd.n1414 gnd 0.009526f
C2559 vdd.n1416 gnd 0.009526f
C2560 vdd.n1417 gnd 0.007668f
C2561 vdd.n1418 gnd 0.009526f
C2562 vdd.n1419 gnd 0.009526f
C2563 vdd.n1421 gnd 0.009526f
C2564 vdd.n1422 gnd 0.009526f
C2565 vdd.n1424 gnd 0.009526f
C2566 vdd.n1425 gnd 0.007668f
C2567 vdd.n1426 gnd 0.009526f
C2568 vdd.n1427 gnd 0.009526f
C2569 vdd.n1429 gnd 0.009526f
C2570 vdd.n1430 gnd 0.007591f
C2571 vdd.n1432 gnd 0.007668f
C2572 vdd.n1433 gnd 0.009526f
C2573 vdd.n1434 gnd 0.009526f
C2574 vdd.n1435 gnd 0.009526f
C2575 vdd.n1436 gnd 0.009526f
C2576 vdd.n1438 gnd 0.009526f
C2577 vdd.n1439 gnd 0.009526f
C2578 vdd.n1440 gnd 0.007668f
C2579 vdd.n1441 gnd 0.009526f
C2580 vdd.n1443 gnd 0.009526f
C2581 vdd.n1444 gnd 0.009526f
C2582 vdd.n1446 gnd 0.009526f
C2583 vdd.n1447 gnd 0.009526f
C2584 vdd.n1448 gnd 0.007668f
C2585 vdd.n1449 gnd 0.009526f
C2586 vdd.n1451 gnd 0.009526f
C2587 vdd.n1452 gnd 0.009526f
C2588 vdd.n1454 gnd 0.009526f
C2589 vdd.n1455 gnd 0.009526f
C2590 vdd.n1456 gnd 0.007668f
C2591 vdd.n1457 gnd 0.009526f
C2592 vdd.n1459 gnd 0.009526f
C2593 vdd.n1460 gnd 0.009526f
C2594 vdd.n1462 gnd 0.009526f
C2595 vdd.n1463 gnd 0.009526f
C2596 vdd.n1464 gnd 0.007668f
C2597 vdd.n1465 gnd 0.009526f
C2598 vdd.n1467 gnd 0.009526f
C2599 vdd.n1468 gnd 0.009526f
C2600 vdd.n1470 gnd 0.009526f
C2601 vdd.n1471 gnd 0.003642f
C2602 vdd.t26 gnd 0.117199f
C2603 vdd.t27 gnd 0.125253f
C2604 vdd.t24 gnd 0.15306f
C2605 vdd.n1472 gnd 0.196201f
C2606 vdd.n1473 gnd 0.165611f
C2607 vdd.n1474 gnd 0.012575f
C2608 vdd.n1475 gnd 0.004025f
C2609 vdd.n1476 gnd 0.007668f
C2610 vdd.n1477 gnd 0.009526f
C2611 vdd.n1478 gnd 0.009526f
C2612 vdd.n1479 gnd 0.009526f
C2613 vdd.n1480 gnd 0.007668f
C2614 vdd.n1481 gnd 0.007668f
C2615 vdd.n1482 gnd 0.007668f
C2616 vdd.n1483 gnd 0.009526f
C2617 vdd.n1484 gnd 0.009526f
C2618 vdd.n1485 gnd 0.009526f
C2619 vdd.n1486 gnd 0.007668f
C2620 vdd.n1487 gnd 0.007668f
C2621 vdd.n1488 gnd 0.007668f
C2622 vdd.n1489 gnd 0.009526f
C2623 vdd.n1490 gnd 0.009526f
C2624 vdd.n1491 gnd 0.009526f
C2625 vdd.n1492 gnd 0.007668f
C2626 vdd.n1493 gnd 0.007668f
C2627 vdd.n1494 gnd 0.007668f
C2628 vdd.n1495 gnd 0.009526f
C2629 vdd.n1496 gnd 0.009526f
C2630 vdd.n1497 gnd 0.009526f
C2631 vdd.n1498 gnd 0.007668f
C2632 vdd.n1499 gnd 0.007668f
C2633 vdd.n1500 gnd 0.007668f
C2634 vdd.n1501 gnd 0.009526f
C2635 vdd.n1502 gnd 0.009526f
C2636 vdd.n1503 gnd 0.009526f
C2637 vdd.n1504 gnd 0.007668f
C2638 vdd.n1505 gnd 0.009526f
C2639 vdd.n1506 gnd 0.009526f
C2640 vdd.n1508 gnd 0.009526f
C2641 vdd.t32 gnd 0.117199f
C2642 vdd.t33 gnd 0.125253f
C2643 vdd.t31 gnd 0.15306f
C2644 vdd.n1509 gnd 0.196201f
C2645 vdd.n1510 gnd 0.165611f
C2646 vdd.n1511 gnd 0.016409f
C2647 vdd.n1512 gnd 0.005214f
C2648 vdd.n1513 gnd 0.009526f
C2649 vdd.n1514 gnd 0.009526f
C2650 vdd.n1515 gnd 0.009526f
C2651 vdd.n1516 gnd 0.007668f
C2652 vdd.n1517 gnd 0.007668f
C2653 vdd.n1518 gnd 0.007668f
C2654 vdd.n1519 gnd 0.009526f
C2655 vdd.n1520 gnd 0.009526f
C2656 vdd.n1521 gnd 0.009526f
C2657 vdd.n1522 gnd 0.007668f
C2658 vdd.n1523 gnd 0.007668f
C2659 vdd.n1524 gnd 0.007668f
C2660 vdd.n1525 gnd 0.009526f
C2661 vdd.n1526 gnd 0.009526f
C2662 vdd.n1527 gnd 0.009526f
C2663 vdd.n1528 gnd 0.007668f
C2664 vdd.n1529 gnd 0.007668f
C2665 vdd.n1530 gnd 0.007668f
C2666 vdd.n1531 gnd 0.009526f
C2667 vdd.n1532 gnd 0.009526f
C2668 vdd.n1533 gnd 0.009526f
C2669 vdd.n1534 gnd 0.007668f
C2670 vdd.n1535 gnd 0.007668f
C2671 vdd.n1536 gnd 0.007668f
C2672 vdd.n1537 gnd 0.009526f
C2673 vdd.n1538 gnd 0.009526f
C2674 vdd.n1539 gnd 0.009526f
C2675 vdd.n1540 gnd 0.007668f
C2676 vdd.n1541 gnd 0.007668f
C2677 vdd.n1542 gnd 0.006402f
C2678 vdd.n1543 gnd 0.009526f
C2679 vdd.n1544 gnd 0.009526f
C2680 vdd.n1545 gnd 0.009526f
C2681 vdd.n1546 gnd 0.006402f
C2682 vdd.n1547 gnd 0.007668f
C2683 vdd.n1548 gnd 0.007668f
C2684 vdd.n1549 gnd 0.009526f
C2685 vdd.n1550 gnd 0.009526f
C2686 vdd.n1551 gnd 0.009526f
C2687 vdd.n1552 gnd 0.007668f
C2688 vdd.n1553 gnd 0.007668f
C2689 vdd.n1554 gnd 0.007668f
C2690 vdd.n1555 gnd 0.009526f
C2691 vdd.n1556 gnd 0.009526f
C2692 vdd.n1557 gnd 0.009526f
C2693 vdd.n1558 gnd 0.007668f
C2694 vdd.n1559 gnd 0.007668f
C2695 vdd.n1560 gnd 0.007668f
C2696 vdd.n1561 gnd 0.009526f
C2697 vdd.n1562 gnd 0.009526f
C2698 vdd.n1563 gnd 0.009526f
C2699 vdd.n1564 gnd 0.007668f
C2700 vdd.n1565 gnd 0.007668f
C2701 vdd.n1566 gnd 0.007668f
C2702 vdd.n1567 gnd 0.009526f
C2703 vdd.n1568 gnd 0.009526f
C2704 vdd.n1569 gnd 0.009526f
C2705 vdd.n1570 gnd 0.007668f
C2706 vdd.n1571 gnd 0.007668f
C2707 vdd.n1572 gnd 0.006364f
C2708 vdd.n1573 gnd 0.0228f
C2709 vdd.n1574 gnd 0.02245f
C2710 vdd.n1575 gnd 0.006364f
C2711 vdd.n1576 gnd 0.02245f
C2712 vdd.n1577 gnd 1.3727f
C2713 vdd.n1578 gnd 0.02245f
C2714 vdd.n1579 gnd 0.006364f
C2715 vdd.n1580 gnd 0.02245f
C2716 vdd.n1581 gnd 0.009526f
C2717 vdd.n1582 gnd 0.009526f
C2718 vdd.n1583 gnd 0.007668f
C2719 vdd.n1584 gnd 0.009526f
C2720 vdd.n1585 gnd 0.910263f
C2721 vdd.n1586 gnd 0.009526f
C2722 vdd.n1587 gnd 0.007668f
C2723 vdd.n1588 gnd 0.009526f
C2724 vdd.n1589 gnd 0.009526f
C2725 vdd.n1590 gnd 0.009526f
C2726 vdd.n1591 gnd 0.007668f
C2727 vdd.n1592 gnd 0.009526f
C2728 vdd.n1593 gnd 0.958941f
C2729 vdd.n1594 gnd 0.009526f
C2730 vdd.n1595 gnd 0.007668f
C2731 vdd.n1596 gnd 0.009526f
C2732 vdd.n1597 gnd 0.009526f
C2733 vdd.n1598 gnd 0.009526f
C2734 vdd.n1599 gnd 0.007668f
C2735 vdd.n1600 gnd 0.009526f
C2736 vdd.t192 gnd 0.486772f
C2737 vdd.n1601 gnd 0.793438f
C2738 vdd.n1602 gnd 0.009526f
C2739 vdd.n1603 gnd 0.007668f
C2740 vdd.n1604 gnd 0.009526f
C2741 vdd.n1605 gnd 0.009526f
C2742 vdd.n1606 gnd 0.009526f
C2743 vdd.n1607 gnd 0.007668f
C2744 vdd.n1608 gnd 0.009526f
C2745 vdd.n1609 gnd 0.627936f
C2746 vdd.n1610 gnd 0.009526f
C2747 vdd.n1611 gnd 0.007668f
C2748 vdd.n1612 gnd 0.009526f
C2749 vdd.n1613 gnd 0.009526f
C2750 vdd.n1614 gnd 0.009526f
C2751 vdd.n1615 gnd 0.007668f
C2752 vdd.n1616 gnd 0.009526f
C2753 vdd.n1617 gnd 0.783703f
C2754 vdd.n1618 gnd 0.511111f
C2755 vdd.n1619 gnd 0.009526f
C2756 vdd.n1620 gnd 0.007668f
C2757 vdd.n1621 gnd 0.009526f
C2758 vdd.n1622 gnd 0.009526f
C2759 vdd.n1623 gnd 0.009526f
C2760 vdd.n1624 gnd 0.007668f
C2761 vdd.n1625 gnd 0.009526f
C2762 vdd.n1626 gnd 0.676613f
C2763 vdd.n1627 gnd 0.009526f
C2764 vdd.n1628 gnd 0.007668f
C2765 vdd.n1629 gnd 0.009526f
C2766 vdd.n1630 gnd 0.009526f
C2767 vdd.n1631 gnd 0.009526f
C2768 vdd.n1632 gnd 0.007668f
C2769 vdd.n1633 gnd 0.009526f
C2770 vdd.t142 gnd 0.486772f
C2771 vdd.n1634 gnd 0.808041f
C2772 vdd.n1635 gnd 0.009526f
C2773 vdd.n1636 gnd 0.007668f
C2774 vdd.n1637 gnd 0.005228f
C2775 vdd.n1638 gnd 0.004851f
C2776 vdd.n1639 gnd 0.002684f
C2777 vdd.n1640 gnd 0.006162f
C2778 vdd.n1641 gnd 0.002607f
C2779 vdd.n1642 gnd 0.00276f
C2780 vdd.n1643 gnd 0.004851f
C2781 vdd.n1644 gnd 0.002607f
C2782 vdd.n1645 gnd 0.006162f
C2783 vdd.n1646 gnd 0.00276f
C2784 vdd.n1647 gnd 0.004851f
C2785 vdd.n1648 gnd 0.002607f
C2786 vdd.n1649 gnd 0.004621f
C2787 vdd.n1650 gnd 0.004635f
C2788 vdd.t162 gnd 0.013238f
C2789 vdd.n1651 gnd 0.029455f
C2790 vdd.n1652 gnd 0.153291f
C2791 vdd.n1653 gnd 0.002607f
C2792 vdd.n1654 gnd 0.00276f
C2793 vdd.n1655 gnd 0.006162f
C2794 vdd.n1656 gnd 0.006162f
C2795 vdd.n1657 gnd 0.00276f
C2796 vdd.n1658 gnd 0.002607f
C2797 vdd.n1659 gnd 0.004851f
C2798 vdd.n1660 gnd 0.004851f
C2799 vdd.n1661 gnd 0.002607f
C2800 vdd.n1662 gnd 0.00276f
C2801 vdd.n1663 gnd 0.006162f
C2802 vdd.n1664 gnd 0.006162f
C2803 vdd.n1665 gnd 0.00276f
C2804 vdd.n1666 gnd 0.002607f
C2805 vdd.n1667 gnd 0.004851f
C2806 vdd.n1668 gnd 0.004851f
C2807 vdd.n1669 gnd 0.002607f
C2808 vdd.n1670 gnd 0.00276f
C2809 vdd.n1671 gnd 0.006162f
C2810 vdd.n1672 gnd 0.006162f
C2811 vdd.n1673 gnd 0.014568f
C2812 vdd.n1674 gnd 0.002684f
C2813 vdd.n1675 gnd 0.002607f
C2814 vdd.n1676 gnd 0.012539f
C2815 vdd.n1677 gnd 0.008754f
C2816 vdd.t182 gnd 0.03067f
C2817 vdd.t214 gnd 0.03067f
C2818 vdd.n1678 gnd 0.210786f
C2819 vdd.n1679 gnd 0.165751f
C2820 vdd.t196 gnd 0.03067f
C2821 vdd.t224 gnd 0.03067f
C2822 vdd.n1680 gnd 0.210786f
C2823 vdd.n1681 gnd 0.13376f
C2824 vdd.t175 gnd 0.03067f
C2825 vdd.t143 gnd 0.03067f
C2826 vdd.n1682 gnd 0.210786f
C2827 vdd.n1683 gnd 0.13376f
C2828 vdd.t189 gnd 0.03067f
C2829 vdd.t149 gnd 0.03067f
C2830 vdd.n1684 gnd 0.210786f
C2831 vdd.n1685 gnd 0.13376f
C2832 vdd.t217 gnd 0.03067f
C2833 vdd.t228 gnd 0.03067f
C2834 vdd.n1686 gnd 0.210786f
C2835 vdd.n1687 gnd 0.13376f
C2836 vdd.n1688 gnd 0.005228f
C2837 vdd.n1689 gnd 0.004851f
C2838 vdd.n1690 gnd 0.002684f
C2839 vdd.n1691 gnd 0.006162f
C2840 vdd.n1692 gnd 0.002607f
C2841 vdd.n1693 gnd 0.00276f
C2842 vdd.n1694 gnd 0.004851f
C2843 vdd.n1695 gnd 0.002607f
C2844 vdd.n1696 gnd 0.006162f
C2845 vdd.n1697 gnd 0.00276f
C2846 vdd.n1698 gnd 0.004851f
C2847 vdd.n1699 gnd 0.002607f
C2848 vdd.n1700 gnd 0.004621f
C2849 vdd.n1701 gnd 0.004635f
C2850 vdd.t153 gnd 0.013238f
C2851 vdd.n1702 gnd 0.029455f
C2852 vdd.n1703 gnd 0.153291f
C2853 vdd.n1704 gnd 0.002607f
C2854 vdd.n1705 gnd 0.00276f
C2855 vdd.n1706 gnd 0.006162f
C2856 vdd.n1707 gnd 0.006162f
C2857 vdd.n1708 gnd 0.00276f
C2858 vdd.n1709 gnd 0.002607f
C2859 vdd.n1710 gnd 0.004851f
C2860 vdd.n1711 gnd 0.004851f
C2861 vdd.n1712 gnd 0.002607f
C2862 vdd.n1713 gnd 0.00276f
C2863 vdd.n1714 gnd 0.006162f
C2864 vdd.n1715 gnd 0.006162f
C2865 vdd.n1716 gnd 0.00276f
C2866 vdd.n1717 gnd 0.002607f
C2867 vdd.n1718 gnd 0.004851f
C2868 vdd.n1719 gnd 0.004851f
C2869 vdd.n1720 gnd 0.002607f
C2870 vdd.n1721 gnd 0.00276f
C2871 vdd.n1722 gnd 0.006162f
C2872 vdd.n1723 gnd 0.006162f
C2873 vdd.n1724 gnd 0.014568f
C2874 vdd.n1725 gnd 0.002684f
C2875 vdd.n1726 gnd 0.002607f
C2876 vdd.n1727 gnd 0.012539f
C2877 vdd.n1728 gnd 0.00848f
C2878 vdd.n1729 gnd 0.099518f
C2879 vdd.n1730 gnd 0.005228f
C2880 vdd.n1731 gnd 0.004851f
C2881 vdd.n1732 gnd 0.002684f
C2882 vdd.n1733 gnd 0.006162f
C2883 vdd.n1734 gnd 0.002607f
C2884 vdd.n1735 gnd 0.00276f
C2885 vdd.n1736 gnd 0.004851f
C2886 vdd.n1737 gnd 0.002607f
C2887 vdd.n1738 gnd 0.006162f
C2888 vdd.n1739 gnd 0.00276f
C2889 vdd.n1740 gnd 0.004851f
C2890 vdd.n1741 gnd 0.002607f
C2891 vdd.n1742 gnd 0.004621f
C2892 vdd.n1743 gnd 0.004635f
C2893 vdd.t212 gnd 0.013238f
C2894 vdd.n1744 gnd 0.029455f
C2895 vdd.n1745 gnd 0.153291f
C2896 vdd.n1746 gnd 0.002607f
C2897 vdd.n1747 gnd 0.00276f
C2898 vdd.n1748 gnd 0.006162f
C2899 vdd.n1749 gnd 0.006162f
C2900 vdd.n1750 gnd 0.00276f
C2901 vdd.n1751 gnd 0.002607f
C2902 vdd.n1752 gnd 0.004851f
C2903 vdd.n1753 gnd 0.004851f
C2904 vdd.n1754 gnd 0.002607f
C2905 vdd.n1755 gnd 0.00276f
C2906 vdd.n1756 gnd 0.006162f
C2907 vdd.n1757 gnd 0.006162f
C2908 vdd.n1758 gnd 0.00276f
C2909 vdd.n1759 gnd 0.002607f
C2910 vdd.n1760 gnd 0.004851f
C2911 vdd.n1761 gnd 0.004851f
C2912 vdd.n1762 gnd 0.002607f
C2913 vdd.n1763 gnd 0.00276f
C2914 vdd.n1764 gnd 0.006162f
C2915 vdd.n1765 gnd 0.006162f
C2916 vdd.n1766 gnd 0.014568f
C2917 vdd.n1767 gnd 0.002684f
C2918 vdd.n1768 gnd 0.002607f
C2919 vdd.n1769 gnd 0.012539f
C2920 vdd.n1770 gnd 0.008754f
C2921 vdd.t184 gnd 0.03067f
C2922 vdd.t137 gnd 0.03067f
C2923 vdd.n1771 gnd 0.210786f
C2924 vdd.n1772 gnd 0.165751f
C2925 vdd.t222 gnd 0.03067f
C2926 vdd.t203 gnd 0.03067f
C2927 vdd.n1773 gnd 0.210786f
C2928 vdd.n1774 gnd 0.13376f
C2929 vdd.t200 gnd 0.03067f
C2930 vdd.t163 gnd 0.03067f
C2931 vdd.n1775 gnd 0.210786f
C2932 vdd.n1776 gnd 0.13376f
C2933 vdd.t157 gnd 0.03067f
C2934 vdd.t201 gnd 0.03067f
C2935 vdd.n1777 gnd 0.210786f
C2936 vdd.n1778 gnd 0.13376f
C2937 vdd.t193 gnd 0.03067f
C2938 vdd.t191 gnd 0.03067f
C2939 vdd.n1779 gnd 0.210786f
C2940 vdd.n1780 gnd 0.13376f
C2941 vdd.n1781 gnd 0.005228f
C2942 vdd.n1782 gnd 0.004851f
C2943 vdd.n1783 gnd 0.002684f
C2944 vdd.n1784 gnd 0.006162f
C2945 vdd.n1785 gnd 0.002607f
C2946 vdd.n1786 gnd 0.00276f
C2947 vdd.n1787 gnd 0.004851f
C2948 vdd.n1788 gnd 0.002607f
C2949 vdd.n1789 gnd 0.006162f
C2950 vdd.n1790 gnd 0.00276f
C2951 vdd.n1791 gnd 0.004851f
C2952 vdd.n1792 gnd 0.002607f
C2953 vdd.n1793 gnd 0.004621f
C2954 vdd.n1794 gnd 0.004635f
C2955 vdd.t141 gnd 0.013238f
C2956 vdd.n1795 gnd 0.029455f
C2957 vdd.n1796 gnd 0.153291f
C2958 vdd.n1797 gnd 0.002607f
C2959 vdd.n1798 gnd 0.00276f
C2960 vdd.n1799 gnd 0.006162f
C2961 vdd.n1800 gnd 0.006162f
C2962 vdd.n1801 gnd 0.00276f
C2963 vdd.n1802 gnd 0.002607f
C2964 vdd.n1803 gnd 0.004851f
C2965 vdd.n1804 gnd 0.004851f
C2966 vdd.n1805 gnd 0.002607f
C2967 vdd.n1806 gnd 0.00276f
C2968 vdd.n1807 gnd 0.006162f
C2969 vdd.n1808 gnd 0.006162f
C2970 vdd.n1809 gnd 0.00276f
C2971 vdd.n1810 gnd 0.002607f
C2972 vdd.n1811 gnd 0.004851f
C2973 vdd.n1812 gnd 0.004851f
C2974 vdd.n1813 gnd 0.002607f
C2975 vdd.n1814 gnd 0.00276f
C2976 vdd.n1815 gnd 0.006162f
C2977 vdd.n1816 gnd 0.006162f
C2978 vdd.n1817 gnd 0.014568f
C2979 vdd.n1818 gnd 0.002684f
C2980 vdd.n1819 gnd 0.002607f
C2981 vdd.n1820 gnd 0.012539f
C2982 vdd.n1821 gnd 0.00848f
C2983 vdd.n1822 gnd 0.059203f
C2984 vdd.n1823 gnd 0.213325f
C2985 vdd.n1824 gnd 0.005228f
C2986 vdd.n1825 gnd 0.004851f
C2987 vdd.n1826 gnd 0.002684f
C2988 vdd.n1827 gnd 0.006162f
C2989 vdd.n1828 gnd 0.002607f
C2990 vdd.n1829 gnd 0.00276f
C2991 vdd.n1830 gnd 0.004851f
C2992 vdd.n1831 gnd 0.002607f
C2993 vdd.n1832 gnd 0.006162f
C2994 vdd.n1833 gnd 0.00276f
C2995 vdd.n1834 gnd 0.004851f
C2996 vdd.n1835 gnd 0.002607f
C2997 vdd.n1836 gnd 0.004621f
C2998 vdd.n1837 gnd 0.004635f
C2999 vdd.t221 gnd 0.013238f
C3000 vdd.n1838 gnd 0.029455f
C3001 vdd.n1839 gnd 0.153291f
C3002 vdd.n1840 gnd 0.002607f
C3003 vdd.n1841 gnd 0.00276f
C3004 vdd.n1842 gnd 0.006162f
C3005 vdd.n1843 gnd 0.006162f
C3006 vdd.n1844 gnd 0.00276f
C3007 vdd.n1845 gnd 0.002607f
C3008 vdd.n1846 gnd 0.004851f
C3009 vdd.n1847 gnd 0.004851f
C3010 vdd.n1848 gnd 0.002607f
C3011 vdd.n1849 gnd 0.00276f
C3012 vdd.n1850 gnd 0.006162f
C3013 vdd.n1851 gnd 0.006162f
C3014 vdd.n1852 gnd 0.00276f
C3015 vdd.n1853 gnd 0.002607f
C3016 vdd.n1854 gnd 0.004851f
C3017 vdd.n1855 gnd 0.004851f
C3018 vdd.n1856 gnd 0.002607f
C3019 vdd.n1857 gnd 0.00276f
C3020 vdd.n1858 gnd 0.006162f
C3021 vdd.n1859 gnd 0.006162f
C3022 vdd.n1860 gnd 0.014568f
C3023 vdd.n1861 gnd 0.002684f
C3024 vdd.n1862 gnd 0.002607f
C3025 vdd.n1863 gnd 0.012539f
C3026 vdd.n1864 gnd 0.008754f
C3027 vdd.t194 gnd 0.03067f
C3028 vdd.t154 gnd 0.03067f
C3029 vdd.n1865 gnd 0.210786f
C3030 vdd.n1866 gnd 0.165751f
C3031 vdd.t229 gnd 0.03067f
C3032 vdd.t209 gnd 0.03067f
C3033 vdd.n1867 gnd 0.210786f
C3034 vdd.n1868 gnd 0.13376f
C3035 vdd.t207 gnd 0.03067f
C3036 vdd.t177 gnd 0.03067f
C3037 vdd.n1869 gnd 0.210786f
C3038 vdd.n1870 gnd 0.13376f
C3039 vdd.t176 gnd 0.03067f
C3040 vdd.t208 gnd 0.03067f
C3041 vdd.n1871 gnd 0.210786f
C3042 vdd.n1872 gnd 0.13376f
C3043 vdd.t199 gnd 0.03067f
C3044 vdd.t198 gnd 0.03067f
C3045 vdd.n1873 gnd 0.210786f
C3046 vdd.n1874 gnd 0.13376f
C3047 vdd.n1875 gnd 0.005228f
C3048 vdd.n1876 gnd 0.004851f
C3049 vdd.n1877 gnd 0.002684f
C3050 vdd.n1878 gnd 0.006162f
C3051 vdd.n1879 gnd 0.002607f
C3052 vdd.n1880 gnd 0.00276f
C3053 vdd.n1881 gnd 0.004851f
C3054 vdd.n1882 gnd 0.002607f
C3055 vdd.n1883 gnd 0.006162f
C3056 vdd.n1884 gnd 0.00276f
C3057 vdd.n1885 gnd 0.004851f
C3058 vdd.n1886 gnd 0.002607f
C3059 vdd.n1887 gnd 0.004621f
C3060 vdd.n1888 gnd 0.004635f
C3061 vdd.t155 gnd 0.013238f
C3062 vdd.n1889 gnd 0.029455f
C3063 vdd.n1890 gnd 0.153291f
C3064 vdd.n1891 gnd 0.002607f
C3065 vdd.n1892 gnd 0.00276f
C3066 vdd.n1893 gnd 0.006162f
C3067 vdd.n1894 gnd 0.006162f
C3068 vdd.n1895 gnd 0.00276f
C3069 vdd.n1896 gnd 0.002607f
C3070 vdd.n1897 gnd 0.004851f
C3071 vdd.n1898 gnd 0.004851f
C3072 vdd.n1899 gnd 0.002607f
C3073 vdd.n1900 gnd 0.00276f
C3074 vdd.n1901 gnd 0.006162f
C3075 vdd.n1902 gnd 0.006162f
C3076 vdd.n1903 gnd 0.00276f
C3077 vdd.n1904 gnd 0.002607f
C3078 vdd.n1905 gnd 0.004851f
C3079 vdd.n1906 gnd 0.004851f
C3080 vdd.n1907 gnd 0.002607f
C3081 vdd.n1908 gnd 0.00276f
C3082 vdd.n1909 gnd 0.006162f
C3083 vdd.n1910 gnd 0.006162f
C3084 vdd.n1911 gnd 0.014568f
C3085 vdd.n1912 gnd 0.002684f
C3086 vdd.n1913 gnd 0.002607f
C3087 vdd.n1914 gnd 0.012539f
C3088 vdd.n1915 gnd 0.00848f
C3089 vdd.n1916 gnd 0.059203f
C3090 vdd.n1917 gnd 0.234451f
C3091 vdd.n1918 gnd 2.22508f
C3092 vdd.n1919 gnd 0.56708f
C3093 vdd.n1920 gnd 0.009494f
C3094 vdd.n1921 gnd 0.009526f
C3095 vdd.n1922 gnd 0.007668f
C3096 vdd.n1923 gnd 0.009526f
C3097 vdd.n1924 gnd 0.773967f
C3098 vdd.n1925 gnd 0.009526f
C3099 vdd.n1926 gnd 0.007668f
C3100 vdd.n1927 gnd 0.009526f
C3101 vdd.n1928 gnd 0.009526f
C3102 vdd.n1929 gnd 0.009526f
C3103 vdd.n1930 gnd 0.007668f
C3104 vdd.n1931 gnd 0.009526f
C3105 vdd.n1932 gnd 0.808041f
C3106 vdd.t202 gnd 0.486772f
C3107 vdd.n1933 gnd 0.608465f
C3108 vdd.n1934 gnd 0.009526f
C3109 vdd.n1935 gnd 0.007668f
C3110 vdd.n1936 gnd 0.009526f
C3111 vdd.n1937 gnd 0.009526f
C3112 vdd.n1938 gnd 0.009526f
C3113 vdd.n1939 gnd 0.007668f
C3114 vdd.n1940 gnd 0.009526f
C3115 vdd.n1941 gnd 0.530581f
C3116 vdd.n1942 gnd 0.009526f
C3117 vdd.n1943 gnd 0.007668f
C3118 vdd.n1944 gnd 0.009526f
C3119 vdd.n1945 gnd 0.009526f
C3120 vdd.n1946 gnd 0.009526f
C3121 vdd.n1947 gnd 0.007668f
C3122 vdd.n1948 gnd 0.009526f
C3123 vdd.n1949 gnd 0.598729f
C3124 vdd.n1950 gnd 0.696084f
C3125 vdd.n1951 gnd 0.009526f
C3126 vdd.n1952 gnd 0.007668f
C3127 vdd.n1953 gnd 0.009526f
C3128 vdd.n1954 gnd 0.009526f
C3129 vdd.n1955 gnd 0.009526f
C3130 vdd.n1956 gnd 0.007668f
C3131 vdd.n1957 gnd 0.009526f
C3132 vdd.n1958 gnd 0.861586f
C3133 vdd.n1959 gnd 0.009526f
C3134 vdd.n1960 gnd 0.007668f
C3135 vdd.n1961 gnd 0.009526f
C3136 vdd.n1962 gnd 0.009526f
C3137 vdd.n1963 gnd 0.02245f
C3138 vdd.n1964 gnd 0.009526f
C3139 vdd.n1965 gnd 0.009526f
C3140 vdd.n1966 gnd 0.007668f
C3141 vdd.n1967 gnd 0.009526f
C3142 vdd.n1968 gnd 0.520846f
C3143 vdd.n1969 gnd 0.973544f
C3144 vdd.n1970 gnd 0.009526f
C3145 vdd.n1971 gnd 0.007668f
C3146 vdd.n1972 gnd 0.009526f
C3147 vdd.n1973 gnd 0.009526f
C3148 vdd.n1974 gnd 0.02245f
C3149 vdd.n1975 gnd 0.006364f
C3150 vdd.n1976 gnd 0.02245f
C3151 vdd.n1977 gnd 1.33862f
C3152 vdd.n1978 gnd 0.02245f
C3153 vdd.n1979 gnd 0.0228f
C3154 vdd.n1980 gnd 0.003642f
C3155 vdd.t19 gnd 0.117199f
C3156 vdd.t18 gnd 0.125253f
C3157 vdd.t16 gnd 0.15306f
C3158 vdd.n1981 gnd 0.196201f
C3159 vdd.n1982 gnd 0.164844f
C3160 vdd.n1983 gnd 0.011808f
C3161 vdd.n1984 gnd 0.004025f
C3162 vdd.n1985 gnd 0.008193f
C3163 vdd.n1986 gnd 0.720431f
C3164 vdd.n1988 gnd 0.007668f
C3165 vdd.n1989 gnd 0.007668f
C3166 vdd.n1990 gnd 0.009526f
C3167 vdd.n1992 gnd 0.009526f
C3168 vdd.n1993 gnd 0.009526f
C3169 vdd.n1994 gnd 0.007668f
C3170 vdd.n1995 gnd 0.007668f
C3171 vdd.n1996 gnd 0.007668f
C3172 vdd.n1997 gnd 0.009526f
C3173 vdd.n1999 gnd 0.009526f
C3174 vdd.n2000 gnd 0.009526f
C3175 vdd.n2001 gnd 0.007668f
C3176 vdd.n2002 gnd 0.007668f
C3177 vdd.n2003 gnd 0.007668f
C3178 vdd.n2004 gnd 0.009526f
C3179 vdd.n2006 gnd 0.009526f
C3180 vdd.n2007 gnd 0.009526f
C3181 vdd.n2008 gnd 0.007668f
C3182 vdd.n2009 gnd 0.007668f
C3183 vdd.n2010 gnd 0.007668f
C3184 vdd.n2011 gnd 0.009526f
C3185 vdd.n2013 gnd 0.009526f
C3186 vdd.n2014 gnd 0.009526f
C3187 vdd.n2015 gnd 0.007668f
C3188 vdd.n2016 gnd 0.009526f
C3189 vdd.n2017 gnd 0.009526f
C3190 vdd.n2018 gnd 0.009526f
C3191 vdd.n2019 gnd 0.015642f
C3192 vdd.n2020 gnd 0.005214f
C3193 vdd.n2021 gnd 0.007668f
C3194 vdd.n2022 gnd 0.009526f
C3195 vdd.n2024 gnd 0.009526f
C3196 vdd.n2025 gnd 0.009526f
C3197 vdd.n2026 gnd 0.007668f
C3198 vdd.n2027 gnd 0.007668f
C3199 vdd.n2028 gnd 0.007668f
C3200 vdd.n2029 gnd 0.009526f
C3201 vdd.n2031 gnd 0.009526f
C3202 vdd.n2032 gnd 0.009526f
C3203 vdd.n2033 gnd 0.007668f
C3204 vdd.n2034 gnd 0.007668f
C3205 vdd.n2035 gnd 0.007668f
C3206 vdd.n2036 gnd 0.009526f
C3207 vdd.n2038 gnd 0.009526f
C3208 vdd.n2039 gnd 0.009526f
C3209 vdd.n2040 gnd 0.007668f
C3210 vdd.n2041 gnd 0.007668f
C3211 vdd.n2042 gnd 0.007668f
C3212 vdd.n2043 gnd 0.009526f
C3213 vdd.n2045 gnd 0.009526f
C3214 vdd.n2046 gnd 0.009526f
C3215 vdd.n2047 gnd 0.007668f
C3216 vdd.n2048 gnd 0.007668f
C3217 vdd.n2049 gnd 0.007668f
C3218 vdd.n2050 gnd 0.009526f
C3219 vdd.n2052 gnd 0.009526f
C3220 vdd.n2053 gnd 0.009526f
C3221 vdd.n2054 gnd 0.007668f
C3222 vdd.n2055 gnd 0.009526f
C3223 vdd.n2056 gnd 0.009526f
C3224 vdd.n2057 gnd 0.009526f
C3225 vdd.n2058 gnd 0.015642f
C3226 vdd.n2059 gnd 0.006402f
C3227 vdd.n2060 gnd 0.007668f
C3228 vdd.n2061 gnd 0.009526f
C3229 vdd.n2063 gnd 0.009526f
C3230 vdd.n2064 gnd 0.009526f
C3231 vdd.n2065 gnd 0.007668f
C3232 vdd.n2066 gnd 0.007668f
C3233 vdd.n2067 gnd 0.007668f
C3234 vdd.n2068 gnd 0.009526f
C3235 vdd.n2070 gnd 0.009526f
C3236 vdd.n2071 gnd 0.009526f
C3237 vdd.n2072 gnd 0.007668f
C3238 vdd.n2073 gnd 0.007668f
C3239 vdd.n2074 gnd 0.007668f
C3240 vdd.n2075 gnd 0.009526f
C3241 vdd.n2077 gnd 0.009526f
C3242 vdd.n2078 gnd 0.009526f
C3243 vdd.n2079 gnd 0.007668f
C3244 vdd.n2080 gnd 0.007668f
C3245 vdd.n2081 gnd 0.007668f
C3246 vdd.n2082 gnd 0.009526f
C3247 vdd.n2084 gnd 0.009526f
C3248 vdd.n2085 gnd 0.007668f
C3249 vdd.n2086 gnd 0.007668f
C3250 vdd.n2087 gnd 0.009526f
C3251 vdd.n2089 gnd 0.009526f
C3252 vdd.n2090 gnd 0.009526f
C3253 vdd.n2091 gnd 0.007668f
C3254 vdd.n2092 gnd 0.008193f
C3255 vdd.n2093 gnd 0.720431f
C3256 vdd.n2094 gnd 0.025963f
C3257 vdd.n2095 gnd 0.006478f
C3258 vdd.n2096 gnd 0.006478f
C3259 vdd.n2097 gnd 0.006478f
C3260 vdd.n2098 gnd 0.006478f
C3261 vdd.n2099 gnd 0.006478f
C3262 vdd.n2100 gnd 0.006478f
C3263 vdd.n2101 gnd 0.006478f
C3264 vdd.n2102 gnd 0.006478f
C3265 vdd.n2103 gnd 0.006478f
C3266 vdd.n2104 gnd 0.006478f
C3267 vdd.n2105 gnd 0.006478f
C3268 vdd.n2106 gnd 0.006478f
C3269 vdd.n2107 gnd 0.006478f
C3270 vdd.n2108 gnd 0.006478f
C3271 vdd.n2109 gnd 0.006478f
C3272 vdd.n2110 gnd 0.006478f
C3273 vdd.n2111 gnd 0.006478f
C3274 vdd.n2112 gnd 0.006478f
C3275 vdd.n2113 gnd 0.006478f
C3276 vdd.n2114 gnd 0.006478f
C3277 vdd.n2115 gnd 0.006478f
C3278 vdd.n2116 gnd 0.006478f
C3279 vdd.n2117 gnd 0.006478f
C3280 vdd.n2118 gnd 0.006478f
C3281 vdd.n2119 gnd 0.006478f
C3282 vdd.n2120 gnd 0.006478f
C3283 vdd.n2121 gnd 0.006478f
C3284 vdd.n2122 gnd 0.006478f
C3285 vdd.n2123 gnd 0.006478f
C3286 vdd.n2124 gnd 0.006478f
C3287 vdd.n2125 gnd 0.006478f
C3288 vdd.n2126 gnd 0.015151f
C3289 vdd.n2127 gnd 0.015151f
C3290 vdd.n2129 gnd 8.304331f
C3291 vdd.n2131 gnd 0.015151f
C3292 vdd.n2132 gnd 0.015151f
C3293 vdd.n2133 gnd 0.01419f
C3294 vdd.n2134 gnd 0.006478f
C3295 vdd.n2135 gnd 0.006478f
C3296 vdd.n2136 gnd 0.66201f
C3297 vdd.n2137 gnd 0.006478f
C3298 vdd.n2138 gnd 0.006478f
C3299 vdd.n2139 gnd 0.006478f
C3300 vdd.n2140 gnd 0.006478f
C3301 vdd.n2141 gnd 0.006478f
C3302 vdd.n2142 gnd 0.559788f
C3303 vdd.n2143 gnd 0.006478f
C3304 vdd.n2144 gnd 0.006478f
C3305 vdd.n2145 gnd 0.006478f
C3306 vdd.n2146 gnd 0.006478f
C3307 vdd.n2147 gnd 0.006478f
C3308 vdd.n2148 gnd 0.66201f
C3309 vdd.n2149 gnd 0.006478f
C3310 vdd.n2150 gnd 0.006478f
C3311 vdd.n2151 gnd 0.006478f
C3312 vdd.n2152 gnd 0.006478f
C3313 vdd.n2153 gnd 0.006478f
C3314 vdd.n2154 gnd 0.647407f
C3315 vdd.n2155 gnd 0.006478f
C3316 vdd.n2156 gnd 0.006478f
C3317 vdd.n2157 gnd 0.006478f
C3318 vdd.n2158 gnd 0.006478f
C3319 vdd.n2159 gnd 0.006478f
C3320 vdd.n2160 gnd 0.66201f
C3321 vdd.n2161 gnd 0.006478f
C3322 vdd.n2162 gnd 0.006478f
C3323 vdd.n2163 gnd 0.006478f
C3324 vdd.n2164 gnd 0.006478f
C3325 vdd.n2165 gnd 0.006478f
C3326 vdd.n2166 gnd 0.530581f
C3327 vdd.n2167 gnd 0.006478f
C3328 vdd.n2168 gnd 0.006478f
C3329 vdd.n2169 gnd 0.005525f
C3330 vdd.n2170 gnd 0.018766f
C3331 vdd.n2171 gnd 0.004192f
C3332 vdd.n2172 gnd 0.006478f
C3333 vdd.n2173 gnd 0.38455f
C3334 vdd.n2174 gnd 0.006478f
C3335 vdd.n2175 gnd 0.006478f
C3336 vdd.n2176 gnd 0.006478f
C3337 vdd.n2177 gnd 0.006478f
C3338 vdd.n2178 gnd 0.006478f
C3339 vdd.n2179 gnd 0.423492f
C3340 vdd.n2180 gnd 0.006478f
C3341 vdd.n2181 gnd 0.006478f
C3342 vdd.n2182 gnd 0.006478f
C3343 vdd.n2183 gnd 0.006478f
C3344 vdd.n2184 gnd 0.006478f
C3345 vdd.n2185 gnd 0.569523f
C3346 vdd.n2186 gnd 0.006478f
C3347 vdd.n2187 gnd 0.006478f
C3348 vdd.n2188 gnd 0.006478f
C3349 vdd.n2189 gnd 0.006478f
C3350 vdd.n2190 gnd 0.006478f
C3351 vdd.n2191 gnd 0.545185f
C3352 vdd.n2192 gnd 0.006478f
C3353 vdd.n2193 gnd 0.006478f
C3354 vdd.n2194 gnd 0.006478f
C3355 vdd.n2195 gnd 0.006478f
C3356 vdd.n2196 gnd 0.006478f
C3357 vdd.n2197 gnd 0.399153f
C3358 vdd.n2198 gnd 0.006478f
C3359 vdd.n2199 gnd 0.006478f
C3360 vdd.n2200 gnd 0.006478f
C3361 vdd.n2201 gnd 0.006478f
C3362 vdd.n2202 gnd 0.006478f
C3363 vdd.n2203 gnd 0.209312f
C3364 vdd.n2204 gnd 0.006478f
C3365 vdd.n2205 gnd 0.006478f
C3366 vdd.n2206 gnd 0.006478f
C3367 vdd.n2207 gnd 0.006478f
C3368 vdd.n2208 gnd 0.006478f
C3369 vdd.n2209 gnd 0.345608f
C3370 vdd.n2210 gnd 0.006478f
C3371 vdd.n2211 gnd 0.006478f
C3372 vdd.n2212 gnd 0.006478f
C3373 vdd.n2213 gnd 0.006478f
C3374 vdd.n2214 gnd 0.006478f
C3375 vdd.n2215 gnd 0.66201f
C3376 vdd.n2216 gnd 0.006478f
C3377 vdd.n2217 gnd 0.006478f
C3378 vdd.n2218 gnd 0.006478f
C3379 vdd.n2219 gnd 0.006478f
C3380 vdd.n2220 gnd 0.006478f
C3381 vdd.n2221 gnd 0.006478f
C3382 vdd.n2222 gnd 0.006478f
C3383 vdd.n2223 gnd 0.496507f
C3384 vdd.n2224 gnd 0.006478f
C3385 vdd.n2225 gnd 0.006478f
C3386 vdd.n2226 gnd 0.006478f
C3387 vdd.n2227 gnd 0.006478f
C3388 vdd.n2228 gnd 0.006478f
C3389 vdd.n2229 gnd 0.006478f
C3390 vdd.n2230 gnd 0.413756f
C3391 vdd.n2231 gnd 0.006478f
C3392 vdd.n2232 gnd 0.006478f
C3393 vdd.n2233 gnd 0.006478f
C3394 vdd.n2234 gnd 0.014994f
C3395 vdd.n2235 gnd 0.014347f
C3396 vdd.n2236 gnd 0.006478f
C3397 vdd.n2237 gnd 0.006478f
C3398 vdd.n2238 gnd 0.005001f
C3399 vdd.n2239 gnd 0.006478f
C3400 vdd.n2240 gnd 0.006478f
C3401 vdd.n2241 gnd 0.004716f
C3402 vdd.n2242 gnd 0.006478f
C3403 vdd.n2243 gnd 0.006478f
C3404 vdd.n2244 gnd 0.006478f
C3405 vdd.n2245 gnd 0.006478f
C3406 vdd.n2246 gnd 0.006478f
C3407 vdd.n2247 gnd 0.006478f
C3408 vdd.n2248 gnd 0.006478f
C3409 vdd.n2249 gnd 0.006478f
C3410 vdd.n2250 gnd 0.006478f
C3411 vdd.n2251 gnd 0.006478f
C3412 vdd.n2252 gnd 0.006478f
C3413 vdd.n2253 gnd 0.006478f
C3414 vdd.n2254 gnd 0.006478f
C3415 vdd.n2255 gnd 0.006478f
C3416 vdd.n2256 gnd 0.006478f
C3417 vdd.n2257 gnd 0.006478f
C3418 vdd.n2258 gnd 0.006478f
C3419 vdd.n2259 gnd 0.006478f
C3420 vdd.n2260 gnd 0.006478f
C3421 vdd.n2261 gnd 0.006478f
C3422 vdd.n2262 gnd 0.006478f
C3423 vdd.n2263 gnd 0.006478f
C3424 vdd.n2264 gnd 0.006478f
C3425 vdd.n2265 gnd 0.006478f
C3426 vdd.n2266 gnd 0.006478f
C3427 vdd.n2267 gnd 0.006478f
C3428 vdd.n2268 gnd 0.006478f
C3429 vdd.n2269 gnd 0.006478f
C3430 vdd.n2270 gnd 0.006478f
C3431 vdd.n2271 gnd 0.006478f
C3432 vdd.n2272 gnd 0.006478f
C3433 vdd.n2273 gnd 0.006478f
C3434 vdd.n2274 gnd 0.006478f
C3435 vdd.n2275 gnd 0.006478f
C3436 vdd.n2276 gnd 0.006478f
C3437 vdd.n2277 gnd 0.006478f
C3438 vdd.n2278 gnd 0.006478f
C3439 vdd.n2279 gnd 0.006478f
C3440 vdd.n2280 gnd 0.006478f
C3441 vdd.n2281 gnd 0.006478f
C3442 vdd.n2282 gnd 0.006478f
C3443 vdd.n2283 gnd 0.006478f
C3444 vdd.n2284 gnd 0.006478f
C3445 vdd.n2285 gnd 0.006478f
C3446 vdd.n2286 gnd 0.006478f
C3447 vdd.n2287 gnd 0.006478f
C3448 vdd.n2288 gnd 0.006478f
C3449 vdd.n2289 gnd 0.006478f
C3450 vdd.n2290 gnd 0.006478f
C3451 vdd.n2291 gnd 0.006478f
C3452 vdd.n2292 gnd 0.006478f
C3453 vdd.n2293 gnd 0.006478f
C3454 vdd.n2294 gnd 0.006478f
C3455 vdd.n2295 gnd 0.006478f
C3456 vdd.n2296 gnd 0.006478f
C3457 vdd.n2297 gnd 0.006478f
C3458 vdd.n2298 gnd 0.006478f
C3459 vdd.n2299 gnd 0.006478f
C3460 vdd.n2300 gnd 0.006478f
C3461 vdd.n2301 gnd 0.006478f
C3462 vdd.n2302 gnd 0.015151f
C3463 vdd.n2303 gnd 0.01419f
C3464 vdd.n2304 gnd 0.01419f
C3465 vdd.n2305 gnd 0.78857f
C3466 vdd.n2306 gnd 0.01419f
C3467 vdd.n2307 gnd 0.015151f
C3468 vdd.n2308 gnd 0.014347f
C3469 vdd.n2309 gnd 0.006478f
C3470 vdd.n2310 gnd 0.006478f
C3471 vdd.n2311 gnd 0.006478f
C3472 vdd.n2312 gnd 0.005001f
C3473 vdd.n2313 gnd 0.009258f
C3474 vdd.n2314 gnd 0.004716f
C3475 vdd.n2315 gnd 0.006478f
C3476 vdd.n2316 gnd 0.006478f
C3477 vdd.n2317 gnd 0.006478f
C3478 vdd.n2318 gnd 0.006478f
C3479 vdd.n2319 gnd 0.006478f
C3480 vdd.n2320 gnd 0.006478f
C3481 vdd.n2321 gnd 0.006478f
C3482 vdd.n2322 gnd 0.006478f
C3483 vdd.n2323 gnd 0.006478f
C3484 vdd.n2324 gnd 0.006478f
C3485 vdd.n2325 gnd 0.006478f
C3486 vdd.n2326 gnd 0.006478f
C3487 vdd.n2327 gnd 0.006478f
C3488 vdd.n2328 gnd 0.006478f
C3489 vdd.n2329 gnd 0.006478f
C3490 vdd.n2330 gnd 0.006478f
C3491 vdd.n2331 gnd 0.006478f
C3492 vdd.n2332 gnd 0.006478f
C3493 vdd.n2333 gnd 0.006478f
C3494 vdd.n2334 gnd 0.006478f
C3495 vdd.n2335 gnd 0.006478f
C3496 vdd.n2336 gnd 0.006478f
C3497 vdd.n2337 gnd 0.006478f
C3498 vdd.n2338 gnd 0.006478f
C3499 vdd.n2339 gnd 0.006478f
C3500 vdd.n2340 gnd 0.006478f
C3501 vdd.n2341 gnd 0.006478f
C3502 vdd.n2342 gnd 0.006478f
C3503 vdd.n2343 gnd 0.006478f
C3504 vdd.n2344 gnd 0.006478f
C3505 vdd.n2345 gnd 0.006478f
C3506 vdd.n2346 gnd 0.006478f
C3507 vdd.n2347 gnd 0.006478f
C3508 vdd.n2348 gnd 0.006478f
C3509 vdd.n2349 gnd 0.006478f
C3510 vdd.n2350 gnd 0.006478f
C3511 vdd.n2351 gnd 0.006478f
C3512 vdd.n2352 gnd 0.006478f
C3513 vdd.n2353 gnd 0.006478f
C3514 vdd.n2354 gnd 0.006478f
C3515 vdd.n2355 gnd 0.006478f
C3516 vdd.n2356 gnd 0.006478f
C3517 vdd.n2357 gnd 0.006478f
C3518 vdd.n2358 gnd 0.006478f
C3519 vdd.n2359 gnd 0.006478f
C3520 vdd.n2360 gnd 0.006478f
C3521 vdd.n2361 gnd 0.006478f
C3522 vdd.n2362 gnd 0.006478f
C3523 vdd.n2363 gnd 0.006478f
C3524 vdd.n2364 gnd 0.006478f
C3525 vdd.n2365 gnd 0.006478f
C3526 vdd.n2366 gnd 0.006478f
C3527 vdd.n2367 gnd 0.006478f
C3528 vdd.n2368 gnd 0.006478f
C3529 vdd.n2369 gnd 0.006478f
C3530 vdd.n2370 gnd 0.006478f
C3531 vdd.n2371 gnd 0.006478f
C3532 vdd.n2372 gnd 0.006478f
C3533 vdd.n2373 gnd 0.006478f
C3534 vdd.n2374 gnd 0.006478f
C3535 vdd.n2375 gnd 0.015151f
C3536 vdd.n2376 gnd 0.015151f
C3537 vdd.n2377 gnd 0.808041f
C3538 vdd.t120 gnd 2.87195f
C3539 vdd.t114 gnd 2.87195f
C3540 vdd.n2410 gnd 0.015151f
C3541 vdd.t129 gnd 0.603597f
C3542 vdd.n2411 gnd 0.006478f
C3543 vdd.n2412 gnd 0.006478f
C3544 vdd.t56 gnd 0.261771f
C3545 vdd.t57 gnd 0.267955f
C3546 vdd.t54 gnd 0.170894f
C3547 vdd.n2413 gnd 0.092359f
C3548 vdd.n2414 gnd 0.052389f
C3549 vdd.n2415 gnd 0.006478f
C3550 vdd.t66 gnd 0.261771f
C3551 vdd.t67 gnd 0.267955f
C3552 vdd.t65 gnd 0.170894f
C3553 vdd.n2416 gnd 0.092359f
C3554 vdd.n2417 gnd 0.052389f
C3555 vdd.n2418 gnd 0.009258f
C3556 vdd.n2419 gnd 0.006478f
C3557 vdd.n2420 gnd 0.006478f
C3558 vdd.n2421 gnd 0.006478f
C3559 vdd.n2422 gnd 0.006478f
C3560 vdd.n2423 gnd 0.006478f
C3561 vdd.n2424 gnd 0.006478f
C3562 vdd.n2425 gnd 0.006478f
C3563 vdd.n2426 gnd 0.006478f
C3564 vdd.n2427 gnd 0.006478f
C3565 vdd.n2428 gnd 0.006478f
C3566 vdd.n2429 gnd 0.006478f
C3567 vdd.n2430 gnd 0.006478f
C3568 vdd.n2431 gnd 0.006478f
C3569 vdd.n2432 gnd 0.006478f
C3570 vdd.n2433 gnd 0.006478f
C3571 vdd.n2434 gnd 0.006478f
C3572 vdd.n2435 gnd 0.006478f
C3573 vdd.n2436 gnd 0.006478f
C3574 vdd.n2437 gnd 0.006478f
C3575 vdd.n2438 gnd 0.006478f
C3576 vdd.n2439 gnd 0.006478f
C3577 vdd.n2440 gnd 0.006478f
C3578 vdd.n2441 gnd 0.006478f
C3579 vdd.n2442 gnd 0.006478f
C3580 vdd.n2443 gnd 0.006478f
C3581 vdd.n2444 gnd 0.006478f
C3582 vdd.n2445 gnd 0.006478f
C3583 vdd.n2446 gnd 0.006478f
C3584 vdd.n2447 gnd 0.006478f
C3585 vdd.n2448 gnd 0.006478f
C3586 vdd.n2449 gnd 0.006478f
C3587 vdd.n2450 gnd 0.006478f
C3588 vdd.n2451 gnd 0.006478f
C3589 vdd.n2452 gnd 0.006478f
C3590 vdd.n2453 gnd 0.006478f
C3591 vdd.n2454 gnd 0.006478f
C3592 vdd.n2455 gnd 0.006478f
C3593 vdd.n2456 gnd 0.006478f
C3594 vdd.n2457 gnd 0.006478f
C3595 vdd.n2458 gnd 0.006478f
C3596 vdd.n2459 gnd 0.006478f
C3597 vdd.n2460 gnd 0.006478f
C3598 vdd.n2461 gnd 0.006478f
C3599 vdd.n2462 gnd 0.006478f
C3600 vdd.n2463 gnd 0.006478f
C3601 vdd.n2464 gnd 0.006478f
C3602 vdd.n2465 gnd 0.006478f
C3603 vdd.n2466 gnd 0.006478f
C3604 vdd.n2467 gnd 0.006478f
C3605 vdd.n2468 gnd 0.006478f
C3606 vdd.n2469 gnd 0.006478f
C3607 vdd.n2470 gnd 0.006478f
C3608 vdd.n2471 gnd 0.006478f
C3609 vdd.n2472 gnd 0.006478f
C3610 vdd.n2473 gnd 0.006478f
C3611 vdd.n2474 gnd 0.006478f
C3612 vdd.n2475 gnd 0.006478f
C3613 vdd.n2476 gnd 0.006478f
C3614 vdd.n2477 gnd 0.004716f
C3615 vdd.n2478 gnd 0.006478f
C3616 vdd.n2479 gnd 0.006478f
C3617 vdd.n2480 gnd 0.005001f
C3618 vdd.n2481 gnd 0.006478f
C3619 vdd.n2482 gnd 0.006478f
C3620 vdd.n2483 gnd 0.015151f
C3621 vdd.n2484 gnd 0.01419f
C3622 vdd.n2485 gnd 0.01419f
C3623 vdd.n2486 gnd 0.006478f
C3624 vdd.n2487 gnd 0.006478f
C3625 vdd.n2488 gnd 0.006478f
C3626 vdd.n2489 gnd 0.006478f
C3627 vdd.n2490 gnd 0.006478f
C3628 vdd.n2491 gnd 0.006478f
C3629 vdd.n2492 gnd 0.006478f
C3630 vdd.n2493 gnd 0.006478f
C3631 vdd.n2494 gnd 0.006478f
C3632 vdd.n2495 gnd 0.006478f
C3633 vdd.n2496 gnd 0.006478f
C3634 vdd.n2497 gnd 0.006478f
C3635 vdd.n2498 gnd 0.006478f
C3636 vdd.n2499 gnd 0.006478f
C3637 vdd.n2500 gnd 0.006478f
C3638 vdd.n2501 gnd 0.006478f
C3639 vdd.n2502 gnd 0.006478f
C3640 vdd.n2503 gnd 0.006478f
C3641 vdd.n2504 gnd 0.006478f
C3642 vdd.n2505 gnd 0.006478f
C3643 vdd.n2506 gnd 0.006478f
C3644 vdd.n2507 gnd 0.006478f
C3645 vdd.n2508 gnd 0.006478f
C3646 vdd.n2509 gnd 0.006478f
C3647 vdd.n2510 gnd 0.006478f
C3648 vdd.n2511 gnd 0.006478f
C3649 vdd.n2512 gnd 0.006478f
C3650 vdd.n2513 gnd 0.006478f
C3651 vdd.n2514 gnd 0.006478f
C3652 vdd.n2515 gnd 0.006478f
C3653 vdd.n2516 gnd 0.006478f
C3654 vdd.n2517 gnd 0.006478f
C3655 vdd.n2518 gnd 0.006478f
C3656 vdd.n2519 gnd 0.006478f
C3657 vdd.n2520 gnd 0.006478f
C3658 vdd.n2521 gnd 0.006478f
C3659 vdd.n2522 gnd 0.006478f
C3660 vdd.n2523 gnd 0.006478f
C3661 vdd.n2524 gnd 0.006478f
C3662 vdd.n2525 gnd 0.006478f
C3663 vdd.n2526 gnd 0.006478f
C3664 vdd.n2527 gnd 0.006478f
C3665 vdd.n2528 gnd 0.006478f
C3666 vdd.n2529 gnd 0.006478f
C3667 vdd.n2530 gnd 0.006478f
C3668 vdd.n2531 gnd 0.006478f
C3669 vdd.n2532 gnd 0.006478f
C3670 vdd.n2533 gnd 0.006478f
C3671 vdd.n2534 gnd 0.006478f
C3672 vdd.n2535 gnd 0.006478f
C3673 vdd.n2536 gnd 0.006478f
C3674 vdd.n2537 gnd 0.006478f
C3675 vdd.n2538 gnd 0.006478f
C3676 vdd.n2539 gnd 0.006478f
C3677 vdd.n2540 gnd 0.006478f
C3678 vdd.n2541 gnd 0.006478f
C3679 vdd.n2542 gnd 0.006478f
C3680 vdd.n2543 gnd 0.006478f
C3681 vdd.n2544 gnd 0.006478f
C3682 vdd.n2545 gnd 0.006478f
C3683 vdd.n2546 gnd 0.006478f
C3684 vdd.n2547 gnd 0.006478f
C3685 vdd.n2548 gnd 0.006478f
C3686 vdd.n2549 gnd 0.006478f
C3687 vdd.n2550 gnd 0.006478f
C3688 vdd.n2551 gnd 0.006478f
C3689 vdd.n2552 gnd 0.006478f
C3690 vdd.n2553 gnd 0.006478f
C3691 vdd.n2554 gnd 0.006478f
C3692 vdd.n2555 gnd 0.006478f
C3693 vdd.n2556 gnd 0.006478f
C3694 vdd.n2557 gnd 0.006478f
C3695 vdd.n2558 gnd 0.006478f
C3696 vdd.n2559 gnd 0.209312f
C3697 vdd.n2560 gnd 0.006478f
C3698 vdd.n2561 gnd 0.006478f
C3699 vdd.n2562 gnd 0.006478f
C3700 vdd.n2563 gnd 0.006478f
C3701 vdd.n2564 gnd 0.006478f
C3702 vdd.n2565 gnd 0.006478f
C3703 vdd.n2566 gnd 0.006478f
C3704 vdd.n2567 gnd 0.006478f
C3705 vdd.n2568 gnd 0.006478f
C3706 vdd.n2569 gnd 0.006478f
C3707 vdd.n2570 gnd 0.006478f
C3708 vdd.n2571 gnd 0.006478f
C3709 vdd.n2572 gnd 0.006478f
C3710 vdd.n2573 gnd 0.006478f
C3711 vdd.n2574 gnd 0.413756f
C3712 vdd.n2575 gnd 0.006478f
C3713 vdd.n2576 gnd 0.006478f
C3714 vdd.n2577 gnd 0.006478f
C3715 vdd.n2578 gnd 0.01419f
C3716 vdd.n2579 gnd 0.01419f
C3717 vdd.n2580 gnd 0.015151f
C3718 vdd.n2581 gnd 0.015151f
C3719 vdd.n2582 gnd 0.006478f
C3720 vdd.n2583 gnd 0.006478f
C3721 vdd.n2584 gnd 0.006478f
C3722 vdd.n2585 gnd 0.005001f
C3723 vdd.n2586 gnd 0.009258f
C3724 vdd.n2587 gnd 0.004716f
C3725 vdd.n2588 gnd 0.006478f
C3726 vdd.n2589 gnd 0.006478f
C3727 vdd.n2590 gnd 0.006478f
C3728 vdd.n2591 gnd 0.006478f
C3729 vdd.n2592 gnd 0.006478f
C3730 vdd.n2593 gnd 0.006478f
C3731 vdd.n2594 gnd 0.006478f
C3732 vdd.n2595 gnd 0.006478f
C3733 vdd.n2596 gnd 0.006478f
C3734 vdd.n2597 gnd 0.006478f
C3735 vdd.n2598 gnd 0.006478f
C3736 vdd.n2599 gnd 0.006478f
C3737 vdd.n2600 gnd 0.006478f
C3738 vdd.n2601 gnd 0.006478f
C3739 vdd.n2602 gnd 0.006478f
C3740 vdd.n2603 gnd 0.006478f
C3741 vdd.n2604 gnd 0.006478f
C3742 vdd.n2605 gnd 0.006478f
C3743 vdd.n2606 gnd 0.006478f
C3744 vdd.n2607 gnd 0.006478f
C3745 vdd.n2608 gnd 0.006478f
C3746 vdd.n2609 gnd 0.006478f
C3747 vdd.n2610 gnd 0.006478f
C3748 vdd.n2611 gnd 0.006478f
C3749 vdd.n2612 gnd 0.006478f
C3750 vdd.n2613 gnd 0.006478f
C3751 vdd.n2614 gnd 0.006478f
C3752 vdd.n2615 gnd 0.006478f
C3753 vdd.n2616 gnd 0.006478f
C3754 vdd.n2617 gnd 0.006478f
C3755 vdd.n2618 gnd 0.006478f
C3756 vdd.n2619 gnd 0.006478f
C3757 vdd.n2620 gnd 0.006478f
C3758 vdd.n2621 gnd 0.006478f
C3759 vdd.n2622 gnd 0.006478f
C3760 vdd.n2623 gnd 0.006478f
C3761 vdd.n2624 gnd 0.006478f
C3762 vdd.n2625 gnd 0.006478f
C3763 vdd.n2626 gnd 0.006478f
C3764 vdd.n2627 gnd 0.006478f
C3765 vdd.n2628 gnd 0.006478f
C3766 vdd.n2629 gnd 0.006478f
C3767 vdd.n2630 gnd 0.006478f
C3768 vdd.n2631 gnd 0.006478f
C3769 vdd.n2632 gnd 0.006478f
C3770 vdd.n2633 gnd 0.006478f
C3771 vdd.n2634 gnd 0.006478f
C3772 vdd.n2635 gnd 0.006478f
C3773 vdd.n2636 gnd 0.006478f
C3774 vdd.n2637 gnd 0.006478f
C3775 vdd.n2638 gnd 0.006478f
C3776 vdd.n2639 gnd 0.006478f
C3777 vdd.n2640 gnd 0.006478f
C3778 vdd.n2641 gnd 0.006478f
C3779 vdd.n2642 gnd 0.006478f
C3780 vdd.n2643 gnd 0.006478f
C3781 vdd.n2644 gnd 0.006478f
C3782 vdd.n2645 gnd 0.006478f
C3783 vdd.n2646 gnd 0.006478f
C3784 vdd.n2647 gnd 0.015151f
C3785 vdd.n2648 gnd 0.015151f
C3786 vdd.n2650 gnd 0.808041f
C3787 vdd.n2652 gnd 0.015151f
C3788 vdd.n2653 gnd 0.015151f
C3789 vdd.n2654 gnd 0.01419f
C3790 vdd.n2655 gnd 0.006478f
C3791 vdd.n2656 gnd 0.006478f
C3792 vdd.n2657 gnd 0.350476f
C3793 vdd.n2658 gnd 0.006478f
C3794 vdd.n2659 gnd 0.006478f
C3795 vdd.n2660 gnd 0.006478f
C3796 vdd.n2661 gnd 0.006478f
C3797 vdd.n2662 gnd 0.006478f
C3798 vdd.n2663 gnd 0.394285f
C3799 vdd.n2664 gnd 0.006478f
C3800 vdd.n2665 gnd 0.006478f
C3801 vdd.n2666 gnd 0.006478f
C3802 vdd.n2667 gnd 0.006478f
C3803 vdd.n2668 gnd 0.006478f
C3804 vdd.n2669 gnd 0.66201f
C3805 vdd.n2670 gnd 0.006478f
C3806 vdd.n2671 gnd 0.006478f
C3807 vdd.n2672 gnd 0.006478f
C3808 vdd.n2673 gnd 0.006478f
C3809 vdd.n2674 gnd 0.006478f
C3810 vdd.n2675 gnd 0.438095f
C3811 vdd.n2676 gnd 0.006478f
C3812 vdd.n2677 gnd 0.006478f
C3813 vdd.n2678 gnd 0.006478f
C3814 vdd.n2679 gnd 0.006478f
C3815 vdd.n2680 gnd 0.006478f
C3816 vdd.n2681 gnd 0.584126f
C3817 vdd.n2682 gnd 0.006478f
C3818 vdd.n2683 gnd 0.006478f
C3819 vdd.n2684 gnd 0.006478f
C3820 vdd.n2685 gnd 0.006478f
C3821 vdd.n2686 gnd 0.006478f
C3822 vdd.n2687 gnd 0.530581f
C3823 vdd.n2688 gnd 0.006478f
C3824 vdd.n2689 gnd 0.006478f
C3825 vdd.n2690 gnd 0.006478f
C3826 vdd.n2691 gnd 0.006478f
C3827 vdd.n2692 gnd 0.006478f
C3828 vdd.n2693 gnd 0.38455f
C3829 vdd.n2694 gnd 0.006478f
C3830 vdd.n2695 gnd 0.006478f
C3831 vdd.n2696 gnd 0.006478f
C3832 vdd.n2697 gnd 0.006478f
C3833 vdd.n2698 gnd 0.006478f
C3834 vdd.n2699 gnd 0.209312f
C3835 vdd.n2700 gnd 0.006478f
C3836 vdd.n2701 gnd 0.006478f
C3837 vdd.n2702 gnd 0.006478f
C3838 vdd.n2703 gnd 0.006478f
C3839 vdd.n2704 gnd 0.006478f
C3840 vdd.n2705 gnd 0.569523f
C3841 vdd.n2706 gnd 0.006478f
C3842 vdd.n2707 gnd 0.006478f
C3843 vdd.n2708 gnd 0.006478f
C3844 vdd.n2709 gnd 0.006478f
C3845 vdd.n2710 gnd 0.006478f
C3846 vdd.n2711 gnd 0.66201f
C3847 vdd.n2712 gnd 0.006478f
C3848 vdd.n2713 gnd 0.006478f
C3849 vdd.n2714 gnd 0.004192f
C3850 vdd.n2715 gnd 0.018766f
C3851 vdd.n2716 gnd 0.005525f
C3852 vdd.n2717 gnd 0.006478f
C3853 vdd.n2718 gnd 0.564655f
C3854 vdd.n2719 gnd 0.006478f
C3855 vdd.n2720 gnd 0.006478f
C3856 vdd.n2721 gnd 0.006478f
C3857 vdd.n2722 gnd 0.006478f
C3858 vdd.n2723 gnd 0.006478f
C3859 vdd.n2724 gnd 0.462433f
C3860 vdd.n2725 gnd 0.006478f
C3861 vdd.n2726 gnd 0.006478f
C3862 vdd.n2727 gnd 0.006478f
C3863 vdd.n2728 gnd 0.006478f
C3864 vdd.n2729 gnd 0.006478f
C3865 vdd.n2730 gnd 0.345608f
C3866 vdd.n2731 gnd 0.006478f
C3867 vdd.n2732 gnd 0.006478f
C3868 vdd.n2733 gnd 0.006478f
C3869 vdd.n2734 gnd 0.006478f
C3870 vdd.n2735 gnd 0.006478f
C3871 vdd.n2736 gnd 0.66201f
C3872 vdd.n2737 gnd 0.006478f
C3873 vdd.n2738 gnd 0.006478f
C3874 vdd.n2739 gnd 0.006478f
C3875 vdd.n2740 gnd 0.006478f
C3876 vdd.n2741 gnd 0.006478f
C3877 vdd.n2742 gnd 0.006478f
C3878 vdd.n2744 gnd 0.006478f
C3879 vdd.n2745 gnd 0.006478f
C3880 vdd.n2747 gnd 0.006478f
C3881 vdd.n2748 gnd 0.006478f
C3882 vdd.n2751 gnd 0.006478f
C3883 vdd.n2752 gnd 0.006478f
C3884 vdd.n2753 gnd 0.006478f
C3885 vdd.n2754 gnd 0.006478f
C3886 vdd.n2756 gnd 0.006478f
C3887 vdd.n2757 gnd 0.006478f
C3888 vdd.n2758 gnd 0.006478f
C3889 vdd.n2759 gnd 0.006478f
C3890 vdd.n2760 gnd 0.006478f
C3891 vdd.n2761 gnd 0.006478f
C3892 vdd.n2763 gnd 0.006478f
C3893 vdd.n2764 gnd 0.006478f
C3894 vdd.n2765 gnd 0.006478f
C3895 vdd.n2766 gnd 0.006478f
C3896 vdd.n2767 gnd 0.006478f
C3897 vdd.n2768 gnd 0.006478f
C3898 vdd.n2770 gnd 0.006478f
C3899 vdd.n2771 gnd 0.006478f
C3900 vdd.n2772 gnd 0.006478f
C3901 vdd.n2773 gnd 0.006478f
C3902 vdd.n2774 gnd 0.006478f
C3903 vdd.n2775 gnd 0.006478f
C3904 vdd.n2777 gnd 0.006478f
C3905 vdd.n2778 gnd 0.015151f
C3906 vdd.n2779 gnd 0.015151f
C3907 vdd.n2780 gnd 0.01419f
C3908 vdd.n2781 gnd 0.006478f
C3909 vdd.n2782 gnd 0.006478f
C3910 vdd.n2783 gnd 0.006478f
C3911 vdd.n2784 gnd 0.006478f
C3912 vdd.n2785 gnd 0.006478f
C3913 vdd.n2786 gnd 0.006478f
C3914 vdd.n2787 gnd 0.66201f
C3915 vdd.n2788 gnd 0.006478f
C3916 vdd.n2789 gnd 0.006478f
C3917 vdd.n2790 gnd 0.006478f
C3918 vdd.n2791 gnd 0.006478f
C3919 vdd.n2792 gnd 0.006478f
C3920 vdd.n2793 gnd 0.433227f
C3921 vdd.n2794 gnd 0.006478f
C3922 vdd.n2795 gnd 0.006478f
C3923 vdd.n2796 gnd 0.006478f
C3924 vdd.n2797 gnd 0.014994f
C3925 vdd.n2799 gnd 0.015151f
C3926 vdd.n2800 gnd 0.014347f
C3927 vdd.n2801 gnd 0.006478f
C3928 vdd.n2802 gnd 0.005001f
C3929 vdd.n2803 gnd 0.006478f
C3930 vdd.n2805 gnd 0.006478f
C3931 vdd.n2806 gnd 0.006478f
C3932 vdd.n2807 gnd 0.006478f
C3933 vdd.n2808 gnd 0.006478f
C3934 vdd.n2809 gnd 0.006478f
C3935 vdd.n2810 gnd 0.006478f
C3936 vdd.n2812 gnd 0.006478f
C3937 vdd.n2813 gnd 0.006478f
C3938 vdd.n2814 gnd 0.006478f
C3939 vdd.n2815 gnd 0.006478f
C3940 vdd.n2816 gnd 0.006478f
C3941 vdd.n2817 gnd 0.006478f
C3942 vdd.n2819 gnd 0.006478f
C3943 vdd.n2820 gnd 0.006478f
C3944 vdd.n2821 gnd 0.006478f
C3945 vdd.n2822 gnd 0.006478f
C3946 vdd.n2823 gnd 0.006478f
C3947 vdd.n2824 gnd 0.006478f
C3948 vdd.n2826 gnd 0.006478f
C3949 vdd.n2827 gnd 0.006478f
C3950 vdd.n2828 gnd 0.006478f
C3951 vdd.n2829 gnd 0.724147f
C3952 vdd.n2830 gnd 0.022247f
C3953 vdd.n2831 gnd 0.006478f
C3954 vdd.n2832 gnd 0.006478f
C3955 vdd.n2834 gnd 0.006478f
C3956 vdd.n2835 gnd 0.006478f
C3957 vdd.n2836 gnd 0.006478f
C3958 vdd.n2837 gnd 0.006478f
C3959 vdd.n2838 gnd 0.006478f
C3960 vdd.n2839 gnd 0.006478f
C3961 vdd.n2841 gnd 0.006478f
C3962 vdd.n2842 gnd 0.006478f
C3963 vdd.n2843 gnd 0.006478f
C3964 vdd.n2844 gnd 0.006478f
C3965 vdd.n2845 gnd 0.006478f
C3966 vdd.n2846 gnd 0.006478f
C3967 vdd.n2848 gnd 0.006478f
C3968 vdd.n2849 gnd 0.006478f
C3969 vdd.n2850 gnd 0.006478f
C3970 vdd.n2851 gnd 0.006478f
C3971 vdd.n2852 gnd 0.006478f
C3972 vdd.n2853 gnd 0.006478f
C3973 vdd.n2855 gnd 0.006478f
C3974 vdd.n2856 gnd 0.006478f
C3975 vdd.n2858 gnd 0.006478f
C3976 vdd.n2859 gnd 0.006478f
C3977 vdd.n2860 gnd 0.015151f
C3978 vdd.n2861 gnd 0.01419f
C3979 vdd.n2862 gnd 0.01419f
C3980 vdd.n2863 gnd 0.934602f
C3981 vdd.n2864 gnd 0.01419f
C3982 vdd.n2865 gnd 0.015151f
C3983 vdd.n2866 gnd 0.014347f
C3984 vdd.n2867 gnd 0.006478f
C3985 vdd.n2868 gnd 0.005001f
C3986 vdd.n2869 gnd 0.006478f
C3987 vdd.n2871 gnd 0.006478f
C3988 vdd.n2872 gnd 0.006478f
C3989 vdd.n2873 gnd 0.006478f
C3990 vdd.n2874 gnd 0.006478f
C3991 vdd.n2875 gnd 0.006478f
C3992 vdd.n2876 gnd 0.006478f
C3993 vdd.n2878 gnd 0.006478f
C3994 vdd.n2879 gnd 0.006478f
C3995 vdd.n2880 gnd 0.006478f
C3996 vdd.n2881 gnd 0.006478f
C3997 vdd.n2882 gnd 0.006478f
C3998 vdd.n2883 gnd 0.006478f
C3999 vdd.n2885 gnd 0.006478f
C4000 vdd.n2886 gnd 0.006478f
C4001 vdd.n2887 gnd 0.006478f
C4002 vdd.n2888 gnd 0.006478f
C4003 vdd.n2889 gnd 0.006478f
C4004 vdd.n2890 gnd 0.006478f
C4005 vdd.n2892 gnd 0.006478f
C4006 vdd.n2893 gnd 0.006478f
C4007 vdd.n2895 gnd 0.006478f
C4008 vdd.n2896 gnd 0.022247f
C4009 vdd.n2897 gnd 0.724147f
C4010 vdd.n2898 gnd 0.008193f
C4011 vdd.n2899 gnd 0.003642f
C4012 vdd.t14 gnd 0.117199f
C4013 vdd.t15 gnd 0.125253f
C4014 vdd.t12 gnd 0.15306f
C4015 vdd.n2900 gnd 0.196201f
C4016 vdd.n2901 gnd 0.164844f
C4017 vdd.n2902 gnd 0.011808f
C4018 vdd.n2903 gnd 0.009526f
C4019 vdd.n2904 gnd 0.004025f
C4020 vdd.n2905 gnd 0.007668f
C4021 vdd.n2906 gnd 0.009526f
C4022 vdd.n2907 gnd 0.009526f
C4023 vdd.n2908 gnd 0.007668f
C4024 vdd.n2909 gnd 0.007668f
C4025 vdd.n2910 gnd 0.009526f
C4026 vdd.n2912 gnd 0.009526f
C4027 vdd.n2913 gnd 0.007668f
C4028 vdd.n2914 gnd 0.007668f
C4029 vdd.n2915 gnd 0.007668f
C4030 vdd.n2916 gnd 0.009526f
C4031 vdd.n2918 gnd 0.009526f
C4032 vdd.n2920 gnd 0.009526f
C4033 vdd.n2921 gnd 0.007668f
C4034 vdd.n2922 gnd 0.007668f
C4035 vdd.n2923 gnd 0.007668f
C4036 vdd.n2924 gnd 0.009526f
C4037 vdd.n2926 gnd 0.009526f
C4038 vdd.n2928 gnd 0.009526f
C4039 vdd.n2929 gnd 0.007668f
C4040 vdd.n2930 gnd 0.007668f
C4041 vdd.n2931 gnd 0.007668f
C4042 vdd.n2932 gnd 0.009526f
C4043 vdd.n2934 gnd 0.009526f
C4044 vdd.n2935 gnd 0.009526f
C4045 vdd.n2936 gnd 0.007668f
C4046 vdd.n2937 gnd 0.007668f
C4047 vdd.n2938 gnd 0.009526f
C4048 vdd.n2939 gnd 0.009526f
C4049 vdd.n2941 gnd 0.009526f
C4050 vdd.n2942 gnd 0.007668f
C4051 vdd.n2943 gnd 0.009526f
C4052 vdd.n2944 gnd 0.009526f
C4053 vdd.n2945 gnd 0.009526f
C4054 vdd.n2946 gnd 0.015642f
C4055 vdd.n2947 gnd 0.005214f
C4056 vdd.n2948 gnd 0.009526f
C4057 vdd.n2950 gnd 0.009526f
C4058 vdd.n2952 gnd 0.009526f
C4059 vdd.n2953 gnd 0.007668f
C4060 vdd.n2954 gnd 0.007668f
C4061 vdd.n2955 gnd 0.007668f
C4062 vdd.n2956 gnd 0.009526f
C4063 vdd.n2958 gnd 0.009526f
C4064 vdd.n2960 gnd 0.009526f
C4065 vdd.n2961 gnd 0.007668f
C4066 vdd.n2962 gnd 0.007668f
C4067 vdd.n2963 gnd 0.007668f
C4068 vdd.n2964 gnd 0.009526f
C4069 vdd.n2966 gnd 0.009526f
C4070 vdd.n2968 gnd 0.009526f
C4071 vdd.n2969 gnd 0.007668f
C4072 vdd.n2970 gnd 0.007668f
C4073 vdd.n2971 gnd 0.007668f
C4074 vdd.n2972 gnd 0.009526f
C4075 vdd.n2974 gnd 0.009526f
C4076 vdd.n2976 gnd 0.009526f
C4077 vdd.n2977 gnd 0.007668f
C4078 vdd.n2978 gnd 0.007668f
C4079 vdd.n2979 gnd 0.007668f
C4080 vdd.n2980 gnd 0.009526f
C4081 vdd.n2982 gnd 0.009526f
C4082 vdd.n2984 gnd 0.009526f
C4083 vdd.n2985 gnd 0.007668f
C4084 vdd.n2986 gnd 0.007668f
C4085 vdd.n2987 gnd 0.006402f
C4086 vdd.n2988 gnd 0.009526f
C4087 vdd.n2990 gnd 0.009526f
C4088 vdd.n2992 gnd 0.009526f
C4089 vdd.n2993 gnd 0.006402f
C4090 vdd.n2994 gnd 0.007668f
C4091 vdd.n2995 gnd 0.007668f
C4092 vdd.n2996 gnd 0.009526f
C4093 vdd.n2998 gnd 0.009526f
C4094 vdd.n3000 gnd 0.009526f
C4095 vdd.n3001 gnd 0.007668f
C4096 vdd.n3002 gnd 0.007668f
C4097 vdd.n3003 gnd 0.007668f
C4098 vdd.n3004 gnd 0.009526f
C4099 vdd.n3006 gnd 0.009526f
C4100 vdd.n3008 gnd 0.009526f
C4101 vdd.n3009 gnd 0.007668f
C4102 vdd.n3010 gnd 0.007668f
C4103 vdd.n3011 gnd 0.007668f
C4104 vdd.n3012 gnd 0.009526f
C4105 vdd.n3014 gnd 0.009526f
C4106 vdd.n3015 gnd 0.009526f
C4107 vdd.n3016 gnd 0.007668f
C4108 vdd.n3017 gnd 0.007668f
C4109 vdd.n3018 gnd 0.009526f
C4110 vdd.n3019 gnd 0.009526f
C4111 vdd.n3020 gnd 0.007668f
C4112 vdd.n3021 gnd 0.007668f
C4113 vdd.n3022 gnd 0.009526f
C4114 vdd.n3023 gnd 0.009526f
C4115 vdd.n3025 gnd 0.009526f
C4116 vdd.n3026 gnd 0.007668f
C4117 vdd.n3027 gnd 0.006364f
C4118 vdd.n3028 gnd 0.0228f
C4119 vdd.n3029 gnd 0.02245f
C4120 vdd.n3030 gnd 0.006364f
C4121 vdd.n3031 gnd 0.02245f
C4122 vdd.n3032 gnd 1.33862f
C4123 vdd.n3033 gnd 0.02245f
C4124 vdd.n3034 gnd 0.006364f
C4125 vdd.n3035 gnd 0.02245f
C4126 vdd.n3036 gnd 0.009526f
C4127 vdd.n3037 gnd 0.009526f
C4128 vdd.n3038 gnd 0.007668f
C4129 vdd.n3039 gnd 0.009526f
C4130 vdd.n3040 gnd 0.973544f
C4131 vdd.n3041 gnd 0.009526f
C4132 vdd.n3042 gnd 0.007668f
C4133 vdd.n3043 gnd 0.009526f
C4134 vdd.n3044 gnd 0.009526f
C4135 vdd.n3045 gnd 0.009526f
C4136 vdd.n3046 gnd 0.007668f
C4137 vdd.n3047 gnd 0.009526f
C4138 vdd.n3048 gnd 0.861586f
C4139 vdd.n3049 gnd 0.009526f
C4140 vdd.n3050 gnd 0.007668f
C4141 vdd.n3051 gnd 0.009526f
C4142 vdd.n3052 gnd 0.009526f
C4143 vdd.n3053 gnd 0.009526f
C4144 vdd.n3054 gnd 0.007668f
C4145 vdd.n3055 gnd 0.009526f
C4146 vdd.t204 gnd 0.486772f
C4147 vdd.n3056 gnd 0.696084f
C4148 vdd.n3057 gnd 0.009526f
C4149 vdd.n3058 gnd 0.007668f
C4150 vdd.n3059 gnd 0.009526f
C4151 vdd.n3060 gnd 0.009526f
C4152 vdd.n3061 gnd 0.009526f
C4153 vdd.n3062 gnd 0.007668f
C4154 vdd.n3063 gnd 0.009526f
C4155 vdd.n3064 gnd 0.530581f
C4156 vdd.n3065 gnd 0.009526f
C4157 vdd.n3066 gnd 0.007668f
C4158 vdd.n3067 gnd 0.009526f
C4159 vdd.n3068 gnd 0.009526f
C4160 vdd.n3069 gnd 0.009526f
C4161 vdd.n3070 gnd 0.007668f
C4162 vdd.n3071 gnd 0.009526f
C4163 vdd.n3072 gnd 0.686348f
C4164 vdd.n3073 gnd 0.608465f
C4165 vdd.n3074 gnd 0.009526f
C4166 vdd.n3075 gnd 0.007668f
C4167 vdd.n3076 gnd 0.009526f
C4168 vdd.n3077 gnd 0.009526f
C4169 vdd.n3078 gnd 0.009526f
C4170 vdd.n3079 gnd 0.007668f
C4171 vdd.n3080 gnd 0.009526f
C4172 vdd.n3081 gnd 0.773967f
C4173 vdd.n3082 gnd 0.009526f
C4174 vdd.n3083 gnd 0.007668f
C4175 vdd.n3084 gnd 0.009526f
C4176 vdd.n3085 gnd 0.009526f
C4177 vdd.n3086 gnd 0.009526f
C4178 vdd.n3087 gnd 0.007668f
C4179 vdd.n3088 gnd 0.007668f
C4180 vdd.n3089 gnd 0.007668f
C4181 vdd.n3090 gnd 0.009526f
C4182 vdd.n3091 gnd 0.009526f
C4183 vdd.n3092 gnd 0.009526f
C4184 vdd.n3093 gnd 0.007668f
C4185 vdd.n3094 gnd 0.007668f
C4186 vdd.n3095 gnd 0.007668f
C4187 vdd.n3096 gnd 0.009526f
C4188 vdd.n3097 gnd 0.009526f
C4189 vdd.n3098 gnd 0.009526f
C4190 vdd.n3099 gnd 0.007668f
C4191 vdd.n3100 gnd 0.007668f
C4192 vdd.n3101 gnd 0.007668f
C4193 vdd.n3102 gnd 0.009526f
C4194 vdd.n3103 gnd 0.009526f
C4195 vdd.n3104 gnd 0.009526f
C4196 vdd.n3105 gnd 0.007668f
C4197 vdd.n3106 gnd 0.007668f
C4198 vdd.n3107 gnd 0.006364f
C4199 vdd.n3108 gnd 0.02245f
C4200 vdd.n3109 gnd 0.0228f
C4201 vdd.n3111 gnd 0.0228f
C4202 vdd.n3112 gnd 0.003642f
C4203 vdd.t23 gnd 0.117199f
C4204 vdd.t22 gnd 0.125253f
C4205 vdd.t20 gnd 0.15306f
C4206 vdd.n3113 gnd 0.196201f
C4207 vdd.n3114 gnd 0.165611f
C4208 vdd.n3115 gnd 0.012575f
C4209 vdd.n3116 gnd 0.004025f
C4210 vdd.n3117 gnd 0.007668f
C4211 vdd.n3118 gnd 0.009526f
C4212 vdd.n3120 gnd 0.009526f
C4213 vdd.n3121 gnd 0.009526f
C4214 vdd.n3122 gnd 0.007668f
C4215 vdd.n3123 gnd 0.007668f
C4216 vdd.n3124 gnd 0.007668f
C4217 vdd.n3125 gnd 0.009526f
C4218 vdd.n3127 gnd 0.009526f
C4219 vdd.n3128 gnd 0.009526f
C4220 vdd.n3129 gnd 0.007668f
C4221 vdd.n3130 gnd 0.007668f
C4222 vdd.n3131 gnd 0.007668f
C4223 vdd.n3132 gnd 0.009526f
C4224 vdd.n3134 gnd 0.009526f
C4225 vdd.n3135 gnd 0.009526f
C4226 vdd.n3136 gnd 0.007668f
C4227 vdd.n3137 gnd 0.007668f
C4228 vdd.n3138 gnd 0.007668f
C4229 vdd.n3139 gnd 0.009526f
C4230 vdd.n3141 gnd 0.009526f
C4231 vdd.n3142 gnd 0.009526f
C4232 vdd.n3143 gnd 0.007668f
C4233 vdd.n3144 gnd 0.007668f
C4234 vdd.n3145 gnd 0.007668f
C4235 vdd.n3146 gnd 0.009526f
C4236 vdd.n3148 gnd 0.009526f
C4237 vdd.n3149 gnd 0.009526f
C4238 vdd.n3150 gnd 0.007668f
C4239 vdd.n3151 gnd 0.009526f
C4240 vdd.n3152 gnd 0.009526f
C4241 vdd.n3153 gnd 0.009526f
C4242 vdd.n3154 gnd 0.016409f
C4243 vdd.n3155 gnd 0.005214f
C4244 vdd.n3156 gnd 0.007668f
C4245 vdd.n3157 gnd 0.009526f
C4246 vdd.n3159 gnd 0.009526f
C4247 vdd.n3160 gnd 0.009526f
C4248 vdd.n3161 gnd 0.007668f
C4249 vdd.n3162 gnd 0.007668f
C4250 vdd.n3163 gnd 0.007668f
C4251 vdd.n3164 gnd 0.009526f
C4252 vdd.n3166 gnd 0.009526f
C4253 vdd.n3167 gnd 0.009526f
C4254 vdd.n3168 gnd 0.007668f
C4255 vdd.n3169 gnd 0.007668f
C4256 vdd.n3170 gnd 0.007668f
C4257 vdd.n3171 gnd 0.009526f
C4258 vdd.n3173 gnd 0.009526f
C4259 vdd.n3174 gnd 0.009526f
C4260 vdd.n3175 gnd 0.007668f
C4261 vdd.n3176 gnd 0.007668f
C4262 vdd.n3177 gnd 0.007668f
C4263 vdd.n3178 gnd 0.009526f
C4264 vdd.n3180 gnd 0.009526f
C4265 vdd.n3181 gnd 0.009526f
C4266 vdd.n3182 gnd 0.007668f
C4267 vdd.n3183 gnd 0.007668f
C4268 vdd.n3184 gnd 0.007668f
C4269 vdd.n3185 gnd 0.009526f
C4270 vdd.n3187 gnd 0.009526f
C4271 vdd.n3188 gnd 0.009526f
C4272 vdd.n3189 gnd 0.007668f
C4273 vdd.n3190 gnd 0.009526f
C4274 vdd.n3191 gnd 0.009526f
C4275 vdd.n3192 gnd 0.009526f
C4276 vdd.n3193 gnd 0.016409f
C4277 vdd.n3194 gnd 0.006402f
C4278 vdd.n3195 gnd 0.007668f
C4279 vdd.n3196 gnd 0.009526f
C4280 vdd.n3198 gnd 0.009526f
C4281 vdd.n3199 gnd 0.009526f
C4282 vdd.n3200 gnd 0.007668f
C4283 vdd.n3201 gnd 0.007668f
C4284 vdd.n3202 gnd 0.007668f
C4285 vdd.n3203 gnd 0.009526f
C4286 vdd.n3205 gnd 0.009526f
C4287 vdd.n3206 gnd 0.009526f
C4288 vdd.n3207 gnd 0.007668f
C4289 vdd.n3208 gnd 0.007668f
C4290 vdd.n3209 gnd 0.007668f
C4291 vdd.n3210 gnd 0.009526f
C4292 vdd.n3212 gnd 0.009526f
C4293 vdd.n3213 gnd 0.009526f
C4294 vdd.n3214 gnd 0.007668f
C4295 vdd.n3215 gnd 0.007668f
C4296 vdd.n3216 gnd 0.007668f
C4297 vdd.n3217 gnd 0.009526f
C4298 vdd.n3219 gnd 0.009526f
C4299 vdd.n3220 gnd 0.009526f
C4300 vdd.n3222 gnd 0.009526f
C4301 vdd.n3223 gnd 0.007668f
C4302 vdd.n3224 gnd 0.007668f
C4303 vdd.n3225 gnd 0.006364f
C4304 vdd.n3226 gnd 0.0228f
C4305 vdd.n3227 gnd 0.02245f
C4306 vdd.n3228 gnd 0.006364f
C4307 vdd.n3229 gnd 0.02245f
C4308 vdd.n3230 gnd 1.3727f
C4309 vdd.n3231 gnd 0.550052f
C4310 vdd.t21 gnd 0.486772f
C4311 vdd.n3232 gnd 0.910263f
C4312 vdd.n3233 gnd 0.009526f
C4313 vdd.n3234 gnd 0.007668f
C4314 vdd.n3235 gnd 0.007668f
C4315 vdd.n3236 gnd 0.007668f
C4316 vdd.n3237 gnd 0.009526f
C4317 vdd.n3238 gnd 0.958941f
C4318 vdd.t151 gnd 0.486772f
C4319 vdd.n3239 gnd 0.501375f
C4320 vdd.n3240 gnd 0.793438f
C4321 vdd.n3241 gnd 0.009526f
C4322 vdd.n3242 gnd 0.007668f
C4323 vdd.n3243 gnd 0.007668f
C4324 vdd.n3244 gnd 0.007668f
C4325 vdd.n3245 gnd 0.009526f
C4326 vdd.n3246 gnd 0.627936f
C4327 vdd.t167 gnd 0.486772f
C4328 vdd.n3247 gnd 0.808041f
C4329 vdd.t187 gnd 0.486772f
C4330 vdd.n3248 gnd 0.511111f
C4331 vdd.n3249 gnd 0.009526f
C4332 vdd.n3250 gnd 0.007668f
C4333 vdd.n3251 gnd 0.007668f
C4334 vdd.n3252 gnd 0.007668f
C4335 vdd.n3253 gnd 0.009526f
C4336 vdd.n3254 gnd 0.676613f
C4337 vdd.n3255 gnd 0.6182f
C4338 vdd.t164 gnd 0.486772f
C4339 vdd.n3256 gnd 0.808041f
C4340 vdd.n3257 gnd 0.009526f
C4341 vdd.n3258 gnd 0.007668f
C4342 vdd.n3259 gnd 0.56708f
C4343 vdd.n3260 gnd 2.21436f
C4344 a_n6972_8799.n0 gnd 4.27785f
C4345 a_n6972_8799.n1 gnd 2.09379f
C4346 a_n6972_8799.n2 gnd 3.51585f
C4347 a_n6972_8799.n3 gnd 0.876714f
C4348 a_n6972_8799.n4 gnd 0.177106f
C4349 a_n6972_8799.n5 gnd 0.207402f
C4350 a_n6972_8799.n6 gnd 0.207402f
C4351 a_n6972_8799.n7 gnd 0.207402f
C4352 a_n6972_8799.n8 gnd 0.177106f
C4353 a_n6972_8799.n9 gnd 0.207402f
C4354 a_n6972_8799.n10 gnd 0.207402f
C4355 a_n6972_8799.n11 gnd 0.207402f
C4356 a_n6972_8799.n12 gnd 0.342106f
C4357 a_n6972_8799.n13 gnd 0.207402f
C4358 a_n6972_8799.n14 gnd 0.207402f
C4359 a_n6972_8799.n15 gnd 0.207402f
C4360 a_n6972_8799.n16 gnd 0.207402f
C4361 a_n6972_8799.n17 gnd 0.207402f
C4362 a_n6972_8799.n18 gnd 0.177106f
C4363 a_n6972_8799.n19 gnd 0.207402f
C4364 a_n6972_8799.n20 gnd 0.207402f
C4365 a_n6972_8799.n21 gnd 0.207402f
C4366 a_n6972_8799.n22 gnd 0.177106f
C4367 a_n6972_8799.n23 gnd 0.207402f
C4368 a_n6972_8799.n24 gnd 0.207402f
C4369 a_n6972_8799.n25 gnd 0.207402f
C4370 a_n6972_8799.n26 gnd 0.342106f
C4371 a_n6972_8799.n27 gnd 0.207402f
C4372 a_n6972_8799.n28 gnd 1.0182f
C4373 a_n6972_8799.n29 gnd 2.48947f
C4374 a_n6972_8799.n30 gnd 1.52009f
C4375 a_n6972_8799.n31 gnd 0.250817f
C4376 a_n6972_8799.n33 gnd 0.007725f
C4377 a_n6972_8799.n34 gnd 0.011676f
C4378 a_n6972_8799.n35 gnd 0.00803f
C4379 a_n6972_8799.n37 gnd 4.01e-19
C4380 a_n6972_8799.n38 gnd 0.008322f
C4381 a_n6972_8799.n39 gnd 0.262385f
C4382 a_n6972_8799.n40 gnd 0.250817f
C4383 a_n6972_8799.n42 gnd 0.007725f
C4384 a_n6972_8799.n43 gnd 0.011676f
C4385 a_n6972_8799.n44 gnd 0.00803f
C4386 a_n6972_8799.n46 gnd 4.01e-19
C4387 a_n6972_8799.n47 gnd 0.008322f
C4388 a_n6972_8799.n48 gnd 0.262385f
C4389 a_n6972_8799.n49 gnd 0.250817f
C4390 a_n6972_8799.n51 gnd 0.007725f
C4391 a_n6972_8799.n52 gnd 0.011676f
C4392 a_n6972_8799.n53 gnd 0.00803f
C4393 a_n6972_8799.n55 gnd 4.01e-19
C4394 a_n6972_8799.n56 gnd 0.008322f
C4395 a_n6972_8799.n57 gnd 0.262385f
C4396 a_n6972_8799.n58 gnd 0.008322f
C4397 a_n6972_8799.n59 gnd 0.262385f
C4398 a_n6972_8799.n60 gnd 4.01e-19
C4399 a_n6972_8799.n62 gnd 0.00803f
C4400 a_n6972_8799.n63 gnd 0.011676f
C4401 a_n6972_8799.n64 gnd 0.007725f
C4402 a_n6972_8799.n66 gnd 0.250817f
C4403 a_n6972_8799.n67 gnd 0.008322f
C4404 a_n6972_8799.n68 gnd 0.262385f
C4405 a_n6972_8799.n69 gnd 4.01e-19
C4406 a_n6972_8799.n71 gnd 0.00803f
C4407 a_n6972_8799.n72 gnd 0.011676f
C4408 a_n6972_8799.n73 gnd 0.007725f
C4409 a_n6972_8799.n75 gnd 0.250817f
C4410 a_n6972_8799.n76 gnd 0.008322f
C4411 a_n6972_8799.n77 gnd 0.262385f
C4412 a_n6972_8799.n78 gnd 4.01e-19
C4413 a_n6972_8799.n80 gnd 0.00803f
C4414 a_n6972_8799.n81 gnd 0.011676f
C4415 a_n6972_8799.n82 gnd 0.007725f
C4416 a_n6972_8799.n84 gnd 0.250817f
C4417 a_n6972_8799.t21 gnd 0.143856f
C4418 a_n6972_8799.t17 gnd 0.143856f
C4419 a_n6972_8799.t27 gnd 0.143856f
C4420 a_n6972_8799.n85 gnd 1.13462f
C4421 a_n6972_8799.t25 gnd 0.143856f
C4422 a_n6972_8799.t6 gnd 0.143856f
C4423 a_n6972_8799.n86 gnd 1.13274f
C4424 a_n6972_8799.t33 gnd 0.143856f
C4425 a_n6972_8799.t22 gnd 0.143856f
C4426 a_n6972_8799.n87 gnd 1.13274f
C4427 a_n6972_8799.t7 gnd 0.143856f
C4428 a_n6972_8799.t30 gnd 0.143856f
C4429 a_n6972_8799.n88 gnd 1.13274f
C4430 a_n6972_8799.t20 gnd 0.111888f
C4431 a_n6972_8799.t35 gnd 0.111888f
C4432 a_n6972_8799.n89 gnd 0.991598f
C4433 a_n6972_8799.t37 gnd 0.111888f
C4434 a_n6972_8799.t8 gnd 0.111888f
C4435 a_n6972_8799.n90 gnd 0.988683f
C4436 a_n6972_8799.t29 gnd 0.111888f
C4437 a_n6972_8799.t24 gnd 0.111888f
C4438 a_n6972_8799.n91 gnd 0.988683f
C4439 a_n6972_8799.t9 gnd 0.111888f
C4440 a_n6972_8799.t0 gnd 0.111888f
C4441 a_n6972_8799.n92 gnd 0.991597f
C4442 a_n6972_8799.t34 gnd 0.111888f
C4443 a_n6972_8799.t36 gnd 0.111888f
C4444 a_n6972_8799.n93 gnd 0.988682f
C4445 a_n6972_8799.t14 gnd 0.111888f
C4446 a_n6972_8799.t12 gnd 0.111888f
C4447 a_n6972_8799.n94 gnd 0.988682f
C4448 a_n6972_8799.t23 gnd 0.111888f
C4449 a_n6972_8799.t13 gnd 0.111888f
C4450 a_n6972_8799.n95 gnd 0.991597f
C4451 a_n6972_8799.t10 gnd 0.111888f
C4452 a_n6972_8799.t18 gnd 0.111888f
C4453 a_n6972_8799.n96 gnd 0.988682f
C4454 a_n6972_8799.t3 gnd 0.111888f
C4455 a_n6972_8799.t2 gnd 0.111888f
C4456 a_n6972_8799.n97 gnd 0.988682f
C4457 a_n6972_8799.t1 gnd 0.111888f
C4458 a_n6972_8799.t32 gnd 0.111888f
C4459 a_n6972_8799.n98 gnd 0.988683f
C4460 a_n6972_8799.t4 gnd 0.111888f
C4461 a_n6972_8799.t28 gnd 0.111888f
C4462 a_n6972_8799.n99 gnd 0.988683f
C4463 a_n6972_8799.t11 gnd 0.111888f
C4464 a_n6972_8799.t15 gnd 0.111888f
C4465 a_n6972_8799.n100 gnd 0.988683f
C4466 a_n6972_8799.t72 gnd 0.596495f
C4467 a_n6972_8799.n101 gnd 0.269967f
C4468 a_n6972_8799.t100 gnd 0.596495f
C4469 a_n6972_8799.t40 gnd 0.596495f
C4470 a_n6972_8799.n102 gnd 0.261131f
C4471 a_n6972_8799.t61 gnd 0.596495f
C4472 a_n6972_8799.n103 gnd 0.272496f
C4473 a_n6972_8799.t62 gnd 0.596495f
C4474 a_n6972_8799.t69 gnd 0.596495f
C4475 a_n6972_8799.n104 gnd 0.265926f
C4476 a_n6972_8799.t99 gnd 0.610514f
C4477 a_n6972_8799.t68 gnd 0.596495f
C4478 a_n6972_8799.n105 gnd 0.272062f
C4479 a_n6972_8799.n106 gnd 0.248651f
C4480 a_n6972_8799.t86 gnd 0.596495f
C4481 a_n6972_8799.n107 gnd 0.26985f
C4482 a_n6972_8799.n108 gnd 0.269982f
C4483 a_n6972_8799.t85 gnd 0.596495f
C4484 a_n6972_8799.n109 gnd 0.266246f
C4485 a_n6972_8799.t60 gnd 0.596495f
C4486 a_n6972_8799.n110 gnd 0.266496f
C4487 a_n6972_8799.n111 gnd 0.272062f
C4488 a_n6972_8799.t48 gnd 0.607324f
C4489 a_n6972_8799.t79 gnd 0.596495f
C4490 a_n6972_8799.n112 gnd 0.269967f
C4491 a_n6972_8799.t110 gnd 0.596495f
C4492 a_n6972_8799.t47 gnd 0.596495f
C4493 a_n6972_8799.n113 gnd 0.261131f
C4494 a_n6972_8799.t66 gnd 0.596495f
C4495 a_n6972_8799.n114 gnd 0.272496f
C4496 a_n6972_8799.t67 gnd 0.596495f
C4497 a_n6972_8799.t74 gnd 0.596495f
C4498 a_n6972_8799.n115 gnd 0.265926f
C4499 a_n6972_8799.t108 gnd 0.610514f
C4500 a_n6972_8799.t73 gnd 0.596495f
C4501 a_n6972_8799.n116 gnd 0.272062f
C4502 a_n6972_8799.n117 gnd 0.248651f
C4503 a_n6972_8799.t98 gnd 0.596495f
C4504 a_n6972_8799.n118 gnd 0.26985f
C4505 a_n6972_8799.n119 gnd 0.269982f
C4506 a_n6972_8799.t94 gnd 0.596495f
C4507 a_n6972_8799.n120 gnd 0.266246f
C4508 a_n6972_8799.t65 gnd 0.596495f
C4509 a_n6972_8799.n121 gnd 0.266496f
C4510 a_n6972_8799.n122 gnd 0.272062f
C4511 a_n6972_8799.t57 gnd 0.607324f
C4512 a_n6972_8799.n123 gnd 0.895502f
C4513 a_n6972_8799.t81 gnd 0.596495f
C4514 a_n6972_8799.n124 gnd 0.269967f
C4515 a_n6972_8799.t55 gnd 0.596495f
C4516 a_n6972_8799.t71 gnd 0.596495f
C4517 a_n6972_8799.n125 gnd 0.261131f
C4518 a_n6972_8799.t104 gnd 0.596495f
C4519 a_n6972_8799.n126 gnd 0.272496f
C4520 a_n6972_8799.t87 gnd 0.596495f
C4521 a_n6972_8799.t41 gnd 0.596495f
C4522 a_n6972_8799.n127 gnd 0.265926f
C4523 a_n6972_8799.t101 gnd 0.610514f
C4524 a_n6972_8799.t52 gnd 0.596495f
C4525 a_n6972_8799.n128 gnd 0.272062f
C4526 a_n6972_8799.n129 gnd 0.248651f
C4527 a_n6972_8799.t75 gnd 0.596495f
C4528 a_n6972_8799.n130 gnd 0.26985f
C4529 a_n6972_8799.n131 gnd 0.269982f
C4530 a_n6972_8799.t107 gnd 0.596495f
C4531 a_n6972_8799.n132 gnd 0.266246f
C4532 a_n6972_8799.t45 gnd 0.596495f
C4533 a_n6972_8799.n133 gnd 0.266496f
C4534 a_n6972_8799.n134 gnd 0.272062f
C4535 a_n6972_8799.t95 gnd 0.607324f
C4536 a_n6972_8799.n135 gnd 1.66315f
C4537 a_n6972_8799.t70 gnd 0.607324f
C4538 a_n6972_8799.t58 gnd 0.596495f
C4539 a_n6972_8799.t103 gnd 0.596495f
C4540 a_n6972_8799.t80 gnd 0.596495f
C4541 a_n6972_8799.n136 gnd 0.266496f
C4542 a_n6972_8799.t78 gnd 0.596495f
C4543 a_n6972_8799.t42 gnd 0.596495f
C4544 a_n6972_8799.t84 gnd 0.596495f
C4545 a_n6972_8799.n137 gnd 0.269982f
C4546 a_n6972_8799.t83 gnd 0.596495f
C4547 a_n6972_8799.t44 gnd 0.596495f
C4548 a_n6972_8799.t43 gnd 0.596495f
C4549 a_n6972_8799.n138 gnd 0.265926f
C4550 a_n6972_8799.t54 gnd 0.610514f
C4551 a_n6972_8799.t97 gnd 0.596495f
C4552 a_n6972_8799.n139 gnd 0.272062f
C4553 a_n6972_8799.n140 gnd 0.248651f
C4554 a_n6972_8799.n141 gnd 0.26985f
C4555 a_n6972_8799.n142 gnd 0.272496f
C4556 a_n6972_8799.n143 gnd 0.266246f
C4557 a_n6972_8799.n144 gnd 0.261131f
C4558 a_n6972_8799.n145 gnd 0.269967f
C4559 a_n6972_8799.n146 gnd 0.272062f
C4560 a_n6972_8799.t77 gnd 0.607324f
C4561 a_n6972_8799.t64 gnd 0.596495f
C4562 a_n6972_8799.t111 gnd 0.596495f
C4563 a_n6972_8799.t90 gnd 0.596495f
C4564 a_n6972_8799.n147 gnd 0.266496f
C4565 a_n6972_8799.t89 gnd 0.596495f
C4566 a_n6972_8799.t49 gnd 0.596495f
C4567 a_n6972_8799.t93 gnd 0.596495f
C4568 a_n6972_8799.n148 gnd 0.269982f
C4569 a_n6972_8799.t92 gnd 0.596495f
C4570 a_n6972_8799.t51 gnd 0.596495f
C4571 a_n6972_8799.t50 gnd 0.596495f
C4572 a_n6972_8799.n149 gnd 0.265926f
C4573 a_n6972_8799.t63 gnd 0.610514f
C4574 a_n6972_8799.t106 gnd 0.596495f
C4575 a_n6972_8799.n150 gnd 0.272062f
C4576 a_n6972_8799.n151 gnd 0.248651f
C4577 a_n6972_8799.n152 gnd 0.26985f
C4578 a_n6972_8799.n153 gnd 0.272496f
C4579 a_n6972_8799.n154 gnd 0.266246f
C4580 a_n6972_8799.n155 gnd 0.261131f
C4581 a_n6972_8799.n156 gnd 0.269967f
C4582 a_n6972_8799.n157 gnd 0.272062f
C4583 a_n6972_8799.n158 gnd 0.895502f
C4584 a_n6972_8799.t96 gnd 0.607324f
C4585 a_n6972_8799.t56 gnd 0.596495f
C4586 a_n6972_8799.t82 gnd 0.596495f
C4587 a_n6972_8799.t46 gnd 0.596495f
C4588 a_n6972_8799.n159 gnd 0.266496f
C4589 a_n6972_8799.t59 gnd 0.596495f
C4590 a_n6972_8799.t109 gnd 0.596495f
C4591 a_n6972_8799.t88 gnd 0.596495f
C4592 a_n6972_8799.n160 gnd 0.269982f
C4593 a_n6972_8799.t105 gnd 0.596495f
C4594 a_n6972_8799.t76 gnd 0.596495f
C4595 a_n6972_8799.t91 gnd 0.596495f
C4596 a_n6972_8799.n161 gnd 0.265926f
C4597 a_n6972_8799.t102 gnd 0.610514f
C4598 a_n6972_8799.t53 gnd 0.596495f
C4599 a_n6972_8799.n162 gnd 0.272062f
C4600 a_n6972_8799.n163 gnd 0.248651f
C4601 a_n6972_8799.n164 gnd 0.26985f
C4602 a_n6972_8799.n165 gnd 0.272496f
C4603 a_n6972_8799.n166 gnd 0.266246f
C4604 a_n6972_8799.n167 gnd 0.261131f
C4605 a_n6972_8799.n168 gnd 0.269967f
C4606 a_n6972_8799.n169 gnd 0.272062f
C4607 a_n6972_8799.n170 gnd 1.15468f
C4608 a_n6972_8799.n171 gnd 13.9136f
C4609 a_n6972_8799.n172 gnd 4.36548f
C4610 a_n6972_8799.n173 gnd 6.31987f
C4611 a_n6972_8799.t39 gnd 0.143856f
C4612 a_n6972_8799.t31 gnd 0.143856f
C4613 a_n6972_8799.n174 gnd 1.13461f
C4614 a_n6972_8799.t16 gnd 0.143856f
C4615 a_n6972_8799.t26 gnd 0.143856f
C4616 a_n6972_8799.n175 gnd 1.13274f
C4617 a_n6972_8799.t38 gnd 0.143856f
C4618 a_n6972_8799.t19 gnd 0.143856f
C4619 a_n6972_8799.n176 gnd 1.13274f
C4620 a_n6972_8799.n177 gnd 3.24672f
C4621 a_n6972_8799.n178 gnd 1.13275f
C4622 a_n6972_8799.t5 gnd 0.143856f
C4623 CSoutput.n0 gnd 0.040934f
C4624 CSoutput.t170 gnd 0.270772f
C4625 CSoutput.n1 gnd 0.122267f
C4626 CSoutput.n2 gnd 0.040934f
C4627 CSoutput.t168 gnd 0.270772f
C4628 CSoutput.n3 gnd 0.032444f
C4629 CSoutput.n4 gnd 0.040934f
C4630 CSoutput.t161 gnd 0.270772f
C4631 CSoutput.n5 gnd 0.027977f
C4632 CSoutput.n6 gnd 0.040934f
C4633 CSoutput.t165 gnd 0.270772f
C4634 CSoutput.t154 gnd 0.270772f
C4635 CSoutput.n7 gnd 0.120935f
C4636 CSoutput.n8 gnd 0.040934f
C4637 CSoutput.t153 gnd 0.270772f
C4638 CSoutput.n9 gnd 0.026674f
C4639 CSoutput.n10 gnd 0.040934f
C4640 CSoutput.t162 gnd 0.270772f
C4641 CSoutput.t167 gnd 0.270772f
C4642 CSoutput.n11 gnd 0.120935f
C4643 CSoutput.n12 gnd 0.040934f
C4644 CSoutput.t173 gnd 0.270772f
C4645 CSoutput.n13 gnd 0.027977f
C4646 CSoutput.n14 gnd 0.040934f
C4647 CSoutput.t155 gnd 0.270772f
C4648 CSoutput.t164 gnd 0.270772f
C4649 CSoutput.n15 gnd 0.120935f
C4650 CSoutput.n16 gnd 0.040934f
C4651 CSoutput.t171 gnd 0.270772f
C4652 CSoutput.n17 gnd 0.02988f
C4653 CSoutput.t158 gnd 0.32358f
C4654 CSoutput.t169 gnd 0.270772f
C4655 CSoutput.n18 gnd 0.154386f
C4656 CSoutput.n19 gnd 0.149808f
C4657 CSoutput.n20 gnd 0.173795f
C4658 CSoutput.n21 gnd 0.040934f
C4659 CSoutput.n22 gnd 0.034164f
C4660 CSoutput.n23 gnd 0.120935f
C4661 CSoutput.n24 gnd 0.032933f
C4662 CSoutput.n25 gnd 0.032444f
C4663 CSoutput.n26 gnd 0.040934f
C4664 CSoutput.n27 gnd 0.040934f
C4665 CSoutput.n28 gnd 0.033902f
C4666 CSoutput.n29 gnd 0.028783f
C4667 CSoutput.n30 gnd 0.123627f
C4668 CSoutput.n31 gnd 0.02918f
C4669 CSoutput.n32 gnd 0.040934f
C4670 CSoutput.n33 gnd 0.040934f
C4671 CSoutput.n34 gnd 0.040934f
C4672 CSoutput.n35 gnd 0.03354f
C4673 CSoutput.n36 gnd 0.120935f
C4674 CSoutput.n37 gnd 0.032077f
C4675 CSoutput.n38 gnd 0.0333f
C4676 CSoutput.n39 gnd 0.040934f
C4677 CSoutput.n40 gnd 0.040934f
C4678 CSoutput.n41 gnd 0.034157f
C4679 CSoutput.n42 gnd 0.03122f
C4680 CSoutput.n43 gnd 0.120935f
C4681 CSoutput.n44 gnd 0.032011f
C4682 CSoutput.n45 gnd 0.040934f
C4683 CSoutput.n46 gnd 0.040934f
C4684 CSoutput.n47 gnd 0.040934f
C4685 CSoutput.n48 gnd 0.032011f
C4686 CSoutput.n49 gnd 0.120935f
C4687 CSoutput.n50 gnd 0.03122f
C4688 CSoutput.n51 gnd 0.034157f
C4689 CSoutput.n52 gnd 0.040934f
C4690 CSoutput.n53 gnd 0.040934f
C4691 CSoutput.n54 gnd 0.0333f
C4692 CSoutput.n55 gnd 0.032077f
C4693 CSoutput.n56 gnd 0.120935f
C4694 CSoutput.n57 gnd 0.03354f
C4695 CSoutput.n58 gnd 0.040934f
C4696 CSoutput.n59 gnd 0.040934f
C4697 CSoutput.n60 gnd 0.040934f
C4698 CSoutput.n61 gnd 0.02918f
C4699 CSoutput.n62 gnd 0.123627f
C4700 CSoutput.n63 gnd 0.028783f
C4701 CSoutput.t157 gnd 0.270772f
C4702 CSoutput.n64 gnd 0.120935f
C4703 CSoutput.n65 gnd 0.033902f
C4704 CSoutput.n66 gnd 0.040934f
C4705 CSoutput.n67 gnd 0.040934f
C4706 CSoutput.n68 gnd 0.040934f
C4707 CSoutput.n69 gnd 0.032933f
C4708 CSoutput.n70 gnd 0.120935f
C4709 CSoutput.n71 gnd 0.034164f
C4710 CSoutput.n72 gnd 0.02988f
C4711 CSoutput.n73 gnd 0.040934f
C4712 CSoutput.n74 gnd 0.040934f
C4713 CSoutput.n75 gnd 0.030988f
C4714 CSoutput.n76 gnd 0.018404f
C4715 CSoutput.t160 gnd 0.304232f
C4716 CSoutput.n77 gnd 0.15113f
C4717 CSoutput.n78 gnd 0.646672f
C4718 CSoutput.t44 gnd 0.05106f
C4719 CSoutput.t33 gnd 0.05106f
C4720 CSoutput.n79 gnd 0.395322f
C4721 CSoutput.t21 gnd 0.05106f
C4722 CSoutput.t1 gnd 0.05106f
C4723 CSoutput.n80 gnd 0.394618f
C4724 CSoutput.n81 gnd 0.400536f
C4725 CSoutput.t30 gnd 0.05106f
C4726 CSoutput.t50 gnd 0.05106f
C4727 CSoutput.n82 gnd 0.394618f
C4728 CSoutput.n83 gnd 0.197367f
C4729 CSoutput.t18 gnd 0.05106f
C4730 CSoutput.t56 gnd 0.05106f
C4731 CSoutput.n84 gnd 0.394618f
C4732 CSoutput.n85 gnd 0.197367f
C4733 CSoutput.t24 gnd 0.05106f
C4734 CSoutput.t60 gnd 0.05106f
C4735 CSoutput.n86 gnd 0.394618f
C4736 CSoutput.n87 gnd 0.197367f
C4737 CSoutput.t57 gnd 0.05106f
C4738 CSoutput.t143 gnd 0.05106f
C4739 CSoutput.n88 gnd 0.394618f
C4740 CSoutput.n89 gnd 0.361926f
C4741 CSoutput.t55 gnd 0.05106f
C4742 CSoutput.t144 gnd 0.05106f
C4743 CSoutput.n90 gnd 0.395322f
C4744 CSoutput.t12 gnd 0.05106f
C4745 CSoutput.t19 gnd 0.05106f
C4746 CSoutput.n91 gnd 0.394618f
C4747 CSoutput.n92 gnd 0.400536f
C4748 CSoutput.t34 gnd 0.05106f
C4749 CSoutput.t45 gnd 0.05106f
C4750 CSoutput.n93 gnd 0.394618f
C4751 CSoutput.n94 gnd 0.197367f
C4752 CSoutput.t5 gnd 0.05106f
C4753 CSoutput.t28 gnd 0.05106f
C4754 CSoutput.n95 gnd 0.394618f
C4755 CSoutput.n96 gnd 0.197367f
C4756 CSoutput.t35 gnd 0.05106f
C4757 CSoutput.t27 gnd 0.05106f
C4758 CSoutput.n97 gnd 0.394618f
C4759 CSoutput.n98 gnd 0.197367f
C4760 CSoutput.t3 gnd 0.05106f
C4761 CSoutput.t31 gnd 0.05106f
C4762 CSoutput.n99 gnd 0.394618f
C4763 CSoutput.n100 gnd 0.294324f
C4764 CSoutput.n101 gnd 0.371141f
C4765 CSoutput.t9 gnd 0.05106f
C4766 CSoutput.t48 gnd 0.05106f
C4767 CSoutput.n102 gnd 0.395322f
C4768 CSoutput.t145 gnd 0.05106f
C4769 CSoutput.t51 gnd 0.05106f
C4770 CSoutput.n103 gnd 0.394618f
C4771 CSoutput.n104 gnd 0.400536f
C4772 CSoutput.t43 gnd 0.05106f
C4773 CSoutput.t150 gnd 0.05106f
C4774 CSoutput.n105 gnd 0.394618f
C4775 CSoutput.n106 gnd 0.197367f
C4776 CSoutput.t142 gnd 0.05106f
C4777 CSoutput.t20 gnd 0.05106f
C4778 CSoutput.n107 gnd 0.394618f
C4779 CSoutput.n108 gnd 0.197367f
C4780 CSoutput.t22 gnd 0.05106f
C4781 CSoutput.t151 gnd 0.05106f
C4782 CSoutput.n109 gnd 0.394618f
C4783 CSoutput.n110 gnd 0.197367f
C4784 CSoutput.t46 gnd 0.05106f
C4785 CSoutput.t146 gnd 0.05106f
C4786 CSoutput.n111 gnd 0.394618f
C4787 CSoutput.n112 gnd 0.294324f
C4788 CSoutput.n113 gnd 0.414841f
C4789 CSoutput.n114 gnd 8.1305f
C4790 CSoutput.n116 gnd 0.724122f
C4791 CSoutput.n117 gnd 0.543091f
C4792 CSoutput.n118 gnd 0.724122f
C4793 CSoutput.n119 gnd 0.724122f
C4794 CSoutput.n120 gnd 1.94956f
C4795 CSoutput.n121 gnd 0.724122f
C4796 CSoutput.n122 gnd 0.724122f
C4797 CSoutput.t163 gnd 0.905152f
C4798 CSoutput.n123 gnd 0.724122f
C4799 CSoutput.n124 gnd 0.724122f
C4800 CSoutput.n128 gnd 0.724122f
C4801 CSoutput.n132 gnd 0.724122f
C4802 CSoutput.n133 gnd 0.724122f
C4803 CSoutput.n135 gnd 0.724122f
C4804 CSoutput.n140 gnd 0.724122f
C4805 CSoutput.n142 gnd 0.724122f
C4806 CSoutput.n143 gnd 0.724122f
C4807 CSoutput.n145 gnd 0.724122f
C4808 CSoutput.n146 gnd 0.724122f
C4809 CSoutput.n148 gnd 0.724122f
C4810 CSoutput.t156 gnd 12.1f
C4811 CSoutput.n150 gnd 0.724122f
C4812 CSoutput.n151 gnd 0.543091f
C4813 CSoutput.n152 gnd 0.724122f
C4814 CSoutput.n153 gnd 0.724122f
C4815 CSoutput.n154 gnd 1.94956f
C4816 CSoutput.n155 gnd 0.724122f
C4817 CSoutput.n156 gnd 0.724122f
C4818 CSoutput.t172 gnd 0.905152f
C4819 CSoutput.n157 gnd 0.724122f
C4820 CSoutput.n158 gnd 0.724122f
C4821 CSoutput.n162 gnd 0.724122f
C4822 CSoutput.n166 gnd 0.724122f
C4823 CSoutput.n167 gnd 0.724122f
C4824 CSoutput.n169 gnd 0.724122f
C4825 CSoutput.n174 gnd 0.724122f
C4826 CSoutput.n176 gnd 0.724122f
C4827 CSoutput.n177 gnd 0.724122f
C4828 CSoutput.n179 gnd 0.724122f
C4829 CSoutput.n180 gnd 0.724122f
C4830 CSoutput.n182 gnd 0.724122f
C4831 CSoutput.n183 gnd 0.543091f
C4832 CSoutput.n185 gnd 0.724122f
C4833 CSoutput.n186 gnd 0.543091f
C4834 CSoutput.n187 gnd 0.724122f
C4835 CSoutput.n188 gnd 0.724122f
C4836 CSoutput.n189 gnd 1.94956f
C4837 CSoutput.n190 gnd 0.724122f
C4838 CSoutput.n191 gnd 0.724122f
C4839 CSoutput.t166 gnd 0.905152f
C4840 CSoutput.n192 gnd 0.724122f
C4841 CSoutput.n193 gnd 1.94956f
C4842 CSoutput.n195 gnd 0.724122f
C4843 CSoutput.n196 gnd 0.724122f
C4844 CSoutput.n198 gnd 0.724122f
C4845 CSoutput.n199 gnd 0.724122f
C4846 CSoutput.t152 gnd 11.9028f
C4847 CSoutput.t159 gnd 12.1f
C4848 CSoutput.n205 gnd 2.27168f
C4849 CSoutput.n206 gnd 9.253981f
C4850 CSoutput.n207 gnd 9.641211f
C4851 CSoutput.n212 gnd 2.46084f
C4852 CSoutput.n218 gnd 0.724122f
C4853 CSoutput.n220 gnd 0.724122f
C4854 CSoutput.n222 gnd 0.724122f
C4855 CSoutput.n224 gnd 0.724122f
C4856 CSoutput.n226 gnd 0.724122f
C4857 CSoutput.n232 gnd 0.724122f
C4858 CSoutput.n239 gnd 1.32848f
C4859 CSoutput.n240 gnd 1.32848f
C4860 CSoutput.n241 gnd 0.724122f
C4861 CSoutput.n242 gnd 0.724122f
C4862 CSoutput.n244 gnd 0.543091f
C4863 CSoutput.n245 gnd 0.465109f
C4864 CSoutput.n247 gnd 0.543091f
C4865 CSoutput.n248 gnd 0.465109f
C4866 CSoutput.n249 gnd 0.543091f
C4867 CSoutput.n251 gnd 0.724122f
C4868 CSoutput.n253 gnd 1.94956f
C4869 CSoutput.n254 gnd 2.27168f
C4870 CSoutput.n255 gnd 8.51128f
C4871 CSoutput.n257 gnd 0.543091f
C4872 CSoutput.n258 gnd 1.39741f
C4873 CSoutput.n259 gnd 0.543091f
C4874 CSoutput.n261 gnd 0.724122f
C4875 CSoutput.n263 gnd 1.94956f
C4876 CSoutput.n264 gnd 4.24645f
C4877 CSoutput.t40 gnd 0.05106f
C4878 CSoutput.t149 gnd 0.05106f
C4879 CSoutput.n265 gnd 0.395322f
C4880 CSoutput.t4 gnd 0.05106f
C4881 CSoutput.t10 gnd 0.05106f
C4882 CSoutput.n266 gnd 0.394618f
C4883 CSoutput.n267 gnd 0.400536f
C4884 CSoutput.t29 gnd 0.05106f
C4885 CSoutput.t148 gnd 0.05106f
C4886 CSoutput.n268 gnd 0.394618f
C4887 CSoutput.n269 gnd 0.197367f
C4888 CSoutput.t54 gnd 0.05106f
C4889 CSoutput.t23 gnd 0.05106f
C4890 CSoutput.n270 gnd 0.394618f
C4891 CSoutput.n271 gnd 0.197367f
C4892 CSoutput.t61 gnd 0.05106f
C4893 CSoutput.t25 gnd 0.05106f
C4894 CSoutput.n272 gnd 0.394618f
C4895 CSoutput.n273 gnd 0.197367f
C4896 CSoutput.t41 gnd 0.05106f
C4897 CSoutput.t38 gnd 0.05106f
C4898 CSoutput.n274 gnd 0.394618f
C4899 CSoutput.n275 gnd 0.361926f
C4900 CSoutput.t42 gnd 0.05106f
C4901 CSoutput.t36 gnd 0.05106f
C4902 CSoutput.n276 gnd 0.395322f
C4903 CSoutput.t147 gnd 0.05106f
C4904 CSoutput.t37 gnd 0.05106f
C4905 CSoutput.n277 gnd 0.394618f
C4906 CSoutput.n278 gnd 0.400536f
C4907 CSoutput.t49 gnd 0.05106f
C4908 CSoutput.t13 gnd 0.05106f
C4909 CSoutput.n279 gnd 0.394618f
C4910 CSoutput.n280 gnd 0.197367f
C4911 CSoutput.t26 gnd 0.05106f
C4912 CSoutput.t58 gnd 0.05106f
C4913 CSoutput.n281 gnd 0.394618f
C4914 CSoutput.n282 gnd 0.197367f
C4915 CSoutput.t15 gnd 0.05106f
C4916 CSoutput.t2 gnd 0.05106f
C4917 CSoutput.n283 gnd 0.394618f
C4918 CSoutput.n284 gnd 0.197367f
C4919 CSoutput.t6 gnd 0.05106f
C4920 CSoutput.t14 gnd 0.05106f
C4921 CSoutput.n285 gnd 0.394618f
C4922 CSoutput.n286 gnd 0.294324f
C4923 CSoutput.n287 gnd 0.371141f
C4924 CSoutput.t16 gnd 0.05106f
C4925 CSoutput.t11 gnd 0.05106f
C4926 CSoutput.n288 gnd 0.395322f
C4927 CSoutput.t7 gnd 0.05106f
C4928 CSoutput.t17 gnd 0.05106f
C4929 CSoutput.n289 gnd 0.394618f
C4930 CSoutput.n290 gnd 0.400536f
C4931 CSoutput.t53 gnd 0.05106f
C4932 CSoutput.t52 gnd 0.05106f
C4933 CSoutput.n291 gnd 0.394618f
C4934 CSoutput.n292 gnd 0.197367f
C4935 CSoutput.t59 gnd 0.05106f
C4936 CSoutput.t8 gnd 0.05106f
C4937 CSoutput.n293 gnd 0.394618f
C4938 CSoutput.n294 gnd 0.197367f
C4939 CSoutput.t0 gnd 0.05106f
C4940 CSoutput.t39 gnd 0.05106f
C4941 CSoutput.n295 gnd 0.394618f
C4942 CSoutput.n296 gnd 0.197367f
C4943 CSoutput.t32 gnd 0.05106f
C4944 CSoutput.t47 gnd 0.05106f
C4945 CSoutput.n297 gnd 0.394616f
C4946 CSoutput.n298 gnd 0.294326f
C4947 CSoutput.n299 gnd 0.414841f
C4948 CSoutput.n300 gnd 11.3858f
C4949 CSoutput.t122 gnd 0.044677f
C4950 CSoutput.t82 gnd 0.044677f
C4951 CSoutput.n301 gnd 0.396106f
C4952 CSoutput.t112 gnd 0.044677f
C4953 CSoutput.t114 gnd 0.044677f
C4954 CSoutput.n302 gnd 0.394785f
C4955 CSoutput.n303 gnd 0.367866f
C4956 CSoutput.t84 gnd 0.044677f
C4957 CSoutput.t93 gnd 0.044677f
C4958 CSoutput.n304 gnd 0.394785f
C4959 CSoutput.n305 gnd 0.18134f
C4960 CSoutput.t104 gnd 0.044677f
C4961 CSoutput.t123 gnd 0.044677f
C4962 CSoutput.n306 gnd 0.394785f
C4963 CSoutput.n307 gnd 0.18134f
C4964 CSoutput.t129 gnd 0.044677f
C4965 CSoutput.t64 gnd 0.044677f
C4966 CSoutput.n308 gnd 0.394785f
C4967 CSoutput.n309 gnd 0.18134f
C4968 CSoutput.t132 gnd 0.044677f
C4969 CSoutput.t136 gnd 0.044677f
C4970 CSoutput.n310 gnd 0.394785f
C4971 CSoutput.n311 gnd 0.18134f
C4972 CSoutput.t118 gnd 0.044677f
C4973 CSoutput.t79 gnd 0.044677f
C4974 CSoutput.n312 gnd 0.394785f
C4975 CSoutput.n313 gnd 0.18134f
C4976 CSoutput.t109 gnd 0.044677f
C4977 CSoutput.t128 gnd 0.044677f
C4978 CSoutput.n314 gnd 0.394785f
C4979 CSoutput.n315 gnd 0.18134f
C4980 CSoutput.t65 gnd 0.044677f
C4981 CSoutput.t99 gnd 0.044677f
C4982 CSoutput.n316 gnd 0.394785f
C4983 CSoutput.n317 gnd 0.18134f
C4984 CSoutput.t103 gnd 0.044677f
C4985 CSoutput.t120 gnd 0.044677f
C4986 CSoutput.n318 gnd 0.394785f
C4987 CSoutput.n319 gnd 0.334429f
C4988 CSoutput.t138 gnd 0.044677f
C4989 CSoutput.t119 gnd 0.044677f
C4990 CSoutput.n320 gnd 0.396106f
C4991 CSoutput.t105 gnd 0.044677f
C4992 CSoutput.t85 gnd 0.044677f
C4993 CSoutput.n321 gnd 0.394785f
C4994 CSoutput.n322 gnd 0.367866f
C4995 CSoutput.t130 gnd 0.044677f
C4996 CSoutput.t66 gnd 0.044677f
C4997 CSoutput.n323 gnd 0.394785f
C4998 CSoutput.n324 gnd 0.18134f
C4999 CSoutput.t73 gnd 0.044677f
C5000 CSoutput.t139 gnd 0.044677f
C5001 CSoutput.n325 gnd 0.394785f
C5002 CSoutput.n326 gnd 0.18134f
C5003 CSoutput.t108 gnd 0.044677f
C5004 CSoutput.t126 gnd 0.044677f
C5005 CSoutput.n327 gnd 0.394785f
C5006 CSoutput.n328 gnd 0.18134f
C5007 CSoutput.t110 gnd 0.044677f
C5008 CSoutput.t113 gnd 0.044677f
C5009 CSoutput.n329 gnd 0.394785f
C5010 CSoutput.n330 gnd 0.18134f
C5011 CSoutput.t135 gnd 0.044677f
C5012 CSoutput.t117 gnd 0.044677f
C5013 CSoutput.n331 gnd 0.394785f
C5014 CSoutput.n332 gnd 0.18134f
C5015 CSoutput.t102 gnd 0.044677f
C5016 CSoutput.t107 gnd 0.044677f
C5017 CSoutput.n333 gnd 0.394785f
C5018 CSoutput.n334 gnd 0.18134f
C5019 CSoutput.t127 gnd 0.044677f
C5020 CSoutput.t87 gnd 0.044677f
C5021 CSoutput.n335 gnd 0.394785f
C5022 CSoutput.n336 gnd 0.18134f
C5023 CSoutput.t72 gnd 0.044677f
C5024 CSoutput.t137 gnd 0.044677f
C5025 CSoutput.n337 gnd 0.394785f
C5026 CSoutput.n338 gnd 0.275314f
C5027 CSoutput.n339 gnd 0.511554f
C5028 CSoutput.n340 gnd 12.1413f
C5029 CSoutput.t71 gnd 0.044677f
C5030 CSoutput.t77 gnd 0.044677f
C5031 CSoutput.n341 gnd 0.396106f
C5032 CSoutput.t134 gnd 0.044677f
C5033 CSoutput.t100 gnd 0.044677f
C5034 CSoutput.n342 gnd 0.394785f
C5035 CSoutput.n343 gnd 0.367866f
C5036 CSoutput.t106 gnd 0.044677f
C5037 CSoutput.t92 gnd 0.044677f
C5038 CSoutput.n344 gnd 0.394785f
C5039 CSoutput.n345 gnd 0.18134f
C5040 CSoutput.t78 gnd 0.044677f
C5041 CSoutput.t88 gnd 0.044677f
C5042 CSoutput.n346 gnd 0.394785f
C5043 CSoutput.n347 gnd 0.18134f
C5044 CSoutput.t75 gnd 0.044677f
C5045 CSoutput.t83 gnd 0.044677f
C5046 CSoutput.n348 gnd 0.394785f
C5047 CSoutput.n349 gnd 0.18134f
C5048 CSoutput.t69 gnd 0.044677f
C5049 CSoutput.t141 gnd 0.044677f
C5050 CSoutput.n350 gnd 0.394785f
C5051 CSoutput.n351 gnd 0.18134f
C5052 CSoutput.t89 gnd 0.044677f
C5053 CSoutput.t96 gnd 0.044677f
C5054 CSoutput.n352 gnd 0.394785f
C5055 CSoutput.n353 gnd 0.18134f
C5056 CSoutput.t62 gnd 0.044677f
C5057 CSoutput.t125 gnd 0.044677f
C5058 CSoutput.n354 gnd 0.394785f
C5059 CSoutput.n355 gnd 0.18134f
C5060 CSoutput.t101 gnd 0.044677f
C5061 CSoutput.t76 gnd 0.044677f
C5062 CSoutput.n356 gnd 0.394785f
C5063 CSoutput.n357 gnd 0.18134f
C5064 CSoutput.t68 gnd 0.044677f
C5065 CSoutput.t115 gnd 0.044677f
C5066 CSoutput.n358 gnd 0.394785f
C5067 CSoutput.n359 gnd 0.334429f
C5068 CSoutput.t97 gnd 0.044677f
C5069 CSoutput.t70 gnd 0.044677f
C5070 CSoutput.n360 gnd 0.396106f
C5071 CSoutput.t111 gnd 0.044677f
C5072 CSoutput.t90 gnd 0.044677f
C5073 CSoutput.n361 gnd 0.394785f
C5074 CSoutput.n362 gnd 0.367866f
C5075 CSoutput.t91 gnd 0.044677f
C5076 CSoutput.t63 gnd 0.044677f
C5077 CSoutput.n363 gnd 0.394785f
C5078 CSoutput.n364 gnd 0.18134f
C5079 CSoutput.t116 gnd 0.044677f
C5080 CSoutput.t94 gnd 0.044677f
C5081 CSoutput.n365 gnd 0.394785f
C5082 CSoutput.n366 gnd 0.18134f
C5083 CSoutput.t80 gnd 0.044677f
C5084 CSoutput.t124 gnd 0.044677f
C5085 CSoutput.n367 gnd 0.394785f
C5086 CSoutput.n368 gnd 0.18134f
C5087 CSoutput.t133 gnd 0.044677f
C5088 CSoutput.t98 gnd 0.044677f
C5089 CSoutput.n369 gnd 0.394785f
C5090 CSoutput.n370 gnd 0.18134f
C5091 CSoutput.t95 gnd 0.044677f
C5092 CSoutput.t67 gnd 0.044677f
C5093 CSoutput.n371 gnd 0.394785f
C5094 CSoutput.n372 gnd 0.18134f
C5095 CSoutput.t121 gnd 0.044677f
C5096 CSoutput.t140 gnd 0.044677f
C5097 CSoutput.n373 gnd 0.394785f
C5098 CSoutput.n374 gnd 0.18134f
C5099 CSoutput.t74 gnd 0.044677f
C5100 CSoutput.t81 gnd 0.044677f
C5101 CSoutput.n375 gnd 0.394785f
C5102 CSoutput.n376 gnd 0.18134f
C5103 CSoutput.t131 gnd 0.044677f
C5104 CSoutput.t86 gnd 0.044677f
C5105 CSoutput.n377 gnd 0.394785f
C5106 CSoutput.n378 gnd 0.275314f
C5107 CSoutput.n379 gnd 0.511554f
C5108 CSoutput.n380 gnd 7.1925f
C5109 CSoutput.n381 gnd 13.316401f
C5110 commonsourceibias.n0 gnd 0.010705f
C5111 commonsourceibias.t117 gnd 0.162096f
C5112 commonsourceibias.t135 gnd 0.149881f
C5113 commonsourceibias.n1 gnd 0.007808f
C5114 commonsourceibias.n2 gnd 0.008022f
C5115 commonsourceibias.t92 gnd 0.149881f
C5116 commonsourceibias.n3 gnd 0.010321f
C5117 commonsourceibias.n4 gnd 0.008022f
C5118 commonsourceibias.t90 gnd 0.149881f
C5119 commonsourceibias.n5 gnd 0.059802f
C5120 commonsourceibias.t127 gnd 0.149881f
C5121 commonsourceibias.n6 gnd 0.007564f
C5122 commonsourceibias.n7 gnd 0.008022f
C5123 commonsourceibias.t145 gnd 0.149881f
C5124 commonsourceibias.n8 gnd 0.010168f
C5125 commonsourceibias.n9 gnd 0.008022f
C5126 commonsourceibias.t83 gnd 0.149881f
C5127 commonsourceibias.n10 gnd 0.059802f
C5128 commonsourceibias.t116 gnd 0.149881f
C5129 commonsourceibias.n11 gnd 0.007348f
C5130 commonsourceibias.n12 gnd 0.008022f
C5131 commonsourceibias.t110 gnd 0.149881f
C5132 commonsourceibias.n13 gnd 0.009997f
C5133 commonsourceibias.n14 gnd 0.010705f
C5134 commonsourceibias.t76 gnd 0.162096f
C5135 commonsourceibias.t24 gnd 0.149881f
C5136 commonsourceibias.n15 gnd 0.007808f
C5137 commonsourceibias.n16 gnd 0.008022f
C5138 commonsourceibias.t64 gnd 0.149881f
C5139 commonsourceibias.n17 gnd 0.010321f
C5140 commonsourceibias.n18 gnd 0.008022f
C5141 commonsourceibias.t74 gnd 0.149881f
C5142 commonsourceibias.n19 gnd 0.059802f
C5143 commonsourceibias.t4 gnd 0.149881f
C5144 commonsourceibias.n20 gnd 0.007564f
C5145 commonsourceibias.n21 gnd 0.008022f
C5146 commonsourceibias.t48 gnd 0.149881f
C5147 commonsourceibias.n22 gnd 0.010168f
C5148 commonsourceibias.n23 gnd 0.008022f
C5149 commonsourceibias.t44 gnd 0.149881f
C5150 commonsourceibias.n24 gnd 0.059802f
C5151 commonsourceibias.t70 gnd 0.149881f
C5152 commonsourceibias.n25 gnd 0.007348f
C5153 commonsourceibias.n26 gnd 0.008022f
C5154 commonsourceibias.t78 gnd 0.149881f
C5155 commonsourceibias.n27 gnd 0.009997f
C5156 commonsourceibias.n28 gnd 0.008022f
C5157 commonsourceibias.t8 gnd 0.149881f
C5158 commonsourceibias.n29 gnd 0.059802f
C5159 commonsourceibias.t40 gnd 0.149881f
C5160 commonsourceibias.n30 gnd 0.007159f
C5161 commonsourceibias.n31 gnd 0.008022f
C5162 commonsourceibias.t46 gnd 0.149881f
C5163 commonsourceibias.n32 gnd 0.009806f
C5164 commonsourceibias.n33 gnd 0.008022f
C5165 commonsourceibias.t0 gnd 0.149881f
C5166 commonsourceibias.n34 gnd 0.059802f
C5167 commonsourceibias.t50 gnd 0.149881f
C5168 commonsourceibias.n35 gnd 0.006995f
C5169 commonsourceibias.n36 gnd 0.008022f
C5170 commonsourceibias.t26 gnd 0.149881f
C5171 commonsourceibias.n37 gnd 0.009595f
C5172 commonsourceibias.n38 gnd 0.008022f
C5173 commonsourceibias.t60 gnd 0.149881f
C5174 commonsourceibias.n39 gnd 0.059802f
C5175 commonsourceibias.t34 gnd 0.149881f
C5176 commonsourceibias.n40 gnd 0.006855f
C5177 commonsourceibias.n41 gnd 0.008022f
C5178 commonsourceibias.t22 gnd 0.149881f
C5179 commonsourceibias.n42 gnd 0.00936f
C5180 commonsourceibias.t54 gnd 0.16664f
C5181 commonsourceibias.t12 gnd 0.149881f
C5182 commonsourceibias.n43 gnd 0.065328f
C5183 commonsourceibias.n44 gnd 0.07169f
C5184 commonsourceibias.n45 gnd 0.033265f
C5185 commonsourceibias.n46 gnd 0.008022f
C5186 commonsourceibias.n47 gnd 0.007808f
C5187 commonsourceibias.n48 gnd 0.01119f
C5188 commonsourceibias.n49 gnd 0.059802f
C5189 commonsourceibias.n50 gnd 0.011182f
C5190 commonsourceibias.n51 gnd 0.008022f
C5191 commonsourceibias.n52 gnd 0.008022f
C5192 commonsourceibias.n53 gnd 0.008022f
C5193 commonsourceibias.n54 gnd 0.010321f
C5194 commonsourceibias.n55 gnd 0.059802f
C5195 commonsourceibias.n56 gnd 0.010563f
C5196 commonsourceibias.n57 gnd 0.010263f
C5197 commonsourceibias.n58 gnd 0.008022f
C5198 commonsourceibias.n59 gnd 0.008022f
C5199 commonsourceibias.n60 gnd 0.008022f
C5200 commonsourceibias.n61 gnd 0.007564f
C5201 commonsourceibias.n62 gnd 0.0112f
C5202 commonsourceibias.n63 gnd 0.059802f
C5203 commonsourceibias.n64 gnd 0.011196f
C5204 commonsourceibias.n65 gnd 0.008022f
C5205 commonsourceibias.n66 gnd 0.008022f
C5206 commonsourceibias.n67 gnd 0.008022f
C5207 commonsourceibias.n68 gnd 0.010168f
C5208 commonsourceibias.n69 gnd 0.059802f
C5209 commonsourceibias.n70 gnd 0.010488f
C5210 commonsourceibias.n71 gnd 0.010338f
C5211 commonsourceibias.n72 gnd 0.008022f
C5212 commonsourceibias.n73 gnd 0.008022f
C5213 commonsourceibias.n74 gnd 0.008022f
C5214 commonsourceibias.n75 gnd 0.007348f
C5215 commonsourceibias.n76 gnd 0.011204f
C5216 commonsourceibias.n77 gnd 0.059802f
C5217 commonsourceibias.n78 gnd 0.011203f
C5218 commonsourceibias.n79 gnd 0.008022f
C5219 commonsourceibias.n80 gnd 0.008022f
C5220 commonsourceibias.n81 gnd 0.008022f
C5221 commonsourceibias.n82 gnd 0.009997f
C5222 commonsourceibias.n83 gnd 0.059802f
C5223 commonsourceibias.n84 gnd 0.010413f
C5224 commonsourceibias.n85 gnd 0.010413f
C5225 commonsourceibias.n86 gnd 0.008022f
C5226 commonsourceibias.n87 gnd 0.008022f
C5227 commonsourceibias.n88 gnd 0.008022f
C5228 commonsourceibias.n89 gnd 0.007159f
C5229 commonsourceibias.n90 gnd 0.011203f
C5230 commonsourceibias.n91 gnd 0.059802f
C5231 commonsourceibias.n92 gnd 0.011204f
C5232 commonsourceibias.n93 gnd 0.008022f
C5233 commonsourceibias.n94 gnd 0.008022f
C5234 commonsourceibias.n95 gnd 0.008022f
C5235 commonsourceibias.n96 gnd 0.009806f
C5236 commonsourceibias.n97 gnd 0.059802f
C5237 commonsourceibias.n98 gnd 0.010338f
C5238 commonsourceibias.n99 gnd 0.010488f
C5239 commonsourceibias.n100 gnd 0.008022f
C5240 commonsourceibias.n101 gnd 0.008022f
C5241 commonsourceibias.n102 gnd 0.008022f
C5242 commonsourceibias.n103 gnd 0.006995f
C5243 commonsourceibias.n104 gnd 0.011196f
C5244 commonsourceibias.n105 gnd 0.059802f
C5245 commonsourceibias.n106 gnd 0.0112f
C5246 commonsourceibias.n107 gnd 0.008022f
C5247 commonsourceibias.n108 gnd 0.008022f
C5248 commonsourceibias.n109 gnd 0.008022f
C5249 commonsourceibias.n110 gnd 0.009595f
C5250 commonsourceibias.n111 gnd 0.059802f
C5251 commonsourceibias.n112 gnd 0.010263f
C5252 commonsourceibias.n113 gnd 0.010563f
C5253 commonsourceibias.n114 gnd 0.008022f
C5254 commonsourceibias.n115 gnd 0.008022f
C5255 commonsourceibias.n116 gnd 0.008022f
C5256 commonsourceibias.n117 gnd 0.006855f
C5257 commonsourceibias.n118 gnd 0.011182f
C5258 commonsourceibias.n119 gnd 0.059802f
C5259 commonsourceibias.n120 gnd 0.01119f
C5260 commonsourceibias.n121 gnd 0.008022f
C5261 commonsourceibias.n122 gnd 0.008022f
C5262 commonsourceibias.n123 gnd 0.008022f
C5263 commonsourceibias.n124 gnd 0.00936f
C5264 commonsourceibias.n125 gnd 0.059802f
C5265 commonsourceibias.n126 gnd 0.009843f
C5266 commonsourceibias.n127 gnd 0.071758f
C5267 commonsourceibias.n128 gnd 0.079928f
C5268 commonsourceibias.t77 gnd 0.017311f
C5269 commonsourceibias.t25 gnd 0.017311f
C5270 commonsourceibias.n129 gnd 0.152968f
C5271 commonsourceibias.n130 gnd 0.132319f
C5272 commonsourceibias.t65 gnd 0.017311f
C5273 commonsourceibias.t75 gnd 0.017311f
C5274 commonsourceibias.n131 gnd 0.152968f
C5275 commonsourceibias.n132 gnd 0.070264f
C5276 commonsourceibias.t5 gnd 0.017311f
C5277 commonsourceibias.t49 gnd 0.017311f
C5278 commonsourceibias.n133 gnd 0.152968f
C5279 commonsourceibias.n134 gnd 0.070264f
C5280 commonsourceibias.t45 gnd 0.017311f
C5281 commonsourceibias.t71 gnd 0.017311f
C5282 commonsourceibias.n135 gnd 0.152968f
C5283 commonsourceibias.n136 gnd 0.070264f
C5284 commonsourceibias.t79 gnd 0.017311f
C5285 commonsourceibias.t9 gnd 0.017311f
C5286 commonsourceibias.n137 gnd 0.152968f
C5287 commonsourceibias.n138 gnd 0.058702f
C5288 commonsourceibias.t13 gnd 0.017311f
C5289 commonsourceibias.t55 gnd 0.017311f
C5290 commonsourceibias.n139 gnd 0.15348f
C5291 commonsourceibias.t35 gnd 0.017311f
C5292 commonsourceibias.t23 gnd 0.017311f
C5293 commonsourceibias.n140 gnd 0.152968f
C5294 commonsourceibias.n141 gnd 0.142538f
C5295 commonsourceibias.t27 gnd 0.017311f
C5296 commonsourceibias.t61 gnd 0.017311f
C5297 commonsourceibias.n142 gnd 0.152968f
C5298 commonsourceibias.n143 gnd 0.070264f
C5299 commonsourceibias.t1 gnd 0.017311f
C5300 commonsourceibias.t51 gnd 0.017311f
C5301 commonsourceibias.n144 gnd 0.152968f
C5302 commonsourceibias.n145 gnd 0.070264f
C5303 commonsourceibias.t41 gnd 0.017311f
C5304 commonsourceibias.t47 gnd 0.017311f
C5305 commonsourceibias.n146 gnd 0.152968f
C5306 commonsourceibias.n147 gnd 0.058702f
C5307 commonsourceibias.n148 gnd 0.071082f
C5308 commonsourceibias.n149 gnd 0.05192f
C5309 commonsourceibias.t131 gnd 0.149881f
C5310 commonsourceibias.n150 gnd 0.059802f
C5311 commonsourceibias.t107 gnd 0.149881f
C5312 commonsourceibias.n151 gnd 0.059802f
C5313 commonsourceibias.n152 gnd 0.008022f
C5314 commonsourceibias.t103 gnd 0.149881f
C5315 commonsourceibias.n153 gnd 0.059802f
C5316 commonsourceibias.n154 gnd 0.008022f
C5317 commonsourceibias.t121 gnd 0.149881f
C5318 commonsourceibias.n155 gnd 0.059802f
C5319 commonsourceibias.n156 gnd 0.008022f
C5320 commonsourceibias.t138 gnd 0.149881f
C5321 commonsourceibias.n157 gnd 0.006995f
C5322 commonsourceibias.n158 gnd 0.008022f
C5323 commonsourceibias.t95 gnd 0.149881f
C5324 commonsourceibias.n159 gnd 0.009595f
C5325 commonsourceibias.n160 gnd 0.008022f
C5326 commonsourceibias.t111 gnd 0.149881f
C5327 commonsourceibias.n161 gnd 0.059802f
C5328 commonsourceibias.t130 gnd 0.149881f
C5329 commonsourceibias.n162 gnd 0.006855f
C5330 commonsourceibias.n163 gnd 0.008022f
C5331 commonsourceibias.t87 gnd 0.149881f
C5332 commonsourceibias.n164 gnd 0.00936f
C5333 commonsourceibias.t119 gnd 0.16664f
C5334 commonsourceibias.t84 gnd 0.149881f
C5335 commonsourceibias.n165 gnd 0.065328f
C5336 commonsourceibias.n166 gnd 0.07169f
C5337 commonsourceibias.n167 gnd 0.033265f
C5338 commonsourceibias.n168 gnd 0.008022f
C5339 commonsourceibias.n169 gnd 0.007808f
C5340 commonsourceibias.n170 gnd 0.01119f
C5341 commonsourceibias.n171 gnd 0.059802f
C5342 commonsourceibias.n172 gnd 0.011182f
C5343 commonsourceibias.n173 gnd 0.008022f
C5344 commonsourceibias.n174 gnd 0.008022f
C5345 commonsourceibias.n175 gnd 0.008022f
C5346 commonsourceibias.n176 gnd 0.010321f
C5347 commonsourceibias.n177 gnd 0.059802f
C5348 commonsourceibias.n178 gnd 0.010563f
C5349 commonsourceibias.n179 gnd 0.010263f
C5350 commonsourceibias.n180 gnd 0.008022f
C5351 commonsourceibias.n181 gnd 0.008022f
C5352 commonsourceibias.n182 gnd 0.008022f
C5353 commonsourceibias.n183 gnd 0.007564f
C5354 commonsourceibias.n184 gnd 0.0112f
C5355 commonsourceibias.n185 gnd 0.059802f
C5356 commonsourceibias.n186 gnd 0.011196f
C5357 commonsourceibias.n187 gnd 0.008022f
C5358 commonsourceibias.n188 gnd 0.008022f
C5359 commonsourceibias.n189 gnd 0.008022f
C5360 commonsourceibias.n190 gnd 0.010168f
C5361 commonsourceibias.n191 gnd 0.059802f
C5362 commonsourceibias.n192 gnd 0.010488f
C5363 commonsourceibias.n193 gnd 0.010338f
C5364 commonsourceibias.n194 gnd 0.008022f
C5365 commonsourceibias.n195 gnd 0.008022f
C5366 commonsourceibias.n196 gnd 0.009806f
C5367 commonsourceibias.n197 gnd 0.007348f
C5368 commonsourceibias.n198 gnd 0.011204f
C5369 commonsourceibias.n199 gnd 0.008022f
C5370 commonsourceibias.n200 gnd 0.008022f
C5371 commonsourceibias.n201 gnd 0.011203f
C5372 commonsourceibias.n202 gnd 0.007159f
C5373 commonsourceibias.n203 gnd 0.009997f
C5374 commonsourceibias.n204 gnd 0.008022f
C5375 commonsourceibias.n205 gnd 0.007008f
C5376 commonsourceibias.n206 gnd 0.010413f
C5377 commonsourceibias.n207 gnd 0.010413f
C5378 commonsourceibias.n208 gnd 0.007008f
C5379 commonsourceibias.n209 gnd 0.008022f
C5380 commonsourceibias.n210 gnd 0.008022f
C5381 commonsourceibias.n211 gnd 0.007159f
C5382 commonsourceibias.n212 gnd 0.011203f
C5383 commonsourceibias.n213 gnd 0.059802f
C5384 commonsourceibias.n214 gnd 0.011204f
C5385 commonsourceibias.n215 gnd 0.008022f
C5386 commonsourceibias.n216 gnd 0.008022f
C5387 commonsourceibias.n217 gnd 0.008022f
C5388 commonsourceibias.n218 gnd 0.009806f
C5389 commonsourceibias.n219 gnd 0.059802f
C5390 commonsourceibias.n220 gnd 0.010338f
C5391 commonsourceibias.n221 gnd 0.010488f
C5392 commonsourceibias.n222 gnd 0.008022f
C5393 commonsourceibias.n223 gnd 0.008022f
C5394 commonsourceibias.n224 gnd 0.008022f
C5395 commonsourceibias.n225 gnd 0.006995f
C5396 commonsourceibias.n226 gnd 0.011196f
C5397 commonsourceibias.n227 gnd 0.059802f
C5398 commonsourceibias.n228 gnd 0.0112f
C5399 commonsourceibias.n229 gnd 0.008022f
C5400 commonsourceibias.n230 gnd 0.008022f
C5401 commonsourceibias.n231 gnd 0.008022f
C5402 commonsourceibias.n232 gnd 0.009595f
C5403 commonsourceibias.n233 gnd 0.059802f
C5404 commonsourceibias.n234 gnd 0.010263f
C5405 commonsourceibias.n235 gnd 0.010563f
C5406 commonsourceibias.n236 gnd 0.008022f
C5407 commonsourceibias.n237 gnd 0.008022f
C5408 commonsourceibias.n238 gnd 0.008022f
C5409 commonsourceibias.n239 gnd 0.006855f
C5410 commonsourceibias.n240 gnd 0.011182f
C5411 commonsourceibias.n241 gnd 0.059802f
C5412 commonsourceibias.n242 gnd 0.01119f
C5413 commonsourceibias.n243 gnd 0.008022f
C5414 commonsourceibias.n244 gnd 0.008022f
C5415 commonsourceibias.n245 gnd 0.008022f
C5416 commonsourceibias.n246 gnd 0.00936f
C5417 commonsourceibias.n247 gnd 0.059802f
C5418 commonsourceibias.n248 gnd 0.009843f
C5419 commonsourceibias.n249 gnd 0.071758f
C5420 commonsourceibias.n250 gnd 0.046883f
C5421 commonsourceibias.n251 gnd 0.010705f
C5422 commonsourceibias.t120 gnd 0.149881f
C5423 commonsourceibias.n252 gnd 0.007808f
C5424 commonsourceibias.n253 gnd 0.008022f
C5425 commonsourceibias.t81 gnd 0.149881f
C5426 commonsourceibias.n254 gnd 0.010321f
C5427 commonsourceibias.n255 gnd 0.008022f
C5428 commonsourceibias.t159 gnd 0.149881f
C5429 commonsourceibias.n256 gnd 0.059802f
C5430 commonsourceibias.t109 gnd 0.149881f
C5431 commonsourceibias.n257 gnd 0.007564f
C5432 commonsourceibias.n258 gnd 0.008022f
C5433 commonsourceibias.t129 gnd 0.149881f
C5434 commonsourceibias.n259 gnd 0.010168f
C5435 commonsourceibias.n260 gnd 0.008022f
C5436 commonsourceibias.t151 gnd 0.149881f
C5437 commonsourceibias.n261 gnd 0.059802f
C5438 commonsourceibias.t100 gnd 0.149881f
C5439 commonsourceibias.n262 gnd 0.007348f
C5440 commonsourceibias.n263 gnd 0.008022f
C5441 commonsourceibias.t96 gnd 0.149881f
C5442 commonsourceibias.n264 gnd 0.009997f
C5443 commonsourceibias.n265 gnd 0.008022f
C5444 commonsourceibias.t113 gnd 0.149881f
C5445 commonsourceibias.n266 gnd 0.059802f
C5446 commonsourceibias.t94 gnd 0.149881f
C5447 commonsourceibias.n267 gnd 0.007159f
C5448 commonsourceibias.n268 gnd 0.008022f
C5449 commonsourceibias.t91 gnd 0.149881f
C5450 commonsourceibias.n269 gnd 0.009806f
C5451 commonsourceibias.n270 gnd 0.008022f
C5452 commonsourceibias.t104 gnd 0.149881f
C5453 commonsourceibias.n271 gnd 0.059802f
C5454 commonsourceibias.t122 gnd 0.149881f
C5455 commonsourceibias.n272 gnd 0.006995f
C5456 commonsourceibias.n273 gnd 0.008022f
C5457 commonsourceibias.t85 gnd 0.149881f
C5458 commonsourceibias.n274 gnd 0.009595f
C5459 commonsourceibias.n275 gnd 0.008022f
C5460 commonsourceibias.t97 gnd 0.149881f
C5461 commonsourceibias.n276 gnd 0.059802f
C5462 commonsourceibias.t112 gnd 0.149881f
C5463 commonsourceibias.n277 gnd 0.006855f
C5464 commonsourceibias.n278 gnd 0.008022f
C5465 commonsourceibias.t157 gnd 0.149881f
C5466 commonsourceibias.n279 gnd 0.00936f
C5467 commonsourceibias.t102 gnd 0.16664f
C5468 commonsourceibias.t152 gnd 0.149881f
C5469 commonsourceibias.n280 gnd 0.065328f
C5470 commonsourceibias.n281 gnd 0.07169f
C5471 commonsourceibias.n282 gnd 0.033265f
C5472 commonsourceibias.n283 gnd 0.008022f
C5473 commonsourceibias.n284 gnd 0.007808f
C5474 commonsourceibias.n285 gnd 0.01119f
C5475 commonsourceibias.n286 gnd 0.059802f
C5476 commonsourceibias.n287 gnd 0.011182f
C5477 commonsourceibias.n288 gnd 0.008022f
C5478 commonsourceibias.n289 gnd 0.008022f
C5479 commonsourceibias.n290 gnd 0.008022f
C5480 commonsourceibias.n291 gnd 0.010321f
C5481 commonsourceibias.n292 gnd 0.059802f
C5482 commonsourceibias.n293 gnd 0.010563f
C5483 commonsourceibias.n294 gnd 0.010263f
C5484 commonsourceibias.n295 gnd 0.008022f
C5485 commonsourceibias.n296 gnd 0.008022f
C5486 commonsourceibias.n297 gnd 0.008022f
C5487 commonsourceibias.n298 gnd 0.007564f
C5488 commonsourceibias.n299 gnd 0.0112f
C5489 commonsourceibias.n300 gnd 0.059802f
C5490 commonsourceibias.n301 gnd 0.011196f
C5491 commonsourceibias.n302 gnd 0.008022f
C5492 commonsourceibias.n303 gnd 0.008022f
C5493 commonsourceibias.n304 gnd 0.008022f
C5494 commonsourceibias.n305 gnd 0.010168f
C5495 commonsourceibias.n306 gnd 0.059802f
C5496 commonsourceibias.n307 gnd 0.010488f
C5497 commonsourceibias.n308 gnd 0.010338f
C5498 commonsourceibias.n309 gnd 0.008022f
C5499 commonsourceibias.n310 gnd 0.008022f
C5500 commonsourceibias.n311 gnd 0.008022f
C5501 commonsourceibias.n312 gnd 0.007348f
C5502 commonsourceibias.n313 gnd 0.011204f
C5503 commonsourceibias.n314 gnd 0.059802f
C5504 commonsourceibias.n315 gnd 0.011203f
C5505 commonsourceibias.n316 gnd 0.008022f
C5506 commonsourceibias.n317 gnd 0.008022f
C5507 commonsourceibias.n318 gnd 0.008022f
C5508 commonsourceibias.n319 gnd 0.009997f
C5509 commonsourceibias.n320 gnd 0.059802f
C5510 commonsourceibias.n321 gnd 0.010413f
C5511 commonsourceibias.n322 gnd 0.010413f
C5512 commonsourceibias.n323 gnd 0.008022f
C5513 commonsourceibias.n324 gnd 0.008022f
C5514 commonsourceibias.n325 gnd 0.008022f
C5515 commonsourceibias.n326 gnd 0.007159f
C5516 commonsourceibias.n327 gnd 0.011203f
C5517 commonsourceibias.n328 gnd 0.059802f
C5518 commonsourceibias.n329 gnd 0.011204f
C5519 commonsourceibias.n330 gnd 0.008022f
C5520 commonsourceibias.n331 gnd 0.008022f
C5521 commonsourceibias.n332 gnd 0.008022f
C5522 commonsourceibias.n333 gnd 0.009806f
C5523 commonsourceibias.n334 gnd 0.059802f
C5524 commonsourceibias.n335 gnd 0.010338f
C5525 commonsourceibias.n336 gnd 0.010488f
C5526 commonsourceibias.n337 gnd 0.008022f
C5527 commonsourceibias.n338 gnd 0.008022f
C5528 commonsourceibias.n339 gnd 0.008022f
C5529 commonsourceibias.n340 gnd 0.006995f
C5530 commonsourceibias.n341 gnd 0.011196f
C5531 commonsourceibias.n342 gnd 0.059802f
C5532 commonsourceibias.n343 gnd 0.0112f
C5533 commonsourceibias.n344 gnd 0.008022f
C5534 commonsourceibias.n345 gnd 0.008022f
C5535 commonsourceibias.n346 gnd 0.008022f
C5536 commonsourceibias.n347 gnd 0.009595f
C5537 commonsourceibias.n348 gnd 0.059802f
C5538 commonsourceibias.n349 gnd 0.010263f
C5539 commonsourceibias.n350 gnd 0.010563f
C5540 commonsourceibias.n351 gnd 0.008022f
C5541 commonsourceibias.n352 gnd 0.008022f
C5542 commonsourceibias.n353 gnd 0.008022f
C5543 commonsourceibias.n354 gnd 0.006855f
C5544 commonsourceibias.n355 gnd 0.011182f
C5545 commonsourceibias.n356 gnd 0.059802f
C5546 commonsourceibias.n357 gnd 0.01119f
C5547 commonsourceibias.n358 gnd 0.008022f
C5548 commonsourceibias.n359 gnd 0.008022f
C5549 commonsourceibias.n360 gnd 0.008022f
C5550 commonsourceibias.n361 gnd 0.00936f
C5551 commonsourceibias.n362 gnd 0.059802f
C5552 commonsourceibias.n363 gnd 0.009843f
C5553 commonsourceibias.t101 gnd 0.162096f
C5554 commonsourceibias.n364 gnd 0.071758f
C5555 commonsourceibias.n365 gnd 0.024957f
C5556 commonsourceibias.n366 gnd 0.404135f
C5557 commonsourceibias.n367 gnd 0.010705f
C5558 commonsourceibias.t140 gnd 0.162096f
C5559 commonsourceibias.t153 gnd 0.149881f
C5560 commonsourceibias.n368 gnd 0.007808f
C5561 commonsourceibias.n369 gnd 0.008022f
C5562 commonsourceibias.t86 gnd 0.149881f
C5563 commonsourceibias.n370 gnd 0.010321f
C5564 commonsourceibias.n371 gnd 0.008022f
C5565 commonsourceibias.t146 gnd 0.149881f
C5566 commonsourceibias.n372 gnd 0.007564f
C5567 commonsourceibias.n373 gnd 0.008022f
C5568 commonsourceibias.t80 gnd 0.149881f
C5569 commonsourceibias.n374 gnd 0.010168f
C5570 commonsourceibias.n375 gnd 0.008022f
C5571 commonsourceibias.t139 gnd 0.149881f
C5572 commonsourceibias.n376 gnd 0.007348f
C5573 commonsourceibias.n377 gnd 0.008022f
C5574 commonsourceibias.t133 gnd 0.149881f
C5575 commonsourceibias.n378 gnd 0.009997f
C5576 commonsourceibias.t17 gnd 0.017311f
C5577 commonsourceibias.t69 gnd 0.017311f
C5578 commonsourceibias.n379 gnd 0.15348f
C5579 commonsourceibias.t67 gnd 0.017311f
C5580 commonsourceibias.t15 gnd 0.017311f
C5581 commonsourceibias.n380 gnd 0.152968f
C5582 commonsourceibias.n381 gnd 0.142538f
C5583 commonsourceibias.t57 gnd 0.017311f
C5584 commonsourceibias.t59 gnd 0.017311f
C5585 commonsourceibias.n382 gnd 0.152968f
C5586 commonsourceibias.n383 gnd 0.070264f
C5587 commonsourceibias.t19 gnd 0.017311f
C5588 commonsourceibias.t63 gnd 0.017311f
C5589 commonsourceibias.n384 gnd 0.152968f
C5590 commonsourceibias.n385 gnd 0.070264f
C5591 commonsourceibias.t29 gnd 0.017311f
C5592 commonsourceibias.t21 gnd 0.017311f
C5593 commonsourceibias.n386 gnd 0.152968f
C5594 commonsourceibias.n387 gnd 0.058702f
C5595 commonsourceibias.n388 gnd 0.010705f
C5596 commonsourceibias.t6 gnd 0.149881f
C5597 commonsourceibias.n389 gnd 0.007808f
C5598 commonsourceibias.n390 gnd 0.008022f
C5599 commonsourceibias.t52 gnd 0.149881f
C5600 commonsourceibias.n391 gnd 0.010321f
C5601 commonsourceibias.n392 gnd 0.008022f
C5602 commonsourceibias.t72 gnd 0.149881f
C5603 commonsourceibias.n393 gnd 0.007564f
C5604 commonsourceibias.n394 gnd 0.008022f
C5605 commonsourceibias.t38 gnd 0.149881f
C5606 commonsourceibias.n395 gnd 0.010168f
C5607 commonsourceibias.n396 gnd 0.008022f
C5608 commonsourceibias.t42 gnd 0.149881f
C5609 commonsourceibias.n397 gnd 0.007348f
C5610 commonsourceibias.n398 gnd 0.008022f
C5611 commonsourceibias.t36 gnd 0.149881f
C5612 commonsourceibias.n399 gnd 0.009997f
C5613 commonsourceibias.n400 gnd 0.008022f
C5614 commonsourceibias.t20 gnd 0.149881f
C5615 commonsourceibias.n401 gnd 0.007159f
C5616 commonsourceibias.n402 gnd 0.008022f
C5617 commonsourceibias.t28 gnd 0.149881f
C5618 commonsourceibias.n403 gnd 0.009806f
C5619 commonsourceibias.n404 gnd 0.008022f
C5620 commonsourceibias.t18 gnd 0.149881f
C5621 commonsourceibias.n405 gnd 0.006995f
C5622 commonsourceibias.n406 gnd 0.008022f
C5623 commonsourceibias.t58 gnd 0.149881f
C5624 commonsourceibias.n407 gnd 0.009595f
C5625 commonsourceibias.n408 gnd 0.008022f
C5626 commonsourceibias.t14 gnd 0.149881f
C5627 commonsourceibias.n409 gnd 0.006855f
C5628 commonsourceibias.n410 gnd 0.008022f
C5629 commonsourceibias.t66 gnd 0.149881f
C5630 commonsourceibias.n411 gnd 0.00936f
C5631 commonsourceibias.t16 gnd 0.16664f
C5632 commonsourceibias.t68 gnd 0.149881f
C5633 commonsourceibias.n412 gnd 0.065328f
C5634 commonsourceibias.n413 gnd 0.07169f
C5635 commonsourceibias.n414 gnd 0.033265f
C5636 commonsourceibias.n415 gnd 0.008022f
C5637 commonsourceibias.n416 gnd 0.007808f
C5638 commonsourceibias.n417 gnd 0.01119f
C5639 commonsourceibias.n418 gnd 0.059802f
C5640 commonsourceibias.n419 gnd 0.011182f
C5641 commonsourceibias.n420 gnd 0.008022f
C5642 commonsourceibias.n421 gnd 0.008022f
C5643 commonsourceibias.n422 gnd 0.008022f
C5644 commonsourceibias.n423 gnd 0.010321f
C5645 commonsourceibias.n424 gnd 0.059802f
C5646 commonsourceibias.n425 gnd 0.010563f
C5647 commonsourceibias.t56 gnd 0.149881f
C5648 commonsourceibias.n426 gnd 0.059802f
C5649 commonsourceibias.n427 gnd 0.010263f
C5650 commonsourceibias.n428 gnd 0.008022f
C5651 commonsourceibias.n429 gnd 0.008022f
C5652 commonsourceibias.n430 gnd 0.008022f
C5653 commonsourceibias.n431 gnd 0.007564f
C5654 commonsourceibias.n432 gnd 0.0112f
C5655 commonsourceibias.n433 gnd 0.059802f
C5656 commonsourceibias.n434 gnd 0.011196f
C5657 commonsourceibias.n435 gnd 0.008022f
C5658 commonsourceibias.n436 gnd 0.008022f
C5659 commonsourceibias.n437 gnd 0.008022f
C5660 commonsourceibias.n438 gnd 0.010168f
C5661 commonsourceibias.n439 gnd 0.059802f
C5662 commonsourceibias.n440 gnd 0.010488f
C5663 commonsourceibias.t62 gnd 0.149881f
C5664 commonsourceibias.n441 gnd 0.059802f
C5665 commonsourceibias.n442 gnd 0.010338f
C5666 commonsourceibias.n443 gnd 0.008022f
C5667 commonsourceibias.n444 gnd 0.008022f
C5668 commonsourceibias.n445 gnd 0.008022f
C5669 commonsourceibias.n446 gnd 0.007348f
C5670 commonsourceibias.n447 gnd 0.011204f
C5671 commonsourceibias.n448 gnd 0.059802f
C5672 commonsourceibias.n449 gnd 0.011203f
C5673 commonsourceibias.n450 gnd 0.008022f
C5674 commonsourceibias.n451 gnd 0.008022f
C5675 commonsourceibias.n452 gnd 0.008022f
C5676 commonsourceibias.n453 gnd 0.009997f
C5677 commonsourceibias.n454 gnd 0.059802f
C5678 commonsourceibias.n455 gnd 0.010413f
C5679 commonsourceibias.t2 gnd 0.149881f
C5680 commonsourceibias.n456 gnd 0.059802f
C5681 commonsourceibias.n457 gnd 0.010413f
C5682 commonsourceibias.n458 gnd 0.008022f
C5683 commonsourceibias.n459 gnd 0.008022f
C5684 commonsourceibias.n460 gnd 0.008022f
C5685 commonsourceibias.n461 gnd 0.007159f
C5686 commonsourceibias.n462 gnd 0.011203f
C5687 commonsourceibias.n463 gnd 0.059802f
C5688 commonsourceibias.n464 gnd 0.011204f
C5689 commonsourceibias.n465 gnd 0.008022f
C5690 commonsourceibias.n466 gnd 0.008022f
C5691 commonsourceibias.n467 gnd 0.008022f
C5692 commonsourceibias.n468 gnd 0.009806f
C5693 commonsourceibias.n469 gnd 0.059802f
C5694 commonsourceibias.n470 gnd 0.010338f
C5695 commonsourceibias.t10 gnd 0.149881f
C5696 commonsourceibias.n471 gnd 0.059802f
C5697 commonsourceibias.n472 gnd 0.010488f
C5698 commonsourceibias.n473 gnd 0.008022f
C5699 commonsourceibias.n474 gnd 0.008022f
C5700 commonsourceibias.n475 gnd 0.008022f
C5701 commonsourceibias.n476 gnd 0.006995f
C5702 commonsourceibias.n477 gnd 0.011196f
C5703 commonsourceibias.n478 gnd 0.059802f
C5704 commonsourceibias.n479 gnd 0.0112f
C5705 commonsourceibias.n480 gnd 0.008022f
C5706 commonsourceibias.n481 gnd 0.008022f
C5707 commonsourceibias.n482 gnd 0.008022f
C5708 commonsourceibias.n483 gnd 0.009595f
C5709 commonsourceibias.n484 gnd 0.059802f
C5710 commonsourceibias.n485 gnd 0.010263f
C5711 commonsourceibias.t30 gnd 0.149881f
C5712 commonsourceibias.n486 gnd 0.059802f
C5713 commonsourceibias.n487 gnd 0.010563f
C5714 commonsourceibias.n488 gnd 0.008022f
C5715 commonsourceibias.n489 gnd 0.008022f
C5716 commonsourceibias.n490 gnd 0.008022f
C5717 commonsourceibias.n491 gnd 0.006855f
C5718 commonsourceibias.n492 gnd 0.011182f
C5719 commonsourceibias.n493 gnd 0.059802f
C5720 commonsourceibias.n494 gnd 0.01119f
C5721 commonsourceibias.n495 gnd 0.008022f
C5722 commonsourceibias.n496 gnd 0.008022f
C5723 commonsourceibias.n497 gnd 0.008022f
C5724 commonsourceibias.n498 gnd 0.00936f
C5725 commonsourceibias.n499 gnd 0.059802f
C5726 commonsourceibias.n500 gnd 0.009843f
C5727 commonsourceibias.t32 gnd 0.162096f
C5728 commonsourceibias.n501 gnd 0.071758f
C5729 commonsourceibias.n502 gnd 0.079928f
C5730 commonsourceibias.t7 gnd 0.017311f
C5731 commonsourceibias.t33 gnd 0.017311f
C5732 commonsourceibias.n503 gnd 0.152968f
C5733 commonsourceibias.n504 gnd 0.132319f
C5734 commonsourceibias.t31 gnd 0.017311f
C5735 commonsourceibias.t53 gnd 0.017311f
C5736 commonsourceibias.n505 gnd 0.152968f
C5737 commonsourceibias.n506 gnd 0.070264f
C5738 commonsourceibias.t39 gnd 0.017311f
C5739 commonsourceibias.t73 gnd 0.017311f
C5740 commonsourceibias.n507 gnd 0.152968f
C5741 commonsourceibias.n508 gnd 0.070264f
C5742 commonsourceibias.t43 gnd 0.017311f
C5743 commonsourceibias.t11 gnd 0.017311f
C5744 commonsourceibias.n509 gnd 0.152968f
C5745 commonsourceibias.n510 gnd 0.070264f
C5746 commonsourceibias.t3 gnd 0.017311f
C5747 commonsourceibias.t37 gnd 0.017311f
C5748 commonsourceibias.n511 gnd 0.152968f
C5749 commonsourceibias.n512 gnd 0.058702f
C5750 commonsourceibias.n513 gnd 0.071082f
C5751 commonsourceibias.n514 gnd 0.05192f
C5752 commonsourceibias.t98 gnd 0.149881f
C5753 commonsourceibias.n515 gnd 0.059802f
C5754 commonsourceibias.n516 gnd 0.008022f
C5755 commonsourceibias.t125 gnd 0.149881f
C5756 commonsourceibias.n517 gnd 0.059802f
C5757 commonsourceibias.n518 gnd 0.008022f
C5758 commonsourceibias.t142 gnd 0.149881f
C5759 commonsourceibias.n519 gnd 0.059802f
C5760 commonsourceibias.n520 gnd 0.008022f
C5761 commonsourceibias.t155 gnd 0.149881f
C5762 commonsourceibias.n521 gnd 0.006995f
C5763 commonsourceibias.n522 gnd 0.008022f
C5764 commonsourceibias.t114 gnd 0.149881f
C5765 commonsourceibias.n523 gnd 0.009595f
C5766 commonsourceibias.n524 gnd 0.008022f
C5767 commonsourceibias.t148 gnd 0.149881f
C5768 commonsourceibias.n525 gnd 0.006855f
C5769 commonsourceibias.n526 gnd 0.008022f
C5770 commonsourceibias.t82 gnd 0.149881f
C5771 commonsourceibias.n527 gnd 0.00936f
C5772 commonsourceibias.t126 gnd 0.16664f
C5773 commonsourceibias.t89 gnd 0.149881f
C5774 commonsourceibias.n528 gnd 0.065328f
C5775 commonsourceibias.n529 gnd 0.07169f
C5776 commonsourceibias.n530 gnd 0.033265f
C5777 commonsourceibias.n531 gnd 0.008022f
C5778 commonsourceibias.n532 gnd 0.007808f
C5779 commonsourceibias.n533 gnd 0.01119f
C5780 commonsourceibias.n534 gnd 0.059802f
C5781 commonsourceibias.n535 gnd 0.011182f
C5782 commonsourceibias.n536 gnd 0.008022f
C5783 commonsourceibias.n537 gnd 0.008022f
C5784 commonsourceibias.n538 gnd 0.008022f
C5785 commonsourceibias.n539 gnd 0.010321f
C5786 commonsourceibias.n540 gnd 0.059802f
C5787 commonsourceibias.n541 gnd 0.010563f
C5788 commonsourceibias.t134 gnd 0.149881f
C5789 commonsourceibias.n542 gnd 0.059802f
C5790 commonsourceibias.n543 gnd 0.010263f
C5791 commonsourceibias.n544 gnd 0.008022f
C5792 commonsourceibias.n545 gnd 0.008022f
C5793 commonsourceibias.n546 gnd 0.008022f
C5794 commonsourceibias.n547 gnd 0.007564f
C5795 commonsourceibias.n548 gnd 0.0112f
C5796 commonsourceibias.n549 gnd 0.059802f
C5797 commonsourceibias.n550 gnd 0.011196f
C5798 commonsourceibias.n551 gnd 0.008022f
C5799 commonsourceibias.n552 gnd 0.008022f
C5800 commonsourceibias.n553 gnd 0.008022f
C5801 commonsourceibias.n554 gnd 0.010168f
C5802 commonsourceibias.n555 gnd 0.059802f
C5803 commonsourceibias.n556 gnd 0.010488f
C5804 commonsourceibias.n557 gnd 0.010338f
C5805 commonsourceibias.n558 gnd 0.008022f
C5806 commonsourceibias.n559 gnd 0.008022f
C5807 commonsourceibias.n560 gnd 0.009806f
C5808 commonsourceibias.n561 gnd 0.007348f
C5809 commonsourceibias.n562 gnd 0.011204f
C5810 commonsourceibias.n563 gnd 0.008022f
C5811 commonsourceibias.n564 gnd 0.008022f
C5812 commonsourceibias.n565 gnd 0.011203f
C5813 commonsourceibias.n566 gnd 0.007159f
C5814 commonsourceibias.n567 gnd 0.009997f
C5815 commonsourceibias.n568 gnd 0.008022f
C5816 commonsourceibias.n569 gnd 0.007008f
C5817 commonsourceibias.n570 gnd 0.010413f
C5818 commonsourceibias.t149 gnd 0.149881f
C5819 commonsourceibias.n571 gnd 0.059802f
C5820 commonsourceibias.n572 gnd 0.010413f
C5821 commonsourceibias.n573 gnd 0.007008f
C5822 commonsourceibias.n574 gnd 0.008022f
C5823 commonsourceibias.n575 gnd 0.008022f
C5824 commonsourceibias.n576 gnd 0.007159f
C5825 commonsourceibias.n577 gnd 0.011203f
C5826 commonsourceibias.n578 gnd 0.059802f
C5827 commonsourceibias.n579 gnd 0.011204f
C5828 commonsourceibias.n580 gnd 0.008022f
C5829 commonsourceibias.n581 gnd 0.008022f
C5830 commonsourceibias.n582 gnd 0.008022f
C5831 commonsourceibias.n583 gnd 0.009806f
C5832 commonsourceibias.n584 gnd 0.059802f
C5833 commonsourceibias.n585 gnd 0.010338f
C5834 commonsourceibias.t156 gnd 0.149881f
C5835 commonsourceibias.n586 gnd 0.059802f
C5836 commonsourceibias.n587 gnd 0.010488f
C5837 commonsourceibias.n588 gnd 0.008022f
C5838 commonsourceibias.n589 gnd 0.008022f
C5839 commonsourceibias.n590 gnd 0.008022f
C5840 commonsourceibias.n591 gnd 0.006995f
C5841 commonsourceibias.n592 gnd 0.011196f
C5842 commonsourceibias.n593 gnd 0.059802f
C5843 commonsourceibias.n594 gnd 0.0112f
C5844 commonsourceibias.n595 gnd 0.008022f
C5845 commonsourceibias.n596 gnd 0.008022f
C5846 commonsourceibias.n597 gnd 0.008022f
C5847 commonsourceibias.n598 gnd 0.009595f
C5848 commonsourceibias.n599 gnd 0.059802f
C5849 commonsourceibias.n600 gnd 0.010263f
C5850 commonsourceibias.t105 gnd 0.149881f
C5851 commonsourceibias.n601 gnd 0.059802f
C5852 commonsourceibias.n602 gnd 0.010563f
C5853 commonsourceibias.n603 gnd 0.008022f
C5854 commonsourceibias.n604 gnd 0.008022f
C5855 commonsourceibias.n605 gnd 0.008022f
C5856 commonsourceibias.n606 gnd 0.006855f
C5857 commonsourceibias.n607 gnd 0.011182f
C5858 commonsourceibias.n608 gnd 0.059802f
C5859 commonsourceibias.n609 gnd 0.01119f
C5860 commonsourceibias.n610 gnd 0.008022f
C5861 commonsourceibias.n611 gnd 0.008022f
C5862 commonsourceibias.n612 gnd 0.008022f
C5863 commonsourceibias.n613 gnd 0.00936f
C5864 commonsourceibias.n614 gnd 0.059802f
C5865 commonsourceibias.n615 gnd 0.009843f
C5866 commonsourceibias.n616 gnd 0.071758f
C5867 commonsourceibias.n617 gnd 0.046883f
C5868 commonsourceibias.n618 gnd 0.010705f
C5869 commonsourceibias.t141 gnd 0.149881f
C5870 commonsourceibias.n619 gnd 0.007808f
C5871 commonsourceibias.n620 gnd 0.008022f
C5872 commonsourceibias.t154 gnd 0.149881f
C5873 commonsourceibias.n621 gnd 0.010321f
C5874 commonsourceibias.n622 gnd 0.008022f
C5875 commonsourceibias.t132 gnd 0.149881f
C5876 commonsourceibias.n623 gnd 0.007564f
C5877 commonsourceibias.n624 gnd 0.008022f
C5878 commonsourceibias.t147 gnd 0.149881f
C5879 commonsourceibias.n625 gnd 0.010168f
C5880 commonsourceibias.n626 gnd 0.008022f
C5881 commonsourceibias.t123 gnd 0.149881f
C5882 commonsourceibias.n627 gnd 0.007348f
C5883 commonsourceibias.n628 gnd 0.008022f
C5884 commonsourceibias.t115 gnd 0.149881f
C5885 commonsourceibias.n629 gnd 0.009997f
C5886 commonsourceibias.n630 gnd 0.008022f
C5887 commonsourceibias.t88 gnd 0.149881f
C5888 commonsourceibias.n631 gnd 0.007159f
C5889 commonsourceibias.n632 gnd 0.008022f
C5890 commonsourceibias.t106 gnd 0.149881f
C5891 commonsourceibias.n633 gnd 0.009806f
C5892 commonsourceibias.n634 gnd 0.008022f
C5893 commonsourceibias.t143 gnd 0.149881f
C5894 commonsourceibias.n635 gnd 0.006995f
C5895 commonsourceibias.n636 gnd 0.008022f
C5896 commonsourceibias.t99 gnd 0.149881f
C5897 commonsourceibias.n637 gnd 0.009595f
C5898 commonsourceibias.n638 gnd 0.008022f
C5899 commonsourceibias.t136 gnd 0.149881f
C5900 commonsourceibias.n639 gnd 0.006855f
C5901 commonsourceibias.n640 gnd 0.008022f
C5902 commonsourceibias.t150 gnd 0.149881f
C5903 commonsourceibias.n641 gnd 0.00936f
C5904 commonsourceibias.t108 gnd 0.16664f
C5905 commonsourceibias.t158 gnd 0.149881f
C5906 commonsourceibias.n642 gnd 0.065328f
C5907 commonsourceibias.n643 gnd 0.07169f
C5908 commonsourceibias.n644 gnd 0.033265f
C5909 commonsourceibias.n645 gnd 0.008022f
C5910 commonsourceibias.n646 gnd 0.007808f
C5911 commonsourceibias.n647 gnd 0.01119f
C5912 commonsourceibias.n648 gnd 0.059802f
C5913 commonsourceibias.n649 gnd 0.011182f
C5914 commonsourceibias.n650 gnd 0.008022f
C5915 commonsourceibias.n651 gnd 0.008022f
C5916 commonsourceibias.n652 gnd 0.008022f
C5917 commonsourceibias.n653 gnd 0.010321f
C5918 commonsourceibias.n654 gnd 0.059802f
C5919 commonsourceibias.n655 gnd 0.010563f
C5920 commonsourceibias.t118 gnd 0.149881f
C5921 commonsourceibias.n656 gnd 0.059802f
C5922 commonsourceibias.n657 gnd 0.010263f
C5923 commonsourceibias.n658 gnd 0.008022f
C5924 commonsourceibias.n659 gnd 0.008022f
C5925 commonsourceibias.n660 gnd 0.008022f
C5926 commonsourceibias.n661 gnd 0.007564f
C5927 commonsourceibias.n662 gnd 0.0112f
C5928 commonsourceibias.n663 gnd 0.059802f
C5929 commonsourceibias.n664 gnd 0.011196f
C5930 commonsourceibias.n665 gnd 0.008022f
C5931 commonsourceibias.n666 gnd 0.008022f
C5932 commonsourceibias.n667 gnd 0.008022f
C5933 commonsourceibias.n668 gnd 0.010168f
C5934 commonsourceibias.n669 gnd 0.059802f
C5935 commonsourceibias.n670 gnd 0.010488f
C5936 commonsourceibias.t128 gnd 0.149881f
C5937 commonsourceibias.n671 gnd 0.059802f
C5938 commonsourceibias.n672 gnd 0.010338f
C5939 commonsourceibias.n673 gnd 0.008022f
C5940 commonsourceibias.n674 gnd 0.008022f
C5941 commonsourceibias.n675 gnd 0.008022f
C5942 commonsourceibias.n676 gnd 0.007348f
C5943 commonsourceibias.n677 gnd 0.011204f
C5944 commonsourceibias.n678 gnd 0.059802f
C5945 commonsourceibias.n679 gnd 0.011203f
C5946 commonsourceibias.n680 gnd 0.008022f
C5947 commonsourceibias.n681 gnd 0.008022f
C5948 commonsourceibias.n682 gnd 0.008022f
C5949 commonsourceibias.n683 gnd 0.009997f
C5950 commonsourceibias.n684 gnd 0.059802f
C5951 commonsourceibias.n685 gnd 0.010413f
C5952 commonsourceibias.t137 gnd 0.149881f
C5953 commonsourceibias.n686 gnd 0.059802f
C5954 commonsourceibias.n687 gnd 0.010413f
C5955 commonsourceibias.n688 gnd 0.008022f
C5956 commonsourceibias.n689 gnd 0.008022f
C5957 commonsourceibias.n690 gnd 0.008022f
C5958 commonsourceibias.n691 gnd 0.007159f
C5959 commonsourceibias.n692 gnd 0.011203f
C5960 commonsourceibias.n693 gnd 0.059802f
C5961 commonsourceibias.n694 gnd 0.011204f
C5962 commonsourceibias.n695 gnd 0.008022f
C5963 commonsourceibias.n696 gnd 0.008022f
C5964 commonsourceibias.n697 gnd 0.008022f
C5965 commonsourceibias.n698 gnd 0.009806f
C5966 commonsourceibias.n699 gnd 0.059802f
C5967 commonsourceibias.n700 gnd 0.010338f
C5968 commonsourceibias.t144 gnd 0.149881f
C5969 commonsourceibias.n701 gnd 0.059802f
C5970 commonsourceibias.n702 gnd 0.010488f
C5971 commonsourceibias.n703 gnd 0.008022f
C5972 commonsourceibias.n704 gnd 0.008022f
C5973 commonsourceibias.n705 gnd 0.008022f
C5974 commonsourceibias.n706 gnd 0.006995f
C5975 commonsourceibias.n707 gnd 0.011196f
C5976 commonsourceibias.n708 gnd 0.059802f
C5977 commonsourceibias.n709 gnd 0.0112f
C5978 commonsourceibias.n710 gnd 0.008022f
C5979 commonsourceibias.n711 gnd 0.008022f
C5980 commonsourceibias.n712 gnd 0.008022f
C5981 commonsourceibias.n713 gnd 0.009595f
C5982 commonsourceibias.n714 gnd 0.059802f
C5983 commonsourceibias.n715 gnd 0.010263f
C5984 commonsourceibias.t93 gnd 0.149881f
C5985 commonsourceibias.n716 gnd 0.059802f
C5986 commonsourceibias.n717 gnd 0.010563f
C5987 commonsourceibias.n718 gnd 0.008022f
C5988 commonsourceibias.n719 gnd 0.008022f
C5989 commonsourceibias.n720 gnd 0.008022f
C5990 commonsourceibias.n721 gnd 0.006855f
C5991 commonsourceibias.n722 gnd 0.011182f
C5992 commonsourceibias.n723 gnd 0.059802f
C5993 commonsourceibias.n724 gnd 0.01119f
C5994 commonsourceibias.n725 gnd 0.008022f
C5995 commonsourceibias.n726 gnd 0.008022f
C5996 commonsourceibias.n727 gnd 0.008022f
C5997 commonsourceibias.n728 gnd 0.00936f
C5998 commonsourceibias.n729 gnd 0.059802f
C5999 commonsourceibias.n730 gnd 0.009843f
C6000 commonsourceibias.t124 gnd 0.162096f
C6001 commonsourceibias.n731 gnd 0.071758f
C6002 commonsourceibias.n732 gnd 0.024957f
C6003 commonsourceibias.n733 gnd 0.221543f
C6004 commonsourceibias.n734 gnd 4.49224f
.ends

