* NGSPICE file created from opamp345.ext - technology: sky130A

.subckt opamp345 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 a_n2140_13878.t15 a_n2408_n452.t19 a_n2408_n452.t20 vdd.t129 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X1 CSoutput.t76 a_n6308_8799.t40 vdd.t159 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X2 a_n2140_13878.t21 a_n2408_n452.t56 vdd.t140 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 vdd.t77 vdd.t75 vdd.t76 vdd.t7 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X4 gnd.t218 gnd.t216 gnd.t217 gnd.t184 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X5 a_n6308_8799.t17 plus.t5 a_n2903_n3924.t30 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X6 gnd.t215 gnd.t212 gnd.t214 gnd.t213 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X7 commonsourceibias.t47 commonsourceibias.t46 gnd.t237 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X8 gnd.t9 commonsourceibias.t48 CSoutput.t1 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X9 gnd.t211 gnd.t209 gnd.t210 gnd.t191 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X10 gnd.t208 gnd.t206 minus.t4 gnd.t207 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X11 output.t3 outputibias.t8 gnd.t287 gnd.t286 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X12 output.t19 CSoutput.t96 vdd.t203 gnd.t101 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X13 CSoutput.t75 a_n6308_8799.t41 vdd.t161 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X14 gnd.t39 commonsourceibias.t49 CSoutput.t9 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X15 a_n2903_n3924.t29 plus.t6 a_n6308_8799.t18 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X16 gnd.t273 commonsourceibias.t44 commonsourceibias.t45 gnd.t64 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X17 a_n2318_8322.t23 a_n2408_n452.t57 a_n6308_8799.t6 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X18 gnd.t285 commonsourceibias.t50 CSoutput.t93 gnd.t64 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 a_n2903_n3924.t35 minus.t5 a_n2408_n452.t40 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X20 outputibias.t7 outputibias.t6 gnd.t13 gnd.t12 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X21 output.t18 CSoutput.t97 vdd.t151 gnd.t100 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X22 a_n2408_n452.t0 minus.t6 a_n2903_n3924.t0 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X23 a_n6308_8799.t15 a_n2408_n452.t58 a_n2318_8322.t22 vdd.t127 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X24 gnd.t264 commonsourceibias.t42 commonsourceibias.t43 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X25 CSoutput.t74 a_n6308_8799.t42 vdd.t175 vdd.t82 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X26 vdd.t176 a_n6308_8799.t43 CSoutput.t73 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X27 a_n2408_n452.t48 minus.t7 a_n2903_n3924.t47 gnd.t270 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X28 a_n6308_8799.t1 a_n2408_n452.t59 a_n2318_8322.t21 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X29 vdd.t74 vdd.t72 vdd.t73 vdd.t7 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X30 CSoutput.t83 commonsourceibias.t51 gnd.t258 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X31 a_n2903_n3924.t52 minus.t8 a_n2408_n452.t53 gnd.t271 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X32 CSoutput.t98 a_n2318_8322.t24 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X33 gnd.t49 commonsourceibias.t40 commonsourceibias.t41 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X34 vdd.t71 vdd.t69 vdd.t70 vdd.t11 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X35 CSoutput.t72 a_n6308_8799.t44 vdd.t199 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X36 vdd.t152 CSoutput.t99 output.t17 gnd.t99 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X37 vdd.t153 CSoutput.t100 output.t16 gnd.t98 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X38 CSoutput.t71 a_n6308_8799.t45 vdd.t200 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X39 CSoutput.t88 commonsourceibias.t52 gnd.t275 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X40 a_n2903_n3924.t33 diffpairibias.t16 gnd.t72 gnd.t71 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X41 CSoutput.t70 a_n6308_8799.t46 vdd.t191 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X42 CSoutput.t24 commonsourceibias.t53 gnd.t221 gnd.t104 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 a_n2903_n3924.t28 plus.t7 a_n6308_8799.t29 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X44 a_n2140_13878.t14 a_n2408_n452.t33 a_n2408_n452.t34 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X45 a_n2408_n452.t28 a_n2408_n452.t27 a_n2140_13878.t13 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X46 CSoutput.t15 commonsourceibias.t54 gnd.t67 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X47 a_n6308_8799.t27 plus.t8 a_n2903_n3924.t27 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X48 a_n6308_8799.t30 plus.t9 a_n2903_n3924.t26 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X49 vdd.t68 vdd.t66 vdd.t67 vdd.t49 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X50 a_n2903_n3924.t25 plus.t10 a_n6308_8799.t26 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X51 a_n2408_n452.t39 minus.t9 a_n2903_n3924.t31 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X52 diffpairibias.t15 diffpairibias.t14 gnd.t279 gnd.t278 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X53 gnd.t205 gnd.t203 gnd.t204 gnd.t191 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X54 a_n6308_8799.t2 a_n2408_n452.t60 a_n2318_8322.t20 vdd.t122 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X55 gnd.t202 gnd.t200 plus.t4 gnd.t201 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X56 gnd.t225 commonsourceibias.t55 CSoutput.t27 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X57 gnd.t21 commonsourceibias.t56 CSoutput.t3 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X58 diffpairibias.t13 diffpairibias.t12 gnd.t110 gnd.t109 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X59 output.t15 CSoutput.t101 vdd.t154 gnd.t97 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X60 gnd.t70 commonsourceibias.t57 CSoutput.t17 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X61 commonsourceibias.t39 commonsourceibias.t38 gnd.t43 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X62 vdd.t155 CSoutput.t102 output.t14 gnd.t96 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X63 CSoutput.t69 a_n6308_8799.t47 vdd.t192 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X64 vdd.t189 a_n6308_8799.t48 CSoutput.t68 vdd.t86 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X65 CSoutput.t67 a_n6308_8799.t49 vdd.t190 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X66 CSoutput.t66 a_n6308_8799.t50 vdd.t142 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X67 gnd.t199 gnd.t197 gnd.t198 gnd.t127 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X68 gnd.t196 gnd.t194 plus.t3 gnd.t195 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X69 gnd.t274 commonsourceibias.t58 CSoutput.t87 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X70 a_n2903_n3924.t24 plus.t11 a_n6308_8799.t38 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X71 commonsourceibias.t37 commonsourceibias.t36 gnd.t103 gnd.t102 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X72 a_n2903_n3924.t55 diffpairibias.t17 gnd.t291 gnd.t290 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X73 gnd.t19 commonsourceibias.t34 commonsourceibias.t35 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X74 vdd.t144 a_n6308_8799.t51 CSoutput.t65 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X75 vdd.t181 a_n6308_8799.t52 CSoutput.t64 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X76 a_n6308_8799.t7 a_n2408_n452.t61 a_n2318_8322.t19 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X77 a_n2408_n452.t14 a_n2408_n452.t13 a_n2140_13878.t12 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X78 a_n2408_n452.t18 a_n2408_n452.t17 a_n2140_13878.t11 vdd.t99 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X79 gnd.t280 commonsourceibias.t32 commonsourceibias.t33 gnd.t79 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X80 commonsourceibias.t31 commonsourceibias.t30 gnd.t246 gnd.t104 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X81 outputibias.t5 outputibias.t4 gnd.t76 gnd.t75 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X82 CSoutput.t63 a_n6308_8799.t53 vdd.t182 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 vdd.t146 a_n6308_8799.t54 CSoutput.t62 vdd.t145 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X84 CSoutput.t94 commonsourceibias.t59 gnd.t288 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 a_n2408_n452.t5 minus.t10 a_n2903_n3924.t5 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X86 vdd.t188 CSoutput.t103 output.t13 gnd.t95 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X87 vdd.t65 vdd.t63 vdd.t64 vdd.t23 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X88 vdd.t62 vdd.t60 vdd.t61 vdd.t53 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X89 CSoutput.t79 commonsourceibias.t60 gnd.t244 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 vdd.t59 vdd.t56 vdd.t58 vdd.t57 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X91 gnd.t268 commonsourceibias.t61 CSoutput.t86 gnd.t79 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X92 gnd.t193 gnd.t190 gnd.t192 gnd.t191 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X93 commonsourceibias.t29 commonsourceibias.t28 gnd.t238 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 CSoutput.t84 commonsourceibias.t62 gnd.t259 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X95 a_n2903_n3924.t6 minus.t11 a_n2408_n452.t6 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X96 CSoutput.t104 a_n2318_8322.t25 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X97 outputibias.t3 outputibias.t2 gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X98 a_n2318_8322.t7 a_n2408_n452.t62 vdd.t137 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X99 vdd.t135 a_n2408_n452.t63 a_n2318_8322.t6 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X100 a_n2408_n452.t12 a_n2408_n452.t11 a_n2140_13878.t10 vdd.t106 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X101 CSoutput.t61 a_n6308_8799.t55 vdd.t148 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X102 a_n2903_n3924.t32 diffpairibias.t18 gnd.t57 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X103 a_n2903_n3924.t40 minus.t12 a_n2408_n452.t42 gnd.t85 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X104 a_n2903_n3924.t4 minus.t13 a_n2408_n452.t4 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X105 commonsourceibias.t27 commonsourceibias.t26 gnd.t243 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X106 vdd.t133 a_n2408_n452.t64 a_n2140_13878.t22 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X107 a_n2408_n452.t54 minus.t14 a_n2903_n3924.t53 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X108 vdd.t55 vdd.t52 vdd.t54 vdd.t53 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X109 a_n2903_n3924.t23 plus.t12 a_n6308_8799.t25 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X110 a_n2903_n3924.t22 plus.t13 a_n6308_8799.t28 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X111 vdd.t149 a_n6308_8799.t56 CSoutput.t60 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X112 a_n2408_n452.t46 minus.t15 a_n2903_n3924.t45 gnd.t269 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X113 gnd.t59 commonsourceibias.t24 commonsourceibias.t25 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X114 gnd.t81 commonsourceibias.t63 CSoutput.t20 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X115 gnd.t189 gnd.t187 plus.t2 gnd.t188 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X116 a_n6308_8799.t32 plus.t14 a_n2903_n3924.t21 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X117 a_n6308_8799.t12 a_n2408_n452.t65 a_n2318_8322.t18 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X118 a_n2318_8322.t5 a_n2408_n452.t66 vdd.t131 vdd.t130 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X119 vdd.t51 vdd.t48 vdd.t50 vdd.t49 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X120 gnd.t281 commonsourceibias.t64 CSoutput.t90 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X121 a_n6308_8799.t21 plus.t15 a_n2903_n3924.t20 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X122 gnd.t219 commonsourceibias.t65 CSoutput.t23 gnd.t28 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X123 vdd.t150 a_n6308_8799.t57 CSoutput.t59 vdd.t145 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X124 a_n2408_n452.t16 a_n2408_n452.t15 a_n2140_13878.t9 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X125 a_n2408_n452.t47 minus.t16 a_n2903_n3924.t46 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X126 diffpairibias.t11 diffpairibias.t10 gnd.t83 gnd.t82 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X127 CSoutput.t58 a_n6308_8799.t58 vdd.t169 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X128 a_n6308_8799.t4 a_n2408_n452.t67 a_n2318_8322.t17 vdd.t129 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X129 gnd.t41 commonsourceibias.t66 CSoutput.t10 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X130 a_n2140_13878.t8 a_n2408_n452.t37 a_n2408_n452.t38 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X131 outputibias.t1 outputibias.t0 gnd.t257 gnd.t256 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X132 vdd.t47 vdd.t45 vdd.t46 vdd.t23 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X133 gnd.t231 commonsourceibias.t67 CSoutput.t77 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X134 a_n2903_n3924.t3 minus.t17 a_n2408_n452.t3 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X135 CSoutput.t105 a_n2318_8322.t27 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X136 a_n2140_13878.t7 a_n2408_n452.t35 a_n2408_n452.t36 vdd.t127 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X137 vdd.t126 a_n2408_n452.t68 a_n2318_8322.t4 vdd.t125 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X138 CSoutput.t12 commonsourceibias.t68 gnd.t62 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X139 gnd.t186 gnd.t183 gnd.t185 gnd.t184 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X140 CSoutput.t106 a_n2318_8322.t26 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X141 a_n2408_n452.t22 a_n2408_n452.t21 a_n2140_13878.t6 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X142 minus.t3 gnd.t180 gnd.t182 gnd.t181 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X143 a_n2903_n3924.t19 plus.t16 a_n6308_8799.t24 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X144 gnd.t179 gnd.t176 gnd.t178 gnd.t177 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X145 a_n2903_n3924.t41 diffpairibias.t19 gnd.t261 gnd.t260 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X146 CSoutput.t11 commonsourceibias.t69 gnd.t55 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X147 CSoutput.t7 commonsourceibias.t70 gnd.t33 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X148 a_n2903_n3924.t39 diffpairibias.t20 gnd.t255 gnd.t254 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X149 vdd.t156 CSoutput.t107 output.t12 gnd.t94 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X150 vdd.t170 a_n6308_8799.t59 CSoutput.t57 vdd.t162 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X151 gnd.t80 commonsourceibias.t71 CSoutput.t19 gnd.t79 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X152 a_n6308_8799.t19 plus.t17 a_n2903_n3924.t18 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X153 CSoutput.t2 commonsourceibias.t72 gnd.t11 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X154 CSoutput.t56 a_n6308_8799.t60 vdd.t167 vdd.t166 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X155 CSoutput.t55 a_n6308_8799.t61 vdd.t168 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X156 a_n2140_13878.t17 a_n2408_n452.t69 vdd.t124 vdd.t123 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X157 gnd.t175 gnd.t173 gnd.t174 gnd.t134 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X158 diffpairibias.t9 diffpairibias.t8 gnd.t230 gnd.t229 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X159 vdd.t121 a_n2408_n452.t70 a_n2140_13878.t16 vdd.t120 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X160 CSoutput.t82 commonsourceibias.t73 gnd.t249 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X161 gnd.t74 commonsourceibias.t74 CSoutput.t18 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X162 a_n2140_13878.t5 a_n2408_n452.t7 a_n2408_n452.t8 vdd.t122 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X163 plus.t1 gnd.t170 gnd.t172 gnd.t171 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X164 gnd.t267 commonsourceibias.t22 commonsourceibias.t23 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 gnd.t37 commonsourceibias.t75 CSoutput.t8 gnd.t28 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X166 a_n2903_n3924.t38 minus.t18 a_n2408_n452.t41 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X167 a_n2318_8322.t16 a_n2408_n452.t71 a_n6308_8799.t10 vdd.t93 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X168 gnd.t226 commonsourceibias.t76 CSoutput.t28 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X169 a_n2408_n452.t2 minus.t19 a_n2903_n3924.t2 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X170 a_n2408_n452.t1 minus.t20 a_n2903_n3924.t1 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X171 diffpairibias.t7 diffpairibias.t6 gnd.t45 gnd.t44 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X172 vdd.t163 a_n6308_8799.t62 CSoutput.t54 vdd.t162 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X173 vdd.t119 a_n2408_n452.t72 a_n2318_8322.t3 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X174 a_n2408_n452.t44 minus.t21 a_n2903_n3924.t43 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X175 gnd.t58 commonsourceibias.t20 commonsourceibias.t21 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X176 CSoutput.t22 commonsourceibias.t77 gnd.t106 gnd.t102 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X177 a_n2903_n3924.t48 minus.t22 a_n2408_n452.t49 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X178 a_n6308_8799.t39 plus.t18 a_n2903_n3924.t17 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X179 gnd.t169 gnd.t167 gnd.t168 gnd.t134 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X180 gnd.t166 gnd.t164 gnd.t165 gnd.t119 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X181 CSoutput.t5 commonsourceibias.t78 gnd.t24 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X182 a_n2903_n3924.t42 minus.t23 a_n2408_n452.t43 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X183 a_n2140_13878.t19 a_n2408_n452.t73 vdd.t98 vdd.t97 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X184 vdd.t165 a_n6308_8799.t63 CSoutput.t53 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X185 vdd.t44 vdd.t42 vdd.t43 vdd.t3 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X186 CSoutput.t52 a_n6308_8799.t64 vdd.t197 vdd.t82 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X187 CSoutput.t51 a_n6308_8799.t65 vdd.t198 vdd.t166 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X188 gnd.t163 gnd.t161 minus.t2 gnd.t162 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X189 gnd.t36 commonsourceibias.t18 commonsourceibias.t19 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X190 gnd.t160 gnd.t157 gnd.t159 gnd.t158 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X191 a_n2318_8322.t15 a_n2408_n452.t74 a_n6308_8799.t13 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X192 vdd.t116 a_n2408_n452.t75 a_n2318_8322.t2 vdd.t115 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X193 CSoutput.t50 a_n6308_8799.t66 vdd.t183 vdd.t166 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X194 CSoutput.t25 commonsourceibias.t79 gnd.t223 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X195 a_n2903_n3924.t37 diffpairibias.t21 gnd.t233 gnd.t232 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X196 output.t11 CSoutput.t108 vdd.t157 gnd.t93 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X197 CSoutput.t49 a_n6308_8799.t67 vdd.t184 vdd.t84 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X198 vdd.t79 a_n6308_8799.t68 CSoutput.t48 vdd.t78 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X199 CSoutput.t4 commonsourceibias.t80 gnd.t22 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X200 vdd.t81 a_n6308_8799.t69 CSoutput.t47 vdd.t80 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X201 vdd.t90 a_n6308_8799.t70 CSoutput.t46 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X202 CSoutput.t109 a_n2318_8322.t25 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X203 CSoutput.t92 commonsourceibias.t81 gnd.t283 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X204 a_n6308_8799.t37 plus.t19 a_n2903_n3924.t16 gnd.t270 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X205 vdd.t41 vdd.t39 vdd.t40 vdd.t19 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X206 gnd.t289 commonsourceibias.t82 CSoutput.t95 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 output.t2 outputibias.t9 gnd.t253 gnd.t252 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X208 output.t10 CSoutput.t110 vdd.t173 gnd.t92 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X209 vdd.t38 vdd.t35 vdd.t37 vdd.t36 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X210 a_n2903_n3924.t15 plus.t20 a_n6308_8799.t35 gnd.t271 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X211 gnd.t156 gnd.t154 gnd.t155 gnd.t123 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X212 a_n2140_13878.t4 a_n2408_n452.t29 a_n2408_n452.t30 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X213 a_n2318_8322.t14 a_n2408_n452.t76 a_n6308_8799.t0 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X214 gnd.t153 gnd.t151 gnd.t152 gnd.t123 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X215 output.t1 outputibias.t10 gnd.t251 gnd.t250 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X216 diffpairibias.t5 diffpairibias.t4 gnd.t263 gnd.t262 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X217 CSoutput.t45 a_n6308_8799.t71 vdd.t92 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X218 vdd.t177 a_n6308_8799.t72 CSoutput.t44 vdd.t80 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X219 gnd.t247 commonsourceibias.t83 CSoutput.t80 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X220 CSoutput.t13 commonsourceibias.t84 gnd.t63 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X221 vdd.t178 a_n6308_8799.t73 CSoutput.t43 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X222 vdd.t34 vdd.t32 vdd.t33 vdd.t3 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X223 CSoutput.t42 a_n6308_8799.t74 vdd.t83 vdd.t82 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X224 a_n2318_8322.t1 a_n2408_n452.t77 vdd.t113 vdd.t112 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X225 gnd.t241 commonsourceibias.t85 CSoutput.t78 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X226 gnd.t29 commonsourceibias.t16 commonsourceibias.t17 gnd.t28 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X227 output.t9 CSoutput.t111 vdd.t174 gnd.t91 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X228 vdd.t31 vdd.t29 vdd.t30 vdd.t15 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X229 gnd.t150 gnd.t147 gnd.t149 gnd.t148 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X230 vdd.t111 a_n2408_n452.t78 a_n2140_13878.t20 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X231 plus.t0 gnd.t144 gnd.t146 gnd.t145 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X232 gnd.t143 gnd.t140 gnd.t142 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X233 CSoutput.t41 a_n6308_8799.t75 vdd.t85 vdd.t84 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X234 vdd.t193 a_n6308_8799.t76 CSoutput.t40 vdd.t80 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X235 vdd.t194 a_n6308_8799.t77 CSoutput.t39 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X236 gnd.t139 gnd.t137 gnd.t138 gnd.t119 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X237 CSoutput.t26 commonsourceibias.t86 gnd.t224 gnd.t102 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X238 a_n2903_n3924.t14 plus.t21 a_n6308_8799.t20 gnd.t85 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X239 CSoutput.t85 commonsourceibias.t87 gnd.t265 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X240 gnd.t136 gnd.t133 gnd.t135 gnd.t134 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X241 vdd.t185 CSoutput.t112 output.t8 gnd.t90 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X242 vdd.t28 vdd.t26 vdd.t27 vdd.t19 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X243 a_n6308_8799.t9 a_n2408_n452.t79 a_n2318_8322.t13 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X244 a_n2318_8322.t12 a_n2408_n452.t80 a_n6308_8799.t3 vdd.t103 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X245 CSoutput.t38 a_n6308_8799.t78 vdd.t171 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X246 a_n2903_n3924.t44 minus.t24 a_n2408_n452.t45 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X247 a_n2140_13878.t23 a_n2408_n452.t81 vdd.t108 vdd.t107 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X248 vdd.t172 a_n6308_8799.t79 CSoutput.t37 vdd.t162 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X249 a_n6308_8799.t36 plus.t22 a_n2903_n3924.t13 gnd.t269 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X250 a_n2408_n452.t52 minus.t25 a_n2903_n3924.t51 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X251 output.t0 outputibias.t11 gnd.t108 gnd.t107 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X252 a_n2318_8322.t11 a_n2408_n452.t82 a_n6308_8799.t14 vdd.t106 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X253 gnd.t132 gnd.t130 minus.t1 gnd.t131 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X254 gnd.t129 gnd.t126 gnd.t128 gnd.t127 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X255 a_n6308_8799.t22 plus.t23 a_n2903_n3924.t12 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X256 CSoutput.t91 commonsourceibias.t88 gnd.t282 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X257 a_n2903_n3924.t54 minus.t26 a_n2408_n452.t55 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X258 vdd.t186 CSoutput.t113 output.t7 gnd.t89 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X259 a_n2140_13878.t3 a_n2408_n452.t9 a_n2408_n452.t10 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X260 commonsourceibias.t15 commonsourceibias.t14 gnd.t220 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X261 output.t6 CSoutput.t114 vdd.t187 gnd.t88 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X262 vdd.t25 vdd.t22 vdd.t24 vdd.t23 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X263 a_n2903_n3924.t11 plus.t24 a_n6308_8799.t33 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X264 gnd.t3 commonsourceibias.t89 CSoutput.t0 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X265 vdd.t21 vdd.t18 vdd.t20 vdd.t19 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X266 gnd.t248 commonsourceibias.t90 CSoutput.t81 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X267 output.t5 CSoutput.t115 vdd.t0 gnd.t87 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X268 vdd.t201 a_n6308_8799.t80 CSoutput.t36 vdd.t86 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X269 gnd.t125 gnd.t122 gnd.t124 gnd.t123 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X270 a_n2903_n3924.t34 diffpairibias.t22 gnd.t78 gnd.t77 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X271 a_n6308_8799.t8 a_n2408_n452.t83 a_n2318_8322.t10 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X272 a_n2408_n452.t32 a_n2408_n452.t31 a_n2140_13878.t2 vdd.t103 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X273 gnd.t65 commonsourceibias.t91 CSoutput.t14 gnd.t64 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X274 commonsourceibias.t13 commonsourceibias.t12 gnd.t272 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 a_n6308_8799.t34 plus.t25 a_n2903_n3924.t10 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X276 vdd.t202 a_n6308_8799.t81 CSoutput.t35 vdd.t78 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X277 CSoutput.t34 a_n6308_8799.t82 vdd.t179 vdd.t84 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X278 vdd.t180 a_n6308_8799.t83 CSoutput.t33 vdd.t145 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X279 diffpairibias.t3 diffpairibias.t2 gnd.t47 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X280 a_n2318_8322.t9 a_n2408_n452.t84 a_n6308_8799.t5 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X281 a_n2903_n3924.t9 plus.t26 a_n6308_8799.t23 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X282 commonsourceibias.t11 commonsourceibias.t10 gnd.t242 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X283 gnd.t69 commonsourceibias.t92 CSoutput.t16 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X284 CSoutput.t116 a_n2318_8322.t24 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X285 diffpairibias.t1 diffpairibias.t0 gnd.t53 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X286 a_n2903_n3924.t8 plus.t27 a_n6308_8799.t31 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X287 CSoutput.t89 commonsourceibias.t93 gnd.t277 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X288 vdd.t1 CSoutput.t117 output.t4 gnd.t86 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X289 vdd.t101 a_n2408_n452.t85 a_n2140_13878.t18 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X290 vdd.t17 vdd.t14 vdd.t16 vdd.t15 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X291 a_n6308_8799.t16 plus.t28 a_n2903_n3924.t7 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X292 vdd.t13 vdd.t10 vdd.t12 vdd.t11 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X293 vdd.t195 a_n6308_8799.t84 CSoutput.t32 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X294 gnd.t121 gnd.t118 gnd.t120 gnd.t119 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X295 a_n2903_n3924.t50 minus.t27 a_n2408_n452.t51 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X296 CSoutput.t6 commonsourceibias.t94 gnd.t26 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X297 CSoutput.t31 a_n6308_8799.t85 vdd.t196 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X298 commonsourceibias.t9 commonsourceibias.t8 gnd.t8 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X299 a_n2318_8322.t8 a_n2408_n452.t86 a_n6308_8799.t11 vdd.t99 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X300 CSoutput.t21 commonsourceibias.t95 gnd.t105 gnd.t104 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X301 a_n2408_n452.t50 minus.t28 a_n2903_n3924.t49 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X302 vdd.t87 a_n6308_8799.t86 CSoutput.t30 vdd.t86 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X303 gnd.t284 commonsourceibias.t6 commonsourceibias.t7 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X304 commonsourceibias.t5 commonsourceibias.t4 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X305 vdd.t9 vdd.t6 vdd.t8 vdd.t7 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X306 a_n2318_8322.t0 a_n2408_n452.t87 vdd.t96 vdd.t95 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X307 a_n2140_13878.t1 a_n2408_n452.t25 a_n2408_n452.t26 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X308 vdd.t88 a_n6308_8799.t87 CSoutput.t29 vdd.t78 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X309 minus.t0 gnd.t115 gnd.t117 gnd.t116 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X310 commonsourceibias.t3 commonsourceibias.t2 gnd.t61 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X311 a_n2408_n452.t24 a_n2408_n452.t23 a_n2140_13878.t0 vdd.t93 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X312 vdd.t5 vdd.t2 vdd.t4 vdd.t3 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X313 gnd.t34 commonsourceibias.t0 commonsourceibias.t1 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X314 a_n2903_n3924.t36 diffpairibias.t23 gnd.t228 gnd.t227 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X315 gnd.t114 gnd.t111 gnd.t113 gnd.t112 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
R0 a_n2408_n452.n95 a_n2408_n452.t73 512.366
R1 a_n2408_n452.n85 a_n2408_n452.t64 512.366
R2 a_n2408_n452.n96 a_n2408_n452.t56 512.366
R3 a_n2408_n452.n93 a_n2408_n452.t81 512.366
R4 a_n2408_n452.n86 a_n2408_n452.t70 512.366
R5 a_n2408_n452.n94 a_n2408_n452.t69 512.366
R6 a_n2408_n452.n91 a_n2408_n452.t77 512.366
R7 a_n2408_n452.n87 a_n2408_n452.t63 512.366
R8 a_n2408_n452.n92 a_n2408_n452.t62 512.366
R9 a_n2408_n452.n89 a_n2408_n452.t66 512.366
R10 a_n2408_n452.n88 a_n2408_n452.t75 512.366
R11 a_n2408_n452.n90 a_n2408_n452.t87 512.366
R12 a_n2408_n452.n36 a_n2408_n452.t86 533.335
R13 a_n2408_n452.n101 a_n2408_n452.t67 512.366
R14 a_n2408_n452.n67 a_n2408_n452.t71 512.366
R15 a_n2408_n452.n100 a_n2408_n452.t61 512.366
R16 a_n2408_n452.n99 a_n2408_n452.t76 512.366
R17 a_n2408_n452.n68 a_n2408_n452.t83 512.366
R18 a_n2408_n452.n98 a_n2408_n452.t84 512.366
R19 a_n2408_n452.n35 a_n2408_n452.t25 533.335
R20 a_n2408_n452.n102 a_n2408_n452.t15 512.366
R21 a_n2408_n452.n65 a_n2408_n452.t9 512.366
R22 a_n2408_n452.n31 a_n2408_n452.t11 533.335
R23 a_n2408_n452.n117 a_n2408_n452.t7 512.366
R24 a_n2408_n452.n66 a_n2408_n452.t31 512.366
R25 a_n2408_n452.n116 a_n2408_n452.t29 512.366
R26 a_n2408_n452.n115 a_n2408_n452.t13 512.366
R27 a_n2408_n452.n49 a_n2408_n452.t17 533.335
R28 a_n2408_n452.n79 a_n2408_n452.t19 512.366
R29 a_n2408_n452.n80 a_n2408_n452.t23 512.366
R30 a_n2408_n452.n81 a_n2408_n452.t37 512.366
R31 a_n2408_n452.n82 a_n2408_n452.t27 512.366
R32 a_n2408_n452.n72 a_n2408_n452.t33 512.366
R33 a_n2408_n452.n83 a_n2408_n452.t21 512.366
R34 a_n2408_n452.n42 a_n2408_n452.t82 533.335
R35 a_n2408_n452.n74 a_n2408_n452.t60 512.366
R36 a_n2408_n452.n75 a_n2408_n452.t80 512.366
R37 a_n2408_n452.n76 a_n2408_n452.t79 512.366
R38 a_n2408_n452.n77 a_n2408_n452.t57 512.366
R39 a_n2408_n452.n73 a_n2408_n452.t65 512.366
R40 a_n2408_n452.n78 a_n2408_n452.t74 512.366
R41 a_n2408_n452.n5 a_n2408_n452.n63 70.1674
R42 a_n2408_n452.n7 a_n2408_n452.n61 70.1674
R43 a_n2408_n452.n9 a_n2408_n452.n59 70.1674
R44 a_n2408_n452.n12 a_n2408_n452.n57 70.1674
R45 a_n2408_n452.n41 a_n2408_n452.n21 70.1674
R46 a_n2408_n452.n34 a_n2408_n452.n24 77.6622
R47 a_n2408_n452.n115 a_n2408_n452.n34 5.97853
R48 a_n2408_n452.n33 a_n2408_n452.n26 77.6622
R49 a_n2408_n452.n26 a_n2408_n452.n32 72.3034
R50 a_n2408_n452.n117 a_n2408_n452.n31 20.9683
R51 a_n2408_n452.n25 a_n2408_n452.n31 70.1674
R52 a_n2408_n452.n64 a_n2408_n452.n65 16.6962
R53 a_n2408_n452.n35 a_n2408_n452.n24 70.1674
R54 a_n2408_n452.n102 a_n2408_n452.n35 20.9683
R55 a_n2408_n452.n24 a_n2408_n452.n64 72.3034
R56 a_n2408_n452.n98 a_n2408_n452.n41 20.9683
R57 a_n2408_n452.n22 a_n2408_n452.n40 72.3034
R58 a_n2408_n452.n40 a_n2408_n452.n68 16.6962
R59 a_n2408_n452.n39 a_n2408_n452.n22 77.6622
R60 a_n2408_n452.n99 a_n2408_n452.n39 5.97853
R61 a_n2408_n452.n38 a_n2408_n452.n20 77.6622
R62 a_n2408_n452.n20 a_n2408_n452.n37 72.3034
R63 a_n2408_n452.n101 a_n2408_n452.n36 20.9683
R64 a_n2408_n452.n23 a_n2408_n452.n36 70.1674
R65 a_n2408_n452.n14 a_n2408_n452.n55 70.1674
R66 a_n2408_n452.n17 a_n2408_n452.n48 70.1674
R67 a_n2408_n452.n78 a_n2408_n452.n48 20.9683
R68 a_n2408_n452.n47 a_n2408_n452.n18 72.3034
R69 a_n2408_n452.n47 a_n2408_n452.n73 16.6962
R70 a_n2408_n452.n18 a_n2408_n452.n46 77.6622
R71 a_n2408_n452.n77 a_n2408_n452.n46 5.97853
R72 a_n2408_n452.n45 a_n2408_n452.n19 77.6622
R73 a_n2408_n452.n19 a_n2408_n452.n44 72.3034
R74 a_n2408_n452.n74 a_n2408_n452.n42 20.9683
R75 a_n2408_n452.n43 a_n2408_n452.n42 70.1674
R76 a_n2408_n452.n83 a_n2408_n452.n55 20.9683
R77 a_n2408_n452.n54 a_n2408_n452.n15 72.3034
R78 a_n2408_n452.n54 a_n2408_n452.n72 16.6962
R79 a_n2408_n452.n15 a_n2408_n452.n53 77.6622
R80 a_n2408_n452.n82 a_n2408_n452.n53 5.97853
R81 a_n2408_n452.n52 a_n2408_n452.n16 77.6622
R82 a_n2408_n452.n16 a_n2408_n452.n51 72.3034
R83 a_n2408_n452.n79 a_n2408_n452.n49 20.9683
R84 a_n2408_n452.n50 a_n2408_n452.n49 70.1674
R85 a_n2408_n452.n90 a_n2408_n452.n57 20.9683
R86 a_n2408_n452.n56 a_n2408_n452.n13 75.0448
R87 a_n2408_n452.n56 a_n2408_n452.n88 11.2134
R88 a_n2408_n452.n13 a_n2408_n452.n89 161.3
R89 a_n2408_n452.n92 a_n2408_n452.n59 20.9683
R90 a_n2408_n452.n58 a_n2408_n452.n10 75.0448
R91 a_n2408_n452.n58 a_n2408_n452.n87 11.2134
R92 a_n2408_n452.n10 a_n2408_n452.n91 161.3
R93 a_n2408_n452.n94 a_n2408_n452.n61 20.9683
R94 a_n2408_n452.n60 a_n2408_n452.n8 75.0448
R95 a_n2408_n452.n60 a_n2408_n452.n86 11.2134
R96 a_n2408_n452.n8 a_n2408_n452.n93 161.3
R97 a_n2408_n452.n96 a_n2408_n452.n63 20.9683
R98 a_n2408_n452.n62 a_n2408_n452.n6 75.0448
R99 a_n2408_n452.n62 a_n2408_n452.n85 11.2134
R100 a_n2408_n452.n6 a_n2408_n452.n95 161.3
R101 a_n2408_n452.n3 a_n2408_n452.n112 81.3764
R102 a_n2408_n452.n4 a_n2408_n452.n106 81.3764
R103 a_n2408_n452.n0 a_n2408_n452.n103 81.3764
R104 a_n2408_n452.n3 a_n2408_n452.n113 80.9324
R105 a_n2408_n452.n2 a_n2408_n452.n114 80.9324
R106 a_n2408_n452.n2 a_n2408_n452.n111 80.9324
R107 a_n2408_n452.n2 a_n2408_n452.n110 80.9324
R108 a_n2408_n452.n1 a_n2408_n452.n109 80.9324
R109 a_n2408_n452.n4 a_n2408_n452.n107 80.9324
R110 a_n2408_n452.n0 a_n2408_n452.n108 80.9324
R111 a_n2408_n452.n0 a_n2408_n452.n105 80.9324
R112 a_n2408_n452.n0 a_n2408_n452.n104 80.9324
R113 a_n2408_n452.n29 a_n2408_n452.t26 74.6477
R114 a_n2408_n452.n27 a_n2408_n452.t18 74.6477
R115 a_n2408_n452.n30 a_n2408_n452.t12 74.2899
R116 a_n2408_n452.n28 a_n2408_n452.t36 74.2897
R117 a_n2408_n452.n29 a_n2408_n452.n119 70.6783
R118 a_n2408_n452.n29 a_n2408_n452.n120 70.6783
R119 a_n2408_n452.n28 a_n2408_n452.n71 70.6783
R120 a_n2408_n452.n27 a_n2408_n452.n70 70.6783
R121 a_n2408_n452.n27 a_n2408_n452.n69 70.6783
R122 a_n2408_n452.n121 a_n2408_n452.n30 70.6782
R123 a_n2408_n452.n95 a_n2408_n452.n85 48.2005
R124 a_n2408_n452.t78 a_n2408_n452.n63 533.335
R125 a_n2408_n452.n93 a_n2408_n452.n86 48.2005
R126 a_n2408_n452.t85 a_n2408_n452.n61 533.335
R127 a_n2408_n452.n91 a_n2408_n452.n87 48.2005
R128 a_n2408_n452.t72 a_n2408_n452.n59 533.335
R129 a_n2408_n452.n89 a_n2408_n452.n88 48.2005
R130 a_n2408_n452.t68 a_n2408_n452.n57 533.335
R131 a_n2408_n452.n100 a_n2408_n452.n99 48.2005
R132 a_n2408_n452.n41 a_n2408_n452.t58 533.335
R133 a_n2408_n452.n116 a_n2408_n452.n115 48.2005
R134 a_n2408_n452.n82 a_n2408_n452.n81 48.2005
R135 a_n2408_n452.t35 a_n2408_n452.n55 533.335
R136 a_n2408_n452.n77 a_n2408_n452.n76 48.2005
R137 a_n2408_n452.t59 a_n2408_n452.n48 533.335
R138 a_n2408_n452.n37 a_n2408_n452.n67 16.6962
R139 a_n2408_n452.n98 a_n2408_n452.n40 27.6507
R140 a_n2408_n452.n102 a_n2408_n452.n64 27.6507
R141 a_n2408_n452.n32 a_n2408_n452.n66 16.6962
R142 a_n2408_n452.n80 a_n2408_n452.n51 16.6962
R143 a_n2408_n452.n83 a_n2408_n452.n54 27.6507
R144 a_n2408_n452.n75 a_n2408_n452.n44 16.6962
R145 a_n2408_n452.n78 a_n2408_n452.n47 27.6507
R146 a_n2408_n452.n38 a_n2408_n452.n67 41.7634
R147 a_n2408_n452.n33 a_n2408_n452.n66 41.7634
R148 a_n2408_n452.n80 a_n2408_n452.n52 41.7634
R149 a_n2408_n452.n75 a_n2408_n452.n45 41.7634
R150 a_n2408_n452.n1 a_n2408_n452.n0 32.6799
R151 a_n2408_n452.n96 a_n2408_n452.n62 35.3134
R152 a_n2408_n452.n94 a_n2408_n452.n60 35.3134
R153 a_n2408_n452.n92 a_n2408_n452.n58 35.3134
R154 a_n2408_n452.n90 a_n2408_n452.n56 35.3134
R155 a_n2408_n452.n24 a_n2408_n452.n2 23.891
R156 a_n2408_n452.n43 a_n2408_n452.n11 12.705
R157 a_n2408_n452.n21 a_n2408_n452.n97 12.5005
R158 a_n2408_n452.n38 a_n2408_n452.n100 5.97853
R159 a_n2408_n452.n39 a_n2408_n452.n68 41.7634
R160 a_n2408_n452.n33 a_n2408_n452.n116 5.97853
R161 a_n2408_n452.n34 a_n2408_n452.n65 41.7634
R162 a_n2408_n452.n81 a_n2408_n452.n52 5.97853
R163 a_n2408_n452.n72 a_n2408_n452.n53 41.7634
R164 a_n2408_n452.n76 a_n2408_n452.n45 5.97853
R165 a_n2408_n452.n73 a_n2408_n452.n46 41.7634
R166 a_n2408_n452.n118 a_n2408_n452.n25 11.1956
R167 a_n2408_n452.n101 a_n2408_n452.n37 27.6507
R168 a_n2408_n452.n117 a_n2408_n452.n32 27.6507
R169 a_n2408_n452.n51 a_n2408_n452.n79 27.6507
R170 a_n2408_n452.n44 a_n2408_n452.n74 27.6507
R171 a_n2408_n452.n84 a_n2408_n452.n28 9.85898
R172 a_n2408_n452.n97 a_n2408_n452.n5 8.73345
R173 a_n2408_n452.n13 a_n2408_n452.n11 8.73345
R174 a_n2408_n452.n84 a_n2408_n452.n14 7.36035
R175 a_n2408_n452.n30 a_n2408_n452.n118 6.01559
R176 a_n2408_n452.n97 a_n2408_n452.n84 5.3452
R177 a_n2408_n452.n24 a_n2408_n452.n23 4.01186
R178 a_n2408_n452.n50 a_n2408_n452.n17 4.01186
R179 a_n2408_n452.n119 a_n2408_n452.t10 3.61217
R180 a_n2408_n452.n119 a_n2408_n452.t16 3.61217
R181 a_n2408_n452.n120 a_n2408_n452.t30 3.61217
R182 a_n2408_n452.n120 a_n2408_n452.t14 3.61217
R183 a_n2408_n452.n71 a_n2408_n452.t34 3.61217
R184 a_n2408_n452.n71 a_n2408_n452.t22 3.61217
R185 a_n2408_n452.n70 a_n2408_n452.t38 3.61217
R186 a_n2408_n452.n70 a_n2408_n452.t28 3.61217
R187 a_n2408_n452.n69 a_n2408_n452.t20 3.61217
R188 a_n2408_n452.n69 a_n2408_n452.t24 3.61217
R189 a_n2408_n452.t8 a_n2408_n452.n121 3.61217
R190 a_n2408_n452.n121 a_n2408_n452.t32 3.61217
R191 a_n2408_n452.n112 a_n2408_n452.t51 2.82907
R192 a_n2408_n452.n112 a_n2408_n452.t50 2.82907
R193 a_n2408_n452.n113 a_n2408_n452.t3 2.82907
R194 a_n2408_n452.n113 a_n2408_n452.t39 2.82907
R195 a_n2408_n452.n114 a_n2408_n452.t43 2.82907
R196 a_n2408_n452.n114 a_n2408_n452.t47 2.82907
R197 a_n2408_n452.n111 a_n2408_n452.t55 2.82907
R198 a_n2408_n452.n111 a_n2408_n452.t44 2.82907
R199 a_n2408_n452.n110 a_n2408_n452.t40 2.82907
R200 a_n2408_n452.n110 a_n2408_n452.t0 2.82907
R201 a_n2408_n452.n109 a_n2408_n452.t42 2.82907
R202 a_n2408_n452.n109 a_n2408_n452.t46 2.82907
R203 a_n2408_n452.n106 a_n2408_n452.t49 2.82907
R204 a_n2408_n452.n106 a_n2408_n452.t2 2.82907
R205 a_n2408_n452.n107 a_n2408_n452.t45 2.82907
R206 a_n2408_n452.n107 a_n2408_n452.t54 2.82907
R207 a_n2408_n452.n108 a_n2408_n452.t41 2.82907
R208 a_n2408_n452.n108 a_n2408_n452.t52 2.82907
R209 a_n2408_n452.n105 a_n2408_n452.t4 2.82907
R210 a_n2408_n452.n105 a_n2408_n452.t1 2.82907
R211 a_n2408_n452.n104 a_n2408_n452.t6 2.82907
R212 a_n2408_n452.n104 a_n2408_n452.t5 2.82907
R213 a_n2408_n452.n103 a_n2408_n452.t53 2.82907
R214 a_n2408_n452.n103 a_n2408_n452.t48 2.82907
R215 a_n2408_n452.n0 a_n2408_n452.n4 1.3324
R216 a_n2408_n452.n118 a_n2408_n452.n11 1.30542
R217 a_n2408_n452.n24 a_n2408_n452.n26 1.09898
R218 a_n2408_n452.n30 a_n2408_n452.n29 1.07378
R219 a_n2408_n452.n28 a_n2408_n452.n27 1.07378
R220 a_n2408_n452.n8 a_n2408_n452.n9 1.04595
R221 a_n2408_n452.n26 a_n2408_n452.n25 0.94747
R222 a_n2408_n452.n2 a_n2408_n452.n3 0.888431
R223 a_n2408_n452.n2 a_n2408_n452.n1 0.888431
R224 a_n2408_n452.n22 a_n2408_n452.n20 0.758076
R225 a_n2408_n452.n22 a_n2408_n452.n21 0.758076
R226 a_n2408_n452.n19 a_n2408_n452.n18 0.758076
R227 a_n2408_n452.n18 a_n2408_n452.n17 0.758076
R228 a_n2408_n452.n16 a_n2408_n452.n15 0.758076
R229 a_n2408_n452.n15 a_n2408_n452.n14 0.758076
R230 a_n2408_n452.n13 a_n2408_n452.n12 0.758076
R231 a_n2408_n452.n10 a_n2408_n452.n9 0.758076
R232 a_n2408_n452.n8 a_n2408_n452.n7 0.758076
R233 a_n2408_n452.n6 a_n2408_n452.n5 0.758076
R234 a_n2408_n452.n10 a_n2408_n452.n12 0.67853
R235 a_n2408_n452.n6 a_n2408_n452.n7 0.67853
R236 a_n2408_n452.n50 a_n2408_n452.n16 0.568682
R237 a_n2408_n452.n43 a_n2408_n452.n19 0.568682
R238 a_n2408_n452.n20 a_n2408_n452.n23 0.568682
R239 a_n2140_13878.n21 a_n2140_13878.n20 98.9632
R240 a_n2140_13878.n2 a_n2140_13878.n0 98.7517
R241 a_n2140_13878.n18 a_n2140_13878.n17 98.6055
R242 a_n2140_13878.n20 a_n2140_13878.n19 98.6055
R243 a_n2140_13878.n6 a_n2140_13878.n5 98.6055
R244 a_n2140_13878.n4 a_n2140_13878.n3 98.6055
R245 a_n2140_13878.n2 a_n2140_13878.n1 98.6055
R246 a_n2140_13878.n16 a_n2140_13878.n15 98.6054
R247 a_n2140_13878.n8 a_n2140_13878.t23 74.6477
R248 a_n2140_13878.n13 a_n2140_13878.t20 74.2899
R249 a_n2140_13878.n10 a_n2140_13878.t19 74.2899
R250 a_n2140_13878.n9 a_n2140_13878.t18 74.2899
R251 a_n2140_13878.n12 a_n2140_13878.n11 70.6783
R252 a_n2140_13878.n8 a_n2140_13878.n7 70.6783
R253 a_n2140_13878.n14 a_n2140_13878.n6 14.2849
R254 a_n2140_13878.n16 a_n2140_13878.n14 11.9339
R255 a_n2140_13878.n14 a_n2140_13878.n13 6.95632
R256 a_n2140_13878.n15 a_n2140_13878.t6 3.61217
R257 a_n2140_13878.n15 a_n2140_13878.t7 3.61217
R258 a_n2140_13878.n17 a_n2140_13878.t13 3.61217
R259 a_n2140_13878.n17 a_n2140_13878.t14 3.61217
R260 a_n2140_13878.n19 a_n2140_13878.t0 3.61217
R261 a_n2140_13878.n19 a_n2140_13878.t8 3.61217
R262 a_n2140_13878.n11 a_n2140_13878.t22 3.61217
R263 a_n2140_13878.n11 a_n2140_13878.t21 3.61217
R264 a_n2140_13878.n7 a_n2140_13878.t16 3.61217
R265 a_n2140_13878.n7 a_n2140_13878.t17 3.61217
R266 a_n2140_13878.n5 a_n2140_13878.t9 3.61217
R267 a_n2140_13878.n5 a_n2140_13878.t1 3.61217
R268 a_n2140_13878.n3 a_n2140_13878.t12 3.61217
R269 a_n2140_13878.n3 a_n2140_13878.t3 3.61217
R270 a_n2140_13878.n1 a_n2140_13878.t2 3.61217
R271 a_n2140_13878.n1 a_n2140_13878.t4 3.61217
R272 a_n2140_13878.n0 a_n2140_13878.t10 3.61217
R273 a_n2140_13878.n0 a_n2140_13878.t5 3.61217
R274 a_n2140_13878.n21 a_n2140_13878.t11 3.61217
R275 a_n2140_13878.t15 a_n2140_13878.n21 3.61217
R276 a_n2140_13878.n9 a_n2140_13878.n8 0.358259
R277 a_n2140_13878.n12 a_n2140_13878.n10 0.358259
R278 a_n2140_13878.n13 a_n2140_13878.n12 0.358259
R279 a_n2140_13878.n20 a_n2140_13878.n18 0.358259
R280 a_n2140_13878.n18 a_n2140_13878.n16 0.358259
R281 a_n2140_13878.n4 a_n2140_13878.n2 0.146627
R282 a_n2140_13878.n6 a_n2140_13878.n4 0.146627
R283 a_n2140_13878.n10 a_n2140_13878.n9 0.101793
R284 vdd.n291 vdd.n255 756.745
R285 vdd.n244 vdd.n208 756.745
R286 vdd.n201 vdd.n165 756.745
R287 vdd.n154 vdd.n118 756.745
R288 vdd.n112 vdd.n76 756.745
R289 vdd.n65 vdd.n29 756.745
R290 vdd.n1468 vdd.n1432 756.745
R291 vdd.n1515 vdd.n1479 756.745
R292 vdd.n1378 vdd.n1342 756.745
R293 vdd.n1425 vdd.n1389 756.745
R294 vdd.n1289 vdd.n1253 756.745
R295 vdd.n1336 vdd.n1300 756.745
R296 vdd.n1043 vdd.t14 640.208
R297 vdd.n771 vdd.t48 640.208
R298 vdd.n1063 vdd.t29 640.208
R299 vdd.n762 vdd.t66 640.208
R300 vdd.n662 vdd.t35 640.208
R301 vdd.n2318 vdd.t60 640.208
R302 vdd.n622 vdd.t69 640.208
R303 vdd.n2315 vdd.t52 640.208
R304 vdd.n589 vdd.t10 640.208
R305 vdd.n833 vdd.t56 640.208
R306 vdd.n1682 vdd.t2 592.009
R307 vdd.n1720 vdd.t32 592.009
R308 vdd.n1616 vdd.t42 592.009
R309 vdd.n1883 vdd.t22 592.009
R310 vdd.n980 vdd.t45 592.009
R311 vdd.n940 vdd.t63 592.009
R312 vdd.n3000 vdd.t75 592.009
R313 vdd.n405 vdd.t72 592.009
R314 vdd.n365 vdd.t6 592.009
R315 vdd.n557 vdd.t26 592.009
R316 vdd.n2896 vdd.t39 592.009
R317 vdd.n2803 vdd.t18 592.009
R318 vdd.n292 vdd.n291 585
R319 vdd.n290 vdd.n257 585
R320 vdd.n289 vdd.n288 585
R321 vdd.n260 vdd.n258 585
R322 vdd.n283 vdd.n282 585
R323 vdd.n281 vdd.n280 585
R324 vdd.n264 vdd.n263 585
R325 vdd.n275 vdd.n274 585
R326 vdd.n273 vdd.n272 585
R327 vdd.n268 vdd.n267 585
R328 vdd.n245 vdd.n244 585
R329 vdd.n243 vdd.n210 585
R330 vdd.n242 vdd.n241 585
R331 vdd.n213 vdd.n211 585
R332 vdd.n236 vdd.n235 585
R333 vdd.n234 vdd.n233 585
R334 vdd.n217 vdd.n216 585
R335 vdd.n228 vdd.n227 585
R336 vdd.n226 vdd.n225 585
R337 vdd.n221 vdd.n220 585
R338 vdd.n202 vdd.n201 585
R339 vdd.n200 vdd.n167 585
R340 vdd.n199 vdd.n198 585
R341 vdd.n170 vdd.n168 585
R342 vdd.n193 vdd.n192 585
R343 vdd.n191 vdd.n190 585
R344 vdd.n174 vdd.n173 585
R345 vdd.n185 vdd.n184 585
R346 vdd.n183 vdd.n182 585
R347 vdd.n178 vdd.n177 585
R348 vdd.n155 vdd.n154 585
R349 vdd.n153 vdd.n120 585
R350 vdd.n152 vdd.n151 585
R351 vdd.n123 vdd.n121 585
R352 vdd.n146 vdd.n145 585
R353 vdd.n144 vdd.n143 585
R354 vdd.n127 vdd.n126 585
R355 vdd.n138 vdd.n137 585
R356 vdd.n136 vdd.n135 585
R357 vdd.n131 vdd.n130 585
R358 vdd.n113 vdd.n112 585
R359 vdd.n111 vdd.n78 585
R360 vdd.n110 vdd.n109 585
R361 vdd.n81 vdd.n79 585
R362 vdd.n104 vdd.n103 585
R363 vdd.n102 vdd.n101 585
R364 vdd.n85 vdd.n84 585
R365 vdd.n96 vdd.n95 585
R366 vdd.n94 vdd.n93 585
R367 vdd.n89 vdd.n88 585
R368 vdd.n66 vdd.n65 585
R369 vdd.n64 vdd.n31 585
R370 vdd.n63 vdd.n62 585
R371 vdd.n34 vdd.n32 585
R372 vdd.n57 vdd.n56 585
R373 vdd.n55 vdd.n54 585
R374 vdd.n38 vdd.n37 585
R375 vdd.n49 vdd.n48 585
R376 vdd.n47 vdd.n46 585
R377 vdd.n42 vdd.n41 585
R378 vdd.n1469 vdd.n1468 585
R379 vdd.n1467 vdd.n1434 585
R380 vdd.n1466 vdd.n1465 585
R381 vdd.n1437 vdd.n1435 585
R382 vdd.n1460 vdd.n1459 585
R383 vdd.n1458 vdd.n1457 585
R384 vdd.n1441 vdd.n1440 585
R385 vdd.n1452 vdd.n1451 585
R386 vdd.n1450 vdd.n1449 585
R387 vdd.n1445 vdd.n1444 585
R388 vdd.n1516 vdd.n1515 585
R389 vdd.n1514 vdd.n1481 585
R390 vdd.n1513 vdd.n1512 585
R391 vdd.n1484 vdd.n1482 585
R392 vdd.n1507 vdd.n1506 585
R393 vdd.n1505 vdd.n1504 585
R394 vdd.n1488 vdd.n1487 585
R395 vdd.n1499 vdd.n1498 585
R396 vdd.n1497 vdd.n1496 585
R397 vdd.n1492 vdd.n1491 585
R398 vdd.n1379 vdd.n1378 585
R399 vdd.n1377 vdd.n1344 585
R400 vdd.n1376 vdd.n1375 585
R401 vdd.n1347 vdd.n1345 585
R402 vdd.n1370 vdd.n1369 585
R403 vdd.n1368 vdd.n1367 585
R404 vdd.n1351 vdd.n1350 585
R405 vdd.n1362 vdd.n1361 585
R406 vdd.n1360 vdd.n1359 585
R407 vdd.n1355 vdd.n1354 585
R408 vdd.n1426 vdd.n1425 585
R409 vdd.n1424 vdd.n1391 585
R410 vdd.n1423 vdd.n1422 585
R411 vdd.n1394 vdd.n1392 585
R412 vdd.n1417 vdd.n1416 585
R413 vdd.n1415 vdd.n1414 585
R414 vdd.n1398 vdd.n1397 585
R415 vdd.n1409 vdd.n1408 585
R416 vdd.n1407 vdd.n1406 585
R417 vdd.n1402 vdd.n1401 585
R418 vdd.n1290 vdd.n1289 585
R419 vdd.n1288 vdd.n1255 585
R420 vdd.n1287 vdd.n1286 585
R421 vdd.n1258 vdd.n1256 585
R422 vdd.n1281 vdd.n1280 585
R423 vdd.n1279 vdd.n1278 585
R424 vdd.n1262 vdd.n1261 585
R425 vdd.n1273 vdd.n1272 585
R426 vdd.n1271 vdd.n1270 585
R427 vdd.n1266 vdd.n1265 585
R428 vdd.n1337 vdd.n1336 585
R429 vdd.n1335 vdd.n1302 585
R430 vdd.n1334 vdd.n1333 585
R431 vdd.n1305 vdd.n1303 585
R432 vdd.n1328 vdd.n1327 585
R433 vdd.n1326 vdd.n1325 585
R434 vdd.n1309 vdd.n1308 585
R435 vdd.n1320 vdd.n1319 585
R436 vdd.n1318 vdd.n1317 585
R437 vdd.n1313 vdd.n1312 585
R438 vdd.n3116 vdd.n330 515.122
R439 vdd.n2998 vdd.n328 515.122
R440 vdd.n515 vdd.n478 515.122
R441 vdd.n2934 vdd.n479 515.122
R442 vdd.n1878 vdd.n1227 515.122
R443 vdd.n1881 vdd.n1880 515.122
R444 vdd.n1589 vdd.n1553 515.122
R445 vdd.n1785 vdd.n1554 515.122
R446 vdd.n269 vdd.t184 329.043
R447 vdd.n222 vdd.t170 329.043
R448 vdd.n179 vdd.t85 329.043
R449 vdd.n132 vdd.t163 329.043
R450 vdd.n90 vdd.t179 329.043
R451 vdd.n43 vdd.t172 329.043
R452 vdd.n1446 vdd.t200 329.043
R453 vdd.n1493 vdd.t146 329.043
R454 vdd.n1356 vdd.t142 329.043
R455 vdd.n1403 vdd.t150 329.043
R456 vdd.n1267 vdd.t171 329.043
R457 vdd.n1314 vdd.t180 329.043
R458 vdd.n1682 vdd.t5 319.788
R459 vdd.n1720 vdd.t34 319.788
R460 vdd.n1616 vdd.t44 319.788
R461 vdd.n1883 vdd.t24 319.788
R462 vdd.n980 vdd.t46 319.788
R463 vdd.n940 vdd.t64 319.788
R464 vdd.n3000 vdd.t76 319.788
R465 vdd.n405 vdd.t73 319.788
R466 vdd.n365 vdd.t8 319.788
R467 vdd.n557 vdd.t28 319.788
R468 vdd.n2896 vdd.t41 319.788
R469 vdd.n2803 vdd.t21 319.788
R470 vdd.n1683 vdd.t4 303.69
R471 vdd.n1721 vdd.t33 303.69
R472 vdd.n1617 vdd.t43 303.69
R473 vdd.n1884 vdd.t25 303.69
R474 vdd.n981 vdd.t47 303.69
R475 vdd.n941 vdd.t65 303.69
R476 vdd.n3001 vdd.t77 303.69
R477 vdd.n406 vdd.t74 303.69
R478 vdd.n366 vdd.t9 303.69
R479 vdd.n558 vdd.t27 303.69
R480 vdd.n2897 vdd.t40 303.69
R481 vdd.n2804 vdd.t20 303.69
R482 vdd.n2550 vdd.n717 291.221
R483 vdd.n2764 vdd.n599 291.221
R484 vdd.n2701 vdd.n596 291.221
R485 vdd.n2482 vdd.n2481 291.221
R486 vdd.n2278 vdd.n759 291.221
R487 vdd.n2209 vdd.n2208 291.221
R488 vdd.n1099 vdd.n1098 291.221
R489 vdd.n2029 vdd.n865 291.221
R490 vdd.n2680 vdd.n597 291.221
R491 vdd.n2767 vdd.n2766 291.221
R492 vdd.n2386 vdd.n2312 291.221
R493 vdd.n2554 vdd.n721 291.221
R494 vdd.n2206 vdd.n769 291.221
R495 vdd.n767 vdd.n741 291.221
R496 vdd.n1177 vdd.n906 291.221
R497 vdd.n2033 vdd.n870 291.221
R498 vdd.n2682 vdd.n597 185
R499 vdd.n2765 vdd.n597 185
R500 vdd.n2684 vdd.n2683 185
R501 vdd.n2683 vdd.n595 185
R502 vdd.n2685 vdd.n629 185
R503 vdd.n2695 vdd.n629 185
R504 vdd.n2686 vdd.n638 185
R505 vdd.n638 vdd.n636 185
R506 vdd.n2688 vdd.n2687 185
R507 vdd.n2689 vdd.n2688 185
R508 vdd.n2641 vdd.n637 185
R509 vdd.n637 vdd.n633 185
R510 vdd.n2640 vdd.n2639 185
R511 vdd.n2639 vdd.n2638 185
R512 vdd.n640 vdd.n639 185
R513 vdd.n641 vdd.n640 185
R514 vdd.n2631 vdd.n2630 185
R515 vdd.n2632 vdd.n2631 185
R516 vdd.n2629 vdd.n650 185
R517 vdd.n650 vdd.n647 185
R518 vdd.n2628 vdd.n2627 185
R519 vdd.n2627 vdd.n2626 185
R520 vdd.n652 vdd.n651 185
R521 vdd.n660 vdd.n652 185
R522 vdd.n2619 vdd.n2618 185
R523 vdd.n2620 vdd.n2619 185
R524 vdd.n2616 vdd.n661 185
R525 vdd.n668 vdd.n661 185
R526 vdd.n2615 vdd.n2614 185
R527 vdd.n2614 vdd.n2613 185
R528 vdd.n664 vdd.n663 185
R529 vdd.n665 vdd.n664 185
R530 vdd.n2606 vdd.n2605 185
R531 vdd.n2607 vdd.n2606 185
R532 vdd.n2604 vdd.n675 185
R533 vdd.n675 vdd.n672 185
R534 vdd.n2603 vdd.n2602 185
R535 vdd.n2602 vdd.n2601 185
R536 vdd.n677 vdd.n676 185
R537 vdd.n685 vdd.n677 185
R538 vdd.n2594 vdd.n2593 185
R539 vdd.n2595 vdd.n2594 185
R540 vdd.n2592 vdd.n686 185
R541 vdd.n691 vdd.n686 185
R542 vdd.n2591 vdd.n2590 185
R543 vdd.n2590 vdd.n2589 185
R544 vdd.n688 vdd.n687 185
R545 vdd.n2461 vdd.n688 185
R546 vdd.n2582 vdd.n2581 185
R547 vdd.n2583 vdd.n2582 185
R548 vdd.n2580 vdd.n698 185
R549 vdd.n698 vdd.n695 185
R550 vdd.n2579 vdd.n2578 185
R551 vdd.n2578 vdd.n2577 185
R552 vdd.n700 vdd.n699 185
R553 vdd.n701 vdd.n700 185
R554 vdd.n2570 vdd.n2569 185
R555 vdd.n2571 vdd.n2570 185
R556 vdd.n2568 vdd.n710 185
R557 vdd.n710 vdd.n707 185
R558 vdd.n2567 vdd.n2566 185
R559 vdd.n2566 vdd.n2565 185
R560 vdd.n712 vdd.n711 185
R561 vdd.n2476 vdd.n712 185
R562 vdd.n2558 vdd.n2557 185
R563 vdd.n2559 vdd.n2558 185
R564 vdd.n2556 vdd.n721 185
R565 vdd.n721 vdd.n718 185
R566 vdd.n2555 vdd.n2554 185
R567 vdd.n723 vdd.n722 185
R568 vdd.n2322 vdd.n2321 185
R569 vdd.n2324 vdd.n2323 185
R570 vdd.n2326 vdd.n2325 185
R571 vdd.n2328 vdd.n2327 185
R572 vdd.n2330 vdd.n2329 185
R573 vdd.n2332 vdd.n2331 185
R574 vdd.n2334 vdd.n2333 185
R575 vdd.n2336 vdd.n2335 185
R576 vdd.n2338 vdd.n2337 185
R577 vdd.n2340 vdd.n2339 185
R578 vdd.n2342 vdd.n2341 185
R579 vdd.n2344 vdd.n2343 185
R580 vdd.n2346 vdd.n2345 185
R581 vdd.n2348 vdd.n2347 185
R582 vdd.n2350 vdd.n2349 185
R583 vdd.n2352 vdd.n2351 185
R584 vdd.n2354 vdd.n2353 185
R585 vdd.n2356 vdd.n2355 185
R586 vdd.n2358 vdd.n2357 185
R587 vdd.n2360 vdd.n2359 185
R588 vdd.n2362 vdd.n2361 185
R589 vdd.n2364 vdd.n2363 185
R590 vdd.n2366 vdd.n2365 185
R591 vdd.n2368 vdd.n2367 185
R592 vdd.n2370 vdd.n2369 185
R593 vdd.n2372 vdd.n2371 185
R594 vdd.n2374 vdd.n2373 185
R595 vdd.n2376 vdd.n2375 185
R596 vdd.n2378 vdd.n2377 185
R597 vdd.n2380 vdd.n2379 185
R598 vdd.n2382 vdd.n2381 185
R599 vdd.n2384 vdd.n2383 185
R600 vdd.n2385 vdd.n2312 185
R601 vdd.n2552 vdd.n2312 185
R602 vdd.n2768 vdd.n2767 185
R603 vdd.n2769 vdd.n588 185
R604 vdd.n2771 vdd.n2770 185
R605 vdd.n2773 vdd.n586 185
R606 vdd.n2775 vdd.n2774 185
R607 vdd.n2776 vdd.n585 185
R608 vdd.n2778 vdd.n2777 185
R609 vdd.n2780 vdd.n583 185
R610 vdd.n2782 vdd.n2781 185
R611 vdd.n2783 vdd.n582 185
R612 vdd.n2785 vdd.n2784 185
R613 vdd.n2787 vdd.n580 185
R614 vdd.n2789 vdd.n2788 185
R615 vdd.n2790 vdd.n579 185
R616 vdd.n2792 vdd.n2791 185
R617 vdd.n2794 vdd.n578 185
R618 vdd.n2795 vdd.n576 185
R619 vdd.n2798 vdd.n2797 185
R620 vdd.n577 vdd.n575 185
R621 vdd.n2654 vdd.n2653 185
R622 vdd.n2656 vdd.n2655 185
R623 vdd.n2658 vdd.n2650 185
R624 vdd.n2660 vdd.n2659 185
R625 vdd.n2661 vdd.n2649 185
R626 vdd.n2663 vdd.n2662 185
R627 vdd.n2665 vdd.n2647 185
R628 vdd.n2667 vdd.n2666 185
R629 vdd.n2668 vdd.n2646 185
R630 vdd.n2670 vdd.n2669 185
R631 vdd.n2672 vdd.n2644 185
R632 vdd.n2674 vdd.n2673 185
R633 vdd.n2675 vdd.n2643 185
R634 vdd.n2677 vdd.n2676 185
R635 vdd.n2679 vdd.n2642 185
R636 vdd.n2681 vdd.n2680 185
R637 vdd.n2680 vdd.n484 185
R638 vdd.n2766 vdd.n592 185
R639 vdd.n2766 vdd.n2765 185
R640 vdd.n2389 vdd.n594 185
R641 vdd.n595 vdd.n594 185
R642 vdd.n2390 vdd.n628 185
R643 vdd.n2695 vdd.n628 185
R644 vdd.n2392 vdd.n2391 185
R645 vdd.n2391 vdd.n636 185
R646 vdd.n2393 vdd.n635 185
R647 vdd.n2689 vdd.n635 185
R648 vdd.n2395 vdd.n2394 185
R649 vdd.n2394 vdd.n633 185
R650 vdd.n2396 vdd.n643 185
R651 vdd.n2638 vdd.n643 185
R652 vdd.n2398 vdd.n2397 185
R653 vdd.n2397 vdd.n641 185
R654 vdd.n2399 vdd.n649 185
R655 vdd.n2632 vdd.n649 185
R656 vdd.n2401 vdd.n2400 185
R657 vdd.n2400 vdd.n647 185
R658 vdd.n2402 vdd.n654 185
R659 vdd.n2626 vdd.n654 185
R660 vdd.n2404 vdd.n2403 185
R661 vdd.n2403 vdd.n660 185
R662 vdd.n2405 vdd.n659 185
R663 vdd.n2620 vdd.n659 185
R664 vdd.n2407 vdd.n2406 185
R665 vdd.n2406 vdd.n668 185
R666 vdd.n2408 vdd.n667 185
R667 vdd.n2613 vdd.n667 185
R668 vdd.n2410 vdd.n2409 185
R669 vdd.n2409 vdd.n665 185
R670 vdd.n2411 vdd.n674 185
R671 vdd.n2607 vdd.n674 185
R672 vdd.n2413 vdd.n2412 185
R673 vdd.n2412 vdd.n672 185
R674 vdd.n2414 vdd.n679 185
R675 vdd.n2601 vdd.n679 185
R676 vdd.n2416 vdd.n2415 185
R677 vdd.n2415 vdd.n685 185
R678 vdd.n2417 vdd.n684 185
R679 vdd.n2595 vdd.n684 185
R680 vdd.n2419 vdd.n2418 185
R681 vdd.n2418 vdd.n691 185
R682 vdd.n2420 vdd.n690 185
R683 vdd.n2589 vdd.n690 185
R684 vdd.n2463 vdd.n2462 185
R685 vdd.n2462 vdd.n2461 185
R686 vdd.n2464 vdd.n697 185
R687 vdd.n2583 vdd.n697 185
R688 vdd.n2466 vdd.n2465 185
R689 vdd.n2465 vdd.n695 185
R690 vdd.n2467 vdd.n703 185
R691 vdd.n2577 vdd.n703 185
R692 vdd.n2469 vdd.n2468 185
R693 vdd.n2468 vdd.n701 185
R694 vdd.n2470 vdd.n709 185
R695 vdd.n2571 vdd.n709 185
R696 vdd.n2472 vdd.n2471 185
R697 vdd.n2471 vdd.n707 185
R698 vdd.n2473 vdd.n714 185
R699 vdd.n2565 vdd.n714 185
R700 vdd.n2475 vdd.n2474 185
R701 vdd.n2476 vdd.n2475 185
R702 vdd.n2388 vdd.n720 185
R703 vdd.n2559 vdd.n720 185
R704 vdd.n2387 vdd.n2386 185
R705 vdd.n2386 vdd.n718 185
R706 vdd.n1878 vdd.n1877 185
R707 vdd.n1879 vdd.n1878 185
R708 vdd.n1228 vdd.n1226 185
R709 vdd.n1870 vdd.n1226 185
R710 vdd.n1873 vdd.n1872 185
R711 vdd.n1872 vdd.n1871 185
R712 vdd.n1231 vdd.n1230 185
R713 vdd.n1232 vdd.n1231 185
R714 vdd.n1859 vdd.n1858 185
R715 vdd.n1860 vdd.n1859 185
R716 vdd.n1240 vdd.n1239 185
R717 vdd.n1851 vdd.n1239 185
R718 vdd.n1854 vdd.n1853 185
R719 vdd.n1853 vdd.n1852 185
R720 vdd.n1243 vdd.n1242 185
R721 vdd.n1250 vdd.n1243 185
R722 vdd.n1842 vdd.n1841 185
R723 vdd.n1843 vdd.n1842 185
R724 vdd.n1252 vdd.n1251 185
R725 vdd.n1251 vdd.n1249 185
R726 vdd.n1837 vdd.n1836 185
R727 vdd.n1836 vdd.n1835 185
R728 vdd.n1525 vdd.n1524 185
R729 vdd.n1526 vdd.n1525 185
R730 vdd.n1826 vdd.n1825 185
R731 vdd.n1827 vdd.n1826 185
R732 vdd.n1533 vdd.n1532 185
R733 vdd.n1817 vdd.n1532 185
R734 vdd.n1820 vdd.n1819 185
R735 vdd.n1819 vdd.n1818 185
R736 vdd.n1536 vdd.n1535 185
R737 vdd.n1542 vdd.n1536 185
R738 vdd.n1808 vdd.n1807 185
R739 vdd.n1809 vdd.n1808 185
R740 vdd.n1544 vdd.n1543 185
R741 vdd.n1800 vdd.n1543 185
R742 vdd.n1803 vdd.n1802 185
R743 vdd.n1802 vdd.n1801 185
R744 vdd.n1547 vdd.n1546 185
R745 vdd.n1548 vdd.n1547 185
R746 vdd.n1791 vdd.n1790 185
R747 vdd.n1792 vdd.n1791 185
R748 vdd.n1555 vdd.n1554 185
R749 vdd.n1590 vdd.n1554 185
R750 vdd.n1786 vdd.n1785 185
R751 vdd.n1558 vdd.n1557 185
R752 vdd.n1782 vdd.n1781 185
R753 vdd.n1783 vdd.n1782 185
R754 vdd.n1592 vdd.n1591 185
R755 vdd.n1777 vdd.n1594 185
R756 vdd.n1776 vdd.n1595 185
R757 vdd.n1775 vdd.n1596 185
R758 vdd.n1598 vdd.n1597 185
R759 vdd.n1771 vdd.n1600 185
R760 vdd.n1770 vdd.n1601 185
R761 vdd.n1769 vdd.n1602 185
R762 vdd.n1604 vdd.n1603 185
R763 vdd.n1765 vdd.n1606 185
R764 vdd.n1764 vdd.n1607 185
R765 vdd.n1763 vdd.n1608 185
R766 vdd.n1610 vdd.n1609 185
R767 vdd.n1759 vdd.n1612 185
R768 vdd.n1758 vdd.n1613 185
R769 vdd.n1757 vdd.n1614 185
R770 vdd.n1618 vdd.n1615 185
R771 vdd.n1753 vdd.n1620 185
R772 vdd.n1752 vdd.n1621 185
R773 vdd.n1751 vdd.n1622 185
R774 vdd.n1624 vdd.n1623 185
R775 vdd.n1747 vdd.n1626 185
R776 vdd.n1746 vdd.n1627 185
R777 vdd.n1745 vdd.n1628 185
R778 vdd.n1630 vdd.n1629 185
R779 vdd.n1741 vdd.n1632 185
R780 vdd.n1740 vdd.n1633 185
R781 vdd.n1739 vdd.n1634 185
R782 vdd.n1636 vdd.n1635 185
R783 vdd.n1735 vdd.n1638 185
R784 vdd.n1734 vdd.n1639 185
R785 vdd.n1733 vdd.n1640 185
R786 vdd.n1642 vdd.n1641 185
R787 vdd.n1729 vdd.n1644 185
R788 vdd.n1728 vdd.n1645 185
R789 vdd.n1727 vdd.n1646 185
R790 vdd.n1648 vdd.n1647 185
R791 vdd.n1723 vdd.n1650 185
R792 vdd.n1722 vdd.n1719 185
R793 vdd.n1718 vdd.n1651 185
R794 vdd.n1653 vdd.n1652 185
R795 vdd.n1714 vdd.n1655 185
R796 vdd.n1713 vdd.n1656 185
R797 vdd.n1712 vdd.n1657 185
R798 vdd.n1659 vdd.n1658 185
R799 vdd.n1708 vdd.n1661 185
R800 vdd.n1707 vdd.n1662 185
R801 vdd.n1706 vdd.n1663 185
R802 vdd.n1665 vdd.n1664 185
R803 vdd.n1702 vdd.n1667 185
R804 vdd.n1701 vdd.n1668 185
R805 vdd.n1700 vdd.n1669 185
R806 vdd.n1671 vdd.n1670 185
R807 vdd.n1696 vdd.n1673 185
R808 vdd.n1695 vdd.n1674 185
R809 vdd.n1694 vdd.n1675 185
R810 vdd.n1677 vdd.n1676 185
R811 vdd.n1690 vdd.n1679 185
R812 vdd.n1689 vdd.n1680 185
R813 vdd.n1688 vdd.n1681 185
R814 vdd.n1685 vdd.n1589 185
R815 vdd.n1783 vdd.n1589 185
R816 vdd.n1882 vdd.n1881 185
R817 vdd.n1886 vdd.n1222 185
R818 vdd.n1221 vdd.n1215 185
R819 vdd.n1219 vdd.n1218 185
R820 vdd.n1217 vdd.n1011 185
R821 vdd.n1890 vdd.n1008 185
R822 vdd.n1892 vdd.n1891 185
R823 vdd.n1894 vdd.n1006 185
R824 vdd.n1896 vdd.n1895 185
R825 vdd.n1897 vdd.n1001 185
R826 vdd.n1899 vdd.n1898 185
R827 vdd.n1901 vdd.n999 185
R828 vdd.n1903 vdd.n1902 185
R829 vdd.n1904 vdd.n994 185
R830 vdd.n1906 vdd.n1905 185
R831 vdd.n1908 vdd.n992 185
R832 vdd.n1910 vdd.n1909 185
R833 vdd.n1911 vdd.n988 185
R834 vdd.n1913 vdd.n1912 185
R835 vdd.n1915 vdd.n985 185
R836 vdd.n1917 vdd.n1916 185
R837 vdd.n986 vdd.n979 185
R838 vdd.n1921 vdd.n983 185
R839 vdd.n1922 vdd.n975 185
R840 vdd.n1924 vdd.n1923 185
R841 vdd.n1926 vdd.n973 185
R842 vdd.n1928 vdd.n1927 185
R843 vdd.n1929 vdd.n968 185
R844 vdd.n1931 vdd.n1930 185
R845 vdd.n1933 vdd.n966 185
R846 vdd.n1935 vdd.n1934 185
R847 vdd.n1936 vdd.n961 185
R848 vdd.n1938 vdd.n1937 185
R849 vdd.n1940 vdd.n959 185
R850 vdd.n1942 vdd.n1941 185
R851 vdd.n1943 vdd.n954 185
R852 vdd.n1945 vdd.n1944 185
R853 vdd.n1947 vdd.n952 185
R854 vdd.n1949 vdd.n1948 185
R855 vdd.n1950 vdd.n948 185
R856 vdd.n1952 vdd.n1951 185
R857 vdd.n1954 vdd.n945 185
R858 vdd.n1956 vdd.n1955 185
R859 vdd.n946 vdd.n939 185
R860 vdd.n1960 vdd.n943 185
R861 vdd.n1961 vdd.n935 185
R862 vdd.n1963 vdd.n1962 185
R863 vdd.n1965 vdd.n933 185
R864 vdd.n1967 vdd.n1966 185
R865 vdd.n1968 vdd.n928 185
R866 vdd.n1970 vdd.n1969 185
R867 vdd.n1972 vdd.n926 185
R868 vdd.n1974 vdd.n1973 185
R869 vdd.n1975 vdd.n921 185
R870 vdd.n1977 vdd.n1976 185
R871 vdd.n1979 vdd.n919 185
R872 vdd.n1981 vdd.n1980 185
R873 vdd.n1982 vdd.n917 185
R874 vdd.n1984 vdd.n1983 185
R875 vdd.n1987 vdd.n1986 185
R876 vdd.n1989 vdd.n1988 185
R877 vdd.n1991 vdd.n915 185
R878 vdd.n1993 vdd.n1992 185
R879 vdd.n1227 vdd.n914 185
R880 vdd.n1880 vdd.n1225 185
R881 vdd.n1880 vdd.n1879 185
R882 vdd.n1235 vdd.n1224 185
R883 vdd.n1870 vdd.n1224 185
R884 vdd.n1869 vdd.n1868 185
R885 vdd.n1871 vdd.n1869 185
R886 vdd.n1234 vdd.n1233 185
R887 vdd.n1233 vdd.n1232 185
R888 vdd.n1862 vdd.n1861 185
R889 vdd.n1861 vdd.n1860 185
R890 vdd.n1238 vdd.n1237 185
R891 vdd.n1851 vdd.n1238 185
R892 vdd.n1850 vdd.n1849 185
R893 vdd.n1852 vdd.n1850 185
R894 vdd.n1245 vdd.n1244 185
R895 vdd.n1250 vdd.n1244 185
R896 vdd.n1845 vdd.n1844 185
R897 vdd.n1844 vdd.n1843 185
R898 vdd.n1248 vdd.n1247 185
R899 vdd.n1249 vdd.n1248 185
R900 vdd.n1834 vdd.n1833 185
R901 vdd.n1835 vdd.n1834 185
R902 vdd.n1528 vdd.n1527 185
R903 vdd.n1527 vdd.n1526 185
R904 vdd.n1829 vdd.n1828 185
R905 vdd.n1828 vdd.n1827 185
R906 vdd.n1531 vdd.n1530 185
R907 vdd.n1817 vdd.n1531 185
R908 vdd.n1816 vdd.n1815 185
R909 vdd.n1818 vdd.n1816 185
R910 vdd.n1538 vdd.n1537 185
R911 vdd.n1542 vdd.n1537 185
R912 vdd.n1811 vdd.n1810 185
R913 vdd.n1810 vdd.n1809 185
R914 vdd.n1541 vdd.n1540 185
R915 vdd.n1800 vdd.n1541 185
R916 vdd.n1799 vdd.n1798 185
R917 vdd.n1801 vdd.n1799 185
R918 vdd.n1550 vdd.n1549 185
R919 vdd.n1549 vdd.n1548 185
R920 vdd.n1794 vdd.n1793 185
R921 vdd.n1793 vdd.n1792 185
R922 vdd.n1553 vdd.n1552 185
R923 vdd.n1590 vdd.n1553 185
R924 vdd.n761 vdd.n759 185
R925 vdd.n2207 vdd.n759 185
R926 vdd.n2129 vdd.n779 185
R927 vdd.n779 vdd.n766 185
R928 vdd.n2131 vdd.n2130 185
R929 vdd.n2132 vdd.n2131 185
R930 vdd.n2128 vdd.n778 185
R931 vdd.n1128 vdd.n778 185
R932 vdd.n2127 vdd.n2126 185
R933 vdd.n2126 vdd.n2125 185
R934 vdd.n781 vdd.n780 185
R935 vdd.n782 vdd.n781 185
R936 vdd.n2116 vdd.n2115 185
R937 vdd.n2117 vdd.n2116 185
R938 vdd.n2114 vdd.n792 185
R939 vdd.n792 vdd.n789 185
R940 vdd.n2113 vdd.n2112 185
R941 vdd.n2112 vdd.n2111 185
R942 vdd.n794 vdd.n793 185
R943 vdd.n795 vdd.n794 185
R944 vdd.n2104 vdd.n2103 185
R945 vdd.n2105 vdd.n2104 185
R946 vdd.n2102 vdd.n803 185
R947 vdd.n808 vdd.n803 185
R948 vdd.n2101 vdd.n2100 185
R949 vdd.n2100 vdd.n2099 185
R950 vdd.n805 vdd.n804 185
R951 vdd.n814 vdd.n805 185
R952 vdd.n2092 vdd.n2091 185
R953 vdd.n2093 vdd.n2092 185
R954 vdd.n2090 vdd.n815 185
R955 vdd.n1149 vdd.n815 185
R956 vdd.n2089 vdd.n2088 185
R957 vdd.n2088 vdd.n2087 185
R958 vdd.n817 vdd.n816 185
R959 vdd.n818 vdd.n817 185
R960 vdd.n2080 vdd.n2079 185
R961 vdd.n2081 vdd.n2080 185
R962 vdd.n2078 vdd.n827 185
R963 vdd.n827 vdd.n824 185
R964 vdd.n2077 vdd.n2076 185
R965 vdd.n2076 vdd.n2075 185
R966 vdd.n829 vdd.n828 185
R967 vdd.n838 vdd.n829 185
R968 vdd.n2067 vdd.n2066 185
R969 vdd.n2068 vdd.n2067 185
R970 vdd.n2065 vdd.n839 185
R971 vdd.n845 vdd.n839 185
R972 vdd.n2064 vdd.n2063 185
R973 vdd.n2063 vdd.n2062 185
R974 vdd.n841 vdd.n840 185
R975 vdd.n842 vdd.n841 185
R976 vdd.n2055 vdd.n2054 185
R977 vdd.n2056 vdd.n2055 185
R978 vdd.n2053 vdd.n852 185
R979 vdd.n852 vdd.n849 185
R980 vdd.n2052 vdd.n2051 185
R981 vdd.n2051 vdd.n2050 185
R982 vdd.n854 vdd.n853 185
R983 vdd.n855 vdd.n854 185
R984 vdd.n2043 vdd.n2042 185
R985 vdd.n2044 vdd.n2043 185
R986 vdd.n2041 vdd.n863 185
R987 vdd.n869 vdd.n863 185
R988 vdd.n2040 vdd.n2039 185
R989 vdd.n2039 vdd.n2038 185
R990 vdd.n865 vdd.n864 185
R991 vdd.n866 vdd.n865 185
R992 vdd.n2029 vdd.n2028 185
R993 vdd.n2027 vdd.n908 185
R994 vdd.n2026 vdd.n907 185
R995 vdd.n2031 vdd.n907 185
R996 vdd.n2025 vdd.n2024 185
R997 vdd.n2023 vdd.n2022 185
R998 vdd.n2021 vdd.n2020 185
R999 vdd.n2019 vdd.n2018 185
R1000 vdd.n2017 vdd.n2016 185
R1001 vdd.n2015 vdd.n2014 185
R1002 vdd.n2013 vdd.n2012 185
R1003 vdd.n2011 vdd.n2010 185
R1004 vdd.n2009 vdd.n2008 185
R1005 vdd.n2007 vdd.n2006 185
R1006 vdd.n2005 vdd.n2004 185
R1007 vdd.n2003 vdd.n2002 185
R1008 vdd.n2001 vdd.n2000 185
R1009 vdd.n1999 vdd.n1998 185
R1010 vdd.n1997 vdd.n1996 185
R1011 vdd.n1065 vdd.n909 185
R1012 vdd.n1067 vdd.n1066 185
R1013 vdd.n1069 vdd.n1068 185
R1014 vdd.n1071 vdd.n1070 185
R1015 vdd.n1073 vdd.n1072 185
R1016 vdd.n1075 vdd.n1074 185
R1017 vdd.n1077 vdd.n1076 185
R1018 vdd.n1079 vdd.n1078 185
R1019 vdd.n1081 vdd.n1080 185
R1020 vdd.n1083 vdd.n1082 185
R1021 vdd.n1085 vdd.n1084 185
R1022 vdd.n1087 vdd.n1086 185
R1023 vdd.n1089 vdd.n1088 185
R1024 vdd.n1091 vdd.n1090 185
R1025 vdd.n1094 vdd.n1093 185
R1026 vdd.n1096 vdd.n1095 185
R1027 vdd.n1098 vdd.n1097 185
R1028 vdd.n2210 vdd.n2209 185
R1029 vdd.n2212 vdd.n2211 185
R1030 vdd.n2214 vdd.n2213 185
R1031 vdd.n2217 vdd.n2216 185
R1032 vdd.n2219 vdd.n2218 185
R1033 vdd.n2221 vdd.n2220 185
R1034 vdd.n2223 vdd.n2222 185
R1035 vdd.n2225 vdd.n2224 185
R1036 vdd.n2227 vdd.n2226 185
R1037 vdd.n2229 vdd.n2228 185
R1038 vdd.n2231 vdd.n2230 185
R1039 vdd.n2233 vdd.n2232 185
R1040 vdd.n2235 vdd.n2234 185
R1041 vdd.n2237 vdd.n2236 185
R1042 vdd.n2239 vdd.n2238 185
R1043 vdd.n2241 vdd.n2240 185
R1044 vdd.n2243 vdd.n2242 185
R1045 vdd.n2245 vdd.n2244 185
R1046 vdd.n2247 vdd.n2246 185
R1047 vdd.n2249 vdd.n2248 185
R1048 vdd.n2251 vdd.n2250 185
R1049 vdd.n2253 vdd.n2252 185
R1050 vdd.n2255 vdd.n2254 185
R1051 vdd.n2257 vdd.n2256 185
R1052 vdd.n2259 vdd.n2258 185
R1053 vdd.n2261 vdd.n2260 185
R1054 vdd.n2263 vdd.n2262 185
R1055 vdd.n2265 vdd.n2264 185
R1056 vdd.n2267 vdd.n2266 185
R1057 vdd.n2269 vdd.n2268 185
R1058 vdd.n2271 vdd.n2270 185
R1059 vdd.n2273 vdd.n2272 185
R1060 vdd.n2275 vdd.n2274 185
R1061 vdd.n2276 vdd.n760 185
R1062 vdd.n2278 vdd.n2277 185
R1063 vdd.n2279 vdd.n2278 185
R1064 vdd.n2208 vdd.n764 185
R1065 vdd.n2208 vdd.n2207 185
R1066 vdd.n1126 vdd.n765 185
R1067 vdd.n766 vdd.n765 185
R1068 vdd.n1127 vdd.n776 185
R1069 vdd.n2132 vdd.n776 185
R1070 vdd.n1130 vdd.n1129 185
R1071 vdd.n1129 vdd.n1128 185
R1072 vdd.n1131 vdd.n783 185
R1073 vdd.n2125 vdd.n783 185
R1074 vdd.n1133 vdd.n1132 185
R1075 vdd.n1132 vdd.n782 185
R1076 vdd.n1134 vdd.n790 185
R1077 vdd.n2117 vdd.n790 185
R1078 vdd.n1136 vdd.n1135 185
R1079 vdd.n1135 vdd.n789 185
R1080 vdd.n1137 vdd.n796 185
R1081 vdd.n2111 vdd.n796 185
R1082 vdd.n1139 vdd.n1138 185
R1083 vdd.n1138 vdd.n795 185
R1084 vdd.n1140 vdd.n801 185
R1085 vdd.n2105 vdd.n801 185
R1086 vdd.n1142 vdd.n1141 185
R1087 vdd.n1141 vdd.n808 185
R1088 vdd.n1143 vdd.n806 185
R1089 vdd.n2099 vdd.n806 185
R1090 vdd.n1145 vdd.n1144 185
R1091 vdd.n1144 vdd.n814 185
R1092 vdd.n1146 vdd.n812 185
R1093 vdd.n2093 vdd.n812 185
R1094 vdd.n1148 vdd.n1147 185
R1095 vdd.n1149 vdd.n1148 185
R1096 vdd.n1125 vdd.n819 185
R1097 vdd.n2087 vdd.n819 185
R1098 vdd.n1124 vdd.n1123 185
R1099 vdd.n1123 vdd.n818 185
R1100 vdd.n1122 vdd.n825 185
R1101 vdd.n2081 vdd.n825 185
R1102 vdd.n1121 vdd.n1120 185
R1103 vdd.n1120 vdd.n824 185
R1104 vdd.n1119 vdd.n830 185
R1105 vdd.n2075 vdd.n830 185
R1106 vdd.n1118 vdd.n1117 185
R1107 vdd.n1117 vdd.n838 185
R1108 vdd.n1116 vdd.n836 185
R1109 vdd.n2068 vdd.n836 185
R1110 vdd.n1115 vdd.n1114 185
R1111 vdd.n1114 vdd.n845 185
R1112 vdd.n1113 vdd.n843 185
R1113 vdd.n2062 vdd.n843 185
R1114 vdd.n1112 vdd.n1111 185
R1115 vdd.n1111 vdd.n842 185
R1116 vdd.n1110 vdd.n850 185
R1117 vdd.n2056 vdd.n850 185
R1118 vdd.n1109 vdd.n1108 185
R1119 vdd.n1108 vdd.n849 185
R1120 vdd.n1107 vdd.n856 185
R1121 vdd.n2050 vdd.n856 185
R1122 vdd.n1106 vdd.n1105 185
R1123 vdd.n1105 vdd.n855 185
R1124 vdd.n1104 vdd.n861 185
R1125 vdd.n2044 vdd.n861 185
R1126 vdd.n1103 vdd.n1102 185
R1127 vdd.n1102 vdd.n869 185
R1128 vdd.n1101 vdd.n867 185
R1129 vdd.n2038 vdd.n867 185
R1130 vdd.n1100 vdd.n1099 185
R1131 vdd.n1099 vdd.n866 185
R1132 vdd.n3116 vdd.n3115 185
R1133 vdd.n3117 vdd.n3116 185
R1134 vdd.n325 vdd.n324 185
R1135 vdd.n3118 vdd.n325 185
R1136 vdd.n3121 vdd.n3120 185
R1137 vdd.n3120 vdd.n3119 185
R1138 vdd.n3122 vdd.n319 185
R1139 vdd.n319 vdd.n318 185
R1140 vdd.n3124 vdd.n3123 185
R1141 vdd.n3125 vdd.n3124 185
R1142 vdd.n314 vdd.n313 185
R1143 vdd.n3126 vdd.n314 185
R1144 vdd.n3129 vdd.n3128 185
R1145 vdd.n3128 vdd.n3127 185
R1146 vdd.n3130 vdd.n309 185
R1147 vdd.n309 vdd.n308 185
R1148 vdd.n3132 vdd.n3131 185
R1149 vdd.n3133 vdd.n3132 185
R1150 vdd.n303 vdd.n301 185
R1151 vdd.n3134 vdd.n303 185
R1152 vdd.n3137 vdd.n3136 185
R1153 vdd.n3136 vdd.n3135 185
R1154 vdd.n302 vdd.n300 185
R1155 vdd.n304 vdd.n302 185
R1156 vdd.n2973 vdd.n2972 185
R1157 vdd.n2974 vdd.n2973 185
R1158 vdd.n458 vdd.n457 185
R1159 vdd.n457 vdd.n456 185
R1160 vdd.n2968 vdd.n2967 185
R1161 vdd.n2967 vdd.n2966 185
R1162 vdd.n461 vdd.n460 185
R1163 vdd.n467 vdd.n461 185
R1164 vdd.n2957 vdd.n2956 185
R1165 vdd.n2958 vdd.n2957 185
R1166 vdd.n469 vdd.n468 185
R1167 vdd.n2949 vdd.n468 185
R1168 vdd.n2952 vdd.n2951 185
R1169 vdd.n2951 vdd.n2950 185
R1170 vdd.n472 vdd.n471 185
R1171 vdd.n473 vdd.n472 185
R1172 vdd.n2940 vdd.n2939 185
R1173 vdd.n2941 vdd.n2940 185
R1174 vdd.n480 vdd.n479 185
R1175 vdd.n516 vdd.n479 185
R1176 vdd.n2935 vdd.n2934 185
R1177 vdd.n483 vdd.n482 185
R1178 vdd.n2931 vdd.n2930 185
R1179 vdd.n2932 vdd.n2931 185
R1180 vdd.n518 vdd.n517 185
R1181 vdd.n522 vdd.n521 185
R1182 vdd.n2926 vdd.n523 185
R1183 vdd.n2925 vdd.n2924 185
R1184 vdd.n2923 vdd.n2922 185
R1185 vdd.n2921 vdd.n2920 185
R1186 vdd.n2919 vdd.n2918 185
R1187 vdd.n2917 vdd.n2916 185
R1188 vdd.n2915 vdd.n2914 185
R1189 vdd.n2913 vdd.n2912 185
R1190 vdd.n2911 vdd.n2910 185
R1191 vdd.n2909 vdd.n2908 185
R1192 vdd.n2907 vdd.n2906 185
R1193 vdd.n2905 vdd.n2904 185
R1194 vdd.n2903 vdd.n2902 185
R1195 vdd.n2901 vdd.n2900 185
R1196 vdd.n2899 vdd.n2898 185
R1197 vdd.n2890 vdd.n536 185
R1198 vdd.n2892 vdd.n2891 185
R1199 vdd.n2889 vdd.n2888 185
R1200 vdd.n2887 vdd.n2886 185
R1201 vdd.n2885 vdd.n2884 185
R1202 vdd.n2883 vdd.n2882 185
R1203 vdd.n2881 vdd.n2880 185
R1204 vdd.n2879 vdd.n2878 185
R1205 vdd.n2877 vdd.n2876 185
R1206 vdd.n2875 vdd.n2874 185
R1207 vdd.n2873 vdd.n2872 185
R1208 vdd.n2871 vdd.n2870 185
R1209 vdd.n2869 vdd.n2868 185
R1210 vdd.n2867 vdd.n2866 185
R1211 vdd.n2865 vdd.n2864 185
R1212 vdd.n2863 vdd.n2862 185
R1213 vdd.n2861 vdd.n2860 185
R1214 vdd.n2859 vdd.n2858 185
R1215 vdd.n2857 vdd.n2856 185
R1216 vdd.n2855 vdd.n2854 185
R1217 vdd.n2853 vdd.n2852 185
R1218 vdd.n2851 vdd.n2850 185
R1219 vdd.n2844 vdd.n556 185
R1220 vdd.n2846 vdd.n2845 185
R1221 vdd.n2843 vdd.n2842 185
R1222 vdd.n2841 vdd.n2840 185
R1223 vdd.n2839 vdd.n2838 185
R1224 vdd.n2837 vdd.n2836 185
R1225 vdd.n2835 vdd.n2834 185
R1226 vdd.n2833 vdd.n2832 185
R1227 vdd.n2831 vdd.n2830 185
R1228 vdd.n2829 vdd.n2828 185
R1229 vdd.n2827 vdd.n2826 185
R1230 vdd.n2825 vdd.n2824 185
R1231 vdd.n2823 vdd.n2822 185
R1232 vdd.n2821 vdd.n2820 185
R1233 vdd.n2819 vdd.n2818 185
R1234 vdd.n2817 vdd.n2816 185
R1235 vdd.n2815 vdd.n2814 185
R1236 vdd.n2813 vdd.n2812 185
R1237 vdd.n2811 vdd.n2810 185
R1238 vdd.n2809 vdd.n2808 185
R1239 vdd.n2807 vdd.n2806 185
R1240 vdd.n2802 vdd.n515 185
R1241 vdd.n2932 vdd.n515 185
R1242 vdd.n2999 vdd.n2998 185
R1243 vdd.n3003 vdd.n440 185
R1244 vdd.n3005 vdd.n3004 185
R1245 vdd.n3007 vdd.n438 185
R1246 vdd.n3009 vdd.n3008 185
R1247 vdd.n3010 vdd.n433 185
R1248 vdd.n3012 vdd.n3011 185
R1249 vdd.n3014 vdd.n431 185
R1250 vdd.n3016 vdd.n3015 185
R1251 vdd.n3017 vdd.n426 185
R1252 vdd.n3019 vdd.n3018 185
R1253 vdd.n3021 vdd.n424 185
R1254 vdd.n3023 vdd.n3022 185
R1255 vdd.n3024 vdd.n419 185
R1256 vdd.n3026 vdd.n3025 185
R1257 vdd.n3028 vdd.n417 185
R1258 vdd.n3030 vdd.n3029 185
R1259 vdd.n3031 vdd.n413 185
R1260 vdd.n3033 vdd.n3032 185
R1261 vdd.n3035 vdd.n410 185
R1262 vdd.n3037 vdd.n3036 185
R1263 vdd.n411 vdd.n404 185
R1264 vdd.n3041 vdd.n408 185
R1265 vdd.n3042 vdd.n400 185
R1266 vdd.n3044 vdd.n3043 185
R1267 vdd.n3046 vdd.n398 185
R1268 vdd.n3048 vdd.n3047 185
R1269 vdd.n3049 vdd.n393 185
R1270 vdd.n3051 vdd.n3050 185
R1271 vdd.n3053 vdd.n391 185
R1272 vdd.n3055 vdd.n3054 185
R1273 vdd.n3056 vdd.n386 185
R1274 vdd.n3058 vdd.n3057 185
R1275 vdd.n3060 vdd.n384 185
R1276 vdd.n3062 vdd.n3061 185
R1277 vdd.n3063 vdd.n379 185
R1278 vdd.n3065 vdd.n3064 185
R1279 vdd.n3067 vdd.n377 185
R1280 vdd.n3069 vdd.n3068 185
R1281 vdd.n3070 vdd.n373 185
R1282 vdd.n3072 vdd.n3071 185
R1283 vdd.n3074 vdd.n370 185
R1284 vdd.n3076 vdd.n3075 185
R1285 vdd.n371 vdd.n364 185
R1286 vdd.n3080 vdd.n368 185
R1287 vdd.n3081 vdd.n360 185
R1288 vdd.n3083 vdd.n3082 185
R1289 vdd.n3085 vdd.n358 185
R1290 vdd.n3087 vdd.n3086 185
R1291 vdd.n3088 vdd.n353 185
R1292 vdd.n3090 vdd.n3089 185
R1293 vdd.n3092 vdd.n351 185
R1294 vdd.n3094 vdd.n3093 185
R1295 vdd.n3095 vdd.n346 185
R1296 vdd.n3097 vdd.n3096 185
R1297 vdd.n3099 vdd.n344 185
R1298 vdd.n3101 vdd.n3100 185
R1299 vdd.n3102 vdd.n338 185
R1300 vdd.n3104 vdd.n3103 185
R1301 vdd.n3106 vdd.n337 185
R1302 vdd.n3107 vdd.n336 185
R1303 vdd.n3110 vdd.n3109 185
R1304 vdd.n3111 vdd.n334 185
R1305 vdd.n3112 vdd.n330 185
R1306 vdd.n2994 vdd.n328 185
R1307 vdd.n3117 vdd.n328 185
R1308 vdd.n2993 vdd.n327 185
R1309 vdd.n3118 vdd.n327 185
R1310 vdd.n2992 vdd.n326 185
R1311 vdd.n3119 vdd.n326 185
R1312 vdd.n446 vdd.n445 185
R1313 vdd.n445 vdd.n318 185
R1314 vdd.n2988 vdd.n317 185
R1315 vdd.n3125 vdd.n317 185
R1316 vdd.n2987 vdd.n316 185
R1317 vdd.n3126 vdd.n316 185
R1318 vdd.n2986 vdd.n315 185
R1319 vdd.n3127 vdd.n315 185
R1320 vdd.n449 vdd.n448 185
R1321 vdd.n448 vdd.n308 185
R1322 vdd.n2982 vdd.n307 185
R1323 vdd.n3133 vdd.n307 185
R1324 vdd.n2981 vdd.n306 185
R1325 vdd.n3134 vdd.n306 185
R1326 vdd.n2980 vdd.n305 185
R1327 vdd.n3135 vdd.n305 185
R1328 vdd.n455 vdd.n451 185
R1329 vdd.n455 vdd.n304 185
R1330 vdd.n2976 vdd.n2975 185
R1331 vdd.n2975 vdd.n2974 185
R1332 vdd.n454 vdd.n453 185
R1333 vdd.n456 vdd.n454 185
R1334 vdd.n2965 vdd.n2964 185
R1335 vdd.n2966 vdd.n2965 185
R1336 vdd.n463 vdd.n462 185
R1337 vdd.n467 vdd.n462 185
R1338 vdd.n2960 vdd.n2959 185
R1339 vdd.n2959 vdd.n2958 185
R1340 vdd.n466 vdd.n465 185
R1341 vdd.n2949 vdd.n466 185
R1342 vdd.n2948 vdd.n2947 185
R1343 vdd.n2950 vdd.n2948 185
R1344 vdd.n475 vdd.n474 185
R1345 vdd.n474 vdd.n473 185
R1346 vdd.n2943 vdd.n2942 185
R1347 vdd.n2942 vdd.n2941 185
R1348 vdd.n478 vdd.n477 185
R1349 vdd.n516 vdd.n478 185
R1350 vdd.n2550 vdd.n2549 185
R1351 vdd.n2548 vdd.n2314 185
R1352 vdd.n2547 vdd.n2313 185
R1353 vdd.n2552 vdd.n2313 185
R1354 vdd.n2546 vdd.n2545 185
R1355 vdd.n2544 vdd.n2543 185
R1356 vdd.n2542 vdd.n2541 185
R1357 vdd.n2540 vdd.n2539 185
R1358 vdd.n2538 vdd.n2537 185
R1359 vdd.n2536 vdd.n2535 185
R1360 vdd.n2534 vdd.n2533 185
R1361 vdd.n2532 vdd.n2531 185
R1362 vdd.n2530 vdd.n2529 185
R1363 vdd.n2528 vdd.n2527 185
R1364 vdd.n2526 vdd.n2525 185
R1365 vdd.n2524 vdd.n2523 185
R1366 vdd.n2522 vdd.n2521 185
R1367 vdd.n2520 vdd.n2519 185
R1368 vdd.n2518 vdd.n2517 185
R1369 vdd.n2516 vdd.n2515 185
R1370 vdd.n2514 vdd.n2513 185
R1371 vdd.n2512 vdd.n2511 185
R1372 vdd.n2510 vdd.n2509 185
R1373 vdd.n2508 vdd.n2507 185
R1374 vdd.n2506 vdd.n2505 185
R1375 vdd.n2504 vdd.n2503 185
R1376 vdd.n2502 vdd.n2501 185
R1377 vdd.n2500 vdd.n2499 185
R1378 vdd.n2498 vdd.n2497 185
R1379 vdd.n2496 vdd.n2495 185
R1380 vdd.n2494 vdd.n2493 185
R1381 vdd.n2492 vdd.n2491 185
R1382 vdd.n2490 vdd.n2489 185
R1383 vdd.n2487 vdd.n2486 185
R1384 vdd.n2485 vdd.n2484 185
R1385 vdd.n2483 vdd.n2482 185
R1386 vdd.n2701 vdd.n2700 185
R1387 vdd.n2703 vdd.n624 185
R1388 vdd.n2705 vdd.n2704 185
R1389 vdd.n2707 vdd.n621 185
R1390 vdd.n2709 vdd.n2708 185
R1391 vdd.n2711 vdd.n619 185
R1392 vdd.n2713 vdd.n2712 185
R1393 vdd.n2714 vdd.n618 185
R1394 vdd.n2716 vdd.n2715 185
R1395 vdd.n2718 vdd.n616 185
R1396 vdd.n2720 vdd.n2719 185
R1397 vdd.n2721 vdd.n615 185
R1398 vdd.n2723 vdd.n2722 185
R1399 vdd.n2725 vdd.n613 185
R1400 vdd.n2727 vdd.n2726 185
R1401 vdd.n2728 vdd.n612 185
R1402 vdd.n2730 vdd.n2729 185
R1403 vdd.n2732 vdd.n520 185
R1404 vdd.n2734 vdd.n2733 185
R1405 vdd.n2736 vdd.n610 185
R1406 vdd.n2738 vdd.n2737 185
R1407 vdd.n2739 vdd.n609 185
R1408 vdd.n2741 vdd.n2740 185
R1409 vdd.n2743 vdd.n607 185
R1410 vdd.n2745 vdd.n2744 185
R1411 vdd.n2746 vdd.n606 185
R1412 vdd.n2748 vdd.n2747 185
R1413 vdd.n2750 vdd.n604 185
R1414 vdd.n2752 vdd.n2751 185
R1415 vdd.n2753 vdd.n603 185
R1416 vdd.n2755 vdd.n2754 185
R1417 vdd.n2757 vdd.n602 185
R1418 vdd.n2758 vdd.n601 185
R1419 vdd.n2761 vdd.n2760 185
R1420 vdd.n2762 vdd.n599 185
R1421 vdd.n599 vdd.n484 185
R1422 vdd.n2699 vdd.n596 185
R1423 vdd.n2765 vdd.n596 185
R1424 vdd.n2698 vdd.n2697 185
R1425 vdd.n2697 vdd.n595 185
R1426 vdd.n2696 vdd.n626 185
R1427 vdd.n2696 vdd.n2695 185
R1428 vdd.n2430 vdd.n627 185
R1429 vdd.n636 vdd.n627 185
R1430 vdd.n2431 vdd.n634 185
R1431 vdd.n2689 vdd.n634 185
R1432 vdd.n2433 vdd.n2432 185
R1433 vdd.n2432 vdd.n633 185
R1434 vdd.n2434 vdd.n642 185
R1435 vdd.n2638 vdd.n642 185
R1436 vdd.n2436 vdd.n2435 185
R1437 vdd.n2435 vdd.n641 185
R1438 vdd.n2437 vdd.n648 185
R1439 vdd.n2632 vdd.n648 185
R1440 vdd.n2439 vdd.n2438 185
R1441 vdd.n2438 vdd.n647 185
R1442 vdd.n2440 vdd.n653 185
R1443 vdd.n2626 vdd.n653 185
R1444 vdd.n2442 vdd.n2441 185
R1445 vdd.n2441 vdd.n660 185
R1446 vdd.n2443 vdd.n658 185
R1447 vdd.n2620 vdd.n658 185
R1448 vdd.n2445 vdd.n2444 185
R1449 vdd.n2444 vdd.n668 185
R1450 vdd.n2446 vdd.n666 185
R1451 vdd.n2613 vdd.n666 185
R1452 vdd.n2448 vdd.n2447 185
R1453 vdd.n2447 vdd.n665 185
R1454 vdd.n2449 vdd.n673 185
R1455 vdd.n2607 vdd.n673 185
R1456 vdd.n2451 vdd.n2450 185
R1457 vdd.n2450 vdd.n672 185
R1458 vdd.n2452 vdd.n678 185
R1459 vdd.n2601 vdd.n678 185
R1460 vdd.n2454 vdd.n2453 185
R1461 vdd.n2453 vdd.n685 185
R1462 vdd.n2455 vdd.n683 185
R1463 vdd.n2595 vdd.n683 185
R1464 vdd.n2457 vdd.n2456 185
R1465 vdd.n2456 vdd.n691 185
R1466 vdd.n2458 vdd.n689 185
R1467 vdd.n2589 vdd.n689 185
R1468 vdd.n2460 vdd.n2459 185
R1469 vdd.n2461 vdd.n2460 185
R1470 vdd.n2429 vdd.n696 185
R1471 vdd.n2583 vdd.n696 185
R1472 vdd.n2428 vdd.n2427 185
R1473 vdd.n2427 vdd.n695 185
R1474 vdd.n2426 vdd.n702 185
R1475 vdd.n2577 vdd.n702 185
R1476 vdd.n2425 vdd.n2424 185
R1477 vdd.n2424 vdd.n701 185
R1478 vdd.n2423 vdd.n708 185
R1479 vdd.n2571 vdd.n708 185
R1480 vdd.n2422 vdd.n2421 185
R1481 vdd.n2421 vdd.n707 185
R1482 vdd.n2317 vdd.n713 185
R1483 vdd.n2565 vdd.n713 185
R1484 vdd.n2478 vdd.n2477 185
R1485 vdd.n2477 vdd.n2476 185
R1486 vdd.n2479 vdd.n719 185
R1487 vdd.n2559 vdd.n719 185
R1488 vdd.n2481 vdd.n2480 185
R1489 vdd.n2481 vdd.n718 185
R1490 vdd.n717 vdd.n716 185
R1491 vdd.n718 vdd.n717 185
R1492 vdd.n2561 vdd.n2560 185
R1493 vdd.n2560 vdd.n2559 185
R1494 vdd.n2562 vdd.n715 185
R1495 vdd.n2476 vdd.n715 185
R1496 vdd.n2564 vdd.n2563 185
R1497 vdd.n2565 vdd.n2564 185
R1498 vdd.n706 vdd.n705 185
R1499 vdd.n707 vdd.n706 185
R1500 vdd.n2573 vdd.n2572 185
R1501 vdd.n2572 vdd.n2571 185
R1502 vdd.n2574 vdd.n704 185
R1503 vdd.n704 vdd.n701 185
R1504 vdd.n2576 vdd.n2575 185
R1505 vdd.n2577 vdd.n2576 185
R1506 vdd.n694 vdd.n693 185
R1507 vdd.n695 vdd.n694 185
R1508 vdd.n2585 vdd.n2584 185
R1509 vdd.n2584 vdd.n2583 185
R1510 vdd.n2586 vdd.n692 185
R1511 vdd.n2461 vdd.n692 185
R1512 vdd.n2588 vdd.n2587 185
R1513 vdd.n2589 vdd.n2588 185
R1514 vdd.n682 vdd.n681 185
R1515 vdd.n691 vdd.n682 185
R1516 vdd.n2597 vdd.n2596 185
R1517 vdd.n2596 vdd.n2595 185
R1518 vdd.n2598 vdd.n680 185
R1519 vdd.n685 vdd.n680 185
R1520 vdd.n2600 vdd.n2599 185
R1521 vdd.n2601 vdd.n2600 185
R1522 vdd.n671 vdd.n670 185
R1523 vdd.n672 vdd.n671 185
R1524 vdd.n2609 vdd.n2608 185
R1525 vdd.n2608 vdd.n2607 185
R1526 vdd.n2610 vdd.n669 185
R1527 vdd.n669 vdd.n665 185
R1528 vdd.n2612 vdd.n2611 185
R1529 vdd.n2613 vdd.n2612 185
R1530 vdd.n657 vdd.n656 185
R1531 vdd.n668 vdd.n657 185
R1532 vdd.n2622 vdd.n2621 185
R1533 vdd.n2621 vdd.n2620 185
R1534 vdd.n2623 vdd.n655 185
R1535 vdd.n660 vdd.n655 185
R1536 vdd.n2625 vdd.n2624 185
R1537 vdd.n2626 vdd.n2625 185
R1538 vdd.n646 vdd.n645 185
R1539 vdd.n647 vdd.n646 185
R1540 vdd.n2634 vdd.n2633 185
R1541 vdd.n2633 vdd.n2632 185
R1542 vdd.n2635 vdd.n644 185
R1543 vdd.n644 vdd.n641 185
R1544 vdd.n2637 vdd.n2636 185
R1545 vdd.n2638 vdd.n2637 185
R1546 vdd.n632 vdd.n631 185
R1547 vdd.n633 vdd.n632 185
R1548 vdd.n2691 vdd.n2690 185
R1549 vdd.n2690 vdd.n2689 185
R1550 vdd.n2692 vdd.n630 185
R1551 vdd.n636 vdd.n630 185
R1552 vdd.n2694 vdd.n2693 185
R1553 vdd.n2695 vdd.n2694 185
R1554 vdd.n600 vdd.n598 185
R1555 vdd.n598 vdd.n595 185
R1556 vdd.n2764 vdd.n2763 185
R1557 vdd.n2765 vdd.n2764 185
R1558 vdd.n2206 vdd.n2205 185
R1559 vdd.n2207 vdd.n2206 185
R1560 vdd.n770 vdd.n768 185
R1561 vdd.n768 vdd.n766 185
R1562 vdd.n2121 vdd.n777 185
R1563 vdd.n2132 vdd.n777 185
R1564 vdd.n2122 vdd.n786 185
R1565 vdd.n1128 vdd.n786 185
R1566 vdd.n2124 vdd.n2123 185
R1567 vdd.n2125 vdd.n2124 185
R1568 vdd.n2120 vdd.n785 185
R1569 vdd.n785 vdd.n782 185
R1570 vdd.n2119 vdd.n2118 185
R1571 vdd.n2118 vdd.n2117 185
R1572 vdd.n788 vdd.n787 185
R1573 vdd.n789 vdd.n788 185
R1574 vdd.n2110 vdd.n2109 185
R1575 vdd.n2111 vdd.n2110 185
R1576 vdd.n2108 vdd.n798 185
R1577 vdd.n798 vdd.n795 185
R1578 vdd.n2107 vdd.n2106 185
R1579 vdd.n2106 vdd.n2105 185
R1580 vdd.n800 vdd.n799 185
R1581 vdd.n808 vdd.n800 185
R1582 vdd.n2098 vdd.n2097 185
R1583 vdd.n2099 vdd.n2098 185
R1584 vdd.n2096 vdd.n809 185
R1585 vdd.n814 vdd.n809 185
R1586 vdd.n2095 vdd.n2094 185
R1587 vdd.n2094 vdd.n2093 185
R1588 vdd.n811 vdd.n810 185
R1589 vdd.n1149 vdd.n811 185
R1590 vdd.n2086 vdd.n2085 185
R1591 vdd.n2087 vdd.n2086 185
R1592 vdd.n2084 vdd.n821 185
R1593 vdd.n821 vdd.n818 185
R1594 vdd.n2083 vdd.n2082 185
R1595 vdd.n2082 vdd.n2081 185
R1596 vdd.n823 vdd.n822 185
R1597 vdd.n824 vdd.n823 185
R1598 vdd.n2074 vdd.n2073 185
R1599 vdd.n2075 vdd.n2074 185
R1600 vdd.n2071 vdd.n832 185
R1601 vdd.n838 vdd.n832 185
R1602 vdd.n2070 vdd.n2069 185
R1603 vdd.n2069 vdd.n2068 185
R1604 vdd.n835 vdd.n834 185
R1605 vdd.n845 vdd.n835 185
R1606 vdd.n2061 vdd.n2060 185
R1607 vdd.n2062 vdd.n2061 185
R1608 vdd.n2059 vdd.n846 185
R1609 vdd.n846 vdd.n842 185
R1610 vdd.n2058 vdd.n2057 185
R1611 vdd.n2057 vdd.n2056 185
R1612 vdd.n848 vdd.n847 185
R1613 vdd.n849 vdd.n848 185
R1614 vdd.n2049 vdd.n2048 185
R1615 vdd.n2050 vdd.n2049 185
R1616 vdd.n2047 vdd.n858 185
R1617 vdd.n858 vdd.n855 185
R1618 vdd.n2046 vdd.n2045 185
R1619 vdd.n2045 vdd.n2044 185
R1620 vdd.n860 vdd.n859 185
R1621 vdd.n869 vdd.n860 185
R1622 vdd.n2037 vdd.n2036 185
R1623 vdd.n2038 vdd.n2037 185
R1624 vdd.n2035 vdd.n870 185
R1625 vdd.n870 vdd.n866 185
R1626 vdd.n2137 vdd.n741 185
R1627 vdd.n2279 vdd.n741 185
R1628 vdd.n2139 vdd.n2138 185
R1629 vdd.n2141 vdd.n2140 185
R1630 vdd.n2143 vdd.n2142 185
R1631 vdd.n2145 vdd.n2144 185
R1632 vdd.n2147 vdd.n2146 185
R1633 vdd.n2149 vdd.n2148 185
R1634 vdd.n2151 vdd.n2150 185
R1635 vdd.n2153 vdd.n2152 185
R1636 vdd.n2155 vdd.n2154 185
R1637 vdd.n2157 vdd.n2156 185
R1638 vdd.n2159 vdd.n2158 185
R1639 vdd.n2161 vdd.n2160 185
R1640 vdd.n2163 vdd.n2162 185
R1641 vdd.n2165 vdd.n2164 185
R1642 vdd.n2167 vdd.n2166 185
R1643 vdd.n2169 vdd.n2168 185
R1644 vdd.n2171 vdd.n2170 185
R1645 vdd.n2173 vdd.n2172 185
R1646 vdd.n2175 vdd.n2174 185
R1647 vdd.n2177 vdd.n2176 185
R1648 vdd.n2179 vdd.n2178 185
R1649 vdd.n2181 vdd.n2180 185
R1650 vdd.n2183 vdd.n2182 185
R1651 vdd.n2185 vdd.n2184 185
R1652 vdd.n2187 vdd.n2186 185
R1653 vdd.n2189 vdd.n2188 185
R1654 vdd.n2191 vdd.n2190 185
R1655 vdd.n2193 vdd.n2192 185
R1656 vdd.n2195 vdd.n2194 185
R1657 vdd.n2197 vdd.n2196 185
R1658 vdd.n2199 vdd.n2198 185
R1659 vdd.n2201 vdd.n2200 185
R1660 vdd.n2203 vdd.n2202 185
R1661 vdd.n2204 vdd.n769 185
R1662 vdd.n2136 vdd.n767 185
R1663 vdd.n2207 vdd.n767 185
R1664 vdd.n2135 vdd.n2134 185
R1665 vdd.n2134 vdd.n766 185
R1666 vdd.n2133 vdd.n774 185
R1667 vdd.n2133 vdd.n2132 185
R1668 vdd.n1046 vdd.n775 185
R1669 vdd.n1128 vdd.n775 185
R1670 vdd.n1047 vdd.n784 185
R1671 vdd.n2125 vdd.n784 185
R1672 vdd.n1049 vdd.n1048 185
R1673 vdd.n1048 vdd.n782 185
R1674 vdd.n1050 vdd.n791 185
R1675 vdd.n2117 vdd.n791 185
R1676 vdd.n1052 vdd.n1051 185
R1677 vdd.n1051 vdd.n789 185
R1678 vdd.n1053 vdd.n797 185
R1679 vdd.n2111 vdd.n797 185
R1680 vdd.n1055 vdd.n1054 185
R1681 vdd.n1054 vdd.n795 185
R1682 vdd.n1056 vdd.n802 185
R1683 vdd.n2105 vdd.n802 185
R1684 vdd.n1058 vdd.n1057 185
R1685 vdd.n1057 vdd.n808 185
R1686 vdd.n1059 vdd.n807 185
R1687 vdd.n2099 vdd.n807 185
R1688 vdd.n1061 vdd.n1060 185
R1689 vdd.n1060 vdd.n814 185
R1690 vdd.n1062 vdd.n813 185
R1691 vdd.n2093 vdd.n813 185
R1692 vdd.n1151 vdd.n1150 185
R1693 vdd.n1150 vdd.n1149 185
R1694 vdd.n1152 vdd.n820 185
R1695 vdd.n2087 vdd.n820 185
R1696 vdd.n1154 vdd.n1153 185
R1697 vdd.n1153 vdd.n818 185
R1698 vdd.n1155 vdd.n826 185
R1699 vdd.n2081 vdd.n826 185
R1700 vdd.n1157 vdd.n1156 185
R1701 vdd.n1156 vdd.n824 185
R1702 vdd.n1158 vdd.n831 185
R1703 vdd.n2075 vdd.n831 185
R1704 vdd.n1160 vdd.n1159 185
R1705 vdd.n1159 vdd.n838 185
R1706 vdd.n1161 vdd.n837 185
R1707 vdd.n2068 vdd.n837 185
R1708 vdd.n1163 vdd.n1162 185
R1709 vdd.n1162 vdd.n845 185
R1710 vdd.n1164 vdd.n844 185
R1711 vdd.n2062 vdd.n844 185
R1712 vdd.n1166 vdd.n1165 185
R1713 vdd.n1165 vdd.n842 185
R1714 vdd.n1167 vdd.n851 185
R1715 vdd.n2056 vdd.n851 185
R1716 vdd.n1169 vdd.n1168 185
R1717 vdd.n1168 vdd.n849 185
R1718 vdd.n1170 vdd.n857 185
R1719 vdd.n2050 vdd.n857 185
R1720 vdd.n1172 vdd.n1171 185
R1721 vdd.n1171 vdd.n855 185
R1722 vdd.n1173 vdd.n862 185
R1723 vdd.n2044 vdd.n862 185
R1724 vdd.n1175 vdd.n1174 185
R1725 vdd.n1174 vdd.n869 185
R1726 vdd.n1176 vdd.n868 185
R1727 vdd.n2038 vdd.n868 185
R1728 vdd.n1178 vdd.n1177 185
R1729 vdd.n1177 vdd.n866 185
R1730 vdd.n2034 vdd.n2033 185
R1731 vdd.n872 vdd.n871 185
R1732 vdd.n1013 vdd.n1012 185
R1733 vdd.n1015 vdd.n1014 185
R1734 vdd.n1017 vdd.n1016 185
R1735 vdd.n1019 vdd.n1018 185
R1736 vdd.n1021 vdd.n1020 185
R1737 vdd.n1023 vdd.n1022 185
R1738 vdd.n1025 vdd.n1024 185
R1739 vdd.n1027 vdd.n1026 185
R1740 vdd.n1029 vdd.n1028 185
R1741 vdd.n1031 vdd.n1030 185
R1742 vdd.n1033 vdd.n1032 185
R1743 vdd.n1035 vdd.n1034 185
R1744 vdd.n1037 vdd.n1036 185
R1745 vdd.n1039 vdd.n1038 185
R1746 vdd.n1041 vdd.n1040 185
R1747 vdd.n1212 vdd.n1042 185
R1748 vdd.n1211 vdd.n1210 185
R1749 vdd.n1209 vdd.n1208 185
R1750 vdd.n1207 vdd.n1206 185
R1751 vdd.n1205 vdd.n1204 185
R1752 vdd.n1203 vdd.n1202 185
R1753 vdd.n1201 vdd.n1200 185
R1754 vdd.n1199 vdd.n1198 185
R1755 vdd.n1197 vdd.n1196 185
R1756 vdd.n1195 vdd.n1194 185
R1757 vdd.n1193 vdd.n1192 185
R1758 vdd.n1191 vdd.n1190 185
R1759 vdd.n1189 vdd.n1188 185
R1760 vdd.n1187 vdd.n1186 185
R1761 vdd.n1185 vdd.n1184 185
R1762 vdd.n1183 vdd.n1182 185
R1763 vdd.n1181 vdd.n1180 185
R1764 vdd.n1179 vdd.n906 185
R1765 vdd.n2031 vdd.n906 185
R1766 vdd.n2031 vdd.n873 179.345
R1767 vdd.n2932 vdd.n484 179.345
R1768 vdd.n291 vdd.n290 171.744
R1769 vdd.n290 vdd.n289 171.744
R1770 vdd.n289 vdd.n258 171.744
R1771 vdd.n282 vdd.n258 171.744
R1772 vdd.n282 vdd.n281 171.744
R1773 vdd.n281 vdd.n263 171.744
R1774 vdd.n274 vdd.n263 171.744
R1775 vdd.n274 vdd.n273 171.744
R1776 vdd.n273 vdd.n267 171.744
R1777 vdd.n244 vdd.n243 171.744
R1778 vdd.n243 vdd.n242 171.744
R1779 vdd.n242 vdd.n211 171.744
R1780 vdd.n235 vdd.n211 171.744
R1781 vdd.n235 vdd.n234 171.744
R1782 vdd.n234 vdd.n216 171.744
R1783 vdd.n227 vdd.n216 171.744
R1784 vdd.n227 vdd.n226 171.744
R1785 vdd.n226 vdd.n220 171.744
R1786 vdd.n201 vdd.n200 171.744
R1787 vdd.n200 vdd.n199 171.744
R1788 vdd.n199 vdd.n168 171.744
R1789 vdd.n192 vdd.n168 171.744
R1790 vdd.n192 vdd.n191 171.744
R1791 vdd.n191 vdd.n173 171.744
R1792 vdd.n184 vdd.n173 171.744
R1793 vdd.n184 vdd.n183 171.744
R1794 vdd.n183 vdd.n177 171.744
R1795 vdd.n154 vdd.n153 171.744
R1796 vdd.n153 vdd.n152 171.744
R1797 vdd.n152 vdd.n121 171.744
R1798 vdd.n145 vdd.n121 171.744
R1799 vdd.n145 vdd.n144 171.744
R1800 vdd.n144 vdd.n126 171.744
R1801 vdd.n137 vdd.n126 171.744
R1802 vdd.n137 vdd.n136 171.744
R1803 vdd.n136 vdd.n130 171.744
R1804 vdd.n112 vdd.n111 171.744
R1805 vdd.n111 vdd.n110 171.744
R1806 vdd.n110 vdd.n79 171.744
R1807 vdd.n103 vdd.n79 171.744
R1808 vdd.n103 vdd.n102 171.744
R1809 vdd.n102 vdd.n84 171.744
R1810 vdd.n95 vdd.n84 171.744
R1811 vdd.n95 vdd.n94 171.744
R1812 vdd.n94 vdd.n88 171.744
R1813 vdd.n65 vdd.n64 171.744
R1814 vdd.n64 vdd.n63 171.744
R1815 vdd.n63 vdd.n32 171.744
R1816 vdd.n56 vdd.n32 171.744
R1817 vdd.n56 vdd.n55 171.744
R1818 vdd.n55 vdd.n37 171.744
R1819 vdd.n48 vdd.n37 171.744
R1820 vdd.n48 vdd.n47 171.744
R1821 vdd.n47 vdd.n41 171.744
R1822 vdd.n1468 vdd.n1467 171.744
R1823 vdd.n1467 vdd.n1466 171.744
R1824 vdd.n1466 vdd.n1435 171.744
R1825 vdd.n1459 vdd.n1435 171.744
R1826 vdd.n1459 vdd.n1458 171.744
R1827 vdd.n1458 vdd.n1440 171.744
R1828 vdd.n1451 vdd.n1440 171.744
R1829 vdd.n1451 vdd.n1450 171.744
R1830 vdd.n1450 vdd.n1444 171.744
R1831 vdd.n1515 vdd.n1514 171.744
R1832 vdd.n1514 vdd.n1513 171.744
R1833 vdd.n1513 vdd.n1482 171.744
R1834 vdd.n1506 vdd.n1482 171.744
R1835 vdd.n1506 vdd.n1505 171.744
R1836 vdd.n1505 vdd.n1487 171.744
R1837 vdd.n1498 vdd.n1487 171.744
R1838 vdd.n1498 vdd.n1497 171.744
R1839 vdd.n1497 vdd.n1491 171.744
R1840 vdd.n1378 vdd.n1377 171.744
R1841 vdd.n1377 vdd.n1376 171.744
R1842 vdd.n1376 vdd.n1345 171.744
R1843 vdd.n1369 vdd.n1345 171.744
R1844 vdd.n1369 vdd.n1368 171.744
R1845 vdd.n1368 vdd.n1350 171.744
R1846 vdd.n1361 vdd.n1350 171.744
R1847 vdd.n1361 vdd.n1360 171.744
R1848 vdd.n1360 vdd.n1354 171.744
R1849 vdd.n1425 vdd.n1424 171.744
R1850 vdd.n1424 vdd.n1423 171.744
R1851 vdd.n1423 vdd.n1392 171.744
R1852 vdd.n1416 vdd.n1392 171.744
R1853 vdd.n1416 vdd.n1415 171.744
R1854 vdd.n1415 vdd.n1397 171.744
R1855 vdd.n1408 vdd.n1397 171.744
R1856 vdd.n1408 vdd.n1407 171.744
R1857 vdd.n1407 vdd.n1401 171.744
R1858 vdd.n1289 vdd.n1288 171.744
R1859 vdd.n1288 vdd.n1287 171.744
R1860 vdd.n1287 vdd.n1256 171.744
R1861 vdd.n1280 vdd.n1256 171.744
R1862 vdd.n1280 vdd.n1279 171.744
R1863 vdd.n1279 vdd.n1261 171.744
R1864 vdd.n1272 vdd.n1261 171.744
R1865 vdd.n1272 vdd.n1271 171.744
R1866 vdd.n1271 vdd.n1265 171.744
R1867 vdd.n1336 vdd.n1335 171.744
R1868 vdd.n1335 vdd.n1334 171.744
R1869 vdd.n1334 vdd.n1303 171.744
R1870 vdd.n1327 vdd.n1303 171.744
R1871 vdd.n1327 vdd.n1326 171.744
R1872 vdd.n1326 vdd.n1308 171.744
R1873 vdd.n1319 vdd.n1308 171.744
R1874 vdd.n1319 vdd.n1318 171.744
R1875 vdd.n1318 vdd.n1312 171.744
R1876 vdd.n3109 vdd.n334 146.341
R1877 vdd.n3107 vdd.n3106 146.341
R1878 vdd.n3104 vdd.n338 146.341
R1879 vdd.n3100 vdd.n3099 146.341
R1880 vdd.n3097 vdd.n346 146.341
R1881 vdd.n3093 vdd.n3092 146.341
R1882 vdd.n3090 vdd.n353 146.341
R1883 vdd.n3086 vdd.n3085 146.341
R1884 vdd.n3083 vdd.n360 146.341
R1885 vdd.n371 vdd.n368 146.341
R1886 vdd.n3075 vdd.n3074 146.341
R1887 vdd.n3072 vdd.n373 146.341
R1888 vdd.n3068 vdd.n3067 146.341
R1889 vdd.n3065 vdd.n379 146.341
R1890 vdd.n3061 vdd.n3060 146.341
R1891 vdd.n3058 vdd.n386 146.341
R1892 vdd.n3054 vdd.n3053 146.341
R1893 vdd.n3051 vdd.n393 146.341
R1894 vdd.n3047 vdd.n3046 146.341
R1895 vdd.n3044 vdd.n400 146.341
R1896 vdd.n411 vdd.n408 146.341
R1897 vdd.n3036 vdd.n3035 146.341
R1898 vdd.n3033 vdd.n413 146.341
R1899 vdd.n3029 vdd.n3028 146.341
R1900 vdd.n3026 vdd.n419 146.341
R1901 vdd.n3022 vdd.n3021 146.341
R1902 vdd.n3019 vdd.n426 146.341
R1903 vdd.n3015 vdd.n3014 146.341
R1904 vdd.n3012 vdd.n433 146.341
R1905 vdd.n3008 vdd.n3007 146.341
R1906 vdd.n3005 vdd.n440 146.341
R1907 vdd.n2942 vdd.n478 146.341
R1908 vdd.n2942 vdd.n474 146.341
R1909 vdd.n2948 vdd.n474 146.341
R1910 vdd.n2948 vdd.n466 146.341
R1911 vdd.n2959 vdd.n466 146.341
R1912 vdd.n2959 vdd.n462 146.341
R1913 vdd.n2965 vdd.n462 146.341
R1914 vdd.n2965 vdd.n454 146.341
R1915 vdd.n2975 vdd.n454 146.341
R1916 vdd.n2975 vdd.n455 146.341
R1917 vdd.n455 vdd.n305 146.341
R1918 vdd.n306 vdd.n305 146.341
R1919 vdd.n307 vdd.n306 146.341
R1920 vdd.n448 vdd.n307 146.341
R1921 vdd.n448 vdd.n315 146.341
R1922 vdd.n316 vdd.n315 146.341
R1923 vdd.n317 vdd.n316 146.341
R1924 vdd.n445 vdd.n317 146.341
R1925 vdd.n445 vdd.n326 146.341
R1926 vdd.n327 vdd.n326 146.341
R1927 vdd.n328 vdd.n327 146.341
R1928 vdd.n2931 vdd.n483 146.341
R1929 vdd.n2931 vdd.n517 146.341
R1930 vdd.n523 vdd.n522 146.341
R1931 vdd.n2924 vdd.n2923 146.341
R1932 vdd.n2920 vdd.n2919 146.341
R1933 vdd.n2916 vdd.n2915 146.341
R1934 vdd.n2912 vdd.n2911 146.341
R1935 vdd.n2908 vdd.n2907 146.341
R1936 vdd.n2904 vdd.n2903 146.341
R1937 vdd.n2900 vdd.n2899 146.341
R1938 vdd.n2891 vdd.n2890 146.341
R1939 vdd.n2888 vdd.n2887 146.341
R1940 vdd.n2884 vdd.n2883 146.341
R1941 vdd.n2880 vdd.n2879 146.341
R1942 vdd.n2876 vdd.n2875 146.341
R1943 vdd.n2872 vdd.n2871 146.341
R1944 vdd.n2868 vdd.n2867 146.341
R1945 vdd.n2864 vdd.n2863 146.341
R1946 vdd.n2860 vdd.n2859 146.341
R1947 vdd.n2856 vdd.n2855 146.341
R1948 vdd.n2852 vdd.n2851 146.341
R1949 vdd.n2845 vdd.n2844 146.341
R1950 vdd.n2842 vdd.n2841 146.341
R1951 vdd.n2838 vdd.n2837 146.341
R1952 vdd.n2834 vdd.n2833 146.341
R1953 vdd.n2830 vdd.n2829 146.341
R1954 vdd.n2826 vdd.n2825 146.341
R1955 vdd.n2822 vdd.n2821 146.341
R1956 vdd.n2818 vdd.n2817 146.341
R1957 vdd.n2814 vdd.n2813 146.341
R1958 vdd.n2810 vdd.n2809 146.341
R1959 vdd.n2806 vdd.n515 146.341
R1960 vdd.n2940 vdd.n479 146.341
R1961 vdd.n2940 vdd.n472 146.341
R1962 vdd.n2951 vdd.n472 146.341
R1963 vdd.n2951 vdd.n468 146.341
R1964 vdd.n2957 vdd.n468 146.341
R1965 vdd.n2957 vdd.n461 146.341
R1966 vdd.n2967 vdd.n461 146.341
R1967 vdd.n2967 vdd.n457 146.341
R1968 vdd.n2973 vdd.n457 146.341
R1969 vdd.n2973 vdd.n302 146.341
R1970 vdd.n3136 vdd.n302 146.341
R1971 vdd.n3136 vdd.n303 146.341
R1972 vdd.n3132 vdd.n303 146.341
R1973 vdd.n3132 vdd.n309 146.341
R1974 vdd.n3128 vdd.n309 146.341
R1975 vdd.n3128 vdd.n314 146.341
R1976 vdd.n3124 vdd.n314 146.341
R1977 vdd.n3124 vdd.n319 146.341
R1978 vdd.n3120 vdd.n319 146.341
R1979 vdd.n3120 vdd.n325 146.341
R1980 vdd.n3116 vdd.n325 146.341
R1981 vdd.n1992 vdd.n1991 146.341
R1982 vdd.n1989 vdd.n1986 146.341
R1983 vdd.n1984 vdd.n917 146.341
R1984 vdd.n1980 vdd.n1979 146.341
R1985 vdd.n1977 vdd.n921 146.341
R1986 vdd.n1973 vdd.n1972 146.341
R1987 vdd.n1970 vdd.n928 146.341
R1988 vdd.n1966 vdd.n1965 146.341
R1989 vdd.n1963 vdd.n935 146.341
R1990 vdd.n946 vdd.n943 146.341
R1991 vdd.n1955 vdd.n1954 146.341
R1992 vdd.n1952 vdd.n948 146.341
R1993 vdd.n1948 vdd.n1947 146.341
R1994 vdd.n1945 vdd.n954 146.341
R1995 vdd.n1941 vdd.n1940 146.341
R1996 vdd.n1938 vdd.n961 146.341
R1997 vdd.n1934 vdd.n1933 146.341
R1998 vdd.n1931 vdd.n968 146.341
R1999 vdd.n1927 vdd.n1926 146.341
R2000 vdd.n1924 vdd.n975 146.341
R2001 vdd.n986 vdd.n983 146.341
R2002 vdd.n1916 vdd.n1915 146.341
R2003 vdd.n1913 vdd.n988 146.341
R2004 vdd.n1909 vdd.n1908 146.341
R2005 vdd.n1906 vdd.n994 146.341
R2006 vdd.n1902 vdd.n1901 146.341
R2007 vdd.n1899 vdd.n1001 146.341
R2008 vdd.n1895 vdd.n1894 146.341
R2009 vdd.n1892 vdd.n1008 146.341
R2010 vdd.n1219 vdd.n1217 146.341
R2011 vdd.n1222 vdd.n1221 146.341
R2012 vdd.n1793 vdd.n1553 146.341
R2013 vdd.n1793 vdd.n1549 146.341
R2014 vdd.n1799 vdd.n1549 146.341
R2015 vdd.n1799 vdd.n1541 146.341
R2016 vdd.n1810 vdd.n1541 146.341
R2017 vdd.n1810 vdd.n1537 146.341
R2018 vdd.n1816 vdd.n1537 146.341
R2019 vdd.n1816 vdd.n1531 146.341
R2020 vdd.n1828 vdd.n1531 146.341
R2021 vdd.n1828 vdd.n1527 146.341
R2022 vdd.n1834 vdd.n1527 146.341
R2023 vdd.n1834 vdd.n1248 146.341
R2024 vdd.n1844 vdd.n1248 146.341
R2025 vdd.n1844 vdd.n1244 146.341
R2026 vdd.n1850 vdd.n1244 146.341
R2027 vdd.n1850 vdd.n1238 146.341
R2028 vdd.n1861 vdd.n1238 146.341
R2029 vdd.n1861 vdd.n1233 146.341
R2030 vdd.n1869 vdd.n1233 146.341
R2031 vdd.n1869 vdd.n1224 146.341
R2032 vdd.n1880 vdd.n1224 146.341
R2033 vdd.n1782 vdd.n1558 146.341
R2034 vdd.n1782 vdd.n1591 146.341
R2035 vdd.n1595 vdd.n1594 146.341
R2036 vdd.n1597 vdd.n1596 146.341
R2037 vdd.n1601 vdd.n1600 146.341
R2038 vdd.n1603 vdd.n1602 146.341
R2039 vdd.n1607 vdd.n1606 146.341
R2040 vdd.n1609 vdd.n1608 146.341
R2041 vdd.n1613 vdd.n1612 146.341
R2042 vdd.n1615 vdd.n1614 146.341
R2043 vdd.n1621 vdd.n1620 146.341
R2044 vdd.n1623 vdd.n1622 146.341
R2045 vdd.n1627 vdd.n1626 146.341
R2046 vdd.n1629 vdd.n1628 146.341
R2047 vdd.n1633 vdd.n1632 146.341
R2048 vdd.n1635 vdd.n1634 146.341
R2049 vdd.n1639 vdd.n1638 146.341
R2050 vdd.n1641 vdd.n1640 146.341
R2051 vdd.n1645 vdd.n1644 146.341
R2052 vdd.n1647 vdd.n1646 146.341
R2053 vdd.n1719 vdd.n1650 146.341
R2054 vdd.n1652 vdd.n1651 146.341
R2055 vdd.n1656 vdd.n1655 146.341
R2056 vdd.n1658 vdd.n1657 146.341
R2057 vdd.n1662 vdd.n1661 146.341
R2058 vdd.n1664 vdd.n1663 146.341
R2059 vdd.n1668 vdd.n1667 146.341
R2060 vdd.n1670 vdd.n1669 146.341
R2061 vdd.n1674 vdd.n1673 146.341
R2062 vdd.n1676 vdd.n1675 146.341
R2063 vdd.n1680 vdd.n1679 146.341
R2064 vdd.n1681 vdd.n1589 146.341
R2065 vdd.n1791 vdd.n1554 146.341
R2066 vdd.n1791 vdd.n1547 146.341
R2067 vdd.n1802 vdd.n1547 146.341
R2068 vdd.n1802 vdd.n1543 146.341
R2069 vdd.n1808 vdd.n1543 146.341
R2070 vdd.n1808 vdd.n1536 146.341
R2071 vdd.n1819 vdd.n1536 146.341
R2072 vdd.n1819 vdd.n1532 146.341
R2073 vdd.n1826 vdd.n1532 146.341
R2074 vdd.n1826 vdd.n1525 146.341
R2075 vdd.n1836 vdd.n1525 146.341
R2076 vdd.n1836 vdd.n1251 146.341
R2077 vdd.n1842 vdd.n1251 146.341
R2078 vdd.n1842 vdd.n1243 146.341
R2079 vdd.n1853 vdd.n1243 146.341
R2080 vdd.n1853 vdd.n1239 146.341
R2081 vdd.n1859 vdd.n1239 146.341
R2082 vdd.n1859 vdd.n1231 146.341
R2083 vdd.n1872 vdd.n1231 146.341
R2084 vdd.n1872 vdd.n1226 146.341
R2085 vdd.n1878 vdd.n1226 146.341
R2086 vdd.n1043 vdd.t17 127.284
R2087 vdd.n771 vdd.t50 127.284
R2088 vdd.n1063 vdd.t31 127.284
R2089 vdd.n762 vdd.t67 127.284
R2090 vdd.n662 vdd.t37 127.284
R2091 vdd.n662 vdd.t38 127.284
R2092 vdd.n2318 vdd.t62 127.284
R2093 vdd.n622 vdd.t70 127.284
R2094 vdd.n2315 vdd.t55 127.284
R2095 vdd.n589 vdd.t12 127.284
R2096 vdd.n833 vdd.t58 127.284
R2097 vdd.n833 vdd.t59 127.284
R2098 vdd.n22 vdd.n20 117.314
R2099 vdd.n17 vdd.n15 117.314
R2100 vdd.n27 vdd.n26 116.927
R2101 vdd.n24 vdd.n23 116.927
R2102 vdd.n22 vdd.n21 116.927
R2103 vdd.n17 vdd.n16 116.927
R2104 vdd.n19 vdd.n18 116.927
R2105 vdd.n27 vdd.n25 116.927
R2106 vdd.n1044 vdd.t16 111.188
R2107 vdd.n772 vdd.t51 111.188
R2108 vdd.n1064 vdd.t30 111.188
R2109 vdd.n763 vdd.t68 111.188
R2110 vdd.n2319 vdd.t61 111.188
R2111 vdd.n623 vdd.t71 111.188
R2112 vdd.n2316 vdd.t54 111.188
R2113 vdd.n590 vdd.t13 111.188
R2114 vdd.n2560 vdd.n717 99.5127
R2115 vdd.n2560 vdd.n715 99.5127
R2116 vdd.n2564 vdd.n715 99.5127
R2117 vdd.n2564 vdd.n706 99.5127
R2118 vdd.n2572 vdd.n706 99.5127
R2119 vdd.n2572 vdd.n704 99.5127
R2120 vdd.n2576 vdd.n704 99.5127
R2121 vdd.n2576 vdd.n694 99.5127
R2122 vdd.n2584 vdd.n694 99.5127
R2123 vdd.n2584 vdd.n692 99.5127
R2124 vdd.n2588 vdd.n692 99.5127
R2125 vdd.n2588 vdd.n682 99.5127
R2126 vdd.n2596 vdd.n682 99.5127
R2127 vdd.n2596 vdd.n680 99.5127
R2128 vdd.n2600 vdd.n680 99.5127
R2129 vdd.n2600 vdd.n671 99.5127
R2130 vdd.n2608 vdd.n671 99.5127
R2131 vdd.n2608 vdd.n669 99.5127
R2132 vdd.n2612 vdd.n669 99.5127
R2133 vdd.n2612 vdd.n657 99.5127
R2134 vdd.n2621 vdd.n657 99.5127
R2135 vdd.n2621 vdd.n655 99.5127
R2136 vdd.n2625 vdd.n655 99.5127
R2137 vdd.n2625 vdd.n646 99.5127
R2138 vdd.n2633 vdd.n646 99.5127
R2139 vdd.n2633 vdd.n644 99.5127
R2140 vdd.n2637 vdd.n644 99.5127
R2141 vdd.n2637 vdd.n632 99.5127
R2142 vdd.n2690 vdd.n632 99.5127
R2143 vdd.n2690 vdd.n630 99.5127
R2144 vdd.n2694 vdd.n630 99.5127
R2145 vdd.n2694 vdd.n598 99.5127
R2146 vdd.n2764 vdd.n598 99.5127
R2147 vdd.n2760 vdd.n599 99.5127
R2148 vdd.n2758 vdd.n2757 99.5127
R2149 vdd.n2755 vdd.n603 99.5127
R2150 vdd.n2751 vdd.n2750 99.5127
R2151 vdd.n2748 vdd.n606 99.5127
R2152 vdd.n2744 vdd.n2743 99.5127
R2153 vdd.n2741 vdd.n609 99.5127
R2154 vdd.n2737 vdd.n2736 99.5127
R2155 vdd.n2734 vdd.n2732 99.5127
R2156 vdd.n2730 vdd.n612 99.5127
R2157 vdd.n2726 vdd.n2725 99.5127
R2158 vdd.n2723 vdd.n615 99.5127
R2159 vdd.n2719 vdd.n2718 99.5127
R2160 vdd.n2716 vdd.n618 99.5127
R2161 vdd.n2712 vdd.n2711 99.5127
R2162 vdd.n2709 vdd.n621 99.5127
R2163 vdd.n2704 vdd.n2703 99.5127
R2164 vdd.n2481 vdd.n719 99.5127
R2165 vdd.n2477 vdd.n719 99.5127
R2166 vdd.n2477 vdd.n713 99.5127
R2167 vdd.n2421 vdd.n713 99.5127
R2168 vdd.n2421 vdd.n708 99.5127
R2169 vdd.n2424 vdd.n708 99.5127
R2170 vdd.n2424 vdd.n702 99.5127
R2171 vdd.n2427 vdd.n702 99.5127
R2172 vdd.n2427 vdd.n696 99.5127
R2173 vdd.n2460 vdd.n696 99.5127
R2174 vdd.n2460 vdd.n689 99.5127
R2175 vdd.n2456 vdd.n689 99.5127
R2176 vdd.n2456 vdd.n683 99.5127
R2177 vdd.n2453 vdd.n683 99.5127
R2178 vdd.n2453 vdd.n678 99.5127
R2179 vdd.n2450 vdd.n678 99.5127
R2180 vdd.n2450 vdd.n673 99.5127
R2181 vdd.n2447 vdd.n673 99.5127
R2182 vdd.n2447 vdd.n666 99.5127
R2183 vdd.n2444 vdd.n666 99.5127
R2184 vdd.n2444 vdd.n658 99.5127
R2185 vdd.n2441 vdd.n658 99.5127
R2186 vdd.n2441 vdd.n653 99.5127
R2187 vdd.n2438 vdd.n653 99.5127
R2188 vdd.n2438 vdd.n648 99.5127
R2189 vdd.n2435 vdd.n648 99.5127
R2190 vdd.n2435 vdd.n642 99.5127
R2191 vdd.n2432 vdd.n642 99.5127
R2192 vdd.n2432 vdd.n634 99.5127
R2193 vdd.n634 vdd.n627 99.5127
R2194 vdd.n2696 vdd.n627 99.5127
R2195 vdd.n2697 vdd.n2696 99.5127
R2196 vdd.n2697 vdd.n596 99.5127
R2197 vdd.n2314 vdd.n2313 99.5127
R2198 vdd.n2545 vdd.n2313 99.5127
R2199 vdd.n2543 vdd.n2542 99.5127
R2200 vdd.n2539 vdd.n2538 99.5127
R2201 vdd.n2535 vdd.n2534 99.5127
R2202 vdd.n2531 vdd.n2530 99.5127
R2203 vdd.n2527 vdd.n2526 99.5127
R2204 vdd.n2523 vdd.n2522 99.5127
R2205 vdd.n2519 vdd.n2518 99.5127
R2206 vdd.n2515 vdd.n2514 99.5127
R2207 vdd.n2511 vdd.n2510 99.5127
R2208 vdd.n2507 vdd.n2506 99.5127
R2209 vdd.n2503 vdd.n2502 99.5127
R2210 vdd.n2499 vdd.n2498 99.5127
R2211 vdd.n2495 vdd.n2494 99.5127
R2212 vdd.n2491 vdd.n2490 99.5127
R2213 vdd.n2486 vdd.n2485 99.5127
R2214 vdd.n2278 vdd.n760 99.5127
R2215 vdd.n2274 vdd.n2273 99.5127
R2216 vdd.n2270 vdd.n2269 99.5127
R2217 vdd.n2266 vdd.n2265 99.5127
R2218 vdd.n2262 vdd.n2261 99.5127
R2219 vdd.n2258 vdd.n2257 99.5127
R2220 vdd.n2254 vdd.n2253 99.5127
R2221 vdd.n2250 vdd.n2249 99.5127
R2222 vdd.n2246 vdd.n2245 99.5127
R2223 vdd.n2242 vdd.n2241 99.5127
R2224 vdd.n2238 vdd.n2237 99.5127
R2225 vdd.n2234 vdd.n2233 99.5127
R2226 vdd.n2230 vdd.n2229 99.5127
R2227 vdd.n2226 vdd.n2225 99.5127
R2228 vdd.n2222 vdd.n2221 99.5127
R2229 vdd.n2218 vdd.n2217 99.5127
R2230 vdd.n2213 vdd.n2212 99.5127
R2231 vdd.n1099 vdd.n867 99.5127
R2232 vdd.n1102 vdd.n867 99.5127
R2233 vdd.n1102 vdd.n861 99.5127
R2234 vdd.n1105 vdd.n861 99.5127
R2235 vdd.n1105 vdd.n856 99.5127
R2236 vdd.n1108 vdd.n856 99.5127
R2237 vdd.n1108 vdd.n850 99.5127
R2238 vdd.n1111 vdd.n850 99.5127
R2239 vdd.n1111 vdd.n843 99.5127
R2240 vdd.n1114 vdd.n843 99.5127
R2241 vdd.n1114 vdd.n836 99.5127
R2242 vdd.n1117 vdd.n836 99.5127
R2243 vdd.n1117 vdd.n830 99.5127
R2244 vdd.n1120 vdd.n830 99.5127
R2245 vdd.n1120 vdd.n825 99.5127
R2246 vdd.n1123 vdd.n825 99.5127
R2247 vdd.n1123 vdd.n819 99.5127
R2248 vdd.n1148 vdd.n819 99.5127
R2249 vdd.n1148 vdd.n812 99.5127
R2250 vdd.n1144 vdd.n812 99.5127
R2251 vdd.n1144 vdd.n806 99.5127
R2252 vdd.n1141 vdd.n806 99.5127
R2253 vdd.n1141 vdd.n801 99.5127
R2254 vdd.n1138 vdd.n801 99.5127
R2255 vdd.n1138 vdd.n796 99.5127
R2256 vdd.n1135 vdd.n796 99.5127
R2257 vdd.n1135 vdd.n790 99.5127
R2258 vdd.n1132 vdd.n790 99.5127
R2259 vdd.n1132 vdd.n783 99.5127
R2260 vdd.n1129 vdd.n783 99.5127
R2261 vdd.n1129 vdd.n776 99.5127
R2262 vdd.n776 vdd.n765 99.5127
R2263 vdd.n2208 vdd.n765 99.5127
R2264 vdd.n908 vdd.n907 99.5127
R2265 vdd.n2024 vdd.n907 99.5127
R2266 vdd.n2022 vdd.n2021 99.5127
R2267 vdd.n2018 vdd.n2017 99.5127
R2268 vdd.n2014 vdd.n2013 99.5127
R2269 vdd.n2010 vdd.n2009 99.5127
R2270 vdd.n2006 vdd.n2005 99.5127
R2271 vdd.n2002 vdd.n2001 99.5127
R2272 vdd.n1998 vdd.n1997 99.5127
R2273 vdd.n1066 vdd.n1065 99.5127
R2274 vdd.n1070 vdd.n1069 99.5127
R2275 vdd.n1074 vdd.n1073 99.5127
R2276 vdd.n1078 vdd.n1077 99.5127
R2277 vdd.n1082 vdd.n1081 99.5127
R2278 vdd.n1086 vdd.n1085 99.5127
R2279 vdd.n1090 vdd.n1089 99.5127
R2280 vdd.n1095 vdd.n1094 99.5127
R2281 vdd.n2039 vdd.n865 99.5127
R2282 vdd.n2039 vdd.n863 99.5127
R2283 vdd.n2043 vdd.n863 99.5127
R2284 vdd.n2043 vdd.n854 99.5127
R2285 vdd.n2051 vdd.n854 99.5127
R2286 vdd.n2051 vdd.n852 99.5127
R2287 vdd.n2055 vdd.n852 99.5127
R2288 vdd.n2055 vdd.n841 99.5127
R2289 vdd.n2063 vdd.n841 99.5127
R2290 vdd.n2063 vdd.n839 99.5127
R2291 vdd.n2067 vdd.n839 99.5127
R2292 vdd.n2067 vdd.n829 99.5127
R2293 vdd.n2076 vdd.n829 99.5127
R2294 vdd.n2076 vdd.n827 99.5127
R2295 vdd.n2080 vdd.n827 99.5127
R2296 vdd.n2080 vdd.n817 99.5127
R2297 vdd.n2088 vdd.n817 99.5127
R2298 vdd.n2088 vdd.n815 99.5127
R2299 vdd.n2092 vdd.n815 99.5127
R2300 vdd.n2092 vdd.n805 99.5127
R2301 vdd.n2100 vdd.n805 99.5127
R2302 vdd.n2100 vdd.n803 99.5127
R2303 vdd.n2104 vdd.n803 99.5127
R2304 vdd.n2104 vdd.n794 99.5127
R2305 vdd.n2112 vdd.n794 99.5127
R2306 vdd.n2112 vdd.n792 99.5127
R2307 vdd.n2116 vdd.n792 99.5127
R2308 vdd.n2116 vdd.n781 99.5127
R2309 vdd.n2126 vdd.n781 99.5127
R2310 vdd.n2126 vdd.n778 99.5127
R2311 vdd.n2131 vdd.n778 99.5127
R2312 vdd.n2131 vdd.n779 99.5127
R2313 vdd.n779 vdd.n759 99.5127
R2314 vdd.n2680 vdd.n2679 99.5127
R2315 vdd.n2677 vdd.n2643 99.5127
R2316 vdd.n2673 vdd.n2672 99.5127
R2317 vdd.n2670 vdd.n2646 99.5127
R2318 vdd.n2666 vdd.n2665 99.5127
R2319 vdd.n2663 vdd.n2649 99.5127
R2320 vdd.n2659 vdd.n2658 99.5127
R2321 vdd.n2656 vdd.n2653 99.5127
R2322 vdd.n2797 vdd.n577 99.5127
R2323 vdd.n2795 vdd.n2794 99.5127
R2324 vdd.n2792 vdd.n579 99.5127
R2325 vdd.n2788 vdd.n2787 99.5127
R2326 vdd.n2785 vdd.n582 99.5127
R2327 vdd.n2781 vdd.n2780 99.5127
R2328 vdd.n2778 vdd.n585 99.5127
R2329 vdd.n2774 vdd.n2773 99.5127
R2330 vdd.n2771 vdd.n588 99.5127
R2331 vdd.n2386 vdd.n720 99.5127
R2332 vdd.n2475 vdd.n720 99.5127
R2333 vdd.n2475 vdd.n714 99.5127
R2334 vdd.n2471 vdd.n714 99.5127
R2335 vdd.n2471 vdd.n709 99.5127
R2336 vdd.n2468 vdd.n709 99.5127
R2337 vdd.n2468 vdd.n703 99.5127
R2338 vdd.n2465 vdd.n703 99.5127
R2339 vdd.n2465 vdd.n697 99.5127
R2340 vdd.n2462 vdd.n697 99.5127
R2341 vdd.n2462 vdd.n690 99.5127
R2342 vdd.n2418 vdd.n690 99.5127
R2343 vdd.n2418 vdd.n684 99.5127
R2344 vdd.n2415 vdd.n684 99.5127
R2345 vdd.n2415 vdd.n679 99.5127
R2346 vdd.n2412 vdd.n679 99.5127
R2347 vdd.n2412 vdd.n674 99.5127
R2348 vdd.n2409 vdd.n674 99.5127
R2349 vdd.n2409 vdd.n667 99.5127
R2350 vdd.n2406 vdd.n667 99.5127
R2351 vdd.n2406 vdd.n659 99.5127
R2352 vdd.n2403 vdd.n659 99.5127
R2353 vdd.n2403 vdd.n654 99.5127
R2354 vdd.n2400 vdd.n654 99.5127
R2355 vdd.n2400 vdd.n649 99.5127
R2356 vdd.n2397 vdd.n649 99.5127
R2357 vdd.n2397 vdd.n643 99.5127
R2358 vdd.n2394 vdd.n643 99.5127
R2359 vdd.n2394 vdd.n635 99.5127
R2360 vdd.n2391 vdd.n635 99.5127
R2361 vdd.n2391 vdd.n628 99.5127
R2362 vdd.n628 vdd.n594 99.5127
R2363 vdd.n2766 vdd.n594 99.5127
R2364 vdd.n2321 vdd.n723 99.5127
R2365 vdd.n2325 vdd.n2324 99.5127
R2366 vdd.n2329 vdd.n2328 99.5127
R2367 vdd.n2333 vdd.n2332 99.5127
R2368 vdd.n2337 vdd.n2336 99.5127
R2369 vdd.n2341 vdd.n2340 99.5127
R2370 vdd.n2345 vdd.n2344 99.5127
R2371 vdd.n2349 vdd.n2348 99.5127
R2372 vdd.n2353 vdd.n2352 99.5127
R2373 vdd.n2357 vdd.n2356 99.5127
R2374 vdd.n2361 vdd.n2360 99.5127
R2375 vdd.n2365 vdd.n2364 99.5127
R2376 vdd.n2369 vdd.n2368 99.5127
R2377 vdd.n2373 vdd.n2372 99.5127
R2378 vdd.n2377 vdd.n2376 99.5127
R2379 vdd.n2381 vdd.n2380 99.5127
R2380 vdd.n2383 vdd.n2312 99.5127
R2381 vdd.n2558 vdd.n721 99.5127
R2382 vdd.n2558 vdd.n712 99.5127
R2383 vdd.n2566 vdd.n712 99.5127
R2384 vdd.n2566 vdd.n710 99.5127
R2385 vdd.n2570 vdd.n710 99.5127
R2386 vdd.n2570 vdd.n700 99.5127
R2387 vdd.n2578 vdd.n700 99.5127
R2388 vdd.n2578 vdd.n698 99.5127
R2389 vdd.n2582 vdd.n698 99.5127
R2390 vdd.n2582 vdd.n688 99.5127
R2391 vdd.n2590 vdd.n688 99.5127
R2392 vdd.n2590 vdd.n686 99.5127
R2393 vdd.n2594 vdd.n686 99.5127
R2394 vdd.n2594 vdd.n677 99.5127
R2395 vdd.n2602 vdd.n677 99.5127
R2396 vdd.n2602 vdd.n675 99.5127
R2397 vdd.n2606 vdd.n675 99.5127
R2398 vdd.n2606 vdd.n664 99.5127
R2399 vdd.n2614 vdd.n664 99.5127
R2400 vdd.n2614 vdd.n661 99.5127
R2401 vdd.n2619 vdd.n661 99.5127
R2402 vdd.n2619 vdd.n652 99.5127
R2403 vdd.n2627 vdd.n652 99.5127
R2404 vdd.n2627 vdd.n650 99.5127
R2405 vdd.n2631 vdd.n650 99.5127
R2406 vdd.n2631 vdd.n640 99.5127
R2407 vdd.n2639 vdd.n640 99.5127
R2408 vdd.n2639 vdd.n637 99.5127
R2409 vdd.n2688 vdd.n637 99.5127
R2410 vdd.n2688 vdd.n638 99.5127
R2411 vdd.n638 vdd.n629 99.5127
R2412 vdd.n2683 vdd.n629 99.5127
R2413 vdd.n2683 vdd.n597 99.5127
R2414 vdd.n2202 vdd.n2201 99.5127
R2415 vdd.n2198 vdd.n2197 99.5127
R2416 vdd.n2194 vdd.n2193 99.5127
R2417 vdd.n2190 vdd.n2189 99.5127
R2418 vdd.n2186 vdd.n2185 99.5127
R2419 vdd.n2182 vdd.n2181 99.5127
R2420 vdd.n2178 vdd.n2177 99.5127
R2421 vdd.n2174 vdd.n2173 99.5127
R2422 vdd.n2170 vdd.n2169 99.5127
R2423 vdd.n2166 vdd.n2165 99.5127
R2424 vdd.n2162 vdd.n2161 99.5127
R2425 vdd.n2158 vdd.n2157 99.5127
R2426 vdd.n2154 vdd.n2153 99.5127
R2427 vdd.n2150 vdd.n2149 99.5127
R2428 vdd.n2146 vdd.n2145 99.5127
R2429 vdd.n2142 vdd.n2141 99.5127
R2430 vdd.n2138 vdd.n741 99.5127
R2431 vdd.n1177 vdd.n868 99.5127
R2432 vdd.n1174 vdd.n868 99.5127
R2433 vdd.n1174 vdd.n862 99.5127
R2434 vdd.n1171 vdd.n862 99.5127
R2435 vdd.n1171 vdd.n857 99.5127
R2436 vdd.n1168 vdd.n857 99.5127
R2437 vdd.n1168 vdd.n851 99.5127
R2438 vdd.n1165 vdd.n851 99.5127
R2439 vdd.n1165 vdd.n844 99.5127
R2440 vdd.n1162 vdd.n844 99.5127
R2441 vdd.n1162 vdd.n837 99.5127
R2442 vdd.n1159 vdd.n837 99.5127
R2443 vdd.n1159 vdd.n831 99.5127
R2444 vdd.n1156 vdd.n831 99.5127
R2445 vdd.n1156 vdd.n826 99.5127
R2446 vdd.n1153 vdd.n826 99.5127
R2447 vdd.n1153 vdd.n820 99.5127
R2448 vdd.n1150 vdd.n820 99.5127
R2449 vdd.n1150 vdd.n813 99.5127
R2450 vdd.n1060 vdd.n813 99.5127
R2451 vdd.n1060 vdd.n807 99.5127
R2452 vdd.n1057 vdd.n807 99.5127
R2453 vdd.n1057 vdd.n802 99.5127
R2454 vdd.n1054 vdd.n802 99.5127
R2455 vdd.n1054 vdd.n797 99.5127
R2456 vdd.n1051 vdd.n797 99.5127
R2457 vdd.n1051 vdd.n791 99.5127
R2458 vdd.n1048 vdd.n791 99.5127
R2459 vdd.n1048 vdd.n784 99.5127
R2460 vdd.n784 vdd.n775 99.5127
R2461 vdd.n2133 vdd.n775 99.5127
R2462 vdd.n2134 vdd.n2133 99.5127
R2463 vdd.n2134 vdd.n767 99.5127
R2464 vdd.n1012 vdd.n872 99.5127
R2465 vdd.n1016 vdd.n1015 99.5127
R2466 vdd.n1020 vdd.n1019 99.5127
R2467 vdd.n1024 vdd.n1023 99.5127
R2468 vdd.n1028 vdd.n1027 99.5127
R2469 vdd.n1032 vdd.n1031 99.5127
R2470 vdd.n1036 vdd.n1035 99.5127
R2471 vdd.n1040 vdd.n1039 99.5127
R2472 vdd.n1210 vdd.n1042 99.5127
R2473 vdd.n1208 vdd.n1207 99.5127
R2474 vdd.n1204 vdd.n1203 99.5127
R2475 vdd.n1200 vdd.n1199 99.5127
R2476 vdd.n1196 vdd.n1195 99.5127
R2477 vdd.n1192 vdd.n1191 99.5127
R2478 vdd.n1188 vdd.n1187 99.5127
R2479 vdd.n1184 vdd.n1183 99.5127
R2480 vdd.n1180 vdd.n906 99.5127
R2481 vdd.n2037 vdd.n870 99.5127
R2482 vdd.n2037 vdd.n860 99.5127
R2483 vdd.n2045 vdd.n860 99.5127
R2484 vdd.n2045 vdd.n858 99.5127
R2485 vdd.n2049 vdd.n858 99.5127
R2486 vdd.n2049 vdd.n848 99.5127
R2487 vdd.n2057 vdd.n848 99.5127
R2488 vdd.n2057 vdd.n846 99.5127
R2489 vdd.n2061 vdd.n846 99.5127
R2490 vdd.n2061 vdd.n835 99.5127
R2491 vdd.n2069 vdd.n835 99.5127
R2492 vdd.n2069 vdd.n832 99.5127
R2493 vdd.n2074 vdd.n832 99.5127
R2494 vdd.n2074 vdd.n823 99.5127
R2495 vdd.n2082 vdd.n823 99.5127
R2496 vdd.n2082 vdd.n821 99.5127
R2497 vdd.n2086 vdd.n821 99.5127
R2498 vdd.n2086 vdd.n811 99.5127
R2499 vdd.n2094 vdd.n811 99.5127
R2500 vdd.n2094 vdd.n809 99.5127
R2501 vdd.n2098 vdd.n809 99.5127
R2502 vdd.n2098 vdd.n800 99.5127
R2503 vdd.n2106 vdd.n800 99.5127
R2504 vdd.n2106 vdd.n798 99.5127
R2505 vdd.n2110 vdd.n798 99.5127
R2506 vdd.n2110 vdd.n788 99.5127
R2507 vdd.n2118 vdd.n788 99.5127
R2508 vdd.n2118 vdd.n785 99.5127
R2509 vdd.n2124 vdd.n785 99.5127
R2510 vdd.n2124 vdd.n786 99.5127
R2511 vdd.n786 vdd.n777 99.5127
R2512 vdd.n777 vdd.n768 99.5127
R2513 vdd.n2206 vdd.n768 99.5127
R2514 vdd.n9 vdd.n7 98.9633
R2515 vdd.n2 vdd.n0 98.9633
R2516 vdd.n9 vdd.n8 98.6055
R2517 vdd.n11 vdd.n10 98.6055
R2518 vdd.n13 vdd.n12 98.6055
R2519 vdd.n6 vdd.n5 98.6055
R2520 vdd.n4 vdd.n3 98.6055
R2521 vdd.n2 vdd.n1 98.6055
R2522 vdd.t184 vdd.n267 85.8723
R2523 vdd.t170 vdd.n220 85.8723
R2524 vdd.t85 vdd.n177 85.8723
R2525 vdd.t163 vdd.n130 85.8723
R2526 vdd.t179 vdd.n88 85.8723
R2527 vdd.t172 vdd.n41 85.8723
R2528 vdd.t200 vdd.n1444 85.8723
R2529 vdd.t146 vdd.n1491 85.8723
R2530 vdd.t142 vdd.n1354 85.8723
R2531 vdd.t150 vdd.n1401 85.8723
R2532 vdd.t171 vdd.n1265 85.8723
R2533 vdd.t180 vdd.n1312 85.8723
R2534 vdd.n2617 vdd.n662 78.546
R2535 vdd.n2072 vdd.n833 78.546
R2536 vdd.n254 vdd.n253 75.1835
R2537 vdd.n252 vdd.n251 75.1835
R2538 vdd.n250 vdd.n249 75.1835
R2539 vdd.n164 vdd.n163 75.1835
R2540 vdd.n162 vdd.n161 75.1835
R2541 vdd.n160 vdd.n159 75.1835
R2542 vdd.n75 vdd.n74 75.1835
R2543 vdd.n73 vdd.n72 75.1835
R2544 vdd.n71 vdd.n70 75.1835
R2545 vdd.n1474 vdd.n1473 75.1835
R2546 vdd.n1476 vdd.n1475 75.1835
R2547 vdd.n1478 vdd.n1477 75.1835
R2548 vdd.n1384 vdd.n1383 75.1835
R2549 vdd.n1386 vdd.n1385 75.1835
R2550 vdd.n1388 vdd.n1387 75.1835
R2551 vdd.n1295 vdd.n1294 75.1835
R2552 vdd.n1297 vdd.n1296 75.1835
R2553 vdd.n1299 vdd.n1298 75.1835
R2554 vdd.n2553 vdd.n2552 72.8958
R2555 vdd.n2552 vdd.n2296 72.8958
R2556 vdd.n2552 vdd.n2297 72.8958
R2557 vdd.n2552 vdd.n2298 72.8958
R2558 vdd.n2552 vdd.n2299 72.8958
R2559 vdd.n2552 vdd.n2300 72.8958
R2560 vdd.n2552 vdd.n2301 72.8958
R2561 vdd.n2552 vdd.n2302 72.8958
R2562 vdd.n2552 vdd.n2303 72.8958
R2563 vdd.n2552 vdd.n2304 72.8958
R2564 vdd.n2552 vdd.n2305 72.8958
R2565 vdd.n2552 vdd.n2306 72.8958
R2566 vdd.n2552 vdd.n2307 72.8958
R2567 vdd.n2552 vdd.n2308 72.8958
R2568 vdd.n2552 vdd.n2309 72.8958
R2569 vdd.n2552 vdd.n2310 72.8958
R2570 vdd.n2552 vdd.n2311 72.8958
R2571 vdd.n593 vdd.n484 72.8958
R2572 vdd.n2772 vdd.n484 72.8958
R2573 vdd.n587 vdd.n484 72.8958
R2574 vdd.n2779 vdd.n484 72.8958
R2575 vdd.n584 vdd.n484 72.8958
R2576 vdd.n2786 vdd.n484 72.8958
R2577 vdd.n581 vdd.n484 72.8958
R2578 vdd.n2793 vdd.n484 72.8958
R2579 vdd.n2796 vdd.n484 72.8958
R2580 vdd.n2652 vdd.n484 72.8958
R2581 vdd.n2657 vdd.n484 72.8958
R2582 vdd.n2651 vdd.n484 72.8958
R2583 vdd.n2664 vdd.n484 72.8958
R2584 vdd.n2648 vdd.n484 72.8958
R2585 vdd.n2671 vdd.n484 72.8958
R2586 vdd.n2645 vdd.n484 72.8958
R2587 vdd.n2678 vdd.n484 72.8958
R2588 vdd.n2031 vdd.n2030 72.8958
R2589 vdd.n2031 vdd.n874 72.8958
R2590 vdd.n2031 vdd.n875 72.8958
R2591 vdd.n2031 vdd.n876 72.8958
R2592 vdd.n2031 vdd.n877 72.8958
R2593 vdd.n2031 vdd.n878 72.8958
R2594 vdd.n2031 vdd.n879 72.8958
R2595 vdd.n2031 vdd.n880 72.8958
R2596 vdd.n2031 vdd.n881 72.8958
R2597 vdd.n2031 vdd.n882 72.8958
R2598 vdd.n2031 vdd.n883 72.8958
R2599 vdd.n2031 vdd.n884 72.8958
R2600 vdd.n2031 vdd.n885 72.8958
R2601 vdd.n2031 vdd.n886 72.8958
R2602 vdd.n2031 vdd.n887 72.8958
R2603 vdd.n2031 vdd.n888 72.8958
R2604 vdd.n2031 vdd.n889 72.8958
R2605 vdd.n2279 vdd.n742 72.8958
R2606 vdd.n2279 vdd.n743 72.8958
R2607 vdd.n2279 vdd.n744 72.8958
R2608 vdd.n2279 vdd.n745 72.8958
R2609 vdd.n2279 vdd.n746 72.8958
R2610 vdd.n2279 vdd.n747 72.8958
R2611 vdd.n2279 vdd.n748 72.8958
R2612 vdd.n2279 vdd.n749 72.8958
R2613 vdd.n2279 vdd.n750 72.8958
R2614 vdd.n2279 vdd.n751 72.8958
R2615 vdd.n2279 vdd.n752 72.8958
R2616 vdd.n2279 vdd.n753 72.8958
R2617 vdd.n2279 vdd.n754 72.8958
R2618 vdd.n2279 vdd.n755 72.8958
R2619 vdd.n2279 vdd.n756 72.8958
R2620 vdd.n2279 vdd.n757 72.8958
R2621 vdd.n2279 vdd.n758 72.8958
R2622 vdd.n2552 vdd.n2551 72.8958
R2623 vdd.n2552 vdd.n2280 72.8958
R2624 vdd.n2552 vdd.n2281 72.8958
R2625 vdd.n2552 vdd.n2282 72.8958
R2626 vdd.n2552 vdd.n2283 72.8958
R2627 vdd.n2552 vdd.n2284 72.8958
R2628 vdd.n2552 vdd.n2285 72.8958
R2629 vdd.n2552 vdd.n2286 72.8958
R2630 vdd.n2552 vdd.n2287 72.8958
R2631 vdd.n2552 vdd.n2288 72.8958
R2632 vdd.n2552 vdd.n2289 72.8958
R2633 vdd.n2552 vdd.n2290 72.8958
R2634 vdd.n2552 vdd.n2291 72.8958
R2635 vdd.n2552 vdd.n2292 72.8958
R2636 vdd.n2552 vdd.n2293 72.8958
R2637 vdd.n2552 vdd.n2294 72.8958
R2638 vdd.n2552 vdd.n2295 72.8958
R2639 vdd.n2702 vdd.n484 72.8958
R2640 vdd.n625 vdd.n484 72.8958
R2641 vdd.n2710 vdd.n484 72.8958
R2642 vdd.n620 vdd.n484 72.8958
R2643 vdd.n2717 vdd.n484 72.8958
R2644 vdd.n617 vdd.n484 72.8958
R2645 vdd.n2724 vdd.n484 72.8958
R2646 vdd.n614 vdd.n484 72.8958
R2647 vdd.n2731 vdd.n484 72.8958
R2648 vdd.n2735 vdd.n484 72.8958
R2649 vdd.n611 vdd.n484 72.8958
R2650 vdd.n2742 vdd.n484 72.8958
R2651 vdd.n608 vdd.n484 72.8958
R2652 vdd.n2749 vdd.n484 72.8958
R2653 vdd.n605 vdd.n484 72.8958
R2654 vdd.n2756 vdd.n484 72.8958
R2655 vdd.n2759 vdd.n484 72.8958
R2656 vdd.n2279 vdd.n740 72.8958
R2657 vdd.n2279 vdd.n739 72.8958
R2658 vdd.n2279 vdd.n738 72.8958
R2659 vdd.n2279 vdd.n737 72.8958
R2660 vdd.n2279 vdd.n736 72.8958
R2661 vdd.n2279 vdd.n735 72.8958
R2662 vdd.n2279 vdd.n734 72.8958
R2663 vdd.n2279 vdd.n733 72.8958
R2664 vdd.n2279 vdd.n732 72.8958
R2665 vdd.n2279 vdd.n731 72.8958
R2666 vdd.n2279 vdd.n730 72.8958
R2667 vdd.n2279 vdd.n729 72.8958
R2668 vdd.n2279 vdd.n728 72.8958
R2669 vdd.n2279 vdd.n727 72.8958
R2670 vdd.n2279 vdd.n726 72.8958
R2671 vdd.n2279 vdd.n725 72.8958
R2672 vdd.n2279 vdd.n724 72.8958
R2673 vdd.n2032 vdd.n2031 72.8958
R2674 vdd.n2031 vdd.n890 72.8958
R2675 vdd.n2031 vdd.n891 72.8958
R2676 vdd.n2031 vdd.n892 72.8958
R2677 vdd.n2031 vdd.n893 72.8958
R2678 vdd.n2031 vdd.n894 72.8958
R2679 vdd.n2031 vdd.n895 72.8958
R2680 vdd.n2031 vdd.n896 72.8958
R2681 vdd.n2031 vdd.n897 72.8958
R2682 vdd.n2031 vdd.n898 72.8958
R2683 vdd.n2031 vdd.n899 72.8958
R2684 vdd.n2031 vdd.n900 72.8958
R2685 vdd.n2031 vdd.n901 72.8958
R2686 vdd.n2031 vdd.n902 72.8958
R2687 vdd.n2031 vdd.n903 72.8958
R2688 vdd.n2031 vdd.n904 72.8958
R2689 vdd.n2031 vdd.n905 72.8958
R2690 vdd.n1784 vdd.n1783 66.2847
R2691 vdd.n1783 vdd.n1559 66.2847
R2692 vdd.n1783 vdd.n1560 66.2847
R2693 vdd.n1783 vdd.n1561 66.2847
R2694 vdd.n1783 vdd.n1562 66.2847
R2695 vdd.n1783 vdd.n1563 66.2847
R2696 vdd.n1783 vdd.n1564 66.2847
R2697 vdd.n1783 vdd.n1565 66.2847
R2698 vdd.n1783 vdd.n1566 66.2847
R2699 vdd.n1783 vdd.n1567 66.2847
R2700 vdd.n1783 vdd.n1568 66.2847
R2701 vdd.n1783 vdd.n1569 66.2847
R2702 vdd.n1783 vdd.n1570 66.2847
R2703 vdd.n1783 vdd.n1571 66.2847
R2704 vdd.n1783 vdd.n1572 66.2847
R2705 vdd.n1783 vdd.n1573 66.2847
R2706 vdd.n1783 vdd.n1574 66.2847
R2707 vdd.n1783 vdd.n1575 66.2847
R2708 vdd.n1783 vdd.n1576 66.2847
R2709 vdd.n1783 vdd.n1577 66.2847
R2710 vdd.n1783 vdd.n1578 66.2847
R2711 vdd.n1783 vdd.n1579 66.2847
R2712 vdd.n1783 vdd.n1580 66.2847
R2713 vdd.n1783 vdd.n1581 66.2847
R2714 vdd.n1783 vdd.n1582 66.2847
R2715 vdd.n1783 vdd.n1583 66.2847
R2716 vdd.n1783 vdd.n1584 66.2847
R2717 vdd.n1783 vdd.n1585 66.2847
R2718 vdd.n1783 vdd.n1586 66.2847
R2719 vdd.n1783 vdd.n1587 66.2847
R2720 vdd.n1783 vdd.n1588 66.2847
R2721 vdd.n1223 vdd.n873 66.2847
R2722 vdd.n1220 vdd.n873 66.2847
R2723 vdd.n1216 vdd.n873 66.2847
R2724 vdd.n1893 vdd.n873 66.2847
R2725 vdd.n1007 vdd.n873 66.2847
R2726 vdd.n1900 vdd.n873 66.2847
R2727 vdd.n1000 vdd.n873 66.2847
R2728 vdd.n1907 vdd.n873 66.2847
R2729 vdd.n993 vdd.n873 66.2847
R2730 vdd.n1914 vdd.n873 66.2847
R2731 vdd.n987 vdd.n873 66.2847
R2732 vdd.n982 vdd.n873 66.2847
R2733 vdd.n1925 vdd.n873 66.2847
R2734 vdd.n974 vdd.n873 66.2847
R2735 vdd.n1932 vdd.n873 66.2847
R2736 vdd.n967 vdd.n873 66.2847
R2737 vdd.n1939 vdd.n873 66.2847
R2738 vdd.n960 vdd.n873 66.2847
R2739 vdd.n1946 vdd.n873 66.2847
R2740 vdd.n953 vdd.n873 66.2847
R2741 vdd.n1953 vdd.n873 66.2847
R2742 vdd.n947 vdd.n873 66.2847
R2743 vdd.n942 vdd.n873 66.2847
R2744 vdd.n1964 vdd.n873 66.2847
R2745 vdd.n934 vdd.n873 66.2847
R2746 vdd.n1971 vdd.n873 66.2847
R2747 vdd.n927 vdd.n873 66.2847
R2748 vdd.n1978 vdd.n873 66.2847
R2749 vdd.n920 vdd.n873 66.2847
R2750 vdd.n1985 vdd.n873 66.2847
R2751 vdd.n1990 vdd.n873 66.2847
R2752 vdd.n916 vdd.n873 66.2847
R2753 vdd.n2933 vdd.n2932 66.2847
R2754 vdd.n2932 vdd.n485 66.2847
R2755 vdd.n2932 vdd.n486 66.2847
R2756 vdd.n2932 vdd.n487 66.2847
R2757 vdd.n2932 vdd.n488 66.2847
R2758 vdd.n2932 vdd.n489 66.2847
R2759 vdd.n2932 vdd.n490 66.2847
R2760 vdd.n2932 vdd.n491 66.2847
R2761 vdd.n2932 vdd.n492 66.2847
R2762 vdd.n2932 vdd.n493 66.2847
R2763 vdd.n2932 vdd.n494 66.2847
R2764 vdd.n2932 vdd.n495 66.2847
R2765 vdd.n2932 vdd.n496 66.2847
R2766 vdd.n2932 vdd.n497 66.2847
R2767 vdd.n2932 vdd.n498 66.2847
R2768 vdd.n2932 vdd.n499 66.2847
R2769 vdd.n2932 vdd.n500 66.2847
R2770 vdd.n2932 vdd.n501 66.2847
R2771 vdd.n2932 vdd.n502 66.2847
R2772 vdd.n2932 vdd.n503 66.2847
R2773 vdd.n2932 vdd.n504 66.2847
R2774 vdd.n2932 vdd.n505 66.2847
R2775 vdd.n2932 vdd.n506 66.2847
R2776 vdd.n2932 vdd.n507 66.2847
R2777 vdd.n2932 vdd.n508 66.2847
R2778 vdd.n2932 vdd.n509 66.2847
R2779 vdd.n2932 vdd.n510 66.2847
R2780 vdd.n2932 vdd.n511 66.2847
R2781 vdd.n2932 vdd.n512 66.2847
R2782 vdd.n2932 vdd.n513 66.2847
R2783 vdd.n2932 vdd.n514 66.2847
R2784 vdd.n2997 vdd.n329 66.2847
R2785 vdd.n3006 vdd.n329 66.2847
R2786 vdd.n439 vdd.n329 66.2847
R2787 vdd.n3013 vdd.n329 66.2847
R2788 vdd.n432 vdd.n329 66.2847
R2789 vdd.n3020 vdd.n329 66.2847
R2790 vdd.n425 vdd.n329 66.2847
R2791 vdd.n3027 vdd.n329 66.2847
R2792 vdd.n418 vdd.n329 66.2847
R2793 vdd.n3034 vdd.n329 66.2847
R2794 vdd.n412 vdd.n329 66.2847
R2795 vdd.n407 vdd.n329 66.2847
R2796 vdd.n3045 vdd.n329 66.2847
R2797 vdd.n399 vdd.n329 66.2847
R2798 vdd.n3052 vdd.n329 66.2847
R2799 vdd.n392 vdd.n329 66.2847
R2800 vdd.n3059 vdd.n329 66.2847
R2801 vdd.n385 vdd.n329 66.2847
R2802 vdd.n3066 vdd.n329 66.2847
R2803 vdd.n378 vdd.n329 66.2847
R2804 vdd.n3073 vdd.n329 66.2847
R2805 vdd.n372 vdd.n329 66.2847
R2806 vdd.n367 vdd.n329 66.2847
R2807 vdd.n3084 vdd.n329 66.2847
R2808 vdd.n359 vdd.n329 66.2847
R2809 vdd.n3091 vdd.n329 66.2847
R2810 vdd.n352 vdd.n329 66.2847
R2811 vdd.n3098 vdd.n329 66.2847
R2812 vdd.n345 vdd.n329 66.2847
R2813 vdd.n3105 vdd.n329 66.2847
R2814 vdd.n3108 vdd.n329 66.2847
R2815 vdd.n333 vdd.n329 66.2847
R2816 vdd.n334 vdd.n333 52.4337
R2817 vdd.n3108 vdd.n3107 52.4337
R2818 vdd.n3105 vdd.n3104 52.4337
R2819 vdd.n3100 vdd.n345 52.4337
R2820 vdd.n3098 vdd.n3097 52.4337
R2821 vdd.n3093 vdd.n352 52.4337
R2822 vdd.n3091 vdd.n3090 52.4337
R2823 vdd.n3086 vdd.n359 52.4337
R2824 vdd.n3084 vdd.n3083 52.4337
R2825 vdd.n368 vdd.n367 52.4337
R2826 vdd.n3075 vdd.n372 52.4337
R2827 vdd.n3073 vdd.n3072 52.4337
R2828 vdd.n3068 vdd.n378 52.4337
R2829 vdd.n3066 vdd.n3065 52.4337
R2830 vdd.n3061 vdd.n385 52.4337
R2831 vdd.n3059 vdd.n3058 52.4337
R2832 vdd.n3054 vdd.n392 52.4337
R2833 vdd.n3052 vdd.n3051 52.4337
R2834 vdd.n3047 vdd.n399 52.4337
R2835 vdd.n3045 vdd.n3044 52.4337
R2836 vdd.n408 vdd.n407 52.4337
R2837 vdd.n3036 vdd.n412 52.4337
R2838 vdd.n3034 vdd.n3033 52.4337
R2839 vdd.n3029 vdd.n418 52.4337
R2840 vdd.n3027 vdd.n3026 52.4337
R2841 vdd.n3022 vdd.n425 52.4337
R2842 vdd.n3020 vdd.n3019 52.4337
R2843 vdd.n3015 vdd.n432 52.4337
R2844 vdd.n3013 vdd.n3012 52.4337
R2845 vdd.n3008 vdd.n439 52.4337
R2846 vdd.n3006 vdd.n3005 52.4337
R2847 vdd.n2998 vdd.n2997 52.4337
R2848 vdd.n2934 vdd.n2933 52.4337
R2849 vdd.n517 vdd.n485 52.4337
R2850 vdd.n523 vdd.n486 52.4337
R2851 vdd.n2923 vdd.n487 52.4337
R2852 vdd.n2919 vdd.n488 52.4337
R2853 vdd.n2915 vdd.n489 52.4337
R2854 vdd.n2911 vdd.n490 52.4337
R2855 vdd.n2907 vdd.n491 52.4337
R2856 vdd.n2903 vdd.n492 52.4337
R2857 vdd.n2899 vdd.n493 52.4337
R2858 vdd.n2891 vdd.n494 52.4337
R2859 vdd.n2887 vdd.n495 52.4337
R2860 vdd.n2883 vdd.n496 52.4337
R2861 vdd.n2879 vdd.n497 52.4337
R2862 vdd.n2875 vdd.n498 52.4337
R2863 vdd.n2871 vdd.n499 52.4337
R2864 vdd.n2867 vdd.n500 52.4337
R2865 vdd.n2863 vdd.n501 52.4337
R2866 vdd.n2859 vdd.n502 52.4337
R2867 vdd.n2855 vdd.n503 52.4337
R2868 vdd.n2851 vdd.n504 52.4337
R2869 vdd.n2845 vdd.n505 52.4337
R2870 vdd.n2841 vdd.n506 52.4337
R2871 vdd.n2837 vdd.n507 52.4337
R2872 vdd.n2833 vdd.n508 52.4337
R2873 vdd.n2829 vdd.n509 52.4337
R2874 vdd.n2825 vdd.n510 52.4337
R2875 vdd.n2821 vdd.n511 52.4337
R2876 vdd.n2817 vdd.n512 52.4337
R2877 vdd.n2813 vdd.n513 52.4337
R2878 vdd.n2809 vdd.n514 52.4337
R2879 vdd.n1992 vdd.n916 52.4337
R2880 vdd.n1990 vdd.n1989 52.4337
R2881 vdd.n1985 vdd.n1984 52.4337
R2882 vdd.n1980 vdd.n920 52.4337
R2883 vdd.n1978 vdd.n1977 52.4337
R2884 vdd.n1973 vdd.n927 52.4337
R2885 vdd.n1971 vdd.n1970 52.4337
R2886 vdd.n1966 vdd.n934 52.4337
R2887 vdd.n1964 vdd.n1963 52.4337
R2888 vdd.n943 vdd.n942 52.4337
R2889 vdd.n1955 vdd.n947 52.4337
R2890 vdd.n1953 vdd.n1952 52.4337
R2891 vdd.n1948 vdd.n953 52.4337
R2892 vdd.n1946 vdd.n1945 52.4337
R2893 vdd.n1941 vdd.n960 52.4337
R2894 vdd.n1939 vdd.n1938 52.4337
R2895 vdd.n1934 vdd.n967 52.4337
R2896 vdd.n1932 vdd.n1931 52.4337
R2897 vdd.n1927 vdd.n974 52.4337
R2898 vdd.n1925 vdd.n1924 52.4337
R2899 vdd.n983 vdd.n982 52.4337
R2900 vdd.n1916 vdd.n987 52.4337
R2901 vdd.n1914 vdd.n1913 52.4337
R2902 vdd.n1909 vdd.n993 52.4337
R2903 vdd.n1907 vdd.n1906 52.4337
R2904 vdd.n1902 vdd.n1000 52.4337
R2905 vdd.n1900 vdd.n1899 52.4337
R2906 vdd.n1895 vdd.n1007 52.4337
R2907 vdd.n1893 vdd.n1892 52.4337
R2908 vdd.n1217 vdd.n1216 52.4337
R2909 vdd.n1221 vdd.n1220 52.4337
R2910 vdd.n1881 vdd.n1223 52.4337
R2911 vdd.n1785 vdd.n1784 52.4337
R2912 vdd.n1591 vdd.n1559 52.4337
R2913 vdd.n1595 vdd.n1560 52.4337
R2914 vdd.n1597 vdd.n1561 52.4337
R2915 vdd.n1601 vdd.n1562 52.4337
R2916 vdd.n1603 vdd.n1563 52.4337
R2917 vdd.n1607 vdd.n1564 52.4337
R2918 vdd.n1609 vdd.n1565 52.4337
R2919 vdd.n1613 vdd.n1566 52.4337
R2920 vdd.n1615 vdd.n1567 52.4337
R2921 vdd.n1621 vdd.n1568 52.4337
R2922 vdd.n1623 vdd.n1569 52.4337
R2923 vdd.n1627 vdd.n1570 52.4337
R2924 vdd.n1629 vdd.n1571 52.4337
R2925 vdd.n1633 vdd.n1572 52.4337
R2926 vdd.n1635 vdd.n1573 52.4337
R2927 vdd.n1639 vdd.n1574 52.4337
R2928 vdd.n1641 vdd.n1575 52.4337
R2929 vdd.n1645 vdd.n1576 52.4337
R2930 vdd.n1647 vdd.n1577 52.4337
R2931 vdd.n1719 vdd.n1578 52.4337
R2932 vdd.n1652 vdd.n1579 52.4337
R2933 vdd.n1656 vdd.n1580 52.4337
R2934 vdd.n1658 vdd.n1581 52.4337
R2935 vdd.n1662 vdd.n1582 52.4337
R2936 vdd.n1664 vdd.n1583 52.4337
R2937 vdd.n1668 vdd.n1584 52.4337
R2938 vdd.n1670 vdd.n1585 52.4337
R2939 vdd.n1674 vdd.n1586 52.4337
R2940 vdd.n1676 vdd.n1587 52.4337
R2941 vdd.n1680 vdd.n1588 52.4337
R2942 vdd.n1784 vdd.n1558 52.4337
R2943 vdd.n1594 vdd.n1559 52.4337
R2944 vdd.n1596 vdd.n1560 52.4337
R2945 vdd.n1600 vdd.n1561 52.4337
R2946 vdd.n1602 vdd.n1562 52.4337
R2947 vdd.n1606 vdd.n1563 52.4337
R2948 vdd.n1608 vdd.n1564 52.4337
R2949 vdd.n1612 vdd.n1565 52.4337
R2950 vdd.n1614 vdd.n1566 52.4337
R2951 vdd.n1620 vdd.n1567 52.4337
R2952 vdd.n1622 vdd.n1568 52.4337
R2953 vdd.n1626 vdd.n1569 52.4337
R2954 vdd.n1628 vdd.n1570 52.4337
R2955 vdd.n1632 vdd.n1571 52.4337
R2956 vdd.n1634 vdd.n1572 52.4337
R2957 vdd.n1638 vdd.n1573 52.4337
R2958 vdd.n1640 vdd.n1574 52.4337
R2959 vdd.n1644 vdd.n1575 52.4337
R2960 vdd.n1646 vdd.n1576 52.4337
R2961 vdd.n1650 vdd.n1577 52.4337
R2962 vdd.n1651 vdd.n1578 52.4337
R2963 vdd.n1655 vdd.n1579 52.4337
R2964 vdd.n1657 vdd.n1580 52.4337
R2965 vdd.n1661 vdd.n1581 52.4337
R2966 vdd.n1663 vdd.n1582 52.4337
R2967 vdd.n1667 vdd.n1583 52.4337
R2968 vdd.n1669 vdd.n1584 52.4337
R2969 vdd.n1673 vdd.n1585 52.4337
R2970 vdd.n1675 vdd.n1586 52.4337
R2971 vdd.n1679 vdd.n1587 52.4337
R2972 vdd.n1681 vdd.n1588 52.4337
R2973 vdd.n1223 vdd.n1222 52.4337
R2974 vdd.n1220 vdd.n1219 52.4337
R2975 vdd.n1216 vdd.n1008 52.4337
R2976 vdd.n1894 vdd.n1893 52.4337
R2977 vdd.n1007 vdd.n1001 52.4337
R2978 vdd.n1901 vdd.n1900 52.4337
R2979 vdd.n1000 vdd.n994 52.4337
R2980 vdd.n1908 vdd.n1907 52.4337
R2981 vdd.n993 vdd.n988 52.4337
R2982 vdd.n1915 vdd.n1914 52.4337
R2983 vdd.n987 vdd.n986 52.4337
R2984 vdd.n982 vdd.n975 52.4337
R2985 vdd.n1926 vdd.n1925 52.4337
R2986 vdd.n974 vdd.n968 52.4337
R2987 vdd.n1933 vdd.n1932 52.4337
R2988 vdd.n967 vdd.n961 52.4337
R2989 vdd.n1940 vdd.n1939 52.4337
R2990 vdd.n960 vdd.n954 52.4337
R2991 vdd.n1947 vdd.n1946 52.4337
R2992 vdd.n953 vdd.n948 52.4337
R2993 vdd.n1954 vdd.n1953 52.4337
R2994 vdd.n947 vdd.n946 52.4337
R2995 vdd.n942 vdd.n935 52.4337
R2996 vdd.n1965 vdd.n1964 52.4337
R2997 vdd.n934 vdd.n928 52.4337
R2998 vdd.n1972 vdd.n1971 52.4337
R2999 vdd.n927 vdd.n921 52.4337
R3000 vdd.n1979 vdd.n1978 52.4337
R3001 vdd.n920 vdd.n917 52.4337
R3002 vdd.n1986 vdd.n1985 52.4337
R3003 vdd.n1991 vdd.n1990 52.4337
R3004 vdd.n1227 vdd.n916 52.4337
R3005 vdd.n2933 vdd.n483 52.4337
R3006 vdd.n522 vdd.n485 52.4337
R3007 vdd.n2924 vdd.n486 52.4337
R3008 vdd.n2920 vdd.n487 52.4337
R3009 vdd.n2916 vdd.n488 52.4337
R3010 vdd.n2912 vdd.n489 52.4337
R3011 vdd.n2908 vdd.n490 52.4337
R3012 vdd.n2904 vdd.n491 52.4337
R3013 vdd.n2900 vdd.n492 52.4337
R3014 vdd.n2890 vdd.n493 52.4337
R3015 vdd.n2888 vdd.n494 52.4337
R3016 vdd.n2884 vdd.n495 52.4337
R3017 vdd.n2880 vdd.n496 52.4337
R3018 vdd.n2876 vdd.n497 52.4337
R3019 vdd.n2872 vdd.n498 52.4337
R3020 vdd.n2868 vdd.n499 52.4337
R3021 vdd.n2864 vdd.n500 52.4337
R3022 vdd.n2860 vdd.n501 52.4337
R3023 vdd.n2856 vdd.n502 52.4337
R3024 vdd.n2852 vdd.n503 52.4337
R3025 vdd.n2844 vdd.n504 52.4337
R3026 vdd.n2842 vdd.n505 52.4337
R3027 vdd.n2838 vdd.n506 52.4337
R3028 vdd.n2834 vdd.n507 52.4337
R3029 vdd.n2830 vdd.n508 52.4337
R3030 vdd.n2826 vdd.n509 52.4337
R3031 vdd.n2822 vdd.n510 52.4337
R3032 vdd.n2818 vdd.n511 52.4337
R3033 vdd.n2814 vdd.n512 52.4337
R3034 vdd.n2810 vdd.n513 52.4337
R3035 vdd.n2806 vdd.n514 52.4337
R3036 vdd.n2997 vdd.n440 52.4337
R3037 vdd.n3007 vdd.n3006 52.4337
R3038 vdd.n439 vdd.n433 52.4337
R3039 vdd.n3014 vdd.n3013 52.4337
R3040 vdd.n432 vdd.n426 52.4337
R3041 vdd.n3021 vdd.n3020 52.4337
R3042 vdd.n425 vdd.n419 52.4337
R3043 vdd.n3028 vdd.n3027 52.4337
R3044 vdd.n418 vdd.n413 52.4337
R3045 vdd.n3035 vdd.n3034 52.4337
R3046 vdd.n412 vdd.n411 52.4337
R3047 vdd.n407 vdd.n400 52.4337
R3048 vdd.n3046 vdd.n3045 52.4337
R3049 vdd.n399 vdd.n393 52.4337
R3050 vdd.n3053 vdd.n3052 52.4337
R3051 vdd.n392 vdd.n386 52.4337
R3052 vdd.n3060 vdd.n3059 52.4337
R3053 vdd.n385 vdd.n379 52.4337
R3054 vdd.n3067 vdd.n3066 52.4337
R3055 vdd.n378 vdd.n373 52.4337
R3056 vdd.n3074 vdd.n3073 52.4337
R3057 vdd.n372 vdd.n371 52.4337
R3058 vdd.n367 vdd.n360 52.4337
R3059 vdd.n3085 vdd.n3084 52.4337
R3060 vdd.n359 vdd.n353 52.4337
R3061 vdd.n3092 vdd.n3091 52.4337
R3062 vdd.n352 vdd.n346 52.4337
R3063 vdd.n3099 vdd.n3098 52.4337
R3064 vdd.n345 vdd.n338 52.4337
R3065 vdd.n3106 vdd.n3105 52.4337
R3066 vdd.n3109 vdd.n3108 52.4337
R3067 vdd.n333 vdd.n330 52.4337
R3068 vdd.t107 vdd.t118 51.4683
R3069 vdd.n250 vdd.n248 42.0461
R3070 vdd.n160 vdd.n158 42.0461
R3071 vdd.n71 vdd.n69 42.0461
R3072 vdd.n1474 vdd.n1472 42.0461
R3073 vdd.n1384 vdd.n1382 42.0461
R3074 vdd.n1295 vdd.n1293 42.0461
R3075 vdd.n296 vdd.n295 41.6884
R3076 vdd.n206 vdd.n205 41.6884
R3077 vdd.n117 vdd.n116 41.6884
R3078 vdd.n1520 vdd.n1519 41.6884
R3079 vdd.n1430 vdd.n1429 41.6884
R3080 vdd.n1341 vdd.n1340 41.6884
R3081 vdd.n1684 vdd.n1683 41.1157
R3082 vdd.n1722 vdd.n1721 41.1157
R3083 vdd.n1618 vdd.n1617 41.1157
R3084 vdd.n3002 vdd.n3001 41.1157
R3085 vdd.n3041 vdd.n406 41.1157
R3086 vdd.n3080 vdd.n366 41.1157
R3087 vdd.n2759 vdd.n2758 39.2114
R3088 vdd.n2756 vdd.n2755 39.2114
R3089 vdd.n2751 vdd.n605 39.2114
R3090 vdd.n2749 vdd.n2748 39.2114
R3091 vdd.n2744 vdd.n608 39.2114
R3092 vdd.n2742 vdd.n2741 39.2114
R3093 vdd.n2737 vdd.n611 39.2114
R3094 vdd.n2735 vdd.n2734 39.2114
R3095 vdd.n2731 vdd.n2730 39.2114
R3096 vdd.n2726 vdd.n614 39.2114
R3097 vdd.n2724 vdd.n2723 39.2114
R3098 vdd.n2719 vdd.n617 39.2114
R3099 vdd.n2717 vdd.n2716 39.2114
R3100 vdd.n2712 vdd.n620 39.2114
R3101 vdd.n2710 vdd.n2709 39.2114
R3102 vdd.n2704 vdd.n625 39.2114
R3103 vdd.n2702 vdd.n2701 39.2114
R3104 vdd.n2551 vdd.n2550 39.2114
R3105 vdd.n2545 vdd.n2280 39.2114
R3106 vdd.n2542 vdd.n2281 39.2114
R3107 vdd.n2538 vdd.n2282 39.2114
R3108 vdd.n2534 vdd.n2283 39.2114
R3109 vdd.n2530 vdd.n2284 39.2114
R3110 vdd.n2526 vdd.n2285 39.2114
R3111 vdd.n2522 vdd.n2286 39.2114
R3112 vdd.n2518 vdd.n2287 39.2114
R3113 vdd.n2514 vdd.n2288 39.2114
R3114 vdd.n2510 vdd.n2289 39.2114
R3115 vdd.n2506 vdd.n2290 39.2114
R3116 vdd.n2502 vdd.n2291 39.2114
R3117 vdd.n2498 vdd.n2292 39.2114
R3118 vdd.n2494 vdd.n2293 39.2114
R3119 vdd.n2490 vdd.n2294 39.2114
R3120 vdd.n2485 vdd.n2295 39.2114
R3121 vdd.n2274 vdd.n758 39.2114
R3122 vdd.n2270 vdd.n757 39.2114
R3123 vdd.n2266 vdd.n756 39.2114
R3124 vdd.n2262 vdd.n755 39.2114
R3125 vdd.n2258 vdd.n754 39.2114
R3126 vdd.n2254 vdd.n753 39.2114
R3127 vdd.n2250 vdd.n752 39.2114
R3128 vdd.n2246 vdd.n751 39.2114
R3129 vdd.n2242 vdd.n750 39.2114
R3130 vdd.n2238 vdd.n749 39.2114
R3131 vdd.n2234 vdd.n748 39.2114
R3132 vdd.n2230 vdd.n747 39.2114
R3133 vdd.n2226 vdd.n746 39.2114
R3134 vdd.n2222 vdd.n745 39.2114
R3135 vdd.n2218 vdd.n744 39.2114
R3136 vdd.n2213 vdd.n743 39.2114
R3137 vdd.n2209 vdd.n742 39.2114
R3138 vdd.n2030 vdd.n2029 39.2114
R3139 vdd.n2024 vdd.n874 39.2114
R3140 vdd.n2021 vdd.n875 39.2114
R3141 vdd.n2017 vdd.n876 39.2114
R3142 vdd.n2013 vdd.n877 39.2114
R3143 vdd.n2009 vdd.n878 39.2114
R3144 vdd.n2005 vdd.n879 39.2114
R3145 vdd.n2001 vdd.n880 39.2114
R3146 vdd.n1997 vdd.n881 39.2114
R3147 vdd.n1066 vdd.n882 39.2114
R3148 vdd.n1070 vdd.n883 39.2114
R3149 vdd.n1074 vdd.n884 39.2114
R3150 vdd.n1078 vdd.n885 39.2114
R3151 vdd.n1082 vdd.n886 39.2114
R3152 vdd.n1086 vdd.n887 39.2114
R3153 vdd.n1090 vdd.n888 39.2114
R3154 vdd.n1095 vdd.n889 39.2114
R3155 vdd.n2678 vdd.n2677 39.2114
R3156 vdd.n2673 vdd.n2645 39.2114
R3157 vdd.n2671 vdd.n2670 39.2114
R3158 vdd.n2666 vdd.n2648 39.2114
R3159 vdd.n2664 vdd.n2663 39.2114
R3160 vdd.n2659 vdd.n2651 39.2114
R3161 vdd.n2657 vdd.n2656 39.2114
R3162 vdd.n2652 vdd.n577 39.2114
R3163 vdd.n2796 vdd.n2795 39.2114
R3164 vdd.n2793 vdd.n2792 39.2114
R3165 vdd.n2788 vdd.n581 39.2114
R3166 vdd.n2786 vdd.n2785 39.2114
R3167 vdd.n2781 vdd.n584 39.2114
R3168 vdd.n2779 vdd.n2778 39.2114
R3169 vdd.n2774 vdd.n587 39.2114
R3170 vdd.n2772 vdd.n2771 39.2114
R3171 vdd.n2767 vdd.n593 39.2114
R3172 vdd.n2554 vdd.n2553 39.2114
R3173 vdd.n2321 vdd.n2296 39.2114
R3174 vdd.n2325 vdd.n2297 39.2114
R3175 vdd.n2329 vdd.n2298 39.2114
R3176 vdd.n2333 vdd.n2299 39.2114
R3177 vdd.n2337 vdd.n2300 39.2114
R3178 vdd.n2341 vdd.n2301 39.2114
R3179 vdd.n2345 vdd.n2302 39.2114
R3180 vdd.n2349 vdd.n2303 39.2114
R3181 vdd.n2353 vdd.n2304 39.2114
R3182 vdd.n2357 vdd.n2305 39.2114
R3183 vdd.n2361 vdd.n2306 39.2114
R3184 vdd.n2365 vdd.n2307 39.2114
R3185 vdd.n2369 vdd.n2308 39.2114
R3186 vdd.n2373 vdd.n2309 39.2114
R3187 vdd.n2377 vdd.n2310 39.2114
R3188 vdd.n2381 vdd.n2311 39.2114
R3189 vdd.n2553 vdd.n723 39.2114
R3190 vdd.n2324 vdd.n2296 39.2114
R3191 vdd.n2328 vdd.n2297 39.2114
R3192 vdd.n2332 vdd.n2298 39.2114
R3193 vdd.n2336 vdd.n2299 39.2114
R3194 vdd.n2340 vdd.n2300 39.2114
R3195 vdd.n2344 vdd.n2301 39.2114
R3196 vdd.n2348 vdd.n2302 39.2114
R3197 vdd.n2352 vdd.n2303 39.2114
R3198 vdd.n2356 vdd.n2304 39.2114
R3199 vdd.n2360 vdd.n2305 39.2114
R3200 vdd.n2364 vdd.n2306 39.2114
R3201 vdd.n2368 vdd.n2307 39.2114
R3202 vdd.n2372 vdd.n2308 39.2114
R3203 vdd.n2376 vdd.n2309 39.2114
R3204 vdd.n2380 vdd.n2310 39.2114
R3205 vdd.n2383 vdd.n2311 39.2114
R3206 vdd.n593 vdd.n588 39.2114
R3207 vdd.n2773 vdd.n2772 39.2114
R3208 vdd.n587 vdd.n585 39.2114
R3209 vdd.n2780 vdd.n2779 39.2114
R3210 vdd.n584 vdd.n582 39.2114
R3211 vdd.n2787 vdd.n2786 39.2114
R3212 vdd.n581 vdd.n579 39.2114
R3213 vdd.n2794 vdd.n2793 39.2114
R3214 vdd.n2797 vdd.n2796 39.2114
R3215 vdd.n2653 vdd.n2652 39.2114
R3216 vdd.n2658 vdd.n2657 39.2114
R3217 vdd.n2651 vdd.n2649 39.2114
R3218 vdd.n2665 vdd.n2664 39.2114
R3219 vdd.n2648 vdd.n2646 39.2114
R3220 vdd.n2672 vdd.n2671 39.2114
R3221 vdd.n2645 vdd.n2643 39.2114
R3222 vdd.n2679 vdd.n2678 39.2114
R3223 vdd.n2030 vdd.n908 39.2114
R3224 vdd.n2022 vdd.n874 39.2114
R3225 vdd.n2018 vdd.n875 39.2114
R3226 vdd.n2014 vdd.n876 39.2114
R3227 vdd.n2010 vdd.n877 39.2114
R3228 vdd.n2006 vdd.n878 39.2114
R3229 vdd.n2002 vdd.n879 39.2114
R3230 vdd.n1998 vdd.n880 39.2114
R3231 vdd.n1065 vdd.n881 39.2114
R3232 vdd.n1069 vdd.n882 39.2114
R3233 vdd.n1073 vdd.n883 39.2114
R3234 vdd.n1077 vdd.n884 39.2114
R3235 vdd.n1081 vdd.n885 39.2114
R3236 vdd.n1085 vdd.n886 39.2114
R3237 vdd.n1089 vdd.n887 39.2114
R3238 vdd.n1094 vdd.n888 39.2114
R3239 vdd.n1098 vdd.n889 39.2114
R3240 vdd.n2212 vdd.n742 39.2114
R3241 vdd.n2217 vdd.n743 39.2114
R3242 vdd.n2221 vdd.n744 39.2114
R3243 vdd.n2225 vdd.n745 39.2114
R3244 vdd.n2229 vdd.n746 39.2114
R3245 vdd.n2233 vdd.n747 39.2114
R3246 vdd.n2237 vdd.n748 39.2114
R3247 vdd.n2241 vdd.n749 39.2114
R3248 vdd.n2245 vdd.n750 39.2114
R3249 vdd.n2249 vdd.n751 39.2114
R3250 vdd.n2253 vdd.n752 39.2114
R3251 vdd.n2257 vdd.n753 39.2114
R3252 vdd.n2261 vdd.n754 39.2114
R3253 vdd.n2265 vdd.n755 39.2114
R3254 vdd.n2269 vdd.n756 39.2114
R3255 vdd.n2273 vdd.n757 39.2114
R3256 vdd.n760 vdd.n758 39.2114
R3257 vdd.n2551 vdd.n2314 39.2114
R3258 vdd.n2543 vdd.n2280 39.2114
R3259 vdd.n2539 vdd.n2281 39.2114
R3260 vdd.n2535 vdd.n2282 39.2114
R3261 vdd.n2531 vdd.n2283 39.2114
R3262 vdd.n2527 vdd.n2284 39.2114
R3263 vdd.n2523 vdd.n2285 39.2114
R3264 vdd.n2519 vdd.n2286 39.2114
R3265 vdd.n2515 vdd.n2287 39.2114
R3266 vdd.n2511 vdd.n2288 39.2114
R3267 vdd.n2507 vdd.n2289 39.2114
R3268 vdd.n2503 vdd.n2290 39.2114
R3269 vdd.n2499 vdd.n2291 39.2114
R3270 vdd.n2495 vdd.n2292 39.2114
R3271 vdd.n2491 vdd.n2293 39.2114
R3272 vdd.n2486 vdd.n2294 39.2114
R3273 vdd.n2482 vdd.n2295 39.2114
R3274 vdd.n2703 vdd.n2702 39.2114
R3275 vdd.n625 vdd.n621 39.2114
R3276 vdd.n2711 vdd.n2710 39.2114
R3277 vdd.n620 vdd.n618 39.2114
R3278 vdd.n2718 vdd.n2717 39.2114
R3279 vdd.n617 vdd.n615 39.2114
R3280 vdd.n2725 vdd.n2724 39.2114
R3281 vdd.n614 vdd.n612 39.2114
R3282 vdd.n2732 vdd.n2731 39.2114
R3283 vdd.n2736 vdd.n2735 39.2114
R3284 vdd.n611 vdd.n609 39.2114
R3285 vdd.n2743 vdd.n2742 39.2114
R3286 vdd.n608 vdd.n606 39.2114
R3287 vdd.n2750 vdd.n2749 39.2114
R3288 vdd.n605 vdd.n603 39.2114
R3289 vdd.n2757 vdd.n2756 39.2114
R3290 vdd.n2760 vdd.n2759 39.2114
R3291 vdd.n769 vdd.n724 39.2114
R3292 vdd.n2201 vdd.n725 39.2114
R3293 vdd.n2197 vdd.n726 39.2114
R3294 vdd.n2193 vdd.n727 39.2114
R3295 vdd.n2189 vdd.n728 39.2114
R3296 vdd.n2185 vdd.n729 39.2114
R3297 vdd.n2181 vdd.n730 39.2114
R3298 vdd.n2177 vdd.n731 39.2114
R3299 vdd.n2173 vdd.n732 39.2114
R3300 vdd.n2169 vdd.n733 39.2114
R3301 vdd.n2165 vdd.n734 39.2114
R3302 vdd.n2161 vdd.n735 39.2114
R3303 vdd.n2157 vdd.n736 39.2114
R3304 vdd.n2153 vdd.n737 39.2114
R3305 vdd.n2149 vdd.n738 39.2114
R3306 vdd.n2145 vdd.n739 39.2114
R3307 vdd.n2141 vdd.n740 39.2114
R3308 vdd.n2033 vdd.n2032 39.2114
R3309 vdd.n1012 vdd.n890 39.2114
R3310 vdd.n1016 vdd.n891 39.2114
R3311 vdd.n1020 vdd.n892 39.2114
R3312 vdd.n1024 vdd.n893 39.2114
R3313 vdd.n1028 vdd.n894 39.2114
R3314 vdd.n1032 vdd.n895 39.2114
R3315 vdd.n1036 vdd.n896 39.2114
R3316 vdd.n1040 vdd.n897 39.2114
R3317 vdd.n1210 vdd.n898 39.2114
R3318 vdd.n1207 vdd.n899 39.2114
R3319 vdd.n1203 vdd.n900 39.2114
R3320 vdd.n1199 vdd.n901 39.2114
R3321 vdd.n1195 vdd.n902 39.2114
R3322 vdd.n1191 vdd.n903 39.2114
R3323 vdd.n1187 vdd.n904 39.2114
R3324 vdd.n1183 vdd.n905 39.2114
R3325 vdd.n2138 vdd.n740 39.2114
R3326 vdd.n2142 vdd.n739 39.2114
R3327 vdd.n2146 vdd.n738 39.2114
R3328 vdd.n2150 vdd.n737 39.2114
R3329 vdd.n2154 vdd.n736 39.2114
R3330 vdd.n2158 vdd.n735 39.2114
R3331 vdd.n2162 vdd.n734 39.2114
R3332 vdd.n2166 vdd.n733 39.2114
R3333 vdd.n2170 vdd.n732 39.2114
R3334 vdd.n2174 vdd.n731 39.2114
R3335 vdd.n2178 vdd.n730 39.2114
R3336 vdd.n2182 vdd.n729 39.2114
R3337 vdd.n2186 vdd.n728 39.2114
R3338 vdd.n2190 vdd.n727 39.2114
R3339 vdd.n2194 vdd.n726 39.2114
R3340 vdd.n2198 vdd.n725 39.2114
R3341 vdd.n2202 vdd.n724 39.2114
R3342 vdd.n2032 vdd.n872 39.2114
R3343 vdd.n1015 vdd.n890 39.2114
R3344 vdd.n1019 vdd.n891 39.2114
R3345 vdd.n1023 vdd.n892 39.2114
R3346 vdd.n1027 vdd.n893 39.2114
R3347 vdd.n1031 vdd.n894 39.2114
R3348 vdd.n1035 vdd.n895 39.2114
R3349 vdd.n1039 vdd.n896 39.2114
R3350 vdd.n1042 vdd.n897 39.2114
R3351 vdd.n1208 vdd.n898 39.2114
R3352 vdd.n1204 vdd.n899 39.2114
R3353 vdd.n1200 vdd.n900 39.2114
R3354 vdd.n1196 vdd.n901 39.2114
R3355 vdd.n1192 vdd.n902 39.2114
R3356 vdd.n1188 vdd.n903 39.2114
R3357 vdd.n1184 vdd.n904 39.2114
R3358 vdd.n1180 vdd.n905 39.2114
R3359 vdd.n1885 vdd.n1884 37.2369
R3360 vdd.n1921 vdd.n981 37.2369
R3361 vdd.n1960 vdd.n941 37.2369
R3362 vdd.n2850 vdd.n558 37.2369
R3363 vdd.n2898 vdd.n2897 37.2369
R3364 vdd.n2805 vdd.n2804 37.2369
R3365 vdd.n2028 vdd.n864 31.0639
R3366 vdd.n2277 vdd.n761 31.0639
R3367 vdd.n2210 vdd.n764 31.0639
R3368 vdd.n1100 vdd.n1097 31.0639
R3369 vdd.n2483 vdd.n2480 31.0639
R3370 vdd.n2700 vdd.n2699 31.0639
R3371 vdd.n2549 vdd.n716 31.0639
R3372 vdd.n2763 vdd.n2762 31.0639
R3373 vdd.n2682 vdd.n2681 31.0639
R3374 vdd.n2768 vdd.n592 31.0639
R3375 vdd.n2387 vdd.n2385 31.0639
R3376 vdd.n2556 vdd.n2555 31.0639
R3377 vdd.n2035 vdd.n2034 31.0639
R3378 vdd.n2205 vdd.n2204 31.0639
R3379 vdd.n2137 vdd.n2136 31.0639
R3380 vdd.n1179 vdd.n1178 31.0639
R3381 vdd.n1045 vdd.n1044 30.449
R3382 vdd.n773 vdd.n772 30.449
R3383 vdd.n1092 vdd.n1064 30.449
R3384 vdd.n2215 vdd.n763 30.449
R3385 vdd.n2320 vdd.n2319 30.449
R3386 vdd.n2706 vdd.n623 30.449
R3387 vdd.n2488 vdd.n2316 30.449
R3388 vdd.n591 vdd.n590 30.449
R3389 vdd.n1783 vdd.n1590 22.6735
R3390 vdd.n1879 vdd.n873 22.6735
R3391 vdd.n2932 vdd.n516 22.6735
R3392 vdd.n3117 vdd.n329 22.6735
R3393 vdd.n1794 vdd.n1552 19.3944
R3394 vdd.n1794 vdd.n1550 19.3944
R3395 vdd.n1798 vdd.n1550 19.3944
R3396 vdd.n1798 vdd.n1540 19.3944
R3397 vdd.n1811 vdd.n1540 19.3944
R3398 vdd.n1811 vdd.n1538 19.3944
R3399 vdd.n1815 vdd.n1538 19.3944
R3400 vdd.n1815 vdd.n1530 19.3944
R3401 vdd.n1829 vdd.n1530 19.3944
R3402 vdd.n1829 vdd.n1528 19.3944
R3403 vdd.n1833 vdd.n1528 19.3944
R3404 vdd.n1833 vdd.n1247 19.3944
R3405 vdd.n1845 vdd.n1247 19.3944
R3406 vdd.n1845 vdd.n1245 19.3944
R3407 vdd.n1849 vdd.n1245 19.3944
R3408 vdd.n1849 vdd.n1237 19.3944
R3409 vdd.n1862 vdd.n1237 19.3944
R3410 vdd.n1862 vdd.n1234 19.3944
R3411 vdd.n1868 vdd.n1234 19.3944
R3412 vdd.n1868 vdd.n1235 19.3944
R3413 vdd.n1235 vdd.n1225 19.3944
R3414 vdd.n1718 vdd.n1653 19.3944
R3415 vdd.n1714 vdd.n1653 19.3944
R3416 vdd.n1714 vdd.n1713 19.3944
R3417 vdd.n1713 vdd.n1712 19.3944
R3418 vdd.n1712 vdd.n1659 19.3944
R3419 vdd.n1708 vdd.n1659 19.3944
R3420 vdd.n1708 vdd.n1707 19.3944
R3421 vdd.n1707 vdd.n1706 19.3944
R3422 vdd.n1706 vdd.n1665 19.3944
R3423 vdd.n1702 vdd.n1665 19.3944
R3424 vdd.n1702 vdd.n1701 19.3944
R3425 vdd.n1701 vdd.n1700 19.3944
R3426 vdd.n1700 vdd.n1671 19.3944
R3427 vdd.n1696 vdd.n1671 19.3944
R3428 vdd.n1696 vdd.n1695 19.3944
R3429 vdd.n1695 vdd.n1694 19.3944
R3430 vdd.n1694 vdd.n1677 19.3944
R3431 vdd.n1690 vdd.n1677 19.3944
R3432 vdd.n1690 vdd.n1689 19.3944
R3433 vdd.n1689 vdd.n1688 19.3944
R3434 vdd.n1753 vdd.n1752 19.3944
R3435 vdd.n1752 vdd.n1751 19.3944
R3436 vdd.n1751 vdd.n1624 19.3944
R3437 vdd.n1747 vdd.n1624 19.3944
R3438 vdd.n1747 vdd.n1746 19.3944
R3439 vdd.n1746 vdd.n1745 19.3944
R3440 vdd.n1745 vdd.n1630 19.3944
R3441 vdd.n1741 vdd.n1630 19.3944
R3442 vdd.n1741 vdd.n1740 19.3944
R3443 vdd.n1740 vdd.n1739 19.3944
R3444 vdd.n1739 vdd.n1636 19.3944
R3445 vdd.n1735 vdd.n1636 19.3944
R3446 vdd.n1735 vdd.n1734 19.3944
R3447 vdd.n1734 vdd.n1733 19.3944
R3448 vdd.n1733 vdd.n1642 19.3944
R3449 vdd.n1729 vdd.n1642 19.3944
R3450 vdd.n1729 vdd.n1728 19.3944
R3451 vdd.n1728 vdd.n1727 19.3944
R3452 vdd.n1727 vdd.n1648 19.3944
R3453 vdd.n1723 vdd.n1648 19.3944
R3454 vdd.n1786 vdd.n1557 19.3944
R3455 vdd.n1781 vdd.n1557 19.3944
R3456 vdd.n1781 vdd.n1592 19.3944
R3457 vdd.n1777 vdd.n1592 19.3944
R3458 vdd.n1777 vdd.n1776 19.3944
R3459 vdd.n1776 vdd.n1775 19.3944
R3460 vdd.n1775 vdd.n1598 19.3944
R3461 vdd.n1771 vdd.n1598 19.3944
R3462 vdd.n1771 vdd.n1770 19.3944
R3463 vdd.n1770 vdd.n1769 19.3944
R3464 vdd.n1769 vdd.n1604 19.3944
R3465 vdd.n1765 vdd.n1604 19.3944
R3466 vdd.n1765 vdd.n1764 19.3944
R3467 vdd.n1764 vdd.n1763 19.3944
R3468 vdd.n1763 vdd.n1610 19.3944
R3469 vdd.n1759 vdd.n1610 19.3944
R3470 vdd.n1759 vdd.n1758 19.3944
R3471 vdd.n1758 vdd.n1757 19.3944
R3472 vdd.n1917 vdd.n979 19.3944
R3473 vdd.n1917 vdd.n985 19.3944
R3474 vdd.n1912 vdd.n985 19.3944
R3475 vdd.n1912 vdd.n1911 19.3944
R3476 vdd.n1911 vdd.n1910 19.3944
R3477 vdd.n1910 vdd.n992 19.3944
R3478 vdd.n1905 vdd.n992 19.3944
R3479 vdd.n1905 vdd.n1904 19.3944
R3480 vdd.n1904 vdd.n1903 19.3944
R3481 vdd.n1903 vdd.n999 19.3944
R3482 vdd.n1898 vdd.n999 19.3944
R3483 vdd.n1898 vdd.n1897 19.3944
R3484 vdd.n1897 vdd.n1896 19.3944
R3485 vdd.n1896 vdd.n1006 19.3944
R3486 vdd.n1891 vdd.n1006 19.3944
R3487 vdd.n1891 vdd.n1890 19.3944
R3488 vdd.n1218 vdd.n1011 19.3944
R3489 vdd.n1886 vdd.n1215 19.3944
R3490 vdd.n1956 vdd.n939 19.3944
R3491 vdd.n1956 vdd.n945 19.3944
R3492 vdd.n1951 vdd.n945 19.3944
R3493 vdd.n1951 vdd.n1950 19.3944
R3494 vdd.n1950 vdd.n1949 19.3944
R3495 vdd.n1949 vdd.n952 19.3944
R3496 vdd.n1944 vdd.n952 19.3944
R3497 vdd.n1944 vdd.n1943 19.3944
R3498 vdd.n1943 vdd.n1942 19.3944
R3499 vdd.n1942 vdd.n959 19.3944
R3500 vdd.n1937 vdd.n959 19.3944
R3501 vdd.n1937 vdd.n1936 19.3944
R3502 vdd.n1936 vdd.n1935 19.3944
R3503 vdd.n1935 vdd.n966 19.3944
R3504 vdd.n1930 vdd.n966 19.3944
R3505 vdd.n1930 vdd.n1929 19.3944
R3506 vdd.n1929 vdd.n1928 19.3944
R3507 vdd.n1928 vdd.n973 19.3944
R3508 vdd.n1923 vdd.n973 19.3944
R3509 vdd.n1923 vdd.n1922 19.3944
R3510 vdd.n1993 vdd.n914 19.3944
R3511 vdd.n1993 vdd.n915 19.3944
R3512 vdd.n1988 vdd.n1987 19.3944
R3513 vdd.n1983 vdd.n1982 19.3944
R3514 vdd.n1982 vdd.n1981 19.3944
R3515 vdd.n1981 vdd.n919 19.3944
R3516 vdd.n1976 vdd.n919 19.3944
R3517 vdd.n1976 vdd.n1975 19.3944
R3518 vdd.n1975 vdd.n1974 19.3944
R3519 vdd.n1974 vdd.n926 19.3944
R3520 vdd.n1969 vdd.n926 19.3944
R3521 vdd.n1969 vdd.n1968 19.3944
R3522 vdd.n1968 vdd.n1967 19.3944
R3523 vdd.n1967 vdd.n933 19.3944
R3524 vdd.n1962 vdd.n933 19.3944
R3525 vdd.n1962 vdd.n1961 19.3944
R3526 vdd.n1790 vdd.n1555 19.3944
R3527 vdd.n1790 vdd.n1546 19.3944
R3528 vdd.n1803 vdd.n1546 19.3944
R3529 vdd.n1803 vdd.n1544 19.3944
R3530 vdd.n1807 vdd.n1544 19.3944
R3531 vdd.n1807 vdd.n1535 19.3944
R3532 vdd.n1820 vdd.n1535 19.3944
R3533 vdd.n1820 vdd.n1533 19.3944
R3534 vdd.n1825 vdd.n1533 19.3944
R3535 vdd.n1825 vdd.n1524 19.3944
R3536 vdd.n1837 vdd.n1524 19.3944
R3537 vdd.n1837 vdd.n1252 19.3944
R3538 vdd.n1841 vdd.n1252 19.3944
R3539 vdd.n1841 vdd.n1242 19.3944
R3540 vdd.n1854 vdd.n1242 19.3944
R3541 vdd.n1854 vdd.n1240 19.3944
R3542 vdd.n1858 vdd.n1240 19.3944
R3543 vdd.n1858 vdd.n1230 19.3944
R3544 vdd.n1873 vdd.n1230 19.3944
R3545 vdd.n1873 vdd.n1228 19.3944
R3546 vdd.n1877 vdd.n1228 19.3944
R3547 vdd.n2943 vdd.n477 19.3944
R3548 vdd.n2943 vdd.n475 19.3944
R3549 vdd.n2947 vdd.n475 19.3944
R3550 vdd.n2947 vdd.n465 19.3944
R3551 vdd.n2960 vdd.n465 19.3944
R3552 vdd.n2960 vdd.n463 19.3944
R3553 vdd.n2964 vdd.n463 19.3944
R3554 vdd.n2964 vdd.n453 19.3944
R3555 vdd.n2976 vdd.n453 19.3944
R3556 vdd.n2976 vdd.n451 19.3944
R3557 vdd.n2980 vdd.n451 19.3944
R3558 vdd.n2981 vdd.n2980 19.3944
R3559 vdd.n2982 vdd.n2981 19.3944
R3560 vdd.n2982 vdd.n449 19.3944
R3561 vdd.n2986 vdd.n449 19.3944
R3562 vdd.n2987 vdd.n2986 19.3944
R3563 vdd.n2988 vdd.n2987 19.3944
R3564 vdd.n2988 vdd.n446 19.3944
R3565 vdd.n2992 vdd.n446 19.3944
R3566 vdd.n2993 vdd.n2992 19.3944
R3567 vdd.n2994 vdd.n2993 19.3944
R3568 vdd.n3037 vdd.n404 19.3944
R3569 vdd.n3037 vdd.n410 19.3944
R3570 vdd.n3032 vdd.n410 19.3944
R3571 vdd.n3032 vdd.n3031 19.3944
R3572 vdd.n3031 vdd.n3030 19.3944
R3573 vdd.n3030 vdd.n417 19.3944
R3574 vdd.n3025 vdd.n417 19.3944
R3575 vdd.n3025 vdd.n3024 19.3944
R3576 vdd.n3024 vdd.n3023 19.3944
R3577 vdd.n3023 vdd.n424 19.3944
R3578 vdd.n3018 vdd.n424 19.3944
R3579 vdd.n3018 vdd.n3017 19.3944
R3580 vdd.n3017 vdd.n3016 19.3944
R3581 vdd.n3016 vdd.n431 19.3944
R3582 vdd.n3011 vdd.n431 19.3944
R3583 vdd.n3011 vdd.n3010 19.3944
R3584 vdd.n3010 vdd.n3009 19.3944
R3585 vdd.n3009 vdd.n438 19.3944
R3586 vdd.n3004 vdd.n438 19.3944
R3587 vdd.n3004 vdd.n3003 19.3944
R3588 vdd.n3076 vdd.n364 19.3944
R3589 vdd.n3076 vdd.n370 19.3944
R3590 vdd.n3071 vdd.n370 19.3944
R3591 vdd.n3071 vdd.n3070 19.3944
R3592 vdd.n3070 vdd.n3069 19.3944
R3593 vdd.n3069 vdd.n377 19.3944
R3594 vdd.n3064 vdd.n377 19.3944
R3595 vdd.n3064 vdd.n3063 19.3944
R3596 vdd.n3063 vdd.n3062 19.3944
R3597 vdd.n3062 vdd.n384 19.3944
R3598 vdd.n3057 vdd.n384 19.3944
R3599 vdd.n3057 vdd.n3056 19.3944
R3600 vdd.n3056 vdd.n3055 19.3944
R3601 vdd.n3055 vdd.n391 19.3944
R3602 vdd.n3050 vdd.n391 19.3944
R3603 vdd.n3050 vdd.n3049 19.3944
R3604 vdd.n3049 vdd.n3048 19.3944
R3605 vdd.n3048 vdd.n398 19.3944
R3606 vdd.n3043 vdd.n398 19.3944
R3607 vdd.n3043 vdd.n3042 19.3944
R3608 vdd.n3112 vdd.n3111 19.3944
R3609 vdd.n3111 vdd.n3110 19.3944
R3610 vdd.n3110 vdd.n336 19.3944
R3611 vdd.n337 vdd.n336 19.3944
R3612 vdd.n3103 vdd.n337 19.3944
R3613 vdd.n3103 vdd.n3102 19.3944
R3614 vdd.n3102 vdd.n3101 19.3944
R3615 vdd.n3101 vdd.n344 19.3944
R3616 vdd.n3096 vdd.n344 19.3944
R3617 vdd.n3096 vdd.n3095 19.3944
R3618 vdd.n3095 vdd.n3094 19.3944
R3619 vdd.n3094 vdd.n351 19.3944
R3620 vdd.n3089 vdd.n351 19.3944
R3621 vdd.n3089 vdd.n3088 19.3944
R3622 vdd.n3088 vdd.n3087 19.3944
R3623 vdd.n3087 vdd.n358 19.3944
R3624 vdd.n3082 vdd.n358 19.3944
R3625 vdd.n3082 vdd.n3081 19.3944
R3626 vdd.n2939 vdd.n480 19.3944
R3627 vdd.n2939 vdd.n471 19.3944
R3628 vdd.n2952 vdd.n471 19.3944
R3629 vdd.n2952 vdd.n469 19.3944
R3630 vdd.n2956 vdd.n469 19.3944
R3631 vdd.n2956 vdd.n460 19.3944
R3632 vdd.n2968 vdd.n460 19.3944
R3633 vdd.n2968 vdd.n458 19.3944
R3634 vdd.n2972 vdd.n458 19.3944
R3635 vdd.n2972 vdd.n300 19.3944
R3636 vdd.n3137 vdd.n300 19.3944
R3637 vdd.n3137 vdd.n301 19.3944
R3638 vdd.n3131 vdd.n301 19.3944
R3639 vdd.n3131 vdd.n3130 19.3944
R3640 vdd.n3130 vdd.n3129 19.3944
R3641 vdd.n3129 vdd.n313 19.3944
R3642 vdd.n3123 vdd.n313 19.3944
R3643 vdd.n3123 vdd.n3122 19.3944
R3644 vdd.n3122 vdd.n3121 19.3944
R3645 vdd.n3121 vdd.n324 19.3944
R3646 vdd.n3115 vdd.n324 19.3944
R3647 vdd.n2892 vdd.n536 19.3944
R3648 vdd.n2892 vdd.n2889 19.3944
R3649 vdd.n2889 vdd.n2886 19.3944
R3650 vdd.n2886 vdd.n2885 19.3944
R3651 vdd.n2885 vdd.n2882 19.3944
R3652 vdd.n2882 vdd.n2881 19.3944
R3653 vdd.n2881 vdd.n2878 19.3944
R3654 vdd.n2878 vdd.n2877 19.3944
R3655 vdd.n2877 vdd.n2874 19.3944
R3656 vdd.n2874 vdd.n2873 19.3944
R3657 vdd.n2873 vdd.n2870 19.3944
R3658 vdd.n2870 vdd.n2869 19.3944
R3659 vdd.n2869 vdd.n2866 19.3944
R3660 vdd.n2866 vdd.n2865 19.3944
R3661 vdd.n2865 vdd.n2862 19.3944
R3662 vdd.n2862 vdd.n2861 19.3944
R3663 vdd.n2861 vdd.n2858 19.3944
R3664 vdd.n2858 vdd.n2857 19.3944
R3665 vdd.n2857 vdd.n2854 19.3944
R3666 vdd.n2854 vdd.n2853 19.3944
R3667 vdd.n2935 vdd.n482 19.3944
R3668 vdd.n2930 vdd.n482 19.3944
R3669 vdd.n521 vdd.n518 19.3944
R3670 vdd.n2926 vdd.n2925 19.3944
R3671 vdd.n2925 vdd.n2922 19.3944
R3672 vdd.n2922 vdd.n2921 19.3944
R3673 vdd.n2921 vdd.n2918 19.3944
R3674 vdd.n2918 vdd.n2917 19.3944
R3675 vdd.n2917 vdd.n2914 19.3944
R3676 vdd.n2914 vdd.n2913 19.3944
R3677 vdd.n2913 vdd.n2910 19.3944
R3678 vdd.n2910 vdd.n2909 19.3944
R3679 vdd.n2909 vdd.n2906 19.3944
R3680 vdd.n2906 vdd.n2905 19.3944
R3681 vdd.n2905 vdd.n2902 19.3944
R3682 vdd.n2902 vdd.n2901 19.3944
R3683 vdd.n2846 vdd.n556 19.3944
R3684 vdd.n2846 vdd.n2843 19.3944
R3685 vdd.n2843 vdd.n2840 19.3944
R3686 vdd.n2840 vdd.n2839 19.3944
R3687 vdd.n2839 vdd.n2836 19.3944
R3688 vdd.n2836 vdd.n2835 19.3944
R3689 vdd.n2835 vdd.n2832 19.3944
R3690 vdd.n2832 vdd.n2831 19.3944
R3691 vdd.n2831 vdd.n2828 19.3944
R3692 vdd.n2828 vdd.n2827 19.3944
R3693 vdd.n2827 vdd.n2824 19.3944
R3694 vdd.n2824 vdd.n2823 19.3944
R3695 vdd.n2823 vdd.n2820 19.3944
R3696 vdd.n2820 vdd.n2819 19.3944
R3697 vdd.n2819 vdd.n2816 19.3944
R3698 vdd.n2816 vdd.n2815 19.3944
R3699 vdd.n2812 vdd.n2811 19.3944
R3700 vdd.n2808 vdd.n2807 19.3944
R3701 vdd.n1722 vdd.n1718 19.0066
R3702 vdd.n1921 vdd.n979 19.0066
R3703 vdd.n3041 vdd.n404 19.0066
R3704 vdd.n2850 vdd.n556 19.0066
R3705 vdd.n1044 vdd.n1043 16.0975
R3706 vdd.n772 vdd.n771 16.0975
R3707 vdd.n1683 vdd.n1682 16.0975
R3708 vdd.n1721 vdd.n1720 16.0975
R3709 vdd.n1617 vdd.n1616 16.0975
R3710 vdd.n1884 vdd.n1883 16.0975
R3711 vdd.n981 vdd.n980 16.0975
R3712 vdd.n941 vdd.n940 16.0975
R3713 vdd.n1064 vdd.n1063 16.0975
R3714 vdd.n763 vdd.n762 16.0975
R3715 vdd.n2319 vdd.n2318 16.0975
R3716 vdd.n3001 vdd.n3000 16.0975
R3717 vdd.n406 vdd.n405 16.0975
R3718 vdd.n366 vdd.n365 16.0975
R3719 vdd.n558 vdd.n557 16.0975
R3720 vdd.n2897 vdd.n2896 16.0975
R3721 vdd.n623 vdd.n622 16.0975
R3722 vdd.n2316 vdd.n2315 16.0975
R3723 vdd.n2804 vdd.n2803 16.0975
R3724 vdd.n590 vdd.n589 16.0975
R3725 vdd.t118 vdd.n2279 15.4182
R3726 vdd.n2552 vdd.t107 15.4182
R3727 vdd.n28 vdd.n27 14.5238
R3728 vdd.n2031 vdd.n866 14.0578
R3729 vdd.n2765 vdd.n484 14.0578
R3730 vdd.n292 vdd.n257 13.1884
R3731 vdd.n245 vdd.n210 13.1884
R3732 vdd.n202 vdd.n167 13.1884
R3733 vdd.n155 vdd.n120 13.1884
R3734 vdd.n113 vdd.n78 13.1884
R3735 vdd.n66 vdd.n31 13.1884
R3736 vdd.n1469 vdd.n1434 13.1884
R3737 vdd.n1516 vdd.n1481 13.1884
R3738 vdd.n1379 vdd.n1344 13.1884
R3739 vdd.n1426 vdd.n1391 13.1884
R3740 vdd.n1290 vdd.n1255 13.1884
R3741 vdd.n1337 vdd.n1302 13.1884
R3742 vdd.n1753 vdd.n1618 12.9944
R3743 vdd.n1757 vdd.n1618 12.9944
R3744 vdd.n1960 vdd.n939 12.9944
R3745 vdd.n1961 vdd.n1960 12.9944
R3746 vdd.n3080 vdd.n364 12.9944
R3747 vdd.n3081 vdd.n3080 12.9944
R3748 vdd.n2898 vdd.n536 12.9944
R3749 vdd.n2901 vdd.n2898 12.9944
R3750 vdd.n293 vdd.n255 12.8005
R3751 vdd.n288 vdd.n259 12.8005
R3752 vdd.n246 vdd.n208 12.8005
R3753 vdd.n241 vdd.n212 12.8005
R3754 vdd.n203 vdd.n165 12.8005
R3755 vdd.n198 vdd.n169 12.8005
R3756 vdd.n156 vdd.n118 12.8005
R3757 vdd.n151 vdd.n122 12.8005
R3758 vdd.n114 vdd.n76 12.8005
R3759 vdd.n109 vdd.n80 12.8005
R3760 vdd.n67 vdd.n29 12.8005
R3761 vdd.n62 vdd.n33 12.8005
R3762 vdd.n1470 vdd.n1432 12.8005
R3763 vdd.n1465 vdd.n1436 12.8005
R3764 vdd.n1517 vdd.n1479 12.8005
R3765 vdd.n1512 vdd.n1483 12.8005
R3766 vdd.n1380 vdd.n1342 12.8005
R3767 vdd.n1375 vdd.n1346 12.8005
R3768 vdd.n1427 vdd.n1389 12.8005
R3769 vdd.n1422 vdd.n1393 12.8005
R3770 vdd.n1291 vdd.n1253 12.8005
R3771 vdd.n1286 vdd.n1257 12.8005
R3772 vdd.n1338 vdd.n1300 12.8005
R3773 vdd.n1333 vdd.n1304 12.8005
R3774 vdd.n287 vdd.n260 12.0247
R3775 vdd.n240 vdd.n213 12.0247
R3776 vdd.n197 vdd.n170 12.0247
R3777 vdd.n150 vdd.n123 12.0247
R3778 vdd.n108 vdd.n81 12.0247
R3779 vdd.n61 vdd.n34 12.0247
R3780 vdd.n1464 vdd.n1437 12.0247
R3781 vdd.n1511 vdd.n1484 12.0247
R3782 vdd.n1374 vdd.n1347 12.0247
R3783 vdd.n1421 vdd.n1394 12.0247
R3784 vdd.n1285 vdd.n1258 12.0247
R3785 vdd.n1332 vdd.n1305 12.0247
R3786 vdd.n1792 vdd.n1548 11.337
R3787 vdd.n1801 vdd.n1548 11.337
R3788 vdd.n1801 vdd.n1800 11.337
R3789 vdd.n1809 vdd.n1542 11.337
R3790 vdd.n1818 vdd.n1817 11.337
R3791 vdd.n1835 vdd.n1526 11.337
R3792 vdd.n1843 vdd.n1249 11.337
R3793 vdd.n1852 vdd.n1851 11.337
R3794 vdd.n1860 vdd.n1232 11.337
R3795 vdd.n1871 vdd.n1232 11.337
R3796 vdd.n1871 vdd.n1870 11.337
R3797 vdd.n2941 vdd.n473 11.337
R3798 vdd.n2950 vdd.n473 11.337
R3799 vdd.n2950 vdd.n2949 11.337
R3800 vdd.n2958 vdd.n467 11.337
R3801 vdd.n2974 vdd.n456 11.337
R3802 vdd.n3135 vdd.n304 11.337
R3803 vdd.n3133 vdd.n308 11.337
R3804 vdd.n3127 vdd.n3126 11.337
R3805 vdd.n3125 vdd.n318 11.337
R3806 vdd.n3119 vdd.n318 11.337
R3807 vdd.n3119 vdd.n3118 11.337
R3808 vdd.n284 vdd.n283 11.249
R3809 vdd.n237 vdd.n236 11.249
R3810 vdd.n194 vdd.n193 11.249
R3811 vdd.n147 vdd.n146 11.249
R3812 vdd.n105 vdd.n104 11.249
R3813 vdd.n58 vdd.n57 11.249
R3814 vdd.n1461 vdd.n1460 11.249
R3815 vdd.n1508 vdd.n1507 11.249
R3816 vdd.n1371 vdd.n1370 11.249
R3817 vdd.n1418 vdd.n1417 11.249
R3818 vdd.n1282 vdd.n1281 11.249
R3819 vdd.n1329 vdd.n1328 11.249
R3820 vdd.n1590 vdd.t3 10.7702
R3821 vdd.t7 vdd.n3117 10.7702
R3822 vdd.n269 vdd.n268 10.7238
R3823 vdd.n222 vdd.n221 10.7238
R3824 vdd.n179 vdd.n178 10.7238
R3825 vdd.n132 vdd.n131 10.7238
R3826 vdd.n90 vdd.n89 10.7238
R3827 vdd.n43 vdd.n42 10.7238
R3828 vdd.n1446 vdd.n1445 10.7238
R3829 vdd.n1493 vdd.n1492 10.7238
R3830 vdd.n1356 vdd.n1355 10.7238
R3831 vdd.n1403 vdd.n1402 10.7238
R3832 vdd.n1267 vdd.n1266 10.7238
R3833 vdd.n1314 vdd.n1313 10.7238
R3834 vdd.n2207 vdd.t136 10.6568
R3835 vdd.t120 vdd.n718 10.6568
R3836 vdd.n2040 vdd.n864 10.6151
R3837 vdd.n2041 vdd.n2040 10.6151
R3838 vdd.n2042 vdd.n2041 10.6151
R3839 vdd.n2042 vdd.n853 10.6151
R3840 vdd.n2052 vdd.n853 10.6151
R3841 vdd.n2053 vdd.n2052 10.6151
R3842 vdd.n2054 vdd.n2053 10.6151
R3843 vdd.n2054 vdd.n840 10.6151
R3844 vdd.n2064 vdd.n840 10.6151
R3845 vdd.n2065 vdd.n2064 10.6151
R3846 vdd.n2066 vdd.n2065 10.6151
R3847 vdd.n2066 vdd.n828 10.6151
R3848 vdd.n2077 vdd.n828 10.6151
R3849 vdd.n2078 vdd.n2077 10.6151
R3850 vdd.n2079 vdd.n2078 10.6151
R3851 vdd.n2079 vdd.n816 10.6151
R3852 vdd.n2089 vdd.n816 10.6151
R3853 vdd.n2090 vdd.n2089 10.6151
R3854 vdd.n2091 vdd.n2090 10.6151
R3855 vdd.n2091 vdd.n804 10.6151
R3856 vdd.n2101 vdd.n804 10.6151
R3857 vdd.n2102 vdd.n2101 10.6151
R3858 vdd.n2103 vdd.n2102 10.6151
R3859 vdd.n2103 vdd.n793 10.6151
R3860 vdd.n2113 vdd.n793 10.6151
R3861 vdd.n2114 vdd.n2113 10.6151
R3862 vdd.n2115 vdd.n2114 10.6151
R3863 vdd.n2115 vdd.n780 10.6151
R3864 vdd.n2127 vdd.n780 10.6151
R3865 vdd.n2128 vdd.n2127 10.6151
R3866 vdd.n2130 vdd.n2128 10.6151
R3867 vdd.n2130 vdd.n2129 10.6151
R3868 vdd.n2129 vdd.n761 10.6151
R3869 vdd.n2277 vdd.n2276 10.6151
R3870 vdd.n2276 vdd.n2275 10.6151
R3871 vdd.n2275 vdd.n2272 10.6151
R3872 vdd.n2272 vdd.n2271 10.6151
R3873 vdd.n2271 vdd.n2268 10.6151
R3874 vdd.n2268 vdd.n2267 10.6151
R3875 vdd.n2267 vdd.n2264 10.6151
R3876 vdd.n2264 vdd.n2263 10.6151
R3877 vdd.n2263 vdd.n2260 10.6151
R3878 vdd.n2260 vdd.n2259 10.6151
R3879 vdd.n2259 vdd.n2256 10.6151
R3880 vdd.n2256 vdd.n2255 10.6151
R3881 vdd.n2255 vdd.n2252 10.6151
R3882 vdd.n2252 vdd.n2251 10.6151
R3883 vdd.n2251 vdd.n2248 10.6151
R3884 vdd.n2248 vdd.n2247 10.6151
R3885 vdd.n2247 vdd.n2244 10.6151
R3886 vdd.n2244 vdd.n2243 10.6151
R3887 vdd.n2243 vdd.n2240 10.6151
R3888 vdd.n2240 vdd.n2239 10.6151
R3889 vdd.n2239 vdd.n2236 10.6151
R3890 vdd.n2236 vdd.n2235 10.6151
R3891 vdd.n2235 vdd.n2232 10.6151
R3892 vdd.n2232 vdd.n2231 10.6151
R3893 vdd.n2231 vdd.n2228 10.6151
R3894 vdd.n2228 vdd.n2227 10.6151
R3895 vdd.n2227 vdd.n2224 10.6151
R3896 vdd.n2224 vdd.n2223 10.6151
R3897 vdd.n2223 vdd.n2220 10.6151
R3898 vdd.n2220 vdd.n2219 10.6151
R3899 vdd.n2219 vdd.n2216 10.6151
R3900 vdd.n2214 vdd.n2211 10.6151
R3901 vdd.n2211 vdd.n2210 10.6151
R3902 vdd.n1101 vdd.n1100 10.6151
R3903 vdd.n1103 vdd.n1101 10.6151
R3904 vdd.n1104 vdd.n1103 10.6151
R3905 vdd.n1106 vdd.n1104 10.6151
R3906 vdd.n1107 vdd.n1106 10.6151
R3907 vdd.n1109 vdd.n1107 10.6151
R3908 vdd.n1110 vdd.n1109 10.6151
R3909 vdd.n1112 vdd.n1110 10.6151
R3910 vdd.n1113 vdd.n1112 10.6151
R3911 vdd.n1115 vdd.n1113 10.6151
R3912 vdd.n1116 vdd.n1115 10.6151
R3913 vdd.n1118 vdd.n1116 10.6151
R3914 vdd.n1119 vdd.n1118 10.6151
R3915 vdd.n1121 vdd.n1119 10.6151
R3916 vdd.n1122 vdd.n1121 10.6151
R3917 vdd.n1124 vdd.n1122 10.6151
R3918 vdd.n1125 vdd.n1124 10.6151
R3919 vdd.n1147 vdd.n1125 10.6151
R3920 vdd.n1147 vdd.n1146 10.6151
R3921 vdd.n1146 vdd.n1145 10.6151
R3922 vdd.n1145 vdd.n1143 10.6151
R3923 vdd.n1143 vdd.n1142 10.6151
R3924 vdd.n1142 vdd.n1140 10.6151
R3925 vdd.n1140 vdd.n1139 10.6151
R3926 vdd.n1139 vdd.n1137 10.6151
R3927 vdd.n1137 vdd.n1136 10.6151
R3928 vdd.n1136 vdd.n1134 10.6151
R3929 vdd.n1134 vdd.n1133 10.6151
R3930 vdd.n1133 vdd.n1131 10.6151
R3931 vdd.n1131 vdd.n1130 10.6151
R3932 vdd.n1130 vdd.n1127 10.6151
R3933 vdd.n1127 vdd.n1126 10.6151
R3934 vdd.n1126 vdd.n764 10.6151
R3935 vdd.n2028 vdd.n2027 10.6151
R3936 vdd.n2027 vdd.n2026 10.6151
R3937 vdd.n2026 vdd.n2025 10.6151
R3938 vdd.n2025 vdd.n2023 10.6151
R3939 vdd.n2023 vdd.n2020 10.6151
R3940 vdd.n2020 vdd.n2019 10.6151
R3941 vdd.n2019 vdd.n2016 10.6151
R3942 vdd.n2016 vdd.n2015 10.6151
R3943 vdd.n2015 vdd.n2012 10.6151
R3944 vdd.n2012 vdd.n2011 10.6151
R3945 vdd.n2011 vdd.n2008 10.6151
R3946 vdd.n2008 vdd.n2007 10.6151
R3947 vdd.n2007 vdd.n2004 10.6151
R3948 vdd.n2004 vdd.n2003 10.6151
R3949 vdd.n2003 vdd.n2000 10.6151
R3950 vdd.n2000 vdd.n1999 10.6151
R3951 vdd.n1999 vdd.n1996 10.6151
R3952 vdd.n1996 vdd.n909 10.6151
R3953 vdd.n1067 vdd.n909 10.6151
R3954 vdd.n1068 vdd.n1067 10.6151
R3955 vdd.n1071 vdd.n1068 10.6151
R3956 vdd.n1072 vdd.n1071 10.6151
R3957 vdd.n1075 vdd.n1072 10.6151
R3958 vdd.n1076 vdd.n1075 10.6151
R3959 vdd.n1079 vdd.n1076 10.6151
R3960 vdd.n1080 vdd.n1079 10.6151
R3961 vdd.n1083 vdd.n1080 10.6151
R3962 vdd.n1084 vdd.n1083 10.6151
R3963 vdd.n1087 vdd.n1084 10.6151
R3964 vdd.n1088 vdd.n1087 10.6151
R3965 vdd.n1091 vdd.n1088 10.6151
R3966 vdd.n1096 vdd.n1093 10.6151
R3967 vdd.n1097 vdd.n1096 10.6151
R3968 vdd.n2480 vdd.n2479 10.6151
R3969 vdd.n2479 vdd.n2478 10.6151
R3970 vdd.n2478 vdd.n2317 10.6151
R3971 vdd.n2422 vdd.n2317 10.6151
R3972 vdd.n2423 vdd.n2422 10.6151
R3973 vdd.n2425 vdd.n2423 10.6151
R3974 vdd.n2426 vdd.n2425 10.6151
R3975 vdd.n2428 vdd.n2426 10.6151
R3976 vdd.n2429 vdd.n2428 10.6151
R3977 vdd.n2459 vdd.n2429 10.6151
R3978 vdd.n2459 vdd.n2458 10.6151
R3979 vdd.n2458 vdd.n2457 10.6151
R3980 vdd.n2457 vdd.n2455 10.6151
R3981 vdd.n2455 vdd.n2454 10.6151
R3982 vdd.n2454 vdd.n2452 10.6151
R3983 vdd.n2452 vdd.n2451 10.6151
R3984 vdd.n2451 vdd.n2449 10.6151
R3985 vdd.n2449 vdd.n2448 10.6151
R3986 vdd.n2448 vdd.n2446 10.6151
R3987 vdd.n2446 vdd.n2445 10.6151
R3988 vdd.n2445 vdd.n2443 10.6151
R3989 vdd.n2443 vdd.n2442 10.6151
R3990 vdd.n2442 vdd.n2440 10.6151
R3991 vdd.n2440 vdd.n2439 10.6151
R3992 vdd.n2439 vdd.n2437 10.6151
R3993 vdd.n2437 vdd.n2436 10.6151
R3994 vdd.n2436 vdd.n2434 10.6151
R3995 vdd.n2434 vdd.n2433 10.6151
R3996 vdd.n2433 vdd.n2431 10.6151
R3997 vdd.n2431 vdd.n2430 10.6151
R3998 vdd.n2430 vdd.n626 10.6151
R3999 vdd.n2698 vdd.n626 10.6151
R4000 vdd.n2699 vdd.n2698 10.6151
R4001 vdd.n2549 vdd.n2548 10.6151
R4002 vdd.n2548 vdd.n2547 10.6151
R4003 vdd.n2547 vdd.n2546 10.6151
R4004 vdd.n2546 vdd.n2544 10.6151
R4005 vdd.n2544 vdd.n2541 10.6151
R4006 vdd.n2541 vdd.n2540 10.6151
R4007 vdd.n2540 vdd.n2537 10.6151
R4008 vdd.n2537 vdd.n2536 10.6151
R4009 vdd.n2536 vdd.n2533 10.6151
R4010 vdd.n2533 vdd.n2532 10.6151
R4011 vdd.n2532 vdd.n2529 10.6151
R4012 vdd.n2529 vdd.n2528 10.6151
R4013 vdd.n2528 vdd.n2525 10.6151
R4014 vdd.n2525 vdd.n2524 10.6151
R4015 vdd.n2524 vdd.n2521 10.6151
R4016 vdd.n2521 vdd.n2520 10.6151
R4017 vdd.n2520 vdd.n2517 10.6151
R4018 vdd.n2517 vdd.n2516 10.6151
R4019 vdd.n2516 vdd.n2513 10.6151
R4020 vdd.n2513 vdd.n2512 10.6151
R4021 vdd.n2512 vdd.n2509 10.6151
R4022 vdd.n2509 vdd.n2508 10.6151
R4023 vdd.n2508 vdd.n2505 10.6151
R4024 vdd.n2505 vdd.n2504 10.6151
R4025 vdd.n2504 vdd.n2501 10.6151
R4026 vdd.n2501 vdd.n2500 10.6151
R4027 vdd.n2500 vdd.n2497 10.6151
R4028 vdd.n2497 vdd.n2496 10.6151
R4029 vdd.n2496 vdd.n2493 10.6151
R4030 vdd.n2493 vdd.n2492 10.6151
R4031 vdd.n2492 vdd.n2489 10.6151
R4032 vdd.n2487 vdd.n2484 10.6151
R4033 vdd.n2484 vdd.n2483 10.6151
R4034 vdd.n2561 vdd.n716 10.6151
R4035 vdd.n2562 vdd.n2561 10.6151
R4036 vdd.n2563 vdd.n2562 10.6151
R4037 vdd.n2563 vdd.n705 10.6151
R4038 vdd.n2573 vdd.n705 10.6151
R4039 vdd.n2574 vdd.n2573 10.6151
R4040 vdd.n2575 vdd.n2574 10.6151
R4041 vdd.n2575 vdd.n693 10.6151
R4042 vdd.n2585 vdd.n693 10.6151
R4043 vdd.n2586 vdd.n2585 10.6151
R4044 vdd.n2587 vdd.n2586 10.6151
R4045 vdd.n2587 vdd.n681 10.6151
R4046 vdd.n2597 vdd.n681 10.6151
R4047 vdd.n2598 vdd.n2597 10.6151
R4048 vdd.n2599 vdd.n2598 10.6151
R4049 vdd.n2599 vdd.n670 10.6151
R4050 vdd.n2609 vdd.n670 10.6151
R4051 vdd.n2610 vdd.n2609 10.6151
R4052 vdd.n2611 vdd.n2610 10.6151
R4053 vdd.n2611 vdd.n656 10.6151
R4054 vdd.n2622 vdd.n656 10.6151
R4055 vdd.n2623 vdd.n2622 10.6151
R4056 vdd.n2624 vdd.n2623 10.6151
R4057 vdd.n2624 vdd.n645 10.6151
R4058 vdd.n2634 vdd.n645 10.6151
R4059 vdd.n2635 vdd.n2634 10.6151
R4060 vdd.n2636 vdd.n2635 10.6151
R4061 vdd.n2636 vdd.n631 10.6151
R4062 vdd.n2691 vdd.n631 10.6151
R4063 vdd.n2692 vdd.n2691 10.6151
R4064 vdd.n2693 vdd.n2692 10.6151
R4065 vdd.n2693 vdd.n600 10.6151
R4066 vdd.n2763 vdd.n600 10.6151
R4067 vdd.n2762 vdd.n2761 10.6151
R4068 vdd.n2761 vdd.n601 10.6151
R4069 vdd.n602 vdd.n601 10.6151
R4070 vdd.n2754 vdd.n602 10.6151
R4071 vdd.n2754 vdd.n2753 10.6151
R4072 vdd.n2753 vdd.n2752 10.6151
R4073 vdd.n2752 vdd.n604 10.6151
R4074 vdd.n2747 vdd.n604 10.6151
R4075 vdd.n2747 vdd.n2746 10.6151
R4076 vdd.n2746 vdd.n2745 10.6151
R4077 vdd.n2745 vdd.n607 10.6151
R4078 vdd.n2740 vdd.n607 10.6151
R4079 vdd.n2740 vdd.n2739 10.6151
R4080 vdd.n2739 vdd.n2738 10.6151
R4081 vdd.n2738 vdd.n610 10.6151
R4082 vdd.n2733 vdd.n610 10.6151
R4083 vdd.n2733 vdd.n520 10.6151
R4084 vdd.n2729 vdd.n520 10.6151
R4085 vdd.n2729 vdd.n2728 10.6151
R4086 vdd.n2728 vdd.n2727 10.6151
R4087 vdd.n2727 vdd.n613 10.6151
R4088 vdd.n2722 vdd.n613 10.6151
R4089 vdd.n2722 vdd.n2721 10.6151
R4090 vdd.n2721 vdd.n2720 10.6151
R4091 vdd.n2720 vdd.n616 10.6151
R4092 vdd.n2715 vdd.n616 10.6151
R4093 vdd.n2715 vdd.n2714 10.6151
R4094 vdd.n2714 vdd.n2713 10.6151
R4095 vdd.n2713 vdd.n619 10.6151
R4096 vdd.n2708 vdd.n619 10.6151
R4097 vdd.n2708 vdd.n2707 10.6151
R4098 vdd.n2705 vdd.n624 10.6151
R4099 vdd.n2700 vdd.n624 10.6151
R4100 vdd.n2681 vdd.n2642 10.6151
R4101 vdd.n2676 vdd.n2642 10.6151
R4102 vdd.n2676 vdd.n2675 10.6151
R4103 vdd.n2675 vdd.n2674 10.6151
R4104 vdd.n2674 vdd.n2644 10.6151
R4105 vdd.n2669 vdd.n2644 10.6151
R4106 vdd.n2669 vdd.n2668 10.6151
R4107 vdd.n2668 vdd.n2667 10.6151
R4108 vdd.n2667 vdd.n2647 10.6151
R4109 vdd.n2662 vdd.n2647 10.6151
R4110 vdd.n2662 vdd.n2661 10.6151
R4111 vdd.n2661 vdd.n2660 10.6151
R4112 vdd.n2660 vdd.n2650 10.6151
R4113 vdd.n2655 vdd.n2650 10.6151
R4114 vdd.n2655 vdd.n2654 10.6151
R4115 vdd.n2654 vdd.n575 10.6151
R4116 vdd.n2798 vdd.n575 10.6151
R4117 vdd.n2798 vdd.n576 10.6151
R4118 vdd.n578 vdd.n576 10.6151
R4119 vdd.n2791 vdd.n578 10.6151
R4120 vdd.n2791 vdd.n2790 10.6151
R4121 vdd.n2790 vdd.n2789 10.6151
R4122 vdd.n2789 vdd.n580 10.6151
R4123 vdd.n2784 vdd.n580 10.6151
R4124 vdd.n2784 vdd.n2783 10.6151
R4125 vdd.n2783 vdd.n2782 10.6151
R4126 vdd.n2782 vdd.n583 10.6151
R4127 vdd.n2777 vdd.n583 10.6151
R4128 vdd.n2777 vdd.n2776 10.6151
R4129 vdd.n2776 vdd.n2775 10.6151
R4130 vdd.n2775 vdd.n586 10.6151
R4131 vdd.n2770 vdd.n2769 10.6151
R4132 vdd.n2769 vdd.n2768 10.6151
R4133 vdd.n2388 vdd.n2387 10.6151
R4134 vdd.n2474 vdd.n2388 10.6151
R4135 vdd.n2474 vdd.n2473 10.6151
R4136 vdd.n2473 vdd.n2472 10.6151
R4137 vdd.n2472 vdd.n2470 10.6151
R4138 vdd.n2470 vdd.n2469 10.6151
R4139 vdd.n2469 vdd.n2467 10.6151
R4140 vdd.n2467 vdd.n2466 10.6151
R4141 vdd.n2466 vdd.n2464 10.6151
R4142 vdd.n2464 vdd.n2463 10.6151
R4143 vdd.n2463 vdd.n2420 10.6151
R4144 vdd.n2420 vdd.n2419 10.6151
R4145 vdd.n2419 vdd.n2417 10.6151
R4146 vdd.n2417 vdd.n2416 10.6151
R4147 vdd.n2416 vdd.n2414 10.6151
R4148 vdd.n2414 vdd.n2413 10.6151
R4149 vdd.n2413 vdd.n2411 10.6151
R4150 vdd.n2411 vdd.n2410 10.6151
R4151 vdd.n2410 vdd.n2408 10.6151
R4152 vdd.n2408 vdd.n2407 10.6151
R4153 vdd.n2407 vdd.n2405 10.6151
R4154 vdd.n2405 vdd.n2404 10.6151
R4155 vdd.n2404 vdd.n2402 10.6151
R4156 vdd.n2402 vdd.n2401 10.6151
R4157 vdd.n2401 vdd.n2399 10.6151
R4158 vdd.n2399 vdd.n2398 10.6151
R4159 vdd.n2398 vdd.n2396 10.6151
R4160 vdd.n2396 vdd.n2395 10.6151
R4161 vdd.n2395 vdd.n2393 10.6151
R4162 vdd.n2393 vdd.n2392 10.6151
R4163 vdd.n2392 vdd.n2390 10.6151
R4164 vdd.n2390 vdd.n2389 10.6151
R4165 vdd.n2389 vdd.n592 10.6151
R4166 vdd.n2555 vdd.n722 10.6151
R4167 vdd.n2322 vdd.n722 10.6151
R4168 vdd.n2323 vdd.n2322 10.6151
R4169 vdd.n2326 vdd.n2323 10.6151
R4170 vdd.n2327 vdd.n2326 10.6151
R4171 vdd.n2330 vdd.n2327 10.6151
R4172 vdd.n2331 vdd.n2330 10.6151
R4173 vdd.n2334 vdd.n2331 10.6151
R4174 vdd.n2335 vdd.n2334 10.6151
R4175 vdd.n2338 vdd.n2335 10.6151
R4176 vdd.n2339 vdd.n2338 10.6151
R4177 vdd.n2342 vdd.n2339 10.6151
R4178 vdd.n2343 vdd.n2342 10.6151
R4179 vdd.n2346 vdd.n2343 10.6151
R4180 vdd.n2347 vdd.n2346 10.6151
R4181 vdd.n2350 vdd.n2347 10.6151
R4182 vdd.n2351 vdd.n2350 10.6151
R4183 vdd.n2354 vdd.n2351 10.6151
R4184 vdd.n2355 vdd.n2354 10.6151
R4185 vdd.n2358 vdd.n2355 10.6151
R4186 vdd.n2359 vdd.n2358 10.6151
R4187 vdd.n2362 vdd.n2359 10.6151
R4188 vdd.n2363 vdd.n2362 10.6151
R4189 vdd.n2366 vdd.n2363 10.6151
R4190 vdd.n2367 vdd.n2366 10.6151
R4191 vdd.n2370 vdd.n2367 10.6151
R4192 vdd.n2371 vdd.n2370 10.6151
R4193 vdd.n2374 vdd.n2371 10.6151
R4194 vdd.n2375 vdd.n2374 10.6151
R4195 vdd.n2378 vdd.n2375 10.6151
R4196 vdd.n2379 vdd.n2378 10.6151
R4197 vdd.n2384 vdd.n2382 10.6151
R4198 vdd.n2385 vdd.n2384 10.6151
R4199 vdd.n2557 vdd.n2556 10.6151
R4200 vdd.n2557 vdd.n711 10.6151
R4201 vdd.n2567 vdd.n711 10.6151
R4202 vdd.n2568 vdd.n2567 10.6151
R4203 vdd.n2569 vdd.n2568 10.6151
R4204 vdd.n2569 vdd.n699 10.6151
R4205 vdd.n2579 vdd.n699 10.6151
R4206 vdd.n2580 vdd.n2579 10.6151
R4207 vdd.n2581 vdd.n2580 10.6151
R4208 vdd.n2581 vdd.n687 10.6151
R4209 vdd.n2591 vdd.n687 10.6151
R4210 vdd.n2592 vdd.n2591 10.6151
R4211 vdd.n2593 vdd.n2592 10.6151
R4212 vdd.n2593 vdd.n676 10.6151
R4213 vdd.n2603 vdd.n676 10.6151
R4214 vdd.n2604 vdd.n2603 10.6151
R4215 vdd.n2605 vdd.n2604 10.6151
R4216 vdd.n2605 vdd.n663 10.6151
R4217 vdd.n2615 vdd.n663 10.6151
R4218 vdd.n2616 vdd.n2615 10.6151
R4219 vdd.n2618 vdd.n651 10.6151
R4220 vdd.n2628 vdd.n651 10.6151
R4221 vdd.n2629 vdd.n2628 10.6151
R4222 vdd.n2630 vdd.n2629 10.6151
R4223 vdd.n2630 vdd.n639 10.6151
R4224 vdd.n2640 vdd.n639 10.6151
R4225 vdd.n2641 vdd.n2640 10.6151
R4226 vdd.n2687 vdd.n2641 10.6151
R4227 vdd.n2687 vdd.n2686 10.6151
R4228 vdd.n2686 vdd.n2685 10.6151
R4229 vdd.n2685 vdd.n2684 10.6151
R4230 vdd.n2684 vdd.n2682 10.6151
R4231 vdd.n2036 vdd.n2035 10.6151
R4232 vdd.n2036 vdd.n859 10.6151
R4233 vdd.n2046 vdd.n859 10.6151
R4234 vdd.n2047 vdd.n2046 10.6151
R4235 vdd.n2048 vdd.n2047 10.6151
R4236 vdd.n2048 vdd.n847 10.6151
R4237 vdd.n2058 vdd.n847 10.6151
R4238 vdd.n2059 vdd.n2058 10.6151
R4239 vdd.n2060 vdd.n2059 10.6151
R4240 vdd.n2060 vdd.n834 10.6151
R4241 vdd.n2070 vdd.n834 10.6151
R4242 vdd.n2071 vdd.n2070 10.6151
R4243 vdd.n2073 vdd.n822 10.6151
R4244 vdd.n2083 vdd.n822 10.6151
R4245 vdd.n2084 vdd.n2083 10.6151
R4246 vdd.n2085 vdd.n2084 10.6151
R4247 vdd.n2085 vdd.n810 10.6151
R4248 vdd.n2095 vdd.n810 10.6151
R4249 vdd.n2096 vdd.n2095 10.6151
R4250 vdd.n2097 vdd.n2096 10.6151
R4251 vdd.n2097 vdd.n799 10.6151
R4252 vdd.n2107 vdd.n799 10.6151
R4253 vdd.n2108 vdd.n2107 10.6151
R4254 vdd.n2109 vdd.n2108 10.6151
R4255 vdd.n2109 vdd.n787 10.6151
R4256 vdd.n2119 vdd.n787 10.6151
R4257 vdd.n2120 vdd.n2119 10.6151
R4258 vdd.n2123 vdd.n2120 10.6151
R4259 vdd.n2123 vdd.n2122 10.6151
R4260 vdd.n2122 vdd.n2121 10.6151
R4261 vdd.n2121 vdd.n770 10.6151
R4262 vdd.n2205 vdd.n770 10.6151
R4263 vdd.n2204 vdd.n2203 10.6151
R4264 vdd.n2203 vdd.n2200 10.6151
R4265 vdd.n2200 vdd.n2199 10.6151
R4266 vdd.n2199 vdd.n2196 10.6151
R4267 vdd.n2196 vdd.n2195 10.6151
R4268 vdd.n2195 vdd.n2192 10.6151
R4269 vdd.n2192 vdd.n2191 10.6151
R4270 vdd.n2191 vdd.n2188 10.6151
R4271 vdd.n2188 vdd.n2187 10.6151
R4272 vdd.n2187 vdd.n2184 10.6151
R4273 vdd.n2184 vdd.n2183 10.6151
R4274 vdd.n2183 vdd.n2180 10.6151
R4275 vdd.n2180 vdd.n2179 10.6151
R4276 vdd.n2179 vdd.n2176 10.6151
R4277 vdd.n2176 vdd.n2175 10.6151
R4278 vdd.n2175 vdd.n2172 10.6151
R4279 vdd.n2172 vdd.n2171 10.6151
R4280 vdd.n2171 vdd.n2168 10.6151
R4281 vdd.n2168 vdd.n2167 10.6151
R4282 vdd.n2167 vdd.n2164 10.6151
R4283 vdd.n2164 vdd.n2163 10.6151
R4284 vdd.n2163 vdd.n2160 10.6151
R4285 vdd.n2160 vdd.n2159 10.6151
R4286 vdd.n2159 vdd.n2156 10.6151
R4287 vdd.n2156 vdd.n2155 10.6151
R4288 vdd.n2155 vdd.n2152 10.6151
R4289 vdd.n2152 vdd.n2151 10.6151
R4290 vdd.n2151 vdd.n2148 10.6151
R4291 vdd.n2148 vdd.n2147 10.6151
R4292 vdd.n2147 vdd.n2144 10.6151
R4293 vdd.n2144 vdd.n2143 10.6151
R4294 vdd.n2140 vdd.n2139 10.6151
R4295 vdd.n2139 vdd.n2137 10.6151
R4296 vdd.n1178 vdd.n1176 10.6151
R4297 vdd.n1176 vdd.n1175 10.6151
R4298 vdd.n1175 vdd.n1173 10.6151
R4299 vdd.n1173 vdd.n1172 10.6151
R4300 vdd.n1172 vdd.n1170 10.6151
R4301 vdd.n1170 vdd.n1169 10.6151
R4302 vdd.n1169 vdd.n1167 10.6151
R4303 vdd.n1167 vdd.n1166 10.6151
R4304 vdd.n1166 vdd.n1164 10.6151
R4305 vdd.n1164 vdd.n1163 10.6151
R4306 vdd.n1163 vdd.n1161 10.6151
R4307 vdd.n1161 vdd.n1160 10.6151
R4308 vdd.n1160 vdd.n1158 10.6151
R4309 vdd.n1158 vdd.n1157 10.6151
R4310 vdd.n1157 vdd.n1155 10.6151
R4311 vdd.n1155 vdd.n1154 10.6151
R4312 vdd.n1154 vdd.n1152 10.6151
R4313 vdd.n1152 vdd.n1151 10.6151
R4314 vdd.n1151 vdd.n1062 10.6151
R4315 vdd.n1062 vdd.n1061 10.6151
R4316 vdd.n1061 vdd.n1059 10.6151
R4317 vdd.n1059 vdd.n1058 10.6151
R4318 vdd.n1058 vdd.n1056 10.6151
R4319 vdd.n1056 vdd.n1055 10.6151
R4320 vdd.n1055 vdd.n1053 10.6151
R4321 vdd.n1053 vdd.n1052 10.6151
R4322 vdd.n1052 vdd.n1050 10.6151
R4323 vdd.n1050 vdd.n1049 10.6151
R4324 vdd.n1049 vdd.n1047 10.6151
R4325 vdd.n1047 vdd.n1046 10.6151
R4326 vdd.n1046 vdd.n774 10.6151
R4327 vdd.n2135 vdd.n774 10.6151
R4328 vdd.n2136 vdd.n2135 10.6151
R4329 vdd.n2034 vdd.n871 10.6151
R4330 vdd.n1013 vdd.n871 10.6151
R4331 vdd.n1014 vdd.n1013 10.6151
R4332 vdd.n1017 vdd.n1014 10.6151
R4333 vdd.n1018 vdd.n1017 10.6151
R4334 vdd.n1021 vdd.n1018 10.6151
R4335 vdd.n1022 vdd.n1021 10.6151
R4336 vdd.n1025 vdd.n1022 10.6151
R4337 vdd.n1026 vdd.n1025 10.6151
R4338 vdd.n1029 vdd.n1026 10.6151
R4339 vdd.n1030 vdd.n1029 10.6151
R4340 vdd.n1033 vdd.n1030 10.6151
R4341 vdd.n1034 vdd.n1033 10.6151
R4342 vdd.n1037 vdd.n1034 10.6151
R4343 vdd.n1038 vdd.n1037 10.6151
R4344 vdd.n1041 vdd.n1038 10.6151
R4345 vdd.n1212 vdd.n1041 10.6151
R4346 vdd.n1212 vdd.n1211 10.6151
R4347 vdd.n1211 vdd.n1209 10.6151
R4348 vdd.n1209 vdd.n1206 10.6151
R4349 vdd.n1206 vdd.n1205 10.6151
R4350 vdd.n1205 vdd.n1202 10.6151
R4351 vdd.n1202 vdd.n1201 10.6151
R4352 vdd.n1201 vdd.n1198 10.6151
R4353 vdd.n1198 vdd.n1197 10.6151
R4354 vdd.n1197 vdd.n1194 10.6151
R4355 vdd.n1194 vdd.n1193 10.6151
R4356 vdd.n1193 vdd.n1190 10.6151
R4357 vdd.n1190 vdd.n1189 10.6151
R4358 vdd.n1189 vdd.n1186 10.6151
R4359 vdd.n1186 vdd.n1185 10.6151
R4360 vdd.n1182 vdd.n1181 10.6151
R4361 vdd.n1181 vdd.n1179 10.6151
R4362 vdd.n280 vdd.n262 10.4732
R4363 vdd.n233 vdd.n215 10.4732
R4364 vdd.n190 vdd.n172 10.4732
R4365 vdd.n143 vdd.n125 10.4732
R4366 vdd.n101 vdd.n83 10.4732
R4367 vdd.n54 vdd.n36 10.4732
R4368 vdd.n1457 vdd.n1439 10.4732
R4369 vdd.n1504 vdd.n1486 10.4732
R4370 vdd.n1367 vdd.n1349 10.4732
R4371 vdd.n1414 vdd.n1396 10.4732
R4372 vdd.n1278 vdd.n1260 10.4732
R4373 vdd.n1325 vdd.n1307 10.4732
R4374 vdd.t166 vdd.n1250 10.3167
R4375 vdd.n2966 vdd.t78 10.3167
R4376 vdd.n1827 vdd.t89 10.09
R4377 vdd.n3134 vdd.t160 10.09
R4378 vdd.n1996 vdd.n1995 9.78206
R4379 vdd.n2928 vdd.n520 9.78206
R4380 vdd.n2799 vdd.n2798 9.78206
R4381 vdd.n1888 vdd.n1212 9.78206
R4382 vdd.n279 vdd.n264 9.69747
R4383 vdd.n232 vdd.n217 9.69747
R4384 vdd.n189 vdd.n174 9.69747
R4385 vdd.n142 vdd.n127 9.69747
R4386 vdd.n100 vdd.n85 9.69747
R4387 vdd.n53 vdd.n38 9.69747
R4388 vdd.n1456 vdd.n1441 9.69747
R4389 vdd.n1503 vdd.n1488 9.69747
R4390 vdd.n1366 vdd.n1351 9.69747
R4391 vdd.n1413 vdd.n1398 9.69747
R4392 vdd.n1277 vdd.n1262 9.69747
R4393 vdd.n1324 vdd.n1309 9.69747
R4394 vdd.n295 vdd.n294 9.45567
R4395 vdd.n248 vdd.n247 9.45567
R4396 vdd.n205 vdd.n204 9.45567
R4397 vdd.n158 vdd.n157 9.45567
R4398 vdd.n116 vdd.n115 9.45567
R4399 vdd.n69 vdd.n68 9.45567
R4400 vdd.n1472 vdd.n1471 9.45567
R4401 vdd.n1519 vdd.n1518 9.45567
R4402 vdd.n1382 vdd.n1381 9.45567
R4403 vdd.n1429 vdd.n1428 9.45567
R4404 vdd.n1293 vdd.n1292 9.45567
R4405 vdd.n1340 vdd.n1339 9.45567
R4406 vdd.n1958 vdd.n939 9.3005
R4407 vdd.n1957 vdd.n1956 9.3005
R4408 vdd.n945 vdd.n944 9.3005
R4409 vdd.n1951 vdd.n949 9.3005
R4410 vdd.n1950 vdd.n950 9.3005
R4411 vdd.n1949 vdd.n951 9.3005
R4412 vdd.n955 vdd.n952 9.3005
R4413 vdd.n1944 vdd.n956 9.3005
R4414 vdd.n1943 vdd.n957 9.3005
R4415 vdd.n1942 vdd.n958 9.3005
R4416 vdd.n962 vdd.n959 9.3005
R4417 vdd.n1937 vdd.n963 9.3005
R4418 vdd.n1936 vdd.n964 9.3005
R4419 vdd.n1935 vdd.n965 9.3005
R4420 vdd.n969 vdd.n966 9.3005
R4421 vdd.n1930 vdd.n970 9.3005
R4422 vdd.n1929 vdd.n971 9.3005
R4423 vdd.n1928 vdd.n972 9.3005
R4424 vdd.n976 vdd.n973 9.3005
R4425 vdd.n1923 vdd.n977 9.3005
R4426 vdd.n1922 vdd.n978 9.3005
R4427 vdd.n1921 vdd.n1920 9.3005
R4428 vdd.n1919 vdd.n979 9.3005
R4429 vdd.n1918 vdd.n1917 9.3005
R4430 vdd.n985 vdd.n984 9.3005
R4431 vdd.n1912 vdd.n989 9.3005
R4432 vdd.n1911 vdd.n990 9.3005
R4433 vdd.n1910 vdd.n991 9.3005
R4434 vdd.n995 vdd.n992 9.3005
R4435 vdd.n1905 vdd.n996 9.3005
R4436 vdd.n1904 vdd.n997 9.3005
R4437 vdd.n1903 vdd.n998 9.3005
R4438 vdd.n1002 vdd.n999 9.3005
R4439 vdd.n1898 vdd.n1003 9.3005
R4440 vdd.n1897 vdd.n1004 9.3005
R4441 vdd.n1896 vdd.n1005 9.3005
R4442 vdd.n1009 vdd.n1006 9.3005
R4443 vdd.n1891 vdd.n1010 9.3005
R4444 vdd.n1960 vdd.n1959 9.3005
R4445 vdd.n1982 vdd.n910 9.3005
R4446 vdd.n1981 vdd.n918 9.3005
R4447 vdd.n922 vdd.n919 9.3005
R4448 vdd.n1976 vdd.n923 9.3005
R4449 vdd.n1975 vdd.n924 9.3005
R4450 vdd.n1974 vdd.n925 9.3005
R4451 vdd.n929 vdd.n926 9.3005
R4452 vdd.n1969 vdd.n930 9.3005
R4453 vdd.n1968 vdd.n931 9.3005
R4454 vdd.n1967 vdd.n932 9.3005
R4455 vdd.n936 vdd.n933 9.3005
R4456 vdd.n1962 vdd.n937 9.3005
R4457 vdd.n1961 vdd.n938 9.3005
R4458 vdd.n1994 vdd.n1993 9.3005
R4459 vdd.n914 vdd.n913 9.3005
R4460 vdd.n1838 vdd.n1837 9.3005
R4461 vdd.n1839 vdd.n1252 9.3005
R4462 vdd.n1841 vdd.n1840 9.3005
R4463 vdd.n1242 vdd.n1241 9.3005
R4464 vdd.n1855 vdd.n1854 9.3005
R4465 vdd.n1856 vdd.n1240 9.3005
R4466 vdd.n1858 vdd.n1857 9.3005
R4467 vdd.n1230 vdd.n1229 9.3005
R4468 vdd.n1874 vdd.n1873 9.3005
R4469 vdd.n1875 vdd.n1228 9.3005
R4470 vdd.n1877 vdd.n1876 9.3005
R4471 vdd.n271 vdd.n270 9.3005
R4472 vdd.n266 vdd.n265 9.3005
R4473 vdd.n277 vdd.n276 9.3005
R4474 vdd.n279 vdd.n278 9.3005
R4475 vdd.n262 vdd.n261 9.3005
R4476 vdd.n285 vdd.n284 9.3005
R4477 vdd.n287 vdd.n286 9.3005
R4478 vdd.n259 vdd.n256 9.3005
R4479 vdd.n294 vdd.n293 9.3005
R4480 vdd.n224 vdd.n223 9.3005
R4481 vdd.n219 vdd.n218 9.3005
R4482 vdd.n230 vdd.n229 9.3005
R4483 vdd.n232 vdd.n231 9.3005
R4484 vdd.n215 vdd.n214 9.3005
R4485 vdd.n238 vdd.n237 9.3005
R4486 vdd.n240 vdd.n239 9.3005
R4487 vdd.n212 vdd.n209 9.3005
R4488 vdd.n247 vdd.n246 9.3005
R4489 vdd.n181 vdd.n180 9.3005
R4490 vdd.n176 vdd.n175 9.3005
R4491 vdd.n187 vdd.n186 9.3005
R4492 vdd.n189 vdd.n188 9.3005
R4493 vdd.n172 vdd.n171 9.3005
R4494 vdd.n195 vdd.n194 9.3005
R4495 vdd.n197 vdd.n196 9.3005
R4496 vdd.n169 vdd.n166 9.3005
R4497 vdd.n204 vdd.n203 9.3005
R4498 vdd.n134 vdd.n133 9.3005
R4499 vdd.n129 vdd.n128 9.3005
R4500 vdd.n140 vdd.n139 9.3005
R4501 vdd.n142 vdd.n141 9.3005
R4502 vdd.n125 vdd.n124 9.3005
R4503 vdd.n148 vdd.n147 9.3005
R4504 vdd.n150 vdd.n149 9.3005
R4505 vdd.n122 vdd.n119 9.3005
R4506 vdd.n157 vdd.n156 9.3005
R4507 vdd.n92 vdd.n91 9.3005
R4508 vdd.n87 vdd.n86 9.3005
R4509 vdd.n98 vdd.n97 9.3005
R4510 vdd.n100 vdd.n99 9.3005
R4511 vdd.n83 vdd.n82 9.3005
R4512 vdd.n106 vdd.n105 9.3005
R4513 vdd.n108 vdd.n107 9.3005
R4514 vdd.n80 vdd.n77 9.3005
R4515 vdd.n115 vdd.n114 9.3005
R4516 vdd.n45 vdd.n44 9.3005
R4517 vdd.n40 vdd.n39 9.3005
R4518 vdd.n51 vdd.n50 9.3005
R4519 vdd.n53 vdd.n52 9.3005
R4520 vdd.n36 vdd.n35 9.3005
R4521 vdd.n59 vdd.n58 9.3005
R4522 vdd.n61 vdd.n60 9.3005
R4523 vdd.n33 vdd.n30 9.3005
R4524 vdd.n68 vdd.n67 9.3005
R4525 vdd.n2850 vdd.n2849 9.3005
R4526 vdd.n2853 vdd.n555 9.3005
R4527 vdd.n2854 vdd.n554 9.3005
R4528 vdd.n2857 vdd.n553 9.3005
R4529 vdd.n2858 vdd.n552 9.3005
R4530 vdd.n2861 vdd.n551 9.3005
R4531 vdd.n2862 vdd.n550 9.3005
R4532 vdd.n2865 vdd.n549 9.3005
R4533 vdd.n2866 vdd.n548 9.3005
R4534 vdd.n2869 vdd.n547 9.3005
R4535 vdd.n2870 vdd.n546 9.3005
R4536 vdd.n2873 vdd.n545 9.3005
R4537 vdd.n2874 vdd.n544 9.3005
R4538 vdd.n2877 vdd.n543 9.3005
R4539 vdd.n2878 vdd.n542 9.3005
R4540 vdd.n2881 vdd.n541 9.3005
R4541 vdd.n2882 vdd.n540 9.3005
R4542 vdd.n2885 vdd.n539 9.3005
R4543 vdd.n2886 vdd.n538 9.3005
R4544 vdd.n2889 vdd.n537 9.3005
R4545 vdd.n2893 vdd.n2892 9.3005
R4546 vdd.n2894 vdd.n536 9.3005
R4547 vdd.n2898 vdd.n2895 9.3005
R4548 vdd.n2901 vdd.n535 9.3005
R4549 vdd.n2902 vdd.n534 9.3005
R4550 vdd.n2905 vdd.n533 9.3005
R4551 vdd.n2906 vdd.n532 9.3005
R4552 vdd.n2909 vdd.n531 9.3005
R4553 vdd.n2910 vdd.n530 9.3005
R4554 vdd.n2913 vdd.n529 9.3005
R4555 vdd.n2914 vdd.n528 9.3005
R4556 vdd.n2917 vdd.n527 9.3005
R4557 vdd.n2918 vdd.n526 9.3005
R4558 vdd.n2921 vdd.n525 9.3005
R4559 vdd.n2922 vdd.n524 9.3005
R4560 vdd.n2925 vdd.n519 9.3005
R4561 vdd.n482 vdd.n481 9.3005
R4562 vdd.n2936 vdd.n2935 9.3005
R4563 vdd.n2939 vdd.n2938 9.3005
R4564 vdd.n471 vdd.n470 9.3005
R4565 vdd.n2953 vdd.n2952 9.3005
R4566 vdd.n2954 vdd.n469 9.3005
R4567 vdd.n2956 vdd.n2955 9.3005
R4568 vdd.n460 vdd.n459 9.3005
R4569 vdd.n2969 vdd.n2968 9.3005
R4570 vdd.n2970 vdd.n458 9.3005
R4571 vdd.n2972 vdd.n2971 9.3005
R4572 vdd.n300 vdd.n298 9.3005
R4573 vdd.n2937 vdd.n480 9.3005
R4574 vdd.n3138 vdd.n3137 9.3005
R4575 vdd.n301 vdd.n299 9.3005
R4576 vdd.n3131 vdd.n310 9.3005
R4577 vdd.n3130 vdd.n311 9.3005
R4578 vdd.n3129 vdd.n312 9.3005
R4579 vdd.n320 vdd.n313 9.3005
R4580 vdd.n3123 vdd.n321 9.3005
R4581 vdd.n3122 vdd.n322 9.3005
R4582 vdd.n3121 vdd.n323 9.3005
R4583 vdd.n331 vdd.n324 9.3005
R4584 vdd.n3115 vdd.n3114 9.3005
R4585 vdd.n3111 vdd.n332 9.3005
R4586 vdd.n3110 vdd.n335 9.3005
R4587 vdd.n339 vdd.n336 9.3005
R4588 vdd.n340 vdd.n337 9.3005
R4589 vdd.n3103 vdd.n341 9.3005
R4590 vdd.n3102 vdd.n342 9.3005
R4591 vdd.n3101 vdd.n343 9.3005
R4592 vdd.n347 vdd.n344 9.3005
R4593 vdd.n3096 vdd.n348 9.3005
R4594 vdd.n3095 vdd.n349 9.3005
R4595 vdd.n3094 vdd.n350 9.3005
R4596 vdd.n354 vdd.n351 9.3005
R4597 vdd.n3089 vdd.n355 9.3005
R4598 vdd.n3088 vdd.n356 9.3005
R4599 vdd.n3087 vdd.n357 9.3005
R4600 vdd.n361 vdd.n358 9.3005
R4601 vdd.n3082 vdd.n362 9.3005
R4602 vdd.n3081 vdd.n363 9.3005
R4603 vdd.n3080 vdd.n3079 9.3005
R4604 vdd.n3078 vdd.n364 9.3005
R4605 vdd.n3077 vdd.n3076 9.3005
R4606 vdd.n370 vdd.n369 9.3005
R4607 vdd.n3071 vdd.n374 9.3005
R4608 vdd.n3070 vdd.n375 9.3005
R4609 vdd.n3069 vdd.n376 9.3005
R4610 vdd.n380 vdd.n377 9.3005
R4611 vdd.n3064 vdd.n381 9.3005
R4612 vdd.n3063 vdd.n382 9.3005
R4613 vdd.n3062 vdd.n383 9.3005
R4614 vdd.n387 vdd.n384 9.3005
R4615 vdd.n3057 vdd.n388 9.3005
R4616 vdd.n3056 vdd.n389 9.3005
R4617 vdd.n3055 vdd.n390 9.3005
R4618 vdd.n394 vdd.n391 9.3005
R4619 vdd.n3050 vdd.n395 9.3005
R4620 vdd.n3049 vdd.n396 9.3005
R4621 vdd.n3048 vdd.n397 9.3005
R4622 vdd.n401 vdd.n398 9.3005
R4623 vdd.n3043 vdd.n402 9.3005
R4624 vdd.n3042 vdd.n403 9.3005
R4625 vdd.n3041 vdd.n3040 9.3005
R4626 vdd.n3039 vdd.n404 9.3005
R4627 vdd.n3038 vdd.n3037 9.3005
R4628 vdd.n410 vdd.n409 9.3005
R4629 vdd.n3032 vdd.n414 9.3005
R4630 vdd.n3031 vdd.n415 9.3005
R4631 vdd.n3030 vdd.n416 9.3005
R4632 vdd.n420 vdd.n417 9.3005
R4633 vdd.n3025 vdd.n421 9.3005
R4634 vdd.n3024 vdd.n422 9.3005
R4635 vdd.n3023 vdd.n423 9.3005
R4636 vdd.n427 vdd.n424 9.3005
R4637 vdd.n3018 vdd.n428 9.3005
R4638 vdd.n3017 vdd.n429 9.3005
R4639 vdd.n3016 vdd.n430 9.3005
R4640 vdd.n434 vdd.n431 9.3005
R4641 vdd.n3011 vdd.n435 9.3005
R4642 vdd.n3010 vdd.n436 9.3005
R4643 vdd.n3009 vdd.n437 9.3005
R4644 vdd.n441 vdd.n438 9.3005
R4645 vdd.n3004 vdd.n442 9.3005
R4646 vdd.n3003 vdd.n443 9.3005
R4647 vdd.n2999 vdd.n2996 9.3005
R4648 vdd.n3113 vdd.n3112 9.3005
R4649 vdd.n2944 vdd.n2943 9.3005
R4650 vdd.n2945 vdd.n475 9.3005
R4651 vdd.n2947 vdd.n2946 9.3005
R4652 vdd.n465 vdd.n464 9.3005
R4653 vdd.n2961 vdd.n2960 9.3005
R4654 vdd.n2962 vdd.n463 9.3005
R4655 vdd.n2964 vdd.n2963 9.3005
R4656 vdd.n453 vdd.n452 9.3005
R4657 vdd.n2977 vdd.n2976 9.3005
R4658 vdd.n2978 vdd.n451 9.3005
R4659 vdd.n2980 vdd.n2979 9.3005
R4660 vdd.n2981 vdd.n450 9.3005
R4661 vdd.n2983 vdd.n2982 9.3005
R4662 vdd.n2984 vdd.n449 9.3005
R4663 vdd.n2986 vdd.n2985 9.3005
R4664 vdd.n2987 vdd.n447 9.3005
R4665 vdd.n2989 vdd.n2988 9.3005
R4666 vdd.n2990 vdd.n446 9.3005
R4667 vdd.n2992 vdd.n2991 9.3005
R4668 vdd.n2993 vdd.n444 9.3005
R4669 vdd.n2995 vdd.n2994 9.3005
R4670 vdd.n477 vdd.n476 9.3005
R4671 vdd.n2802 vdd.n2801 9.3005
R4672 vdd.n2807 vdd.n2800 9.3005
R4673 vdd.n2816 vdd.n572 9.3005
R4674 vdd.n2819 vdd.n571 9.3005
R4675 vdd.n2820 vdd.n570 9.3005
R4676 vdd.n2823 vdd.n569 9.3005
R4677 vdd.n2824 vdd.n568 9.3005
R4678 vdd.n2827 vdd.n567 9.3005
R4679 vdd.n2828 vdd.n566 9.3005
R4680 vdd.n2831 vdd.n565 9.3005
R4681 vdd.n2832 vdd.n564 9.3005
R4682 vdd.n2835 vdd.n563 9.3005
R4683 vdd.n2836 vdd.n562 9.3005
R4684 vdd.n2839 vdd.n561 9.3005
R4685 vdd.n2840 vdd.n560 9.3005
R4686 vdd.n2843 vdd.n559 9.3005
R4687 vdd.n2847 vdd.n2846 9.3005
R4688 vdd.n2848 vdd.n556 9.3005
R4689 vdd.n1887 vdd.n1886 9.3005
R4690 vdd.n1882 vdd.n1214 9.3005
R4691 vdd.n1795 vdd.n1794 9.3005
R4692 vdd.n1796 vdd.n1550 9.3005
R4693 vdd.n1798 vdd.n1797 9.3005
R4694 vdd.n1540 vdd.n1539 9.3005
R4695 vdd.n1812 vdd.n1811 9.3005
R4696 vdd.n1813 vdd.n1538 9.3005
R4697 vdd.n1815 vdd.n1814 9.3005
R4698 vdd.n1530 vdd.n1529 9.3005
R4699 vdd.n1830 vdd.n1829 9.3005
R4700 vdd.n1831 vdd.n1528 9.3005
R4701 vdd.n1833 vdd.n1832 9.3005
R4702 vdd.n1247 vdd.n1246 9.3005
R4703 vdd.n1846 vdd.n1845 9.3005
R4704 vdd.n1847 vdd.n1245 9.3005
R4705 vdd.n1849 vdd.n1848 9.3005
R4706 vdd.n1237 vdd.n1236 9.3005
R4707 vdd.n1863 vdd.n1862 9.3005
R4708 vdd.n1864 vdd.n1234 9.3005
R4709 vdd.n1868 vdd.n1867 9.3005
R4710 vdd.n1866 vdd.n1235 9.3005
R4711 vdd.n1865 vdd.n1225 9.3005
R4712 vdd.n1552 vdd.n1551 9.3005
R4713 vdd.n1688 vdd.n1687 9.3005
R4714 vdd.n1689 vdd.n1678 9.3005
R4715 vdd.n1691 vdd.n1690 9.3005
R4716 vdd.n1692 vdd.n1677 9.3005
R4717 vdd.n1694 vdd.n1693 9.3005
R4718 vdd.n1695 vdd.n1672 9.3005
R4719 vdd.n1697 vdd.n1696 9.3005
R4720 vdd.n1698 vdd.n1671 9.3005
R4721 vdd.n1700 vdd.n1699 9.3005
R4722 vdd.n1701 vdd.n1666 9.3005
R4723 vdd.n1703 vdd.n1702 9.3005
R4724 vdd.n1704 vdd.n1665 9.3005
R4725 vdd.n1706 vdd.n1705 9.3005
R4726 vdd.n1707 vdd.n1660 9.3005
R4727 vdd.n1709 vdd.n1708 9.3005
R4728 vdd.n1710 vdd.n1659 9.3005
R4729 vdd.n1712 vdd.n1711 9.3005
R4730 vdd.n1713 vdd.n1654 9.3005
R4731 vdd.n1715 vdd.n1714 9.3005
R4732 vdd.n1716 vdd.n1653 9.3005
R4733 vdd.n1718 vdd.n1717 9.3005
R4734 vdd.n1722 vdd.n1649 9.3005
R4735 vdd.n1724 vdd.n1723 9.3005
R4736 vdd.n1725 vdd.n1648 9.3005
R4737 vdd.n1727 vdd.n1726 9.3005
R4738 vdd.n1728 vdd.n1643 9.3005
R4739 vdd.n1730 vdd.n1729 9.3005
R4740 vdd.n1731 vdd.n1642 9.3005
R4741 vdd.n1733 vdd.n1732 9.3005
R4742 vdd.n1734 vdd.n1637 9.3005
R4743 vdd.n1736 vdd.n1735 9.3005
R4744 vdd.n1737 vdd.n1636 9.3005
R4745 vdd.n1739 vdd.n1738 9.3005
R4746 vdd.n1740 vdd.n1631 9.3005
R4747 vdd.n1742 vdd.n1741 9.3005
R4748 vdd.n1743 vdd.n1630 9.3005
R4749 vdd.n1745 vdd.n1744 9.3005
R4750 vdd.n1746 vdd.n1625 9.3005
R4751 vdd.n1748 vdd.n1747 9.3005
R4752 vdd.n1749 vdd.n1624 9.3005
R4753 vdd.n1751 vdd.n1750 9.3005
R4754 vdd.n1752 vdd.n1619 9.3005
R4755 vdd.n1754 vdd.n1753 9.3005
R4756 vdd.n1755 vdd.n1618 9.3005
R4757 vdd.n1757 vdd.n1756 9.3005
R4758 vdd.n1758 vdd.n1611 9.3005
R4759 vdd.n1760 vdd.n1759 9.3005
R4760 vdd.n1761 vdd.n1610 9.3005
R4761 vdd.n1763 vdd.n1762 9.3005
R4762 vdd.n1764 vdd.n1605 9.3005
R4763 vdd.n1766 vdd.n1765 9.3005
R4764 vdd.n1767 vdd.n1604 9.3005
R4765 vdd.n1769 vdd.n1768 9.3005
R4766 vdd.n1770 vdd.n1599 9.3005
R4767 vdd.n1772 vdd.n1771 9.3005
R4768 vdd.n1773 vdd.n1598 9.3005
R4769 vdd.n1775 vdd.n1774 9.3005
R4770 vdd.n1776 vdd.n1593 9.3005
R4771 vdd.n1778 vdd.n1777 9.3005
R4772 vdd.n1779 vdd.n1592 9.3005
R4773 vdd.n1781 vdd.n1780 9.3005
R4774 vdd.n1557 vdd.n1556 9.3005
R4775 vdd.n1787 vdd.n1786 9.3005
R4776 vdd.n1686 vdd.n1685 9.3005
R4777 vdd.n1790 vdd.n1789 9.3005
R4778 vdd.n1546 vdd.n1545 9.3005
R4779 vdd.n1804 vdd.n1803 9.3005
R4780 vdd.n1805 vdd.n1544 9.3005
R4781 vdd.n1807 vdd.n1806 9.3005
R4782 vdd.n1535 vdd.n1534 9.3005
R4783 vdd.n1821 vdd.n1820 9.3005
R4784 vdd.n1822 vdd.n1533 9.3005
R4785 vdd.n1825 vdd.n1824 9.3005
R4786 vdd.n1823 vdd.n1524 9.3005
R4787 vdd.n1788 vdd.n1555 9.3005
R4788 vdd.n1448 vdd.n1447 9.3005
R4789 vdd.n1443 vdd.n1442 9.3005
R4790 vdd.n1454 vdd.n1453 9.3005
R4791 vdd.n1456 vdd.n1455 9.3005
R4792 vdd.n1439 vdd.n1438 9.3005
R4793 vdd.n1462 vdd.n1461 9.3005
R4794 vdd.n1464 vdd.n1463 9.3005
R4795 vdd.n1436 vdd.n1433 9.3005
R4796 vdd.n1471 vdd.n1470 9.3005
R4797 vdd.n1495 vdd.n1494 9.3005
R4798 vdd.n1490 vdd.n1489 9.3005
R4799 vdd.n1501 vdd.n1500 9.3005
R4800 vdd.n1503 vdd.n1502 9.3005
R4801 vdd.n1486 vdd.n1485 9.3005
R4802 vdd.n1509 vdd.n1508 9.3005
R4803 vdd.n1511 vdd.n1510 9.3005
R4804 vdd.n1483 vdd.n1480 9.3005
R4805 vdd.n1518 vdd.n1517 9.3005
R4806 vdd.n1358 vdd.n1357 9.3005
R4807 vdd.n1353 vdd.n1352 9.3005
R4808 vdd.n1364 vdd.n1363 9.3005
R4809 vdd.n1366 vdd.n1365 9.3005
R4810 vdd.n1349 vdd.n1348 9.3005
R4811 vdd.n1372 vdd.n1371 9.3005
R4812 vdd.n1374 vdd.n1373 9.3005
R4813 vdd.n1346 vdd.n1343 9.3005
R4814 vdd.n1381 vdd.n1380 9.3005
R4815 vdd.n1405 vdd.n1404 9.3005
R4816 vdd.n1400 vdd.n1399 9.3005
R4817 vdd.n1411 vdd.n1410 9.3005
R4818 vdd.n1413 vdd.n1412 9.3005
R4819 vdd.n1396 vdd.n1395 9.3005
R4820 vdd.n1419 vdd.n1418 9.3005
R4821 vdd.n1421 vdd.n1420 9.3005
R4822 vdd.n1393 vdd.n1390 9.3005
R4823 vdd.n1428 vdd.n1427 9.3005
R4824 vdd.n1269 vdd.n1268 9.3005
R4825 vdd.n1264 vdd.n1263 9.3005
R4826 vdd.n1275 vdd.n1274 9.3005
R4827 vdd.n1277 vdd.n1276 9.3005
R4828 vdd.n1260 vdd.n1259 9.3005
R4829 vdd.n1283 vdd.n1282 9.3005
R4830 vdd.n1285 vdd.n1284 9.3005
R4831 vdd.n1257 vdd.n1254 9.3005
R4832 vdd.n1292 vdd.n1291 9.3005
R4833 vdd.n1316 vdd.n1315 9.3005
R4834 vdd.n1311 vdd.n1310 9.3005
R4835 vdd.n1322 vdd.n1321 9.3005
R4836 vdd.n1324 vdd.n1323 9.3005
R4837 vdd.n1307 vdd.n1306 9.3005
R4838 vdd.n1330 vdd.n1329 9.3005
R4839 vdd.n1332 vdd.n1331 9.3005
R4840 vdd.n1304 vdd.n1301 9.3005
R4841 vdd.n1339 vdd.n1338 9.3005
R4842 vdd.n1800 vdd.t145 8.95635
R4843 vdd.t84 vdd.n3125 8.95635
R4844 vdd.n276 vdd.n275 8.92171
R4845 vdd.n229 vdd.n228 8.92171
R4846 vdd.n186 vdd.n185 8.92171
R4847 vdd.n139 vdd.n138 8.92171
R4848 vdd.n97 vdd.n96 8.92171
R4849 vdd.n50 vdd.n49 8.92171
R4850 vdd.n1453 vdd.n1452 8.92171
R4851 vdd.n1500 vdd.n1499 8.92171
R4852 vdd.n1363 vdd.n1362 8.92171
R4853 vdd.n1410 vdd.n1409 8.92171
R4854 vdd.n1274 vdd.n1273 8.92171
R4855 vdd.n1321 vdd.n1320 8.92171
R4856 vdd.n207 vdd.n117 8.81535
R4857 vdd.n1431 vdd.n1341 8.81535
R4858 vdd.n1827 vdd.t158 8.72962
R4859 vdd.t164 vdd.n3134 8.72962
R4860 vdd.n1250 vdd.t86 8.50289
R4861 vdd.n1879 vdd.t23 8.50289
R4862 vdd.n516 vdd.t19 8.50289
R4863 vdd.n2966 vdd.t147 8.50289
R4864 vdd.n28 vdd.n14 8.42249
R4865 vdd.n3140 vdd.n3139 8.16225
R4866 vdd.n1523 vdd.n1522 8.16225
R4867 vdd.n272 vdd.n266 8.14595
R4868 vdd.n225 vdd.n219 8.14595
R4869 vdd.n182 vdd.n176 8.14595
R4870 vdd.n135 vdd.n129 8.14595
R4871 vdd.n93 vdd.n87 8.14595
R4872 vdd.n46 vdd.n40 8.14595
R4873 vdd.n1449 vdd.n1443 8.14595
R4874 vdd.n1496 vdd.n1490 8.14595
R4875 vdd.n1359 vdd.n1353 8.14595
R4876 vdd.n1406 vdd.n1400 8.14595
R4877 vdd.n1270 vdd.n1264 8.14595
R4878 vdd.n1317 vdd.n1311 8.14595
R4879 vdd.n2038 vdd.n866 7.70933
R4880 vdd.n2038 vdd.n869 7.70933
R4881 vdd.n2044 vdd.n855 7.70933
R4882 vdd.n2050 vdd.n855 7.70933
R4883 vdd.n2050 vdd.n849 7.70933
R4884 vdd.n2056 vdd.n849 7.70933
R4885 vdd.n2062 vdd.n842 7.70933
R4886 vdd.n2062 vdd.n845 7.70933
R4887 vdd.n2068 vdd.n838 7.70933
R4888 vdd.n2075 vdd.n824 7.70933
R4889 vdd.n2081 vdd.n824 7.70933
R4890 vdd.n2087 vdd.n818 7.70933
R4891 vdd.n2093 vdd.n814 7.70933
R4892 vdd.n2099 vdd.n808 7.70933
R4893 vdd.n2111 vdd.n795 7.70933
R4894 vdd.n2117 vdd.n789 7.70933
R4895 vdd.n2117 vdd.n782 7.70933
R4896 vdd.n2125 vdd.n782 7.70933
R4897 vdd.n2207 vdd.n766 7.70933
R4898 vdd.n2559 vdd.n718 7.70933
R4899 vdd.n2571 vdd.n707 7.70933
R4900 vdd.n2571 vdd.n701 7.70933
R4901 vdd.n2577 vdd.n701 7.70933
R4902 vdd.n2583 vdd.n695 7.70933
R4903 vdd.n2589 vdd.n691 7.70933
R4904 vdd.n2595 vdd.n685 7.70933
R4905 vdd.n2607 vdd.n672 7.70933
R4906 vdd.n2613 vdd.n665 7.70933
R4907 vdd.n2613 vdd.n668 7.70933
R4908 vdd.n2620 vdd.n660 7.70933
R4909 vdd.n2626 vdd.n647 7.70933
R4910 vdd.n2632 vdd.n647 7.70933
R4911 vdd.n2638 vdd.n641 7.70933
R4912 vdd.n2638 vdd.n633 7.70933
R4913 vdd.n2689 vdd.n633 7.70933
R4914 vdd.n2689 vdd.n636 7.70933
R4915 vdd.n2695 vdd.n595 7.70933
R4916 vdd.n2765 vdd.n595 7.70933
R4917 vdd.n2618 vdd.n2617 7.49318
R4918 vdd.n2072 vdd.n2071 7.49318
R4919 vdd.n271 vdd.n268 7.3702
R4920 vdd.n224 vdd.n221 7.3702
R4921 vdd.n181 vdd.n178 7.3702
R4922 vdd.n134 vdd.n131 7.3702
R4923 vdd.n92 vdd.n89 7.3702
R4924 vdd.n45 vdd.n42 7.3702
R4925 vdd.n1448 vdd.n1445 7.3702
R4926 vdd.n1495 vdd.n1492 7.3702
R4927 vdd.n1358 vdd.n1355 7.3702
R4928 vdd.n1405 vdd.n1402 7.3702
R4929 vdd.n1269 vdd.n1266 7.3702
R4930 vdd.n1316 vdd.n1313 7.3702
R4931 vdd.n2056 vdd.t106 7.36923
R4932 vdd.t127 vdd.n641 7.36923
R4933 vdd.n2132 vdd.t134 7.25587
R4934 vdd.n2476 vdd.t123 7.25587
R4935 vdd.n1723 vdd.n1722 6.98232
R4936 vdd.n1922 vdd.n1921 6.98232
R4937 vdd.n3042 vdd.n3041 6.98232
R4938 vdd.n2853 vdd.n2850 6.98232
R4939 vdd.n1860 vdd.t141 6.68904
R4940 vdd.n2949 vdd.t162 6.68904
R4941 vdd.t143 vdd.n1249 6.46231
R4942 vdd.n2974 vdd.t82 6.46231
R4943 vdd.n1818 vdd.t91 6.23558
R4944 vdd.t80 vdd.n308 6.23558
R4945 vdd.n3140 vdd.n297 6.22547
R4946 vdd.n1522 vdd.n1521 6.22547
R4947 vdd.t95 vdd.n795 5.89549
R4948 vdd.n2583 vdd.t132 5.89549
R4949 vdd.n272 vdd.n271 5.81868
R4950 vdd.n225 vdd.n224 5.81868
R4951 vdd.n182 vdd.n181 5.81868
R4952 vdd.n135 vdd.n134 5.81868
R4953 vdd.n93 vdd.n92 5.81868
R4954 vdd.n46 vdd.n45 5.81868
R4955 vdd.n1449 vdd.n1448 5.81868
R4956 vdd.n1496 vdd.n1495 5.81868
R4957 vdd.n1359 vdd.n1358 5.81868
R4958 vdd.n1406 vdd.n1405 5.81868
R4959 vdd.n1270 vdd.n1269 5.81868
R4960 vdd.n1317 vdd.n1316 5.81868
R4961 vdd.n2215 vdd.n2214 5.77611
R4962 vdd.n1093 vdd.n1092 5.77611
R4963 vdd.n2488 vdd.n2487 5.77611
R4964 vdd.n2706 vdd.n2705 5.77611
R4965 vdd.n2770 vdd.n591 5.77611
R4966 vdd.n2382 vdd.n2320 5.77611
R4967 vdd.n2140 vdd.n773 5.77611
R4968 vdd.n1182 vdd.n1045 5.77611
R4969 vdd.n1685 vdd.n1684 5.62474
R4970 vdd.n1885 vdd.n1882 5.62474
R4971 vdd.n3002 vdd.n2999 5.62474
R4972 vdd.n2805 vdd.n2802 5.62474
R4973 vdd.t109 vdd.n818 5.55539
R4974 vdd.n2087 vdd.t138 5.55539
R4975 vdd.t128 vdd.n672 5.55539
R4976 vdd.n2607 vdd.t114 5.55539
R4977 vdd.n838 vdd.t57 5.44203
R4978 vdd.n2620 vdd.t36 5.44203
R4979 vdd.n2044 vdd.t15 5.32866
R4980 vdd.n1128 vdd.t49 5.32866
R4981 vdd.n2565 vdd.t53 5.32866
R4982 vdd.n636 vdd.t11 5.32866
R4983 vdd.n1542 vdd.t91 5.10193
R4984 vdd.n3127 vdd.t80 5.10193
R4985 vdd.n275 vdd.n266 5.04292
R4986 vdd.n228 vdd.n219 5.04292
R4987 vdd.n185 vdd.n176 5.04292
R4988 vdd.n138 vdd.n129 5.04292
R4989 vdd.n96 vdd.n87 5.04292
R4990 vdd.n49 vdd.n40 5.04292
R4991 vdd.n1452 vdd.n1443 5.04292
R4992 vdd.n1499 vdd.n1490 5.04292
R4993 vdd.n1362 vdd.n1353 5.04292
R4994 vdd.n1409 vdd.n1400 5.04292
R4995 vdd.n1273 vdd.n1264 5.04292
R4996 vdd.n1320 vdd.n1311 5.04292
R4997 vdd.n2093 vdd.t130 4.98857
R4998 vdd.n685 vdd.t110 4.98857
R4999 vdd.n1835 vdd.t143 4.8752
R5000 vdd.t105 vdd.t115 4.8752
R5001 vdd.t94 vdd.t125 4.8752
R5002 vdd.t97 vdd.t99 4.8752
R5003 vdd.t139 vdd.t93 4.8752
R5004 vdd.t82 vdd.n304 4.8752
R5005 vdd.n2216 vdd.n2215 4.83952
R5006 vdd.n1092 vdd.n1091 4.83952
R5007 vdd.n2489 vdd.n2488 4.83952
R5008 vdd.n2707 vdd.n2706 4.83952
R5009 vdd.n591 vdd.n586 4.83952
R5010 vdd.n2379 vdd.n2320 4.83952
R5011 vdd.n2143 vdd.n773 4.83952
R5012 vdd.n1185 vdd.n1045 4.83952
R5013 vdd.n1890 vdd.n1889 4.74817
R5014 vdd.n1218 vdd.n1213 4.74817
R5015 vdd.n915 vdd.n912 4.74817
R5016 vdd.n1983 vdd.n911 4.74817
R5017 vdd.n1988 vdd.n912 4.74817
R5018 vdd.n1987 vdd.n911 4.74817
R5019 vdd.n2930 vdd.n2929 4.74817
R5020 vdd.n2927 vdd.n2926 4.74817
R5021 vdd.n2927 vdd.n521 4.74817
R5022 vdd.n2929 vdd.n518 4.74817
R5023 vdd.n2812 vdd.n573 4.74817
R5024 vdd.n2808 vdd.n574 4.74817
R5025 vdd.n2811 vdd.n574 4.74817
R5026 vdd.n2815 vdd.n573 4.74817
R5027 vdd.n1889 vdd.n1011 4.74817
R5028 vdd.n1215 vdd.n1213 4.74817
R5029 vdd.n297 vdd.n296 4.7074
R5030 vdd.n207 vdd.n206 4.7074
R5031 vdd.n1521 vdd.n1520 4.7074
R5032 vdd.n1431 vdd.n1430 4.7074
R5033 vdd.n1851 vdd.t141 4.64847
R5034 vdd.n2068 vdd.t122 4.64847
R5035 vdd.n808 vdd.t117 4.64847
R5036 vdd.n2589 vdd.t129 4.64847
R5037 vdd.n660 vdd.t102 4.64847
R5038 vdd.n2958 vdd.t162 4.64847
R5039 vdd.n276 vdd.n264 4.26717
R5040 vdd.n229 vdd.n217 4.26717
R5041 vdd.n186 vdd.n174 4.26717
R5042 vdd.n139 vdd.n127 4.26717
R5043 vdd.n97 vdd.n85 4.26717
R5044 vdd.n50 vdd.n38 4.26717
R5045 vdd.n1453 vdd.n1441 4.26717
R5046 vdd.n1500 vdd.n1488 4.26717
R5047 vdd.n1363 vdd.n1351 4.26717
R5048 vdd.n1410 vdd.n1398 4.26717
R5049 vdd.n1274 vdd.n1262 4.26717
R5050 vdd.n1321 vdd.n1309 4.26717
R5051 vdd.n297 vdd.n207 4.10845
R5052 vdd.n1521 vdd.n1431 4.10845
R5053 vdd.n253 vdd.t161 4.06363
R5054 vdd.n253 vdd.t81 4.06363
R5055 vdd.n251 vdd.t197 4.06363
R5056 vdd.n251 vdd.t165 4.06363
R5057 vdd.n249 vdd.t190 4.06363
R5058 vdd.n249 vdd.t202 4.06363
R5059 vdd.n163 vdd.t191 4.06363
R5060 vdd.n163 vdd.t193 4.06363
R5061 vdd.n161 vdd.t83 4.06363
R5062 vdd.n161 vdd.t178 4.06363
R5063 vdd.n159 vdd.t148 4.06363
R5064 vdd.n159 vdd.t88 4.06363
R5065 vdd.n74 vdd.t196 4.06363
R5066 vdd.n74 vdd.t177 4.06363
R5067 vdd.n72 vdd.t175 4.06363
R5068 vdd.n72 vdd.t181 4.06363
R5069 vdd.n70 vdd.t192 4.06363
R5070 vdd.n70 vdd.t79 4.06363
R5071 vdd.n1473 vdd.t167 4.06363
R5072 vdd.n1473 vdd.t201 4.06363
R5073 vdd.n1475 vdd.t159 4.06363
R5074 vdd.n1475 vdd.t144 4.06363
R5075 vdd.n1477 vdd.t182 4.06363
R5076 vdd.n1477 vdd.t90 4.06363
R5077 vdd.n1383 vdd.t198 4.06363
R5078 vdd.n1383 vdd.t87 4.06363
R5079 vdd.n1385 vdd.t199 4.06363
R5080 vdd.n1385 vdd.t149 4.06363
R5081 vdd.n1387 vdd.t169 4.06363
R5082 vdd.n1387 vdd.t194 4.06363
R5083 vdd.n1294 vdd.t183 4.06363
R5084 vdd.n1294 vdd.t189 4.06363
R5085 vdd.n1296 vdd.t168 4.06363
R5086 vdd.n1296 vdd.t176 4.06363
R5087 vdd.n1298 vdd.t92 4.06363
R5088 vdd.n1298 vdd.t195 4.06363
R5089 vdd.n26 vdd.t0 3.9605
R5090 vdd.n26 vdd.t1 3.9605
R5091 vdd.n23 vdd.t154 3.9605
R5092 vdd.n23 vdd.t185 3.9605
R5093 vdd.n21 vdd.t173 3.9605
R5094 vdd.n21 vdd.t156 3.9605
R5095 vdd.n20 vdd.t151 3.9605
R5096 vdd.n20 vdd.t152 3.9605
R5097 vdd.n15 vdd.t157 3.9605
R5098 vdd.n15 vdd.t153 3.9605
R5099 vdd.n16 vdd.t203 3.9605
R5100 vdd.n16 vdd.t186 3.9605
R5101 vdd.n18 vdd.t174 3.9605
R5102 vdd.n18 vdd.t155 3.9605
R5103 vdd.n25 vdd.t187 3.9605
R5104 vdd.n25 vdd.t188 3.9605
R5105 vdd.n2125 vdd.t112 3.85492
R5106 vdd.n1128 vdd.t112 3.85492
R5107 vdd.n2565 vdd.t100 3.85492
R5108 vdd.t100 vdd.n707 3.85492
R5109 vdd.n7 vdd.t140 3.61217
R5110 vdd.n7 vdd.t111 3.61217
R5111 vdd.n8 vdd.t98 3.61217
R5112 vdd.n8 vdd.t133 3.61217
R5113 vdd.n10 vdd.t124 3.61217
R5114 vdd.n10 vdd.t101 3.61217
R5115 vdd.n12 vdd.t108 3.61217
R5116 vdd.n12 vdd.t121 3.61217
R5117 vdd.n5 vdd.t137 3.61217
R5118 vdd.n5 vdd.t119 3.61217
R5119 vdd.n3 vdd.t113 3.61217
R5120 vdd.n3 vdd.t135 3.61217
R5121 vdd.n1 vdd.t96 3.61217
R5122 vdd.n1 vdd.t126 3.61217
R5123 vdd.n0 vdd.t131 3.61217
R5124 vdd.n0 vdd.t116 3.61217
R5125 vdd.n280 vdd.n279 3.49141
R5126 vdd.n233 vdd.n232 3.49141
R5127 vdd.n190 vdd.n189 3.49141
R5128 vdd.n143 vdd.n142 3.49141
R5129 vdd.n101 vdd.n100 3.49141
R5130 vdd.n54 vdd.n53 3.49141
R5131 vdd.n1457 vdd.n1456 3.49141
R5132 vdd.n1504 vdd.n1503 3.49141
R5133 vdd.n1367 vdd.n1366 3.49141
R5134 vdd.n1414 vdd.n1413 3.49141
R5135 vdd.n1278 vdd.n1277 3.49141
R5136 vdd.n1325 vdd.n1324 3.49141
R5137 vdd.n2279 vdd.t136 3.40145
R5138 vdd.n2552 vdd.t120 3.40145
R5139 vdd.n2617 vdd.n2616 3.12245
R5140 vdd.n2073 vdd.n2072 3.12245
R5141 vdd.n845 vdd.t122 3.06136
R5142 vdd.n2105 vdd.t117 3.06136
R5143 vdd.n2461 vdd.t129 3.06136
R5144 vdd.n2626 vdd.t102 3.06136
R5145 vdd.n1852 vdd.t86 2.83463
R5146 vdd.n1870 vdd.t23 2.83463
R5147 vdd.n2941 vdd.t19 2.83463
R5148 vdd.n467 vdd.t147 2.83463
R5149 vdd.n1149 vdd.t130 2.72126
R5150 vdd.n2601 vdd.t110 2.72126
R5151 vdd.n283 vdd.n262 2.71565
R5152 vdd.n236 vdd.n215 2.71565
R5153 vdd.n193 vdd.n172 2.71565
R5154 vdd.n146 vdd.n125 2.71565
R5155 vdd.n104 vdd.n83 2.71565
R5156 vdd.n57 vdd.n36 2.71565
R5157 vdd.n1460 vdd.n1439 2.71565
R5158 vdd.n1507 vdd.n1486 2.71565
R5159 vdd.n1370 vdd.n1349 2.71565
R5160 vdd.n1417 vdd.n1396 2.71565
R5161 vdd.n1281 vdd.n1260 2.71565
R5162 vdd.n1328 vdd.n1307 2.71565
R5163 vdd.t158 vdd.n1526 2.6079
R5164 vdd.n3135 vdd.t164 2.6079
R5165 vdd.t125 vdd.n789 2.49453
R5166 vdd.n2577 vdd.t97 2.49453
R5167 vdd.n270 vdd.n269 2.4129
R5168 vdd.n223 vdd.n222 2.4129
R5169 vdd.n180 vdd.n179 2.4129
R5170 vdd.n133 vdd.n132 2.4129
R5171 vdd.n91 vdd.n90 2.4129
R5172 vdd.n44 vdd.n43 2.4129
R5173 vdd.n1447 vdd.n1446 2.4129
R5174 vdd.n1494 vdd.n1493 2.4129
R5175 vdd.n1357 vdd.n1356 2.4129
R5176 vdd.n1404 vdd.n1403 2.4129
R5177 vdd.n1268 vdd.n1267 2.4129
R5178 vdd.n1315 vdd.n1314 2.4129
R5179 vdd.n1809 vdd.t145 2.38117
R5180 vdd.n869 vdd.t15 2.38117
R5181 vdd.n2132 vdd.t49 2.38117
R5182 vdd.n2476 vdd.t53 2.38117
R5183 vdd.n2695 vdd.t11 2.38117
R5184 vdd.n3126 vdd.t84 2.38117
R5185 vdd.n1995 vdd.n912 2.27742
R5186 vdd.n1995 vdd.n911 2.27742
R5187 vdd.n2928 vdd.n2927 2.27742
R5188 vdd.n2929 vdd.n2928 2.27742
R5189 vdd.n2799 vdd.n574 2.27742
R5190 vdd.n2799 vdd.n573 2.27742
R5191 vdd.n1889 vdd.n1888 2.27742
R5192 vdd.n1888 vdd.n1213 2.27742
R5193 vdd.n2081 vdd.t109 2.15444
R5194 vdd.n1149 vdd.t138 2.15444
R5195 vdd.n2601 vdd.t128 2.15444
R5196 vdd.t114 vdd.n665 2.15444
R5197 vdd.n284 vdd.n260 1.93989
R5198 vdd.n237 vdd.n213 1.93989
R5199 vdd.n194 vdd.n170 1.93989
R5200 vdd.n147 vdd.n123 1.93989
R5201 vdd.n105 vdd.n81 1.93989
R5202 vdd.n58 vdd.n34 1.93989
R5203 vdd.n1461 vdd.n1437 1.93989
R5204 vdd.n1508 vdd.n1484 1.93989
R5205 vdd.n1371 vdd.n1347 1.93989
R5206 vdd.n1418 vdd.n1394 1.93989
R5207 vdd.n1282 vdd.n1258 1.93989
R5208 vdd.n1329 vdd.n1305 1.93989
R5209 vdd.n2105 vdd.t95 1.81434
R5210 vdd.n2461 vdd.t132 1.81434
R5211 vdd.n2099 vdd.t115 1.58761
R5212 vdd.n691 vdd.t139 1.58761
R5213 vdd.n1817 vdd.t89 1.24752
R5214 vdd.n2075 vdd.t103 1.24752
R5215 vdd.n814 vdd.t105 1.24752
R5216 vdd.n2595 vdd.t93 1.24752
R5217 vdd.n668 vdd.t104 1.24752
R5218 vdd.t160 vdd.n3133 1.24752
R5219 vdd.n295 vdd.n255 1.16414
R5220 vdd.n288 vdd.n287 1.16414
R5221 vdd.n248 vdd.n208 1.16414
R5222 vdd.n241 vdd.n240 1.16414
R5223 vdd.n205 vdd.n165 1.16414
R5224 vdd.n198 vdd.n197 1.16414
R5225 vdd.n158 vdd.n118 1.16414
R5226 vdd.n151 vdd.n150 1.16414
R5227 vdd.n116 vdd.n76 1.16414
R5228 vdd.n109 vdd.n108 1.16414
R5229 vdd.n69 vdd.n29 1.16414
R5230 vdd.n62 vdd.n61 1.16414
R5231 vdd.n1472 vdd.n1432 1.16414
R5232 vdd.n1465 vdd.n1464 1.16414
R5233 vdd.n1519 vdd.n1479 1.16414
R5234 vdd.n1512 vdd.n1511 1.16414
R5235 vdd.n1382 vdd.n1342 1.16414
R5236 vdd.n1375 vdd.n1374 1.16414
R5237 vdd.n1429 vdd.n1389 1.16414
R5238 vdd.n1422 vdd.n1421 1.16414
R5239 vdd.n1293 vdd.n1253 1.16414
R5240 vdd.n1286 vdd.n1285 1.16414
R5241 vdd.n1340 vdd.n1300 1.16414
R5242 vdd.n1333 vdd.n1332 1.16414
R5243 vdd.n1843 vdd.t166 1.02079
R5244 vdd.t57 vdd.t103 1.02079
R5245 vdd.t104 vdd.t36 1.02079
R5246 vdd.t78 vdd.n456 1.02079
R5247 vdd.n1688 vdd.n1684 0.970197
R5248 vdd.n1886 vdd.n1885 0.970197
R5249 vdd.n3003 vdd.n3002 0.970197
R5250 vdd.n2807 vdd.n2805 0.970197
R5251 vdd.n1522 vdd.n28 0.852297
R5252 vdd vdd.n3140 0.844463
R5253 vdd.n1792 vdd.t3 0.567326
R5254 vdd.n3118 vdd.t7 0.567326
R5255 vdd.n1876 vdd.n913 0.537085
R5256 vdd.n2937 vdd.n2936 0.537085
R5257 vdd.n3114 vdd.n3113 0.537085
R5258 vdd.n2996 vdd.n2995 0.537085
R5259 vdd.n2801 vdd.n476 0.537085
R5260 vdd.n1865 vdd.n1214 0.537085
R5261 vdd.n1686 vdd.n1551 0.537085
R5262 vdd.n1788 vdd.n1787 0.537085
R5263 vdd.n4 vdd.n2 0.459552
R5264 vdd.n11 vdd.n9 0.459552
R5265 vdd.t134 vdd.n766 0.453961
R5266 vdd.n2559 vdd.t123 0.453961
R5267 vdd.n293 vdd.n292 0.388379
R5268 vdd.n259 vdd.n257 0.388379
R5269 vdd.n246 vdd.n245 0.388379
R5270 vdd.n212 vdd.n210 0.388379
R5271 vdd.n203 vdd.n202 0.388379
R5272 vdd.n169 vdd.n167 0.388379
R5273 vdd.n156 vdd.n155 0.388379
R5274 vdd.n122 vdd.n120 0.388379
R5275 vdd.n114 vdd.n113 0.388379
R5276 vdd.n80 vdd.n78 0.388379
R5277 vdd.n67 vdd.n66 0.388379
R5278 vdd.n33 vdd.n31 0.388379
R5279 vdd.n1470 vdd.n1469 0.388379
R5280 vdd.n1436 vdd.n1434 0.388379
R5281 vdd.n1517 vdd.n1516 0.388379
R5282 vdd.n1483 vdd.n1481 0.388379
R5283 vdd.n1380 vdd.n1379 0.388379
R5284 vdd.n1346 vdd.n1344 0.388379
R5285 vdd.n1427 vdd.n1426 0.388379
R5286 vdd.n1393 vdd.n1391 0.388379
R5287 vdd.n1291 vdd.n1290 0.388379
R5288 vdd.n1257 vdd.n1255 0.388379
R5289 vdd.n1338 vdd.n1337 0.388379
R5290 vdd.n1304 vdd.n1302 0.388379
R5291 vdd.n19 vdd.n17 0.387128
R5292 vdd.n24 vdd.n22 0.387128
R5293 vdd.n6 vdd.n4 0.358259
R5294 vdd.n13 vdd.n11 0.358259
R5295 vdd.n252 vdd.n250 0.358259
R5296 vdd.n254 vdd.n252 0.358259
R5297 vdd.n296 vdd.n254 0.358259
R5298 vdd.n162 vdd.n160 0.358259
R5299 vdd.n164 vdd.n162 0.358259
R5300 vdd.n206 vdd.n164 0.358259
R5301 vdd.n73 vdd.n71 0.358259
R5302 vdd.n75 vdd.n73 0.358259
R5303 vdd.n117 vdd.n75 0.358259
R5304 vdd.n1520 vdd.n1478 0.358259
R5305 vdd.n1478 vdd.n1476 0.358259
R5306 vdd.n1476 vdd.n1474 0.358259
R5307 vdd.n1430 vdd.n1388 0.358259
R5308 vdd.n1388 vdd.n1386 0.358259
R5309 vdd.n1386 vdd.n1384 0.358259
R5310 vdd.n1341 vdd.n1299 0.358259
R5311 vdd.n1299 vdd.n1297 0.358259
R5312 vdd.n1297 vdd.n1295 0.358259
R5313 vdd.t106 vdd.n842 0.340595
R5314 vdd.n2111 vdd.t94 0.340595
R5315 vdd.t99 vdd.n695 0.340595
R5316 vdd.n2632 vdd.t127 0.340595
R5317 vdd.n14 vdd.n6 0.334552
R5318 vdd.n14 vdd.n13 0.334552
R5319 vdd.n27 vdd.n19 0.21707
R5320 vdd.n27 vdd.n24 0.21707
R5321 vdd.n294 vdd.n256 0.155672
R5322 vdd.n286 vdd.n256 0.155672
R5323 vdd.n286 vdd.n285 0.155672
R5324 vdd.n285 vdd.n261 0.155672
R5325 vdd.n278 vdd.n261 0.155672
R5326 vdd.n278 vdd.n277 0.155672
R5327 vdd.n277 vdd.n265 0.155672
R5328 vdd.n270 vdd.n265 0.155672
R5329 vdd.n247 vdd.n209 0.155672
R5330 vdd.n239 vdd.n209 0.155672
R5331 vdd.n239 vdd.n238 0.155672
R5332 vdd.n238 vdd.n214 0.155672
R5333 vdd.n231 vdd.n214 0.155672
R5334 vdd.n231 vdd.n230 0.155672
R5335 vdd.n230 vdd.n218 0.155672
R5336 vdd.n223 vdd.n218 0.155672
R5337 vdd.n204 vdd.n166 0.155672
R5338 vdd.n196 vdd.n166 0.155672
R5339 vdd.n196 vdd.n195 0.155672
R5340 vdd.n195 vdd.n171 0.155672
R5341 vdd.n188 vdd.n171 0.155672
R5342 vdd.n188 vdd.n187 0.155672
R5343 vdd.n187 vdd.n175 0.155672
R5344 vdd.n180 vdd.n175 0.155672
R5345 vdd.n157 vdd.n119 0.155672
R5346 vdd.n149 vdd.n119 0.155672
R5347 vdd.n149 vdd.n148 0.155672
R5348 vdd.n148 vdd.n124 0.155672
R5349 vdd.n141 vdd.n124 0.155672
R5350 vdd.n141 vdd.n140 0.155672
R5351 vdd.n140 vdd.n128 0.155672
R5352 vdd.n133 vdd.n128 0.155672
R5353 vdd.n115 vdd.n77 0.155672
R5354 vdd.n107 vdd.n77 0.155672
R5355 vdd.n107 vdd.n106 0.155672
R5356 vdd.n106 vdd.n82 0.155672
R5357 vdd.n99 vdd.n82 0.155672
R5358 vdd.n99 vdd.n98 0.155672
R5359 vdd.n98 vdd.n86 0.155672
R5360 vdd.n91 vdd.n86 0.155672
R5361 vdd.n68 vdd.n30 0.155672
R5362 vdd.n60 vdd.n30 0.155672
R5363 vdd.n60 vdd.n59 0.155672
R5364 vdd.n59 vdd.n35 0.155672
R5365 vdd.n52 vdd.n35 0.155672
R5366 vdd.n52 vdd.n51 0.155672
R5367 vdd.n51 vdd.n39 0.155672
R5368 vdd.n44 vdd.n39 0.155672
R5369 vdd.n1471 vdd.n1433 0.155672
R5370 vdd.n1463 vdd.n1433 0.155672
R5371 vdd.n1463 vdd.n1462 0.155672
R5372 vdd.n1462 vdd.n1438 0.155672
R5373 vdd.n1455 vdd.n1438 0.155672
R5374 vdd.n1455 vdd.n1454 0.155672
R5375 vdd.n1454 vdd.n1442 0.155672
R5376 vdd.n1447 vdd.n1442 0.155672
R5377 vdd.n1518 vdd.n1480 0.155672
R5378 vdd.n1510 vdd.n1480 0.155672
R5379 vdd.n1510 vdd.n1509 0.155672
R5380 vdd.n1509 vdd.n1485 0.155672
R5381 vdd.n1502 vdd.n1485 0.155672
R5382 vdd.n1502 vdd.n1501 0.155672
R5383 vdd.n1501 vdd.n1489 0.155672
R5384 vdd.n1494 vdd.n1489 0.155672
R5385 vdd.n1381 vdd.n1343 0.155672
R5386 vdd.n1373 vdd.n1343 0.155672
R5387 vdd.n1373 vdd.n1372 0.155672
R5388 vdd.n1372 vdd.n1348 0.155672
R5389 vdd.n1365 vdd.n1348 0.155672
R5390 vdd.n1365 vdd.n1364 0.155672
R5391 vdd.n1364 vdd.n1352 0.155672
R5392 vdd.n1357 vdd.n1352 0.155672
R5393 vdd.n1428 vdd.n1390 0.155672
R5394 vdd.n1420 vdd.n1390 0.155672
R5395 vdd.n1420 vdd.n1419 0.155672
R5396 vdd.n1419 vdd.n1395 0.155672
R5397 vdd.n1412 vdd.n1395 0.155672
R5398 vdd.n1412 vdd.n1411 0.155672
R5399 vdd.n1411 vdd.n1399 0.155672
R5400 vdd.n1404 vdd.n1399 0.155672
R5401 vdd.n1292 vdd.n1254 0.155672
R5402 vdd.n1284 vdd.n1254 0.155672
R5403 vdd.n1284 vdd.n1283 0.155672
R5404 vdd.n1283 vdd.n1259 0.155672
R5405 vdd.n1276 vdd.n1259 0.155672
R5406 vdd.n1276 vdd.n1275 0.155672
R5407 vdd.n1275 vdd.n1263 0.155672
R5408 vdd.n1268 vdd.n1263 0.155672
R5409 vdd.n1339 vdd.n1301 0.155672
R5410 vdd.n1331 vdd.n1301 0.155672
R5411 vdd.n1331 vdd.n1330 0.155672
R5412 vdd.n1330 vdd.n1306 0.155672
R5413 vdd.n1323 vdd.n1306 0.155672
R5414 vdd.n1323 vdd.n1322 0.155672
R5415 vdd.n1322 vdd.n1310 0.155672
R5416 vdd.n1315 vdd.n1310 0.155672
R5417 vdd.n918 vdd.n910 0.152939
R5418 vdd.n922 vdd.n918 0.152939
R5419 vdd.n923 vdd.n922 0.152939
R5420 vdd.n924 vdd.n923 0.152939
R5421 vdd.n925 vdd.n924 0.152939
R5422 vdd.n929 vdd.n925 0.152939
R5423 vdd.n930 vdd.n929 0.152939
R5424 vdd.n931 vdd.n930 0.152939
R5425 vdd.n932 vdd.n931 0.152939
R5426 vdd.n936 vdd.n932 0.152939
R5427 vdd.n937 vdd.n936 0.152939
R5428 vdd.n938 vdd.n937 0.152939
R5429 vdd.n1959 vdd.n938 0.152939
R5430 vdd.n1959 vdd.n1958 0.152939
R5431 vdd.n1958 vdd.n1957 0.152939
R5432 vdd.n1957 vdd.n944 0.152939
R5433 vdd.n949 vdd.n944 0.152939
R5434 vdd.n950 vdd.n949 0.152939
R5435 vdd.n951 vdd.n950 0.152939
R5436 vdd.n955 vdd.n951 0.152939
R5437 vdd.n956 vdd.n955 0.152939
R5438 vdd.n957 vdd.n956 0.152939
R5439 vdd.n958 vdd.n957 0.152939
R5440 vdd.n962 vdd.n958 0.152939
R5441 vdd.n963 vdd.n962 0.152939
R5442 vdd.n964 vdd.n963 0.152939
R5443 vdd.n965 vdd.n964 0.152939
R5444 vdd.n969 vdd.n965 0.152939
R5445 vdd.n970 vdd.n969 0.152939
R5446 vdd.n971 vdd.n970 0.152939
R5447 vdd.n972 vdd.n971 0.152939
R5448 vdd.n976 vdd.n972 0.152939
R5449 vdd.n977 vdd.n976 0.152939
R5450 vdd.n978 vdd.n977 0.152939
R5451 vdd.n1920 vdd.n978 0.152939
R5452 vdd.n1920 vdd.n1919 0.152939
R5453 vdd.n1919 vdd.n1918 0.152939
R5454 vdd.n1918 vdd.n984 0.152939
R5455 vdd.n989 vdd.n984 0.152939
R5456 vdd.n990 vdd.n989 0.152939
R5457 vdd.n991 vdd.n990 0.152939
R5458 vdd.n995 vdd.n991 0.152939
R5459 vdd.n996 vdd.n995 0.152939
R5460 vdd.n997 vdd.n996 0.152939
R5461 vdd.n998 vdd.n997 0.152939
R5462 vdd.n1002 vdd.n998 0.152939
R5463 vdd.n1003 vdd.n1002 0.152939
R5464 vdd.n1004 vdd.n1003 0.152939
R5465 vdd.n1005 vdd.n1004 0.152939
R5466 vdd.n1009 vdd.n1005 0.152939
R5467 vdd.n1010 vdd.n1009 0.152939
R5468 vdd.n1994 vdd.n913 0.152939
R5469 vdd.n1839 vdd.n1838 0.152939
R5470 vdd.n1840 vdd.n1839 0.152939
R5471 vdd.n1840 vdd.n1241 0.152939
R5472 vdd.n1855 vdd.n1241 0.152939
R5473 vdd.n1856 vdd.n1855 0.152939
R5474 vdd.n1857 vdd.n1856 0.152939
R5475 vdd.n1857 vdd.n1229 0.152939
R5476 vdd.n1874 vdd.n1229 0.152939
R5477 vdd.n1875 vdd.n1874 0.152939
R5478 vdd.n1876 vdd.n1875 0.152939
R5479 vdd.n524 vdd.n519 0.152939
R5480 vdd.n525 vdd.n524 0.152939
R5481 vdd.n526 vdd.n525 0.152939
R5482 vdd.n527 vdd.n526 0.152939
R5483 vdd.n528 vdd.n527 0.152939
R5484 vdd.n529 vdd.n528 0.152939
R5485 vdd.n530 vdd.n529 0.152939
R5486 vdd.n531 vdd.n530 0.152939
R5487 vdd.n532 vdd.n531 0.152939
R5488 vdd.n533 vdd.n532 0.152939
R5489 vdd.n534 vdd.n533 0.152939
R5490 vdd.n535 vdd.n534 0.152939
R5491 vdd.n2895 vdd.n535 0.152939
R5492 vdd.n2895 vdd.n2894 0.152939
R5493 vdd.n2894 vdd.n2893 0.152939
R5494 vdd.n2893 vdd.n537 0.152939
R5495 vdd.n538 vdd.n537 0.152939
R5496 vdd.n539 vdd.n538 0.152939
R5497 vdd.n540 vdd.n539 0.152939
R5498 vdd.n541 vdd.n540 0.152939
R5499 vdd.n542 vdd.n541 0.152939
R5500 vdd.n543 vdd.n542 0.152939
R5501 vdd.n544 vdd.n543 0.152939
R5502 vdd.n545 vdd.n544 0.152939
R5503 vdd.n546 vdd.n545 0.152939
R5504 vdd.n547 vdd.n546 0.152939
R5505 vdd.n548 vdd.n547 0.152939
R5506 vdd.n549 vdd.n548 0.152939
R5507 vdd.n550 vdd.n549 0.152939
R5508 vdd.n551 vdd.n550 0.152939
R5509 vdd.n552 vdd.n551 0.152939
R5510 vdd.n553 vdd.n552 0.152939
R5511 vdd.n554 vdd.n553 0.152939
R5512 vdd.n555 vdd.n554 0.152939
R5513 vdd.n2849 vdd.n555 0.152939
R5514 vdd.n2849 vdd.n2848 0.152939
R5515 vdd.n2848 vdd.n2847 0.152939
R5516 vdd.n2847 vdd.n559 0.152939
R5517 vdd.n560 vdd.n559 0.152939
R5518 vdd.n561 vdd.n560 0.152939
R5519 vdd.n562 vdd.n561 0.152939
R5520 vdd.n563 vdd.n562 0.152939
R5521 vdd.n564 vdd.n563 0.152939
R5522 vdd.n565 vdd.n564 0.152939
R5523 vdd.n566 vdd.n565 0.152939
R5524 vdd.n567 vdd.n566 0.152939
R5525 vdd.n568 vdd.n567 0.152939
R5526 vdd.n569 vdd.n568 0.152939
R5527 vdd.n570 vdd.n569 0.152939
R5528 vdd.n571 vdd.n570 0.152939
R5529 vdd.n572 vdd.n571 0.152939
R5530 vdd.n2936 vdd.n481 0.152939
R5531 vdd.n2938 vdd.n2937 0.152939
R5532 vdd.n2938 vdd.n470 0.152939
R5533 vdd.n2953 vdd.n470 0.152939
R5534 vdd.n2954 vdd.n2953 0.152939
R5535 vdd.n2955 vdd.n2954 0.152939
R5536 vdd.n2955 vdd.n459 0.152939
R5537 vdd.n2969 vdd.n459 0.152939
R5538 vdd.n2970 vdd.n2969 0.152939
R5539 vdd.n2971 vdd.n2970 0.152939
R5540 vdd.n2971 vdd.n298 0.152939
R5541 vdd.n3138 vdd.n299 0.152939
R5542 vdd.n310 vdd.n299 0.152939
R5543 vdd.n311 vdd.n310 0.152939
R5544 vdd.n312 vdd.n311 0.152939
R5545 vdd.n320 vdd.n312 0.152939
R5546 vdd.n321 vdd.n320 0.152939
R5547 vdd.n322 vdd.n321 0.152939
R5548 vdd.n323 vdd.n322 0.152939
R5549 vdd.n331 vdd.n323 0.152939
R5550 vdd.n3114 vdd.n331 0.152939
R5551 vdd.n3113 vdd.n332 0.152939
R5552 vdd.n335 vdd.n332 0.152939
R5553 vdd.n339 vdd.n335 0.152939
R5554 vdd.n340 vdd.n339 0.152939
R5555 vdd.n341 vdd.n340 0.152939
R5556 vdd.n342 vdd.n341 0.152939
R5557 vdd.n343 vdd.n342 0.152939
R5558 vdd.n347 vdd.n343 0.152939
R5559 vdd.n348 vdd.n347 0.152939
R5560 vdd.n349 vdd.n348 0.152939
R5561 vdd.n350 vdd.n349 0.152939
R5562 vdd.n354 vdd.n350 0.152939
R5563 vdd.n355 vdd.n354 0.152939
R5564 vdd.n356 vdd.n355 0.152939
R5565 vdd.n357 vdd.n356 0.152939
R5566 vdd.n361 vdd.n357 0.152939
R5567 vdd.n362 vdd.n361 0.152939
R5568 vdd.n363 vdd.n362 0.152939
R5569 vdd.n3079 vdd.n363 0.152939
R5570 vdd.n3079 vdd.n3078 0.152939
R5571 vdd.n3078 vdd.n3077 0.152939
R5572 vdd.n3077 vdd.n369 0.152939
R5573 vdd.n374 vdd.n369 0.152939
R5574 vdd.n375 vdd.n374 0.152939
R5575 vdd.n376 vdd.n375 0.152939
R5576 vdd.n380 vdd.n376 0.152939
R5577 vdd.n381 vdd.n380 0.152939
R5578 vdd.n382 vdd.n381 0.152939
R5579 vdd.n383 vdd.n382 0.152939
R5580 vdd.n387 vdd.n383 0.152939
R5581 vdd.n388 vdd.n387 0.152939
R5582 vdd.n389 vdd.n388 0.152939
R5583 vdd.n390 vdd.n389 0.152939
R5584 vdd.n394 vdd.n390 0.152939
R5585 vdd.n395 vdd.n394 0.152939
R5586 vdd.n396 vdd.n395 0.152939
R5587 vdd.n397 vdd.n396 0.152939
R5588 vdd.n401 vdd.n397 0.152939
R5589 vdd.n402 vdd.n401 0.152939
R5590 vdd.n403 vdd.n402 0.152939
R5591 vdd.n3040 vdd.n403 0.152939
R5592 vdd.n3040 vdd.n3039 0.152939
R5593 vdd.n3039 vdd.n3038 0.152939
R5594 vdd.n3038 vdd.n409 0.152939
R5595 vdd.n414 vdd.n409 0.152939
R5596 vdd.n415 vdd.n414 0.152939
R5597 vdd.n416 vdd.n415 0.152939
R5598 vdd.n420 vdd.n416 0.152939
R5599 vdd.n421 vdd.n420 0.152939
R5600 vdd.n422 vdd.n421 0.152939
R5601 vdd.n423 vdd.n422 0.152939
R5602 vdd.n427 vdd.n423 0.152939
R5603 vdd.n428 vdd.n427 0.152939
R5604 vdd.n429 vdd.n428 0.152939
R5605 vdd.n430 vdd.n429 0.152939
R5606 vdd.n434 vdd.n430 0.152939
R5607 vdd.n435 vdd.n434 0.152939
R5608 vdd.n436 vdd.n435 0.152939
R5609 vdd.n437 vdd.n436 0.152939
R5610 vdd.n441 vdd.n437 0.152939
R5611 vdd.n442 vdd.n441 0.152939
R5612 vdd.n443 vdd.n442 0.152939
R5613 vdd.n2996 vdd.n443 0.152939
R5614 vdd.n2944 vdd.n476 0.152939
R5615 vdd.n2945 vdd.n2944 0.152939
R5616 vdd.n2946 vdd.n2945 0.152939
R5617 vdd.n2946 vdd.n464 0.152939
R5618 vdd.n2961 vdd.n464 0.152939
R5619 vdd.n2962 vdd.n2961 0.152939
R5620 vdd.n2963 vdd.n2962 0.152939
R5621 vdd.n2963 vdd.n452 0.152939
R5622 vdd.n2977 vdd.n452 0.152939
R5623 vdd.n2978 vdd.n2977 0.152939
R5624 vdd.n2979 vdd.n2978 0.152939
R5625 vdd.n2979 vdd.n450 0.152939
R5626 vdd.n2983 vdd.n450 0.152939
R5627 vdd.n2984 vdd.n2983 0.152939
R5628 vdd.n2985 vdd.n2984 0.152939
R5629 vdd.n2985 vdd.n447 0.152939
R5630 vdd.n2989 vdd.n447 0.152939
R5631 vdd.n2990 vdd.n2989 0.152939
R5632 vdd.n2991 vdd.n2990 0.152939
R5633 vdd.n2991 vdd.n444 0.152939
R5634 vdd.n2995 vdd.n444 0.152939
R5635 vdd.n2801 vdd.n2800 0.152939
R5636 vdd.n1887 vdd.n1214 0.152939
R5637 vdd.n1795 vdd.n1551 0.152939
R5638 vdd.n1796 vdd.n1795 0.152939
R5639 vdd.n1797 vdd.n1796 0.152939
R5640 vdd.n1797 vdd.n1539 0.152939
R5641 vdd.n1812 vdd.n1539 0.152939
R5642 vdd.n1813 vdd.n1812 0.152939
R5643 vdd.n1814 vdd.n1813 0.152939
R5644 vdd.n1814 vdd.n1529 0.152939
R5645 vdd.n1830 vdd.n1529 0.152939
R5646 vdd.n1831 vdd.n1830 0.152939
R5647 vdd.n1832 vdd.n1831 0.152939
R5648 vdd.n1832 vdd.n1246 0.152939
R5649 vdd.n1846 vdd.n1246 0.152939
R5650 vdd.n1847 vdd.n1846 0.152939
R5651 vdd.n1848 vdd.n1847 0.152939
R5652 vdd.n1848 vdd.n1236 0.152939
R5653 vdd.n1863 vdd.n1236 0.152939
R5654 vdd.n1864 vdd.n1863 0.152939
R5655 vdd.n1867 vdd.n1864 0.152939
R5656 vdd.n1867 vdd.n1866 0.152939
R5657 vdd.n1866 vdd.n1865 0.152939
R5658 vdd.n1787 vdd.n1556 0.152939
R5659 vdd.n1780 vdd.n1556 0.152939
R5660 vdd.n1780 vdd.n1779 0.152939
R5661 vdd.n1779 vdd.n1778 0.152939
R5662 vdd.n1778 vdd.n1593 0.152939
R5663 vdd.n1774 vdd.n1593 0.152939
R5664 vdd.n1774 vdd.n1773 0.152939
R5665 vdd.n1773 vdd.n1772 0.152939
R5666 vdd.n1772 vdd.n1599 0.152939
R5667 vdd.n1768 vdd.n1599 0.152939
R5668 vdd.n1768 vdd.n1767 0.152939
R5669 vdd.n1767 vdd.n1766 0.152939
R5670 vdd.n1766 vdd.n1605 0.152939
R5671 vdd.n1762 vdd.n1605 0.152939
R5672 vdd.n1762 vdd.n1761 0.152939
R5673 vdd.n1761 vdd.n1760 0.152939
R5674 vdd.n1760 vdd.n1611 0.152939
R5675 vdd.n1756 vdd.n1611 0.152939
R5676 vdd.n1756 vdd.n1755 0.152939
R5677 vdd.n1755 vdd.n1754 0.152939
R5678 vdd.n1754 vdd.n1619 0.152939
R5679 vdd.n1750 vdd.n1619 0.152939
R5680 vdd.n1750 vdd.n1749 0.152939
R5681 vdd.n1749 vdd.n1748 0.152939
R5682 vdd.n1748 vdd.n1625 0.152939
R5683 vdd.n1744 vdd.n1625 0.152939
R5684 vdd.n1744 vdd.n1743 0.152939
R5685 vdd.n1743 vdd.n1742 0.152939
R5686 vdd.n1742 vdd.n1631 0.152939
R5687 vdd.n1738 vdd.n1631 0.152939
R5688 vdd.n1738 vdd.n1737 0.152939
R5689 vdd.n1737 vdd.n1736 0.152939
R5690 vdd.n1736 vdd.n1637 0.152939
R5691 vdd.n1732 vdd.n1637 0.152939
R5692 vdd.n1732 vdd.n1731 0.152939
R5693 vdd.n1731 vdd.n1730 0.152939
R5694 vdd.n1730 vdd.n1643 0.152939
R5695 vdd.n1726 vdd.n1643 0.152939
R5696 vdd.n1726 vdd.n1725 0.152939
R5697 vdd.n1725 vdd.n1724 0.152939
R5698 vdd.n1724 vdd.n1649 0.152939
R5699 vdd.n1717 vdd.n1649 0.152939
R5700 vdd.n1717 vdd.n1716 0.152939
R5701 vdd.n1716 vdd.n1715 0.152939
R5702 vdd.n1715 vdd.n1654 0.152939
R5703 vdd.n1711 vdd.n1654 0.152939
R5704 vdd.n1711 vdd.n1710 0.152939
R5705 vdd.n1710 vdd.n1709 0.152939
R5706 vdd.n1709 vdd.n1660 0.152939
R5707 vdd.n1705 vdd.n1660 0.152939
R5708 vdd.n1705 vdd.n1704 0.152939
R5709 vdd.n1704 vdd.n1703 0.152939
R5710 vdd.n1703 vdd.n1666 0.152939
R5711 vdd.n1699 vdd.n1666 0.152939
R5712 vdd.n1699 vdd.n1698 0.152939
R5713 vdd.n1698 vdd.n1697 0.152939
R5714 vdd.n1697 vdd.n1672 0.152939
R5715 vdd.n1693 vdd.n1672 0.152939
R5716 vdd.n1693 vdd.n1692 0.152939
R5717 vdd.n1692 vdd.n1691 0.152939
R5718 vdd.n1691 vdd.n1678 0.152939
R5719 vdd.n1687 vdd.n1678 0.152939
R5720 vdd.n1687 vdd.n1686 0.152939
R5721 vdd.n1789 vdd.n1788 0.152939
R5722 vdd.n1789 vdd.n1545 0.152939
R5723 vdd.n1804 vdd.n1545 0.152939
R5724 vdd.n1805 vdd.n1804 0.152939
R5725 vdd.n1806 vdd.n1805 0.152939
R5726 vdd.n1806 vdd.n1534 0.152939
R5727 vdd.n1821 vdd.n1534 0.152939
R5728 vdd.n1822 vdd.n1821 0.152939
R5729 vdd.n1824 vdd.n1822 0.152939
R5730 vdd.n1824 vdd.n1823 0.152939
R5731 vdd.n1995 vdd.n1994 0.110256
R5732 vdd.n2928 vdd.n481 0.110256
R5733 vdd.n2800 vdd.n2799 0.110256
R5734 vdd.n1888 vdd.n1887 0.110256
R5735 vdd.n1838 vdd.n1523 0.0695946
R5736 vdd.n3139 vdd.n298 0.0695946
R5737 vdd.n3139 vdd.n3138 0.0695946
R5738 vdd.n1823 vdd.n1523 0.0695946
R5739 vdd.n1995 vdd.n910 0.0431829
R5740 vdd.n1888 vdd.n1010 0.0431829
R5741 vdd.n2928 vdd.n519 0.0431829
R5742 vdd.n2799 vdd.n572 0.0431829
R5743 vdd vdd.n28 0.00833333
R5744 a_n6308_8799.n99 a_n6308_8799.t67 485.149
R5745 a_n6308_8799.n106 a_n6308_8799.t75 485.149
R5746 a_n6308_8799.n114 a_n6308_8799.t82 485.149
R5747 a_n6308_8799.n75 a_n6308_8799.t54 485.149
R5748 a_n6308_8799.n82 a_n6308_8799.t57 485.149
R5749 a_n6308_8799.n90 a_n6308_8799.t83 485.149
R5750 a_n6308_8799.n25 a_n6308_8799.t59 485.135
R5751 a_n6308_8799.n103 a_n6308_8799.t49 464.166
R5752 a_n6308_8799.n97 a_n6308_8799.t81 464.166
R5753 a_n6308_8799.n102 a_n6308_8799.t64 464.166
R5754 a_n6308_8799.n101 a_n6308_8799.t63 464.166
R5755 a_n6308_8799.n98 a_n6308_8799.t41 464.166
R5756 a_n6308_8799.n100 a_n6308_8799.t69 464.166
R5757 a_n6308_8799.n30 a_n6308_8799.t62 485.135
R5758 a_n6308_8799.n110 a_n6308_8799.t55 464.166
R5759 a_n6308_8799.n104 a_n6308_8799.t87 464.166
R5760 a_n6308_8799.n109 a_n6308_8799.t74 464.166
R5761 a_n6308_8799.n108 a_n6308_8799.t73 464.166
R5762 a_n6308_8799.n105 a_n6308_8799.t46 464.166
R5763 a_n6308_8799.n107 a_n6308_8799.t76 464.166
R5764 a_n6308_8799.n35 a_n6308_8799.t79 485.135
R5765 a_n6308_8799.n118 a_n6308_8799.t47 464.166
R5766 a_n6308_8799.n112 a_n6308_8799.t68 464.166
R5767 a_n6308_8799.n117 a_n6308_8799.t42 464.166
R5768 a_n6308_8799.n116 a_n6308_8799.t52 464.166
R5769 a_n6308_8799.n113 a_n6308_8799.t85 464.166
R5770 a_n6308_8799.n115 a_n6308_8799.t72 464.166
R5771 a_n6308_8799.n76 a_n6308_8799.t53 464.166
R5772 a_n6308_8799.n77 a_n6308_8799.t70 464.166
R5773 a_n6308_8799.n78 a_n6308_8799.t40 464.166
R5774 a_n6308_8799.n79 a_n6308_8799.t51 464.166
R5775 a_n6308_8799.n74 a_n6308_8799.t60 464.166
R5776 a_n6308_8799.n80 a_n6308_8799.t80 464.166
R5777 a_n6308_8799.n83 a_n6308_8799.t58 464.166
R5778 a_n6308_8799.n84 a_n6308_8799.t77 464.166
R5779 a_n6308_8799.n85 a_n6308_8799.t44 464.166
R5780 a_n6308_8799.n86 a_n6308_8799.t56 464.166
R5781 a_n6308_8799.n81 a_n6308_8799.t65 464.166
R5782 a_n6308_8799.n87 a_n6308_8799.t86 464.166
R5783 a_n6308_8799.n91 a_n6308_8799.t71 464.166
R5784 a_n6308_8799.n92 a_n6308_8799.t84 464.166
R5785 a_n6308_8799.n93 a_n6308_8799.t61 464.166
R5786 a_n6308_8799.n94 a_n6308_8799.t43 464.166
R5787 a_n6308_8799.n89 a_n6308_8799.t66 464.166
R5788 a_n6308_8799.n95 a_n6308_8799.t48 464.166
R5789 a_n6308_8799.n20 a_n6308_8799.n29 72.3034
R5790 a_n6308_8799.n29 a_n6308_8799.n98 16.6962
R5791 a_n6308_8799.n28 a_n6308_8799.n20 77.6622
R5792 a_n6308_8799.n101 a_n6308_8799.n28 5.97853
R5793 a_n6308_8799.n27 a_n6308_8799.n19 77.6622
R5794 a_n6308_8799.n19 a_n6308_8799.n26 72.3034
R5795 a_n6308_8799.n103 a_n6308_8799.n25 20.9683
R5796 a_n6308_8799.n21 a_n6308_8799.n25 70.1674
R5797 a_n6308_8799.n17 a_n6308_8799.n34 72.3034
R5798 a_n6308_8799.n34 a_n6308_8799.n105 16.6962
R5799 a_n6308_8799.n33 a_n6308_8799.n17 77.6622
R5800 a_n6308_8799.n108 a_n6308_8799.n33 5.97853
R5801 a_n6308_8799.n32 a_n6308_8799.n16 77.6622
R5802 a_n6308_8799.n16 a_n6308_8799.n31 72.3034
R5803 a_n6308_8799.n110 a_n6308_8799.n30 20.9683
R5804 a_n6308_8799.n18 a_n6308_8799.n30 70.1674
R5805 a_n6308_8799.n14 a_n6308_8799.n39 72.3034
R5806 a_n6308_8799.n39 a_n6308_8799.n113 16.6962
R5807 a_n6308_8799.n38 a_n6308_8799.n14 77.6622
R5808 a_n6308_8799.n116 a_n6308_8799.n38 5.97853
R5809 a_n6308_8799.n37 a_n6308_8799.n13 77.6622
R5810 a_n6308_8799.n13 a_n6308_8799.n36 72.3034
R5811 a_n6308_8799.n118 a_n6308_8799.n35 20.9683
R5812 a_n6308_8799.n15 a_n6308_8799.n35 70.1674
R5813 a_n6308_8799.n11 a_n6308_8799.n44 70.1674
R5814 a_n6308_8799.n80 a_n6308_8799.n44 20.9683
R5815 a_n6308_8799.n43 a_n6308_8799.n11 72.3034
R5816 a_n6308_8799.n43 a_n6308_8799.n74 16.6962
R5817 a_n6308_8799.n10 a_n6308_8799.n42 77.6622
R5818 a_n6308_8799.n79 a_n6308_8799.n42 5.97853
R5819 a_n6308_8799.n41 a_n6308_8799.n10 77.6622
R5820 a_n6308_8799.n40 a_n6308_8799.n77 16.6962
R5821 a_n6308_8799.n40 a_n6308_8799.n12 72.3034
R5822 a_n6308_8799.n8 a_n6308_8799.n49 70.1674
R5823 a_n6308_8799.n87 a_n6308_8799.n49 20.9683
R5824 a_n6308_8799.n48 a_n6308_8799.n8 72.3034
R5825 a_n6308_8799.n48 a_n6308_8799.n81 16.6962
R5826 a_n6308_8799.n7 a_n6308_8799.n47 77.6622
R5827 a_n6308_8799.n86 a_n6308_8799.n47 5.97853
R5828 a_n6308_8799.n46 a_n6308_8799.n7 77.6622
R5829 a_n6308_8799.n45 a_n6308_8799.n84 16.6962
R5830 a_n6308_8799.n45 a_n6308_8799.n9 72.3034
R5831 a_n6308_8799.n5 a_n6308_8799.n54 70.1674
R5832 a_n6308_8799.n95 a_n6308_8799.n54 20.9683
R5833 a_n6308_8799.n53 a_n6308_8799.n5 72.3034
R5834 a_n6308_8799.n53 a_n6308_8799.n89 16.6962
R5835 a_n6308_8799.n4 a_n6308_8799.n52 77.6622
R5836 a_n6308_8799.n94 a_n6308_8799.n52 5.97853
R5837 a_n6308_8799.n51 a_n6308_8799.n4 77.6622
R5838 a_n6308_8799.n50 a_n6308_8799.n92 16.6962
R5839 a_n6308_8799.n50 a_n6308_8799.n6 72.3034
R5840 a_n6308_8799.n23 a_n6308_8799.n55 98.9633
R5841 a_n6308_8799.n22 a_n6308_8799.n57 98.9631
R5842 a_n6308_8799.n24 a_n6308_8799.n123 98.6055
R5843 a_n6308_8799.n23 a_n6308_8799.n56 98.6055
R5844 a_n6308_8799.n22 a_n6308_8799.n58 98.6055
R5845 a_n6308_8799.n22 a_n6308_8799.n59 98.6055
R5846 a_n6308_8799.n61 a_n6308_8799.n60 98.6055
R5847 a_n6308_8799.n124 a_n6308_8799.n24 98.6054
R5848 a_n6308_8799.n1 a_n6308_8799.n62 81.3764
R5849 a_n6308_8799.n3 a_n6308_8799.n68 81.3764
R5850 a_n6308_8799.n0 a_n6308_8799.n65 81.3764
R5851 a_n6308_8799.n2 a_n6308_8799.n71 80.9324
R5852 a_n6308_8799.n2 a_n6308_8799.n72 80.9324
R5853 a_n6308_8799.n1 a_n6308_8799.n73 80.9324
R5854 a_n6308_8799.n1 a_n6308_8799.n64 80.9324
R5855 a_n6308_8799.n1 a_n6308_8799.n63 80.9324
R5856 a_n6308_8799.n3 a_n6308_8799.n69 80.9324
R5857 a_n6308_8799.n0 a_n6308_8799.n70 80.9324
R5858 a_n6308_8799.n0 a_n6308_8799.n67 80.9324
R5859 a_n6308_8799.n0 a_n6308_8799.n66 80.9324
R5860 a_n6308_8799.n20 a_n6308_8799.n99 70.4033
R5861 a_n6308_8799.n17 a_n6308_8799.n106 70.4033
R5862 a_n6308_8799.n14 a_n6308_8799.n114 70.4033
R5863 a_n6308_8799.n75 a_n6308_8799.n12 70.4033
R5864 a_n6308_8799.n82 a_n6308_8799.n9 70.4033
R5865 a_n6308_8799.n90 a_n6308_8799.n6 70.4033
R5866 a_n6308_8799.n102 a_n6308_8799.n101 48.2005
R5867 a_n6308_8799.n109 a_n6308_8799.n108 48.2005
R5868 a_n6308_8799.n117 a_n6308_8799.n116 48.2005
R5869 a_n6308_8799.n79 a_n6308_8799.n78 48.2005
R5870 a_n6308_8799.t45 a_n6308_8799.n44 485.135
R5871 a_n6308_8799.n86 a_n6308_8799.n85 48.2005
R5872 a_n6308_8799.t50 a_n6308_8799.n49 485.135
R5873 a_n6308_8799.n94 a_n6308_8799.n93 48.2005
R5874 a_n6308_8799.t78 a_n6308_8799.n54 485.135
R5875 a_n6308_8799.n26 a_n6308_8799.n97 16.6962
R5876 a_n6308_8799.n100 a_n6308_8799.n29 27.6507
R5877 a_n6308_8799.n31 a_n6308_8799.n104 16.6962
R5878 a_n6308_8799.n107 a_n6308_8799.n34 27.6507
R5879 a_n6308_8799.n36 a_n6308_8799.n112 16.6962
R5880 a_n6308_8799.n115 a_n6308_8799.n39 27.6507
R5881 a_n6308_8799.n80 a_n6308_8799.n43 27.6507
R5882 a_n6308_8799.n87 a_n6308_8799.n48 27.6507
R5883 a_n6308_8799.n95 a_n6308_8799.n53 27.6507
R5884 a_n6308_8799.n27 a_n6308_8799.n97 41.7634
R5885 a_n6308_8799.n32 a_n6308_8799.n104 41.7634
R5886 a_n6308_8799.n37 a_n6308_8799.n112 41.7634
R5887 a_n6308_8799.n77 a_n6308_8799.n41 41.7634
R5888 a_n6308_8799.n84 a_n6308_8799.n46 41.7634
R5889 a_n6308_8799.n92 a_n6308_8799.n51 41.7634
R5890 a_n6308_8799.n2 a_n6308_8799.n0 33.4185
R5891 a_n6308_8799.n122 a_n6308_8799.n61 32.0088
R5892 a_n6308_8799.n100 a_n6308_8799.n99 20.9576
R5893 a_n6308_8799.n107 a_n6308_8799.n106 20.9576
R5894 a_n6308_8799.n115 a_n6308_8799.n114 20.9576
R5895 a_n6308_8799.n76 a_n6308_8799.n75 20.9576
R5896 a_n6308_8799.n83 a_n6308_8799.n82 20.9576
R5897 a_n6308_8799.n91 a_n6308_8799.n90 20.9576
R5898 a_n6308_8799.n24 a_n6308_8799.n122 18.5874
R5899 a_n6308_8799.n27 a_n6308_8799.n102 5.97853
R5900 a_n6308_8799.n28 a_n6308_8799.n98 41.7634
R5901 a_n6308_8799.n32 a_n6308_8799.n109 5.97853
R5902 a_n6308_8799.n33 a_n6308_8799.n105 41.7634
R5903 a_n6308_8799.n37 a_n6308_8799.n117 5.97853
R5904 a_n6308_8799.n38 a_n6308_8799.n113 41.7634
R5905 a_n6308_8799.n78 a_n6308_8799.n41 5.97853
R5906 a_n6308_8799.n74 a_n6308_8799.n42 41.7634
R5907 a_n6308_8799.n85 a_n6308_8799.n46 5.97853
R5908 a_n6308_8799.n81 a_n6308_8799.n47 41.7634
R5909 a_n6308_8799.n93 a_n6308_8799.n51 5.97853
R5910 a_n6308_8799.n89 a_n6308_8799.n52 41.7634
R5911 a_n6308_8799.n121 a_n6308_8799.n1 12.3339
R5912 a_n6308_8799.n122 a_n6308_8799.n121 11.4887
R5913 a_n6308_8799.n103 a_n6308_8799.n26 27.6507
R5914 a_n6308_8799.n110 a_n6308_8799.n31 27.6507
R5915 a_n6308_8799.n118 a_n6308_8799.n36 27.6507
R5916 a_n6308_8799.n40 a_n6308_8799.n76 27.6507
R5917 a_n6308_8799.n45 a_n6308_8799.n83 27.6507
R5918 a_n6308_8799.n50 a_n6308_8799.n91 27.6507
R5919 a_n6308_8799.n111 a_n6308_8799.n21 9.05164
R5920 a_n6308_8799.n88 a_n6308_8799.n11 9.05164
R5921 a_n6308_8799.n120 a_n6308_8799.n96 7.00615
R5922 a_n6308_8799.n120 a_n6308_8799.n119 6.58471
R5923 a_n6308_8799.n111 a_n6308_8799.n18 4.94368
R5924 a_n6308_8799.n119 a_n6308_8799.n15 4.94368
R5925 a_n6308_8799.n88 a_n6308_8799.n8 4.94368
R5926 a_n6308_8799.n96 a_n6308_8799.n5 4.94368
R5927 a_n6308_8799.n119 a_n6308_8799.n111 4.10845
R5928 a_n6308_8799.n96 a_n6308_8799.n88 4.10845
R5929 a_n6308_8799.n123 a_n6308_8799.t5 3.61217
R5930 a_n6308_8799.n123 a_n6308_8799.t15 3.61217
R5931 a_n6308_8799.n56 a_n6308_8799.t10 3.61217
R5932 a_n6308_8799.n56 a_n6308_8799.t7 3.61217
R5933 a_n6308_8799.n55 a_n6308_8799.t11 3.61217
R5934 a_n6308_8799.n55 a_n6308_8799.t4 3.61217
R5935 a_n6308_8799.n57 a_n6308_8799.t13 3.61217
R5936 a_n6308_8799.n57 a_n6308_8799.t1 3.61217
R5937 a_n6308_8799.n58 a_n6308_8799.t6 3.61217
R5938 a_n6308_8799.n58 a_n6308_8799.t12 3.61217
R5939 a_n6308_8799.n59 a_n6308_8799.t3 3.61217
R5940 a_n6308_8799.n59 a_n6308_8799.t9 3.61217
R5941 a_n6308_8799.n60 a_n6308_8799.t14 3.61217
R5942 a_n6308_8799.n60 a_n6308_8799.t2 3.61217
R5943 a_n6308_8799.t0 a_n6308_8799.n124 3.61217
R5944 a_n6308_8799.n124 a_n6308_8799.t8 3.61217
R5945 a_n6308_8799.n121 a_n6308_8799.n120 3.4105
R5946 a_n6308_8799.n71 a_n6308_8799.t26 2.82907
R5947 a_n6308_8799.n71 a_n6308_8799.t27 2.82907
R5948 a_n6308_8799.n72 a_n6308_8799.t25 2.82907
R5949 a_n6308_8799.n72 a_n6308_8799.t16 2.82907
R5950 a_n6308_8799.n73 a_n6308_8799.t29 2.82907
R5951 a_n6308_8799.n73 a_n6308_8799.t32 2.82907
R5952 a_n6308_8799.n64 a_n6308_8799.t31 2.82907
R5953 a_n6308_8799.n64 a_n6308_8799.t30 2.82907
R5954 a_n6308_8799.n63 a_n6308_8799.t23 2.82907
R5955 a_n6308_8799.n63 a_n6308_8799.t34 2.82907
R5956 a_n6308_8799.n62 a_n6308_8799.t35 2.82907
R5957 a_n6308_8799.n62 a_n6308_8799.t37 2.82907
R5958 a_n6308_8799.n68 a_n6308_8799.t28 2.82907
R5959 a_n6308_8799.n68 a_n6308_8799.t21 2.82907
R5960 a_n6308_8799.n69 a_n6308_8799.t33 2.82907
R5961 a_n6308_8799.n69 a_n6308_8799.t39 2.82907
R5962 a_n6308_8799.n70 a_n6308_8799.t18 2.82907
R5963 a_n6308_8799.n70 a_n6308_8799.t22 2.82907
R5964 a_n6308_8799.n67 a_n6308_8799.t38 2.82907
R5965 a_n6308_8799.n67 a_n6308_8799.t17 2.82907
R5966 a_n6308_8799.n66 a_n6308_8799.t24 2.82907
R5967 a_n6308_8799.n66 a_n6308_8799.t19 2.82907
R5968 a_n6308_8799.n65 a_n6308_8799.t20 2.82907
R5969 a_n6308_8799.n65 a_n6308_8799.t36 2.82907
R5970 a_n6308_8799.n1 a_n6308_8799.n2 1.77636
R5971 a_n6308_8799.n0 a_n6308_8799.n3 1.3324
R5972 a_n6308_8799.n20 a_n6308_8799.n19 1.13686
R5973 a_n6308_8799.n17 a_n6308_8799.n16 1.13686
R5974 a_n6308_8799.n14 a_n6308_8799.n13 1.13686
R5975 a_n6308_8799.n11 a_n6308_8799.n10 1.13686
R5976 a_n6308_8799.n8 a_n6308_8799.n7 1.13686
R5977 a_n6308_8799.n5 a_n6308_8799.n4 1.13686
R5978 a_n6308_8799.n24 a_n6308_8799.n23 0.716017
R5979 a_n6308_8799.n61 a_n6308_8799.n22 0.716017
R5980 a_n6308_8799.n4 a_n6308_8799.n6 0.568682
R5981 a_n6308_8799.n7 a_n6308_8799.n9 0.568682
R5982 a_n6308_8799.n10 a_n6308_8799.n12 0.568682
R5983 a_n6308_8799.n13 a_n6308_8799.n15 0.568682
R5984 a_n6308_8799.n16 a_n6308_8799.n18 0.568682
R5985 a_n6308_8799.n19 a_n6308_8799.n21 0.568682
R5986 CSoutput.n19 CSoutput.t97 184.661
R5987 CSoutput.n78 CSoutput.n77 165.8
R5988 CSoutput.n76 CSoutput.n0 165.8
R5989 CSoutput.n75 CSoutput.n74 165.8
R5990 CSoutput.n73 CSoutput.n72 165.8
R5991 CSoutput.n71 CSoutput.n2 165.8
R5992 CSoutput.n69 CSoutput.n68 165.8
R5993 CSoutput.n67 CSoutput.n3 165.8
R5994 CSoutput.n66 CSoutput.n65 165.8
R5995 CSoutput.n63 CSoutput.n4 165.8
R5996 CSoutput.n61 CSoutput.n60 165.8
R5997 CSoutput.n59 CSoutput.n5 165.8
R5998 CSoutput.n58 CSoutput.n57 165.8
R5999 CSoutput.n55 CSoutput.n6 165.8
R6000 CSoutput.n54 CSoutput.n53 165.8
R6001 CSoutput.n52 CSoutput.n51 165.8
R6002 CSoutput.n50 CSoutput.n8 165.8
R6003 CSoutput.n48 CSoutput.n47 165.8
R6004 CSoutput.n46 CSoutput.n9 165.8
R6005 CSoutput.n45 CSoutput.n44 165.8
R6006 CSoutput.n42 CSoutput.n10 165.8
R6007 CSoutput.n41 CSoutput.n40 165.8
R6008 CSoutput.n39 CSoutput.n38 165.8
R6009 CSoutput.n37 CSoutput.n12 165.8
R6010 CSoutput.n35 CSoutput.n34 165.8
R6011 CSoutput.n33 CSoutput.n13 165.8
R6012 CSoutput.n32 CSoutput.n31 165.8
R6013 CSoutput.n29 CSoutput.n14 165.8
R6014 CSoutput.n28 CSoutput.n27 165.8
R6015 CSoutput.n26 CSoutput.n25 165.8
R6016 CSoutput.n24 CSoutput.n16 165.8
R6017 CSoutput.n22 CSoutput.n21 165.8
R6018 CSoutput.n20 CSoutput.n17 165.8
R6019 CSoutput.n77 CSoutput.t100 162.194
R6020 CSoutput.n18 CSoutput.t99 120.501
R6021 CSoutput.n23 CSoutput.t110 120.501
R6022 CSoutput.n15 CSoutput.t107 120.501
R6023 CSoutput.n30 CSoutput.t101 120.501
R6024 CSoutput.n36 CSoutput.t112 120.501
R6025 CSoutput.n11 CSoutput.t114 120.501
R6026 CSoutput.n43 CSoutput.t103 120.501
R6027 CSoutput.n49 CSoutput.t115 120.501
R6028 CSoutput.n7 CSoutput.t117 120.501
R6029 CSoutput.n56 CSoutput.t111 120.501
R6030 CSoutput.n62 CSoutput.t102 120.501
R6031 CSoutput.n64 CSoutput.t96 120.501
R6032 CSoutput.n70 CSoutput.t113 120.501
R6033 CSoutput.n1 CSoutput.t108 120.501
R6034 CSoutput.n270 CSoutput.n268 103.469
R6035 CSoutput.n262 CSoutput.n260 103.469
R6036 CSoutput.n255 CSoutput.n253 103.469
R6037 CSoutput.n96 CSoutput.n94 103.469
R6038 CSoutput.n88 CSoutput.n86 103.469
R6039 CSoutput.n81 CSoutput.n79 103.469
R6040 CSoutput.n272 CSoutput.n271 103.111
R6041 CSoutput.n270 CSoutput.n269 103.111
R6042 CSoutput.n266 CSoutput.n265 103.111
R6043 CSoutput.n264 CSoutput.n263 103.111
R6044 CSoutput.n262 CSoutput.n261 103.111
R6045 CSoutput.n259 CSoutput.n258 103.111
R6046 CSoutput.n257 CSoutput.n256 103.111
R6047 CSoutput.n255 CSoutput.n254 103.111
R6048 CSoutput.n96 CSoutput.n95 103.111
R6049 CSoutput.n98 CSoutput.n97 103.111
R6050 CSoutput.n100 CSoutput.n99 103.111
R6051 CSoutput.n88 CSoutput.n87 103.111
R6052 CSoutput.n90 CSoutput.n89 103.111
R6053 CSoutput.n92 CSoutput.n91 103.111
R6054 CSoutput.n81 CSoutput.n80 103.111
R6055 CSoutput.n83 CSoutput.n82 103.111
R6056 CSoutput.n85 CSoutput.n84 103.111
R6057 CSoutput.n274 CSoutput.n273 103.111
R6058 CSoutput.n290 CSoutput.n288 81.5057
R6059 CSoutput.n279 CSoutput.n277 81.5057
R6060 CSoutput.n314 CSoutput.n312 81.5057
R6061 CSoutput.n303 CSoutput.n301 81.5057
R6062 CSoutput.n298 CSoutput.n297 80.9324
R6063 CSoutput.n296 CSoutput.n295 80.9324
R6064 CSoutput.n294 CSoutput.n293 80.9324
R6065 CSoutput.n292 CSoutput.n291 80.9324
R6066 CSoutput.n290 CSoutput.n289 80.9324
R6067 CSoutput.n287 CSoutput.n286 80.9324
R6068 CSoutput.n285 CSoutput.n284 80.9324
R6069 CSoutput.n283 CSoutput.n282 80.9324
R6070 CSoutput.n281 CSoutput.n280 80.9324
R6071 CSoutput.n279 CSoutput.n278 80.9324
R6072 CSoutput.n314 CSoutput.n313 80.9324
R6073 CSoutput.n316 CSoutput.n315 80.9324
R6074 CSoutput.n318 CSoutput.n317 80.9324
R6075 CSoutput.n320 CSoutput.n319 80.9324
R6076 CSoutput.n322 CSoutput.n321 80.9324
R6077 CSoutput.n303 CSoutput.n302 80.9324
R6078 CSoutput.n305 CSoutput.n304 80.9324
R6079 CSoutput.n307 CSoutput.n306 80.9324
R6080 CSoutput.n309 CSoutput.n308 80.9324
R6081 CSoutput.n311 CSoutput.n310 80.9324
R6082 CSoutput.n25 CSoutput.n24 48.1486
R6083 CSoutput.n69 CSoutput.n3 48.1486
R6084 CSoutput.n38 CSoutput.n37 48.1486
R6085 CSoutput.n42 CSoutput.n41 48.1486
R6086 CSoutput.n51 CSoutput.n50 48.1486
R6087 CSoutput.n55 CSoutput.n54 48.1486
R6088 CSoutput.n22 CSoutput.n17 46.462
R6089 CSoutput.n72 CSoutput.n71 46.462
R6090 CSoutput.n20 CSoutput.n19 44.9055
R6091 CSoutput.n29 CSoutput.n28 43.7635
R6092 CSoutput.n65 CSoutput.n63 43.7635
R6093 CSoutput.n35 CSoutput.n13 41.7396
R6094 CSoutput.n57 CSoutput.n5 41.7396
R6095 CSoutput.n44 CSoutput.n9 37.0171
R6096 CSoutput.n48 CSoutput.n9 37.0171
R6097 CSoutput.n76 CSoutput.n75 34.9932
R6098 CSoutput.n31 CSoutput.n13 32.2947
R6099 CSoutput.n61 CSoutput.n5 32.2947
R6100 CSoutput.n30 CSoutput.n29 29.6014
R6101 CSoutput.n63 CSoutput.n62 29.6014
R6102 CSoutput.n19 CSoutput.n18 28.4085
R6103 CSoutput.n18 CSoutput.n17 25.1176
R6104 CSoutput.n72 CSoutput.n1 25.1176
R6105 CSoutput.n43 CSoutput.n42 22.0922
R6106 CSoutput.n50 CSoutput.n49 22.0922
R6107 CSoutput.n77 CSoutput.n76 21.8586
R6108 CSoutput.n37 CSoutput.n36 18.9681
R6109 CSoutput.n56 CSoutput.n55 18.9681
R6110 CSoutput.n25 CSoutput.n15 17.6292
R6111 CSoutput.n64 CSoutput.n3 17.6292
R6112 CSoutput.n24 CSoutput.n23 15.844
R6113 CSoutput.n70 CSoutput.n69 15.844
R6114 CSoutput.n38 CSoutput.n11 14.5051
R6115 CSoutput.n54 CSoutput.n7 14.5051
R6116 CSoutput.n325 CSoutput.n78 11.6139
R6117 CSoutput.n41 CSoutput.n11 11.3811
R6118 CSoutput.n51 CSoutput.n7 11.3811
R6119 CSoutput.n23 CSoutput.n22 10.0422
R6120 CSoutput.n71 CSoutput.n70 10.0422
R6121 CSoutput.n267 CSoutput.n259 9.25285
R6122 CSoutput.n93 CSoutput.n85 9.25285
R6123 CSoutput.n299 CSoutput.n287 8.97993
R6124 CSoutput.n323 CSoutput.n311 8.97993
R6125 CSoutput.n300 CSoutput.n276 8.82427
R6126 CSoutput.n28 CSoutput.n15 8.25698
R6127 CSoutput.n65 CSoutput.n64 8.25698
R6128 CSoutput.n300 CSoutput.n299 7.89345
R6129 CSoutput.n324 CSoutput.n323 7.89345
R6130 CSoutput.n276 CSoutput.n275 7.12641
R6131 CSoutput.n102 CSoutput.n101 7.12641
R6132 CSoutput.n36 CSoutput.n35 6.91809
R6133 CSoutput.n57 CSoutput.n56 6.91809
R6134 CSoutput.n299 CSoutput.n298 5.25266
R6135 CSoutput.n323 CSoutput.n322 5.25266
R6136 CSoutput.n325 CSoutput.n102 5.23183
R6137 CSoutput.n275 CSoutput.n274 5.1449
R6138 CSoutput.n267 CSoutput.n266 5.1449
R6139 CSoutput.n101 CSoutput.n100 5.1449
R6140 CSoutput.n93 CSoutput.n92 5.1449
R6141 CSoutput.n193 CSoutput.n146 4.5005
R6142 CSoutput.n162 CSoutput.n146 4.5005
R6143 CSoutput.n157 CSoutput.n141 4.5005
R6144 CSoutput.n157 CSoutput.n143 4.5005
R6145 CSoutput.n157 CSoutput.n140 4.5005
R6146 CSoutput.n157 CSoutput.n144 4.5005
R6147 CSoutput.n157 CSoutput.n139 4.5005
R6148 CSoutput.n157 CSoutput.t104 4.5005
R6149 CSoutput.n157 CSoutput.n138 4.5005
R6150 CSoutput.n157 CSoutput.n145 4.5005
R6151 CSoutput.n157 CSoutput.n146 4.5005
R6152 CSoutput.n155 CSoutput.n141 4.5005
R6153 CSoutput.n155 CSoutput.n143 4.5005
R6154 CSoutput.n155 CSoutput.n140 4.5005
R6155 CSoutput.n155 CSoutput.n144 4.5005
R6156 CSoutput.n155 CSoutput.n139 4.5005
R6157 CSoutput.n155 CSoutput.t104 4.5005
R6158 CSoutput.n155 CSoutput.n138 4.5005
R6159 CSoutput.n155 CSoutput.n145 4.5005
R6160 CSoutput.n155 CSoutput.n146 4.5005
R6161 CSoutput.n154 CSoutput.n141 4.5005
R6162 CSoutput.n154 CSoutput.n143 4.5005
R6163 CSoutput.n154 CSoutput.n140 4.5005
R6164 CSoutput.n154 CSoutput.n144 4.5005
R6165 CSoutput.n154 CSoutput.n139 4.5005
R6166 CSoutput.n154 CSoutput.t104 4.5005
R6167 CSoutput.n154 CSoutput.n138 4.5005
R6168 CSoutput.n154 CSoutput.n145 4.5005
R6169 CSoutput.n154 CSoutput.n146 4.5005
R6170 CSoutput.n239 CSoutput.n141 4.5005
R6171 CSoutput.n239 CSoutput.n143 4.5005
R6172 CSoutput.n239 CSoutput.n140 4.5005
R6173 CSoutput.n239 CSoutput.n144 4.5005
R6174 CSoutput.n239 CSoutput.n139 4.5005
R6175 CSoutput.n239 CSoutput.t104 4.5005
R6176 CSoutput.n239 CSoutput.n138 4.5005
R6177 CSoutput.n239 CSoutput.n145 4.5005
R6178 CSoutput.n239 CSoutput.n146 4.5005
R6179 CSoutput.n237 CSoutput.n141 4.5005
R6180 CSoutput.n237 CSoutput.n143 4.5005
R6181 CSoutput.n237 CSoutput.n140 4.5005
R6182 CSoutput.n237 CSoutput.n144 4.5005
R6183 CSoutput.n237 CSoutput.n139 4.5005
R6184 CSoutput.n237 CSoutput.t104 4.5005
R6185 CSoutput.n237 CSoutput.n138 4.5005
R6186 CSoutput.n237 CSoutput.n145 4.5005
R6187 CSoutput.n235 CSoutput.n141 4.5005
R6188 CSoutput.n235 CSoutput.n143 4.5005
R6189 CSoutput.n235 CSoutput.n140 4.5005
R6190 CSoutput.n235 CSoutput.n144 4.5005
R6191 CSoutput.n235 CSoutput.n139 4.5005
R6192 CSoutput.n235 CSoutput.t104 4.5005
R6193 CSoutput.n235 CSoutput.n138 4.5005
R6194 CSoutput.n235 CSoutput.n145 4.5005
R6195 CSoutput.n165 CSoutput.n141 4.5005
R6196 CSoutput.n165 CSoutput.n143 4.5005
R6197 CSoutput.n165 CSoutput.n140 4.5005
R6198 CSoutput.n165 CSoutput.n144 4.5005
R6199 CSoutput.n165 CSoutput.n139 4.5005
R6200 CSoutput.n165 CSoutput.t104 4.5005
R6201 CSoutput.n165 CSoutput.n138 4.5005
R6202 CSoutput.n165 CSoutput.n145 4.5005
R6203 CSoutput.n165 CSoutput.n146 4.5005
R6204 CSoutput.n164 CSoutput.n141 4.5005
R6205 CSoutput.n164 CSoutput.n143 4.5005
R6206 CSoutput.n164 CSoutput.n140 4.5005
R6207 CSoutput.n164 CSoutput.n144 4.5005
R6208 CSoutput.n164 CSoutput.n139 4.5005
R6209 CSoutput.n164 CSoutput.t104 4.5005
R6210 CSoutput.n164 CSoutput.n138 4.5005
R6211 CSoutput.n164 CSoutput.n145 4.5005
R6212 CSoutput.n164 CSoutput.n146 4.5005
R6213 CSoutput.n168 CSoutput.n141 4.5005
R6214 CSoutput.n168 CSoutput.n143 4.5005
R6215 CSoutput.n168 CSoutput.n140 4.5005
R6216 CSoutput.n168 CSoutput.n144 4.5005
R6217 CSoutput.n168 CSoutput.n139 4.5005
R6218 CSoutput.n168 CSoutput.t104 4.5005
R6219 CSoutput.n168 CSoutput.n138 4.5005
R6220 CSoutput.n168 CSoutput.n145 4.5005
R6221 CSoutput.n168 CSoutput.n146 4.5005
R6222 CSoutput.n167 CSoutput.n141 4.5005
R6223 CSoutput.n167 CSoutput.n143 4.5005
R6224 CSoutput.n167 CSoutput.n140 4.5005
R6225 CSoutput.n167 CSoutput.n144 4.5005
R6226 CSoutput.n167 CSoutput.n139 4.5005
R6227 CSoutput.n167 CSoutput.t104 4.5005
R6228 CSoutput.n167 CSoutput.n138 4.5005
R6229 CSoutput.n167 CSoutput.n145 4.5005
R6230 CSoutput.n167 CSoutput.n146 4.5005
R6231 CSoutput.n150 CSoutput.n141 4.5005
R6232 CSoutput.n150 CSoutput.n143 4.5005
R6233 CSoutput.n150 CSoutput.n140 4.5005
R6234 CSoutput.n150 CSoutput.n144 4.5005
R6235 CSoutput.n150 CSoutput.n139 4.5005
R6236 CSoutput.n150 CSoutput.t104 4.5005
R6237 CSoutput.n150 CSoutput.n138 4.5005
R6238 CSoutput.n150 CSoutput.n145 4.5005
R6239 CSoutput.n150 CSoutput.n146 4.5005
R6240 CSoutput.n242 CSoutput.n141 4.5005
R6241 CSoutput.n242 CSoutput.n143 4.5005
R6242 CSoutput.n242 CSoutput.n140 4.5005
R6243 CSoutput.n242 CSoutput.n144 4.5005
R6244 CSoutput.n242 CSoutput.n139 4.5005
R6245 CSoutput.n242 CSoutput.t104 4.5005
R6246 CSoutput.n242 CSoutput.n138 4.5005
R6247 CSoutput.n242 CSoutput.n145 4.5005
R6248 CSoutput.n242 CSoutput.n146 4.5005
R6249 CSoutput.n229 CSoutput.n200 4.5005
R6250 CSoutput.n229 CSoutput.n206 4.5005
R6251 CSoutput.n187 CSoutput.n176 4.5005
R6252 CSoutput.n187 CSoutput.n178 4.5005
R6253 CSoutput.n187 CSoutput.n175 4.5005
R6254 CSoutput.n187 CSoutput.n179 4.5005
R6255 CSoutput.n187 CSoutput.n174 4.5005
R6256 CSoutput.n187 CSoutput.t98 4.5005
R6257 CSoutput.n187 CSoutput.n173 4.5005
R6258 CSoutput.n187 CSoutput.n180 4.5005
R6259 CSoutput.n229 CSoutput.n187 4.5005
R6260 CSoutput.n208 CSoutput.n176 4.5005
R6261 CSoutput.n208 CSoutput.n178 4.5005
R6262 CSoutput.n208 CSoutput.n175 4.5005
R6263 CSoutput.n208 CSoutput.n179 4.5005
R6264 CSoutput.n208 CSoutput.n174 4.5005
R6265 CSoutput.n208 CSoutput.t98 4.5005
R6266 CSoutput.n208 CSoutput.n173 4.5005
R6267 CSoutput.n208 CSoutput.n180 4.5005
R6268 CSoutput.n229 CSoutput.n208 4.5005
R6269 CSoutput.n186 CSoutput.n176 4.5005
R6270 CSoutput.n186 CSoutput.n178 4.5005
R6271 CSoutput.n186 CSoutput.n175 4.5005
R6272 CSoutput.n186 CSoutput.n179 4.5005
R6273 CSoutput.n186 CSoutput.n174 4.5005
R6274 CSoutput.n186 CSoutput.t98 4.5005
R6275 CSoutput.n186 CSoutput.n173 4.5005
R6276 CSoutput.n186 CSoutput.n180 4.5005
R6277 CSoutput.n229 CSoutput.n186 4.5005
R6278 CSoutput.n210 CSoutput.n176 4.5005
R6279 CSoutput.n210 CSoutput.n178 4.5005
R6280 CSoutput.n210 CSoutput.n175 4.5005
R6281 CSoutput.n210 CSoutput.n179 4.5005
R6282 CSoutput.n210 CSoutput.n174 4.5005
R6283 CSoutput.n210 CSoutput.t98 4.5005
R6284 CSoutput.n210 CSoutput.n173 4.5005
R6285 CSoutput.n210 CSoutput.n180 4.5005
R6286 CSoutput.n229 CSoutput.n210 4.5005
R6287 CSoutput.n176 CSoutput.n171 4.5005
R6288 CSoutput.n178 CSoutput.n171 4.5005
R6289 CSoutput.n175 CSoutput.n171 4.5005
R6290 CSoutput.n179 CSoutput.n171 4.5005
R6291 CSoutput.n174 CSoutput.n171 4.5005
R6292 CSoutput.t98 CSoutput.n171 4.5005
R6293 CSoutput.n173 CSoutput.n171 4.5005
R6294 CSoutput.n180 CSoutput.n171 4.5005
R6295 CSoutput.n232 CSoutput.n176 4.5005
R6296 CSoutput.n232 CSoutput.n178 4.5005
R6297 CSoutput.n232 CSoutput.n175 4.5005
R6298 CSoutput.n232 CSoutput.n179 4.5005
R6299 CSoutput.n232 CSoutput.n174 4.5005
R6300 CSoutput.n232 CSoutput.t98 4.5005
R6301 CSoutput.n232 CSoutput.n173 4.5005
R6302 CSoutput.n232 CSoutput.n180 4.5005
R6303 CSoutput.n230 CSoutput.n176 4.5005
R6304 CSoutput.n230 CSoutput.n178 4.5005
R6305 CSoutput.n230 CSoutput.n175 4.5005
R6306 CSoutput.n230 CSoutput.n179 4.5005
R6307 CSoutput.n230 CSoutput.n174 4.5005
R6308 CSoutput.n230 CSoutput.t98 4.5005
R6309 CSoutput.n230 CSoutput.n173 4.5005
R6310 CSoutput.n230 CSoutput.n180 4.5005
R6311 CSoutput.n230 CSoutput.n229 4.5005
R6312 CSoutput.n212 CSoutput.n176 4.5005
R6313 CSoutput.n212 CSoutput.n178 4.5005
R6314 CSoutput.n212 CSoutput.n175 4.5005
R6315 CSoutput.n212 CSoutput.n179 4.5005
R6316 CSoutput.n212 CSoutput.n174 4.5005
R6317 CSoutput.n212 CSoutput.t98 4.5005
R6318 CSoutput.n212 CSoutput.n173 4.5005
R6319 CSoutput.n212 CSoutput.n180 4.5005
R6320 CSoutput.n229 CSoutput.n212 4.5005
R6321 CSoutput.n184 CSoutput.n176 4.5005
R6322 CSoutput.n184 CSoutput.n178 4.5005
R6323 CSoutput.n184 CSoutput.n175 4.5005
R6324 CSoutput.n184 CSoutput.n179 4.5005
R6325 CSoutput.n184 CSoutput.n174 4.5005
R6326 CSoutput.n184 CSoutput.t98 4.5005
R6327 CSoutput.n184 CSoutput.n173 4.5005
R6328 CSoutput.n184 CSoutput.n180 4.5005
R6329 CSoutput.n229 CSoutput.n184 4.5005
R6330 CSoutput.n214 CSoutput.n176 4.5005
R6331 CSoutput.n214 CSoutput.n178 4.5005
R6332 CSoutput.n214 CSoutput.n175 4.5005
R6333 CSoutput.n214 CSoutput.n179 4.5005
R6334 CSoutput.n214 CSoutput.n174 4.5005
R6335 CSoutput.n214 CSoutput.t98 4.5005
R6336 CSoutput.n214 CSoutput.n173 4.5005
R6337 CSoutput.n214 CSoutput.n180 4.5005
R6338 CSoutput.n229 CSoutput.n214 4.5005
R6339 CSoutput.n183 CSoutput.n176 4.5005
R6340 CSoutput.n183 CSoutput.n178 4.5005
R6341 CSoutput.n183 CSoutput.n175 4.5005
R6342 CSoutput.n183 CSoutput.n179 4.5005
R6343 CSoutput.n183 CSoutput.n174 4.5005
R6344 CSoutput.n183 CSoutput.t98 4.5005
R6345 CSoutput.n183 CSoutput.n173 4.5005
R6346 CSoutput.n183 CSoutput.n180 4.5005
R6347 CSoutput.n229 CSoutput.n183 4.5005
R6348 CSoutput.n228 CSoutput.n176 4.5005
R6349 CSoutput.n228 CSoutput.n178 4.5005
R6350 CSoutput.n228 CSoutput.n175 4.5005
R6351 CSoutput.n228 CSoutput.n179 4.5005
R6352 CSoutput.n228 CSoutput.n174 4.5005
R6353 CSoutput.n228 CSoutput.t98 4.5005
R6354 CSoutput.n228 CSoutput.n173 4.5005
R6355 CSoutput.n228 CSoutput.n180 4.5005
R6356 CSoutput.n229 CSoutput.n228 4.5005
R6357 CSoutput.n227 CSoutput.n112 4.5005
R6358 CSoutput.n128 CSoutput.n112 4.5005
R6359 CSoutput.n123 CSoutput.n107 4.5005
R6360 CSoutput.n123 CSoutput.n109 4.5005
R6361 CSoutput.n123 CSoutput.n106 4.5005
R6362 CSoutput.n123 CSoutput.n110 4.5005
R6363 CSoutput.n123 CSoutput.n105 4.5005
R6364 CSoutput.n123 CSoutput.t116 4.5005
R6365 CSoutput.n123 CSoutput.n104 4.5005
R6366 CSoutput.n123 CSoutput.n111 4.5005
R6367 CSoutput.n123 CSoutput.n112 4.5005
R6368 CSoutput.n121 CSoutput.n107 4.5005
R6369 CSoutput.n121 CSoutput.n109 4.5005
R6370 CSoutput.n121 CSoutput.n106 4.5005
R6371 CSoutput.n121 CSoutput.n110 4.5005
R6372 CSoutput.n121 CSoutput.n105 4.5005
R6373 CSoutput.n121 CSoutput.t116 4.5005
R6374 CSoutput.n121 CSoutput.n104 4.5005
R6375 CSoutput.n121 CSoutput.n111 4.5005
R6376 CSoutput.n121 CSoutput.n112 4.5005
R6377 CSoutput.n120 CSoutput.n107 4.5005
R6378 CSoutput.n120 CSoutput.n109 4.5005
R6379 CSoutput.n120 CSoutput.n106 4.5005
R6380 CSoutput.n120 CSoutput.n110 4.5005
R6381 CSoutput.n120 CSoutput.n105 4.5005
R6382 CSoutput.n120 CSoutput.t116 4.5005
R6383 CSoutput.n120 CSoutput.n104 4.5005
R6384 CSoutput.n120 CSoutput.n111 4.5005
R6385 CSoutput.n120 CSoutput.n112 4.5005
R6386 CSoutput.n249 CSoutput.n107 4.5005
R6387 CSoutput.n249 CSoutput.n109 4.5005
R6388 CSoutput.n249 CSoutput.n106 4.5005
R6389 CSoutput.n249 CSoutput.n110 4.5005
R6390 CSoutput.n249 CSoutput.n105 4.5005
R6391 CSoutput.n249 CSoutput.t116 4.5005
R6392 CSoutput.n249 CSoutput.n104 4.5005
R6393 CSoutput.n249 CSoutput.n111 4.5005
R6394 CSoutput.n249 CSoutput.n112 4.5005
R6395 CSoutput.n247 CSoutput.n107 4.5005
R6396 CSoutput.n247 CSoutput.n109 4.5005
R6397 CSoutput.n247 CSoutput.n106 4.5005
R6398 CSoutput.n247 CSoutput.n110 4.5005
R6399 CSoutput.n247 CSoutput.n105 4.5005
R6400 CSoutput.n247 CSoutput.t116 4.5005
R6401 CSoutput.n247 CSoutput.n104 4.5005
R6402 CSoutput.n247 CSoutput.n111 4.5005
R6403 CSoutput.n245 CSoutput.n107 4.5005
R6404 CSoutput.n245 CSoutput.n109 4.5005
R6405 CSoutput.n245 CSoutput.n106 4.5005
R6406 CSoutput.n245 CSoutput.n110 4.5005
R6407 CSoutput.n245 CSoutput.n105 4.5005
R6408 CSoutput.n245 CSoutput.t116 4.5005
R6409 CSoutput.n245 CSoutput.n104 4.5005
R6410 CSoutput.n245 CSoutput.n111 4.5005
R6411 CSoutput.n131 CSoutput.n107 4.5005
R6412 CSoutput.n131 CSoutput.n109 4.5005
R6413 CSoutput.n131 CSoutput.n106 4.5005
R6414 CSoutput.n131 CSoutput.n110 4.5005
R6415 CSoutput.n131 CSoutput.n105 4.5005
R6416 CSoutput.n131 CSoutput.t116 4.5005
R6417 CSoutput.n131 CSoutput.n104 4.5005
R6418 CSoutput.n131 CSoutput.n111 4.5005
R6419 CSoutput.n131 CSoutput.n112 4.5005
R6420 CSoutput.n130 CSoutput.n107 4.5005
R6421 CSoutput.n130 CSoutput.n109 4.5005
R6422 CSoutput.n130 CSoutput.n106 4.5005
R6423 CSoutput.n130 CSoutput.n110 4.5005
R6424 CSoutput.n130 CSoutput.n105 4.5005
R6425 CSoutput.n130 CSoutput.t116 4.5005
R6426 CSoutput.n130 CSoutput.n104 4.5005
R6427 CSoutput.n130 CSoutput.n111 4.5005
R6428 CSoutput.n130 CSoutput.n112 4.5005
R6429 CSoutput.n134 CSoutput.n107 4.5005
R6430 CSoutput.n134 CSoutput.n109 4.5005
R6431 CSoutput.n134 CSoutput.n106 4.5005
R6432 CSoutput.n134 CSoutput.n110 4.5005
R6433 CSoutput.n134 CSoutput.n105 4.5005
R6434 CSoutput.n134 CSoutput.t116 4.5005
R6435 CSoutput.n134 CSoutput.n104 4.5005
R6436 CSoutput.n134 CSoutput.n111 4.5005
R6437 CSoutput.n134 CSoutput.n112 4.5005
R6438 CSoutput.n133 CSoutput.n107 4.5005
R6439 CSoutput.n133 CSoutput.n109 4.5005
R6440 CSoutput.n133 CSoutput.n106 4.5005
R6441 CSoutput.n133 CSoutput.n110 4.5005
R6442 CSoutput.n133 CSoutput.n105 4.5005
R6443 CSoutput.n133 CSoutput.t116 4.5005
R6444 CSoutput.n133 CSoutput.n104 4.5005
R6445 CSoutput.n133 CSoutput.n111 4.5005
R6446 CSoutput.n133 CSoutput.n112 4.5005
R6447 CSoutput.n116 CSoutput.n107 4.5005
R6448 CSoutput.n116 CSoutput.n109 4.5005
R6449 CSoutput.n116 CSoutput.n106 4.5005
R6450 CSoutput.n116 CSoutput.n110 4.5005
R6451 CSoutput.n116 CSoutput.n105 4.5005
R6452 CSoutput.n116 CSoutput.t116 4.5005
R6453 CSoutput.n116 CSoutput.n104 4.5005
R6454 CSoutput.n116 CSoutput.n111 4.5005
R6455 CSoutput.n116 CSoutput.n112 4.5005
R6456 CSoutput.n252 CSoutput.n107 4.5005
R6457 CSoutput.n252 CSoutput.n109 4.5005
R6458 CSoutput.n252 CSoutput.n106 4.5005
R6459 CSoutput.n252 CSoutput.n110 4.5005
R6460 CSoutput.n252 CSoutput.n105 4.5005
R6461 CSoutput.n252 CSoutput.t116 4.5005
R6462 CSoutput.n252 CSoutput.n104 4.5005
R6463 CSoutput.n252 CSoutput.n111 4.5005
R6464 CSoutput.n252 CSoutput.n112 4.5005
R6465 CSoutput.n275 CSoutput.n267 4.10845
R6466 CSoutput.n101 CSoutput.n93 4.10845
R6467 CSoutput.n273 CSoutput.t47 4.06363
R6468 CSoutput.n273 CSoutput.t49 4.06363
R6469 CSoutput.n271 CSoutput.t53 4.06363
R6470 CSoutput.n271 CSoutput.t75 4.06363
R6471 CSoutput.n269 CSoutput.t35 4.06363
R6472 CSoutput.n269 CSoutput.t52 4.06363
R6473 CSoutput.n268 CSoutput.t57 4.06363
R6474 CSoutput.n268 CSoutput.t67 4.06363
R6475 CSoutput.n265 CSoutput.t40 4.06363
R6476 CSoutput.n265 CSoutput.t41 4.06363
R6477 CSoutput.n263 CSoutput.t43 4.06363
R6478 CSoutput.n263 CSoutput.t70 4.06363
R6479 CSoutput.n261 CSoutput.t29 4.06363
R6480 CSoutput.n261 CSoutput.t42 4.06363
R6481 CSoutput.n260 CSoutput.t54 4.06363
R6482 CSoutput.n260 CSoutput.t61 4.06363
R6483 CSoutput.n258 CSoutput.t44 4.06363
R6484 CSoutput.n258 CSoutput.t34 4.06363
R6485 CSoutput.n256 CSoutput.t64 4.06363
R6486 CSoutput.n256 CSoutput.t31 4.06363
R6487 CSoutput.n254 CSoutput.t48 4.06363
R6488 CSoutput.n254 CSoutput.t74 4.06363
R6489 CSoutput.n253 CSoutput.t37 4.06363
R6490 CSoutput.n253 CSoutput.t69 4.06363
R6491 CSoutput.n94 CSoutput.t36 4.06363
R6492 CSoutput.n94 CSoutput.t71 4.06363
R6493 CSoutput.n95 CSoutput.t65 4.06363
R6494 CSoutput.n95 CSoutput.t56 4.06363
R6495 CSoutput.n97 CSoutput.t46 4.06363
R6496 CSoutput.n97 CSoutput.t76 4.06363
R6497 CSoutput.n99 CSoutput.t62 4.06363
R6498 CSoutput.n99 CSoutput.t63 4.06363
R6499 CSoutput.n86 CSoutput.t30 4.06363
R6500 CSoutput.n86 CSoutput.t66 4.06363
R6501 CSoutput.n87 CSoutput.t60 4.06363
R6502 CSoutput.n87 CSoutput.t51 4.06363
R6503 CSoutput.n89 CSoutput.t39 4.06363
R6504 CSoutput.n89 CSoutput.t72 4.06363
R6505 CSoutput.n91 CSoutput.t59 4.06363
R6506 CSoutput.n91 CSoutput.t58 4.06363
R6507 CSoutput.n79 CSoutput.t68 4.06363
R6508 CSoutput.n79 CSoutput.t38 4.06363
R6509 CSoutput.n80 CSoutput.t73 4.06363
R6510 CSoutput.n80 CSoutput.t50 4.06363
R6511 CSoutput.n82 CSoutput.t32 4.06363
R6512 CSoutput.n82 CSoutput.t55 4.06363
R6513 CSoutput.n84 CSoutput.t33 4.06363
R6514 CSoutput.n84 CSoutput.t45 4.06363
R6515 CSoutput.n44 CSoutput.n43 3.79402
R6516 CSoutput.n49 CSoutput.n48 3.79402
R6517 CSoutput.n325 CSoutput.n324 3.57343
R6518 CSoutput.n297 CSoutput.t17 2.82907
R6519 CSoutput.n297 CSoutput.t15 2.82907
R6520 CSoutput.n295 CSoutput.t87 2.82907
R6521 CSoutput.n295 CSoutput.t12 2.82907
R6522 CSoutput.n293 CSoutput.t14 2.82907
R6523 CSoutput.n293 CSoutput.t79 2.82907
R6524 CSoutput.n291 CSoutput.t10 2.82907
R6525 CSoutput.n291 CSoutput.t22 2.82907
R6526 CSoutput.n289 CSoutput.t9 2.82907
R6527 CSoutput.n289 CSoutput.t21 2.82907
R6528 CSoutput.n288 CSoutput.t86 2.82907
R6529 CSoutput.n288 CSoutput.t2 2.82907
R6530 CSoutput.n286 CSoutput.t90 2.82907
R6531 CSoutput.n286 CSoutput.t84 2.82907
R6532 CSoutput.n284 CSoutput.t77 2.82907
R6533 CSoutput.n284 CSoutput.t5 2.82907
R6534 CSoutput.n282 CSoutput.t93 2.82907
R6535 CSoutput.n282 CSoutput.t11 2.82907
R6536 CSoutput.n280 CSoutput.t28 2.82907
R6537 CSoutput.n280 CSoutput.t26 2.82907
R6538 CSoutput.n278 CSoutput.t27 2.82907
R6539 CSoutput.n278 CSoutput.t24 2.82907
R6540 CSoutput.n277 CSoutput.t19 2.82907
R6541 CSoutput.n277 CSoutput.t92 2.82907
R6542 CSoutput.n312 CSoutput.t78 2.82907
R6543 CSoutput.n312 CSoutput.t82 2.82907
R6544 CSoutput.n313 CSoutput.t3 2.82907
R6545 CSoutput.n313 CSoutput.t89 2.82907
R6546 CSoutput.n315 CSoutput.t0 2.82907
R6547 CSoutput.n315 CSoutput.t25 2.82907
R6548 CSoutput.n317 CSoutput.t18 2.82907
R6549 CSoutput.n317 CSoutput.t85 2.82907
R6550 CSoutput.n319 CSoutput.t95 2.82907
R6551 CSoutput.n319 CSoutput.t7 2.82907
R6552 CSoutput.n321 CSoutput.t23 2.82907
R6553 CSoutput.n321 CSoutput.t88 2.82907
R6554 CSoutput.n301 CSoutput.t16 2.82907
R6555 CSoutput.n301 CSoutput.t13 2.82907
R6556 CSoutput.n302 CSoutput.t20 2.82907
R6557 CSoutput.n302 CSoutput.t83 2.82907
R6558 CSoutput.n304 CSoutput.t1 2.82907
R6559 CSoutput.n304 CSoutput.t91 2.82907
R6560 CSoutput.n306 CSoutput.t80 2.82907
R6561 CSoutput.n306 CSoutput.t6 2.82907
R6562 CSoutput.n308 CSoutput.t81 2.82907
R6563 CSoutput.n308 CSoutput.t4 2.82907
R6564 CSoutput.n310 CSoutput.t8 2.82907
R6565 CSoutput.n310 CSoutput.t94 2.82907
R6566 CSoutput.n324 CSoutput.n300 2.75627
R6567 CSoutput.n75 CSoutput.n1 2.45513
R6568 CSoutput.n193 CSoutput.n191 2.251
R6569 CSoutput.n193 CSoutput.n190 2.251
R6570 CSoutput.n193 CSoutput.n189 2.251
R6571 CSoutput.n193 CSoutput.n188 2.251
R6572 CSoutput.n162 CSoutput.n161 2.251
R6573 CSoutput.n162 CSoutput.n160 2.251
R6574 CSoutput.n162 CSoutput.n159 2.251
R6575 CSoutput.n162 CSoutput.n158 2.251
R6576 CSoutput.n235 CSoutput.n234 2.251
R6577 CSoutput.n200 CSoutput.n198 2.251
R6578 CSoutput.n200 CSoutput.n197 2.251
R6579 CSoutput.n200 CSoutput.n196 2.251
R6580 CSoutput.n218 CSoutput.n200 2.251
R6581 CSoutput.n206 CSoutput.n205 2.251
R6582 CSoutput.n206 CSoutput.n204 2.251
R6583 CSoutput.n206 CSoutput.n203 2.251
R6584 CSoutput.n206 CSoutput.n202 2.251
R6585 CSoutput.n232 CSoutput.n172 2.251
R6586 CSoutput.n227 CSoutput.n225 2.251
R6587 CSoutput.n227 CSoutput.n224 2.251
R6588 CSoutput.n227 CSoutput.n223 2.251
R6589 CSoutput.n227 CSoutput.n222 2.251
R6590 CSoutput.n128 CSoutput.n127 2.251
R6591 CSoutput.n128 CSoutput.n126 2.251
R6592 CSoutput.n128 CSoutput.n125 2.251
R6593 CSoutput.n128 CSoutput.n124 2.251
R6594 CSoutput.n245 CSoutput.n244 2.251
R6595 CSoutput.n162 CSoutput.n142 2.2505
R6596 CSoutput.n157 CSoutput.n142 2.2505
R6597 CSoutput.n155 CSoutput.n142 2.2505
R6598 CSoutput.n154 CSoutput.n142 2.2505
R6599 CSoutput.n239 CSoutput.n142 2.2505
R6600 CSoutput.n237 CSoutput.n142 2.2505
R6601 CSoutput.n235 CSoutput.n142 2.2505
R6602 CSoutput.n165 CSoutput.n142 2.2505
R6603 CSoutput.n164 CSoutput.n142 2.2505
R6604 CSoutput.n168 CSoutput.n142 2.2505
R6605 CSoutput.n167 CSoutput.n142 2.2505
R6606 CSoutput.n150 CSoutput.n142 2.2505
R6607 CSoutput.n242 CSoutput.n142 2.2505
R6608 CSoutput.n242 CSoutput.n241 2.2505
R6609 CSoutput.n206 CSoutput.n177 2.2505
R6610 CSoutput.n187 CSoutput.n177 2.2505
R6611 CSoutput.n208 CSoutput.n177 2.2505
R6612 CSoutput.n186 CSoutput.n177 2.2505
R6613 CSoutput.n210 CSoutput.n177 2.2505
R6614 CSoutput.n177 CSoutput.n171 2.2505
R6615 CSoutput.n232 CSoutput.n177 2.2505
R6616 CSoutput.n230 CSoutput.n177 2.2505
R6617 CSoutput.n212 CSoutput.n177 2.2505
R6618 CSoutput.n184 CSoutput.n177 2.2505
R6619 CSoutput.n214 CSoutput.n177 2.2505
R6620 CSoutput.n183 CSoutput.n177 2.2505
R6621 CSoutput.n228 CSoutput.n177 2.2505
R6622 CSoutput.n228 CSoutput.n181 2.2505
R6623 CSoutput.n128 CSoutput.n108 2.2505
R6624 CSoutput.n123 CSoutput.n108 2.2505
R6625 CSoutput.n121 CSoutput.n108 2.2505
R6626 CSoutput.n120 CSoutput.n108 2.2505
R6627 CSoutput.n249 CSoutput.n108 2.2505
R6628 CSoutput.n247 CSoutput.n108 2.2505
R6629 CSoutput.n245 CSoutput.n108 2.2505
R6630 CSoutput.n131 CSoutput.n108 2.2505
R6631 CSoutput.n130 CSoutput.n108 2.2505
R6632 CSoutput.n134 CSoutput.n108 2.2505
R6633 CSoutput.n133 CSoutput.n108 2.2505
R6634 CSoutput.n116 CSoutput.n108 2.2505
R6635 CSoutput.n252 CSoutput.n108 2.2505
R6636 CSoutput.n252 CSoutput.n251 2.2505
R6637 CSoutput.n170 CSoutput.n163 2.25024
R6638 CSoutput.n170 CSoutput.n156 2.25024
R6639 CSoutput.n238 CSoutput.n170 2.25024
R6640 CSoutput.n170 CSoutput.n166 2.25024
R6641 CSoutput.n170 CSoutput.n169 2.25024
R6642 CSoutput.n170 CSoutput.n137 2.25024
R6643 CSoutput.n220 CSoutput.n217 2.25024
R6644 CSoutput.n220 CSoutput.n216 2.25024
R6645 CSoutput.n220 CSoutput.n215 2.25024
R6646 CSoutput.n220 CSoutput.n182 2.25024
R6647 CSoutput.n220 CSoutput.n219 2.25024
R6648 CSoutput.n221 CSoutput.n220 2.25024
R6649 CSoutput.n136 CSoutput.n129 2.25024
R6650 CSoutput.n136 CSoutput.n122 2.25024
R6651 CSoutput.n248 CSoutput.n136 2.25024
R6652 CSoutput.n136 CSoutput.n132 2.25024
R6653 CSoutput.n136 CSoutput.n135 2.25024
R6654 CSoutput.n136 CSoutput.n103 2.25024
R6655 CSoutput.n276 CSoutput.n102 2.15937
R6656 CSoutput.n237 CSoutput.n147 1.50111
R6657 CSoutput.n185 CSoutput.n171 1.50111
R6658 CSoutput.n247 CSoutput.n113 1.50111
R6659 CSoutput.n193 CSoutput.n192 1.501
R6660 CSoutput.n200 CSoutput.n199 1.501
R6661 CSoutput.n227 CSoutput.n226 1.501
R6662 CSoutput.n241 CSoutput.n152 1.12536
R6663 CSoutput.n241 CSoutput.n153 1.12536
R6664 CSoutput.n241 CSoutput.n240 1.12536
R6665 CSoutput.n201 CSoutput.n181 1.12536
R6666 CSoutput.n207 CSoutput.n181 1.12536
R6667 CSoutput.n209 CSoutput.n181 1.12536
R6668 CSoutput.n251 CSoutput.n118 1.12536
R6669 CSoutput.n251 CSoutput.n119 1.12536
R6670 CSoutput.n251 CSoutput.n250 1.12536
R6671 CSoutput.n241 CSoutput.n148 1.12536
R6672 CSoutput.n241 CSoutput.n149 1.12536
R6673 CSoutput.n241 CSoutput.n151 1.12536
R6674 CSoutput.n231 CSoutput.n181 1.12536
R6675 CSoutput.n211 CSoutput.n181 1.12536
R6676 CSoutput.n213 CSoutput.n181 1.12536
R6677 CSoutput.n251 CSoutput.n114 1.12536
R6678 CSoutput.n251 CSoutput.n115 1.12536
R6679 CSoutput.n251 CSoutput.n117 1.12536
R6680 CSoutput.n31 CSoutput.n30 0.669944
R6681 CSoutput.n62 CSoutput.n61 0.669944
R6682 CSoutput.n292 CSoutput.n290 0.573776
R6683 CSoutput.n294 CSoutput.n292 0.573776
R6684 CSoutput.n296 CSoutput.n294 0.573776
R6685 CSoutput.n298 CSoutput.n296 0.573776
R6686 CSoutput.n281 CSoutput.n279 0.573776
R6687 CSoutput.n283 CSoutput.n281 0.573776
R6688 CSoutput.n285 CSoutput.n283 0.573776
R6689 CSoutput.n287 CSoutput.n285 0.573776
R6690 CSoutput.n322 CSoutput.n320 0.573776
R6691 CSoutput.n320 CSoutput.n318 0.573776
R6692 CSoutput.n318 CSoutput.n316 0.573776
R6693 CSoutput.n316 CSoutput.n314 0.573776
R6694 CSoutput.n311 CSoutput.n309 0.573776
R6695 CSoutput.n309 CSoutput.n307 0.573776
R6696 CSoutput.n307 CSoutput.n305 0.573776
R6697 CSoutput.n305 CSoutput.n303 0.573776
R6698 CSoutput.n325 CSoutput.n252 0.53442
R6699 CSoutput.n272 CSoutput.n270 0.358259
R6700 CSoutput.n274 CSoutput.n272 0.358259
R6701 CSoutput.n264 CSoutput.n262 0.358259
R6702 CSoutput.n266 CSoutput.n264 0.358259
R6703 CSoutput.n257 CSoutput.n255 0.358259
R6704 CSoutput.n259 CSoutput.n257 0.358259
R6705 CSoutput.n100 CSoutput.n98 0.358259
R6706 CSoutput.n98 CSoutput.n96 0.358259
R6707 CSoutput.n92 CSoutput.n90 0.358259
R6708 CSoutput.n90 CSoutput.n88 0.358259
R6709 CSoutput.n85 CSoutput.n83 0.358259
R6710 CSoutput.n83 CSoutput.n81 0.358259
R6711 CSoutput.n21 CSoutput.n20 0.169105
R6712 CSoutput.n21 CSoutput.n16 0.169105
R6713 CSoutput.n26 CSoutput.n16 0.169105
R6714 CSoutput.n27 CSoutput.n26 0.169105
R6715 CSoutput.n27 CSoutput.n14 0.169105
R6716 CSoutput.n32 CSoutput.n14 0.169105
R6717 CSoutput.n33 CSoutput.n32 0.169105
R6718 CSoutput.n34 CSoutput.n33 0.169105
R6719 CSoutput.n34 CSoutput.n12 0.169105
R6720 CSoutput.n39 CSoutput.n12 0.169105
R6721 CSoutput.n40 CSoutput.n39 0.169105
R6722 CSoutput.n40 CSoutput.n10 0.169105
R6723 CSoutput.n45 CSoutput.n10 0.169105
R6724 CSoutput.n46 CSoutput.n45 0.169105
R6725 CSoutput.n47 CSoutput.n46 0.169105
R6726 CSoutput.n47 CSoutput.n8 0.169105
R6727 CSoutput.n52 CSoutput.n8 0.169105
R6728 CSoutput.n53 CSoutput.n52 0.169105
R6729 CSoutput.n53 CSoutput.n6 0.169105
R6730 CSoutput.n58 CSoutput.n6 0.169105
R6731 CSoutput.n59 CSoutput.n58 0.169105
R6732 CSoutput.n60 CSoutput.n59 0.169105
R6733 CSoutput.n60 CSoutput.n4 0.169105
R6734 CSoutput.n66 CSoutput.n4 0.169105
R6735 CSoutput.n67 CSoutput.n66 0.169105
R6736 CSoutput.n68 CSoutput.n67 0.169105
R6737 CSoutput.n68 CSoutput.n2 0.169105
R6738 CSoutput.n73 CSoutput.n2 0.169105
R6739 CSoutput.n74 CSoutput.n73 0.169105
R6740 CSoutput.n74 CSoutput.n0 0.169105
R6741 CSoutput.n78 CSoutput.n0 0.169105
R6742 CSoutput.n195 CSoutput.n194 0.0910737
R6743 CSoutput.n246 CSoutput.n243 0.0723685
R6744 CSoutput.n200 CSoutput.n195 0.0522944
R6745 CSoutput.n243 CSoutput.n242 0.0499135
R6746 CSoutput.n194 CSoutput.n193 0.0499135
R6747 CSoutput.n228 CSoutput.n227 0.0464294
R6748 CSoutput.n236 CSoutput.n233 0.0391444
R6749 CSoutput.n195 CSoutput.t106 0.023435
R6750 CSoutput.n243 CSoutput.t105 0.02262
R6751 CSoutput.n194 CSoutput.t109 0.02262
R6752 CSoutput CSoutput.n325 0.0052
R6753 CSoutput.n165 CSoutput.n148 0.00365111
R6754 CSoutput.n168 CSoutput.n149 0.00365111
R6755 CSoutput.n151 CSoutput.n150 0.00365111
R6756 CSoutput.n193 CSoutput.n152 0.00365111
R6757 CSoutput.n157 CSoutput.n153 0.00365111
R6758 CSoutput.n240 CSoutput.n154 0.00365111
R6759 CSoutput.n231 CSoutput.n230 0.00365111
R6760 CSoutput.n211 CSoutput.n184 0.00365111
R6761 CSoutput.n213 CSoutput.n183 0.00365111
R6762 CSoutput.n201 CSoutput.n200 0.00365111
R6763 CSoutput.n207 CSoutput.n187 0.00365111
R6764 CSoutput.n209 CSoutput.n186 0.00365111
R6765 CSoutput.n131 CSoutput.n114 0.00365111
R6766 CSoutput.n134 CSoutput.n115 0.00365111
R6767 CSoutput.n117 CSoutput.n116 0.00365111
R6768 CSoutput.n227 CSoutput.n118 0.00365111
R6769 CSoutput.n123 CSoutput.n119 0.00365111
R6770 CSoutput.n250 CSoutput.n120 0.00365111
R6771 CSoutput.n162 CSoutput.n152 0.00340054
R6772 CSoutput.n155 CSoutput.n153 0.00340054
R6773 CSoutput.n240 CSoutput.n239 0.00340054
R6774 CSoutput.n235 CSoutput.n148 0.00340054
R6775 CSoutput.n164 CSoutput.n149 0.00340054
R6776 CSoutput.n167 CSoutput.n151 0.00340054
R6777 CSoutput.n206 CSoutput.n201 0.00340054
R6778 CSoutput.n208 CSoutput.n207 0.00340054
R6779 CSoutput.n210 CSoutput.n209 0.00340054
R6780 CSoutput.n232 CSoutput.n231 0.00340054
R6781 CSoutput.n212 CSoutput.n211 0.00340054
R6782 CSoutput.n214 CSoutput.n213 0.00340054
R6783 CSoutput.n128 CSoutput.n118 0.00340054
R6784 CSoutput.n121 CSoutput.n119 0.00340054
R6785 CSoutput.n250 CSoutput.n249 0.00340054
R6786 CSoutput.n245 CSoutput.n114 0.00340054
R6787 CSoutput.n130 CSoutput.n115 0.00340054
R6788 CSoutput.n133 CSoutput.n117 0.00340054
R6789 CSoutput.n163 CSoutput.n157 0.00252698
R6790 CSoutput.n156 CSoutput.n154 0.00252698
R6791 CSoutput.n238 CSoutput.n237 0.00252698
R6792 CSoutput.n166 CSoutput.n164 0.00252698
R6793 CSoutput.n169 CSoutput.n167 0.00252698
R6794 CSoutput.n242 CSoutput.n137 0.00252698
R6795 CSoutput.n163 CSoutput.n162 0.00252698
R6796 CSoutput.n156 CSoutput.n155 0.00252698
R6797 CSoutput.n239 CSoutput.n238 0.00252698
R6798 CSoutput.n166 CSoutput.n165 0.00252698
R6799 CSoutput.n169 CSoutput.n168 0.00252698
R6800 CSoutput.n150 CSoutput.n137 0.00252698
R6801 CSoutput.n217 CSoutput.n187 0.00252698
R6802 CSoutput.n216 CSoutput.n186 0.00252698
R6803 CSoutput.n215 CSoutput.n171 0.00252698
R6804 CSoutput.n212 CSoutput.n182 0.00252698
R6805 CSoutput.n219 CSoutput.n214 0.00252698
R6806 CSoutput.n228 CSoutput.n221 0.00252698
R6807 CSoutput.n217 CSoutput.n206 0.00252698
R6808 CSoutput.n216 CSoutput.n208 0.00252698
R6809 CSoutput.n215 CSoutput.n210 0.00252698
R6810 CSoutput.n230 CSoutput.n182 0.00252698
R6811 CSoutput.n219 CSoutput.n184 0.00252698
R6812 CSoutput.n221 CSoutput.n183 0.00252698
R6813 CSoutput.n129 CSoutput.n123 0.00252698
R6814 CSoutput.n122 CSoutput.n120 0.00252698
R6815 CSoutput.n248 CSoutput.n247 0.00252698
R6816 CSoutput.n132 CSoutput.n130 0.00252698
R6817 CSoutput.n135 CSoutput.n133 0.00252698
R6818 CSoutput.n252 CSoutput.n103 0.00252698
R6819 CSoutput.n129 CSoutput.n128 0.00252698
R6820 CSoutput.n122 CSoutput.n121 0.00252698
R6821 CSoutput.n249 CSoutput.n248 0.00252698
R6822 CSoutput.n132 CSoutput.n131 0.00252698
R6823 CSoutput.n135 CSoutput.n134 0.00252698
R6824 CSoutput.n116 CSoutput.n103 0.00252698
R6825 CSoutput.n237 CSoutput.n236 0.0020275
R6826 CSoutput.n236 CSoutput.n235 0.0020275
R6827 CSoutput.n233 CSoutput.n171 0.0020275
R6828 CSoutput.n233 CSoutput.n232 0.0020275
R6829 CSoutput.n247 CSoutput.n246 0.0020275
R6830 CSoutput.n246 CSoutput.n245 0.0020275
R6831 CSoutput.n147 CSoutput.n146 0.00166668
R6832 CSoutput.n229 CSoutput.n185 0.00166668
R6833 CSoutput.n113 CSoutput.n112 0.00166668
R6834 CSoutput.n251 CSoutput.n113 0.00133328
R6835 CSoutput.n185 CSoutput.n181 0.00133328
R6836 CSoutput.n241 CSoutput.n147 0.00133328
R6837 CSoutput.n244 CSoutput.n136 0.001
R6838 CSoutput.n222 CSoutput.n136 0.001
R6839 CSoutput.n124 CSoutput.n104 0.001
R6840 CSoutput.n223 CSoutput.n104 0.001
R6841 CSoutput.n125 CSoutput.n105 0.001
R6842 CSoutput.n224 CSoutput.n105 0.001
R6843 CSoutput.n126 CSoutput.n106 0.001
R6844 CSoutput.n225 CSoutput.n106 0.001
R6845 CSoutput.n127 CSoutput.n107 0.001
R6846 CSoutput.n226 CSoutput.n107 0.001
R6847 CSoutput.n220 CSoutput.n172 0.001
R6848 CSoutput.n220 CSoutput.n218 0.001
R6849 CSoutput.n202 CSoutput.n173 0.001
R6850 CSoutput.n196 CSoutput.n173 0.001
R6851 CSoutput.n203 CSoutput.n174 0.001
R6852 CSoutput.n197 CSoutput.n174 0.001
R6853 CSoutput.n204 CSoutput.n175 0.001
R6854 CSoutput.n198 CSoutput.n175 0.001
R6855 CSoutput.n205 CSoutput.n176 0.001
R6856 CSoutput.n199 CSoutput.n176 0.001
R6857 CSoutput.n234 CSoutput.n170 0.001
R6858 CSoutput.n188 CSoutput.n170 0.001
R6859 CSoutput.n158 CSoutput.n138 0.001
R6860 CSoutput.n189 CSoutput.n138 0.001
R6861 CSoutput.n159 CSoutput.n139 0.001
R6862 CSoutput.n190 CSoutput.n139 0.001
R6863 CSoutput.n160 CSoutput.n140 0.001
R6864 CSoutput.n191 CSoutput.n140 0.001
R6865 CSoutput.n161 CSoutput.n141 0.001
R6866 CSoutput.n192 CSoutput.n141 0.001
R6867 CSoutput.n192 CSoutput.n142 0.001
R6868 CSoutput.n191 CSoutput.n143 0.001
R6869 CSoutput.n190 CSoutput.n144 0.001
R6870 CSoutput.n189 CSoutput.t104 0.001
R6871 CSoutput.n188 CSoutput.n145 0.001
R6872 CSoutput.n161 CSoutput.n143 0.001
R6873 CSoutput.n160 CSoutput.n144 0.001
R6874 CSoutput.n159 CSoutput.t104 0.001
R6875 CSoutput.n158 CSoutput.n145 0.001
R6876 CSoutput.n234 CSoutput.n146 0.001
R6877 CSoutput.n199 CSoutput.n177 0.001
R6878 CSoutput.n198 CSoutput.n178 0.001
R6879 CSoutput.n197 CSoutput.n179 0.001
R6880 CSoutput.n196 CSoutput.t98 0.001
R6881 CSoutput.n218 CSoutput.n180 0.001
R6882 CSoutput.n205 CSoutput.n178 0.001
R6883 CSoutput.n204 CSoutput.n179 0.001
R6884 CSoutput.n203 CSoutput.t98 0.001
R6885 CSoutput.n202 CSoutput.n180 0.001
R6886 CSoutput.n229 CSoutput.n172 0.001
R6887 CSoutput.n226 CSoutput.n108 0.001
R6888 CSoutput.n225 CSoutput.n109 0.001
R6889 CSoutput.n224 CSoutput.n110 0.001
R6890 CSoutput.n223 CSoutput.t116 0.001
R6891 CSoutput.n222 CSoutput.n111 0.001
R6892 CSoutput.n127 CSoutput.n109 0.001
R6893 CSoutput.n126 CSoutput.n110 0.001
R6894 CSoutput.n125 CSoutput.t116 0.001
R6895 CSoutput.n124 CSoutput.n111 0.001
R6896 CSoutput.n244 CSoutput.n112 0.001
R6897 gnd.n6424 gnd.n383 1323.14
R6898 gnd.n4483 gnd.n4482 939.716
R6899 gnd.n6719 gnd.n84 838.452
R6900 gnd.n6882 gnd.n80 838.452
R6901 gnd.n3552 gnd.n1214 838.452
R6902 gnd.n3471 gnd.n1216 838.452
R6903 gnd.n4276 gnd.n1083 838.452
R6904 gnd.n2158 gnd.n1081 838.452
R6905 gnd.n2271 gnd.n829 838.452
R6906 gnd.n2334 gnd.n2272 838.452
R6907 gnd.n6880 gnd.n86 819.232
R6908 gnd.n154 gnd.n82 819.232
R6909 gnd.n3883 gnd.n1213 819.232
R6910 gnd.n4129 gnd.n1217 819.232
R6911 gnd.n4278 gnd.n1078 819.232
R6912 gnd.n2669 gnd.n1080 819.232
R6913 gnd.n4404 gnd.n4403 819.232
R6914 gnd.n4480 gnd.n833 819.232
R6915 gnd.n2204 gnd.n1088 771.183
R6916 gnd.n4147 gnd.n1191 771.183
R6917 gnd.n2087 gnd.n2054 771.183
R6918 gnd.n3585 gnd.n1193 771.183
R6919 gnd.n5876 gnd.n798 766.379
R6920 gnd.n5792 gnd.n800 766.379
R6921 gnd.n4992 gnd.n4895 766.379
R6922 gnd.n4988 gnd.n4893 766.379
R6923 gnd.n5873 gnd.n4485 756.769
R6924 gnd.n5842 gnd.n801 756.769
R6925 gnd.n5159 gnd.n4802 756.769
R6926 gnd.n5157 gnd.n4805 756.769
R6927 gnd.n6066 gnd.n596 689.5
R6928 gnd.n6423 gnd.n384 689.5
R6929 gnd.n6637 gnd.n6635 689.5
R6930 gnd.n2463 gnd.n764 689.5
R6931 gnd.n599 gnd.n596 585
R6932 gnd.n6064 gnd.n596 585
R6933 gnd.n6062 gnd.n6061 585
R6934 gnd.n6063 gnd.n6062 585
R6935 gnd.n6060 gnd.n598 585
R6936 gnd.n598 gnd.n597 585
R6937 gnd.n6059 gnd.n6058 585
R6938 gnd.n6058 gnd.n6057 585
R6939 gnd.n604 gnd.n603 585
R6940 gnd.n6056 gnd.n604 585
R6941 gnd.n6054 gnd.n6053 585
R6942 gnd.n6055 gnd.n6054 585
R6943 gnd.n6052 gnd.n606 585
R6944 gnd.n606 gnd.n605 585
R6945 gnd.n6051 gnd.n6050 585
R6946 gnd.n6050 gnd.n6049 585
R6947 gnd.n612 gnd.n611 585
R6948 gnd.n6048 gnd.n612 585
R6949 gnd.n6046 gnd.n6045 585
R6950 gnd.n6047 gnd.n6046 585
R6951 gnd.n6044 gnd.n614 585
R6952 gnd.n614 gnd.n613 585
R6953 gnd.n6043 gnd.n6042 585
R6954 gnd.n6042 gnd.n6041 585
R6955 gnd.n620 gnd.n619 585
R6956 gnd.n6040 gnd.n620 585
R6957 gnd.n6038 gnd.n6037 585
R6958 gnd.n6039 gnd.n6038 585
R6959 gnd.n6036 gnd.n622 585
R6960 gnd.n622 gnd.n621 585
R6961 gnd.n6035 gnd.n6034 585
R6962 gnd.n6034 gnd.n6033 585
R6963 gnd.n628 gnd.n627 585
R6964 gnd.n6032 gnd.n628 585
R6965 gnd.n6030 gnd.n6029 585
R6966 gnd.n6031 gnd.n6030 585
R6967 gnd.n6028 gnd.n630 585
R6968 gnd.n630 gnd.n629 585
R6969 gnd.n6027 gnd.n6026 585
R6970 gnd.n6026 gnd.n6025 585
R6971 gnd.n636 gnd.n635 585
R6972 gnd.n6024 gnd.n636 585
R6973 gnd.n6022 gnd.n6021 585
R6974 gnd.n6023 gnd.n6022 585
R6975 gnd.n6020 gnd.n638 585
R6976 gnd.n638 gnd.n637 585
R6977 gnd.n6019 gnd.n6018 585
R6978 gnd.n6018 gnd.n6017 585
R6979 gnd.n644 gnd.n643 585
R6980 gnd.n6016 gnd.n644 585
R6981 gnd.n6014 gnd.n6013 585
R6982 gnd.n6015 gnd.n6014 585
R6983 gnd.n6012 gnd.n646 585
R6984 gnd.n646 gnd.n645 585
R6985 gnd.n6011 gnd.n6010 585
R6986 gnd.n6010 gnd.n6009 585
R6987 gnd.n652 gnd.n651 585
R6988 gnd.n6008 gnd.n652 585
R6989 gnd.n6006 gnd.n6005 585
R6990 gnd.n6007 gnd.n6006 585
R6991 gnd.n6004 gnd.n654 585
R6992 gnd.n654 gnd.n653 585
R6993 gnd.n6003 gnd.n6002 585
R6994 gnd.n6002 gnd.n6001 585
R6995 gnd.n660 gnd.n659 585
R6996 gnd.n6000 gnd.n660 585
R6997 gnd.n5998 gnd.n5997 585
R6998 gnd.n5999 gnd.n5998 585
R6999 gnd.n5996 gnd.n662 585
R7000 gnd.n662 gnd.n661 585
R7001 gnd.n5995 gnd.n5994 585
R7002 gnd.n5994 gnd.n5993 585
R7003 gnd.n668 gnd.n667 585
R7004 gnd.n5992 gnd.n668 585
R7005 gnd.n5990 gnd.n5989 585
R7006 gnd.n5991 gnd.n5990 585
R7007 gnd.n5988 gnd.n670 585
R7008 gnd.n670 gnd.n669 585
R7009 gnd.n5987 gnd.n5986 585
R7010 gnd.n5986 gnd.n5985 585
R7011 gnd.n676 gnd.n675 585
R7012 gnd.n5984 gnd.n676 585
R7013 gnd.n5982 gnd.n5981 585
R7014 gnd.n5983 gnd.n5982 585
R7015 gnd.n5980 gnd.n678 585
R7016 gnd.n678 gnd.n677 585
R7017 gnd.n5979 gnd.n5978 585
R7018 gnd.n5978 gnd.n5977 585
R7019 gnd.n684 gnd.n683 585
R7020 gnd.n5976 gnd.n684 585
R7021 gnd.n5974 gnd.n5973 585
R7022 gnd.n5975 gnd.n5974 585
R7023 gnd.n5972 gnd.n686 585
R7024 gnd.n686 gnd.n685 585
R7025 gnd.n5971 gnd.n5970 585
R7026 gnd.n5970 gnd.n5969 585
R7027 gnd.n692 gnd.n691 585
R7028 gnd.n5968 gnd.n692 585
R7029 gnd.n5966 gnd.n5965 585
R7030 gnd.n5967 gnd.n5966 585
R7031 gnd.n5964 gnd.n694 585
R7032 gnd.n694 gnd.n693 585
R7033 gnd.n5963 gnd.n5962 585
R7034 gnd.n5962 gnd.n5961 585
R7035 gnd.n700 gnd.n699 585
R7036 gnd.n5960 gnd.n700 585
R7037 gnd.n5958 gnd.n5957 585
R7038 gnd.n5959 gnd.n5958 585
R7039 gnd.n5956 gnd.n702 585
R7040 gnd.n702 gnd.n701 585
R7041 gnd.n5955 gnd.n5954 585
R7042 gnd.n5954 gnd.n5953 585
R7043 gnd.n708 gnd.n707 585
R7044 gnd.n5952 gnd.n708 585
R7045 gnd.n5950 gnd.n5949 585
R7046 gnd.n5951 gnd.n5950 585
R7047 gnd.n5948 gnd.n710 585
R7048 gnd.n710 gnd.n709 585
R7049 gnd.n5947 gnd.n5946 585
R7050 gnd.n5946 gnd.n5945 585
R7051 gnd.n716 gnd.n715 585
R7052 gnd.n5944 gnd.n716 585
R7053 gnd.n5942 gnd.n5941 585
R7054 gnd.n5943 gnd.n5942 585
R7055 gnd.n5940 gnd.n718 585
R7056 gnd.n718 gnd.n717 585
R7057 gnd.n5939 gnd.n5938 585
R7058 gnd.n5938 gnd.n5937 585
R7059 gnd.n724 gnd.n723 585
R7060 gnd.n5936 gnd.n724 585
R7061 gnd.n5934 gnd.n5933 585
R7062 gnd.n5935 gnd.n5934 585
R7063 gnd.n5932 gnd.n726 585
R7064 gnd.n726 gnd.n725 585
R7065 gnd.n5931 gnd.n5930 585
R7066 gnd.n5930 gnd.n5929 585
R7067 gnd.n732 gnd.n731 585
R7068 gnd.n5928 gnd.n732 585
R7069 gnd.n5926 gnd.n5925 585
R7070 gnd.n5927 gnd.n5926 585
R7071 gnd.n5924 gnd.n734 585
R7072 gnd.n734 gnd.n733 585
R7073 gnd.n5923 gnd.n5922 585
R7074 gnd.n5922 gnd.n5921 585
R7075 gnd.n740 gnd.n739 585
R7076 gnd.n5920 gnd.n740 585
R7077 gnd.n5918 gnd.n5917 585
R7078 gnd.n5919 gnd.n5918 585
R7079 gnd.n5916 gnd.n742 585
R7080 gnd.n742 gnd.n741 585
R7081 gnd.n5915 gnd.n5914 585
R7082 gnd.n5914 gnd.n5913 585
R7083 gnd.n748 gnd.n747 585
R7084 gnd.n5912 gnd.n748 585
R7085 gnd.n5910 gnd.n5909 585
R7086 gnd.n5911 gnd.n5910 585
R7087 gnd.n5908 gnd.n750 585
R7088 gnd.n750 gnd.n749 585
R7089 gnd.n5907 gnd.n5906 585
R7090 gnd.n5906 gnd.n5905 585
R7091 gnd.n756 gnd.n755 585
R7092 gnd.n5904 gnd.n756 585
R7093 gnd.n5902 gnd.n5901 585
R7094 gnd.n5903 gnd.n5902 585
R7095 gnd.n5900 gnd.n758 585
R7096 gnd.n758 gnd.n757 585
R7097 gnd.n5899 gnd.n5898 585
R7098 gnd.n5898 gnd.n5897 585
R7099 gnd.n6067 gnd.n6066 585
R7100 gnd.n6066 gnd.n6065 585
R7101 gnd.n594 gnd.n593 585
R7102 gnd.n593 gnd.n592 585
R7103 gnd.n6072 gnd.n6071 585
R7104 gnd.n6073 gnd.n6072 585
R7105 gnd.n591 gnd.n590 585
R7106 gnd.n6074 gnd.n591 585
R7107 gnd.n6077 gnd.n6076 585
R7108 gnd.n6076 gnd.n6075 585
R7109 gnd.n588 gnd.n587 585
R7110 gnd.n587 gnd.n586 585
R7111 gnd.n6082 gnd.n6081 585
R7112 gnd.n6083 gnd.n6082 585
R7113 gnd.n585 gnd.n584 585
R7114 gnd.n6084 gnd.n585 585
R7115 gnd.n6087 gnd.n6086 585
R7116 gnd.n6086 gnd.n6085 585
R7117 gnd.n582 gnd.n581 585
R7118 gnd.n581 gnd.n580 585
R7119 gnd.n6092 gnd.n6091 585
R7120 gnd.n6093 gnd.n6092 585
R7121 gnd.n579 gnd.n578 585
R7122 gnd.n6094 gnd.n579 585
R7123 gnd.n6097 gnd.n6096 585
R7124 gnd.n6096 gnd.n6095 585
R7125 gnd.n576 gnd.n575 585
R7126 gnd.n575 gnd.n574 585
R7127 gnd.n6102 gnd.n6101 585
R7128 gnd.n6103 gnd.n6102 585
R7129 gnd.n573 gnd.n572 585
R7130 gnd.n6104 gnd.n573 585
R7131 gnd.n6107 gnd.n6106 585
R7132 gnd.n6106 gnd.n6105 585
R7133 gnd.n570 gnd.n569 585
R7134 gnd.n569 gnd.n568 585
R7135 gnd.n6112 gnd.n6111 585
R7136 gnd.n6113 gnd.n6112 585
R7137 gnd.n567 gnd.n566 585
R7138 gnd.n6114 gnd.n567 585
R7139 gnd.n6117 gnd.n6116 585
R7140 gnd.n6116 gnd.n6115 585
R7141 gnd.n564 gnd.n563 585
R7142 gnd.n563 gnd.n562 585
R7143 gnd.n6122 gnd.n6121 585
R7144 gnd.n6123 gnd.n6122 585
R7145 gnd.n561 gnd.n560 585
R7146 gnd.n6124 gnd.n561 585
R7147 gnd.n6127 gnd.n6126 585
R7148 gnd.n6126 gnd.n6125 585
R7149 gnd.n558 gnd.n557 585
R7150 gnd.n557 gnd.n556 585
R7151 gnd.n6132 gnd.n6131 585
R7152 gnd.n6133 gnd.n6132 585
R7153 gnd.n555 gnd.n554 585
R7154 gnd.n6134 gnd.n555 585
R7155 gnd.n6137 gnd.n6136 585
R7156 gnd.n6136 gnd.n6135 585
R7157 gnd.n552 gnd.n551 585
R7158 gnd.n551 gnd.n550 585
R7159 gnd.n6142 gnd.n6141 585
R7160 gnd.n6143 gnd.n6142 585
R7161 gnd.n549 gnd.n548 585
R7162 gnd.n6144 gnd.n549 585
R7163 gnd.n6147 gnd.n6146 585
R7164 gnd.n6146 gnd.n6145 585
R7165 gnd.n546 gnd.n545 585
R7166 gnd.n545 gnd.n544 585
R7167 gnd.n6152 gnd.n6151 585
R7168 gnd.n6153 gnd.n6152 585
R7169 gnd.n543 gnd.n542 585
R7170 gnd.n6154 gnd.n543 585
R7171 gnd.n6157 gnd.n6156 585
R7172 gnd.n6156 gnd.n6155 585
R7173 gnd.n540 gnd.n539 585
R7174 gnd.n539 gnd.n538 585
R7175 gnd.n6162 gnd.n6161 585
R7176 gnd.n6163 gnd.n6162 585
R7177 gnd.n537 gnd.n536 585
R7178 gnd.n6164 gnd.n537 585
R7179 gnd.n6167 gnd.n6166 585
R7180 gnd.n6166 gnd.n6165 585
R7181 gnd.n534 gnd.n533 585
R7182 gnd.n533 gnd.n532 585
R7183 gnd.n6172 gnd.n6171 585
R7184 gnd.n6173 gnd.n6172 585
R7185 gnd.n531 gnd.n530 585
R7186 gnd.n6174 gnd.n531 585
R7187 gnd.n6177 gnd.n6176 585
R7188 gnd.n6176 gnd.n6175 585
R7189 gnd.n528 gnd.n527 585
R7190 gnd.n527 gnd.n526 585
R7191 gnd.n6182 gnd.n6181 585
R7192 gnd.n6183 gnd.n6182 585
R7193 gnd.n525 gnd.n524 585
R7194 gnd.n6184 gnd.n525 585
R7195 gnd.n6187 gnd.n6186 585
R7196 gnd.n6186 gnd.n6185 585
R7197 gnd.n522 gnd.n521 585
R7198 gnd.n521 gnd.n520 585
R7199 gnd.n6192 gnd.n6191 585
R7200 gnd.n6193 gnd.n6192 585
R7201 gnd.n519 gnd.n518 585
R7202 gnd.n6194 gnd.n519 585
R7203 gnd.n6197 gnd.n6196 585
R7204 gnd.n6196 gnd.n6195 585
R7205 gnd.n516 gnd.n515 585
R7206 gnd.n515 gnd.n514 585
R7207 gnd.n6202 gnd.n6201 585
R7208 gnd.n6203 gnd.n6202 585
R7209 gnd.n513 gnd.n512 585
R7210 gnd.n6204 gnd.n513 585
R7211 gnd.n6207 gnd.n6206 585
R7212 gnd.n6206 gnd.n6205 585
R7213 gnd.n510 gnd.n509 585
R7214 gnd.n509 gnd.n508 585
R7215 gnd.n6212 gnd.n6211 585
R7216 gnd.n6213 gnd.n6212 585
R7217 gnd.n507 gnd.n506 585
R7218 gnd.n6214 gnd.n507 585
R7219 gnd.n6217 gnd.n6216 585
R7220 gnd.n6216 gnd.n6215 585
R7221 gnd.n504 gnd.n503 585
R7222 gnd.n503 gnd.n502 585
R7223 gnd.n6222 gnd.n6221 585
R7224 gnd.n6223 gnd.n6222 585
R7225 gnd.n501 gnd.n500 585
R7226 gnd.n6224 gnd.n501 585
R7227 gnd.n6227 gnd.n6226 585
R7228 gnd.n6226 gnd.n6225 585
R7229 gnd.n498 gnd.n497 585
R7230 gnd.n497 gnd.n496 585
R7231 gnd.n6232 gnd.n6231 585
R7232 gnd.n6233 gnd.n6232 585
R7233 gnd.n495 gnd.n494 585
R7234 gnd.n6234 gnd.n495 585
R7235 gnd.n6237 gnd.n6236 585
R7236 gnd.n6236 gnd.n6235 585
R7237 gnd.n492 gnd.n491 585
R7238 gnd.n491 gnd.n490 585
R7239 gnd.n6242 gnd.n6241 585
R7240 gnd.n6243 gnd.n6242 585
R7241 gnd.n489 gnd.n488 585
R7242 gnd.n6244 gnd.n489 585
R7243 gnd.n6247 gnd.n6246 585
R7244 gnd.n6246 gnd.n6245 585
R7245 gnd.n486 gnd.n485 585
R7246 gnd.n485 gnd.n484 585
R7247 gnd.n6252 gnd.n6251 585
R7248 gnd.n6253 gnd.n6252 585
R7249 gnd.n483 gnd.n482 585
R7250 gnd.n6254 gnd.n483 585
R7251 gnd.n6257 gnd.n6256 585
R7252 gnd.n6256 gnd.n6255 585
R7253 gnd.n480 gnd.n479 585
R7254 gnd.n479 gnd.n478 585
R7255 gnd.n6262 gnd.n6261 585
R7256 gnd.n6263 gnd.n6262 585
R7257 gnd.n477 gnd.n476 585
R7258 gnd.n6264 gnd.n477 585
R7259 gnd.n6267 gnd.n6266 585
R7260 gnd.n6266 gnd.n6265 585
R7261 gnd.n474 gnd.n473 585
R7262 gnd.n473 gnd.n472 585
R7263 gnd.n6272 gnd.n6271 585
R7264 gnd.n6273 gnd.n6272 585
R7265 gnd.n471 gnd.n470 585
R7266 gnd.n6274 gnd.n471 585
R7267 gnd.n6277 gnd.n6276 585
R7268 gnd.n6276 gnd.n6275 585
R7269 gnd.n468 gnd.n467 585
R7270 gnd.n467 gnd.n466 585
R7271 gnd.n6282 gnd.n6281 585
R7272 gnd.n6283 gnd.n6282 585
R7273 gnd.n465 gnd.n464 585
R7274 gnd.n6284 gnd.n465 585
R7275 gnd.n6287 gnd.n6286 585
R7276 gnd.n6286 gnd.n6285 585
R7277 gnd.n462 gnd.n461 585
R7278 gnd.n461 gnd.n460 585
R7279 gnd.n6292 gnd.n6291 585
R7280 gnd.n6293 gnd.n6292 585
R7281 gnd.n459 gnd.n458 585
R7282 gnd.n6294 gnd.n459 585
R7283 gnd.n6297 gnd.n6296 585
R7284 gnd.n6296 gnd.n6295 585
R7285 gnd.n456 gnd.n455 585
R7286 gnd.n455 gnd.n454 585
R7287 gnd.n6302 gnd.n6301 585
R7288 gnd.n6303 gnd.n6302 585
R7289 gnd.n453 gnd.n452 585
R7290 gnd.n6304 gnd.n453 585
R7291 gnd.n6307 gnd.n6306 585
R7292 gnd.n6306 gnd.n6305 585
R7293 gnd.n450 gnd.n449 585
R7294 gnd.n449 gnd.n448 585
R7295 gnd.n6312 gnd.n6311 585
R7296 gnd.n6313 gnd.n6312 585
R7297 gnd.n447 gnd.n446 585
R7298 gnd.n6314 gnd.n447 585
R7299 gnd.n6317 gnd.n6316 585
R7300 gnd.n6316 gnd.n6315 585
R7301 gnd.n444 gnd.n443 585
R7302 gnd.n443 gnd.n442 585
R7303 gnd.n6322 gnd.n6321 585
R7304 gnd.n6323 gnd.n6322 585
R7305 gnd.n441 gnd.n440 585
R7306 gnd.n6324 gnd.n441 585
R7307 gnd.n6327 gnd.n6326 585
R7308 gnd.n6326 gnd.n6325 585
R7309 gnd.n438 gnd.n437 585
R7310 gnd.n437 gnd.n436 585
R7311 gnd.n6332 gnd.n6331 585
R7312 gnd.n6333 gnd.n6332 585
R7313 gnd.n435 gnd.n434 585
R7314 gnd.n6334 gnd.n435 585
R7315 gnd.n6337 gnd.n6336 585
R7316 gnd.n6336 gnd.n6335 585
R7317 gnd.n432 gnd.n431 585
R7318 gnd.n431 gnd.n430 585
R7319 gnd.n6342 gnd.n6341 585
R7320 gnd.n6343 gnd.n6342 585
R7321 gnd.n429 gnd.n428 585
R7322 gnd.n6344 gnd.n429 585
R7323 gnd.n6347 gnd.n6346 585
R7324 gnd.n6346 gnd.n6345 585
R7325 gnd.n426 gnd.n425 585
R7326 gnd.n425 gnd.n424 585
R7327 gnd.n6352 gnd.n6351 585
R7328 gnd.n6353 gnd.n6352 585
R7329 gnd.n423 gnd.n422 585
R7330 gnd.n6354 gnd.n423 585
R7331 gnd.n6357 gnd.n6356 585
R7332 gnd.n6356 gnd.n6355 585
R7333 gnd.n420 gnd.n419 585
R7334 gnd.n419 gnd.n418 585
R7335 gnd.n6362 gnd.n6361 585
R7336 gnd.n6363 gnd.n6362 585
R7337 gnd.n417 gnd.n416 585
R7338 gnd.n6364 gnd.n417 585
R7339 gnd.n6367 gnd.n6366 585
R7340 gnd.n6366 gnd.n6365 585
R7341 gnd.n414 gnd.n413 585
R7342 gnd.n413 gnd.n412 585
R7343 gnd.n6372 gnd.n6371 585
R7344 gnd.n6373 gnd.n6372 585
R7345 gnd.n411 gnd.n410 585
R7346 gnd.n6374 gnd.n411 585
R7347 gnd.n6377 gnd.n6376 585
R7348 gnd.n6376 gnd.n6375 585
R7349 gnd.n408 gnd.n407 585
R7350 gnd.n407 gnd.n406 585
R7351 gnd.n6382 gnd.n6381 585
R7352 gnd.n6383 gnd.n6382 585
R7353 gnd.n405 gnd.n404 585
R7354 gnd.n6384 gnd.n405 585
R7355 gnd.n6387 gnd.n6386 585
R7356 gnd.n6386 gnd.n6385 585
R7357 gnd.n402 gnd.n401 585
R7358 gnd.n401 gnd.n400 585
R7359 gnd.n6392 gnd.n6391 585
R7360 gnd.n6393 gnd.n6392 585
R7361 gnd.n399 gnd.n398 585
R7362 gnd.n6394 gnd.n399 585
R7363 gnd.n6397 gnd.n6396 585
R7364 gnd.n6396 gnd.n6395 585
R7365 gnd.n396 gnd.n395 585
R7366 gnd.n395 gnd.n394 585
R7367 gnd.n6402 gnd.n6401 585
R7368 gnd.n6403 gnd.n6402 585
R7369 gnd.n393 gnd.n392 585
R7370 gnd.n6404 gnd.n393 585
R7371 gnd.n6407 gnd.n6406 585
R7372 gnd.n6406 gnd.n6405 585
R7373 gnd.n390 gnd.n389 585
R7374 gnd.n389 gnd.n388 585
R7375 gnd.n6413 gnd.n6412 585
R7376 gnd.n6414 gnd.n6413 585
R7377 gnd.n387 gnd.n386 585
R7378 gnd.n6415 gnd.n387 585
R7379 gnd.n6418 gnd.n6417 585
R7380 gnd.n6417 gnd.n6416 585
R7381 gnd.n6419 gnd.n384 585
R7382 gnd.n384 gnd.n383 585
R7383 gnd.n259 gnd.n258 585
R7384 gnd.n6626 gnd.n258 585
R7385 gnd.n6629 gnd.n6628 585
R7386 gnd.n6628 gnd.n6627 585
R7387 gnd.n262 gnd.n261 585
R7388 gnd.n6625 gnd.n262 585
R7389 gnd.n6623 gnd.n6622 585
R7390 gnd.n6624 gnd.n6623 585
R7391 gnd.n265 gnd.n264 585
R7392 gnd.n264 gnd.n263 585
R7393 gnd.n6618 gnd.n6617 585
R7394 gnd.n6617 gnd.n6616 585
R7395 gnd.n268 gnd.n267 585
R7396 gnd.n6615 gnd.n268 585
R7397 gnd.n6613 gnd.n6612 585
R7398 gnd.n6614 gnd.n6613 585
R7399 gnd.n271 gnd.n270 585
R7400 gnd.n270 gnd.n269 585
R7401 gnd.n6608 gnd.n6607 585
R7402 gnd.n6607 gnd.n6606 585
R7403 gnd.n274 gnd.n273 585
R7404 gnd.n6605 gnd.n274 585
R7405 gnd.n6603 gnd.n6602 585
R7406 gnd.n6604 gnd.n6603 585
R7407 gnd.n277 gnd.n276 585
R7408 gnd.n276 gnd.n275 585
R7409 gnd.n6598 gnd.n6597 585
R7410 gnd.n6597 gnd.n6596 585
R7411 gnd.n280 gnd.n279 585
R7412 gnd.n6595 gnd.n280 585
R7413 gnd.n6593 gnd.n6592 585
R7414 gnd.n6594 gnd.n6593 585
R7415 gnd.n283 gnd.n282 585
R7416 gnd.n282 gnd.n281 585
R7417 gnd.n6588 gnd.n6587 585
R7418 gnd.n6587 gnd.n6586 585
R7419 gnd.n286 gnd.n285 585
R7420 gnd.n6585 gnd.n286 585
R7421 gnd.n6583 gnd.n6582 585
R7422 gnd.n6584 gnd.n6583 585
R7423 gnd.n289 gnd.n288 585
R7424 gnd.n288 gnd.n287 585
R7425 gnd.n6578 gnd.n6577 585
R7426 gnd.n6577 gnd.n6576 585
R7427 gnd.n292 gnd.n291 585
R7428 gnd.n6575 gnd.n292 585
R7429 gnd.n6573 gnd.n6572 585
R7430 gnd.n6574 gnd.n6573 585
R7431 gnd.n295 gnd.n294 585
R7432 gnd.n294 gnd.n293 585
R7433 gnd.n6568 gnd.n6567 585
R7434 gnd.n6567 gnd.n6566 585
R7435 gnd.n298 gnd.n297 585
R7436 gnd.n6565 gnd.n298 585
R7437 gnd.n6563 gnd.n6562 585
R7438 gnd.n6564 gnd.n6563 585
R7439 gnd.n301 gnd.n300 585
R7440 gnd.n300 gnd.n299 585
R7441 gnd.n6558 gnd.n6557 585
R7442 gnd.n6557 gnd.n6556 585
R7443 gnd.n304 gnd.n303 585
R7444 gnd.n6555 gnd.n304 585
R7445 gnd.n6553 gnd.n6552 585
R7446 gnd.n6554 gnd.n6553 585
R7447 gnd.n307 gnd.n306 585
R7448 gnd.n306 gnd.n305 585
R7449 gnd.n6548 gnd.n6547 585
R7450 gnd.n6547 gnd.n6546 585
R7451 gnd.n310 gnd.n309 585
R7452 gnd.n6545 gnd.n310 585
R7453 gnd.n6543 gnd.n6542 585
R7454 gnd.n6544 gnd.n6543 585
R7455 gnd.n313 gnd.n312 585
R7456 gnd.n312 gnd.n311 585
R7457 gnd.n6538 gnd.n6537 585
R7458 gnd.n6537 gnd.n6536 585
R7459 gnd.n316 gnd.n315 585
R7460 gnd.n6535 gnd.n316 585
R7461 gnd.n6533 gnd.n6532 585
R7462 gnd.n6534 gnd.n6533 585
R7463 gnd.n319 gnd.n318 585
R7464 gnd.n318 gnd.n317 585
R7465 gnd.n6528 gnd.n6527 585
R7466 gnd.n6527 gnd.n6526 585
R7467 gnd.n322 gnd.n321 585
R7468 gnd.n6525 gnd.n322 585
R7469 gnd.n6523 gnd.n6522 585
R7470 gnd.n6524 gnd.n6523 585
R7471 gnd.n325 gnd.n324 585
R7472 gnd.n324 gnd.n323 585
R7473 gnd.n6518 gnd.n6517 585
R7474 gnd.n6517 gnd.n6516 585
R7475 gnd.n328 gnd.n327 585
R7476 gnd.n6515 gnd.n328 585
R7477 gnd.n6513 gnd.n6512 585
R7478 gnd.n6514 gnd.n6513 585
R7479 gnd.n331 gnd.n330 585
R7480 gnd.n330 gnd.n329 585
R7481 gnd.n6508 gnd.n6507 585
R7482 gnd.n6507 gnd.n6506 585
R7483 gnd.n334 gnd.n333 585
R7484 gnd.n6505 gnd.n334 585
R7485 gnd.n6503 gnd.n6502 585
R7486 gnd.n6504 gnd.n6503 585
R7487 gnd.n337 gnd.n336 585
R7488 gnd.n336 gnd.n335 585
R7489 gnd.n6498 gnd.n6497 585
R7490 gnd.n6497 gnd.n6496 585
R7491 gnd.n340 gnd.n339 585
R7492 gnd.n6495 gnd.n340 585
R7493 gnd.n6493 gnd.n6492 585
R7494 gnd.n6494 gnd.n6493 585
R7495 gnd.n343 gnd.n342 585
R7496 gnd.n342 gnd.n341 585
R7497 gnd.n6488 gnd.n6487 585
R7498 gnd.n6487 gnd.n6486 585
R7499 gnd.n346 gnd.n345 585
R7500 gnd.n6485 gnd.n346 585
R7501 gnd.n6483 gnd.n6482 585
R7502 gnd.n6484 gnd.n6483 585
R7503 gnd.n349 gnd.n348 585
R7504 gnd.n348 gnd.n347 585
R7505 gnd.n6478 gnd.n6477 585
R7506 gnd.n6477 gnd.n6476 585
R7507 gnd.n352 gnd.n351 585
R7508 gnd.n6475 gnd.n352 585
R7509 gnd.n6473 gnd.n6472 585
R7510 gnd.n6474 gnd.n6473 585
R7511 gnd.n355 gnd.n354 585
R7512 gnd.n354 gnd.n353 585
R7513 gnd.n6468 gnd.n6467 585
R7514 gnd.n6467 gnd.n6466 585
R7515 gnd.n358 gnd.n357 585
R7516 gnd.n6465 gnd.n358 585
R7517 gnd.n6463 gnd.n6462 585
R7518 gnd.n6464 gnd.n6463 585
R7519 gnd.n361 gnd.n360 585
R7520 gnd.n360 gnd.n359 585
R7521 gnd.n6458 gnd.n6457 585
R7522 gnd.n6457 gnd.n6456 585
R7523 gnd.n364 gnd.n363 585
R7524 gnd.n6455 gnd.n364 585
R7525 gnd.n6453 gnd.n6452 585
R7526 gnd.n6454 gnd.n6453 585
R7527 gnd.n367 gnd.n366 585
R7528 gnd.n366 gnd.n365 585
R7529 gnd.n6448 gnd.n6447 585
R7530 gnd.n6447 gnd.n6446 585
R7531 gnd.n370 gnd.n369 585
R7532 gnd.n6445 gnd.n370 585
R7533 gnd.n6443 gnd.n6442 585
R7534 gnd.n6444 gnd.n6443 585
R7535 gnd.n373 gnd.n372 585
R7536 gnd.n372 gnd.n371 585
R7537 gnd.n6438 gnd.n6437 585
R7538 gnd.n6437 gnd.n6436 585
R7539 gnd.n376 gnd.n375 585
R7540 gnd.n6435 gnd.n376 585
R7541 gnd.n6433 gnd.n6432 585
R7542 gnd.n6434 gnd.n6433 585
R7543 gnd.n379 gnd.n378 585
R7544 gnd.n378 gnd.n377 585
R7545 gnd.n6428 gnd.n6427 585
R7546 gnd.n6427 gnd.n6426 585
R7547 gnd.n382 gnd.n381 585
R7548 gnd.n6425 gnd.n382 585
R7549 gnd.n6423 gnd.n6422 585
R7550 gnd.n6424 gnd.n6423 585
R7551 gnd.n4276 gnd.n4275 585
R7552 gnd.n4277 gnd.n4276 585
R7553 gnd.n1068 gnd.n1067 585
R7554 gnd.n2662 gnd.n1068 585
R7555 gnd.n4285 gnd.n4284 585
R7556 gnd.n4284 gnd.n4283 585
R7557 gnd.n4286 gnd.n1062 585
R7558 gnd.n2543 gnd.n1062 585
R7559 gnd.n4288 gnd.n4287 585
R7560 gnd.n4289 gnd.n4288 585
R7561 gnd.n1047 gnd.n1046 585
R7562 gnd.n2534 gnd.n1047 585
R7563 gnd.n4297 gnd.n4296 585
R7564 gnd.n4296 gnd.n4295 585
R7565 gnd.n4298 gnd.n1041 585
R7566 gnd.n2554 gnd.n1041 585
R7567 gnd.n4300 gnd.n4299 585
R7568 gnd.n4301 gnd.n4300 585
R7569 gnd.n1025 gnd.n1024 585
R7570 gnd.n2526 gnd.n1025 585
R7571 gnd.n4309 gnd.n4308 585
R7572 gnd.n4308 gnd.n4307 585
R7573 gnd.n4310 gnd.n1019 585
R7574 gnd.n2518 gnd.n1019 585
R7575 gnd.n4312 gnd.n4311 585
R7576 gnd.n4313 gnd.n4312 585
R7577 gnd.n1005 gnd.n1004 585
R7578 gnd.n2510 gnd.n1005 585
R7579 gnd.n4321 gnd.n4320 585
R7580 gnd.n4320 gnd.n4319 585
R7581 gnd.n4322 gnd.n999 585
R7582 gnd.n2502 gnd.n999 585
R7583 gnd.n4324 gnd.n4323 585
R7584 gnd.n4325 gnd.n4324 585
R7585 gnd.n986 gnd.n985 585
R7586 gnd.n2445 gnd.n986 585
R7587 gnd.n4334 gnd.n4333 585
R7588 gnd.n4333 gnd.n4332 585
R7589 gnd.n4335 gnd.n981 585
R7590 gnd.n2453 gnd.n981 585
R7591 gnd.n4337 gnd.n4336 585
R7592 gnd.n4338 gnd.n4337 585
R7593 gnd.n970 gnd.n969 585
R7594 gnd.n2431 gnd.n970 585
R7595 gnd.n4347 gnd.n4346 585
R7596 gnd.n4346 gnd.n4345 585
R7597 gnd.n4348 gnd.n962 585
R7598 gnd.n962 gnd.n960 585
R7599 gnd.n4350 gnd.n4349 585
R7600 gnd.n4351 gnd.n4350 585
R7601 gnd.n963 gnd.n961 585
R7602 gnd.n2420 gnd.n961 585
R7603 gnd.n946 gnd.n945 585
R7604 gnd.n949 gnd.n946 585
R7605 gnd.n4361 gnd.n4360 585
R7606 gnd.n4360 gnd.n4359 585
R7607 gnd.n4362 gnd.n940 585
R7608 gnd.n940 gnd.n939 585
R7609 gnd.n4364 gnd.n4363 585
R7610 gnd.n4365 gnd.n4364 585
R7611 gnd.n925 gnd.n924 585
R7612 gnd.n936 gnd.n925 585
R7613 gnd.n4373 gnd.n4372 585
R7614 gnd.n4372 gnd.n4371 585
R7615 gnd.n4374 gnd.n919 585
R7616 gnd.n926 gnd.n919 585
R7617 gnd.n4376 gnd.n4375 585
R7618 gnd.n4377 gnd.n4376 585
R7619 gnd.n906 gnd.n905 585
R7620 gnd.n909 gnd.n906 585
R7621 gnd.n4385 gnd.n4384 585
R7622 gnd.n4384 gnd.n4383 585
R7623 gnd.n4386 gnd.n900 585
R7624 gnd.n900 gnd.n898 585
R7625 gnd.n4388 gnd.n4387 585
R7626 gnd.n4389 gnd.n4388 585
R7627 gnd.n901 gnd.n899 585
R7628 gnd.n899 gnd.n886 585
R7629 gnd.n2339 gnd.n887 585
R7630 gnd.n4395 gnd.n887 585
R7631 gnd.n2275 gnd.n2273 585
R7632 gnd.n2273 gnd.n884 585
R7633 gnd.n2344 gnd.n2343 585
R7634 gnd.n2351 gnd.n2344 585
R7635 gnd.n2274 gnd.n2272 585
R7636 gnd.n2272 gnd.n830 585
R7637 gnd.n2335 gnd.n2334 585
R7638 gnd.n2333 gnd.n2332 585
R7639 gnd.n2331 gnd.n2330 585
R7640 gnd.n2329 gnd.n2328 585
R7641 gnd.n2327 gnd.n2326 585
R7642 gnd.n2325 gnd.n2324 585
R7643 gnd.n2323 gnd.n2322 585
R7644 gnd.n2321 gnd.n2320 585
R7645 gnd.n2319 gnd.n2318 585
R7646 gnd.n2317 gnd.n2316 585
R7647 gnd.n2315 gnd.n2314 585
R7648 gnd.n2313 gnd.n2312 585
R7649 gnd.n2311 gnd.n2310 585
R7650 gnd.n2309 gnd.n2308 585
R7651 gnd.n2307 gnd.n2306 585
R7652 gnd.n2305 gnd.n2304 585
R7653 gnd.n2303 gnd.n2302 585
R7654 gnd.n2294 gnd.n2291 585
R7655 gnd.n2298 gnd.n829 585
R7656 gnd.n4482 gnd.n829 585
R7657 gnd.n2159 gnd.n2158 585
R7658 gnd.n2156 gnd.n2150 585
R7659 gnd.n2166 gnd.n2147 585
R7660 gnd.n2167 gnd.n2145 585
R7661 gnd.n2144 gnd.n2137 585
R7662 gnd.n2174 gnd.n2136 585
R7663 gnd.n2175 gnd.n2135 585
R7664 gnd.n2133 gnd.n2125 585
R7665 gnd.n2182 gnd.n2124 585
R7666 gnd.n2183 gnd.n2122 585
R7667 gnd.n2121 gnd.n2114 585
R7668 gnd.n2190 gnd.n2113 585
R7669 gnd.n2191 gnd.n2112 585
R7670 gnd.n2110 gnd.n2103 585
R7671 gnd.n2198 gnd.n2102 585
R7672 gnd.n2199 gnd.n2100 585
R7673 gnd.n2099 gnd.n2095 585
R7674 gnd.n2097 gnd.n2096 585
R7675 gnd.n1085 gnd.n1083 585
R7676 gnd.n1996 gnd.n1083 585
R7677 gnd.n2032 gnd.n1081 585
R7678 gnd.n4277 gnd.n1081 585
R7679 gnd.n2661 gnd.n2660 585
R7680 gnd.n2662 gnd.n2661 585
R7681 gnd.n2031 gnd.n1071 585
R7682 gnd.n4283 gnd.n1071 585
R7683 gnd.n2546 gnd.n2544 585
R7684 gnd.n2544 gnd.n2543 585
R7685 gnd.n2547 gnd.n1060 585
R7686 gnd.n4289 gnd.n1060 585
R7687 gnd.n2548 gnd.n2226 585
R7688 gnd.n2534 gnd.n2226 585
R7689 gnd.n2223 gnd.n1049 585
R7690 gnd.n4295 gnd.n1049 585
R7691 gnd.n2553 gnd.n2552 585
R7692 gnd.n2554 gnd.n2553 585
R7693 gnd.n2222 gnd.n1039 585
R7694 gnd.n4301 gnd.n1039 585
R7695 gnd.n2525 gnd.n2524 585
R7696 gnd.n2526 gnd.n2525 585
R7697 gnd.n2232 gnd.n1028 585
R7698 gnd.n4307 gnd.n1028 585
R7699 gnd.n2520 gnd.n2519 585
R7700 gnd.n2519 gnd.n2518 585
R7701 gnd.n2234 gnd.n1018 585
R7702 gnd.n4313 gnd.n1018 585
R7703 gnd.n2509 gnd.n2508 585
R7704 gnd.n2510 gnd.n2509 585
R7705 gnd.n2239 gnd.n1007 585
R7706 gnd.n4319 gnd.n1007 585
R7707 gnd.n2504 gnd.n2503 585
R7708 gnd.n2503 gnd.n2502 585
R7709 gnd.n2241 gnd.n997 585
R7710 gnd.n4325 gnd.n997 585
R7711 gnd.n2447 gnd.n2446 585
R7712 gnd.n2446 gnd.n2445 585
R7713 gnd.n2250 gnd.n989 585
R7714 gnd.n4332 gnd.n989 585
R7715 gnd.n2452 gnd.n2451 585
R7716 gnd.n2453 gnd.n2452 585
R7717 gnd.n2249 gnd.n980 585
R7718 gnd.n4338 gnd.n980 585
R7719 gnd.n2430 gnd.n2429 585
R7720 gnd.n2431 gnd.n2430 585
R7721 gnd.n2257 gnd.n972 585
R7722 gnd.n4345 gnd.n972 585
R7723 gnd.n2425 gnd.n2424 585
R7724 gnd.n2424 gnd.n960 585
R7725 gnd.n2423 gnd.n959 585
R7726 gnd.n4351 gnd.n959 585
R7727 gnd.n2422 gnd.n2421 585
R7728 gnd.n2421 gnd.n2420 585
R7729 gnd.n2380 gnd.n2259 585
R7730 gnd.n2380 gnd.n949 585
R7731 gnd.n2376 gnd.n948 585
R7732 gnd.n4359 gnd.n948 585
R7733 gnd.n2375 gnd.n2374 585
R7734 gnd.n2374 gnd.n939 585
R7735 gnd.n2373 gnd.n938 585
R7736 gnd.n4365 gnd.n938 585
R7737 gnd.n2262 gnd.n2261 585
R7738 gnd.n2261 gnd.n936 585
R7739 gnd.n2369 gnd.n928 585
R7740 gnd.n4371 gnd.n928 585
R7741 gnd.n2368 gnd.n2367 585
R7742 gnd.n2367 gnd.n926 585
R7743 gnd.n2366 gnd.n918 585
R7744 gnd.n4377 gnd.n918 585
R7745 gnd.n2265 gnd.n2264 585
R7746 gnd.n2264 gnd.n909 585
R7747 gnd.n2362 gnd.n908 585
R7748 gnd.n4383 gnd.n908 585
R7749 gnd.n2361 gnd.n2360 585
R7750 gnd.n2360 gnd.n898 585
R7751 gnd.n2359 gnd.n897 585
R7752 gnd.n4389 gnd.n897 585
R7753 gnd.n2268 gnd.n2267 585
R7754 gnd.n2267 gnd.n886 585
R7755 gnd.n2355 gnd.n885 585
R7756 gnd.n4395 gnd.n885 585
R7757 gnd.n2354 gnd.n2353 585
R7758 gnd.n2353 gnd.n884 585
R7759 gnd.n2352 gnd.n2270 585
R7760 gnd.n2352 gnd.n2351 585
R7761 gnd.n2296 gnd.n2271 585
R7762 gnd.n2271 gnd.n830 585
R7763 gnd.n6785 gnd.n84 585
R7764 gnd.n6881 gnd.n84 585
R7765 gnd.n6786 gnd.n6717 585
R7766 gnd.n6717 gnd.n81 585
R7767 gnd.n6787 gnd.n163 585
R7768 gnd.n6801 gnd.n163 585
R7769 gnd.n175 gnd.n173 585
R7770 gnd.n173 gnd.n161 585
R7771 gnd.n6792 gnd.n6791 585
R7772 gnd.n6793 gnd.n6792 585
R7773 gnd.n174 gnd.n172 585
R7774 gnd.n172 gnd.n170 585
R7775 gnd.n6713 gnd.n6712 585
R7776 gnd.n6712 gnd.n6711 585
R7777 gnd.n178 gnd.n177 585
R7778 gnd.n188 gnd.n178 585
R7779 gnd.n6702 gnd.n6701 585
R7780 gnd.n6703 gnd.n6702 585
R7781 gnd.n190 gnd.n189 585
R7782 gnd.n189 gnd.n186 585
R7783 gnd.n6697 gnd.n6696 585
R7784 gnd.n6696 gnd.n6695 585
R7785 gnd.n193 gnd.n192 585
R7786 gnd.n194 gnd.n193 585
R7787 gnd.n6686 gnd.n6685 585
R7788 gnd.n6687 gnd.n6686 585
R7789 gnd.n205 gnd.n204 585
R7790 gnd.n204 gnd.n202 585
R7791 gnd.n6681 gnd.n6680 585
R7792 gnd.n6680 gnd.n6679 585
R7793 gnd.n208 gnd.n207 585
R7794 gnd.n224 gnd.n208 585
R7795 gnd.n6670 gnd.n6669 585
R7796 gnd.n6671 gnd.n6670 585
R7797 gnd.n226 gnd.n225 585
R7798 gnd.n225 gnd.n222 585
R7799 gnd.n6665 gnd.n6664 585
R7800 gnd.n6664 gnd.n6663 585
R7801 gnd.n229 gnd.n228 585
R7802 gnd.n230 gnd.n229 585
R7803 gnd.n6656 gnd.n6655 585
R7804 gnd.n6657 gnd.n6656 585
R7805 gnd.n239 gnd.n238 585
R7806 gnd.n3966 gnd.n238 585
R7807 gnd.n6651 gnd.n6650 585
R7808 gnd.n6650 gnd.n6649 585
R7809 gnd.n243 gnd.n242 585
R7810 gnd.n6644 gnd.n243 585
R7811 gnd.n4098 gnd.n4096 585
R7812 gnd.n4096 gnd.n4095 585
R7813 gnd.n4099 gnd.n1250 585
R7814 gnd.n3972 gnd.n1250 585
R7815 gnd.n4100 gnd.n1249 585
R7816 gnd.n4086 gnd.n1249 585
R7817 gnd.n1273 gnd.n1247 585
R7818 gnd.n1274 gnd.n1273 585
R7819 gnd.n4104 gnd.n1246 585
R7820 gnd.n4080 gnd.n1246 585
R7821 gnd.n4105 gnd.n1245 585
R7822 gnd.n4061 gnd.n1245 585
R7823 gnd.n4106 gnd.n1244 585
R7824 gnd.n1281 gnd.n1244 585
R7825 gnd.n1292 gnd.n1242 585
R7826 gnd.n4052 gnd.n1292 585
R7827 gnd.n4110 gnd.n1241 585
R7828 gnd.n1302 gnd.n1241 585
R7829 gnd.n4111 gnd.n1240 585
R7830 gnd.n4041 gnd.n1240 585
R7831 gnd.n4112 gnd.n1239 585
R7832 gnd.n4029 gnd.n1239 585
R7833 gnd.n1309 gnd.n1237 585
R7834 gnd.n1310 gnd.n1309 585
R7835 gnd.n4116 gnd.n1236 585
R7836 gnd.n4020 gnd.n1236 585
R7837 gnd.n4117 gnd.n1235 585
R7838 gnd.n3992 gnd.n1235 585
R7839 gnd.n4118 gnd.n1234 585
R7840 gnd.n4010 gnd.n1234 585
R7841 gnd.n1231 gnd.n1229 585
R7842 gnd.n3899 gnd.n1229 585
R7843 gnd.n4123 gnd.n4122 585
R7844 gnd.n4124 gnd.n4123 585
R7845 gnd.n1230 gnd.n1228 585
R7846 gnd.n3890 gnd.n1228 585
R7847 gnd.n3467 gnd.n1216 585
R7848 gnd.n4130 gnd.n1216 585
R7849 gnd.n3471 gnd.n3470 585
R7850 gnd.n3473 gnd.n3464 585
R7851 gnd.n3476 gnd.n3475 585
R7852 gnd.n3457 gnd.n3456 585
R7853 gnd.n3490 gnd.n3489 585
R7854 gnd.n3492 gnd.n3455 585
R7855 gnd.n3495 gnd.n3494 585
R7856 gnd.n3448 gnd.n3447 585
R7857 gnd.n3509 gnd.n3508 585
R7858 gnd.n3511 gnd.n3446 585
R7859 gnd.n3514 gnd.n3513 585
R7860 gnd.n3439 gnd.n3438 585
R7861 gnd.n3528 gnd.n3527 585
R7862 gnd.n3530 gnd.n3437 585
R7863 gnd.n3533 gnd.n3532 585
R7864 gnd.n3430 gnd.n3429 585
R7865 gnd.n3549 gnd.n3548 585
R7866 gnd.n3551 gnd.n3428 585
R7867 gnd.n3553 gnd.n3552 585
R7868 gnd.n3552 gnd.n1204 585
R7869 gnd.n6756 gnd.n80 585
R7870 gnd.n6757 gnd.n6755 585
R7871 gnd.n6758 gnd.n6751 585
R7872 gnd.n6749 gnd.n6747 585
R7873 gnd.n6762 gnd.n6746 585
R7874 gnd.n6763 gnd.n6744 585
R7875 gnd.n6764 gnd.n6743 585
R7876 gnd.n6741 gnd.n6739 585
R7877 gnd.n6768 gnd.n6738 585
R7878 gnd.n6769 gnd.n6736 585
R7879 gnd.n6770 gnd.n6735 585
R7880 gnd.n6733 gnd.n6731 585
R7881 gnd.n6774 gnd.n6730 585
R7882 gnd.n6775 gnd.n6728 585
R7883 gnd.n6776 gnd.n6727 585
R7884 gnd.n6725 gnd.n6723 585
R7885 gnd.n6780 gnd.n6722 585
R7886 gnd.n6781 gnd.n6720 585
R7887 gnd.n6782 gnd.n6719 585
R7888 gnd.n6719 gnd.n83 585
R7889 gnd.n6883 gnd.n6882 585
R7890 gnd.n6882 gnd.n6881 585
R7891 gnd.n79 gnd.n77 585
R7892 gnd.n81 gnd.n79 585
R7893 gnd.n6887 gnd.n76 585
R7894 gnd.n6801 gnd.n76 585
R7895 gnd.n6888 gnd.n75 585
R7896 gnd.n161 gnd.n75 585
R7897 gnd.n6889 gnd.n74 585
R7898 gnd.n6793 gnd.n74 585
R7899 gnd.n169 gnd.n72 585
R7900 gnd.n170 gnd.n169 585
R7901 gnd.n6893 gnd.n71 585
R7902 gnd.n6711 gnd.n71 585
R7903 gnd.n6894 gnd.n70 585
R7904 gnd.n188 gnd.n70 585
R7905 gnd.n6895 gnd.n69 585
R7906 gnd.n6703 gnd.n69 585
R7907 gnd.n185 gnd.n67 585
R7908 gnd.n186 gnd.n185 585
R7909 gnd.n6899 gnd.n66 585
R7910 gnd.n6695 gnd.n66 585
R7911 gnd.n6900 gnd.n65 585
R7912 gnd.n194 gnd.n65 585
R7913 gnd.n6901 gnd.n64 585
R7914 gnd.n6687 gnd.n64 585
R7915 gnd.n201 gnd.n62 585
R7916 gnd.n202 gnd.n201 585
R7917 gnd.n6905 gnd.n61 585
R7918 gnd.n6679 gnd.n61 585
R7919 gnd.n6906 gnd.n60 585
R7920 gnd.n224 gnd.n60 585
R7921 gnd.n6907 gnd.n59 585
R7922 gnd.n6671 gnd.n59 585
R7923 gnd.n221 gnd.n57 585
R7924 gnd.n222 gnd.n221 585
R7925 gnd.n6911 gnd.n56 585
R7926 gnd.n6663 gnd.n56 585
R7927 gnd.n6912 gnd.n55 585
R7928 gnd.n230 gnd.n55 585
R7929 gnd.n6913 gnd.n54 585
R7930 gnd.n6657 gnd.n54 585
R7931 gnd.n3965 gnd.n52 585
R7932 gnd.n3966 gnd.n3965 585
R7933 gnd.n1255 gnd.n245 585
R7934 gnd.n6649 gnd.n245 585
R7935 gnd.n1256 gnd.n250 585
R7936 gnd.n6644 gnd.n250 585
R7937 gnd.n4094 gnd.n4093 585
R7938 gnd.n4095 gnd.n4094 585
R7939 gnd.n1254 gnd.n1253 585
R7940 gnd.n3972 gnd.n1253 585
R7941 gnd.n4088 gnd.n4087 585
R7942 gnd.n4087 gnd.n4086 585
R7943 gnd.n1259 gnd.n1258 585
R7944 gnd.n1274 gnd.n1259 585
R7945 gnd.n1285 gnd.n1272 585
R7946 gnd.n4080 gnd.n1272 585
R7947 gnd.n4060 gnd.n4059 585
R7948 gnd.n4061 gnd.n4060 585
R7949 gnd.n1284 gnd.n1283 585
R7950 gnd.n1283 gnd.n1281 585
R7951 gnd.n4054 gnd.n4053 585
R7952 gnd.n4053 gnd.n4052 585
R7953 gnd.n1288 gnd.n1287 585
R7954 gnd.n1302 gnd.n1288 585
R7955 gnd.n1314 gnd.n1301 585
R7956 gnd.n4041 gnd.n1301 585
R7957 gnd.n4028 gnd.n4027 585
R7958 gnd.n4029 gnd.n4028 585
R7959 gnd.n1313 gnd.n1312 585
R7960 gnd.n1312 gnd.n1310 585
R7961 gnd.n4022 gnd.n4021 585
R7962 gnd.n4021 gnd.n4020 585
R7963 gnd.n1317 gnd.n1316 585
R7964 gnd.n3992 gnd.n1317 585
R7965 gnd.n1332 gnd.n1327 585
R7966 gnd.n4010 gnd.n1327 585
R7967 gnd.n3898 gnd.n3897 585
R7968 gnd.n3899 gnd.n3898 585
R7969 gnd.n1331 gnd.n1226 585
R7970 gnd.n4124 gnd.n1226 585
R7971 gnd.n3892 gnd.n3891 585
R7972 gnd.n3891 gnd.n3890 585
R7973 gnd.n1334 gnd.n1214 585
R7974 gnd.n4130 gnd.n1214 585
R7975 gnd.n5877 gnd.n5876 585
R7976 gnd.n5876 gnd.n5875 585
R7977 gnd.n5878 gnd.n793 585
R7978 gnd.n5785 gnd.n793 585
R7979 gnd.n5880 gnd.n5879 585
R7980 gnd.n5881 gnd.n5880 585
R7981 gnd.n794 gnd.n792 585
R7982 gnd.n792 gnd.n788 585
R7983 gnd.n775 gnd.n774 585
R7984 gnd.n779 gnd.n775 585
R7985 gnd.n5891 gnd.n5890 585
R7986 gnd.n5890 gnd.n5889 585
R7987 gnd.n5892 gnd.n769 585
R7988 gnd.n5774 gnd.n769 585
R7989 gnd.n5894 gnd.n5893 585
R7990 gnd.n5895 gnd.n5894 585
R7991 gnd.n770 gnd.n768 585
R7992 gnd.n5768 gnd.n768 585
R7993 gnd.n5749 gnd.n4586 585
R7994 gnd.n4586 gnd.n4585 585
R7995 gnd.n5751 gnd.n5750 585
R7996 gnd.n5752 gnd.n5751 585
R7997 gnd.n4587 gnd.n4584 585
R7998 gnd.n4584 gnd.n4580 585
R7999 gnd.n5456 gnd.n5455 585
R8000 gnd.n5455 gnd.n5454 585
R8001 gnd.n4594 gnd.n4593 585
R8002 gnd.n4603 gnd.n4594 585
R8003 gnd.n5445 gnd.n5444 585
R8004 gnd.n5444 gnd.n5443 585
R8005 gnd.n4601 gnd.n4600 585
R8006 gnd.n5431 gnd.n4601 585
R8007 gnd.n5406 gnd.n4618 585
R8008 gnd.n5399 gnd.n4618 585
R8009 gnd.n5408 gnd.n5407 585
R8010 gnd.n5409 gnd.n5408 585
R8011 gnd.n4619 gnd.n4617 585
R8012 gnd.n4627 gnd.n4617 585
R8013 gnd.n5382 gnd.n4639 585
R8014 gnd.n4639 gnd.n4626 585
R8015 gnd.n5384 gnd.n5383 585
R8016 gnd.n5385 gnd.n5384 585
R8017 gnd.n4640 gnd.n4638 585
R8018 gnd.n4638 gnd.n4634 585
R8019 gnd.n5370 gnd.n5369 585
R8020 gnd.n5369 gnd.n5368 585
R8021 gnd.n4645 gnd.n4644 585
R8022 gnd.n4649 gnd.n4645 585
R8023 gnd.n5354 gnd.n5353 585
R8024 gnd.n5355 gnd.n5354 585
R8025 gnd.n4659 gnd.n4658 585
R8026 gnd.n5345 gnd.n4658 585
R8027 gnd.n5319 gnd.n4674 585
R8028 gnd.n4674 gnd.n4666 585
R8029 gnd.n5321 gnd.n5320 585
R8030 gnd.n5322 gnd.n5321 585
R8031 gnd.n4675 gnd.n4673 585
R8032 gnd.n4679 gnd.n4673 585
R8033 gnd.n5300 gnd.n5299 585
R8034 gnd.n5301 gnd.n5300 585
R8035 gnd.n4691 gnd.n4690 585
R8036 gnd.n4690 gnd.n4686 585
R8037 gnd.n5290 gnd.n5289 585
R8038 gnd.n5291 gnd.n5290 585
R8039 gnd.n4699 gnd.n4698 585
R8040 gnd.n4703 gnd.n4698 585
R8041 gnd.n5268 gnd.n4715 585
R8042 gnd.n5059 gnd.n4715 585
R8043 gnd.n5270 gnd.n5269 585
R8044 gnd.n5271 gnd.n5270 585
R8045 gnd.n4716 gnd.n4714 585
R8046 gnd.n4714 gnd.n4710 585
R8047 gnd.n5259 gnd.n5258 585
R8048 gnd.n5260 gnd.n5259 585
R8049 gnd.n4724 gnd.n4723 585
R8050 gnd.n4729 gnd.n4723 585
R8051 gnd.n5237 gnd.n4741 585
R8052 gnd.n4741 gnd.n4728 585
R8053 gnd.n5239 gnd.n5238 585
R8054 gnd.n5240 gnd.n5239 585
R8055 gnd.n4742 gnd.n4740 585
R8056 gnd.n4740 gnd.n4736 585
R8057 gnd.n5228 gnd.n5227 585
R8058 gnd.n5229 gnd.n5228 585
R8059 gnd.n4750 gnd.n4749 585
R8060 gnd.n5112 gnd.n4749 585
R8061 gnd.n5206 gnd.n4766 585
R8062 gnd.n4766 gnd.n4754 585
R8063 gnd.n5208 gnd.n5207 585
R8064 gnd.n5209 gnd.n5208 585
R8065 gnd.n4767 gnd.n4765 585
R8066 gnd.n4765 gnd.n4761 585
R8067 gnd.n5197 gnd.n5196 585
R8068 gnd.n5198 gnd.n5197 585
R8069 gnd.n4774 gnd.n4773 585
R8070 gnd.n4779 gnd.n4773 585
R8071 gnd.n5175 gnd.n4792 585
R8072 gnd.n4792 gnd.n4778 585
R8073 gnd.n5177 gnd.n5176 585
R8074 gnd.n5178 gnd.n5177 585
R8075 gnd.n4793 gnd.n4791 585
R8076 gnd.n4791 gnd.n4787 585
R8077 gnd.n5166 gnd.n5165 585
R8078 gnd.n5167 gnd.n5166 585
R8079 gnd.n4800 gnd.n4799 585
R8080 gnd.n4804 gnd.n4799 585
R8081 gnd.n5143 gnd.n4821 585
R8082 gnd.n4821 gnd.n4803 585
R8083 gnd.n5145 gnd.n5144 585
R8084 gnd.n5146 gnd.n5145 585
R8085 gnd.n4822 gnd.n4820 585
R8086 gnd.n4820 gnd.n4811 585
R8087 gnd.n5138 gnd.n5137 585
R8088 gnd.n5137 gnd.n5136 585
R8089 gnd.n4869 gnd.n4868 585
R8090 gnd.n4870 gnd.n4869 585
R8091 gnd.n5023 gnd.n5022 585
R8092 gnd.n5024 gnd.n5023 585
R8093 gnd.n4879 gnd.n4878 585
R8094 gnd.n4878 gnd.n4877 585
R8095 gnd.n5018 gnd.n5017 585
R8096 gnd.n5017 gnd.n5016 585
R8097 gnd.n4882 gnd.n4881 585
R8098 gnd.n4883 gnd.n4882 585
R8099 gnd.n5007 gnd.n5006 585
R8100 gnd.n5008 gnd.n5007 585
R8101 gnd.n4890 gnd.n4889 585
R8102 gnd.n4999 gnd.n4889 585
R8103 gnd.n5002 gnd.n5001 585
R8104 gnd.n5001 gnd.n5000 585
R8105 gnd.n4893 gnd.n4892 585
R8106 gnd.n4894 gnd.n4893 585
R8107 gnd.n4988 gnd.n4987 585
R8108 gnd.n4986 gnd.n4912 585
R8109 gnd.n4985 gnd.n4911 585
R8110 gnd.n4990 gnd.n4911 585
R8111 gnd.n4984 gnd.n4983 585
R8112 gnd.n4982 gnd.n4981 585
R8113 gnd.n4980 gnd.n4979 585
R8114 gnd.n4978 gnd.n4977 585
R8115 gnd.n4976 gnd.n4975 585
R8116 gnd.n4974 gnd.n4973 585
R8117 gnd.n4972 gnd.n4971 585
R8118 gnd.n4970 gnd.n4969 585
R8119 gnd.n4968 gnd.n4967 585
R8120 gnd.n4966 gnd.n4965 585
R8121 gnd.n4964 gnd.n4963 585
R8122 gnd.n4962 gnd.n4961 585
R8123 gnd.n4960 gnd.n4959 585
R8124 gnd.n4958 gnd.n4957 585
R8125 gnd.n4956 gnd.n4955 585
R8126 gnd.n4954 gnd.n4953 585
R8127 gnd.n4952 gnd.n4951 585
R8128 gnd.n4950 gnd.n4949 585
R8129 gnd.n4948 gnd.n4947 585
R8130 gnd.n4946 gnd.n4945 585
R8131 gnd.n4944 gnd.n4943 585
R8132 gnd.n4942 gnd.n4941 585
R8133 gnd.n4899 gnd.n4898 585
R8134 gnd.n4993 gnd.n4992 585
R8135 gnd.n5793 gnd.n5792 585
R8136 gnd.n5794 gnd.n4562 585
R8137 gnd.n5796 gnd.n5795 585
R8138 gnd.n5798 gnd.n4561 585
R8139 gnd.n5800 gnd.n5799 585
R8140 gnd.n5801 gnd.n4552 585
R8141 gnd.n5803 gnd.n5802 585
R8142 gnd.n5805 gnd.n4550 585
R8143 gnd.n5807 gnd.n5806 585
R8144 gnd.n5808 gnd.n4545 585
R8145 gnd.n5810 gnd.n5809 585
R8146 gnd.n5812 gnd.n4543 585
R8147 gnd.n5814 gnd.n5813 585
R8148 gnd.n5815 gnd.n4538 585
R8149 gnd.n5817 gnd.n5816 585
R8150 gnd.n5819 gnd.n4536 585
R8151 gnd.n5821 gnd.n5820 585
R8152 gnd.n5822 gnd.n4531 585
R8153 gnd.n5824 gnd.n5823 585
R8154 gnd.n5826 gnd.n4529 585
R8155 gnd.n5828 gnd.n5827 585
R8156 gnd.n5829 gnd.n4524 585
R8157 gnd.n5831 gnd.n5830 585
R8158 gnd.n5833 gnd.n4522 585
R8159 gnd.n5835 gnd.n5834 585
R8160 gnd.n5836 gnd.n4520 585
R8161 gnd.n5837 gnd.n798 585
R8162 gnd.n4483 gnd.n798 585
R8163 gnd.n5788 gnd.n800 585
R8164 gnd.n5875 gnd.n800 585
R8165 gnd.n5787 gnd.n5786 585
R8166 gnd.n5786 gnd.n5785 585
R8167 gnd.n5784 gnd.n790 585
R8168 gnd.n5881 gnd.n790 585
R8169 gnd.n5778 gnd.n4567 585
R8170 gnd.n5778 gnd.n788 585
R8171 gnd.n5780 gnd.n5779 585
R8172 gnd.n5779 gnd.n779 585
R8173 gnd.n5777 gnd.n777 585
R8174 gnd.n5889 gnd.n777 585
R8175 gnd.n5776 gnd.n5775 585
R8176 gnd.n5775 gnd.n5774 585
R8177 gnd.n4569 gnd.n766 585
R8178 gnd.n5895 gnd.n766 585
R8179 gnd.n5770 gnd.n5769 585
R8180 gnd.n5769 gnd.n5768 585
R8181 gnd.n4572 gnd.n4571 585
R8182 gnd.n4585 gnd.n4572 585
R8183 gnd.n5420 gnd.n4582 585
R8184 gnd.n5752 gnd.n4582 585
R8185 gnd.n5422 gnd.n5421 585
R8186 gnd.n5421 gnd.n4580 585
R8187 gnd.n5423 gnd.n4596 585
R8188 gnd.n5454 gnd.n4596 585
R8189 gnd.n5425 gnd.n5424 585
R8190 gnd.n5424 gnd.n4603 585
R8191 gnd.n5426 gnd.n4602 585
R8192 gnd.n5443 gnd.n4602 585
R8193 gnd.n5428 gnd.n5427 585
R8194 gnd.n5431 gnd.n5428 585
R8195 gnd.n4612 gnd.n4611 585
R8196 gnd.n5399 gnd.n4611 585
R8197 gnd.n5411 gnd.n5410 585
R8198 gnd.n5410 gnd.n5409 585
R8199 gnd.n4615 gnd.n4614 585
R8200 gnd.n4627 gnd.n4615 585
R8201 gnd.n5335 gnd.n5334 585
R8202 gnd.n5334 gnd.n4626 585
R8203 gnd.n5336 gnd.n4636 585
R8204 gnd.n5385 gnd.n4636 585
R8205 gnd.n5338 gnd.n5337 585
R8206 gnd.n5337 gnd.n4634 585
R8207 gnd.n5339 gnd.n4646 585
R8208 gnd.n5368 gnd.n4646 585
R8209 gnd.n5341 gnd.n5340 585
R8210 gnd.n5340 gnd.n4649 585
R8211 gnd.n5342 gnd.n4656 585
R8212 gnd.n5355 gnd.n4656 585
R8213 gnd.n5344 gnd.n5343 585
R8214 gnd.n5345 gnd.n5344 585
R8215 gnd.n4668 gnd.n4667 585
R8216 gnd.n4667 gnd.n4666 585
R8217 gnd.n5324 gnd.n5323 585
R8218 gnd.n5323 gnd.n5322 585
R8219 gnd.n4671 gnd.n4670 585
R8220 gnd.n4679 gnd.n4671 585
R8221 gnd.n5051 gnd.n4688 585
R8222 gnd.n5301 gnd.n4688 585
R8223 gnd.n5054 gnd.n5053 585
R8224 gnd.n5053 gnd.n4686 585
R8225 gnd.n5055 gnd.n4697 585
R8226 gnd.n5291 gnd.n4697 585
R8227 gnd.n5058 gnd.n5057 585
R8228 gnd.n5058 gnd.n4703 585
R8229 gnd.n5061 gnd.n5060 585
R8230 gnd.n5060 gnd.n5059 585
R8231 gnd.n5062 gnd.n4712 585
R8232 gnd.n5271 gnd.n4712 585
R8233 gnd.n5050 gnd.n5049 585
R8234 gnd.n5049 gnd.n4710 585
R8235 gnd.n5102 gnd.n4722 585
R8236 gnd.n5260 gnd.n4722 585
R8237 gnd.n5104 gnd.n5103 585
R8238 gnd.n5104 gnd.n4729 585
R8239 gnd.n5106 gnd.n5105 585
R8240 gnd.n5105 gnd.n4728 585
R8241 gnd.n5107 gnd.n4738 585
R8242 gnd.n5240 gnd.n4738 585
R8243 gnd.n5109 gnd.n5108 585
R8244 gnd.n5108 gnd.n4736 585
R8245 gnd.n5110 gnd.n4748 585
R8246 gnd.n5229 gnd.n4748 585
R8247 gnd.n5113 gnd.n5111 585
R8248 gnd.n5113 gnd.n5112 585
R8249 gnd.n5115 gnd.n5114 585
R8250 gnd.n5114 gnd.n4754 585
R8251 gnd.n5116 gnd.n4763 585
R8252 gnd.n5209 gnd.n4763 585
R8253 gnd.n5118 gnd.n5117 585
R8254 gnd.n5117 gnd.n4761 585
R8255 gnd.n5119 gnd.n4772 585
R8256 gnd.n5198 gnd.n4772 585
R8257 gnd.n5121 gnd.n5120 585
R8258 gnd.n5121 gnd.n4779 585
R8259 gnd.n5123 gnd.n5122 585
R8260 gnd.n5122 gnd.n4778 585
R8261 gnd.n5124 gnd.n4789 585
R8262 gnd.n5178 gnd.n4789 585
R8263 gnd.n5126 gnd.n5125 585
R8264 gnd.n5125 gnd.n4787 585
R8265 gnd.n5127 gnd.n4798 585
R8266 gnd.n5167 gnd.n4798 585
R8267 gnd.n5129 gnd.n5128 585
R8268 gnd.n5129 gnd.n4804 585
R8269 gnd.n5131 gnd.n5130 585
R8270 gnd.n5130 gnd.n4803 585
R8271 gnd.n5132 gnd.n4819 585
R8272 gnd.n5146 gnd.n4819 585
R8273 gnd.n5133 gnd.n4872 585
R8274 gnd.n4872 gnd.n4811 585
R8275 gnd.n5135 gnd.n5134 585
R8276 gnd.n5136 gnd.n5135 585
R8277 gnd.n4873 gnd.n4871 585
R8278 gnd.n4871 gnd.n4870 585
R8279 gnd.n5026 gnd.n5025 585
R8280 gnd.n5025 gnd.n5024 585
R8281 gnd.n4876 gnd.n4875 585
R8282 gnd.n4877 gnd.n4876 585
R8283 gnd.n5015 gnd.n5014 585
R8284 gnd.n5016 gnd.n5015 585
R8285 gnd.n4885 gnd.n4884 585
R8286 gnd.n4884 gnd.n4883 585
R8287 gnd.n5010 gnd.n5009 585
R8288 gnd.n5009 gnd.n5008 585
R8289 gnd.n4888 gnd.n4887 585
R8290 gnd.n4999 gnd.n4888 585
R8291 gnd.n4998 gnd.n4997 585
R8292 gnd.n5000 gnd.n4998 585
R8293 gnd.n4896 gnd.n4895 585
R8294 gnd.n4895 gnd.n4894 585
R8295 gnd.n5873 gnd.n5872 585
R8296 gnd.n5874 gnd.n5873 585
R8297 gnd.n4486 gnd.n4484 585
R8298 gnd.n4484 gnd.n799 585
R8299 gnd.n787 gnd.n786 585
R8300 gnd.n791 gnd.n787 585
R8301 gnd.n5884 gnd.n5883 585
R8302 gnd.n5883 gnd.n5882 585
R8303 gnd.n5885 gnd.n781 585
R8304 gnd.n5737 gnd.n781 585
R8305 gnd.n5887 gnd.n5886 585
R8306 gnd.n5888 gnd.n5887 585
R8307 gnd.n782 gnd.n780 585
R8308 gnd.n780 gnd.n776 585
R8309 gnd.n5763 gnd.n5762 585
R8310 gnd.n5762 gnd.n767 585
R8311 gnd.n5764 gnd.n4575 585
R8312 gnd.n4575 gnd.n765 585
R8313 gnd.n5766 gnd.n5765 585
R8314 gnd.n5767 gnd.n5766 585
R8315 gnd.n4576 gnd.n4574 585
R8316 gnd.n4583 gnd.n4574 585
R8317 gnd.n5755 gnd.n5754 585
R8318 gnd.n5754 gnd.n5753 585
R8319 gnd.n4579 gnd.n4578 585
R8320 gnd.n5453 gnd.n4579 585
R8321 gnd.n5439 gnd.n4605 585
R8322 gnd.n4605 gnd.n4595 585
R8323 gnd.n5441 gnd.n5440 585
R8324 gnd.n5442 gnd.n5441 585
R8325 gnd.n4606 gnd.n4604 585
R8326 gnd.n5430 gnd.n4604 585
R8327 gnd.n5434 gnd.n5433 585
R8328 gnd.n5433 gnd.n5432 585
R8329 gnd.n4609 gnd.n4608 585
R8330 gnd.n5400 gnd.n4609 585
R8331 gnd.n5393 gnd.n4629 585
R8332 gnd.n4629 gnd.n4616 585
R8333 gnd.n5395 gnd.n5394 585
R8334 gnd.n5396 gnd.n5395 585
R8335 gnd.n4630 gnd.n4628 585
R8336 gnd.n4637 gnd.n4628 585
R8337 gnd.n5388 gnd.n5387 585
R8338 gnd.n5387 gnd.n5386 585
R8339 gnd.n4633 gnd.n4632 585
R8340 gnd.n5367 gnd.n4633 585
R8341 gnd.n5363 gnd.n5362 585
R8342 gnd.n5364 gnd.n5363 585
R8343 gnd.n4651 gnd.n4650 585
R8344 gnd.n4657 gnd.n4650 585
R8345 gnd.n5358 gnd.n5357 585
R8346 gnd.n5357 gnd.n5356 585
R8347 gnd.n4654 gnd.n4653 585
R8348 gnd.n5346 gnd.n4654 585
R8349 gnd.n5309 gnd.n4681 585
R8350 gnd.n4681 gnd.n4672 585
R8351 gnd.n5311 gnd.n5310 585
R8352 gnd.n5312 gnd.n5311 585
R8353 gnd.n4682 gnd.n4680 585
R8354 gnd.n4689 gnd.n4680 585
R8355 gnd.n5304 gnd.n5303 585
R8356 gnd.n5303 gnd.n5302 585
R8357 gnd.n4685 gnd.n4684 585
R8358 gnd.n5292 gnd.n4685 585
R8359 gnd.n5279 gnd.n4705 585
R8360 gnd.n4705 gnd.n4696 585
R8361 gnd.n5281 gnd.n5280 585
R8362 gnd.n5282 gnd.n5281 585
R8363 gnd.n4706 gnd.n4704 585
R8364 gnd.n4713 gnd.n4704 585
R8365 gnd.n5274 gnd.n5273 585
R8366 gnd.n5273 gnd.n5272 585
R8367 gnd.n4709 gnd.n4708 585
R8368 gnd.n5261 gnd.n4709 585
R8369 gnd.n5248 gnd.n4731 585
R8370 gnd.n4731 gnd.n4721 585
R8371 gnd.n5250 gnd.n5249 585
R8372 gnd.n5251 gnd.n5250 585
R8373 gnd.n4732 gnd.n4730 585
R8374 gnd.n4739 gnd.n4730 585
R8375 gnd.n5243 gnd.n5242 585
R8376 gnd.n5242 gnd.n5241 585
R8377 gnd.n4735 gnd.n4734 585
R8378 gnd.n5230 gnd.n4735 585
R8379 gnd.n5217 gnd.n4756 585
R8380 gnd.n4756 gnd.n4747 585
R8381 gnd.n5219 gnd.n5218 585
R8382 gnd.n5220 gnd.n5219 585
R8383 gnd.n4757 gnd.n4755 585
R8384 gnd.n4764 gnd.n4755 585
R8385 gnd.n5212 gnd.n5211 585
R8386 gnd.n5211 gnd.n5210 585
R8387 gnd.n4760 gnd.n4759 585
R8388 gnd.n5199 gnd.n4760 585
R8389 gnd.n5186 gnd.n4782 585
R8390 gnd.n4782 gnd.n4781 585
R8391 gnd.n5188 gnd.n5187 585
R8392 gnd.n5189 gnd.n5188 585
R8393 gnd.n4783 gnd.n4780 585
R8394 gnd.n4790 gnd.n4780 585
R8395 gnd.n5181 gnd.n5180 585
R8396 gnd.n5180 gnd.n5179 585
R8397 gnd.n4786 gnd.n4785 585
R8398 gnd.n5168 gnd.n4786 585
R8399 gnd.n5155 gnd.n4807 585
R8400 gnd.n4807 gnd.n4806 585
R8401 gnd.n5157 gnd.n5156 585
R8402 gnd.n5158 gnd.n5157 585
R8403 gnd.n5151 gnd.n4805 585
R8404 gnd.n5150 gnd.n5149 585
R8405 gnd.n4810 gnd.n4809 585
R8406 gnd.n5147 gnd.n4810 585
R8407 gnd.n4832 gnd.n4831 585
R8408 gnd.n4835 gnd.n4834 585
R8409 gnd.n4833 gnd.n4828 585
R8410 gnd.n4840 gnd.n4839 585
R8411 gnd.n4842 gnd.n4841 585
R8412 gnd.n4845 gnd.n4844 585
R8413 gnd.n4843 gnd.n4826 585
R8414 gnd.n4850 gnd.n4849 585
R8415 gnd.n4852 gnd.n4851 585
R8416 gnd.n4855 gnd.n4854 585
R8417 gnd.n4853 gnd.n4824 585
R8418 gnd.n4860 gnd.n4859 585
R8419 gnd.n4864 gnd.n4861 585
R8420 gnd.n4865 gnd.n4802 585
R8421 gnd.n5842 gnd.n5841 585
R8422 gnd.n5844 gnd.n4515 585
R8423 gnd.n5846 gnd.n5845 585
R8424 gnd.n5847 gnd.n4508 585
R8425 gnd.n5849 gnd.n5848 585
R8426 gnd.n5851 gnd.n4506 585
R8427 gnd.n5853 gnd.n5852 585
R8428 gnd.n5854 gnd.n4501 585
R8429 gnd.n5856 gnd.n5855 585
R8430 gnd.n5858 gnd.n4499 585
R8431 gnd.n5860 gnd.n5859 585
R8432 gnd.n5861 gnd.n4494 585
R8433 gnd.n5863 gnd.n5862 585
R8434 gnd.n5865 gnd.n4492 585
R8435 gnd.n5867 gnd.n5866 585
R8436 gnd.n5868 gnd.n4490 585
R8437 gnd.n5869 gnd.n4485 585
R8438 gnd.n4485 gnd.n4483 585
R8439 gnd.n5731 gnd.n801 585
R8440 gnd.n5874 gnd.n801 585
R8441 gnd.n5733 gnd.n5732 585
R8442 gnd.n5733 gnd.n799 585
R8443 gnd.n5735 gnd.n5734 585
R8444 gnd.n5734 gnd.n791 585
R8445 gnd.n5736 gnd.n789 585
R8446 gnd.n5882 gnd.n789 585
R8447 gnd.n5739 gnd.n5738 585
R8448 gnd.n5738 gnd.n5737 585
R8449 gnd.n5740 gnd.n778 585
R8450 gnd.n5888 gnd.n778 585
R8451 gnd.n5742 gnd.n5741 585
R8452 gnd.n5742 gnd.n776 585
R8453 gnd.n5743 gnd.n5466 585
R8454 gnd.n5743 gnd.n767 585
R8455 gnd.n5745 gnd.n5744 585
R8456 gnd.n5744 gnd.n765 585
R8457 gnd.n5746 gnd.n4573 585
R8458 gnd.n5767 gnd.n4573 585
R8459 gnd.n5463 gnd.n5462 585
R8460 gnd.n5462 gnd.n4583 585
R8461 gnd.n5461 gnd.n4581 585
R8462 gnd.n5753 gnd.n4581 585
R8463 gnd.n5452 gnd.n4591 585
R8464 gnd.n5453 gnd.n5452 585
R8465 gnd.n5451 gnd.n5450 585
R8466 gnd.n5451 gnd.n4595 585
R8467 gnd.n5449 gnd.n4597 585
R8468 gnd.n5442 gnd.n4597 585
R8469 gnd.n5429 gnd.n4598 585
R8470 gnd.n5430 gnd.n5429 585
R8471 gnd.n5403 gnd.n4610 585
R8472 gnd.n5432 gnd.n4610 585
R8473 gnd.n5402 gnd.n5401 585
R8474 gnd.n5401 gnd.n5400 585
R8475 gnd.n5398 gnd.n4623 585
R8476 gnd.n5398 gnd.n4616 585
R8477 gnd.n5397 gnd.n4625 585
R8478 gnd.n5397 gnd.n5396 585
R8479 gnd.n5376 gnd.n4624 585
R8480 gnd.n4637 gnd.n4624 585
R8481 gnd.n5375 gnd.n4635 585
R8482 gnd.n5386 gnd.n4635 585
R8483 gnd.n5366 gnd.n4642 585
R8484 gnd.n5367 gnd.n5366 585
R8485 gnd.n5365 gnd.n4648 585
R8486 gnd.n5365 gnd.n5364 585
R8487 gnd.n5350 gnd.n4647 585
R8488 gnd.n4657 gnd.n4647 585
R8489 gnd.n5349 gnd.n4655 585
R8490 gnd.n5356 gnd.n4655 585
R8491 gnd.n5348 gnd.n5347 585
R8492 gnd.n5347 gnd.n5346 585
R8493 gnd.n4665 gnd.n4662 585
R8494 gnd.n4672 gnd.n4665 585
R8495 gnd.n5314 gnd.n5313 585
R8496 gnd.n5313 gnd.n5312 585
R8497 gnd.n4678 gnd.n4677 585
R8498 gnd.n4689 gnd.n4678 585
R8499 gnd.n5295 gnd.n4687 585
R8500 gnd.n5302 gnd.n4687 585
R8501 gnd.n5294 gnd.n5293 585
R8502 gnd.n5293 gnd.n5292 585
R8503 gnd.n4695 gnd.n4693 585
R8504 gnd.n4696 gnd.n4695 585
R8505 gnd.n5284 gnd.n5283 585
R8506 gnd.n5283 gnd.n5282 585
R8507 gnd.n4702 gnd.n4701 585
R8508 gnd.n4713 gnd.n4702 585
R8509 gnd.n5264 gnd.n4711 585
R8510 gnd.n5272 gnd.n4711 585
R8511 gnd.n5263 gnd.n5262 585
R8512 gnd.n5262 gnd.n5261 585
R8513 gnd.n4720 gnd.n4718 585
R8514 gnd.n4721 gnd.n4720 585
R8515 gnd.n5253 gnd.n5252 585
R8516 gnd.n5252 gnd.n5251 585
R8517 gnd.n4727 gnd.n4726 585
R8518 gnd.n4739 gnd.n4727 585
R8519 gnd.n5233 gnd.n4737 585
R8520 gnd.n5241 gnd.n4737 585
R8521 gnd.n5232 gnd.n5231 585
R8522 gnd.n5231 gnd.n5230 585
R8523 gnd.n4746 gnd.n4744 585
R8524 gnd.n4747 gnd.n4746 585
R8525 gnd.n5222 gnd.n5221 585
R8526 gnd.n5221 gnd.n5220 585
R8527 gnd.n4753 gnd.n4752 585
R8528 gnd.n4764 gnd.n4753 585
R8529 gnd.n5202 gnd.n4762 585
R8530 gnd.n5210 gnd.n4762 585
R8531 gnd.n5201 gnd.n5200 585
R8532 gnd.n5200 gnd.n5199 585
R8533 gnd.n4771 gnd.n4769 585
R8534 gnd.n4781 gnd.n4771 585
R8535 gnd.n5191 gnd.n5190 585
R8536 gnd.n5190 gnd.n5189 585
R8537 gnd.n4777 gnd.n4776 585
R8538 gnd.n4790 gnd.n4777 585
R8539 gnd.n5171 gnd.n4788 585
R8540 gnd.n5179 gnd.n4788 585
R8541 gnd.n5170 gnd.n5169 585
R8542 gnd.n5169 gnd.n5168 585
R8543 gnd.n4797 gnd.n4795 585
R8544 gnd.n4806 gnd.n4797 585
R8545 gnd.n5160 gnd.n5159 585
R8546 gnd.n5159 gnd.n5158 585
R8547 gnd.n4279 gnd.n4278 585
R8548 gnd.n4278 gnd.n4277 585
R8549 gnd.n4280 gnd.n1073 585
R8550 gnd.n2662 gnd.n1073 585
R8551 gnd.n4282 gnd.n4281 585
R8552 gnd.n4283 gnd.n4282 585
R8553 gnd.n1057 gnd.n1056 585
R8554 gnd.n2543 gnd.n1057 585
R8555 gnd.n4291 gnd.n4290 585
R8556 gnd.n4290 gnd.n4289 585
R8557 gnd.n4292 gnd.n1051 585
R8558 gnd.n2534 gnd.n1051 585
R8559 gnd.n4294 gnd.n4293 585
R8560 gnd.n4295 gnd.n4294 585
R8561 gnd.n1036 gnd.n1035 585
R8562 gnd.n2554 gnd.n1036 585
R8563 gnd.n4303 gnd.n4302 585
R8564 gnd.n4302 gnd.n4301 585
R8565 gnd.n4304 gnd.n1030 585
R8566 gnd.n2526 gnd.n1030 585
R8567 gnd.n4306 gnd.n4305 585
R8568 gnd.n4307 gnd.n4306 585
R8569 gnd.n1015 gnd.n1014 585
R8570 gnd.n2518 gnd.n1015 585
R8571 gnd.n4315 gnd.n4314 585
R8572 gnd.n4314 gnd.n4313 585
R8573 gnd.n4316 gnd.n1009 585
R8574 gnd.n2510 gnd.n1009 585
R8575 gnd.n4318 gnd.n4317 585
R8576 gnd.n4319 gnd.n4318 585
R8577 gnd.n994 gnd.n993 585
R8578 gnd.n2502 gnd.n994 585
R8579 gnd.n4327 gnd.n4326 585
R8580 gnd.n4326 gnd.n4325 585
R8581 gnd.n4328 gnd.n991 585
R8582 gnd.n2445 gnd.n991 585
R8583 gnd.n4331 gnd.n4330 585
R8584 gnd.n4332 gnd.n4331 585
R8585 gnd.n992 gnd.n977 585
R8586 gnd.n2453 gnd.n977 585
R8587 gnd.n4340 gnd.n4339 585
R8588 gnd.n4339 gnd.n4338 585
R8589 gnd.n4341 gnd.n974 585
R8590 gnd.n2431 gnd.n974 585
R8591 gnd.n4344 gnd.n4343 585
R8592 gnd.n4345 gnd.n4344 585
R8593 gnd.n975 gnd.n956 585
R8594 gnd.n960 gnd.n956 585
R8595 gnd.n4353 gnd.n4352 585
R8596 gnd.n4352 gnd.n4351 585
R8597 gnd.n4354 gnd.n954 585
R8598 gnd.n2420 gnd.n954 585
R8599 gnd.n4356 gnd.n950 585
R8600 gnd.n950 gnd.n949 585
R8601 gnd.n4358 gnd.n4357 585
R8602 gnd.n4359 gnd.n4358 585
R8603 gnd.n935 gnd.n934 585
R8604 gnd.n939 gnd.n935 585
R8605 gnd.n4367 gnd.n4366 585
R8606 gnd.n4366 gnd.n4365 585
R8607 gnd.n4368 gnd.n929 585
R8608 gnd.n936 gnd.n929 585
R8609 gnd.n4370 gnd.n4369 585
R8610 gnd.n4371 gnd.n4370 585
R8611 gnd.n916 gnd.n915 585
R8612 gnd.n926 gnd.n916 585
R8613 gnd.n4379 gnd.n4378 585
R8614 gnd.n4378 gnd.n4377 585
R8615 gnd.n4380 gnd.n910 585
R8616 gnd.n910 gnd.n909 585
R8617 gnd.n4382 gnd.n4381 585
R8618 gnd.n4383 gnd.n4382 585
R8619 gnd.n895 gnd.n894 585
R8620 gnd.n898 gnd.n895 585
R8621 gnd.n4391 gnd.n4390 585
R8622 gnd.n4390 gnd.n4389 585
R8623 gnd.n4392 gnd.n889 585
R8624 gnd.n889 gnd.n886 585
R8625 gnd.n4394 gnd.n4393 585
R8626 gnd.n4395 gnd.n4394 585
R8627 gnd.n890 gnd.n888 585
R8628 gnd.n888 gnd.n884 585
R8629 gnd.n2350 gnd.n2349 585
R8630 gnd.n2351 gnd.n2350 585
R8631 gnd.n2345 gnd.n833 585
R8632 gnd.n833 gnd.n830 585
R8633 gnd.n4480 gnd.n4479 585
R8634 gnd.n4478 gnd.n832 585
R8635 gnd.n4477 gnd.n831 585
R8636 gnd.n4482 gnd.n831 585
R8637 gnd.n4476 gnd.n4475 585
R8638 gnd.n4474 gnd.n4473 585
R8639 gnd.n4472 gnd.n4471 585
R8640 gnd.n4470 gnd.n4469 585
R8641 gnd.n4468 gnd.n4467 585
R8642 gnd.n4466 gnd.n4465 585
R8643 gnd.n4464 gnd.n4463 585
R8644 gnd.n4462 gnd.n4461 585
R8645 gnd.n4460 gnd.n4459 585
R8646 gnd.n4458 gnd.n4457 585
R8647 gnd.n4456 gnd.n4455 585
R8648 gnd.n4454 gnd.n4453 585
R8649 gnd.n4452 gnd.n4451 585
R8650 gnd.n4450 gnd.n4449 585
R8651 gnd.n4448 gnd.n4447 585
R8652 gnd.n4445 gnd.n4444 585
R8653 gnd.n4443 gnd.n4442 585
R8654 gnd.n4441 gnd.n4440 585
R8655 gnd.n4439 gnd.n4438 585
R8656 gnd.n4437 gnd.n4436 585
R8657 gnd.n4435 gnd.n4434 585
R8658 gnd.n4433 gnd.n4432 585
R8659 gnd.n4431 gnd.n4430 585
R8660 gnd.n4429 gnd.n4428 585
R8661 gnd.n4427 gnd.n4426 585
R8662 gnd.n4425 gnd.n4424 585
R8663 gnd.n4423 gnd.n4422 585
R8664 gnd.n4421 gnd.n4420 585
R8665 gnd.n4419 gnd.n4418 585
R8666 gnd.n4417 gnd.n4416 585
R8667 gnd.n4415 gnd.n4414 585
R8668 gnd.n4413 gnd.n4412 585
R8669 gnd.n4411 gnd.n4410 585
R8670 gnd.n4409 gnd.n872 585
R8671 gnd.n876 gnd.n873 585
R8672 gnd.n4405 gnd.n4404 585
R8673 gnd.n2669 gnd.n2668 585
R8674 gnd.n2671 gnd.n2026 585
R8675 gnd.n2673 gnd.n2672 585
R8676 gnd.n2674 gnd.n2019 585
R8677 gnd.n2676 gnd.n2675 585
R8678 gnd.n2678 gnd.n2017 585
R8679 gnd.n2680 gnd.n2679 585
R8680 gnd.n2681 gnd.n2012 585
R8681 gnd.n2683 gnd.n2682 585
R8682 gnd.n2685 gnd.n2010 585
R8683 gnd.n2687 gnd.n2686 585
R8684 gnd.n2688 gnd.n2005 585
R8685 gnd.n2690 gnd.n2689 585
R8686 gnd.n2692 gnd.n2003 585
R8687 gnd.n2694 gnd.n2693 585
R8688 gnd.n2695 gnd.n1998 585
R8689 gnd.n2697 gnd.n2696 585
R8690 gnd.n2699 gnd.n1997 585
R8691 gnd.n2700 gnd.n1940 585
R8692 gnd.n2703 gnd.n2702 585
R8693 gnd.n1941 gnd.n1933 585
R8694 gnd.n1969 gnd.n1934 585
R8695 gnd.n1971 gnd.n1970 585
R8696 gnd.n1973 gnd.n1972 585
R8697 gnd.n1975 gnd.n1974 585
R8698 gnd.n1977 gnd.n1976 585
R8699 gnd.n1979 gnd.n1978 585
R8700 gnd.n1981 gnd.n1980 585
R8701 gnd.n1983 gnd.n1982 585
R8702 gnd.n1985 gnd.n1984 585
R8703 gnd.n1987 gnd.n1986 585
R8704 gnd.n1989 gnd.n1988 585
R8705 gnd.n1991 gnd.n1990 585
R8706 gnd.n1992 gnd.n1951 585
R8707 gnd.n1994 gnd.n1993 585
R8708 gnd.n1952 gnd.n1950 585
R8709 gnd.n1953 gnd.n1078 585
R8710 gnd.n1996 gnd.n1078 585
R8711 gnd.n2665 gnd.n1080 585
R8712 gnd.n4277 gnd.n1080 585
R8713 gnd.n2664 gnd.n2663 585
R8714 gnd.n2663 gnd.n2662 585
R8715 gnd.n2030 gnd.n1070 585
R8716 gnd.n4283 gnd.n1070 585
R8717 gnd.n2542 gnd.n2541 585
R8718 gnd.n2543 gnd.n2542 585
R8719 gnd.n2227 gnd.n1059 585
R8720 gnd.n4289 gnd.n1059 585
R8721 gnd.n2536 gnd.n2535 585
R8722 gnd.n2535 gnd.n2534 585
R8723 gnd.n2533 gnd.n1048 585
R8724 gnd.n4295 gnd.n1048 585
R8725 gnd.n2532 gnd.n2221 585
R8726 gnd.n2554 gnd.n2221 585
R8727 gnd.n2229 gnd.n1038 585
R8728 gnd.n4301 gnd.n1038 585
R8729 gnd.n2528 gnd.n2527 585
R8730 gnd.n2527 gnd.n2526 585
R8731 gnd.n2231 gnd.n1027 585
R8732 gnd.n4307 gnd.n1027 585
R8733 gnd.n2517 gnd.n2516 585
R8734 gnd.n2518 gnd.n2517 585
R8735 gnd.n2236 gnd.n1017 585
R8736 gnd.n4313 gnd.n1017 585
R8737 gnd.n2512 gnd.n2511 585
R8738 gnd.n2511 gnd.n2510 585
R8739 gnd.n2238 gnd.n1006 585
R8740 gnd.n4319 gnd.n1006 585
R8741 gnd.n2441 gnd.n2242 585
R8742 gnd.n2502 gnd.n2242 585
R8743 gnd.n2442 gnd.n996 585
R8744 gnd.n4325 gnd.n996 585
R8745 gnd.n2444 gnd.n2443 585
R8746 gnd.n2445 gnd.n2444 585
R8747 gnd.n2252 gnd.n988 585
R8748 gnd.n4332 gnd.n988 585
R8749 gnd.n2435 gnd.n2248 585
R8750 gnd.n2453 gnd.n2248 585
R8751 gnd.n2434 gnd.n979 585
R8752 gnd.n4338 gnd.n979 585
R8753 gnd.n2433 gnd.n2432 585
R8754 gnd.n2432 gnd.n2431 585
R8755 gnd.n2254 gnd.n971 585
R8756 gnd.n4345 gnd.n971 585
R8757 gnd.n2416 gnd.n2415 585
R8758 gnd.n2415 gnd.n960 585
R8759 gnd.n2417 gnd.n958 585
R8760 gnd.n4351 gnd.n958 585
R8761 gnd.n2419 gnd.n2418 585
R8762 gnd.n2420 gnd.n2419 585
R8763 gnd.n2382 gnd.n2381 585
R8764 gnd.n2381 gnd.n949 585
R8765 gnd.n2408 gnd.n947 585
R8766 gnd.n4359 gnd.n947 585
R8767 gnd.n2407 gnd.n2406 585
R8768 gnd.n2406 gnd.n939 585
R8769 gnd.n2405 gnd.n937 585
R8770 gnd.n4365 gnd.n937 585
R8771 gnd.n2385 gnd.n2384 585
R8772 gnd.n2384 gnd.n936 585
R8773 gnd.n2401 gnd.n927 585
R8774 gnd.n4371 gnd.n927 585
R8775 gnd.n2400 gnd.n2399 585
R8776 gnd.n2399 gnd.n926 585
R8777 gnd.n2398 gnd.n917 585
R8778 gnd.n4377 gnd.n917 585
R8779 gnd.n2388 gnd.n2387 585
R8780 gnd.n2387 gnd.n909 585
R8781 gnd.n2394 gnd.n907 585
R8782 gnd.n4383 gnd.n907 585
R8783 gnd.n2393 gnd.n2392 585
R8784 gnd.n2392 gnd.n898 585
R8785 gnd.n2391 gnd.n896 585
R8786 gnd.n4389 gnd.n896 585
R8787 gnd.n883 gnd.n881 585
R8788 gnd.n886 gnd.n883 585
R8789 gnd.n4397 gnd.n4396 585
R8790 gnd.n4396 gnd.n4395 585
R8791 gnd.n882 gnd.n879 585
R8792 gnd.n884 gnd.n882 585
R8793 gnd.n4401 gnd.n878 585
R8794 gnd.n2351 gnd.n878 585
R8795 gnd.n4403 gnd.n4402 585
R8796 gnd.n4403 gnd.n830 585
R8797 gnd.n6880 gnd.n6879 585
R8798 gnd.n6881 gnd.n6880 585
R8799 gnd.n87 gnd.n85 585
R8800 gnd.n85 gnd.n81 585
R8801 gnd.n6800 gnd.n6799 585
R8802 gnd.n6801 gnd.n6800 585
R8803 gnd.n165 gnd.n164 585
R8804 gnd.n164 gnd.n161 585
R8805 gnd.n6795 gnd.n6794 585
R8806 gnd.n6794 gnd.n6793 585
R8807 gnd.n168 gnd.n167 585
R8808 gnd.n170 gnd.n168 585
R8809 gnd.n6710 gnd.n6709 585
R8810 gnd.n6711 gnd.n6710 585
R8811 gnd.n181 gnd.n180 585
R8812 gnd.n188 gnd.n180 585
R8813 gnd.n6705 gnd.n6704 585
R8814 gnd.n6704 gnd.n6703 585
R8815 gnd.n184 gnd.n183 585
R8816 gnd.n186 gnd.n184 585
R8817 gnd.n6694 gnd.n6693 585
R8818 gnd.n6695 gnd.n6694 585
R8819 gnd.n197 gnd.n196 585
R8820 gnd.n196 gnd.n194 585
R8821 gnd.n6689 gnd.n6688 585
R8822 gnd.n6688 gnd.n6687 585
R8823 gnd.n200 gnd.n199 585
R8824 gnd.n202 gnd.n200 585
R8825 gnd.n6678 gnd.n6677 585
R8826 gnd.n6679 gnd.n6678 585
R8827 gnd.n211 gnd.n210 585
R8828 gnd.n224 gnd.n210 585
R8829 gnd.n6673 gnd.n6672 585
R8830 gnd.n6672 gnd.n6671 585
R8831 gnd.n220 gnd.n219 585
R8832 gnd.n222 gnd.n220 585
R8833 gnd.n6662 gnd.n6661 585
R8834 gnd.n6663 gnd.n6662 585
R8835 gnd.n6660 gnd.n6659 585
R8836 gnd.n6659 gnd.n230 585
R8837 gnd.n6658 gnd.n235 585
R8838 gnd.n6658 gnd.n6657 585
R8839 gnd.n234 gnd.n233 585
R8840 gnd.n3966 gnd.n233 585
R8841 gnd.n6648 gnd.n6647 585
R8842 gnd.n6649 gnd.n6648 585
R8843 gnd.n6646 gnd.n6645 585
R8844 gnd.n6645 gnd.n6644 585
R8845 gnd.n1264 gnd.n247 585
R8846 gnd.n4095 gnd.n247 585
R8847 gnd.n1266 gnd.n1265 585
R8848 gnd.n3972 gnd.n1266 585
R8849 gnd.n4085 gnd.n4084 585
R8850 gnd.n4086 gnd.n4085 585
R8851 gnd.n4083 gnd.n1263 585
R8852 gnd.n1274 gnd.n1263 585
R8853 gnd.n4082 gnd.n4081 585
R8854 gnd.n4081 gnd.n4080 585
R8855 gnd.n1269 gnd.n1267 585
R8856 gnd.n4061 gnd.n1269 585
R8857 gnd.n4049 gnd.n1294 585
R8858 gnd.n1294 gnd.n1281 585
R8859 gnd.n4051 gnd.n4050 585
R8860 gnd.n4052 gnd.n4051 585
R8861 gnd.n1295 gnd.n1293 585
R8862 gnd.n1302 gnd.n1293 585
R8863 gnd.n4043 gnd.n4042 585
R8864 gnd.n4042 gnd.n4041 585
R8865 gnd.n1298 gnd.n1297 585
R8866 gnd.n4029 gnd.n1298 585
R8867 gnd.n4017 gnd.n1322 585
R8868 gnd.n1322 gnd.n1310 585
R8869 gnd.n4019 gnd.n4018 585
R8870 gnd.n4020 gnd.n4019 585
R8871 gnd.n1323 gnd.n1321 585
R8872 gnd.n3992 gnd.n1321 585
R8873 gnd.n4012 gnd.n4011 585
R8874 gnd.n4011 gnd.n4010 585
R8875 gnd.n1223 gnd.n1222 585
R8876 gnd.n3899 gnd.n1223 585
R8877 gnd.n4126 gnd.n4125 585
R8878 gnd.n4125 gnd.n4124 585
R8879 gnd.n4127 gnd.n1218 585
R8880 gnd.n3890 gnd.n1218 585
R8881 gnd.n4129 gnd.n4128 585
R8882 gnd.n4130 gnd.n4129 585
R8883 gnd.n3789 gnd.n1217 585
R8884 gnd.n3794 gnd.n3792 585
R8885 gnd.n3795 gnd.n3788 585
R8886 gnd.n3795 gnd.n1204 585
R8887 gnd.n3798 gnd.n3797 585
R8888 gnd.n3786 gnd.n3785 585
R8889 gnd.n3803 gnd.n3802 585
R8890 gnd.n3805 gnd.n3784 585
R8891 gnd.n3808 gnd.n3807 585
R8892 gnd.n3782 gnd.n3781 585
R8893 gnd.n3813 gnd.n3812 585
R8894 gnd.n3815 gnd.n3780 585
R8895 gnd.n3818 gnd.n3817 585
R8896 gnd.n3778 gnd.n3777 585
R8897 gnd.n3824 gnd.n3823 585
R8898 gnd.n3826 gnd.n3776 585
R8899 gnd.n3827 gnd.n1360 585
R8900 gnd.n1358 gnd.n1357 585
R8901 gnd.n3837 gnd.n3836 585
R8902 gnd.n3839 gnd.n1356 585
R8903 gnd.n3842 gnd.n3841 585
R8904 gnd.n1354 gnd.n1353 585
R8905 gnd.n3847 gnd.n3846 585
R8906 gnd.n3849 gnd.n1352 585
R8907 gnd.n3852 gnd.n3851 585
R8908 gnd.n1350 gnd.n1349 585
R8909 gnd.n3857 gnd.n3856 585
R8910 gnd.n3859 gnd.n1348 585
R8911 gnd.n3862 gnd.n3861 585
R8912 gnd.n1346 gnd.n1345 585
R8913 gnd.n3867 gnd.n3866 585
R8914 gnd.n3869 gnd.n1344 585
R8915 gnd.n3872 gnd.n3871 585
R8916 gnd.n1342 gnd.n1341 585
R8917 gnd.n3878 gnd.n3877 585
R8918 gnd.n3880 gnd.n1340 585
R8919 gnd.n3881 gnd.n1339 585
R8920 gnd.n3884 gnd.n3883 585
R8921 gnd.n155 gnd.n154 585
R8922 gnd.n6809 gnd.n150 585
R8923 gnd.n6811 gnd.n6810 585
R8924 gnd.n6813 gnd.n148 585
R8925 gnd.n6815 gnd.n6814 585
R8926 gnd.n6816 gnd.n143 585
R8927 gnd.n6818 gnd.n6817 585
R8928 gnd.n6820 gnd.n141 585
R8929 gnd.n6822 gnd.n6821 585
R8930 gnd.n6823 gnd.n136 585
R8931 gnd.n6825 gnd.n6824 585
R8932 gnd.n6827 gnd.n134 585
R8933 gnd.n6829 gnd.n6828 585
R8934 gnd.n6830 gnd.n129 585
R8935 gnd.n6832 gnd.n6831 585
R8936 gnd.n6834 gnd.n127 585
R8937 gnd.n6836 gnd.n6835 585
R8938 gnd.n6837 gnd.n122 585
R8939 gnd.n6839 gnd.n6838 585
R8940 gnd.n6841 gnd.n120 585
R8941 gnd.n6843 gnd.n6842 585
R8942 gnd.n6847 gnd.n115 585
R8943 gnd.n6849 gnd.n6848 585
R8944 gnd.n6851 gnd.n113 585
R8945 gnd.n6853 gnd.n6852 585
R8946 gnd.n6854 gnd.n108 585
R8947 gnd.n6856 gnd.n6855 585
R8948 gnd.n6858 gnd.n106 585
R8949 gnd.n6860 gnd.n6859 585
R8950 gnd.n6861 gnd.n101 585
R8951 gnd.n6863 gnd.n6862 585
R8952 gnd.n6865 gnd.n99 585
R8953 gnd.n6867 gnd.n6866 585
R8954 gnd.n6868 gnd.n94 585
R8955 gnd.n6870 gnd.n6869 585
R8956 gnd.n6872 gnd.n92 585
R8957 gnd.n6874 gnd.n6873 585
R8958 gnd.n6875 gnd.n90 585
R8959 gnd.n6876 gnd.n86 585
R8960 gnd.n86 gnd.n83 585
R8961 gnd.n6805 gnd.n82 585
R8962 gnd.n6881 gnd.n82 585
R8963 gnd.n6804 gnd.n6803 585
R8964 gnd.n6803 gnd.n81 585
R8965 gnd.n6802 gnd.n159 585
R8966 gnd.n6802 gnd.n6801 585
R8967 gnd.n3939 gnd.n160 585
R8968 gnd.n161 gnd.n160 585
R8969 gnd.n3940 gnd.n171 585
R8970 gnd.n6793 gnd.n171 585
R8971 gnd.n3942 gnd.n3941 585
R8972 gnd.n3941 gnd.n170 585
R8973 gnd.n3943 gnd.n179 585
R8974 gnd.n6711 gnd.n179 585
R8975 gnd.n3945 gnd.n3944 585
R8976 gnd.n3944 gnd.n188 585
R8977 gnd.n3946 gnd.n187 585
R8978 gnd.n6703 gnd.n187 585
R8979 gnd.n3948 gnd.n3947 585
R8980 gnd.n3947 gnd.n186 585
R8981 gnd.n3949 gnd.n195 585
R8982 gnd.n6695 gnd.n195 585
R8983 gnd.n3951 gnd.n3950 585
R8984 gnd.n3950 gnd.n194 585
R8985 gnd.n3952 gnd.n203 585
R8986 gnd.n6687 gnd.n203 585
R8987 gnd.n3954 gnd.n3953 585
R8988 gnd.n3953 gnd.n202 585
R8989 gnd.n3955 gnd.n209 585
R8990 gnd.n6679 gnd.n209 585
R8991 gnd.n3957 gnd.n3956 585
R8992 gnd.n3956 gnd.n224 585
R8993 gnd.n3958 gnd.n223 585
R8994 gnd.n6671 gnd.n223 585
R8995 gnd.n3960 gnd.n3959 585
R8996 gnd.n3959 gnd.n222 585
R8997 gnd.n3961 gnd.n231 585
R8998 gnd.n6663 gnd.n231 585
R8999 gnd.n3963 gnd.n3962 585
R9000 gnd.n3962 gnd.n230 585
R9001 gnd.n3964 gnd.n237 585
R9002 gnd.n6657 gnd.n237 585
R9003 gnd.n3968 gnd.n3967 585
R9004 gnd.n3967 gnd.n3966 585
R9005 gnd.n3969 gnd.n244 585
R9006 gnd.n6649 gnd.n244 585
R9007 gnd.n3970 gnd.n249 585
R9008 gnd.n6644 gnd.n249 585
R9009 gnd.n3971 gnd.n1252 585
R9010 gnd.n4095 gnd.n1252 585
R9011 gnd.n3974 gnd.n3973 585
R9012 gnd.n3973 gnd.n3972 585
R9013 gnd.n3975 gnd.n1261 585
R9014 gnd.n4086 gnd.n1261 585
R9015 gnd.n3977 gnd.n3976 585
R9016 gnd.n3976 gnd.n1274 585
R9017 gnd.n3978 gnd.n1271 585
R9018 gnd.n4080 gnd.n1271 585
R9019 gnd.n3979 gnd.n1282 585
R9020 gnd.n4061 gnd.n1282 585
R9021 gnd.n3981 gnd.n3980 585
R9022 gnd.n3980 gnd.n1281 585
R9023 gnd.n3982 gnd.n1290 585
R9024 gnd.n4052 gnd.n1290 585
R9025 gnd.n3984 gnd.n3983 585
R9026 gnd.n3983 gnd.n1302 585
R9027 gnd.n3985 gnd.n1300 585
R9028 gnd.n4041 gnd.n1300 585
R9029 gnd.n3986 gnd.n1311 585
R9030 gnd.n4029 gnd.n1311 585
R9031 gnd.n3988 gnd.n3987 585
R9032 gnd.n3987 gnd.n1310 585
R9033 gnd.n3989 gnd.n1319 585
R9034 gnd.n4020 gnd.n1319 585
R9035 gnd.n3991 gnd.n3990 585
R9036 gnd.n3992 gnd.n3991 585
R9037 gnd.n1328 gnd.n1326 585
R9038 gnd.n4010 gnd.n1326 585
R9039 gnd.n3901 gnd.n3900 585
R9040 gnd.n3900 gnd.n3899 585
R9041 gnd.n1330 gnd.n1225 585
R9042 gnd.n4124 gnd.n1225 585
R9043 gnd.n3889 gnd.n3888 585
R9044 gnd.n3890 gnd.n3889 585
R9045 gnd.n1335 gnd.n1213 585
R9046 gnd.n4130 gnd.n1213 585
R9047 gnd.n3703 gnd.n3702 585
R9048 gnd.n3704 gnd.n3703 585
R9049 gnd.n3617 gnd.n1403 585
R9050 gnd.n1410 gnd.n1403 585
R9051 gnd.n3616 gnd.n3615 585
R9052 gnd.n3615 gnd.n3614 585
R9053 gnd.n1406 gnd.n1405 585
R9054 gnd.n3388 gnd.n1406 585
R9055 gnd.n3377 gnd.n1455 585
R9056 gnd.n1455 gnd.n1449 585
R9057 gnd.n3379 gnd.n3378 585
R9058 gnd.n3380 gnd.n3379 585
R9059 gnd.n3376 gnd.n1454 585
R9060 gnd.n3371 gnd.n1454 585
R9061 gnd.n3375 gnd.n3374 585
R9062 gnd.n3374 gnd.n3373 585
R9063 gnd.n1457 gnd.n1456 585
R9064 gnd.n3358 gnd.n1457 585
R9065 gnd.n3333 gnd.n3332 585
R9066 gnd.n3332 gnd.n1468 585
R9067 gnd.n3334 gnd.n1477 585
R9068 gnd.n3347 gnd.n1477 585
R9069 gnd.n3335 gnd.n1487 585
R9070 gnd.n1487 gnd.n1476 585
R9071 gnd.n3337 gnd.n3336 585
R9072 gnd.n3338 gnd.n3337 585
R9073 gnd.n3331 gnd.n1486 585
R9074 gnd.n3326 gnd.n1486 585
R9075 gnd.n3330 gnd.n3329 585
R9076 gnd.n3329 gnd.n3328 585
R9077 gnd.n1489 gnd.n1488 585
R9078 gnd.n3312 gnd.n1489 585
R9079 gnd.n3301 gnd.n1504 585
R9080 gnd.n1504 gnd.n1498 585
R9081 gnd.n3303 gnd.n3302 585
R9082 gnd.n3304 gnd.n3303 585
R9083 gnd.n3300 gnd.n1503 585
R9084 gnd.n1510 gnd.n1503 585
R9085 gnd.n3299 gnd.n3298 585
R9086 gnd.n3298 gnd.n3297 585
R9087 gnd.n1506 gnd.n1505 585
R9088 gnd.n3177 gnd.n1506 585
R9089 gnd.n3284 gnd.n3283 585
R9090 gnd.n3285 gnd.n3284 585
R9091 gnd.n3282 gnd.n1521 585
R9092 gnd.n1521 gnd.n1517 585
R9093 gnd.n3281 gnd.n3280 585
R9094 gnd.n3280 gnd.n3279 585
R9095 gnd.n1523 gnd.n1522 585
R9096 gnd.n3186 gnd.n1523 585
R9097 gnd.n3253 gnd.n3252 585
R9098 gnd.n3254 gnd.n3253 585
R9099 gnd.n3251 gnd.n1534 585
R9100 gnd.n1534 gnd.n1531 585
R9101 gnd.n3250 gnd.n3249 585
R9102 gnd.n3249 gnd.n3248 585
R9103 gnd.n1536 gnd.n1535 585
R9104 gnd.n3193 gnd.n1536 585
R9105 gnd.n3233 gnd.n3232 585
R9106 gnd.n3234 gnd.n3233 585
R9107 gnd.n3231 gnd.n1547 585
R9108 gnd.n3226 gnd.n1547 585
R9109 gnd.n3230 gnd.n3229 585
R9110 gnd.n3229 gnd.n3228 585
R9111 gnd.n1549 gnd.n1548 585
R9112 gnd.n1561 gnd.n1549 585
R9113 gnd.n3163 gnd.n3162 585
R9114 gnd.n3163 gnd.n1560 585
R9115 gnd.n3167 gnd.n3166 585
R9116 gnd.n3166 gnd.n3165 585
R9117 gnd.n3168 gnd.n1567 585
R9118 gnd.n3206 gnd.n1567 585
R9119 gnd.n3169 gnd.n1576 585
R9120 gnd.n3094 gnd.n1576 585
R9121 gnd.n3171 gnd.n3170 585
R9122 gnd.n3172 gnd.n3171 585
R9123 gnd.n3161 gnd.n1575 585
R9124 gnd.n3155 gnd.n1575 585
R9125 gnd.n3160 gnd.n3159 585
R9126 gnd.n3159 gnd.n3158 585
R9127 gnd.n1578 gnd.n1577 585
R9128 gnd.n3144 gnd.n1578 585
R9129 gnd.n3134 gnd.n1595 585
R9130 gnd.n1595 gnd.n1587 585
R9131 gnd.n3136 gnd.n3135 585
R9132 gnd.n3137 gnd.n3136 585
R9133 gnd.n3133 gnd.n1594 585
R9134 gnd.n1599 gnd.n1594 585
R9135 gnd.n3132 gnd.n3131 585
R9136 gnd.n3131 gnd.n3130 585
R9137 gnd.n1597 gnd.n1596 585
R9138 gnd.n3085 gnd.n1597 585
R9139 gnd.n3118 gnd.n3117 585
R9140 gnd.n3119 gnd.n3118 585
R9141 gnd.n3116 gnd.n1610 585
R9142 gnd.n1610 gnd.n1606 585
R9143 gnd.n3115 gnd.n3114 585
R9144 gnd.n3114 gnd.n3113 585
R9145 gnd.n1612 gnd.n1611 585
R9146 gnd.n3075 gnd.n1612 585
R9147 gnd.n3060 gnd.n3059 585
R9148 gnd.n3059 gnd.n1622 585
R9149 gnd.n3061 gnd.n1632 585
R9150 gnd.n3044 gnd.n1632 585
R9151 gnd.n3063 gnd.n3062 585
R9152 gnd.n3064 gnd.n3063 585
R9153 gnd.n3058 gnd.n1631 585
R9154 gnd.n1631 gnd.n1628 585
R9155 gnd.n3057 gnd.n3056 585
R9156 gnd.n3056 gnd.n3055 585
R9157 gnd.n1634 gnd.n1633 585
R9158 gnd.n3035 gnd.n1634 585
R9159 gnd.n3020 gnd.n3019 585
R9160 gnd.n3019 gnd.n1645 585
R9161 gnd.n3021 gnd.n1655 585
R9162 gnd.n3008 gnd.n1655 585
R9163 gnd.n3023 gnd.n3022 585
R9164 gnd.n3024 gnd.n3023 585
R9165 gnd.n3018 gnd.n1654 585
R9166 gnd.n1654 gnd.n1651 585
R9167 gnd.n3017 gnd.n3016 585
R9168 gnd.n3016 gnd.n3015 585
R9169 gnd.n1657 gnd.n1656 585
R9170 gnd.n1670 gnd.n1657 585
R9171 gnd.n2992 gnd.n2991 585
R9172 gnd.n2993 gnd.n2992 585
R9173 gnd.n2990 gnd.n1672 585
R9174 gnd.n2985 gnd.n1672 585
R9175 gnd.n2989 gnd.n2988 585
R9176 gnd.n2988 gnd.n2987 585
R9177 gnd.n1674 gnd.n1673 585
R9178 gnd.n2972 gnd.n1674 585
R9179 gnd.n2960 gnd.n1692 585
R9180 gnd.n1692 gnd.n1684 585
R9181 gnd.n2962 gnd.n2961 585
R9182 gnd.n2963 gnd.n2962 585
R9183 gnd.n2959 gnd.n1691 585
R9184 gnd.n2903 gnd.n1691 585
R9185 gnd.n2958 gnd.n2957 585
R9186 gnd.n2957 gnd.n2956 585
R9187 gnd.n1694 gnd.n1693 585
R9188 gnd.n2931 gnd.n1694 585
R9189 gnd.n2944 gnd.n2943 585
R9190 gnd.n2945 gnd.n2944 585
R9191 gnd.n2942 gnd.n1705 585
R9192 gnd.n2937 gnd.n1705 585
R9193 gnd.n2941 gnd.n2940 585
R9194 gnd.n2940 gnd.n2939 585
R9195 gnd.n1707 gnd.n1706 585
R9196 gnd.n2926 gnd.n1707 585
R9197 gnd.n2877 gnd.n2874 585
R9198 gnd.n2877 gnd.n2876 585
R9199 gnd.n2878 gnd.n2873 585
R9200 gnd.n2878 gnd.n1721 585
R9201 gnd.n2880 gnd.n2879 585
R9202 gnd.n2879 gnd.n1720 585
R9203 gnd.n2881 gnd.n1733 585
R9204 gnd.n2861 gnd.n1733 585
R9205 gnd.n2883 gnd.n2882 585
R9206 gnd.n2884 gnd.n2883 585
R9207 gnd.n2872 gnd.n1732 585
R9208 gnd.n2867 gnd.n1732 585
R9209 gnd.n2871 gnd.n2870 585
R9210 gnd.n2870 gnd.n2869 585
R9211 gnd.n1735 gnd.n1734 585
R9212 gnd.n2852 gnd.n1735 585
R9213 gnd.n1757 gnd.n1756 585
R9214 gnd.n2827 gnd.n1757 585
R9215 gnd.n2831 gnd.n2830 585
R9216 gnd.n2830 gnd.n2829 585
R9217 gnd.n2832 gnd.n1746 585
R9218 gnd.n2843 gnd.n1746 585
R9219 gnd.n2833 gnd.n1754 585
R9220 gnd.n1758 gnd.n1754 585
R9221 gnd.n2835 gnd.n2834 585
R9222 gnd.n2836 gnd.n2835 585
R9223 gnd.n1755 gnd.n1753 585
R9224 gnd.n2809 gnd.n1753 585
R9225 gnd.n2795 gnd.n1778 585
R9226 gnd.n1778 gnd.n1768 585
R9227 gnd.n2797 gnd.n2796 585
R9228 gnd.n2798 gnd.n2797 585
R9229 gnd.n2794 gnd.n1777 585
R9230 gnd.n1777 gnd.n1774 585
R9231 gnd.n2793 gnd.n2792 585
R9232 gnd.n2792 gnd.n2791 585
R9233 gnd.n1780 gnd.n1779 585
R9234 gnd.n1863 gnd.n1780 585
R9235 gnd.n2778 gnd.n2777 585
R9236 gnd.n2779 gnd.n2778 585
R9237 gnd.n2776 gnd.n1792 585
R9238 gnd.n1792 gnd.n1789 585
R9239 gnd.n2774 gnd.n2773 585
R9240 gnd.n1814 gnd.n1813 585
R9241 gnd.n2770 gnd.n2769 585
R9242 gnd.n2771 gnd.n2770 585
R9243 gnd.n2768 gnd.n1850 585
R9244 gnd.n2767 gnd.n2766 585
R9245 gnd.n2765 gnd.n2764 585
R9246 gnd.n2763 gnd.n2762 585
R9247 gnd.n2761 gnd.n2760 585
R9248 gnd.n2759 gnd.n2758 585
R9249 gnd.n2757 gnd.n2756 585
R9250 gnd.n2755 gnd.n2754 585
R9251 gnd.n2753 gnd.n2752 585
R9252 gnd.n2751 gnd.n2750 585
R9253 gnd.n2749 gnd.n2748 585
R9254 gnd.n2747 gnd.n2746 585
R9255 gnd.n2745 gnd.n2744 585
R9256 gnd.n2743 gnd.n2742 585
R9257 gnd.n2741 gnd.n2740 585
R9258 gnd.n2739 gnd.n2738 585
R9259 gnd.n2737 gnd.n2736 585
R9260 gnd.n2735 gnd.n2734 585
R9261 gnd.n2733 gnd.n2732 585
R9262 gnd.n2731 gnd.n2730 585
R9263 gnd.n2729 gnd.n2728 585
R9264 gnd.n2727 gnd.n2726 585
R9265 gnd.n2725 gnd.n2724 585
R9266 gnd.n2723 gnd.n2722 585
R9267 gnd.n2721 gnd.n2720 585
R9268 gnd.n2719 gnd.n2718 585
R9269 gnd.n2717 gnd.n2716 585
R9270 gnd.n2715 gnd.n2714 585
R9271 gnd.n2713 gnd.n2712 585
R9272 gnd.n2711 gnd.n2710 585
R9273 gnd.n2709 gnd.n1932 585
R9274 gnd.n1931 gnd.n1930 585
R9275 gnd.n1929 gnd.n1928 585
R9276 gnd.n1926 gnd.n1925 585
R9277 gnd.n1924 gnd.n1923 585
R9278 gnd.n1922 gnd.n1921 585
R9279 gnd.n1920 gnd.n1919 585
R9280 gnd.n1918 gnd.n1917 585
R9281 gnd.n1916 gnd.n1915 585
R9282 gnd.n1914 gnd.n1913 585
R9283 gnd.n1912 gnd.n1911 585
R9284 gnd.n1910 gnd.n1909 585
R9285 gnd.n1908 gnd.n1907 585
R9286 gnd.n1906 gnd.n1905 585
R9287 gnd.n1904 gnd.n1903 585
R9288 gnd.n1902 gnd.n1901 585
R9289 gnd.n1900 gnd.n1899 585
R9290 gnd.n1898 gnd.n1897 585
R9291 gnd.n1896 gnd.n1895 585
R9292 gnd.n1894 gnd.n1893 585
R9293 gnd.n1892 gnd.n1891 585
R9294 gnd.n1890 gnd.n1889 585
R9295 gnd.n1888 gnd.n1887 585
R9296 gnd.n1886 gnd.n1885 585
R9297 gnd.n1884 gnd.n1883 585
R9298 gnd.n1882 gnd.n1881 585
R9299 gnd.n1880 gnd.n1879 585
R9300 gnd.n1878 gnd.n1877 585
R9301 gnd.n1876 gnd.n1875 585
R9302 gnd.n1874 gnd.n1873 585
R9303 gnd.n1872 gnd.n1871 585
R9304 gnd.n1870 gnd.n1869 585
R9305 gnd.n3707 gnd.n3706 585
R9306 gnd.n3709 gnd.n3708 585
R9307 gnd.n3711 gnd.n3710 585
R9308 gnd.n3713 gnd.n3712 585
R9309 gnd.n3715 gnd.n3714 585
R9310 gnd.n3717 gnd.n3716 585
R9311 gnd.n3719 gnd.n3718 585
R9312 gnd.n3721 gnd.n3720 585
R9313 gnd.n3723 gnd.n3722 585
R9314 gnd.n3725 gnd.n3724 585
R9315 gnd.n3727 gnd.n3726 585
R9316 gnd.n3729 gnd.n3728 585
R9317 gnd.n3731 gnd.n3730 585
R9318 gnd.n3733 gnd.n3732 585
R9319 gnd.n3735 gnd.n3734 585
R9320 gnd.n3737 gnd.n3736 585
R9321 gnd.n3739 gnd.n3738 585
R9322 gnd.n3741 gnd.n3740 585
R9323 gnd.n3743 gnd.n3742 585
R9324 gnd.n3745 gnd.n3744 585
R9325 gnd.n3747 gnd.n3746 585
R9326 gnd.n3749 gnd.n3748 585
R9327 gnd.n3751 gnd.n3750 585
R9328 gnd.n3753 gnd.n3752 585
R9329 gnd.n3755 gnd.n3754 585
R9330 gnd.n3757 gnd.n3756 585
R9331 gnd.n3759 gnd.n3758 585
R9332 gnd.n3761 gnd.n3760 585
R9333 gnd.n3763 gnd.n3762 585
R9334 gnd.n3765 gnd.n1397 585
R9335 gnd.n3767 gnd.n3766 585
R9336 gnd.n3769 gnd.n1361 585
R9337 gnd.n3771 gnd.n3770 585
R9338 gnd.n3774 gnd.n3773 585
R9339 gnd.n1364 gnd.n1362 585
R9340 gnd.n3640 gnd.n3639 585
R9341 gnd.n3642 gnd.n3641 585
R9342 gnd.n3645 gnd.n3644 585
R9343 gnd.n3647 gnd.n3646 585
R9344 gnd.n3649 gnd.n3648 585
R9345 gnd.n3651 gnd.n3650 585
R9346 gnd.n3653 gnd.n3652 585
R9347 gnd.n3655 gnd.n3654 585
R9348 gnd.n3657 gnd.n3656 585
R9349 gnd.n3659 gnd.n3658 585
R9350 gnd.n3661 gnd.n3660 585
R9351 gnd.n3663 gnd.n3662 585
R9352 gnd.n3665 gnd.n3664 585
R9353 gnd.n3667 gnd.n3666 585
R9354 gnd.n3669 gnd.n3668 585
R9355 gnd.n3671 gnd.n3670 585
R9356 gnd.n3673 gnd.n3672 585
R9357 gnd.n3675 gnd.n3674 585
R9358 gnd.n3677 gnd.n3676 585
R9359 gnd.n3679 gnd.n3678 585
R9360 gnd.n3681 gnd.n3680 585
R9361 gnd.n3683 gnd.n3682 585
R9362 gnd.n3685 gnd.n3684 585
R9363 gnd.n3687 gnd.n3686 585
R9364 gnd.n3689 gnd.n3688 585
R9365 gnd.n3691 gnd.n3690 585
R9366 gnd.n3693 gnd.n3692 585
R9367 gnd.n3695 gnd.n3694 585
R9368 gnd.n3697 gnd.n3696 585
R9369 gnd.n3699 gnd.n3698 585
R9370 gnd.n3700 gnd.n1404 585
R9371 gnd.n3705 gnd.n1400 585
R9372 gnd.n3705 gnd.n3704 585
R9373 gnd.n3384 gnd.n1401 585
R9374 gnd.n1410 gnd.n1401 585
R9375 gnd.n3385 gnd.n1408 585
R9376 gnd.n3614 gnd.n1408 585
R9377 gnd.n3387 gnd.n3386 585
R9378 gnd.n3388 gnd.n3387 585
R9379 gnd.n3383 gnd.n1450 585
R9380 gnd.n1450 gnd.n1449 585
R9381 gnd.n3382 gnd.n3381 585
R9382 gnd.n3381 gnd.n3380 585
R9383 gnd.n1452 gnd.n1451 585
R9384 gnd.n3371 gnd.n1452 585
R9385 gnd.n3342 gnd.n1459 585
R9386 gnd.n3373 gnd.n1459 585
R9387 gnd.n3343 gnd.n1469 585
R9388 gnd.n3358 gnd.n1469 585
R9389 gnd.n3344 gnd.n1481 585
R9390 gnd.n1481 gnd.n1468 585
R9391 gnd.n3346 gnd.n3345 585
R9392 gnd.n3347 gnd.n3346 585
R9393 gnd.n3341 gnd.n1480 585
R9394 gnd.n1480 gnd.n1476 585
R9395 gnd.n3340 gnd.n3339 585
R9396 gnd.n3339 gnd.n3338 585
R9397 gnd.n1483 gnd.n1482 585
R9398 gnd.n3326 gnd.n1483 585
R9399 gnd.n3308 gnd.n1490 585
R9400 gnd.n3328 gnd.n1490 585
R9401 gnd.n3310 gnd.n3309 585
R9402 gnd.n3312 gnd.n3310 585
R9403 gnd.n3307 gnd.n1500 585
R9404 gnd.n1500 gnd.n1498 585
R9405 gnd.n3306 gnd.n3305 585
R9406 gnd.n3305 gnd.n3304 585
R9407 gnd.n1502 gnd.n1501 585
R9408 gnd.n1510 gnd.n1502 585
R9409 gnd.n3176 gnd.n1508 585
R9410 gnd.n3297 gnd.n1508 585
R9411 gnd.n3179 gnd.n3178 585
R9412 gnd.n3178 gnd.n3177 585
R9413 gnd.n3180 gnd.n1519 585
R9414 gnd.n3285 gnd.n1519 585
R9415 gnd.n3182 gnd.n3181 585
R9416 gnd.n3181 gnd.n1517 585
R9417 gnd.n3183 gnd.n1524 585
R9418 gnd.n3279 gnd.n1524 585
R9419 gnd.n3188 gnd.n3187 585
R9420 gnd.n3187 gnd.n3186 585
R9421 gnd.n3189 gnd.n1532 585
R9422 gnd.n3254 gnd.n1532 585
R9423 gnd.n3191 gnd.n3190 585
R9424 gnd.n3190 gnd.n1531 585
R9425 gnd.n3192 gnd.n1538 585
R9426 gnd.n3248 gnd.n1538 585
R9427 gnd.n3195 gnd.n3194 585
R9428 gnd.n3194 gnd.n3193 585
R9429 gnd.n3196 gnd.n1545 585
R9430 gnd.n3234 gnd.n1545 585
R9431 gnd.n3197 gnd.n1552 585
R9432 gnd.n3226 gnd.n1552 585
R9433 gnd.n3198 gnd.n1551 585
R9434 gnd.n3228 gnd.n1551 585
R9435 gnd.n3200 gnd.n3199 585
R9436 gnd.n3200 gnd.n1561 585
R9437 gnd.n3202 gnd.n3201 585
R9438 gnd.n3201 gnd.n1560 585
R9439 gnd.n3203 gnd.n1570 585
R9440 gnd.n3165 gnd.n1570 585
R9441 gnd.n3205 gnd.n3204 585
R9442 gnd.n3206 gnd.n3205 585
R9443 gnd.n3175 gnd.n1569 585
R9444 gnd.n3094 gnd.n1569 585
R9445 gnd.n3174 gnd.n3173 585
R9446 gnd.n3173 gnd.n3172 585
R9447 gnd.n1572 gnd.n1571 585
R9448 gnd.n3155 gnd.n1572 585
R9449 gnd.n3141 gnd.n1580 585
R9450 gnd.n3158 gnd.n1580 585
R9451 gnd.n3143 gnd.n3142 585
R9452 gnd.n3144 gnd.n3143 585
R9453 gnd.n3140 gnd.n1589 585
R9454 gnd.n1589 gnd.n1587 585
R9455 gnd.n3139 gnd.n3138 585
R9456 gnd.n3138 gnd.n3137 585
R9457 gnd.n1591 gnd.n1590 585
R9458 gnd.n1599 gnd.n1591 585
R9459 gnd.n3082 gnd.n1598 585
R9460 gnd.n3130 gnd.n1598 585
R9461 gnd.n3084 gnd.n3083 585
R9462 gnd.n3085 gnd.n3084 585
R9463 gnd.n3081 gnd.n1608 585
R9464 gnd.n3119 gnd.n1608 585
R9465 gnd.n3080 gnd.n3079 585
R9466 gnd.n3079 gnd.n1606 585
R9467 gnd.n3078 gnd.n1614 585
R9468 gnd.n3113 gnd.n1614 585
R9469 gnd.n3077 gnd.n3076 585
R9470 gnd.n3076 gnd.n3075 585
R9471 gnd.n1621 gnd.n1620 585
R9472 gnd.n1622 gnd.n1621 585
R9473 gnd.n3043 gnd.n3042 585
R9474 gnd.n3044 gnd.n3043 585
R9475 gnd.n3041 gnd.n1629 585
R9476 gnd.n3064 gnd.n1629 585
R9477 gnd.n3040 gnd.n3039 585
R9478 gnd.n3039 gnd.n1628 585
R9479 gnd.n3038 gnd.n1636 585
R9480 gnd.n3055 gnd.n1636 585
R9481 gnd.n3037 gnd.n3036 585
R9482 gnd.n3036 gnd.n3035 585
R9483 gnd.n1644 gnd.n1643 585
R9484 gnd.n1645 gnd.n1644 585
R9485 gnd.n3010 gnd.n3009 585
R9486 gnd.n3009 gnd.n3008 585
R9487 gnd.n3011 gnd.n1652 585
R9488 gnd.n3024 gnd.n1652 585
R9489 gnd.n3012 gnd.n1660 585
R9490 gnd.n1660 gnd.n1651 585
R9491 gnd.n3014 gnd.n3013 585
R9492 gnd.n3015 gnd.n3014 585
R9493 gnd.n1661 gnd.n1659 585
R9494 gnd.n1670 gnd.n1659 585
R9495 gnd.n2967 gnd.n1669 585
R9496 gnd.n2993 gnd.n1669 585
R9497 gnd.n2968 gnd.n1677 585
R9498 gnd.n2985 gnd.n1677 585
R9499 gnd.n2969 gnd.n1676 585
R9500 gnd.n2987 gnd.n1676 585
R9501 gnd.n2971 gnd.n2970 585
R9502 gnd.n2972 gnd.n2971 585
R9503 gnd.n2966 gnd.n1686 585
R9504 gnd.n1686 gnd.n1684 585
R9505 gnd.n2965 gnd.n2964 585
R9506 gnd.n2964 gnd.n2963 585
R9507 gnd.n1688 gnd.n1687 585
R9508 gnd.n2903 gnd.n1688 585
R9509 gnd.n2930 gnd.n1696 585
R9510 gnd.n2956 gnd.n1696 585
R9511 gnd.n2933 gnd.n2932 585
R9512 gnd.n2932 gnd.n2931 585
R9513 gnd.n2934 gnd.n1703 585
R9514 gnd.n2945 gnd.n1703 585
R9515 gnd.n2936 gnd.n2935 585
R9516 gnd.n2937 gnd.n2936 585
R9517 gnd.n2929 gnd.n1709 585
R9518 gnd.n2939 gnd.n1709 585
R9519 gnd.n2928 gnd.n2927 585
R9520 gnd.n2927 gnd.n2926 585
R9521 gnd.n1712 gnd.n1711 585
R9522 gnd.n2876 gnd.n1712 585
R9523 gnd.n2858 gnd.n2857 585
R9524 gnd.n2858 gnd.n1721 585
R9525 gnd.n2859 gnd.n2856 585
R9526 gnd.n2859 gnd.n1720 585
R9527 gnd.n2863 gnd.n2862 585
R9528 gnd.n2862 gnd.n2861 585
R9529 gnd.n2864 gnd.n1730 585
R9530 gnd.n2884 gnd.n1730 585
R9531 gnd.n2866 gnd.n2865 585
R9532 gnd.n2867 gnd.n2866 585
R9533 gnd.n2855 gnd.n1737 585
R9534 gnd.n2869 gnd.n1737 585
R9535 gnd.n2854 gnd.n2853 585
R9536 gnd.n2853 gnd.n2852 585
R9537 gnd.n1739 gnd.n1738 585
R9538 gnd.n2827 gnd.n1739 585
R9539 gnd.n2840 gnd.n1748 585
R9540 gnd.n2829 gnd.n1748 585
R9541 gnd.n2842 gnd.n2841 585
R9542 gnd.n2843 gnd.n2842 585
R9543 gnd.n2839 gnd.n1747 585
R9544 gnd.n1758 gnd.n1747 585
R9545 gnd.n2838 gnd.n2837 585
R9546 gnd.n2837 gnd.n2836 585
R9547 gnd.n1750 gnd.n1749 585
R9548 gnd.n2809 gnd.n1750 585
R9549 gnd.n1857 gnd.n1856 585
R9550 gnd.n1856 gnd.n1768 585
R9551 gnd.n1858 gnd.n1775 585
R9552 gnd.n2798 gnd.n1775 585
R9553 gnd.n1860 gnd.n1859 585
R9554 gnd.n1859 gnd.n1774 585
R9555 gnd.n1861 gnd.n1782 585
R9556 gnd.n2791 gnd.n1782 585
R9557 gnd.n1865 gnd.n1864 585
R9558 gnd.n1864 gnd.n1863 585
R9559 gnd.n1866 gnd.n1790 585
R9560 gnd.n2779 gnd.n1790 585
R9561 gnd.n1868 gnd.n1867 585
R9562 gnd.n1868 gnd.n1789 585
R9563 gnd.n764 gnd.n763 585
R9564 gnd.n957 gnd.n764 585
R9565 gnd.n6635 gnd.n6634 585
R9566 gnd.n6635 gnd.n232 585
R9567 gnd.n6637 gnd.n257 585
R9568 gnd.n6637 gnd.n6636 585
R9569 gnd.n6639 gnd.n6638 585
R9570 gnd.n6638 gnd.n236 585
R9571 gnd.n6640 gnd.n252 585
R9572 gnd.n252 gnd.n246 585
R9573 gnd.n6642 gnd.n6641 585
R9574 gnd.n6643 gnd.n6642 585
R9575 gnd.n253 gnd.n251 585
R9576 gnd.n251 gnd.n248 585
R9577 gnd.n4071 gnd.n4070 585
R9578 gnd.n4070 gnd.n1251 585
R9579 gnd.n4075 gnd.n4069 585
R9580 gnd.n4069 gnd.n1262 585
R9581 gnd.n4076 gnd.n1276 585
R9582 gnd.n1276 gnd.n1260 585
R9583 gnd.n4078 gnd.n4077 585
R9584 gnd.n4079 gnd.n4078 585
R9585 gnd.n1277 gnd.n1275 585
R9586 gnd.n1275 gnd.n1270 585
R9587 gnd.n4064 gnd.n4063 585
R9588 gnd.n4063 gnd.n4062 585
R9589 gnd.n1280 gnd.n1279 585
R9590 gnd.n1291 gnd.n1280 585
R9591 gnd.n4037 gnd.n1304 585
R9592 gnd.n1304 gnd.n1289 585
R9593 gnd.n4039 gnd.n4038 585
R9594 gnd.n4040 gnd.n4039 585
R9595 gnd.n1305 gnd.n1303 585
R9596 gnd.n1303 gnd.n1299 585
R9597 gnd.n4032 gnd.n4031 585
R9598 gnd.n4031 gnd.n4030 585
R9599 gnd.n1308 gnd.n1307 585
R9600 gnd.n1320 gnd.n1308 585
R9601 gnd.n4006 gnd.n3994 585
R9602 gnd.n3994 gnd.n1318 585
R9603 gnd.n4008 gnd.n4007 585
R9604 gnd.n4009 gnd.n4008 585
R9605 gnd.n3995 gnd.n3993 585
R9606 gnd.n3993 gnd.n1325 585
R9607 gnd.n4001 gnd.n4000 585
R9608 gnd.n4000 gnd.n1227 585
R9609 gnd.n3999 gnd.n3998 585
R9610 gnd.n3999 gnd.n1224 585
R9611 gnd.n1211 gnd.n1210 585
R9612 gnd.n1215 gnd.n1211 585
R9613 gnd.n4133 gnd.n4132 585
R9614 gnd.n4132 gnd.n4131 585
R9615 gnd.n4134 gnd.n1205 585
R9616 gnd.n1212 gnd.n1205 585
R9617 gnd.n4136 gnd.n4135 585
R9618 gnd.n4137 gnd.n4136 585
R9619 gnd.n1202 gnd.n1201 585
R9620 gnd.n4138 gnd.n1202 585
R9621 gnd.n4141 gnd.n4140 585
R9622 gnd.n4140 gnd.n4139 585
R9623 gnd.n4142 gnd.n1196 585
R9624 gnd.n1196 gnd.n1194 585
R9625 gnd.n4144 gnd.n4143 585
R9626 gnd.n4145 gnd.n4144 585
R9627 gnd.n1197 gnd.n1195 585
R9628 gnd.n1195 gnd.n1192 585
R9629 gnd.n1434 gnd.n1433 585
R9630 gnd.n3593 gnd.n1434 585
R9631 gnd.n3597 gnd.n3596 585
R9632 gnd.n3596 gnd.n3595 585
R9633 gnd.n3598 gnd.n1424 585
R9634 gnd.n1435 gnd.n1424 585
R9635 gnd.n3600 gnd.n3599 585
R9636 gnd.n3601 gnd.n3600 585
R9637 gnd.n1425 gnd.n1418 585
R9638 gnd.n3603 gnd.n1418 585
R9639 gnd.n3606 gnd.n1417 585
R9640 gnd.n3606 gnd.n3605 585
R9641 gnd.n3608 gnd.n3607 585
R9642 gnd.n3607 gnd.n1365 585
R9643 gnd.n3609 gnd.n1412 585
R9644 gnd.n1412 gnd.n1402 585
R9645 gnd.n3611 gnd.n3610 585
R9646 gnd.n3612 gnd.n3611 585
R9647 gnd.n1413 gnd.n1411 585
R9648 gnd.n1411 gnd.n1407 585
R9649 gnd.n3367 gnd.n1463 585
R9650 gnd.n1463 gnd.n1462 585
R9651 gnd.n3369 gnd.n3368 585
R9652 gnd.n3370 gnd.n3369 585
R9653 gnd.n1464 gnd.n1461 585
R9654 gnd.n1461 gnd.n1458 585
R9655 gnd.n3361 gnd.n3360 585
R9656 gnd.n3360 gnd.n3359 585
R9657 gnd.n1467 gnd.n1466 585
R9658 gnd.n3347 gnd.n1467 585
R9659 gnd.n3322 gnd.n1493 585
R9660 gnd.n1493 gnd.n1485 585
R9661 gnd.n3324 gnd.n3323 585
R9662 gnd.n3325 gnd.n3324 585
R9663 gnd.n1494 gnd.n1492 585
R9664 gnd.n3311 gnd.n1492 585
R9665 gnd.n3317 gnd.n3316 585
R9666 gnd.n3316 gnd.n3315 585
R9667 gnd.n1497 gnd.n1496 585
R9668 gnd.n1509 gnd.n1497 585
R9669 gnd.n3295 gnd.n3294 585
R9670 gnd.n3296 gnd.n3295 585
R9671 gnd.n1513 gnd.n1512 585
R9672 gnd.n1520 gnd.n1512 585
R9673 gnd.n3290 gnd.n3289 585
R9674 gnd.n3289 gnd.n3288 585
R9675 gnd.n1516 gnd.n1515 585
R9676 gnd.n3184 gnd.n1516 585
R9677 gnd.n3242 gnd.n1540 585
R9678 gnd.n1540 gnd.n1533 585
R9679 gnd.n3244 gnd.n3243 585
R9680 gnd.n3245 gnd.n3244 585
R9681 gnd.n1541 gnd.n1539 585
R9682 gnd.n1539 gnd.n1537 585
R9683 gnd.n3237 gnd.n3236 585
R9684 gnd.n3236 gnd.n3235 585
R9685 gnd.n1544 gnd.n1543 585
R9686 gnd.n3227 gnd.n1544 585
R9687 gnd.n3213 gnd.n3212 585
R9688 gnd.n3214 gnd.n3213 585
R9689 gnd.n1563 gnd.n1562 585
R9690 gnd.n3164 gnd.n1562 585
R9691 gnd.n3208 gnd.n3207 585
R9692 gnd.n3207 gnd.n3206 585
R9693 gnd.n1566 gnd.n1565 585
R9694 gnd.n1574 gnd.n1566 585
R9695 gnd.n3153 gnd.n3152 585
R9696 gnd.n3154 gnd.n3153 585
R9697 gnd.n1583 gnd.n1582 585
R9698 gnd.n1582 gnd.n1579 585
R9699 gnd.n3148 gnd.n3147 585
R9700 gnd.n3147 gnd.n3146 585
R9701 gnd.n1586 gnd.n1585 585
R9702 gnd.n1592 gnd.n1586 585
R9703 gnd.n3128 gnd.n3127 585
R9704 gnd.n3129 gnd.n3128 585
R9705 gnd.n1602 gnd.n1601 585
R9706 gnd.n1609 gnd.n1601 585
R9707 gnd.n3123 gnd.n3122 585
R9708 gnd.n3122 gnd.n3121 585
R9709 gnd.n1605 gnd.n1604 585
R9710 gnd.n1613 gnd.n1605 585
R9711 gnd.n3072 gnd.n3071 585
R9712 gnd.n3073 gnd.n3072 585
R9713 gnd.n1624 gnd.n1623 585
R9714 gnd.n1642 gnd.n1623 585
R9715 gnd.n3067 gnd.n3066 585
R9716 gnd.n3066 gnd.n3065 585
R9717 gnd.n1627 gnd.n1626 585
R9718 gnd.n1635 gnd.n1627 585
R9719 gnd.n3032 gnd.n3031 585
R9720 gnd.n3033 gnd.n3032 585
R9721 gnd.n1647 gnd.n1646 585
R9722 gnd.n1662 gnd.n1646 585
R9723 gnd.n3027 gnd.n3026 585
R9724 gnd.n3026 gnd.n3025 585
R9725 gnd.n1650 gnd.n1649 585
R9726 gnd.n3015 gnd.n1650 585
R9727 gnd.n2981 gnd.n1679 585
R9728 gnd.n1679 gnd.n1671 585
R9729 gnd.n2983 gnd.n2982 585
R9730 gnd.n2984 gnd.n2983 585
R9731 gnd.n1680 gnd.n1678 585
R9732 gnd.n1678 gnd.n1675 585
R9733 gnd.n2976 gnd.n2975 585
R9734 gnd.n2975 gnd.n2974 585
R9735 gnd.n1683 gnd.n1682 585
R9736 gnd.n1689 gnd.n1683 585
R9737 gnd.n2954 gnd.n2953 585
R9738 gnd.n2955 gnd.n2954 585
R9739 gnd.n1698 gnd.n1697 585
R9740 gnd.n1704 gnd.n1697 585
R9741 gnd.n2949 gnd.n2948 585
R9742 gnd.n2948 gnd.n2947 585
R9743 gnd.n1701 gnd.n1700 585
R9744 gnd.n1708 gnd.n1701 585
R9745 gnd.n2892 gnd.n1723 585
R9746 gnd.n1723 gnd.n1713 585
R9747 gnd.n2894 gnd.n2893 585
R9748 gnd.n2895 gnd.n2894 585
R9749 gnd.n1724 gnd.n1722 585
R9750 gnd.n2860 gnd.n1722 585
R9751 gnd.n2887 gnd.n2886 585
R9752 gnd.n2886 gnd.n2885 585
R9753 gnd.n1727 gnd.n1726 585
R9754 gnd.n2868 gnd.n1727 585
R9755 gnd.n2850 gnd.n2849 585
R9756 gnd.n2851 gnd.n2850 585
R9757 gnd.n1742 gnd.n1741 585
R9758 gnd.n2828 gnd.n1741 585
R9759 gnd.n2845 gnd.n2844 585
R9760 gnd.n2844 gnd.n2843 585
R9761 gnd.n1745 gnd.n1744 585
R9762 gnd.n1752 gnd.n1745 585
R9763 gnd.n2807 gnd.n2806 585
R9764 gnd.n2808 gnd.n2807 585
R9765 gnd.n1770 gnd.n1769 585
R9766 gnd.n1776 gnd.n1769 585
R9767 gnd.n2802 gnd.n2801 585
R9768 gnd.n2801 gnd.n2800 585
R9769 gnd.n1773 gnd.n1772 585
R9770 gnd.n1781 gnd.n1773 585
R9771 gnd.n2615 gnd.n2614 585
R9772 gnd.n2615 gnd.n1791 585
R9773 gnd.n2619 gnd.n2618 585
R9774 gnd.n2618 gnd.n2617 585
R9775 gnd.n2620 gnd.n2063 585
R9776 gnd.n2063 gnd.n1849 585
R9777 gnd.n2622 gnd.n2621 585
R9778 gnd.n2623 gnd.n2622 585
R9779 gnd.n2064 gnd.n2062 585
R9780 gnd.n2062 gnd.n2061 585
R9781 gnd.n2607 gnd.n2606 585
R9782 gnd.n2606 gnd.n2605 585
R9783 gnd.n2067 gnd.n2066 585
R9784 gnd.n2602 gnd.n2067 585
R9785 gnd.n2597 gnd.n2596 585
R9786 gnd.n2598 gnd.n2597 585
R9787 gnd.n2070 gnd.n2069 585
R9788 gnd.n2588 gnd.n2069 585
R9789 gnd.n2592 gnd.n2591 585
R9790 gnd.n2591 gnd.n2590 585
R9791 gnd.n2073 gnd.n2072 585
R9792 gnd.n2586 gnd.n2073 585
R9793 gnd.n2584 gnd.n2583 585
R9794 gnd.n2585 gnd.n2584 585
R9795 gnd.n2208 gnd.n2207 585
R9796 gnd.n2576 gnd.n2207 585
R9797 gnd.n2579 gnd.n2578 585
R9798 gnd.n2578 gnd.n2577 585
R9799 gnd.n2574 gnd.n2210 585
R9800 gnd.n2575 gnd.n2574 585
R9801 gnd.n2573 gnd.n2571 585
R9802 gnd.n2573 gnd.n2572 585
R9803 gnd.n2212 gnd.n2211 585
R9804 gnd.n2211 gnd.n1082 585
R9805 gnd.n2567 gnd.n2566 585
R9806 gnd.n2566 gnd.n1079 585
R9807 gnd.n2565 gnd.n2214 585
R9808 gnd.n2565 gnd.n1072 585
R9809 gnd.n2564 gnd.n2563 585
R9810 gnd.n2564 gnd.n1069 585
R9811 gnd.n2216 gnd.n2215 585
R9812 gnd.n2215 gnd.n1061 585
R9813 gnd.n2559 gnd.n2558 585
R9814 gnd.n2558 gnd.n1058 585
R9815 gnd.n2557 gnd.n2218 585
R9816 gnd.n2557 gnd.n1050 585
R9817 gnd.n2556 gnd.n2220 585
R9818 gnd.n2556 gnd.n2555 585
R9819 gnd.n2489 gnd.n2219 585
R9820 gnd.n2219 gnd.n1040 585
R9821 gnd.n2491 gnd.n2490 585
R9822 gnd.n2490 gnd.n1037 585
R9823 gnd.n2492 gnd.n2482 585
R9824 gnd.n2482 gnd.n1029 585
R9825 gnd.n2494 gnd.n2493 585
R9826 gnd.n2494 gnd.n1026 585
R9827 gnd.n2495 gnd.n2481 585
R9828 gnd.n2495 gnd.n2235 585
R9829 gnd.n2497 gnd.n2496 585
R9830 gnd.n2496 gnd.n1016 585
R9831 gnd.n2498 gnd.n2244 585
R9832 gnd.n2244 gnd.n1008 585
R9833 gnd.n2500 gnd.n2499 585
R9834 gnd.n2501 gnd.n2500 585
R9835 gnd.n2245 gnd.n2243 585
R9836 gnd.n2243 gnd.n998 585
R9837 gnd.n2475 gnd.n2474 585
R9838 gnd.n2474 gnd.n995 585
R9839 gnd.n2473 gnd.n2247 585
R9840 gnd.n2473 gnd.n990 585
R9841 gnd.n2472 gnd.n2471 585
R9842 gnd.n2472 gnd.n987 585
R9843 gnd.n2456 gnd.n2455 585
R9844 gnd.n2455 gnd.n2454 585
R9845 gnd.n2466 gnd.n2465 585
R9846 gnd.n2465 gnd.n978 585
R9847 gnd.n2464 gnd.n2458 585
R9848 gnd.n2464 gnd.n973 585
R9849 gnd.n2463 gnd.n2461 585
R9850 gnd.n2463 gnd.n2462 585
R9851 gnd.n4148 gnd.n4147 585
R9852 gnd.n4147 gnd.n4146 585
R9853 gnd.n4149 gnd.n1189 585
R9854 gnd.n3592 gnd.n1189 585
R9855 gnd.n4150 gnd.n1188 585
R9856 gnd.n3594 gnd.n1188 585
R9857 gnd.n1436 gnd.n1186 585
R9858 gnd.n1437 gnd.n1436 585
R9859 gnd.n4154 gnd.n1185 585
R9860 gnd.n1423 gnd.n1185 585
R9861 gnd.n4155 gnd.n1184 585
R9862 gnd.n3602 gnd.n1184 585
R9863 gnd.n4156 gnd.n1183 585
R9864 gnd.n3604 gnd.n1183 585
R9865 gnd.n1419 gnd.n1181 585
R9866 gnd.n1420 gnd.n1419 585
R9867 gnd.n4160 gnd.n1180 585
R9868 gnd.n3399 gnd.n1180 585
R9869 gnd.n4161 gnd.n1179 585
R9870 gnd.n3397 gnd.n1179 585
R9871 gnd.n4162 gnd.n1178 585
R9872 gnd.n3613 gnd.n1178 585
R9873 gnd.n3389 gnd.n1176 585
R9874 gnd.n3390 gnd.n3389 585
R9875 gnd.n4166 gnd.n1175 585
R9876 gnd.n1453 gnd.n1175 585
R9877 gnd.n4167 gnd.n1174 585
R9878 gnd.n3372 gnd.n1174 585
R9879 gnd.n4168 gnd.n1173 585
R9880 gnd.n3357 gnd.n1173 585
R9881 gnd.n1478 gnd.n1171 585
R9882 gnd.n1479 gnd.n1478 585
R9883 gnd.n4172 gnd.n1170 585
R9884 gnd.n3348 gnd.n1170 585
R9885 gnd.n4173 gnd.n1169 585
R9886 gnd.n1484 gnd.n1169 585
R9887 gnd.n4174 gnd.n1168 585
R9888 gnd.n3327 gnd.n1168 585
R9889 gnd.n3313 gnd.n1166 585
R9890 gnd.n3314 gnd.n3313 585
R9891 gnd.n4178 gnd.n1165 585
R9892 gnd.n3263 gnd.n1165 585
R9893 gnd.n4179 gnd.n1164 585
R9894 gnd.n1511 gnd.n1164 585
R9895 gnd.n4180 gnd.n1163 585
R9896 gnd.n1507 gnd.n1163 585
R9897 gnd.n3286 gnd.n1161 585
R9898 gnd.n3287 gnd.n3286 585
R9899 gnd.n4184 gnd.n1160 585
R9900 gnd.n3278 gnd.n1160 585
R9901 gnd.n4185 gnd.n1159 585
R9902 gnd.n3185 gnd.n1159 585
R9903 gnd.n4186 gnd.n1158 585
R9904 gnd.n3255 gnd.n1158 585
R9905 gnd.n3246 gnd.n1156 585
R9906 gnd.n3247 gnd.n3246 585
R9907 gnd.n4190 gnd.n1155 585
R9908 gnd.n1546 gnd.n1155 585
R9909 gnd.n4191 gnd.n1154 585
R9910 gnd.n3225 gnd.n1154 585
R9911 gnd.n4192 gnd.n1153 585
R9912 gnd.n1550 gnd.n1153 585
R9913 gnd.n3215 gnd.n1151 585
R9914 gnd.n3216 gnd.n3215 585
R9915 gnd.n4196 gnd.n1150 585
R9916 gnd.n1568 gnd.n1150 585
R9917 gnd.n4197 gnd.n1149 585
R9918 gnd.n3095 gnd.n1149 585
R9919 gnd.n4198 gnd.n1148 585
R9920 gnd.n1573 gnd.n1148 585
R9921 gnd.n3156 gnd.n1146 585
R9922 gnd.n3157 gnd.n3156 585
R9923 gnd.n4202 gnd.n1145 585
R9924 gnd.n3145 gnd.n1145 585
R9925 gnd.n4203 gnd.n1144 585
R9926 gnd.n1593 gnd.n1144 585
R9927 gnd.n4204 gnd.n1143 585
R9928 gnd.n1600 gnd.n1143 585
R9929 gnd.n3086 gnd.n1141 585
R9930 gnd.n3087 gnd.n3086 585
R9931 gnd.n4208 gnd.n1140 585
R9932 gnd.n3120 gnd.n1140 585
R9933 gnd.n4209 gnd.n1139 585
R9934 gnd.n3112 gnd.n1139 585
R9935 gnd.n4210 gnd.n1138 585
R9936 gnd.n3074 gnd.n1138 585
R9937 gnd.n3045 gnd.n1136 585
R9938 gnd.n3046 gnd.n3045 585
R9939 gnd.n4214 gnd.n1135 585
R9940 gnd.n1630 gnd.n1135 585
R9941 gnd.n4215 gnd.n1134 585
R9942 gnd.n3054 gnd.n1134 585
R9943 gnd.n4216 gnd.n1133 585
R9944 gnd.n3034 gnd.n1133 585
R9945 gnd.n3006 gnd.n1131 585
R9946 gnd.n3007 gnd.n3006 585
R9947 gnd.n4220 gnd.n1130 585
R9948 gnd.n1653 gnd.n1130 585
R9949 gnd.n4221 gnd.n1129 585
R9950 gnd.n2998 gnd.n1129 585
R9951 gnd.n4222 gnd.n1128 585
R9952 gnd.n1658 gnd.n1128 585
R9953 gnd.n2994 gnd.n1126 585
R9954 gnd.n2995 gnd.n2994 585
R9955 gnd.n4226 gnd.n1125 585
R9956 gnd.n2986 gnd.n1125 585
R9957 gnd.n4227 gnd.n1124 585
R9958 gnd.n2973 gnd.n1124 585
R9959 gnd.n4228 gnd.n1123 585
R9960 gnd.n1690 gnd.n1123 585
R9961 gnd.n2904 gnd.n1121 585
R9962 gnd.n2905 gnd.n2904 585
R9963 gnd.n4232 gnd.n1120 585
R9964 gnd.n1695 gnd.n1120 585
R9965 gnd.n4233 gnd.n1119 585
R9966 gnd.n2946 gnd.n1119 585
R9967 gnd.n4234 gnd.n1118 585
R9968 gnd.n2938 gnd.n1118 585
R9969 gnd.n2924 gnd.n1116 585
R9970 gnd.n2925 gnd.n2924 585
R9971 gnd.n4238 gnd.n1115 585
R9972 gnd.n2875 gnd.n1115 585
R9973 gnd.n4239 gnd.n1114 585
R9974 gnd.n2896 gnd.n1114 585
R9975 gnd.n4240 gnd.n1113 585
R9976 gnd.n1731 gnd.n1113 585
R9977 gnd.n1728 gnd.n1111 585
R9978 gnd.n1729 gnd.n1728 585
R9979 gnd.n4244 gnd.n1110 585
R9980 gnd.n1736 gnd.n1110 585
R9981 gnd.n4245 gnd.n1109 585
R9982 gnd.n1740 gnd.n1109 585
R9983 gnd.n4246 gnd.n1108 585
R9984 gnd.n2826 gnd.n1108 585
R9985 gnd.n1759 gnd.n1106 585
R9986 gnd.n1760 gnd.n1759 585
R9987 gnd.n4250 gnd.n1105 585
R9988 gnd.n1751 gnd.n1105 585
R9989 gnd.n4251 gnd.n1104 585
R9990 gnd.n2810 gnd.n1104 585
R9991 gnd.n4252 gnd.n1103 585
R9992 gnd.n2799 gnd.n1103 585
R9993 gnd.n2789 gnd.n1101 585
R9994 gnd.n2790 gnd.n2789 585
R9995 gnd.n4256 gnd.n1100 585
R9996 gnd.n1862 gnd.n1100 585
R9997 gnd.n4257 gnd.n1099 585
R9998 gnd.n2780 gnd.n1099 585
R9999 gnd.n4258 gnd.n1098 585
R10000 gnd.n2616 gnd.n1098 585
R10001 gnd.n1815 gnd.n1096 585
R10002 gnd.n1816 gnd.n1815 585
R10003 gnd.n4262 gnd.n1095 585
R10004 gnd.n2624 gnd.n1095 585
R10005 gnd.n4263 gnd.n1094 585
R10006 gnd.n2604 gnd.n1094 585
R10007 gnd.n4264 gnd.n1093 585
R10008 gnd.n2603 gnd.n1093 585
R10009 gnd.n2600 gnd.n1091 585
R10010 gnd.n2601 gnd.n2600 585
R10011 gnd.n4268 gnd.n1090 585
R10012 gnd.n2068 gnd.n1090 585
R10013 gnd.n4269 gnd.n1089 585
R10014 gnd.n2589 gnd.n1089 585
R10015 gnd.n4270 gnd.n1088 585
R10016 gnd.n2587 gnd.n1088 585
R10017 gnd.n2204 gnd.n2203 585
R10018 gnd.n2202 gnd.n2090 585
R10019 gnd.n2092 gnd.n2089 585
R10020 gnd.n2206 gnd.n2089 585
R10021 gnd.n2195 gnd.n2105 585
R10022 gnd.n2194 gnd.n2106 585
R10023 gnd.n2108 gnd.n2107 585
R10024 gnd.n2187 gnd.n2116 585
R10025 gnd.n2186 gnd.n2117 585
R10026 gnd.n2127 gnd.n2118 585
R10027 gnd.n2179 gnd.n2128 585
R10028 gnd.n2178 gnd.n2129 585
R10029 gnd.n2131 gnd.n2130 585
R10030 gnd.n2171 gnd.n2139 585
R10031 gnd.n2170 gnd.n2140 585
R10032 gnd.n2152 gnd.n2141 585
R10033 gnd.n2163 gnd.n2153 585
R10034 gnd.n2162 gnd.n2155 585
R10035 gnd.n2154 gnd.n2036 585
R10036 gnd.n2655 gnd.n2037 585
R10037 gnd.n2654 gnd.n2038 585
R10038 gnd.n2653 gnd.n2039 585
R10039 gnd.n2083 gnd.n2040 585
R10040 gnd.n2649 gnd.n2042 585
R10041 gnd.n2648 gnd.n2043 585
R10042 gnd.n2647 gnd.n2044 585
R10043 gnd.n2644 gnd.n2049 585
R10044 gnd.n2643 gnd.n2050 585
R10045 gnd.n2642 gnd.n2051 585
R10046 gnd.n2087 gnd.n2052 585
R10047 gnd.n1440 gnd.n1193 585
R10048 gnd.n4146 gnd.n1193 585
R10049 gnd.n3591 gnd.n3590 585
R10050 gnd.n3592 gnd.n3591 585
R10051 gnd.n1439 gnd.n1438 585
R10052 gnd.n3594 gnd.n1438 585
R10053 gnd.n3410 gnd.n3409 585
R10054 gnd.n3409 gnd.n1437 585
R10055 gnd.n3408 gnd.n3407 585
R10056 gnd.n3408 gnd.n1423 585
R10057 gnd.n3406 gnd.n1422 585
R10058 gnd.n3602 gnd.n1422 585
R10059 gnd.n1442 gnd.n1421 585
R10060 gnd.n3604 gnd.n1421 585
R10061 gnd.n3402 gnd.n3401 585
R10062 gnd.n3401 gnd.n1420 585
R10063 gnd.n3400 gnd.n1444 585
R10064 gnd.n3400 gnd.n3399 585
R10065 gnd.n3398 gnd.n3396 585
R10066 gnd.n3398 gnd.n3397 585
R10067 gnd.n1445 gnd.n1409 585
R10068 gnd.n3613 gnd.n1409 585
R10069 gnd.n3392 gnd.n3391 585
R10070 gnd.n3391 gnd.n3390 585
R10071 gnd.n1448 gnd.n1447 585
R10072 gnd.n1453 gnd.n1448 585
R10073 gnd.n1472 gnd.n1460 585
R10074 gnd.n3372 gnd.n1460 585
R10075 gnd.n3356 gnd.n3355 585
R10076 gnd.n3357 gnd.n3356 585
R10077 gnd.n1471 gnd.n1470 585
R10078 gnd.n1479 gnd.n1470 585
R10079 gnd.n3350 gnd.n3349 585
R10080 gnd.n3349 gnd.n3348 585
R10081 gnd.n1475 gnd.n1474 585
R10082 gnd.n1484 gnd.n1475 585
R10083 gnd.n3266 gnd.n1491 585
R10084 gnd.n3327 gnd.n1491 585
R10085 gnd.n3265 gnd.n1499 585
R10086 gnd.n3314 gnd.n1499 585
R10087 gnd.n3270 gnd.n3264 585
R10088 gnd.n3264 gnd.n3263 585
R10089 gnd.n3271 gnd.n3262 585
R10090 gnd.n3262 gnd.n1511 585
R10091 gnd.n3272 gnd.n3261 585
R10092 gnd.n3261 gnd.n1507 585
R10093 gnd.n1527 gnd.n1518 585
R10094 gnd.n3287 gnd.n1518 585
R10095 gnd.n3277 gnd.n3276 585
R10096 gnd.n3278 gnd.n3277 585
R10097 gnd.n1526 gnd.n1525 585
R10098 gnd.n3185 gnd.n1525 585
R10099 gnd.n3257 gnd.n3256 585
R10100 gnd.n3256 gnd.n3255 585
R10101 gnd.n1530 gnd.n1529 585
R10102 gnd.n3247 gnd.n1530 585
R10103 gnd.n1556 gnd.n1554 585
R10104 gnd.n1554 gnd.n1546 585
R10105 gnd.n3224 gnd.n3223 585
R10106 gnd.n3225 gnd.n3224 585
R10107 gnd.n1555 gnd.n1553 585
R10108 gnd.n1553 gnd.n1550 585
R10109 gnd.n3218 gnd.n3217 585
R10110 gnd.n3217 gnd.n3216 585
R10111 gnd.n1559 gnd.n1558 585
R10112 gnd.n1568 gnd.n1559 585
R10113 gnd.n3098 gnd.n3096 585
R10114 gnd.n3096 gnd.n3095 585
R10115 gnd.n3099 gnd.n3093 585
R10116 gnd.n3093 gnd.n1573 585
R10117 gnd.n3100 gnd.n1581 585
R10118 gnd.n3157 gnd.n1581 585
R10119 gnd.n3091 gnd.n1588 585
R10120 gnd.n3145 gnd.n1588 585
R10121 gnd.n3104 gnd.n3090 585
R10122 gnd.n3090 gnd.n1593 585
R10123 gnd.n3105 gnd.n3089 585
R10124 gnd.n3089 gnd.n1600 585
R10125 gnd.n3106 gnd.n3088 585
R10126 gnd.n3088 gnd.n3087 585
R10127 gnd.n1617 gnd.n1607 585
R10128 gnd.n3120 gnd.n1607 585
R10129 gnd.n3111 gnd.n3110 585
R10130 gnd.n3112 gnd.n3111 585
R10131 gnd.n1616 gnd.n1615 585
R10132 gnd.n3074 gnd.n1615 585
R10133 gnd.n3048 gnd.n3047 585
R10134 gnd.n3047 gnd.n3046 585
R10135 gnd.n1640 gnd.n1638 585
R10136 gnd.n1638 gnd.n1630 585
R10137 gnd.n3053 gnd.n3052 585
R10138 gnd.n3054 gnd.n3053 585
R10139 gnd.n1639 gnd.n1637 585
R10140 gnd.n3034 gnd.n1637 585
R10141 gnd.n3005 gnd.n3004 585
R10142 gnd.n3007 gnd.n3005 585
R10143 gnd.n1664 gnd.n1663 585
R10144 gnd.n1663 gnd.n1653 585
R10145 gnd.n3000 gnd.n2999 585
R10146 gnd.n2999 gnd.n2998 585
R10147 gnd.n2997 gnd.n1666 585
R10148 gnd.n2997 gnd.n1658 585
R10149 gnd.n2996 gnd.n1668 585
R10150 gnd.n2996 gnd.n2995 585
R10151 gnd.n2911 gnd.n1667 585
R10152 gnd.n2986 gnd.n1667 585
R10153 gnd.n2912 gnd.n1685 585
R10154 gnd.n2973 gnd.n1685 585
R10155 gnd.n2908 gnd.n2907 585
R10156 gnd.n2907 gnd.n1690 585
R10157 gnd.n2916 gnd.n2906 585
R10158 gnd.n2906 gnd.n2905 585
R10159 gnd.n2917 gnd.n2902 585
R10160 gnd.n2902 gnd.n1695 585
R10161 gnd.n2918 gnd.n1702 585
R10162 gnd.n2946 gnd.n1702 585
R10163 gnd.n1716 gnd.n1710 585
R10164 gnd.n2938 gnd.n1710 585
R10165 gnd.n2923 gnd.n2922 585
R10166 gnd.n2925 gnd.n2923 585
R10167 gnd.n1715 gnd.n1714 585
R10168 gnd.n2875 gnd.n1714 585
R10169 gnd.n2898 gnd.n2897 585
R10170 gnd.n2897 gnd.n2896 585
R10171 gnd.n1719 gnd.n1718 585
R10172 gnd.n1731 gnd.n1719 585
R10173 gnd.n2819 gnd.n2818 585
R10174 gnd.n2818 gnd.n1729 585
R10175 gnd.n2820 gnd.n2817 585
R10176 gnd.n2817 gnd.n1736 585
R10177 gnd.n1764 gnd.n1762 585
R10178 gnd.n1762 gnd.n1740 585
R10179 gnd.n2825 gnd.n2824 585
R10180 gnd.n2826 gnd.n2825 585
R10181 gnd.n1763 gnd.n1761 585
R10182 gnd.n1761 gnd.n1760 585
R10183 gnd.n2813 gnd.n2812 585
R10184 gnd.n2812 gnd.n1751 585
R10185 gnd.n2811 gnd.n1766 585
R10186 gnd.n2811 gnd.n2810 585
R10187 gnd.n1785 gnd.n1767 585
R10188 gnd.n2799 gnd.n1767 585
R10189 gnd.n2788 gnd.n2787 585
R10190 gnd.n2790 gnd.n2788 585
R10191 gnd.n1784 gnd.n1783 585
R10192 gnd.n1862 gnd.n1783 585
R10193 gnd.n2782 gnd.n2781 585
R10194 gnd.n2781 gnd.n2780 585
R10195 gnd.n1788 gnd.n1787 585
R10196 gnd.n2616 gnd.n1788 585
R10197 gnd.n2627 gnd.n2626 585
R10198 gnd.n2626 gnd.n1816 585
R10199 gnd.n2630 gnd.n2625 585
R10200 gnd.n2625 gnd.n2624 585
R10201 gnd.n2631 gnd.n2060 585
R10202 gnd.n2604 gnd.n2060 585
R10203 gnd.n2632 gnd.n2059 585
R10204 gnd.n2603 gnd.n2059 585
R10205 gnd.n2599 gnd.n2057 585
R10206 gnd.n2601 gnd.n2599 585
R10207 gnd.n2636 gnd.n2056 585
R10208 gnd.n2068 gnd.n2056 585
R10209 gnd.n2637 gnd.n2055 585
R10210 gnd.n2589 gnd.n2055 585
R10211 gnd.n2638 gnd.n2054 585
R10212 gnd.n2587 gnd.n2054 585
R10213 gnd.n3586 gnd.n3585 585
R10214 gnd.n3585 gnd.n1203 585
R10215 gnd.n3584 gnd.n3414 585
R10216 gnd.n3582 gnd.n3581 585
R10217 gnd.n3416 gnd.n3415 585
R10218 gnd.n3577 gnd.n3573 585
R10219 gnd.n3571 gnd.n3418 585
R10220 gnd.n3569 gnd.n3568 585
R10221 gnd.n3420 gnd.n3419 585
R10222 gnd.n3564 gnd.n3563 585
R10223 gnd.n3561 gnd.n3422 585
R10224 gnd.n3559 gnd.n3558 585
R10225 gnd.n3424 gnd.n3423 585
R10226 gnd.n3544 gnd.n3543 585
R10227 gnd.n3545 gnd.n3541 585
R10228 gnd.n3539 gnd.n3433 585
R10229 gnd.n3538 gnd.n3537 585
R10230 gnd.n3522 gnd.n3435 585
R10231 gnd.n3524 gnd.n3523 585
R10232 gnd.n3520 gnd.n3442 585
R10233 gnd.n3519 gnd.n3518 585
R10234 gnd.n3503 gnd.n3444 585
R10235 gnd.n3505 gnd.n3504 585
R10236 gnd.n3501 gnd.n3451 585
R10237 gnd.n3500 gnd.n3499 585
R10238 gnd.n3484 gnd.n3453 585
R10239 gnd.n3486 gnd.n3485 585
R10240 gnd.n3482 gnd.n3460 585
R10241 gnd.n3481 gnd.n3480 585
R10242 gnd.n3462 gnd.n1191 585
R10243 gnd.n3703 gnd.n1404 482.89
R10244 gnd.n3706 gnd.n3705 482.89
R10245 gnd.n1869 gnd.n1868 482.89
R10246 gnd.n2773 gnd.n1792 482.89
R10247 gnd.n1854 gnd.t183 443.966
R10248 gnd.n1398 gnd.t197 443.966
R10249 gnd.n1851 gnd.t216 443.966
R10250 gnd.n3637 gnd.t126 443.966
R10251 gnd.n6065 gnd.n6064 422.406
R10252 gnd.n2045 gnd.t176 371.625
R10253 gnd.n6752 gnd.t164 371.625
R10254 gnd.n3426 gnd.t154 371.625
R10255 gnd.n2148 gnd.t173 371.625
R10256 gnd.n3830 gnd.t151 371.625
R10257 gnd.n1337 gnd.t122 371.625
R10258 gnd.n156 gnd.t118 371.625
R10259 gnd.n6844 gnd.t137 371.625
R10260 gnd.n852 gnd.t209 371.625
R10261 gnd.n874 gnd.t203 371.625
R10262 gnd.n2292 gnd.t190 371.625
R10263 gnd.n2024 gnd.t133 371.625
R10264 gnd.n1935 gnd.t167 371.625
R10265 gnd.n3574 gnd.t157 371.625
R10266 gnd.n4862 gnd.t111 323.425
R10267 gnd.n4513 gnd.t140 323.425
R10268 gnd.n5717 gnd.n5691 289.615
R10269 gnd.n5685 gnd.n5659 289.615
R10270 gnd.n5653 gnd.n5627 289.615
R10271 gnd.n5622 gnd.n5596 289.615
R10272 gnd.n5590 gnd.n5564 289.615
R10273 gnd.n5558 gnd.n5532 289.615
R10274 gnd.n5526 gnd.n5500 289.615
R10275 gnd.n5495 gnd.n5469 289.615
R10276 gnd.n4936 gnd.t212 279.217
R10277 gnd.n4557 gnd.t147 279.217
R10278 gnd.n1799 gnd.t202 260.649
R10279 gnd.n3629 gnd.t132 260.649
R10280 gnd.n2772 gnd.n2771 256.663
R10281 gnd.n2771 gnd.n1817 256.663
R10282 gnd.n2771 gnd.n1818 256.663
R10283 gnd.n2771 gnd.n1819 256.663
R10284 gnd.n2771 gnd.n1820 256.663
R10285 gnd.n2771 gnd.n1821 256.663
R10286 gnd.n2771 gnd.n1822 256.663
R10287 gnd.n2771 gnd.n1823 256.663
R10288 gnd.n2771 gnd.n1824 256.663
R10289 gnd.n2771 gnd.n1825 256.663
R10290 gnd.n2771 gnd.n1826 256.663
R10291 gnd.n2771 gnd.n1827 256.663
R10292 gnd.n2771 gnd.n1828 256.663
R10293 gnd.n2771 gnd.n1829 256.663
R10294 gnd.n2771 gnd.n1830 256.663
R10295 gnd.n2771 gnd.n1831 256.663
R10296 gnd.n2711 gnd.n2708 256.663
R10297 gnd.n2771 gnd.n1832 256.663
R10298 gnd.n2771 gnd.n1833 256.663
R10299 gnd.n2771 gnd.n1834 256.663
R10300 gnd.n2771 gnd.n1835 256.663
R10301 gnd.n2771 gnd.n1836 256.663
R10302 gnd.n2771 gnd.n1837 256.663
R10303 gnd.n2771 gnd.n1838 256.663
R10304 gnd.n2771 gnd.n1839 256.663
R10305 gnd.n2771 gnd.n1840 256.663
R10306 gnd.n2771 gnd.n1841 256.663
R10307 gnd.n2771 gnd.n1842 256.663
R10308 gnd.n2771 gnd.n1843 256.663
R10309 gnd.n2771 gnd.n1844 256.663
R10310 gnd.n2771 gnd.n1845 256.663
R10311 gnd.n2771 gnd.n1846 256.663
R10312 gnd.n2771 gnd.n1847 256.663
R10313 gnd.n2771 gnd.n1848 256.663
R10314 gnd.n3771 gnd.n1382 256.663
R10315 gnd.n3771 gnd.n1383 256.663
R10316 gnd.n3771 gnd.n1384 256.663
R10317 gnd.n3771 gnd.n1385 256.663
R10318 gnd.n3771 gnd.n1386 256.663
R10319 gnd.n3771 gnd.n1387 256.663
R10320 gnd.n3771 gnd.n1388 256.663
R10321 gnd.n3771 gnd.n1389 256.663
R10322 gnd.n3771 gnd.n1390 256.663
R10323 gnd.n3771 gnd.n1391 256.663
R10324 gnd.n3771 gnd.n1392 256.663
R10325 gnd.n3771 gnd.n1393 256.663
R10326 gnd.n3771 gnd.n1394 256.663
R10327 gnd.n3771 gnd.n1395 256.663
R10328 gnd.n3771 gnd.n1396 256.663
R10329 gnd.n3771 gnd.n3768 256.663
R10330 gnd.n3774 gnd.n1363 256.663
R10331 gnd.n3772 gnd.n3771 256.663
R10332 gnd.n3771 gnd.n1381 256.663
R10333 gnd.n3771 gnd.n1380 256.663
R10334 gnd.n3771 gnd.n1379 256.663
R10335 gnd.n3771 gnd.n1378 256.663
R10336 gnd.n3771 gnd.n1377 256.663
R10337 gnd.n3771 gnd.n1376 256.663
R10338 gnd.n3771 gnd.n1375 256.663
R10339 gnd.n3771 gnd.n1374 256.663
R10340 gnd.n3771 gnd.n1373 256.663
R10341 gnd.n3771 gnd.n1372 256.663
R10342 gnd.n3771 gnd.n1371 256.663
R10343 gnd.n3771 gnd.n1370 256.663
R10344 gnd.n3771 gnd.n1369 256.663
R10345 gnd.n3771 gnd.n1368 256.663
R10346 gnd.n3771 gnd.n1367 256.663
R10347 gnd.n3771 gnd.n1366 256.663
R10348 gnd.n4482 gnd.n820 242.672
R10349 gnd.n4482 gnd.n821 242.672
R10350 gnd.n4482 gnd.n822 242.672
R10351 gnd.n4482 gnd.n823 242.672
R10352 gnd.n4482 gnd.n824 242.672
R10353 gnd.n4482 gnd.n825 242.672
R10354 gnd.n4482 gnd.n826 242.672
R10355 gnd.n4482 gnd.n827 242.672
R10356 gnd.n4482 gnd.n828 242.672
R10357 gnd.n2157 gnd.n1996 242.672
R10358 gnd.n2146 gnd.n1996 242.672
R10359 gnd.n2143 gnd.n1996 242.672
R10360 gnd.n2134 gnd.n1996 242.672
R10361 gnd.n2123 gnd.n1996 242.672
R10362 gnd.n2120 gnd.n1996 242.672
R10363 gnd.n2111 gnd.n1996 242.672
R10364 gnd.n2101 gnd.n1996 242.672
R10365 gnd.n2098 gnd.n1996 242.672
R10366 gnd.n3472 gnd.n1204 242.672
R10367 gnd.n3474 gnd.n1204 242.672
R10368 gnd.n3491 gnd.n1204 242.672
R10369 gnd.n3493 gnd.n1204 242.672
R10370 gnd.n3510 gnd.n1204 242.672
R10371 gnd.n3512 gnd.n1204 242.672
R10372 gnd.n3529 gnd.n1204 242.672
R10373 gnd.n3531 gnd.n1204 242.672
R10374 gnd.n3550 gnd.n1204 242.672
R10375 gnd.n6754 gnd.n83 242.672
R10376 gnd.n6750 gnd.n83 242.672
R10377 gnd.n6745 gnd.n83 242.672
R10378 gnd.n6742 gnd.n83 242.672
R10379 gnd.n6737 gnd.n83 242.672
R10380 gnd.n6734 gnd.n83 242.672
R10381 gnd.n6729 gnd.n83 242.672
R10382 gnd.n6726 gnd.n83 242.672
R10383 gnd.n6721 gnd.n83 242.672
R10384 gnd.n4990 gnd.n4989 242.672
R10385 gnd.n4990 gnd.n4900 242.672
R10386 gnd.n4990 gnd.n4901 242.672
R10387 gnd.n4990 gnd.n4902 242.672
R10388 gnd.n4990 gnd.n4903 242.672
R10389 gnd.n4990 gnd.n4904 242.672
R10390 gnd.n4990 gnd.n4905 242.672
R10391 gnd.n4990 gnd.n4906 242.672
R10392 gnd.n4990 gnd.n4907 242.672
R10393 gnd.n4990 gnd.n4908 242.672
R10394 gnd.n4990 gnd.n4909 242.672
R10395 gnd.n4990 gnd.n4910 242.672
R10396 gnd.n4991 gnd.n4990 242.672
R10397 gnd.n5791 gnd.n4483 242.672
R10398 gnd.n5797 gnd.n4483 242.672
R10399 gnd.n4560 gnd.n4483 242.672
R10400 gnd.n5804 gnd.n4483 242.672
R10401 gnd.n4551 gnd.n4483 242.672
R10402 gnd.n5811 gnd.n4483 242.672
R10403 gnd.n4544 gnd.n4483 242.672
R10404 gnd.n5818 gnd.n4483 242.672
R10405 gnd.n4537 gnd.n4483 242.672
R10406 gnd.n5825 gnd.n4483 242.672
R10407 gnd.n4530 gnd.n4483 242.672
R10408 gnd.n5832 gnd.n4483 242.672
R10409 gnd.n4523 gnd.n4483 242.672
R10410 gnd.n5148 gnd.n5147 242.672
R10411 gnd.n5147 gnd.n4812 242.672
R10412 gnd.n5147 gnd.n4813 242.672
R10413 gnd.n5147 gnd.n4814 242.672
R10414 gnd.n5147 gnd.n4815 242.672
R10415 gnd.n5147 gnd.n4816 242.672
R10416 gnd.n5147 gnd.n4817 242.672
R10417 gnd.n5147 gnd.n4818 242.672
R10418 gnd.n5843 gnd.n4483 242.672
R10419 gnd.n4516 gnd.n4483 242.672
R10420 gnd.n5850 gnd.n4483 242.672
R10421 gnd.n4507 gnd.n4483 242.672
R10422 gnd.n5857 gnd.n4483 242.672
R10423 gnd.n4500 gnd.n4483 242.672
R10424 gnd.n5864 gnd.n4483 242.672
R10425 gnd.n4493 gnd.n4483 242.672
R10426 gnd.n4482 gnd.n4481 242.672
R10427 gnd.n4482 gnd.n802 242.672
R10428 gnd.n4482 gnd.n803 242.672
R10429 gnd.n4482 gnd.n804 242.672
R10430 gnd.n4482 gnd.n805 242.672
R10431 gnd.n4482 gnd.n806 242.672
R10432 gnd.n4482 gnd.n807 242.672
R10433 gnd.n4482 gnd.n808 242.672
R10434 gnd.n4482 gnd.n809 242.672
R10435 gnd.n4482 gnd.n810 242.672
R10436 gnd.n4482 gnd.n811 242.672
R10437 gnd.n4482 gnd.n812 242.672
R10438 gnd.n4482 gnd.n813 242.672
R10439 gnd.n4482 gnd.n814 242.672
R10440 gnd.n4482 gnd.n815 242.672
R10441 gnd.n4482 gnd.n816 242.672
R10442 gnd.n4482 gnd.n817 242.672
R10443 gnd.n4482 gnd.n818 242.672
R10444 gnd.n4482 gnd.n819 242.672
R10445 gnd.n2670 gnd.n1996 242.672
R10446 gnd.n2027 gnd.n1996 242.672
R10447 gnd.n2677 gnd.n1996 242.672
R10448 gnd.n2018 gnd.n1996 242.672
R10449 gnd.n2684 gnd.n1996 242.672
R10450 gnd.n2011 gnd.n1996 242.672
R10451 gnd.n2691 gnd.n1996 242.672
R10452 gnd.n2004 gnd.n1996 242.672
R10453 gnd.n2698 gnd.n1996 242.672
R10454 gnd.n2701 gnd.n1996 242.672
R10455 gnd.n1996 gnd.n1942 242.672
R10456 gnd.n2707 gnd.n1937 242.672
R10457 gnd.n1996 gnd.n1943 242.672
R10458 gnd.n1996 gnd.n1944 242.672
R10459 gnd.n1996 gnd.n1945 242.672
R10460 gnd.n1996 gnd.n1946 242.672
R10461 gnd.n1996 gnd.n1947 242.672
R10462 gnd.n1996 gnd.n1948 242.672
R10463 gnd.n1996 gnd.n1949 242.672
R10464 gnd.n1996 gnd.n1995 242.672
R10465 gnd.n3793 gnd.n1204 242.672
R10466 gnd.n3796 gnd.n1204 242.672
R10467 gnd.n3804 gnd.n1204 242.672
R10468 gnd.n3806 gnd.n1204 242.672
R10469 gnd.n3814 gnd.n1204 242.672
R10470 gnd.n3816 gnd.n1204 242.672
R10471 gnd.n3825 gnd.n1204 242.672
R10472 gnd.n3828 gnd.n1204 242.672
R10473 gnd.n3832 gnd.n3829 242.672
R10474 gnd.n3775 gnd.n1204 242.672
R10475 gnd.n3838 gnd.n1204 242.672
R10476 gnd.n3840 gnd.n1204 242.672
R10477 gnd.n3848 gnd.n1204 242.672
R10478 gnd.n3850 gnd.n1204 242.672
R10479 gnd.n3858 gnd.n1204 242.672
R10480 gnd.n3860 gnd.n1204 242.672
R10481 gnd.n3868 gnd.n1204 242.672
R10482 gnd.n3870 gnd.n1204 242.672
R10483 gnd.n3879 gnd.n1204 242.672
R10484 gnd.n3882 gnd.n1204 242.672
R10485 gnd.n153 gnd.n83 242.672
R10486 gnd.n6812 gnd.n83 242.672
R10487 gnd.n149 gnd.n83 242.672
R10488 gnd.n6819 gnd.n83 242.672
R10489 gnd.n142 gnd.n83 242.672
R10490 gnd.n6826 gnd.n83 242.672
R10491 gnd.n135 gnd.n83 242.672
R10492 gnd.n6833 gnd.n83 242.672
R10493 gnd.n128 gnd.n83 242.672
R10494 gnd.n6840 gnd.n83 242.672
R10495 gnd.n121 gnd.n83 242.672
R10496 gnd.n6850 gnd.n83 242.672
R10497 gnd.n114 gnd.n83 242.672
R10498 gnd.n6857 gnd.n83 242.672
R10499 gnd.n107 gnd.n83 242.672
R10500 gnd.n6864 gnd.n83 242.672
R10501 gnd.n100 gnd.n83 242.672
R10502 gnd.n6871 gnd.n83 242.672
R10503 gnd.n93 gnd.n83 242.672
R10504 gnd.n2206 gnd.n2205 242.672
R10505 gnd.n2206 gnd.n2074 242.672
R10506 gnd.n2206 gnd.n2075 242.672
R10507 gnd.n2206 gnd.n2076 242.672
R10508 gnd.n2206 gnd.n2077 242.672
R10509 gnd.n2206 gnd.n2078 242.672
R10510 gnd.n2206 gnd.n2079 242.672
R10511 gnd.n2206 gnd.n2080 242.672
R10512 gnd.n2206 gnd.n2081 242.672
R10513 gnd.n2206 gnd.n2082 242.672
R10514 gnd.n2206 gnd.n2084 242.672
R10515 gnd.n2206 gnd.n2085 242.672
R10516 gnd.n2206 gnd.n2086 242.672
R10517 gnd.n2206 gnd.n2088 242.672
R10518 gnd.n3583 gnd.n1203 242.672
R10519 gnd.n3572 gnd.n1203 242.672
R10520 gnd.n3570 gnd.n1203 242.672
R10521 gnd.n3562 gnd.n1203 242.672
R10522 gnd.n3560 gnd.n1203 242.672
R10523 gnd.n3542 gnd.n1203 242.672
R10524 gnd.n3540 gnd.n1203 242.672
R10525 gnd.n3434 gnd.n1203 242.672
R10526 gnd.n3521 gnd.n1203 242.672
R10527 gnd.n3443 gnd.n1203 242.672
R10528 gnd.n3502 gnd.n1203 242.672
R10529 gnd.n3452 gnd.n1203 242.672
R10530 gnd.n3483 gnd.n1203 242.672
R10531 gnd.n3461 gnd.n1203 242.672
R10532 gnd.n90 gnd.n86 240.244
R10533 gnd.n6873 gnd.n6872 240.244
R10534 gnd.n6870 gnd.n94 240.244
R10535 gnd.n6866 gnd.n6865 240.244
R10536 gnd.n6863 gnd.n101 240.244
R10537 gnd.n6859 gnd.n6858 240.244
R10538 gnd.n6856 gnd.n108 240.244
R10539 gnd.n6852 gnd.n6851 240.244
R10540 gnd.n6849 gnd.n115 240.244
R10541 gnd.n6842 gnd.n6841 240.244
R10542 gnd.n6839 gnd.n122 240.244
R10543 gnd.n6835 gnd.n6834 240.244
R10544 gnd.n6832 gnd.n129 240.244
R10545 gnd.n6828 gnd.n6827 240.244
R10546 gnd.n6825 gnd.n136 240.244
R10547 gnd.n6821 gnd.n6820 240.244
R10548 gnd.n6818 gnd.n143 240.244
R10549 gnd.n6814 gnd.n6813 240.244
R10550 gnd.n6811 gnd.n150 240.244
R10551 gnd.n3889 gnd.n1213 240.244
R10552 gnd.n3889 gnd.n1225 240.244
R10553 gnd.n3900 gnd.n1225 240.244
R10554 gnd.n3900 gnd.n1326 240.244
R10555 gnd.n3991 gnd.n1326 240.244
R10556 gnd.n3991 gnd.n1319 240.244
R10557 gnd.n3987 gnd.n1319 240.244
R10558 gnd.n3987 gnd.n1311 240.244
R10559 gnd.n1311 gnd.n1300 240.244
R10560 gnd.n3983 gnd.n1300 240.244
R10561 gnd.n3983 gnd.n1290 240.244
R10562 gnd.n3980 gnd.n1290 240.244
R10563 gnd.n3980 gnd.n1282 240.244
R10564 gnd.n1282 gnd.n1271 240.244
R10565 gnd.n3976 gnd.n1271 240.244
R10566 gnd.n3976 gnd.n1261 240.244
R10567 gnd.n3973 gnd.n1261 240.244
R10568 gnd.n3973 gnd.n1252 240.244
R10569 gnd.n1252 gnd.n249 240.244
R10570 gnd.n249 gnd.n244 240.244
R10571 gnd.n3967 gnd.n244 240.244
R10572 gnd.n3967 gnd.n237 240.244
R10573 gnd.n3962 gnd.n237 240.244
R10574 gnd.n3962 gnd.n231 240.244
R10575 gnd.n3959 gnd.n231 240.244
R10576 gnd.n3959 gnd.n223 240.244
R10577 gnd.n3956 gnd.n223 240.244
R10578 gnd.n3956 gnd.n209 240.244
R10579 gnd.n3953 gnd.n209 240.244
R10580 gnd.n3953 gnd.n203 240.244
R10581 gnd.n3950 gnd.n203 240.244
R10582 gnd.n3950 gnd.n195 240.244
R10583 gnd.n3947 gnd.n195 240.244
R10584 gnd.n3947 gnd.n187 240.244
R10585 gnd.n3944 gnd.n187 240.244
R10586 gnd.n3944 gnd.n179 240.244
R10587 gnd.n3941 gnd.n179 240.244
R10588 gnd.n3941 gnd.n171 240.244
R10589 gnd.n171 gnd.n160 240.244
R10590 gnd.n6802 gnd.n160 240.244
R10591 gnd.n6803 gnd.n6802 240.244
R10592 gnd.n6803 gnd.n82 240.244
R10593 gnd.n3795 gnd.n3794 240.244
R10594 gnd.n3797 gnd.n3795 240.244
R10595 gnd.n3803 gnd.n3785 240.244
R10596 gnd.n3807 gnd.n3805 240.244
R10597 gnd.n3813 gnd.n3781 240.244
R10598 gnd.n3817 gnd.n3815 240.244
R10599 gnd.n3824 gnd.n3777 240.244
R10600 gnd.n3827 gnd.n3826 240.244
R10601 gnd.n3837 gnd.n1357 240.244
R10602 gnd.n3841 gnd.n3839 240.244
R10603 gnd.n3847 gnd.n1353 240.244
R10604 gnd.n3851 gnd.n3849 240.244
R10605 gnd.n3857 gnd.n1349 240.244
R10606 gnd.n3861 gnd.n3859 240.244
R10607 gnd.n3867 gnd.n1345 240.244
R10608 gnd.n3871 gnd.n3869 240.244
R10609 gnd.n3878 gnd.n1341 240.244
R10610 gnd.n3881 gnd.n3880 240.244
R10611 gnd.n4129 gnd.n1218 240.244
R10612 gnd.n4125 gnd.n1218 240.244
R10613 gnd.n4125 gnd.n1223 240.244
R10614 gnd.n4011 gnd.n1223 240.244
R10615 gnd.n4011 gnd.n1321 240.244
R10616 gnd.n4019 gnd.n1321 240.244
R10617 gnd.n4019 gnd.n1322 240.244
R10618 gnd.n1322 gnd.n1298 240.244
R10619 gnd.n4042 gnd.n1298 240.244
R10620 gnd.n4042 gnd.n1293 240.244
R10621 gnd.n4051 gnd.n1293 240.244
R10622 gnd.n4051 gnd.n1294 240.244
R10623 gnd.n1294 gnd.n1269 240.244
R10624 gnd.n4081 gnd.n1269 240.244
R10625 gnd.n4081 gnd.n1263 240.244
R10626 gnd.n4085 gnd.n1263 240.244
R10627 gnd.n4085 gnd.n1266 240.244
R10628 gnd.n1266 gnd.n247 240.244
R10629 gnd.n6645 gnd.n247 240.244
R10630 gnd.n6648 gnd.n6645 240.244
R10631 gnd.n6648 gnd.n233 240.244
R10632 gnd.n6658 gnd.n233 240.244
R10633 gnd.n6659 gnd.n6658 240.244
R10634 gnd.n6662 gnd.n6659 240.244
R10635 gnd.n6662 gnd.n220 240.244
R10636 gnd.n6672 gnd.n220 240.244
R10637 gnd.n6672 gnd.n210 240.244
R10638 gnd.n6678 gnd.n210 240.244
R10639 gnd.n6678 gnd.n200 240.244
R10640 gnd.n6688 gnd.n200 240.244
R10641 gnd.n6688 gnd.n196 240.244
R10642 gnd.n6694 gnd.n196 240.244
R10643 gnd.n6694 gnd.n184 240.244
R10644 gnd.n6704 gnd.n184 240.244
R10645 gnd.n6704 gnd.n180 240.244
R10646 gnd.n6710 gnd.n180 240.244
R10647 gnd.n6710 gnd.n168 240.244
R10648 gnd.n6794 gnd.n168 240.244
R10649 gnd.n6794 gnd.n164 240.244
R10650 gnd.n6800 gnd.n164 240.244
R10651 gnd.n6800 gnd.n85 240.244
R10652 gnd.n6880 gnd.n85 240.244
R10653 gnd.n1950 gnd.n1078 240.244
R10654 gnd.n1994 gnd.n1951 240.244
R10655 gnd.n1990 gnd.n1989 240.244
R10656 gnd.n1986 gnd.n1985 240.244
R10657 gnd.n1982 gnd.n1981 240.244
R10658 gnd.n1978 gnd.n1977 240.244
R10659 gnd.n1974 gnd.n1973 240.244
R10660 gnd.n1970 gnd.n1969 240.244
R10661 gnd.n2702 gnd.n1941 240.244
R10662 gnd.n2700 gnd.n2699 240.244
R10663 gnd.n2697 gnd.n1998 240.244
R10664 gnd.n2693 gnd.n2692 240.244
R10665 gnd.n2690 gnd.n2005 240.244
R10666 gnd.n2686 gnd.n2685 240.244
R10667 gnd.n2683 gnd.n2012 240.244
R10668 gnd.n2679 gnd.n2678 240.244
R10669 gnd.n2676 gnd.n2019 240.244
R10670 gnd.n2672 gnd.n2671 240.244
R10671 gnd.n4403 gnd.n878 240.244
R10672 gnd.n882 gnd.n878 240.244
R10673 gnd.n4396 gnd.n882 240.244
R10674 gnd.n4396 gnd.n883 240.244
R10675 gnd.n896 gnd.n883 240.244
R10676 gnd.n2392 gnd.n896 240.244
R10677 gnd.n2392 gnd.n907 240.244
R10678 gnd.n2387 gnd.n907 240.244
R10679 gnd.n2387 gnd.n917 240.244
R10680 gnd.n2399 gnd.n917 240.244
R10681 gnd.n2399 gnd.n927 240.244
R10682 gnd.n2384 gnd.n927 240.244
R10683 gnd.n2384 gnd.n937 240.244
R10684 gnd.n2406 gnd.n937 240.244
R10685 gnd.n2406 gnd.n947 240.244
R10686 gnd.n2381 gnd.n947 240.244
R10687 gnd.n2419 gnd.n2381 240.244
R10688 gnd.n2419 gnd.n958 240.244
R10689 gnd.n2415 gnd.n958 240.244
R10690 gnd.n2415 gnd.n971 240.244
R10691 gnd.n2432 gnd.n971 240.244
R10692 gnd.n2432 gnd.n979 240.244
R10693 gnd.n2248 gnd.n979 240.244
R10694 gnd.n2248 gnd.n988 240.244
R10695 gnd.n2444 gnd.n988 240.244
R10696 gnd.n2444 gnd.n996 240.244
R10697 gnd.n2242 gnd.n996 240.244
R10698 gnd.n2242 gnd.n1006 240.244
R10699 gnd.n2511 gnd.n1006 240.244
R10700 gnd.n2511 gnd.n1017 240.244
R10701 gnd.n2517 gnd.n1017 240.244
R10702 gnd.n2517 gnd.n1027 240.244
R10703 gnd.n2527 gnd.n1027 240.244
R10704 gnd.n2527 gnd.n1038 240.244
R10705 gnd.n2221 gnd.n1038 240.244
R10706 gnd.n2221 gnd.n1048 240.244
R10707 gnd.n2535 gnd.n1048 240.244
R10708 gnd.n2535 gnd.n1059 240.244
R10709 gnd.n2542 gnd.n1059 240.244
R10710 gnd.n2542 gnd.n1070 240.244
R10711 gnd.n2663 gnd.n1070 240.244
R10712 gnd.n2663 gnd.n1080 240.244
R10713 gnd.n832 gnd.n831 240.244
R10714 gnd.n4475 gnd.n831 240.244
R10715 gnd.n4473 gnd.n4472 240.244
R10716 gnd.n4469 gnd.n4468 240.244
R10717 gnd.n4465 gnd.n4464 240.244
R10718 gnd.n4461 gnd.n4460 240.244
R10719 gnd.n4457 gnd.n4456 240.244
R10720 gnd.n4453 gnd.n4452 240.244
R10721 gnd.n4449 gnd.n4448 240.244
R10722 gnd.n4444 gnd.n4443 240.244
R10723 gnd.n4440 gnd.n4439 240.244
R10724 gnd.n4436 gnd.n4435 240.244
R10725 gnd.n4432 gnd.n4431 240.244
R10726 gnd.n4428 gnd.n4427 240.244
R10727 gnd.n4424 gnd.n4423 240.244
R10728 gnd.n4420 gnd.n4419 240.244
R10729 gnd.n4416 gnd.n4415 240.244
R10730 gnd.n4412 gnd.n4411 240.244
R10731 gnd.n873 gnd.n872 240.244
R10732 gnd.n2350 gnd.n833 240.244
R10733 gnd.n2350 gnd.n888 240.244
R10734 gnd.n4394 gnd.n888 240.244
R10735 gnd.n4394 gnd.n889 240.244
R10736 gnd.n4390 gnd.n889 240.244
R10737 gnd.n4390 gnd.n895 240.244
R10738 gnd.n4382 gnd.n895 240.244
R10739 gnd.n4382 gnd.n910 240.244
R10740 gnd.n4378 gnd.n910 240.244
R10741 gnd.n4378 gnd.n916 240.244
R10742 gnd.n4370 gnd.n916 240.244
R10743 gnd.n4370 gnd.n929 240.244
R10744 gnd.n4366 gnd.n929 240.244
R10745 gnd.n4366 gnd.n935 240.244
R10746 gnd.n4358 gnd.n935 240.244
R10747 gnd.n4358 gnd.n950 240.244
R10748 gnd.n954 gnd.n950 240.244
R10749 gnd.n4352 gnd.n954 240.244
R10750 gnd.n4352 gnd.n956 240.244
R10751 gnd.n4344 gnd.n956 240.244
R10752 gnd.n4344 gnd.n974 240.244
R10753 gnd.n4339 gnd.n974 240.244
R10754 gnd.n4339 gnd.n977 240.244
R10755 gnd.n4331 gnd.n977 240.244
R10756 gnd.n4331 gnd.n991 240.244
R10757 gnd.n4326 gnd.n991 240.244
R10758 gnd.n4326 gnd.n994 240.244
R10759 gnd.n4318 gnd.n994 240.244
R10760 gnd.n4318 gnd.n1009 240.244
R10761 gnd.n4314 gnd.n1009 240.244
R10762 gnd.n4314 gnd.n1015 240.244
R10763 gnd.n4306 gnd.n1015 240.244
R10764 gnd.n4306 gnd.n1030 240.244
R10765 gnd.n4302 gnd.n1030 240.244
R10766 gnd.n4302 gnd.n1036 240.244
R10767 gnd.n4294 gnd.n1036 240.244
R10768 gnd.n4294 gnd.n1051 240.244
R10769 gnd.n4290 gnd.n1051 240.244
R10770 gnd.n4290 gnd.n1057 240.244
R10771 gnd.n4282 gnd.n1057 240.244
R10772 gnd.n4282 gnd.n1073 240.244
R10773 gnd.n4278 gnd.n1073 240.244
R10774 gnd.n4490 gnd.n4485 240.244
R10775 gnd.n5866 gnd.n5865 240.244
R10776 gnd.n5863 gnd.n4494 240.244
R10777 gnd.n5859 gnd.n5858 240.244
R10778 gnd.n5856 gnd.n4501 240.244
R10779 gnd.n5852 gnd.n5851 240.244
R10780 gnd.n5849 gnd.n4508 240.244
R10781 gnd.n5845 gnd.n5844 240.244
R10782 gnd.n5159 gnd.n4797 240.244
R10783 gnd.n5169 gnd.n4797 240.244
R10784 gnd.n5169 gnd.n4788 240.244
R10785 gnd.n4788 gnd.n4777 240.244
R10786 gnd.n5190 gnd.n4777 240.244
R10787 gnd.n5190 gnd.n4771 240.244
R10788 gnd.n5200 gnd.n4771 240.244
R10789 gnd.n5200 gnd.n4762 240.244
R10790 gnd.n4762 gnd.n4753 240.244
R10791 gnd.n5221 gnd.n4753 240.244
R10792 gnd.n5221 gnd.n4746 240.244
R10793 gnd.n5231 gnd.n4746 240.244
R10794 gnd.n5231 gnd.n4737 240.244
R10795 gnd.n4737 gnd.n4727 240.244
R10796 gnd.n5252 gnd.n4727 240.244
R10797 gnd.n5252 gnd.n4720 240.244
R10798 gnd.n5262 gnd.n4720 240.244
R10799 gnd.n5262 gnd.n4711 240.244
R10800 gnd.n4711 gnd.n4702 240.244
R10801 gnd.n5283 gnd.n4702 240.244
R10802 gnd.n5283 gnd.n4695 240.244
R10803 gnd.n5293 gnd.n4695 240.244
R10804 gnd.n5293 gnd.n4687 240.244
R10805 gnd.n4687 gnd.n4678 240.244
R10806 gnd.n5313 gnd.n4678 240.244
R10807 gnd.n5313 gnd.n4665 240.244
R10808 gnd.n5347 gnd.n4665 240.244
R10809 gnd.n5347 gnd.n4655 240.244
R10810 gnd.n4655 gnd.n4647 240.244
R10811 gnd.n5365 gnd.n4647 240.244
R10812 gnd.n5366 gnd.n5365 240.244
R10813 gnd.n5366 gnd.n4635 240.244
R10814 gnd.n4635 gnd.n4624 240.244
R10815 gnd.n5397 gnd.n4624 240.244
R10816 gnd.n5398 gnd.n5397 240.244
R10817 gnd.n5401 gnd.n5398 240.244
R10818 gnd.n5401 gnd.n4610 240.244
R10819 gnd.n5429 gnd.n4610 240.244
R10820 gnd.n5429 gnd.n4597 240.244
R10821 gnd.n5451 gnd.n4597 240.244
R10822 gnd.n5452 gnd.n5451 240.244
R10823 gnd.n5452 gnd.n4581 240.244
R10824 gnd.n5462 gnd.n4581 240.244
R10825 gnd.n5462 gnd.n4573 240.244
R10826 gnd.n5744 gnd.n4573 240.244
R10827 gnd.n5744 gnd.n5743 240.244
R10828 gnd.n5743 gnd.n5742 240.244
R10829 gnd.n5742 gnd.n778 240.244
R10830 gnd.n5738 gnd.n778 240.244
R10831 gnd.n5738 gnd.n789 240.244
R10832 gnd.n5734 gnd.n789 240.244
R10833 gnd.n5734 gnd.n5733 240.244
R10834 gnd.n5733 gnd.n801 240.244
R10835 gnd.n5149 gnd.n4810 240.244
R10836 gnd.n4831 gnd.n4810 240.244
R10837 gnd.n4834 gnd.n4833 240.244
R10838 gnd.n4841 gnd.n4840 240.244
R10839 gnd.n4844 gnd.n4843 240.244
R10840 gnd.n4851 gnd.n4850 240.244
R10841 gnd.n4854 gnd.n4853 240.244
R10842 gnd.n4861 gnd.n4860 240.244
R10843 gnd.n5157 gnd.n4807 240.244
R10844 gnd.n4807 gnd.n4786 240.244
R10845 gnd.n5180 gnd.n4786 240.244
R10846 gnd.n5180 gnd.n4780 240.244
R10847 gnd.n5188 gnd.n4780 240.244
R10848 gnd.n5188 gnd.n4782 240.244
R10849 gnd.n4782 gnd.n4760 240.244
R10850 gnd.n5211 gnd.n4760 240.244
R10851 gnd.n5211 gnd.n4755 240.244
R10852 gnd.n5219 gnd.n4755 240.244
R10853 gnd.n5219 gnd.n4756 240.244
R10854 gnd.n4756 gnd.n4735 240.244
R10855 gnd.n5242 gnd.n4735 240.244
R10856 gnd.n5242 gnd.n4730 240.244
R10857 gnd.n5250 gnd.n4730 240.244
R10858 gnd.n5250 gnd.n4731 240.244
R10859 gnd.n4731 gnd.n4709 240.244
R10860 gnd.n5273 gnd.n4709 240.244
R10861 gnd.n5273 gnd.n4704 240.244
R10862 gnd.n5281 gnd.n4704 240.244
R10863 gnd.n5281 gnd.n4705 240.244
R10864 gnd.n4705 gnd.n4685 240.244
R10865 gnd.n5303 gnd.n4685 240.244
R10866 gnd.n5303 gnd.n4680 240.244
R10867 gnd.n5311 gnd.n4680 240.244
R10868 gnd.n5311 gnd.n4681 240.244
R10869 gnd.n4681 gnd.n4654 240.244
R10870 gnd.n5357 gnd.n4654 240.244
R10871 gnd.n5357 gnd.n4650 240.244
R10872 gnd.n5363 gnd.n4650 240.244
R10873 gnd.n5363 gnd.n4633 240.244
R10874 gnd.n5387 gnd.n4633 240.244
R10875 gnd.n5387 gnd.n4628 240.244
R10876 gnd.n5395 gnd.n4628 240.244
R10877 gnd.n5395 gnd.n4629 240.244
R10878 gnd.n4629 gnd.n4609 240.244
R10879 gnd.n5433 gnd.n4609 240.244
R10880 gnd.n5433 gnd.n4604 240.244
R10881 gnd.n5441 gnd.n4604 240.244
R10882 gnd.n5441 gnd.n4605 240.244
R10883 gnd.n4605 gnd.n4579 240.244
R10884 gnd.n5754 gnd.n4579 240.244
R10885 gnd.n5754 gnd.n4574 240.244
R10886 gnd.n5766 gnd.n4574 240.244
R10887 gnd.n5766 gnd.n4575 240.244
R10888 gnd.n5762 gnd.n4575 240.244
R10889 gnd.n5762 gnd.n780 240.244
R10890 gnd.n5887 gnd.n780 240.244
R10891 gnd.n5887 gnd.n781 240.244
R10892 gnd.n5883 gnd.n781 240.244
R10893 gnd.n5883 gnd.n787 240.244
R10894 gnd.n4484 gnd.n787 240.244
R10895 gnd.n5873 gnd.n4484 240.244
R10896 gnd.n4520 gnd.n798 240.244
R10897 gnd.n5834 gnd.n5833 240.244
R10898 gnd.n5831 gnd.n4524 240.244
R10899 gnd.n5827 gnd.n5826 240.244
R10900 gnd.n5824 gnd.n4531 240.244
R10901 gnd.n5820 gnd.n5819 240.244
R10902 gnd.n5817 gnd.n4538 240.244
R10903 gnd.n5813 gnd.n5812 240.244
R10904 gnd.n5810 gnd.n4545 240.244
R10905 gnd.n5806 gnd.n5805 240.244
R10906 gnd.n5803 gnd.n4552 240.244
R10907 gnd.n5799 gnd.n5798 240.244
R10908 gnd.n5796 gnd.n4562 240.244
R10909 gnd.n4998 gnd.n4895 240.244
R10910 gnd.n4998 gnd.n4888 240.244
R10911 gnd.n5009 gnd.n4888 240.244
R10912 gnd.n5009 gnd.n4884 240.244
R10913 gnd.n5015 gnd.n4884 240.244
R10914 gnd.n5015 gnd.n4876 240.244
R10915 gnd.n5025 gnd.n4876 240.244
R10916 gnd.n5025 gnd.n4871 240.244
R10917 gnd.n5135 gnd.n4871 240.244
R10918 gnd.n5135 gnd.n4872 240.244
R10919 gnd.n4872 gnd.n4819 240.244
R10920 gnd.n5130 gnd.n4819 240.244
R10921 gnd.n5130 gnd.n5129 240.244
R10922 gnd.n5129 gnd.n4798 240.244
R10923 gnd.n5125 gnd.n4798 240.244
R10924 gnd.n5125 gnd.n4789 240.244
R10925 gnd.n5122 gnd.n4789 240.244
R10926 gnd.n5122 gnd.n5121 240.244
R10927 gnd.n5121 gnd.n4772 240.244
R10928 gnd.n5117 gnd.n4772 240.244
R10929 gnd.n5117 gnd.n4763 240.244
R10930 gnd.n5114 gnd.n4763 240.244
R10931 gnd.n5114 gnd.n5113 240.244
R10932 gnd.n5113 gnd.n4748 240.244
R10933 gnd.n5108 gnd.n4748 240.244
R10934 gnd.n5108 gnd.n4738 240.244
R10935 gnd.n5105 gnd.n4738 240.244
R10936 gnd.n5105 gnd.n5104 240.244
R10937 gnd.n5104 gnd.n4722 240.244
R10938 gnd.n5049 gnd.n4722 240.244
R10939 gnd.n5049 gnd.n4712 240.244
R10940 gnd.n5060 gnd.n4712 240.244
R10941 gnd.n5060 gnd.n5058 240.244
R10942 gnd.n5058 gnd.n4697 240.244
R10943 gnd.n5053 gnd.n4697 240.244
R10944 gnd.n5053 gnd.n4688 240.244
R10945 gnd.n4688 gnd.n4671 240.244
R10946 gnd.n5323 gnd.n4671 240.244
R10947 gnd.n5323 gnd.n4667 240.244
R10948 gnd.n5344 gnd.n4667 240.244
R10949 gnd.n5344 gnd.n4656 240.244
R10950 gnd.n5340 gnd.n4656 240.244
R10951 gnd.n5340 gnd.n4646 240.244
R10952 gnd.n5337 gnd.n4646 240.244
R10953 gnd.n5337 gnd.n4636 240.244
R10954 gnd.n5334 gnd.n4636 240.244
R10955 gnd.n5334 gnd.n4615 240.244
R10956 gnd.n5410 gnd.n4615 240.244
R10957 gnd.n5410 gnd.n4611 240.244
R10958 gnd.n5428 gnd.n4611 240.244
R10959 gnd.n5428 gnd.n4602 240.244
R10960 gnd.n5424 gnd.n4602 240.244
R10961 gnd.n5424 gnd.n4596 240.244
R10962 gnd.n5421 gnd.n4596 240.244
R10963 gnd.n5421 gnd.n4582 240.244
R10964 gnd.n4582 gnd.n4572 240.244
R10965 gnd.n5769 gnd.n4572 240.244
R10966 gnd.n5769 gnd.n766 240.244
R10967 gnd.n5775 gnd.n766 240.244
R10968 gnd.n5775 gnd.n777 240.244
R10969 gnd.n5779 gnd.n777 240.244
R10970 gnd.n5779 gnd.n5778 240.244
R10971 gnd.n5778 gnd.n790 240.244
R10972 gnd.n5786 gnd.n790 240.244
R10973 gnd.n5786 gnd.n800 240.244
R10974 gnd.n4912 gnd.n4911 240.244
R10975 gnd.n4983 gnd.n4911 240.244
R10976 gnd.n4981 gnd.n4980 240.244
R10977 gnd.n4977 gnd.n4976 240.244
R10978 gnd.n4973 gnd.n4972 240.244
R10979 gnd.n4969 gnd.n4968 240.244
R10980 gnd.n4965 gnd.n4964 240.244
R10981 gnd.n4961 gnd.n4960 240.244
R10982 gnd.n4957 gnd.n4956 240.244
R10983 gnd.n4953 gnd.n4952 240.244
R10984 gnd.n4949 gnd.n4948 240.244
R10985 gnd.n4945 gnd.n4944 240.244
R10986 gnd.n4941 gnd.n4899 240.244
R10987 gnd.n5001 gnd.n4893 240.244
R10988 gnd.n5001 gnd.n4889 240.244
R10989 gnd.n5007 gnd.n4889 240.244
R10990 gnd.n5007 gnd.n4882 240.244
R10991 gnd.n5017 gnd.n4882 240.244
R10992 gnd.n5017 gnd.n4878 240.244
R10993 gnd.n5023 gnd.n4878 240.244
R10994 gnd.n5023 gnd.n4869 240.244
R10995 gnd.n5137 gnd.n4869 240.244
R10996 gnd.n5137 gnd.n4820 240.244
R10997 gnd.n5145 gnd.n4820 240.244
R10998 gnd.n5145 gnd.n4821 240.244
R10999 gnd.n4821 gnd.n4799 240.244
R11000 gnd.n5166 gnd.n4799 240.244
R11001 gnd.n5166 gnd.n4791 240.244
R11002 gnd.n5177 gnd.n4791 240.244
R11003 gnd.n5177 gnd.n4792 240.244
R11004 gnd.n4792 gnd.n4773 240.244
R11005 gnd.n5197 gnd.n4773 240.244
R11006 gnd.n5197 gnd.n4765 240.244
R11007 gnd.n5208 gnd.n4765 240.244
R11008 gnd.n5208 gnd.n4766 240.244
R11009 gnd.n4766 gnd.n4749 240.244
R11010 gnd.n5228 gnd.n4749 240.244
R11011 gnd.n5228 gnd.n4740 240.244
R11012 gnd.n5239 gnd.n4740 240.244
R11013 gnd.n5239 gnd.n4741 240.244
R11014 gnd.n4741 gnd.n4723 240.244
R11015 gnd.n5259 gnd.n4723 240.244
R11016 gnd.n5259 gnd.n4714 240.244
R11017 gnd.n5270 gnd.n4714 240.244
R11018 gnd.n5270 gnd.n4715 240.244
R11019 gnd.n4715 gnd.n4698 240.244
R11020 gnd.n5290 gnd.n4698 240.244
R11021 gnd.n5290 gnd.n4690 240.244
R11022 gnd.n5300 gnd.n4690 240.244
R11023 gnd.n5300 gnd.n4673 240.244
R11024 gnd.n5321 gnd.n4673 240.244
R11025 gnd.n5321 gnd.n4674 240.244
R11026 gnd.n4674 gnd.n4658 240.244
R11027 gnd.n5354 gnd.n4658 240.244
R11028 gnd.n5354 gnd.n4645 240.244
R11029 gnd.n5369 gnd.n4645 240.244
R11030 gnd.n5369 gnd.n4638 240.244
R11031 gnd.n5384 gnd.n4638 240.244
R11032 gnd.n5384 gnd.n4639 240.244
R11033 gnd.n4639 gnd.n4617 240.244
R11034 gnd.n5408 gnd.n4617 240.244
R11035 gnd.n5408 gnd.n4618 240.244
R11036 gnd.n4618 gnd.n4601 240.244
R11037 gnd.n5444 gnd.n4601 240.244
R11038 gnd.n5444 gnd.n4594 240.244
R11039 gnd.n5455 gnd.n4594 240.244
R11040 gnd.n5455 gnd.n4584 240.244
R11041 gnd.n5751 gnd.n4584 240.244
R11042 gnd.n5751 gnd.n4586 240.244
R11043 gnd.n4586 gnd.n768 240.244
R11044 gnd.n5894 gnd.n768 240.244
R11045 gnd.n5894 gnd.n769 240.244
R11046 gnd.n5890 gnd.n769 240.244
R11047 gnd.n5890 gnd.n775 240.244
R11048 gnd.n792 gnd.n775 240.244
R11049 gnd.n5880 gnd.n792 240.244
R11050 gnd.n5880 gnd.n793 240.244
R11051 gnd.n5876 gnd.n793 240.244
R11052 gnd.n6720 gnd.n6719 240.244
R11053 gnd.n6725 gnd.n6722 240.244
R11054 gnd.n6728 gnd.n6727 240.244
R11055 gnd.n6733 gnd.n6730 240.244
R11056 gnd.n6736 gnd.n6735 240.244
R11057 gnd.n6741 gnd.n6738 240.244
R11058 gnd.n6744 gnd.n6743 240.244
R11059 gnd.n6749 gnd.n6746 240.244
R11060 gnd.n6755 gnd.n6751 240.244
R11061 gnd.n3891 gnd.n1214 240.244
R11062 gnd.n3891 gnd.n1226 240.244
R11063 gnd.n3898 gnd.n1226 240.244
R11064 gnd.n3898 gnd.n1327 240.244
R11065 gnd.n1327 gnd.n1317 240.244
R11066 gnd.n4021 gnd.n1317 240.244
R11067 gnd.n4021 gnd.n1312 240.244
R11068 gnd.n4028 gnd.n1312 240.244
R11069 gnd.n4028 gnd.n1301 240.244
R11070 gnd.n1301 gnd.n1288 240.244
R11071 gnd.n4053 gnd.n1288 240.244
R11072 gnd.n4053 gnd.n1283 240.244
R11073 gnd.n4060 gnd.n1283 240.244
R11074 gnd.n4060 gnd.n1272 240.244
R11075 gnd.n1272 gnd.n1259 240.244
R11076 gnd.n4087 gnd.n1259 240.244
R11077 gnd.n4087 gnd.n1253 240.244
R11078 gnd.n4094 gnd.n1253 240.244
R11079 gnd.n4094 gnd.n250 240.244
R11080 gnd.n250 gnd.n245 240.244
R11081 gnd.n3965 gnd.n245 240.244
R11082 gnd.n3965 gnd.n54 240.244
R11083 gnd.n55 gnd.n54 240.244
R11084 gnd.n56 gnd.n55 240.244
R11085 gnd.n221 gnd.n56 240.244
R11086 gnd.n221 gnd.n59 240.244
R11087 gnd.n60 gnd.n59 240.244
R11088 gnd.n61 gnd.n60 240.244
R11089 gnd.n201 gnd.n61 240.244
R11090 gnd.n201 gnd.n64 240.244
R11091 gnd.n65 gnd.n64 240.244
R11092 gnd.n66 gnd.n65 240.244
R11093 gnd.n185 gnd.n66 240.244
R11094 gnd.n185 gnd.n69 240.244
R11095 gnd.n70 gnd.n69 240.244
R11096 gnd.n71 gnd.n70 240.244
R11097 gnd.n169 gnd.n71 240.244
R11098 gnd.n169 gnd.n74 240.244
R11099 gnd.n75 gnd.n74 240.244
R11100 gnd.n76 gnd.n75 240.244
R11101 gnd.n79 gnd.n76 240.244
R11102 gnd.n6882 gnd.n79 240.244
R11103 gnd.n3475 gnd.n3473 240.244
R11104 gnd.n3490 gnd.n3456 240.244
R11105 gnd.n3494 gnd.n3492 240.244
R11106 gnd.n3509 gnd.n3447 240.244
R11107 gnd.n3513 gnd.n3511 240.244
R11108 gnd.n3528 gnd.n3438 240.244
R11109 gnd.n3532 gnd.n3530 240.244
R11110 gnd.n3549 gnd.n3429 240.244
R11111 gnd.n3552 gnd.n3551 240.244
R11112 gnd.n1228 gnd.n1216 240.244
R11113 gnd.n4123 gnd.n1228 240.244
R11114 gnd.n4123 gnd.n1229 240.244
R11115 gnd.n1234 gnd.n1229 240.244
R11116 gnd.n1235 gnd.n1234 240.244
R11117 gnd.n1236 gnd.n1235 240.244
R11118 gnd.n1309 gnd.n1236 240.244
R11119 gnd.n1309 gnd.n1239 240.244
R11120 gnd.n1240 gnd.n1239 240.244
R11121 gnd.n1241 gnd.n1240 240.244
R11122 gnd.n1292 gnd.n1241 240.244
R11123 gnd.n1292 gnd.n1244 240.244
R11124 gnd.n1245 gnd.n1244 240.244
R11125 gnd.n1246 gnd.n1245 240.244
R11126 gnd.n1273 gnd.n1246 240.244
R11127 gnd.n1273 gnd.n1249 240.244
R11128 gnd.n1250 gnd.n1249 240.244
R11129 gnd.n4096 gnd.n1250 240.244
R11130 gnd.n4096 gnd.n243 240.244
R11131 gnd.n6650 gnd.n243 240.244
R11132 gnd.n6650 gnd.n238 240.244
R11133 gnd.n6656 gnd.n238 240.244
R11134 gnd.n6656 gnd.n229 240.244
R11135 gnd.n6664 gnd.n229 240.244
R11136 gnd.n6664 gnd.n225 240.244
R11137 gnd.n6670 gnd.n225 240.244
R11138 gnd.n6670 gnd.n208 240.244
R11139 gnd.n6680 gnd.n208 240.244
R11140 gnd.n6680 gnd.n204 240.244
R11141 gnd.n6686 gnd.n204 240.244
R11142 gnd.n6686 gnd.n193 240.244
R11143 gnd.n6696 gnd.n193 240.244
R11144 gnd.n6696 gnd.n189 240.244
R11145 gnd.n6702 gnd.n189 240.244
R11146 gnd.n6702 gnd.n178 240.244
R11147 gnd.n6712 gnd.n178 240.244
R11148 gnd.n6712 gnd.n172 240.244
R11149 gnd.n6792 gnd.n172 240.244
R11150 gnd.n6792 gnd.n173 240.244
R11151 gnd.n173 gnd.n163 240.244
R11152 gnd.n6717 gnd.n163 240.244
R11153 gnd.n6717 gnd.n84 240.244
R11154 gnd.n2097 gnd.n1083 240.244
R11155 gnd.n2100 gnd.n2099 240.244
R11156 gnd.n2110 gnd.n2102 240.244
R11157 gnd.n2113 gnd.n2112 240.244
R11158 gnd.n2122 gnd.n2121 240.244
R11159 gnd.n2133 gnd.n2124 240.244
R11160 gnd.n2136 gnd.n2135 240.244
R11161 gnd.n2145 gnd.n2144 240.244
R11162 gnd.n2156 gnd.n2147 240.244
R11163 gnd.n2352 gnd.n2271 240.244
R11164 gnd.n2353 gnd.n2352 240.244
R11165 gnd.n2353 gnd.n885 240.244
R11166 gnd.n2267 gnd.n885 240.244
R11167 gnd.n2267 gnd.n897 240.244
R11168 gnd.n2360 gnd.n897 240.244
R11169 gnd.n2360 gnd.n908 240.244
R11170 gnd.n2264 gnd.n908 240.244
R11171 gnd.n2264 gnd.n918 240.244
R11172 gnd.n2367 gnd.n918 240.244
R11173 gnd.n2367 gnd.n928 240.244
R11174 gnd.n2261 gnd.n928 240.244
R11175 gnd.n2261 gnd.n938 240.244
R11176 gnd.n2374 gnd.n938 240.244
R11177 gnd.n2374 gnd.n948 240.244
R11178 gnd.n2380 gnd.n948 240.244
R11179 gnd.n2421 gnd.n2380 240.244
R11180 gnd.n2421 gnd.n959 240.244
R11181 gnd.n2424 gnd.n959 240.244
R11182 gnd.n2424 gnd.n972 240.244
R11183 gnd.n2430 gnd.n972 240.244
R11184 gnd.n2430 gnd.n980 240.244
R11185 gnd.n2452 gnd.n980 240.244
R11186 gnd.n2452 gnd.n989 240.244
R11187 gnd.n2446 gnd.n989 240.244
R11188 gnd.n2446 gnd.n997 240.244
R11189 gnd.n2503 gnd.n997 240.244
R11190 gnd.n2503 gnd.n1007 240.244
R11191 gnd.n2509 gnd.n1007 240.244
R11192 gnd.n2509 gnd.n1018 240.244
R11193 gnd.n2519 gnd.n1018 240.244
R11194 gnd.n2519 gnd.n1028 240.244
R11195 gnd.n2525 gnd.n1028 240.244
R11196 gnd.n2525 gnd.n1039 240.244
R11197 gnd.n2553 gnd.n1039 240.244
R11198 gnd.n2553 gnd.n1049 240.244
R11199 gnd.n2226 gnd.n1049 240.244
R11200 gnd.n2226 gnd.n1060 240.244
R11201 gnd.n2544 gnd.n1060 240.244
R11202 gnd.n2544 gnd.n1071 240.244
R11203 gnd.n2661 gnd.n1071 240.244
R11204 gnd.n2661 gnd.n1081 240.244
R11205 gnd.n2332 gnd.n2331 240.244
R11206 gnd.n2328 gnd.n2327 240.244
R11207 gnd.n2324 gnd.n2323 240.244
R11208 gnd.n2320 gnd.n2319 240.244
R11209 gnd.n2316 gnd.n2315 240.244
R11210 gnd.n2312 gnd.n2311 240.244
R11211 gnd.n2308 gnd.n2307 240.244
R11212 gnd.n2304 gnd.n2303 240.244
R11213 gnd.n2291 gnd.n829 240.244
R11214 gnd.n2344 gnd.n2272 240.244
R11215 gnd.n2344 gnd.n2273 240.244
R11216 gnd.n2273 gnd.n887 240.244
R11217 gnd.n899 gnd.n887 240.244
R11218 gnd.n4388 gnd.n899 240.244
R11219 gnd.n4388 gnd.n900 240.244
R11220 gnd.n4384 gnd.n900 240.244
R11221 gnd.n4384 gnd.n906 240.244
R11222 gnd.n4376 gnd.n906 240.244
R11223 gnd.n4376 gnd.n919 240.244
R11224 gnd.n4372 gnd.n919 240.244
R11225 gnd.n4372 gnd.n925 240.244
R11226 gnd.n4364 gnd.n925 240.244
R11227 gnd.n4364 gnd.n940 240.244
R11228 gnd.n4360 gnd.n940 240.244
R11229 gnd.n4360 gnd.n946 240.244
R11230 gnd.n961 gnd.n946 240.244
R11231 gnd.n4350 gnd.n961 240.244
R11232 gnd.n4350 gnd.n962 240.244
R11233 gnd.n4346 gnd.n962 240.244
R11234 gnd.n4346 gnd.n970 240.244
R11235 gnd.n4337 gnd.n970 240.244
R11236 gnd.n4337 gnd.n981 240.244
R11237 gnd.n4333 gnd.n981 240.244
R11238 gnd.n4333 gnd.n986 240.244
R11239 gnd.n4324 gnd.n986 240.244
R11240 gnd.n4324 gnd.n999 240.244
R11241 gnd.n4320 gnd.n999 240.244
R11242 gnd.n4320 gnd.n1005 240.244
R11243 gnd.n4312 gnd.n1005 240.244
R11244 gnd.n4312 gnd.n1019 240.244
R11245 gnd.n4308 gnd.n1019 240.244
R11246 gnd.n4308 gnd.n1025 240.244
R11247 gnd.n4300 gnd.n1025 240.244
R11248 gnd.n4300 gnd.n1041 240.244
R11249 gnd.n4296 gnd.n1041 240.244
R11250 gnd.n4296 gnd.n1047 240.244
R11251 gnd.n4288 gnd.n1047 240.244
R11252 gnd.n4288 gnd.n1062 240.244
R11253 gnd.n4284 gnd.n1062 240.244
R11254 gnd.n4284 gnd.n1068 240.244
R11255 gnd.n4276 gnd.n1068 240.244
R11256 gnd.n6066 gnd.n593 240.244
R11257 gnd.n6072 gnd.n593 240.244
R11258 gnd.n6072 gnd.n591 240.244
R11259 gnd.n6076 gnd.n591 240.244
R11260 gnd.n6076 gnd.n587 240.244
R11261 gnd.n6082 gnd.n587 240.244
R11262 gnd.n6082 gnd.n585 240.244
R11263 gnd.n6086 gnd.n585 240.244
R11264 gnd.n6086 gnd.n581 240.244
R11265 gnd.n6092 gnd.n581 240.244
R11266 gnd.n6092 gnd.n579 240.244
R11267 gnd.n6096 gnd.n579 240.244
R11268 gnd.n6096 gnd.n575 240.244
R11269 gnd.n6102 gnd.n575 240.244
R11270 gnd.n6102 gnd.n573 240.244
R11271 gnd.n6106 gnd.n573 240.244
R11272 gnd.n6106 gnd.n569 240.244
R11273 gnd.n6112 gnd.n569 240.244
R11274 gnd.n6112 gnd.n567 240.244
R11275 gnd.n6116 gnd.n567 240.244
R11276 gnd.n6116 gnd.n563 240.244
R11277 gnd.n6122 gnd.n563 240.244
R11278 gnd.n6122 gnd.n561 240.244
R11279 gnd.n6126 gnd.n561 240.244
R11280 gnd.n6126 gnd.n557 240.244
R11281 gnd.n6132 gnd.n557 240.244
R11282 gnd.n6132 gnd.n555 240.244
R11283 gnd.n6136 gnd.n555 240.244
R11284 gnd.n6136 gnd.n551 240.244
R11285 gnd.n6142 gnd.n551 240.244
R11286 gnd.n6142 gnd.n549 240.244
R11287 gnd.n6146 gnd.n549 240.244
R11288 gnd.n6146 gnd.n545 240.244
R11289 gnd.n6152 gnd.n545 240.244
R11290 gnd.n6152 gnd.n543 240.244
R11291 gnd.n6156 gnd.n543 240.244
R11292 gnd.n6156 gnd.n539 240.244
R11293 gnd.n6162 gnd.n539 240.244
R11294 gnd.n6162 gnd.n537 240.244
R11295 gnd.n6166 gnd.n537 240.244
R11296 gnd.n6166 gnd.n533 240.244
R11297 gnd.n6172 gnd.n533 240.244
R11298 gnd.n6172 gnd.n531 240.244
R11299 gnd.n6176 gnd.n531 240.244
R11300 gnd.n6176 gnd.n527 240.244
R11301 gnd.n6182 gnd.n527 240.244
R11302 gnd.n6182 gnd.n525 240.244
R11303 gnd.n6186 gnd.n525 240.244
R11304 gnd.n6186 gnd.n521 240.244
R11305 gnd.n6192 gnd.n521 240.244
R11306 gnd.n6192 gnd.n519 240.244
R11307 gnd.n6196 gnd.n519 240.244
R11308 gnd.n6196 gnd.n515 240.244
R11309 gnd.n6202 gnd.n515 240.244
R11310 gnd.n6202 gnd.n513 240.244
R11311 gnd.n6206 gnd.n513 240.244
R11312 gnd.n6206 gnd.n509 240.244
R11313 gnd.n6212 gnd.n509 240.244
R11314 gnd.n6212 gnd.n507 240.244
R11315 gnd.n6216 gnd.n507 240.244
R11316 gnd.n6216 gnd.n503 240.244
R11317 gnd.n6222 gnd.n503 240.244
R11318 gnd.n6222 gnd.n501 240.244
R11319 gnd.n6226 gnd.n501 240.244
R11320 gnd.n6226 gnd.n497 240.244
R11321 gnd.n6232 gnd.n497 240.244
R11322 gnd.n6232 gnd.n495 240.244
R11323 gnd.n6236 gnd.n495 240.244
R11324 gnd.n6236 gnd.n491 240.244
R11325 gnd.n6242 gnd.n491 240.244
R11326 gnd.n6242 gnd.n489 240.244
R11327 gnd.n6246 gnd.n489 240.244
R11328 gnd.n6246 gnd.n485 240.244
R11329 gnd.n6252 gnd.n485 240.244
R11330 gnd.n6252 gnd.n483 240.244
R11331 gnd.n6256 gnd.n483 240.244
R11332 gnd.n6256 gnd.n479 240.244
R11333 gnd.n6262 gnd.n479 240.244
R11334 gnd.n6262 gnd.n477 240.244
R11335 gnd.n6266 gnd.n477 240.244
R11336 gnd.n6266 gnd.n473 240.244
R11337 gnd.n6272 gnd.n473 240.244
R11338 gnd.n6272 gnd.n471 240.244
R11339 gnd.n6276 gnd.n471 240.244
R11340 gnd.n6276 gnd.n467 240.244
R11341 gnd.n6282 gnd.n467 240.244
R11342 gnd.n6282 gnd.n465 240.244
R11343 gnd.n6286 gnd.n465 240.244
R11344 gnd.n6286 gnd.n461 240.244
R11345 gnd.n6292 gnd.n461 240.244
R11346 gnd.n6292 gnd.n459 240.244
R11347 gnd.n6296 gnd.n459 240.244
R11348 gnd.n6296 gnd.n455 240.244
R11349 gnd.n6302 gnd.n455 240.244
R11350 gnd.n6302 gnd.n453 240.244
R11351 gnd.n6306 gnd.n453 240.244
R11352 gnd.n6306 gnd.n449 240.244
R11353 gnd.n6312 gnd.n449 240.244
R11354 gnd.n6312 gnd.n447 240.244
R11355 gnd.n6316 gnd.n447 240.244
R11356 gnd.n6316 gnd.n443 240.244
R11357 gnd.n6322 gnd.n443 240.244
R11358 gnd.n6322 gnd.n441 240.244
R11359 gnd.n6326 gnd.n441 240.244
R11360 gnd.n6326 gnd.n437 240.244
R11361 gnd.n6332 gnd.n437 240.244
R11362 gnd.n6332 gnd.n435 240.244
R11363 gnd.n6336 gnd.n435 240.244
R11364 gnd.n6336 gnd.n431 240.244
R11365 gnd.n6342 gnd.n431 240.244
R11366 gnd.n6342 gnd.n429 240.244
R11367 gnd.n6346 gnd.n429 240.244
R11368 gnd.n6346 gnd.n425 240.244
R11369 gnd.n6352 gnd.n425 240.244
R11370 gnd.n6352 gnd.n423 240.244
R11371 gnd.n6356 gnd.n423 240.244
R11372 gnd.n6356 gnd.n419 240.244
R11373 gnd.n6362 gnd.n419 240.244
R11374 gnd.n6362 gnd.n417 240.244
R11375 gnd.n6366 gnd.n417 240.244
R11376 gnd.n6366 gnd.n413 240.244
R11377 gnd.n6372 gnd.n413 240.244
R11378 gnd.n6372 gnd.n411 240.244
R11379 gnd.n6376 gnd.n411 240.244
R11380 gnd.n6376 gnd.n407 240.244
R11381 gnd.n6382 gnd.n407 240.244
R11382 gnd.n6382 gnd.n405 240.244
R11383 gnd.n6386 gnd.n405 240.244
R11384 gnd.n6386 gnd.n401 240.244
R11385 gnd.n6392 gnd.n401 240.244
R11386 gnd.n6392 gnd.n399 240.244
R11387 gnd.n6396 gnd.n399 240.244
R11388 gnd.n6396 gnd.n395 240.244
R11389 gnd.n6402 gnd.n395 240.244
R11390 gnd.n6402 gnd.n393 240.244
R11391 gnd.n6406 gnd.n393 240.244
R11392 gnd.n6406 gnd.n389 240.244
R11393 gnd.n6413 gnd.n389 240.244
R11394 gnd.n6413 gnd.n387 240.244
R11395 gnd.n6417 gnd.n387 240.244
R11396 gnd.n6417 gnd.n384 240.244
R11397 gnd.n6423 gnd.n382 240.244
R11398 gnd.n6427 gnd.n382 240.244
R11399 gnd.n6427 gnd.n378 240.244
R11400 gnd.n6433 gnd.n378 240.244
R11401 gnd.n6433 gnd.n376 240.244
R11402 gnd.n6437 gnd.n376 240.244
R11403 gnd.n6437 gnd.n372 240.244
R11404 gnd.n6443 gnd.n372 240.244
R11405 gnd.n6443 gnd.n370 240.244
R11406 gnd.n6447 gnd.n370 240.244
R11407 gnd.n6447 gnd.n366 240.244
R11408 gnd.n6453 gnd.n366 240.244
R11409 gnd.n6453 gnd.n364 240.244
R11410 gnd.n6457 gnd.n364 240.244
R11411 gnd.n6457 gnd.n360 240.244
R11412 gnd.n6463 gnd.n360 240.244
R11413 gnd.n6463 gnd.n358 240.244
R11414 gnd.n6467 gnd.n358 240.244
R11415 gnd.n6467 gnd.n354 240.244
R11416 gnd.n6473 gnd.n354 240.244
R11417 gnd.n6473 gnd.n352 240.244
R11418 gnd.n6477 gnd.n352 240.244
R11419 gnd.n6477 gnd.n348 240.244
R11420 gnd.n6483 gnd.n348 240.244
R11421 gnd.n6483 gnd.n346 240.244
R11422 gnd.n6487 gnd.n346 240.244
R11423 gnd.n6487 gnd.n342 240.244
R11424 gnd.n6493 gnd.n342 240.244
R11425 gnd.n6493 gnd.n340 240.244
R11426 gnd.n6497 gnd.n340 240.244
R11427 gnd.n6497 gnd.n336 240.244
R11428 gnd.n6503 gnd.n336 240.244
R11429 gnd.n6503 gnd.n334 240.244
R11430 gnd.n6507 gnd.n334 240.244
R11431 gnd.n6507 gnd.n330 240.244
R11432 gnd.n6513 gnd.n330 240.244
R11433 gnd.n6513 gnd.n328 240.244
R11434 gnd.n6517 gnd.n328 240.244
R11435 gnd.n6517 gnd.n324 240.244
R11436 gnd.n6523 gnd.n324 240.244
R11437 gnd.n6523 gnd.n322 240.244
R11438 gnd.n6527 gnd.n322 240.244
R11439 gnd.n6527 gnd.n318 240.244
R11440 gnd.n6533 gnd.n318 240.244
R11441 gnd.n6533 gnd.n316 240.244
R11442 gnd.n6537 gnd.n316 240.244
R11443 gnd.n6537 gnd.n312 240.244
R11444 gnd.n6543 gnd.n312 240.244
R11445 gnd.n6543 gnd.n310 240.244
R11446 gnd.n6547 gnd.n310 240.244
R11447 gnd.n6547 gnd.n306 240.244
R11448 gnd.n6553 gnd.n306 240.244
R11449 gnd.n6553 gnd.n304 240.244
R11450 gnd.n6557 gnd.n304 240.244
R11451 gnd.n6557 gnd.n300 240.244
R11452 gnd.n6563 gnd.n300 240.244
R11453 gnd.n6563 gnd.n298 240.244
R11454 gnd.n6567 gnd.n298 240.244
R11455 gnd.n6567 gnd.n294 240.244
R11456 gnd.n6573 gnd.n294 240.244
R11457 gnd.n6573 gnd.n292 240.244
R11458 gnd.n6577 gnd.n292 240.244
R11459 gnd.n6577 gnd.n288 240.244
R11460 gnd.n6583 gnd.n288 240.244
R11461 gnd.n6583 gnd.n286 240.244
R11462 gnd.n6587 gnd.n286 240.244
R11463 gnd.n6587 gnd.n282 240.244
R11464 gnd.n6593 gnd.n282 240.244
R11465 gnd.n6593 gnd.n280 240.244
R11466 gnd.n6597 gnd.n280 240.244
R11467 gnd.n6597 gnd.n276 240.244
R11468 gnd.n6603 gnd.n276 240.244
R11469 gnd.n6603 gnd.n274 240.244
R11470 gnd.n6607 gnd.n274 240.244
R11471 gnd.n6607 gnd.n270 240.244
R11472 gnd.n6613 gnd.n270 240.244
R11473 gnd.n6613 gnd.n268 240.244
R11474 gnd.n6617 gnd.n268 240.244
R11475 gnd.n6617 gnd.n264 240.244
R11476 gnd.n6623 gnd.n264 240.244
R11477 gnd.n6623 gnd.n262 240.244
R11478 gnd.n6628 gnd.n262 240.244
R11479 gnd.n6628 gnd.n258 240.244
R11480 gnd.n6635 gnd.n258 240.244
R11481 gnd.n2464 gnd.n2463 240.244
R11482 gnd.n2465 gnd.n2464 240.244
R11483 gnd.n2465 gnd.n2455 240.244
R11484 gnd.n2472 gnd.n2455 240.244
R11485 gnd.n2473 gnd.n2472 240.244
R11486 gnd.n2474 gnd.n2473 240.244
R11487 gnd.n2474 gnd.n2243 240.244
R11488 gnd.n2500 gnd.n2243 240.244
R11489 gnd.n2500 gnd.n2244 240.244
R11490 gnd.n2496 gnd.n2244 240.244
R11491 gnd.n2496 gnd.n2495 240.244
R11492 gnd.n2495 gnd.n2494 240.244
R11493 gnd.n2494 gnd.n2482 240.244
R11494 gnd.n2490 gnd.n2482 240.244
R11495 gnd.n2490 gnd.n2219 240.244
R11496 gnd.n2556 gnd.n2219 240.244
R11497 gnd.n2557 gnd.n2556 240.244
R11498 gnd.n2558 gnd.n2557 240.244
R11499 gnd.n2558 gnd.n2215 240.244
R11500 gnd.n2564 gnd.n2215 240.244
R11501 gnd.n2565 gnd.n2564 240.244
R11502 gnd.n2566 gnd.n2565 240.244
R11503 gnd.n2566 gnd.n2211 240.244
R11504 gnd.n2573 gnd.n2211 240.244
R11505 gnd.n2574 gnd.n2573 240.244
R11506 gnd.n2578 gnd.n2574 240.244
R11507 gnd.n2578 gnd.n2207 240.244
R11508 gnd.n2584 gnd.n2207 240.244
R11509 gnd.n2584 gnd.n2073 240.244
R11510 gnd.n2591 gnd.n2073 240.244
R11511 gnd.n2591 gnd.n2069 240.244
R11512 gnd.n2597 gnd.n2069 240.244
R11513 gnd.n2597 gnd.n2067 240.244
R11514 gnd.n2606 gnd.n2067 240.244
R11515 gnd.n2606 gnd.n2062 240.244
R11516 gnd.n2622 gnd.n2062 240.244
R11517 gnd.n2622 gnd.n2063 240.244
R11518 gnd.n2618 gnd.n2063 240.244
R11519 gnd.n2618 gnd.n2615 240.244
R11520 gnd.n2615 gnd.n1773 240.244
R11521 gnd.n2801 gnd.n1773 240.244
R11522 gnd.n2801 gnd.n1769 240.244
R11523 gnd.n2807 gnd.n1769 240.244
R11524 gnd.n2807 gnd.n1745 240.244
R11525 gnd.n2844 gnd.n1745 240.244
R11526 gnd.n2844 gnd.n1741 240.244
R11527 gnd.n2850 gnd.n1741 240.244
R11528 gnd.n2850 gnd.n1727 240.244
R11529 gnd.n2886 gnd.n1727 240.244
R11530 gnd.n2886 gnd.n1722 240.244
R11531 gnd.n2894 gnd.n1722 240.244
R11532 gnd.n2894 gnd.n1723 240.244
R11533 gnd.n1723 gnd.n1701 240.244
R11534 gnd.n2948 gnd.n1701 240.244
R11535 gnd.n2948 gnd.n1697 240.244
R11536 gnd.n2954 gnd.n1697 240.244
R11537 gnd.n2954 gnd.n1683 240.244
R11538 gnd.n2975 gnd.n1683 240.244
R11539 gnd.n2975 gnd.n1678 240.244
R11540 gnd.n2983 gnd.n1678 240.244
R11541 gnd.n2983 gnd.n1679 240.244
R11542 gnd.n1679 gnd.n1650 240.244
R11543 gnd.n3026 gnd.n1650 240.244
R11544 gnd.n3026 gnd.n1646 240.244
R11545 gnd.n3032 gnd.n1646 240.244
R11546 gnd.n3032 gnd.n1627 240.244
R11547 gnd.n3066 gnd.n1627 240.244
R11548 gnd.n3066 gnd.n1623 240.244
R11549 gnd.n3072 gnd.n1623 240.244
R11550 gnd.n3072 gnd.n1605 240.244
R11551 gnd.n3122 gnd.n1605 240.244
R11552 gnd.n3122 gnd.n1601 240.244
R11553 gnd.n3128 gnd.n1601 240.244
R11554 gnd.n3128 gnd.n1586 240.244
R11555 gnd.n3147 gnd.n1586 240.244
R11556 gnd.n3147 gnd.n1582 240.244
R11557 gnd.n3153 gnd.n1582 240.244
R11558 gnd.n3153 gnd.n1566 240.244
R11559 gnd.n3207 gnd.n1566 240.244
R11560 gnd.n3207 gnd.n1562 240.244
R11561 gnd.n3213 gnd.n1562 240.244
R11562 gnd.n3213 gnd.n1544 240.244
R11563 gnd.n3236 gnd.n1544 240.244
R11564 gnd.n3236 gnd.n1539 240.244
R11565 gnd.n3244 gnd.n1539 240.244
R11566 gnd.n3244 gnd.n1540 240.244
R11567 gnd.n1540 gnd.n1516 240.244
R11568 gnd.n3289 gnd.n1516 240.244
R11569 gnd.n3289 gnd.n1512 240.244
R11570 gnd.n3295 gnd.n1512 240.244
R11571 gnd.n3295 gnd.n1497 240.244
R11572 gnd.n3316 gnd.n1497 240.244
R11573 gnd.n3316 gnd.n1492 240.244
R11574 gnd.n3324 gnd.n1492 240.244
R11575 gnd.n3324 gnd.n1493 240.244
R11576 gnd.n1493 gnd.n1467 240.244
R11577 gnd.n3360 gnd.n1467 240.244
R11578 gnd.n3360 gnd.n1461 240.244
R11579 gnd.n3369 gnd.n1461 240.244
R11580 gnd.n3369 gnd.n1463 240.244
R11581 gnd.n1463 gnd.n1411 240.244
R11582 gnd.n3611 gnd.n1411 240.244
R11583 gnd.n3611 gnd.n1412 240.244
R11584 gnd.n3607 gnd.n1412 240.244
R11585 gnd.n3607 gnd.n3606 240.244
R11586 gnd.n3606 gnd.n1418 240.244
R11587 gnd.n3600 gnd.n1418 240.244
R11588 gnd.n3600 gnd.n1424 240.244
R11589 gnd.n3596 gnd.n1424 240.244
R11590 gnd.n3596 gnd.n1434 240.244
R11591 gnd.n1434 gnd.n1195 240.244
R11592 gnd.n4144 gnd.n1195 240.244
R11593 gnd.n4144 gnd.n1196 240.244
R11594 gnd.n4140 gnd.n1196 240.244
R11595 gnd.n4140 gnd.n1202 240.244
R11596 gnd.n4136 gnd.n1202 240.244
R11597 gnd.n4136 gnd.n1205 240.244
R11598 gnd.n4132 gnd.n1205 240.244
R11599 gnd.n4132 gnd.n1211 240.244
R11600 gnd.n3999 gnd.n1211 240.244
R11601 gnd.n4000 gnd.n3999 240.244
R11602 gnd.n4000 gnd.n3993 240.244
R11603 gnd.n4008 gnd.n3993 240.244
R11604 gnd.n4008 gnd.n3994 240.244
R11605 gnd.n3994 gnd.n1308 240.244
R11606 gnd.n4031 gnd.n1308 240.244
R11607 gnd.n4031 gnd.n1303 240.244
R11608 gnd.n4039 gnd.n1303 240.244
R11609 gnd.n4039 gnd.n1304 240.244
R11610 gnd.n1304 gnd.n1280 240.244
R11611 gnd.n4063 gnd.n1280 240.244
R11612 gnd.n4063 gnd.n1275 240.244
R11613 gnd.n4078 gnd.n1275 240.244
R11614 gnd.n4078 gnd.n1276 240.244
R11615 gnd.n4069 gnd.n1276 240.244
R11616 gnd.n4070 gnd.n4069 240.244
R11617 gnd.n4070 gnd.n251 240.244
R11618 gnd.n6642 gnd.n251 240.244
R11619 gnd.n6642 gnd.n252 240.244
R11620 gnd.n6638 gnd.n252 240.244
R11621 gnd.n6638 gnd.n6637 240.244
R11622 gnd.n6062 gnd.n596 240.244
R11623 gnd.n6062 gnd.n598 240.244
R11624 gnd.n6058 gnd.n598 240.244
R11625 gnd.n6058 gnd.n604 240.244
R11626 gnd.n6054 gnd.n604 240.244
R11627 gnd.n6054 gnd.n606 240.244
R11628 gnd.n6050 gnd.n606 240.244
R11629 gnd.n6050 gnd.n612 240.244
R11630 gnd.n6046 gnd.n612 240.244
R11631 gnd.n6046 gnd.n614 240.244
R11632 gnd.n6042 gnd.n614 240.244
R11633 gnd.n6042 gnd.n620 240.244
R11634 gnd.n6038 gnd.n620 240.244
R11635 gnd.n6038 gnd.n622 240.244
R11636 gnd.n6034 gnd.n622 240.244
R11637 gnd.n6034 gnd.n628 240.244
R11638 gnd.n6030 gnd.n628 240.244
R11639 gnd.n6030 gnd.n630 240.244
R11640 gnd.n6026 gnd.n630 240.244
R11641 gnd.n6026 gnd.n636 240.244
R11642 gnd.n6022 gnd.n636 240.244
R11643 gnd.n6022 gnd.n638 240.244
R11644 gnd.n6018 gnd.n638 240.244
R11645 gnd.n6018 gnd.n644 240.244
R11646 gnd.n6014 gnd.n644 240.244
R11647 gnd.n6014 gnd.n646 240.244
R11648 gnd.n6010 gnd.n646 240.244
R11649 gnd.n6010 gnd.n652 240.244
R11650 gnd.n6006 gnd.n652 240.244
R11651 gnd.n6006 gnd.n654 240.244
R11652 gnd.n6002 gnd.n654 240.244
R11653 gnd.n6002 gnd.n660 240.244
R11654 gnd.n5998 gnd.n660 240.244
R11655 gnd.n5998 gnd.n662 240.244
R11656 gnd.n5994 gnd.n662 240.244
R11657 gnd.n5994 gnd.n668 240.244
R11658 gnd.n5990 gnd.n668 240.244
R11659 gnd.n5990 gnd.n670 240.244
R11660 gnd.n5986 gnd.n670 240.244
R11661 gnd.n5986 gnd.n676 240.244
R11662 gnd.n5982 gnd.n676 240.244
R11663 gnd.n5982 gnd.n678 240.244
R11664 gnd.n5978 gnd.n678 240.244
R11665 gnd.n5978 gnd.n684 240.244
R11666 gnd.n5974 gnd.n684 240.244
R11667 gnd.n5974 gnd.n686 240.244
R11668 gnd.n5970 gnd.n686 240.244
R11669 gnd.n5970 gnd.n692 240.244
R11670 gnd.n5966 gnd.n692 240.244
R11671 gnd.n5966 gnd.n694 240.244
R11672 gnd.n5962 gnd.n694 240.244
R11673 gnd.n5962 gnd.n700 240.244
R11674 gnd.n5958 gnd.n700 240.244
R11675 gnd.n5958 gnd.n702 240.244
R11676 gnd.n5954 gnd.n702 240.244
R11677 gnd.n5954 gnd.n708 240.244
R11678 gnd.n5950 gnd.n708 240.244
R11679 gnd.n5950 gnd.n710 240.244
R11680 gnd.n5946 gnd.n710 240.244
R11681 gnd.n5946 gnd.n716 240.244
R11682 gnd.n5942 gnd.n716 240.244
R11683 gnd.n5942 gnd.n718 240.244
R11684 gnd.n5938 gnd.n718 240.244
R11685 gnd.n5938 gnd.n724 240.244
R11686 gnd.n5934 gnd.n724 240.244
R11687 gnd.n5934 gnd.n726 240.244
R11688 gnd.n5930 gnd.n726 240.244
R11689 gnd.n5930 gnd.n732 240.244
R11690 gnd.n5926 gnd.n732 240.244
R11691 gnd.n5926 gnd.n734 240.244
R11692 gnd.n5922 gnd.n734 240.244
R11693 gnd.n5922 gnd.n740 240.244
R11694 gnd.n5918 gnd.n740 240.244
R11695 gnd.n5918 gnd.n742 240.244
R11696 gnd.n5914 gnd.n742 240.244
R11697 gnd.n5914 gnd.n748 240.244
R11698 gnd.n5910 gnd.n748 240.244
R11699 gnd.n5910 gnd.n750 240.244
R11700 gnd.n5906 gnd.n750 240.244
R11701 gnd.n5906 gnd.n756 240.244
R11702 gnd.n5902 gnd.n756 240.244
R11703 gnd.n5902 gnd.n758 240.244
R11704 gnd.n5898 gnd.n758 240.244
R11705 gnd.n5898 gnd.n764 240.244
R11706 gnd.n1089 gnd.n1088 240.244
R11707 gnd.n1090 gnd.n1089 240.244
R11708 gnd.n2600 gnd.n1090 240.244
R11709 gnd.n2600 gnd.n1093 240.244
R11710 gnd.n1094 gnd.n1093 240.244
R11711 gnd.n1095 gnd.n1094 240.244
R11712 gnd.n1815 gnd.n1095 240.244
R11713 gnd.n1815 gnd.n1098 240.244
R11714 gnd.n1099 gnd.n1098 240.244
R11715 gnd.n1100 gnd.n1099 240.244
R11716 gnd.n2789 gnd.n1100 240.244
R11717 gnd.n2789 gnd.n1103 240.244
R11718 gnd.n1104 gnd.n1103 240.244
R11719 gnd.n1105 gnd.n1104 240.244
R11720 gnd.n1759 gnd.n1105 240.244
R11721 gnd.n1759 gnd.n1108 240.244
R11722 gnd.n1109 gnd.n1108 240.244
R11723 gnd.n1110 gnd.n1109 240.244
R11724 gnd.n1728 gnd.n1110 240.244
R11725 gnd.n1728 gnd.n1113 240.244
R11726 gnd.n1114 gnd.n1113 240.244
R11727 gnd.n1115 gnd.n1114 240.244
R11728 gnd.n2924 gnd.n1115 240.244
R11729 gnd.n2924 gnd.n1118 240.244
R11730 gnd.n1119 gnd.n1118 240.244
R11731 gnd.n1120 gnd.n1119 240.244
R11732 gnd.n2904 gnd.n1120 240.244
R11733 gnd.n2904 gnd.n1123 240.244
R11734 gnd.n1124 gnd.n1123 240.244
R11735 gnd.n1125 gnd.n1124 240.244
R11736 gnd.n2994 gnd.n1125 240.244
R11737 gnd.n2994 gnd.n1128 240.244
R11738 gnd.n1129 gnd.n1128 240.244
R11739 gnd.n1130 gnd.n1129 240.244
R11740 gnd.n3006 gnd.n1130 240.244
R11741 gnd.n3006 gnd.n1133 240.244
R11742 gnd.n1134 gnd.n1133 240.244
R11743 gnd.n1135 gnd.n1134 240.244
R11744 gnd.n3045 gnd.n1135 240.244
R11745 gnd.n3045 gnd.n1138 240.244
R11746 gnd.n1139 gnd.n1138 240.244
R11747 gnd.n1140 gnd.n1139 240.244
R11748 gnd.n3086 gnd.n1140 240.244
R11749 gnd.n3086 gnd.n1143 240.244
R11750 gnd.n1144 gnd.n1143 240.244
R11751 gnd.n1145 gnd.n1144 240.244
R11752 gnd.n3156 gnd.n1145 240.244
R11753 gnd.n3156 gnd.n1148 240.244
R11754 gnd.n1149 gnd.n1148 240.244
R11755 gnd.n1150 gnd.n1149 240.244
R11756 gnd.n3215 gnd.n1150 240.244
R11757 gnd.n3215 gnd.n1153 240.244
R11758 gnd.n1154 gnd.n1153 240.244
R11759 gnd.n1155 gnd.n1154 240.244
R11760 gnd.n3246 gnd.n1155 240.244
R11761 gnd.n3246 gnd.n1158 240.244
R11762 gnd.n1159 gnd.n1158 240.244
R11763 gnd.n1160 gnd.n1159 240.244
R11764 gnd.n3286 gnd.n1160 240.244
R11765 gnd.n3286 gnd.n1163 240.244
R11766 gnd.n1164 gnd.n1163 240.244
R11767 gnd.n1165 gnd.n1164 240.244
R11768 gnd.n3313 gnd.n1165 240.244
R11769 gnd.n3313 gnd.n1168 240.244
R11770 gnd.n1169 gnd.n1168 240.244
R11771 gnd.n1170 gnd.n1169 240.244
R11772 gnd.n1478 gnd.n1170 240.244
R11773 gnd.n1478 gnd.n1173 240.244
R11774 gnd.n1174 gnd.n1173 240.244
R11775 gnd.n1175 gnd.n1174 240.244
R11776 gnd.n3389 gnd.n1175 240.244
R11777 gnd.n3389 gnd.n1178 240.244
R11778 gnd.n1179 gnd.n1178 240.244
R11779 gnd.n1180 gnd.n1179 240.244
R11780 gnd.n1419 gnd.n1180 240.244
R11781 gnd.n1419 gnd.n1183 240.244
R11782 gnd.n1184 gnd.n1183 240.244
R11783 gnd.n1185 gnd.n1184 240.244
R11784 gnd.n1436 gnd.n1185 240.244
R11785 gnd.n1436 gnd.n1188 240.244
R11786 gnd.n1189 gnd.n1188 240.244
R11787 gnd.n4147 gnd.n1189 240.244
R11788 gnd.n2090 gnd.n2089 240.244
R11789 gnd.n2105 gnd.n2089 240.244
R11790 gnd.n2107 gnd.n2106 240.244
R11791 gnd.n2117 gnd.n2116 240.244
R11792 gnd.n2128 gnd.n2127 240.244
R11793 gnd.n2130 gnd.n2129 240.244
R11794 gnd.n2140 gnd.n2139 240.244
R11795 gnd.n2153 gnd.n2152 240.244
R11796 gnd.n2155 gnd.n2154 240.244
R11797 gnd.n2038 gnd.n2037 240.244
R11798 gnd.n2083 gnd.n2039 240.244
R11799 gnd.n2043 gnd.n2042 240.244
R11800 gnd.n2049 gnd.n2044 240.244
R11801 gnd.n2051 gnd.n2050 240.244
R11802 gnd.n2055 gnd.n2054 240.244
R11803 gnd.n2056 gnd.n2055 240.244
R11804 gnd.n2599 gnd.n2056 240.244
R11805 gnd.n2599 gnd.n2059 240.244
R11806 gnd.n2060 gnd.n2059 240.244
R11807 gnd.n2625 gnd.n2060 240.244
R11808 gnd.n2626 gnd.n2625 240.244
R11809 gnd.n2626 gnd.n1788 240.244
R11810 gnd.n2781 gnd.n1788 240.244
R11811 gnd.n2781 gnd.n1783 240.244
R11812 gnd.n2788 gnd.n1783 240.244
R11813 gnd.n2788 gnd.n1767 240.244
R11814 gnd.n2811 gnd.n1767 240.244
R11815 gnd.n2812 gnd.n2811 240.244
R11816 gnd.n2812 gnd.n1761 240.244
R11817 gnd.n2825 gnd.n1761 240.244
R11818 gnd.n2825 gnd.n1762 240.244
R11819 gnd.n2817 gnd.n1762 240.244
R11820 gnd.n2818 gnd.n2817 240.244
R11821 gnd.n2818 gnd.n1719 240.244
R11822 gnd.n2897 gnd.n1719 240.244
R11823 gnd.n2897 gnd.n1714 240.244
R11824 gnd.n2923 gnd.n1714 240.244
R11825 gnd.n2923 gnd.n1710 240.244
R11826 gnd.n1710 gnd.n1702 240.244
R11827 gnd.n2902 gnd.n1702 240.244
R11828 gnd.n2906 gnd.n2902 240.244
R11829 gnd.n2907 gnd.n2906 240.244
R11830 gnd.n2907 gnd.n1685 240.244
R11831 gnd.n1685 gnd.n1667 240.244
R11832 gnd.n2996 gnd.n1667 240.244
R11833 gnd.n2997 gnd.n2996 240.244
R11834 gnd.n2999 gnd.n2997 240.244
R11835 gnd.n2999 gnd.n1663 240.244
R11836 gnd.n3005 gnd.n1663 240.244
R11837 gnd.n3005 gnd.n1637 240.244
R11838 gnd.n3053 gnd.n1637 240.244
R11839 gnd.n3053 gnd.n1638 240.244
R11840 gnd.n3047 gnd.n1638 240.244
R11841 gnd.n3047 gnd.n1615 240.244
R11842 gnd.n3111 gnd.n1615 240.244
R11843 gnd.n3111 gnd.n1607 240.244
R11844 gnd.n3088 gnd.n1607 240.244
R11845 gnd.n3089 gnd.n3088 240.244
R11846 gnd.n3090 gnd.n3089 240.244
R11847 gnd.n3090 gnd.n1588 240.244
R11848 gnd.n1588 gnd.n1581 240.244
R11849 gnd.n3093 gnd.n1581 240.244
R11850 gnd.n3096 gnd.n3093 240.244
R11851 gnd.n3096 gnd.n1559 240.244
R11852 gnd.n3217 gnd.n1559 240.244
R11853 gnd.n3217 gnd.n1553 240.244
R11854 gnd.n3224 gnd.n1553 240.244
R11855 gnd.n3224 gnd.n1554 240.244
R11856 gnd.n1554 gnd.n1530 240.244
R11857 gnd.n3256 gnd.n1530 240.244
R11858 gnd.n3256 gnd.n1525 240.244
R11859 gnd.n3277 gnd.n1525 240.244
R11860 gnd.n3277 gnd.n1518 240.244
R11861 gnd.n3261 gnd.n1518 240.244
R11862 gnd.n3262 gnd.n3261 240.244
R11863 gnd.n3264 gnd.n3262 240.244
R11864 gnd.n3264 gnd.n1499 240.244
R11865 gnd.n1499 gnd.n1491 240.244
R11866 gnd.n1491 gnd.n1475 240.244
R11867 gnd.n3349 gnd.n1475 240.244
R11868 gnd.n3349 gnd.n1470 240.244
R11869 gnd.n3356 gnd.n1470 240.244
R11870 gnd.n3356 gnd.n1460 240.244
R11871 gnd.n1460 gnd.n1448 240.244
R11872 gnd.n3391 gnd.n1448 240.244
R11873 gnd.n3391 gnd.n1409 240.244
R11874 gnd.n3398 gnd.n1409 240.244
R11875 gnd.n3400 gnd.n3398 240.244
R11876 gnd.n3401 gnd.n3400 240.244
R11877 gnd.n3401 gnd.n1421 240.244
R11878 gnd.n1422 gnd.n1421 240.244
R11879 gnd.n3408 gnd.n1422 240.244
R11880 gnd.n3409 gnd.n3408 240.244
R11881 gnd.n3409 gnd.n1438 240.244
R11882 gnd.n3591 gnd.n1438 240.244
R11883 gnd.n3591 gnd.n1193 240.244
R11884 gnd.n3482 gnd.n3481 240.244
R11885 gnd.n3485 gnd.n3484 240.244
R11886 gnd.n3501 gnd.n3500 240.244
R11887 gnd.n3504 gnd.n3503 240.244
R11888 gnd.n3520 gnd.n3519 240.244
R11889 gnd.n3523 gnd.n3522 240.244
R11890 gnd.n3539 gnd.n3538 240.244
R11891 gnd.n3543 gnd.n3541 240.244
R11892 gnd.n3559 gnd.n3423 240.244
R11893 gnd.n3563 gnd.n3561 240.244
R11894 gnd.n3569 gnd.n3419 240.244
R11895 gnd.n3573 gnd.n3571 240.244
R11896 gnd.n3582 gnd.n3415 240.244
R11897 gnd.n3585 gnd.n3584 240.244
R11898 gnd.n1799 gnd.n1798 240.132
R11899 gnd.n3629 gnd.n3628 240.132
R11900 gnd.n6065 gnd.n592 225.874
R11901 gnd.n6073 gnd.n592 225.874
R11902 gnd.n6074 gnd.n6073 225.874
R11903 gnd.n6075 gnd.n6074 225.874
R11904 gnd.n6075 gnd.n586 225.874
R11905 gnd.n6083 gnd.n586 225.874
R11906 gnd.n6084 gnd.n6083 225.874
R11907 gnd.n6085 gnd.n6084 225.874
R11908 gnd.n6085 gnd.n580 225.874
R11909 gnd.n6093 gnd.n580 225.874
R11910 gnd.n6094 gnd.n6093 225.874
R11911 gnd.n6095 gnd.n6094 225.874
R11912 gnd.n6095 gnd.n574 225.874
R11913 gnd.n6103 gnd.n574 225.874
R11914 gnd.n6104 gnd.n6103 225.874
R11915 gnd.n6105 gnd.n6104 225.874
R11916 gnd.n6105 gnd.n568 225.874
R11917 gnd.n6113 gnd.n568 225.874
R11918 gnd.n6114 gnd.n6113 225.874
R11919 gnd.n6115 gnd.n6114 225.874
R11920 gnd.n6115 gnd.n562 225.874
R11921 gnd.n6123 gnd.n562 225.874
R11922 gnd.n6124 gnd.n6123 225.874
R11923 gnd.n6125 gnd.n6124 225.874
R11924 gnd.n6125 gnd.n556 225.874
R11925 gnd.n6133 gnd.n556 225.874
R11926 gnd.n6134 gnd.n6133 225.874
R11927 gnd.n6135 gnd.n6134 225.874
R11928 gnd.n6135 gnd.n550 225.874
R11929 gnd.n6143 gnd.n550 225.874
R11930 gnd.n6144 gnd.n6143 225.874
R11931 gnd.n6145 gnd.n6144 225.874
R11932 gnd.n6145 gnd.n544 225.874
R11933 gnd.n6153 gnd.n544 225.874
R11934 gnd.n6154 gnd.n6153 225.874
R11935 gnd.n6155 gnd.n6154 225.874
R11936 gnd.n6155 gnd.n538 225.874
R11937 gnd.n6163 gnd.n538 225.874
R11938 gnd.n6164 gnd.n6163 225.874
R11939 gnd.n6165 gnd.n6164 225.874
R11940 gnd.n6165 gnd.n532 225.874
R11941 gnd.n6173 gnd.n532 225.874
R11942 gnd.n6174 gnd.n6173 225.874
R11943 gnd.n6175 gnd.n6174 225.874
R11944 gnd.n6175 gnd.n526 225.874
R11945 gnd.n6183 gnd.n526 225.874
R11946 gnd.n6184 gnd.n6183 225.874
R11947 gnd.n6185 gnd.n6184 225.874
R11948 gnd.n6185 gnd.n520 225.874
R11949 gnd.n6193 gnd.n520 225.874
R11950 gnd.n6194 gnd.n6193 225.874
R11951 gnd.n6195 gnd.n6194 225.874
R11952 gnd.n6195 gnd.n514 225.874
R11953 gnd.n6203 gnd.n514 225.874
R11954 gnd.n6204 gnd.n6203 225.874
R11955 gnd.n6205 gnd.n6204 225.874
R11956 gnd.n6205 gnd.n508 225.874
R11957 gnd.n6213 gnd.n508 225.874
R11958 gnd.n6214 gnd.n6213 225.874
R11959 gnd.n6215 gnd.n6214 225.874
R11960 gnd.n6215 gnd.n502 225.874
R11961 gnd.n6223 gnd.n502 225.874
R11962 gnd.n6224 gnd.n6223 225.874
R11963 gnd.n6225 gnd.n6224 225.874
R11964 gnd.n6225 gnd.n496 225.874
R11965 gnd.n6233 gnd.n496 225.874
R11966 gnd.n6234 gnd.n6233 225.874
R11967 gnd.n6235 gnd.n6234 225.874
R11968 gnd.n6235 gnd.n490 225.874
R11969 gnd.n6243 gnd.n490 225.874
R11970 gnd.n6244 gnd.n6243 225.874
R11971 gnd.n6245 gnd.n6244 225.874
R11972 gnd.n6245 gnd.n484 225.874
R11973 gnd.n6253 gnd.n484 225.874
R11974 gnd.n6254 gnd.n6253 225.874
R11975 gnd.n6255 gnd.n6254 225.874
R11976 gnd.n6255 gnd.n478 225.874
R11977 gnd.n6263 gnd.n478 225.874
R11978 gnd.n6264 gnd.n6263 225.874
R11979 gnd.n6265 gnd.n6264 225.874
R11980 gnd.n6265 gnd.n472 225.874
R11981 gnd.n6273 gnd.n472 225.874
R11982 gnd.n6274 gnd.n6273 225.874
R11983 gnd.n6275 gnd.n6274 225.874
R11984 gnd.n6275 gnd.n466 225.874
R11985 gnd.n6283 gnd.n466 225.874
R11986 gnd.n6284 gnd.n6283 225.874
R11987 gnd.n6285 gnd.n6284 225.874
R11988 gnd.n6285 gnd.n460 225.874
R11989 gnd.n6293 gnd.n460 225.874
R11990 gnd.n6294 gnd.n6293 225.874
R11991 gnd.n6295 gnd.n6294 225.874
R11992 gnd.n6295 gnd.n454 225.874
R11993 gnd.n6303 gnd.n454 225.874
R11994 gnd.n6304 gnd.n6303 225.874
R11995 gnd.n6305 gnd.n6304 225.874
R11996 gnd.n6305 gnd.n448 225.874
R11997 gnd.n6313 gnd.n448 225.874
R11998 gnd.n6314 gnd.n6313 225.874
R11999 gnd.n6315 gnd.n6314 225.874
R12000 gnd.n6315 gnd.n442 225.874
R12001 gnd.n6323 gnd.n442 225.874
R12002 gnd.n6324 gnd.n6323 225.874
R12003 gnd.n6325 gnd.n6324 225.874
R12004 gnd.n6325 gnd.n436 225.874
R12005 gnd.n6333 gnd.n436 225.874
R12006 gnd.n6334 gnd.n6333 225.874
R12007 gnd.n6335 gnd.n6334 225.874
R12008 gnd.n6335 gnd.n430 225.874
R12009 gnd.n6343 gnd.n430 225.874
R12010 gnd.n6344 gnd.n6343 225.874
R12011 gnd.n6345 gnd.n6344 225.874
R12012 gnd.n6345 gnd.n424 225.874
R12013 gnd.n6353 gnd.n424 225.874
R12014 gnd.n6354 gnd.n6353 225.874
R12015 gnd.n6355 gnd.n6354 225.874
R12016 gnd.n6355 gnd.n418 225.874
R12017 gnd.n6363 gnd.n418 225.874
R12018 gnd.n6364 gnd.n6363 225.874
R12019 gnd.n6365 gnd.n6364 225.874
R12020 gnd.n6365 gnd.n412 225.874
R12021 gnd.n6373 gnd.n412 225.874
R12022 gnd.n6374 gnd.n6373 225.874
R12023 gnd.n6375 gnd.n6374 225.874
R12024 gnd.n6375 gnd.n406 225.874
R12025 gnd.n6383 gnd.n406 225.874
R12026 gnd.n6384 gnd.n6383 225.874
R12027 gnd.n6385 gnd.n6384 225.874
R12028 gnd.n6385 gnd.n400 225.874
R12029 gnd.n6393 gnd.n400 225.874
R12030 gnd.n6394 gnd.n6393 225.874
R12031 gnd.n6395 gnd.n6394 225.874
R12032 gnd.n6395 gnd.n394 225.874
R12033 gnd.n6403 gnd.n394 225.874
R12034 gnd.n6404 gnd.n6403 225.874
R12035 gnd.n6405 gnd.n6404 225.874
R12036 gnd.n6405 gnd.n388 225.874
R12037 gnd.n6414 gnd.n388 225.874
R12038 gnd.n6415 gnd.n6414 225.874
R12039 gnd.n6416 gnd.n6415 225.874
R12040 gnd.n6416 gnd.n383 225.874
R12041 gnd.n4936 gnd.t215 224.174
R12042 gnd.n4557 gnd.t149 224.174
R12043 gnd.n3829 gnd.n3828 199.319
R12044 gnd.n3829 gnd.n3775 199.319
R12045 gnd.n1943 gnd.n1937 199.319
R12046 gnd.n1942 gnd.n1937 199.319
R12047 gnd.n1800 gnd.n1797 186.49
R12048 gnd.n3630 gnd.n3627 186.49
R12049 gnd.n5718 gnd.n5717 185
R12050 gnd.n5716 gnd.n5715 185
R12051 gnd.n5695 gnd.n5694 185
R12052 gnd.n5710 gnd.n5709 185
R12053 gnd.n5708 gnd.n5707 185
R12054 gnd.n5699 gnd.n5698 185
R12055 gnd.n5702 gnd.n5701 185
R12056 gnd.n5686 gnd.n5685 185
R12057 gnd.n5684 gnd.n5683 185
R12058 gnd.n5663 gnd.n5662 185
R12059 gnd.n5678 gnd.n5677 185
R12060 gnd.n5676 gnd.n5675 185
R12061 gnd.n5667 gnd.n5666 185
R12062 gnd.n5670 gnd.n5669 185
R12063 gnd.n5654 gnd.n5653 185
R12064 gnd.n5652 gnd.n5651 185
R12065 gnd.n5631 gnd.n5630 185
R12066 gnd.n5646 gnd.n5645 185
R12067 gnd.n5644 gnd.n5643 185
R12068 gnd.n5635 gnd.n5634 185
R12069 gnd.n5638 gnd.n5637 185
R12070 gnd.n5623 gnd.n5622 185
R12071 gnd.n5621 gnd.n5620 185
R12072 gnd.n5600 gnd.n5599 185
R12073 gnd.n5615 gnd.n5614 185
R12074 gnd.n5613 gnd.n5612 185
R12075 gnd.n5604 gnd.n5603 185
R12076 gnd.n5607 gnd.n5606 185
R12077 gnd.n5591 gnd.n5590 185
R12078 gnd.n5589 gnd.n5588 185
R12079 gnd.n5568 gnd.n5567 185
R12080 gnd.n5583 gnd.n5582 185
R12081 gnd.n5581 gnd.n5580 185
R12082 gnd.n5572 gnd.n5571 185
R12083 gnd.n5575 gnd.n5574 185
R12084 gnd.n5559 gnd.n5558 185
R12085 gnd.n5557 gnd.n5556 185
R12086 gnd.n5536 gnd.n5535 185
R12087 gnd.n5551 gnd.n5550 185
R12088 gnd.n5549 gnd.n5548 185
R12089 gnd.n5540 gnd.n5539 185
R12090 gnd.n5543 gnd.n5542 185
R12091 gnd.n5527 gnd.n5526 185
R12092 gnd.n5525 gnd.n5524 185
R12093 gnd.n5504 gnd.n5503 185
R12094 gnd.n5519 gnd.n5518 185
R12095 gnd.n5517 gnd.n5516 185
R12096 gnd.n5508 gnd.n5507 185
R12097 gnd.n5511 gnd.n5510 185
R12098 gnd.n5496 gnd.n5495 185
R12099 gnd.n5494 gnd.n5493 185
R12100 gnd.n5473 gnd.n5472 185
R12101 gnd.n5488 gnd.n5487 185
R12102 gnd.n5486 gnd.n5485 185
R12103 gnd.n5477 gnd.n5476 185
R12104 gnd.n5480 gnd.n5479 185
R12105 gnd.n4937 gnd.t214 178.987
R12106 gnd.n4558 gnd.t150 178.987
R12107 gnd.n1 gnd.t233 170.774
R12108 gnd.n7 gnd.t57 170.103
R12109 gnd.n6 gnd.t78 170.103
R12110 gnd.n5 gnd.t255 170.103
R12111 gnd.n4 gnd.t228 170.103
R12112 gnd.n3 gnd.t261 170.103
R12113 gnd.n2 gnd.t72 170.103
R12114 gnd.n1 gnd.t291 170.103
R12115 gnd.n3698 gnd.n3697 163.367
R12116 gnd.n3694 gnd.n3693 163.367
R12117 gnd.n3690 gnd.n3689 163.367
R12118 gnd.n3686 gnd.n3685 163.367
R12119 gnd.n3682 gnd.n3681 163.367
R12120 gnd.n3678 gnd.n3677 163.367
R12121 gnd.n3674 gnd.n3673 163.367
R12122 gnd.n3670 gnd.n3669 163.367
R12123 gnd.n3666 gnd.n3665 163.367
R12124 gnd.n3662 gnd.n3661 163.367
R12125 gnd.n3658 gnd.n3657 163.367
R12126 gnd.n3654 gnd.n3653 163.367
R12127 gnd.n3650 gnd.n3649 163.367
R12128 gnd.n3646 gnd.n3645 163.367
R12129 gnd.n3641 gnd.n3640 163.367
R12130 gnd.n3773 gnd.n1364 163.367
R12131 gnd.n3770 gnd.n3769 163.367
R12132 gnd.n3767 gnd.n1397 163.367
R12133 gnd.n3762 gnd.n3761 163.367
R12134 gnd.n3758 gnd.n3757 163.367
R12135 gnd.n3754 gnd.n3753 163.367
R12136 gnd.n3750 gnd.n3749 163.367
R12137 gnd.n3746 gnd.n3745 163.367
R12138 gnd.n3742 gnd.n3741 163.367
R12139 gnd.n3738 gnd.n3737 163.367
R12140 gnd.n3734 gnd.n3733 163.367
R12141 gnd.n3730 gnd.n3729 163.367
R12142 gnd.n3726 gnd.n3725 163.367
R12143 gnd.n3722 gnd.n3721 163.367
R12144 gnd.n3718 gnd.n3717 163.367
R12145 gnd.n3714 gnd.n3713 163.367
R12146 gnd.n3710 gnd.n3709 163.367
R12147 gnd.n1868 gnd.n1790 163.367
R12148 gnd.n1864 gnd.n1790 163.367
R12149 gnd.n1864 gnd.n1782 163.367
R12150 gnd.n1859 gnd.n1782 163.367
R12151 gnd.n1859 gnd.n1775 163.367
R12152 gnd.n1856 gnd.n1775 163.367
R12153 gnd.n1856 gnd.n1750 163.367
R12154 gnd.n2837 gnd.n1750 163.367
R12155 gnd.n2837 gnd.n1747 163.367
R12156 gnd.n2842 gnd.n1747 163.367
R12157 gnd.n2842 gnd.n1748 163.367
R12158 gnd.n1748 gnd.n1739 163.367
R12159 gnd.n2853 gnd.n1739 163.367
R12160 gnd.n2853 gnd.n1737 163.367
R12161 gnd.n2866 gnd.n1737 163.367
R12162 gnd.n2866 gnd.n1730 163.367
R12163 gnd.n2862 gnd.n1730 163.367
R12164 gnd.n2862 gnd.n2859 163.367
R12165 gnd.n2859 gnd.n2858 163.367
R12166 gnd.n2858 gnd.n1712 163.367
R12167 gnd.n2927 gnd.n1712 163.367
R12168 gnd.n2927 gnd.n1709 163.367
R12169 gnd.n2936 gnd.n1709 163.367
R12170 gnd.n2936 gnd.n1703 163.367
R12171 gnd.n2932 gnd.n1703 163.367
R12172 gnd.n2932 gnd.n1696 163.367
R12173 gnd.n1696 gnd.n1688 163.367
R12174 gnd.n2964 gnd.n1688 163.367
R12175 gnd.n2964 gnd.n1686 163.367
R12176 gnd.n2971 gnd.n1686 163.367
R12177 gnd.n2971 gnd.n1676 163.367
R12178 gnd.n1677 gnd.n1676 163.367
R12179 gnd.n1677 gnd.n1669 163.367
R12180 gnd.n1669 gnd.n1659 163.367
R12181 gnd.n3014 gnd.n1659 163.367
R12182 gnd.n3014 gnd.n1660 163.367
R12183 gnd.n1660 gnd.n1652 163.367
R12184 gnd.n3009 gnd.n1652 163.367
R12185 gnd.n3009 gnd.n1644 163.367
R12186 gnd.n3036 gnd.n1644 163.367
R12187 gnd.n3036 gnd.n1636 163.367
R12188 gnd.n3039 gnd.n1636 163.367
R12189 gnd.n3039 gnd.n1629 163.367
R12190 gnd.n3043 gnd.n1629 163.367
R12191 gnd.n3043 gnd.n1621 163.367
R12192 gnd.n3076 gnd.n1621 163.367
R12193 gnd.n3076 gnd.n1614 163.367
R12194 gnd.n3079 gnd.n1614 163.367
R12195 gnd.n3079 gnd.n1608 163.367
R12196 gnd.n3084 gnd.n1608 163.367
R12197 gnd.n3084 gnd.n1598 163.367
R12198 gnd.n1598 gnd.n1591 163.367
R12199 gnd.n3138 gnd.n1591 163.367
R12200 gnd.n3138 gnd.n1589 163.367
R12201 gnd.n3143 gnd.n1589 163.367
R12202 gnd.n3143 gnd.n1580 163.367
R12203 gnd.n1580 gnd.n1572 163.367
R12204 gnd.n3173 gnd.n1572 163.367
R12205 gnd.n3173 gnd.n1569 163.367
R12206 gnd.n3205 gnd.n1569 163.367
R12207 gnd.n3205 gnd.n1570 163.367
R12208 gnd.n3201 gnd.n1570 163.367
R12209 gnd.n3201 gnd.n3200 163.367
R12210 gnd.n3200 gnd.n1551 163.367
R12211 gnd.n1552 gnd.n1551 163.367
R12212 gnd.n1552 gnd.n1545 163.367
R12213 gnd.n3194 gnd.n1545 163.367
R12214 gnd.n3194 gnd.n1538 163.367
R12215 gnd.n3190 gnd.n1538 163.367
R12216 gnd.n3190 gnd.n1532 163.367
R12217 gnd.n3187 gnd.n1532 163.367
R12218 gnd.n3187 gnd.n1524 163.367
R12219 gnd.n3181 gnd.n1524 163.367
R12220 gnd.n3181 gnd.n1519 163.367
R12221 gnd.n3178 gnd.n1519 163.367
R12222 gnd.n3178 gnd.n1508 163.367
R12223 gnd.n1508 gnd.n1502 163.367
R12224 gnd.n3305 gnd.n1502 163.367
R12225 gnd.n3305 gnd.n1500 163.367
R12226 gnd.n3310 gnd.n1500 163.367
R12227 gnd.n3310 gnd.n1490 163.367
R12228 gnd.n1490 gnd.n1483 163.367
R12229 gnd.n3339 gnd.n1483 163.367
R12230 gnd.n3339 gnd.n1480 163.367
R12231 gnd.n3346 gnd.n1480 163.367
R12232 gnd.n3346 gnd.n1481 163.367
R12233 gnd.n1481 gnd.n1469 163.367
R12234 gnd.n1469 gnd.n1459 163.367
R12235 gnd.n1459 gnd.n1452 163.367
R12236 gnd.n3381 gnd.n1452 163.367
R12237 gnd.n3381 gnd.n1450 163.367
R12238 gnd.n3387 gnd.n1450 163.367
R12239 gnd.n3387 gnd.n1408 163.367
R12240 gnd.n1408 gnd.n1401 163.367
R12241 gnd.n3705 gnd.n1401 163.367
R12242 gnd.n2770 gnd.n1814 163.367
R12243 gnd.n2770 gnd.n1850 163.367
R12244 gnd.n2766 gnd.n2765 163.367
R12245 gnd.n2762 gnd.n2761 163.367
R12246 gnd.n2758 gnd.n2757 163.367
R12247 gnd.n2754 gnd.n2753 163.367
R12248 gnd.n2750 gnd.n2749 163.367
R12249 gnd.n2746 gnd.n2745 163.367
R12250 gnd.n2742 gnd.n2741 163.367
R12251 gnd.n2738 gnd.n2737 163.367
R12252 gnd.n2734 gnd.n2733 163.367
R12253 gnd.n2730 gnd.n2729 163.367
R12254 gnd.n2726 gnd.n2725 163.367
R12255 gnd.n2722 gnd.n2721 163.367
R12256 gnd.n2718 gnd.n2717 163.367
R12257 gnd.n2714 gnd.n2713 163.367
R12258 gnd.n2710 gnd.n2709 163.367
R12259 gnd.n1930 gnd.n1929 163.367
R12260 gnd.n1925 gnd.n1924 163.367
R12261 gnd.n1921 gnd.n1920 163.367
R12262 gnd.n1917 gnd.n1916 163.367
R12263 gnd.n1913 gnd.n1912 163.367
R12264 gnd.n1909 gnd.n1908 163.367
R12265 gnd.n1905 gnd.n1904 163.367
R12266 gnd.n1901 gnd.n1900 163.367
R12267 gnd.n1897 gnd.n1896 163.367
R12268 gnd.n1893 gnd.n1892 163.367
R12269 gnd.n1889 gnd.n1888 163.367
R12270 gnd.n1885 gnd.n1884 163.367
R12271 gnd.n1881 gnd.n1880 163.367
R12272 gnd.n1877 gnd.n1876 163.367
R12273 gnd.n1873 gnd.n1872 163.367
R12274 gnd.n2778 gnd.n1792 163.367
R12275 gnd.n2778 gnd.n1780 163.367
R12276 gnd.n2792 gnd.n1780 163.367
R12277 gnd.n2792 gnd.n1777 163.367
R12278 gnd.n2797 gnd.n1777 163.367
R12279 gnd.n2797 gnd.n1778 163.367
R12280 gnd.n1778 gnd.n1753 163.367
R12281 gnd.n2835 gnd.n1753 163.367
R12282 gnd.n2835 gnd.n1754 163.367
R12283 gnd.n1754 gnd.n1746 163.367
R12284 gnd.n2830 gnd.n1746 163.367
R12285 gnd.n2830 gnd.n1757 163.367
R12286 gnd.n1757 gnd.n1735 163.367
R12287 gnd.n2870 gnd.n1735 163.367
R12288 gnd.n2870 gnd.n1732 163.367
R12289 gnd.n2883 gnd.n1732 163.367
R12290 gnd.n2883 gnd.n1733 163.367
R12291 gnd.n2879 gnd.n1733 163.367
R12292 gnd.n2879 gnd.n2878 163.367
R12293 gnd.n2878 gnd.n2877 163.367
R12294 gnd.n2877 gnd.n1707 163.367
R12295 gnd.n2940 gnd.n1707 163.367
R12296 gnd.n2940 gnd.n1705 163.367
R12297 gnd.n2944 gnd.n1705 163.367
R12298 gnd.n2944 gnd.n1694 163.367
R12299 gnd.n2957 gnd.n1694 163.367
R12300 gnd.n2957 gnd.n1691 163.367
R12301 gnd.n2962 gnd.n1691 163.367
R12302 gnd.n2962 gnd.n1692 163.367
R12303 gnd.n1692 gnd.n1674 163.367
R12304 gnd.n2988 gnd.n1674 163.367
R12305 gnd.n2988 gnd.n1672 163.367
R12306 gnd.n2992 gnd.n1672 163.367
R12307 gnd.n2992 gnd.n1657 163.367
R12308 gnd.n3016 gnd.n1657 163.367
R12309 gnd.n3016 gnd.n1654 163.367
R12310 gnd.n3023 gnd.n1654 163.367
R12311 gnd.n3023 gnd.n1655 163.367
R12312 gnd.n3019 gnd.n1655 163.367
R12313 gnd.n3019 gnd.n1634 163.367
R12314 gnd.n3056 gnd.n1634 163.367
R12315 gnd.n3056 gnd.n1631 163.367
R12316 gnd.n3063 gnd.n1631 163.367
R12317 gnd.n3063 gnd.n1632 163.367
R12318 gnd.n3059 gnd.n1632 163.367
R12319 gnd.n3059 gnd.n1612 163.367
R12320 gnd.n3114 gnd.n1612 163.367
R12321 gnd.n3114 gnd.n1610 163.367
R12322 gnd.n3118 gnd.n1610 163.367
R12323 gnd.n3118 gnd.n1597 163.367
R12324 gnd.n3131 gnd.n1597 163.367
R12325 gnd.n3131 gnd.n1594 163.367
R12326 gnd.n3136 gnd.n1594 163.367
R12327 gnd.n3136 gnd.n1595 163.367
R12328 gnd.n1595 gnd.n1578 163.367
R12329 gnd.n3159 gnd.n1578 163.367
R12330 gnd.n3159 gnd.n1575 163.367
R12331 gnd.n3171 gnd.n1575 163.367
R12332 gnd.n3171 gnd.n1576 163.367
R12333 gnd.n1576 gnd.n1567 163.367
R12334 gnd.n3166 gnd.n1567 163.367
R12335 gnd.n3166 gnd.n3163 163.367
R12336 gnd.n3163 gnd.n1549 163.367
R12337 gnd.n3229 gnd.n1549 163.367
R12338 gnd.n3229 gnd.n1547 163.367
R12339 gnd.n3233 gnd.n1547 163.367
R12340 gnd.n3233 gnd.n1536 163.367
R12341 gnd.n3249 gnd.n1536 163.367
R12342 gnd.n3249 gnd.n1534 163.367
R12343 gnd.n3253 gnd.n1534 163.367
R12344 gnd.n3253 gnd.n1523 163.367
R12345 gnd.n3280 gnd.n1523 163.367
R12346 gnd.n3280 gnd.n1521 163.367
R12347 gnd.n3284 gnd.n1521 163.367
R12348 gnd.n3284 gnd.n1506 163.367
R12349 gnd.n3298 gnd.n1506 163.367
R12350 gnd.n3298 gnd.n1503 163.367
R12351 gnd.n3303 gnd.n1503 163.367
R12352 gnd.n3303 gnd.n1504 163.367
R12353 gnd.n1504 gnd.n1489 163.367
R12354 gnd.n3329 gnd.n1489 163.367
R12355 gnd.n3329 gnd.n1486 163.367
R12356 gnd.n3337 gnd.n1486 163.367
R12357 gnd.n3337 gnd.n1487 163.367
R12358 gnd.n1487 gnd.n1477 163.367
R12359 gnd.n3332 gnd.n1477 163.367
R12360 gnd.n3332 gnd.n1457 163.367
R12361 gnd.n3374 gnd.n1457 163.367
R12362 gnd.n3374 gnd.n1454 163.367
R12363 gnd.n3379 gnd.n1454 163.367
R12364 gnd.n3379 gnd.n1455 163.367
R12365 gnd.n1455 gnd.n1406 163.367
R12366 gnd.n3615 gnd.n1406 163.367
R12367 gnd.n3615 gnd.n1403 163.367
R12368 gnd.n3703 gnd.n1403 163.367
R12369 gnd.n3636 gnd.n3635 156.462
R12370 gnd.n5658 gnd.n5626 153.042
R12371 gnd.n5722 gnd.n5721 152.079
R12372 gnd.n5690 gnd.n5689 152.079
R12373 gnd.n5658 gnd.n5657 152.079
R12374 gnd.n1805 gnd.n1804 152
R12375 gnd.n1806 gnd.n1795 152
R12376 gnd.n1808 gnd.n1807 152
R12377 gnd.n1810 gnd.n1793 152
R12378 gnd.n1812 gnd.n1811 152
R12379 gnd.n3634 gnd.n3618 152
R12380 gnd.n3626 gnd.n3619 152
R12381 gnd.n3625 gnd.n3624 152
R12382 gnd.n3623 gnd.n3620 152
R12383 gnd.n3621 gnd.t130 150.546
R12384 gnd.t287 gnd.n5700 147.661
R12385 gnd.t253 gnd.n5668 147.661
R12386 gnd.t251 gnd.n5636 147.661
R12387 gnd.t108 gnd.n5605 147.661
R12388 gnd.t76 gnd.n5573 147.661
R12389 gnd.t13 gnd.n5541 147.661
R12390 gnd.t257 gnd.n5509 147.661
R12391 gnd.t5 gnd.n5478 147.661
R12392 gnd.n3772 gnd.n1363 143.351
R12393 gnd.n2708 gnd.n1831 143.351
R12394 gnd.n2708 gnd.n1832 143.351
R12395 gnd.n1802 gnd.t187 130.484
R12396 gnd.n6425 gnd.n6424 127.204
R12397 gnd.n6426 gnd.n6425 127.204
R12398 gnd.n6426 gnd.n377 127.204
R12399 gnd.n6434 gnd.n377 127.204
R12400 gnd.n6435 gnd.n6434 127.204
R12401 gnd.n6436 gnd.n6435 127.204
R12402 gnd.n6436 gnd.n371 127.204
R12403 gnd.n6444 gnd.n371 127.204
R12404 gnd.n6445 gnd.n6444 127.204
R12405 gnd.n6446 gnd.n6445 127.204
R12406 gnd.n6446 gnd.n365 127.204
R12407 gnd.n6454 gnd.n365 127.204
R12408 gnd.n6455 gnd.n6454 127.204
R12409 gnd.n6456 gnd.n6455 127.204
R12410 gnd.n6456 gnd.n359 127.204
R12411 gnd.n6464 gnd.n359 127.204
R12412 gnd.n6465 gnd.n6464 127.204
R12413 gnd.n6466 gnd.n6465 127.204
R12414 gnd.n6466 gnd.n353 127.204
R12415 gnd.n6474 gnd.n353 127.204
R12416 gnd.n6475 gnd.n6474 127.204
R12417 gnd.n6476 gnd.n6475 127.204
R12418 gnd.n6476 gnd.n347 127.204
R12419 gnd.n6484 gnd.n347 127.204
R12420 gnd.n6485 gnd.n6484 127.204
R12421 gnd.n6486 gnd.n6485 127.204
R12422 gnd.n6486 gnd.n341 127.204
R12423 gnd.n6494 gnd.n341 127.204
R12424 gnd.n6495 gnd.n6494 127.204
R12425 gnd.n6496 gnd.n6495 127.204
R12426 gnd.n6496 gnd.n335 127.204
R12427 gnd.n6504 gnd.n335 127.204
R12428 gnd.n6505 gnd.n6504 127.204
R12429 gnd.n6506 gnd.n6505 127.204
R12430 gnd.n6506 gnd.n329 127.204
R12431 gnd.n6514 gnd.n329 127.204
R12432 gnd.n6515 gnd.n6514 127.204
R12433 gnd.n6516 gnd.n6515 127.204
R12434 gnd.n6516 gnd.n323 127.204
R12435 gnd.n6524 gnd.n323 127.204
R12436 gnd.n6525 gnd.n6524 127.204
R12437 gnd.n6526 gnd.n6525 127.204
R12438 gnd.n6526 gnd.n317 127.204
R12439 gnd.n6534 gnd.n317 127.204
R12440 gnd.n6535 gnd.n6534 127.204
R12441 gnd.n6536 gnd.n6535 127.204
R12442 gnd.n6536 gnd.n311 127.204
R12443 gnd.n6544 gnd.n311 127.204
R12444 gnd.n6545 gnd.n6544 127.204
R12445 gnd.n6546 gnd.n6545 127.204
R12446 gnd.n6546 gnd.n305 127.204
R12447 gnd.n6554 gnd.n305 127.204
R12448 gnd.n6555 gnd.n6554 127.204
R12449 gnd.n6556 gnd.n6555 127.204
R12450 gnd.n6556 gnd.n299 127.204
R12451 gnd.n6564 gnd.n299 127.204
R12452 gnd.n6565 gnd.n6564 127.204
R12453 gnd.n6566 gnd.n6565 127.204
R12454 gnd.n6566 gnd.n293 127.204
R12455 gnd.n6574 gnd.n293 127.204
R12456 gnd.n6575 gnd.n6574 127.204
R12457 gnd.n6576 gnd.n6575 127.204
R12458 gnd.n6576 gnd.n287 127.204
R12459 gnd.n6584 gnd.n287 127.204
R12460 gnd.n6585 gnd.n6584 127.204
R12461 gnd.n6586 gnd.n6585 127.204
R12462 gnd.n6586 gnd.n281 127.204
R12463 gnd.n6594 gnd.n281 127.204
R12464 gnd.n6595 gnd.n6594 127.204
R12465 gnd.n6596 gnd.n6595 127.204
R12466 gnd.n6596 gnd.n275 127.204
R12467 gnd.n6604 gnd.n275 127.204
R12468 gnd.n6605 gnd.n6604 127.204
R12469 gnd.n6606 gnd.n6605 127.204
R12470 gnd.n6606 gnd.n269 127.204
R12471 gnd.n6614 gnd.n269 127.204
R12472 gnd.n6615 gnd.n6614 127.204
R12473 gnd.n6616 gnd.n6615 127.204
R12474 gnd.n6616 gnd.n263 127.204
R12475 gnd.n6624 gnd.n263 127.204
R12476 gnd.n6625 gnd.n6624 127.204
R12477 gnd.n6627 gnd.n6625 127.204
R12478 gnd.n6627 gnd.n6626 127.204
R12479 gnd.n1811 gnd.t200 126.766
R12480 gnd.n1809 gnd.t144 126.766
R12481 gnd.n1795 gnd.t194 126.766
R12482 gnd.n1803 gnd.t170 126.766
R12483 gnd.n3622 gnd.t115 126.766
R12484 gnd.n3624 gnd.t206 126.766
R12485 gnd.n3633 gnd.t180 126.766
R12486 gnd.n3635 gnd.t161 126.766
R12487 gnd.n5717 gnd.n5716 104.615
R12488 gnd.n5716 gnd.n5694 104.615
R12489 gnd.n5709 gnd.n5694 104.615
R12490 gnd.n5709 gnd.n5708 104.615
R12491 gnd.n5708 gnd.n5698 104.615
R12492 gnd.n5701 gnd.n5698 104.615
R12493 gnd.n5685 gnd.n5684 104.615
R12494 gnd.n5684 gnd.n5662 104.615
R12495 gnd.n5677 gnd.n5662 104.615
R12496 gnd.n5677 gnd.n5676 104.615
R12497 gnd.n5676 gnd.n5666 104.615
R12498 gnd.n5669 gnd.n5666 104.615
R12499 gnd.n5653 gnd.n5652 104.615
R12500 gnd.n5652 gnd.n5630 104.615
R12501 gnd.n5645 gnd.n5630 104.615
R12502 gnd.n5645 gnd.n5644 104.615
R12503 gnd.n5644 gnd.n5634 104.615
R12504 gnd.n5637 gnd.n5634 104.615
R12505 gnd.n5622 gnd.n5621 104.615
R12506 gnd.n5621 gnd.n5599 104.615
R12507 gnd.n5614 gnd.n5599 104.615
R12508 gnd.n5614 gnd.n5613 104.615
R12509 gnd.n5613 gnd.n5603 104.615
R12510 gnd.n5606 gnd.n5603 104.615
R12511 gnd.n5590 gnd.n5589 104.615
R12512 gnd.n5589 gnd.n5567 104.615
R12513 gnd.n5582 gnd.n5567 104.615
R12514 gnd.n5582 gnd.n5581 104.615
R12515 gnd.n5581 gnd.n5571 104.615
R12516 gnd.n5574 gnd.n5571 104.615
R12517 gnd.n5558 gnd.n5557 104.615
R12518 gnd.n5557 gnd.n5535 104.615
R12519 gnd.n5550 gnd.n5535 104.615
R12520 gnd.n5550 gnd.n5549 104.615
R12521 gnd.n5549 gnd.n5539 104.615
R12522 gnd.n5542 gnd.n5539 104.615
R12523 gnd.n5526 gnd.n5525 104.615
R12524 gnd.n5525 gnd.n5503 104.615
R12525 gnd.n5518 gnd.n5503 104.615
R12526 gnd.n5518 gnd.n5517 104.615
R12527 gnd.n5517 gnd.n5507 104.615
R12528 gnd.n5510 gnd.n5507 104.615
R12529 gnd.n5495 gnd.n5494 104.615
R12530 gnd.n5494 gnd.n5472 104.615
R12531 gnd.n5487 gnd.n5472 104.615
R12532 gnd.n5487 gnd.n5486 104.615
R12533 gnd.n5486 gnd.n5476 104.615
R12534 gnd.n5479 gnd.n5476 104.615
R12535 gnd.n4862 gnd.t114 100.632
R12536 gnd.n4513 gnd.t142 100.632
R12537 gnd.n6873 gnd.n93 99.6594
R12538 gnd.n6871 gnd.n6870 99.6594
R12539 gnd.n6866 gnd.n100 99.6594
R12540 gnd.n6864 gnd.n6863 99.6594
R12541 gnd.n6859 gnd.n107 99.6594
R12542 gnd.n6857 gnd.n6856 99.6594
R12543 gnd.n6852 gnd.n114 99.6594
R12544 gnd.n6850 gnd.n6849 99.6594
R12545 gnd.n6842 gnd.n121 99.6594
R12546 gnd.n6840 gnd.n6839 99.6594
R12547 gnd.n6835 gnd.n128 99.6594
R12548 gnd.n6833 gnd.n6832 99.6594
R12549 gnd.n6828 gnd.n135 99.6594
R12550 gnd.n6826 gnd.n6825 99.6594
R12551 gnd.n6821 gnd.n142 99.6594
R12552 gnd.n6819 gnd.n6818 99.6594
R12553 gnd.n6814 gnd.n149 99.6594
R12554 gnd.n6812 gnd.n6811 99.6594
R12555 gnd.n154 gnd.n153 99.6594
R12556 gnd.n3793 gnd.n1217 99.6594
R12557 gnd.n3797 gnd.n3796 99.6594
R12558 gnd.n3804 gnd.n3803 99.6594
R12559 gnd.n3807 gnd.n3806 99.6594
R12560 gnd.n3814 gnd.n3813 99.6594
R12561 gnd.n3817 gnd.n3816 99.6594
R12562 gnd.n3825 gnd.n3824 99.6594
R12563 gnd.n3828 gnd.n3827 99.6594
R12564 gnd.n3838 gnd.n3837 99.6594
R12565 gnd.n3841 gnd.n3840 99.6594
R12566 gnd.n3848 gnd.n3847 99.6594
R12567 gnd.n3851 gnd.n3850 99.6594
R12568 gnd.n3858 gnd.n3857 99.6594
R12569 gnd.n3861 gnd.n3860 99.6594
R12570 gnd.n3868 gnd.n3867 99.6594
R12571 gnd.n3871 gnd.n3870 99.6594
R12572 gnd.n3879 gnd.n3878 99.6594
R12573 gnd.n3882 gnd.n3881 99.6594
R12574 gnd.n1995 gnd.n1994 99.6594
R12575 gnd.n1990 gnd.n1949 99.6594
R12576 gnd.n1986 gnd.n1948 99.6594
R12577 gnd.n1982 gnd.n1947 99.6594
R12578 gnd.n1978 gnd.n1946 99.6594
R12579 gnd.n1974 gnd.n1945 99.6594
R12580 gnd.n1970 gnd.n1944 99.6594
R12581 gnd.n1942 gnd.n1941 99.6594
R12582 gnd.n2701 gnd.n2700 99.6594
R12583 gnd.n2698 gnd.n2697 99.6594
R12584 gnd.n2693 gnd.n2004 99.6594
R12585 gnd.n2691 gnd.n2690 99.6594
R12586 gnd.n2686 gnd.n2011 99.6594
R12587 gnd.n2684 gnd.n2683 99.6594
R12588 gnd.n2679 gnd.n2018 99.6594
R12589 gnd.n2677 gnd.n2676 99.6594
R12590 gnd.n2672 gnd.n2027 99.6594
R12591 gnd.n2670 gnd.n2669 99.6594
R12592 gnd.n4481 gnd.n4480 99.6594
R12593 gnd.n4475 gnd.n802 99.6594
R12594 gnd.n4472 gnd.n803 99.6594
R12595 gnd.n4468 gnd.n804 99.6594
R12596 gnd.n4464 gnd.n805 99.6594
R12597 gnd.n4460 gnd.n806 99.6594
R12598 gnd.n4456 gnd.n807 99.6594
R12599 gnd.n4452 gnd.n808 99.6594
R12600 gnd.n4448 gnd.n809 99.6594
R12601 gnd.n4443 gnd.n810 99.6594
R12602 gnd.n4439 gnd.n811 99.6594
R12603 gnd.n4435 gnd.n812 99.6594
R12604 gnd.n4431 gnd.n813 99.6594
R12605 gnd.n4427 gnd.n814 99.6594
R12606 gnd.n4423 gnd.n815 99.6594
R12607 gnd.n4419 gnd.n816 99.6594
R12608 gnd.n4415 gnd.n817 99.6594
R12609 gnd.n4411 gnd.n818 99.6594
R12610 gnd.n873 gnd.n819 99.6594
R12611 gnd.n5866 gnd.n4493 99.6594
R12612 gnd.n5864 gnd.n5863 99.6594
R12613 gnd.n5859 gnd.n4500 99.6594
R12614 gnd.n5857 gnd.n5856 99.6594
R12615 gnd.n5852 gnd.n4507 99.6594
R12616 gnd.n5850 gnd.n5849 99.6594
R12617 gnd.n5845 gnd.n4516 99.6594
R12618 gnd.n5843 gnd.n5842 99.6594
R12619 gnd.n5148 gnd.n4805 99.6594
R12620 gnd.n4831 gnd.n4812 99.6594
R12621 gnd.n4833 gnd.n4813 99.6594
R12622 gnd.n4841 gnd.n4814 99.6594
R12623 gnd.n4843 gnd.n4815 99.6594
R12624 gnd.n4851 gnd.n4816 99.6594
R12625 gnd.n4853 gnd.n4817 99.6594
R12626 gnd.n4861 gnd.n4818 99.6594
R12627 gnd.n5834 gnd.n4523 99.6594
R12628 gnd.n5832 gnd.n5831 99.6594
R12629 gnd.n5827 gnd.n4530 99.6594
R12630 gnd.n5825 gnd.n5824 99.6594
R12631 gnd.n5820 gnd.n4537 99.6594
R12632 gnd.n5818 gnd.n5817 99.6594
R12633 gnd.n5813 gnd.n4544 99.6594
R12634 gnd.n5811 gnd.n5810 99.6594
R12635 gnd.n5806 gnd.n4551 99.6594
R12636 gnd.n5804 gnd.n5803 99.6594
R12637 gnd.n5799 gnd.n4560 99.6594
R12638 gnd.n5797 gnd.n5796 99.6594
R12639 gnd.n5792 gnd.n5791 99.6594
R12640 gnd.n4989 gnd.n4988 99.6594
R12641 gnd.n4983 gnd.n4900 99.6594
R12642 gnd.n4980 gnd.n4901 99.6594
R12643 gnd.n4976 gnd.n4902 99.6594
R12644 gnd.n4972 gnd.n4903 99.6594
R12645 gnd.n4968 gnd.n4904 99.6594
R12646 gnd.n4964 gnd.n4905 99.6594
R12647 gnd.n4960 gnd.n4906 99.6594
R12648 gnd.n4956 gnd.n4907 99.6594
R12649 gnd.n4952 gnd.n4908 99.6594
R12650 gnd.n4948 gnd.n4909 99.6594
R12651 gnd.n4944 gnd.n4910 99.6594
R12652 gnd.n4991 gnd.n4899 99.6594
R12653 gnd.n6722 gnd.n6721 99.6594
R12654 gnd.n6727 gnd.n6726 99.6594
R12655 gnd.n6730 gnd.n6729 99.6594
R12656 gnd.n6735 gnd.n6734 99.6594
R12657 gnd.n6738 gnd.n6737 99.6594
R12658 gnd.n6743 gnd.n6742 99.6594
R12659 gnd.n6746 gnd.n6745 99.6594
R12660 gnd.n6751 gnd.n6750 99.6594
R12661 gnd.n6754 gnd.n80 99.6594
R12662 gnd.n3472 gnd.n3471 99.6594
R12663 gnd.n3475 gnd.n3474 99.6594
R12664 gnd.n3491 gnd.n3490 99.6594
R12665 gnd.n3494 gnd.n3493 99.6594
R12666 gnd.n3510 gnd.n3509 99.6594
R12667 gnd.n3513 gnd.n3512 99.6594
R12668 gnd.n3529 gnd.n3528 99.6594
R12669 gnd.n3532 gnd.n3531 99.6594
R12670 gnd.n3550 gnd.n3549 99.6594
R12671 gnd.n2099 gnd.n2098 99.6594
R12672 gnd.n2102 gnd.n2101 99.6594
R12673 gnd.n2112 gnd.n2111 99.6594
R12674 gnd.n2121 gnd.n2120 99.6594
R12675 gnd.n2124 gnd.n2123 99.6594
R12676 gnd.n2135 gnd.n2134 99.6594
R12677 gnd.n2144 gnd.n2143 99.6594
R12678 gnd.n2147 gnd.n2146 99.6594
R12679 gnd.n2158 gnd.n2157 99.6594
R12680 gnd.n2334 gnd.n820 99.6594
R12681 gnd.n2331 gnd.n821 99.6594
R12682 gnd.n2327 gnd.n822 99.6594
R12683 gnd.n2323 gnd.n823 99.6594
R12684 gnd.n2319 gnd.n824 99.6594
R12685 gnd.n2315 gnd.n825 99.6594
R12686 gnd.n2311 gnd.n826 99.6594
R12687 gnd.n2307 gnd.n827 99.6594
R12688 gnd.n2303 gnd.n828 99.6594
R12689 gnd.n2332 gnd.n820 99.6594
R12690 gnd.n2328 gnd.n821 99.6594
R12691 gnd.n2324 gnd.n822 99.6594
R12692 gnd.n2320 gnd.n823 99.6594
R12693 gnd.n2316 gnd.n824 99.6594
R12694 gnd.n2312 gnd.n825 99.6594
R12695 gnd.n2308 gnd.n826 99.6594
R12696 gnd.n2304 gnd.n827 99.6594
R12697 gnd.n2291 gnd.n828 99.6594
R12698 gnd.n2157 gnd.n2156 99.6594
R12699 gnd.n2146 gnd.n2145 99.6594
R12700 gnd.n2143 gnd.n2136 99.6594
R12701 gnd.n2134 gnd.n2133 99.6594
R12702 gnd.n2123 gnd.n2122 99.6594
R12703 gnd.n2120 gnd.n2113 99.6594
R12704 gnd.n2111 gnd.n2110 99.6594
R12705 gnd.n2101 gnd.n2100 99.6594
R12706 gnd.n2098 gnd.n2097 99.6594
R12707 gnd.n3473 gnd.n3472 99.6594
R12708 gnd.n3474 gnd.n3456 99.6594
R12709 gnd.n3492 gnd.n3491 99.6594
R12710 gnd.n3493 gnd.n3447 99.6594
R12711 gnd.n3511 gnd.n3510 99.6594
R12712 gnd.n3512 gnd.n3438 99.6594
R12713 gnd.n3530 gnd.n3529 99.6594
R12714 gnd.n3531 gnd.n3429 99.6594
R12715 gnd.n3551 gnd.n3550 99.6594
R12716 gnd.n6755 gnd.n6754 99.6594
R12717 gnd.n6750 gnd.n6749 99.6594
R12718 gnd.n6745 gnd.n6744 99.6594
R12719 gnd.n6742 gnd.n6741 99.6594
R12720 gnd.n6737 gnd.n6736 99.6594
R12721 gnd.n6734 gnd.n6733 99.6594
R12722 gnd.n6729 gnd.n6728 99.6594
R12723 gnd.n6726 gnd.n6725 99.6594
R12724 gnd.n6721 gnd.n6720 99.6594
R12725 gnd.n4989 gnd.n4912 99.6594
R12726 gnd.n4981 gnd.n4900 99.6594
R12727 gnd.n4977 gnd.n4901 99.6594
R12728 gnd.n4973 gnd.n4902 99.6594
R12729 gnd.n4969 gnd.n4903 99.6594
R12730 gnd.n4965 gnd.n4904 99.6594
R12731 gnd.n4961 gnd.n4905 99.6594
R12732 gnd.n4957 gnd.n4906 99.6594
R12733 gnd.n4953 gnd.n4907 99.6594
R12734 gnd.n4949 gnd.n4908 99.6594
R12735 gnd.n4945 gnd.n4909 99.6594
R12736 gnd.n4941 gnd.n4910 99.6594
R12737 gnd.n4992 gnd.n4991 99.6594
R12738 gnd.n5791 gnd.n4562 99.6594
R12739 gnd.n5798 gnd.n5797 99.6594
R12740 gnd.n4560 gnd.n4552 99.6594
R12741 gnd.n5805 gnd.n5804 99.6594
R12742 gnd.n4551 gnd.n4545 99.6594
R12743 gnd.n5812 gnd.n5811 99.6594
R12744 gnd.n4544 gnd.n4538 99.6594
R12745 gnd.n5819 gnd.n5818 99.6594
R12746 gnd.n4537 gnd.n4531 99.6594
R12747 gnd.n5826 gnd.n5825 99.6594
R12748 gnd.n4530 gnd.n4524 99.6594
R12749 gnd.n5833 gnd.n5832 99.6594
R12750 gnd.n4523 gnd.n4520 99.6594
R12751 gnd.n5149 gnd.n5148 99.6594
R12752 gnd.n4834 gnd.n4812 99.6594
R12753 gnd.n4840 gnd.n4813 99.6594
R12754 gnd.n4844 gnd.n4814 99.6594
R12755 gnd.n4850 gnd.n4815 99.6594
R12756 gnd.n4854 gnd.n4816 99.6594
R12757 gnd.n4860 gnd.n4817 99.6594
R12758 gnd.n4818 gnd.n4802 99.6594
R12759 gnd.n5844 gnd.n5843 99.6594
R12760 gnd.n4516 gnd.n4508 99.6594
R12761 gnd.n5851 gnd.n5850 99.6594
R12762 gnd.n4507 gnd.n4501 99.6594
R12763 gnd.n5858 gnd.n5857 99.6594
R12764 gnd.n4500 gnd.n4494 99.6594
R12765 gnd.n5865 gnd.n5864 99.6594
R12766 gnd.n4493 gnd.n4490 99.6594
R12767 gnd.n4481 gnd.n832 99.6594
R12768 gnd.n4473 gnd.n802 99.6594
R12769 gnd.n4469 gnd.n803 99.6594
R12770 gnd.n4465 gnd.n804 99.6594
R12771 gnd.n4461 gnd.n805 99.6594
R12772 gnd.n4457 gnd.n806 99.6594
R12773 gnd.n4453 gnd.n807 99.6594
R12774 gnd.n4449 gnd.n808 99.6594
R12775 gnd.n4444 gnd.n809 99.6594
R12776 gnd.n4440 gnd.n810 99.6594
R12777 gnd.n4436 gnd.n811 99.6594
R12778 gnd.n4432 gnd.n812 99.6594
R12779 gnd.n4428 gnd.n813 99.6594
R12780 gnd.n4424 gnd.n814 99.6594
R12781 gnd.n4420 gnd.n815 99.6594
R12782 gnd.n4416 gnd.n816 99.6594
R12783 gnd.n4412 gnd.n817 99.6594
R12784 gnd.n872 gnd.n818 99.6594
R12785 gnd.n4404 gnd.n819 99.6594
R12786 gnd.n2671 gnd.n2670 99.6594
R12787 gnd.n2027 gnd.n2019 99.6594
R12788 gnd.n2678 gnd.n2677 99.6594
R12789 gnd.n2018 gnd.n2012 99.6594
R12790 gnd.n2685 gnd.n2684 99.6594
R12791 gnd.n2011 gnd.n2005 99.6594
R12792 gnd.n2692 gnd.n2691 99.6594
R12793 gnd.n2004 gnd.n1998 99.6594
R12794 gnd.n2699 gnd.n2698 99.6594
R12795 gnd.n2702 gnd.n2701 99.6594
R12796 gnd.n1969 gnd.n1943 99.6594
R12797 gnd.n1973 gnd.n1944 99.6594
R12798 gnd.n1977 gnd.n1945 99.6594
R12799 gnd.n1981 gnd.n1946 99.6594
R12800 gnd.n1985 gnd.n1947 99.6594
R12801 gnd.n1989 gnd.n1948 99.6594
R12802 gnd.n1951 gnd.n1949 99.6594
R12803 gnd.n1995 gnd.n1950 99.6594
R12804 gnd.n3794 gnd.n3793 99.6594
R12805 gnd.n3796 gnd.n3785 99.6594
R12806 gnd.n3805 gnd.n3804 99.6594
R12807 gnd.n3806 gnd.n3781 99.6594
R12808 gnd.n3815 gnd.n3814 99.6594
R12809 gnd.n3816 gnd.n3777 99.6594
R12810 gnd.n3826 gnd.n3825 99.6594
R12811 gnd.n3775 gnd.n1357 99.6594
R12812 gnd.n3839 gnd.n3838 99.6594
R12813 gnd.n3840 gnd.n1353 99.6594
R12814 gnd.n3849 gnd.n3848 99.6594
R12815 gnd.n3850 gnd.n1349 99.6594
R12816 gnd.n3859 gnd.n3858 99.6594
R12817 gnd.n3860 gnd.n1345 99.6594
R12818 gnd.n3869 gnd.n3868 99.6594
R12819 gnd.n3870 gnd.n1341 99.6594
R12820 gnd.n3880 gnd.n3879 99.6594
R12821 gnd.n3883 gnd.n3882 99.6594
R12822 gnd.n153 gnd.n150 99.6594
R12823 gnd.n6813 gnd.n6812 99.6594
R12824 gnd.n149 gnd.n143 99.6594
R12825 gnd.n6820 gnd.n6819 99.6594
R12826 gnd.n142 gnd.n136 99.6594
R12827 gnd.n6827 gnd.n6826 99.6594
R12828 gnd.n135 gnd.n129 99.6594
R12829 gnd.n6834 gnd.n6833 99.6594
R12830 gnd.n128 gnd.n122 99.6594
R12831 gnd.n6841 gnd.n6840 99.6594
R12832 gnd.n121 gnd.n115 99.6594
R12833 gnd.n6851 gnd.n6850 99.6594
R12834 gnd.n114 gnd.n108 99.6594
R12835 gnd.n6858 gnd.n6857 99.6594
R12836 gnd.n107 gnd.n101 99.6594
R12837 gnd.n6865 gnd.n6864 99.6594
R12838 gnd.n100 gnd.n94 99.6594
R12839 gnd.n6872 gnd.n6871 99.6594
R12840 gnd.n93 gnd.n90 99.6594
R12841 gnd.n2205 gnd.n2204 99.6594
R12842 gnd.n2105 gnd.n2074 99.6594
R12843 gnd.n2107 gnd.n2075 99.6594
R12844 gnd.n2117 gnd.n2076 99.6594
R12845 gnd.n2128 gnd.n2077 99.6594
R12846 gnd.n2130 gnd.n2078 99.6594
R12847 gnd.n2140 gnd.n2079 99.6594
R12848 gnd.n2153 gnd.n2080 99.6594
R12849 gnd.n2154 gnd.n2081 99.6594
R12850 gnd.n2082 gnd.n2038 99.6594
R12851 gnd.n2084 gnd.n2083 99.6594
R12852 gnd.n2085 gnd.n2043 99.6594
R12853 gnd.n2086 gnd.n2049 99.6594
R12854 gnd.n2088 gnd.n2051 99.6594
R12855 gnd.n2205 gnd.n2090 99.6594
R12856 gnd.n2106 gnd.n2074 99.6594
R12857 gnd.n2116 gnd.n2075 99.6594
R12858 gnd.n2127 gnd.n2076 99.6594
R12859 gnd.n2129 gnd.n2077 99.6594
R12860 gnd.n2139 gnd.n2078 99.6594
R12861 gnd.n2152 gnd.n2079 99.6594
R12862 gnd.n2155 gnd.n2080 99.6594
R12863 gnd.n2081 gnd.n2037 99.6594
R12864 gnd.n2082 gnd.n2039 99.6594
R12865 gnd.n2084 gnd.n2042 99.6594
R12866 gnd.n2085 gnd.n2044 99.6594
R12867 gnd.n2086 gnd.n2050 99.6594
R12868 gnd.n2088 gnd.n2087 99.6594
R12869 gnd.n3481 gnd.n3461 99.6594
R12870 gnd.n3485 gnd.n3483 99.6594
R12871 gnd.n3500 gnd.n3452 99.6594
R12872 gnd.n3504 gnd.n3502 99.6594
R12873 gnd.n3519 gnd.n3443 99.6594
R12874 gnd.n3523 gnd.n3521 99.6594
R12875 gnd.n3538 gnd.n3434 99.6594
R12876 gnd.n3541 gnd.n3540 99.6594
R12877 gnd.n3542 gnd.n3423 99.6594
R12878 gnd.n3561 gnd.n3560 99.6594
R12879 gnd.n3562 gnd.n3419 99.6594
R12880 gnd.n3571 gnd.n3570 99.6594
R12881 gnd.n3572 gnd.n3415 99.6594
R12882 gnd.n3584 gnd.n3583 99.6594
R12883 gnd.n3583 gnd.n3582 99.6594
R12884 gnd.n3573 gnd.n3572 99.6594
R12885 gnd.n3570 gnd.n3569 99.6594
R12886 gnd.n3563 gnd.n3562 99.6594
R12887 gnd.n3560 gnd.n3559 99.6594
R12888 gnd.n3543 gnd.n3542 99.6594
R12889 gnd.n3540 gnd.n3539 99.6594
R12890 gnd.n3522 gnd.n3434 99.6594
R12891 gnd.n3521 gnd.n3520 99.6594
R12892 gnd.n3503 gnd.n3443 99.6594
R12893 gnd.n3502 gnd.n3501 99.6594
R12894 gnd.n3484 gnd.n3452 99.6594
R12895 gnd.n3483 gnd.n3482 99.6594
R12896 gnd.n3461 gnd.n1191 99.6594
R12897 gnd.n2045 gnd.t179 98.63
R12898 gnd.n6752 gnd.t165 98.63
R12899 gnd.n3426 gnd.t156 98.63
R12900 gnd.n2148 gnd.t174 98.63
R12901 gnd.n3830 gnd.t153 98.63
R12902 gnd.n1337 gnd.t125 98.63
R12903 gnd.n156 gnd.t120 98.63
R12904 gnd.n6844 gnd.t138 98.63
R12905 gnd.n852 gnd.t211 98.63
R12906 gnd.n874 gnd.t205 98.63
R12907 gnd.n2292 gnd.t193 98.63
R12908 gnd.n2024 gnd.t135 98.63
R12909 gnd.n1935 gnd.t168 98.63
R12910 gnd.n3574 gnd.t159 98.63
R12911 gnd.n1854 gnd.t186 92.8196
R12912 gnd.n1398 gnd.t198 92.8196
R12913 gnd.n1851 gnd.t218 92.8118
R12914 gnd.n3637 gnd.t128 92.8118
R12915 gnd.n1802 gnd.n1801 81.8399
R12916 gnd.n3832 gnd.n3774 78.9125
R12917 gnd.n2711 gnd.n2707 78.9125
R12918 gnd.n6626 gnd.n162 76.3231
R12919 gnd.n4863 gnd.t113 74.8376
R12920 gnd.n4514 gnd.t143 74.8376
R12921 gnd.n1855 gnd.t185 72.8438
R12922 gnd.n1399 gnd.t199 72.8438
R12923 gnd.n1803 gnd.n1796 72.8411
R12924 gnd.n1809 gnd.n1794 72.8411
R12925 gnd.n3633 gnd.n3632 72.8411
R12926 gnd.n2046 gnd.t178 72.836
R12927 gnd.n1852 gnd.t217 72.836
R12928 gnd.n3638 gnd.t129 72.836
R12929 gnd.n6753 gnd.t166 72.836
R12930 gnd.n3427 gnd.t155 72.836
R12931 gnd.n2149 gnd.t175 72.836
R12932 gnd.n3831 gnd.t152 72.836
R12933 gnd.n1338 gnd.t124 72.836
R12934 gnd.n157 gnd.t121 72.836
R12935 gnd.n6845 gnd.t139 72.836
R12936 gnd.n853 gnd.t210 72.836
R12937 gnd.n875 gnd.t204 72.836
R12938 gnd.n2293 gnd.t192 72.836
R12939 gnd.n2025 gnd.t136 72.836
R12940 gnd.n1936 gnd.t169 72.836
R12941 gnd.n3575 gnd.t160 72.836
R12942 gnd.n3698 gnd.n1366 71.676
R12943 gnd.n3694 gnd.n1367 71.676
R12944 gnd.n3690 gnd.n1368 71.676
R12945 gnd.n3686 gnd.n1369 71.676
R12946 gnd.n3682 gnd.n1370 71.676
R12947 gnd.n3678 gnd.n1371 71.676
R12948 gnd.n3674 gnd.n1372 71.676
R12949 gnd.n3670 gnd.n1373 71.676
R12950 gnd.n3666 gnd.n1374 71.676
R12951 gnd.n3662 gnd.n1375 71.676
R12952 gnd.n3658 gnd.n1376 71.676
R12953 gnd.n3654 gnd.n1377 71.676
R12954 gnd.n3650 gnd.n1378 71.676
R12955 gnd.n3646 gnd.n1379 71.676
R12956 gnd.n3641 gnd.n1380 71.676
R12957 gnd.n1381 gnd.n1364 71.676
R12958 gnd.n3770 gnd.n1363 71.676
R12959 gnd.n3768 gnd.n3767 71.676
R12960 gnd.n3762 gnd.n1396 71.676
R12961 gnd.n3758 gnd.n1395 71.676
R12962 gnd.n3754 gnd.n1394 71.676
R12963 gnd.n3750 gnd.n1393 71.676
R12964 gnd.n3746 gnd.n1392 71.676
R12965 gnd.n3742 gnd.n1391 71.676
R12966 gnd.n3738 gnd.n1390 71.676
R12967 gnd.n3734 gnd.n1389 71.676
R12968 gnd.n3730 gnd.n1388 71.676
R12969 gnd.n3726 gnd.n1387 71.676
R12970 gnd.n3722 gnd.n1386 71.676
R12971 gnd.n3718 gnd.n1385 71.676
R12972 gnd.n3714 gnd.n1384 71.676
R12973 gnd.n3710 gnd.n1383 71.676
R12974 gnd.n3706 gnd.n1382 71.676
R12975 gnd.n2773 gnd.n2772 71.676
R12976 gnd.n1850 gnd.n1817 71.676
R12977 gnd.n2765 gnd.n1818 71.676
R12978 gnd.n2761 gnd.n1819 71.676
R12979 gnd.n2757 gnd.n1820 71.676
R12980 gnd.n2753 gnd.n1821 71.676
R12981 gnd.n2749 gnd.n1822 71.676
R12982 gnd.n2745 gnd.n1823 71.676
R12983 gnd.n2741 gnd.n1824 71.676
R12984 gnd.n2737 gnd.n1825 71.676
R12985 gnd.n2733 gnd.n1826 71.676
R12986 gnd.n2729 gnd.n1827 71.676
R12987 gnd.n2725 gnd.n1828 71.676
R12988 gnd.n2721 gnd.n1829 71.676
R12989 gnd.n2717 gnd.n1830 71.676
R12990 gnd.n2713 gnd.n1831 71.676
R12991 gnd.n2709 gnd.n1833 71.676
R12992 gnd.n1929 gnd.n1834 71.676
R12993 gnd.n1924 gnd.n1835 71.676
R12994 gnd.n1920 gnd.n1836 71.676
R12995 gnd.n1916 gnd.n1837 71.676
R12996 gnd.n1912 gnd.n1838 71.676
R12997 gnd.n1908 gnd.n1839 71.676
R12998 gnd.n1904 gnd.n1840 71.676
R12999 gnd.n1900 gnd.n1841 71.676
R13000 gnd.n1896 gnd.n1842 71.676
R13001 gnd.n1892 gnd.n1843 71.676
R13002 gnd.n1888 gnd.n1844 71.676
R13003 gnd.n1884 gnd.n1845 71.676
R13004 gnd.n1880 gnd.n1846 71.676
R13005 gnd.n1876 gnd.n1847 71.676
R13006 gnd.n1872 gnd.n1848 71.676
R13007 gnd.n2772 gnd.n1814 71.676
R13008 gnd.n2766 gnd.n1817 71.676
R13009 gnd.n2762 gnd.n1818 71.676
R13010 gnd.n2758 gnd.n1819 71.676
R13011 gnd.n2754 gnd.n1820 71.676
R13012 gnd.n2750 gnd.n1821 71.676
R13013 gnd.n2746 gnd.n1822 71.676
R13014 gnd.n2742 gnd.n1823 71.676
R13015 gnd.n2738 gnd.n1824 71.676
R13016 gnd.n2734 gnd.n1825 71.676
R13017 gnd.n2730 gnd.n1826 71.676
R13018 gnd.n2726 gnd.n1827 71.676
R13019 gnd.n2722 gnd.n1828 71.676
R13020 gnd.n2718 gnd.n1829 71.676
R13021 gnd.n2714 gnd.n1830 71.676
R13022 gnd.n2710 gnd.n1832 71.676
R13023 gnd.n1930 gnd.n1833 71.676
R13024 gnd.n1925 gnd.n1834 71.676
R13025 gnd.n1921 gnd.n1835 71.676
R13026 gnd.n1917 gnd.n1836 71.676
R13027 gnd.n1913 gnd.n1837 71.676
R13028 gnd.n1909 gnd.n1838 71.676
R13029 gnd.n1905 gnd.n1839 71.676
R13030 gnd.n1901 gnd.n1840 71.676
R13031 gnd.n1897 gnd.n1841 71.676
R13032 gnd.n1893 gnd.n1842 71.676
R13033 gnd.n1889 gnd.n1843 71.676
R13034 gnd.n1885 gnd.n1844 71.676
R13035 gnd.n1881 gnd.n1845 71.676
R13036 gnd.n1877 gnd.n1846 71.676
R13037 gnd.n1873 gnd.n1847 71.676
R13038 gnd.n1869 gnd.n1848 71.676
R13039 gnd.n3709 gnd.n1382 71.676
R13040 gnd.n3713 gnd.n1383 71.676
R13041 gnd.n3717 gnd.n1384 71.676
R13042 gnd.n3721 gnd.n1385 71.676
R13043 gnd.n3725 gnd.n1386 71.676
R13044 gnd.n3729 gnd.n1387 71.676
R13045 gnd.n3733 gnd.n1388 71.676
R13046 gnd.n3737 gnd.n1389 71.676
R13047 gnd.n3741 gnd.n1390 71.676
R13048 gnd.n3745 gnd.n1391 71.676
R13049 gnd.n3749 gnd.n1392 71.676
R13050 gnd.n3753 gnd.n1393 71.676
R13051 gnd.n3757 gnd.n1394 71.676
R13052 gnd.n3761 gnd.n1395 71.676
R13053 gnd.n1397 gnd.n1396 71.676
R13054 gnd.n3769 gnd.n3768 71.676
R13055 gnd.n3773 gnd.n3772 71.676
R13056 gnd.n3640 gnd.n1381 71.676
R13057 gnd.n3645 gnd.n1380 71.676
R13058 gnd.n3649 gnd.n1379 71.676
R13059 gnd.n3653 gnd.n1378 71.676
R13060 gnd.n3657 gnd.n1377 71.676
R13061 gnd.n3661 gnd.n1376 71.676
R13062 gnd.n3665 gnd.n1375 71.676
R13063 gnd.n3669 gnd.n1374 71.676
R13064 gnd.n3673 gnd.n1373 71.676
R13065 gnd.n3677 gnd.n1372 71.676
R13066 gnd.n3681 gnd.n1371 71.676
R13067 gnd.n3685 gnd.n1370 71.676
R13068 gnd.n3689 gnd.n1369 71.676
R13069 gnd.n3693 gnd.n1368 71.676
R13070 gnd.n3697 gnd.n1367 71.676
R13071 gnd.n1404 gnd.n1366 71.676
R13072 gnd.n8 gnd.t279 69.1507
R13073 gnd.n14 gnd.t53 68.4792
R13074 gnd.n13 gnd.t230 68.4792
R13075 gnd.n12 gnd.t83 68.4792
R13076 gnd.n11 gnd.t45 68.4792
R13077 gnd.n10 gnd.t47 68.4792
R13078 gnd.n9 gnd.t110 68.4792
R13079 gnd.n8 gnd.t263 68.4792
R13080 gnd.n4990 gnd.n4894 64.369
R13081 gnd.n4482 gnd.n830 63.0944
R13082 gnd.n6881 gnd.n83 63.0944
R13083 gnd.n1927 gnd.n1855 59.5399
R13084 gnd.n3764 gnd.n1399 59.5399
R13085 gnd.n1853 gnd.n1852 59.5399
R13086 gnd.n3643 gnd.n3638 59.5399
R13087 gnd.n2775 gnd.n1812 59.1804
R13088 gnd.n5874 gnd.n4483 57.3586
R13089 gnd.n5088 gnd.t61 56.607
R13090 gnd.n40 gnd.t280 56.607
R13091 gnd.n5065 gnd.t249 56.407
R13092 gnd.n5076 gnd.t63 56.407
R13093 gnd.n17 gnd.t268 56.407
R13094 gnd.n28 gnd.t80 56.407
R13095 gnd.n5097 gnd.t29 55.8337
R13096 gnd.n5074 gnd.t219 55.8337
R13097 gnd.n5085 gnd.t37 55.8337
R13098 gnd.n49 gnd.t237 55.8337
R13099 gnd.n26 gnd.t67 55.8337
R13100 gnd.n37 gnd.t259 55.8337
R13101 gnd.n1800 gnd.n1799 54.358
R13102 gnd.n3630 gnd.n3629 54.358
R13103 gnd.n5088 gnd.n5087 53.0052
R13104 gnd.n5090 gnd.n5089 53.0052
R13105 gnd.n5092 gnd.n5091 53.0052
R13106 gnd.n5094 gnd.n5093 53.0052
R13107 gnd.n5096 gnd.n5095 53.0052
R13108 gnd.n5065 gnd.n5064 53.0052
R13109 gnd.n5067 gnd.n5066 53.0052
R13110 gnd.n5069 gnd.n5068 53.0052
R13111 gnd.n5071 gnd.n5070 53.0052
R13112 gnd.n5073 gnd.n5072 53.0052
R13113 gnd.n5076 gnd.n5075 53.0052
R13114 gnd.n5078 gnd.n5077 53.0052
R13115 gnd.n5080 gnd.n5079 53.0052
R13116 gnd.n5082 gnd.n5081 53.0052
R13117 gnd.n5084 gnd.n5083 53.0052
R13118 gnd.n48 gnd.n47 53.0052
R13119 gnd.n46 gnd.n45 53.0052
R13120 gnd.n44 gnd.n43 53.0052
R13121 gnd.n42 gnd.n41 53.0052
R13122 gnd.n40 gnd.n39 53.0052
R13123 gnd.n25 gnd.n24 53.0052
R13124 gnd.n23 gnd.n22 53.0052
R13125 gnd.n21 gnd.n20 53.0052
R13126 gnd.n19 gnd.n18 53.0052
R13127 gnd.n17 gnd.n16 53.0052
R13128 gnd.n36 gnd.n35 53.0052
R13129 gnd.n34 gnd.n33 53.0052
R13130 gnd.n32 gnd.n31 53.0052
R13131 gnd.n30 gnd.n29 53.0052
R13132 gnd.n28 gnd.n27 53.0052
R13133 gnd.n3621 gnd.n3620 52.4801
R13134 gnd.n5701 gnd.t287 52.3082
R13135 gnd.n5669 gnd.t253 52.3082
R13136 gnd.n5637 gnd.t251 52.3082
R13137 gnd.n5606 gnd.t108 52.3082
R13138 gnd.n5574 gnd.t76 52.3082
R13139 gnd.n5542 gnd.t13 52.3082
R13140 gnd.n5510 gnd.t257 52.3082
R13141 gnd.n5479 gnd.t5 52.3082
R13142 gnd.n5531 gnd.n5499 51.4173
R13143 gnd.n5595 gnd.n5594 50.455
R13144 gnd.n5563 gnd.n5562 50.455
R13145 gnd.n5531 gnd.n5530 50.455
R13146 gnd.n4937 gnd.n4936 45.1884
R13147 gnd.n4558 gnd.n4557 45.1884
R13148 gnd.n3701 gnd.n3636 44.3322
R13149 gnd.n1803 gnd.n1802 44.3189
R13150 gnd.n2047 gnd.n2046 42.2793
R13151 gnd.n4938 gnd.n4937 42.2793
R13152 gnd.n4559 gnd.n4558 42.2793
R13153 gnd.n4864 gnd.n4863 42.2793
R13154 gnd.n4515 gnd.n4514 42.2793
R13155 gnd.n6757 gnd.n6753 42.2793
R13156 gnd.n3428 gnd.n3427 42.2793
R13157 gnd.n2150 gnd.n2149 42.2793
R13158 gnd.n1339 gnd.n1338 42.2793
R13159 gnd.n6809 gnd.n157 42.2793
R13160 gnd.n6846 gnd.n6845 42.2793
R13161 gnd.n4446 gnd.n853 42.2793
R13162 gnd.n876 gnd.n875 42.2793
R13163 gnd.n2294 gnd.n2293 42.2793
R13164 gnd.n2026 gnd.n2025 42.2793
R13165 gnd.n3576 gnd.n3575 42.2793
R13166 gnd.n1801 gnd.n1800 41.6274
R13167 gnd.n3631 gnd.n3630 41.6274
R13168 gnd.n1810 gnd.n1809 40.8975
R13169 gnd.n3634 gnd.n3633 40.8975
R13170 gnd.n3832 gnd.n3831 36.9518
R13171 gnd.n2707 gnd.n1936 36.9518
R13172 gnd.n6064 gnd.n6063 36.5879
R13173 gnd.n6063 gnd.n597 36.5879
R13174 gnd.n6057 gnd.n597 36.5879
R13175 gnd.n6057 gnd.n6056 36.5879
R13176 gnd.n6056 gnd.n6055 36.5879
R13177 gnd.n6055 gnd.n605 36.5879
R13178 gnd.n6049 gnd.n605 36.5879
R13179 gnd.n6049 gnd.n6048 36.5879
R13180 gnd.n6048 gnd.n6047 36.5879
R13181 gnd.n6047 gnd.n613 36.5879
R13182 gnd.n6041 gnd.n613 36.5879
R13183 gnd.n6041 gnd.n6040 36.5879
R13184 gnd.n6040 gnd.n6039 36.5879
R13185 gnd.n6039 gnd.n621 36.5879
R13186 gnd.n6033 gnd.n621 36.5879
R13187 gnd.n6033 gnd.n6032 36.5879
R13188 gnd.n6032 gnd.n6031 36.5879
R13189 gnd.n6031 gnd.n629 36.5879
R13190 gnd.n6025 gnd.n629 36.5879
R13191 gnd.n6025 gnd.n6024 36.5879
R13192 gnd.n6024 gnd.n6023 36.5879
R13193 gnd.n6023 gnd.n637 36.5879
R13194 gnd.n6017 gnd.n637 36.5879
R13195 gnd.n6017 gnd.n6016 36.5879
R13196 gnd.n6016 gnd.n6015 36.5879
R13197 gnd.n6015 gnd.n645 36.5879
R13198 gnd.n6009 gnd.n645 36.5879
R13199 gnd.n6009 gnd.n6008 36.5879
R13200 gnd.n6008 gnd.n6007 36.5879
R13201 gnd.n6007 gnd.n653 36.5879
R13202 gnd.n6001 gnd.n653 36.5879
R13203 gnd.n6001 gnd.n6000 36.5879
R13204 gnd.n6000 gnd.n5999 36.5879
R13205 gnd.n5999 gnd.n661 36.5879
R13206 gnd.n5993 gnd.n661 36.5879
R13207 gnd.n5993 gnd.n5992 36.5879
R13208 gnd.n5992 gnd.n5991 36.5879
R13209 gnd.n5991 gnd.n669 36.5879
R13210 gnd.n5985 gnd.n669 36.5879
R13211 gnd.n5985 gnd.n5984 36.5879
R13212 gnd.n5984 gnd.n5983 36.5879
R13213 gnd.n5983 gnd.n677 36.5879
R13214 gnd.n5977 gnd.n677 36.5879
R13215 gnd.n5977 gnd.n5976 36.5879
R13216 gnd.n5976 gnd.n5975 36.5879
R13217 gnd.n5975 gnd.n685 36.5879
R13218 gnd.n5969 gnd.n685 36.5879
R13219 gnd.n5969 gnd.n5968 36.5879
R13220 gnd.n5968 gnd.n5967 36.5879
R13221 gnd.n5967 gnd.n693 36.5879
R13222 gnd.n5961 gnd.n693 36.5879
R13223 gnd.n5961 gnd.n5960 36.5879
R13224 gnd.n5960 gnd.n5959 36.5879
R13225 gnd.n5959 gnd.n701 36.5879
R13226 gnd.n5953 gnd.n701 36.5879
R13227 gnd.n5953 gnd.n5952 36.5879
R13228 gnd.n5952 gnd.n5951 36.5879
R13229 gnd.n5951 gnd.n709 36.5879
R13230 gnd.n5945 gnd.n709 36.5879
R13231 gnd.n5945 gnd.n5944 36.5879
R13232 gnd.n5944 gnd.n5943 36.5879
R13233 gnd.n5943 gnd.n717 36.5879
R13234 gnd.n5937 gnd.n717 36.5879
R13235 gnd.n5937 gnd.n5936 36.5879
R13236 gnd.n5936 gnd.n5935 36.5879
R13237 gnd.n5935 gnd.n725 36.5879
R13238 gnd.n5929 gnd.n725 36.5879
R13239 gnd.n5929 gnd.n5928 36.5879
R13240 gnd.n5928 gnd.n5927 36.5879
R13241 gnd.n5927 gnd.n733 36.5879
R13242 gnd.n5921 gnd.n733 36.5879
R13243 gnd.n5921 gnd.n5920 36.5879
R13244 gnd.n5920 gnd.n5919 36.5879
R13245 gnd.n5919 gnd.n741 36.5879
R13246 gnd.n5913 gnd.n741 36.5879
R13247 gnd.n5913 gnd.n5912 36.5879
R13248 gnd.n5912 gnd.n5911 36.5879
R13249 gnd.n5911 gnd.n749 36.5879
R13250 gnd.n5905 gnd.n749 36.5879
R13251 gnd.n5905 gnd.n5904 36.5879
R13252 gnd.n5904 gnd.n5903 36.5879
R13253 gnd.n5903 gnd.n757 36.5879
R13254 gnd.n5897 gnd.n757 36.5879
R13255 gnd.n1809 gnd.n1808 35.055
R13256 gnd.n1804 gnd.n1803 35.055
R13257 gnd.n3623 gnd.n3622 35.055
R13258 gnd.n3633 gnd.n3619 35.055
R13259 gnd.n5000 gnd.n4894 31.8661
R13260 gnd.n5000 gnd.n4999 31.8661
R13261 gnd.n5008 gnd.n4883 31.8661
R13262 gnd.n5016 gnd.n4883 31.8661
R13263 gnd.n5016 gnd.n4877 31.8661
R13264 gnd.n5024 gnd.n4877 31.8661
R13265 gnd.n5024 gnd.n4870 31.8661
R13266 gnd.n5136 gnd.n4870 31.8661
R13267 gnd.n5146 gnd.n4803 31.8661
R13268 gnd.n2351 gnd.n830 31.8661
R13269 gnd.n4395 gnd.n884 31.8661
R13270 gnd.n4395 gnd.n886 31.8661
R13271 gnd.n4389 gnd.n886 31.8661
R13272 gnd.n4389 gnd.n898 31.8661
R13273 gnd.n4383 gnd.n909 31.8661
R13274 gnd.n4377 gnd.n909 31.8661
R13275 gnd.n4371 gnd.n926 31.8661
R13276 gnd.n4365 gnd.n936 31.8661
R13277 gnd.n4365 gnd.n939 31.8661
R13278 gnd.n4359 gnd.n949 31.8661
R13279 gnd.n2420 gnd.n949 31.8661
R13280 gnd.n4351 gnd.n960 31.8661
R13281 gnd.n2572 gnd.n1082 31.8661
R13282 gnd.n2577 gnd.n2575 31.8661
R13283 gnd.n2577 gnd.n2576 31.8661
R13284 gnd.n2586 gnd.n2585 31.8661
R13285 gnd.n4145 gnd.n1194 31.8661
R13286 gnd.n4139 gnd.n4138 31.8661
R13287 gnd.n4138 gnd.n4137 31.8661
R13288 gnd.n4131 gnd.n1212 31.8661
R13289 gnd.n6663 gnd.n230 31.8661
R13290 gnd.n6671 gnd.n222 31.8661
R13291 gnd.n6671 gnd.n224 31.8661
R13292 gnd.n6679 gnd.n202 31.8661
R13293 gnd.n6687 gnd.n202 31.8661
R13294 gnd.n6695 gnd.n194 31.8661
R13295 gnd.n6703 gnd.n186 31.8661
R13296 gnd.n6703 gnd.n188 31.8661
R13297 gnd.n6711 gnd.n170 31.8661
R13298 gnd.n6793 gnd.n170 31.8661
R13299 gnd.n6793 gnd.n161 31.8661
R13300 gnd.n6801 gnd.n161 31.8661
R13301 gnd.n6881 gnd.n81 31.8661
R13302 gnd.n3707 gnd.n1400 31.3761
R13303 gnd.n1870 gnd.n1867 31.3761
R13304 gnd.n926 gnd.t7 30.9101
R13305 gnd.n6695 gnd.t48 30.9101
R13306 gnd.n2046 gnd.n2045 25.7944
R13307 gnd.n4863 gnd.n4862 25.7944
R13308 gnd.n4514 gnd.n4513 25.7944
R13309 gnd.n6753 gnd.n6752 25.7944
R13310 gnd.n3427 gnd.n3426 25.7944
R13311 gnd.n2149 gnd.n2148 25.7944
R13312 gnd.n3831 gnd.n3830 25.7944
R13313 gnd.n1338 gnd.n1337 25.7944
R13314 gnd.n157 gnd.n156 25.7944
R13315 gnd.n6845 gnd.n6844 25.7944
R13316 gnd.n853 gnd.n852 25.7944
R13317 gnd.n875 gnd.n874 25.7944
R13318 gnd.n2293 gnd.n2292 25.7944
R13319 gnd.n2025 gnd.n2024 25.7944
R13320 gnd.n1936 gnd.n1935 25.7944
R13321 gnd.n3575 gnd.n3574 25.7944
R13322 gnd.n5158 gnd.n4804 24.8557
R13323 gnd.n5168 gnd.n4787 24.8557
R13324 gnd.n4790 gnd.n4778 24.8557
R13325 gnd.n5189 gnd.n4779 24.8557
R13326 gnd.n5199 gnd.n4761 24.8557
R13327 gnd.n5210 gnd.n5209 24.8557
R13328 gnd.n5229 gnd.n4747 24.8557
R13329 gnd.n5230 gnd.n4736 24.8557
R13330 gnd.n5241 gnd.n5240 24.8557
R13331 gnd.n5251 gnd.n4729 24.8557
R13332 gnd.n5260 gnd.n4721 24.8557
R13333 gnd.n5272 gnd.n5271 24.8557
R13334 gnd.n5059 gnd.n4713 24.8557
R13335 gnd.n5282 gnd.n4703 24.8557
R13336 gnd.n5291 gnd.n4696 24.8557
R13337 gnd.n4689 gnd.n4679 24.8557
R13338 gnd.n4672 gnd.n4666 24.8557
R13339 gnd.n5346 gnd.n5345 24.8557
R13340 gnd.n5356 gnd.n5355 24.8557
R13341 gnd.n4657 gnd.n4649 24.8557
R13342 gnd.n5367 gnd.n4634 24.8557
R13343 gnd.n5386 gnd.n5385 24.8557
R13344 gnd.n5396 gnd.n4627 24.8557
R13345 gnd.n5409 gnd.n4616 24.8557
R13346 gnd.n5400 gnd.n5399 24.8557
R13347 gnd.n5432 gnd.n5431 24.8557
R13348 gnd.n5442 gnd.n4603 24.8557
R13349 gnd.n5454 gnd.n4595 24.8557
R13350 gnd.n5753 gnd.n5752 24.8557
R13351 gnd.n5768 gnd.n5767 24.8557
R13352 gnd.n5889 gnd.n776 24.8557
R13353 gnd.n5888 gnd.n779 24.8557
R13354 gnd.n5737 gnd.n788 24.8557
R13355 gnd.n5875 gnd.n799 24.8557
R13356 gnd.n5179 gnd.t4 23.2624
R13357 gnd.n4806 gnd.t112 22.6251
R13358 gnd.n4371 gnd.t35 21.9878
R13359 gnd.t23 gnd.n194 21.9878
R13360 gnd.n5897 gnd.n5896 21.9529
R13361 gnd.t107 gnd.n4811 21.3504
R13362 gnd.t73 gnd.n957 21.0318
R13363 gnd.n2431 gnd.n973 21.0318
R13364 gnd.n4338 gnd.n978 21.0318
R13365 gnd.n2454 gnd.n2453 21.0318
R13366 gnd.n4332 gnd.n987 21.0318
R13367 gnd.n4325 gnd.n995 21.0318
R13368 gnd.n2502 gnd.n998 21.0318
R13369 gnd.n2510 gnd.n1008 21.0318
R13370 gnd.n4313 gnd.n1016 21.0318
R13371 gnd.n2518 gnd.n2235 21.0318
R13372 gnd.n4307 gnd.n1026 21.0318
R13373 gnd.n4301 gnd.n1037 21.0318
R13374 gnd.n2554 gnd.n1040 21.0318
R13375 gnd.n2534 gnd.n1050 21.0318
R13376 gnd.n4289 gnd.n1058 21.0318
R13377 gnd.n2543 gnd.n1061 21.0318
R13378 gnd.n4283 gnd.n1069 21.0318
R13379 gnd.n4277 gnd.n1079 21.0318
R13380 gnd.n4130 gnd.n1215 21.0318
R13381 gnd.n4124 gnd.n1227 21.0318
R13382 gnd.n3899 gnd.n1325 21.0318
R13383 gnd.n4010 gnd.n4009 21.0318
R13384 gnd.n3992 gnd.n1318 21.0318
R13385 gnd.n4030 gnd.n1310 21.0318
R13386 gnd.n4029 gnd.n1299 21.0318
R13387 gnd.n1302 gnd.n1289 21.0318
R13388 gnd.n4052 gnd.n1291 21.0318
R13389 gnd.n4062 gnd.n1281 21.0318
R13390 gnd.n4061 gnd.n1270 21.0318
R13391 gnd.n1274 gnd.n1260 21.0318
R13392 gnd.n4086 gnd.n1262 21.0318
R13393 gnd.n4095 gnd.n248 21.0318
R13394 gnd.n6644 gnd.n6643 21.0318
R13395 gnd.n6649 gnd.n246 21.0318
R13396 gnd.n3966 gnd.n236 21.0318
R13397 gnd.n232 gnd.t54 21.0318
R13398 gnd.t89 gnd.n4580 20.7131
R13399 gnd.n4359 gnd.t0 20.7131
R13400 gnd.t222 gnd.n990 20.7131
R13401 gnd.t40 gnd.n1251 20.7131
R13402 gnd.n224 gnd.t18 20.7131
R13403 gnd.n2572 gnd.n1996 20.3945
R13404 gnd.n1212 gnd.n1204 20.3945
R13405 gnd.t91 gnd.n4626 20.0758
R13406 gnd.n4383 gnd.t28 20.0758
R13407 gnd.t68 gnd.n1029 20.0758
R13408 gnd.t10 gnd.n4040 20.0758
R13409 gnd.n188 gnd.t66 20.0758
R13410 gnd.n1855 gnd.n1854 19.9763
R13411 gnd.n1399 gnd.n1398 19.9763
R13412 gnd.n1852 gnd.n1851 19.9763
R13413 gnd.n3638 gnd.n3637 19.9763
R13414 gnd.n1797 gnd.t172 19.8005
R13415 gnd.n1797 gnd.t189 19.8005
R13416 gnd.n1798 gnd.t146 19.8005
R13417 gnd.n1798 gnd.t196 19.8005
R13418 gnd.n3627 gnd.t182 19.8005
R13419 gnd.n3627 gnd.t163 19.8005
R13420 gnd.n3628 gnd.t117 19.8005
R13421 gnd.n3628 gnd.t208 19.8005
R13422 gnd.n1794 gnd.n1793 19.5087
R13423 gnd.n1807 gnd.n1794 19.5087
R13424 gnd.n1805 gnd.n1796 19.5087
R13425 gnd.n3632 gnd.n3626 19.5087
R13426 gnd.n5322 gnd.t95 19.4385
R13427 gnd.n2638 gnd.n2637 19.3944
R13428 gnd.n2637 gnd.n2636 19.3944
R13429 gnd.n2636 gnd.n2057 19.3944
R13430 gnd.n2632 gnd.n2057 19.3944
R13431 gnd.n2632 gnd.n2631 19.3944
R13432 gnd.n2631 gnd.n2630 19.3944
R13433 gnd.n2630 gnd.n2627 19.3944
R13434 gnd.n2627 gnd.n1787 19.3944
R13435 gnd.n2782 gnd.n1787 19.3944
R13436 gnd.n2782 gnd.n1784 19.3944
R13437 gnd.n2787 gnd.n1784 19.3944
R13438 gnd.n2787 gnd.n1785 19.3944
R13439 gnd.n1785 gnd.n1766 19.3944
R13440 gnd.n2813 gnd.n1766 19.3944
R13441 gnd.n2813 gnd.n1763 19.3944
R13442 gnd.n2824 gnd.n1763 19.3944
R13443 gnd.n2824 gnd.n1764 19.3944
R13444 gnd.n2820 gnd.n1764 19.3944
R13445 gnd.n2820 gnd.n2819 19.3944
R13446 gnd.n2819 gnd.n1718 19.3944
R13447 gnd.n2898 gnd.n1718 19.3944
R13448 gnd.n2898 gnd.n1715 19.3944
R13449 gnd.n2922 gnd.n1715 19.3944
R13450 gnd.n2922 gnd.n1716 19.3944
R13451 gnd.n2918 gnd.n1716 19.3944
R13452 gnd.n2918 gnd.n2917 19.3944
R13453 gnd.n2917 gnd.n2916 19.3944
R13454 gnd.n2916 gnd.n2908 19.3944
R13455 gnd.n2912 gnd.n2908 19.3944
R13456 gnd.n2912 gnd.n2911 19.3944
R13457 gnd.n2911 gnd.n1668 19.3944
R13458 gnd.n1668 gnd.n1666 19.3944
R13459 gnd.n3000 gnd.n1666 19.3944
R13460 gnd.n3000 gnd.n1664 19.3944
R13461 gnd.n3004 gnd.n1664 19.3944
R13462 gnd.n3004 gnd.n1639 19.3944
R13463 gnd.n3052 gnd.n1639 19.3944
R13464 gnd.n3052 gnd.n1640 19.3944
R13465 gnd.n3048 gnd.n1640 19.3944
R13466 gnd.n3048 gnd.n1616 19.3944
R13467 gnd.n3110 gnd.n1616 19.3944
R13468 gnd.n3110 gnd.n1617 19.3944
R13469 gnd.n3106 gnd.n1617 19.3944
R13470 gnd.n3106 gnd.n3105 19.3944
R13471 gnd.n3105 gnd.n3104 19.3944
R13472 gnd.n3104 gnd.n3091 19.3944
R13473 gnd.n3100 gnd.n3091 19.3944
R13474 gnd.n3100 gnd.n3099 19.3944
R13475 gnd.n3099 gnd.n3098 19.3944
R13476 gnd.n3098 gnd.n1558 19.3944
R13477 gnd.n3218 gnd.n1558 19.3944
R13478 gnd.n3218 gnd.n1555 19.3944
R13479 gnd.n3223 gnd.n1555 19.3944
R13480 gnd.n3223 gnd.n1556 19.3944
R13481 gnd.n1556 gnd.n1529 19.3944
R13482 gnd.n3257 gnd.n1529 19.3944
R13483 gnd.n3257 gnd.n1526 19.3944
R13484 gnd.n3276 gnd.n1526 19.3944
R13485 gnd.n3276 gnd.n1527 19.3944
R13486 gnd.n3272 gnd.n1527 19.3944
R13487 gnd.n3272 gnd.n3271 19.3944
R13488 gnd.n3271 gnd.n3270 19.3944
R13489 gnd.n3270 gnd.n3265 19.3944
R13490 gnd.n3266 gnd.n3265 19.3944
R13491 gnd.n3266 gnd.n1474 19.3944
R13492 gnd.n3350 gnd.n1474 19.3944
R13493 gnd.n3350 gnd.n1471 19.3944
R13494 gnd.n3355 gnd.n1471 19.3944
R13495 gnd.n3355 gnd.n1472 19.3944
R13496 gnd.n1472 gnd.n1447 19.3944
R13497 gnd.n3392 gnd.n1447 19.3944
R13498 gnd.n3392 gnd.n1445 19.3944
R13499 gnd.n3396 gnd.n1445 19.3944
R13500 gnd.n3396 gnd.n1444 19.3944
R13501 gnd.n3402 gnd.n1444 19.3944
R13502 gnd.n3402 gnd.n1442 19.3944
R13503 gnd.n3406 gnd.n1442 19.3944
R13504 gnd.n3407 gnd.n3406 19.3944
R13505 gnd.n3410 gnd.n3407 19.3944
R13506 gnd.n3410 gnd.n1439 19.3944
R13507 gnd.n3590 gnd.n1439 19.3944
R13508 gnd.n3590 gnd.n1440 19.3944
R13509 gnd.n2644 gnd.n2643 19.3944
R13510 gnd.n2643 gnd.n2642 19.3944
R13511 gnd.n2642 gnd.n2052 19.3944
R13512 gnd.n2203 gnd.n2202 19.3944
R13513 gnd.n2202 gnd.n2092 19.3944
R13514 gnd.n2195 gnd.n2092 19.3944
R13515 gnd.n2195 gnd.n2194 19.3944
R13516 gnd.n2194 gnd.n2108 19.3944
R13517 gnd.n2187 gnd.n2108 19.3944
R13518 gnd.n2187 gnd.n2186 19.3944
R13519 gnd.n2186 gnd.n2118 19.3944
R13520 gnd.n2179 gnd.n2118 19.3944
R13521 gnd.n2179 gnd.n2178 19.3944
R13522 gnd.n2178 gnd.n2131 19.3944
R13523 gnd.n2171 gnd.n2131 19.3944
R13524 gnd.n2171 gnd.n2170 19.3944
R13525 gnd.n2170 gnd.n2141 19.3944
R13526 gnd.n2163 gnd.n2141 19.3944
R13527 gnd.n2163 gnd.n2162 19.3944
R13528 gnd.n2162 gnd.n2036 19.3944
R13529 gnd.n2655 gnd.n2036 19.3944
R13530 gnd.n2655 gnd.n2654 19.3944
R13531 gnd.n2654 gnd.n2653 19.3944
R13532 gnd.n2653 gnd.n2040 19.3944
R13533 gnd.n2649 gnd.n2040 19.3944
R13534 gnd.n2649 gnd.n2648 19.3944
R13535 gnd.n2648 gnd.n2647 19.3944
R13536 gnd.n4987 gnd.n4986 19.3944
R13537 gnd.n4986 gnd.n4985 19.3944
R13538 gnd.n4985 gnd.n4984 19.3944
R13539 gnd.n4984 gnd.n4982 19.3944
R13540 gnd.n4982 gnd.n4979 19.3944
R13541 gnd.n4979 gnd.n4978 19.3944
R13542 gnd.n4978 gnd.n4975 19.3944
R13543 gnd.n4975 gnd.n4974 19.3944
R13544 gnd.n4974 gnd.n4971 19.3944
R13545 gnd.n4971 gnd.n4970 19.3944
R13546 gnd.n4970 gnd.n4967 19.3944
R13547 gnd.n4967 gnd.n4966 19.3944
R13548 gnd.n4966 gnd.n4963 19.3944
R13549 gnd.n4963 gnd.n4962 19.3944
R13550 gnd.n4962 gnd.n4959 19.3944
R13551 gnd.n4959 gnd.n4958 19.3944
R13552 gnd.n4958 gnd.n4955 19.3944
R13553 gnd.n4955 gnd.n4954 19.3944
R13554 gnd.n4954 gnd.n4951 19.3944
R13555 gnd.n4951 gnd.n4950 19.3944
R13556 gnd.n4950 gnd.n4947 19.3944
R13557 gnd.n4947 gnd.n4946 19.3944
R13558 gnd.n4943 gnd.n4942 19.3944
R13559 gnd.n4942 gnd.n4898 19.3944
R13560 gnd.n4993 gnd.n4898 19.3944
R13561 gnd.n5795 gnd.n4561 19.3944
R13562 gnd.n5795 gnd.n5794 19.3944
R13563 gnd.n5794 gnd.n5793 19.3944
R13564 gnd.n5837 gnd.n5836 19.3944
R13565 gnd.n5836 gnd.n5835 19.3944
R13566 gnd.n5835 gnd.n4522 19.3944
R13567 gnd.n5830 gnd.n4522 19.3944
R13568 gnd.n5830 gnd.n5829 19.3944
R13569 gnd.n5829 gnd.n5828 19.3944
R13570 gnd.n5828 gnd.n4529 19.3944
R13571 gnd.n5823 gnd.n4529 19.3944
R13572 gnd.n5823 gnd.n5822 19.3944
R13573 gnd.n5822 gnd.n5821 19.3944
R13574 gnd.n5821 gnd.n4536 19.3944
R13575 gnd.n5816 gnd.n4536 19.3944
R13576 gnd.n5816 gnd.n5815 19.3944
R13577 gnd.n5815 gnd.n5814 19.3944
R13578 gnd.n5814 gnd.n4543 19.3944
R13579 gnd.n5809 gnd.n4543 19.3944
R13580 gnd.n5809 gnd.n5808 19.3944
R13581 gnd.n5808 gnd.n5807 19.3944
R13582 gnd.n5807 gnd.n4550 19.3944
R13583 gnd.n5802 gnd.n4550 19.3944
R13584 gnd.n5802 gnd.n5801 19.3944
R13585 gnd.n5801 gnd.n5800 19.3944
R13586 gnd.n5160 gnd.n4795 19.3944
R13587 gnd.n5170 gnd.n4795 19.3944
R13588 gnd.n5171 gnd.n5170 19.3944
R13589 gnd.n5171 gnd.n4776 19.3944
R13590 gnd.n5191 gnd.n4776 19.3944
R13591 gnd.n5191 gnd.n4769 19.3944
R13592 gnd.n5201 gnd.n4769 19.3944
R13593 gnd.n5202 gnd.n5201 19.3944
R13594 gnd.n5202 gnd.n4752 19.3944
R13595 gnd.n5222 gnd.n4752 19.3944
R13596 gnd.n5222 gnd.n4744 19.3944
R13597 gnd.n5232 gnd.n4744 19.3944
R13598 gnd.n5233 gnd.n5232 19.3944
R13599 gnd.n5233 gnd.n4726 19.3944
R13600 gnd.n5253 gnd.n4726 19.3944
R13601 gnd.n5253 gnd.n4718 19.3944
R13602 gnd.n5263 gnd.n4718 19.3944
R13603 gnd.n5264 gnd.n5263 19.3944
R13604 gnd.n5264 gnd.n4701 19.3944
R13605 gnd.n5284 gnd.n4701 19.3944
R13606 gnd.n5284 gnd.n4693 19.3944
R13607 gnd.n5294 gnd.n4693 19.3944
R13608 gnd.n5295 gnd.n5294 19.3944
R13609 gnd.n5295 gnd.n4677 19.3944
R13610 gnd.n5314 gnd.n4677 19.3944
R13611 gnd.n5314 gnd.n4662 19.3944
R13612 gnd.n5348 gnd.n4662 19.3944
R13613 gnd.n5349 gnd.n5348 19.3944
R13614 gnd.n5350 gnd.n5349 19.3944
R13615 gnd.n5350 gnd.n4648 19.3944
R13616 gnd.n4648 gnd.n4642 19.3944
R13617 gnd.n5375 gnd.n4642 19.3944
R13618 gnd.n5376 gnd.n5375 19.3944
R13619 gnd.n5376 gnd.n4625 19.3944
R13620 gnd.n4625 gnd.n4623 19.3944
R13621 gnd.n5402 gnd.n4623 19.3944
R13622 gnd.n5403 gnd.n5402 19.3944
R13623 gnd.n5403 gnd.n4598 19.3944
R13624 gnd.n5449 gnd.n4598 19.3944
R13625 gnd.n5450 gnd.n5449 19.3944
R13626 gnd.n5450 gnd.n4591 19.3944
R13627 gnd.n5461 gnd.n4591 19.3944
R13628 gnd.n5463 gnd.n5461 19.3944
R13629 gnd.n5746 gnd.n5463 19.3944
R13630 gnd.n5746 gnd.n5745 19.3944
R13631 gnd.n5745 gnd.n5466 19.3944
R13632 gnd.n5741 gnd.n5466 19.3944
R13633 gnd.n5741 gnd.n5740 19.3944
R13634 gnd.n5740 gnd.n5739 19.3944
R13635 gnd.n5739 gnd.n5736 19.3944
R13636 gnd.n5736 gnd.n5735 19.3944
R13637 gnd.n5735 gnd.n5732 19.3944
R13638 gnd.n5732 gnd.n5731 19.3944
R13639 gnd.n5151 gnd.n5150 19.3944
R13640 gnd.n5150 gnd.n4809 19.3944
R13641 gnd.n4832 gnd.n4809 19.3944
R13642 gnd.n4835 gnd.n4832 19.3944
R13643 gnd.n4835 gnd.n4828 19.3944
R13644 gnd.n4839 gnd.n4828 19.3944
R13645 gnd.n4842 gnd.n4839 19.3944
R13646 gnd.n4845 gnd.n4842 19.3944
R13647 gnd.n4845 gnd.n4826 19.3944
R13648 gnd.n4849 gnd.n4826 19.3944
R13649 gnd.n4852 gnd.n4849 19.3944
R13650 gnd.n4855 gnd.n4852 19.3944
R13651 gnd.n4855 gnd.n4824 19.3944
R13652 gnd.n4859 gnd.n4824 19.3944
R13653 gnd.n5156 gnd.n5155 19.3944
R13654 gnd.n5155 gnd.n4785 19.3944
R13655 gnd.n5181 gnd.n4785 19.3944
R13656 gnd.n5181 gnd.n4783 19.3944
R13657 gnd.n5187 gnd.n4783 19.3944
R13658 gnd.n5187 gnd.n5186 19.3944
R13659 gnd.n5186 gnd.n4759 19.3944
R13660 gnd.n5212 gnd.n4759 19.3944
R13661 gnd.n5212 gnd.n4757 19.3944
R13662 gnd.n5218 gnd.n4757 19.3944
R13663 gnd.n5218 gnd.n5217 19.3944
R13664 gnd.n5217 gnd.n4734 19.3944
R13665 gnd.n5243 gnd.n4734 19.3944
R13666 gnd.n5243 gnd.n4732 19.3944
R13667 gnd.n5249 gnd.n4732 19.3944
R13668 gnd.n5249 gnd.n5248 19.3944
R13669 gnd.n5248 gnd.n4708 19.3944
R13670 gnd.n5274 gnd.n4708 19.3944
R13671 gnd.n5274 gnd.n4706 19.3944
R13672 gnd.n5280 gnd.n4706 19.3944
R13673 gnd.n5280 gnd.n5279 19.3944
R13674 gnd.n5279 gnd.n4684 19.3944
R13675 gnd.n5304 gnd.n4684 19.3944
R13676 gnd.n5304 gnd.n4682 19.3944
R13677 gnd.n5310 gnd.n4682 19.3944
R13678 gnd.n5310 gnd.n5309 19.3944
R13679 gnd.n5309 gnd.n4653 19.3944
R13680 gnd.n5358 gnd.n4653 19.3944
R13681 gnd.n5358 gnd.n4651 19.3944
R13682 gnd.n5362 gnd.n4651 19.3944
R13683 gnd.n5362 gnd.n4632 19.3944
R13684 gnd.n5388 gnd.n4632 19.3944
R13685 gnd.n5388 gnd.n4630 19.3944
R13686 gnd.n5394 gnd.n4630 19.3944
R13687 gnd.n5394 gnd.n5393 19.3944
R13688 gnd.n5393 gnd.n4608 19.3944
R13689 gnd.n5434 gnd.n4608 19.3944
R13690 gnd.n5434 gnd.n4606 19.3944
R13691 gnd.n5440 gnd.n4606 19.3944
R13692 gnd.n5440 gnd.n5439 19.3944
R13693 gnd.n5439 gnd.n4578 19.3944
R13694 gnd.n5755 gnd.n4578 19.3944
R13695 gnd.n5755 gnd.n4576 19.3944
R13696 gnd.n5765 gnd.n4576 19.3944
R13697 gnd.n5765 gnd.n5764 19.3944
R13698 gnd.n5764 gnd.n5763 19.3944
R13699 gnd.n5763 gnd.n782 19.3944
R13700 gnd.n5886 gnd.n782 19.3944
R13701 gnd.n5886 gnd.n5885 19.3944
R13702 gnd.n5885 gnd.n5884 19.3944
R13703 gnd.n5884 gnd.n786 19.3944
R13704 gnd.n4486 gnd.n786 19.3944
R13705 gnd.n5872 gnd.n4486 19.3944
R13706 gnd.n5869 gnd.n5868 19.3944
R13707 gnd.n5868 gnd.n5867 19.3944
R13708 gnd.n5867 gnd.n4492 19.3944
R13709 gnd.n5862 gnd.n4492 19.3944
R13710 gnd.n5862 gnd.n5861 19.3944
R13711 gnd.n5861 gnd.n5860 19.3944
R13712 gnd.n5860 gnd.n4499 19.3944
R13713 gnd.n5855 gnd.n4499 19.3944
R13714 gnd.n5855 gnd.n5854 19.3944
R13715 gnd.n5854 gnd.n5853 19.3944
R13716 gnd.n5853 gnd.n4506 19.3944
R13717 gnd.n5848 gnd.n4506 19.3944
R13718 gnd.n5848 gnd.n5847 19.3944
R13719 gnd.n5847 gnd.n5846 19.3944
R13720 gnd.n4997 gnd.n4896 19.3944
R13721 gnd.n4997 gnd.n4887 19.3944
R13722 gnd.n5010 gnd.n4887 19.3944
R13723 gnd.n5010 gnd.n4885 19.3944
R13724 gnd.n5014 gnd.n4885 19.3944
R13725 gnd.n5014 gnd.n4875 19.3944
R13726 gnd.n5026 gnd.n4875 19.3944
R13727 gnd.n5026 gnd.n4873 19.3944
R13728 gnd.n5134 gnd.n4873 19.3944
R13729 gnd.n5134 gnd.n5133 19.3944
R13730 gnd.n5133 gnd.n5132 19.3944
R13731 gnd.n5132 gnd.n5131 19.3944
R13732 gnd.n5131 gnd.n5128 19.3944
R13733 gnd.n5128 gnd.n5127 19.3944
R13734 gnd.n5127 gnd.n5126 19.3944
R13735 gnd.n5126 gnd.n5124 19.3944
R13736 gnd.n5124 gnd.n5123 19.3944
R13737 gnd.n5123 gnd.n5120 19.3944
R13738 gnd.n5120 gnd.n5119 19.3944
R13739 gnd.n5119 gnd.n5118 19.3944
R13740 gnd.n5118 gnd.n5116 19.3944
R13741 gnd.n5116 gnd.n5115 19.3944
R13742 gnd.n5115 gnd.n5111 19.3944
R13743 gnd.n5111 gnd.n5110 19.3944
R13744 gnd.n5110 gnd.n5109 19.3944
R13745 gnd.n5109 gnd.n5107 19.3944
R13746 gnd.n5107 gnd.n5106 19.3944
R13747 gnd.n5106 gnd.n5103 19.3944
R13748 gnd.n5103 gnd.n5102 19.3944
R13749 gnd.n5062 gnd.n5050 19.3944
R13750 gnd.n5061 gnd.n5057 19.3944
R13751 gnd.n5055 gnd.n5054 19.3944
R13752 gnd.n5051 gnd.n4670 19.3944
R13753 gnd.n5324 gnd.n4670 19.3944
R13754 gnd.n5324 gnd.n4668 19.3944
R13755 gnd.n5343 gnd.n4668 19.3944
R13756 gnd.n5343 gnd.n5342 19.3944
R13757 gnd.n5342 gnd.n5341 19.3944
R13758 gnd.n5341 gnd.n5339 19.3944
R13759 gnd.n5339 gnd.n5338 19.3944
R13760 gnd.n5338 gnd.n5336 19.3944
R13761 gnd.n5336 gnd.n5335 19.3944
R13762 gnd.n5335 gnd.n4614 19.3944
R13763 gnd.n5411 gnd.n4614 19.3944
R13764 gnd.n5411 gnd.n4612 19.3944
R13765 gnd.n5427 gnd.n4612 19.3944
R13766 gnd.n5427 gnd.n5426 19.3944
R13767 gnd.n5426 gnd.n5425 19.3944
R13768 gnd.n5425 gnd.n5423 19.3944
R13769 gnd.n5423 gnd.n5422 19.3944
R13770 gnd.n5422 gnd.n5420 19.3944
R13771 gnd.n5420 gnd.n4571 19.3944
R13772 gnd.n5770 gnd.n4571 19.3944
R13773 gnd.n5770 gnd.n4569 19.3944
R13774 gnd.n5776 gnd.n4569 19.3944
R13775 gnd.n5777 gnd.n5776 19.3944
R13776 gnd.n5780 gnd.n5777 19.3944
R13777 gnd.n5780 gnd.n4567 19.3944
R13778 gnd.n5784 gnd.n4567 19.3944
R13779 gnd.n5787 gnd.n5784 19.3944
R13780 gnd.n5788 gnd.n5787 19.3944
R13781 gnd.n5002 gnd.n4892 19.3944
R13782 gnd.n5002 gnd.n4890 19.3944
R13783 gnd.n5006 gnd.n4890 19.3944
R13784 gnd.n5006 gnd.n4881 19.3944
R13785 gnd.n5018 gnd.n4881 19.3944
R13786 gnd.n5018 gnd.n4879 19.3944
R13787 gnd.n5022 gnd.n4879 19.3944
R13788 gnd.n5022 gnd.n4868 19.3944
R13789 gnd.n5138 gnd.n4868 19.3944
R13790 gnd.n5138 gnd.n4822 19.3944
R13791 gnd.n5144 gnd.n4822 19.3944
R13792 gnd.n5144 gnd.n5143 19.3944
R13793 gnd.n5143 gnd.n4800 19.3944
R13794 gnd.n5165 gnd.n4800 19.3944
R13795 gnd.n5165 gnd.n4793 19.3944
R13796 gnd.n5176 gnd.n4793 19.3944
R13797 gnd.n5176 gnd.n5175 19.3944
R13798 gnd.n5175 gnd.n4774 19.3944
R13799 gnd.n5196 gnd.n4774 19.3944
R13800 gnd.n5196 gnd.n4767 19.3944
R13801 gnd.n5207 gnd.n4767 19.3944
R13802 gnd.n5207 gnd.n5206 19.3944
R13803 gnd.n5206 gnd.n4750 19.3944
R13804 gnd.n5227 gnd.n4750 19.3944
R13805 gnd.n5227 gnd.n4742 19.3944
R13806 gnd.n5238 gnd.n4742 19.3944
R13807 gnd.n5238 gnd.n5237 19.3944
R13808 gnd.n5237 gnd.n4724 19.3944
R13809 gnd.n5258 gnd.n4724 19.3944
R13810 gnd.n5258 gnd.n4716 19.3944
R13811 gnd.n5269 gnd.n4716 19.3944
R13812 gnd.n5269 gnd.n5268 19.3944
R13813 gnd.n5268 gnd.n4699 19.3944
R13814 gnd.n5289 gnd.n4699 19.3944
R13815 gnd.n5289 gnd.n4691 19.3944
R13816 gnd.n5299 gnd.n4691 19.3944
R13817 gnd.n5299 gnd.n4675 19.3944
R13818 gnd.n5320 gnd.n4675 19.3944
R13819 gnd.n5320 gnd.n5319 19.3944
R13820 gnd.n5319 gnd.n4659 19.3944
R13821 gnd.n5353 gnd.n4659 19.3944
R13822 gnd.n5353 gnd.n4644 19.3944
R13823 gnd.n5370 gnd.n4644 19.3944
R13824 gnd.n5370 gnd.n4640 19.3944
R13825 gnd.n5383 gnd.n4640 19.3944
R13826 gnd.n5383 gnd.n5382 19.3944
R13827 gnd.n5382 gnd.n4619 19.3944
R13828 gnd.n5407 gnd.n4619 19.3944
R13829 gnd.n5407 gnd.n5406 19.3944
R13830 gnd.n5406 gnd.n4600 19.3944
R13831 gnd.n5445 gnd.n4600 19.3944
R13832 gnd.n5445 gnd.n4593 19.3944
R13833 gnd.n5456 gnd.n4593 19.3944
R13834 gnd.n5456 gnd.n4587 19.3944
R13835 gnd.n5750 gnd.n4587 19.3944
R13836 gnd.n5750 gnd.n5749 19.3944
R13837 gnd.n5749 gnd.n770 19.3944
R13838 gnd.n5893 gnd.n770 19.3944
R13839 gnd.n5893 gnd.n5892 19.3944
R13840 gnd.n5892 gnd.n5891 19.3944
R13841 gnd.n5891 gnd.n774 19.3944
R13842 gnd.n794 gnd.n774 19.3944
R13843 gnd.n5879 gnd.n794 19.3944
R13844 gnd.n5879 gnd.n5878 19.3944
R13845 gnd.n5878 gnd.n5877 19.3944
R13846 gnd.n3892 gnd.n1334 19.3944
R13847 gnd.n3892 gnd.n1331 19.3944
R13848 gnd.n3897 gnd.n1331 19.3944
R13849 gnd.n3897 gnd.n1332 19.3944
R13850 gnd.n1332 gnd.n1316 19.3944
R13851 gnd.n4022 gnd.n1316 19.3944
R13852 gnd.n4022 gnd.n1313 19.3944
R13853 gnd.n4027 gnd.n1313 19.3944
R13854 gnd.n4027 gnd.n1314 19.3944
R13855 gnd.n1314 gnd.n1287 19.3944
R13856 gnd.n4054 gnd.n1287 19.3944
R13857 gnd.n4054 gnd.n1284 19.3944
R13858 gnd.n4059 gnd.n1284 19.3944
R13859 gnd.n4059 gnd.n1285 19.3944
R13860 gnd.n1285 gnd.n1258 19.3944
R13861 gnd.n4088 gnd.n1258 19.3944
R13862 gnd.n4088 gnd.n1254 19.3944
R13863 gnd.n4093 gnd.n1254 19.3944
R13864 gnd.n4093 gnd.n1256 19.3944
R13865 gnd.n1256 gnd.n1255 19.3944
R13866 gnd.n1255 gnd.n52 19.3944
R13867 gnd.n6913 gnd.n52 19.3944
R13868 gnd.n6913 gnd.n6912 19.3944
R13869 gnd.n6912 gnd.n6911 19.3944
R13870 gnd.n6911 gnd.n57 19.3944
R13871 gnd.n6907 gnd.n57 19.3944
R13872 gnd.n6907 gnd.n6906 19.3944
R13873 gnd.n6906 gnd.n6905 19.3944
R13874 gnd.n6905 gnd.n62 19.3944
R13875 gnd.n6901 gnd.n62 19.3944
R13876 gnd.n6901 gnd.n6900 19.3944
R13877 gnd.n6900 gnd.n6899 19.3944
R13878 gnd.n6899 gnd.n67 19.3944
R13879 gnd.n6895 gnd.n67 19.3944
R13880 gnd.n6895 gnd.n6894 19.3944
R13881 gnd.n6894 gnd.n6893 19.3944
R13882 gnd.n6893 gnd.n72 19.3944
R13883 gnd.n6889 gnd.n72 19.3944
R13884 gnd.n6889 gnd.n6888 19.3944
R13885 gnd.n6888 gnd.n6887 19.3944
R13886 gnd.n6887 gnd.n77 19.3944
R13887 gnd.n6883 gnd.n77 19.3944
R13888 gnd.n6782 gnd.n6781 19.3944
R13889 gnd.n6781 gnd.n6780 19.3944
R13890 gnd.n6780 gnd.n6723 19.3944
R13891 gnd.n6776 gnd.n6723 19.3944
R13892 gnd.n6776 gnd.n6775 19.3944
R13893 gnd.n6775 gnd.n6774 19.3944
R13894 gnd.n6774 gnd.n6731 19.3944
R13895 gnd.n6770 gnd.n6731 19.3944
R13896 gnd.n6770 gnd.n6769 19.3944
R13897 gnd.n6769 gnd.n6768 19.3944
R13898 gnd.n6768 gnd.n6739 19.3944
R13899 gnd.n6764 gnd.n6739 19.3944
R13900 gnd.n6764 gnd.n6763 19.3944
R13901 gnd.n6763 gnd.n6762 19.3944
R13902 gnd.n6762 gnd.n6747 19.3944
R13903 gnd.n6758 gnd.n6747 19.3944
R13904 gnd.n3470 gnd.n3464 19.3944
R13905 gnd.n3476 gnd.n3464 19.3944
R13906 gnd.n3476 gnd.n3457 19.3944
R13907 gnd.n3489 gnd.n3457 19.3944
R13908 gnd.n3489 gnd.n3455 19.3944
R13909 gnd.n3495 gnd.n3455 19.3944
R13910 gnd.n3495 gnd.n3448 19.3944
R13911 gnd.n3508 gnd.n3448 19.3944
R13912 gnd.n3508 gnd.n3446 19.3944
R13913 gnd.n3514 gnd.n3446 19.3944
R13914 gnd.n3514 gnd.n3439 19.3944
R13915 gnd.n3527 gnd.n3439 19.3944
R13916 gnd.n3527 gnd.n3437 19.3944
R13917 gnd.n3533 gnd.n3437 19.3944
R13918 gnd.n3533 gnd.n3430 19.3944
R13919 gnd.n3548 gnd.n3430 19.3944
R13920 gnd.n3467 gnd.n1230 19.3944
R13921 gnd.n4122 gnd.n1230 19.3944
R13922 gnd.n4122 gnd.n1231 19.3944
R13923 gnd.n4118 gnd.n1231 19.3944
R13924 gnd.n4118 gnd.n4117 19.3944
R13925 gnd.n4117 gnd.n4116 19.3944
R13926 gnd.n4116 gnd.n1237 19.3944
R13927 gnd.n4112 gnd.n1237 19.3944
R13928 gnd.n4112 gnd.n4111 19.3944
R13929 gnd.n4111 gnd.n4110 19.3944
R13930 gnd.n4110 gnd.n1242 19.3944
R13931 gnd.n4106 gnd.n1242 19.3944
R13932 gnd.n4106 gnd.n4105 19.3944
R13933 gnd.n4105 gnd.n4104 19.3944
R13934 gnd.n4104 gnd.n1247 19.3944
R13935 gnd.n4100 gnd.n1247 19.3944
R13936 gnd.n4100 gnd.n4099 19.3944
R13937 gnd.n4099 gnd.n4098 19.3944
R13938 gnd.n4098 gnd.n242 19.3944
R13939 gnd.n6651 gnd.n242 19.3944
R13940 gnd.n6651 gnd.n239 19.3944
R13941 gnd.n6655 gnd.n239 19.3944
R13942 gnd.n6655 gnd.n228 19.3944
R13943 gnd.n6665 gnd.n228 19.3944
R13944 gnd.n6665 gnd.n226 19.3944
R13945 gnd.n6669 gnd.n226 19.3944
R13946 gnd.n6669 gnd.n207 19.3944
R13947 gnd.n6681 gnd.n207 19.3944
R13948 gnd.n6681 gnd.n205 19.3944
R13949 gnd.n6685 gnd.n205 19.3944
R13950 gnd.n6685 gnd.n192 19.3944
R13951 gnd.n6697 gnd.n192 19.3944
R13952 gnd.n6697 gnd.n190 19.3944
R13953 gnd.n6701 gnd.n190 19.3944
R13954 gnd.n6701 gnd.n177 19.3944
R13955 gnd.n6713 gnd.n177 19.3944
R13956 gnd.n6713 gnd.n174 19.3944
R13957 gnd.n6791 gnd.n174 19.3944
R13958 gnd.n6791 gnd.n175 19.3944
R13959 gnd.n6787 gnd.n175 19.3944
R13960 gnd.n6787 gnd.n6786 19.3944
R13961 gnd.n6786 gnd.n6785 19.3944
R13962 gnd.n2096 gnd.n1085 19.3944
R13963 gnd.n2096 gnd.n2095 19.3944
R13964 gnd.n2199 gnd.n2095 19.3944
R13965 gnd.n2199 gnd.n2198 19.3944
R13966 gnd.n2198 gnd.n2103 19.3944
R13967 gnd.n2191 gnd.n2103 19.3944
R13968 gnd.n2191 gnd.n2190 19.3944
R13969 gnd.n2190 gnd.n2114 19.3944
R13970 gnd.n2183 gnd.n2114 19.3944
R13971 gnd.n2183 gnd.n2182 19.3944
R13972 gnd.n2182 gnd.n2125 19.3944
R13973 gnd.n2175 gnd.n2125 19.3944
R13974 gnd.n2175 gnd.n2174 19.3944
R13975 gnd.n2174 gnd.n2137 19.3944
R13976 gnd.n2167 gnd.n2137 19.3944
R13977 gnd.n2167 gnd.n2166 19.3944
R13978 gnd.n2461 gnd.n2458 19.3944
R13979 gnd.n2466 gnd.n2458 19.3944
R13980 gnd.n2466 gnd.n2456 19.3944
R13981 gnd.n2471 gnd.n2456 19.3944
R13982 gnd.n2471 gnd.n2247 19.3944
R13983 gnd.n2475 gnd.n2247 19.3944
R13984 gnd.n2475 gnd.n2245 19.3944
R13985 gnd.n2499 gnd.n2245 19.3944
R13986 gnd.n2499 gnd.n2498 19.3944
R13987 gnd.n2498 gnd.n2497 19.3944
R13988 gnd.n2497 gnd.n2481 19.3944
R13989 gnd.n2493 gnd.n2481 19.3944
R13990 gnd.n2493 gnd.n2492 19.3944
R13991 gnd.n2492 gnd.n2491 19.3944
R13992 gnd.n2491 gnd.n2489 19.3944
R13993 gnd.n2489 gnd.n2220 19.3944
R13994 gnd.n2220 gnd.n2218 19.3944
R13995 gnd.n2559 gnd.n2218 19.3944
R13996 gnd.n2559 gnd.n2216 19.3944
R13997 gnd.n2563 gnd.n2216 19.3944
R13998 gnd.n2563 gnd.n2214 19.3944
R13999 gnd.n2567 gnd.n2214 19.3944
R14000 gnd.n2567 gnd.n2212 19.3944
R14001 gnd.n2571 gnd.n2212 19.3944
R14002 gnd.n2571 gnd.n2210 19.3944
R14003 gnd.n2579 gnd.n2210 19.3944
R14004 gnd.n2579 gnd.n2208 19.3944
R14005 gnd.n2583 gnd.n2208 19.3944
R14006 gnd.n2583 gnd.n2072 19.3944
R14007 gnd.n2592 gnd.n2072 19.3944
R14008 gnd.n2592 gnd.n2070 19.3944
R14009 gnd.n2596 gnd.n2070 19.3944
R14010 gnd.n2596 gnd.n2066 19.3944
R14011 gnd.n2607 gnd.n2066 19.3944
R14012 gnd.n2607 gnd.n2064 19.3944
R14013 gnd.n2621 gnd.n2064 19.3944
R14014 gnd.n2621 gnd.n2620 19.3944
R14015 gnd.n2620 gnd.n2619 19.3944
R14016 gnd.n2619 gnd.n2614 19.3944
R14017 gnd.n2614 gnd.n1772 19.3944
R14018 gnd.n2802 gnd.n1772 19.3944
R14019 gnd.n2802 gnd.n1770 19.3944
R14020 gnd.n2806 gnd.n1770 19.3944
R14021 gnd.n2806 gnd.n1744 19.3944
R14022 gnd.n2845 gnd.n1744 19.3944
R14023 gnd.n2845 gnd.n1742 19.3944
R14024 gnd.n2849 gnd.n1742 19.3944
R14025 gnd.n2849 gnd.n1726 19.3944
R14026 gnd.n2887 gnd.n1726 19.3944
R14027 gnd.n2887 gnd.n1724 19.3944
R14028 gnd.n2893 gnd.n1724 19.3944
R14029 gnd.n2893 gnd.n2892 19.3944
R14030 gnd.n2892 gnd.n1700 19.3944
R14031 gnd.n2949 gnd.n1700 19.3944
R14032 gnd.n2949 gnd.n1698 19.3944
R14033 gnd.n2953 gnd.n1698 19.3944
R14034 gnd.n2953 gnd.n1682 19.3944
R14035 gnd.n2976 gnd.n1682 19.3944
R14036 gnd.n2976 gnd.n1680 19.3944
R14037 gnd.n2982 gnd.n1680 19.3944
R14038 gnd.n2982 gnd.n2981 19.3944
R14039 gnd.n2981 gnd.n1649 19.3944
R14040 gnd.n3027 gnd.n1649 19.3944
R14041 gnd.n3027 gnd.n1647 19.3944
R14042 gnd.n3031 gnd.n1647 19.3944
R14043 gnd.n3031 gnd.n1626 19.3944
R14044 gnd.n3067 gnd.n1626 19.3944
R14045 gnd.n3067 gnd.n1624 19.3944
R14046 gnd.n3071 gnd.n1624 19.3944
R14047 gnd.n3071 gnd.n1604 19.3944
R14048 gnd.n3123 gnd.n1604 19.3944
R14049 gnd.n3123 gnd.n1602 19.3944
R14050 gnd.n3127 gnd.n1602 19.3944
R14051 gnd.n3127 gnd.n1585 19.3944
R14052 gnd.n3148 gnd.n1585 19.3944
R14053 gnd.n3148 gnd.n1583 19.3944
R14054 gnd.n3152 gnd.n1583 19.3944
R14055 gnd.n3152 gnd.n1565 19.3944
R14056 gnd.n3208 gnd.n1565 19.3944
R14057 gnd.n3208 gnd.n1563 19.3944
R14058 gnd.n3212 gnd.n1563 19.3944
R14059 gnd.n3212 gnd.n1543 19.3944
R14060 gnd.n3237 gnd.n1543 19.3944
R14061 gnd.n3237 gnd.n1541 19.3944
R14062 gnd.n3243 gnd.n1541 19.3944
R14063 gnd.n3243 gnd.n3242 19.3944
R14064 gnd.n3242 gnd.n1515 19.3944
R14065 gnd.n3290 gnd.n1515 19.3944
R14066 gnd.n3290 gnd.n1513 19.3944
R14067 gnd.n3294 gnd.n1513 19.3944
R14068 gnd.n3294 gnd.n1496 19.3944
R14069 gnd.n3317 gnd.n1496 19.3944
R14070 gnd.n3317 gnd.n1494 19.3944
R14071 gnd.n3323 gnd.n1494 19.3944
R14072 gnd.n3323 gnd.n3322 19.3944
R14073 gnd.n3322 gnd.n1466 19.3944
R14074 gnd.n3361 gnd.n1466 19.3944
R14075 gnd.n3361 gnd.n1464 19.3944
R14076 gnd.n3368 gnd.n1464 19.3944
R14077 gnd.n3368 gnd.n3367 19.3944
R14078 gnd.n3367 gnd.n1413 19.3944
R14079 gnd.n3610 gnd.n1413 19.3944
R14080 gnd.n3610 gnd.n3609 19.3944
R14081 gnd.n3609 gnd.n3608 19.3944
R14082 gnd.n3608 gnd.n1417 19.3944
R14083 gnd.n1425 gnd.n1417 19.3944
R14084 gnd.n3599 gnd.n1425 19.3944
R14085 gnd.n3599 gnd.n3598 19.3944
R14086 gnd.n3598 gnd.n3597 19.3944
R14087 gnd.n3597 gnd.n1433 19.3944
R14088 gnd.n1433 gnd.n1197 19.3944
R14089 gnd.n4143 gnd.n1197 19.3944
R14090 gnd.n4143 gnd.n4142 19.3944
R14091 gnd.n4142 gnd.n4141 19.3944
R14092 gnd.n4141 gnd.n1201 19.3944
R14093 gnd.n4135 gnd.n1201 19.3944
R14094 gnd.n4135 gnd.n4134 19.3944
R14095 gnd.n4134 gnd.n4133 19.3944
R14096 gnd.n4133 gnd.n1210 19.3944
R14097 gnd.n3998 gnd.n1210 19.3944
R14098 gnd.n4001 gnd.n3998 19.3944
R14099 gnd.n4001 gnd.n3995 19.3944
R14100 gnd.n4007 gnd.n3995 19.3944
R14101 gnd.n4007 gnd.n4006 19.3944
R14102 gnd.n4006 gnd.n1307 19.3944
R14103 gnd.n4032 gnd.n1307 19.3944
R14104 gnd.n4032 gnd.n1305 19.3944
R14105 gnd.n4038 gnd.n1305 19.3944
R14106 gnd.n4038 gnd.n4037 19.3944
R14107 gnd.n4037 gnd.n1279 19.3944
R14108 gnd.n4064 gnd.n1279 19.3944
R14109 gnd.n4064 gnd.n1277 19.3944
R14110 gnd.n4077 gnd.n1277 19.3944
R14111 gnd.n4077 gnd.n4076 19.3944
R14112 gnd.n4076 gnd.n4075 19.3944
R14113 gnd.n4075 gnd.n4071 19.3944
R14114 gnd.n4071 gnd.n253 19.3944
R14115 gnd.n6641 gnd.n253 19.3944
R14116 gnd.n6641 gnd.n6640 19.3944
R14117 gnd.n6640 gnd.n6639 19.3944
R14118 gnd.n6639 gnd.n257 19.3944
R14119 gnd.n6422 gnd.n381 19.3944
R14120 gnd.n6428 gnd.n381 19.3944
R14121 gnd.n6428 gnd.n379 19.3944
R14122 gnd.n6432 gnd.n379 19.3944
R14123 gnd.n6432 gnd.n375 19.3944
R14124 gnd.n6438 gnd.n375 19.3944
R14125 gnd.n6438 gnd.n373 19.3944
R14126 gnd.n6442 gnd.n373 19.3944
R14127 gnd.n6442 gnd.n369 19.3944
R14128 gnd.n6448 gnd.n369 19.3944
R14129 gnd.n6448 gnd.n367 19.3944
R14130 gnd.n6452 gnd.n367 19.3944
R14131 gnd.n6452 gnd.n363 19.3944
R14132 gnd.n6458 gnd.n363 19.3944
R14133 gnd.n6458 gnd.n361 19.3944
R14134 gnd.n6462 gnd.n361 19.3944
R14135 gnd.n6462 gnd.n357 19.3944
R14136 gnd.n6468 gnd.n357 19.3944
R14137 gnd.n6468 gnd.n355 19.3944
R14138 gnd.n6472 gnd.n355 19.3944
R14139 gnd.n6472 gnd.n351 19.3944
R14140 gnd.n6478 gnd.n351 19.3944
R14141 gnd.n6478 gnd.n349 19.3944
R14142 gnd.n6482 gnd.n349 19.3944
R14143 gnd.n6482 gnd.n345 19.3944
R14144 gnd.n6488 gnd.n345 19.3944
R14145 gnd.n6488 gnd.n343 19.3944
R14146 gnd.n6492 gnd.n343 19.3944
R14147 gnd.n6492 gnd.n339 19.3944
R14148 gnd.n6498 gnd.n339 19.3944
R14149 gnd.n6498 gnd.n337 19.3944
R14150 gnd.n6502 gnd.n337 19.3944
R14151 gnd.n6502 gnd.n333 19.3944
R14152 gnd.n6508 gnd.n333 19.3944
R14153 gnd.n6508 gnd.n331 19.3944
R14154 gnd.n6512 gnd.n331 19.3944
R14155 gnd.n6512 gnd.n327 19.3944
R14156 gnd.n6518 gnd.n327 19.3944
R14157 gnd.n6518 gnd.n325 19.3944
R14158 gnd.n6522 gnd.n325 19.3944
R14159 gnd.n6522 gnd.n321 19.3944
R14160 gnd.n6528 gnd.n321 19.3944
R14161 gnd.n6528 gnd.n319 19.3944
R14162 gnd.n6532 gnd.n319 19.3944
R14163 gnd.n6532 gnd.n315 19.3944
R14164 gnd.n6538 gnd.n315 19.3944
R14165 gnd.n6538 gnd.n313 19.3944
R14166 gnd.n6542 gnd.n313 19.3944
R14167 gnd.n6542 gnd.n309 19.3944
R14168 gnd.n6548 gnd.n309 19.3944
R14169 gnd.n6548 gnd.n307 19.3944
R14170 gnd.n6552 gnd.n307 19.3944
R14171 gnd.n6552 gnd.n303 19.3944
R14172 gnd.n6558 gnd.n303 19.3944
R14173 gnd.n6558 gnd.n301 19.3944
R14174 gnd.n6562 gnd.n301 19.3944
R14175 gnd.n6562 gnd.n297 19.3944
R14176 gnd.n6568 gnd.n297 19.3944
R14177 gnd.n6568 gnd.n295 19.3944
R14178 gnd.n6572 gnd.n295 19.3944
R14179 gnd.n6572 gnd.n291 19.3944
R14180 gnd.n6578 gnd.n291 19.3944
R14181 gnd.n6578 gnd.n289 19.3944
R14182 gnd.n6582 gnd.n289 19.3944
R14183 gnd.n6582 gnd.n285 19.3944
R14184 gnd.n6588 gnd.n285 19.3944
R14185 gnd.n6588 gnd.n283 19.3944
R14186 gnd.n6592 gnd.n283 19.3944
R14187 gnd.n6592 gnd.n279 19.3944
R14188 gnd.n6598 gnd.n279 19.3944
R14189 gnd.n6598 gnd.n277 19.3944
R14190 gnd.n6602 gnd.n277 19.3944
R14191 gnd.n6602 gnd.n273 19.3944
R14192 gnd.n6608 gnd.n273 19.3944
R14193 gnd.n6608 gnd.n271 19.3944
R14194 gnd.n6612 gnd.n271 19.3944
R14195 gnd.n6612 gnd.n267 19.3944
R14196 gnd.n6618 gnd.n267 19.3944
R14197 gnd.n6618 gnd.n265 19.3944
R14198 gnd.n6622 gnd.n265 19.3944
R14199 gnd.n6622 gnd.n261 19.3944
R14200 gnd.n6629 gnd.n261 19.3944
R14201 gnd.n6629 gnd.n259 19.3944
R14202 gnd.n6634 gnd.n259 19.3944
R14203 gnd.n6067 gnd.n594 19.3944
R14204 gnd.n6071 gnd.n594 19.3944
R14205 gnd.n6071 gnd.n590 19.3944
R14206 gnd.n6077 gnd.n590 19.3944
R14207 gnd.n6077 gnd.n588 19.3944
R14208 gnd.n6081 gnd.n588 19.3944
R14209 gnd.n6081 gnd.n584 19.3944
R14210 gnd.n6087 gnd.n584 19.3944
R14211 gnd.n6087 gnd.n582 19.3944
R14212 gnd.n6091 gnd.n582 19.3944
R14213 gnd.n6091 gnd.n578 19.3944
R14214 gnd.n6097 gnd.n578 19.3944
R14215 gnd.n6097 gnd.n576 19.3944
R14216 gnd.n6101 gnd.n576 19.3944
R14217 gnd.n6101 gnd.n572 19.3944
R14218 gnd.n6107 gnd.n572 19.3944
R14219 gnd.n6107 gnd.n570 19.3944
R14220 gnd.n6111 gnd.n570 19.3944
R14221 gnd.n6111 gnd.n566 19.3944
R14222 gnd.n6117 gnd.n566 19.3944
R14223 gnd.n6117 gnd.n564 19.3944
R14224 gnd.n6121 gnd.n564 19.3944
R14225 gnd.n6121 gnd.n560 19.3944
R14226 gnd.n6127 gnd.n560 19.3944
R14227 gnd.n6127 gnd.n558 19.3944
R14228 gnd.n6131 gnd.n558 19.3944
R14229 gnd.n6131 gnd.n554 19.3944
R14230 gnd.n6137 gnd.n554 19.3944
R14231 gnd.n6137 gnd.n552 19.3944
R14232 gnd.n6141 gnd.n552 19.3944
R14233 gnd.n6141 gnd.n548 19.3944
R14234 gnd.n6147 gnd.n548 19.3944
R14235 gnd.n6147 gnd.n546 19.3944
R14236 gnd.n6151 gnd.n546 19.3944
R14237 gnd.n6151 gnd.n542 19.3944
R14238 gnd.n6157 gnd.n542 19.3944
R14239 gnd.n6157 gnd.n540 19.3944
R14240 gnd.n6161 gnd.n540 19.3944
R14241 gnd.n6161 gnd.n536 19.3944
R14242 gnd.n6167 gnd.n536 19.3944
R14243 gnd.n6167 gnd.n534 19.3944
R14244 gnd.n6171 gnd.n534 19.3944
R14245 gnd.n6171 gnd.n530 19.3944
R14246 gnd.n6177 gnd.n530 19.3944
R14247 gnd.n6177 gnd.n528 19.3944
R14248 gnd.n6181 gnd.n528 19.3944
R14249 gnd.n6181 gnd.n524 19.3944
R14250 gnd.n6187 gnd.n524 19.3944
R14251 gnd.n6187 gnd.n522 19.3944
R14252 gnd.n6191 gnd.n522 19.3944
R14253 gnd.n6191 gnd.n518 19.3944
R14254 gnd.n6197 gnd.n518 19.3944
R14255 gnd.n6197 gnd.n516 19.3944
R14256 gnd.n6201 gnd.n516 19.3944
R14257 gnd.n6201 gnd.n512 19.3944
R14258 gnd.n6207 gnd.n512 19.3944
R14259 gnd.n6207 gnd.n510 19.3944
R14260 gnd.n6211 gnd.n510 19.3944
R14261 gnd.n6211 gnd.n506 19.3944
R14262 gnd.n6217 gnd.n506 19.3944
R14263 gnd.n6217 gnd.n504 19.3944
R14264 gnd.n6221 gnd.n504 19.3944
R14265 gnd.n6221 gnd.n500 19.3944
R14266 gnd.n6227 gnd.n500 19.3944
R14267 gnd.n6227 gnd.n498 19.3944
R14268 gnd.n6231 gnd.n498 19.3944
R14269 gnd.n6231 gnd.n494 19.3944
R14270 gnd.n6237 gnd.n494 19.3944
R14271 gnd.n6237 gnd.n492 19.3944
R14272 gnd.n6241 gnd.n492 19.3944
R14273 gnd.n6241 gnd.n488 19.3944
R14274 gnd.n6247 gnd.n488 19.3944
R14275 gnd.n6247 gnd.n486 19.3944
R14276 gnd.n6251 gnd.n486 19.3944
R14277 gnd.n6251 gnd.n482 19.3944
R14278 gnd.n6257 gnd.n482 19.3944
R14279 gnd.n6257 gnd.n480 19.3944
R14280 gnd.n6261 gnd.n480 19.3944
R14281 gnd.n6261 gnd.n476 19.3944
R14282 gnd.n6267 gnd.n476 19.3944
R14283 gnd.n6267 gnd.n474 19.3944
R14284 gnd.n6271 gnd.n474 19.3944
R14285 gnd.n6271 gnd.n470 19.3944
R14286 gnd.n6277 gnd.n470 19.3944
R14287 gnd.n6277 gnd.n468 19.3944
R14288 gnd.n6281 gnd.n468 19.3944
R14289 gnd.n6281 gnd.n464 19.3944
R14290 gnd.n6287 gnd.n464 19.3944
R14291 gnd.n6287 gnd.n462 19.3944
R14292 gnd.n6291 gnd.n462 19.3944
R14293 gnd.n6291 gnd.n458 19.3944
R14294 gnd.n6297 gnd.n458 19.3944
R14295 gnd.n6297 gnd.n456 19.3944
R14296 gnd.n6301 gnd.n456 19.3944
R14297 gnd.n6301 gnd.n452 19.3944
R14298 gnd.n6307 gnd.n452 19.3944
R14299 gnd.n6307 gnd.n450 19.3944
R14300 gnd.n6311 gnd.n450 19.3944
R14301 gnd.n6311 gnd.n446 19.3944
R14302 gnd.n6317 gnd.n446 19.3944
R14303 gnd.n6317 gnd.n444 19.3944
R14304 gnd.n6321 gnd.n444 19.3944
R14305 gnd.n6321 gnd.n440 19.3944
R14306 gnd.n6327 gnd.n440 19.3944
R14307 gnd.n6327 gnd.n438 19.3944
R14308 gnd.n6331 gnd.n438 19.3944
R14309 gnd.n6331 gnd.n434 19.3944
R14310 gnd.n6337 gnd.n434 19.3944
R14311 gnd.n6337 gnd.n432 19.3944
R14312 gnd.n6341 gnd.n432 19.3944
R14313 gnd.n6341 gnd.n428 19.3944
R14314 gnd.n6347 gnd.n428 19.3944
R14315 gnd.n6347 gnd.n426 19.3944
R14316 gnd.n6351 gnd.n426 19.3944
R14317 gnd.n6351 gnd.n422 19.3944
R14318 gnd.n6357 gnd.n422 19.3944
R14319 gnd.n6357 gnd.n420 19.3944
R14320 gnd.n6361 gnd.n420 19.3944
R14321 gnd.n6361 gnd.n416 19.3944
R14322 gnd.n6367 gnd.n416 19.3944
R14323 gnd.n6367 gnd.n414 19.3944
R14324 gnd.n6371 gnd.n414 19.3944
R14325 gnd.n6371 gnd.n410 19.3944
R14326 gnd.n6377 gnd.n410 19.3944
R14327 gnd.n6377 gnd.n408 19.3944
R14328 gnd.n6381 gnd.n408 19.3944
R14329 gnd.n6381 gnd.n404 19.3944
R14330 gnd.n6387 gnd.n404 19.3944
R14331 gnd.n6387 gnd.n402 19.3944
R14332 gnd.n6391 gnd.n402 19.3944
R14333 gnd.n6391 gnd.n398 19.3944
R14334 gnd.n6397 gnd.n398 19.3944
R14335 gnd.n6397 gnd.n396 19.3944
R14336 gnd.n6401 gnd.n396 19.3944
R14337 gnd.n6401 gnd.n392 19.3944
R14338 gnd.n6407 gnd.n392 19.3944
R14339 gnd.n6407 gnd.n390 19.3944
R14340 gnd.n6412 gnd.n390 19.3944
R14341 gnd.n6412 gnd.n386 19.3944
R14342 gnd.n6418 gnd.n386 19.3944
R14343 gnd.n6419 gnd.n6418 19.3944
R14344 gnd.n3792 gnd.n3789 19.3944
R14345 gnd.n3792 gnd.n3788 19.3944
R14346 gnd.n3798 gnd.n3788 19.3944
R14347 gnd.n3798 gnd.n3786 19.3944
R14348 gnd.n3802 gnd.n3786 19.3944
R14349 gnd.n3802 gnd.n3784 19.3944
R14350 gnd.n3808 gnd.n3784 19.3944
R14351 gnd.n3808 gnd.n3782 19.3944
R14352 gnd.n3812 gnd.n3782 19.3944
R14353 gnd.n3812 gnd.n3780 19.3944
R14354 gnd.n3818 gnd.n3780 19.3944
R14355 gnd.n3818 gnd.n3778 19.3944
R14356 gnd.n3823 gnd.n3778 19.3944
R14357 gnd.n3823 gnd.n3776 19.3944
R14358 gnd.n3776 gnd.n1360 19.3944
R14359 gnd.n3836 gnd.n1358 19.3944
R14360 gnd.n3836 gnd.n1356 19.3944
R14361 gnd.n3842 gnd.n1356 19.3944
R14362 gnd.n3842 gnd.n1354 19.3944
R14363 gnd.n3846 gnd.n1354 19.3944
R14364 gnd.n3846 gnd.n1352 19.3944
R14365 gnd.n3852 gnd.n1352 19.3944
R14366 gnd.n3852 gnd.n1350 19.3944
R14367 gnd.n3856 gnd.n1350 19.3944
R14368 gnd.n3856 gnd.n1348 19.3944
R14369 gnd.n3862 gnd.n1348 19.3944
R14370 gnd.n3862 gnd.n1346 19.3944
R14371 gnd.n3866 gnd.n1346 19.3944
R14372 gnd.n3866 gnd.n1344 19.3944
R14373 gnd.n3872 gnd.n1344 19.3944
R14374 gnd.n3872 gnd.n1342 19.3944
R14375 gnd.n3877 gnd.n1342 19.3944
R14376 gnd.n3877 gnd.n1340 19.3944
R14377 gnd.n3888 gnd.n1335 19.3944
R14378 gnd.n3888 gnd.n1330 19.3944
R14379 gnd.n3901 gnd.n1330 19.3944
R14380 gnd.n3901 gnd.n1328 19.3944
R14381 gnd.n3990 gnd.n1328 19.3944
R14382 gnd.n3990 gnd.n3989 19.3944
R14383 gnd.n3989 gnd.n3988 19.3944
R14384 gnd.n3988 gnd.n3986 19.3944
R14385 gnd.n3986 gnd.n3985 19.3944
R14386 gnd.n3985 gnd.n3984 19.3944
R14387 gnd.n3984 gnd.n3982 19.3944
R14388 gnd.n3982 gnd.n3981 19.3944
R14389 gnd.n3981 gnd.n3979 19.3944
R14390 gnd.n3979 gnd.n3978 19.3944
R14391 gnd.n3978 gnd.n3977 19.3944
R14392 gnd.n3977 gnd.n3975 19.3944
R14393 gnd.n3975 gnd.n3974 19.3944
R14394 gnd.n3974 gnd.n3971 19.3944
R14395 gnd.n3971 gnd.n3970 19.3944
R14396 gnd.n3970 gnd.n3969 19.3944
R14397 gnd.n3969 gnd.n3968 19.3944
R14398 gnd.n3968 gnd.n3964 19.3944
R14399 gnd.n3964 gnd.n3963 19.3944
R14400 gnd.n3963 gnd.n3961 19.3944
R14401 gnd.n3961 gnd.n3960 19.3944
R14402 gnd.n3960 gnd.n3958 19.3944
R14403 gnd.n3958 gnd.n3957 19.3944
R14404 gnd.n3957 gnd.n3955 19.3944
R14405 gnd.n3955 gnd.n3954 19.3944
R14406 gnd.n3954 gnd.n3952 19.3944
R14407 gnd.n3952 gnd.n3951 19.3944
R14408 gnd.n3951 gnd.n3949 19.3944
R14409 gnd.n3949 gnd.n3948 19.3944
R14410 gnd.n3948 gnd.n3946 19.3944
R14411 gnd.n3946 gnd.n3945 19.3944
R14412 gnd.n3945 gnd.n3943 19.3944
R14413 gnd.n3943 gnd.n3942 19.3944
R14414 gnd.n3942 gnd.n3940 19.3944
R14415 gnd.n3940 gnd.n3939 19.3944
R14416 gnd.n3939 gnd.n159 19.3944
R14417 gnd.n6804 gnd.n159 19.3944
R14418 gnd.n6805 gnd.n6804 19.3944
R14419 gnd.n6843 gnd.n120 19.3944
R14420 gnd.n6838 gnd.n120 19.3944
R14421 gnd.n6838 gnd.n6837 19.3944
R14422 gnd.n6837 gnd.n6836 19.3944
R14423 gnd.n6836 gnd.n127 19.3944
R14424 gnd.n6831 gnd.n127 19.3944
R14425 gnd.n6831 gnd.n6830 19.3944
R14426 gnd.n6830 gnd.n6829 19.3944
R14427 gnd.n6829 gnd.n134 19.3944
R14428 gnd.n6824 gnd.n134 19.3944
R14429 gnd.n6824 gnd.n6823 19.3944
R14430 gnd.n6823 gnd.n6822 19.3944
R14431 gnd.n6822 gnd.n141 19.3944
R14432 gnd.n6817 gnd.n141 19.3944
R14433 gnd.n6817 gnd.n6816 19.3944
R14434 gnd.n6816 gnd.n6815 19.3944
R14435 gnd.n6815 gnd.n148 19.3944
R14436 gnd.n6810 gnd.n148 19.3944
R14437 gnd.n6876 gnd.n6875 19.3944
R14438 gnd.n6875 gnd.n6874 19.3944
R14439 gnd.n6874 gnd.n92 19.3944
R14440 gnd.n6869 gnd.n92 19.3944
R14441 gnd.n6869 gnd.n6868 19.3944
R14442 gnd.n6868 gnd.n6867 19.3944
R14443 gnd.n6867 gnd.n99 19.3944
R14444 gnd.n6862 gnd.n99 19.3944
R14445 gnd.n6862 gnd.n6861 19.3944
R14446 gnd.n6861 gnd.n6860 19.3944
R14447 gnd.n6860 gnd.n106 19.3944
R14448 gnd.n6855 gnd.n106 19.3944
R14449 gnd.n6855 gnd.n6854 19.3944
R14450 gnd.n6854 gnd.n6853 19.3944
R14451 gnd.n6853 gnd.n113 19.3944
R14452 gnd.n6848 gnd.n113 19.3944
R14453 gnd.n6848 gnd.n6847 19.3944
R14454 gnd.n4128 gnd.n4127 19.3944
R14455 gnd.n4127 gnd.n4126 19.3944
R14456 gnd.n4126 gnd.n1222 19.3944
R14457 gnd.n4012 gnd.n1222 19.3944
R14458 gnd.n4012 gnd.n1323 19.3944
R14459 gnd.n4018 gnd.n1323 19.3944
R14460 gnd.n4018 gnd.n4017 19.3944
R14461 gnd.n4017 gnd.n1297 19.3944
R14462 gnd.n4043 gnd.n1297 19.3944
R14463 gnd.n4043 gnd.n1295 19.3944
R14464 gnd.n4050 gnd.n1295 19.3944
R14465 gnd.n4050 gnd.n4049 19.3944
R14466 gnd.n4049 gnd.n1267 19.3944
R14467 gnd.n4082 gnd.n1267 19.3944
R14468 gnd.n4083 gnd.n4082 19.3944
R14469 gnd.n4084 gnd.n4083 19.3944
R14470 gnd.n1265 gnd.n1264 19.3944
R14471 gnd.n6647 gnd.n6646 19.3944
R14472 gnd.n235 gnd.n234 19.3944
R14473 gnd.n6661 gnd.n6660 19.3944
R14474 gnd.n6673 gnd.n219 19.3944
R14475 gnd.n6673 gnd.n211 19.3944
R14476 gnd.n6677 gnd.n211 19.3944
R14477 gnd.n6677 gnd.n199 19.3944
R14478 gnd.n6689 gnd.n199 19.3944
R14479 gnd.n6689 gnd.n197 19.3944
R14480 gnd.n6693 gnd.n197 19.3944
R14481 gnd.n6693 gnd.n183 19.3944
R14482 gnd.n6705 gnd.n183 19.3944
R14483 gnd.n6705 gnd.n181 19.3944
R14484 gnd.n6709 gnd.n181 19.3944
R14485 gnd.n6709 gnd.n167 19.3944
R14486 gnd.n6795 gnd.n167 19.3944
R14487 gnd.n6795 gnd.n165 19.3944
R14488 gnd.n6799 gnd.n165 19.3944
R14489 gnd.n6799 gnd.n87 19.3944
R14490 gnd.n6879 gnd.n87 19.3944
R14491 gnd.n4479 gnd.n4478 19.3944
R14492 gnd.n4478 gnd.n4477 19.3944
R14493 gnd.n4477 gnd.n4476 19.3944
R14494 gnd.n4476 gnd.n4474 19.3944
R14495 gnd.n4474 gnd.n4471 19.3944
R14496 gnd.n4471 gnd.n4470 19.3944
R14497 gnd.n4470 gnd.n4467 19.3944
R14498 gnd.n4467 gnd.n4466 19.3944
R14499 gnd.n4466 gnd.n4463 19.3944
R14500 gnd.n4463 gnd.n4462 19.3944
R14501 gnd.n4462 gnd.n4459 19.3944
R14502 gnd.n4459 gnd.n4458 19.3944
R14503 gnd.n4458 gnd.n4455 19.3944
R14504 gnd.n4455 gnd.n4454 19.3944
R14505 gnd.n4454 gnd.n4451 19.3944
R14506 gnd.n4451 gnd.n4450 19.3944
R14507 gnd.n4450 gnd.n4447 19.3944
R14508 gnd.n4445 gnd.n4442 19.3944
R14509 gnd.n4442 gnd.n4441 19.3944
R14510 gnd.n4441 gnd.n4438 19.3944
R14511 gnd.n4438 gnd.n4437 19.3944
R14512 gnd.n4437 gnd.n4434 19.3944
R14513 gnd.n4434 gnd.n4433 19.3944
R14514 gnd.n4433 gnd.n4430 19.3944
R14515 gnd.n4430 gnd.n4429 19.3944
R14516 gnd.n4429 gnd.n4426 19.3944
R14517 gnd.n4426 gnd.n4425 19.3944
R14518 gnd.n4425 gnd.n4422 19.3944
R14519 gnd.n4422 gnd.n4421 19.3944
R14520 gnd.n4421 gnd.n4418 19.3944
R14521 gnd.n4418 gnd.n4417 19.3944
R14522 gnd.n4417 gnd.n4414 19.3944
R14523 gnd.n4414 gnd.n4413 19.3944
R14524 gnd.n4413 gnd.n4410 19.3944
R14525 gnd.n4410 gnd.n4409 19.3944
R14526 gnd.n2343 gnd.n2274 19.3944
R14527 gnd.n2343 gnd.n2275 19.3944
R14528 gnd.n2339 gnd.n2275 19.3944
R14529 gnd.n2339 gnd.n901 19.3944
R14530 gnd.n4387 gnd.n901 19.3944
R14531 gnd.n4387 gnd.n4386 19.3944
R14532 gnd.n4386 gnd.n4385 19.3944
R14533 gnd.n4385 gnd.n905 19.3944
R14534 gnd.n4375 gnd.n905 19.3944
R14535 gnd.n4375 gnd.n4374 19.3944
R14536 gnd.n4374 gnd.n4373 19.3944
R14537 gnd.n4373 gnd.n924 19.3944
R14538 gnd.n4363 gnd.n924 19.3944
R14539 gnd.n4363 gnd.n4362 19.3944
R14540 gnd.n4362 gnd.n4361 19.3944
R14541 gnd.n4361 gnd.n945 19.3944
R14542 gnd.n963 gnd.n945 19.3944
R14543 gnd.n4349 gnd.n963 19.3944
R14544 gnd.n4349 gnd.n4348 19.3944
R14545 gnd.n4348 gnd.n4347 19.3944
R14546 gnd.n4347 gnd.n969 19.3944
R14547 gnd.n4336 gnd.n969 19.3944
R14548 gnd.n4336 gnd.n4335 19.3944
R14549 gnd.n4335 gnd.n4334 19.3944
R14550 gnd.n4334 gnd.n985 19.3944
R14551 gnd.n4323 gnd.n985 19.3944
R14552 gnd.n4323 gnd.n4322 19.3944
R14553 gnd.n4322 gnd.n4321 19.3944
R14554 gnd.n4321 gnd.n1004 19.3944
R14555 gnd.n4311 gnd.n1004 19.3944
R14556 gnd.n4311 gnd.n4310 19.3944
R14557 gnd.n4310 gnd.n4309 19.3944
R14558 gnd.n4309 gnd.n1024 19.3944
R14559 gnd.n4299 gnd.n1024 19.3944
R14560 gnd.n4299 gnd.n4298 19.3944
R14561 gnd.n4298 gnd.n4297 19.3944
R14562 gnd.n4297 gnd.n1046 19.3944
R14563 gnd.n4287 gnd.n1046 19.3944
R14564 gnd.n4287 gnd.n4286 19.3944
R14565 gnd.n4286 gnd.n4285 19.3944
R14566 gnd.n4285 gnd.n1067 19.3944
R14567 gnd.n4275 gnd.n1067 19.3944
R14568 gnd.n2335 gnd.n2333 19.3944
R14569 gnd.n2333 gnd.n2330 19.3944
R14570 gnd.n2330 gnd.n2329 19.3944
R14571 gnd.n2329 gnd.n2326 19.3944
R14572 gnd.n2326 gnd.n2325 19.3944
R14573 gnd.n2325 gnd.n2322 19.3944
R14574 gnd.n2322 gnd.n2321 19.3944
R14575 gnd.n2321 gnd.n2318 19.3944
R14576 gnd.n2318 gnd.n2317 19.3944
R14577 gnd.n2317 gnd.n2314 19.3944
R14578 gnd.n2314 gnd.n2313 19.3944
R14579 gnd.n2313 gnd.n2310 19.3944
R14580 gnd.n2310 gnd.n2309 19.3944
R14581 gnd.n2309 gnd.n2306 19.3944
R14582 gnd.n2306 gnd.n2305 19.3944
R14583 gnd.n2305 gnd.n2302 19.3944
R14584 gnd.n2296 gnd.n2270 19.3944
R14585 gnd.n2354 gnd.n2270 19.3944
R14586 gnd.n2355 gnd.n2354 19.3944
R14587 gnd.n2355 gnd.n2268 19.3944
R14588 gnd.n2359 gnd.n2268 19.3944
R14589 gnd.n2361 gnd.n2359 19.3944
R14590 gnd.n2362 gnd.n2361 19.3944
R14591 gnd.n2362 gnd.n2265 19.3944
R14592 gnd.n2366 gnd.n2265 19.3944
R14593 gnd.n2368 gnd.n2366 19.3944
R14594 gnd.n2369 gnd.n2368 19.3944
R14595 gnd.n2369 gnd.n2262 19.3944
R14596 gnd.n2373 gnd.n2262 19.3944
R14597 gnd.n2375 gnd.n2373 19.3944
R14598 gnd.n2376 gnd.n2375 19.3944
R14599 gnd.n2376 gnd.n2259 19.3944
R14600 gnd.n2422 gnd.n2259 19.3944
R14601 gnd.n2423 gnd.n2422 19.3944
R14602 gnd.n2425 gnd.n2423 19.3944
R14603 gnd.n2425 gnd.n2257 19.3944
R14604 gnd.n2429 gnd.n2257 19.3944
R14605 gnd.n2429 gnd.n2249 19.3944
R14606 gnd.n2451 gnd.n2249 19.3944
R14607 gnd.n2451 gnd.n2250 19.3944
R14608 gnd.n2447 gnd.n2250 19.3944
R14609 gnd.n2447 gnd.n2241 19.3944
R14610 gnd.n2504 gnd.n2241 19.3944
R14611 gnd.n2504 gnd.n2239 19.3944
R14612 gnd.n2508 gnd.n2239 19.3944
R14613 gnd.n2508 gnd.n2234 19.3944
R14614 gnd.n2520 gnd.n2234 19.3944
R14615 gnd.n2520 gnd.n2232 19.3944
R14616 gnd.n2524 gnd.n2232 19.3944
R14617 gnd.n2524 gnd.n2222 19.3944
R14618 gnd.n2552 gnd.n2222 19.3944
R14619 gnd.n2552 gnd.n2223 19.3944
R14620 gnd.n2548 gnd.n2223 19.3944
R14621 gnd.n2548 gnd.n2547 19.3944
R14622 gnd.n2547 gnd.n2546 19.3944
R14623 gnd.n2546 gnd.n2031 19.3944
R14624 gnd.n2660 gnd.n2031 19.3944
R14625 gnd.n2660 gnd.n2032 19.3944
R14626 gnd.n4402 gnd.n4401 19.3944
R14627 gnd.n4401 gnd.n879 19.3944
R14628 gnd.n4397 gnd.n879 19.3944
R14629 gnd.n4397 gnd.n881 19.3944
R14630 gnd.n2391 gnd.n881 19.3944
R14631 gnd.n2393 gnd.n2391 19.3944
R14632 gnd.n2394 gnd.n2393 19.3944
R14633 gnd.n2394 gnd.n2388 19.3944
R14634 gnd.n2398 gnd.n2388 19.3944
R14635 gnd.n2400 gnd.n2398 19.3944
R14636 gnd.n2401 gnd.n2400 19.3944
R14637 gnd.n2401 gnd.n2385 19.3944
R14638 gnd.n2405 gnd.n2385 19.3944
R14639 gnd.n2407 gnd.n2405 19.3944
R14640 gnd.n2408 gnd.n2407 19.3944
R14641 gnd.n2408 gnd.n2382 19.3944
R14642 gnd.n2418 gnd.n2382 19.3944
R14643 gnd.n2418 gnd.n2417 19.3944
R14644 gnd.n2417 gnd.n2416 19.3944
R14645 gnd.n2416 gnd.n2254 19.3944
R14646 gnd.n2433 gnd.n2254 19.3944
R14647 gnd.n2434 gnd.n2433 19.3944
R14648 gnd.n2435 gnd.n2434 19.3944
R14649 gnd.n2435 gnd.n2252 19.3944
R14650 gnd.n2443 gnd.n2252 19.3944
R14651 gnd.n2443 gnd.n2442 19.3944
R14652 gnd.n2442 gnd.n2441 19.3944
R14653 gnd.n2441 gnd.n2238 19.3944
R14654 gnd.n2512 gnd.n2238 19.3944
R14655 gnd.n2512 gnd.n2236 19.3944
R14656 gnd.n2516 gnd.n2236 19.3944
R14657 gnd.n2516 gnd.n2231 19.3944
R14658 gnd.n2528 gnd.n2231 19.3944
R14659 gnd.n2528 gnd.n2229 19.3944
R14660 gnd.n2532 gnd.n2229 19.3944
R14661 gnd.n2533 gnd.n2532 19.3944
R14662 gnd.n2536 gnd.n2533 19.3944
R14663 gnd.n2536 gnd.n2227 19.3944
R14664 gnd.n2541 gnd.n2227 19.3944
R14665 gnd.n2541 gnd.n2030 19.3944
R14666 gnd.n2664 gnd.n2030 19.3944
R14667 gnd.n2665 gnd.n2664 19.3944
R14668 gnd.n2703 gnd.n1933 19.3944
R14669 gnd.n2703 gnd.n1940 19.3944
R14670 gnd.n1997 gnd.n1940 19.3944
R14671 gnd.n2696 gnd.n1997 19.3944
R14672 gnd.n2696 gnd.n2695 19.3944
R14673 gnd.n2695 gnd.n2694 19.3944
R14674 gnd.n2694 gnd.n2003 19.3944
R14675 gnd.n2689 gnd.n2003 19.3944
R14676 gnd.n2689 gnd.n2688 19.3944
R14677 gnd.n2688 gnd.n2687 19.3944
R14678 gnd.n2687 gnd.n2010 19.3944
R14679 gnd.n2682 gnd.n2010 19.3944
R14680 gnd.n2682 gnd.n2681 19.3944
R14681 gnd.n2681 gnd.n2680 19.3944
R14682 gnd.n2680 gnd.n2017 19.3944
R14683 gnd.n2675 gnd.n2017 19.3944
R14684 gnd.n2675 gnd.n2674 19.3944
R14685 gnd.n2674 gnd.n2673 19.3944
R14686 gnd.n1953 gnd.n1952 19.3944
R14687 gnd.n1993 gnd.n1952 19.3944
R14688 gnd.n1993 gnd.n1992 19.3944
R14689 gnd.n1992 gnd.n1991 19.3944
R14690 gnd.n1991 gnd.n1988 19.3944
R14691 gnd.n1988 gnd.n1987 19.3944
R14692 gnd.n1987 gnd.n1984 19.3944
R14693 gnd.n1984 gnd.n1983 19.3944
R14694 gnd.n1983 gnd.n1980 19.3944
R14695 gnd.n1980 gnd.n1979 19.3944
R14696 gnd.n1979 gnd.n1976 19.3944
R14697 gnd.n1976 gnd.n1975 19.3944
R14698 gnd.n1975 gnd.n1972 19.3944
R14699 gnd.n1972 gnd.n1971 19.3944
R14700 gnd.n1971 gnd.n1934 19.3944
R14701 gnd.n2349 gnd.n2345 19.3944
R14702 gnd.n2349 gnd.n890 19.3944
R14703 gnd.n4393 gnd.n890 19.3944
R14704 gnd.n4393 gnd.n4392 19.3944
R14705 gnd.n4392 gnd.n4391 19.3944
R14706 gnd.n4391 gnd.n894 19.3944
R14707 gnd.n4381 gnd.n894 19.3944
R14708 gnd.n4381 gnd.n4380 19.3944
R14709 gnd.n4380 gnd.n4379 19.3944
R14710 gnd.n4379 gnd.n915 19.3944
R14711 gnd.n4369 gnd.n915 19.3944
R14712 gnd.n4369 gnd.n4368 19.3944
R14713 gnd.n4368 gnd.n4367 19.3944
R14714 gnd.n4367 gnd.n934 19.3944
R14715 gnd.n4357 gnd.n934 19.3944
R14716 gnd.n4357 gnd.n4356 19.3944
R14717 gnd.n4354 gnd.n4353 19.3944
R14718 gnd.n4343 gnd.n975 19.3944
R14719 gnd.n4341 gnd.n4340 19.3944
R14720 gnd.n4330 gnd.n992 19.3944
R14721 gnd.n4328 gnd.n4327 19.3944
R14722 gnd.n4327 gnd.n993 19.3944
R14723 gnd.n4317 gnd.n993 19.3944
R14724 gnd.n4317 gnd.n4316 19.3944
R14725 gnd.n4316 gnd.n4315 19.3944
R14726 gnd.n4315 gnd.n1014 19.3944
R14727 gnd.n4305 gnd.n1014 19.3944
R14728 gnd.n4305 gnd.n4304 19.3944
R14729 gnd.n4304 gnd.n4303 19.3944
R14730 gnd.n4303 gnd.n1035 19.3944
R14731 gnd.n4293 gnd.n1035 19.3944
R14732 gnd.n4293 gnd.n4292 19.3944
R14733 gnd.n4292 gnd.n4291 19.3944
R14734 gnd.n4291 gnd.n1056 19.3944
R14735 gnd.n4281 gnd.n1056 19.3944
R14736 gnd.n4281 gnd.n4280 19.3944
R14737 gnd.n4280 gnd.n4279 19.3944
R14738 gnd.n6061 gnd.n599 19.3944
R14739 gnd.n6061 gnd.n6060 19.3944
R14740 gnd.n6060 gnd.n6059 19.3944
R14741 gnd.n6059 gnd.n603 19.3944
R14742 gnd.n6053 gnd.n603 19.3944
R14743 gnd.n6053 gnd.n6052 19.3944
R14744 gnd.n6052 gnd.n6051 19.3944
R14745 gnd.n6051 gnd.n611 19.3944
R14746 gnd.n6045 gnd.n611 19.3944
R14747 gnd.n6045 gnd.n6044 19.3944
R14748 gnd.n6044 gnd.n6043 19.3944
R14749 gnd.n6043 gnd.n619 19.3944
R14750 gnd.n6037 gnd.n619 19.3944
R14751 gnd.n6037 gnd.n6036 19.3944
R14752 gnd.n6036 gnd.n6035 19.3944
R14753 gnd.n6035 gnd.n627 19.3944
R14754 gnd.n6029 gnd.n627 19.3944
R14755 gnd.n6029 gnd.n6028 19.3944
R14756 gnd.n6028 gnd.n6027 19.3944
R14757 gnd.n6027 gnd.n635 19.3944
R14758 gnd.n6021 gnd.n635 19.3944
R14759 gnd.n6021 gnd.n6020 19.3944
R14760 gnd.n6020 gnd.n6019 19.3944
R14761 gnd.n6019 gnd.n643 19.3944
R14762 gnd.n6013 gnd.n643 19.3944
R14763 gnd.n6013 gnd.n6012 19.3944
R14764 gnd.n6012 gnd.n6011 19.3944
R14765 gnd.n6011 gnd.n651 19.3944
R14766 gnd.n6005 gnd.n651 19.3944
R14767 gnd.n6005 gnd.n6004 19.3944
R14768 gnd.n6004 gnd.n6003 19.3944
R14769 gnd.n6003 gnd.n659 19.3944
R14770 gnd.n5997 gnd.n659 19.3944
R14771 gnd.n5997 gnd.n5996 19.3944
R14772 gnd.n5996 gnd.n5995 19.3944
R14773 gnd.n5995 gnd.n667 19.3944
R14774 gnd.n5989 gnd.n667 19.3944
R14775 gnd.n5989 gnd.n5988 19.3944
R14776 gnd.n5988 gnd.n5987 19.3944
R14777 gnd.n5987 gnd.n675 19.3944
R14778 gnd.n5981 gnd.n675 19.3944
R14779 gnd.n5981 gnd.n5980 19.3944
R14780 gnd.n5980 gnd.n5979 19.3944
R14781 gnd.n5979 gnd.n683 19.3944
R14782 gnd.n5973 gnd.n683 19.3944
R14783 gnd.n5973 gnd.n5972 19.3944
R14784 gnd.n5972 gnd.n5971 19.3944
R14785 gnd.n5971 gnd.n691 19.3944
R14786 gnd.n5965 gnd.n691 19.3944
R14787 gnd.n5965 gnd.n5964 19.3944
R14788 gnd.n5964 gnd.n5963 19.3944
R14789 gnd.n5963 gnd.n699 19.3944
R14790 gnd.n5957 gnd.n699 19.3944
R14791 gnd.n5957 gnd.n5956 19.3944
R14792 gnd.n5956 gnd.n5955 19.3944
R14793 gnd.n5955 gnd.n707 19.3944
R14794 gnd.n5949 gnd.n707 19.3944
R14795 gnd.n5949 gnd.n5948 19.3944
R14796 gnd.n5948 gnd.n5947 19.3944
R14797 gnd.n5947 gnd.n715 19.3944
R14798 gnd.n5941 gnd.n715 19.3944
R14799 gnd.n5941 gnd.n5940 19.3944
R14800 gnd.n5940 gnd.n5939 19.3944
R14801 gnd.n5939 gnd.n723 19.3944
R14802 gnd.n5933 gnd.n723 19.3944
R14803 gnd.n5933 gnd.n5932 19.3944
R14804 gnd.n5932 gnd.n5931 19.3944
R14805 gnd.n5931 gnd.n731 19.3944
R14806 gnd.n5925 gnd.n731 19.3944
R14807 gnd.n5925 gnd.n5924 19.3944
R14808 gnd.n5924 gnd.n5923 19.3944
R14809 gnd.n5923 gnd.n739 19.3944
R14810 gnd.n5917 gnd.n739 19.3944
R14811 gnd.n5917 gnd.n5916 19.3944
R14812 gnd.n5916 gnd.n5915 19.3944
R14813 gnd.n5915 gnd.n747 19.3944
R14814 gnd.n5909 gnd.n747 19.3944
R14815 gnd.n5909 gnd.n5908 19.3944
R14816 gnd.n5908 gnd.n5907 19.3944
R14817 gnd.n5907 gnd.n755 19.3944
R14818 gnd.n5901 gnd.n755 19.3944
R14819 gnd.n5901 gnd.n5900 19.3944
R14820 gnd.n5900 gnd.n5899 19.3944
R14821 gnd.n5899 gnd.n763 19.3944
R14822 gnd.n4270 gnd.n4269 19.3944
R14823 gnd.n4269 gnd.n4268 19.3944
R14824 gnd.n4268 gnd.n1091 19.3944
R14825 gnd.n4264 gnd.n1091 19.3944
R14826 gnd.n4264 gnd.n4263 19.3944
R14827 gnd.n4263 gnd.n4262 19.3944
R14828 gnd.n4262 gnd.n1096 19.3944
R14829 gnd.n4258 gnd.n1096 19.3944
R14830 gnd.n4258 gnd.n4257 19.3944
R14831 gnd.n4257 gnd.n4256 19.3944
R14832 gnd.n4256 gnd.n1101 19.3944
R14833 gnd.n4252 gnd.n1101 19.3944
R14834 gnd.n4252 gnd.n4251 19.3944
R14835 gnd.n4251 gnd.n4250 19.3944
R14836 gnd.n4250 gnd.n1106 19.3944
R14837 gnd.n4246 gnd.n1106 19.3944
R14838 gnd.n4246 gnd.n4245 19.3944
R14839 gnd.n4245 gnd.n4244 19.3944
R14840 gnd.n4244 gnd.n1111 19.3944
R14841 gnd.n4240 gnd.n1111 19.3944
R14842 gnd.n4240 gnd.n4239 19.3944
R14843 gnd.n4239 gnd.n4238 19.3944
R14844 gnd.n4238 gnd.n1116 19.3944
R14845 gnd.n4234 gnd.n1116 19.3944
R14846 gnd.n4234 gnd.n4233 19.3944
R14847 gnd.n4233 gnd.n4232 19.3944
R14848 gnd.n4232 gnd.n1121 19.3944
R14849 gnd.n4228 gnd.n1121 19.3944
R14850 gnd.n4228 gnd.n4227 19.3944
R14851 gnd.n4227 gnd.n4226 19.3944
R14852 gnd.n4226 gnd.n1126 19.3944
R14853 gnd.n4222 gnd.n1126 19.3944
R14854 gnd.n4222 gnd.n4221 19.3944
R14855 gnd.n4221 gnd.n4220 19.3944
R14856 gnd.n4220 gnd.n1131 19.3944
R14857 gnd.n4216 gnd.n1131 19.3944
R14858 gnd.n4216 gnd.n4215 19.3944
R14859 gnd.n4215 gnd.n4214 19.3944
R14860 gnd.n4214 gnd.n1136 19.3944
R14861 gnd.n4210 gnd.n1136 19.3944
R14862 gnd.n4210 gnd.n4209 19.3944
R14863 gnd.n4209 gnd.n4208 19.3944
R14864 gnd.n4208 gnd.n1141 19.3944
R14865 gnd.n4204 gnd.n1141 19.3944
R14866 gnd.n4204 gnd.n4203 19.3944
R14867 gnd.n4203 gnd.n4202 19.3944
R14868 gnd.n4202 gnd.n1146 19.3944
R14869 gnd.n4198 gnd.n1146 19.3944
R14870 gnd.n4198 gnd.n4197 19.3944
R14871 gnd.n4197 gnd.n4196 19.3944
R14872 gnd.n4196 gnd.n1151 19.3944
R14873 gnd.n4192 gnd.n1151 19.3944
R14874 gnd.n4192 gnd.n4191 19.3944
R14875 gnd.n4191 gnd.n4190 19.3944
R14876 gnd.n4190 gnd.n1156 19.3944
R14877 gnd.n4186 gnd.n1156 19.3944
R14878 gnd.n4186 gnd.n4185 19.3944
R14879 gnd.n4185 gnd.n4184 19.3944
R14880 gnd.n4184 gnd.n1161 19.3944
R14881 gnd.n4180 gnd.n1161 19.3944
R14882 gnd.n4180 gnd.n4179 19.3944
R14883 gnd.n4179 gnd.n4178 19.3944
R14884 gnd.n4178 gnd.n1166 19.3944
R14885 gnd.n4174 gnd.n1166 19.3944
R14886 gnd.n4174 gnd.n4173 19.3944
R14887 gnd.n4173 gnd.n4172 19.3944
R14888 gnd.n4172 gnd.n1171 19.3944
R14889 gnd.n4168 gnd.n1171 19.3944
R14890 gnd.n4168 gnd.n4167 19.3944
R14891 gnd.n4167 gnd.n4166 19.3944
R14892 gnd.n4166 gnd.n1176 19.3944
R14893 gnd.n4162 gnd.n1176 19.3944
R14894 gnd.n4162 gnd.n4161 19.3944
R14895 gnd.n4161 gnd.n4160 19.3944
R14896 gnd.n4160 gnd.n1181 19.3944
R14897 gnd.n4156 gnd.n1181 19.3944
R14898 gnd.n4156 gnd.n4155 19.3944
R14899 gnd.n4155 gnd.n4154 19.3944
R14900 gnd.n4154 gnd.n1186 19.3944
R14901 gnd.n4150 gnd.n1186 19.3944
R14902 gnd.n4150 gnd.n4149 19.3944
R14903 gnd.n4149 gnd.n4148 19.3944
R14904 gnd.n3581 gnd.n3416 19.3944
R14905 gnd.n3581 gnd.n3414 19.3944
R14906 gnd.n3586 gnd.n3414 19.3944
R14907 gnd.n3480 gnd.n3462 19.3944
R14908 gnd.n3480 gnd.n3460 19.3944
R14909 gnd.n3486 gnd.n3460 19.3944
R14910 gnd.n3486 gnd.n3453 19.3944
R14911 gnd.n3499 gnd.n3453 19.3944
R14912 gnd.n3499 gnd.n3451 19.3944
R14913 gnd.n3505 gnd.n3451 19.3944
R14914 gnd.n3505 gnd.n3444 19.3944
R14915 gnd.n3518 gnd.n3444 19.3944
R14916 gnd.n3518 gnd.n3442 19.3944
R14917 gnd.n3524 gnd.n3442 19.3944
R14918 gnd.n3524 gnd.n3435 19.3944
R14919 gnd.n3537 gnd.n3435 19.3944
R14920 gnd.n3537 gnd.n3433 19.3944
R14921 gnd.n3545 gnd.n3433 19.3944
R14922 gnd.n3545 gnd.n3544 19.3944
R14923 gnd.n3544 gnd.n3424 19.3944
R14924 gnd.n3558 gnd.n3424 19.3944
R14925 gnd.n3558 gnd.n3422 19.3944
R14926 gnd.n3564 gnd.n3422 19.3944
R14927 gnd.n3564 gnd.n3420 19.3944
R14928 gnd.n3568 gnd.n3420 19.3944
R14929 gnd.n3568 gnd.n3418 19.3944
R14930 gnd.n3577 gnd.n3418 19.3944
R14931 gnd.n2776 gnd.n2775 19.2005
R14932 gnd.n3702 gnd.n3701 19.2005
R14933 gnd.t97 gnd.n4710 18.8012
R14934 gnd.n5302 gnd.t252 18.8012
R14935 gnd.n5147 gnd.n5146 18.4825
R14936 gnd.n3832 gnd.n1360 18.4247
R14937 gnd.n2707 gnd.n1934 18.4247
R14938 gnd.n6758 gnd.n6757 18.2308
R14939 gnd.n3548 gnd.n3428 18.2308
R14940 gnd.n2166 gnd.n2150 18.2308
R14941 gnd.n2302 gnd.n2294 18.2308
R14942 gnd.t99 gnd.n4754 18.1639
R14943 gnd.n5896 gnd.n5895 17.8452
R14944 gnd.n4781 gnd.t100 17.5266
R14945 gnd.n4739 gnd.t94 16.8893
R14946 gnd.n2351 gnd.t191 16.8893
R14947 gnd.n2662 gnd.t134 16.8893
R14948 gnd.n3890 gnd.t123 16.8893
R14949 gnd.t119 gnd.n81 16.8893
R14950 gnd.n5008 gnd.t213 16.2519
R14951 gnd.n5292 gnd.t88 16.2519
R14952 gnd.n2576 gnd.n2206 15.9333
R14953 gnd.n2585 gnd.n2206 15.9333
R14954 gnd.n2587 gnd.n2586 15.9333
R14955 gnd.n2590 gnd.n2587 15.9333
R14956 gnd.n2590 gnd.n2589 15.9333
R14957 gnd.n2589 gnd.n2588 15.9333
R14958 gnd.n2598 gnd.n2068 15.9333
R14959 gnd.n2601 gnd.n2598 15.9333
R14960 gnd.n2602 gnd.n2601 15.9333
R14961 gnd.n2603 gnd.n2602 15.9333
R14962 gnd.n2605 gnd.n2603 15.9333
R14963 gnd.n2605 gnd.n2604 15.9333
R14964 gnd.n2604 gnd.n2061 15.9333
R14965 gnd.n2624 gnd.n2061 15.9333
R14966 gnd.n2623 gnd.n1816 15.9333
R14967 gnd.n2616 gnd.n1849 15.9333
R14968 gnd.n1862 gnd.n1791 15.9333
R14969 gnd.n2808 gnd.n1751 15.9333
R14970 gnd.n2851 gnd.n1740 15.9333
R14971 gnd.n2885 gnd.n1729 15.9333
R14972 gnd.n2896 gnd.n2895 15.9333
R14973 gnd.n2925 gnd.n1708 15.9333
R14974 gnd.n3015 gnd.n1658 15.9333
R14975 gnd.n3034 gnd.n1635 15.9333
R14976 gnd.n1642 gnd.n1630 15.9333
R14977 gnd.n3074 gnd.n1613 15.9333
R14978 gnd.n3121 gnd.n3120 15.9333
R14979 gnd.n3129 gnd.n1600 15.9333
R14980 gnd.n3146 gnd.n3145 15.9333
R14981 gnd.n3206 gnd.n1568 15.9333
R14982 gnd.n3288 gnd.n3287 15.9333
R14983 gnd.n3296 gnd.n1511 15.9333
R14984 gnd.n3315 gnd.n3314 15.9333
R14985 gnd.n3325 gnd.n1484 15.9333
R14986 gnd.n3347 gnd.n1479 15.9333
R14987 gnd.n3613 gnd.n3612 15.9333
R14988 gnd.n3399 gnd.n1402 15.9333
R14989 gnd.n3399 gnd.n1365 15.9333
R14990 gnd.n3605 gnd.n1420 15.9333
R14991 gnd.n3604 gnd.n3603 15.9333
R14992 gnd.n3603 gnd.n3602 15.9333
R14993 gnd.n3602 gnd.n3601 15.9333
R14994 gnd.n3601 gnd.n1423 15.9333
R14995 gnd.n1435 gnd.n1423 15.9333
R14996 gnd.n1437 gnd.n1435 15.9333
R14997 gnd.n3595 gnd.n1437 15.9333
R14998 gnd.n3595 gnd.n3594 15.9333
R14999 gnd.n3593 gnd.n3592 15.9333
R15000 gnd.n3592 gnd.n1192 15.9333
R15001 gnd.n4146 gnd.n1192 15.9333
R15002 gnd.n4146 gnd.n4145 15.9333
R15003 gnd.n1203 gnd.n1194 15.9333
R15004 gnd.n4139 gnd.n1203 15.9333
R15005 gnd.n5702 gnd.n5700 15.6674
R15006 gnd.n5670 gnd.n5668 15.6674
R15007 gnd.n5638 gnd.n5636 15.6674
R15008 gnd.n5607 gnd.n5605 15.6674
R15009 gnd.n5575 gnd.n5573 15.6674
R15010 gnd.n5543 gnd.n5541 15.6674
R15011 gnd.n5511 gnd.n5509 15.6674
R15012 gnd.n5480 gnd.n5478 15.6674
R15013 gnd.n4999 gnd.t213 15.6146
R15014 gnd.t148 gnd.n5881 15.6146
R15015 gnd.n5785 gnd.t141 15.6146
R15016 gnd.t177 gnd.n2068 15.6146
R15017 gnd.n3594 gnd.t158 15.6146
R15018 gnd.n2926 gnd.n1713 15.296
R15019 gnd.n2945 gnd.n1704 15.296
R15020 gnd.n2905 gnd.t32 15.296
R15021 gnd.n3075 gnd.n3073 15.296
R15022 gnd.n3119 gnd.n1609 15.296
R15023 gnd.n3247 gnd.t239 15.296
R15024 gnd.n3186 gnd.n1533 15.296
R15025 gnd.n3285 gnd.n1520 15.296
R15026 gnd.n1462 gnd.t127 15.296
R15027 gnd.n3622 gnd.n3621 15.0827
R15028 gnd.n1801 gnd.n1796 15.0481
R15029 gnd.n3632 gnd.n3631 15.0481
R15030 gnd.n5430 gnd.t101 14.9773
R15031 gnd.t191 gnd.n884 14.9773
R15032 gnd.n2771 gnd.n1816 14.9773
R15033 gnd.t201 gnd.n2616 14.6587
R15034 gnd.n2852 gnd.n1736 14.6587
R15035 gnd.n2986 gnd.n2985 14.6587
R15036 gnd.n1561 gnd.n1550 14.6587
R15037 gnd.n3327 gnd.n3326 14.6587
R15038 gnd.t131 gnd.n1458 14.6587
R15039 gnd.n3373 gnd.n3372 14.6587
R15040 gnd.t75 gnd.n4583 14.34
R15041 gnd.t98 gnd.n767 14.34
R15042 gnd.n2810 gnd.t171 14.0214
R15043 gnd.n2860 gnd.n1720 14.0214
R15044 gnd.n2903 gnd.n1689 14.0214
R15045 gnd.n3065 gnd.n3064 14.0214
R15046 gnd.n1599 gnd.n1592 14.0214
R15047 gnd.n3248 gnd.n1537 14.0214
R15048 gnd.n1510 gnd.n1509 14.0214
R15049 gnd.n3614 gnd.n1407 14.0214
R15050 gnd.n5112 gnd.t250 13.7027
R15051 gnd.n1662 gnd.t260 13.7027
R15052 gnd.n3154 gnd.t44 13.7027
R15053 gnd.n4865 gnd.n4864 13.5763
R15054 gnd.n5841 gnd.n4515 13.5763
R15055 gnd.n1340 gnd.n1339 13.5763
R15056 gnd.n6810 gnd.n6809 13.5763
R15057 gnd.n4409 gnd.n876 13.5763
R15058 gnd.n2673 gnd.n2026 13.5763
R15059 gnd.n5147 gnd.n4811 13.384
R15060 gnd.n2790 gnd.n1774 13.384
R15061 gnd.n2884 gnd.n1731 13.384
R15062 gnd.n1690 gnd.n1684 13.384
R15063 gnd.t51 gnd.n2973 13.384
R15064 gnd.n3225 gnd.t14 13.384
R15065 gnd.n3234 gnd.n1546 13.384
R15066 gnd.n3263 gnd.n1498 13.384
R15067 gnd.n3390 gnd.n1449 13.384
R15068 gnd.n1812 gnd.n1793 13.1884
R15069 gnd.n1807 gnd.n1806 13.1884
R15070 gnd.n1806 gnd.n1805 13.1884
R15071 gnd.n3625 gnd.n3620 13.1884
R15072 gnd.n3626 gnd.n3625 13.1884
R15073 gnd.n1808 gnd.n1795 13.146
R15074 gnd.n1804 gnd.n1795 13.146
R15075 gnd.n3624 gnd.n3623 13.146
R15076 gnd.n3624 gnd.n3619 13.146
R15077 gnd.n2826 gnd.t290 13.0654
R15078 gnd.n3348 gnd.t229 13.0654
R15079 gnd.n5703 gnd.n5699 12.8005
R15080 gnd.n5671 gnd.n5667 12.8005
R15081 gnd.n5639 gnd.n5635 12.8005
R15082 gnd.n5608 gnd.n5604 12.8005
R15083 gnd.n5576 gnd.n5572 12.8005
R15084 gnd.n5544 gnd.n5540 12.8005
R15085 gnd.n5512 gnd.n5508 12.8005
R15086 gnd.n5481 gnd.n5477 12.8005
R15087 gnd.n2798 gnd.n1776 12.7467
R15088 gnd.n2843 gnd.t188 12.7467
R15089 gnd.n2868 gnd.n2867 12.7467
R15090 gnd.n3035 gnd.n3033 12.7467
R15091 gnd.n3144 gnd.n1579 12.7467
R15092 gnd.n3312 gnd.n3311 12.7467
R15093 gnd.n4864 gnd.n4859 12.4126
R15094 gnd.n5846 gnd.n4515 12.4126
R15095 gnd.n3884 gnd.n1339 12.4126
R15096 gnd.n6809 gnd.n155 12.4126
R15097 gnd.n4405 gnd.n876 12.4126
R15098 gnd.n2668 gnd.n2026 12.4126
R15099 gnd.n2775 gnd.n2774 12.1761
R15100 gnd.n3701 gnd.n3700 12.1761
R15101 gnd.n2780 gnd.n2779 12.1094
R15102 gnd.t145 gnd.n1781 12.1094
R15103 gnd.n2875 gnd.n1721 12.1094
R15104 gnd.n2956 gnd.n1695 12.1094
R15105 gnd.n3255 gnd.n1531 12.1094
R15106 gnd.n3297 gnd.n1507 12.1094
R15107 gnd.n3397 gnd.n1410 12.1094
R15108 gnd.n5707 gnd.n5706 12.0247
R15109 gnd.n5675 gnd.n5674 12.0247
R15110 gnd.n5643 gnd.n5642 12.0247
R15111 gnd.n5612 gnd.n5611 12.0247
R15112 gnd.n5580 gnd.n5579 12.0247
R15113 gnd.n5548 gnd.n5547 12.0247
R15114 gnd.n5516 gnd.n5515 12.0247
R15115 gnd.n5485 gnd.n5484 12.0247
R15116 gnd.t28 gnd.n898 11.7908
R15117 gnd.n4295 gnd.t60 11.7908
R15118 gnd.n4020 gnd.t79 11.7908
R15119 gnd.n6711 gnd.t66 11.7908
R15120 gnd.n2575 gnd.n1996 11.4721
R15121 gnd.n2836 gnd.n1752 11.4721
R15122 gnd.n2828 gnd.n2827 11.4721
R15123 gnd.n2995 gnd.t235 11.4721
R15124 gnd.n2993 gnd.n1671 11.4721
R15125 gnd.n3025 gnd.n3024 11.4721
R15126 gnd.n3172 gnd.n1574 11.4721
R15127 gnd.n3164 gnd.n1560 11.4721
R15128 gnd.n3216 gnd.t17 11.4721
R15129 gnd.n3338 gnd.n1485 11.4721
R15130 gnd.n3359 gnd.n3358 11.4721
R15131 gnd.n4137 gnd.n1204 11.4721
R15132 gnd.n5710 gnd.n5697 11.249
R15133 gnd.n5678 gnd.n5665 11.249
R15134 gnd.n5646 gnd.n5633 11.249
R15135 gnd.n5615 gnd.n5602 11.249
R15136 gnd.n5583 gnd.n5570 11.249
R15137 gnd.n5551 gnd.n5538 11.249
R15138 gnd.n5519 gnd.n5506 11.249
R15139 gnd.n5488 gnd.n5475 11.249
R15140 gnd.n5220 gnd.t250 11.1535
R15141 gnd.t0 gnd.n939 11.1535
R15142 gnd.n4319 gnd.t20 11.1535
R15143 gnd.n2624 gnd.t232 11.1535
R15144 gnd.n2972 gnd.t109 11.1535
R15145 gnd.t254 gnd.n3226 11.1535
R15146 gnd.t52 gnd.n3604 11.1535
R15147 gnd.n4080 gnd.t104 11.1535
R15148 gnd.n6679 gnd.t18 11.1535
R15149 gnd.n2462 gnd.n960 10.8348
R15150 gnd.n4345 gnd.n973 10.8348
R15151 gnd.n2431 gnd.n978 10.8348
R15152 gnd.n2453 gnd.n987 10.8348
R15153 gnd.n4332 gnd.n990 10.8348
R15154 gnd.n2445 gnd.n995 10.8348
R15155 gnd.n4325 gnd.n998 10.8348
R15156 gnd.n2502 gnd.n2501 10.8348
R15157 gnd.n4319 gnd.n1008 10.8348
R15158 gnd.n2510 gnd.n1016 10.8348
R15159 gnd.n2518 gnd.n1026 10.8348
R15160 gnd.n4307 gnd.n1029 10.8348
R15161 gnd.n2526 gnd.n1037 10.8348
R15162 gnd.n4301 gnd.n1040 10.8348
R15163 gnd.n2555 gnd.n2554 10.8348
R15164 gnd.n4295 gnd.n1050 10.8348
R15165 gnd.n2534 gnd.n1058 10.8348
R15166 gnd.n4289 gnd.n1061 10.8348
R15167 gnd.n2543 gnd.n1069 10.8348
R15168 gnd.n4283 gnd.n1072 10.8348
R15169 gnd.n2662 gnd.n1079 10.8348
R15170 gnd.n4277 gnd.n1082 10.8348
R15171 gnd.n2939 gnd.n2938 10.8348
R15172 gnd.n2938 gnd.n2937 10.8348
R15173 gnd.n3113 gnd.n3112 10.8348
R15174 gnd.n3112 gnd.n1606 10.8348
R15175 gnd.n3279 gnd.n3278 10.8348
R15176 gnd.n3278 gnd.n1517 10.8348
R15177 gnd.n4131 gnd.n4130 10.8348
R15178 gnd.n3890 gnd.n1215 10.8348
R15179 gnd.n4124 gnd.n1224 10.8348
R15180 gnd.n3899 gnd.n1227 10.8348
R15181 gnd.n4010 gnd.n1325 10.8348
R15182 gnd.n4009 gnd.n3992 10.8348
R15183 gnd.n4020 gnd.n1318 10.8348
R15184 gnd.n1320 gnd.n1310 10.8348
R15185 gnd.n4030 gnd.n4029 10.8348
R15186 gnd.n4041 gnd.n1299 10.8348
R15187 gnd.n4040 gnd.n1302 10.8348
R15188 gnd.n4052 gnd.n1289 10.8348
R15189 gnd.n4062 gnd.n4061 10.8348
R15190 gnd.n4080 gnd.n1270 10.8348
R15191 gnd.n4079 gnd.n1274 10.8348
R15192 gnd.n4086 gnd.n1260 10.8348
R15193 gnd.n3972 gnd.n1262 10.8348
R15194 gnd.n4095 gnd.n1251 10.8348
R15195 gnd.n6644 gnd.n248 10.8348
R15196 gnd.n3966 gnd.n246 10.8348
R15197 gnd.n6657 gnd.n236 10.8348
R15198 gnd.n6636 gnd.n230 10.8348
R15199 gnd.n3766 gnd.n1361 10.6151
R15200 gnd.n3766 gnd.n3765 10.6151
R15201 gnd.n3763 gnd.n3760 10.6151
R15202 gnd.n3760 gnd.n3759 10.6151
R15203 gnd.n3759 gnd.n3756 10.6151
R15204 gnd.n3756 gnd.n3755 10.6151
R15205 gnd.n3755 gnd.n3752 10.6151
R15206 gnd.n3752 gnd.n3751 10.6151
R15207 gnd.n3751 gnd.n3748 10.6151
R15208 gnd.n3748 gnd.n3747 10.6151
R15209 gnd.n3747 gnd.n3744 10.6151
R15210 gnd.n3744 gnd.n3743 10.6151
R15211 gnd.n3743 gnd.n3740 10.6151
R15212 gnd.n3740 gnd.n3739 10.6151
R15213 gnd.n3739 gnd.n3736 10.6151
R15214 gnd.n3736 gnd.n3735 10.6151
R15215 gnd.n3735 gnd.n3732 10.6151
R15216 gnd.n3732 gnd.n3731 10.6151
R15217 gnd.n3731 gnd.n3728 10.6151
R15218 gnd.n3728 gnd.n3727 10.6151
R15219 gnd.n3727 gnd.n3724 10.6151
R15220 gnd.n3724 gnd.n3723 10.6151
R15221 gnd.n3723 gnd.n3720 10.6151
R15222 gnd.n3720 gnd.n3719 10.6151
R15223 gnd.n3719 gnd.n3716 10.6151
R15224 gnd.n3716 gnd.n3715 10.6151
R15225 gnd.n3715 gnd.n3712 10.6151
R15226 gnd.n3712 gnd.n3711 10.6151
R15227 gnd.n3711 gnd.n3708 10.6151
R15228 gnd.n3708 gnd.n3707 10.6151
R15229 gnd.n1867 gnd.n1866 10.6151
R15230 gnd.n1866 gnd.n1865 10.6151
R15231 gnd.n1865 gnd.n1861 10.6151
R15232 gnd.n1861 gnd.n1860 10.6151
R15233 gnd.n1860 gnd.n1858 10.6151
R15234 gnd.n1858 gnd.n1857 10.6151
R15235 gnd.n1857 gnd.n1749 10.6151
R15236 gnd.n2838 gnd.n1749 10.6151
R15237 gnd.n2839 gnd.n2838 10.6151
R15238 gnd.n2841 gnd.n2839 10.6151
R15239 gnd.n2841 gnd.n2840 10.6151
R15240 gnd.n2840 gnd.n1738 10.6151
R15241 gnd.n2854 gnd.n1738 10.6151
R15242 gnd.n2855 gnd.n2854 10.6151
R15243 gnd.n2865 gnd.n2855 10.6151
R15244 gnd.n2865 gnd.n2864 10.6151
R15245 gnd.n2864 gnd.n2863 10.6151
R15246 gnd.n2863 gnd.n2856 10.6151
R15247 gnd.n2857 gnd.n2856 10.6151
R15248 gnd.n2857 gnd.n1711 10.6151
R15249 gnd.n2928 gnd.n1711 10.6151
R15250 gnd.n2929 gnd.n2928 10.6151
R15251 gnd.n2935 gnd.n2929 10.6151
R15252 gnd.n2935 gnd.n2934 10.6151
R15253 gnd.n2934 gnd.n2933 10.6151
R15254 gnd.n2933 gnd.n2930 10.6151
R15255 gnd.n2930 gnd.n1687 10.6151
R15256 gnd.n2965 gnd.n1687 10.6151
R15257 gnd.n2966 gnd.n2965 10.6151
R15258 gnd.n2970 gnd.n2966 10.6151
R15259 gnd.n2970 gnd.n2969 10.6151
R15260 gnd.n2969 gnd.n2968 10.6151
R15261 gnd.n2968 gnd.n2967 10.6151
R15262 gnd.n2967 gnd.n1661 10.6151
R15263 gnd.n3013 gnd.n1661 10.6151
R15264 gnd.n3013 gnd.n3012 10.6151
R15265 gnd.n3012 gnd.n3011 10.6151
R15266 gnd.n3011 gnd.n3010 10.6151
R15267 gnd.n3010 gnd.n1643 10.6151
R15268 gnd.n3037 gnd.n1643 10.6151
R15269 gnd.n3038 gnd.n3037 10.6151
R15270 gnd.n3040 gnd.n3038 10.6151
R15271 gnd.n3041 gnd.n3040 10.6151
R15272 gnd.n3042 gnd.n3041 10.6151
R15273 gnd.n3042 gnd.n1620 10.6151
R15274 gnd.n3077 gnd.n1620 10.6151
R15275 gnd.n3078 gnd.n3077 10.6151
R15276 gnd.n3080 gnd.n3078 10.6151
R15277 gnd.n3081 gnd.n3080 10.6151
R15278 gnd.n3083 gnd.n3081 10.6151
R15279 gnd.n3083 gnd.n3082 10.6151
R15280 gnd.n3082 gnd.n1590 10.6151
R15281 gnd.n3139 gnd.n1590 10.6151
R15282 gnd.n3140 gnd.n3139 10.6151
R15283 gnd.n3142 gnd.n3140 10.6151
R15284 gnd.n3142 gnd.n3141 10.6151
R15285 gnd.n3141 gnd.n1571 10.6151
R15286 gnd.n3174 gnd.n1571 10.6151
R15287 gnd.n3175 gnd.n3174 10.6151
R15288 gnd.n3204 gnd.n3175 10.6151
R15289 gnd.n3204 gnd.n3203 10.6151
R15290 gnd.n3203 gnd.n3202 10.6151
R15291 gnd.n3202 gnd.n3199 10.6151
R15292 gnd.n3199 gnd.n3198 10.6151
R15293 gnd.n3198 gnd.n3197 10.6151
R15294 gnd.n3197 gnd.n3196 10.6151
R15295 gnd.n3196 gnd.n3195 10.6151
R15296 gnd.n3195 gnd.n3192 10.6151
R15297 gnd.n3192 gnd.n3191 10.6151
R15298 gnd.n3191 gnd.n3189 10.6151
R15299 gnd.n3189 gnd.n3188 10.6151
R15300 gnd.n3188 gnd.n3183 10.6151
R15301 gnd.n3183 gnd.n3182 10.6151
R15302 gnd.n3182 gnd.n3180 10.6151
R15303 gnd.n3180 gnd.n3179 10.6151
R15304 gnd.n3179 gnd.n3176 10.6151
R15305 gnd.n3176 gnd.n1501 10.6151
R15306 gnd.n3306 gnd.n1501 10.6151
R15307 gnd.n3307 gnd.n3306 10.6151
R15308 gnd.n3309 gnd.n3307 10.6151
R15309 gnd.n3309 gnd.n3308 10.6151
R15310 gnd.n3308 gnd.n1482 10.6151
R15311 gnd.n3340 gnd.n1482 10.6151
R15312 gnd.n3341 gnd.n3340 10.6151
R15313 gnd.n3345 gnd.n3341 10.6151
R15314 gnd.n3345 gnd.n3344 10.6151
R15315 gnd.n3344 gnd.n3343 10.6151
R15316 gnd.n3343 gnd.n3342 10.6151
R15317 gnd.n3342 gnd.n1451 10.6151
R15318 gnd.n3382 gnd.n1451 10.6151
R15319 gnd.n3383 gnd.n3382 10.6151
R15320 gnd.n3386 gnd.n3383 10.6151
R15321 gnd.n3386 gnd.n3385 10.6151
R15322 gnd.n3385 gnd.n3384 10.6151
R15323 gnd.n3384 gnd.n1400 10.6151
R15324 gnd.n1932 gnd.n1931 10.6151
R15325 gnd.n1931 gnd.n1928 10.6151
R15326 gnd.n1926 gnd.n1923 10.6151
R15327 gnd.n1923 gnd.n1922 10.6151
R15328 gnd.n1922 gnd.n1919 10.6151
R15329 gnd.n1919 gnd.n1918 10.6151
R15330 gnd.n1918 gnd.n1915 10.6151
R15331 gnd.n1915 gnd.n1914 10.6151
R15332 gnd.n1914 gnd.n1911 10.6151
R15333 gnd.n1911 gnd.n1910 10.6151
R15334 gnd.n1910 gnd.n1907 10.6151
R15335 gnd.n1907 gnd.n1906 10.6151
R15336 gnd.n1906 gnd.n1903 10.6151
R15337 gnd.n1903 gnd.n1902 10.6151
R15338 gnd.n1902 gnd.n1899 10.6151
R15339 gnd.n1899 gnd.n1898 10.6151
R15340 gnd.n1898 gnd.n1895 10.6151
R15341 gnd.n1895 gnd.n1894 10.6151
R15342 gnd.n1894 gnd.n1891 10.6151
R15343 gnd.n1891 gnd.n1890 10.6151
R15344 gnd.n1890 gnd.n1887 10.6151
R15345 gnd.n1887 gnd.n1886 10.6151
R15346 gnd.n1886 gnd.n1883 10.6151
R15347 gnd.n1883 gnd.n1882 10.6151
R15348 gnd.n1882 gnd.n1879 10.6151
R15349 gnd.n1879 gnd.n1878 10.6151
R15350 gnd.n1878 gnd.n1875 10.6151
R15351 gnd.n1875 gnd.n1874 10.6151
R15352 gnd.n1874 gnd.n1871 10.6151
R15353 gnd.n1871 gnd.n1870 10.6151
R15354 gnd.n2774 gnd.n1813 10.6151
R15355 gnd.n2769 gnd.n1813 10.6151
R15356 gnd.n2769 gnd.n2768 10.6151
R15357 gnd.n2768 gnd.n2767 10.6151
R15358 gnd.n2767 gnd.n2764 10.6151
R15359 gnd.n2764 gnd.n2763 10.6151
R15360 gnd.n2763 gnd.n2760 10.6151
R15361 gnd.n2760 gnd.n2759 10.6151
R15362 gnd.n2759 gnd.n2756 10.6151
R15363 gnd.n2756 gnd.n2755 10.6151
R15364 gnd.n2755 gnd.n2752 10.6151
R15365 gnd.n2752 gnd.n2751 10.6151
R15366 gnd.n2751 gnd.n2748 10.6151
R15367 gnd.n2748 gnd.n2747 10.6151
R15368 gnd.n2747 gnd.n2744 10.6151
R15369 gnd.n2744 gnd.n2743 10.6151
R15370 gnd.n2743 gnd.n2740 10.6151
R15371 gnd.n2740 gnd.n2739 10.6151
R15372 gnd.n2739 gnd.n2736 10.6151
R15373 gnd.n2736 gnd.n2735 10.6151
R15374 gnd.n2735 gnd.n2732 10.6151
R15375 gnd.n2732 gnd.n2731 10.6151
R15376 gnd.n2731 gnd.n2728 10.6151
R15377 gnd.n2728 gnd.n2727 10.6151
R15378 gnd.n2727 gnd.n2724 10.6151
R15379 gnd.n2724 gnd.n2723 10.6151
R15380 gnd.n2723 gnd.n2720 10.6151
R15381 gnd.n2720 gnd.n2719 10.6151
R15382 gnd.n2716 gnd.n2715 10.6151
R15383 gnd.n2715 gnd.n2712 10.6151
R15384 gnd.n3700 gnd.n3699 10.6151
R15385 gnd.n3699 gnd.n3696 10.6151
R15386 gnd.n3696 gnd.n3695 10.6151
R15387 gnd.n3695 gnd.n3692 10.6151
R15388 gnd.n3692 gnd.n3691 10.6151
R15389 gnd.n3691 gnd.n3688 10.6151
R15390 gnd.n3688 gnd.n3687 10.6151
R15391 gnd.n3687 gnd.n3684 10.6151
R15392 gnd.n3684 gnd.n3683 10.6151
R15393 gnd.n3683 gnd.n3680 10.6151
R15394 gnd.n3680 gnd.n3679 10.6151
R15395 gnd.n3679 gnd.n3676 10.6151
R15396 gnd.n3676 gnd.n3675 10.6151
R15397 gnd.n3675 gnd.n3672 10.6151
R15398 gnd.n3672 gnd.n3671 10.6151
R15399 gnd.n3671 gnd.n3668 10.6151
R15400 gnd.n3668 gnd.n3667 10.6151
R15401 gnd.n3667 gnd.n3664 10.6151
R15402 gnd.n3664 gnd.n3663 10.6151
R15403 gnd.n3663 gnd.n3660 10.6151
R15404 gnd.n3660 gnd.n3659 10.6151
R15405 gnd.n3659 gnd.n3656 10.6151
R15406 gnd.n3656 gnd.n3655 10.6151
R15407 gnd.n3655 gnd.n3652 10.6151
R15408 gnd.n3652 gnd.n3651 10.6151
R15409 gnd.n3651 gnd.n3648 10.6151
R15410 gnd.n3648 gnd.n3647 10.6151
R15411 gnd.n3647 gnd.n3644 10.6151
R15412 gnd.n3642 gnd.n3639 10.6151
R15413 gnd.n3639 gnd.n1362 10.6151
R15414 gnd.n2777 gnd.n2776 10.6151
R15415 gnd.n2777 gnd.n1779 10.6151
R15416 gnd.n2793 gnd.n1779 10.6151
R15417 gnd.n2794 gnd.n2793 10.6151
R15418 gnd.n2796 gnd.n2794 10.6151
R15419 gnd.n2796 gnd.n2795 10.6151
R15420 gnd.n2795 gnd.n1755 10.6151
R15421 gnd.n2834 gnd.n1755 10.6151
R15422 gnd.n2834 gnd.n2833 10.6151
R15423 gnd.n2833 gnd.n2832 10.6151
R15424 gnd.n2832 gnd.n2831 10.6151
R15425 gnd.n2831 gnd.n1756 10.6151
R15426 gnd.n1756 gnd.n1734 10.6151
R15427 gnd.n2871 gnd.n1734 10.6151
R15428 gnd.n2872 gnd.n2871 10.6151
R15429 gnd.n2882 gnd.n2872 10.6151
R15430 gnd.n2882 gnd.n2881 10.6151
R15431 gnd.n2881 gnd.n2880 10.6151
R15432 gnd.n2880 gnd.n2873 10.6151
R15433 gnd.n2874 gnd.n2873 10.6151
R15434 gnd.n2874 gnd.n1706 10.6151
R15435 gnd.n2941 gnd.n1706 10.6151
R15436 gnd.n2942 gnd.n2941 10.6151
R15437 gnd.n2943 gnd.n2942 10.6151
R15438 gnd.n2943 gnd.n1693 10.6151
R15439 gnd.n2958 gnd.n1693 10.6151
R15440 gnd.n2959 gnd.n2958 10.6151
R15441 gnd.n2961 gnd.n2959 10.6151
R15442 gnd.n2961 gnd.n2960 10.6151
R15443 gnd.n2960 gnd.n1673 10.6151
R15444 gnd.n2989 gnd.n1673 10.6151
R15445 gnd.n2990 gnd.n2989 10.6151
R15446 gnd.n2991 gnd.n2990 10.6151
R15447 gnd.n2991 gnd.n1656 10.6151
R15448 gnd.n3017 gnd.n1656 10.6151
R15449 gnd.n3018 gnd.n3017 10.6151
R15450 gnd.n3022 gnd.n3018 10.6151
R15451 gnd.n3022 gnd.n3021 10.6151
R15452 gnd.n3021 gnd.n3020 10.6151
R15453 gnd.n3020 gnd.n1633 10.6151
R15454 gnd.n3057 gnd.n1633 10.6151
R15455 gnd.n3058 gnd.n3057 10.6151
R15456 gnd.n3062 gnd.n3058 10.6151
R15457 gnd.n3062 gnd.n3061 10.6151
R15458 gnd.n3061 gnd.n3060 10.6151
R15459 gnd.n3060 gnd.n1611 10.6151
R15460 gnd.n3115 gnd.n1611 10.6151
R15461 gnd.n3116 gnd.n3115 10.6151
R15462 gnd.n3117 gnd.n3116 10.6151
R15463 gnd.n3117 gnd.n1596 10.6151
R15464 gnd.n3132 gnd.n1596 10.6151
R15465 gnd.n3133 gnd.n3132 10.6151
R15466 gnd.n3135 gnd.n3133 10.6151
R15467 gnd.n3135 gnd.n3134 10.6151
R15468 gnd.n3134 gnd.n1577 10.6151
R15469 gnd.n3160 gnd.n1577 10.6151
R15470 gnd.n3161 gnd.n3160 10.6151
R15471 gnd.n3170 gnd.n3161 10.6151
R15472 gnd.n3170 gnd.n3169 10.6151
R15473 gnd.n3169 gnd.n3168 10.6151
R15474 gnd.n3168 gnd.n3167 10.6151
R15475 gnd.n3167 gnd.n3162 10.6151
R15476 gnd.n3162 gnd.n1548 10.6151
R15477 gnd.n3230 gnd.n1548 10.6151
R15478 gnd.n3231 gnd.n3230 10.6151
R15479 gnd.n3232 gnd.n3231 10.6151
R15480 gnd.n3232 gnd.n1535 10.6151
R15481 gnd.n3250 gnd.n1535 10.6151
R15482 gnd.n3251 gnd.n3250 10.6151
R15483 gnd.n3252 gnd.n3251 10.6151
R15484 gnd.n3252 gnd.n1522 10.6151
R15485 gnd.n3281 gnd.n1522 10.6151
R15486 gnd.n3282 gnd.n3281 10.6151
R15487 gnd.n3283 gnd.n3282 10.6151
R15488 gnd.n3283 gnd.n1505 10.6151
R15489 gnd.n3299 gnd.n1505 10.6151
R15490 gnd.n3300 gnd.n3299 10.6151
R15491 gnd.n3302 gnd.n3300 10.6151
R15492 gnd.n3302 gnd.n3301 10.6151
R15493 gnd.n3301 gnd.n1488 10.6151
R15494 gnd.n3330 gnd.n1488 10.6151
R15495 gnd.n3331 gnd.n3330 10.6151
R15496 gnd.n3336 gnd.n3331 10.6151
R15497 gnd.n3336 gnd.n3335 10.6151
R15498 gnd.n3335 gnd.n3334 10.6151
R15499 gnd.n3334 gnd.n3333 10.6151
R15500 gnd.n3333 gnd.n1456 10.6151
R15501 gnd.n3375 gnd.n1456 10.6151
R15502 gnd.n3376 gnd.n3375 10.6151
R15503 gnd.n3378 gnd.n3376 10.6151
R15504 gnd.n3378 gnd.n3377 10.6151
R15505 gnd.n3377 gnd.n1405 10.6151
R15506 gnd.n3616 gnd.n1405 10.6151
R15507 gnd.n3617 gnd.n3616 10.6151
R15508 gnd.n3702 gnd.n3617 10.6151
R15509 gnd.n5136 gnd.t107 10.5161
R15510 gnd.n4585 gnd.t75 10.5161
R15511 gnd.n5774 gnd.t98 10.5161
R15512 gnd.n4351 gnd.n957 10.5161
R15513 gnd.n2462 gnd.t25 10.5161
R15514 gnd.n4345 gnd.t25 10.5161
R15515 gnd.n4338 gnd.t2 10.5161
R15516 gnd.n2947 gnd.t71 10.5161
R15517 gnd.t82 gnd.n3184 10.5161
R15518 gnd.n6649 gnd.t102 10.5161
R15519 gnd.n6657 gnd.t64 10.5161
R15520 gnd.n6636 gnd.t64 10.5161
R15521 gnd.n6663 gnd.n232 10.5161
R15522 gnd.n5711 gnd.n5695 10.4732
R15523 gnd.n5679 gnd.n5663 10.4732
R15524 gnd.n5647 gnd.n5631 10.4732
R15525 gnd.n5616 gnd.n5600 10.4732
R15526 gnd.n5584 gnd.n5568 10.4732
R15527 gnd.n5552 gnd.n5536 10.4732
R15528 gnd.n5520 gnd.n5504 10.4732
R15529 gnd.n5489 gnd.n5473 10.4732
R15530 gnd.n1758 gnd.n1752 10.1975
R15531 gnd.n1671 gnd.n1670 10.1975
R15532 gnd.n3025 gnd.n1651 10.1975
R15533 gnd.n3094 gnd.n1574 10.1975
R15534 gnd.n3165 gnd.n3164 10.1975
R15535 gnd.n3359 gnd.n1468 10.1975
R15536 gnd.n1420 gnd.t162 10.1975
R15537 gnd.n5443 gnd.t101 9.87883
R15538 gnd.n936 gnd.t35 9.87883
R15539 gnd.n2501 gnd.t20 9.87883
R15540 gnd.n4313 gnd.t42 9.87883
R15541 gnd.t38 gnd.n1281 9.87883
R15542 gnd.t104 gnd.n4079 9.87883
R15543 gnd.n6687 gnd.t23 9.87883
R15544 gnd.n5715 gnd.n5714 9.69747
R15545 gnd.n5683 gnd.n5682 9.69747
R15546 gnd.n5651 gnd.n5650 9.69747
R15547 gnd.n5620 gnd.n5619 9.69747
R15548 gnd.n5588 gnd.n5587 9.69747
R15549 gnd.n5556 gnd.n5555 9.69747
R15550 gnd.n5524 gnd.n5523 9.69747
R15551 gnd.n5493 gnd.n5492 9.69747
R15552 gnd.n6916 gnd.n50 9.6512
R15553 gnd.n2780 gnd.n1789 9.56018
R15554 gnd.n2876 gnd.n2875 9.56018
R15555 gnd.n2931 gnd.n1695 9.56018
R15556 gnd.n2998 gnd.t16 9.56018
R15557 gnd.n3046 gnd.n1622 9.56018
R15558 gnd.n3087 gnd.n3085 9.56018
R15559 gnd.n3095 gnd.t27 9.56018
R15560 gnd.n3255 gnd.n3254 9.56018
R15561 gnd.n3177 gnd.n1507 9.56018
R15562 gnd.n4273 gnd.n1085 9.45599
R15563 gnd.n3470 gnd.n3469 9.45599
R15564 gnd.n5721 gnd.n5720 9.45567
R15565 gnd.n5689 gnd.n5688 9.45567
R15566 gnd.n5657 gnd.n5656 9.45567
R15567 gnd.n5626 gnd.n5625 9.45567
R15568 gnd.n5594 gnd.n5593 9.45567
R15569 gnd.n5562 gnd.n5561 9.45567
R15570 gnd.n5530 gnd.n5529 9.45567
R15571 gnd.n5499 gnd.n5498 9.45567
R15572 gnd.n5099 gnd.n5098 9.39724
R15573 gnd.n5720 gnd.n5719 9.3005
R15574 gnd.n5693 gnd.n5692 9.3005
R15575 gnd.n5714 gnd.n5713 9.3005
R15576 gnd.n5712 gnd.n5711 9.3005
R15577 gnd.n5697 gnd.n5696 9.3005
R15578 gnd.n5706 gnd.n5705 9.3005
R15579 gnd.n5704 gnd.n5703 9.3005
R15580 gnd.n5688 gnd.n5687 9.3005
R15581 gnd.n5661 gnd.n5660 9.3005
R15582 gnd.n5682 gnd.n5681 9.3005
R15583 gnd.n5680 gnd.n5679 9.3005
R15584 gnd.n5665 gnd.n5664 9.3005
R15585 gnd.n5674 gnd.n5673 9.3005
R15586 gnd.n5672 gnd.n5671 9.3005
R15587 gnd.n5656 gnd.n5655 9.3005
R15588 gnd.n5629 gnd.n5628 9.3005
R15589 gnd.n5650 gnd.n5649 9.3005
R15590 gnd.n5648 gnd.n5647 9.3005
R15591 gnd.n5633 gnd.n5632 9.3005
R15592 gnd.n5642 gnd.n5641 9.3005
R15593 gnd.n5640 gnd.n5639 9.3005
R15594 gnd.n5625 gnd.n5624 9.3005
R15595 gnd.n5598 gnd.n5597 9.3005
R15596 gnd.n5619 gnd.n5618 9.3005
R15597 gnd.n5617 gnd.n5616 9.3005
R15598 gnd.n5602 gnd.n5601 9.3005
R15599 gnd.n5611 gnd.n5610 9.3005
R15600 gnd.n5609 gnd.n5608 9.3005
R15601 gnd.n5593 gnd.n5592 9.3005
R15602 gnd.n5566 gnd.n5565 9.3005
R15603 gnd.n5587 gnd.n5586 9.3005
R15604 gnd.n5585 gnd.n5584 9.3005
R15605 gnd.n5570 gnd.n5569 9.3005
R15606 gnd.n5579 gnd.n5578 9.3005
R15607 gnd.n5577 gnd.n5576 9.3005
R15608 gnd.n5561 gnd.n5560 9.3005
R15609 gnd.n5534 gnd.n5533 9.3005
R15610 gnd.n5555 gnd.n5554 9.3005
R15611 gnd.n5553 gnd.n5552 9.3005
R15612 gnd.n5538 gnd.n5537 9.3005
R15613 gnd.n5547 gnd.n5546 9.3005
R15614 gnd.n5545 gnd.n5544 9.3005
R15615 gnd.n5529 gnd.n5528 9.3005
R15616 gnd.n5502 gnd.n5501 9.3005
R15617 gnd.n5523 gnd.n5522 9.3005
R15618 gnd.n5521 gnd.n5520 9.3005
R15619 gnd.n5506 gnd.n5505 9.3005
R15620 gnd.n5515 gnd.n5514 9.3005
R15621 gnd.n5513 gnd.n5512 9.3005
R15622 gnd.n5498 gnd.n5497 9.3005
R15623 gnd.n5471 gnd.n5470 9.3005
R15624 gnd.n5492 gnd.n5491 9.3005
R15625 gnd.n5490 gnd.n5489 9.3005
R15626 gnd.n5475 gnd.n5474 9.3005
R15627 gnd.n5484 gnd.n5483 9.3005
R15628 gnd.n5482 gnd.n5481 9.3005
R15629 gnd.n5868 gnd.n4489 9.3005
R15630 gnd.n5867 gnd.n4491 9.3005
R15631 gnd.n4495 gnd.n4492 9.3005
R15632 gnd.n5862 gnd.n4496 9.3005
R15633 gnd.n5861 gnd.n4497 9.3005
R15634 gnd.n5860 gnd.n4498 9.3005
R15635 gnd.n4502 gnd.n4499 9.3005
R15636 gnd.n5855 gnd.n4503 9.3005
R15637 gnd.n5854 gnd.n4504 9.3005
R15638 gnd.n5853 gnd.n4505 9.3005
R15639 gnd.n4509 gnd.n4506 9.3005
R15640 gnd.n5848 gnd.n4510 9.3005
R15641 gnd.n5847 gnd.n4511 9.3005
R15642 gnd.n5846 gnd.n4512 9.3005
R15643 gnd.n4517 gnd.n4515 9.3005
R15644 gnd.n5841 gnd.n5840 9.3005
R15645 gnd.n5870 gnd.n5869 9.3005
R15646 gnd.n5155 gnd.n5154 9.3005
R15647 gnd.n4785 gnd.n4784 9.3005
R15648 gnd.n5182 gnd.n5181 9.3005
R15649 gnd.n5183 gnd.n4783 9.3005
R15650 gnd.n5187 gnd.n5184 9.3005
R15651 gnd.n5186 gnd.n5185 9.3005
R15652 gnd.n4759 gnd.n4758 9.3005
R15653 gnd.n5213 gnd.n5212 9.3005
R15654 gnd.n5214 gnd.n4757 9.3005
R15655 gnd.n5218 gnd.n5215 9.3005
R15656 gnd.n5217 gnd.n5216 9.3005
R15657 gnd.n4734 gnd.n4733 9.3005
R15658 gnd.n5244 gnd.n5243 9.3005
R15659 gnd.n5245 gnd.n4732 9.3005
R15660 gnd.n5249 gnd.n5246 9.3005
R15661 gnd.n5248 gnd.n5247 9.3005
R15662 gnd.n4708 gnd.n4707 9.3005
R15663 gnd.n5275 gnd.n5274 9.3005
R15664 gnd.n5276 gnd.n4706 9.3005
R15665 gnd.n5280 gnd.n5277 9.3005
R15666 gnd.n5279 gnd.n5278 9.3005
R15667 gnd.n4684 gnd.n4683 9.3005
R15668 gnd.n5305 gnd.n5304 9.3005
R15669 gnd.n5306 gnd.n4682 9.3005
R15670 gnd.n5310 gnd.n5307 9.3005
R15671 gnd.n5309 gnd.n5308 9.3005
R15672 gnd.n4653 gnd.n4652 9.3005
R15673 gnd.n5359 gnd.n5358 9.3005
R15674 gnd.n5360 gnd.n4651 9.3005
R15675 gnd.n5362 gnd.n5361 9.3005
R15676 gnd.n4632 gnd.n4631 9.3005
R15677 gnd.n5389 gnd.n5388 9.3005
R15678 gnd.n5390 gnd.n4630 9.3005
R15679 gnd.n5394 gnd.n5391 9.3005
R15680 gnd.n5393 gnd.n5392 9.3005
R15681 gnd.n4608 gnd.n4607 9.3005
R15682 gnd.n5435 gnd.n5434 9.3005
R15683 gnd.n5436 gnd.n4606 9.3005
R15684 gnd.n5440 gnd.n5437 9.3005
R15685 gnd.n5439 gnd.n5438 9.3005
R15686 gnd.n4578 gnd.n4577 9.3005
R15687 gnd.n5756 gnd.n5755 9.3005
R15688 gnd.n5757 gnd.n4576 9.3005
R15689 gnd.n5765 gnd.n5758 9.3005
R15690 gnd.n5764 gnd.n5759 9.3005
R15691 gnd.n5763 gnd.n5761 9.3005
R15692 gnd.n5760 gnd.n782 9.3005
R15693 gnd.n5886 gnd.n783 9.3005
R15694 gnd.n5885 gnd.n784 9.3005
R15695 gnd.n5884 gnd.n785 9.3005
R15696 gnd.n4487 gnd.n786 9.3005
R15697 gnd.n4488 gnd.n4486 9.3005
R15698 gnd.n5872 gnd.n5871 9.3005
R15699 gnd.n5156 gnd.n5153 9.3005
R15700 gnd.n4864 gnd.n4823 9.3005
R15701 gnd.n4859 gnd.n4858 9.3005
R15702 gnd.n4857 gnd.n4824 9.3005
R15703 gnd.n4856 gnd.n4855 9.3005
R15704 gnd.n4852 gnd.n4825 9.3005
R15705 gnd.n4849 gnd.n4848 9.3005
R15706 gnd.n4847 gnd.n4826 9.3005
R15707 gnd.n4846 gnd.n4845 9.3005
R15708 gnd.n4842 gnd.n4827 9.3005
R15709 gnd.n4839 gnd.n4838 9.3005
R15710 gnd.n4837 gnd.n4828 9.3005
R15711 gnd.n4836 gnd.n4835 9.3005
R15712 gnd.n4832 gnd.n4830 9.3005
R15713 gnd.n4829 gnd.n4809 9.3005
R15714 gnd.n5150 gnd.n4808 9.3005
R15715 gnd.n5152 gnd.n5151 9.3005
R15716 gnd.n4866 gnd.n4865 9.3005
R15717 gnd.n5163 gnd.n4795 9.3005
R15718 gnd.n5170 gnd.n4796 9.3005
R15719 gnd.n5172 gnd.n5171 9.3005
R15720 gnd.n5173 gnd.n4776 9.3005
R15721 gnd.n5192 gnd.n5191 9.3005
R15722 gnd.n5194 gnd.n4769 9.3005
R15723 gnd.n5201 gnd.n4770 9.3005
R15724 gnd.n5203 gnd.n5202 9.3005
R15725 gnd.n5204 gnd.n4752 9.3005
R15726 gnd.n5223 gnd.n5222 9.3005
R15727 gnd.n5225 gnd.n4744 9.3005
R15728 gnd.n5232 gnd.n4745 9.3005
R15729 gnd.n5234 gnd.n5233 9.3005
R15730 gnd.n5235 gnd.n4726 9.3005
R15731 gnd.n5254 gnd.n5253 9.3005
R15732 gnd.n5256 gnd.n4718 9.3005
R15733 gnd.n5263 gnd.n4719 9.3005
R15734 gnd.n5265 gnd.n5264 9.3005
R15735 gnd.n5266 gnd.n4701 9.3005
R15736 gnd.n5285 gnd.n5284 9.3005
R15737 gnd.n5287 gnd.n4693 9.3005
R15738 gnd.n5294 gnd.n4694 9.3005
R15739 gnd.n5296 gnd.n5295 9.3005
R15740 gnd.n5297 gnd.n4677 9.3005
R15741 gnd.n5315 gnd.n5314 9.3005
R15742 gnd.n5317 gnd.n4662 9.3005
R15743 gnd.n5348 gnd.n4664 9.3005
R15744 gnd.n5349 gnd.n4660 9.3005
R15745 gnd.n5351 gnd.n5350 9.3005
R15746 gnd.n4648 gnd.n4643 9.3005
R15747 gnd.n5372 gnd.n4642 9.3005
R15748 gnd.n5375 gnd.n5374 9.3005
R15749 gnd.n5377 gnd.n5376 9.3005
R15750 gnd.n5380 gnd.n4625 9.3005
R15751 gnd.n5378 gnd.n4623 9.3005
R15752 gnd.n5402 gnd.n4621 9.3005
R15753 gnd.n5404 gnd.n5403 9.3005
R15754 gnd.n4599 gnd.n4598 9.3005
R15755 gnd.n5449 gnd.n5448 9.3005
R15756 gnd.n5450 gnd.n4592 9.3005
R15757 gnd.n5458 gnd.n4591 9.3005
R15758 gnd.n5461 gnd.n5460 9.3005
R15759 gnd.n5463 gnd.n4589 9.3005
R15760 gnd.n5747 gnd.n5746 9.3005
R15761 gnd.n5745 gnd.n5464 9.3005
R15762 gnd.n5466 gnd.n5465 9.3005
R15763 gnd.n5741 gnd.n5467 9.3005
R15764 gnd.n5740 gnd.n5468 9.3005
R15765 gnd.n5739 gnd.n5726 9.3005
R15766 gnd.n5736 gnd.n5728 9.3005
R15767 gnd.n5735 gnd.n5729 9.3005
R15768 gnd.n5732 gnd.n5730 9.3005
R15769 gnd.n5731 gnd.n4518 9.3005
R15770 gnd.n5161 gnd.n5160 9.3005
R15771 gnd.n5836 gnd.n4519 9.3005
R15772 gnd.n5835 gnd.n4521 9.3005
R15773 gnd.n4525 gnd.n4522 9.3005
R15774 gnd.n5830 gnd.n4526 9.3005
R15775 gnd.n5829 gnd.n4527 9.3005
R15776 gnd.n5828 gnd.n4528 9.3005
R15777 gnd.n4532 gnd.n4529 9.3005
R15778 gnd.n5823 gnd.n4533 9.3005
R15779 gnd.n5822 gnd.n4534 9.3005
R15780 gnd.n5821 gnd.n4535 9.3005
R15781 gnd.n4539 gnd.n4536 9.3005
R15782 gnd.n5816 gnd.n4540 9.3005
R15783 gnd.n5815 gnd.n4541 9.3005
R15784 gnd.n5814 gnd.n4542 9.3005
R15785 gnd.n4546 gnd.n4543 9.3005
R15786 gnd.n5809 gnd.n4547 9.3005
R15787 gnd.n5808 gnd.n4548 9.3005
R15788 gnd.n5807 gnd.n4549 9.3005
R15789 gnd.n4553 gnd.n4550 9.3005
R15790 gnd.n5802 gnd.n4554 9.3005
R15791 gnd.n5801 gnd.n4555 9.3005
R15792 gnd.n5800 gnd.n4556 9.3005
R15793 gnd.n4563 gnd.n4561 9.3005
R15794 gnd.n5795 gnd.n4564 9.3005
R15795 gnd.n5794 gnd.n4565 9.3005
R15796 gnd.n5793 gnd.n5790 9.3005
R15797 gnd.n5838 gnd.n5837 9.3005
R15798 gnd.n4670 gnd.n4669 9.3005
R15799 gnd.n5325 gnd.n5324 9.3005
R15800 gnd.n5326 gnd.n4668 9.3005
R15801 gnd.n5343 gnd.n5327 9.3005
R15802 gnd.n5342 gnd.n5328 9.3005
R15803 gnd.n5341 gnd.n5329 9.3005
R15804 gnd.n5339 gnd.n5330 9.3005
R15805 gnd.n5338 gnd.n5331 9.3005
R15806 gnd.n5336 gnd.n5332 9.3005
R15807 gnd.n5335 gnd.n5333 9.3005
R15808 gnd.n4614 gnd.n4613 9.3005
R15809 gnd.n5412 gnd.n5411 9.3005
R15810 gnd.n5413 gnd.n4612 9.3005
R15811 gnd.n5427 gnd.n5414 9.3005
R15812 gnd.n5426 gnd.n5415 9.3005
R15813 gnd.n5425 gnd.n5416 9.3005
R15814 gnd.n5423 gnd.n5417 9.3005
R15815 gnd.n5422 gnd.n5418 9.3005
R15816 gnd.n5420 gnd.n5419 9.3005
R15817 gnd.n4571 gnd.n4570 9.3005
R15818 gnd.n5771 gnd.n5770 9.3005
R15819 gnd.n5772 gnd.n4569 9.3005
R15820 gnd.n5776 gnd.n5773 9.3005
R15821 gnd.n5777 gnd.n4568 9.3005
R15822 gnd.n5781 gnd.n5780 9.3005
R15823 gnd.n5782 gnd.n4567 9.3005
R15824 gnd.n5784 gnd.n5783 9.3005
R15825 gnd.n5787 gnd.n4566 9.3005
R15826 gnd.n5789 gnd.n5788 9.3005
R15827 gnd.n4997 gnd.n4996 9.3005
R15828 gnd.n4887 gnd.n4886 9.3005
R15829 gnd.n5011 gnd.n5010 9.3005
R15830 gnd.n5012 gnd.n4885 9.3005
R15831 gnd.n5014 gnd.n5013 9.3005
R15832 gnd.n4875 gnd.n4874 9.3005
R15833 gnd.n5027 gnd.n5026 9.3005
R15834 gnd.n5028 gnd.n4873 9.3005
R15835 gnd.n5134 gnd.n5029 9.3005
R15836 gnd.n5133 gnd.n5030 9.3005
R15837 gnd.n5132 gnd.n5031 9.3005
R15838 gnd.n5131 gnd.n5032 9.3005
R15839 gnd.n5128 gnd.n5033 9.3005
R15840 gnd.n5127 gnd.n5034 9.3005
R15841 gnd.n5126 gnd.n5035 9.3005
R15842 gnd.n5124 gnd.n5036 9.3005
R15843 gnd.n5123 gnd.n5037 9.3005
R15844 gnd.n5120 gnd.n5038 9.3005
R15845 gnd.n5119 gnd.n5039 9.3005
R15846 gnd.n5118 gnd.n5040 9.3005
R15847 gnd.n5116 gnd.n5041 9.3005
R15848 gnd.n5115 gnd.n5042 9.3005
R15849 gnd.n5111 gnd.n5043 9.3005
R15850 gnd.n5110 gnd.n5044 9.3005
R15851 gnd.n5109 gnd.n5045 9.3005
R15852 gnd.n5107 gnd.n5046 9.3005
R15853 gnd.n5106 gnd.n5047 9.3005
R15854 gnd.n5103 gnd.n5048 9.3005
R15855 gnd.n4995 gnd.n4896 9.3005
R15856 gnd.n4898 gnd.n4897 9.3005
R15857 gnd.n4942 gnd.n4940 9.3005
R15858 gnd.n4943 gnd.n4939 9.3005
R15859 gnd.n4946 gnd.n4935 9.3005
R15860 gnd.n4947 gnd.n4934 9.3005
R15861 gnd.n4950 gnd.n4933 9.3005
R15862 gnd.n4951 gnd.n4932 9.3005
R15863 gnd.n4954 gnd.n4931 9.3005
R15864 gnd.n4955 gnd.n4930 9.3005
R15865 gnd.n4958 gnd.n4929 9.3005
R15866 gnd.n4959 gnd.n4928 9.3005
R15867 gnd.n4962 gnd.n4927 9.3005
R15868 gnd.n4963 gnd.n4926 9.3005
R15869 gnd.n4966 gnd.n4925 9.3005
R15870 gnd.n4967 gnd.n4924 9.3005
R15871 gnd.n4970 gnd.n4923 9.3005
R15872 gnd.n4971 gnd.n4922 9.3005
R15873 gnd.n4974 gnd.n4921 9.3005
R15874 gnd.n4975 gnd.n4920 9.3005
R15875 gnd.n4978 gnd.n4919 9.3005
R15876 gnd.n4979 gnd.n4918 9.3005
R15877 gnd.n4982 gnd.n4917 9.3005
R15878 gnd.n4984 gnd.n4916 9.3005
R15879 gnd.n4985 gnd.n4915 9.3005
R15880 gnd.n4986 gnd.n4914 9.3005
R15881 gnd.n4987 gnd.n4913 9.3005
R15882 gnd.n4994 gnd.n4993 9.3005
R15883 gnd.n5003 gnd.n5002 9.3005
R15884 gnd.n5004 gnd.n4890 9.3005
R15885 gnd.n5006 gnd.n5005 9.3005
R15886 gnd.n4881 gnd.n4880 9.3005
R15887 gnd.n5019 gnd.n5018 9.3005
R15888 gnd.n5020 gnd.n4879 9.3005
R15889 gnd.n5022 gnd.n5021 9.3005
R15890 gnd.n4868 gnd.n4867 9.3005
R15891 gnd.n5139 gnd.n5138 9.3005
R15892 gnd.n5140 gnd.n4822 9.3005
R15893 gnd.n5144 gnd.n5142 9.3005
R15894 gnd.n5143 gnd.n4801 9.3005
R15895 gnd.n5162 gnd.n4800 9.3005
R15896 gnd.n5165 gnd.n5164 9.3005
R15897 gnd.n4794 gnd.n4793 9.3005
R15898 gnd.n5176 gnd.n5174 9.3005
R15899 gnd.n5175 gnd.n4775 9.3005
R15900 gnd.n5193 gnd.n4774 9.3005
R15901 gnd.n5196 gnd.n5195 9.3005
R15902 gnd.n4768 gnd.n4767 9.3005
R15903 gnd.n5207 gnd.n5205 9.3005
R15904 gnd.n5206 gnd.n4751 9.3005
R15905 gnd.n5224 gnd.n4750 9.3005
R15906 gnd.n5227 gnd.n5226 9.3005
R15907 gnd.n4743 gnd.n4742 9.3005
R15908 gnd.n5238 gnd.n5236 9.3005
R15909 gnd.n5237 gnd.n4725 9.3005
R15910 gnd.n5255 gnd.n4724 9.3005
R15911 gnd.n5258 gnd.n5257 9.3005
R15912 gnd.n4717 gnd.n4716 9.3005
R15913 gnd.n5269 gnd.n5267 9.3005
R15914 gnd.n5268 gnd.n4700 9.3005
R15915 gnd.n5286 gnd.n4699 9.3005
R15916 gnd.n5289 gnd.n5288 9.3005
R15917 gnd.n4692 gnd.n4691 9.3005
R15918 gnd.n5299 gnd.n5298 9.3005
R15919 gnd.n4676 gnd.n4675 9.3005
R15920 gnd.n5320 gnd.n5316 9.3005
R15921 gnd.n5319 gnd.n5318 9.3005
R15922 gnd.n4663 gnd.n4659 9.3005
R15923 gnd.n5353 gnd.n5352 9.3005
R15924 gnd.n4661 gnd.n4644 9.3005
R15925 gnd.n5371 gnd.n5370 9.3005
R15926 gnd.n5373 gnd.n4640 9.3005
R15927 gnd.n5383 gnd.n4641 9.3005
R15928 gnd.n5382 gnd.n5381 9.3005
R15929 gnd.n5379 gnd.n4619 9.3005
R15930 gnd.n5407 gnd.n4620 9.3005
R15931 gnd.n5406 gnd.n5405 9.3005
R15932 gnd.n4622 gnd.n4600 9.3005
R15933 gnd.n5446 gnd.n5445 9.3005
R15934 gnd.n5447 gnd.n4593 9.3005
R15935 gnd.n5457 gnd.n5456 9.3005
R15936 gnd.n5459 gnd.n4587 9.3005
R15937 gnd.n5750 gnd.n4588 9.3005
R15938 gnd.n5749 gnd.n5748 9.3005
R15939 gnd.n4590 gnd.n770 9.3005
R15940 gnd.n5893 gnd.n771 9.3005
R15941 gnd.n5892 gnd.n772 9.3005
R15942 gnd.n5891 gnd.n773 9.3005
R15943 gnd.n5725 gnd.n774 9.3005
R15944 gnd.n5727 gnd.n794 9.3005
R15945 gnd.n5879 gnd.n795 9.3005
R15946 gnd.n5878 gnd.n796 9.3005
R15947 gnd.n5877 gnd.n797 9.3005
R15948 gnd.n4892 gnd.n4891 9.3005
R15949 gnd.n6068 gnd.n6067 9.3005
R15950 gnd.n6069 gnd.n594 9.3005
R15951 gnd.n6071 gnd.n6070 9.3005
R15952 gnd.n590 gnd.n589 9.3005
R15953 gnd.n6078 gnd.n6077 9.3005
R15954 gnd.n6079 gnd.n588 9.3005
R15955 gnd.n6081 gnd.n6080 9.3005
R15956 gnd.n584 gnd.n583 9.3005
R15957 gnd.n6088 gnd.n6087 9.3005
R15958 gnd.n6089 gnd.n582 9.3005
R15959 gnd.n6091 gnd.n6090 9.3005
R15960 gnd.n578 gnd.n577 9.3005
R15961 gnd.n6098 gnd.n6097 9.3005
R15962 gnd.n6099 gnd.n576 9.3005
R15963 gnd.n6101 gnd.n6100 9.3005
R15964 gnd.n572 gnd.n571 9.3005
R15965 gnd.n6108 gnd.n6107 9.3005
R15966 gnd.n6109 gnd.n570 9.3005
R15967 gnd.n6111 gnd.n6110 9.3005
R15968 gnd.n566 gnd.n565 9.3005
R15969 gnd.n6118 gnd.n6117 9.3005
R15970 gnd.n6119 gnd.n564 9.3005
R15971 gnd.n6121 gnd.n6120 9.3005
R15972 gnd.n560 gnd.n559 9.3005
R15973 gnd.n6128 gnd.n6127 9.3005
R15974 gnd.n6129 gnd.n558 9.3005
R15975 gnd.n6131 gnd.n6130 9.3005
R15976 gnd.n554 gnd.n553 9.3005
R15977 gnd.n6138 gnd.n6137 9.3005
R15978 gnd.n6139 gnd.n552 9.3005
R15979 gnd.n6141 gnd.n6140 9.3005
R15980 gnd.n548 gnd.n547 9.3005
R15981 gnd.n6148 gnd.n6147 9.3005
R15982 gnd.n6149 gnd.n546 9.3005
R15983 gnd.n6151 gnd.n6150 9.3005
R15984 gnd.n542 gnd.n541 9.3005
R15985 gnd.n6158 gnd.n6157 9.3005
R15986 gnd.n6159 gnd.n540 9.3005
R15987 gnd.n6161 gnd.n6160 9.3005
R15988 gnd.n536 gnd.n535 9.3005
R15989 gnd.n6168 gnd.n6167 9.3005
R15990 gnd.n6169 gnd.n534 9.3005
R15991 gnd.n6171 gnd.n6170 9.3005
R15992 gnd.n530 gnd.n529 9.3005
R15993 gnd.n6178 gnd.n6177 9.3005
R15994 gnd.n6179 gnd.n528 9.3005
R15995 gnd.n6181 gnd.n6180 9.3005
R15996 gnd.n524 gnd.n523 9.3005
R15997 gnd.n6188 gnd.n6187 9.3005
R15998 gnd.n6189 gnd.n522 9.3005
R15999 gnd.n6191 gnd.n6190 9.3005
R16000 gnd.n518 gnd.n517 9.3005
R16001 gnd.n6198 gnd.n6197 9.3005
R16002 gnd.n6199 gnd.n516 9.3005
R16003 gnd.n6201 gnd.n6200 9.3005
R16004 gnd.n512 gnd.n511 9.3005
R16005 gnd.n6208 gnd.n6207 9.3005
R16006 gnd.n6209 gnd.n510 9.3005
R16007 gnd.n6211 gnd.n6210 9.3005
R16008 gnd.n506 gnd.n505 9.3005
R16009 gnd.n6218 gnd.n6217 9.3005
R16010 gnd.n6219 gnd.n504 9.3005
R16011 gnd.n6221 gnd.n6220 9.3005
R16012 gnd.n500 gnd.n499 9.3005
R16013 gnd.n6228 gnd.n6227 9.3005
R16014 gnd.n6229 gnd.n498 9.3005
R16015 gnd.n6231 gnd.n6230 9.3005
R16016 gnd.n494 gnd.n493 9.3005
R16017 gnd.n6238 gnd.n6237 9.3005
R16018 gnd.n6239 gnd.n492 9.3005
R16019 gnd.n6241 gnd.n6240 9.3005
R16020 gnd.n488 gnd.n487 9.3005
R16021 gnd.n6248 gnd.n6247 9.3005
R16022 gnd.n6249 gnd.n486 9.3005
R16023 gnd.n6251 gnd.n6250 9.3005
R16024 gnd.n482 gnd.n481 9.3005
R16025 gnd.n6258 gnd.n6257 9.3005
R16026 gnd.n6259 gnd.n480 9.3005
R16027 gnd.n6261 gnd.n6260 9.3005
R16028 gnd.n476 gnd.n475 9.3005
R16029 gnd.n6268 gnd.n6267 9.3005
R16030 gnd.n6269 gnd.n474 9.3005
R16031 gnd.n6271 gnd.n6270 9.3005
R16032 gnd.n470 gnd.n469 9.3005
R16033 gnd.n6278 gnd.n6277 9.3005
R16034 gnd.n6279 gnd.n468 9.3005
R16035 gnd.n6281 gnd.n6280 9.3005
R16036 gnd.n464 gnd.n463 9.3005
R16037 gnd.n6288 gnd.n6287 9.3005
R16038 gnd.n6289 gnd.n462 9.3005
R16039 gnd.n6291 gnd.n6290 9.3005
R16040 gnd.n458 gnd.n457 9.3005
R16041 gnd.n6298 gnd.n6297 9.3005
R16042 gnd.n6299 gnd.n456 9.3005
R16043 gnd.n6301 gnd.n6300 9.3005
R16044 gnd.n452 gnd.n451 9.3005
R16045 gnd.n6308 gnd.n6307 9.3005
R16046 gnd.n6309 gnd.n450 9.3005
R16047 gnd.n6311 gnd.n6310 9.3005
R16048 gnd.n446 gnd.n445 9.3005
R16049 gnd.n6318 gnd.n6317 9.3005
R16050 gnd.n6319 gnd.n444 9.3005
R16051 gnd.n6321 gnd.n6320 9.3005
R16052 gnd.n440 gnd.n439 9.3005
R16053 gnd.n6328 gnd.n6327 9.3005
R16054 gnd.n6329 gnd.n438 9.3005
R16055 gnd.n6331 gnd.n6330 9.3005
R16056 gnd.n434 gnd.n433 9.3005
R16057 gnd.n6338 gnd.n6337 9.3005
R16058 gnd.n6339 gnd.n432 9.3005
R16059 gnd.n6341 gnd.n6340 9.3005
R16060 gnd.n428 gnd.n427 9.3005
R16061 gnd.n6348 gnd.n6347 9.3005
R16062 gnd.n6349 gnd.n426 9.3005
R16063 gnd.n6351 gnd.n6350 9.3005
R16064 gnd.n422 gnd.n421 9.3005
R16065 gnd.n6358 gnd.n6357 9.3005
R16066 gnd.n6359 gnd.n420 9.3005
R16067 gnd.n6361 gnd.n6360 9.3005
R16068 gnd.n416 gnd.n415 9.3005
R16069 gnd.n6368 gnd.n6367 9.3005
R16070 gnd.n6369 gnd.n414 9.3005
R16071 gnd.n6371 gnd.n6370 9.3005
R16072 gnd.n410 gnd.n409 9.3005
R16073 gnd.n6378 gnd.n6377 9.3005
R16074 gnd.n6379 gnd.n408 9.3005
R16075 gnd.n6381 gnd.n6380 9.3005
R16076 gnd.n404 gnd.n403 9.3005
R16077 gnd.n6388 gnd.n6387 9.3005
R16078 gnd.n6389 gnd.n402 9.3005
R16079 gnd.n6391 gnd.n6390 9.3005
R16080 gnd.n398 gnd.n397 9.3005
R16081 gnd.n6398 gnd.n6397 9.3005
R16082 gnd.n6399 gnd.n396 9.3005
R16083 gnd.n6401 gnd.n6400 9.3005
R16084 gnd.n392 gnd.n391 9.3005
R16085 gnd.n6408 gnd.n6407 9.3005
R16086 gnd.n6409 gnd.n390 9.3005
R16087 gnd.n6412 gnd.n6411 9.3005
R16088 gnd.n6410 gnd.n386 9.3005
R16089 gnd.n6418 gnd.n385 9.3005
R16090 gnd.n6420 gnd.n6419 9.3005
R16091 gnd.n381 gnd.n380 9.3005
R16092 gnd.n6429 gnd.n6428 9.3005
R16093 gnd.n6430 gnd.n379 9.3005
R16094 gnd.n6432 gnd.n6431 9.3005
R16095 gnd.n375 gnd.n374 9.3005
R16096 gnd.n6439 gnd.n6438 9.3005
R16097 gnd.n6440 gnd.n373 9.3005
R16098 gnd.n6442 gnd.n6441 9.3005
R16099 gnd.n369 gnd.n368 9.3005
R16100 gnd.n6449 gnd.n6448 9.3005
R16101 gnd.n6450 gnd.n367 9.3005
R16102 gnd.n6452 gnd.n6451 9.3005
R16103 gnd.n363 gnd.n362 9.3005
R16104 gnd.n6459 gnd.n6458 9.3005
R16105 gnd.n6460 gnd.n361 9.3005
R16106 gnd.n6462 gnd.n6461 9.3005
R16107 gnd.n357 gnd.n356 9.3005
R16108 gnd.n6469 gnd.n6468 9.3005
R16109 gnd.n6470 gnd.n355 9.3005
R16110 gnd.n6472 gnd.n6471 9.3005
R16111 gnd.n351 gnd.n350 9.3005
R16112 gnd.n6479 gnd.n6478 9.3005
R16113 gnd.n6480 gnd.n349 9.3005
R16114 gnd.n6482 gnd.n6481 9.3005
R16115 gnd.n345 gnd.n344 9.3005
R16116 gnd.n6489 gnd.n6488 9.3005
R16117 gnd.n6490 gnd.n343 9.3005
R16118 gnd.n6492 gnd.n6491 9.3005
R16119 gnd.n339 gnd.n338 9.3005
R16120 gnd.n6499 gnd.n6498 9.3005
R16121 gnd.n6500 gnd.n337 9.3005
R16122 gnd.n6502 gnd.n6501 9.3005
R16123 gnd.n333 gnd.n332 9.3005
R16124 gnd.n6509 gnd.n6508 9.3005
R16125 gnd.n6510 gnd.n331 9.3005
R16126 gnd.n6512 gnd.n6511 9.3005
R16127 gnd.n327 gnd.n326 9.3005
R16128 gnd.n6519 gnd.n6518 9.3005
R16129 gnd.n6520 gnd.n325 9.3005
R16130 gnd.n6522 gnd.n6521 9.3005
R16131 gnd.n321 gnd.n320 9.3005
R16132 gnd.n6529 gnd.n6528 9.3005
R16133 gnd.n6530 gnd.n319 9.3005
R16134 gnd.n6532 gnd.n6531 9.3005
R16135 gnd.n315 gnd.n314 9.3005
R16136 gnd.n6539 gnd.n6538 9.3005
R16137 gnd.n6540 gnd.n313 9.3005
R16138 gnd.n6542 gnd.n6541 9.3005
R16139 gnd.n309 gnd.n308 9.3005
R16140 gnd.n6549 gnd.n6548 9.3005
R16141 gnd.n6550 gnd.n307 9.3005
R16142 gnd.n6552 gnd.n6551 9.3005
R16143 gnd.n303 gnd.n302 9.3005
R16144 gnd.n6559 gnd.n6558 9.3005
R16145 gnd.n6560 gnd.n301 9.3005
R16146 gnd.n6562 gnd.n6561 9.3005
R16147 gnd.n297 gnd.n296 9.3005
R16148 gnd.n6569 gnd.n6568 9.3005
R16149 gnd.n6570 gnd.n295 9.3005
R16150 gnd.n6572 gnd.n6571 9.3005
R16151 gnd.n291 gnd.n290 9.3005
R16152 gnd.n6579 gnd.n6578 9.3005
R16153 gnd.n6580 gnd.n289 9.3005
R16154 gnd.n6582 gnd.n6581 9.3005
R16155 gnd.n285 gnd.n284 9.3005
R16156 gnd.n6589 gnd.n6588 9.3005
R16157 gnd.n6590 gnd.n283 9.3005
R16158 gnd.n6592 gnd.n6591 9.3005
R16159 gnd.n279 gnd.n278 9.3005
R16160 gnd.n6599 gnd.n6598 9.3005
R16161 gnd.n6600 gnd.n277 9.3005
R16162 gnd.n6602 gnd.n6601 9.3005
R16163 gnd.n273 gnd.n272 9.3005
R16164 gnd.n6609 gnd.n6608 9.3005
R16165 gnd.n6610 gnd.n271 9.3005
R16166 gnd.n6612 gnd.n6611 9.3005
R16167 gnd.n267 gnd.n266 9.3005
R16168 gnd.n6619 gnd.n6618 9.3005
R16169 gnd.n6620 gnd.n265 9.3005
R16170 gnd.n6622 gnd.n6621 9.3005
R16171 gnd.n261 gnd.n260 9.3005
R16172 gnd.n6630 gnd.n6629 9.3005
R16173 gnd.n6631 gnd.n259 9.3005
R16174 gnd.n6634 gnd.n6633 9.3005
R16175 gnd.n6422 gnd.n6421 9.3005
R16176 gnd.n6875 gnd.n89 9.3005
R16177 gnd.n6874 gnd.n91 9.3005
R16178 gnd.n95 gnd.n92 9.3005
R16179 gnd.n6869 gnd.n96 9.3005
R16180 gnd.n6868 gnd.n97 9.3005
R16181 gnd.n6867 gnd.n98 9.3005
R16182 gnd.n102 gnd.n99 9.3005
R16183 gnd.n6862 gnd.n103 9.3005
R16184 gnd.n6861 gnd.n104 9.3005
R16185 gnd.n6860 gnd.n105 9.3005
R16186 gnd.n109 gnd.n106 9.3005
R16187 gnd.n6855 gnd.n110 9.3005
R16188 gnd.n6854 gnd.n111 9.3005
R16189 gnd.n6853 gnd.n112 9.3005
R16190 gnd.n116 gnd.n113 9.3005
R16191 gnd.n6848 gnd.n117 9.3005
R16192 gnd.n6847 gnd.n118 9.3005
R16193 gnd.n6843 gnd.n119 9.3005
R16194 gnd.n123 gnd.n120 9.3005
R16195 gnd.n6838 gnd.n124 9.3005
R16196 gnd.n6837 gnd.n125 9.3005
R16197 gnd.n6836 gnd.n126 9.3005
R16198 gnd.n130 gnd.n127 9.3005
R16199 gnd.n6831 gnd.n131 9.3005
R16200 gnd.n6830 gnd.n132 9.3005
R16201 gnd.n6829 gnd.n133 9.3005
R16202 gnd.n137 gnd.n134 9.3005
R16203 gnd.n6824 gnd.n138 9.3005
R16204 gnd.n6823 gnd.n139 9.3005
R16205 gnd.n6822 gnd.n140 9.3005
R16206 gnd.n144 gnd.n141 9.3005
R16207 gnd.n6817 gnd.n145 9.3005
R16208 gnd.n6816 gnd.n146 9.3005
R16209 gnd.n6815 gnd.n147 9.3005
R16210 gnd.n151 gnd.n148 9.3005
R16211 gnd.n6810 gnd.n152 9.3005
R16212 gnd.n6809 gnd.n6808 9.3005
R16213 gnd.n6807 gnd.n155 9.3005
R16214 gnd.n6877 gnd.n6876 9.3005
R16215 gnd.n3888 gnd.n3887 9.3005
R16216 gnd.n1330 gnd.n1329 9.3005
R16217 gnd.n3902 gnd.n3901 9.3005
R16218 gnd.n3903 gnd.n1328 9.3005
R16219 gnd.n3990 gnd.n3904 9.3005
R16220 gnd.n3989 gnd.n3905 9.3005
R16221 gnd.n3988 gnd.n3906 9.3005
R16222 gnd.n3986 gnd.n3907 9.3005
R16223 gnd.n3985 gnd.n3908 9.3005
R16224 gnd.n3984 gnd.n3909 9.3005
R16225 gnd.n3982 gnd.n3910 9.3005
R16226 gnd.n3981 gnd.n3911 9.3005
R16227 gnd.n3979 gnd.n3912 9.3005
R16228 gnd.n3978 gnd.n3913 9.3005
R16229 gnd.n3977 gnd.n3914 9.3005
R16230 gnd.n3975 gnd.n3915 9.3005
R16231 gnd.n3974 gnd.n3916 9.3005
R16232 gnd.n3971 gnd.n3917 9.3005
R16233 gnd.n3970 gnd.n3918 9.3005
R16234 gnd.n3969 gnd.n3919 9.3005
R16235 gnd.n3968 gnd.n240 9.3005
R16236 gnd.n3964 gnd.n3920 9.3005
R16237 gnd.n3963 gnd.n3921 9.3005
R16238 gnd.n3961 gnd.n3922 9.3005
R16239 gnd.n3960 gnd.n3923 9.3005
R16240 gnd.n3958 gnd.n3924 9.3005
R16241 gnd.n3957 gnd.n3925 9.3005
R16242 gnd.n3955 gnd.n3926 9.3005
R16243 gnd.n3954 gnd.n3927 9.3005
R16244 gnd.n3952 gnd.n3928 9.3005
R16245 gnd.n3951 gnd.n3929 9.3005
R16246 gnd.n3949 gnd.n3930 9.3005
R16247 gnd.n3948 gnd.n3931 9.3005
R16248 gnd.n3946 gnd.n3932 9.3005
R16249 gnd.n3945 gnd.n3933 9.3005
R16250 gnd.n3943 gnd.n3934 9.3005
R16251 gnd.n3942 gnd.n3935 9.3005
R16252 gnd.n3940 gnd.n3936 9.3005
R16253 gnd.n3939 gnd.n3938 9.3005
R16254 gnd.n3937 gnd.n159 9.3005
R16255 gnd.n6804 gnd.n158 9.3005
R16256 gnd.n6806 gnd.n6805 9.3005
R16257 gnd.n3886 gnd.n1335 9.3005
R16258 gnd.n3875 gnd.n1340 9.3005
R16259 gnd.n3877 gnd.n3876 9.3005
R16260 gnd.n3874 gnd.n1342 9.3005
R16261 gnd.n3873 gnd.n3872 9.3005
R16262 gnd.n1344 gnd.n1343 9.3005
R16263 gnd.n3866 gnd.n3865 9.3005
R16264 gnd.n3864 gnd.n1346 9.3005
R16265 gnd.n3863 gnd.n3862 9.3005
R16266 gnd.n1348 gnd.n1347 9.3005
R16267 gnd.n3856 gnd.n3855 9.3005
R16268 gnd.n3854 gnd.n1350 9.3005
R16269 gnd.n3853 gnd.n3852 9.3005
R16270 gnd.n1352 gnd.n1351 9.3005
R16271 gnd.n3846 gnd.n3845 9.3005
R16272 gnd.n3844 gnd.n1354 9.3005
R16273 gnd.n3843 gnd.n3842 9.3005
R16274 gnd.n1356 gnd.n1355 9.3005
R16275 gnd.n3836 gnd.n3835 9.3005
R16276 gnd.n3834 gnd.n1358 9.3005
R16277 gnd.n1360 gnd.n1359 9.3005
R16278 gnd.n3821 gnd.n3776 9.3005
R16279 gnd.n3823 gnd.n3822 9.3005
R16280 gnd.n3820 gnd.n3778 9.3005
R16281 gnd.n3819 gnd.n3818 9.3005
R16282 gnd.n3780 gnd.n3779 9.3005
R16283 gnd.n3812 gnd.n3811 9.3005
R16284 gnd.n3810 gnd.n3782 9.3005
R16285 gnd.n3809 gnd.n3808 9.3005
R16286 gnd.n3784 gnd.n3783 9.3005
R16287 gnd.n3802 gnd.n3801 9.3005
R16288 gnd.n3800 gnd.n3786 9.3005
R16289 gnd.n3799 gnd.n3798 9.3005
R16290 gnd.n3788 gnd.n3787 9.3005
R16291 gnd.n3792 gnd.n3791 9.3005
R16292 gnd.n3790 gnd.n3789 9.3005
R16293 gnd.n1339 gnd.n1336 9.3005
R16294 gnd.n3885 gnd.n3884 9.3005
R16295 gnd.n4127 gnd.n1220 9.3005
R16296 gnd.n4126 gnd.n1221 9.3005
R16297 gnd.n1324 gnd.n1222 9.3005
R16298 gnd.n4013 gnd.n4012 9.3005
R16299 gnd.n4014 gnd.n1323 9.3005
R16300 gnd.n4018 gnd.n4015 9.3005
R16301 gnd.n4017 gnd.n4016 9.3005
R16302 gnd.n1297 gnd.n1296 9.3005
R16303 gnd.n4044 gnd.n4043 9.3005
R16304 gnd.n4045 gnd.n1295 9.3005
R16305 gnd.n4050 gnd.n4046 9.3005
R16306 gnd.n4049 gnd.n4048 9.3005
R16307 gnd.n4047 gnd.n1267 9.3005
R16308 gnd.n4082 gnd.n1268 9.3005
R16309 gnd.n4083 gnd.n212 9.3005
R16310 gnd.n6675 gnd.n211 9.3005
R16311 gnd.n6677 gnd.n6676 9.3005
R16312 gnd.n199 gnd.n198 9.3005
R16313 gnd.n6690 gnd.n6689 9.3005
R16314 gnd.n6691 gnd.n197 9.3005
R16315 gnd.n6693 gnd.n6692 9.3005
R16316 gnd.n183 gnd.n182 9.3005
R16317 gnd.n6706 gnd.n6705 9.3005
R16318 gnd.n6707 gnd.n181 9.3005
R16319 gnd.n6709 gnd.n6708 9.3005
R16320 gnd.n167 gnd.n166 9.3005
R16321 gnd.n6796 gnd.n6795 9.3005
R16322 gnd.n6797 gnd.n165 9.3005
R16323 gnd.n6799 gnd.n6798 9.3005
R16324 gnd.n88 gnd.n87 9.3005
R16325 gnd.n6879 gnd.n6878 9.3005
R16326 gnd.n4128 gnd.n1219 9.3005
R16327 gnd.n6674 gnd.n6673 9.3005
R16328 gnd.n4075 gnd.n4074 9.3005
R16329 gnd.n4073 gnd.n4071 9.3005
R16330 gnd.n4072 gnd.n253 9.3005
R16331 gnd.n6641 gnd.n254 9.3005
R16332 gnd.n6640 gnd.n255 9.3005
R16333 gnd.n6639 gnd.n256 9.3005
R16334 gnd.n6632 gnd.n257 9.3005
R16335 gnd.n2477 gnd.n2245 9.3005
R16336 gnd.n2499 gnd.n2478 9.3005
R16337 gnd.n2498 gnd.n2479 9.3005
R16338 gnd.n2497 gnd.n2480 9.3005
R16339 gnd.n2483 gnd.n2481 9.3005
R16340 gnd.n2493 gnd.n2484 9.3005
R16341 gnd.n2492 gnd.n2485 9.3005
R16342 gnd.n2491 gnd.n2486 9.3005
R16343 gnd.n2489 gnd.n2488 9.3005
R16344 gnd.n2487 gnd.n2220 9.3005
R16345 gnd.n2218 gnd.n2217 9.3005
R16346 gnd.n2560 gnd.n2559 9.3005
R16347 gnd.n2561 gnd.n2216 9.3005
R16348 gnd.n2563 gnd.n2562 9.3005
R16349 gnd.n2214 gnd.n2213 9.3005
R16350 gnd.n2568 gnd.n2567 9.3005
R16351 gnd.n2569 gnd.n2212 9.3005
R16352 gnd.n2571 gnd.n2570 9.3005
R16353 gnd.n2210 gnd.n2209 9.3005
R16354 gnd.n2580 gnd.n2579 9.3005
R16355 gnd.n2581 gnd.n2208 9.3005
R16356 gnd.n2583 gnd.n2582 9.3005
R16357 gnd.n2072 gnd.n2071 9.3005
R16358 gnd.n2593 gnd.n2592 9.3005
R16359 gnd.n2594 gnd.n2070 9.3005
R16360 gnd.n2596 gnd.n2595 9.3005
R16361 gnd.n2066 gnd.n2065 9.3005
R16362 gnd.n2608 gnd.n2607 9.3005
R16363 gnd.n2609 gnd.n2064 9.3005
R16364 gnd.n2621 gnd.n2610 9.3005
R16365 gnd.n2620 gnd.n2611 9.3005
R16366 gnd.n2619 gnd.n2612 9.3005
R16367 gnd.n2614 gnd.n2613 9.3005
R16368 gnd.n1772 gnd.n1771 9.3005
R16369 gnd.n2803 gnd.n2802 9.3005
R16370 gnd.n2804 gnd.n1770 9.3005
R16371 gnd.n2806 gnd.n2805 9.3005
R16372 gnd.n1744 gnd.n1743 9.3005
R16373 gnd.n2846 gnd.n2845 9.3005
R16374 gnd.n2847 gnd.n1742 9.3005
R16375 gnd.n2849 gnd.n2848 9.3005
R16376 gnd.n1726 gnd.n1725 9.3005
R16377 gnd.n2888 gnd.n2887 9.3005
R16378 gnd.n2889 gnd.n1724 9.3005
R16379 gnd.n2893 gnd.n2890 9.3005
R16380 gnd.n2892 gnd.n2891 9.3005
R16381 gnd.n1700 gnd.n1699 9.3005
R16382 gnd.n2950 gnd.n2949 9.3005
R16383 gnd.n2951 gnd.n1698 9.3005
R16384 gnd.n2953 gnd.n2952 9.3005
R16385 gnd.n1682 gnd.n1681 9.3005
R16386 gnd.n2977 gnd.n2976 9.3005
R16387 gnd.n2978 gnd.n1680 9.3005
R16388 gnd.n2982 gnd.n2979 9.3005
R16389 gnd.n2981 gnd.n2980 9.3005
R16390 gnd.n1649 gnd.n1648 9.3005
R16391 gnd.n3028 gnd.n3027 9.3005
R16392 gnd.n3029 gnd.n1647 9.3005
R16393 gnd.n3031 gnd.n3030 9.3005
R16394 gnd.n1626 gnd.n1625 9.3005
R16395 gnd.n3068 gnd.n3067 9.3005
R16396 gnd.n3069 gnd.n1624 9.3005
R16397 gnd.n3071 gnd.n3070 9.3005
R16398 gnd.n1604 gnd.n1603 9.3005
R16399 gnd.n3124 gnd.n3123 9.3005
R16400 gnd.n3125 gnd.n1602 9.3005
R16401 gnd.n3127 gnd.n3126 9.3005
R16402 gnd.n1585 gnd.n1584 9.3005
R16403 gnd.n3149 gnd.n3148 9.3005
R16404 gnd.n3150 gnd.n1583 9.3005
R16405 gnd.n3152 gnd.n3151 9.3005
R16406 gnd.n1565 gnd.n1564 9.3005
R16407 gnd.n3209 gnd.n3208 9.3005
R16408 gnd.n3210 gnd.n1563 9.3005
R16409 gnd.n3212 gnd.n3211 9.3005
R16410 gnd.n1543 gnd.n1542 9.3005
R16411 gnd.n3238 gnd.n3237 9.3005
R16412 gnd.n3239 gnd.n1541 9.3005
R16413 gnd.n3243 gnd.n3240 9.3005
R16414 gnd.n3242 gnd.n3241 9.3005
R16415 gnd.n1515 gnd.n1514 9.3005
R16416 gnd.n3291 gnd.n3290 9.3005
R16417 gnd.n3292 gnd.n1513 9.3005
R16418 gnd.n3294 gnd.n3293 9.3005
R16419 gnd.n1496 gnd.n1495 9.3005
R16420 gnd.n3318 gnd.n3317 9.3005
R16421 gnd.n3319 gnd.n1494 9.3005
R16422 gnd.n3323 gnd.n3320 9.3005
R16423 gnd.n3322 gnd.n3321 9.3005
R16424 gnd.n1466 gnd.n1465 9.3005
R16425 gnd.n3362 gnd.n3361 9.3005
R16426 gnd.n3363 gnd.n1464 9.3005
R16427 gnd.n3368 gnd.n3364 9.3005
R16428 gnd.n3367 gnd.n3366 9.3005
R16429 gnd.n3365 gnd.n1413 9.3005
R16430 gnd.n3610 gnd.n1414 9.3005
R16431 gnd.n3609 gnd.n1415 9.3005
R16432 gnd.n3608 gnd.n1416 9.3005
R16433 gnd.n1426 gnd.n1417 9.3005
R16434 gnd.n1427 gnd.n1425 9.3005
R16435 gnd.n3599 gnd.n1428 9.3005
R16436 gnd.n3598 gnd.n1429 9.3005
R16437 gnd.n3597 gnd.n1430 9.3005
R16438 gnd.n1433 gnd.n1432 9.3005
R16439 gnd.n1431 gnd.n1197 9.3005
R16440 gnd.n4143 gnd.n1198 9.3005
R16441 gnd.n4142 gnd.n1199 9.3005
R16442 gnd.n4141 gnd.n1200 9.3005
R16443 gnd.n1206 gnd.n1201 9.3005
R16444 gnd.n4135 gnd.n1207 9.3005
R16445 gnd.n4134 gnd.n1208 9.3005
R16446 gnd.n4133 gnd.n1209 9.3005
R16447 gnd.n3996 gnd.n1210 9.3005
R16448 gnd.n3998 gnd.n3997 9.3005
R16449 gnd.n4002 gnd.n4001 9.3005
R16450 gnd.n4003 gnd.n3995 9.3005
R16451 gnd.n4007 gnd.n4004 9.3005
R16452 gnd.n4006 gnd.n4005 9.3005
R16453 gnd.n1307 gnd.n1306 9.3005
R16454 gnd.n4033 gnd.n4032 9.3005
R16455 gnd.n4034 gnd.n1305 9.3005
R16456 gnd.n4038 gnd.n4035 9.3005
R16457 gnd.n4037 gnd.n4036 9.3005
R16458 gnd.n1279 gnd.n1278 9.3005
R16459 gnd.n4065 gnd.n4064 9.3005
R16460 gnd.n4066 gnd.n1277 9.3005
R16461 gnd.n4077 gnd.n4067 9.3005
R16462 gnd.n4076 gnd.n4068 9.3005
R16463 gnd.n2429 gnd.n2428 9.3005
R16464 gnd.n2295 gnd.n2270 9.3005
R16465 gnd.n2354 gnd.n2269 9.3005
R16466 gnd.n2356 gnd.n2355 9.3005
R16467 gnd.n2357 gnd.n2268 9.3005
R16468 gnd.n2359 gnd.n2358 9.3005
R16469 gnd.n2361 gnd.n2266 9.3005
R16470 gnd.n2363 gnd.n2362 9.3005
R16471 gnd.n2364 gnd.n2265 9.3005
R16472 gnd.n2366 gnd.n2365 9.3005
R16473 gnd.n2368 gnd.n2263 9.3005
R16474 gnd.n2370 gnd.n2369 9.3005
R16475 gnd.n2371 gnd.n2262 9.3005
R16476 gnd.n2373 gnd.n2372 9.3005
R16477 gnd.n2375 gnd.n2260 9.3005
R16478 gnd.n2377 gnd.n2376 9.3005
R16479 gnd.n2378 gnd.n2259 9.3005
R16480 gnd.n2422 gnd.n2379 9.3005
R16481 gnd.n2423 gnd.n2258 9.3005
R16482 gnd.n2426 gnd.n2425 9.3005
R16483 gnd.n2427 gnd.n2257 9.3005
R16484 gnd.n2297 gnd.n2296 9.3005
R16485 gnd.n2302 gnd.n2301 9.3005
R16486 gnd.n2305 gnd.n2290 9.3005
R16487 gnd.n2306 gnd.n2289 9.3005
R16488 gnd.n2309 gnd.n2288 9.3005
R16489 gnd.n2310 gnd.n2287 9.3005
R16490 gnd.n2313 gnd.n2286 9.3005
R16491 gnd.n2314 gnd.n2285 9.3005
R16492 gnd.n2317 gnd.n2284 9.3005
R16493 gnd.n2318 gnd.n2283 9.3005
R16494 gnd.n2321 gnd.n2282 9.3005
R16495 gnd.n2322 gnd.n2281 9.3005
R16496 gnd.n2325 gnd.n2280 9.3005
R16497 gnd.n2326 gnd.n2279 9.3005
R16498 gnd.n2329 gnd.n2278 9.3005
R16499 gnd.n2330 gnd.n2277 9.3005
R16500 gnd.n2333 gnd.n2276 9.3005
R16501 gnd.n2336 gnd.n2335 9.3005
R16502 gnd.n2300 gnd.n2294 9.3005
R16503 gnd.n2299 gnd.n2298 9.3005
R16504 gnd.n2343 gnd.n2342 9.3005
R16505 gnd.n2341 gnd.n2275 9.3005
R16506 gnd.n2340 gnd.n2339 9.3005
R16507 gnd.n2338 gnd.n901 9.3005
R16508 gnd.n4387 gnd.n902 9.3005
R16509 gnd.n4386 gnd.n903 9.3005
R16510 gnd.n4385 gnd.n904 9.3005
R16511 gnd.n920 gnd.n905 9.3005
R16512 gnd.n4375 gnd.n921 9.3005
R16513 gnd.n4374 gnd.n922 9.3005
R16514 gnd.n4373 gnd.n923 9.3005
R16515 gnd.n941 gnd.n924 9.3005
R16516 gnd.n4363 gnd.n942 9.3005
R16517 gnd.n4362 gnd.n943 9.3005
R16518 gnd.n4361 gnd.n944 9.3005
R16519 gnd.n964 gnd.n945 9.3005
R16520 gnd.n965 gnd.n963 9.3005
R16521 gnd.n4349 gnd.n966 9.3005
R16522 gnd.n4348 gnd.n967 9.3005
R16523 gnd.n4347 gnd.n968 9.3005
R16524 gnd.n2255 gnd.n969 9.3005
R16525 gnd.n4336 gnd.n982 9.3005
R16526 gnd.n4335 gnd.n983 9.3005
R16527 gnd.n4334 gnd.n984 9.3005
R16528 gnd.n1000 gnd.n985 9.3005
R16529 gnd.n4323 gnd.n1001 9.3005
R16530 gnd.n4322 gnd.n1002 9.3005
R16531 gnd.n4321 gnd.n1003 9.3005
R16532 gnd.n1020 gnd.n1004 9.3005
R16533 gnd.n4311 gnd.n1021 9.3005
R16534 gnd.n4310 gnd.n1022 9.3005
R16535 gnd.n4309 gnd.n1023 9.3005
R16536 gnd.n1042 gnd.n1024 9.3005
R16537 gnd.n4299 gnd.n1043 9.3005
R16538 gnd.n4298 gnd.n1044 9.3005
R16539 gnd.n4297 gnd.n1045 9.3005
R16540 gnd.n1063 gnd.n1046 9.3005
R16541 gnd.n4287 gnd.n1064 9.3005
R16542 gnd.n4286 gnd.n1065 9.3005
R16543 gnd.n4285 gnd.n1066 9.3005
R16544 gnd.n1084 gnd.n1067 9.3005
R16545 gnd.n4275 gnd.n4274 9.3005
R16546 gnd.n2337 gnd.n2274 9.3005
R16547 gnd.n1938 gnd.n1934 9.3005
R16548 gnd.n1971 gnd.n1968 9.3005
R16549 gnd.n1972 gnd.n1967 9.3005
R16550 gnd.n1975 gnd.n1966 9.3005
R16551 gnd.n1976 gnd.n1965 9.3005
R16552 gnd.n1979 gnd.n1964 9.3005
R16553 gnd.n1980 gnd.n1963 9.3005
R16554 gnd.n1983 gnd.n1962 9.3005
R16555 gnd.n1984 gnd.n1961 9.3005
R16556 gnd.n1987 gnd.n1960 9.3005
R16557 gnd.n1988 gnd.n1959 9.3005
R16558 gnd.n1991 gnd.n1958 9.3005
R16559 gnd.n1992 gnd.n1957 9.3005
R16560 gnd.n1993 gnd.n1956 9.3005
R16561 gnd.n1955 gnd.n1952 9.3005
R16562 gnd.n1954 gnd.n1953 9.3005
R16563 gnd.n2704 gnd.n2703 9.3005
R16564 gnd.n1940 gnd.n1939 9.3005
R16565 gnd.n1999 gnd.n1997 9.3005
R16566 gnd.n2696 gnd.n2000 9.3005
R16567 gnd.n2695 gnd.n2001 9.3005
R16568 gnd.n2694 gnd.n2002 9.3005
R16569 gnd.n2006 gnd.n2003 9.3005
R16570 gnd.n2689 gnd.n2007 9.3005
R16571 gnd.n2688 gnd.n2008 9.3005
R16572 gnd.n2687 gnd.n2009 9.3005
R16573 gnd.n2013 gnd.n2010 9.3005
R16574 gnd.n2682 gnd.n2014 9.3005
R16575 gnd.n2681 gnd.n2015 9.3005
R16576 gnd.n2680 gnd.n2016 9.3005
R16577 gnd.n2020 gnd.n2017 9.3005
R16578 gnd.n2675 gnd.n2021 9.3005
R16579 gnd.n2674 gnd.n2022 9.3005
R16580 gnd.n2673 gnd.n2023 9.3005
R16581 gnd.n2028 gnd.n2026 9.3005
R16582 gnd.n2668 gnd.n2667 9.3005
R16583 gnd.n2705 gnd.n1933 9.3005
R16584 gnd.n4401 gnd.n4400 9.3005
R16585 gnd.n4399 gnd.n879 9.3005
R16586 gnd.n4398 gnd.n4397 9.3005
R16587 gnd.n881 gnd.n880 9.3005
R16588 gnd.n2391 gnd.n2390 9.3005
R16589 gnd.n2393 gnd.n2389 9.3005
R16590 gnd.n2395 gnd.n2394 9.3005
R16591 gnd.n2396 gnd.n2388 9.3005
R16592 gnd.n2398 gnd.n2397 9.3005
R16593 gnd.n2400 gnd.n2386 9.3005
R16594 gnd.n2402 gnd.n2401 9.3005
R16595 gnd.n2403 gnd.n2385 9.3005
R16596 gnd.n2405 gnd.n2404 9.3005
R16597 gnd.n2407 gnd.n2383 9.3005
R16598 gnd.n2409 gnd.n2408 9.3005
R16599 gnd.n2410 gnd.n2382 9.3005
R16600 gnd.n2418 gnd.n2411 9.3005
R16601 gnd.n2417 gnd.n2412 9.3005
R16602 gnd.n2416 gnd.n2414 9.3005
R16603 gnd.n2413 gnd.n2254 9.3005
R16604 gnd.n2433 gnd.n2256 9.3005
R16605 gnd.n2434 gnd.n2253 9.3005
R16606 gnd.n2436 gnd.n2435 9.3005
R16607 gnd.n2437 gnd.n2252 9.3005
R16608 gnd.n2443 gnd.n2438 9.3005
R16609 gnd.n2442 gnd.n2439 9.3005
R16610 gnd.n2441 gnd.n2440 9.3005
R16611 gnd.n2238 gnd.n2237 9.3005
R16612 gnd.n2513 gnd.n2512 9.3005
R16613 gnd.n2514 gnd.n2236 9.3005
R16614 gnd.n2516 gnd.n2515 9.3005
R16615 gnd.n2231 gnd.n2230 9.3005
R16616 gnd.n2529 gnd.n2528 9.3005
R16617 gnd.n2530 gnd.n2229 9.3005
R16618 gnd.n2532 gnd.n2531 9.3005
R16619 gnd.n2533 gnd.n2228 9.3005
R16620 gnd.n2537 gnd.n2536 9.3005
R16621 gnd.n2538 gnd.n2227 9.3005
R16622 gnd.n2541 gnd.n2540 9.3005
R16623 gnd.n2539 gnd.n2030 9.3005
R16624 gnd.n2664 gnd.n2029 9.3005
R16625 gnd.n2666 gnd.n2665 9.3005
R16626 gnd.n4402 gnd.n877 9.3005
R16627 gnd.n4409 gnd.n4408 9.3005
R16628 gnd.n4410 gnd.n871 9.3005
R16629 gnd.n4413 gnd.n870 9.3005
R16630 gnd.n4414 gnd.n869 9.3005
R16631 gnd.n4417 gnd.n868 9.3005
R16632 gnd.n4418 gnd.n867 9.3005
R16633 gnd.n4421 gnd.n866 9.3005
R16634 gnd.n4422 gnd.n865 9.3005
R16635 gnd.n4425 gnd.n864 9.3005
R16636 gnd.n4426 gnd.n863 9.3005
R16637 gnd.n4429 gnd.n862 9.3005
R16638 gnd.n4430 gnd.n861 9.3005
R16639 gnd.n4433 gnd.n860 9.3005
R16640 gnd.n4434 gnd.n859 9.3005
R16641 gnd.n4437 gnd.n858 9.3005
R16642 gnd.n4438 gnd.n857 9.3005
R16643 gnd.n4441 gnd.n856 9.3005
R16644 gnd.n4442 gnd.n855 9.3005
R16645 gnd.n4445 gnd.n854 9.3005
R16646 gnd.n4447 gnd.n851 9.3005
R16647 gnd.n4450 gnd.n850 9.3005
R16648 gnd.n4451 gnd.n849 9.3005
R16649 gnd.n4454 gnd.n848 9.3005
R16650 gnd.n4455 gnd.n847 9.3005
R16651 gnd.n4458 gnd.n846 9.3005
R16652 gnd.n4459 gnd.n845 9.3005
R16653 gnd.n4462 gnd.n844 9.3005
R16654 gnd.n4463 gnd.n843 9.3005
R16655 gnd.n4466 gnd.n842 9.3005
R16656 gnd.n4467 gnd.n841 9.3005
R16657 gnd.n4470 gnd.n840 9.3005
R16658 gnd.n4471 gnd.n839 9.3005
R16659 gnd.n4474 gnd.n838 9.3005
R16660 gnd.n4476 gnd.n837 9.3005
R16661 gnd.n4477 gnd.n836 9.3005
R16662 gnd.n4478 gnd.n835 9.3005
R16663 gnd.n4479 gnd.n834 9.3005
R16664 gnd.n4407 gnd.n876 9.3005
R16665 gnd.n4406 gnd.n4405 9.3005
R16666 gnd.n2349 gnd.n2348 9.3005
R16667 gnd.n2347 gnd.n890 9.3005
R16668 gnd.n4393 gnd.n891 9.3005
R16669 gnd.n4392 gnd.n892 9.3005
R16670 gnd.n4391 gnd.n893 9.3005
R16671 gnd.n911 gnd.n894 9.3005
R16672 gnd.n4381 gnd.n912 9.3005
R16673 gnd.n4380 gnd.n913 9.3005
R16674 gnd.n4379 gnd.n914 9.3005
R16675 gnd.n930 gnd.n915 9.3005
R16676 gnd.n4369 gnd.n931 9.3005
R16677 gnd.n4368 gnd.n932 9.3005
R16678 gnd.n4367 gnd.n933 9.3005
R16679 gnd.n951 gnd.n934 9.3005
R16680 gnd.n4357 gnd.n952 9.3005
R16681 gnd.n1010 gnd.n993 9.3005
R16682 gnd.n4317 gnd.n1011 9.3005
R16683 gnd.n4316 gnd.n1012 9.3005
R16684 gnd.n4315 gnd.n1013 9.3005
R16685 gnd.n1031 gnd.n1014 9.3005
R16686 gnd.n4305 gnd.n1032 9.3005
R16687 gnd.n4304 gnd.n1033 9.3005
R16688 gnd.n4303 gnd.n1034 9.3005
R16689 gnd.n1052 gnd.n1035 9.3005
R16690 gnd.n4293 gnd.n1053 9.3005
R16691 gnd.n4292 gnd.n1054 9.3005
R16692 gnd.n4291 gnd.n1055 9.3005
R16693 gnd.n1074 gnd.n1056 9.3005
R16694 gnd.n4281 gnd.n1075 9.3005
R16695 gnd.n4280 gnd.n1076 9.3005
R16696 gnd.n4279 gnd.n1077 9.3005
R16697 gnd.n2346 gnd.n2345 9.3005
R16698 gnd.n4327 gnd.n953 9.3005
R16699 gnd.n2458 gnd.n2457 9.3005
R16700 gnd.n2467 gnd.n2466 9.3005
R16701 gnd.n2469 gnd.n2456 9.3005
R16702 gnd.n2471 gnd.n2470 9.3005
R16703 gnd.n2247 gnd.n2246 9.3005
R16704 gnd.n2476 gnd.n2475 9.3005
R16705 gnd.n2461 gnd.n2460 9.3005
R16706 gnd.n5899 gnd.n762 9.3005
R16707 gnd.n5900 gnd.n761 9.3005
R16708 gnd.n5901 gnd.n760 9.3005
R16709 gnd.n759 gnd.n755 9.3005
R16710 gnd.n5907 gnd.n754 9.3005
R16711 gnd.n5908 gnd.n753 9.3005
R16712 gnd.n5909 gnd.n752 9.3005
R16713 gnd.n751 gnd.n747 9.3005
R16714 gnd.n5915 gnd.n746 9.3005
R16715 gnd.n5916 gnd.n745 9.3005
R16716 gnd.n5917 gnd.n744 9.3005
R16717 gnd.n743 gnd.n739 9.3005
R16718 gnd.n5923 gnd.n738 9.3005
R16719 gnd.n5924 gnd.n737 9.3005
R16720 gnd.n5925 gnd.n736 9.3005
R16721 gnd.n735 gnd.n731 9.3005
R16722 gnd.n5931 gnd.n730 9.3005
R16723 gnd.n5932 gnd.n729 9.3005
R16724 gnd.n5933 gnd.n728 9.3005
R16725 gnd.n727 gnd.n723 9.3005
R16726 gnd.n5939 gnd.n722 9.3005
R16727 gnd.n5940 gnd.n721 9.3005
R16728 gnd.n5941 gnd.n720 9.3005
R16729 gnd.n719 gnd.n715 9.3005
R16730 gnd.n5947 gnd.n714 9.3005
R16731 gnd.n5948 gnd.n713 9.3005
R16732 gnd.n5949 gnd.n712 9.3005
R16733 gnd.n711 gnd.n707 9.3005
R16734 gnd.n5955 gnd.n706 9.3005
R16735 gnd.n5956 gnd.n705 9.3005
R16736 gnd.n5957 gnd.n704 9.3005
R16737 gnd.n703 gnd.n699 9.3005
R16738 gnd.n5963 gnd.n698 9.3005
R16739 gnd.n5964 gnd.n697 9.3005
R16740 gnd.n5965 gnd.n696 9.3005
R16741 gnd.n695 gnd.n691 9.3005
R16742 gnd.n5971 gnd.n690 9.3005
R16743 gnd.n5972 gnd.n689 9.3005
R16744 gnd.n5973 gnd.n688 9.3005
R16745 gnd.n687 gnd.n683 9.3005
R16746 gnd.n5979 gnd.n682 9.3005
R16747 gnd.n5980 gnd.n681 9.3005
R16748 gnd.n5981 gnd.n680 9.3005
R16749 gnd.n679 gnd.n675 9.3005
R16750 gnd.n5987 gnd.n674 9.3005
R16751 gnd.n5988 gnd.n673 9.3005
R16752 gnd.n5989 gnd.n672 9.3005
R16753 gnd.n671 gnd.n667 9.3005
R16754 gnd.n5995 gnd.n666 9.3005
R16755 gnd.n5996 gnd.n665 9.3005
R16756 gnd.n5997 gnd.n664 9.3005
R16757 gnd.n663 gnd.n659 9.3005
R16758 gnd.n6003 gnd.n658 9.3005
R16759 gnd.n6004 gnd.n657 9.3005
R16760 gnd.n6005 gnd.n656 9.3005
R16761 gnd.n655 gnd.n651 9.3005
R16762 gnd.n6011 gnd.n650 9.3005
R16763 gnd.n6012 gnd.n649 9.3005
R16764 gnd.n6013 gnd.n648 9.3005
R16765 gnd.n647 gnd.n643 9.3005
R16766 gnd.n6019 gnd.n642 9.3005
R16767 gnd.n6020 gnd.n641 9.3005
R16768 gnd.n6021 gnd.n640 9.3005
R16769 gnd.n639 gnd.n635 9.3005
R16770 gnd.n6027 gnd.n634 9.3005
R16771 gnd.n6028 gnd.n633 9.3005
R16772 gnd.n6029 gnd.n632 9.3005
R16773 gnd.n631 gnd.n627 9.3005
R16774 gnd.n6035 gnd.n626 9.3005
R16775 gnd.n6036 gnd.n625 9.3005
R16776 gnd.n6037 gnd.n624 9.3005
R16777 gnd.n623 gnd.n619 9.3005
R16778 gnd.n6043 gnd.n618 9.3005
R16779 gnd.n6044 gnd.n617 9.3005
R16780 gnd.n6045 gnd.n616 9.3005
R16781 gnd.n615 gnd.n611 9.3005
R16782 gnd.n6051 gnd.n610 9.3005
R16783 gnd.n6052 gnd.n609 9.3005
R16784 gnd.n6053 gnd.n608 9.3005
R16785 gnd.n607 gnd.n603 9.3005
R16786 gnd.n6059 gnd.n602 9.3005
R16787 gnd.n6060 gnd.n601 9.3005
R16788 gnd.n6061 gnd.n600 9.3005
R16789 gnd.n599 gnd.n595 9.3005
R16790 gnd.n2459 gnd.n763 9.3005
R16791 gnd.n3480 gnd.n3479 9.3005
R16792 gnd.n3460 gnd.n3458 9.3005
R16793 gnd.n3487 gnd.n3486 9.3005
R16794 gnd.n3454 gnd.n3453 9.3005
R16795 gnd.n3499 gnd.n3498 9.3005
R16796 gnd.n3451 gnd.n3449 9.3005
R16797 gnd.n3506 gnd.n3505 9.3005
R16798 gnd.n3445 gnd.n3444 9.3005
R16799 gnd.n3518 gnd.n3517 9.3005
R16800 gnd.n3442 gnd.n3440 9.3005
R16801 gnd.n3525 gnd.n3524 9.3005
R16802 gnd.n3436 gnd.n3435 9.3005
R16803 gnd.n3537 gnd.n3536 9.3005
R16804 gnd.n3433 gnd.n3431 9.3005
R16805 gnd.n3546 gnd.n3545 9.3005
R16806 gnd.n3544 gnd.n3425 9.3005
R16807 gnd.n3555 gnd.n3424 9.3005
R16808 gnd.n3558 gnd.n3557 9.3005
R16809 gnd.n3463 gnd.n3462 9.3005
R16810 gnd.n3548 gnd.n3547 9.3005
R16811 gnd.n3535 gnd.n3430 9.3005
R16812 gnd.n3534 gnd.n3533 9.3005
R16813 gnd.n3441 gnd.n3437 9.3005
R16814 gnd.n3527 gnd.n3526 9.3005
R16815 gnd.n3516 gnd.n3439 9.3005
R16816 gnd.n3515 gnd.n3514 9.3005
R16817 gnd.n3450 gnd.n3446 9.3005
R16818 gnd.n3508 gnd.n3507 9.3005
R16819 gnd.n3497 gnd.n3448 9.3005
R16820 gnd.n3496 gnd.n3495 9.3005
R16821 gnd.n3459 gnd.n3455 9.3005
R16822 gnd.n3489 gnd.n3488 9.3005
R16823 gnd.n3478 gnd.n3457 9.3005
R16824 gnd.n3477 gnd.n3476 9.3005
R16825 gnd.n3465 gnd.n3464 9.3005
R16826 gnd.n3432 gnd.n3428 9.3005
R16827 gnd.n3554 gnd.n3553 9.3005
R16828 gnd.n3422 gnd.n3421 9.3005
R16829 gnd.n3565 gnd.n3564 9.3005
R16830 gnd.n3566 gnd.n3420 9.3005
R16831 gnd.n3568 gnd.n3567 9.3005
R16832 gnd.n3418 gnd.n3417 9.3005
R16833 gnd.n3578 gnd.n3577 9.3005
R16834 gnd.n3579 gnd.n3416 9.3005
R16835 gnd.n3581 gnd.n3580 9.3005
R16836 gnd.n3414 gnd.n3413 9.3005
R16837 gnd.n3587 gnd.n3586 9.3005
R16838 gnd.n2637 gnd.n2053 9.3005
R16839 gnd.n2636 gnd.n2635 9.3005
R16840 gnd.n2634 gnd.n2057 9.3005
R16841 gnd.n2633 gnd.n2632 9.3005
R16842 gnd.n2631 gnd.n2058 9.3005
R16843 gnd.n2630 gnd.n2629 9.3005
R16844 gnd.n2628 gnd.n2627 9.3005
R16845 gnd.n1787 gnd.n1786 9.3005
R16846 gnd.n2783 gnd.n2782 9.3005
R16847 gnd.n2784 gnd.n1784 9.3005
R16848 gnd.n2787 gnd.n2786 9.3005
R16849 gnd.n2785 gnd.n1785 9.3005
R16850 gnd.n1766 gnd.n1765 9.3005
R16851 gnd.n2814 gnd.n2813 9.3005
R16852 gnd.n2815 gnd.n1763 9.3005
R16853 gnd.n2824 gnd.n2823 9.3005
R16854 gnd.n2822 gnd.n1764 9.3005
R16855 gnd.n2821 gnd.n2820 9.3005
R16856 gnd.n2819 gnd.n2816 9.3005
R16857 gnd.n1718 gnd.n1717 9.3005
R16858 gnd.n2899 gnd.n2898 9.3005
R16859 gnd.n2900 gnd.n1715 9.3005
R16860 gnd.n2922 gnd.n2921 9.3005
R16861 gnd.n2920 gnd.n1716 9.3005
R16862 gnd.n2919 gnd.n2918 9.3005
R16863 gnd.n2917 gnd.n2901 9.3005
R16864 gnd.n2916 gnd.n2915 9.3005
R16865 gnd.n2914 gnd.n2908 9.3005
R16866 gnd.n2913 gnd.n2912 9.3005
R16867 gnd.n2911 gnd.n2910 9.3005
R16868 gnd.n2909 gnd.n1668 9.3005
R16869 gnd.n1666 gnd.n1665 9.3005
R16870 gnd.n3001 gnd.n3000 9.3005
R16871 gnd.n3002 gnd.n1664 9.3005
R16872 gnd.n3004 gnd.n3003 9.3005
R16873 gnd.n1641 gnd.n1639 9.3005
R16874 gnd.n3052 gnd.n3051 9.3005
R16875 gnd.n3050 gnd.n1640 9.3005
R16876 gnd.n3049 gnd.n3048 9.3005
R16877 gnd.n1618 gnd.n1616 9.3005
R16878 gnd.n3110 gnd.n3109 9.3005
R16879 gnd.n3108 gnd.n1617 9.3005
R16880 gnd.n3107 gnd.n3106 9.3005
R16881 gnd.n3105 gnd.n1619 9.3005
R16882 gnd.n3104 gnd.n3103 9.3005
R16883 gnd.n3102 gnd.n3091 9.3005
R16884 gnd.n3101 gnd.n3100 9.3005
R16885 gnd.n3099 gnd.n3092 9.3005
R16886 gnd.n3098 gnd.n3097 9.3005
R16887 gnd.n1558 gnd.n1557 9.3005
R16888 gnd.n3219 gnd.n3218 9.3005
R16889 gnd.n3220 gnd.n1555 9.3005
R16890 gnd.n3223 gnd.n3222 9.3005
R16891 gnd.n3221 gnd.n1556 9.3005
R16892 gnd.n1529 gnd.n1528 9.3005
R16893 gnd.n3258 gnd.n3257 9.3005
R16894 gnd.n3259 gnd.n1526 9.3005
R16895 gnd.n3276 gnd.n3275 9.3005
R16896 gnd.n3274 gnd.n1527 9.3005
R16897 gnd.n3273 gnd.n3272 9.3005
R16898 gnd.n3271 gnd.n3260 9.3005
R16899 gnd.n3270 gnd.n3269 9.3005
R16900 gnd.n3268 gnd.n3265 9.3005
R16901 gnd.n3267 gnd.n3266 9.3005
R16902 gnd.n1474 gnd.n1473 9.3005
R16903 gnd.n3351 gnd.n3350 9.3005
R16904 gnd.n3352 gnd.n1471 9.3005
R16905 gnd.n3355 gnd.n3354 9.3005
R16906 gnd.n3353 gnd.n1472 9.3005
R16907 gnd.n1447 gnd.n1446 9.3005
R16908 gnd.n3393 gnd.n3392 9.3005
R16909 gnd.n3394 gnd.n1445 9.3005
R16910 gnd.n3396 gnd.n3395 9.3005
R16911 gnd.n1444 gnd.n1443 9.3005
R16912 gnd.n3403 gnd.n3402 9.3005
R16913 gnd.n3404 gnd.n1442 9.3005
R16914 gnd.n3406 gnd.n3405 9.3005
R16915 gnd.n3407 gnd.n1441 9.3005
R16916 gnd.n3411 gnd.n3410 9.3005
R16917 gnd.n3412 gnd.n1439 9.3005
R16918 gnd.n3590 gnd.n3589 9.3005
R16919 gnd.n3588 gnd.n1440 9.3005
R16920 gnd.n2639 gnd.n2638 9.3005
R16921 gnd.n2642 gnd.n2641 9.3005
R16922 gnd.n2643 gnd.n2048 9.3005
R16923 gnd.n2645 gnd.n2644 9.3005
R16924 gnd.n2647 gnd.n2646 9.3005
R16925 gnd.n2648 gnd.n2041 9.3005
R16926 gnd.n2650 gnd.n2649 9.3005
R16927 gnd.n2651 gnd.n2040 9.3005
R16928 gnd.n2653 gnd.n2652 9.3005
R16929 gnd.n2654 gnd.n2034 9.3005
R16930 gnd.n2640 gnd.n2052 9.3005
R16931 gnd.n2251 gnd.n2249 9.3005
R16932 gnd.n2451 gnd.n2450 9.3005
R16933 gnd.n2449 gnd.n2250 9.3005
R16934 gnd.n2448 gnd.n2447 9.3005
R16935 gnd.n2241 gnd.n2240 9.3005
R16936 gnd.n2505 gnd.n2504 9.3005
R16937 gnd.n2506 gnd.n2239 9.3005
R16938 gnd.n2508 gnd.n2507 9.3005
R16939 gnd.n2234 gnd.n2233 9.3005
R16940 gnd.n2521 gnd.n2520 9.3005
R16941 gnd.n2522 gnd.n2232 9.3005
R16942 gnd.n2524 gnd.n2523 9.3005
R16943 gnd.n2224 gnd.n2222 9.3005
R16944 gnd.n2552 gnd.n2551 9.3005
R16945 gnd.n2550 gnd.n2223 9.3005
R16946 gnd.n2549 gnd.n2548 9.3005
R16947 gnd.n2547 gnd.n2225 9.3005
R16948 gnd.n2546 gnd.n2545 9.3005
R16949 gnd.n2033 gnd.n2031 9.3005
R16950 gnd.n2660 gnd.n2659 9.3005
R16951 gnd.n2658 gnd.n2032 9.3005
R16952 gnd.n2656 gnd.n2655 9.3005
R16953 gnd.n2036 gnd.n2035 9.3005
R16954 gnd.n2162 gnd.n2161 9.3005
R16955 gnd.n2164 gnd.n2163 9.3005
R16956 gnd.n2142 gnd.n2141 9.3005
R16957 gnd.n2170 gnd.n2169 9.3005
R16958 gnd.n2172 gnd.n2171 9.3005
R16959 gnd.n2132 gnd.n2131 9.3005
R16960 gnd.n2178 gnd.n2177 9.3005
R16961 gnd.n2180 gnd.n2179 9.3005
R16962 gnd.n2119 gnd.n2118 9.3005
R16963 gnd.n2186 gnd.n2185 9.3005
R16964 gnd.n2188 gnd.n2187 9.3005
R16965 gnd.n2109 gnd.n2108 9.3005
R16966 gnd.n2194 gnd.n2193 9.3005
R16967 gnd.n2196 gnd.n2195 9.3005
R16968 gnd.n2094 gnd.n2092 9.3005
R16969 gnd.n2202 gnd.n2201 9.3005
R16970 gnd.n2203 gnd.n2091 9.3005
R16971 gnd.n2096 gnd.n1086 9.3005
R16972 gnd.n2095 gnd.n2093 9.3005
R16973 gnd.n2200 gnd.n2199 9.3005
R16974 gnd.n2198 gnd.n2197 9.3005
R16975 gnd.n2104 gnd.n2103 9.3005
R16976 gnd.n2192 gnd.n2191 9.3005
R16977 gnd.n2190 gnd.n2189 9.3005
R16978 gnd.n2115 gnd.n2114 9.3005
R16979 gnd.n2184 gnd.n2183 9.3005
R16980 gnd.n2182 gnd.n2181 9.3005
R16981 gnd.n2126 gnd.n2125 9.3005
R16982 gnd.n2176 gnd.n2175 9.3005
R16983 gnd.n2174 gnd.n2173 9.3005
R16984 gnd.n2138 gnd.n2137 9.3005
R16985 gnd.n2168 gnd.n2167 9.3005
R16986 gnd.n2166 gnd.n2165 9.3005
R16987 gnd.n2151 gnd.n2150 9.3005
R16988 gnd.n2160 gnd.n2159 9.3005
R16989 gnd.n4269 gnd.n1087 9.3005
R16990 gnd.n4268 gnd.n4267 9.3005
R16991 gnd.n4266 gnd.n1091 9.3005
R16992 gnd.n4265 gnd.n4264 9.3005
R16993 gnd.n4263 gnd.n1092 9.3005
R16994 gnd.n4262 gnd.n4261 9.3005
R16995 gnd.n4260 gnd.n1096 9.3005
R16996 gnd.n4259 gnd.n4258 9.3005
R16997 gnd.n4257 gnd.n1097 9.3005
R16998 gnd.n4256 gnd.n4255 9.3005
R16999 gnd.n4254 gnd.n1101 9.3005
R17000 gnd.n4253 gnd.n4252 9.3005
R17001 gnd.n4251 gnd.n1102 9.3005
R17002 gnd.n4250 gnd.n4249 9.3005
R17003 gnd.n4248 gnd.n1106 9.3005
R17004 gnd.n4247 gnd.n4246 9.3005
R17005 gnd.n4245 gnd.n1107 9.3005
R17006 gnd.n4244 gnd.n4243 9.3005
R17007 gnd.n4242 gnd.n1111 9.3005
R17008 gnd.n4241 gnd.n4240 9.3005
R17009 gnd.n4239 gnd.n1112 9.3005
R17010 gnd.n4238 gnd.n4237 9.3005
R17011 gnd.n4236 gnd.n1116 9.3005
R17012 gnd.n4235 gnd.n4234 9.3005
R17013 gnd.n4233 gnd.n1117 9.3005
R17014 gnd.n4232 gnd.n4231 9.3005
R17015 gnd.n4230 gnd.n1121 9.3005
R17016 gnd.n4229 gnd.n4228 9.3005
R17017 gnd.n4227 gnd.n1122 9.3005
R17018 gnd.n4226 gnd.n4225 9.3005
R17019 gnd.n4224 gnd.n1126 9.3005
R17020 gnd.n4223 gnd.n4222 9.3005
R17021 gnd.n4221 gnd.n1127 9.3005
R17022 gnd.n4220 gnd.n4219 9.3005
R17023 gnd.n4218 gnd.n1131 9.3005
R17024 gnd.n4217 gnd.n4216 9.3005
R17025 gnd.n4215 gnd.n1132 9.3005
R17026 gnd.n4214 gnd.n4213 9.3005
R17027 gnd.n4212 gnd.n1136 9.3005
R17028 gnd.n4211 gnd.n4210 9.3005
R17029 gnd.n4209 gnd.n1137 9.3005
R17030 gnd.n4208 gnd.n4207 9.3005
R17031 gnd.n4206 gnd.n1141 9.3005
R17032 gnd.n4205 gnd.n4204 9.3005
R17033 gnd.n4203 gnd.n1142 9.3005
R17034 gnd.n4202 gnd.n4201 9.3005
R17035 gnd.n4200 gnd.n1146 9.3005
R17036 gnd.n4199 gnd.n4198 9.3005
R17037 gnd.n4197 gnd.n1147 9.3005
R17038 gnd.n4196 gnd.n4195 9.3005
R17039 gnd.n4194 gnd.n1151 9.3005
R17040 gnd.n4193 gnd.n4192 9.3005
R17041 gnd.n4191 gnd.n1152 9.3005
R17042 gnd.n4190 gnd.n4189 9.3005
R17043 gnd.n4188 gnd.n1156 9.3005
R17044 gnd.n4187 gnd.n4186 9.3005
R17045 gnd.n4185 gnd.n1157 9.3005
R17046 gnd.n4184 gnd.n4183 9.3005
R17047 gnd.n4182 gnd.n1161 9.3005
R17048 gnd.n4181 gnd.n4180 9.3005
R17049 gnd.n4179 gnd.n1162 9.3005
R17050 gnd.n4178 gnd.n4177 9.3005
R17051 gnd.n4176 gnd.n1166 9.3005
R17052 gnd.n4175 gnd.n4174 9.3005
R17053 gnd.n4173 gnd.n1167 9.3005
R17054 gnd.n4172 gnd.n4171 9.3005
R17055 gnd.n4170 gnd.n1171 9.3005
R17056 gnd.n4169 gnd.n4168 9.3005
R17057 gnd.n4167 gnd.n1172 9.3005
R17058 gnd.n4166 gnd.n4165 9.3005
R17059 gnd.n4164 gnd.n1176 9.3005
R17060 gnd.n4163 gnd.n4162 9.3005
R17061 gnd.n4161 gnd.n1177 9.3005
R17062 gnd.n4160 gnd.n4159 9.3005
R17063 gnd.n4158 gnd.n1181 9.3005
R17064 gnd.n4157 gnd.n4156 9.3005
R17065 gnd.n4155 gnd.n1182 9.3005
R17066 gnd.n4154 gnd.n4153 9.3005
R17067 gnd.n4152 gnd.n1186 9.3005
R17068 gnd.n4151 gnd.n4150 9.3005
R17069 gnd.n4149 gnd.n1187 9.3005
R17070 gnd.n4148 gnd.n1190 9.3005
R17071 gnd.n4271 gnd.n4270 9.3005
R17072 gnd.n1232 gnd.n1230 9.3005
R17073 gnd.n4122 gnd.n4121 9.3005
R17074 gnd.n4120 gnd.n1231 9.3005
R17075 gnd.n4119 gnd.n4118 9.3005
R17076 gnd.n4117 gnd.n1233 9.3005
R17077 gnd.n4116 gnd.n4115 9.3005
R17078 gnd.n4114 gnd.n1237 9.3005
R17079 gnd.n4113 gnd.n4112 9.3005
R17080 gnd.n4111 gnd.n1238 9.3005
R17081 gnd.n4110 gnd.n4109 9.3005
R17082 gnd.n4108 gnd.n1242 9.3005
R17083 gnd.n4107 gnd.n4106 9.3005
R17084 gnd.n4105 gnd.n1243 9.3005
R17085 gnd.n4104 gnd.n4103 9.3005
R17086 gnd.n4102 gnd.n1247 9.3005
R17087 gnd.n4101 gnd.n4100 9.3005
R17088 gnd.n4099 gnd.n1248 9.3005
R17089 gnd.n4098 gnd.n4097 9.3005
R17090 gnd.n242 gnd.n241 9.3005
R17091 gnd.n6652 gnd.n6651 9.3005
R17092 gnd.n6653 gnd.n239 9.3005
R17093 gnd.n6655 gnd.n6654 9.3005
R17094 gnd.n228 gnd.n227 9.3005
R17095 gnd.n6666 gnd.n6665 9.3005
R17096 gnd.n6667 gnd.n226 9.3005
R17097 gnd.n6669 gnd.n6668 9.3005
R17098 gnd.n207 gnd.n206 9.3005
R17099 gnd.n6682 gnd.n6681 9.3005
R17100 gnd.n6683 gnd.n205 9.3005
R17101 gnd.n6685 gnd.n6684 9.3005
R17102 gnd.n192 gnd.n191 9.3005
R17103 gnd.n6698 gnd.n6697 9.3005
R17104 gnd.n6699 gnd.n190 9.3005
R17105 gnd.n6701 gnd.n6700 9.3005
R17106 gnd.n177 gnd.n176 9.3005
R17107 gnd.n6714 gnd.n6713 9.3005
R17108 gnd.n6715 gnd.n174 9.3005
R17109 gnd.n6791 gnd.n6790 9.3005
R17110 gnd.n6789 gnd.n175 9.3005
R17111 gnd.n6788 gnd.n6787 9.3005
R17112 gnd.n6786 gnd.n6716 9.3005
R17113 gnd.n6785 gnd.n6784 9.3005
R17114 gnd.n3468 gnd.n3467 9.3005
R17115 gnd.n6781 gnd.n6718 9.3005
R17116 gnd.n6780 gnd.n6779 9.3005
R17117 gnd.n6778 gnd.n6723 9.3005
R17118 gnd.n6777 gnd.n6776 9.3005
R17119 gnd.n6775 gnd.n6724 9.3005
R17120 gnd.n6774 gnd.n6773 9.3005
R17121 gnd.n6772 gnd.n6731 9.3005
R17122 gnd.n6771 gnd.n6770 9.3005
R17123 gnd.n6769 gnd.n6732 9.3005
R17124 gnd.n6768 gnd.n6767 9.3005
R17125 gnd.n6766 gnd.n6739 9.3005
R17126 gnd.n6765 gnd.n6764 9.3005
R17127 gnd.n6763 gnd.n6740 9.3005
R17128 gnd.n6762 gnd.n6761 9.3005
R17129 gnd.n6760 gnd.n6747 9.3005
R17130 gnd.n6759 gnd.n6758 9.3005
R17131 gnd.n6757 gnd.n6748 9.3005
R17132 gnd.n6756 gnd.n78 9.3005
R17133 gnd.n6783 gnd.n6782 9.3005
R17134 gnd.n3893 gnd.n3892 9.3005
R17135 gnd.n3894 gnd.n1331 9.3005
R17136 gnd.n3897 gnd.n3896 9.3005
R17137 gnd.n3895 gnd.n1332 9.3005
R17138 gnd.n1316 gnd.n1315 9.3005
R17139 gnd.n4023 gnd.n4022 9.3005
R17140 gnd.n4024 gnd.n1313 9.3005
R17141 gnd.n4027 gnd.n4026 9.3005
R17142 gnd.n4025 gnd.n1314 9.3005
R17143 gnd.n1287 gnd.n1286 9.3005
R17144 gnd.n4055 gnd.n4054 9.3005
R17145 gnd.n4056 gnd.n1284 9.3005
R17146 gnd.n4059 gnd.n4058 9.3005
R17147 gnd.n4057 gnd.n1285 9.3005
R17148 gnd.n1258 gnd.n1257 9.3005
R17149 gnd.n4089 gnd.n4088 9.3005
R17150 gnd.n4090 gnd.n1254 9.3005
R17151 gnd.n4093 gnd.n4092 9.3005
R17152 gnd.n4091 gnd.n1256 9.3005
R17153 gnd.n1255 gnd.n51 9.3005
R17154 gnd.n6915 gnd.n52 9.3005
R17155 gnd.n6914 gnd.n6913 9.3005
R17156 gnd.n6912 gnd.n53 9.3005
R17157 gnd.n6911 gnd.n6910 9.3005
R17158 gnd.n6909 gnd.n57 9.3005
R17159 gnd.n6908 gnd.n6907 9.3005
R17160 gnd.n6906 gnd.n58 9.3005
R17161 gnd.n6905 gnd.n6904 9.3005
R17162 gnd.n6903 gnd.n62 9.3005
R17163 gnd.n6902 gnd.n6901 9.3005
R17164 gnd.n6900 gnd.n63 9.3005
R17165 gnd.n6899 gnd.n6898 9.3005
R17166 gnd.n6897 gnd.n67 9.3005
R17167 gnd.n6896 gnd.n6895 9.3005
R17168 gnd.n6894 gnd.n68 9.3005
R17169 gnd.n6893 gnd.n6892 9.3005
R17170 gnd.n6891 gnd.n72 9.3005
R17171 gnd.n6890 gnd.n6889 9.3005
R17172 gnd.n6888 gnd.n73 9.3005
R17173 gnd.n6887 gnd.n6886 9.3005
R17174 gnd.n6885 gnd.n77 9.3005
R17175 gnd.n6884 gnd.n6883 9.3005
R17176 gnd.n1334 gnd.n1333 9.3005
R17177 gnd.n5368 gnd.t86 9.24152
R17178 gnd.n5882 gnd.t148 9.24152
R17179 gnd.t141 gnd.n791 9.24152
R17180 gnd.n2555 gnd.t60 9.24152
R17181 gnd.t79 gnd.n1320 9.24152
R17182 gnd.t12 gnd.t86 8.92286
R17183 gnd.n2800 gnd.t195 8.92286
R17184 gnd.n1776 gnd.n1768 8.92286
R17185 gnd.t85 gnd.n2828 8.92286
R17186 gnd.n2987 gnd.n1675 8.92286
R17187 gnd.n3033 gnd.n1645 8.92286
R17188 gnd.n3158 gnd.n1579 8.92286
R17189 gnd.n3228 gnd.n3227 8.92286
R17190 gnd.n1485 gnd.t15 8.92286
R17191 gnd.n3371 gnd.n3370 8.92286
R17192 gnd.n3704 gnd.t181 8.92286
R17193 gnd.n5718 gnd.n5693 8.92171
R17194 gnd.n5686 gnd.n5661 8.92171
R17195 gnd.n5654 gnd.n5629 8.92171
R17196 gnd.n5623 gnd.n5598 8.92171
R17197 gnd.n5591 gnd.n5566 8.92171
R17198 gnd.n5559 gnd.n5534 8.92171
R17199 gnd.n5527 gnd.n5502 8.92171
R17200 gnd.n5496 gnd.n5471 8.92171
R17201 gnd.n3636 gnd.n3618 8.72777
R17202 gnd.t88 gnd.n4686 8.60421
R17203 gnd.n5086 gnd.n5074 8.43467
R17204 gnd.n38 gnd.n26 8.43467
R17205 gnd.n2428 gnd.n0 8.41456
R17206 gnd.n6916 gnd.n6915 8.41456
R17207 gnd.n2963 gnd.n1690 8.28555
R17208 gnd.n3054 gnd.n1628 8.28555
R17209 gnd.n3137 gnd.n1593 8.28555
R17210 gnd.n3193 gnd.n1546 8.28555
R17211 gnd.n5719 gnd.n5691 8.14595
R17212 gnd.n5687 gnd.n5659 8.14595
R17213 gnd.n5655 gnd.n5627 8.14595
R17214 gnd.n5624 gnd.n5596 8.14595
R17215 gnd.n5592 gnd.n5564 8.14595
R17216 gnd.n5560 gnd.n5532 8.14595
R17217 gnd.n5528 gnd.n5500 8.14595
R17218 gnd.n5497 gnd.n5469 8.14595
R17219 gnd.n5724 gnd.n5723 7.97301
R17220 gnd.t94 gnd.n4728 7.9669
R17221 gnd.n162 gnd.t119 7.9669
R17222 gnd.n6757 gnd.n6756 7.75808
R17223 gnd.n3553 gnd.n3428 7.75808
R17224 gnd.n2159 gnd.n2150 7.75808
R17225 gnd.n2298 gnd.n2294 7.75808
R17226 gnd.n2791 gnd.n1781 7.64824
R17227 gnd.n2963 gnd.n1689 7.64824
R17228 gnd.t50 gnd.n3007 7.64824
R17229 gnd.n3055 gnd.t245 7.64824
R17230 gnd.n3065 gnd.n1628 7.64824
R17231 gnd.n3137 gnd.n1592 7.64824
R17232 gnd.t270 gnd.n1587 7.64824
R17233 gnd.n3157 gnd.t30 7.64824
R17234 gnd.n3193 gnd.n1537 7.64824
R17235 gnd.n5198 gnd.t100 7.32958
R17236 gnd.n2791 gnd.t278 7.32958
R17237 gnd.t56 gnd.n3388 7.32958
R17238 gnd.n1811 gnd.n1810 7.30353
R17239 gnd.n3635 gnd.n3634 7.30353
R17240 gnd.n5158 gnd.n4803 7.01093
R17241 gnd.n4806 gnd.n4804 7.01093
R17242 gnd.n5168 gnd.n5167 7.01093
R17243 gnd.n5179 gnd.n4787 7.01093
R17244 gnd.n5178 gnd.n4790 7.01093
R17245 gnd.n5189 gnd.n4778 7.01093
R17246 gnd.n4781 gnd.n4779 7.01093
R17247 gnd.n5199 gnd.n5198 7.01093
R17248 gnd.n5210 gnd.n4761 7.01093
R17249 gnd.n5209 gnd.n4764 7.01093
R17250 gnd.n5220 gnd.n4754 7.01093
R17251 gnd.n5112 gnd.n4747 7.01093
R17252 gnd.n5241 gnd.n4736 7.01093
R17253 gnd.n5240 gnd.n4739 7.01093
R17254 gnd.n5251 gnd.n4728 7.01093
R17255 gnd.n4729 gnd.n4721 7.01093
R17256 gnd.n5272 gnd.n4710 7.01093
R17257 gnd.n5271 gnd.n4713 7.01093
R17258 gnd.n4703 gnd.n4696 7.01093
R17259 gnd.n5292 gnd.n5291 7.01093
R17260 gnd.n5302 gnd.n4686 7.01093
R17261 gnd.n5301 gnd.n4689 7.01093
R17262 gnd.n5312 gnd.n4679 7.01093
R17263 gnd.n5322 gnd.n4672 7.01093
R17264 gnd.n5346 gnd.n4666 7.01093
R17265 gnd.n5355 gnd.n4657 7.01093
R17266 gnd.n5364 gnd.n4649 7.01093
R17267 gnd.n5368 gnd.n5367 7.01093
R17268 gnd.n5386 gnd.n4634 7.01093
R17269 gnd.n5385 gnd.n4637 7.01093
R17270 gnd.n5396 gnd.n4626 7.01093
R17271 gnd.n4627 gnd.n4616 7.01093
R17272 gnd.n5431 gnd.n5430 7.01093
R17273 gnd.n5443 gnd.n5442 7.01093
R17274 gnd.n4603 gnd.n4595 7.01093
R17275 gnd.n5454 gnd.n5453 7.01093
R17276 gnd.n5753 gnd.n4580 7.01093
R17277 gnd.n5752 gnd.n4583 7.01093
R17278 gnd.n5768 gnd.n765 7.01093
R17279 gnd.n5896 gnd.n765 7.01093
R17280 gnd.n5895 gnd.n767 7.01093
R17281 gnd.n5774 gnd.n776 7.01093
R17282 gnd.n5889 gnd.n5888 7.01093
R17283 gnd.n5737 gnd.n779 7.01093
R17284 gnd.n5882 gnd.n788 7.01093
R17285 gnd.n5881 gnd.n791 7.01093
R17286 gnd.n5785 gnd.n799 7.01093
R17287 gnd.n5875 gnd.n5874 7.01093
R17288 gnd.n2810 gnd.n1768 7.01093
R17289 gnd.n2869 gnd.n1736 7.01093
R17290 gnd.t269 gnd.n2868 7.01093
R17291 gnd.n2987 gnd.n2986 7.01093
R17292 gnd.n3008 gnd.t50 7.01093
R17293 gnd.n3007 gnd.n1645 7.01093
R17294 gnd.n3158 gnd.n3157 7.01093
R17295 gnd.t30 gnd.n3155 7.01093
R17296 gnd.n3228 gnd.n1550 7.01093
R17297 gnd.n3311 gnd.t240 7.01093
R17298 gnd.n3328 gnd.n3327 7.01093
R17299 gnd.n3372 gnd.n3371 7.01093
R17300 gnd.n6801 gnd.n162 7.01093
R17301 gnd.n4764 gnd.t99 6.69227
R17302 gnd.n5364 gnd.t12 6.69227
R17303 gnd.n5767 gnd.t93 6.69227
R17304 gnd.t262 gnd.n1731 6.69227
R17305 gnd.n3263 gnd.t77 6.69227
R17306 gnd.n3765 gnd.n3764 6.5566
R17307 gnd.n1928 gnd.n1927 6.5566
R17308 gnd.n2716 gnd.n1853 6.5566
R17309 gnd.n3643 gnd.n3642 6.5566
R17310 gnd.n2617 gnd.n1789 6.37362
R17311 gnd.t195 gnd.t184 6.37362
R17312 gnd.n2931 gnd.n1704 6.37362
R17313 gnd.n3015 gnd.t16 6.37362
R17314 gnd.n3073 gnd.n1622 6.37362
R17315 gnd.n3085 gnd.n1609 6.37362
R17316 gnd.n3206 gnd.t27 6.37362
R17317 gnd.n3254 gnd.n1533 6.37362
R17318 gnd.n3370 gnd.t116 6.37362
R17319 gnd.n3380 gnd.t116 6.37362
R17320 gnd.n3704 gnd.n1402 6.37362
R17321 gnd.n2644 gnd.n2047 6.20656
R17322 gnd.n6846 gnd.n6843 6.20656
R17323 gnd.n4446 gnd.n4445 6.20656
R17324 gnd.n3576 gnd.n3416 6.20656
R17325 gnd.t256 gnd.n5260 6.05496
R17326 gnd.n5261 gnd.t97 6.05496
R17327 gnd.t252 gnd.n5301 6.05496
R17328 gnd.n5400 gnd.t96 6.05496
R17329 gnd.t234 gnd.t46 6.05496
R17330 gnd.t271 gnd.t227 6.05496
R17331 gnd.n5721 gnd.n5691 5.81868
R17332 gnd.n5689 gnd.n5659 5.81868
R17333 gnd.n5657 gnd.n5627 5.81868
R17334 gnd.n5626 gnd.n5596 5.81868
R17335 gnd.n5594 gnd.n5564 5.81868
R17336 gnd.n5562 gnd.n5532 5.81868
R17337 gnd.n5530 gnd.n5500 5.81868
R17338 gnd.n5499 gnd.n5469 5.81868
R17339 gnd.n1760 gnd.n1758 5.73631
R17340 gnd.n2829 gnd.n2826 5.73631
R17341 gnd.n1670 gnd.n1658 5.73631
R17342 gnd.n2998 gnd.n1651 5.73631
R17343 gnd.t245 gnd.n3054 5.73631
R17344 gnd.n1593 gnd.t270 5.73631
R17345 gnd.n3095 gnd.n3094 5.73631
R17346 gnd.n3165 gnd.n1568 5.73631
R17347 gnd.n3348 gnd.n1476 5.73631
R17348 gnd.n1479 gnd.n1468 5.73631
R17349 gnd.n3774 gnd.n1361 5.62001
R17350 gnd.n2711 gnd.n1932 5.62001
R17351 gnd.n2712 gnd.n2711 5.62001
R17352 gnd.n3774 gnd.n1362 5.62001
R17353 gnd.n4943 gnd.n4938 5.4308
R17354 gnd.n4561 gnd.n4559 5.4308
R17355 gnd.n5312 gnd.t95 5.41765
R17356 gnd.n5356 gnd.t87 5.41765
R17357 gnd.n5432 gnd.t286 5.41765
R17358 gnd.t71 gnd.n2946 5.41765
R17359 gnd.n3185 gnd.t82 5.41765
R17360 gnd.t84 gnd.n2860 5.09899
R17361 gnd.n2939 gnd.n1708 5.09899
R17362 gnd.n3113 gnd.n1613 5.09899
R17363 gnd.n3121 gnd.n1606 5.09899
R17364 gnd.n3288 gnd.n1517 5.09899
R17365 gnd.n1509 gnd.t31 5.09899
R17366 gnd.n5719 gnd.n5718 5.04292
R17367 gnd.n5687 gnd.n5686 5.04292
R17368 gnd.n5655 gnd.n5654 5.04292
R17369 gnd.n5624 gnd.n5623 5.04292
R17370 gnd.n5592 gnd.n5591 5.04292
R17371 gnd.n5560 gnd.n5559 5.04292
R17372 gnd.n5528 gnd.n5527 5.04292
R17373 gnd.n5497 gnd.n5496 5.04292
R17374 gnd.n5098 gnd.n5097 4.82753
R17375 gnd.n50 gnd.n49 4.82753
R17376 gnd.n5282 gnd.t90 4.78034
R17377 gnd.n4637 gnd.t91 4.78034
R17378 gnd.t232 gnd.n2623 4.78034
R17379 gnd.n3771 gnd.t162 4.78034
R17380 gnd.n3605 gnd.t52 4.78034
R17381 gnd.n5102 gnd.n5101 4.74817
R17382 gnd.n5063 gnd.n5061 4.74817
R17383 gnd.n5056 gnd.n5055 4.74817
R17384 gnd.n5052 gnd.n5051 4.74817
R17385 gnd.n5101 gnd.n5050 4.74817
R17386 gnd.n5063 gnd.n5062 4.74817
R17387 gnd.n5057 gnd.n5056 4.74817
R17388 gnd.n5054 gnd.n5052 4.74817
R17389 gnd.n1265 gnd.n218 4.74817
R17390 gnd.n6646 gnd.n217 4.74817
R17391 gnd.n234 gnd.n216 4.74817
R17392 gnd.n6660 gnd.n215 4.74817
R17393 gnd.n219 gnd.n214 4.74817
R17394 gnd.n4084 gnd.n218 4.74817
R17395 gnd.n1264 gnd.n217 4.74817
R17396 gnd.n6647 gnd.n216 4.74817
R17397 gnd.n235 gnd.n215 4.74817
R17398 gnd.n6661 gnd.n214 4.74817
R17399 gnd.n4355 gnd.n4354 4.74817
R17400 gnd.n975 gnd.n955 4.74817
R17401 gnd.n4342 gnd.n4341 4.74817
R17402 gnd.n992 gnd.n976 4.74817
R17403 gnd.n4329 gnd.n4328 4.74817
R17404 gnd.n4356 gnd.n4355 4.74817
R17405 gnd.n4353 gnd.n955 4.74817
R17406 gnd.n4343 gnd.n4342 4.74817
R17407 gnd.n4340 gnd.n976 4.74817
R17408 gnd.n4330 gnd.n4329 4.74817
R17409 gnd.n5086 gnd.n5085 4.7074
R17410 gnd.n38 gnd.n37 4.7074
R17411 gnd.n5098 gnd.n5086 4.65959
R17412 gnd.n50 gnd.n38 4.65959
R17413 gnd.n3833 gnd.n3832 4.6132
R17414 gnd.n2707 gnd.n2706 4.6132
R17415 gnd.n2836 gnd.n1751 4.46168
R17416 gnd.n2827 gnd.n1740 4.46168
R17417 gnd.n2984 gnd.t235 4.46168
R17418 gnd.n2995 gnd.n2993 4.46168
R17419 gnd.n3024 gnd.n1653 4.46168
R17420 gnd.n3172 gnd.n1573 4.46168
R17421 gnd.n3216 gnd.n1560 4.46168
R17422 gnd.t17 gnd.n3214 4.46168
R17423 gnd.n3338 gnd.n1484 4.46168
R17424 gnd.n3358 gnd.n3357 4.46168
R17425 gnd.t207 gnd.n1407 4.46168
R17426 gnd.n3631 gnd.n3618 4.46111
R17427 gnd.n5704 gnd.n5700 4.38594
R17428 gnd.n5672 gnd.n5668 4.38594
R17429 gnd.n5640 gnd.n5636 4.38594
R17430 gnd.n5609 gnd.n5605 4.38594
R17431 gnd.n5577 gnd.n5573 4.38594
R17432 gnd.n5545 gnd.n5541 4.38594
R17433 gnd.n5513 gnd.n5509 4.38594
R17434 gnd.n5482 gnd.n5478 4.38594
R17435 gnd.n5715 gnd.n5693 4.26717
R17436 gnd.n5683 gnd.n5661 4.26717
R17437 gnd.n5651 gnd.n5629 4.26717
R17438 gnd.n5620 gnd.n5598 4.26717
R17439 gnd.n5588 gnd.n5566 4.26717
R17440 gnd.n5556 gnd.n5534 4.26717
R17441 gnd.n5524 gnd.n5502 4.26717
R17442 gnd.n5493 gnd.n5471 4.26717
R17443 gnd.n5230 gnd.t92 4.14303
R17444 gnd.n5453 gnd.t89 4.14303
R17445 gnd.t134 gnd.n1072 4.14303
R17446 gnd.t123 gnd.n1224 4.14303
R17447 gnd.n5723 gnd.n5722 4.08274
R17448 gnd.n3764 gnd.n3763 4.05904
R17449 gnd.n1927 gnd.n1926 4.05904
R17450 gnd.n2719 gnd.n1853 4.05904
R17451 gnd.n3644 gnd.n3643 4.05904
R17452 gnd.n15 gnd.n7 3.99943
R17453 gnd.n2779 gnd.n1791 3.82437
R17454 gnd.n2895 gnd.n1721 3.82437
R17455 gnd.n2937 gnd.t276 3.82437
R17456 gnd.n2956 gnd.n2955 3.82437
R17457 gnd.n3044 gnd.n1642 3.82437
R17458 gnd.n3046 gnd.t234 3.82437
R17459 gnd.n3087 gnd.t271 3.82437
R17460 gnd.n3130 gnd.n3129 3.82437
R17461 gnd.n3245 gnd.n1531 3.82437
R17462 gnd.n3279 gnd.t266 3.82437
R17463 gnd.n3297 gnd.n3296 3.82437
R17464 gnd.n3612 gnd.n1410 3.82437
R17465 gnd.n5723 gnd.n5595 3.70378
R17466 gnd.n5100 gnd.n5099 3.65935
R17467 gnd.n15 gnd.n14 3.60163
R17468 gnd.n5714 gnd.n5695 3.49141
R17469 gnd.n5682 gnd.n5663 3.49141
R17470 gnd.n5650 gnd.n5631 3.49141
R17471 gnd.n5619 gnd.n5600 3.49141
R17472 gnd.n5587 gnd.n5568 3.49141
R17473 gnd.n5555 gnd.n5536 3.49141
R17474 gnd.n5523 gnd.n5504 3.49141
R17475 gnd.n5492 gnd.n5473 3.49141
R17476 gnd.n2799 gnd.n2798 3.18706
R17477 gnd.n1760 gnd.t188 3.18706
R17478 gnd.n2867 gnd.n1729 3.18706
R17479 gnd.n2876 gnd.t6 3.18706
R17480 gnd.t6 gnd.n1713 3.18706
R17481 gnd.n2973 gnd.n2972 3.18706
R17482 gnd.n3035 gnd.n3034 3.18706
R17483 gnd.n3145 gnd.n3144 3.18706
R17484 gnd.n3226 gnd.n3225 3.18706
R17485 gnd.t236 gnd.n1520 3.18706
R17486 gnd.n3177 gnd.t236 3.18706
R17487 gnd.n3314 gnd.n3312 3.18706
R17488 gnd.n3380 gnd.n1453 3.18706
R17489 gnd.n3388 gnd.t207 3.18706
R17490 gnd.t92 gnd.n5229 2.8684
R17491 gnd.n2843 gnd.t290 2.8684
R17492 gnd.t229 gnd.n3347 2.8684
R17493 gnd.n5087 gnd.t43 2.82907
R17494 gnd.n5087 gnd.t267 2.82907
R17495 gnd.n5089 gnd.t238 2.82907
R17496 gnd.n5089 gnd.t34 2.82907
R17497 gnd.n5091 gnd.t272 2.82907
R17498 gnd.n5091 gnd.t284 2.82907
R17499 gnd.n5093 gnd.t1 2.82907
R17500 gnd.n5093 gnd.t264 2.82907
R17501 gnd.n5095 gnd.t8 2.82907
R17502 gnd.n5095 gnd.t36 2.82907
R17503 gnd.n5064 gnd.t277 2.82907
R17504 gnd.n5064 gnd.t241 2.82907
R17505 gnd.n5066 gnd.t223 2.82907
R17506 gnd.n5066 gnd.t21 2.82907
R17507 gnd.n5068 gnd.t265 2.82907
R17508 gnd.n5068 gnd.t3 2.82907
R17509 gnd.n5070 gnd.t33 2.82907
R17510 gnd.n5070 gnd.t74 2.82907
R17511 gnd.n5072 gnd.t275 2.82907
R17512 gnd.n5072 gnd.t289 2.82907
R17513 gnd.n5075 gnd.t258 2.82907
R17514 gnd.n5075 gnd.t69 2.82907
R17515 gnd.n5077 gnd.t282 2.82907
R17516 gnd.n5077 gnd.t81 2.82907
R17517 gnd.n5079 gnd.t26 2.82907
R17518 gnd.n5079 gnd.t9 2.82907
R17519 gnd.n5081 gnd.t22 2.82907
R17520 gnd.n5081 gnd.t247 2.82907
R17521 gnd.n5083 gnd.t288 2.82907
R17522 gnd.n5083 gnd.t248 2.82907
R17523 gnd.n47 gnd.t242 2.82907
R17524 gnd.n47 gnd.t49 2.82907
R17525 gnd.n45 gnd.t243 2.82907
R17526 gnd.n45 gnd.t19 2.82907
R17527 gnd.n43 gnd.t103 2.82907
R17528 gnd.n43 gnd.t273 2.82907
R17529 gnd.n41 gnd.t246 2.82907
R17530 gnd.n41 gnd.t58 2.82907
R17531 gnd.n39 gnd.t220 2.82907
R17532 gnd.n39 gnd.t59 2.82907
R17533 gnd.n24 gnd.t62 2.82907
R17534 gnd.n24 gnd.t70 2.82907
R17535 gnd.n22 gnd.t244 2.82907
R17536 gnd.n22 gnd.t274 2.82907
R17537 gnd.n20 gnd.t106 2.82907
R17538 gnd.n20 gnd.t65 2.82907
R17539 gnd.n18 gnd.t105 2.82907
R17540 gnd.n18 gnd.t41 2.82907
R17541 gnd.n16 gnd.t11 2.82907
R17542 gnd.n16 gnd.t39 2.82907
R17543 gnd.n35 gnd.t24 2.82907
R17544 gnd.n35 gnd.t281 2.82907
R17545 gnd.n33 gnd.t55 2.82907
R17546 gnd.n33 gnd.t231 2.82907
R17547 gnd.n31 gnd.t224 2.82907
R17548 gnd.n31 gnd.t285 2.82907
R17549 gnd.n29 gnd.t221 2.82907
R17550 gnd.n29 gnd.t226 2.82907
R17551 gnd.n27 gnd.t283 2.82907
R17552 gnd.n27 gnd.t225 2.82907
R17553 gnd.n5711 gnd.n5710 2.71565
R17554 gnd.n5679 gnd.n5678 2.71565
R17555 gnd.n5647 gnd.n5646 2.71565
R17556 gnd.n5616 gnd.n5615 2.71565
R17557 gnd.n5584 gnd.n5583 2.71565
R17558 gnd.n5552 gnd.n5551 2.71565
R17559 gnd.n5520 gnd.n5519 2.71565
R17560 gnd.n5489 gnd.n5488 2.71565
R17561 gnd.n2800 gnd.n1774 2.54975
R17562 gnd.n2885 gnd.n2884 2.54975
R17563 gnd.n2861 gnd.t84 2.54975
R17564 gnd.n2974 gnd.n1684 2.54975
R17565 gnd.n2974 gnd.t51 2.54975
R17566 gnd.n3055 gnd.n1635 2.54975
R17567 gnd.n3146 gnd.n1587 2.54975
R17568 gnd.n3235 gnd.t14 2.54975
R17569 gnd.n3235 gnd.n3234 2.54975
R17570 gnd.n3304 gnd.t31 2.54975
R17571 gnd.n3315 gnd.n1498 2.54975
R17572 gnd.n1462 gnd.n1449 2.54975
R17573 gnd.n5101 gnd.n5100 2.27742
R17574 gnd.n5100 gnd.n5063 2.27742
R17575 gnd.n5100 gnd.n5056 2.27742
R17576 gnd.n5100 gnd.n5052 2.27742
R17577 gnd.n6674 gnd.n218 2.27742
R17578 gnd.n6674 gnd.n217 2.27742
R17579 gnd.n6674 gnd.n216 2.27742
R17580 gnd.n6674 gnd.n215 2.27742
R17581 gnd.n6674 gnd.n214 2.27742
R17582 gnd.n4355 gnd.n953 2.27742
R17583 gnd.n955 gnd.n953 2.27742
R17584 gnd.n4342 gnd.n953 2.27742
R17585 gnd.n976 gnd.n953 2.27742
R17586 gnd.n4329 gnd.n953 2.27742
R17587 gnd.n5167 gnd.t112 2.23109
R17588 gnd.n5059 gnd.t90 2.23109
R17589 gnd.t260 gnd.n1653 2.23109
R17590 gnd.t46 gnd.n3044 2.23109
R17591 gnd.n3130 gnd.t227 2.23109
R17592 gnd.t44 gnd.n1573 2.23109
R17593 gnd.n5707 gnd.n5697 1.93989
R17594 gnd.n5675 gnd.n5665 1.93989
R17595 gnd.n5643 gnd.n5633 1.93989
R17596 gnd.n5612 gnd.n5602 1.93989
R17597 gnd.n5580 gnd.n5570 1.93989
R17598 gnd.n5548 gnd.n5538 1.93989
R17599 gnd.n5516 gnd.n5506 1.93989
R17600 gnd.n5485 gnd.n5475 1.93989
R17601 gnd.n1863 gnd.n1862 1.91244
R17602 gnd.n1863 gnd.t145 1.91244
R17603 gnd.n2869 gnd.t269 1.91244
R17604 gnd.n2896 gnd.n1720 1.91244
R17605 gnd.n2905 gnd.n2903 1.91244
R17606 gnd.n3064 gnd.n1630 1.91244
R17607 gnd.n1600 gnd.n1599 1.91244
R17608 gnd.n3248 gnd.n3247 1.91244
R17609 gnd.n1511 gnd.n1510 1.91244
R17610 gnd.n3328 gnd.t240 1.91244
R17611 gnd.n3614 gnd.n3613 1.91244
R17612 gnd.t4 gnd.n5178 1.59378
R17613 gnd.n5345 gnd.t87 1.59378
R17614 gnd.n5399 gnd.t286 1.59378
R17615 gnd.n2861 gnd.t262 1.59378
R17616 gnd.t109 gnd.n1675 1.59378
R17617 gnd.n3227 gnd.t254 1.59378
R17618 gnd.n3304 gnd.t77 1.59378
R17619 gnd.n2617 gnd.t201 1.27512
R17620 gnd.n2809 gnd.n2808 1.27512
R17621 gnd.n2829 gnd.t85 1.27512
R17622 gnd.n2852 gnd.n2851 1.27512
R17623 gnd.n2947 gnd.t276 1.27512
R17624 gnd.n2985 gnd.n2984 1.27512
R17625 gnd.n3008 gnd.n1662 1.27512
R17626 gnd.n3155 gnd.n3154 1.27512
R17627 gnd.n3214 gnd.n1561 1.27512
R17628 gnd.n3184 gnd.t266 1.27512
R17629 gnd.n3326 gnd.n3325 1.27512
R17630 gnd.t15 gnd.n1476 1.27512
R17631 gnd.n3357 gnd.t131 1.27512
R17632 gnd.n3373 gnd.n1458 1.27512
R17633 gnd.n4946 gnd.n4938 1.16414
R17634 gnd.n5800 gnd.n4559 1.16414
R17635 gnd.n5706 gnd.n5699 1.16414
R17636 gnd.n5674 gnd.n5667 1.16414
R17637 gnd.n5642 gnd.n5635 1.16414
R17638 gnd.n5611 gnd.n5604 1.16414
R17639 gnd.n5579 gnd.n5572 1.16414
R17640 gnd.n5547 gnd.n5540 1.16414
R17641 gnd.n5515 gnd.n5508 1.16414
R17642 gnd.n5484 gnd.n5477 1.16414
R17643 gnd.n3832 gnd.n1358 0.970197
R17644 gnd.n2707 gnd.n1933 0.970197
R17645 gnd.n5690 gnd.n5658 0.962709
R17646 gnd.n5722 gnd.n5690 0.962709
R17647 gnd.n5563 gnd.n5531 0.962709
R17648 gnd.n5595 gnd.n5563 0.962709
R17649 gnd.n5261 gnd.t256 0.956468
R17650 gnd.n5409 gnd.t96 0.956468
R17651 gnd.n4377 gnd.t7 0.956468
R17652 gnd.n2235 gnd.t42 0.956468
R17653 gnd.n2526 gnd.t68 0.956468
R17654 gnd.n2771 gnd.n1849 0.956468
R17655 gnd.t278 gnd.n2790 0.956468
R17656 gnd.n3390 gnd.t56 0.956468
R17657 gnd.n3771 gnd.n1365 0.956468
R17658 gnd.n4041 gnd.t10 0.956468
R17659 gnd.n1291 gnd.t38 0.956468
R17660 gnd.t48 gnd.n186 0.956468
R17661 gnd.n5094 gnd.n5092 0.773756
R17662 gnd.n46 gnd.n44 0.773756
R17663 gnd.n5097 gnd.n5096 0.773756
R17664 gnd.n5096 gnd.n5094 0.773756
R17665 gnd.n5092 gnd.n5090 0.773756
R17666 gnd.n5090 gnd.n5088 0.773756
R17667 gnd.n42 gnd.n40 0.773756
R17668 gnd.n44 gnd.n42 0.773756
R17669 gnd.n48 gnd.n46 0.773756
R17670 gnd.n49 gnd.n48 0.773756
R17671 gnd.n2 gnd.n1 0.672012
R17672 gnd.n3 gnd.n2 0.672012
R17673 gnd.n4 gnd.n3 0.672012
R17674 gnd.n5 gnd.n4 0.672012
R17675 gnd.n6 gnd.n5 0.672012
R17676 gnd.n7 gnd.n6 0.672012
R17677 gnd.n9 gnd.n8 0.672012
R17678 gnd.n10 gnd.n9 0.672012
R17679 gnd.n11 gnd.n10 0.672012
R17680 gnd.n12 gnd.n11 0.672012
R17681 gnd.n13 gnd.n12 0.672012
R17682 gnd.n14 gnd.n13 0.672012
R17683 gnd.t184 gnd.n2799 0.637812
R17684 gnd.t171 gnd.n2809 0.637812
R17685 gnd.n2926 gnd.n2925 0.637812
R17686 gnd.n2946 gnd.n2945 0.637812
R17687 gnd.n2955 gnd.t32 0.637812
R17688 gnd.n3075 gnd.n3074 0.637812
R17689 gnd.n3120 gnd.n3119 0.637812
R17690 gnd.t239 gnd.n3245 0.637812
R17691 gnd.n3186 gnd.n3185 0.637812
R17692 gnd.n3287 gnd.n3285 0.637812
R17693 gnd.t127 gnd.n1453 0.637812
R17694 gnd.n3397 gnd.t181 0.637812
R17695 gnd.n5074 gnd.n5073 0.573776
R17696 gnd.n5073 gnd.n5071 0.573776
R17697 gnd.n5071 gnd.n5069 0.573776
R17698 gnd.n5069 gnd.n5067 0.573776
R17699 gnd.n5067 gnd.n5065 0.573776
R17700 gnd.n5085 gnd.n5084 0.573776
R17701 gnd.n5084 gnd.n5082 0.573776
R17702 gnd.n5082 gnd.n5080 0.573776
R17703 gnd.n5080 gnd.n5078 0.573776
R17704 gnd.n5078 gnd.n5076 0.573776
R17705 gnd.n19 gnd.n17 0.573776
R17706 gnd.n21 gnd.n19 0.573776
R17707 gnd.n23 gnd.n21 0.573776
R17708 gnd.n25 gnd.n23 0.573776
R17709 gnd.n26 gnd.n25 0.573776
R17710 gnd.n30 gnd.n28 0.573776
R17711 gnd.n32 gnd.n30 0.573776
R17712 gnd.n34 gnd.n32 0.573776
R17713 gnd.n36 gnd.n34 0.573776
R17714 gnd.n37 gnd.n36 0.573776
R17715 gnd gnd.n0 0.551497
R17716 gnd.n6674 gnd.n213 0.5435
R17717 gnd.n2468 gnd.n953 0.5435
R17718 gnd.n2299 gnd.n2297 0.532512
R17719 gnd.n2337 gnd.n2336 0.532512
R17720 gnd.n6784 gnd.n6783 0.532512
R17721 gnd.n6884 gnd.n78 0.532512
R17722 gnd.n4272 gnd.n4271 0.523366
R17723 gnd.n3466 gnd.n1190 0.523366
R17724 gnd.n6878 gnd.n6877 0.520317
R17725 gnd.n6807 gnd.n6806 0.520317
R17726 gnd.n3886 gnd.n3885 0.520317
R17727 gnd.n3790 gnd.n1219 0.520317
R17728 gnd.n1954 gnd.n1077 0.520317
R17729 gnd.n2667 gnd.n2666 0.520317
R17730 gnd.n4406 gnd.n877 0.520317
R17731 gnd.n2346 gnd.n834 0.520317
R17732 gnd.n3588 gnd.n3587 0.489829
R17733 gnd.n2640 gnd.n2639 0.489829
R17734 gnd.n5790 gnd.n5789 0.486781
R17735 gnd.n4995 gnd.n4994 0.48678
R17736 gnd.n5871 gnd.n5870 0.480683
R17737 gnd.n5153 gnd.n5152 0.480683
R17738 gnd.n6917 gnd.n6916 0.470187
R17739 gnd.n6068 gnd.n595 0.438
R17740 gnd.n6421 gnd.n6420 0.438
R17741 gnd.n6633 gnd.n6632 0.438
R17742 gnd.n2460 gnd.n2459 0.438
R17743 gnd.n4274 gnd.n4273 0.432431
R17744 gnd.n3469 gnd.n3468 0.432431
R17745 gnd.n2647 gnd.n2047 0.388379
R17746 gnd.n5703 gnd.n5702 0.388379
R17747 gnd.n5671 gnd.n5670 0.388379
R17748 gnd.n5639 gnd.n5638 0.388379
R17749 gnd.n5608 gnd.n5607 0.388379
R17750 gnd.n5576 gnd.n5575 0.388379
R17751 gnd.n5544 gnd.n5543 0.388379
R17752 gnd.n5512 gnd.n5511 0.388379
R17753 gnd.n5481 gnd.n5480 0.388379
R17754 gnd.n6847 gnd.n6846 0.388379
R17755 gnd.n4447 gnd.n4446 0.388379
R17756 gnd.n3577 gnd.n3576 0.388379
R17757 gnd.n6917 gnd.n15 0.374463
R17758 gnd.n4585 gnd.t93 0.319156
R17759 gnd.n2420 gnd.t73 0.319156
R17760 gnd.n2454 gnd.t2 0.319156
R17761 gnd.n2445 gnd.t222 0.319156
R17762 gnd.n2588 gnd.t177 0.319156
R17763 gnd.t158 gnd.n3593 0.319156
R17764 gnd.n3972 gnd.t40 0.319156
R17765 gnd.n6643 gnd.t102 0.319156
R17766 gnd.t54 gnd.n222 0.319156
R17767 gnd.n4913 gnd.n4891 0.311721
R17768 gnd.n2658 gnd.n2657 0.302329
R17769 gnd.n3556 gnd.n1333 0.302329
R17770 gnd gnd.n6917 0.295112
R17771 gnd.n5840 gnd.n5839 0.268793
R17772 gnd.n5839 gnd.n5838 0.241354
R17773 gnd.n3833 gnd.n1359 0.229039
R17774 gnd.n3834 gnd.n3833 0.229039
R17775 gnd.n2706 gnd.n1938 0.229039
R17776 gnd.n2706 gnd.n2705 0.229039
R17777 gnd.n5141 gnd.n4866 0.206293
R17778 gnd.n5720 gnd.n5692 0.155672
R17779 gnd.n5713 gnd.n5692 0.155672
R17780 gnd.n5713 gnd.n5712 0.155672
R17781 gnd.n5712 gnd.n5696 0.155672
R17782 gnd.n5705 gnd.n5696 0.155672
R17783 gnd.n5705 gnd.n5704 0.155672
R17784 gnd.n5688 gnd.n5660 0.155672
R17785 gnd.n5681 gnd.n5660 0.155672
R17786 gnd.n5681 gnd.n5680 0.155672
R17787 gnd.n5680 gnd.n5664 0.155672
R17788 gnd.n5673 gnd.n5664 0.155672
R17789 gnd.n5673 gnd.n5672 0.155672
R17790 gnd.n5656 gnd.n5628 0.155672
R17791 gnd.n5649 gnd.n5628 0.155672
R17792 gnd.n5649 gnd.n5648 0.155672
R17793 gnd.n5648 gnd.n5632 0.155672
R17794 gnd.n5641 gnd.n5632 0.155672
R17795 gnd.n5641 gnd.n5640 0.155672
R17796 gnd.n5625 gnd.n5597 0.155672
R17797 gnd.n5618 gnd.n5597 0.155672
R17798 gnd.n5618 gnd.n5617 0.155672
R17799 gnd.n5617 gnd.n5601 0.155672
R17800 gnd.n5610 gnd.n5601 0.155672
R17801 gnd.n5610 gnd.n5609 0.155672
R17802 gnd.n5593 gnd.n5565 0.155672
R17803 gnd.n5586 gnd.n5565 0.155672
R17804 gnd.n5586 gnd.n5585 0.155672
R17805 gnd.n5585 gnd.n5569 0.155672
R17806 gnd.n5578 gnd.n5569 0.155672
R17807 gnd.n5578 gnd.n5577 0.155672
R17808 gnd.n5561 gnd.n5533 0.155672
R17809 gnd.n5554 gnd.n5533 0.155672
R17810 gnd.n5554 gnd.n5553 0.155672
R17811 gnd.n5553 gnd.n5537 0.155672
R17812 gnd.n5546 gnd.n5537 0.155672
R17813 gnd.n5546 gnd.n5545 0.155672
R17814 gnd.n5529 gnd.n5501 0.155672
R17815 gnd.n5522 gnd.n5501 0.155672
R17816 gnd.n5522 gnd.n5521 0.155672
R17817 gnd.n5521 gnd.n5505 0.155672
R17818 gnd.n5514 gnd.n5505 0.155672
R17819 gnd.n5514 gnd.n5513 0.155672
R17820 gnd.n5498 gnd.n5470 0.155672
R17821 gnd.n5491 gnd.n5470 0.155672
R17822 gnd.n5491 gnd.n5490 0.155672
R17823 gnd.n5490 gnd.n5474 0.155672
R17824 gnd.n5483 gnd.n5474 0.155672
R17825 gnd.n5483 gnd.n5482 0.155672
R17826 gnd.n5870 gnd.n4489 0.152939
R17827 gnd.n4491 gnd.n4489 0.152939
R17828 gnd.n4495 gnd.n4491 0.152939
R17829 gnd.n4496 gnd.n4495 0.152939
R17830 gnd.n4497 gnd.n4496 0.152939
R17831 gnd.n4498 gnd.n4497 0.152939
R17832 gnd.n4502 gnd.n4498 0.152939
R17833 gnd.n4503 gnd.n4502 0.152939
R17834 gnd.n4504 gnd.n4503 0.152939
R17835 gnd.n4505 gnd.n4504 0.152939
R17836 gnd.n4509 gnd.n4505 0.152939
R17837 gnd.n4510 gnd.n4509 0.152939
R17838 gnd.n4511 gnd.n4510 0.152939
R17839 gnd.n4512 gnd.n4511 0.152939
R17840 gnd.n4517 gnd.n4512 0.152939
R17841 gnd.n5840 gnd.n4517 0.152939
R17842 gnd.n5154 gnd.n5153 0.152939
R17843 gnd.n5154 gnd.n4784 0.152939
R17844 gnd.n5182 gnd.n4784 0.152939
R17845 gnd.n5183 gnd.n5182 0.152939
R17846 gnd.n5184 gnd.n5183 0.152939
R17847 gnd.n5185 gnd.n5184 0.152939
R17848 gnd.n5185 gnd.n4758 0.152939
R17849 gnd.n5213 gnd.n4758 0.152939
R17850 gnd.n5214 gnd.n5213 0.152939
R17851 gnd.n5215 gnd.n5214 0.152939
R17852 gnd.n5216 gnd.n5215 0.152939
R17853 gnd.n5216 gnd.n4733 0.152939
R17854 gnd.n5244 gnd.n4733 0.152939
R17855 gnd.n5245 gnd.n5244 0.152939
R17856 gnd.n5246 gnd.n5245 0.152939
R17857 gnd.n5247 gnd.n5246 0.152939
R17858 gnd.n5247 gnd.n4707 0.152939
R17859 gnd.n5275 gnd.n4707 0.152939
R17860 gnd.n5276 gnd.n5275 0.152939
R17861 gnd.n5277 gnd.n5276 0.152939
R17862 gnd.n5278 gnd.n5277 0.152939
R17863 gnd.n5278 gnd.n4683 0.152939
R17864 gnd.n5305 gnd.n4683 0.152939
R17865 gnd.n5306 gnd.n5305 0.152939
R17866 gnd.n5307 gnd.n5306 0.152939
R17867 gnd.n5308 gnd.n5307 0.152939
R17868 gnd.n5308 gnd.n4652 0.152939
R17869 gnd.n5359 gnd.n4652 0.152939
R17870 gnd.n5360 gnd.n5359 0.152939
R17871 gnd.n5361 gnd.n5360 0.152939
R17872 gnd.n5361 gnd.n4631 0.152939
R17873 gnd.n5389 gnd.n4631 0.152939
R17874 gnd.n5390 gnd.n5389 0.152939
R17875 gnd.n5391 gnd.n5390 0.152939
R17876 gnd.n5392 gnd.n5391 0.152939
R17877 gnd.n5392 gnd.n4607 0.152939
R17878 gnd.n5435 gnd.n4607 0.152939
R17879 gnd.n5436 gnd.n5435 0.152939
R17880 gnd.n5437 gnd.n5436 0.152939
R17881 gnd.n5438 gnd.n5437 0.152939
R17882 gnd.n5438 gnd.n4577 0.152939
R17883 gnd.n5756 gnd.n4577 0.152939
R17884 gnd.n5757 gnd.n5756 0.152939
R17885 gnd.n5758 gnd.n5757 0.152939
R17886 gnd.n5759 gnd.n5758 0.152939
R17887 gnd.n5761 gnd.n5759 0.152939
R17888 gnd.n5761 gnd.n5760 0.152939
R17889 gnd.n5760 gnd.n783 0.152939
R17890 gnd.n784 gnd.n783 0.152939
R17891 gnd.n785 gnd.n784 0.152939
R17892 gnd.n4487 gnd.n785 0.152939
R17893 gnd.n4488 gnd.n4487 0.152939
R17894 gnd.n5871 gnd.n4488 0.152939
R17895 gnd.n5152 gnd.n4808 0.152939
R17896 gnd.n4829 gnd.n4808 0.152939
R17897 gnd.n4830 gnd.n4829 0.152939
R17898 gnd.n4836 gnd.n4830 0.152939
R17899 gnd.n4837 gnd.n4836 0.152939
R17900 gnd.n4838 gnd.n4837 0.152939
R17901 gnd.n4838 gnd.n4827 0.152939
R17902 gnd.n4846 gnd.n4827 0.152939
R17903 gnd.n4847 gnd.n4846 0.152939
R17904 gnd.n4848 gnd.n4847 0.152939
R17905 gnd.n4848 gnd.n4825 0.152939
R17906 gnd.n4856 gnd.n4825 0.152939
R17907 gnd.n4857 gnd.n4856 0.152939
R17908 gnd.n4858 gnd.n4857 0.152939
R17909 gnd.n4858 gnd.n4823 0.152939
R17910 gnd.n4866 gnd.n4823 0.152939
R17911 gnd.n5838 gnd.n4519 0.152939
R17912 gnd.n4521 gnd.n4519 0.152939
R17913 gnd.n4525 gnd.n4521 0.152939
R17914 gnd.n4526 gnd.n4525 0.152939
R17915 gnd.n4527 gnd.n4526 0.152939
R17916 gnd.n4528 gnd.n4527 0.152939
R17917 gnd.n4532 gnd.n4528 0.152939
R17918 gnd.n4533 gnd.n4532 0.152939
R17919 gnd.n4534 gnd.n4533 0.152939
R17920 gnd.n4535 gnd.n4534 0.152939
R17921 gnd.n4539 gnd.n4535 0.152939
R17922 gnd.n4540 gnd.n4539 0.152939
R17923 gnd.n4541 gnd.n4540 0.152939
R17924 gnd.n4542 gnd.n4541 0.152939
R17925 gnd.n4546 gnd.n4542 0.152939
R17926 gnd.n4547 gnd.n4546 0.152939
R17927 gnd.n4548 gnd.n4547 0.152939
R17928 gnd.n4549 gnd.n4548 0.152939
R17929 gnd.n4553 gnd.n4549 0.152939
R17930 gnd.n4554 gnd.n4553 0.152939
R17931 gnd.n4555 gnd.n4554 0.152939
R17932 gnd.n4556 gnd.n4555 0.152939
R17933 gnd.n4563 gnd.n4556 0.152939
R17934 gnd.n4564 gnd.n4563 0.152939
R17935 gnd.n4565 gnd.n4564 0.152939
R17936 gnd.n5790 gnd.n4565 0.152939
R17937 gnd.n5325 gnd.n4669 0.152939
R17938 gnd.n5326 gnd.n5325 0.152939
R17939 gnd.n5327 gnd.n5326 0.152939
R17940 gnd.n5328 gnd.n5327 0.152939
R17941 gnd.n5329 gnd.n5328 0.152939
R17942 gnd.n5330 gnd.n5329 0.152939
R17943 gnd.n5331 gnd.n5330 0.152939
R17944 gnd.n5332 gnd.n5331 0.152939
R17945 gnd.n5333 gnd.n5332 0.152939
R17946 gnd.n5333 gnd.n4613 0.152939
R17947 gnd.n5412 gnd.n4613 0.152939
R17948 gnd.n5413 gnd.n5412 0.152939
R17949 gnd.n5414 gnd.n5413 0.152939
R17950 gnd.n5415 gnd.n5414 0.152939
R17951 gnd.n5416 gnd.n5415 0.152939
R17952 gnd.n5417 gnd.n5416 0.152939
R17953 gnd.n5418 gnd.n5417 0.152939
R17954 gnd.n5419 gnd.n5418 0.152939
R17955 gnd.n5419 gnd.n4570 0.152939
R17956 gnd.n5771 gnd.n4570 0.152939
R17957 gnd.n5772 gnd.n5771 0.152939
R17958 gnd.n5773 gnd.n5772 0.152939
R17959 gnd.n5773 gnd.n4568 0.152939
R17960 gnd.n5781 gnd.n4568 0.152939
R17961 gnd.n5782 gnd.n5781 0.152939
R17962 gnd.n5783 gnd.n5782 0.152939
R17963 gnd.n5783 gnd.n4566 0.152939
R17964 gnd.n5789 gnd.n4566 0.152939
R17965 gnd.n4996 gnd.n4995 0.152939
R17966 gnd.n4996 gnd.n4886 0.152939
R17967 gnd.n5011 gnd.n4886 0.152939
R17968 gnd.n5012 gnd.n5011 0.152939
R17969 gnd.n5013 gnd.n5012 0.152939
R17970 gnd.n5013 gnd.n4874 0.152939
R17971 gnd.n5027 gnd.n4874 0.152939
R17972 gnd.n5028 gnd.n5027 0.152939
R17973 gnd.n5029 gnd.n5028 0.152939
R17974 gnd.n5030 gnd.n5029 0.152939
R17975 gnd.n5031 gnd.n5030 0.152939
R17976 gnd.n5032 gnd.n5031 0.152939
R17977 gnd.n5033 gnd.n5032 0.152939
R17978 gnd.n5034 gnd.n5033 0.152939
R17979 gnd.n5035 gnd.n5034 0.152939
R17980 gnd.n5036 gnd.n5035 0.152939
R17981 gnd.n5037 gnd.n5036 0.152939
R17982 gnd.n5038 gnd.n5037 0.152939
R17983 gnd.n5039 gnd.n5038 0.152939
R17984 gnd.n5040 gnd.n5039 0.152939
R17985 gnd.n5041 gnd.n5040 0.152939
R17986 gnd.n5042 gnd.n5041 0.152939
R17987 gnd.n5043 gnd.n5042 0.152939
R17988 gnd.n5044 gnd.n5043 0.152939
R17989 gnd.n5045 gnd.n5044 0.152939
R17990 gnd.n5046 gnd.n5045 0.152939
R17991 gnd.n5047 gnd.n5046 0.152939
R17992 gnd.n5048 gnd.n5047 0.152939
R17993 gnd.n4914 gnd.n4913 0.152939
R17994 gnd.n4915 gnd.n4914 0.152939
R17995 gnd.n4916 gnd.n4915 0.152939
R17996 gnd.n4917 gnd.n4916 0.152939
R17997 gnd.n4918 gnd.n4917 0.152939
R17998 gnd.n4919 gnd.n4918 0.152939
R17999 gnd.n4920 gnd.n4919 0.152939
R18000 gnd.n4921 gnd.n4920 0.152939
R18001 gnd.n4922 gnd.n4921 0.152939
R18002 gnd.n4923 gnd.n4922 0.152939
R18003 gnd.n4924 gnd.n4923 0.152939
R18004 gnd.n4925 gnd.n4924 0.152939
R18005 gnd.n4926 gnd.n4925 0.152939
R18006 gnd.n4927 gnd.n4926 0.152939
R18007 gnd.n4928 gnd.n4927 0.152939
R18008 gnd.n4929 gnd.n4928 0.152939
R18009 gnd.n4930 gnd.n4929 0.152939
R18010 gnd.n4931 gnd.n4930 0.152939
R18011 gnd.n4932 gnd.n4931 0.152939
R18012 gnd.n4933 gnd.n4932 0.152939
R18013 gnd.n4934 gnd.n4933 0.152939
R18014 gnd.n4935 gnd.n4934 0.152939
R18015 gnd.n4939 gnd.n4935 0.152939
R18016 gnd.n4940 gnd.n4939 0.152939
R18017 gnd.n4940 gnd.n4897 0.152939
R18018 gnd.n4994 gnd.n4897 0.152939
R18019 gnd.n6069 gnd.n6068 0.152939
R18020 gnd.n6070 gnd.n6069 0.152939
R18021 gnd.n6070 gnd.n589 0.152939
R18022 gnd.n6078 gnd.n589 0.152939
R18023 gnd.n6079 gnd.n6078 0.152939
R18024 gnd.n6080 gnd.n6079 0.152939
R18025 gnd.n6080 gnd.n583 0.152939
R18026 gnd.n6088 gnd.n583 0.152939
R18027 gnd.n6089 gnd.n6088 0.152939
R18028 gnd.n6090 gnd.n6089 0.152939
R18029 gnd.n6090 gnd.n577 0.152939
R18030 gnd.n6098 gnd.n577 0.152939
R18031 gnd.n6099 gnd.n6098 0.152939
R18032 gnd.n6100 gnd.n6099 0.152939
R18033 gnd.n6100 gnd.n571 0.152939
R18034 gnd.n6108 gnd.n571 0.152939
R18035 gnd.n6109 gnd.n6108 0.152939
R18036 gnd.n6110 gnd.n6109 0.152939
R18037 gnd.n6110 gnd.n565 0.152939
R18038 gnd.n6118 gnd.n565 0.152939
R18039 gnd.n6119 gnd.n6118 0.152939
R18040 gnd.n6120 gnd.n6119 0.152939
R18041 gnd.n6120 gnd.n559 0.152939
R18042 gnd.n6128 gnd.n559 0.152939
R18043 gnd.n6129 gnd.n6128 0.152939
R18044 gnd.n6130 gnd.n6129 0.152939
R18045 gnd.n6130 gnd.n553 0.152939
R18046 gnd.n6138 gnd.n553 0.152939
R18047 gnd.n6139 gnd.n6138 0.152939
R18048 gnd.n6140 gnd.n6139 0.152939
R18049 gnd.n6140 gnd.n547 0.152939
R18050 gnd.n6148 gnd.n547 0.152939
R18051 gnd.n6149 gnd.n6148 0.152939
R18052 gnd.n6150 gnd.n6149 0.152939
R18053 gnd.n6150 gnd.n541 0.152939
R18054 gnd.n6158 gnd.n541 0.152939
R18055 gnd.n6159 gnd.n6158 0.152939
R18056 gnd.n6160 gnd.n6159 0.152939
R18057 gnd.n6160 gnd.n535 0.152939
R18058 gnd.n6168 gnd.n535 0.152939
R18059 gnd.n6169 gnd.n6168 0.152939
R18060 gnd.n6170 gnd.n6169 0.152939
R18061 gnd.n6170 gnd.n529 0.152939
R18062 gnd.n6178 gnd.n529 0.152939
R18063 gnd.n6179 gnd.n6178 0.152939
R18064 gnd.n6180 gnd.n6179 0.152939
R18065 gnd.n6180 gnd.n523 0.152939
R18066 gnd.n6188 gnd.n523 0.152939
R18067 gnd.n6189 gnd.n6188 0.152939
R18068 gnd.n6190 gnd.n6189 0.152939
R18069 gnd.n6190 gnd.n517 0.152939
R18070 gnd.n6198 gnd.n517 0.152939
R18071 gnd.n6199 gnd.n6198 0.152939
R18072 gnd.n6200 gnd.n6199 0.152939
R18073 gnd.n6200 gnd.n511 0.152939
R18074 gnd.n6208 gnd.n511 0.152939
R18075 gnd.n6209 gnd.n6208 0.152939
R18076 gnd.n6210 gnd.n6209 0.152939
R18077 gnd.n6210 gnd.n505 0.152939
R18078 gnd.n6218 gnd.n505 0.152939
R18079 gnd.n6219 gnd.n6218 0.152939
R18080 gnd.n6220 gnd.n6219 0.152939
R18081 gnd.n6220 gnd.n499 0.152939
R18082 gnd.n6228 gnd.n499 0.152939
R18083 gnd.n6229 gnd.n6228 0.152939
R18084 gnd.n6230 gnd.n6229 0.152939
R18085 gnd.n6230 gnd.n493 0.152939
R18086 gnd.n6238 gnd.n493 0.152939
R18087 gnd.n6239 gnd.n6238 0.152939
R18088 gnd.n6240 gnd.n6239 0.152939
R18089 gnd.n6240 gnd.n487 0.152939
R18090 gnd.n6248 gnd.n487 0.152939
R18091 gnd.n6249 gnd.n6248 0.152939
R18092 gnd.n6250 gnd.n6249 0.152939
R18093 gnd.n6250 gnd.n481 0.152939
R18094 gnd.n6258 gnd.n481 0.152939
R18095 gnd.n6259 gnd.n6258 0.152939
R18096 gnd.n6260 gnd.n6259 0.152939
R18097 gnd.n6260 gnd.n475 0.152939
R18098 gnd.n6268 gnd.n475 0.152939
R18099 gnd.n6269 gnd.n6268 0.152939
R18100 gnd.n6270 gnd.n6269 0.152939
R18101 gnd.n6270 gnd.n469 0.152939
R18102 gnd.n6278 gnd.n469 0.152939
R18103 gnd.n6279 gnd.n6278 0.152939
R18104 gnd.n6280 gnd.n6279 0.152939
R18105 gnd.n6280 gnd.n463 0.152939
R18106 gnd.n6288 gnd.n463 0.152939
R18107 gnd.n6289 gnd.n6288 0.152939
R18108 gnd.n6290 gnd.n6289 0.152939
R18109 gnd.n6290 gnd.n457 0.152939
R18110 gnd.n6298 gnd.n457 0.152939
R18111 gnd.n6299 gnd.n6298 0.152939
R18112 gnd.n6300 gnd.n6299 0.152939
R18113 gnd.n6300 gnd.n451 0.152939
R18114 gnd.n6308 gnd.n451 0.152939
R18115 gnd.n6309 gnd.n6308 0.152939
R18116 gnd.n6310 gnd.n6309 0.152939
R18117 gnd.n6310 gnd.n445 0.152939
R18118 gnd.n6318 gnd.n445 0.152939
R18119 gnd.n6319 gnd.n6318 0.152939
R18120 gnd.n6320 gnd.n6319 0.152939
R18121 gnd.n6320 gnd.n439 0.152939
R18122 gnd.n6328 gnd.n439 0.152939
R18123 gnd.n6329 gnd.n6328 0.152939
R18124 gnd.n6330 gnd.n6329 0.152939
R18125 gnd.n6330 gnd.n433 0.152939
R18126 gnd.n6338 gnd.n433 0.152939
R18127 gnd.n6339 gnd.n6338 0.152939
R18128 gnd.n6340 gnd.n6339 0.152939
R18129 gnd.n6340 gnd.n427 0.152939
R18130 gnd.n6348 gnd.n427 0.152939
R18131 gnd.n6349 gnd.n6348 0.152939
R18132 gnd.n6350 gnd.n6349 0.152939
R18133 gnd.n6350 gnd.n421 0.152939
R18134 gnd.n6358 gnd.n421 0.152939
R18135 gnd.n6359 gnd.n6358 0.152939
R18136 gnd.n6360 gnd.n6359 0.152939
R18137 gnd.n6360 gnd.n415 0.152939
R18138 gnd.n6368 gnd.n415 0.152939
R18139 gnd.n6369 gnd.n6368 0.152939
R18140 gnd.n6370 gnd.n6369 0.152939
R18141 gnd.n6370 gnd.n409 0.152939
R18142 gnd.n6378 gnd.n409 0.152939
R18143 gnd.n6379 gnd.n6378 0.152939
R18144 gnd.n6380 gnd.n6379 0.152939
R18145 gnd.n6380 gnd.n403 0.152939
R18146 gnd.n6388 gnd.n403 0.152939
R18147 gnd.n6389 gnd.n6388 0.152939
R18148 gnd.n6390 gnd.n6389 0.152939
R18149 gnd.n6390 gnd.n397 0.152939
R18150 gnd.n6398 gnd.n397 0.152939
R18151 gnd.n6399 gnd.n6398 0.152939
R18152 gnd.n6400 gnd.n6399 0.152939
R18153 gnd.n6400 gnd.n391 0.152939
R18154 gnd.n6408 gnd.n391 0.152939
R18155 gnd.n6409 gnd.n6408 0.152939
R18156 gnd.n6411 gnd.n6409 0.152939
R18157 gnd.n6411 gnd.n6410 0.152939
R18158 gnd.n6410 gnd.n385 0.152939
R18159 gnd.n6420 gnd.n385 0.152939
R18160 gnd.n6421 gnd.n380 0.152939
R18161 gnd.n6429 gnd.n380 0.152939
R18162 gnd.n6430 gnd.n6429 0.152939
R18163 gnd.n6431 gnd.n6430 0.152939
R18164 gnd.n6431 gnd.n374 0.152939
R18165 gnd.n6439 gnd.n374 0.152939
R18166 gnd.n6440 gnd.n6439 0.152939
R18167 gnd.n6441 gnd.n6440 0.152939
R18168 gnd.n6441 gnd.n368 0.152939
R18169 gnd.n6449 gnd.n368 0.152939
R18170 gnd.n6450 gnd.n6449 0.152939
R18171 gnd.n6451 gnd.n6450 0.152939
R18172 gnd.n6451 gnd.n362 0.152939
R18173 gnd.n6459 gnd.n362 0.152939
R18174 gnd.n6460 gnd.n6459 0.152939
R18175 gnd.n6461 gnd.n6460 0.152939
R18176 gnd.n6461 gnd.n356 0.152939
R18177 gnd.n6469 gnd.n356 0.152939
R18178 gnd.n6470 gnd.n6469 0.152939
R18179 gnd.n6471 gnd.n6470 0.152939
R18180 gnd.n6471 gnd.n350 0.152939
R18181 gnd.n6479 gnd.n350 0.152939
R18182 gnd.n6480 gnd.n6479 0.152939
R18183 gnd.n6481 gnd.n6480 0.152939
R18184 gnd.n6481 gnd.n344 0.152939
R18185 gnd.n6489 gnd.n344 0.152939
R18186 gnd.n6490 gnd.n6489 0.152939
R18187 gnd.n6491 gnd.n6490 0.152939
R18188 gnd.n6491 gnd.n338 0.152939
R18189 gnd.n6499 gnd.n338 0.152939
R18190 gnd.n6500 gnd.n6499 0.152939
R18191 gnd.n6501 gnd.n6500 0.152939
R18192 gnd.n6501 gnd.n332 0.152939
R18193 gnd.n6509 gnd.n332 0.152939
R18194 gnd.n6510 gnd.n6509 0.152939
R18195 gnd.n6511 gnd.n6510 0.152939
R18196 gnd.n6511 gnd.n326 0.152939
R18197 gnd.n6519 gnd.n326 0.152939
R18198 gnd.n6520 gnd.n6519 0.152939
R18199 gnd.n6521 gnd.n6520 0.152939
R18200 gnd.n6521 gnd.n320 0.152939
R18201 gnd.n6529 gnd.n320 0.152939
R18202 gnd.n6530 gnd.n6529 0.152939
R18203 gnd.n6531 gnd.n6530 0.152939
R18204 gnd.n6531 gnd.n314 0.152939
R18205 gnd.n6539 gnd.n314 0.152939
R18206 gnd.n6540 gnd.n6539 0.152939
R18207 gnd.n6541 gnd.n6540 0.152939
R18208 gnd.n6541 gnd.n308 0.152939
R18209 gnd.n6549 gnd.n308 0.152939
R18210 gnd.n6550 gnd.n6549 0.152939
R18211 gnd.n6551 gnd.n6550 0.152939
R18212 gnd.n6551 gnd.n302 0.152939
R18213 gnd.n6559 gnd.n302 0.152939
R18214 gnd.n6560 gnd.n6559 0.152939
R18215 gnd.n6561 gnd.n6560 0.152939
R18216 gnd.n6561 gnd.n296 0.152939
R18217 gnd.n6569 gnd.n296 0.152939
R18218 gnd.n6570 gnd.n6569 0.152939
R18219 gnd.n6571 gnd.n6570 0.152939
R18220 gnd.n6571 gnd.n290 0.152939
R18221 gnd.n6579 gnd.n290 0.152939
R18222 gnd.n6580 gnd.n6579 0.152939
R18223 gnd.n6581 gnd.n6580 0.152939
R18224 gnd.n6581 gnd.n284 0.152939
R18225 gnd.n6589 gnd.n284 0.152939
R18226 gnd.n6590 gnd.n6589 0.152939
R18227 gnd.n6591 gnd.n6590 0.152939
R18228 gnd.n6591 gnd.n278 0.152939
R18229 gnd.n6599 gnd.n278 0.152939
R18230 gnd.n6600 gnd.n6599 0.152939
R18231 gnd.n6601 gnd.n6600 0.152939
R18232 gnd.n6601 gnd.n272 0.152939
R18233 gnd.n6609 gnd.n272 0.152939
R18234 gnd.n6610 gnd.n6609 0.152939
R18235 gnd.n6611 gnd.n6610 0.152939
R18236 gnd.n6611 gnd.n266 0.152939
R18237 gnd.n6619 gnd.n266 0.152939
R18238 gnd.n6620 gnd.n6619 0.152939
R18239 gnd.n6621 gnd.n6620 0.152939
R18240 gnd.n6621 gnd.n260 0.152939
R18241 gnd.n6630 gnd.n260 0.152939
R18242 gnd.n6631 gnd.n6630 0.152939
R18243 gnd.n6633 gnd.n6631 0.152939
R18244 gnd.n6675 gnd.n6674 0.152939
R18245 gnd.n6676 gnd.n6675 0.152939
R18246 gnd.n6676 gnd.n198 0.152939
R18247 gnd.n6690 gnd.n198 0.152939
R18248 gnd.n6691 gnd.n6690 0.152939
R18249 gnd.n6692 gnd.n6691 0.152939
R18250 gnd.n6692 gnd.n182 0.152939
R18251 gnd.n6706 gnd.n182 0.152939
R18252 gnd.n6707 gnd.n6706 0.152939
R18253 gnd.n6708 gnd.n6707 0.152939
R18254 gnd.n6708 gnd.n166 0.152939
R18255 gnd.n6796 gnd.n166 0.152939
R18256 gnd.n6797 gnd.n6796 0.152939
R18257 gnd.n6798 gnd.n6797 0.152939
R18258 gnd.n6798 gnd.n88 0.152939
R18259 gnd.n6878 gnd.n88 0.152939
R18260 gnd.n6877 gnd.n89 0.152939
R18261 gnd.n91 gnd.n89 0.152939
R18262 gnd.n95 gnd.n91 0.152939
R18263 gnd.n96 gnd.n95 0.152939
R18264 gnd.n97 gnd.n96 0.152939
R18265 gnd.n98 gnd.n97 0.152939
R18266 gnd.n102 gnd.n98 0.152939
R18267 gnd.n103 gnd.n102 0.152939
R18268 gnd.n104 gnd.n103 0.152939
R18269 gnd.n105 gnd.n104 0.152939
R18270 gnd.n109 gnd.n105 0.152939
R18271 gnd.n110 gnd.n109 0.152939
R18272 gnd.n111 gnd.n110 0.152939
R18273 gnd.n112 gnd.n111 0.152939
R18274 gnd.n116 gnd.n112 0.152939
R18275 gnd.n117 gnd.n116 0.152939
R18276 gnd.n118 gnd.n117 0.152939
R18277 gnd.n119 gnd.n118 0.152939
R18278 gnd.n123 gnd.n119 0.152939
R18279 gnd.n124 gnd.n123 0.152939
R18280 gnd.n125 gnd.n124 0.152939
R18281 gnd.n126 gnd.n125 0.152939
R18282 gnd.n130 gnd.n126 0.152939
R18283 gnd.n131 gnd.n130 0.152939
R18284 gnd.n132 gnd.n131 0.152939
R18285 gnd.n133 gnd.n132 0.152939
R18286 gnd.n137 gnd.n133 0.152939
R18287 gnd.n138 gnd.n137 0.152939
R18288 gnd.n139 gnd.n138 0.152939
R18289 gnd.n140 gnd.n139 0.152939
R18290 gnd.n144 gnd.n140 0.152939
R18291 gnd.n145 gnd.n144 0.152939
R18292 gnd.n146 gnd.n145 0.152939
R18293 gnd.n147 gnd.n146 0.152939
R18294 gnd.n151 gnd.n147 0.152939
R18295 gnd.n152 gnd.n151 0.152939
R18296 gnd.n6808 gnd.n152 0.152939
R18297 gnd.n6808 gnd.n6807 0.152939
R18298 gnd.n3887 gnd.n3886 0.152939
R18299 gnd.n3887 gnd.n1329 0.152939
R18300 gnd.n3902 gnd.n1329 0.152939
R18301 gnd.n3903 gnd.n3902 0.152939
R18302 gnd.n3904 gnd.n3903 0.152939
R18303 gnd.n3905 gnd.n3904 0.152939
R18304 gnd.n3906 gnd.n3905 0.152939
R18305 gnd.n3907 gnd.n3906 0.152939
R18306 gnd.n3908 gnd.n3907 0.152939
R18307 gnd.n3909 gnd.n3908 0.152939
R18308 gnd.n3910 gnd.n3909 0.152939
R18309 gnd.n3911 gnd.n3910 0.152939
R18310 gnd.n3912 gnd.n3911 0.152939
R18311 gnd.n3913 gnd.n3912 0.152939
R18312 gnd.n3914 gnd.n3913 0.152939
R18313 gnd.n3915 gnd.n3914 0.152939
R18314 gnd.n3916 gnd.n3915 0.152939
R18315 gnd.n3917 gnd.n3916 0.152939
R18316 gnd.n3918 gnd.n3917 0.152939
R18317 gnd.n3919 gnd.n3918 0.152939
R18318 gnd.n3919 gnd.n240 0.152939
R18319 gnd.n3920 gnd.n240 0.152939
R18320 gnd.n3921 gnd.n3920 0.152939
R18321 gnd.n3922 gnd.n3921 0.152939
R18322 gnd.n3923 gnd.n3922 0.152939
R18323 gnd.n3924 gnd.n3923 0.152939
R18324 gnd.n3925 gnd.n3924 0.152939
R18325 gnd.n3926 gnd.n3925 0.152939
R18326 gnd.n3927 gnd.n3926 0.152939
R18327 gnd.n3928 gnd.n3927 0.152939
R18328 gnd.n3929 gnd.n3928 0.152939
R18329 gnd.n3930 gnd.n3929 0.152939
R18330 gnd.n3931 gnd.n3930 0.152939
R18331 gnd.n3932 gnd.n3931 0.152939
R18332 gnd.n3933 gnd.n3932 0.152939
R18333 gnd.n3934 gnd.n3933 0.152939
R18334 gnd.n3935 gnd.n3934 0.152939
R18335 gnd.n3936 gnd.n3935 0.152939
R18336 gnd.n3938 gnd.n3936 0.152939
R18337 gnd.n3938 gnd.n3937 0.152939
R18338 gnd.n3937 gnd.n158 0.152939
R18339 gnd.n6806 gnd.n158 0.152939
R18340 gnd.n3791 gnd.n3790 0.152939
R18341 gnd.n3791 gnd.n3787 0.152939
R18342 gnd.n3799 gnd.n3787 0.152939
R18343 gnd.n3800 gnd.n3799 0.152939
R18344 gnd.n3801 gnd.n3800 0.152939
R18345 gnd.n3801 gnd.n3783 0.152939
R18346 gnd.n3809 gnd.n3783 0.152939
R18347 gnd.n3810 gnd.n3809 0.152939
R18348 gnd.n3811 gnd.n3810 0.152939
R18349 gnd.n3811 gnd.n3779 0.152939
R18350 gnd.n3819 gnd.n3779 0.152939
R18351 gnd.n3820 gnd.n3819 0.152939
R18352 gnd.n3822 gnd.n3820 0.152939
R18353 gnd.n3822 gnd.n3821 0.152939
R18354 gnd.n3821 gnd.n1359 0.152939
R18355 gnd.n3835 gnd.n3834 0.152939
R18356 gnd.n3835 gnd.n1355 0.152939
R18357 gnd.n3843 gnd.n1355 0.152939
R18358 gnd.n3844 gnd.n3843 0.152939
R18359 gnd.n3845 gnd.n3844 0.152939
R18360 gnd.n3845 gnd.n1351 0.152939
R18361 gnd.n3853 gnd.n1351 0.152939
R18362 gnd.n3854 gnd.n3853 0.152939
R18363 gnd.n3855 gnd.n3854 0.152939
R18364 gnd.n3855 gnd.n1347 0.152939
R18365 gnd.n3863 gnd.n1347 0.152939
R18366 gnd.n3864 gnd.n3863 0.152939
R18367 gnd.n3865 gnd.n3864 0.152939
R18368 gnd.n3865 gnd.n1343 0.152939
R18369 gnd.n3873 gnd.n1343 0.152939
R18370 gnd.n3874 gnd.n3873 0.152939
R18371 gnd.n3876 gnd.n3874 0.152939
R18372 gnd.n3876 gnd.n3875 0.152939
R18373 gnd.n3875 gnd.n1336 0.152939
R18374 gnd.n3885 gnd.n1336 0.152939
R18375 gnd.n1220 gnd.n1219 0.152939
R18376 gnd.n1221 gnd.n1220 0.152939
R18377 gnd.n1324 gnd.n1221 0.152939
R18378 gnd.n4013 gnd.n1324 0.152939
R18379 gnd.n4014 gnd.n4013 0.152939
R18380 gnd.n4015 gnd.n4014 0.152939
R18381 gnd.n4016 gnd.n4015 0.152939
R18382 gnd.n4016 gnd.n1296 0.152939
R18383 gnd.n4044 gnd.n1296 0.152939
R18384 gnd.n4045 gnd.n4044 0.152939
R18385 gnd.n4046 gnd.n4045 0.152939
R18386 gnd.n4048 gnd.n4046 0.152939
R18387 gnd.n4048 gnd.n4047 0.152939
R18388 gnd.n4047 gnd.n1268 0.152939
R18389 gnd.n1268 gnd.n212 0.152939
R18390 gnd.n6674 gnd.n212 0.152939
R18391 gnd.n4074 gnd.n4068 0.152939
R18392 gnd.n4074 gnd.n4073 0.152939
R18393 gnd.n4073 gnd.n4072 0.152939
R18394 gnd.n4072 gnd.n254 0.152939
R18395 gnd.n256 gnd.n255 0.152939
R18396 gnd.n6632 gnd.n256 0.152939
R18397 gnd.n2477 gnd.n2476 0.152939
R18398 gnd.n2478 gnd.n2477 0.152939
R18399 gnd.n2479 gnd.n2478 0.152939
R18400 gnd.n2480 gnd.n2479 0.152939
R18401 gnd.n2483 gnd.n2480 0.152939
R18402 gnd.n2484 gnd.n2483 0.152939
R18403 gnd.n2485 gnd.n2484 0.152939
R18404 gnd.n2486 gnd.n2485 0.152939
R18405 gnd.n2488 gnd.n2486 0.152939
R18406 gnd.n2488 gnd.n2487 0.152939
R18407 gnd.n2487 gnd.n2217 0.152939
R18408 gnd.n2560 gnd.n2217 0.152939
R18409 gnd.n2561 gnd.n2560 0.152939
R18410 gnd.n2562 gnd.n2561 0.152939
R18411 gnd.n2562 gnd.n2213 0.152939
R18412 gnd.n2568 gnd.n2213 0.152939
R18413 gnd.n2569 gnd.n2568 0.152939
R18414 gnd.n2570 gnd.n2569 0.152939
R18415 gnd.n2570 gnd.n2209 0.152939
R18416 gnd.n2580 gnd.n2209 0.152939
R18417 gnd.n2581 gnd.n2580 0.152939
R18418 gnd.n2582 gnd.n2581 0.152939
R18419 gnd.n2582 gnd.n2071 0.152939
R18420 gnd.n2593 gnd.n2071 0.152939
R18421 gnd.n2594 gnd.n2593 0.152939
R18422 gnd.n2595 gnd.n2594 0.152939
R18423 gnd.n2595 gnd.n2065 0.152939
R18424 gnd.n2608 gnd.n2065 0.152939
R18425 gnd.n2609 gnd.n2608 0.152939
R18426 gnd.n2610 gnd.n2609 0.152939
R18427 gnd.n2611 gnd.n2610 0.152939
R18428 gnd.n2612 gnd.n2611 0.152939
R18429 gnd.n2613 gnd.n2612 0.152939
R18430 gnd.n2613 gnd.n1771 0.152939
R18431 gnd.n2803 gnd.n1771 0.152939
R18432 gnd.n2804 gnd.n2803 0.152939
R18433 gnd.n2805 gnd.n2804 0.152939
R18434 gnd.n2805 gnd.n1743 0.152939
R18435 gnd.n2846 gnd.n1743 0.152939
R18436 gnd.n2847 gnd.n2846 0.152939
R18437 gnd.n2848 gnd.n2847 0.152939
R18438 gnd.n2848 gnd.n1725 0.152939
R18439 gnd.n2888 gnd.n1725 0.152939
R18440 gnd.n2889 gnd.n2888 0.152939
R18441 gnd.n2890 gnd.n2889 0.152939
R18442 gnd.n2891 gnd.n2890 0.152939
R18443 gnd.n2891 gnd.n1699 0.152939
R18444 gnd.n2950 gnd.n1699 0.152939
R18445 gnd.n2951 gnd.n2950 0.152939
R18446 gnd.n2952 gnd.n2951 0.152939
R18447 gnd.n2952 gnd.n1681 0.152939
R18448 gnd.n2977 gnd.n1681 0.152939
R18449 gnd.n2978 gnd.n2977 0.152939
R18450 gnd.n2979 gnd.n2978 0.152939
R18451 gnd.n2980 gnd.n2979 0.152939
R18452 gnd.n2980 gnd.n1648 0.152939
R18453 gnd.n3028 gnd.n1648 0.152939
R18454 gnd.n3029 gnd.n3028 0.152939
R18455 gnd.n3030 gnd.n3029 0.152939
R18456 gnd.n3030 gnd.n1625 0.152939
R18457 gnd.n3068 gnd.n1625 0.152939
R18458 gnd.n3069 gnd.n3068 0.152939
R18459 gnd.n3070 gnd.n3069 0.152939
R18460 gnd.n3070 gnd.n1603 0.152939
R18461 gnd.n3124 gnd.n1603 0.152939
R18462 gnd.n3125 gnd.n3124 0.152939
R18463 gnd.n3126 gnd.n3125 0.152939
R18464 gnd.n3126 gnd.n1584 0.152939
R18465 gnd.n3149 gnd.n1584 0.152939
R18466 gnd.n3150 gnd.n3149 0.152939
R18467 gnd.n3151 gnd.n3150 0.152939
R18468 gnd.n3151 gnd.n1564 0.152939
R18469 gnd.n3209 gnd.n1564 0.152939
R18470 gnd.n3210 gnd.n3209 0.152939
R18471 gnd.n3211 gnd.n3210 0.152939
R18472 gnd.n3211 gnd.n1542 0.152939
R18473 gnd.n3238 gnd.n1542 0.152939
R18474 gnd.n3239 gnd.n3238 0.152939
R18475 gnd.n3240 gnd.n3239 0.152939
R18476 gnd.n3241 gnd.n3240 0.152939
R18477 gnd.n3241 gnd.n1514 0.152939
R18478 gnd.n3291 gnd.n1514 0.152939
R18479 gnd.n3292 gnd.n3291 0.152939
R18480 gnd.n3293 gnd.n3292 0.152939
R18481 gnd.n3293 gnd.n1495 0.152939
R18482 gnd.n3318 gnd.n1495 0.152939
R18483 gnd.n3319 gnd.n3318 0.152939
R18484 gnd.n3320 gnd.n3319 0.152939
R18485 gnd.n3321 gnd.n3320 0.152939
R18486 gnd.n3321 gnd.n1465 0.152939
R18487 gnd.n3362 gnd.n1465 0.152939
R18488 gnd.n3363 gnd.n3362 0.152939
R18489 gnd.n3364 gnd.n3363 0.152939
R18490 gnd.n3366 gnd.n3364 0.152939
R18491 gnd.n3366 gnd.n3365 0.152939
R18492 gnd.n3365 gnd.n1414 0.152939
R18493 gnd.n1415 gnd.n1414 0.152939
R18494 gnd.n1416 gnd.n1415 0.152939
R18495 gnd.n1426 gnd.n1416 0.152939
R18496 gnd.n1427 gnd.n1426 0.152939
R18497 gnd.n1428 gnd.n1427 0.152939
R18498 gnd.n1429 gnd.n1428 0.152939
R18499 gnd.n1430 gnd.n1429 0.152939
R18500 gnd.n1432 gnd.n1430 0.152939
R18501 gnd.n1432 gnd.n1431 0.152939
R18502 gnd.n1431 gnd.n1198 0.152939
R18503 gnd.n1199 gnd.n1198 0.152939
R18504 gnd.n1200 gnd.n1199 0.152939
R18505 gnd.n1206 gnd.n1200 0.152939
R18506 gnd.n1207 gnd.n1206 0.152939
R18507 gnd.n1208 gnd.n1207 0.152939
R18508 gnd.n1209 gnd.n1208 0.152939
R18509 gnd.n3996 gnd.n1209 0.152939
R18510 gnd.n3997 gnd.n3996 0.152939
R18511 gnd.n4002 gnd.n3997 0.152939
R18512 gnd.n4003 gnd.n4002 0.152939
R18513 gnd.n4004 gnd.n4003 0.152939
R18514 gnd.n4005 gnd.n4004 0.152939
R18515 gnd.n4005 gnd.n1306 0.152939
R18516 gnd.n4033 gnd.n1306 0.152939
R18517 gnd.n4034 gnd.n4033 0.152939
R18518 gnd.n4035 gnd.n4034 0.152939
R18519 gnd.n4036 gnd.n4035 0.152939
R18520 gnd.n4036 gnd.n1278 0.152939
R18521 gnd.n4065 gnd.n1278 0.152939
R18522 gnd.n4066 gnd.n4065 0.152939
R18523 gnd.n4067 gnd.n4066 0.152939
R18524 gnd.n4068 gnd.n4067 0.152939
R18525 gnd.n2297 gnd.n2295 0.152939
R18526 gnd.n2295 gnd.n2269 0.152939
R18527 gnd.n2356 gnd.n2269 0.152939
R18528 gnd.n2357 gnd.n2356 0.152939
R18529 gnd.n2358 gnd.n2357 0.152939
R18530 gnd.n2358 gnd.n2266 0.152939
R18531 gnd.n2363 gnd.n2266 0.152939
R18532 gnd.n2364 gnd.n2363 0.152939
R18533 gnd.n2365 gnd.n2364 0.152939
R18534 gnd.n2365 gnd.n2263 0.152939
R18535 gnd.n2370 gnd.n2263 0.152939
R18536 gnd.n2371 gnd.n2370 0.152939
R18537 gnd.n2372 gnd.n2371 0.152939
R18538 gnd.n2372 gnd.n2260 0.152939
R18539 gnd.n2377 gnd.n2260 0.152939
R18540 gnd.n2378 gnd.n2377 0.152939
R18541 gnd.n2379 gnd.n2378 0.152939
R18542 gnd.n2379 gnd.n2258 0.152939
R18543 gnd.n2426 gnd.n2258 0.152939
R18544 gnd.n2427 gnd.n2426 0.152939
R18545 gnd.n2336 gnd.n2276 0.152939
R18546 gnd.n2277 gnd.n2276 0.152939
R18547 gnd.n2278 gnd.n2277 0.152939
R18548 gnd.n2279 gnd.n2278 0.152939
R18549 gnd.n2280 gnd.n2279 0.152939
R18550 gnd.n2281 gnd.n2280 0.152939
R18551 gnd.n2282 gnd.n2281 0.152939
R18552 gnd.n2283 gnd.n2282 0.152939
R18553 gnd.n2284 gnd.n2283 0.152939
R18554 gnd.n2285 gnd.n2284 0.152939
R18555 gnd.n2286 gnd.n2285 0.152939
R18556 gnd.n2287 gnd.n2286 0.152939
R18557 gnd.n2288 gnd.n2287 0.152939
R18558 gnd.n2289 gnd.n2288 0.152939
R18559 gnd.n2290 gnd.n2289 0.152939
R18560 gnd.n2301 gnd.n2290 0.152939
R18561 gnd.n2301 gnd.n2300 0.152939
R18562 gnd.n2300 gnd.n2299 0.152939
R18563 gnd.n2342 gnd.n2337 0.152939
R18564 gnd.n2342 gnd.n2341 0.152939
R18565 gnd.n2341 gnd.n2340 0.152939
R18566 gnd.n2340 gnd.n2338 0.152939
R18567 gnd.n2338 gnd.n902 0.152939
R18568 gnd.n903 gnd.n902 0.152939
R18569 gnd.n904 gnd.n903 0.152939
R18570 gnd.n920 gnd.n904 0.152939
R18571 gnd.n921 gnd.n920 0.152939
R18572 gnd.n922 gnd.n921 0.152939
R18573 gnd.n923 gnd.n922 0.152939
R18574 gnd.n941 gnd.n923 0.152939
R18575 gnd.n942 gnd.n941 0.152939
R18576 gnd.n943 gnd.n942 0.152939
R18577 gnd.n944 gnd.n943 0.152939
R18578 gnd.n964 gnd.n944 0.152939
R18579 gnd.n965 gnd.n964 0.152939
R18580 gnd.n966 gnd.n965 0.152939
R18581 gnd.n967 gnd.n966 0.152939
R18582 gnd.n968 gnd.n967 0.152939
R18583 gnd.n2255 gnd.n968 0.152939
R18584 gnd.n2255 gnd.n982 0.152939
R18585 gnd.n983 gnd.n982 0.152939
R18586 gnd.n984 gnd.n983 0.152939
R18587 gnd.n1000 gnd.n984 0.152939
R18588 gnd.n1001 gnd.n1000 0.152939
R18589 gnd.n1002 gnd.n1001 0.152939
R18590 gnd.n1003 gnd.n1002 0.152939
R18591 gnd.n1020 gnd.n1003 0.152939
R18592 gnd.n1021 gnd.n1020 0.152939
R18593 gnd.n1022 gnd.n1021 0.152939
R18594 gnd.n1023 gnd.n1022 0.152939
R18595 gnd.n1042 gnd.n1023 0.152939
R18596 gnd.n1043 gnd.n1042 0.152939
R18597 gnd.n1044 gnd.n1043 0.152939
R18598 gnd.n1045 gnd.n1044 0.152939
R18599 gnd.n1063 gnd.n1045 0.152939
R18600 gnd.n1064 gnd.n1063 0.152939
R18601 gnd.n1065 gnd.n1064 0.152939
R18602 gnd.n1066 gnd.n1065 0.152939
R18603 gnd.n1084 gnd.n1066 0.152939
R18604 gnd.n4274 gnd.n1084 0.152939
R18605 gnd.n1010 gnd.n953 0.152939
R18606 gnd.n1011 gnd.n1010 0.152939
R18607 gnd.n1012 gnd.n1011 0.152939
R18608 gnd.n1013 gnd.n1012 0.152939
R18609 gnd.n1031 gnd.n1013 0.152939
R18610 gnd.n1032 gnd.n1031 0.152939
R18611 gnd.n1033 gnd.n1032 0.152939
R18612 gnd.n1034 gnd.n1033 0.152939
R18613 gnd.n1052 gnd.n1034 0.152939
R18614 gnd.n1053 gnd.n1052 0.152939
R18615 gnd.n1054 gnd.n1053 0.152939
R18616 gnd.n1055 gnd.n1054 0.152939
R18617 gnd.n1074 gnd.n1055 0.152939
R18618 gnd.n1075 gnd.n1074 0.152939
R18619 gnd.n1076 gnd.n1075 0.152939
R18620 gnd.n1077 gnd.n1076 0.152939
R18621 gnd.n1955 gnd.n1954 0.152939
R18622 gnd.n1956 gnd.n1955 0.152939
R18623 gnd.n1957 gnd.n1956 0.152939
R18624 gnd.n1958 gnd.n1957 0.152939
R18625 gnd.n1959 gnd.n1958 0.152939
R18626 gnd.n1960 gnd.n1959 0.152939
R18627 gnd.n1961 gnd.n1960 0.152939
R18628 gnd.n1962 gnd.n1961 0.152939
R18629 gnd.n1963 gnd.n1962 0.152939
R18630 gnd.n1964 gnd.n1963 0.152939
R18631 gnd.n1965 gnd.n1964 0.152939
R18632 gnd.n1966 gnd.n1965 0.152939
R18633 gnd.n1967 gnd.n1966 0.152939
R18634 gnd.n1968 gnd.n1967 0.152939
R18635 gnd.n1968 gnd.n1938 0.152939
R18636 gnd.n2705 gnd.n2704 0.152939
R18637 gnd.n2704 gnd.n1939 0.152939
R18638 gnd.n1999 gnd.n1939 0.152939
R18639 gnd.n2000 gnd.n1999 0.152939
R18640 gnd.n2001 gnd.n2000 0.152939
R18641 gnd.n2002 gnd.n2001 0.152939
R18642 gnd.n2006 gnd.n2002 0.152939
R18643 gnd.n2007 gnd.n2006 0.152939
R18644 gnd.n2008 gnd.n2007 0.152939
R18645 gnd.n2009 gnd.n2008 0.152939
R18646 gnd.n2013 gnd.n2009 0.152939
R18647 gnd.n2014 gnd.n2013 0.152939
R18648 gnd.n2015 gnd.n2014 0.152939
R18649 gnd.n2016 gnd.n2015 0.152939
R18650 gnd.n2020 gnd.n2016 0.152939
R18651 gnd.n2021 gnd.n2020 0.152939
R18652 gnd.n2022 gnd.n2021 0.152939
R18653 gnd.n2023 gnd.n2022 0.152939
R18654 gnd.n2028 gnd.n2023 0.152939
R18655 gnd.n2667 gnd.n2028 0.152939
R18656 gnd.n4400 gnd.n877 0.152939
R18657 gnd.n4400 gnd.n4399 0.152939
R18658 gnd.n4399 gnd.n4398 0.152939
R18659 gnd.n4398 gnd.n880 0.152939
R18660 gnd.n2390 gnd.n880 0.152939
R18661 gnd.n2390 gnd.n2389 0.152939
R18662 gnd.n2395 gnd.n2389 0.152939
R18663 gnd.n2396 gnd.n2395 0.152939
R18664 gnd.n2397 gnd.n2396 0.152939
R18665 gnd.n2397 gnd.n2386 0.152939
R18666 gnd.n2402 gnd.n2386 0.152939
R18667 gnd.n2403 gnd.n2402 0.152939
R18668 gnd.n2404 gnd.n2403 0.152939
R18669 gnd.n2404 gnd.n2383 0.152939
R18670 gnd.n2409 gnd.n2383 0.152939
R18671 gnd.n2410 gnd.n2409 0.152939
R18672 gnd.n2411 gnd.n2410 0.152939
R18673 gnd.n2412 gnd.n2411 0.152939
R18674 gnd.n2414 gnd.n2412 0.152939
R18675 gnd.n2414 gnd.n2413 0.152939
R18676 gnd.n2413 gnd.n2256 0.152939
R18677 gnd.n2256 gnd.n2253 0.152939
R18678 gnd.n2436 gnd.n2253 0.152939
R18679 gnd.n2437 gnd.n2436 0.152939
R18680 gnd.n2438 gnd.n2437 0.152939
R18681 gnd.n2439 gnd.n2438 0.152939
R18682 gnd.n2440 gnd.n2439 0.152939
R18683 gnd.n2440 gnd.n2237 0.152939
R18684 gnd.n2513 gnd.n2237 0.152939
R18685 gnd.n2514 gnd.n2513 0.152939
R18686 gnd.n2515 gnd.n2514 0.152939
R18687 gnd.n2515 gnd.n2230 0.152939
R18688 gnd.n2529 gnd.n2230 0.152939
R18689 gnd.n2530 gnd.n2529 0.152939
R18690 gnd.n2531 gnd.n2530 0.152939
R18691 gnd.n2531 gnd.n2228 0.152939
R18692 gnd.n2537 gnd.n2228 0.152939
R18693 gnd.n2538 gnd.n2537 0.152939
R18694 gnd.n2540 gnd.n2538 0.152939
R18695 gnd.n2540 gnd.n2539 0.152939
R18696 gnd.n2539 gnd.n2029 0.152939
R18697 gnd.n2666 gnd.n2029 0.152939
R18698 gnd.n835 gnd.n834 0.152939
R18699 gnd.n836 gnd.n835 0.152939
R18700 gnd.n837 gnd.n836 0.152939
R18701 gnd.n838 gnd.n837 0.152939
R18702 gnd.n839 gnd.n838 0.152939
R18703 gnd.n840 gnd.n839 0.152939
R18704 gnd.n841 gnd.n840 0.152939
R18705 gnd.n842 gnd.n841 0.152939
R18706 gnd.n843 gnd.n842 0.152939
R18707 gnd.n844 gnd.n843 0.152939
R18708 gnd.n845 gnd.n844 0.152939
R18709 gnd.n846 gnd.n845 0.152939
R18710 gnd.n847 gnd.n846 0.152939
R18711 gnd.n848 gnd.n847 0.152939
R18712 gnd.n849 gnd.n848 0.152939
R18713 gnd.n850 gnd.n849 0.152939
R18714 gnd.n851 gnd.n850 0.152939
R18715 gnd.n854 gnd.n851 0.152939
R18716 gnd.n855 gnd.n854 0.152939
R18717 gnd.n856 gnd.n855 0.152939
R18718 gnd.n857 gnd.n856 0.152939
R18719 gnd.n858 gnd.n857 0.152939
R18720 gnd.n859 gnd.n858 0.152939
R18721 gnd.n860 gnd.n859 0.152939
R18722 gnd.n861 gnd.n860 0.152939
R18723 gnd.n862 gnd.n861 0.152939
R18724 gnd.n863 gnd.n862 0.152939
R18725 gnd.n864 gnd.n863 0.152939
R18726 gnd.n865 gnd.n864 0.152939
R18727 gnd.n866 gnd.n865 0.152939
R18728 gnd.n867 gnd.n866 0.152939
R18729 gnd.n868 gnd.n867 0.152939
R18730 gnd.n869 gnd.n868 0.152939
R18731 gnd.n870 gnd.n869 0.152939
R18732 gnd.n871 gnd.n870 0.152939
R18733 gnd.n4408 gnd.n871 0.152939
R18734 gnd.n4408 gnd.n4407 0.152939
R18735 gnd.n4407 gnd.n4406 0.152939
R18736 gnd.n2348 gnd.n2346 0.152939
R18737 gnd.n2348 gnd.n2347 0.152939
R18738 gnd.n2347 gnd.n891 0.152939
R18739 gnd.n892 gnd.n891 0.152939
R18740 gnd.n893 gnd.n892 0.152939
R18741 gnd.n911 gnd.n893 0.152939
R18742 gnd.n912 gnd.n911 0.152939
R18743 gnd.n913 gnd.n912 0.152939
R18744 gnd.n914 gnd.n913 0.152939
R18745 gnd.n930 gnd.n914 0.152939
R18746 gnd.n931 gnd.n930 0.152939
R18747 gnd.n932 gnd.n931 0.152939
R18748 gnd.n933 gnd.n932 0.152939
R18749 gnd.n951 gnd.n933 0.152939
R18750 gnd.n952 gnd.n951 0.152939
R18751 gnd.n953 gnd.n952 0.152939
R18752 gnd.n2460 gnd.n2457 0.152939
R18753 gnd.n2467 gnd.n2457 0.152939
R18754 gnd.n2470 gnd.n2469 0.152939
R18755 gnd.n2470 gnd.n2246 0.152939
R18756 gnd.n2476 gnd.n2246 0.152939
R18757 gnd.n600 gnd.n595 0.152939
R18758 gnd.n601 gnd.n600 0.152939
R18759 gnd.n602 gnd.n601 0.152939
R18760 gnd.n607 gnd.n602 0.152939
R18761 gnd.n608 gnd.n607 0.152939
R18762 gnd.n609 gnd.n608 0.152939
R18763 gnd.n610 gnd.n609 0.152939
R18764 gnd.n615 gnd.n610 0.152939
R18765 gnd.n616 gnd.n615 0.152939
R18766 gnd.n617 gnd.n616 0.152939
R18767 gnd.n618 gnd.n617 0.152939
R18768 gnd.n623 gnd.n618 0.152939
R18769 gnd.n624 gnd.n623 0.152939
R18770 gnd.n625 gnd.n624 0.152939
R18771 gnd.n626 gnd.n625 0.152939
R18772 gnd.n631 gnd.n626 0.152939
R18773 gnd.n632 gnd.n631 0.152939
R18774 gnd.n633 gnd.n632 0.152939
R18775 gnd.n634 gnd.n633 0.152939
R18776 gnd.n639 gnd.n634 0.152939
R18777 gnd.n640 gnd.n639 0.152939
R18778 gnd.n641 gnd.n640 0.152939
R18779 gnd.n642 gnd.n641 0.152939
R18780 gnd.n647 gnd.n642 0.152939
R18781 gnd.n648 gnd.n647 0.152939
R18782 gnd.n649 gnd.n648 0.152939
R18783 gnd.n650 gnd.n649 0.152939
R18784 gnd.n655 gnd.n650 0.152939
R18785 gnd.n656 gnd.n655 0.152939
R18786 gnd.n657 gnd.n656 0.152939
R18787 gnd.n658 gnd.n657 0.152939
R18788 gnd.n663 gnd.n658 0.152939
R18789 gnd.n664 gnd.n663 0.152939
R18790 gnd.n665 gnd.n664 0.152939
R18791 gnd.n666 gnd.n665 0.152939
R18792 gnd.n671 gnd.n666 0.152939
R18793 gnd.n672 gnd.n671 0.152939
R18794 gnd.n673 gnd.n672 0.152939
R18795 gnd.n674 gnd.n673 0.152939
R18796 gnd.n679 gnd.n674 0.152939
R18797 gnd.n680 gnd.n679 0.152939
R18798 gnd.n681 gnd.n680 0.152939
R18799 gnd.n682 gnd.n681 0.152939
R18800 gnd.n687 gnd.n682 0.152939
R18801 gnd.n688 gnd.n687 0.152939
R18802 gnd.n689 gnd.n688 0.152939
R18803 gnd.n690 gnd.n689 0.152939
R18804 gnd.n695 gnd.n690 0.152939
R18805 gnd.n696 gnd.n695 0.152939
R18806 gnd.n697 gnd.n696 0.152939
R18807 gnd.n698 gnd.n697 0.152939
R18808 gnd.n703 gnd.n698 0.152939
R18809 gnd.n704 gnd.n703 0.152939
R18810 gnd.n705 gnd.n704 0.152939
R18811 gnd.n706 gnd.n705 0.152939
R18812 gnd.n711 gnd.n706 0.152939
R18813 gnd.n712 gnd.n711 0.152939
R18814 gnd.n713 gnd.n712 0.152939
R18815 gnd.n714 gnd.n713 0.152939
R18816 gnd.n719 gnd.n714 0.152939
R18817 gnd.n720 gnd.n719 0.152939
R18818 gnd.n721 gnd.n720 0.152939
R18819 gnd.n722 gnd.n721 0.152939
R18820 gnd.n727 gnd.n722 0.152939
R18821 gnd.n728 gnd.n727 0.152939
R18822 gnd.n729 gnd.n728 0.152939
R18823 gnd.n730 gnd.n729 0.152939
R18824 gnd.n735 gnd.n730 0.152939
R18825 gnd.n736 gnd.n735 0.152939
R18826 gnd.n737 gnd.n736 0.152939
R18827 gnd.n738 gnd.n737 0.152939
R18828 gnd.n743 gnd.n738 0.152939
R18829 gnd.n744 gnd.n743 0.152939
R18830 gnd.n745 gnd.n744 0.152939
R18831 gnd.n746 gnd.n745 0.152939
R18832 gnd.n751 gnd.n746 0.152939
R18833 gnd.n752 gnd.n751 0.152939
R18834 gnd.n753 gnd.n752 0.152939
R18835 gnd.n754 gnd.n753 0.152939
R18836 gnd.n759 gnd.n754 0.152939
R18837 gnd.n760 gnd.n759 0.152939
R18838 gnd.n761 gnd.n760 0.152939
R18839 gnd.n762 gnd.n761 0.152939
R18840 gnd.n2459 gnd.n762 0.152939
R18841 gnd.n3565 gnd.n3421 0.152939
R18842 gnd.n3566 gnd.n3565 0.152939
R18843 gnd.n3567 gnd.n3566 0.152939
R18844 gnd.n3567 gnd.n3417 0.152939
R18845 gnd.n3578 gnd.n3417 0.152939
R18846 gnd.n3579 gnd.n3578 0.152939
R18847 gnd.n3580 gnd.n3579 0.152939
R18848 gnd.n3580 gnd.n3413 0.152939
R18849 gnd.n3587 gnd.n3413 0.152939
R18850 gnd.n2639 gnd.n2053 0.152939
R18851 gnd.n2635 gnd.n2053 0.152939
R18852 gnd.n2635 gnd.n2634 0.152939
R18853 gnd.n2634 gnd.n2633 0.152939
R18854 gnd.n2633 gnd.n2058 0.152939
R18855 gnd.n2629 gnd.n2058 0.152939
R18856 gnd.n2629 gnd.n2628 0.152939
R18857 gnd.n2628 gnd.n1786 0.152939
R18858 gnd.n2783 gnd.n1786 0.152939
R18859 gnd.n2784 gnd.n2783 0.152939
R18860 gnd.n2786 gnd.n2784 0.152939
R18861 gnd.n2786 gnd.n2785 0.152939
R18862 gnd.n2785 gnd.n1765 0.152939
R18863 gnd.n2814 gnd.n1765 0.152939
R18864 gnd.n2815 gnd.n2814 0.152939
R18865 gnd.n2823 gnd.n2815 0.152939
R18866 gnd.n2823 gnd.n2822 0.152939
R18867 gnd.n2822 gnd.n2821 0.152939
R18868 gnd.n2821 gnd.n2816 0.152939
R18869 gnd.n2816 gnd.n1717 0.152939
R18870 gnd.n2899 gnd.n1717 0.152939
R18871 gnd.n2900 gnd.n2899 0.152939
R18872 gnd.n2921 gnd.n2900 0.152939
R18873 gnd.n2921 gnd.n2920 0.152939
R18874 gnd.n2920 gnd.n2919 0.152939
R18875 gnd.n2919 gnd.n2901 0.152939
R18876 gnd.n2915 gnd.n2901 0.152939
R18877 gnd.n2915 gnd.n2914 0.152939
R18878 gnd.n2914 gnd.n2913 0.152939
R18879 gnd.n2913 gnd.n2910 0.152939
R18880 gnd.n2910 gnd.n2909 0.152939
R18881 gnd.n2909 gnd.n1665 0.152939
R18882 gnd.n3001 gnd.n1665 0.152939
R18883 gnd.n3002 gnd.n3001 0.152939
R18884 gnd.n3003 gnd.n3002 0.152939
R18885 gnd.n3003 gnd.n1641 0.152939
R18886 gnd.n3051 gnd.n1641 0.152939
R18887 gnd.n3051 gnd.n3050 0.152939
R18888 gnd.n3050 gnd.n3049 0.152939
R18889 gnd.n3049 gnd.n1618 0.152939
R18890 gnd.n3109 gnd.n1618 0.152939
R18891 gnd.n3109 gnd.n3108 0.152939
R18892 gnd.n3108 gnd.n3107 0.152939
R18893 gnd.n3107 gnd.n1619 0.152939
R18894 gnd.n3103 gnd.n1619 0.152939
R18895 gnd.n3103 gnd.n3102 0.152939
R18896 gnd.n3102 gnd.n3101 0.152939
R18897 gnd.n3101 gnd.n3092 0.152939
R18898 gnd.n3097 gnd.n3092 0.152939
R18899 gnd.n3097 gnd.n1557 0.152939
R18900 gnd.n3219 gnd.n1557 0.152939
R18901 gnd.n3220 gnd.n3219 0.152939
R18902 gnd.n3222 gnd.n3220 0.152939
R18903 gnd.n3222 gnd.n3221 0.152939
R18904 gnd.n3221 gnd.n1528 0.152939
R18905 gnd.n3258 gnd.n1528 0.152939
R18906 gnd.n3259 gnd.n3258 0.152939
R18907 gnd.n3275 gnd.n3259 0.152939
R18908 gnd.n3275 gnd.n3274 0.152939
R18909 gnd.n3274 gnd.n3273 0.152939
R18910 gnd.n3273 gnd.n3260 0.152939
R18911 gnd.n3269 gnd.n3260 0.152939
R18912 gnd.n3269 gnd.n3268 0.152939
R18913 gnd.n3268 gnd.n3267 0.152939
R18914 gnd.n3267 gnd.n1473 0.152939
R18915 gnd.n3351 gnd.n1473 0.152939
R18916 gnd.n3352 gnd.n3351 0.152939
R18917 gnd.n3354 gnd.n3352 0.152939
R18918 gnd.n3354 gnd.n3353 0.152939
R18919 gnd.n3353 gnd.n1446 0.152939
R18920 gnd.n3393 gnd.n1446 0.152939
R18921 gnd.n3394 gnd.n3393 0.152939
R18922 gnd.n3395 gnd.n3394 0.152939
R18923 gnd.n3395 gnd.n1443 0.152939
R18924 gnd.n3403 gnd.n1443 0.152939
R18925 gnd.n3404 gnd.n3403 0.152939
R18926 gnd.n3405 gnd.n3404 0.152939
R18927 gnd.n3405 gnd.n1441 0.152939
R18928 gnd.n3411 gnd.n1441 0.152939
R18929 gnd.n3412 gnd.n3411 0.152939
R18930 gnd.n3589 gnd.n3412 0.152939
R18931 gnd.n3589 gnd.n3588 0.152939
R18932 gnd.n2652 gnd.n2034 0.152939
R18933 gnd.n2652 gnd.n2651 0.152939
R18934 gnd.n2651 gnd.n2650 0.152939
R18935 gnd.n2650 gnd.n2041 0.152939
R18936 gnd.n2646 gnd.n2041 0.152939
R18937 gnd.n2646 gnd.n2645 0.152939
R18938 gnd.n2645 gnd.n2048 0.152939
R18939 gnd.n2641 gnd.n2048 0.152939
R18940 gnd.n2641 gnd.n2640 0.152939
R18941 gnd.n2450 gnd.n2251 0.152939
R18942 gnd.n2450 gnd.n2449 0.152939
R18943 gnd.n2449 gnd.n2448 0.152939
R18944 gnd.n2448 gnd.n2240 0.152939
R18945 gnd.n2505 gnd.n2240 0.152939
R18946 gnd.n2506 gnd.n2505 0.152939
R18947 gnd.n2507 gnd.n2506 0.152939
R18948 gnd.n2507 gnd.n2233 0.152939
R18949 gnd.n2521 gnd.n2233 0.152939
R18950 gnd.n2522 gnd.n2521 0.152939
R18951 gnd.n2523 gnd.n2522 0.152939
R18952 gnd.n2523 gnd.n2224 0.152939
R18953 gnd.n2551 gnd.n2224 0.152939
R18954 gnd.n2551 gnd.n2550 0.152939
R18955 gnd.n2550 gnd.n2549 0.152939
R18956 gnd.n2549 gnd.n2225 0.152939
R18957 gnd.n2545 gnd.n2225 0.152939
R18958 gnd.n2545 gnd.n2033 0.152939
R18959 gnd.n2659 gnd.n2033 0.152939
R18960 gnd.n2659 gnd.n2658 0.152939
R18961 gnd.n4271 gnd.n1087 0.152939
R18962 gnd.n4267 gnd.n1087 0.152939
R18963 gnd.n4267 gnd.n4266 0.152939
R18964 gnd.n4266 gnd.n4265 0.152939
R18965 gnd.n4265 gnd.n1092 0.152939
R18966 gnd.n4261 gnd.n1092 0.152939
R18967 gnd.n4261 gnd.n4260 0.152939
R18968 gnd.n4260 gnd.n4259 0.152939
R18969 gnd.n4259 gnd.n1097 0.152939
R18970 gnd.n4255 gnd.n1097 0.152939
R18971 gnd.n4255 gnd.n4254 0.152939
R18972 gnd.n4254 gnd.n4253 0.152939
R18973 gnd.n4253 gnd.n1102 0.152939
R18974 gnd.n4249 gnd.n1102 0.152939
R18975 gnd.n4249 gnd.n4248 0.152939
R18976 gnd.n4248 gnd.n4247 0.152939
R18977 gnd.n4247 gnd.n1107 0.152939
R18978 gnd.n4243 gnd.n1107 0.152939
R18979 gnd.n4243 gnd.n4242 0.152939
R18980 gnd.n4242 gnd.n4241 0.152939
R18981 gnd.n4241 gnd.n1112 0.152939
R18982 gnd.n4237 gnd.n1112 0.152939
R18983 gnd.n4237 gnd.n4236 0.152939
R18984 gnd.n4236 gnd.n4235 0.152939
R18985 gnd.n4235 gnd.n1117 0.152939
R18986 gnd.n4231 gnd.n1117 0.152939
R18987 gnd.n4231 gnd.n4230 0.152939
R18988 gnd.n4230 gnd.n4229 0.152939
R18989 gnd.n4229 gnd.n1122 0.152939
R18990 gnd.n4225 gnd.n1122 0.152939
R18991 gnd.n4225 gnd.n4224 0.152939
R18992 gnd.n4224 gnd.n4223 0.152939
R18993 gnd.n4223 gnd.n1127 0.152939
R18994 gnd.n4219 gnd.n1127 0.152939
R18995 gnd.n4219 gnd.n4218 0.152939
R18996 gnd.n4218 gnd.n4217 0.152939
R18997 gnd.n4217 gnd.n1132 0.152939
R18998 gnd.n4213 gnd.n1132 0.152939
R18999 gnd.n4213 gnd.n4212 0.152939
R19000 gnd.n4212 gnd.n4211 0.152939
R19001 gnd.n4211 gnd.n1137 0.152939
R19002 gnd.n4207 gnd.n1137 0.152939
R19003 gnd.n4207 gnd.n4206 0.152939
R19004 gnd.n4206 gnd.n4205 0.152939
R19005 gnd.n4205 gnd.n1142 0.152939
R19006 gnd.n4201 gnd.n1142 0.152939
R19007 gnd.n4201 gnd.n4200 0.152939
R19008 gnd.n4200 gnd.n4199 0.152939
R19009 gnd.n4199 gnd.n1147 0.152939
R19010 gnd.n4195 gnd.n1147 0.152939
R19011 gnd.n4195 gnd.n4194 0.152939
R19012 gnd.n4194 gnd.n4193 0.152939
R19013 gnd.n4193 gnd.n1152 0.152939
R19014 gnd.n4189 gnd.n1152 0.152939
R19015 gnd.n4189 gnd.n4188 0.152939
R19016 gnd.n4188 gnd.n4187 0.152939
R19017 gnd.n4187 gnd.n1157 0.152939
R19018 gnd.n4183 gnd.n1157 0.152939
R19019 gnd.n4183 gnd.n4182 0.152939
R19020 gnd.n4182 gnd.n4181 0.152939
R19021 gnd.n4181 gnd.n1162 0.152939
R19022 gnd.n4177 gnd.n1162 0.152939
R19023 gnd.n4177 gnd.n4176 0.152939
R19024 gnd.n4176 gnd.n4175 0.152939
R19025 gnd.n4175 gnd.n1167 0.152939
R19026 gnd.n4171 gnd.n1167 0.152939
R19027 gnd.n4171 gnd.n4170 0.152939
R19028 gnd.n4170 gnd.n4169 0.152939
R19029 gnd.n4169 gnd.n1172 0.152939
R19030 gnd.n4165 gnd.n1172 0.152939
R19031 gnd.n4165 gnd.n4164 0.152939
R19032 gnd.n4164 gnd.n4163 0.152939
R19033 gnd.n4163 gnd.n1177 0.152939
R19034 gnd.n4159 gnd.n1177 0.152939
R19035 gnd.n4159 gnd.n4158 0.152939
R19036 gnd.n4158 gnd.n4157 0.152939
R19037 gnd.n4157 gnd.n1182 0.152939
R19038 gnd.n4153 gnd.n1182 0.152939
R19039 gnd.n4153 gnd.n4152 0.152939
R19040 gnd.n4152 gnd.n4151 0.152939
R19041 gnd.n4151 gnd.n1187 0.152939
R19042 gnd.n1190 gnd.n1187 0.152939
R19043 gnd.n3468 gnd.n1232 0.152939
R19044 gnd.n4121 gnd.n1232 0.152939
R19045 gnd.n4121 gnd.n4120 0.152939
R19046 gnd.n4120 gnd.n4119 0.152939
R19047 gnd.n4119 gnd.n1233 0.152939
R19048 gnd.n4115 gnd.n1233 0.152939
R19049 gnd.n4115 gnd.n4114 0.152939
R19050 gnd.n4114 gnd.n4113 0.152939
R19051 gnd.n4113 gnd.n1238 0.152939
R19052 gnd.n4109 gnd.n1238 0.152939
R19053 gnd.n4109 gnd.n4108 0.152939
R19054 gnd.n4108 gnd.n4107 0.152939
R19055 gnd.n4107 gnd.n1243 0.152939
R19056 gnd.n4103 gnd.n1243 0.152939
R19057 gnd.n4103 gnd.n4102 0.152939
R19058 gnd.n4102 gnd.n4101 0.152939
R19059 gnd.n4101 gnd.n1248 0.152939
R19060 gnd.n4097 gnd.n1248 0.152939
R19061 gnd.n4097 gnd.n241 0.152939
R19062 gnd.n6652 gnd.n241 0.152939
R19063 gnd.n6653 gnd.n6652 0.152939
R19064 gnd.n6654 gnd.n6653 0.152939
R19065 gnd.n6654 gnd.n227 0.152939
R19066 gnd.n6666 gnd.n227 0.152939
R19067 gnd.n6667 gnd.n6666 0.152939
R19068 gnd.n6668 gnd.n6667 0.152939
R19069 gnd.n6668 gnd.n206 0.152939
R19070 gnd.n6682 gnd.n206 0.152939
R19071 gnd.n6683 gnd.n6682 0.152939
R19072 gnd.n6684 gnd.n6683 0.152939
R19073 gnd.n6684 gnd.n191 0.152939
R19074 gnd.n6698 gnd.n191 0.152939
R19075 gnd.n6699 gnd.n6698 0.152939
R19076 gnd.n6700 gnd.n6699 0.152939
R19077 gnd.n6700 gnd.n176 0.152939
R19078 gnd.n6714 gnd.n176 0.152939
R19079 gnd.n6715 gnd.n6714 0.152939
R19080 gnd.n6790 gnd.n6715 0.152939
R19081 gnd.n6790 gnd.n6789 0.152939
R19082 gnd.n6789 gnd.n6788 0.152939
R19083 gnd.n6788 gnd.n6716 0.152939
R19084 gnd.n6784 gnd.n6716 0.152939
R19085 gnd.n6783 gnd.n6718 0.152939
R19086 gnd.n6779 gnd.n6718 0.152939
R19087 gnd.n6779 gnd.n6778 0.152939
R19088 gnd.n6778 gnd.n6777 0.152939
R19089 gnd.n6777 gnd.n6724 0.152939
R19090 gnd.n6773 gnd.n6724 0.152939
R19091 gnd.n6773 gnd.n6772 0.152939
R19092 gnd.n6772 gnd.n6771 0.152939
R19093 gnd.n6771 gnd.n6732 0.152939
R19094 gnd.n6767 gnd.n6732 0.152939
R19095 gnd.n6767 gnd.n6766 0.152939
R19096 gnd.n6766 gnd.n6765 0.152939
R19097 gnd.n6765 gnd.n6740 0.152939
R19098 gnd.n6761 gnd.n6740 0.152939
R19099 gnd.n6761 gnd.n6760 0.152939
R19100 gnd.n6760 gnd.n6759 0.152939
R19101 gnd.n6759 gnd.n6748 0.152939
R19102 gnd.n6748 gnd.n78 0.152939
R19103 gnd.n3893 gnd.n1333 0.152939
R19104 gnd.n3894 gnd.n3893 0.152939
R19105 gnd.n3896 gnd.n3894 0.152939
R19106 gnd.n3896 gnd.n3895 0.152939
R19107 gnd.n3895 gnd.n1315 0.152939
R19108 gnd.n4023 gnd.n1315 0.152939
R19109 gnd.n4024 gnd.n4023 0.152939
R19110 gnd.n4026 gnd.n4024 0.152939
R19111 gnd.n4026 gnd.n4025 0.152939
R19112 gnd.n4025 gnd.n1286 0.152939
R19113 gnd.n4055 gnd.n1286 0.152939
R19114 gnd.n4056 gnd.n4055 0.152939
R19115 gnd.n4058 gnd.n4056 0.152939
R19116 gnd.n4058 gnd.n4057 0.152939
R19117 gnd.n4057 gnd.n1257 0.152939
R19118 gnd.n4089 gnd.n1257 0.152939
R19119 gnd.n4090 gnd.n4089 0.152939
R19120 gnd.n4092 gnd.n4090 0.152939
R19121 gnd.n4092 gnd.n4091 0.152939
R19122 gnd.n4091 gnd.n51 0.152939
R19123 gnd.n6915 gnd.n51 0.152939
R19124 gnd.n6915 gnd.n6914 0.152939
R19125 gnd.n6914 gnd.n53 0.152939
R19126 gnd.n6910 gnd.n53 0.152939
R19127 gnd.n6910 gnd.n6909 0.152939
R19128 gnd.n6909 gnd.n6908 0.152939
R19129 gnd.n6908 gnd.n58 0.152939
R19130 gnd.n6904 gnd.n58 0.152939
R19131 gnd.n6904 gnd.n6903 0.152939
R19132 gnd.n6903 gnd.n6902 0.152939
R19133 gnd.n6902 gnd.n63 0.152939
R19134 gnd.n6898 gnd.n63 0.152939
R19135 gnd.n6898 gnd.n6897 0.152939
R19136 gnd.n6897 gnd.n6896 0.152939
R19137 gnd.n6896 gnd.n68 0.152939
R19138 gnd.n6892 gnd.n68 0.152939
R19139 gnd.n6892 gnd.n6891 0.152939
R19140 gnd.n6891 gnd.n6890 0.152939
R19141 gnd.n6890 gnd.n73 0.152939
R19142 gnd.n6886 gnd.n73 0.152939
R19143 gnd.n6886 gnd.n6885 0.152939
R19144 gnd.n6885 gnd.n6884 0.152939
R19145 gnd.n3556 gnd.n3421 0.151415
R19146 gnd.n2657 gnd.n2034 0.151415
R19147 gnd.n2428 gnd.n2427 0.145814
R19148 gnd.n2428 gnd.n2251 0.145814
R19149 gnd.n5099 gnd.n0 0.127478
R19150 gnd.n254 gnd.n213 0.108732
R19151 gnd.n2469 gnd.n2468 0.108732
R19152 gnd.n5100 gnd.n4669 0.0767195
R19153 gnd.n5100 gnd.n5048 0.0767195
R19154 gnd.n4273 gnd.n4272 0.063
R19155 gnd.n3469 gnd.n3466 0.063
R19156 gnd.n5839 gnd.n4518 0.0477147
R19157 gnd.n255 gnd.n213 0.0447073
R19158 gnd.n2468 gnd.n2467 0.0447073
R19159 gnd.n5003 gnd.n4891 0.0442063
R19160 gnd.n5004 gnd.n5003 0.0442063
R19161 gnd.n5005 gnd.n5004 0.0442063
R19162 gnd.n5005 gnd.n4880 0.0442063
R19163 gnd.n5019 gnd.n4880 0.0442063
R19164 gnd.n5020 gnd.n5019 0.0442063
R19165 gnd.n5021 gnd.n5020 0.0442063
R19166 gnd.n5021 gnd.n4867 0.0442063
R19167 gnd.n5139 gnd.n4867 0.0442063
R19168 gnd.n5140 gnd.n5139 0.0442063
R19169 gnd.n5142 gnd.n4801 0.0344674
R19170 gnd.n3557 gnd.n3555 0.0344674
R19171 gnd.n2656 gnd.n2035 0.0344674
R19172 gnd.n5162 gnd.n5161 0.0269946
R19173 gnd.n5164 gnd.n5163 0.0269946
R19174 gnd.n4796 gnd.n4794 0.0269946
R19175 gnd.n5174 gnd.n5172 0.0269946
R19176 gnd.n5173 gnd.n4775 0.0269946
R19177 gnd.n5193 gnd.n5192 0.0269946
R19178 gnd.n5195 gnd.n5194 0.0269946
R19179 gnd.n4770 gnd.n4768 0.0269946
R19180 gnd.n5205 gnd.n5203 0.0269946
R19181 gnd.n5204 gnd.n4751 0.0269946
R19182 gnd.n5224 gnd.n5223 0.0269946
R19183 gnd.n5226 gnd.n5225 0.0269946
R19184 gnd.n4745 gnd.n4743 0.0269946
R19185 gnd.n5236 gnd.n5234 0.0269946
R19186 gnd.n5235 gnd.n4725 0.0269946
R19187 gnd.n5255 gnd.n5254 0.0269946
R19188 gnd.n5257 gnd.n5256 0.0269946
R19189 gnd.n4719 gnd.n4717 0.0269946
R19190 gnd.n5267 gnd.n5265 0.0269946
R19191 gnd.n5266 gnd.n4700 0.0269946
R19192 gnd.n5286 gnd.n5285 0.0269946
R19193 gnd.n5288 gnd.n5287 0.0269946
R19194 gnd.n4694 gnd.n4692 0.0269946
R19195 gnd.n5298 gnd.n5296 0.0269946
R19196 gnd.n5297 gnd.n4676 0.0269946
R19197 gnd.n5316 gnd.n5315 0.0269946
R19198 gnd.n5318 gnd.n5317 0.0269946
R19199 gnd.n4664 gnd.n4663 0.0269946
R19200 gnd.n5352 gnd.n4660 0.0269946
R19201 gnd.n5351 gnd.n4661 0.0269946
R19202 gnd.n5371 gnd.n4643 0.0269946
R19203 gnd.n5373 gnd.n5372 0.0269946
R19204 gnd.n5374 gnd.n4641 0.0269946
R19205 gnd.n5381 gnd.n5377 0.0269946
R19206 gnd.n5380 gnd.n5379 0.0269946
R19207 gnd.n5378 gnd.n4620 0.0269946
R19208 gnd.n5405 gnd.n4621 0.0269946
R19209 gnd.n5404 gnd.n4622 0.0269946
R19210 gnd.n5446 gnd.n4599 0.0269946
R19211 gnd.n5448 gnd.n5447 0.0269946
R19212 gnd.n5457 gnd.n4592 0.0269946
R19213 gnd.n5459 gnd.n5458 0.0269946
R19214 gnd.n5460 gnd.n4588 0.0269946
R19215 gnd.n5748 gnd.n4589 0.0269946
R19216 gnd.n5747 gnd.n4590 0.0269946
R19217 gnd.n5464 gnd.n771 0.0269946
R19218 gnd.n5465 gnd.n772 0.0269946
R19219 gnd.n5467 gnd.n773 0.0269946
R19220 gnd.n5727 gnd.n5726 0.0269946
R19221 gnd.n5728 gnd.n795 0.0269946
R19222 gnd.n5729 gnd.n796 0.0269946
R19223 gnd.n5730 gnd.n797 0.0269946
R19224 gnd.n3466 gnd.n3465 0.0246168
R19225 gnd.n4272 gnd.n1086 0.0246168
R19226 gnd.n5142 gnd.n5141 0.0202011
R19227 gnd.n3465 gnd.n3463 0.0174837
R19228 gnd.n3477 gnd.n3463 0.0174837
R19229 gnd.n3479 gnd.n3477 0.0174837
R19230 gnd.n3479 gnd.n3478 0.0174837
R19231 gnd.n3478 gnd.n3458 0.0174837
R19232 gnd.n3488 gnd.n3458 0.0174837
R19233 gnd.n3488 gnd.n3487 0.0174837
R19234 gnd.n3487 gnd.n3459 0.0174837
R19235 gnd.n3459 gnd.n3454 0.0174837
R19236 gnd.n3496 gnd.n3454 0.0174837
R19237 gnd.n3498 gnd.n3496 0.0174837
R19238 gnd.n3498 gnd.n3497 0.0174837
R19239 gnd.n3497 gnd.n3449 0.0174837
R19240 gnd.n3507 gnd.n3449 0.0174837
R19241 gnd.n3507 gnd.n3506 0.0174837
R19242 gnd.n3506 gnd.n3450 0.0174837
R19243 gnd.n3450 gnd.n3445 0.0174837
R19244 gnd.n3515 gnd.n3445 0.0174837
R19245 gnd.n3517 gnd.n3515 0.0174837
R19246 gnd.n3517 gnd.n3516 0.0174837
R19247 gnd.n3516 gnd.n3440 0.0174837
R19248 gnd.n3526 gnd.n3440 0.0174837
R19249 gnd.n3526 gnd.n3525 0.0174837
R19250 gnd.n3525 gnd.n3441 0.0174837
R19251 gnd.n3441 gnd.n3436 0.0174837
R19252 gnd.n3534 gnd.n3436 0.0174837
R19253 gnd.n3536 gnd.n3534 0.0174837
R19254 gnd.n3536 gnd.n3535 0.0174837
R19255 gnd.n3535 gnd.n3431 0.0174837
R19256 gnd.n3547 gnd.n3431 0.0174837
R19257 gnd.n3547 gnd.n3546 0.0174837
R19258 gnd.n3546 gnd.n3432 0.0174837
R19259 gnd.n3432 gnd.n3425 0.0174837
R19260 gnd.n3554 gnd.n3425 0.0174837
R19261 gnd.n3555 gnd.n3554 0.0174837
R19262 gnd.n2091 gnd.n1086 0.0174837
R19263 gnd.n2093 gnd.n2091 0.0174837
R19264 gnd.n2201 gnd.n2093 0.0174837
R19265 gnd.n2201 gnd.n2200 0.0174837
R19266 gnd.n2200 gnd.n2094 0.0174837
R19267 gnd.n2197 gnd.n2094 0.0174837
R19268 gnd.n2197 gnd.n2196 0.0174837
R19269 gnd.n2196 gnd.n2104 0.0174837
R19270 gnd.n2193 gnd.n2104 0.0174837
R19271 gnd.n2193 gnd.n2192 0.0174837
R19272 gnd.n2192 gnd.n2109 0.0174837
R19273 gnd.n2189 gnd.n2109 0.0174837
R19274 gnd.n2189 gnd.n2188 0.0174837
R19275 gnd.n2188 gnd.n2115 0.0174837
R19276 gnd.n2185 gnd.n2115 0.0174837
R19277 gnd.n2185 gnd.n2184 0.0174837
R19278 gnd.n2184 gnd.n2119 0.0174837
R19279 gnd.n2181 gnd.n2119 0.0174837
R19280 gnd.n2181 gnd.n2180 0.0174837
R19281 gnd.n2180 gnd.n2126 0.0174837
R19282 gnd.n2177 gnd.n2126 0.0174837
R19283 gnd.n2177 gnd.n2176 0.0174837
R19284 gnd.n2176 gnd.n2132 0.0174837
R19285 gnd.n2173 gnd.n2132 0.0174837
R19286 gnd.n2173 gnd.n2172 0.0174837
R19287 gnd.n2172 gnd.n2138 0.0174837
R19288 gnd.n2169 gnd.n2138 0.0174837
R19289 gnd.n2169 gnd.n2168 0.0174837
R19290 gnd.n2168 gnd.n2142 0.0174837
R19291 gnd.n2165 gnd.n2142 0.0174837
R19292 gnd.n2165 gnd.n2164 0.0174837
R19293 gnd.n2164 gnd.n2151 0.0174837
R19294 gnd.n2161 gnd.n2151 0.0174837
R19295 gnd.n2161 gnd.n2160 0.0174837
R19296 gnd.n2160 gnd.n2035 0.0174837
R19297 gnd.n5141 gnd.n5140 0.0148637
R19298 gnd.n5724 gnd.n5468 0.0144266
R19299 gnd.n5725 gnd.n5724 0.0130679
R19300 gnd.n5161 gnd.n4801 0.00797283
R19301 gnd.n5163 gnd.n5162 0.00797283
R19302 gnd.n5164 gnd.n4796 0.00797283
R19303 gnd.n5172 gnd.n4794 0.00797283
R19304 gnd.n5174 gnd.n5173 0.00797283
R19305 gnd.n5192 gnd.n4775 0.00797283
R19306 gnd.n5194 gnd.n5193 0.00797283
R19307 gnd.n5195 gnd.n4770 0.00797283
R19308 gnd.n5203 gnd.n4768 0.00797283
R19309 gnd.n5205 gnd.n5204 0.00797283
R19310 gnd.n5223 gnd.n4751 0.00797283
R19311 gnd.n5225 gnd.n5224 0.00797283
R19312 gnd.n5226 gnd.n4745 0.00797283
R19313 gnd.n5234 gnd.n4743 0.00797283
R19314 gnd.n5236 gnd.n5235 0.00797283
R19315 gnd.n5254 gnd.n4725 0.00797283
R19316 gnd.n5256 gnd.n5255 0.00797283
R19317 gnd.n5257 gnd.n4719 0.00797283
R19318 gnd.n5265 gnd.n4717 0.00797283
R19319 gnd.n5267 gnd.n5266 0.00797283
R19320 gnd.n5285 gnd.n4700 0.00797283
R19321 gnd.n5287 gnd.n5286 0.00797283
R19322 gnd.n5288 gnd.n4694 0.00797283
R19323 gnd.n5296 gnd.n4692 0.00797283
R19324 gnd.n5298 gnd.n5297 0.00797283
R19325 gnd.n5315 gnd.n4676 0.00797283
R19326 gnd.n5317 gnd.n5316 0.00797283
R19327 gnd.n5318 gnd.n4664 0.00797283
R19328 gnd.n4663 gnd.n4660 0.00797283
R19329 gnd.n5352 gnd.n5351 0.00797283
R19330 gnd.n4661 gnd.n4643 0.00797283
R19331 gnd.n5372 gnd.n5371 0.00797283
R19332 gnd.n5374 gnd.n5373 0.00797283
R19333 gnd.n5377 gnd.n4641 0.00797283
R19334 gnd.n5381 gnd.n5380 0.00797283
R19335 gnd.n5379 gnd.n5378 0.00797283
R19336 gnd.n4621 gnd.n4620 0.00797283
R19337 gnd.n5405 gnd.n5404 0.00797283
R19338 gnd.n4622 gnd.n4599 0.00797283
R19339 gnd.n5448 gnd.n5446 0.00797283
R19340 gnd.n5447 gnd.n4592 0.00797283
R19341 gnd.n5458 gnd.n5457 0.00797283
R19342 gnd.n5460 gnd.n5459 0.00797283
R19343 gnd.n4589 gnd.n4588 0.00797283
R19344 gnd.n5748 gnd.n5747 0.00797283
R19345 gnd.n5464 gnd.n4590 0.00797283
R19346 gnd.n5465 gnd.n771 0.00797283
R19347 gnd.n5467 gnd.n772 0.00797283
R19348 gnd.n5468 gnd.n773 0.00797283
R19349 gnd.n5726 gnd.n5725 0.00797283
R19350 gnd.n5728 gnd.n5727 0.00797283
R19351 gnd.n5729 gnd.n795 0.00797283
R19352 gnd.n5730 gnd.n796 0.00797283
R19353 gnd.n4518 gnd.n797 0.00797283
R19354 gnd.n6653 gnd.n240 0.00614909
R19355 gnd.n2256 gnd.n2255 0.00614909
R19356 gnd.n3557 gnd.n3556 0.000839674
R19357 gnd.n2657 gnd.n2656 0.000839674
R19358 plus.n53 plus.t20 323.478
R19359 plus.n11 plus.t15 323.478
R19360 plus.n52 plus.t19 297.12
R19361 plus.n56 plus.t26 297.12
R19362 plus.n58 plus.t25 297.12
R19363 plus.n62 plus.t27 297.12
R19364 plus.n64 plus.t9 297.12
R19365 plus.n68 plus.t7 297.12
R19366 plus.n70 plus.t14 297.12
R19367 plus.n74 plus.t12 297.12
R19368 plus.n76 plus.t28 297.12
R19369 plus.n80 plus.t10 297.12
R19370 plus.n82 plus.t8 297.12
R19371 plus.n40 plus.t21 297.12
R19372 plus.n38 plus.t22 297.12
R19373 plus.n2 plus.t16 297.12
R19374 plus.n32 plus.t17 297.12
R19375 plus.n4 plus.t11 297.12
R19376 plus.n26 plus.t5 297.12
R19377 plus.n6 plus.t6 297.12
R19378 plus.n20 plus.t23 297.12
R19379 plus.n8 plus.t24 297.12
R19380 plus.n14 plus.t18 297.12
R19381 plus.n10 plus.t13 297.12
R19382 plus.n86 plus.t2 243.97
R19383 plus.n86 plus.n85 223.454
R19384 plus.n88 plus.n87 223.454
R19385 plus.n83 plus.n82 161.3
R19386 plus.n81 plus.n42 161.3
R19387 plus.n80 plus.n79 161.3
R19388 plus.n78 plus.n43 161.3
R19389 plus.n77 plus.n76 161.3
R19390 plus.n75 plus.n44 161.3
R19391 plus.n74 plus.n73 161.3
R19392 plus.n72 plus.n45 161.3
R19393 plus.n71 plus.n70 161.3
R19394 plus.n69 plus.n46 161.3
R19395 plus.n68 plus.n67 161.3
R19396 plus.n66 plus.n47 161.3
R19397 plus.n65 plus.n64 161.3
R19398 plus.n63 plus.n48 161.3
R19399 plus.n62 plus.n61 161.3
R19400 plus.n60 plus.n49 161.3
R19401 plus.n59 plus.n58 161.3
R19402 plus.n57 plus.n50 161.3
R19403 plus.n56 plus.n55 161.3
R19404 plus.n54 plus.n51 161.3
R19405 plus.n13 plus.n12 161.3
R19406 plus.n14 plus.n9 161.3
R19407 plus.n16 plus.n15 161.3
R19408 plus.n17 plus.n8 161.3
R19409 plus.n19 plus.n18 161.3
R19410 plus.n20 plus.n7 161.3
R19411 plus.n22 plus.n21 161.3
R19412 plus.n23 plus.n6 161.3
R19413 plus.n25 plus.n24 161.3
R19414 plus.n26 plus.n5 161.3
R19415 plus.n28 plus.n27 161.3
R19416 plus.n29 plus.n4 161.3
R19417 plus.n31 plus.n30 161.3
R19418 plus.n32 plus.n3 161.3
R19419 plus.n34 plus.n33 161.3
R19420 plus.n35 plus.n2 161.3
R19421 plus.n37 plus.n36 161.3
R19422 plus.n38 plus.n1 161.3
R19423 plus.n39 plus.n0 161.3
R19424 plus.n41 plus.n40 161.3
R19425 plus.n82 plus.n81 46.0096
R19426 plus.n40 plus.n39 46.0096
R19427 plus.n54 plus.n53 45.0871
R19428 plus.n12 plus.n11 45.0871
R19429 plus.n52 plus.n51 41.6278
R19430 plus.n80 plus.n43 41.6278
R19431 plus.n38 plus.n37 41.6278
R19432 plus.n13 plus.n10 41.6278
R19433 plus.n57 plus.n56 37.246
R19434 plus.n76 plus.n75 37.246
R19435 plus.n33 plus.n2 37.246
R19436 plus.n15 plus.n14 37.246
R19437 plus.n84 plus.n83 33.1766
R19438 plus.n58 plus.n49 32.8641
R19439 plus.n74 plus.n45 32.8641
R19440 plus.n32 plus.n31 32.8641
R19441 plus.n19 plus.n8 32.8641
R19442 plus.n63 plus.n62 28.4823
R19443 plus.n70 plus.n69 28.4823
R19444 plus.n27 plus.n4 28.4823
R19445 plus.n21 plus.n20 28.4823
R19446 plus.n64 plus.n47 24.1005
R19447 plus.n68 plus.n47 24.1005
R19448 plus.n26 plus.n25 24.1005
R19449 plus.n25 plus.n6 24.1005
R19450 plus.n85 plus.t3 19.8005
R19451 plus.n85 plus.t1 19.8005
R19452 plus.n87 plus.t4 19.8005
R19453 plus.n87 plus.t0 19.8005
R19454 plus.n64 plus.n63 19.7187
R19455 plus.n69 plus.n68 19.7187
R19456 plus.n27 plus.n26 19.7187
R19457 plus.n21 plus.n6 19.7187
R19458 plus.n62 plus.n49 15.3369
R19459 plus.n70 plus.n45 15.3369
R19460 plus.n31 plus.n4 15.3369
R19461 plus.n20 plus.n19 15.3369
R19462 plus plus.n89 14.2409
R19463 plus.n53 plus.n52 14.1472
R19464 plus.n11 plus.n10 14.1472
R19465 plus.n84 plus.n41 11.8774
R19466 plus.n58 plus.n57 10.955
R19467 plus.n75 plus.n74 10.955
R19468 plus.n33 plus.n32 10.955
R19469 plus.n15 plus.n8 10.955
R19470 plus.n56 plus.n51 6.57323
R19471 plus.n76 plus.n43 6.57323
R19472 plus.n37 plus.n2 6.57323
R19473 plus.n14 plus.n13 6.57323
R19474 plus.n89 plus.n88 5.40567
R19475 plus.n81 plus.n80 2.19141
R19476 plus.n39 plus.n38 2.19141
R19477 plus.n89 plus.n84 1.188
R19478 plus.n88 plus.n86 0.716017
R19479 plus.n55 plus.n54 0.189894
R19480 plus.n55 plus.n50 0.189894
R19481 plus.n59 plus.n50 0.189894
R19482 plus.n60 plus.n59 0.189894
R19483 plus.n61 plus.n60 0.189894
R19484 plus.n61 plus.n48 0.189894
R19485 plus.n65 plus.n48 0.189894
R19486 plus.n66 plus.n65 0.189894
R19487 plus.n67 plus.n66 0.189894
R19488 plus.n67 plus.n46 0.189894
R19489 plus.n71 plus.n46 0.189894
R19490 plus.n72 plus.n71 0.189894
R19491 plus.n73 plus.n72 0.189894
R19492 plus.n73 plus.n44 0.189894
R19493 plus.n77 plus.n44 0.189894
R19494 plus.n78 plus.n77 0.189894
R19495 plus.n79 plus.n78 0.189894
R19496 plus.n79 plus.n42 0.189894
R19497 plus.n83 plus.n42 0.189894
R19498 plus.n41 plus.n0 0.189894
R19499 plus.n1 plus.n0 0.189894
R19500 plus.n36 plus.n1 0.189894
R19501 plus.n36 plus.n35 0.189894
R19502 plus.n35 plus.n34 0.189894
R19503 plus.n34 plus.n3 0.189894
R19504 plus.n30 plus.n3 0.189894
R19505 plus.n30 plus.n29 0.189894
R19506 plus.n29 plus.n28 0.189894
R19507 plus.n28 plus.n5 0.189894
R19508 plus.n24 plus.n5 0.189894
R19509 plus.n24 plus.n23 0.189894
R19510 plus.n23 plus.n22 0.189894
R19511 plus.n22 plus.n7 0.189894
R19512 plus.n18 plus.n7 0.189894
R19513 plus.n18 plus.n17 0.189894
R19514 plus.n17 plus.n16 0.189894
R19515 plus.n16 plus.n9 0.189894
R19516 plus.n12 plus.n9 0.189894
R19517 a_n2903_n3924.n30 a_n2903_n3924.t37 214.643
R19518 a_n2903_n3924.n37 a_n2903_n3924.t32 214.321
R19519 a_n2903_n3924.n36 a_n2903_n3924.t34 214.321
R19520 a_n2903_n3924.n35 a_n2903_n3924.t39 214.321
R19521 a_n2903_n3924.n34 a_n2903_n3924.t36 214.321
R19522 a_n2903_n3924.n33 a_n2903_n3924.t41 214.321
R19523 a_n2903_n3924.n32 a_n2903_n3924.t33 214.321
R19524 a_n2903_n3924.n31 a_n2903_n3924.t55 214.321
R19525 a_n2903_n3924.n13 a_n2903_n3924.t15 55.8337
R19526 a_n2903_n3924.n14 a_n2903_n3924.t49 55.8337
R19527 a_n2903_n3924.n25 a_n2903_n3924.t40 55.8337
R19528 a_n2903_n3924.n2 a_n2903_n3924.t27 55.8335
R19529 a_n2903_n3924.n39 a_n2903_n3924.t2 55.8335
R19530 a_n2903_n3924.n50 a_n2903_n3924.t52 55.8335
R19531 a_n2903_n3924.n51 a_n2903_n3924.t20 55.8335
R19532 a_n2903_n3924.n28 a_n2903_n3924.t14 55.8335
R19533 a_n2903_n3924.n57 a_n2903_n3924.n56 53.0054
R19534 a_n2903_n3924.n4 a_n2903_n3924.n3 53.0052
R19535 a_n2903_n3924.n6 a_n2903_n3924.n5 53.0052
R19536 a_n2903_n3924.n8 a_n2903_n3924.n7 53.0052
R19537 a_n2903_n3924.n10 a_n2903_n3924.n9 53.0052
R19538 a_n2903_n3924.n12 a_n2903_n3924.n11 53.0052
R19539 a_n2903_n3924.n16 a_n2903_n3924.n15 53.0052
R19540 a_n2903_n3924.n18 a_n2903_n3924.n17 53.0052
R19541 a_n2903_n3924.n20 a_n2903_n3924.n19 53.0052
R19542 a_n2903_n3924.n22 a_n2903_n3924.n21 53.0052
R19543 a_n2903_n3924.n24 a_n2903_n3924.n23 53.0052
R19544 a_n2903_n3924.n41 a_n2903_n3924.n40 53.0051
R19545 a_n2903_n3924.n43 a_n2903_n3924.n42 53.0051
R19546 a_n2903_n3924.n45 a_n2903_n3924.n44 53.0051
R19547 a_n2903_n3924.n47 a_n2903_n3924.n46 53.0051
R19548 a_n2903_n3924.n49 a_n2903_n3924.n48 53.0051
R19549 a_n2903_n3924.n53 a_n2903_n3924.n52 53.0051
R19550 a_n2903_n3924.n55 a_n2903_n3924.n54 53.0051
R19551 a_n2903_n3924.n1 a_n2903_n3924.n0 53.0051
R19552 a_n2903_n3924.n27 a_n2903_n3924.n26 53.0051
R19553 a_n2903_n3924.n29 a_n2903_n3924.n25 12.1986
R19554 a_n2903_n3924.n38 a_n2903_n3924.n2 12.1986
R19555 a_n2903_n3924.n29 a_n2903_n3924.n28 5.11903
R19556 a_n2903_n3924.n39 a_n2903_n3924.n38 5.11903
R19557 a_n2903_n3924.n40 a_n2903_n3924.t53 2.82907
R19558 a_n2903_n3924.n40 a_n2903_n3924.t48 2.82907
R19559 a_n2903_n3924.n42 a_n2903_n3924.t51 2.82907
R19560 a_n2903_n3924.n42 a_n2903_n3924.t44 2.82907
R19561 a_n2903_n3924.n44 a_n2903_n3924.t1 2.82907
R19562 a_n2903_n3924.n44 a_n2903_n3924.t38 2.82907
R19563 a_n2903_n3924.n46 a_n2903_n3924.t5 2.82907
R19564 a_n2903_n3924.n46 a_n2903_n3924.t4 2.82907
R19565 a_n2903_n3924.n48 a_n2903_n3924.t47 2.82907
R19566 a_n2903_n3924.n48 a_n2903_n3924.t6 2.82907
R19567 a_n2903_n3924.n52 a_n2903_n3924.t17 2.82907
R19568 a_n2903_n3924.n52 a_n2903_n3924.t22 2.82907
R19569 a_n2903_n3924.n54 a_n2903_n3924.t12 2.82907
R19570 a_n2903_n3924.n54 a_n2903_n3924.t11 2.82907
R19571 a_n2903_n3924.n0 a_n2903_n3924.t18 2.82907
R19572 a_n2903_n3924.n0 a_n2903_n3924.t24 2.82907
R19573 a_n2903_n3924.n26 a_n2903_n3924.t13 2.82907
R19574 a_n2903_n3924.n26 a_n2903_n3924.t19 2.82907
R19575 a_n2903_n3924.n3 a_n2903_n3924.t7 2.82907
R19576 a_n2903_n3924.n3 a_n2903_n3924.t25 2.82907
R19577 a_n2903_n3924.n5 a_n2903_n3924.t21 2.82907
R19578 a_n2903_n3924.n5 a_n2903_n3924.t23 2.82907
R19579 a_n2903_n3924.n7 a_n2903_n3924.t26 2.82907
R19580 a_n2903_n3924.n7 a_n2903_n3924.t28 2.82907
R19581 a_n2903_n3924.n9 a_n2903_n3924.t10 2.82907
R19582 a_n2903_n3924.n9 a_n2903_n3924.t8 2.82907
R19583 a_n2903_n3924.n11 a_n2903_n3924.t16 2.82907
R19584 a_n2903_n3924.n11 a_n2903_n3924.t9 2.82907
R19585 a_n2903_n3924.n15 a_n2903_n3924.t31 2.82907
R19586 a_n2903_n3924.n15 a_n2903_n3924.t50 2.82907
R19587 a_n2903_n3924.n17 a_n2903_n3924.t46 2.82907
R19588 a_n2903_n3924.n17 a_n2903_n3924.t3 2.82907
R19589 a_n2903_n3924.n19 a_n2903_n3924.t43 2.82907
R19590 a_n2903_n3924.n19 a_n2903_n3924.t42 2.82907
R19591 a_n2903_n3924.n21 a_n2903_n3924.t0 2.82907
R19592 a_n2903_n3924.n21 a_n2903_n3924.t54 2.82907
R19593 a_n2903_n3924.n23 a_n2903_n3924.t45 2.82907
R19594 a_n2903_n3924.n23 a_n2903_n3924.t35 2.82907
R19595 a_n2903_n3924.t30 a_n2903_n3924.n57 2.82907
R19596 a_n2903_n3924.n57 a_n2903_n3924.t29 2.82907
R19597 a_n2903_n3924.n38 a_n2903_n3924.n37 2.16406
R19598 a_n2903_n3924.n30 a_n2903_n3924.n29 1.95694
R19599 a_n2903_n3924.n32 a_n2903_n3924.n31 0.672012
R19600 a_n2903_n3924.n33 a_n2903_n3924.n32 0.672012
R19601 a_n2903_n3924.n34 a_n2903_n3924.n33 0.672012
R19602 a_n2903_n3924.n35 a_n2903_n3924.n34 0.672012
R19603 a_n2903_n3924.n36 a_n2903_n3924.n35 0.672012
R19604 a_n2903_n3924.n37 a_n2903_n3924.n36 0.672012
R19605 a_n2903_n3924.n25 a_n2903_n3924.n24 0.444466
R19606 a_n2903_n3924.n24 a_n2903_n3924.n22 0.444466
R19607 a_n2903_n3924.n22 a_n2903_n3924.n20 0.444466
R19608 a_n2903_n3924.n20 a_n2903_n3924.n18 0.444466
R19609 a_n2903_n3924.n18 a_n2903_n3924.n16 0.444466
R19610 a_n2903_n3924.n16 a_n2903_n3924.n14 0.444466
R19611 a_n2903_n3924.n13 a_n2903_n3924.n12 0.444466
R19612 a_n2903_n3924.n12 a_n2903_n3924.n10 0.444466
R19613 a_n2903_n3924.n10 a_n2903_n3924.n8 0.444466
R19614 a_n2903_n3924.n8 a_n2903_n3924.n6 0.444466
R19615 a_n2903_n3924.n6 a_n2903_n3924.n4 0.444466
R19616 a_n2903_n3924.n4 a_n2903_n3924.n2 0.444466
R19617 a_n2903_n3924.n28 a_n2903_n3924.n27 0.444466
R19618 a_n2903_n3924.n27 a_n2903_n3924.n1 0.444466
R19619 a_n2903_n3924.n56 a_n2903_n3924.n1 0.444466
R19620 a_n2903_n3924.n56 a_n2903_n3924.n55 0.444466
R19621 a_n2903_n3924.n55 a_n2903_n3924.n53 0.444466
R19622 a_n2903_n3924.n53 a_n2903_n3924.n51 0.444466
R19623 a_n2903_n3924.n50 a_n2903_n3924.n49 0.444466
R19624 a_n2903_n3924.n49 a_n2903_n3924.n47 0.444466
R19625 a_n2903_n3924.n47 a_n2903_n3924.n45 0.444466
R19626 a_n2903_n3924.n45 a_n2903_n3924.n43 0.444466
R19627 a_n2903_n3924.n43 a_n2903_n3924.n41 0.444466
R19628 a_n2903_n3924.n41 a_n2903_n3924.n39 0.444466
R19629 a_n2903_n3924.n31 a_n2903_n3924.n30 0.350064
R19630 a_n2903_n3924.n14 a_n2903_n3924.n13 0.235414
R19631 a_n2903_n3924.n51 a_n2903_n3924.n50 0.235414
R19632 commonsourceibias.n25 commonsourceibias.t46 230.006
R19633 commonsourceibias.n91 commonsourceibias.t62 230.006
R19634 commonsourceibias.n154 commonsourceibias.t54 230.006
R19635 commonsourceibias.n258 commonsourceibias.t16 230.006
R19636 commonsourceibias.n217 commonsourceibias.t75 230.006
R19637 commonsourceibias.n355 commonsourceibias.t65 230.006
R19638 commonsourceibias.n70 commonsourceibias.t32 207.983
R19639 commonsourceibias.n136 commonsourceibias.t71 207.983
R19640 commonsourceibias.n199 commonsourceibias.t61 207.983
R19641 commonsourceibias.n304 commonsourceibias.t2 207.983
R19642 commonsourceibias.n338 commonsourceibias.t84 207.983
R19643 commonsourceibias.n401 commonsourceibias.t73 207.983
R19644 commonsourceibias.n10 commonsourceibias.t14 168.701
R19645 commonsourceibias.n63 commonsourceibias.t24 168.701
R19646 commonsourceibias.n57 commonsourceibias.t30 168.701
R19647 commonsourceibias.n16 commonsourceibias.t20 168.701
R19648 commonsourceibias.n49 commonsourceibias.t36 168.701
R19649 commonsourceibias.n43 commonsourceibias.t44 168.701
R19650 commonsourceibias.n19 commonsourceibias.t26 168.701
R19651 commonsourceibias.n21 commonsourceibias.t34 168.701
R19652 commonsourceibias.n23 commonsourceibias.t10 168.701
R19653 commonsourceibias.n26 commonsourceibias.t40 168.701
R19654 commonsourceibias.n1 commonsourceibias.t81 168.701
R19655 commonsourceibias.n129 commonsourceibias.t55 168.701
R19656 commonsourceibias.n123 commonsourceibias.t53 168.701
R19657 commonsourceibias.n7 commonsourceibias.t76 168.701
R19658 commonsourceibias.n115 commonsourceibias.t86 168.701
R19659 commonsourceibias.n109 commonsourceibias.t50 168.701
R19660 commonsourceibias.n85 commonsourceibias.t69 168.701
R19661 commonsourceibias.n87 commonsourceibias.t67 168.701
R19662 commonsourceibias.n89 commonsourceibias.t78 168.701
R19663 commonsourceibias.n92 commonsourceibias.t64 168.701
R19664 commonsourceibias.n155 commonsourceibias.t57 168.701
R19665 commonsourceibias.n152 commonsourceibias.t68 168.701
R19666 commonsourceibias.n150 commonsourceibias.t58 168.701
R19667 commonsourceibias.n148 commonsourceibias.t60 168.701
R19668 commonsourceibias.n172 commonsourceibias.t91 168.701
R19669 commonsourceibias.n178 commonsourceibias.t77 168.701
R19670 commonsourceibias.n145 commonsourceibias.t66 168.701
R19671 commonsourceibias.n186 commonsourceibias.t95 168.701
R19672 commonsourceibias.n192 commonsourceibias.t49 168.701
R19673 commonsourceibias.n139 commonsourceibias.t72 168.701
R19674 commonsourceibias.n259 commonsourceibias.t8 168.701
R19675 commonsourceibias.n256 commonsourceibias.t18 168.701
R19676 commonsourceibias.n254 commonsourceibias.t4 168.701
R19677 commonsourceibias.n252 commonsourceibias.t42 168.701
R19678 commonsourceibias.n276 commonsourceibias.t12 168.701
R19679 commonsourceibias.n282 commonsourceibias.t6 168.701
R19680 commonsourceibias.n284 commonsourceibias.t28 168.701
R19681 commonsourceibias.n291 commonsourceibias.t0 168.701
R19682 commonsourceibias.n297 commonsourceibias.t38 168.701
R19683 commonsourceibias.n244 commonsourceibias.t22 168.701
R19684 commonsourceibias.n203 commonsourceibias.t92 168.701
R19685 commonsourceibias.n331 commonsourceibias.t51 168.701
R19686 commonsourceibias.n325 commonsourceibias.t63 168.701
R19687 commonsourceibias.n318 commonsourceibias.t88 168.701
R19688 commonsourceibias.n316 commonsourceibias.t48 168.701
R19689 commonsourceibias.n218 commonsourceibias.t59 168.701
R19690 commonsourceibias.n215 commonsourceibias.t90 168.701
R19691 commonsourceibias.n213 commonsourceibias.t80 168.701
R19692 commonsourceibias.n211 commonsourceibias.t83 168.701
R19693 commonsourceibias.n235 commonsourceibias.t94 168.701
R19694 commonsourceibias.n356 commonsourceibias.t52 168.701
R19695 commonsourceibias.n353 commonsourceibias.t82 168.701
R19696 commonsourceibias.n351 commonsourceibias.t70 168.701
R19697 commonsourceibias.n349 commonsourceibias.t74 168.701
R19698 commonsourceibias.n373 commonsourceibias.t87 168.701
R19699 commonsourceibias.n379 commonsourceibias.t89 168.701
R19700 commonsourceibias.n381 commonsourceibias.t79 168.701
R19701 commonsourceibias.n388 commonsourceibias.t56 168.701
R19702 commonsourceibias.n394 commonsourceibias.t93 168.701
R19703 commonsourceibias.n341 commonsourceibias.t85 168.701
R19704 commonsourceibias.n27 commonsourceibias.n24 161.3
R19705 commonsourceibias.n29 commonsourceibias.n28 161.3
R19706 commonsourceibias.n31 commonsourceibias.n30 161.3
R19707 commonsourceibias.n32 commonsourceibias.n22 161.3
R19708 commonsourceibias.n34 commonsourceibias.n33 161.3
R19709 commonsourceibias.n36 commonsourceibias.n35 161.3
R19710 commonsourceibias.n37 commonsourceibias.n20 161.3
R19711 commonsourceibias.n39 commonsourceibias.n38 161.3
R19712 commonsourceibias.n41 commonsourceibias.n40 161.3
R19713 commonsourceibias.n42 commonsourceibias.n18 161.3
R19714 commonsourceibias.n45 commonsourceibias.n44 161.3
R19715 commonsourceibias.n46 commonsourceibias.n17 161.3
R19716 commonsourceibias.n48 commonsourceibias.n47 161.3
R19717 commonsourceibias.n50 commonsourceibias.n15 161.3
R19718 commonsourceibias.n52 commonsourceibias.n51 161.3
R19719 commonsourceibias.n53 commonsourceibias.n14 161.3
R19720 commonsourceibias.n55 commonsourceibias.n54 161.3
R19721 commonsourceibias.n56 commonsourceibias.n13 161.3
R19722 commonsourceibias.n59 commonsourceibias.n58 161.3
R19723 commonsourceibias.n60 commonsourceibias.n12 161.3
R19724 commonsourceibias.n62 commonsourceibias.n61 161.3
R19725 commonsourceibias.n64 commonsourceibias.n11 161.3
R19726 commonsourceibias.n66 commonsourceibias.n65 161.3
R19727 commonsourceibias.n68 commonsourceibias.n67 161.3
R19728 commonsourceibias.n69 commonsourceibias.n9 161.3
R19729 commonsourceibias.n93 commonsourceibias.n90 161.3
R19730 commonsourceibias.n95 commonsourceibias.n94 161.3
R19731 commonsourceibias.n97 commonsourceibias.n96 161.3
R19732 commonsourceibias.n98 commonsourceibias.n88 161.3
R19733 commonsourceibias.n100 commonsourceibias.n99 161.3
R19734 commonsourceibias.n102 commonsourceibias.n101 161.3
R19735 commonsourceibias.n103 commonsourceibias.n86 161.3
R19736 commonsourceibias.n105 commonsourceibias.n104 161.3
R19737 commonsourceibias.n107 commonsourceibias.n106 161.3
R19738 commonsourceibias.n108 commonsourceibias.n84 161.3
R19739 commonsourceibias.n111 commonsourceibias.n110 161.3
R19740 commonsourceibias.n112 commonsourceibias.n8 161.3
R19741 commonsourceibias.n114 commonsourceibias.n113 161.3
R19742 commonsourceibias.n116 commonsourceibias.n6 161.3
R19743 commonsourceibias.n118 commonsourceibias.n117 161.3
R19744 commonsourceibias.n119 commonsourceibias.n5 161.3
R19745 commonsourceibias.n121 commonsourceibias.n120 161.3
R19746 commonsourceibias.n122 commonsourceibias.n4 161.3
R19747 commonsourceibias.n125 commonsourceibias.n124 161.3
R19748 commonsourceibias.n126 commonsourceibias.n3 161.3
R19749 commonsourceibias.n128 commonsourceibias.n127 161.3
R19750 commonsourceibias.n130 commonsourceibias.n2 161.3
R19751 commonsourceibias.n132 commonsourceibias.n131 161.3
R19752 commonsourceibias.n134 commonsourceibias.n133 161.3
R19753 commonsourceibias.n135 commonsourceibias.n0 161.3
R19754 commonsourceibias.n198 commonsourceibias.n138 161.3
R19755 commonsourceibias.n197 commonsourceibias.n196 161.3
R19756 commonsourceibias.n195 commonsourceibias.n194 161.3
R19757 commonsourceibias.n193 commonsourceibias.n140 161.3
R19758 commonsourceibias.n191 commonsourceibias.n190 161.3
R19759 commonsourceibias.n189 commonsourceibias.n141 161.3
R19760 commonsourceibias.n188 commonsourceibias.n187 161.3
R19761 commonsourceibias.n185 commonsourceibias.n142 161.3
R19762 commonsourceibias.n184 commonsourceibias.n183 161.3
R19763 commonsourceibias.n182 commonsourceibias.n143 161.3
R19764 commonsourceibias.n181 commonsourceibias.n180 161.3
R19765 commonsourceibias.n179 commonsourceibias.n144 161.3
R19766 commonsourceibias.n177 commonsourceibias.n176 161.3
R19767 commonsourceibias.n175 commonsourceibias.n146 161.3
R19768 commonsourceibias.n174 commonsourceibias.n173 161.3
R19769 commonsourceibias.n171 commonsourceibias.n147 161.3
R19770 commonsourceibias.n170 commonsourceibias.n169 161.3
R19771 commonsourceibias.n168 commonsourceibias.n167 161.3
R19772 commonsourceibias.n166 commonsourceibias.n149 161.3
R19773 commonsourceibias.n165 commonsourceibias.n164 161.3
R19774 commonsourceibias.n163 commonsourceibias.n162 161.3
R19775 commonsourceibias.n161 commonsourceibias.n151 161.3
R19776 commonsourceibias.n160 commonsourceibias.n159 161.3
R19777 commonsourceibias.n158 commonsourceibias.n157 161.3
R19778 commonsourceibias.n156 commonsourceibias.n153 161.3
R19779 commonsourceibias.n303 commonsourceibias.n243 161.3
R19780 commonsourceibias.n302 commonsourceibias.n301 161.3
R19781 commonsourceibias.n300 commonsourceibias.n299 161.3
R19782 commonsourceibias.n298 commonsourceibias.n245 161.3
R19783 commonsourceibias.n296 commonsourceibias.n295 161.3
R19784 commonsourceibias.n294 commonsourceibias.n246 161.3
R19785 commonsourceibias.n293 commonsourceibias.n292 161.3
R19786 commonsourceibias.n290 commonsourceibias.n247 161.3
R19787 commonsourceibias.n289 commonsourceibias.n288 161.3
R19788 commonsourceibias.n287 commonsourceibias.n248 161.3
R19789 commonsourceibias.n286 commonsourceibias.n285 161.3
R19790 commonsourceibias.n283 commonsourceibias.n249 161.3
R19791 commonsourceibias.n281 commonsourceibias.n280 161.3
R19792 commonsourceibias.n279 commonsourceibias.n250 161.3
R19793 commonsourceibias.n278 commonsourceibias.n277 161.3
R19794 commonsourceibias.n275 commonsourceibias.n251 161.3
R19795 commonsourceibias.n274 commonsourceibias.n273 161.3
R19796 commonsourceibias.n272 commonsourceibias.n271 161.3
R19797 commonsourceibias.n270 commonsourceibias.n253 161.3
R19798 commonsourceibias.n269 commonsourceibias.n268 161.3
R19799 commonsourceibias.n267 commonsourceibias.n266 161.3
R19800 commonsourceibias.n265 commonsourceibias.n255 161.3
R19801 commonsourceibias.n264 commonsourceibias.n263 161.3
R19802 commonsourceibias.n262 commonsourceibias.n261 161.3
R19803 commonsourceibias.n260 commonsourceibias.n257 161.3
R19804 commonsourceibias.n237 commonsourceibias.n236 161.3
R19805 commonsourceibias.n234 commonsourceibias.n210 161.3
R19806 commonsourceibias.n233 commonsourceibias.n232 161.3
R19807 commonsourceibias.n231 commonsourceibias.n230 161.3
R19808 commonsourceibias.n229 commonsourceibias.n212 161.3
R19809 commonsourceibias.n228 commonsourceibias.n227 161.3
R19810 commonsourceibias.n226 commonsourceibias.n225 161.3
R19811 commonsourceibias.n224 commonsourceibias.n214 161.3
R19812 commonsourceibias.n223 commonsourceibias.n222 161.3
R19813 commonsourceibias.n221 commonsourceibias.n220 161.3
R19814 commonsourceibias.n219 commonsourceibias.n216 161.3
R19815 commonsourceibias.n313 commonsourceibias.n209 161.3
R19816 commonsourceibias.n337 commonsourceibias.n202 161.3
R19817 commonsourceibias.n336 commonsourceibias.n335 161.3
R19818 commonsourceibias.n334 commonsourceibias.n333 161.3
R19819 commonsourceibias.n332 commonsourceibias.n204 161.3
R19820 commonsourceibias.n330 commonsourceibias.n329 161.3
R19821 commonsourceibias.n328 commonsourceibias.n205 161.3
R19822 commonsourceibias.n327 commonsourceibias.n326 161.3
R19823 commonsourceibias.n324 commonsourceibias.n206 161.3
R19824 commonsourceibias.n323 commonsourceibias.n322 161.3
R19825 commonsourceibias.n321 commonsourceibias.n207 161.3
R19826 commonsourceibias.n320 commonsourceibias.n319 161.3
R19827 commonsourceibias.n317 commonsourceibias.n208 161.3
R19828 commonsourceibias.n315 commonsourceibias.n314 161.3
R19829 commonsourceibias.n400 commonsourceibias.n340 161.3
R19830 commonsourceibias.n399 commonsourceibias.n398 161.3
R19831 commonsourceibias.n397 commonsourceibias.n396 161.3
R19832 commonsourceibias.n395 commonsourceibias.n342 161.3
R19833 commonsourceibias.n393 commonsourceibias.n392 161.3
R19834 commonsourceibias.n391 commonsourceibias.n343 161.3
R19835 commonsourceibias.n390 commonsourceibias.n389 161.3
R19836 commonsourceibias.n387 commonsourceibias.n344 161.3
R19837 commonsourceibias.n386 commonsourceibias.n385 161.3
R19838 commonsourceibias.n384 commonsourceibias.n345 161.3
R19839 commonsourceibias.n383 commonsourceibias.n382 161.3
R19840 commonsourceibias.n380 commonsourceibias.n346 161.3
R19841 commonsourceibias.n378 commonsourceibias.n377 161.3
R19842 commonsourceibias.n376 commonsourceibias.n347 161.3
R19843 commonsourceibias.n375 commonsourceibias.n374 161.3
R19844 commonsourceibias.n372 commonsourceibias.n348 161.3
R19845 commonsourceibias.n371 commonsourceibias.n370 161.3
R19846 commonsourceibias.n369 commonsourceibias.n368 161.3
R19847 commonsourceibias.n367 commonsourceibias.n350 161.3
R19848 commonsourceibias.n366 commonsourceibias.n365 161.3
R19849 commonsourceibias.n364 commonsourceibias.n363 161.3
R19850 commonsourceibias.n362 commonsourceibias.n352 161.3
R19851 commonsourceibias.n361 commonsourceibias.n360 161.3
R19852 commonsourceibias.n359 commonsourceibias.n358 161.3
R19853 commonsourceibias.n357 commonsourceibias.n354 161.3
R19854 commonsourceibias.n80 commonsourceibias.n78 81.5057
R19855 commonsourceibias.n240 commonsourceibias.n238 81.5057
R19856 commonsourceibias.n80 commonsourceibias.n79 80.9324
R19857 commonsourceibias.n82 commonsourceibias.n81 80.9324
R19858 commonsourceibias.n77 commonsourceibias.n76 80.9324
R19859 commonsourceibias.n75 commonsourceibias.n74 80.9324
R19860 commonsourceibias.n73 commonsourceibias.n72 80.9324
R19861 commonsourceibias.n307 commonsourceibias.n306 80.9324
R19862 commonsourceibias.n309 commonsourceibias.n308 80.9324
R19863 commonsourceibias.n311 commonsourceibias.n310 80.9324
R19864 commonsourceibias.n242 commonsourceibias.n241 80.9324
R19865 commonsourceibias.n240 commonsourceibias.n239 80.9324
R19866 commonsourceibias.n71 commonsourceibias.n70 80.6037
R19867 commonsourceibias.n137 commonsourceibias.n136 80.6037
R19868 commonsourceibias.n200 commonsourceibias.n199 80.6037
R19869 commonsourceibias.n305 commonsourceibias.n304 80.6037
R19870 commonsourceibias.n339 commonsourceibias.n338 80.6037
R19871 commonsourceibias.n402 commonsourceibias.n401 80.6037
R19872 commonsourceibias.n65 commonsourceibias.n64 56.5617
R19873 commonsourceibias.n51 commonsourceibias.n50 56.5617
R19874 commonsourceibias.n42 commonsourceibias.n41 56.5617
R19875 commonsourceibias.n28 commonsourceibias.n27 56.5617
R19876 commonsourceibias.n131 commonsourceibias.n130 56.5617
R19877 commonsourceibias.n117 commonsourceibias.n116 56.5617
R19878 commonsourceibias.n108 commonsourceibias.n107 56.5617
R19879 commonsourceibias.n94 commonsourceibias.n93 56.5617
R19880 commonsourceibias.n157 commonsourceibias.n156 56.5617
R19881 commonsourceibias.n171 commonsourceibias.n170 56.5617
R19882 commonsourceibias.n180 commonsourceibias.n179 56.5617
R19883 commonsourceibias.n194 commonsourceibias.n193 56.5617
R19884 commonsourceibias.n261 commonsourceibias.n260 56.5617
R19885 commonsourceibias.n275 commonsourceibias.n274 56.5617
R19886 commonsourceibias.n285 commonsourceibias.n283 56.5617
R19887 commonsourceibias.n299 commonsourceibias.n298 56.5617
R19888 commonsourceibias.n333 commonsourceibias.n332 56.5617
R19889 commonsourceibias.n319 commonsourceibias.n317 56.5617
R19890 commonsourceibias.n220 commonsourceibias.n219 56.5617
R19891 commonsourceibias.n234 commonsourceibias.n233 56.5617
R19892 commonsourceibias.n358 commonsourceibias.n357 56.5617
R19893 commonsourceibias.n372 commonsourceibias.n371 56.5617
R19894 commonsourceibias.n382 commonsourceibias.n380 56.5617
R19895 commonsourceibias.n396 commonsourceibias.n395 56.5617
R19896 commonsourceibias.n56 commonsourceibias.n55 56.0773
R19897 commonsourceibias.n37 commonsourceibias.n36 56.0773
R19898 commonsourceibias.n122 commonsourceibias.n121 56.0773
R19899 commonsourceibias.n103 commonsourceibias.n102 56.0773
R19900 commonsourceibias.n166 commonsourceibias.n165 56.0773
R19901 commonsourceibias.n185 commonsourceibias.n184 56.0773
R19902 commonsourceibias.n270 commonsourceibias.n269 56.0773
R19903 commonsourceibias.n290 commonsourceibias.n289 56.0773
R19904 commonsourceibias.n324 commonsourceibias.n323 56.0773
R19905 commonsourceibias.n229 commonsourceibias.n228 56.0773
R19906 commonsourceibias.n367 commonsourceibias.n366 56.0773
R19907 commonsourceibias.n387 commonsourceibias.n386 56.0773
R19908 commonsourceibias.n70 commonsourceibias.n69 46.0096
R19909 commonsourceibias.n136 commonsourceibias.n135 46.0096
R19910 commonsourceibias.n199 commonsourceibias.n198 46.0096
R19911 commonsourceibias.n304 commonsourceibias.n303 46.0096
R19912 commonsourceibias.n338 commonsourceibias.n337 46.0096
R19913 commonsourceibias.n401 commonsourceibias.n400 46.0096
R19914 commonsourceibias.n58 commonsourceibias.n12 41.5458
R19915 commonsourceibias.n33 commonsourceibias.n32 41.5458
R19916 commonsourceibias.n124 commonsourceibias.n3 41.5458
R19917 commonsourceibias.n99 commonsourceibias.n98 41.5458
R19918 commonsourceibias.n162 commonsourceibias.n161 41.5458
R19919 commonsourceibias.n187 commonsourceibias.n141 41.5458
R19920 commonsourceibias.n266 commonsourceibias.n265 41.5458
R19921 commonsourceibias.n292 commonsourceibias.n246 41.5458
R19922 commonsourceibias.n326 commonsourceibias.n205 41.5458
R19923 commonsourceibias.n225 commonsourceibias.n224 41.5458
R19924 commonsourceibias.n363 commonsourceibias.n362 41.5458
R19925 commonsourceibias.n389 commonsourceibias.n343 41.5458
R19926 commonsourceibias.n48 commonsourceibias.n17 40.577
R19927 commonsourceibias.n44 commonsourceibias.n17 40.577
R19928 commonsourceibias.n114 commonsourceibias.n8 40.577
R19929 commonsourceibias.n110 commonsourceibias.n8 40.577
R19930 commonsourceibias.n173 commonsourceibias.n146 40.577
R19931 commonsourceibias.n177 commonsourceibias.n146 40.577
R19932 commonsourceibias.n277 commonsourceibias.n250 40.577
R19933 commonsourceibias.n281 commonsourceibias.n250 40.577
R19934 commonsourceibias.n315 commonsourceibias.n209 40.577
R19935 commonsourceibias.n236 commonsourceibias.n209 40.577
R19936 commonsourceibias.n374 commonsourceibias.n347 40.577
R19937 commonsourceibias.n378 commonsourceibias.n347 40.577
R19938 commonsourceibias.n62 commonsourceibias.n12 39.6083
R19939 commonsourceibias.n32 commonsourceibias.n31 39.6083
R19940 commonsourceibias.n128 commonsourceibias.n3 39.6083
R19941 commonsourceibias.n98 commonsourceibias.n97 39.6083
R19942 commonsourceibias.n161 commonsourceibias.n160 39.6083
R19943 commonsourceibias.n191 commonsourceibias.n141 39.6083
R19944 commonsourceibias.n265 commonsourceibias.n264 39.6083
R19945 commonsourceibias.n296 commonsourceibias.n246 39.6083
R19946 commonsourceibias.n330 commonsourceibias.n205 39.6083
R19947 commonsourceibias.n224 commonsourceibias.n223 39.6083
R19948 commonsourceibias.n362 commonsourceibias.n361 39.6083
R19949 commonsourceibias.n393 commonsourceibias.n343 39.6083
R19950 commonsourceibias.n26 commonsourceibias.n25 33.0515
R19951 commonsourceibias.n92 commonsourceibias.n91 33.0515
R19952 commonsourceibias.n155 commonsourceibias.n154 33.0515
R19953 commonsourceibias.n259 commonsourceibias.n258 33.0515
R19954 commonsourceibias.n218 commonsourceibias.n217 33.0515
R19955 commonsourceibias.n356 commonsourceibias.n355 33.0515
R19956 commonsourceibias.n25 commonsourceibias.n24 28.5514
R19957 commonsourceibias.n91 commonsourceibias.n90 28.5514
R19958 commonsourceibias.n154 commonsourceibias.n153 28.5514
R19959 commonsourceibias.n258 commonsourceibias.n257 28.5514
R19960 commonsourceibias.n217 commonsourceibias.n216 28.5514
R19961 commonsourceibias.n355 commonsourceibias.n354 28.5514
R19962 commonsourceibias.n69 commonsourceibias.n68 26.0455
R19963 commonsourceibias.n135 commonsourceibias.n134 26.0455
R19964 commonsourceibias.n198 commonsourceibias.n197 26.0455
R19965 commonsourceibias.n303 commonsourceibias.n302 26.0455
R19966 commonsourceibias.n337 commonsourceibias.n336 26.0455
R19967 commonsourceibias.n400 commonsourceibias.n399 26.0455
R19968 commonsourceibias.n55 commonsourceibias.n14 25.0767
R19969 commonsourceibias.n38 commonsourceibias.n37 25.0767
R19970 commonsourceibias.n121 commonsourceibias.n5 25.0767
R19971 commonsourceibias.n104 commonsourceibias.n103 25.0767
R19972 commonsourceibias.n167 commonsourceibias.n166 25.0767
R19973 commonsourceibias.n184 commonsourceibias.n143 25.0767
R19974 commonsourceibias.n271 commonsourceibias.n270 25.0767
R19975 commonsourceibias.n289 commonsourceibias.n248 25.0767
R19976 commonsourceibias.n323 commonsourceibias.n207 25.0767
R19977 commonsourceibias.n230 commonsourceibias.n229 25.0767
R19978 commonsourceibias.n368 commonsourceibias.n367 25.0767
R19979 commonsourceibias.n386 commonsourceibias.n345 25.0767
R19980 commonsourceibias.n51 commonsourceibias.n16 24.3464
R19981 commonsourceibias.n41 commonsourceibias.n19 24.3464
R19982 commonsourceibias.n117 commonsourceibias.n7 24.3464
R19983 commonsourceibias.n107 commonsourceibias.n85 24.3464
R19984 commonsourceibias.n170 commonsourceibias.n148 24.3464
R19985 commonsourceibias.n180 commonsourceibias.n145 24.3464
R19986 commonsourceibias.n274 commonsourceibias.n252 24.3464
R19987 commonsourceibias.n285 commonsourceibias.n284 24.3464
R19988 commonsourceibias.n319 commonsourceibias.n318 24.3464
R19989 commonsourceibias.n233 commonsourceibias.n211 24.3464
R19990 commonsourceibias.n371 commonsourceibias.n349 24.3464
R19991 commonsourceibias.n382 commonsourceibias.n381 24.3464
R19992 commonsourceibias.n65 commonsourceibias.n10 23.8546
R19993 commonsourceibias.n27 commonsourceibias.n26 23.8546
R19994 commonsourceibias.n131 commonsourceibias.n1 23.8546
R19995 commonsourceibias.n93 commonsourceibias.n92 23.8546
R19996 commonsourceibias.n156 commonsourceibias.n155 23.8546
R19997 commonsourceibias.n194 commonsourceibias.n139 23.8546
R19998 commonsourceibias.n260 commonsourceibias.n259 23.8546
R19999 commonsourceibias.n299 commonsourceibias.n244 23.8546
R20000 commonsourceibias.n333 commonsourceibias.n203 23.8546
R20001 commonsourceibias.n219 commonsourceibias.n218 23.8546
R20002 commonsourceibias.n357 commonsourceibias.n356 23.8546
R20003 commonsourceibias.n396 commonsourceibias.n341 23.8546
R20004 commonsourceibias.n64 commonsourceibias.n63 16.9689
R20005 commonsourceibias.n28 commonsourceibias.n23 16.9689
R20006 commonsourceibias.n130 commonsourceibias.n129 16.9689
R20007 commonsourceibias.n94 commonsourceibias.n89 16.9689
R20008 commonsourceibias.n157 commonsourceibias.n152 16.9689
R20009 commonsourceibias.n193 commonsourceibias.n192 16.9689
R20010 commonsourceibias.n261 commonsourceibias.n256 16.9689
R20011 commonsourceibias.n298 commonsourceibias.n297 16.9689
R20012 commonsourceibias.n332 commonsourceibias.n331 16.9689
R20013 commonsourceibias.n220 commonsourceibias.n215 16.9689
R20014 commonsourceibias.n358 commonsourceibias.n353 16.9689
R20015 commonsourceibias.n395 commonsourceibias.n394 16.9689
R20016 commonsourceibias.n50 commonsourceibias.n49 16.477
R20017 commonsourceibias.n43 commonsourceibias.n42 16.477
R20018 commonsourceibias.n116 commonsourceibias.n115 16.477
R20019 commonsourceibias.n109 commonsourceibias.n108 16.477
R20020 commonsourceibias.n172 commonsourceibias.n171 16.477
R20021 commonsourceibias.n179 commonsourceibias.n178 16.477
R20022 commonsourceibias.n276 commonsourceibias.n275 16.477
R20023 commonsourceibias.n283 commonsourceibias.n282 16.477
R20024 commonsourceibias.n317 commonsourceibias.n316 16.477
R20025 commonsourceibias.n235 commonsourceibias.n234 16.477
R20026 commonsourceibias.n373 commonsourceibias.n372 16.477
R20027 commonsourceibias.n380 commonsourceibias.n379 16.477
R20028 commonsourceibias.n57 commonsourceibias.n56 15.9852
R20029 commonsourceibias.n36 commonsourceibias.n21 15.9852
R20030 commonsourceibias.n123 commonsourceibias.n122 15.9852
R20031 commonsourceibias.n102 commonsourceibias.n87 15.9852
R20032 commonsourceibias.n165 commonsourceibias.n150 15.9852
R20033 commonsourceibias.n186 commonsourceibias.n185 15.9852
R20034 commonsourceibias.n269 commonsourceibias.n254 15.9852
R20035 commonsourceibias.n291 commonsourceibias.n290 15.9852
R20036 commonsourceibias.n325 commonsourceibias.n324 15.9852
R20037 commonsourceibias.n228 commonsourceibias.n213 15.9852
R20038 commonsourceibias.n366 commonsourceibias.n351 15.9852
R20039 commonsourceibias.n388 commonsourceibias.n387 15.9852
R20040 commonsourceibias.n73 commonsourceibias.n71 13.2057
R20041 commonsourceibias.n307 commonsourceibias.n305 13.2057
R20042 commonsourceibias.n404 commonsourceibias.n201 11.9876
R20043 commonsourceibias.n404 commonsourceibias.n403 10.3347
R20044 commonsourceibias.n112 commonsourceibias.n83 9.50363
R20045 commonsourceibias.n313 commonsourceibias.n312 9.50363
R20046 commonsourceibias.n201 commonsourceibias.n137 8.732
R20047 commonsourceibias.n403 commonsourceibias.n339 8.732
R20048 commonsourceibias.n58 commonsourceibias.n57 8.60764
R20049 commonsourceibias.n33 commonsourceibias.n21 8.60764
R20050 commonsourceibias.n124 commonsourceibias.n123 8.60764
R20051 commonsourceibias.n99 commonsourceibias.n87 8.60764
R20052 commonsourceibias.n162 commonsourceibias.n150 8.60764
R20053 commonsourceibias.n187 commonsourceibias.n186 8.60764
R20054 commonsourceibias.n266 commonsourceibias.n254 8.60764
R20055 commonsourceibias.n292 commonsourceibias.n291 8.60764
R20056 commonsourceibias.n326 commonsourceibias.n325 8.60764
R20057 commonsourceibias.n225 commonsourceibias.n213 8.60764
R20058 commonsourceibias.n363 commonsourceibias.n351 8.60764
R20059 commonsourceibias.n389 commonsourceibias.n388 8.60764
R20060 commonsourceibias.n49 commonsourceibias.n48 8.11581
R20061 commonsourceibias.n44 commonsourceibias.n43 8.11581
R20062 commonsourceibias.n115 commonsourceibias.n114 8.11581
R20063 commonsourceibias.n110 commonsourceibias.n109 8.11581
R20064 commonsourceibias.n173 commonsourceibias.n172 8.11581
R20065 commonsourceibias.n178 commonsourceibias.n177 8.11581
R20066 commonsourceibias.n277 commonsourceibias.n276 8.11581
R20067 commonsourceibias.n282 commonsourceibias.n281 8.11581
R20068 commonsourceibias.n316 commonsourceibias.n315 8.11581
R20069 commonsourceibias.n236 commonsourceibias.n235 8.11581
R20070 commonsourceibias.n374 commonsourceibias.n373 8.11581
R20071 commonsourceibias.n379 commonsourceibias.n378 8.11581
R20072 commonsourceibias.n63 commonsourceibias.n62 7.62397
R20073 commonsourceibias.n31 commonsourceibias.n23 7.62397
R20074 commonsourceibias.n129 commonsourceibias.n128 7.62397
R20075 commonsourceibias.n97 commonsourceibias.n89 7.62397
R20076 commonsourceibias.n160 commonsourceibias.n152 7.62397
R20077 commonsourceibias.n192 commonsourceibias.n191 7.62397
R20078 commonsourceibias.n264 commonsourceibias.n256 7.62397
R20079 commonsourceibias.n297 commonsourceibias.n296 7.62397
R20080 commonsourceibias.n331 commonsourceibias.n330 7.62397
R20081 commonsourceibias.n223 commonsourceibias.n215 7.62397
R20082 commonsourceibias.n361 commonsourceibias.n353 7.62397
R20083 commonsourceibias.n394 commonsourceibias.n393 7.62397
R20084 commonsourceibias.n201 commonsourceibias.n200 5.00473
R20085 commonsourceibias.n403 commonsourceibias.n402 5.00473
R20086 commonsourceibias commonsourceibias.n404 3.87639
R20087 commonsourceibias.n78 commonsourceibias.t41 2.82907
R20088 commonsourceibias.n78 commonsourceibias.t47 2.82907
R20089 commonsourceibias.n79 commonsourceibias.t35 2.82907
R20090 commonsourceibias.n79 commonsourceibias.t11 2.82907
R20091 commonsourceibias.n81 commonsourceibias.t45 2.82907
R20092 commonsourceibias.n81 commonsourceibias.t27 2.82907
R20093 commonsourceibias.n76 commonsourceibias.t21 2.82907
R20094 commonsourceibias.n76 commonsourceibias.t37 2.82907
R20095 commonsourceibias.n74 commonsourceibias.t25 2.82907
R20096 commonsourceibias.n74 commonsourceibias.t31 2.82907
R20097 commonsourceibias.n72 commonsourceibias.t33 2.82907
R20098 commonsourceibias.n72 commonsourceibias.t15 2.82907
R20099 commonsourceibias.n306 commonsourceibias.t23 2.82907
R20100 commonsourceibias.n306 commonsourceibias.t3 2.82907
R20101 commonsourceibias.n308 commonsourceibias.t1 2.82907
R20102 commonsourceibias.n308 commonsourceibias.t39 2.82907
R20103 commonsourceibias.n310 commonsourceibias.t7 2.82907
R20104 commonsourceibias.n310 commonsourceibias.t29 2.82907
R20105 commonsourceibias.n241 commonsourceibias.t43 2.82907
R20106 commonsourceibias.n241 commonsourceibias.t13 2.82907
R20107 commonsourceibias.n239 commonsourceibias.t19 2.82907
R20108 commonsourceibias.n239 commonsourceibias.t5 2.82907
R20109 commonsourceibias.n238 commonsourceibias.t17 2.82907
R20110 commonsourceibias.n238 commonsourceibias.t9 2.82907
R20111 commonsourceibias.n68 commonsourceibias.n10 0.738255
R20112 commonsourceibias.n134 commonsourceibias.n1 0.738255
R20113 commonsourceibias.n197 commonsourceibias.n139 0.738255
R20114 commonsourceibias.n302 commonsourceibias.n244 0.738255
R20115 commonsourceibias.n336 commonsourceibias.n203 0.738255
R20116 commonsourceibias.n399 commonsourceibias.n341 0.738255
R20117 commonsourceibias.n75 commonsourceibias.n73 0.573776
R20118 commonsourceibias.n77 commonsourceibias.n75 0.573776
R20119 commonsourceibias.n82 commonsourceibias.n80 0.573776
R20120 commonsourceibias.n242 commonsourceibias.n240 0.573776
R20121 commonsourceibias.n311 commonsourceibias.n309 0.573776
R20122 commonsourceibias.n309 commonsourceibias.n307 0.573776
R20123 commonsourceibias.n83 commonsourceibias.n77 0.287138
R20124 commonsourceibias.n83 commonsourceibias.n82 0.287138
R20125 commonsourceibias.n312 commonsourceibias.n242 0.287138
R20126 commonsourceibias.n312 commonsourceibias.n311 0.287138
R20127 commonsourceibias.n71 commonsourceibias.n9 0.285035
R20128 commonsourceibias.n137 commonsourceibias.n0 0.285035
R20129 commonsourceibias.n200 commonsourceibias.n138 0.285035
R20130 commonsourceibias.n305 commonsourceibias.n243 0.285035
R20131 commonsourceibias.n339 commonsourceibias.n202 0.285035
R20132 commonsourceibias.n402 commonsourceibias.n340 0.285035
R20133 commonsourceibias.n16 commonsourceibias.n14 0.246418
R20134 commonsourceibias.n38 commonsourceibias.n19 0.246418
R20135 commonsourceibias.n7 commonsourceibias.n5 0.246418
R20136 commonsourceibias.n104 commonsourceibias.n85 0.246418
R20137 commonsourceibias.n167 commonsourceibias.n148 0.246418
R20138 commonsourceibias.n145 commonsourceibias.n143 0.246418
R20139 commonsourceibias.n271 commonsourceibias.n252 0.246418
R20140 commonsourceibias.n284 commonsourceibias.n248 0.246418
R20141 commonsourceibias.n318 commonsourceibias.n207 0.246418
R20142 commonsourceibias.n230 commonsourceibias.n211 0.246418
R20143 commonsourceibias.n368 commonsourceibias.n349 0.246418
R20144 commonsourceibias.n381 commonsourceibias.n345 0.246418
R20145 commonsourceibias.n67 commonsourceibias.n9 0.189894
R20146 commonsourceibias.n67 commonsourceibias.n66 0.189894
R20147 commonsourceibias.n66 commonsourceibias.n11 0.189894
R20148 commonsourceibias.n61 commonsourceibias.n11 0.189894
R20149 commonsourceibias.n61 commonsourceibias.n60 0.189894
R20150 commonsourceibias.n60 commonsourceibias.n59 0.189894
R20151 commonsourceibias.n59 commonsourceibias.n13 0.189894
R20152 commonsourceibias.n54 commonsourceibias.n13 0.189894
R20153 commonsourceibias.n54 commonsourceibias.n53 0.189894
R20154 commonsourceibias.n53 commonsourceibias.n52 0.189894
R20155 commonsourceibias.n52 commonsourceibias.n15 0.189894
R20156 commonsourceibias.n47 commonsourceibias.n15 0.189894
R20157 commonsourceibias.n47 commonsourceibias.n46 0.189894
R20158 commonsourceibias.n46 commonsourceibias.n45 0.189894
R20159 commonsourceibias.n45 commonsourceibias.n18 0.189894
R20160 commonsourceibias.n40 commonsourceibias.n18 0.189894
R20161 commonsourceibias.n40 commonsourceibias.n39 0.189894
R20162 commonsourceibias.n39 commonsourceibias.n20 0.189894
R20163 commonsourceibias.n35 commonsourceibias.n20 0.189894
R20164 commonsourceibias.n35 commonsourceibias.n34 0.189894
R20165 commonsourceibias.n34 commonsourceibias.n22 0.189894
R20166 commonsourceibias.n30 commonsourceibias.n22 0.189894
R20167 commonsourceibias.n30 commonsourceibias.n29 0.189894
R20168 commonsourceibias.n29 commonsourceibias.n24 0.189894
R20169 commonsourceibias.n111 commonsourceibias.n84 0.189894
R20170 commonsourceibias.n106 commonsourceibias.n84 0.189894
R20171 commonsourceibias.n106 commonsourceibias.n105 0.189894
R20172 commonsourceibias.n105 commonsourceibias.n86 0.189894
R20173 commonsourceibias.n101 commonsourceibias.n86 0.189894
R20174 commonsourceibias.n101 commonsourceibias.n100 0.189894
R20175 commonsourceibias.n100 commonsourceibias.n88 0.189894
R20176 commonsourceibias.n96 commonsourceibias.n88 0.189894
R20177 commonsourceibias.n96 commonsourceibias.n95 0.189894
R20178 commonsourceibias.n95 commonsourceibias.n90 0.189894
R20179 commonsourceibias.n133 commonsourceibias.n0 0.189894
R20180 commonsourceibias.n133 commonsourceibias.n132 0.189894
R20181 commonsourceibias.n132 commonsourceibias.n2 0.189894
R20182 commonsourceibias.n127 commonsourceibias.n2 0.189894
R20183 commonsourceibias.n127 commonsourceibias.n126 0.189894
R20184 commonsourceibias.n126 commonsourceibias.n125 0.189894
R20185 commonsourceibias.n125 commonsourceibias.n4 0.189894
R20186 commonsourceibias.n120 commonsourceibias.n4 0.189894
R20187 commonsourceibias.n120 commonsourceibias.n119 0.189894
R20188 commonsourceibias.n119 commonsourceibias.n118 0.189894
R20189 commonsourceibias.n118 commonsourceibias.n6 0.189894
R20190 commonsourceibias.n113 commonsourceibias.n6 0.189894
R20191 commonsourceibias.n196 commonsourceibias.n138 0.189894
R20192 commonsourceibias.n196 commonsourceibias.n195 0.189894
R20193 commonsourceibias.n195 commonsourceibias.n140 0.189894
R20194 commonsourceibias.n190 commonsourceibias.n140 0.189894
R20195 commonsourceibias.n190 commonsourceibias.n189 0.189894
R20196 commonsourceibias.n189 commonsourceibias.n188 0.189894
R20197 commonsourceibias.n188 commonsourceibias.n142 0.189894
R20198 commonsourceibias.n183 commonsourceibias.n142 0.189894
R20199 commonsourceibias.n183 commonsourceibias.n182 0.189894
R20200 commonsourceibias.n182 commonsourceibias.n181 0.189894
R20201 commonsourceibias.n181 commonsourceibias.n144 0.189894
R20202 commonsourceibias.n176 commonsourceibias.n144 0.189894
R20203 commonsourceibias.n176 commonsourceibias.n175 0.189894
R20204 commonsourceibias.n175 commonsourceibias.n174 0.189894
R20205 commonsourceibias.n174 commonsourceibias.n147 0.189894
R20206 commonsourceibias.n169 commonsourceibias.n147 0.189894
R20207 commonsourceibias.n169 commonsourceibias.n168 0.189894
R20208 commonsourceibias.n168 commonsourceibias.n149 0.189894
R20209 commonsourceibias.n164 commonsourceibias.n149 0.189894
R20210 commonsourceibias.n164 commonsourceibias.n163 0.189894
R20211 commonsourceibias.n163 commonsourceibias.n151 0.189894
R20212 commonsourceibias.n159 commonsourceibias.n151 0.189894
R20213 commonsourceibias.n159 commonsourceibias.n158 0.189894
R20214 commonsourceibias.n158 commonsourceibias.n153 0.189894
R20215 commonsourceibias.n262 commonsourceibias.n257 0.189894
R20216 commonsourceibias.n263 commonsourceibias.n262 0.189894
R20217 commonsourceibias.n263 commonsourceibias.n255 0.189894
R20218 commonsourceibias.n267 commonsourceibias.n255 0.189894
R20219 commonsourceibias.n268 commonsourceibias.n267 0.189894
R20220 commonsourceibias.n268 commonsourceibias.n253 0.189894
R20221 commonsourceibias.n272 commonsourceibias.n253 0.189894
R20222 commonsourceibias.n273 commonsourceibias.n272 0.189894
R20223 commonsourceibias.n273 commonsourceibias.n251 0.189894
R20224 commonsourceibias.n278 commonsourceibias.n251 0.189894
R20225 commonsourceibias.n279 commonsourceibias.n278 0.189894
R20226 commonsourceibias.n280 commonsourceibias.n279 0.189894
R20227 commonsourceibias.n280 commonsourceibias.n249 0.189894
R20228 commonsourceibias.n286 commonsourceibias.n249 0.189894
R20229 commonsourceibias.n287 commonsourceibias.n286 0.189894
R20230 commonsourceibias.n288 commonsourceibias.n287 0.189894
R20231 commonsourceibias.n288 commonsourceibias.n247 0.189894
R20232 commonsourceibias.n293 commonsourceibias.n247 0.189894
R20233 commonsourceibias.n294 commonsourceibias.n293 0.189894
R20234 commonsourceibias.n295 commonsourceibias.n294 0.189894
R20235 commonsourceibias.n295 commonsourceibias.n245 0.189894
R20236 commonsourceibias.n300 commonsourceibias.n245 0.189894
R20237 commonsourceibias.n301 commonsourceibias.n300 0.189894
R20238 commonsourceibias.n301 commonsourceibias.n243 0.189894
R20239 commonsourceibias.n221 commonsourceibias.n216 0.189894
R20240 commonsourceibias.n222 commonsourceibias.n221 0.189894
R20241 commonsourceibias.n222 commonsourceibias.n214 0.189894
R20242 commonsourceibias.n226 commonsourceibias.n214 0.189894
R20243 commonsourceibias.n227 commonsourceibias.n226 0.189894
R20244 commonsourceibias.n227 commonsourceibias.n212 0.189894
R20245 commonsourceibias.n231 commonsourceibias.n212 0.189894
R20246 commonsourceibias.n232 commonsourceibias.n231 0.189894
R20247 commonsourceibias.n232 commonsourceibias.n210 0.189894
R20248 commonsourceibias.n237 commonsourceibias.n210 0.189894
R20249 commonsourceibias.n314 commonsourceibias.n208 0.189894
R20250 commonsourceibias.n320 commonsourceibias.n208 0.189894
R20251 commonsourceibias.n321 commonsourceibias.n320 0.189894
R20252 commonsourceibias.n322 commonsourceibias.n321 0.189894
R20253 commonsourceibias.n322 commonsourceibias.n206 0.189894
R20254 commonsourceibias.n327 commonsourceibias.n206 0.189894
R20255 commonsourceibias.n328 commonsourceibias.n327 0.189894
R20256 commonsourceibias.n329 commonsourceibias.n328 0.189894
R20257 commonsourceibias.n329 commonsourceibias.n204 0.189894
R20258 commonsourceibias.n334 commonsourceibias.n204 0.189894
R20259 commonsourceibias.n335 commonsourceibias.n334 0.189894
R20260 commonsourceibias.n335 commonsourceibias.n202 0.189894
R20261 commonsourceibias.n359 commonsourceibias.n354 0.189894
R20262 commonsourceibias.n360 commonsourceibias.n359 0.189894
R20263 commonsourceibias.n360 commonsourceibias.n352 0.189894
R20264 commonsourceibias.n364 commonsourceibias.n352 0.189894
R20265 commonsourceibias.n365 commonsourceibias.n364 0.189894
R20266 commonsourceibias.n365 commonsourceibias.n350 0.189894
R20267 commonsourceibias.n369 commonsourceibias.n350 0.189894
R20268 commonsourceibias.n370 commonsourceibias.n369 0.189894
R20269 commonsourceibias.n370 commonsourceibias.n348 0.189894
R20270 commonsourceibias.n375 commonsourceibias.n348 0.189894
R20271 commonsourceibias.n376 commonsourceibias.n375 0.189894
R20272 commonsourceibias.n377 commonsourceibias.n376 0.189894
R20273 commonsourceibias.n377 commonsourceibias.n346 0.189894
R20274 commonsourceibias.n383 commonsourceibias.n346 0.189894
R20275 commonsourceibias.n384 commonsourceibias.n383 0.189894
R20276 commonsourceibias.n385 commonsourceibias.n384 0.189894
R20277 commonsourceibias.n385 commonsourceibias.n344 0.189894
R20278 commonsourceibias.n390 commonsourceibias.n344 0.189894
R20279 commonsourceibias.n391 commonsourceibias.n390 0.189894
R20280 commonsourceibias.n392 commonsourceibias.n391 0.189894
R20281 commonsourceibias.n392 commonsourceibias.n342 0.189894
R20282 commonsourceibias.n397 commonsourceibias.n342 0.189894
R20283 commonsourceibias.n398 commonsourceibias.n397 0.189894
R20284 commonsourceibias.n398 commonsourceibias.n340 0.189894
R20285 commonsourceibias.n112 commonsourceibias.n111 0.170955
R20286 commonsourceibias.n113 commonsourceibias.n112 0.170955
R20287 commonsourceibias.n313 commonsourceibias.n237 0.170955
R20288 commonsourceibias.n314 commonsourceibias.n313 0.170955
R20289 minus.n53 minus.t28 323.478
R20290 minus.n11 minus.t8 323.478
R20291 minus.n82 minus.t12 297.12
R20292 minus.n80 minus.t15 297.12
R20293 minus.n44 minus.t5 297.12
R20294 minus.n74 minus.t6 297.12
R20295 minus.n46 minus.t26 297.12
R20296 minus.n68 minus.t21 297.12
R20297 minus.n48 minus.t23 297.12
R20298 minus.n62 minus.t16 297.12
R20299 minus.n50 minus.t17 297.12
R20300 minus.n56 minus.t9 297.12
R20301 minus.n52 minus.t27 297.12
R20302 minus.n10 minus.t7 297.12
R20303 minus.n14 minus.t11 297.12
R20304 minus.n16 minus.t10 297.12
R20305 minus.n20 minus.t13 297.12
R20306 minus.n22 minus.t20 297.12
R20307 minus.n26 minus.t18 297.12
R20308 minus.n28 minus.t25 297.12
R20309 minus.n32 minus.t24 297.12
R20310 minus.n34 minus.t14 297.12
R20311 minus.n38 minus.t22 297.12
R20312 minus.n40 minus.t19 297.12
R20313 minus.n88 minus.t2 243.255
R20314 minus.n87 minus.n85 224.169
R20315 minus.n87 minus.n86 223.454
R20316 minus.n55 minus.n54 161.3
R20317 minus.n56 minus.n51 161.3
R20318 minus.n58 minus.n57 161.3
R20319 minus.n59 minus.n50 161.3
R20320 minus.n61 minus.n60 161.3
R20321 minus.n62 minus.n49 161.3
R20322 minus.n64 minus.n63 161.3
R20323 minus.n65 minus.n48 161.3
R20324 minus.n67 minus.n66 161.3
R20325 minus.n68 minus.n47 161.3
R20326 minus.n70 minus.n69 161.3
R20327 minus.n71 minus.n46 161.3
R20328 minus.n73 minus.n72 161.3
R20329 minus.n74 minus.n45 161.3
R20330 minus.n76 minus.n75 161.3
R20331 minus.n77 minus.n44 161.3
R20332 minus.n79 minus.n78 161.3
R20333 minus.n80 minus.n43 161.3
R20334 minus.n81 minus.n42 161.3
R20335 minus.n83 minus.n82 161.3
R20336 minus.n41 minus.n40 161.3
R20337 minus.n39 minus.n0 161.3
R20338 minus.n38 minus.n37 161.3
R20339 minus.n36 minus.n1 161.3
R20340 minus.n35 minus.n34 161.3
R20341 minus.n33 minus.n2 161.3
R20342 minus.n32 minus.n31 161.3
R20343 minus.n30 minus.n3 161.3
R20344 minus.n29 minus.n28 161.3
R20345 minus.n27 minus.n4 161.3
R20346 minus.n26 minus.n25 161.3
R20347 minus.n24 minus.n5 161.3
R20348 minus.n23 minus.n22 161.3
R20349 minus.n21 minus.n6 161.3
R20350 minus.n20 minus.n19 161.3
R20351 minus.n18 minus.n7 161.3
R20352 minus.n17 minus.n16 161.3
R20353 minus.n15 minus.n8 161.3
R20354 minus.n14 minus.n13 161.3
R20355 minus.n12 minus.n9 161.3
R20356 minus.n82 minus.n81 46.0096
R20357 minus.n40 minus.n39 46.0096
R20358 minus.n12 minus.n11 45.0871
R20359 minus.n54 minus.n53 45.0871
R20360 minus.n80 minus.n79 41.6278
R20361 minus.n55 minus.n52 41.6278
R20362 minus.n10 minus.n9 41.6278
R20363 minus.n38 minus.n1 41.6278
R20364 minus.n75 minus.n44 37.246
R20365 minus.n57 minus.n56 37.246
R20366 minus.n15 minus.n14 37.246
R20367 minus.n34 minus.n33 37.246
R20368 minus.n84 minus.n83 33.3925
R20369 minus.n74 minus.n73 32.8641
R20370 minus.n61 minus.n50 32.8641
R20371 minus.n16 minus.n7 32.8641
R20372 minus.n32 minus.n3 32.8641
R20373 minus.n69 minus.n46 28.4823
R20374 minus.n63 minus.n62 28.4823
R20375 minus.n21 minus.n20 28.4823
R20376 minus.n28 minus.n27 28.4823
R20377 minus.n68 minus.n67 24.1005
R20378 minus.n67 minus.n48 24.1005
R20379 minus.n22 minus.n5 24.1005
R20380 minus.n26 minus.n5 24.1005
R20381 minus.n86 minus.t4 19.8005
R20382 minus.n86 minus.t3 19.8005
R20383 minus.n85 minus.t1 19.8005
R20384 minus.n85 minus.t0 19.8005
R20385 minus.n69 minus.n68 19.7187
R20386 minus.n63 minus.n48 19.7187
R20387 minus.n22 minus.n21 19.7187
R20388 minus.n27 minus.n26 19.7187
R20389 minus.n73 minus.n46 15.3369
R20390 minus.n62 minus.n61 15.3369
R20391 minus.n20 minus.n7 15.3369
R20392 minus.n28 minus.n3 15.3369
R20393 minus.n53 minus.n52 14.1472
R20394 minus.n11 minus.n10 14.1472
R20395 minus.n84 minus.n41 12.0933
R20396 minus minus.n89 11.0787
R20397 minus.n75 minus.n74 10.955
R20398 minus.n57 minus.n50 10.955
R20399 minus.n16 minus.n15 10.955
R20400 minus.n33 minus.n32 10.955
R20401 minus.n79 minus.n44 6.57323
R20402 minus.n56 minus.n55 6.57323
R20403 minus.n14 minus.n9 6.57323
R20404 minus.n34 minus.n1 6.57323
R20405 minus.n89 minus.n88 4.80222
R20406 minus.n81 minus.n80 2.19141
R20407 minus.n39 minus.n38 2.19141
R20408 minus.n89 minus.n84 0.972091
R20409 minus.n88 minus.n87 0.716017
R20410 minus.n83 minus.n42 0.189894
R20411 minus.n43 minus.n42 0.189894
R20412 minus.n78 minus.n43 0.189894
R20413 minus.n78 minus.n77 0.189894
R20414 minus.n77 minus.n76 0.189894
R20415 minus.n76 minus.n45 0.189894
R20416 minus.n72 minus.n45 0.189894
R20417 minus.n72 minus.n71 0.189894
R20418 minus.n71 minus.n70 0.189894
R20419 minus.n70 minus.n47 0.189894
R20420 minus.n66 minus.n47 0.189894
R20421 minus.n66 minus.n65 0.189894
R20422 minus.n65 minus.n64 0.189894
R20423 minus.n64 minus.n49 0.189894
R20424 minus.n60 minus.n49 0.189894
R20425 minus.n60 minus.n59 0.189894
R20426 minus.n59 minus.n58 0.189894
R20427 minus.n58 minus.n51 0.189894
R20428 minus.n54 minus.n51 0.189894
R20429 minus.n13 minus.n12 0.189894
R20430 minus.n13 minus.n8 0.189894
R20431 minus.n17 minus.n8 0.189894
R20432 minus.n18 minus.n17 0.189894
R20433 minus.n19 minus.n18 0.189894
R20434 minus.n19 minus.n6 0.189894
R20435 minus.n23 minus.n6 0.189894
R20436 minus.n24 minus.n23 0.189894
R20437 minus.n25 minus.n24 0.189894
R20438 minus.n25 minus.n4 0.189894
R20439 minus.n29 minus.n4 0.189894
R20440 minus.n30 minus.n29 0.189894
R20441 minus.n31 minus.n30 0.189894
R20442 minus.n31 minus.n2 0.189894
R20443 minus.n35 minus.n2 0.189894
R20444 minus.n36 minus.n35 0.189894
R20445 minus.n37 minus.n36 0.189894
R20446 minus.n37 minus.n0 0.189894
R20447 minus.n41 minus.n0 0.189894
R20448 outputibias.n27 outputibias.n1 289.615
R20449 outputibias.n58 outputibias.n32 289.615
R20450 outputibias.n90 outputibias.n64 289.615
R20451 outputibias.n122 outputibias.n96 289.615
R20452 outputibias.n28 outputibias.n27 185
R20453 outputibias.n26 outputibias.n25 185
R20454 outputibias.n5 outputibias.n4 185
R20455 outputibias.n20 outputibias.n19 185
R20456 outputibias.n18 outputibias.n17 185
R20457 outputibias.n9 outputibias.n8 185
R20458 outputibias.n12 outputibias.n11 185
R20459 outputibias.n59 outputibias.n58 185
R20460 outputibias.n57 outputibias.n56 185
R20461 outputibias.n36 outputibias.n35 185
R20462 outputibias.n51 outputibias.n50 185
R20463 outputibias.n49 outputibias.n48 185
R20464 outputibias.n40 outputibias.n39 185
R20465 outputibias.n43 outputibias.n42 185
R20466 outputibias.n91 outputibias.n90 185
R20467 outputibias.n89 outputibias.n88 185
R20468 outputibias.n68 outputibias.n67 185
R20469 outputibias.n83 outputibias.n82 185
R20470 outputibias.n81 outputibias.n80 185
R20471 outputibias.n72 outputibias.n71 185
R20472 outputibias.n75 outputibias.n74 185
R20473 outputibias.n123 outputibias.n122 185
R20474 outputibias.n121 outputibias.n120 185
R20475 outputibias.n100 outputibias.n99 185
R20476 outputibias.n115 outputibias.n114 185
R20477 outputibias.n113 outputibias.n112 185
R20478 outputibias.n104 outputibias.n103 185
R20479 outputibias.n107 outputibias.n106 185
R20480 outputibias.n0 outputibias.t8 178.945
R20481 outputibias.n133 outputibias.t10 177.018
R20482 outputibias.n132 outputibias.t11 177.018
R20483 outputibias.n0 outputibias.t9 177.018
R20484 outputibias.t5 outputibias.n10 147.661
R20485 outputibias.t7 outputibias.n41 147.661
R20486 outputibias.t1 outputibias.n73 147.661
R20487 outputibias.t3 outputibias.n105 147.661
R20488 outputibias.n128 outputibias.t4 132.363
R20489 outputibias.n128 outputibias.t6 130.436
R20490 outputibias.n129 outputibias.t0 130.436
R20491 outputibias.n130 outputibias.t2 130.436
R20492 outputibias.n27 outputibias.n26 104.615
R20493 outputibias.n26 outputibias.n4 104.615
R20494 outputibias.n19 outputibias.n4 104.615
R20495 outputibias.n19 outputibias.n18 104.615
R20496 outputibias.n18 outputibias.n8 104.615
R20497 outputibias.n11 outputibias.n8 104.615
R20498 outputibias.n58 outputibias.n57 104.615
R20499 outputibias.n57 outputibias.n35 104.615
R20500 outputibias.n50 outputibias.n35 104.615
R20501 outputibias.n50 outputibias.n49 104.615
R20502 outputibias.n49 outputibias.n39 104.615
R20503 outputibias.n42 outputibias.n39 104.615
R20504 outputibias.n90 outputibias.n89 104.615
R20505 outputibias.n89 outputibias.n67 104.615
R20506 outputibias.n82 outputibias.n67 104.615
R20507 outputibias.n82 outputibias.n81 104.615
R20508 outputibias.n81 outputibias.n71 104.615
R20509 outputibias.n74 outputibias.n71 104.615
R20510 outputibias.n122 outputibias.n121 104.615
R20511 outputibias.n121 outputibias.n99 104.615
R20512 outputibias.n114 outputibias.n99 104.615
R20513 outputibias.n114 outputibias.n113 104.615
R20514 outputibias.n113 outputibias.n103 104.615
R20515 outputibias.n106 outputibias.n103 104.615
R20516 outputibias.n63 outputibias.n31 95.6354
R20517 outputibias.n63 outputibias.n62 94.6732
R20518 outputibias.n95 outputibias.n94 94.6732
R20519 outputibias.n127 outputibias.n126 94.6732
R20520 outputibias.n11 outputibias.t5 52.3082
R20521 outputibias.n42 outputibias.t7 52.3082
R20522 outputibias.n74 outputibias.t1 52.3082
R20523 outputibias.n106 outputibias.t3 52.3082
R20524 outputibias.n12 outputibias.n10 15.6674
R20525 outputibias.n43 outputibias.n41 15.6674
R20526 outputibias.n75 outputibias.n73 15.6674
R20527 outputibias.n107 outputibias.n105 15.6674
R20528 outputibias.n13 outputibias.n9 12.8005
R20529 outputibias.n44 outputibias.n40 12.8005
R20530 outputibias.n76 outputibias.n72 12.8005
R20531 outputibias.n108 outputibias.n104 12.8005
R20532 outputibias.n17 outputibias.n16 12.0247
R20533 outputibias.n48 outputibias.n47 12.0247
R20534 outputibias.n80 outputibias.n79 12.0247
R20535 outputibias.n112 outputibias.n111 12.0247
R20536 outputibias.n20 outputibias.n7 11.249
R20537 outputibias.n51 outputibias.n38 11.249
R20538 outputibias.n83 outputibias.n70 11.249
R20539 outputibias.n115 outputibias.n102 11.249
R20540 outputibias.n21 outputibias.n5 10.4732
R20541 outputibias.n52 outputibias.n36 10.4732
R20542 outputibias.n84 outputibias.n68 10.4732
R20543 outputibias.n116 outputibias.n100 10.4732
R20544 outputibias.n25 outputibias.n24 9.69747
R20545 outputibias.n56 outputibias.n55 9.69747
R20546 outputibias.n88 outputibias.n87 9.69747
R20547 outputibias.n120 outputibias.n119 9.69747
R20548 outputibias.n31 outputibias.n30 9.45567
R20549 outputibias.n62 outputibias.n61 9.45567
R20550 outputibias.n94 outputibias.n93 9.45567
R20551 outputibias.n126 outputibias.n125 9.45567
R20552 outputibias.n30 outputibias.n29 9.3005
R20553 outputibias.n3 outputibias.n2 9.3005
R20554 outputibias.n24 outputibias.n23 9.3005
R20555 outputibias.n22 outputibias.n21 9.3005
R20556 outputibias.n7 outputibias.n6 9.3005
R20557 outputibias.n16 outputibias.n15 9.3005
R20558 outputibias.n14 outputibias.n13 9.3005
R20559 outputibias.n61 outputibias.n60 9.3005
R20560 outputibias.n34 outputibias.n33 9.3005
R20561 outputibias.n55 outputibias.n54 9.3005
R20562 outputibias.n53 outputibias.n52 9.3005
R20563 outputibias.n38 outputibias.n37 9.3005
R20564 outputibias.n47 outputibias.n46 9.3005
R20565 outputibias.n45 outputibias.n44 9.3005
R20566 outputibias.n93 outputibias.n92 9.3005
R20567 outputibias.n66 outputibias.n65 9.3005
R20568 outputibias.n87 outputibias.n86 9.3005
R20569 outputibias.n85 outputibias.n84 9.3005
R20570 outputibias.n70 outputibias.n69 9.3005
R20571 outputibias.n79 outputibias.n78 9.3005
R20572 outputibias.n77 outputibias.n76 9.3005
R20573 outputibias.n125 outputibias.n124 9.3005
R20574 outputibias.n98 outputibias.n97 9.3005
R20575 outputibias.n119 outputibias.n118 9.3005
R20576 outputibias.n117 outputibias.n116 9.3005
R20577 outputibias.n102 outputibias.n101 9.3005
R20578 outputibias.n111 outputibias.n110 9.3005
R20579 outputibias.n109 outputibias.n108 9.3005
R20580 outputibias.n28 outputibias.n3 8.92171
R20581 outputibias.n59 outputibias.n34 8.92171
R20582 outputibias.n91 outputibias.n66 8.92171
R20583 outputibias.n123 outputibias.n98 8.92171
R20584 outputibias.n29 outputibias.n1 8.14595
R20585 outputibias.n60 outputibias.n32 8.14595
R20586 outputibias.n92 outputibias.n64 8.14595
R20587 outputibias.n124 outputibias.n96 8.14595
R20588 outputibias.n31 outputibias.n1 5.81868
R20589 outputibias.n62 outputibias.n32 5.81868
R20590 outputibias.n94 outputibias.n64 5.81868
R20591 outputibias.n126 outputibias.n96 5.81868
R20592 outputibias.n131 outputibias.n130 5.20947
R20593 outputibias.n29 outputibias.n28 5.04292
R20594 outputibias.n60 outputibias.n59 5.04292
R20595 outputibias.n92 outputibias.n91 5.04292
R20596 outputibias.n124 outputibias.n123 5.04292
R20597 outputibias.n131 outputibias.n127 4.42209
R20598 outputibias.n14 outputibias.n10 4.38594
R20599 outputibias.n45 outputibias.n41 4.38594
R20600 outputibias.n77 outputibias.n73 4.38594
R20601 outputibias.n109 outputibias.n105 4.38594
R20602 outputibias.n132 outputibias.n131 4.28454
R20603 outputibias.n25 outputibias.n3 4.26717
R20604 outputibias.n56 outputibias.n34 4.26717
R20605 outputibias.n88 outputibias.n66 4.26717
R20606 outputibias.n120 outputibias.n98 4.26717
R20607 outputibias.n24 outputibias.n5 3.49141
R20608 outputibias.n55 outputibias.n36 3.49141
R20609 outputibias.n87 outputibias.n68 3.49141
R20610 outputibias.n119 outputibias.n100 3.49141
R20611 outputibias.n21 outputibias.n20 2.71565
R20612 outputibias.n52 outputibias.n51 2.71565
R20613 outputibias.n84 outputibias.n83 2.71565
R20614 outputibias.n116 outputibias.n115 2.71565
R20615 outputibias.n17 outputibias.n7 1.93989
R20616 outputibias.n48 outputibias.n38 1.93989
R20617 outputibias.n80 outputibias.n70 1.93989
R20618 outputibias.n112 outputibias.n102 1.93989
R20619 outputibias.n130 outputibias.n129 1.9266
R20620 outputibias.n129 outputibias.n128 1.9266
R20621 outputibias.n133 outputibias.n132 1.92658
R20622 outputibias.n134 outputibias.n133 1.29913
R20623 outputibias.n16 outputibias.n9 1.16414
R20624 outputibias.n47 outputibias.n40 1.16414
R20625 outputibias.n79 outputibias.n72 1.16414
R20626 outputibias.n111 outputibias.n104 1.16414
R20627 outputibias.n127 outputibias.n95 0.962709
R20628 outputibias.n95 outputibias.n63 0.962709
R20629 outputibias.n13 outputibias.n12 0.388379
R20630 outputibias.n44 outputibias.n43 0.388379
R20631 outputibias.n76 outputibias.n75 0.388379
R20632 outputibias.n108 outputibias.n107 0.388379
R20633 outputibias.n134 outputibias.n0 0.337251
R20634 outputibias outputibias.n134 0.302375
R20635 outputibias.n30 outputibias.n2 0.155672
R20636 outputibias.n23 outputibias.n2 0.155672
R20637 outputibias.n23 outputibias.n22 0.155672
R20638 outputibias.n22 outputibias.n6 0.155672
R20639 outputibias.n15 outputibias.n6 0.155672
R20640 outputibias.n15 outputibias.n14 0.155672
R20641 outputibias.n61 outputibias.n33 0.155672
R20642 outputibias.n54 outputibias.n33 0.155672
R20643 outputibias.n54 outputibias.n53 0.155672
R20644 outputibias.n53 outputibias.n37 0.155672
R20645 outputibias.n46 outputibias.n37 0.155672
R20646 outputibias.n46 outputibias.n45 0.155672
R20647 outputibias.n93 outputibias.n65 0.155672
R20648 outputibias.n86 outputibias.n65 0.155672
R20649 outputibias.n86 outputibias.n85 0.155672
R20650 outputibias.n85 outputibias.n69 0.155672
R20651 outputibias.n78 outputibias.n69 0.155672
R20652 outputibias.n78 outputibias.n77 0.155672
R20653 outputibias.n125 outputibias.n97 0.155672
R20654 outputibias.n118 outputibias.n97 0.155672
R20655 outputibias.n118 outputibias.n117 0.155672
R20656 outputibias.n117 outputibias.n101 0.155672
R20657 outputibias.n110 outputibias.n101 0.155672
R20658 outputibias.n110 outputibias.n109 0.155672
R20659 output.n41 output.n15 289.615
R20660 output.n72 output.n46 289.615
R20661 output.n104 output.n78 289.615
R20662 output.n136 output.n110 289.615
R20663 output.n77 output.n45 197.26
R20664 output.n77 output.n76 196.298
R20665 output.n109 output.n108 196.298
R20666 output.n141 output.n140 196.298
R20667 output.n42 output.n41 185
R20668 output.n40 output.n39 185
R20669 output.n19 output.n18 185
R20670 output.n34 output.n33 185
R20671 output.n32 output.n31 185
R20672 output.n23 output.n22 185
R20673 output.n26 output.n25 185
R20674 output.n73 output.n72 185
R20675 output.n71 output.n70 185
R20676 output.n50 output.n49 185
R20677 output.n65 output.n64 185
R20678 output.n63 output.n62 185
R20679 output.n54 output.n53 185
R20680 output.n57 output.n56 185
R20681 output.n105 output.n104 185
R20682 output.n103 output.n102 185
R20683 output.n82 output.n81 185
R20684 output.n97 output.n96 185
R20685 output.n95 output.n94 185
R20686 output.n86 output.n85 185
R20687 output.n89 output.n88 185
R20688 output.n137 output.n136 185
R20689 output.n135 output.n134 185
R20690 output.n114 output.n113 185
R20691 output.n129 output.n128 185
R20692 output.n127 output.n126 185
R20693 output.n118 output.n117 185
R20694 output.n121 output.n120 185
R20695 output.t3 output.n24 147.661
R20696 output.t2 output.n55 147.661
R20697 output.t1 output.n87 147.661
R20698 output.t0 output.n119 147.661
R20699 output.n41 output.n40 104.615
R20700 output.n40 output.n18 104.615
R20701 output.n33 output.n18 104.615
R20702 output.n33 output.n32 104.615
R20703 output.n32 output.n22 104.615
R20704 output.n25 output.n22 104.615
R20705 output.n72 output.n71 104.615
R20706 output.n71 output.n49 104.615
R20707 output.n64 output.n49 104.615
R20708 output.n64 output.n63 104.615
R20709 output.n63 output.n53 104.615
R20710 output.n56 output.n53 104.615
R20711 output.n104 output.n103 104.615
R20712 output.n103 output.n81 104.615
R20713 output.n96 output.n81 104.615
R20714 output.n96 output.n95 104.615
R20715 output.n95 output.n85 104.615
R20716 output.n88 output.n85 104.615
R20717 output.n136 output.n135 104.615
R20718 output.n135 output.n113 104.615
R20719 output.n128 output.n113 104.615
R20720 output.n128 output.n127 104.615
R20721 output.n127 output.n117 104.615
R20722 output.n120 output.n117 104.615
R20723 output.n1 output.t16 77.056
R20724 output.n14 output.t18 76.6694
R20725 output.n1 output.n0 72.7095
R20726 output.n3 output.n2 72.7095
R20727 output.n5 output.n4 72.7095
R20728 output.n7 output.n6 72.7095
R20729 output.n9 output.n8 72.7095
R20730 output.n11 output.n10 72.7095
R20731 output.n13 output.n12 72.7095
R20732 output.n25 output.t3 52.3082
R20733 output.n56 output.t2 52.3082
R20734 output.n88 output.t1 52.3082
R20735 output.n120 output.t0 52.3082
R20736 output.n26 output.n24 15.6674
R20737 output.n57 output.n55 15.6674
R20738 output.n89 output.n87 15.6674
R20739 output.n121 output.n119 15.6674
R20740 output.n27 output.n23 12.8005
R20741 output.n58 output.n54 12.8005
R20742 output.n90 output.n86 12.8005
R20743 output.n122 output.n118 12.8005
R20744 output.n31 output.n30 12.0247
R20745 output.n62 output.n61 12.0247
R20746 output.n94 output.n93 12.0247
R20747 output.n126 output.n125 12.0247
R20748 output.n34 output.n21 11.249
R20749 output.n65 output.n52 11.249
R20750 output.n97 output.n84 11.249
R20751 output.n129 output.n116 11.249
R20752 output.n35 output.n19 10.4732
R20753 output.n66 output.n50 10.4732
R20754 output.n98 output.n82 10.4732
R20755 output.n130 output.n114 10.4732
R20756 output.n39 output.n38 9.69747
R20757 output.n70 output.n69 9.69747
R20758 output.n102 output.n101 9.69747
R20759 output.n134 output.n133 9.69747
R20760 output.n45 output.n44 9.45567
R20761 output.n76 output.n75 9.45567
R20762 output.n108 output.n107 9.45567
R20763 output.n140 output.n139 9.45567
R20764 output.n44 output.n43 9.3005
R20765 output.n17 output.n16 9.3005
R20766 output.n38 output.n37 9.3005
R20767 output.n36 output.n35 9.3005
R20768 output.n21 output.n20 9.3005
R20769 output.n30 output.n29 9.3005
R20770 output.n28 output.n27 9.3005
R20771 output.n75 output.n74 9.3005
R20772 output.n48 output.n47 9.3005
R20773 output.n69 output.n68 9.3005
R20774 output.n67 output.n66 9.3005
R20775 output.n52 output.n51 9.3005
R20776 output.n61 output.n60 9.3005
R20777 output.n59 output.n58 9.3005
R20778 output.n107 output.n106 9.3005
R20779 output.n80 output.n79 9.3005
R20780 output.n101 output.n100 9.3005
R20781 output.n99 output.n98 9.3005
R20782 output.n84 output.n83 9.3005
R20783 output.n93 output.n92 9.3005
R20784 output.n91 output.n90 9.3005
R20785 output.n139 output.n138 9.3005
R20786 output.n112 output.n111 9.3005
R20787 output.n133 output.n132 9.3005
R20788 output.n131 output.n130 9.3005
R20789 output.n116 output.n115 9.3005
R20790 output.n125 output.n124 9.3005
R20791 output.n123 output.n122 9.3005
R20792 output.n42 output.n17 8.92171
R20793 output.n73 output.n48 8.92171
R20794 output.n105 output.n80 8.92171
R20795 output.n137 output.n112 8.92171
R20796 output output.n141 8.15037
R20797 output.n43 output.n15 8.14595
R20798 output.n74 output.n46 8.14595
R20799 output.n106 output.n78 8.14595
R20800 output.n138 output.n110 8.14595
R20801 output.n45 output.n15 5.81868
R20802 output.n76 output.n46 5.81868
R20803 output.n108 output.n78 5.81868
R20804 output.n140 output.n110 5.81868
R20805 output.n43 output.n42 5.04292
R20806 output.n74 output.n73 5.04292
R20807 output.n106 output.n105 5.04292
R20808 output.n138 output.n137 5.04292
R20809 output.n28 output.n24 4.38594
R20810 output.n59 output.n55 4.38594
R20811 output.n91 output.n87 4.38594
R20812 output.n123 output.n119 4.38594
R20813 output.n39 output.n17 4.26717
R20814 output.n70 output.n48 4.26717
R20815 output.n102 output.n80 4.26717
R20816 output.n134 output.n112 4.26717
R20817 output.n0 output.t7 3.9605
R20818 output.n0 output.t11 3.9605
R20819 output.n2 output.t14 3.9605
R20820 output.n2 output.t19 3.9605
R20821 output.n4 output.t4 3.9605
R20822 output.n4 output.t9 3.9605
R20823 output.n6 output.t13 3.9605
R20824 output.n6 output.t5 3.9605
R20825 output.n8 output.t8 3.9605
R20826 output.n8 output.t6 3.9605
R20827 output.n10 output.t12 3.9605
R20828 output.n10 output.t15 3.9605
R20829 output.n12 output.t17 3.9605
R20830 output.n12 output.t10 3.9605
R20831 output.n38 output.n19 3.49141
R20832 output.n69 output.n50 3.49141
R20833 output.n101 output.n82 3.49141
R20834 output.n133 output.n114 3.49141
R20835 output.n35 output.n34 2.71565
R20836 output.n66 output.n65 2.71565
R20837 output.n98 output.n97 2.71565
R20838 output.n130 output.n129 2.71565
R20839 output.n31 output.n21 1.93989
R20840 output.n62 output.n52 1.93989
R20841 output.n94 output.n84 1.93989
R20842 output.n126 output.n116 1.93989
R20843 output.n30 output.n23 1.16414
R20844 output.n61 output.n54 1.16414
R20845 output.n93 output.n86 1.16414
R20846 output.n125 output.n118 1.16414
R20847 output.n141 output.n109 0.962709
R20848 output.n109 output.n77 0.962709
R20849 output.n27 output.n26 0.388379
R20850 output.n58 output.n57 0.388379
R20851 output.n90 output.n89 0.388379
R20852 output.n122 output.n121 0.388379
R20853 output.n14 output.n13 0.387128
R20854 output.n13 output.n11 0.387128
R20855 output.n11 output.n9 0.387128
R20856 output.n9 output.n7 0.387128
R20857 output.n7 output.n5 0.387128
R20858 output.n5 output.n3 0.387128
R20859 output.n3 output.n1 0.387128
R20860 output.n44 output.n16 0.155672
R20861 output.n37 output.n16 0.155672
R20862 output.n37 output.n36 0.155672
R20863 output.n36 output.n20 0.155672
R20864 output.n29 output.n20 0.155672
R20865 output.n29 output.n28 0.155672
R20866 output.n75 output.n47 0.155672
R20867 output.n68 output.n47 0.155672
R20868 output.n68 output.n67 0.155672
R20869 output.n67 output.n51 0.155672
R20870 output.n60 output.n51 0.155672
R20871 output.n60 output.n59 0.155672
R20872 output.n107 output.n79 0.155672
R20873 output.n100 output.n79 0.155672
R20874 output.n100 output.n99 0.155672
R20875 output.n99 output.n83 0.155672
R20876 output.n92 output.n83 0.155672
R20877 output.n92 output.n91 0.155672
R20878 output.n139 output.n111 0.155672
R20879 output.n132 output.n111 0.155672
R20880 output.n132 output.n131 0.155672
R20881 output.n131 output.n115 0.155672
R20882 output.n124 output.n115 0.155672
R20883 output.n124 output.n123 0.155672
R20884 output output.n14 0.126227
R20885 a_n2318_8322.n8 a_n2318_8322.t3 74.6477
R20886 a_n2318_8322.n1 a_n2318_8322.t22 74.6477
R20887 a_n2318_8322.n20 a_n2318_8322.t21 74.6474
R20888 a_n2318_8322.n16 a_n2318_8322.t11 74.2899
R20889 a_n2318_8322.n9 a_n2318_8322.t1 74.2899
R20890 a_n2318_8322.n10 a_n2318_8322.t4 74.2899
R20891 a_n2318_8322.n13 a_n2318_8322.t5 74.2899
R20892 a_n2318_8322.n6 a_n2318_8322.t8 74.2899
R20893 a_n2318_8322.n20 a_n2318_8322.n19 70.6783
R20894 a_n2318_8322.n18 a_n2318_8322.n17 70.6783
R20895 a_n2318_8322.n8 a_n2318_8322.n7 70.6783
R20896 a_n2318_8322.n12 a_n2318_8322.n11 70.6783
R20897 a_n2318_8322.n1 a_n2318_8322.n0 70.6783
R20898 a_n2318_8322.n3 a_n2318_8322.n2 70.6783
R20899 a_n2318_8322.n5 a_n2318_8322.n4 70.6783
R20900 a_n2318_8322.n22 a_n2318_8322.n21 70.6782
R20901 a_n2318_8322.n14 a_n2318_8322.n6 23.4712
R20902 a_n2318_8322.n15 a_n2318_8322.t26 9.69317
R20903 a_n2318_8322.n14 a_n2318_8322.n13 6.95632
R20904 a_n2318_8322.n16 a_n2318_8322.n15 6.19447
R20905 a_n2318_8322.n15 a_n2318_8322.n14 5.3452
R20906 a_n2318_8322.n19 a_n2318_8322.t18 3.61217
R20907 a_n2318_8322.n19 a_n2318_8322.t15 3.61217
R20908 a_n2318_8322.n17 a_n2318_8322.t20 3.61217
R20909 a_n2318_8322.n17 a_n2318_8322.t12 3.61217
R20910 a_n2318_8322.n7 a_n2318_8322.t6 3.61217
R20911 a_n2318_8322.n7 a_n2318_8322.t7 3.61217
R20912 a_n2318_8322.n11 a_n2318_8322.t2 3.61217
R20913 a_n2318_8322.n11 a_n2318_8322.t0 3.61217
R20914 a_n2318_8322.n0 a_n2318_8322.t10 3.61217
R20915 a_n2318_8322.n0 a_n2318_8322.t9 3.61217
R20916 a_n2318_8322.n2 a_n2318_8322.t19 3.61217
R20917 a_n2318_8322.n2 a_n2318_8322.t14 3.61217
R20918 a_n2318_8322.n4 a_n2318_8322.t17 3.61217
R20919 a_n2318_8322.n4 a_n2318_8322.t16 3.61217
R20920 a_n2318_8322.n22 a_n2318_8322.t13 3.61217
R20921 a_n2318_8322.t23 a_n2318_8322.n22 3.61217
R20922 a_n2318_8322.n13 a_n2318_8322.n12 0.358259
R20923 a_n2318_8322.n12 a_n2318_8322.n10 0.358259
R20924 a_n2318_8322.n9 a_n2318_8322.n8 0.358259
R20925 a_n2318_8322.n6 a_n2318_8322.n5 0.358259
R20926 a_n2318_8322.n5 a_n2318_8322.n3 0.358259
R20927 a_n2318_8322.n3 a_n2318_8322.n1 0.358259
R20928 a_n2318_8322.n18 a_n2318_8322.n16 0.358259
R20929 a_n2318_8322.n21 a_n2318_8322.n18 0.358259
R20930 a_n2318_8322.n21 a_n2318_8322.n20 0.358259
R20931 a_n2318_8322.n10 a_n2318_8322.n9 0.101793
R20932 a_n2318_8322.t27 a_n2318_8322.t24 0.0788333
R20933 a_n2318_8322.t25 a_n2318_8322.t27 0.0631667
R20934 a_n2318_8322.t26 a_n2318_8322.t25 0.0471944
R20935 a_n2318_8322.t26 a_n2318_8322.t24 0.0453889
R20936 diffpairibias.n0 diffpairibias.t18 436.822
R20937 diffpairibias.n21 diffpairibias.t19 435.479
R20938 diffpairibias.n20 diffpairibias.t16 435.479
R20939 diffpairibias.n19 diffpairibias.t17 435.479
R20940 diffpairibias.n18 diffpairibias.t21 435.479
R20941 diffpairibias.n0 diffpairibias.t22 435.479
R20942 diffpairibias.n1 diffpairibias.t20 435.479
R20943 diffpairibias.n2 diffpairibias.t23 435.479
R20944 diffpairibias.n10 diffpairibias.t0 377.536
R20945 diffpairibias.n10 diffpairibias.t8 376.193
R20946 diffpairibias.n11 diffpairibias.t10 376.193
R20947 diffpairibias.n12 diffpairibias.t6 376.193
R20948 diffpairibias.n13 diffpairibias.t2 376.193
R20949 diffpairibias.n14 diffpairibias.t12 376.193
R20950 diffpairibias.n15 diffpairibias.t4 376.193
R20951 diffpairibias.n16 diffpairibias.t14 376.193
R20952 diffpairibias.n3 diffpairibias.t1 113.368
R20953 diffpairibias.n3 diffpairibias.t9 112.698
R20954 diffpairibias.n4 diffpairibias.t11 112.698
R20955 diffpairibias.n5 diffpairibias.t7 112.698
R20956 diffpairibias.n6 diffpairibias.t3 112.698
R20957 diffpairibias.n7 diffpairibias.t13 112.698
R20958 diffpairibias.n8 diffpairibias.t5 112.698
R20959 diffpairibias.n9 diffpairibias.t15 112.698
R20960 diffpairibias.n17 diffpairibias.n16 4.77242
R20961 diffpairibias.n17 diffpairibias.n9 4.30807
R20962 diffpairibias.n18 diffpairibias.n17 4.13945
R20963 diffpairibias.n16 diffpairibias.n15 1.34352
R20964 diffpairibias.n15 diffpairibias.n14 1.34352
R20965 diffpairibias.n14 diffpairibias.n13 1.34352
R20966 diffpairibias.n13 diffpairibias.n12 1.34352
R20967 diffpairibias.n12 diffpairibias.n11 1.34352
R20968 diffpairibias.n11 diffpairibias.n10 1.34352
R20969 diffpairibias.n2 diffpairibias.n1 1.34352
R20970 diffpairibias.n1 diffpairibias.n0 1.34352
R20971 diffpairibias.n19 diffpairibias.n18 1.34352
R20972 diffpairibias.n20 diffpairibias.n19 1.34352
R20973 diffpairibias.n21 diffpairibias.n20 1.34352
R20974 diffpairibias.n22 diffpairibias.n21 0.862419
R20975 diffpairibias diffpairibias.n22 0.684875
R20976 diffpairibias.n9 diffpairibias.n8 0.672012
R20977 diffpairibias.n8 diffpairibias.n7 0.672012
R20978 diffpairibias.n7 diffpairibias.n6 0.672012
R20979 diffpairibias.n6 diffpairibias.n5 0.672012
R20980 diffpairibias.n5 diffpairibias.n4 0.672012
R20981 diffpairibias.n4 diffpairibias.n3 0.672012
R20982 diffpairibias.n22 diffpairibias.n2 0.190907
C0 CSoutput output 6.13571f
C1 CSoutput outputibias 0.032386f
C2 vdd CSoutput 67.965996f
C3 commonsourceibias output 0.006808f
C4 minus diffpairibias 4.33e-19
C5 CSoutput minus 2.38478f
C6 vdd plus 0.072414f
C7 plus diffpairibias 4.56e-19
C8 commonsourceibias outputibias 0.003832f
C9 vdd commonsourceibias 0.004218f
C10 CSoutput plus 0.854911f
C11 commonsourceibias diffpairibias 0.052851f
C12 CSoutput commonsourceibias 29.0223f
C13 minus plus 9.21292f
C14 minus commonsourceibias 0.460263f
C15 plus commonsourceibias 0.41508f
C16 output outputibias 2.34152f
C17 vdd output 7.23429f
C18 diffpairibias gnd 48.96854f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.118437p
C22 plus gnd 35.013f
C23 minus gnd 27.43066f
C24 CSoutput gnd 88.48306f
C25 vdd gnd 0.379974p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 a_n2318_8322.t24 gnd 39.618103f
C74 a_n2318_8322.t26 gnd 27.7211f
C75 a_n2318_8322.t27 gnd 19.739399f
C76 a_n2318_8322.t25 gnd 39.618103f
C77 a_n2318_8322.t13 gnd 0.09582f
C78 a_n2318_8322.t22 gnd 0.89721f
C79 a_n2318_8322.t10 gnd 0.09582f
C80 a_n2318_8322.t9 gnd 0.09582f
C81 a_n2318_8322.n0 gnd 0.674956f
C82 a_n2318_8322.n1 gnd 0.754164f
C83 a_n2318_8322.t19 gnd 0.09582f
C84 a_n2318_8322.t14 gnd 0.09582f
C85 a_n2318_8322.n2 gnd 0.674956f
C86 a_n2318_8322.n3 gnd 0.383181f
C87 a_n2318_8322.t17 gnd 0.09582f
C88 a_n2318_8322.t16 gnd 0.09582f
C89 a_n2318_8322.n4 gnd 0.674956f
C90 a_n2318_8322.n5 gnd 0.383181f
C91 a_n2318_8322.t8 gnd 0.895423f
C92 a_n2318_8322.n6 gnd 1.5519f
C93 a_n2318_8322.t3 gnd 0.89721f
C94 a_n2318_8322.t6 gnd 0.09582f
C95 a_n2318_8322.t7 gnd 0.09582f
C96 a_n2318_8322.n7 gnd 0.674956f
C97 a_n2318_8322.n8 gnd 0.754164f
C98 a_n2318_8322.t1 gnd 0.895423f
C99 a_n2318_8322.n9 gnd 0.379506f
C100 a_n2318_8322.t4 gnd 0.895423f
C101 a_n2318_8322.n10 gnd 0.379506f
C102 a_n2318_8322.t2 gnd 0.09582f
C103 a_n2318_8322.t0 gnd 0.09582f
C104 a_n2318_8322.n11 gnd 0.674956f
C105 a_n2318_8322.n12 gnd 0.383181f
C106 a_n2318_8322.t5 gnd 0.895423f
C107 a_n2318_8322.n13 gnd 1.07467f
C108 a_n2318_8322.n14 gnd 1.82686f
C109 a_n2318_8322.n15 gnd 3.12946f
C110 a_n2318_8322.t11 gnd 0.895423f
C111 a_n2318_8322.n16 gnd 0.881475f
C112 a_n2318_8322.t20 gnd 0.09582f
C113 a_n2318_8322.t12 gnd 0.09582f
C114 a_n2318_8322.n17 gnd 0.674956f
C115 a_n2318_8322.n18 gnd 0.383181f
C116 a_n2318_8322.t21 gnd 0.897208f
C117 a_n2318_8322.t18 gnd 0.09582f
C118 a_n2318_8322.t15 gnd 0.09582f
C119 a_n2318_8322.n19 gnd 0.674956f
C120 a_n2318_8322.n20 gnd 0.754166f
C121 a_n2318_8322.n21 gnd 0.383179f
C122 a_n2318_8322.n22 gnd 0.674958f
C123 a_n2318_8322.t23 gnd 0.09582f
C124 output.t16 gnd 0.464308f
C125 output.t7 gnd 0.044422f
C126 output.t11 gnd 0.044422f
C127 output.n0 gnd 0.364624f
C128 output.n1 gnd 0.614102f
C129 output.t14 gnd 0.044422f
C130 output.t19 gnd 0.044422f
C131 output.n2 gnd 0.364624f
C132 output.n3 gnd 0.350265f
C133 output.t4 gnd 0.044422f
C134 output.t9 gnd 0.044422f
C135 output.n4 gnd 0.364624f
C136 output.n5 gnd 0.350265f
C137 output.t13 gnd 0.044422f
C138 output.t5 gnd 0.044422f
C139 output.n6 gnd 0.364624f
C140 output.n7 gnd 0.350265f
C141 output.t8 gnd 0.044422f
C142 output.t6 gnd 0.044422f
C143 output.n8 gnd 0.364624f
C144 output.n9 gnd 0.350265f
C145 output.t12 gnd 0.044422f
C146 output.t15 gnd 0.044422f
C147 output.n10 gnd 0.364624f
C148 output.n11 gnd 0.350265f
C149 output.t17 gnd 0.044422f
C150 output.t10 gnd 0.044422f
C151 output.n12 gnd 0.364624f
C152 output.n13 gnd 0.350265f
C153 output.t18 gnd 0.462979f
C154 output.n14 gnd 0.28994f
C155 output.n15 gnd 0.015803f
C156 output.n16 gnd 0.011243f
C157 output.n17 gnd 0.006041f
C158 output.n18 gnd 0.01428f
C159 output.n19 gnd 0.006397f
C160 output.n20 gnd 0.011243f
C161 output.n21 gnd 0.006041f
C162 output.n22 gnd 0.01428f
C163 output.n23 gnd 0.006397f
C164 output.n24 gnd 0.048111f
C165 output.t3 gnd 0.023274f
C166 output.n25 gnd 0.01071f
C167 output.n26 gnd 0.008435f
C168 output.n27 gnd 0.006041f
C169 output.n28 gnd 0.267512f
C170 output.n29 gnd 0.011243f
C171 output.n30 gnd 0.006041f
C172 output.n31 gnd 0.006397f
C173 output.n32 gnd 0.01428f
C174 output.n33 gnd 0.01428f
C175 output.n34 gnd 0.006397f
C176 output.n35 gnd 0.006041f
C177 output.n36 gnd 0.011243f
C178 output.n37 gnd 0.011243f
C179 output.n38 gnd 0.006041f
C180 output.n39 gnd 0.006397f
C181 output.n40 gnd 0.01428f
C182 output.n41 gnd 0.030913f
C183 output.n42 gnd 0.006397f
C184 output.n43 gnd 0.006041f
C185 output.n44 gnd 0.025987f
C186 output.n45 gnd 0.097665f
C187 output.n46 gnd 0.015803f
C188 output.n47 gnd 0.011243f
C189 output.n48 gnd 0.006041f
C190 output.n49 gnd 0.01428f
C191 output.n50 gnd 0.006397f
C192 output.n51 gnd 0.011243f
C193 output.n52 gnd 0.006041f
C194 output.n53 gnd 0.01428f
C195 output.n54 gnd 0.006397f
C196 output.n55 gnd 0.048111f
C197 output.t2 gnd 0.023274f
C198 output.n56 gnd 0.01071f
C199 output.n57 gnd 0.008435f
C200 output.n58 gnd 0.006041f
C201 output.n59 gnd 0.267512f
C202 output.n60 gnd 0.011243f
C203 output.n61 gnd 0.006041f
C204 output.n62 gnd 0.006397f
C205 output.n63 gnd 0.01428f
C206 output.n64 gnd 0.01428f
C207 output.n65 gnd 0.006397f
C208 output.n66 gnd 0.006041f
C209 output.n67 gnd 0.011243f
C210 output.n68 gnd 0.011243f
C211 output.n69 gnd 0.006041f
C212 output.n70 gnd 0.006397f
C213 output.n71 gnd 0.01428f
C214 output.n72 gnd 0.030913f
C215 output.n73 gnd 0.006397f
C216 output.n74 gnd 0.006041f
C217 output.n75 gnd 0.025987f
C218 output.n76 gnd 0.09306f
C219 output.n77 gnd 1.65264f
C220 output.n78 gnd 0.015803f
C221 output.n79 gnd 0.011243f
C222 output.n80 gnd 0.006041f
C223 output.n81 gnd 0.01428f
C224 output.n82 gnd 0.006397f
C225 output.n83 gnd 0.011243f
C226 output.n84 gnd 0.006041f
C227 output.n85 gnd 0.01428f
C228 output.n86 gnd 0.006397f
C229 output.n87 gnd 0.048111f
C230 output.t1 gnd 0.023274f
C231 output.n88 gnd 0.01071f
C232 output.n89 gnd 0.008435f
C233 output.n90 gnd 0.006041f
C234 output.n91 gnd 0.267512f
C235 output.n92 gnd 0.011243f
C236 output.n93 gnd 0.006041f
C237 output.n94 gnd 0.006397f
C238 output.n95 gnd 0.01428f
C239 output.n96 gnd 0.01428f
C240 output.n97 gnd 0.006397f
C241 output.n98 gnd 0.006041f
C242 output.n99 gnd 0.011243f
C243 output.n100 gnd 0.011243f
C244 output.n101 gnd 0.006041f
C245 output.n102 gnd 0.006397f
C246 output.n103 gnd 0.01428f
C247 output.n104 gnd 0.030913f
C248 output.n105 gnd 0.006397f
C249 output.n106 gnd 0.006041f
C250 output.n107 gnd 0.025987f
C251 output.n108 gnd 0.09306f
C252 output.n109 gnd 0.713089f
C253 output.n110 gnd 0.015803f
C254 output.n111 gnd 0.011243f
C255 output.n112 gnd 0.006041f
C256 output.n113 gnd 0.01428f
C257 output.n114 gnd 0.006397f
C258 output.n115 gnd 0.011243f
C259 output.n116 gnd 0.006041f
C260 output.n117 gnd 0.01428f
C261 output.n118 gnd 0.006397f
C262 output.n119 gnd 0.048111f
C263 output.t0 gnd 0.023274f
C264 output.n120 gnd 0.01071f
C265 output.n121 gnd 0.008435f
C266 output.n122 gnd 0.006041f
C267 output.n123 gnd 0.267512f
C268 output.n124 gnd 0.011243f
C269 output.n125 gnd 0.006041f
C270 output.n126 gnd 0.006397f
C271 output.n127 gnd 0.01428f
C272 output.n128 gnd 0.01428f
C273 output.n129 gnd 0.006397f
C274 output.n130 gnd 0.006041f
C275 output.n131 gnd 0.011243f
C276 output.n132 gnd 0.011243f
C277 output.n133 gnd 0.006041f
C278 output.n134 gnd 0.006397f
C279 output.n135 gnd 0.01428f
C280 output.n136 gnd 0.030913f
C281 output.n137 gnd 0.006397f
C282 output.n138 gnd 0.006041f
C283 output.n139 gnd 0.025987f
C284 output.n140 gnd 0.09306f
C285 output.n141 gnd 1.67353f
C286 outputibias.t9 gnd 0.11477f
C287 outputibias.t8 gnd 0.115567f
C288 outputibias.n0 gnd 0.130108f
C289 outputibias.n1 gnd 0.001372f
C290 outputibias.n2 gnd 9.76e-19
C291 outputibias.n3 gnd 5.24e-19
C292 outputibias.n4 gnd 0.001239f
C293 outputibias.n5 gnd 5.55e-19
C294 outputibias.n6 gnd 9.76e-19
C295 outputibias.n7 gnd 5.24e-19
C296 outputibias.n8 gnd 0.001239f
C297 outputibias.n9 gnd 5.55e-19
C298 outputibias.n10 gnd 0.004176f
C299 outputibias.t5 gnd 0.00202f
C300 outputibias.n11 gnd 9.3e-19
C301 outputibias.n12 gnd 7.32e-19
C302 outputibias.n13 gnd 5.24e-19
C303 outputibias.n14 gnd 0.02322f
C304 outputibias.n15 gnd 9.76e-19
C305 outputibias.n16 gnd 5.24e-19
C306 outputibias.n17 gnd 5.55e-19
C307 outputibias.n18 gnd 0.001239f
C308 outputibias.n19 gnd 0.001239f
C309 outputibias.n20 gnd 5.55e-19
C310 outputibias.n21 gnd 5.24e-19
C311 outputibias.n22 gnd 9.76e-19
C312 outputibias.n23 gnd 9.76e-19
C313 outputibias.n24 gnd 5.24e-19
C314 outputibias.n25 gnd 5.55e-19
C315 outputibias.n26 gnd 0.001239f
C316 outputibias.n27 gnd 0.002683f
C317 outputibias.n28 gnd 5.55e-19
C318 outputibias.n29 gnd 5.24e-19
C319 outputibias.n30 gnd 0.002256f
C320 outputibias.n31 gnd 0.005781f
C321 outputibias.n32 gnd 0.001372f
C322 outputibias.n33 gnd 9.76e-19
C323 outputibias.n34 gnd 5.24e-19
C324 outputibias.n35 gnd 0.001239f
C325 outputibias.n36 gnd 5.55e-19
C326 outputibias.n37 gnd 9.76e-19
C327 outputibias.n38 gnd 5.24e-19
C328 outputibias.n39 gnd 0.001239f
C329 outputibias.n40 gnd 5.55e-19
C330 outputibias.n41 gnd 0.004176f
C331 outputibias.t7 gnd 0.00202f
C332 outputibias.n42 gnd 9.3e-19
C333 outputibias.n43 gnd 7.32e-19
C334 outputibias.n44 gnd 5.24e-19
C335 outputibias.n45 gnd 0.02322f
C336 outputibias.n46 gnd 9.76e-19
C337 outputibias.n47 gnd 5.24e-19
C338 outputibias.n48 gnd 5.55e-19
C339 outputibias.n49 gnd 0.001239f
C340 outputibias.n50 gnd 0.001239f
C341 outputibias.n51 gnd 5.55e-19
C342 outputibias.n52 gnd 5.24e-19
C343 outputibias.n53 gnd 9.76e-19
C344 outputibias.n54 gnd 9.76e-19
C345 outputibias.n55 gnd 5.24e-19
C346 outputibias.n56 gnd 5.55e-19
C347 outputibias.n57 gnd 0.001239f
C348 outputibias.n58 gnd 0.002683f
C349 outputibias.n59 gnd 5.55e-19
C350 outputibias.n60 gnd 5.24e-19
C351 outputibias.n61 gnd 0.002256f
C352 outputibias.n62 gnd 0.005197f
C353 outputibias.n63 gnd 0.121892f
C354 outputibias.n64 gnd 0.001372f
C355 outputibias.n65 gnd 9.76e-19
C356 outputibias.n66 gnd 5.24e-19
C357 outputibias.n67 gnd 0.001239f
C358 outputibias.n68 gnd 5.55e-19
C359 outputibias.n69 gnd 9.76e-19
C360 outputibias.n70 gnd 5.24e-19
C361 outputibias.n71 gnd 0.001239f
C362 outputibias.n72 gnd 5.55e-19
C363 outputibias.n73 gnd 0.004176f
C364 outputibias.t1 gnd 0.00202f
C365 outputibias.n74 gnd 9.3e-19
C366 outputibias.n75 gnd 7.32e-19
C367 outputibias.n76 gnd 5.24e-19
C368 outputibias.n77 gnd 0.02322f
C369 outputibias.n78 gnd 9.76e-19
C370 outputibias.n79 gnd 5.24e-19
C371 outputibias.n80 gnd 5.55e-19
C372 outputibias.n81 gnd 0.001239f
C373 outputibias.n82 gnd 0.001239f
C374 outputibias.n83 gnd 5.55e-19
C375 outputibias.n84 gnd 5.24e-19
C376 outputibias.n85 gnd 9.76e-19
C377 outputibias.n86 gnd 9.76e-19
C378 outputibias.n87 gnd 5.24e-19
C379 outputibias.n88 gnd 5.55e-19
C380 outputibias.n89 gnd 0.001239f
C381 outputibias.n90 gnd 0.002683f
C382 outputibias.n91 gnd 5.55e-19
C383 outputibias.n92 gnd 5.24e-19
C384 outputibias.n93 gnd 0.002256f
C385 outputibias.n94 gnd 0.005197f
C386 outputibias.n95 gnd 0.064513f
C387 outputibias.n96 gnd 0.001372f
C388 outputibias.n97 gnd 9.76e-19
C389 outputibias.n98 gnd 5.24e-19
C390 outputibias.n99 gnd 0.001239f
C391 outputibias.n100 gnd 5.55e-19
C392 outputibias.n101 gnd 9.76e-19
C393 outputibias.n102 gnd 5.24e-19
C394 outputibias.n103 gnd 0.001239f
C395 outputibias.n104 gnd 5.55e-19
C396 outputibias.n105 gnd 0.004176f
C397 outputibias.t3 gnd 0.00202f
C398 outputibias.n106 gnd 9.3e-19
C399 outputibias.n107 gnd 7.32e-19
C400 outputibias.n108 gnd 5.24e-19
C401 outputibias.n109 gnd 0.02322f
C402 outputibias.n110 gnd 9.76e-19
C403 outputibias.n111 gnd 5.24e-19
C404 outputibias.n112 gnd 5.55e-19
C405 outputibias.n113 gnd 0.001239f
C406 outputibias.n114 gnd 0.001239f
C407 outputibias.n115 gnd 5.55e-19
C408 outputibias.n116 gnd 5.24e-19
C409 outputibias.n117 gnd 9.76e-19
C410 outputibias.n118 gnd 9.76e-19
C411 outputibias.n119 gnd 5.24e-19
C412 outputibias.n120 gnd 5.55e-19
C413 outputibias.n121 gnd 0.001239f
C414 outputibias.n122 gnd 0.002683f
C415 outputibias.n123 gnd 5.55e-19
C416 outputibias.n124 gnd 5.24e-19
C417 outputibias.n125 gnd 0.002256f
C418 outputibias.n126 gnd 0.005197f
C419 outputibias.n127 gnd 0.084814f
C420 outputibias.t2 gnd 0.108319f
C421 outputibias.t0 gnd 0.108319f
C422 outputibias.t6 gnd 0.108319f
C423 outputibias.t4 gnd 0.109238f
C424 outputibias.n128 gnd 0.134674f
C425 outputibias.n129 gnd 0.07244f
C426 outputibias.n130 gnd 0.079818f
C427 outputibias.n131 gnd 0.164901f
C428 outputibias.t11 gnd 0.11477f
C429 outputibias.n132 gnd 0.067481f
C430 outputibias.t10 gnd 0.11477f
C431 outputibias.n133 gnd 0.065115f
C432 outputibias.n134 gnd 0.029159f
C433 minus.n0 gnd 0.033059f
C434 minus.n1 gnd 0.007502f
C435 minus.n2 gnd 0.033059f
C436 minus.n3 gnd 0.007502f
C437 minus.n4 gnd 0.033059f
C438 minus.n5 gnd 0.007502f
C439 minus.n6 gnd 0.033059f
C440 minus.n7 gnd 0.007502f
C441 minus.n8 gnd 0.033059f
C442 minus.n9 gnd 0.007502f
C443 minus.t8 gnd 0.484567f
C444 minus.t7 gnd 0.467594f
C445 minus.n10 gnd 0.214486f
C446 minus.n11 gnd 0.192507f
C447 minus.n12 gnd 0.142322f
C448 minus.n13 gnd 0.033059f
C449 minus.t11 gnd 0.467594f
C450 minus.n14 gnd 0.20772f
C451 minus.n15 gnd 0.007502f
C452 minus.t10 gnd 0.467594f
C453 minus.n16 gnd 0.20772f
C454 minus.n17 gnd 0.033059f
C455 minus.n18 gnd 0.033059f
C456 minus.n19 gnd 0.033059f
C457 minus.t13 gnd 0.467594f
C458 minus.n20 gnd 0.20772f
C459 minus.n21 gnd 0.007502f
C460 minus.t20 gnd 0.467594f
C461 minus.n22 gnd 0.20772f
C462 minus.n23 gnd 0.033059f
C463 minus.n24 gnd 0.033059f
C464 minus.n25 gnd 0.033059f
C465 minus.t18 gnd 0.467594f
C466 minus.n26 gnd 0.20772f
C467 minus.n27 gnd 0.007502f
C468 minus.t25 gnd 0.467594f
C469 minus.n28 gnd 0.20772f
C470 minus.n29 gnd 0.033059f
C471 minus.n30 gnd 0.033059f
C472 minus.n31 gnd 0.033059f
C473 minus.t24 gnd 0.467594f
C474 minus.n32 gnd 0.20772f
C475 minus.n33 gnd 0.007502f
C476 minus.t14 gnd 0.467594f
C477 minus.n34 gnd 0.20772f
C478 minus.n35 gnd 0.033059f
C479 minus.n36 gnd 0.033059f
C480 minus.n37 gnd 0.033059f
C481 minus.t22 gnd 0.467594f
C482 minus.n38 gnd 0.20772f
C483 minus.n39 gnd 0.007502f
C484 minus.t19 gnd 0.467594f
C485 minus.n40 gnd 0.208026f
C486 minus.n41 gnd 0.38286f
C487 minus.n42 gnd 0.033059f
C488 minus.t12 gnd 0.467594f
C489 minus.t15 gnd 0.467594f
C490 minus.n43 gnd 0.033059f
C491 minus.t5 gnd 0.467594f
C492 minus.n44 gnd 0.20772f
C493 minus.n45 gnd 0.033059f
C494 minus.t6 gnd 0.467594f
C495 minus.t26 gnd 0.467594f
C496 minus.n46 gnd 0.20772f
C497 minus.n47 gnd 0.033059f
C498 minus.t21 gnd 0.467594f
C499 minus.t23 gnd 0.467594f
C500 minus.n48 gnd 0.20772f
C501 minus.n49 gnd 0.033059f
C502 minus.t16 gnd 0.467594f
C503 minus.t17 gnd 0.467594f
C504 minus.n50 gnd 0.20772f
C505 minus.n51 gnd 0.033059f
C506 minus.t9 gnd 0.467594f
C507 minus.t27 gnd 0.467594f
C508 minus.n52 gnd 0.214486f
C509 minus.t28 gnd 0.484567f
C510 minus.n53 gnd 0.192507f
C511 minus.n54 gnd 0.142322f
C512 minus.n55 gnd 0.007502f
C513 minus.n56 gnd 0.20772f
C514 minus.n57 gnd 0.007502f
C515 minus.n58 gnd 0.033059f
C516 minus.n59 gnd 0.033059f
C517 minus.n60 gnd 0.033059f
C518 minus.n61 gnd 0.007502f
C519 minus.n62 gnd 0.20772f
C520 minus.n63 gnd 0.007502f
C521 minus.n64 gnd 0.033059f
C522 minus.n65 gnd 0.033059f
C523 minus.n66 gnd 0.033059f
C524 minus.n67 gnd 0.007502f
C525 minus.n68 gnd 0.20772f
C526 minus.n69 gnd 0.007502f
C527 minus.n70 gnd 0.033059f
C528 minus.n71 gnd 0.033059f
C529 minus.n72 gnd 0.033059f
C530 minus.n73 gnd 0.007502f
C531 minus.n74 gnd 0.20772f
C532 minus.n75 gnd 0.007502f
C533 minus.n76 gnd 0.033059f
C534 minus.n77 gnd 0.033059f
C535 minus.n78 gnd 0.033059f
C536 minus.n79 gnd 0.007502f
C537 minus.n80 gnd 0.20772f
C538 minus.n81 gnd 0.007502f
C539 minus.n82 gnd 0.208026f
C540 minus.n83 gnd 1.10752f
C541 minus.n84 gnd 1.65019f
C542 minus.t1 gnd 0.010191f
C543 minus.t0 gnd 0.010191f
C544 minus.n85 gnd 0.033511f
C545 minus.t4 gnd 0.010191f
C546 minus.t3 gnd 0.010191f
C547 minus.n86 gnd 0.033052f
C548 minus.n87 gnd 0.282084f
C549 minus.t2 gnd 0.056723f
C550 minus.n88 gnd 0.15393f
C551 minus.n89 gnd 1.77478f
C552 commonsourceibias.n0 gnd 0.010301f
C553 commonsourceibias.t71 gnd 0.155981f
C554 commonsourceibias.t81 gnd 0.144227f
C555 commonsourceibias.n1 gnd 0.057546f
C556 commonsourceibias.n2 gnd 0.00772f
C557 commonsourceibias.t55 gnd 0.144227f
C558 commonsourceibias.n3 gnd 0.006245f
C559 commonsourceibias.n4 gnd 0.00772f
C560 commonsourceibias.t53 gnd 0.144227f
C561 commonsourceibias.n5 gnd 0.007453f
C562 commonsourceibias.n6 gnd 0.00772f
C563 commonsourceibias.t76 gnd 0.144227f
C564 commonsourceibias.n7 gnd 0.057546f
C565 commonsourceibias.t86 gnd 0.144227f
C566 commonsourceibias.n8 gnd 0.006235f
C567 commonsourceibias.n9 gnd 0.010301f
C568 commonsourceibias.t32 gnd 0.155981f
C569 commonsourceibias.t14 gnd 0.144227f
C570 commonsourceibias.n10 gnd 0.057546f
C571 commonsourceibias.n11 gnd 0.00772f
C572 commonsourceibias.t24 gnd 0.144227f
C573 commonsourceibias.n12 gnd 0.006245f
C574 commonsourceibias.n13 gnd 0.00772f
C575 commonsourceibias.t30 gnd 0.144227f
C576 commonsourceibias.n14 gnd 0.007453f
C577 commonsourceibias.n15 gnd 0.00772f
C578 commonsourceibias.t20 gnd 0.144227f
C579 commonsourceibias.n16 gnd 0.057546f
C580 commonsourceibias.t36 gnd 0.144227f
C581 commonsourceibias.n17 gnd 0.006235f
C582 commonsourceibias.n18 gnd 0.00772f
C583 commonsourceibias.t44 gnd 0.144227f
C584 commonsourceibias.t26 gnd 0.144227f
C585 commonsourceibias.n19 gnd 0.057546f
C586 commonsourceibias.n20 gnd 0.00772f
C587 commonsourceibias.t34 gnd 0.144227f
C588 commonsourceibias.n21 gnd 0.057546f
C589 commonsourceibias.n22 gnd 0.00772f
C590 commonsourceibias.t10 gnd 0.144227f
C591 commonsourceibias.n23 gnd 0.057546f
C592 commonsourceibias.n24 gnd 0.038863f
C593 commonsourceibias.t40 gnd 0.144227f
C594 commonsourceibias.t46 gnd 0.162743f
C595 commonsourceibias.n25 gnd 0.066782f
C596 commonsourceibias.n26 gnd 0.069137f
C597 commonsourceibias.n27 gnd 0.009515f
C598 commonsourceibias.n28 gnd 0.010526f
C599 commonsourceibias.n29 gnd 0.00772f
C600 commonsourceibias.n30 gnd 0.00772f
C601 commonsourceibias.n31 gnd 0.010457f
C602 commonsourceibias.n32 gnd 0.006245f
C603 commonsourceibias.n33 gnd 0.010587f
C604 commonsourceibias.n34 gnd 0.00772f
C605 commonsourceibias.n35 gnd 0.00772f
C606 commonsourceibias.n36 gnd 0.010651f
C607 commonsourceibias.n37 gnd 0.009185f
C608 commonsourceibias.n38 gnd 0.007453f
C609 commonsourceibias.n39 gnd 0.00772f
C610 commonsourceibias.n40 gnd 0.00772f
C611 commonsourceibias.n41 gnd 0.009442f
C612 commonsourceibias.n42 gnd 0.010598f
C613 commonsourceibias.n43 gnd 0.057546f
C614 commonsourceibias.n44 gnd 0.010527f
C615 commonsourceibias.n45 gnd 0.00772f
C616 commonsourceibias.n46 gnd 0.00772f
C617 commonsourceibias.n47 gnd 0.00772f
C618 commonsourceibias.n48 gnd 0.010527f
C619 commonsourceibias.n49 gnd 0.057546f
C620 commonsourceibias.n50 gnd 0.010598f
C621 commonsourceibias.n51 gnd 0.009442f
C622 commonsourceibias.n52 gnd 0.00772f
C623 commonsourceibias.n53 gnd 0.00772f
C624 commonsourceibias.n54 gnd 0.00772f
C625 commonsourceibias.n55 gnd 0.009185f
C626 commonsourceibias.n56 gnd 0.010651f
C627 commonsourceibias.n57 gnd 0.057546f
C628 commonsourceibias.n58 gnd 0.010587f
C629 commonsourceibias.n59 gnd 0.00772f
C630 commonsourceibias.n60 gnd 0.00772f
C631 commonsourceibias.n61 gnd 0.00772f
C632 commonsourceibias.n62 gnd 0.010457f
C633 commonsourceibias.n63 gnd 0.057546f
C634 commonsourceibias.n64 gnd 0.010526f
C635 commonsourceibias.n65 gnd 0.009515f
C636 commonsourceibias.n66 gnd 0.00772f
C637 commonsourceibias.n67 gnd 0.00772f
C638 commonsourceibias.n68 gnd 0.007831f
C639 commonsourceibias.n69 gnd 0.008096f
C640 commonsourceibias.n70 gnd 0.068855f
C641 commonsourceibias.n71 gnd 0.076384f
C642 commonsourceibias.t33 gnd 0.016658f
C643 commonsourceibias.t15 gnd 0.016658f
C644 commonsourceibias.n72 gnd 0.147197f
C645 commonsourceibias.n73 gnd 0.12719f
C646 commonsourceibias.t25 gnd 0.016658f
C647 commonsourceibias.t31 gnd 0.016658f
C648 commonsourceibias.n74 gnd 0.147197f
C649 commonsourceibias.n75 gnd 0.067614f
C650 commonsourceibias.t21 gnd 0.016658f
C651 commonsourceibias.t37 gnd 0.016658f
C652 commonsourceibias.n76 gnd 0.147197f
C653 commonsourceibias.n77 gnd 0.056488f
C654 commonsourceibias.t41 gnd 0.016658f
C655 commonsourceibias.t47 gnd 0.016658f
C656 commonsourceibias.n78 gnd 0.14769f
C657 commonsourceibias.t35 gnd 0.016658f
C658 commonsourceibias.t11 gnd 0.016658f
C659 commonsourceibias.n79 gnd 0.147197f
C660 commonsourceibias.n80 gnd 0.13716f
C661 commonsourceibias.t45 gnd 0.016658f
C662 commonsourceibias.t27 gnd 0.016658f
C663 commonsourceibias.n81 gnd 0.147197f
C664 commonsourceibias.n82 gnd 0.056488f
C665 commonsourceibias.n83 gnd 0.068401f
C666 commonsourceibias.n84 gnd 0.00772f
C667 commonsourceibias.t50 gnd 0.144227f
C668 commonsourceibias.t69 gnd 0.144227f
C669 commonsourceibias.n85 gnd 0.057546f
C670 commonsourceibias.n86 gnd 0.00772f
C671 commonsourceibias.t67 gnd 0.144227f
C672 commonsourceibias.n87 gnd 0.057546f
C673 commonsourceibias.n88 gnd 0.00772f
C674 commonsourceibias.t78 gnd 0.144227f
C675 commonsourceibias.n89 gnd 0.057546f
C676 commonsourceibias.n90 gnd 0.038863f
C677 commonsourceibias.t64 gnd 0.144227f
C678 commonsourceibias.t62 gnd 0.162743f
C679 commonsourceibias.n91 gnd 0.066782f
C680 commonsourceibias.n92 gnd 0.069137f
C681 commonsourceibias.n93 gnd 0.009515f
C682 commonsourceibias.n94 gnd 0.010526f
C683 commonsourceibias.n95 gnd 0.00772f
C684 commonsourceibias.n96 gnd 0.00772f
C685 commonsourceibias.n97 gnd 0.010457f
C686 commonsourceibias.n98 gnd 0.006245f
C687 commonsourceibias.n99 gnd 0.010587f
C688 commonsourceibias.n100 gnd 0.00772f
C689 commonsourceibias.n101 gnd 0.00772f
C690 commonsourceibias.n102 gnd 0.010651f
C691 commonsourceibias.n103 gnd 0.009185f
C692 commonsourceibias.n104 gnd 0.007453f
C693 commonsourceibias.n105 gnd 0.00772f
C694 commonsourceibias.n106 gnd 0.00772f
C695 commonsourceibias.n107 gnd 0.009442f
C696 commonsourceibias.n108 gnd 0.010598f
C697 commonsourceibias.n109 gnd 0.057546f
C698 commonsourceibias.n110 gnd 0.010527f
C699 commonsourceibias.n111 gnd 0.007683f
C700 commonsourceibias.n112 gnd 0.055804f
C701 commonsourceibias.n113 gnd 0.007683f
C702 commonsourceibias.n114 gnd 0.010527f
C703 commonsourceibias.n115 gnd 0.057546f
C704 commonsourceibias.n116 gnd 0.010598f
C705 commonsourceibias.n117 gnd 0.009442f
C706 commonsourceibias.n118 gnd 0.00772f
C707 commonsourceibias.n119 gnd 0.00772f
C708 commonsourceibias.n120 gnd 0.00772f
C709 commonsourceibias.n121 gnd 0.009185f
C710 commonsourceibias.n122 gnd 0.010651f
C711 commonsourceibias.n123 gnd 0.057546f
C712 commonsourceibias.n124 gnd 0.010587f
C713 commonsourceibias.n125 gnd 0.00772f
C714 commonsourceibias.n126 gnd 0.00772f
C715 commonsourceibias.n127 gnd 0.00772f
C716 commonsourceibias.n128 gnd 0.010457f
C717 commonsourceibias.n129 gnd 0.057546f
C718 commonsourceibias.n130 gnd 0.010526f
C719 commonsourceibias.n131 gnd 0.009515f
C720 commonsourceibias.n132 gnd 0.00772f
C721 commonsourceibias.n133 gnd 0.00772f
C722 commonsourceibias.n134 gnd 0.007831f
C723 commonsourceibias.n135 gnd 0.008096f
C724 commonsourceibias.n136 gnd 0.068855f
C725 commonsourceibias.n137 gnd 0.04456f
C726 commonsourceibias.n138 gnd 0.010301f
C727 commonsourceibias.t72 gnd 0.144227f
C728 commonsourceibias.n139 gnd 0.057546f
C729 commonsourceibias.n140 gnd 0.00772f
C730 commonsourceibias.t49 gnd 0.144227f
C731 commonsourceibias.n141 gnd 0.006245f
C732 commonsourceibias.n142 gnd 0.00772f
C733 commonsourceibias.t95 gnd 0.144227f
C734 commonsourceibias.n143 gnd 0.007453f
C735 commonsourceibias.n144 gnd 0.00772f
C736 commonsourceibias.t66 gnd 0.144227f
C737 commonsourceibias.n145 gnd 0.057546f
C738 commonsourceibias.t77 gnd 0.144227f
C739 commonsourceibias.n146 gnd 0.006235f
C740 commonsourceibias.n147 gnd 0.00772f
C741 commonsourceibias.t91 gnd 0.144227f
C742 commonsourceibias.t60 gnd 0.144227f
C743 commonsourceibias.n148 gnd 0.057546f
C744 commonsourceibias.n149 gnd 0.00772f
C745 commonsourceibias.t58 gnd 0.144227f
C746 commonsourceibias.n150 gnd 0.057546f
C747 commonsourceibias.n151 gnd 0.00772f
C748 commonsourceibias.t68 gnd 0.144227f
C749 commonsourceibias.n152 gnd 0.057546f
C750 commonsourceibias.n153 gnd 0.038863f
C751 commonsourceibias.t57 gnd 0.144227f
C752 commonsourceibias.t54 gnd 0.162743f
C753 commonsourceibias.n154 gnd 0.066782f
C754 commonsourceibias.n155 gnd 0.069137f
C755 commonsourceibias.n156 gnd 0.009515f
C756 commonsourceibias.n157 gnd 0.010526f
C757 commonsourceibias.n158 gnd 0.00772f
C758 commonsourceibias.n159 gnd 0.00772f
C759 commonsourceibias.n160 gnd 0.010457f
C760 commonsourceibias.n161 gnd 0.006245f
C761 commonsourceibias.n162 gnd 0.010587f
C762 commonsourceibias.n163 gnd 0.00772f
C763 commonsourceibias.n164 gnd 0.00772f
C764 commonsourceibias.n165 gnd 0.010651f
C765 commonsourceibias.n166 gnd 0.009185f
C766 commonsourceibias.n167 gnd 0.007453f
C767 commonsourceibias.n168 gnd 0.00772f
C768 commonsourceibias.n169 gnd 0.00772f
C769 commonsourceibias.n170 gnd 0.009442f
C770 commonsourceibias.n171 gnd 0.010598f
C771 commonsourceibias.n172 gnd 0.057546f
C772 commonsourceibias.n173 gnd 0.010527f
C773 commonsourceibias.n174 gnd 0.00772f
C774 commonsourceibias.n175 gnd 0.00772f
C775 commonsourceibias.n176 gnd 0.00772f
C776 commonsourceibias.n177 gnd 0.010527f
C777 commonsourceibias.n178 gnd 0.057546f
C778 commonsourceibias.n179 gnd 0.010598f
C779 commonsourceibias.n180 gnd 0.009442f
C780 commonsourceibias.n181 gnd 0.00772f
C781 commonsourceibias.n182 gnd 0.00772f
C782 commonsourceibias.n183 gnd 0.00772f
C783 commonsourceibias.n184 gnd 0.009185f
C784 commonsourceibias.n185 gnd 0.010651f
C785 commonsourceibias.n186 gnd 0.057546f
C786 commonsourceibias.n187 gnd 0.010587f
C787 commonsourceibias.n188 gnd 0.00772f
C788 commonsourceibias.n189 gnd 0.00772f
C789 commonsourceibias.n190 gnd 0.00772f
C790 commonsourceibias.n191 gnd 0.010457f
C791 commonsourceibias.n192 gnd 0.057546f
C792 commonsourceibias.n193 gnd 0.010526f
C793 commonsourceibias.n194 gnd 0.009515f
C794 commonsourceibias.n195 gnd 0.00772f
C795 commonsourceibias.n196 gnd 0.00772f
C796 commonsourceibias.n197 gnd 0.007831f
C797 commonsourceibias.n198 gnd 0.008096f
C798 commonsourceibias.t61 gnd 0.155981f
C799 commonsourceibias.n199 gnd 0.068855f
C800 commonsourceibias.n200 gnd 0.023432f
C801 commonsourceibias.n201 gnd 0.388694f
C802 commonsourceibias.n202 gnd 0.010301f
C803 commonsourceibias.t84 gnd 0.155981f
C804 commonsourceibias.t92 gnd 0.144227f
C805 commonsourceibias.n203 gnd 0.057546f
C806 commonsourceibias.n204 gnd 0.00772f
C807 commonsourceibias.t51 gnd 0.144227f
C808 commonsourceibias.n205 gnd 0.006245f
C809 commonsourceibias.n206 gnd 0.00772f
C810 commonsourceibias.t63 gnd 0.144227f
C811 commonsourceibias.n207 gnd 0.007453f
C812 commonsourceibias.n208 gnd 0.00772f
C813 commonsourceibias.t48 gnd 0.144227f
C814 commonsourceibias.n209 gnd 0.006235f
C815 commonsourceibias.n210 gnd 0.00772f
C816 commonsourceibias.t94 gnd 0.144227f
C817 commonsourceibias.t83 gnd 0.144227f
C818 commonsourceibias.n211 gnd 0.057546f
C819 commonsourceibias.n212 gnd 0.00772f
C820 commonsourceibias.t80 gnd 0.144227f
C821 commonsourceibias.n213 gnd 0.057546f
C822 commonsourceibias.n214 gnd 0.00772f
C823 commonsourceibias.t90 gnd 0.144227f
C824 commonsourceibias.n215 gnd 0.057546f
C825 commonsourceibias.n216 gnd 0.038863f
C826 commonsourceibias.t59 gnd 0.144227f
C827 commonsourceibias.t75 gnd 0.162743f
C828 commonsourceibias.n217 gnd 0.066782f
C829 commonsourceibias.n218 gnd 0.069137f
C830 commonsourceibias.n219 gnd 0.009515f
C831 commonsourceibias.n220 gnd 0.010526f
C832 commonsourceibias.n221 gnd 0.00772f
C833 commonsourceibias.n222 gnd 0.00772f
C834 commonsourceibias.n223 gnd 0.010457f
C835 commonsourceibias.n224 gnd 0.006245f
C836 commonsourceibias.n225 gnd 0.010587f
C837 commonsourceibias.n226 gnd 0.00772f
C838 commonsourceibias.n227 gnd 0.00772f
C839 commonsourceibias.n228 gnd 0.010651f
C840 commonsourceibias.n229 gnd 0.009185f
C841 commonsourceibias.n230 gnd 0.007453f
C842 commonsourceibias.n231 gnd 0.00772f
C843 commonsourceibias.n232 gnd 0.00772f
C844 commonsourceibias.n233 gnd 0.009442f
C845 commonsourceibias.n234 gnd 0.010598f
C846 commonsourceibias.n235 gnd 0.057546f
C847 commonsourceibias.n236 gnd 0.010527f
C848 commonsourceibias.n237 gnd 0.007683f
C849 commonsourceibias.t17 gnd 0.016658f
C850 commonsourceibias.t9 gnd 0.016658f
C851 commonsourceibias.n238 gnd 0.14769f
C852 commonsourceibias.t19 gnd 0.016658f
C853 commonsourceibias.t5 gnd 0.016658f
C854 commonsourceibias.n239 gnd 0.147197f
C855 commonsourceibias.n240 gnd 0.13716f
C856 commonsourceibias.t43 gnd 0.016658f
C857 commonsourceibias.t13 gnd 0.016658f
C858 commonsourceibias.n241 gnd 0.147197f
C859 commonsourceibias.n242 gnd 0.056488f
C860 commonsourceibias.n243 gnd 0.010301f
C861 commonsourceibias.t22 gnd 0.144227f
C862 commonsourceibias.n244 gnd 0.057546f
C863 commonsourceibias.n245 gnd 0.00772f
C864 commonsourceibias.t38 gnd 0.144227f
C865 commonsourceibias.n246 gnd 0.006245f
C866 commonsourceibias.n247 gnd 0.00772f
C867 commonsourceibias.t0 gnd 0.144227f
C868 commonsourceibias.n248 gnd 0.007453f
C869 commonsourceibias.n249 gnd 0.00772f
C870 commonsourceibias.t6 gnd 0.144227f
C871 commonsourceibias.n250 gnd 0.006235f
C872 commonsourceibias.n251 gnd 0.00772f
C873 commonsourceibias.t12 gnd 0.144227f
C874 commonsourceibias.t42 gnd 0.144227f
C875 commonsourceibias.n252 gnd 0.057546f
C876 commonsourceibias.n253 gnd 0.00772f
C877 commonsourceibias.t4 gnd 0.144227f
C878 commonsourceibias.n254 gnd 0.057546f
C879 commonsourceibias.n255 gnd 0.00772f
C880 commonsourceibias.t18 gnd 0.144227f
C881 commonsourceibias.n256 gnd 0.057546f
C882 commonsourceibias.n257 gnd 0.038863f
C883 commonsourceibias.t8 gnd 0.144227f
C884 commonsourceibias.t16 gnd 0.162743f
C885 commonsourceibias.n258 gnd 0.066782f
C886 commonsourceibias.n259 gnd 0.069137f
C887 commonsourceibias.n260 gnd 0.009515f
C888 commonsourceibias.n261 gnd 0.010526f
C889 commonsourceibias.n262 gnd 0.00772f
C890 commonsourceibias.n263 gnd 0.00772f
C891 commonsourceibias.n264 gnd 0.010457f
C892 commonsourceibias.n265 gnd 0.006245f
C893 commonsourceibias.n266 gnd 0.010587f
C894 commonsourceibias.n267 gnd 0.00772f
C895 commonsourceibias.n268 gnd 0.00772f
C896 commonsourceibias.n269 gnd 0.010651f
C897 commonsourceibias.n270 gnd 0.009185f
C898 commonsourceibias.n271 gnd 0.007453f
C899 commonsourceibias.n272 gnd 0.00772f
C900 commonsourceibias.n273 gnd 0.00772f
C901 commonsourceibias.n274 gnd 0.009442f
C902 commonsourceibias.n275 gnd 0.010598f
C903 commonsourceibias.n276 gnd 0.057546f
C904 commonsourceibias.n277 gnd 0.010527f
C905 commonsourceibias.n278 gnd 0.00772f
C906 commonsourceibias.n279 gnd 0.00772f
C907 commonsourceibias.n280 gnd 0.00772f
C908 commonsourceibias.n281 gnd 0.010527f
C909 commonsourceibias.n282 gnd 0.057546f
C910 commonsourceibias.n283 gnd 0.010598f
C911 commonsourceibias.t28 gnd 0.144227f
C912 commonsourceibias.n284 gnd 0.057546f
C913 commonsourceibias.n285 gnd 0.009442f
C914 commonsourceibias.n286 gnd 0.00772f
C915 commonsourceibias.n287 gnd 0.00772f
C916 commonsourceibias.n288 gnd 0.00772f
C917 commonsourceibias.n289 gnd 0.009185f
C918 commonsourceibias.n290 gnd 0.010651f
C919 commonsourceibias.n291 gnd 0.057546f
C920 commonsourceibias.n292 gnd 0.010587f
C921 commonsourceibias.n293 gnd 0.00772f
C922 commonsourceibias.n294 gnd 0.00772f
C923 commonsourceibias.n295 gnd 0.00772f
C924 commonsourceibias.n296 gnd 0.010457f
C925 commonsourceibias.n297 gnd 0.057546f
C926 commonsourceibias.n298 gnd 0.010526f
C927 commonsourceibias.n299 gnd 0.009515f
C928 commonsourceibias.n300 gnd 0.00772f
C929 commonsourceibias.n301 gnd 0.00772f
C930 commonsourceibias.n302 gnd 0.007831f
C931 commonsourceibias.n303 gnd 0.008096f
C932 commonsourceibias.t2 gnd 0.155981f
C933 commonsourceibias.n304 gnd 0.068855f
C934 commonsourceibias.n305 gnd 0.076384f
C935 commonsourceibias.t23 gnd 0.016658f
C936 commonsourceibias.t3 gnd 0.016658f
C937 commonsourceibias.n306 gnd 0.147197f
C938 commonsourceibias.n307 gnd 0.12719f
C939 commonsourceibias.t1 gnd 0.016658f
C940 commonsourceibias.t39 gnd 0.016658f
C941 commonsourceibias.n308 gnd 0.147197f
C942 commonsourceibias.n309 gnd 0.067614f
C943 commonsourceibias.t7 gnd 0.016658f
C944 commonsourceibias.t29 gnd 0.016658f
C945 commonsourceibias.n310 gnd 0.147197f
C946 commonsourceibias.n311 gnd 0.056488f
C947 commonsourceibias.n312 gnd 0.068401f
C948 commonsourceibias.n313 gnd 0.055804f
C949 commonsourceibias.n314 gnd 0.007683f
C950 commonsourceibias.n315 gnd 0.010527f
C951 commonsourceibias.n316 gnd 0.057546f
C952 commonsourceibias.n317 gnd 0.010598f
C953 commonsourceibias.t88 gnd 0.144227f
C954 commonsourceibias.n318 gnd 0.057546f
C955 commonsourceibias.n319 gnd 0.009442f
C956 commonsourceibias.n320 gnd 0.00772f
C957 commonsourceibias.n321 gnd 0.00772f
C958 commonsourceibias.n322 gnd 0.00772f
C959 commonsourceibias.n323 gnd 0.009185f
C960 commonsourceibias.n324 gnd 0.010651f
C961 commonsourceibias.n325 gnd 0.057546f
C962 commonsourceibias.n326 gnd 0.010587f
C963 commonsourceibias.n327 gnd 0.00772f
C964 commonsourceibias.n328 gnd 0.00772f
C965 commonsourceibias.n329 gnd 0.00772f
C966 commonsourceibias.n330 gnd 0.010457f
C967 commonsourceibias.n331 gnd 0.057546f
C968 commonsourceibias.n332 gnd 0.010526f
C969 commonsourceibias.n333 gnd 0.009515f
C970 commonsourceibias.n334 gnd 0.00772f
C971 commonsourceibias.n335 gnd 0.00772f
C972 commonsourceibias.n336 gnd 0.007831f
C973 commonsourceibias.n337 gnd 0.008096f
C974 commonsourceibias.n338 gnd 0.068855f
C975 commonsourceibias.n339 gnd 0.04456f
C976 commonsourceibias.n340 gnd 0.010301f
C977 commonsourceibias.t85 gnd 0.144227f
C978 commonsourceibias.n341 gnd 0.057546f
C979 commonsourceibias.n342 gnd 0.00772f
C980 commonsourceibias.t93 gnd 0.144227f
C981 commonsourceibias.n343 gnd 0.006245f
C982 commonsourceibias.n344 gnd 0.00772f
C983 commonsourceibias.t56 gnd 0.144227f
C984 commonsourceibias.n345 gnd 0.007453f
C985 commonsourceibias.n346 gnd 0.00772f
C986 commonsourceibias.t89 gnd 0.144227f
C987 commonsourceibias.n347 gnd 0.006235f
C988 commonsourceibias.n348 gnd 0.00772f
C989 commonsourceibias.t87 gnd 0.144227f
C990 commonsourceibias.t74 gnd 0.144227f
C991 commonsourceibias.n349 gnd 0.057546f
C992 commonsourceibias.n350 gnd 0.00772f
C993 commonsourceibias.t70 gnd 0.144227f
C994 commonsourceibias.n351 gnd 0.057546f
C995 commonsourceibias.n352 gnd 0.00772f
C996 commonsourceibias.t82 gnd 0.144227f
C997 commonsourceibias.n353 gnd 0.057546f
C998 commonsourceibias.n354 gnd 0.038863f
C999 commonsourceibias.t52 gnd 0.144227f
C1000 commonsourceibias.t65 gnd 0.162743f
C1001 commonsourceibias.n355 gnd 0.066782f
C1002 commonsourceibias.n356 gnd 0.069137f
C1003 commonsourceibias.n357 gnd 0.009515f
C1004 commonsourceibias.n358 gnd 0.010526f
C1005 commonsourceibias.n359 gnd 0.00772f
C1006 commonsourceibias.n360 gnd 0.00772f
C1007 commonsourceibias.n361 gnd 0.010457f
C1008 commonsourceibias.n362 gnd 0.006245f
C1009 commonsourceibias.n363 gnd 0.010587f
C1010 commonsourceibias.n364 gnd 0.00772f
C1011 commonsourceibias.n365 gnd 0.00772f
C1012 commonsourceibias.n366 gnd 0.010651f
C1013 commonsourceibias.n367 gnd 0.009185f
C1014 commonsourceibias.n368 gnd 0.007453f
C1015 commonsourceibias.n369 gnd 0.00772f
C1016 commonsourceibias.n370 gnd 0.00772f
C1017 commonsourceibias.n371 gnd 0.009442f
C1018 commonsourceibias.n372 gnd 0.010598f
C1019 commonsourceibias.n373 gnd 0.057546f
C1020 commonsourceibias.n374 gnd 0.010527f
C1021 commonsourceibias.n375 gnd 0.00772f
C1022 commonsourceibias.n376 gnd 0.00772f
C1023 commonsourceibias.n377 gnd 0.00772f
C1024 commonsourceibias.n378 gnd 0.010527f
C1025 commonsourceibias.n379 gnd 0.057546f
C1026 commonsourceibias.n380 gnd 0.010598f
C1027 commonsourceibias.t79 gnd 0.144227f
C1028 commonsourceibias.n381 gnd 0.057546f
C1029 commonsourceibias.n382 gnd 0.009442f
C1030 commonsourceibias.n383 gnd 0.00772f
C1031 commonsourceibias.n384 gnd 0.00772f
C1032 commonsourceibias.n385 gnd 0.00772f
C1033 commonsourceibias.n386 gnd 0.009185f
C1034 commonsourceibias.n387 gnd 0.010651f
C1035 commonsourceibias.n388 gnd 0.057546f
C1036 commonsourceibias.n389 gnd 0.010587f
C1037 commonsourceibias.n390 gnd 0.00772f
C1038 commonsourceibias.n391 gnd 0.00772f
C1039 commonsourceibias.n392 gnd 0.00772f
C1040 commonsourceibias.n393 gnd 0.010457f
C1041 commonsourceibias.n394 gnd 0.057546f
C1042 commonsourceibias.n395 gnd 0.010526f
C1043 commonsourceibias.n396 gnd 0.009515f
C1044 commonsourceibias.n397 gnd 0.00772f
C1045 commonsourceibias.n398 gnd 0.00772f
C1046 commonsourceibias.n399 gnd 0.007831f
C1047 commonsourceibias.n400 gnd 0.008096f
C1048 commonsourceibias.t73 gnd 0.155981f
C1049 commonsourceibias.n401 gnd 0.068855f
C1050 commonsourceibias.n402 gnd 0.023432f
C1051 commonsourceibias.n403 gnd 0.212991f
C1052 commonsourceibias.n404 gnd 4.01312f
C1053 a_n2903_n3924.t18 gnd 0.102925f
C1054 a_n2903_n3924.t24 gnd 0.102925f
C1055 a_n2903_n3924.n0 gnd 0.840607f
C1056 a_n2903_n3924.n1 gnd 0.382272f
C1057 a_n2903_n3924.t27 gnd 1.06972f
C1058 a_n2903_n3924.n2 gnd 0.962269f
C1059 a_n2903_n3924.t7 gnd 0.102925f
C1060 a_n2903_n3924.t25 gnd 0.102925f
C1061 a_n2903_n3924.n3 gnd 0.840609f
C1062 a_n2903_n3924.n4 gnd 0.382271f
C1063 a_n2903_n3924.t21 gnd 0.102925f
C1064 a_n2903_n3924.t23 gnd 0.102925f
C1065 a_n2903_n3924.n5 gnd 0.840609f
C1066 a_n2903_n3924.n6 gnd 0.382271f
C1067 a_n2903_n3924.t26 gnd 0.102925f
C1068 a_n2903_n3924.t28 gnd 0.102925f
C1069 a_n2903_n3924.n7 gnd 0.840609f
C1070 a_n2903_n3924.n8 gnd 0.382271f
C1071 a_n2903_n3924.t10 gnd 0.102925f
C1072 a_n2903_n3924.t8 gnd 0.102925f
C1073 a_n2903_n3924.n9 gnd 0.840609f
C1074 a_n2903_n3924.n10 gnd 0.382271f
C1075 a_n2903_n3924.t16 gnd 0.102925f
C1076 a_n2903_n3924.t9 gnd 0.102925f
C1077 a_n2903_n3924.n11 gnd 0.840609f
C1078 a_n2903_n3924.n12 gnd 0.382271f
C1079 a_n2903_n3924.t15 gnd 1.06972f
C1080 a_n2903_n3924.n13 gnd 0.383728f
C1081 a_n2903_n3924.t49 gnd 1.06972f
C1082 a_n2903_n3924.n14 gnd 0.383728f
C1083 a_n2903_n3924.t31 gnd 0.102925f
C1084 a_n2903_n3924.t50 gnd 0.102925f
C1085 a_n2903_n3924.n15 gnd 0.840609f
C1086 a_n2903_n3924.n16 gnd 0.382271f
C1087 a_n2903_n3924.t46 gnd 0.102925f
C1088 a_n2903_n3924.t3 gnd 0.102925f
C1089 a_n2903_n3924.n17 gnd 0.840609f
C1090 a_n2903_n3924.n18 gnd 0.382271f
C1091 a_n2903_n3924.t43 gnd 0.102925f
C1092 a_n2903_n3924.t42 gnd 0.102925f
C1093 a_n2903_n3924.n19 gnd 0.840609f
C1094 a_n2903_n3924.n20 gnd 0.382271f
C1095 a_n2903_n3924.t0 gnd 0.102925f
C1096 a_n2903_n3924.t54 gnd 0.102925f
C1097 a_n2903_n3924.n21 gnd 0.840609f
C1098 a_n2903_n3924.n22 gnd 0.382271f
C1099 a_n2903_n3924.t45 gnd 0.102925f
C1100 a_n2903_n3924.t35 gnd 0.102925f
C1101 a_n2903_n3924.n23 gnd 0.840609f
C1102 a_n2903_n3924.n24 gnd 0.382271f
C1103 a_n2903_n3924.t40 gnd 1.06972f
C1104 a_n2903_n3924.n25 gnd 0.962265f
C1105 a_n2903_n3924.t13 gnd 0.102925f
C1106 a_n2903_n3924.t19 gnd 0.102925f
C1107 a_n2903_n3924.n26 gnd 0.840607f
C1108 a_n2903_n3924.n27 gnd 0.382272f
C1109 a_n2903_n3924.t14 gnd 1.06972f
C1110 a_n2903_n3924.n28 gnd 0.625684f
C1111 a_n2903_n3924.n29 gnd 0.965474f
C1112 a_n2903_n3924.t37 gnd 1.32974f
C1113 a_n2903_n3924.n30 gnd 0.928343f
C1114 a_n2903_n3924.t55 gnd 1.3291f
C1115 a_n2903_n3924.n31 gnd 0.76636f
C1116 a_n2903_n3924.t33 gnd 1.3291f
C1117 a_n2903_n3924.n32 gnd 0.936111f
C1118 a_n2903_n3924.t41 gnd 1.3291f
C1119 a_n2903_n3924.n33 gnd 0.936111f
C1120 a_n2903_n3924.t36 gnd 1.3291f
C1121 a_n2903_n3924.n34 gnd 0.936111f
C1122 a_n2903_n3924.t39 gnd 1.3291f
C1123 a_n2903_n3924.n35 gnd 0.936111f
C1124 a_n2903_n3924.t34 gnd 1.3291f
C1125 a_n2903_n3924.n36 gnd 0.936111f
C1126 a_n2903_n3924.t32 gnd 1.3291f
C1127 a_n2903_n3924.n37 gnd 1.25723f
C1128 a_n2903_n3924.n38 gnd 1.02539f
C1129 a_n2903_n3924.t2 gnd 1.06972f
C1130 a_n2903_n3924.n39 gnd 0.625684f
C1131 a_n2903_n3924.t53 gnd 0.102925f
C1132 a_n2903_n3924.t48 gnd 0.102925f
C1133 a_n2903_n3924.n40 gnd 0.840607f
C1134 a_n2903_n3924.n41 gnd 0.382272f
C1135 a_n2903_n3924.t51 gnd 0.102925f
C1136 a_n2903_n3924.t44 gnd 0.102925f
C1137 a_n2903_n3924.n42 gnd 0.840607f
C1138 a_n2903_n3924.n43 gnd 0.382272f
C1139 a_n2903_n3924.t1 gnd 0.102925f
C1140 a_n2903_n3924.t38 gnd 0.102925f
C1141 a_n2903_n3924.n44 gnd 0.840607f
C1142 a_n2903_n3924.n45 gnd 0.382272f
C1143 a_n2903_n3924.t5 gnd 0.102925f
C1144 a_n2903_n3924.t4 gnd 0.102925f
C1145 a_n2903_n3924.n46 gnd 0.840607f
C1146 a_n2903_n3924.n47 gnd 0.382272f
C1147 a_n2903_n3924.t47 gnd 0.102925f
C1148 a_n2903_n3924.t6 gnd 0.102925f
C1149 a_n2903_n3924.n48 gnd 0.840607f
C1150 a_n2903_n3924.n49 gnd 0.382272f
C1151 a_n2903_n3924.t52 gnd 1.06972f
C1152 a_n2903_n3924.n50 gnd 0.383732f
C1153 a_n2903_n3924.t20 gnd 1.06972f
C1154 a_n2903_n3924.n51 gnd 0.383732f
C1155 a_n2903_n3924.t17 gnd 0.102925f
C1156 a_n2903_n3924.t22 gnd 0.102925f
C1157 a_n2903_n3924.n52 gnd 0.840607f
C1158 a_n2903_n3924.n53 gnd 0.382272f
C1159 a_n2903_n3924.t12 gnd 0.102925f
C1160 a_n2903_n3924.t11 gnd 0.102925f
C1161 a_n2903_n3924.n54 gnd 0.840607f
C1162 a_n2903_n3924.n55 gnd 0.382272f
C1163 a_n2903_n3924.n56 gnd 0.382275f
C1164 a_n2903_n3924.t29 gnd 0.102925f
C1165 a_n2903_n3924.n57 gnd 0.840604f
C1166 a_n2903_n3924.t30 gnd 0.102925f
C1167 plus.n0 gnd 0.02427f
C1168 plus.t21 gnd 0.343283f
C1169 plus.n1 gnd 0.02427f
C1170 plus.t22 gnd 0.343283f
C1171 plus.t16 gnd 0.343283f
C1172 plus.n2 gnd 0.152497f
C1173 plus.n3 gnd 0.02427f
C1174 plus.t17 gnd 0.343283f
C1175 plus.t11 gnd 0.343283f
C1176 plus.n4 gnd 0.152497f
C1177 plus.n5 gnd 0.02427f
C1178 plus.t5 gnd 0.343283f
C1179 plus.t6 gnd 0.343283f
C1180 plus.n6 gnd 0.152497f
C1181 plus.n7 gnd 0.02427f
C1182 plus.t23 gnd 0.343283f
C1183 plus.t24 gnd 0.343283f
C1184 plus.n8 gnd 0.152497f
C1185 plus.n9 gnd 0.02427f
C1186 plus.t18 gnd 0.343283f
C1187 plus.t13 gnd 0.343283f
C1188 plus.n10 gnd 0.157464f
C1189 plus.t15 gnd 0.355744f
C1190 plus.n11 gnd 0.141329f
C1191 plus.n12 gnd 0.104486f
C1192 plus.n13 gnd 0.005507f
C1193 plus.n14 gnd 0.152497f
C1194 plus.n15 gnd 0.005507f
C1195 plus.n16 gnd 0.02427f
C1196 plus.n17 gnd 0.02427f
C1197 plus.n18 gnd 0.02427f
C1198 plus.n19 gnd 0.005507f
C1199 plus.n20 gnd 0.152497f
C1200 plus.n21 gnd 0.005507f
C1201 plus.n22 gnd 0.02427f
C1202 plus.n23 gnd 0.02427f
C1203 plus.n24 gnd 0.02427f
C1204 plus.n25 gnd 0.005507f
C1205 plus.n26 gnd 0.152497f
C1206 plus.n27 gnd 0.005507f
C1207 plus.n28 gnd 0.02427f
C1208 plus.n29 gnd 0.02427f
C1209 plus.n30 gnd 0.02427f
C1210 plus.n31 gnd 0.005507f
C1211 plus.n32 gnd 0.152497f
C1212 plus.n33 gnd 0.005507f
C1213 plus.n34 gnd 0.02427f
C1214 plus.n35 gnd 0.02427f
C1215 plus.n36 gnd 0.02427f
C1216 plus.n37 gnd 0.005507f
C1217 plus.n38 gnd 0.152497f
C1218 plus.n39 gnd 0.005507f
C1219 plus.n40 gnd 0.152722f
C1220 plus.n41 gnd 0.274825f
C1221 plus.n42 gnd 0.02427f
C1222 plus.n43 gnd 0.005507f
C1223 plus.t10 gnd 0.343283f
C1224 plus.n44 gnd 0.02427f
C1225 plus.n45 gnd 0.005507f
C1226 plus.t12 gnd 0.343283f
C1227 plus.n46 gnd 0.02427f
C1228 plus.n47 gnd 0.005507f
C1229 plus.t7 gnd 0.343283f
C1230 plus.n48 gnd 0.02427f
C1231 plus.n49 gnd 0.005507f
C1232 plus.t27 gnd 0.343283f
C1233 plus.n50 gnd 0.02427f
C1234 plus.n51 gnd 0.005507f
C1235 plus.t26 gnd 0.343283f
C1236 plus.t20 gnd 0.355744f
C1237 plus.t19 gnd 0.343283f
C1238 plus.n52 gnd 0.157464f
C1239 plus.n53 gnd 0.141329f
C1240 plus.n54 gnd 0.104486f
C1241 plus.n55 gnd 0.02427f
C1242 plus.n56 gnd 0.152497f
C1243 plus.n57 gnd 0.005507f
C1244 plus.t25 gnd 0.343283f
C1245 plus.n58 gnd 0.152497f
C1246 plus.n59 gnd 0.02427f
C1247 plus.n60 gnd 0.02427f
C1248 plus.n61 gnd 0.02427f
C1249 plus.n62 gnd 0.152497f
C1250 plus.n63 gnd 0.005507f
C1251 plus.t9 gnd 0.343283f
C1252 plus.n64 gnd 0.152497f
C1253 plus.n65 gnd 0.02427f
C1254 plus.n66 gnd 0.02427f
C1255 plus.n67 gnd 0.02427f
C1256 plus.n68 gnd 0.152497f
C1257 plus.n69 gnd 0.005507f
C1258 plus.t14 gnd 0.343283f
C1259 plus.n70 gnd 0.152497f
C1260 plus.n71 gnd 0.02427f
C1261 plus.n72 gnd 0.02427f
C1262 plus.n73 gnd 0.02427f
C1263 plus.n74 gnd 0.152497f
C1264 plus.n75 gnd 0.005507f
C1265 plus.t28 gnd 0.343283f
C1266 plus.n76 gnd 0.152497f
C1267 plus.n77 gnd 0.02427f
C1268 plus.n78 gnd 0.02427f
C1269 plus.n79 gnd 0.02427f
C1270 plus.n80 gnd 0.152497f
C1271 plus.n81 gnd 0.005507f
C1272 plus.t8 gnd 0.343283f
C1273 plus.n82 gnd 0.152722f
C1274 plus.n83 gnd 0.803355f
C1275 plus.n84 gnd 1.20187f
C1276 plus.t2 gnd 0.041898f
C1277 plus.t3 gnd 0.007482f
C1278 plus.t1 gnd 0.007482f
C1279 plus.n85 gnd 0.024265f
C1280 plus.n86 gnd 0.188372f
C1281 plus.t4 gnd 0.007482f
C1282 plus.t0 gnd 0.007482f
C1283 plus.n87 gnd 0.024265f
C1284 plus.n88 gnd 0.141396f
C1285 plus.n89 gnd 2.59439f
C1286 CSoutput.n0 gnd 0.036233f
C1287 CSoutput.t108 gnd 0.239676f
C1288 CSoutput.n1 gnd 0.108226f
C1289 CSoutput.n2 gnd 0.036233f
C1290 CSoutput.t113 gnd 0.239676f
C1291 CSoutput.n3 gnd 0.028718f
C1292 CSoutput.n4 gnd 0.036233f
C1293 CSoutput.t102 gnd 0.239676f
C1294 CSoutput.n5 gnd 0.024764f
C1295 CSoutput.n6 gnd 0.036233f
C1296 CSoutput.t111 gnd 0.239676f
C1297 CSoutput.t117 gnd 0.239676f
C1298 CSoutput.n7 gnd 0.107046f
C1299 CSoutput.n8 gnd 0.036233f
C1300 CSoutput.t115 gnd 0.239676f
C1301 CSoutput.n9 gnd 0.023611f
C1302 CSoutput.n10 gnd 0.036233f
C1303 CSoutput.t103 gnd 0.239676f
C1304 CSoutput.t114 gnd 0.239676f
C1305 CSoutput.n11 gnd 0.107046f
C1306 CSoutput.n12 gnd 0.036233f
C1307 CSoutput.t112 gnd 0.239676f
C1308 CSoutput.n13 gnd 0.024764f
C1309 CSoutput.n14 gnd 0.036233f
C1310 CSoutput.t101 gnd 0.239676f
C1311 CSoutput.t107 gnd 0.239676f
C1312 CSoutput.n15 gnd 0.107046f
C1313 CSoutput.n16 gnd 0.036233f
C1314 CSoutput.t110 gnd 0.239676f
C1315 CSoutput.n17 gnd 0.026449f
C1316 CSoutput.t97 gnd 0.286419f
C1317 CSoutput.t99 gnd 0.239676f
C1318 CSoutput.n18 gnd 0.136656f
C1319 CSoutput.n19 gnd 0.132604f
C1320 CSoutput.n20 gnd 0.153836f
C1321 CSoutput.n21 gnd 0.036233f
C1322 CSoutput.n22 gnd 0.030241f
C1323 CSoutput.n23 gnd 0.107046f
C1324 CSoutput.n24 gnd 0.029151f
C1325 CSoutput.n25 gnd 0.028718f
C1326 CSoutput.n26 gnd 0.036233f
C1327 CSoutput.n27 gnd 0.036233f
C1328 CSoutput.n28 gnd 0.030008f
C1329 CSoutput.n29 gnd 0.025478f
C1330 CSoutput.n30 gnd 0.109429f
C1331 CSoutput.n31 gnd 0.025829f
C1332 CSoutput.n32 gnd 0.036233f
C1333 CSoutput.n33 gnd 0.036233f
C1334 CSoutput.n34 gnd 0.036233f
C1335 CSoutput.n35 gnd 0.029689f
C1336 CSoutput.n36 gnd 0.107046f
C1337 CSoutput.n37 gnd 0.028393f
C1338 CSoutput.n38 gnd 0.029476f
C1339 CSoutput.n39 gnd 0.036233f
C1340 CSoutput.n40 gnd 0.036233f
C1341 CSoutput.n41 gnd 0.030235f
C1342 CSoutput.n42 gnd 0.027635f
C1343 CSoutput.n43 gnd 0.107046f
C1344 CSoutput.n44 gnd 0.028335f
C1345 CSoutput.n45 gnd 0.036233f
C1346 CSoutput.n46 gnd 0.036233f
C1347 CSoutput.n47 gnd 0.036233f
C1348 CSoutput.n48 gnd 0.028335f
C1349 CSoutput.n49 gnd 0.107046f
C1350 CSoutput.n50 gnd 0.027635f
C1351 CSoutput.n51 gnd 0.030235f
C1352 CSoutput.n52 gnd 0.036233f
C1353 CSoutput.n53 gnd 0.036233f
C1354 CSoutput.n54 gnd 0.029476f
C1355 CSoutput.n55 gnd 0.028393f
C1356 CSoutput.n56 gnd 0.107046f
C1357 CSoutput.n57 gnd 0.029689f
C1358 CSoutput.n58 gnd 0.036233f
C1359 CSoutput.n59 gnd 0.036233f
C1360 CSoutput.n60 gnd 0.036233f
C1361 CSoutput.n61 gnd 0.025829f
C1362 CSoutput.n62 gnd 0.109429f
C1363 CSoutput.n63 gnd 0.025478f
C1364 CSoutput.t96 gnd 0.239676f
C1365 CSoutput.n64 gnd 0.107046f
C1366 CSoutput.n65 gnd 0.030008f
C1367 CSoutput.n66 gnd 0.036233f
C1368 CSoutput.n67 gnd 0.036233f
C1369 CSoutput.n68 gnd 0.036233f
C1370 CSoutput.n69 gnd 0.029151f
C1371 CSoutput.n70 gnd 0.107046f
C1372 CSoutput.n71 gnd 0.030241f
C1373 CSoutput.n72 gnd 0.026449f
C1374 CSoutput.n73 gnd 0.036233f
C1375 CSoutput.n74 gnd 0.036233f
C1376 CSoutput.n75 gnd 0.027429f
C1377 CSoutput.n76 gnd 0.01629f
C1378 CSoutput.t100 gnd 0.269293f
C1379 CSoutput.n77 gnd 0.133774f
C1380 CSoutput.n78 gnd 0.572406f
C1381 CSoutput.t68 gnd 0.045196f
C1382 CSoutput.t38 gnd 0.045196f
C1383 CSoutput.n79 gnd 0.349923f
C1384 CSoutput.t73 gnd 0.045196f
C1385 CSoutput.t50 gnd 0.045196f
C1386 CSoutput.n80 gnd 0.349299f
C1387 CSoutput.n81 gnd 0.354538f
C1388 CSoutput.t32 gnd 0.045196f
C1389 CSoutput.t55 gnd 0.045196f
C1390 CSoutput.n82 gnd 0.349299f
C1391 CSoutput.n83 gnd 0.174701f
C1392 CSoutput.t33 gnd 0.045196f
C1393 CSoutput.t45 gnd 0.045196f
C1394 CSoutput.n84 gnd 0.349299f
C1395 CSoutput.n85 gnd 0.320362f
C1396 CSoutput.t30 gnd 0.045196f
C1397 CSoutput.t66 gnd 0.045196f
C1398 CSoutput.n86 gnd 0.349923f
C1399 CSoutput.t60 gnd 0.045196f
C1400 CSoutput.t51 gnd 0.045196f
C1401 CSoutput.n87 gnd 0.349299f
C1402 CSoutput.n88 gnd 0.354538f
C1403 CSoutput.t39 gnd 0.045196f
C1404 CSoutput.t72 gnd 0.045196f
C1405 CSoutput.n89 gnd 0.349299f
C1406 CSoutput.n90 gnd 0.174701f
C1407 CSoutput.t59 gnd 0.045196f
C1408 CSoutput.t58 gnd 0.045196f
C1409 CSoutput.n91 gnd 0.349299f
C1410 CSoutput.n92 gnd 0.260523f
C1411 CSoutput.n93 gnd 0.328518f
C1412 CSoutput.t36 gnd 0.045196f
C1413 CSoutput.t71 gnd 0.045196f
C1414 CSoutput.n94 gnd 0.349923f
C1415 CSoutput.t65 gnd 0.045196f
C1416 CSoutput.t56 gnd 0.045196f
C1417 CSoutput.n95 gnd 0.349299f
C1418 CSoutput.n96 gnd 0.354538f
C1419 CSoutput.t46 gnd 0.045196f
C1420 CSoutput.t76 gnd 0.045196f
C1421 CSoutput.n97 gnd 0.349299f
C1422 CSoutput.n98 gnd 0.174701f
C1423 CSoutput.t62 gnd 0.045196f
C1424 CSoutput.t63 gnd 0.045196f
C1425 CSoutput.n99 gnd 0.349299f
C1426 CSoutput.n100 gnd 0.260523f
C1427 CSoutput.n101 gnd 0.367199f
C1428 CSoutput.n102 gnd 6.22684f
C1429 CSoutput.n104 gnd 0.640962f
C1430 CSoutput.n105 gnd 0.480721f
C1431 CSoutput.n106 gnd 0.640962f
C1432 CSoutput.n107 gnd 0.640962f
C1433 CSoutput.n108 gnd 1.72567f
C1434 CSoutput.n109 gnd 0.640962f
C1435 CSoutput.n110 gnd 0.640962f
C1436 CSoutput.t116 gnd 0.801202f
C1437 CSoutput.n111 gnd 0.640962f
C1438 CSoutput.n112 gnd 0.640962f
C1439 CSoutput.n116 gnd 0.640962f
C1440 CSoutput.n120 gnd 0.640962f
C1441 CSoutput.n121 gnd 0.640962f
C1442 CSoutput.n123 gnd 0.640962f
C1443 CSoutput.n128 gnd 0.640962f
C1444 CSoutput.n130 gnd 0.640962f
C1445 CSoutput.n131 gnd 0.640962f
C1446 CSoutput.n133 gnd 0.640962f
C1447 CSoutput.n134 gnd 0.640962f
C1448 CSoutput.n136 gnd 0.640962f
C1449 CSoutput.t105 gnd 10.710401f
C1450 CSoutput.n138 gnd 0.640962f
C1451 CSoutput.n139 gnd 0.480721f
C1452 CSoutput.n140 gnd 0.640962f
C1453 CSoutput.n141 gnd 0.640962f
C1454 CSoutput.n142 gnd 1.72567f
C1455 CSoutput.n143 gnd 0.640962f
C1456 CSoutput.n144 gnd 0.640962f
C1457 CSoutput.t104 gnd 0.801202f
C1458 CSoutput.n145 gnd 0.640962f
C1459 CSoutput.n146 gnd 0.640962f
C1460 CSoutput.n150 gnd 0.640962f
C1461 CSoutput.n154 gnd 0.640962f
C1462 CSoutput.n155 gnd 0.640962f
C1463 CSoutput.n157 gnd 0.640962f
C1464 CSoutput.n162 gnd 0.640962f
C1465 CSoutput.n164 gnd 0.640962f
C1466 CSoutput.n165 gnd 0.640962f
C1467 CSoutput.n167 gnd 0.640962f
C1468 CSoutput.n168 gnd 0.640962f
C1469 CSoutput.n170 gnd 0.640962f
C1470 CSoutput.n171 gnd 0.480721f
C1471 CSoutput.n173 gnd 0.640962f
C1472 CSoutput.n174 gnd 0.480721f
C1473 CSoutput.n175 gnd 0.640962f
C1474 CSoutput.n176 gnd 0.640962f
C1475 CSoutput.n177 gnd 1.72567f
C1476 CSoutput.n178 gnd 0.640962f
C1477 CSoutput.n179 gnd 0.640962f
C1478 CSoutput.t98 gnd 0.801202f
C1479 CSoutput.n180 gnd 0.640962f
C1480 CSoutput.n181 gnd 1.72567f
C1481 CSoutput.n183 gnd 0.640962f
C1482 CSoutput.n184 gnd 0.640962f
C1483 CSoutput.n186 gnd 0.640962f
C1484 CSoutput.n187 gnd 0.640962f
C1485 CSoutput.t106 gnd 10.535901f
C1486 CSoutput.t109 gnd 10.710401f
C1487 CSoutput.n193 gnd 2.01079f
C1488 CSoutput.n194 gnd 8.19123f
C1489 CSoutput.n195 gnd 8.53399f
C1490 CSoutput.n200 gnd 2.17823f
C1491 CSoutput.n206 gnd 0.640962f
C1492 CSoutput.n208 gnd 0.640962f
C1493 CSoutput.n210 gnd 0.640962f
C1494 CSoutput.n212 gnd 0.640962f
C1495 CSoutput.n214 gnd 0.640962f
C1496 CSoutput.n220 gnd 0.640962f
C1497 CSoutput.n227 gnd 1.17592f
C1498 CSoutput.n228 gnd 1.17592f
C1499 CSoutput.n229 gnd 0.640962f
C1500 CSoutput.n230 gnd 0.640962f
C1501 CSoutput.n232 gnd 0.480721f
C1502 CSoutput.n233 gnd 0.411695f
C1503 CSoutput.n235 gnd 0.480721f
C1504 CSoutput.n236 gnd 0.411695f
C1505 CSoutput.n237 gnd 0.480721f
C1506 CSoutput.n239 gnd 0.640962f
C1507 CSoutput.n241 gnd 1.72567f
C1508 CSoutput.n242 gnd 2.01079f
C1509 CSoutput.n243 gnd 7.53383f
C1510 CSoutput.n245 gnd 0.480721f
C1511 CSoutput.n246 gnd 1.23693f
C1512 CSoutput.n247 gnd 0.480721f
C1513 CSoutput.n249 gnd 0.640962f
C1514 CSoutput.n251 gnd 1.72567f
C1515 CSoutput.n252 gnd 3.75878f
C1516 CSoutput.t37 gnd 0.045196f
C1517 CSoutput.t69 gnd 0.045196f
C1518 CSoutput.n253 gnd 0.349923f
C1519 CSoutput.t48 gnd 0.045196f
C1520 CSoutput.t74 gnd 0.045196f
C1521 CSoutput.n254 gnd 0.349299f
C1522 CSoutput.n255 gnd 0.354538f
C1523 CSoutput.t64 gnd 0.045196f
C1524 CSoutput.t31 gnd 0.045196f
C1525 CSoutput.n256 gnd 0.349299f
C1526 CSoutput.n257 gnd 0.174701f
C1527 CSoutput.t44 gnd 0.045196f
C1528 CSoutput.t34 gnd 0.045196f
C1529 CSoutput.n258 gnd 0.349299f
C1530 CSoutput.n259 gnd 0.320362f
C1531 CSoutput.t54 gnd 0.045196f
C1532 CSoutput.t61 gnd 0.045196f
C1533 CSoutput.n260 gnd 0.349923f
C1534 CSoutput.t29 gnd 0.045196f
C1535 CSoutput.t42 gnd 0.045196f
C1536 CSoutput.n261 gnd 0.349299f
C1537 CSoutput.n262 gnd 0.354538f
C1538 CSoutput.t43 gnd 0.045196f
C1539 CSoutput.t70 gnd 0.045196f
C1540 CSoutput.n263 gnd 0.349299f
C1541 CSoutput.n264 gnd 0.174701f
C1542 CSoutput.t40 gnd 0.045196f
C1543 CSoutput.t41 gnd 0.045196f
C1544 CSoutput.n265 gnd 0.349299f
C1545 CSoutput.n266 gnd 0.260523f
C1546 CSoutput.n267 gnd 0.328518f
C1547 CSoutput.t57 gnd 0.045196f
C1548 CSoutput.t67 gnd 0.045196f
C1549 CSoutput.n268 gnd 0.349923f
C1550 CSoutput.t35 gnd 0.045196f
C1551 CSoutput.t52 gnd 0.045196f
C1552 CSoutput.n269 gnd 0.349299f
C1553 CSoutput.n270 gnd 0.354538f
C1554 CSoutput.t53 gnd 0.045196f
C1555 CSoutput.t75 gnd 0.045196f
C1556 CSoutput.n271 gnd 0.349299f
C1557 CSoutput.n272 gnd 0.174701f
C1558 CSoutput.t47 gnd 0.045196f
C1559 CSoutput.t49 gnd 0.045196f
C1560 CSoutput.n273 gnd 0.349297f
C1561 CSoutput.n274 gnd 0.260525f
C1562 CSoutput.n275 gnd 0.367199f
C1563 CSoutput.n276 gnd 9.133111f
C1564 CSoutput.t19 gnd 0.039547f
C1565 CSoutput.t92 gnd 0.039547f
C1566 CSoutput.n277 gnd 0.350616f
C1567 CSoutput.t27 gnd 0.039547f
C1568 CSoutput.t24 gnd 0.039547f
C1569 CSoutput.n278 gnd 0.349447f
C1570 CSoutput.n279 gnd 0.325619f
C1571 CSoutput.t28 gnd 0.039547f
C1572 CSoutput.t26 gnd 0.039547f
C1573 CSoutput.n280 gnd 0.349447f
C1574 CSoutput.n281 gnd 0.160515f
C1575 CSoutput.t93 gnd 0.039547f
C1576 CSoutput.t11 gnd 0.039547f
C1577 CSoutput.n282 gnd 0.349447f
C1578 CSoutput.n283 gnd 0.160515f
C1579 CSoutput.t77 gnd 0.039547f
C1580 CSoutput.t5 gnd 0.039547f
C1581 CSoutput.n284 gnd 0.349447f
C1582 CSoutput.n285 gnd 0.160515f
C1583 CSoutput.t90 gnd 0.039547f
C1584 CSoutput.t84 gnd 0.039547f
C1585 CSoutput.n286 gnd 0.349447f
C1586 CSoutput.n287 gnd 0.296022f
C1587 CSoutput.t86 gnd 0.039547f
C1588 CSoutput.t2 gnd 0.039547f
C1589 CSoutput.n288 gnd 0.350616f
C1590 CSoutput.t9 gnd 0.039547f
C1591 CSoutput.t21 gnd 0.039547f
C1592 CSoutput.n289 gnd 0.349447f
C1593 CSoutput.n290 gnd 0.325619f
C1594 CSoutput.t10 gnd 0.039547f
C1595 CSoutput.t22 gnd 0.039547f
C1596 CSoutput.n291 gnd 0.349447f
C1597 CSoutput.n292 gnd 0.160515f
C1598 CSoutput.t14 gnd 0.039547f
C1599 CSoutput.t79 gnd 0.039547f
C1600 CSoutput.n293 gnd 0.349447f
C1601 CSoutput.n294 gnd 0.160515f
C1602 CSoutput.t87 gnd 0.039547f
C1603 CSoutput.t12 gnd 0.039547f
C1604 CSoutput.n295 gnd 0.349447f
C1605 CSoutput.n296 gnd 0.160515f
C1606 CSoutput.t17 gnd 0.039547f
C1607 CSoutput.t15 gnd 0.039547f
C1608 CSoutput.n297 gnd 0.349447f
C1609 CSoutput.n298 gnd 0.243696f
C1610 CSoutput.n299 gnd 0.452806f
C1611 CSoutput.n300 gnd 9.50622f
C1612 CSoutput.t16 gnd 0.039547f
C1613 CSoutput.t13 gnd 0.039547f
C1614 CSoutput.n301 gnd 0.350616f
C1615 CSoutput.t20 gnd 0.039547f
C1616 CSoutput.t83 gnd 0.039547f
C1617 CSoutput.n302 gnd 0.349447f
C1618 CSoutput.n303 gnd 0.325619f
C1619 CSoutput.t1 gnd 0.039547f
C1620 CSoutput.t91 gnd 0.039547f
C1621 CSoutput.n304 gnd 0.349447f
C1622 CSoutput.n305 gnd 0.160515f
C1623 CSoutput.t80 gnd 0.039547f
C1624 CSoutput.t6 gnd 0.039547f
C1625 CSoutput.n306 gnd 0.349447f
C1626 CSoutput.n307 gnd 0.160515f
C1627 CSoutput.t81 gnd 0.039547f
C1628 CSoutput.t4 gnd 0.039547f
C1629 CSoutput.n308 gnd 0.349447f
C1630 CSoutput.n309 gnd 0.160515f
C1631 CSoutput.t8 gnd 0.039547f
C1632 CSoutput.t94 gnd 0.039547f
C1633 CSoutput.n310 gnd 0.349447f
C1634 CSoutput.n311 gnd 0.296022f
C1635 CSoutput.t78 gnd 0.039547f
C1636 CSoutput.t82 gnd 0.039547f
C1637 CSoutput.n312 gnd 0.350616f
C1638 CSoutput.t3 gnd 0.039547f
C1639 CSoutput.t89 gnd 0.039547f
C1640 CSoutput.n313 gnd 0.349447f
C1641 CSoutput.n314 gnd 0.325619f
C1642 CSoutput.t0 gnd 0.039547f
C1643 CSoutput.t25 gnd 0.039547f
C1644 CSoutput.n315 gnd 0.349447f
C1645 CSoutput.n316 gnd 0.160515f
C1646 CSoutput.t18 gnd 0.039547f
C1647 CSoutput.t85 gnd 0.039547f
C1648 CSoutput.n317 gnd 0.349447f
C1649 CSoutput.n318 gnd 0.160515f
C1650 CSoutput.t95 gnd 0.039547f
C1651 CSoutput.t7 gnd 0.039547f
C1652 CSoutput.n319 gnd 0.349447f
C1653 CSoutput.n320 gnd 0.160515f
C1654 CSoutput.t23 gnd 0.039547f
C1655 CSoutput.t88 gnd 0.039547f
C1656 CSoutput.n321 gnd 0.349447f
C1657 CSoutput.n322 gnd 0.243696f
C1658 CSoutput.n323 gnd 0.452806f
C1659 CSoutput.n324 gnd 5.27357f
C1660 CSoutput.n325 gnd 11.6641f
C1661 a_n6308_8799.n0 gnd 3.87851f
C1662 a_n6308_8799.n1 gnd 1.93319f
C1663 a_n6308_8799.n2 gnd 3.26499f
C1664 a_n6308_8799.n3 gnd 0.795133f
C1665 a_n6308_8799.n4 gnd 0.209403f
C1666 a_n6308_8799.n5 gnd 0.288684f
C1667 a_n6308_8799.n6 gnd 0.219028f
C1668 a_n6308_8799.n7 gnd 0.209403f
C1669 a_n6308_8799.n8 gnd 0.288684f
C1670 a_n6308_8799.n9 gnd 0.219028f
C1671 a_n6308_8799.n10 gnd 0.209403f
C1672 a_n6308_8799.n11 gnd 0.454941f
C1673 a_n6308_8799.n12 gnd 0.219028f
C1674 a_n6308_8799.n13 gnd 0.209403f
C1675 a_n6308_8799.n14 gnd 0.323729f
C1676 a_n6308_8799.n15 gnd 0.183982f
C1677 a_n6308_8799.n16 gnd 0.209403f
C1678 a_n6308_8799.n17 gnd 0.323729f
C1679 a_n6308_8799.n18 gnd 0.183982f
C1680 a_n6308_8799.n19 gnd 0.209403f
C1681 a_n6308_8799.n20 gnd 0.323729f
C1682 a_n6308_8799.n21 gnd 0.350239f
C1683 a_n6308_8799.n22 gnd 1.53476f
C1684 a_n6308_8799.n23 gnd 1.02802f
C1685 a_n6308_8799.n24 gnd 2.53883f
C1686 a_n6308_8799.n25 gnd 0.252102f
C1687 a_n6308_8799.n26 gnd 0.004706f
C1688 a_n6308_8799.n27 gnd 0.010179f
C1689 a_n6308_8799.n28 gnd 0.010179f
C1690 a_n6308_8799.n29 gnd 0.004706f
C1691 a_n6308_8799.n30 gnd 0.252102f
C1692 a_n6308_8799.n31 gnd 0.004706f
C1693 a_n6308_8799.n32 gnd 0.010179f
C1694 a_n6308_8799.n33 gnd 0.010179f
C1695 a_n6308_8799.n34 gnd 0.004706f
C1696 a_n6308_8799.n35 gnd 0.252102f
C1697 a_n6308_8799.n36 gnd 0.004706f
C1698 a_n6308_8799.n37 gnd 0.010179f
C1699 a_n6308_8799.n38 gnd 0.010179f
C1700 a_n6308_8799.n39 gnd 0.004706f
C1701 a_n6308_8799.n40 gnd 0.004706f
C1702 a_n6308_8799.n41 gnd 0.010179f
C1703 a_n6308_8799.n42 gnd 0.010179f
C1704 a_n6308_8799.n43 gnd 0.004706f
C1705 a_n6308_8799.n44 gnd 0.252102f
C1706 a_n6308_8799.n45 gnd 0.004706f
C1707 a_n6308_8799.n46 gnd 0.010179f
C1708 a_n6308_8799.n47 gnd 0.010179f
C1709 a_n6308_8799.n48 gnd 0.004706f
C1710 a_n6308_8799.n49 gnd 0.252102f
C1711 a_n6308_8799.n50 gnd 0.004706f
C1712 a_n6308_8799.n51 gnd 0.010179f
C1713 a_n6308_8799.n52 gnd 0.010179f
C1714 a_n6308_8799.n53 gnd 0.004706f
C1715 a_n6308_8799.n54 gnd 0.252102f
C1716 a_n6308_8799.t8 gnd 0.145244f
C1717 a_n6308_8799.t11 gnd 0.145244f
C1718 a_n6308_8799.t4 gnd 0.145244f
C1719 a_n6308_8799.n55 gnd 1.14557f
C1720 a_n6308_8799.t10 gnd 0.145244f
C1721 a_n6308_8799.t7 gnd 0.145244f
C1722 a_n6308_8799.n56 gnd 1.14368f
C1723 a_n6308_8799.t13 gnd 0.145244f
C1724 a_n6308_8799.t1 gnd 0.145244f
C1725 a_n6308_8799.n57 gnd 1.14556f
C1726 a_n6308_8799.t6 gnd 0.145244f
C1727 a_n6308_8799.t12 gnd 0.145244f
C1728 a_n6308_8799.n58 gnd 1.14368f
C1729 a_n6308_8799.t3 gnd 0.145244f
C1730 a_n6308_8799.t9 gnd 0.145244f
C1731 a_n6308_8799.n59 gnd 1.14368f
C1732 a_n6308_8799.t14 gnd 0.145244f
C1733 a_n6308_8799.t2 gnd 0.145244f
C1734 a_n6308_8799.n60 gnd 1.14368f
C1735 a_n6308_8799.n61 gnd 3.2457f
C1736 a_n6308_8799.t35 gnd 0.112968f
C1737 a_n6308_8799.t37 gnd 0.112968f
C1738 a_n6308_8799.n62 gnd 1.00044f
C1739 a_n6308_8799.t23 gnd 0.112968f
C1740 a_n6308_8799.t34 gnd 0.112968f
C1741 a_n6308_8799.n63 gnd 0.998224f
C1742 a_n6308_8799.t31 gnd 0.112968f
C1743 a_n6308_8799.t30 gnd 0.112968f
C1744 a_n6308_8799.n64 gnd 0.998224f
C1745 a_n6308_8799.t20 gnd 0.112968f
C1746 a_n6308_8799.t36 gnd 0.112968f
C1747 a_n6308_8799.n65 gnd 1.00044f
C1748 a_n6308_8799.t24 gnd 0.112968f
C1749 a_n6308_8799.t19 gnd 0.112968f
C1750 a_n6308_8799.n66 gnd 0.998223f
C1751 a_n6308_8799.t38 gnd 0.112968f
C1752 a_n6308_8799.t17 gnd 0.112968f
C1753 a_n6308_8799.n67 gnd 0.998223f
C1754 a_n6308_8799.t28 gnd 0.112968f
C1755 a_n6308_8799.t21 gnd 0.112968f
C1756 a_n6308_8799.n68 gnd 1.00044f
C1757 a_n6308_8799.t33 gnd 0.112968f
C1758 a_n6308_8799.t39 gnd 0.112968f
C1759 a_n6308_8799.n69 gnd 0.998223f
C1760 a_n6308_8799.t18 gnd 0.112968f
C1761 a_n6308_8799.t22 gnd 0.112968f
C1762 a_n6308_8799.n70 gnd 0.998223f
C1763 a_n6308_8799.t26 gnd 0.112968f
C1764 a_n6308_8799.t27 gnd 0.112968f
C1765 a_n6308_8799.n71 gnd 0.998224f
C1766 a_n6308_8799.t25 gnd 0.112968f
C1767 a_n6308_8799.t16 gnd 0.112968f
C1768 a_n6308_8799.n72 gnd 0.998224f
C1769 a_n6308_8799.t29 gnd 0.112968f
C1770 a_n6308_8799.t32 gnd 0.112968f
C1771 a_n6308_8799.n73 gnd 0.998224f
C1772 a_n6308_8799.t60 gnd 0.602251f
C1773 a_n6308_8799.n74 gnd 0.270677f
C1774 a_n6308_8799.t40 gnd 0.602251f
C1775 a_n6308_8799.t53 gnd 0.602251f
C1776 a_n6308_8799.t54 gnd 0.61365f
C1777 a_n6308_8799.n75 gnd 0.252473f
C1778 a_n6308_8799.n76 gnd 0.273084f
C1779 a_n6308_8799.t70 gnd 0.602251f
C1780 a_n6308_8799.n77 gnd 0.270677f
C1781 a_n6308_8799.n78 gnd 0.266233f
C1782 a_n6308_8799.t51 gnd 0.602251f
C1783 a_n6308_8799.n79 gnd 0.266233f
C1784 a_n6308_8799.t80 gnd 0.602251f
C1785 a_n6308_8799.n80 gnd 0.273084f
C1786 a_n6308_8799.t45 gnd 0.613639f
C1787 a_n6308_8799.t65 gnd 0.602251f
C1788 a_n6308_8799.n81 gnd 0.270677f
C1789 a_n6308_8799.t44 gnd 0.602251f
C1790 a_n6308_8799.t58 gnd 0.602251f
C1791 a_n6308_8799.t57 gnd 0.61365f
C1792 a_n6308_8799.n82 gnd 0.252473f
C1793 a_n6308_8799.n83 gnd 0.273084f
C1794 a_n6308_8799.t77 gnd 0.602251f
C1795 a_n6308_8799.n84 gnd 0.270677f
C1796 a_n6308_8799.n85 gnd 0.266233f
C1797 a_n6308_8799.t56 gnd 0.602251f
C1798 a_n6308_8799.n86 gnd 0.266233f
C1799 a_n6308_8799.t86 gnd 0.602251f
C1800 a_n6308_8799.n87 gnd 0.273084f
C1801 a_n6308_8799.t50 gnd 0.613639f
C1802 a_n6308_8799.n88 gnd 0.905765f
C1803 a_n6308_8799.t66 gnd 0.602251f
C1804 a_n6308_8799.n89 gnd 0.270677f
C1805 a_n6308_8799.t61 gnd 0.602251f
C1806 a_n6308_8799.t71 gnd 0.602251f
C1807 a_n6308_8799.t83 gnd 0.61365f
C1808 a_n6308_8799.n90 gnd 0.252473f
C1809 a_n6308_8799.n91 gnd 0.273084f
C1810 a_n6308_8799.t84 gnd 0.602251f
C1811 a_n6308_8799.n92 gnd 0.270677f
C1812 a_n6308_8799.n93 gnd 0.266233f
C1813 a_n6308_8799.t43 gnd 0.602251f
C1814 a_n6308_8799.n94 gnd 0.266233f
C1815 a_n6308_8799.t48 gnd 0.602251f
C1816 a_n6308_8799.n95 gnd 0.273084f
C1817 a_n6308_8799.t78 gnd 0.613639f
C1818 a_n6308_8799.n96 gnd 1.63199f
C1819 a_n6308_8799.t59 gnd 0.613639f
C1820 a_n6308_8799.t49 gnd 0.602251f
C1821 a_n6308_8799.t81 gnd 0.602251f
C1822 a_n6308_8799.n97 gnd 0.270677f
C1823 a_n6308_8799.t64 gnd 0.602251f
C1824 a_n6308_8799.t63 gnd 0.602251f
C1825 a_n6308_8799.t41 gnd 0.602251f
C1826 a_n6308_8799.n98 gnd 0.270677f
C1827 a_n6308_8799.t67 gnd 0.61365f
C1828 a_n6308_8799.n99 gnd 0.252473f
C1829 a_n6308_8799.t69 gnd 0.602251f
C1830 a_n6308_8799.n100 gnd 0.273084f
C1831 a_n6308_8799.n101 gnd 0.266233f
C1832 a_n6308_8799.n102 gnd 0.266233f
C1833 a_n6308_8799.n103 gnd 0.273084f
C1834 a_n6308_8799.t62 gnd 0.613639f
C1835 a_n6308_8799.t55 gnd 0.602251f
C1836 a_n6308_8799.t87 gnd 0.602251f
C1837 a_n6308_8799.n104 gnd 0.270677f
C1838 a_n6308_8799.t74 gnd 0.602251f
C1839 a_n6308_8799.t73 gnd 0.602251f
C1840 a_n6308_8799.t46 gnd 0.602251f
C1841 a_n6308_8799.n105 gnd 0.270677f
C1842 a_n6308_8799.t75 gnd 0.61365f
C1843 a_n6308_8799.n106 gnd 0.252473f
C1844 a_n6308_8799.t76 gnd 0.602251f
C1845 a_n6308_8799.n107 gnd 0.273084f
C1846 a_n6308_8799.n108 gnd 0.266233f
C1847 a_n6308_8799.n109 gnd 0.266233f
C1848 a_n6308_8799.n110 gnd 0.273084f
C1849 a_n6308_8799.n111 gnd 0.905765f
C1850 a_n6308_8799.t79 gnd 0.613639f
C1851 a_n6308_8799.t47 gnd 0.602251f
C1852 a_n6308_8799.t68 gnd 0.602251f
C1853 a_n6308_8799.n112 gnd 0.270677f
C1854 a_n6308_8799.t42 gnd 0.602251f
C1855 a_n6308_8799.t52 gnd 0.602251f
C1856 a_n6308_8799.t85 gnd 0.602251f
C1857 a_n6308_8799.n113 gnd 0.270677f
C1858 a_n6308_8799.t82 gnd 0.61365f
C1859 a_n6308_8799.n114 gnd 0.252473f
C1860 a_n6308_8799.t72 gnd 0.602251f
C1861 a_n6308_8799.n115 gnd 0.273084f
C1862 a_n6308_8799.n116 gnd 0.266233f
C1863 a_n6308_8799.n117 gnd 0.266233f
C1864 a_n6308_8799.n118 gnd 0.273084f
C1865 a_n6308_8799.n119 gnd 1.19577f
C1866 a_n6308_8799.n120 gnd 14.0664f
C1867 a_n6308_8799.n121 gnd 4.4076f
C1868 a_n6308_8799.n122 gnd 6.38788f
C1869 a_n6308_8799.t5 gnd 0.145244f
C1870 a_n6308_8799.t15 gnd 0.145244f
C1871 a_n6308_8799.n123 gnd 1.14368f
C1872 a_n6308_8799.n124 gnd 1.14368f
C1873 a_n6308_8799.t0 gnd 0.145244f
C1874 vdd.t131 gnd 0.03154f
C1875 vdd.t116 gnd 0.03154f
C1876 vdd.n0 gnd 0.248764f
C1877 vdd.t96 gnd 0.03154f
C1878 vdd.t126 gnd 0.03154f
C1879 vdd.n1 gnd 0.248353f
C1880 vdd.n2 gnd 0.229029f
C1881 vdd.t113 gnd 0.03154f
C1882 vdd.t135 gnd 0.03154f
C1883 vdd.n3 gnd 0.248353f
C1884 vdd.n4 gnd 0.115828f
C1885 vdd.t137 gnd 0.03154f
C1886 vdd.t119 gnd 0.03154f
C1887 vdd.n5 gnd 0.248353f
C1888 vdd.n6 gnd 0.108683f
C1889 vdd.t140 gnd 0.03154f
C1890 vdd.t111 gnd 0.03154f
C1891 vdd.n7 gnd 0.248764f
C1892 vdd.t98 gnd 0.03154f
C1893 vdd.t133 gnd 0.03154f
C1894 vdd.n8 gnd 0.248353f
C1895 vdd.n9 gnd 0.229029f
C1896 vdd.t124 gnd 0.03154f
C1897 vdd.t101 gnd 0.03154f
C1898 vdd.n10 gnd 0.248353f
C1899 vdd.n11 gnd 0.115828f
C1900 vdd.t108 gnd 0.03154f
C1901 vdd.t121 gnd 0.03154f
C1902 vdd.n12 gnd 0.248353f
C1903 vdd.n13 gnd 0.108683f
C1904 vdd.n14 gnd 0.076837f
C1905 vdd.t157 gnd 0.017522f
C1906 vdd.t153 gnd 0.017522f
C1907 vdd.n15 gnd 0.161286f
C1908 vdd.t203 gnd 0.017522f
C1909 vdd.t186 gnd 0.017522f
C1910 vdd.n16 gnd 0.160814f
C1911 vdd.n17 gnd 0.279867f
C1912 vdd.t174 gnd 0.017522f
C1913 vdd.t155 gnd 0.017522f
C1914 vdd.n18 gnd 0.160814f
C1915 vdd.n19 gnd 0.115785f
C1916 vdd.t151 gnd 0.017522f
C1917 vdd.t152 gnd 0.017522f
C1918 vdd.n20 gnd 0.161286f
C1919 vdd.t173 gnd 0.017522f
C1920 vdd.t156 gnd 0.017522f
C1921 vdd.n21 gnd 0.160814f
C1922 vdd.n22 gnd 0.279867f
C1923 vdd.t154 gnd 0.017522f
C1924 vdd.t185 gnd 0.017522f
C1925 vdd.n23 gnd 0.160814f
C1926 vdd.n24 gnd 0.115785f
C1927 vdd.t187 gnd 0.017522f
C1928 vdd.t188 gnd 0.017522f
C1929 vdd.n25 gnd 0.160814f
C1930 vdd.t0 gnd 0.017522f
C1931 vdd.t1 gnd 0.017522f
C1932 vdd.n26 gnd 0.160814f
C1933 vdd.n27 gnd 18.334099f
C1934 vdd.n28 gnd 6.69557f
C1935 vdd.n29 gnd 0.004779f
C1936 vdd.n30 gnd 0.004435f
C1937 vdd.n31 gnd 0.002453f
C1938 vdd.n32 gnd 0.005633f
C1939 vdd.n33 gnd 0.002383f
C1940 vdd.n34 gnd 0.002523f
C1941 vdd.n35 gnd 0.004435f
C1942 vdd.n36 gnd 0.002383f
C1943 vdd.n37 gnd 0.005633f
C1944 vdd.n38 gnd 0.002523f
C1945 vdd.n39 gnd 0.004435f
C1946 vdd.n40 gnd 0.002383f
C1947 vdd.n41 gnd 0.004224f
C1948 vdd.n42 gnd 0.004237f
C1949 vdd.t172 gnd 0.012101f
C1950 vdd.n43 gnd 0.026925f
C1951 vdd.n44 gnd 0.140125f
C1952 vdd.n45 gnd 0.002383f
C1953 vdd.n46 gnd 0.002523f
C1954 vdd.n47 gnd 0.005633f
C1955 vdd.n48 gnd 0.005633f
C1956 vdd.n49 gnd 0.002523f
C1957 vdd.n50 gnd 0.002383f
C1958 vdd.n51 gnd 0.004435f
C1959 vdd.n52 gnd 0.004435f
C1960 vdd.n53 gnd 0.002383f
C1961 vdd.n54 gnd 0.002523f
C1962 vdd.n55 gnd 0.005633f
C1963 vdd.n56 gnd 0.005633f
C1964 vdd.n57 gnd 0.002523f
C1965 vdd.n58 gnd 0.002383f
C1966 vdd.n59 gnd 0.004435f
C1967 vdd.n60 gnd 0.004435f
C1968 vdd.n61 gnd 0.002383f
C1969 vdd.n62 gnd 0.002523f
C1970 vdd.n63 gnd 0.005633f
C1971 vdd.n64 gnd 0.005633f
C1972 vdd.n65 gnd 0.013317f
C1973 vdd.n66 gnd 0.002453f
C1974 vdd.n67 gnd 0.002383f
C1975 vdd.n68 gnd 0.011462f
C1976 vdd.n69 gnd 0.008002f
C1977 vdd.t192 gnd 0.028036f
C1978 vdd.t79 gnd 0.028036f
C1979 vdd.n70 gnd 0.192681f
C1980 vdd.n71 gnd 0.151515f
C1981 vdd.t175 gnd 0.028036f
C1982 vdd.t181 gnd 0.028036f
C1983 vdd.n72 gnd 0.192681f
C1984 vdd.n73 gnd 0.122271f
C1985 vdd.t196 gnd 0.028036f
C1986 vdd.t177 gnd 0.028036f
C1987 vdd.n74 gnd 0.192681f
C1988 vdd.n75 gnd 0.122271f
C1989 vdd.n76 gnd 0.004779f
C1990 vdd.n77 gnd 0.004435f
C1991 vdd.n78 gnd 0.002453f
C1992 vdd.n79 gnd 0.005633f
C1993 vdd.n80 gnd 0.002383f
C1994 vdd.n81 gnd 0.002523f
C1995 vdd.n82 gnd 0.004435f
C1996 vdd.n83 gnd 0.002383f
C1997 vdd.n84 gnd 0.005633f
C1998 vdd.n85 gnd 0.002523f
C1999 vdd.n86 gnd 0.004435f
C2000 vdd.n87 gnd 0.002383f
C2001 vdd.n88 gnd 0.004224f
C2002 vdd.n89 gnd 0.004237f
C2003 vdd.t179 gnd 0.012101f
C2004 vdd.n90 gnd 0.026925f
C2005 vdd.n91 gnd 0.140125f
C2006 vdd.n92 gnd 0.002383f
C2007 vdd.n93 gnd 0.002523f
C2008 vdd.n94 gnd 0.005633f
C2009 vdd.n95 gnd 0.005633f
C2010 vdd.n96 gnd 0.002523f
C2011 vdd.n97 gnd 0.002383f
C2012 vdd.n98 gnd 0.004435f
C2013 vdd.n99 gnd 0.004435f
C2014 vdd.n100 gnd 0.002383f
C2015 vdd.n101 gnd 0.002523f
C2016 vdd.n102 gnd 0.005633f
C2017 vdd.n103 gnd 0.005633f
C2018 vdd.n104 gnd 0.002523f
C2019 vdd.n105 gnd 0.002383f
C2020 vdd.n106 gnd 0.004435f
C2021 vdd.n107 gnd 0.004435f
C2022 vdd.n108 gnd 0.002383f
C2023 vdd.n109 gnd 0.002523f
C2024 vdd.n110 gnd 0.005633f
C2025 vdd.n111 gnd 0.005633f
C2026 vdd.n112 gnd 0.013317f
C2027 vdd.n113 gnd 0.002453f
C2028 vdd.n114 gnd 0.002383f
C2029 vdd.n115 gnd 0.011462f
C2030 vdd.n116 gnd 0.007751f
C2031 vdd.n117 gnd 0.090971f
C2032 vdd.n118 gnd 0.004779f
C2033 vdd.n119 gnd 0.004435f
C2034 vdd.n120 gnd 0.002453f
C2035 vdd.n121 gnd 0.005633f
C2036 vdd.n122 gnd 0.002383f
C2037 vdd.n123 gnd 0.002523f
C2038 vdd.n124 gnd 0.004435f
C2039 vdd.n125 gnd 0.002383f
C2040 vdd.n126 gnd 0.005633f
C2041 vdd.n127 gnd 0.002523f
C2042 vdd.n128 gnd 0.004435f
C2043 vdd.n129 gnd 0.002383f
C2044 vdd.n130 gnd 0.004224f
C2045 vdd.n131 gnd 0.004237f
C2046 vdd.t163 gnd 0.012101f
C2047 vdd.n132 gnd 0.026925f
C2048 vdd.n133 gnd 0.140125f
C2049 vdd.n134 gnd 0.002383f
C2050 vdd.n135 gnd 0.002523f
C2051 vdd.n136 gnd 0.005633f
C2052 vdd.n137 gnd 0.005633f
C2053 vdd.n138 gnd 0.002523f
C2054 vdd.n139 gnd 0.002383f
C2055 vdd.n140 gnd 0.004435f
C2056 vdd.n141 gnd 0.004435f
C2057 vdd.n142 gnd 0.002383f
C2058 vdd.n143 gnd 0.002523f
C2059 vdd.n144 gnd 0.005633f
C2060 vdd.n145 gnd 0.005633f
C2061 vdd.n146 gnd 0.002523f
C2062 vdd.n147 gnd 0.002383f
C2063 vdd.n148 gnd 0.004435f
C2064 vdd.n149 gnd 0.004435f
C2065 vdd.n150 gnd 0.002383f
C2066 vdd.n151 gnd 0.002523f
C2067 vdd.n152 gnd 0.005633f
C2068 vdd.n153 gnd 0.005633f
C2069 vdd.n154 gnd 0.013317f
C2070 vdd.n155 gnd 0.002453f
C2071 vdd.n156 gnd 0.002383f
C2072 vdd.n157 gnd 0.011462f
C2073 vdd.n158 gnd 0.008002f
C2074 vdd.t148 gnd 0.028036f
C2075 vdd.t88 gnd 0.028036f
C2076 vdd.n159 gnd 0.192681f
C2077 vdd.n160 gnd 0.151515f
C2078 vdd.t83 gnd 0.028036f
C2079 vdd.t178 gnd 0.028036f
C2080 vdd.n161 gnd 0.192681f
C2081 vdd.n162 gnd 0.122271f
C2082 vdd.t191 gnd 0.028036f
C2083 vdd.t193 gnd 0.028036f
C2084 vdd.n163 gnd 0.192681f
C2085 vdd.n164 gnd 0.122271f
C2086 vdd.n165 gnd 0.004779f
C2087 vdd.n166 gnd 0.004435f
C2088 vdd.n167 gnd 0.002453f
C2089 vdd.n168 gnd 0.005633f
C2090 vdd.n169 gnd 0.002383f
C2091 vdd.n170 gnd 0.002523f
C2092 vdd.n171 gnd 0.004435f
C2093 vdd.n172 gnd 0.002383f
C2094 vdd.n173 gnd 0.005633f
C2095 vdd.n174 gnd 0.002523f
C2096 vdd.n175 gnd 0.004435f
C2097 vdd.n176 gnd 0.002383f
C2098 vdd.n177 gnd 0.004224f
C2099 vdd.n178 gnd 0.004237f
C2100 vdd.t85 gnd 0.012101f
C2101 vdd.n179 gnd 0.026925f
C2102 vdd.n180 gnd 0.140125f
C2103 vdd.n181 gnd 0.002383f
C2104 vdd.n182 gnd 0.002523f
C2105 vdd.n183 gnd 0.005633f
C2106 vdd.n184 gnd 0.005633f
C2107 vdd.n185 gnd 0.002523f
C2108 vdd.n186 gnd 0.002383f
C2109 vdd.n187 gnd 0.004435f
C2110 vdd.n188 gnd 0.004435f
C2111 vdd.n189 gnd 0.002383f
C2112 vdd.n190 gnd 0.002523f
C2113 vdd.n191 gnd 0.005633f
C2114 vdd.n192 gnd 0.005633f
C2115 vdd.n193 gnd 0.002523f
C2116 vdd.n194 gnd 0.002383f
C2117 vdd.n195 gnd 0.004435f
C2118 vdd.n196 gnd 0.004435f
C2119 vdd.n197 gnd 0.002383f
C2120 vdd.n198 gnd 0.002523f
C2121 vdd.n199 gnd 0.005633f
C2122 vdd.n200 gnd 0.005633f
C2123 vdd.n201 gnd 0.013317f
C2124 vdd.n202 gnd 0.002453f
C2125 vdd.n203 gnd 0.002383f
C2126 vdd.n204 gnd 0.011462f
C2127 vdd.n205 gnd 0.007751f
C2128 vdd.n206 gnd 0.054118f
C2129 vdd.n207 gnd 0.195002f
C2130 vdd.n208 gnd 0.004779f
C2131 vdd.n209 gnd 0.004435f
C2132 vdd.n210 gnd 0.002453f
C2133 vdd.n211 gnd 0.005633f
C2134 vdd.n212 gnd 0.002383f
C2135 vdd.n213 gnd 0.002523f
C2136 vdd.n214 gnd 0.004435f
C2137 vdd.n215 gnd 0.002383f
C2138 vdd.n216 gnd 0.005633f
C2139 vdd.n217 gnd 0.002523f
C2140 vdd.n218 gnd 0.004435f
C2141 vdd.n219 gnd 0.002383f
C2142 vdd.n220 gnd 0.004224f
C2143 vdd.n221 gnd 0.004237f
C2144 vdd.t170 gnd 0.012101f
C2145 vdd.n222 gnd 0.026925f
C2146 vdd.n223 gnd 0.140125f
C2147 vdd.n224 gnd 0.002383f
C2148 vdd.n225 gnd 0.002523f
C2149 vdd.n226 gnd 0.005633f
C2150 vdd.n227 gnd 0.005633f
C2151 vdd.n228 gnd 0.002523f
C2152 vdd.n229 gnd 0.002383f
C2153 vdd.n230 gnd 0.004435f
C2154 vdd.n231 gnd 0.004435f
C2155 vdd.n232 gnd 0.002383f
C2156 vdd.n233 gnd 0.002523f
C2157 vdd.n234 gnd 0.005633f
C2158 vdd.n235 gnd 0.005633f
C2159 vdd.n236 gnd 0.002523f
C2160 vdd.n237 gnd 0.002383f
C2161 vdd.n238 gnd 0.004435f
C2162 vdd.n239 gnd 0.004435f
C2163 vdd.n240 gnd 0.002383f
C2164 vdd.n241 gnd 0.002523f
C2165 vdd.n242 gnd 0.005633f
C2166 vdd.n243 gnd 0.005633f
C2167 vdd.n244 gnd 0.013317f
C2168 vdd.n245 gnd 0.002453f
C2169 vdd.n246 gnd 0.002383f
C2170 vdd.n247 gnd 0.011462f
C2171 vdd.n248 gnd 0.008002f
C2172 vdd.t190 gnd 0.028036f
C2173 vdd.t202 gnd 0.028036f
C2174 vdd.n249 gnd 0.192681f
C2175 vdd.n250 gnd 0.151515f
C2176 vdd.t197 gnd 0.028036f
C2177 vdd.t165 gnd 0.028036f
C2178 vdd.n251 gnd 0.192681f
C2179 vdd.n252 gnd 0.122271f
C2180 vdd.t161 gnd 0.028036f
C2181 vdd.t81 gnd 0.028036f
C2182 vdd.n253 gnd 0.192681f
C2183 vdd.n254 gnd 0.122271f
C2184 vdd.n255 gnd 0.004779f
C2185 vdd.n256 gnd 0.004435f
C2186 vdd.n257 gnd 0.002453f
C2187 vdd.n258 gnd 0.005633f
C2188 vdd.n259 gnd 0.002383f
C2189 vdd.n260 gnd 0.002523f
C2190 vdd.n261 gnd 0.004435f
C2191 vdd.n262 gnd 0.002383f
C2192 vdd.n263 gnd 0.005633f
C2193 vdd.n264 gnd 0.002523f
C2194 vdd.n265 gnd 0.004435f
C2195 vdd.n266 gnd 0.002383f
C2196 vdd.n267 gnd 0.004224f
C2197 vdd.n268 gnd 0.004237f
C2198 vdd.t184 gnd 0.012101f
C2199 vdd.n269 gnd 0.026925f
C2200 vdd.n270 gnd 0.140125f
C2201 vdd.n271 gnd 0.002383f
C2202 vdd.n272 gnd 0.002523f
C2203 vdd.n273 gnd 0.005633f
C2204 vdd.n274 gnd 0.005633f
C2205 vdd.n275 gnd 0.002523f
C2206 vdd.n276 gnd 0.002383f
C2207 vdd.n277 gnd 0.004435f
C2208 vdd.n278 gnd 0.004435f
C2209 vdd.n279 gnd 0.002383f
C2210 vdd.n280 gnd 0.002523f
C2211 vdd.n281 gnd 0.005633f
C2212 vdd.n282 gnd 0.005633f
C2213 vdd.n283 gnd 0.002523f
C2214 vdd.n284 gnd 0.002383f
C2215 vdd.n285 gnd 0.004435f
C2216 vdd.n286 gnd 0.004435f
C2217 vdd.n287 gnd 0.002383f
C2218 vdd.n288 gnd 0.002523f
C2219 vdd.n289 gnd 0.005633f
C2220 vdd.n290 gnd 0.005633f
C2221 vdd.n291 gnd 0.013317f
C2222 vdd.n292 gnd 0.002453f
C2223 vdd.n293 gnd 0.002383f
C2224 vdd.n294 gnd 0.011462f
C2225 vdd.n295 gnd 0.007751f
C2226 vdd.n296 gnd 0.054118f
C2227 vdd.n297 gnd 0.211067f
C2228 vdd.n298 gnd 0.006693f
C2229 vdd.n299 gnd 0.008708f
C2230 vdd.n300 gnd 0.007009f
C2231 vdd.n301 gnd 0.007009f
C2232 vdd.n302 gnd 0.008708f
C2233 vdd.n303 gnd 0.008708f
C2234 vdd.n304 gnd 0.636297f
C2235 vdd.n305 gnd 0.008708f
C2236 vdd.n306 gnd 0.008708f
C2237 vdd.n307 gnd 0.008708f
C2238 vdd.n308 gnd 0.689692f
C2239 vdd.n309 gnd 0.008708f
C2240 vdd.n310 gnd 0.008708f
C2241 vdd.n311 gnd 0.008708f
C2242 vdd.n312 gnd 0.008708f
C2243 vdd.n313 gnd 0.007009f
C2244 vdd.n314 gnd 0.008708f
C2245 vdd.t80 gnd 0.444963f
C2246 vdd.n315 gnd 0.008708f
C2247 vdd.n316 gnd 0.008708f
C2248 vdd.n317 gnd 0.008708f
C2249 vdd.n318 gnd 0.889925f
C2250 vdd.n319 gnd 0.008708f
C2251 vdd.n320 gnd 0.008708f
C2252 vdd.n321 gnd 0.008708f
C2253 vdd.n322 gnd 0.008708f
C2254 vdd.n323 gnd 0.008708f
C2255 vdd.n324 gnd 0.007009f
C2256 vdd.n325 gnd 0.008708f
C2257 vdd.n326 gnd 0.008708f
C2258 vdd.n327 gnd 0.008708f
C2259 vdd.n328 gnd 0.021222f
C2260 vdd.n329 gnd 2.12692f
C2261 vdd.n330 gnd 0.021709f
C2262 vdd.n331 gnd 0.008708f
C2263 vdd.n332 gnd 0.008708f
C2264 vdd.n334 gnd 0.008708f
C2265 vdd.n335 gnd 0.008708f
C2266 vdd.n336 gnd 0.007009f
C2267 vdd.n337 gnd 0.007009f
C2268 vdd.n338 gnd 0.008708f
C2269 vdd.n339 gnd 0.008708f
C2270 vdd.n340 gnd 0.008708f
C2271 vdd.n341 gnd 0.008708f
C2272 vdd.n342 gnd 0.008708f
C2273 vdd.n343 gnd 0.008708f
C2274 vdd.n344 gnd 0.007009f
C2275 vdd.n346 gnd 0.008708f
C2276 vdd.n347 gnd 0.008708f
C2277 vdd.n348 gnd 0.008708f
C2278 vdd.n349 gnd 0.008708f
C2279 vdd.n350 gnd 0.008708f
C2280 vdd.n351 gnd 0.007009f
C2281 vdd.n353 gnd 0.008708f
C2282 vdd.n354 gnd 0.008708f
C2283 vdd.n355 gnd 0.008708f
C2284 vdd.n356 gnd 0.008708f
C2285 vdd.n357 gnd 0.008708f
C2286 vdd.n358 gnd 0.007009f
C2287 vdd.n360 gnd 0.008708f
C2288 vdd.n361 gnd 0.008708f
C2289 vdd.n362 gnd 0.008708f
C2290 vdd.n363 gnd 0.008708f
C2291 vdd.n364 gnd 0.005852f
C2292 vdd.t9 gnd 0.107132f
C2293 vdd.t8 gnd 0.114495f
C2294 vdd.t6 gnd 0.139914f
C2295 vdd.n365 gnd 0.179349f
C2296 vdd.n366 gnd 0.151387f
C2297 vdd.n368 gnd 0.008708f
C2298 vdd.n369 gnd 0.008708f
C2299 vdd.n370 gnd 0.007009f
C2300 vdd.n371 gnd 0.008708f
C2301 vdd.n373 gnd 0.008708f
C2302 vdd.n374 gnd 0.008708f
C2303 vdd.n375 gnd 0.008708f
C2304 vdd.n376 gnd 0.008708f
C2305 vdd.n377 gnd 0.007009f
C2306 vdd.n379 gnd 0.008708f
C2307 vdd.n380 gnd 0.008708f
C2308 vdd.n381 gnd 0.008708f
C2309 vdd.n382 gnd 0.008708f
C2310 vdd.n383 gnd 0.008708f
C2311 vdd.n384 gnd 0.007009f
C2312 vdd.n386 gnd 0.008708f
C2313 vdd.n387 gnd 0.008708f
C2314 vdd.n388 gnd 0.008708f
C2315 vdd.n389 gnd 0.008708f
C2316 vdd.n390 gnd 0.008708f
C2317 vdd.n391 gnd 0.007009f
C2318 vdd.n393 gnd 0.008708f
C2319 vdd.n394 gnd 0.008708f
C2320 vdd.n395 gnd 0.008708f
C2321 vdd.n396 gnd 0.008708f
C2322 vdd.n397 gnd 0.008708f
C2323 vdd.n398 gnd 0.007009f
C2324 vdd.n400 gnd 0.008708f
C2325 vdd.n401 gnd 0.008708f
C2326 vdd.n402 gnd 0.008708f
C2327 vdd.n403 gnd 0.008708f
C2328 vdd.n404 gnd 0.006939f
C2329 vdd.t74 gnd 0.107132f
C2330 vdd.t73 gnd 0.114495f
C2331 vdd.t72 gnd 0.139914f
C2332 vdd.n405 gnd 0.179349f
C2333 vdd.n406 gnd 0.151387f
C2334 vdd.n408 gnd 0.008708f
C2335 vdd.n409 gnd 0.008708f
C2336 vdd.n410 gnd 0.007009f
C2337 vdd.n411 gnd 0.008708f
C2338 vdd.n413 gnd 0.008708f
C2339 vdd.n414 gnd 0.008708f
C2340 vdd.n415 gnd 0.008708f
C2341 vdd.n416 gnd 0.008708f
C2342 vdd.n417 gnd 0.007009f
C2343 vdd.n419 gnd 0.008708f
C2344 vdd.n420 gnd 0.008708f
C2345 vdd.n421 gnd 0.008708f
C2346 vdd.n422 gnd 0.008708f
C2347 vdd.n423 gnd 0.008708f
C2348 vdd.n424 gnd 0.007009f
C2349 vdd.n426 gnd 0.008708f
C2350 vdd.n427 gnd 0.008708f
C2351 vdd.n428 gnd 0.008708f
C2352 vdd.n429 gnd 0.008708f
C2353 vdd.n430 gnd 0.008708f
C2354 vdd.n431 gnd 0.007009f
C2355 vdd.n433 gnd 0.008708f
C2356 vdd.n434 gnd 0.008708f
C2357 vdd.n435 gnd 0.008708f
C2358 vdd.n436 gnd 0.008708f
C2359 vdd.n437 gnd 0.008708f
C2360 vdd.n438 gnd 0.007009f
C2361 vdd.n440 gnd 0.008708f
C2362 vdd.n441 gnd 0.008708f
C2363 vdd.n442 gnd 0.008708f
C2364 vdd.n443 gnd 0.008708f
C2365 vdd.n444 gnd 0.008708f
C2366 vdd.n445 gnd 0.008708f
C2367 vdd.n446 gnd 0.007009f
C2368 vdd.n447 gnd 0.008708f
C2369 vdd.n448 gnd 0.008708f
C2370 vdd.n449 gnd 0.007009f
C2371 vdd.n450 gnd 0.008708f
C2372 vdd.n451 gnd 0.007009f
C2373 vdd.n452 gnd 0.008708f
C2374 vdd.n453 gnd 0.007009f
C2375 vdd.n454 gnd 0.008708f
C2376 vdd.n455 gnd 0.008708f
C2377 vdd.n456 gnd 0.485009f
C2378 vdd.t82 gnd 0.444963f
C2379 vdd.n457 gnd 0.008708f
C2380 vdd.n458 gnd 0.007009f
C2381 vdd.n459 gnd 0.008708f
C2382 vdd.n460 gnd 0.007009f
C2383 vdd.n461 gnd 0.008708f
C2384 vdd.t147 gnd 0.444963f
C2385 vdd.n462 gnd 0.008708f
C2386 vdd.n463 gnd 0.007009f
C2387 vdd.n464 gnd 0.008708f
C2388 vdd.n465 gnd 0.007009f
C2389 vdd.n466 gnd 0.008708f
C2390 vdd.t162 gnd 0.444963f
C2391 vdd.n467 gnd 0.556203f
C2392 vdd.n468 gnd 0.008708f
C2393 vdd.n469 gnd 0.007009f
C2394 vdd.n470 gnd 0.008708f
C2395 vdd.n471 gnd 0.007009f
C2396 vdd.n472 gnd 0.008708f
C2397 vdd.n473 gnd 0.889925f
C2398 vdd.n474 gnd 0.008708f
C2399 vdd.n475 gnd 0.007009f
C2400 vdd.n476 gnd 0.021222f
C2401 vdd.n477 gnd 0.005817f
C2402 vdd.n478 gnd 0.021222f
C2403 vdd.t19 gnd 0.444963f
C2404 vdd.n479 gnd 0.021222f
C2405 vdd.n480 gnd 0.005817f
C2406 vdd.n481 gnd 0.007489f
C2407 vdd.n482 gnd 0.007009f
C2408 vdd.n483 gnd 0.008708f
C2409 vdd.n484 gnd 7.59106f
C2410 vdd.n515 gnd 0.021709f
C2411 vdd.n516 gnd 1.22365f
C2412 vdd.n517 gnd 0.008708f
C2413 vdd.n518 gnd 0.007009f
C2414 vdd.n519 gnd 0.005573f
C2415 vdd.n520 gnd 0.020337f
C2416 vdd.n521 gnd 0.007009f
C2417 vdd.n522 gnd 0.008708f
C2418 vdd.n523 gnd 0.008708f
C2419 vdd.n524 gnd 0.008708f
C2420 vdd.n525 gnd 0.008708f
C2421 vdd.n526 gnd 0.008708f
C2422 vdd.n527 gnd 0.008708f
C2423 vdd.n528 gnd 0.008708f
C2424 vdd.n529 gnd 0.008708f
C2425 vdd.n530 gnd 0.008708f
C2426 vdd.n531 gnd 0.008708f
C2427 vdd.n532 gnd 0.008708f
C2428 vdd.n533 gnd 0.008708f
C2429 vdd.n534 gnd 0.008708f
C2430 vdd.n535 gnd 0.008708f
C2431 vdd.n536 gnd 0.005852f
C2432 vdd.n537 gnd 0.008708f
C2433 vdd.n538 gnd 0.008708f
C2434 vdd.n539 gnd 0.008708f
C2435 vdd.n540 gnd 0.008708f
C2436 vdd.n541 gnd 0.008708f
C2437 vdd.n542 gnd 0.008708f
C2438 vdd.n543 gnd 0.008708f
C2439 vdd.n544 gnd 0.008708f
C2440 vdd.n545 gnd 0.008708f
C2441 vdd.n546 gnd 0.008708f
C2442 vdd.n547 gnd 0.008708f
C2443 vdd.n548 gnd 0.008708f
C2444 vdd.n549 gnd 0.008708f
C2445 vdd.n550 gnd 0.008708f
C2446 vdd.n551 gnd 0.008708f
C2447 vdd.n552 gnd 0.008708f
C2448 vdd.n553 gnd 0.008708f
C2449 vdd.n554 gnd 0.008708f
C2450 vdd.n555 gnd 0.008708f
C2451 vdd.n556 gnd 0.006939f
C2452 vdd.t27 gnd 0.107132f
C2453 vdd.t28 gnd 0.114495f
C2454 vdd.t26 gnd 0.139914f
C2455 vdd.n557 gnd 0.179349f
C2456 vdd.n558 gnd 0.150686f
C2457 vdd.n559 gnd 0.008708f
C2458 vdd.n560 gnd 0.008708f
C2459 vdd.n561 gnd 0.008708f
C2460 vdd.n562 gnd 0.008708f
C2461 vdd.n563 gnd 0.008708f
C2462 vdd.n564 gnd 0.008708f
C2463 vdd.n565 gnd 0.008708f
C2464 vdd.n566 gnd 0.008708f
C2465 vdd.n567 gnd 0.008708f
C2466 vdd.n568 gnd 0.008708f
C2467 vdd.n569 gnd 0.008708f
C2468 vdd.n570 gnd 0.008708f
C2469 vdd.n571 gnd 0.008708f
C2470 vdd.n572 gnd 0.005573f
C2471 vdd.n575 gnd 0.005922f
C2472 vdd.n576 gnd 0.005922f
C2473 vdd.n577 gnd 0.005922f
C2474 vdd.n578 gnd 0.005922f
C2475 vdd.n579 gnd 0.005922f
C2476 vdd.n580 gnd 0.005922f
C2477 vdd.n582 gnd 0.005922f
C2478 vdd.n583 gnd 0.005922f
C2479 vdd.n585 gnd 0.005922f
C2480 vdd.n586 gnd 0.004311f
C2481 vdd.n588 gnd 0.005922f
C2482 vdd.t13 gnd 0.239287f
C2483 vdd.t12 gnd 0.24494f
C2484 vdd.t10 gnd 0.156216f
C2485 vdd.n589 gnd 0.084426f
C2486 vdd.n590 gnd 0.047889f
C2487 vdd.n591 gnd 0.008463f
C2488 vdd.n592 gnd 0.013707f
C2489 vdd.n594 gnd 0.005922f
C2490 vdd.n595 gnd 0.605149f
C2491 vdd.n596 gnd 0.012971f
C2492 vdd.n597 gnd 0.012971f
C2493 vdd.n598 gnd 0.005922f
C2494 vdd.n599 gnd 0.01385f
C2495 vdd.n600 gnd 0.005922f
C2496 vdd.n601 gnd 0.005922f
C2497 vdd.n602 gnd 0.005922f
C2498 vdd.n603 gnd 0.005922f
C2499 vdd.n604 gnd 0.005922f
C2500 vdd.n606 gnd 0.005922f
C2501 vdd.n607 gnd 0.005922f
C2502 vdd.n609 gnd 0.005922f
C2503 vdd.n610 gnd 0.005922f
C2504 vdd.n612 gnd 0.005922f
C2505 vdd.n613 gnd 0.005922f
C2506 vdd.n615 gnd 0.005922f
C2507 vdd.n616 gnd 0.005922f
C2508 vdd.n618 gnd 0.005922f
C2509 vdd.n619 gnd 0.005922f
C2510 vdd.n621 gnd 0.005922f
C2511 vdd.t71 gnd 0.239287f
C2512 vdd.t70 gnd 0.24494f
C2513 vdd.t69 gnd 0.156216f
C2514 vdd.n622 gnd 0.084426f
C2515 vdd.n623 gnd 0.047889f
C2516 vdd.n624 gnd 0.005922f
C2517 vdd.n626 gnd 0.005922f
C2518 vdd.n627 gnd 0.005922f
C2519 vdd.t11 gnd 0.302575f
C2520 vdd.n628 gnd 0.005922f
C2521 vdd.n629 gnd 0.005922f
C2522 vdd.n630 gnd 0.005922f
C2523 vdd.n631 gnd 0.005922f
C2524 vdd.n632 gnd 0.005922f
C2525 vdd.n633 gnd 0.605149f
C2526 vdd.n634 gnd 0.005922f
C2527 vdd.n635 gnd 0.005922f
C2528 vdd.n636 gnd 0.511707f
C2529 vdd.n637 gnd 0.005922f
C2530 vdd.n638 gnd 0.005922f
C2531 vdd.n639 gnd 0.005922f
C2532 vdd.n640 gnd 0.005922f
C2533 vdd.n641 gnd 0.5918f
C2534 vdd.n642 gnd 0.005922f
C2535 vdd.n643 gnd 0.005922f
C2536 vdd.n644 gnd 0.005922f
C2537 vdd.n645 gnd 0.005922f
C2538 vdd.n646 gnd 0.005922f
C2539 vdd.n647 gnd 0.605149f
C2540 vdd.n648 gnd 0.005922f
C2541 vdd.n649 gnd 0.005922f
C2542 vdd.t127 gnd 0.302575f
C2543 vdd.n650 gnd 0.005922f
C2544 vdd.n651 gnd 0.005922f
C2545 vdd.n652 gnd 0.005922f
C2546 vdd.t102 gnd 0.302575f
C2547 vdd.n653 gnd 0.005922f
C2548 vdd.n654 gnd 0.005922f
C2549 vdd.n655 gnd 0.005922f
C2550 vdd.n656 gnd 0.005922f
C2551 vdd.n657 gnd 0.005922f
C2552 vdd.t36 gnd 0.253629f
C2553 vdd.n658 gnd 0.005922f
C2554 vdd.n659 gnd 0.005922f
C2555 vdd.n660 gnd 0.485009f
C2556 vdd.n661 gnd 0.005922f
C2557 vdd.t37 gnd 0.24494f
C2558 vdd.t35 gnd 0.156216f
C2559 vdd.t38 gnd 0.24494f
C2560 vdd.n662 gnd 0.137666f
C2561 vdd.n663 gnd 0.005922f
C2562 vdd.n664 gnd 0.005922f
C2563 vdd.n665 gnd 0.387117f
C2564 vdd.n666 gnd 0.005922f
C2565 vdd.n667 gnd 0.005922f
C2566 vdd.t104 gnd 0.088992f
C2567 vdd.n668 gnd 0.35152f
C2568 vdd.n669 gnd 0.005922f
C2569 vdd.n670 gnd 0.005922f
C2570 vdd.n671 gnd 0.005922f
C2571 vdd.n672 gnd 0.520606f
C2572 vdd.n673 gnd 0.005922f
C2573 vdd.n674 gnd 0.005922f
C2574 vdd.t114 gnd 0.302575f
C2575 vdd.n675 gnd 0.005922f
C2576 vdd.n676 gnd 0.005922f
C2577 vdd.n677 gnd 0.005922f
C2578 vdd.t110 gnd 0.302575f
C2579 vdd.n678 gnd 0.005922f
C2580 vdd.n679 gnd 0.005922f
C2581 vdd.t128 gnd 0.302575f
C2582 vdd.n680 gnd 0.005922f
C2583 vdd.n681 gnd 0.005922f
C2584 vdd.n682 gnd 0.005922f
C2585 vdd.t93 gnd 0.24028f
C2586 vdd.n683 gnd 0.005922f
C2587 vdd.n684 gnd 0.005922f
C2588 vdd.n685 gnd 0.498358f
C2589 vdd.n686 gnd 0.005922f
C2590 vdd.n687 gnd 0.005922f
C2591 vdd.n688 gnd 0.005922f
C2592 vdd.t129 gnd 0.302575f
C2593 vdd.n689 gnd 0.005922f
C2594 vdd.n690 gnd 0.005922f
C2595 vdd.t139 gnd 0.253629f
C2596 vdd.n691 gnd 0.364869f
C2597 vdd.n692 gnd 0.005922f
C2598 vdd.n693 gnd 0.005922f
C2599 vdd.n694 gnd 0.005922f
C2600 vdd.n695 gnd 0.315923f
C2601 vdd.n696 gnd 0.005922f
C2602 vdd.n697 gnd 0.005922f
C2603 vdd.t132 gnd 0.302575f
C2604 vdd.n698 gnd 0.005922f
C2605 vdd.n699 gnd 0.005922f
C2606 vdd.n700 gnd 0.005922f
C2607 vdd.n701 gnd 0.605149f
C2608 vdd.n702 gnd 0.005922f
C2609 vdd.n703 gnd 0.005922f
C2610 vdd.t99 gnd 0.204683f
C2611 vdd.t97 gnd 0.289226f
C2612 vdd.n704 gnd 0.005922f
C2613 vdd.n705 gnd 0.005922f
C2614 vdd.n706 gnd 0.005922f
C2615 vdd.n707 gnd 0.453862f
C2616 vdd.n708 gnd 0.005922f
C2617 vdd.n709 gnd 0.005922f
C2618 vdd.n710 gnd 0.005922f
C2619 vdd.n711 gnd 0.005922f
C2620 vdd.n712 gnd 0.005922f
C2621 vdd.t53 gnd 0.302575f
C2622 vdd.n713 gnd 0.005922f
C2623 vdd.n714 gnd 0.005922f
C2624 vdd.t100 gnd 0.302575f
C2625 vdd.n715 gnd 0.005922f
C2626 vdd.n716 gnd 0.012971f
C2627 vdd.n717 gnd 0.012971f
C2628 vdd.n718 gnd 0.720839f
C2629 vdd.n719 gnd 0.005922f
C2630 vdd.n720 gnd 0.005922f
C2631 vdd.t123 gnd 0.302575f
C2632 vdd.n721 gnd 0.012971f
C2633 vdd.n722 gnd 0.005922f
C2634 vdd.n723 gnd 0.005922f
C2635 vdd.t136 gnd 0.551754f
C2636 vdd.n741 gnd 0.01385f
C2637 vdd.n759 gnd 0.012971f
C2638 vdd.n760 gnd 0.005922f
C2639 vdd.n761 gnd 0.012971f
C2640 vdd.t68 gnd 0.239287f
C2641 vdd.t67 gnd 0.24494f
C2642 vdd.t66 gnd 0.156216f
C2643 vdd.n762 gnd 0.084426f
C2644 vdd.n763 gnd 0.047889f
C2645 vdd.n764 gnd 0.013707f
C2646 vdd.n765 gnd 0.005922f
C2647 vdd.n766 gnd 0.320373f
C2648 vdd.n767 gnd 0.012971f
C2649 vdd.n768 gnd 0.005922f
C2650 vdd.n769 gnd 0.01385f
C2651 vdd.n770 gnd 0.005922f
C2652 vdd.t51 gnd 0.239287f
C2653 vdd.t50 gnd 0.24494f
C2654 vdd.t48 gnd 0.156216f
C2655 vdd.n771 gnd 0.084426f
C2656 vdd.n772 gnd 0.047889f
C2657 vdd.n773 gnd 0.008463f
C2658 vdd.n774 gnd 0.005922f
C2659 vdd.n775 gnd 0.005922f
C2660 vdd.t49 gnd 0.302575f
C2661 vdd.n776 gnd 0.005922f
C2662 vdd.t134 gnd 0.302575f
C2663 vdd.n777 gnd 0.005922f
C2664 vdd.n778 gnd 0.005922f
C2665 vdd.n779 gnd 0.005922f
C2666 vdd.n780 gnd 0.005922f
C2667 vdd.n781 gnd 0.005922f
C2668 vdd.n782 gnd 0.605149f
C2669 vdd.n783 gnd 0.005922f
C2670 vdd.n784 gnd 0.005922f
C2671 vdd.t112 gnd 0.302575f
C2672 vdd.n785 gnd 0.005922f
C2673 vdd.n786 gnd 0.005922f
C2674 vdd.n787 gnd 0.005922f
C2675 vdd.n788 gnd 0.005922f
C2676 vdd.n789 gnd 0.400466f
C2677 vdd.n790 gnd 0.005922f
C2678 vdd.n791 gnd 0.005922f
C2679 vdd.n792 gnd 0.005922f
C2680 vdd.n793 gnd 0.005922f
C2681 vdd.n794 gnd 0.005922f
C2682 vdd.n795 gnd 0.533955f
C2683 vdd.n796 gnd 0.005922f
C2684 vdd.n797 gnd 0.005922f
C2685 vdd.t125 gnd 0.289226f
C2686 vdd.t94 gnd 0.204683f
C2687 vdd.n798 gnd 0.005922f
C2688 vdd.n799 gnd 0.005922f
C2689 vdd.n800 gnd 0.005922f
C2690 vdd.t117 gnd 0.302575f
C2691 vdd.n801 gnd 0.005922f
C2692 vdd.n802 gnd 0.005922f
C2693 vdd.t95 gnd 0.302575f
C2694 vdd.n803 gnd 0.005922f
C2695 vdd.n804 gnd 0.005922f
C2696 vdd.n805 gnd 0.005922f
C2697 vdd.t115 gnd 0.253629f
C2698 vdd.n806 gnd 0.005922f
C2699 vdd.n807 gnd 0.005922f
C2700 vdd.n808 gnd 0.485009f
C2701 vdd.n809 gnd 0.005922f
C2702 vdd.n810 gnd 0.005922f
C2703 vdd.n811 gnd 0.005922f
C2704 vdd.t130 gnd 0.302575f
C2705 vdd.n812 gnd 0.005922f
C2706 vdd.n813 gnd 0.005922f
C2707 vdd.t105 gnd 0.24028f
C2708 vdd.n814 gnd 0.35152f
C2709 vdd.n815 gnd 0.005922f
C2710 vdd.n816 gnd 0.005922f
C2711 vdd.n817 gnd 0.005922f
C2712 vdd.n818 gnd 0.520606f
C2713 vdd.n819 gnd 0.005922f
C2714 vdd.n820 gnd 0.005922f
C2715 vdd.t138 gnd 0.302575f
C2716 vdd.n821 gnd 0.005922f
C2717 vdd.n822 gnd 0.005922f
C2718 vdd.n823 gnd 0.005922f
C2719 vdd.n824 gnd 0.605149f
C2720 vdd.n825 gnd 0.005922f
C2721 vdd.n826 gnd 0.005922f
C2722 vdd.t109 gnd 0.302575f
C2723 vdd.n827 gnd 0.005922f
C2724 vdd.n828 gnd 0.005922f
C2725 vdd.n829 gnd 0.005922f
C2726 vdd.t103 gnd 0.088992f
C2727 vdd.n830 gnd 0.005922f
C2728 vdd.n831 gnd 0.005922f
C2729 vdd.n832 gnd 0.005922f
C2730 vdd.t58 gnd 0.24494f
C2731 vdd.t56 gnd 0.156216f
C2732 vdd.t59 gnd 0.24494f
C2733 vdd.n833 gnd 0.137666f
C2734 vdd.n834 gnd 0.005922f
C2735 vdd.n835 gnd 0.005922f
C2736 vdd.t122 gnd 0.302575f
C2737 vdd.n836 gnd 0.005922f
C2738 vdd.n837 gnd 0.005922f
C2739 vdd.t57 gnd 0.253629f
C2740 vdd.n838 gnd 0.516157f
C2741 vdd.n839 gnd 0.005922f
C2742 vdd.n840 gnd 0.005922f
C2743 vdd.n841 gnd 0.005922f
C2744 vdd.n842 gnd 0.315923f
C2745 vdd.n843 gnd 0.005922f
C2746 vdd.n844 gnd 0.005922f
C2747 vdd.n845 gnd 0.422714f
C2748 vdd.n846 gnd 0.005922f
C2749 vdd.n847 gnd 0.005922f
C2750 vdd.n848 gnd 0.005922f
C2751 vdd.n849 gnd 0.605149f
C2752 vdd.n850 gnd 0.005922f
C2753 vdd.n851 gnd 0.005922f
C2754 vdd.t106 gnd 0.302575f
C2755 vdd.n852 gnd 0.005922f
C2756 vdd.n853 gnd 0.005922f
C2757 vdd.n854 gnd 0.005922f
C2758 vdd.n855 gnd 0.605149f
C2759 vdd.n856 gnd 0.005922f
C2760 vdd.n857 gnd 0.005922f
C2761 vdd.n858 gnd 0.005922f
C2762 vdd.n859 gnd 0.005922f
C2763 vdd.n860 gnd 0.005922f
C2764 vdd.t15 gnd 0.302575f
C2765 vdd.n861 gnd 0.005922f
C2766 vdd.n862 gnd 0.005922f
C2767 vdd.n863 gnd 0.005922f
C2768 vdd.n864 gnd 0.012971f
C2769 vdd.n865 gnd 0.012971f
C2770 vdd.n866 gnd 0.854328f
C2771 vdd.n867 gnd 0.005922f
C2772 vdd.n868 gnd 0.005922f
C2773 vdd.n869 gnd 0.396017f
C2774 vdd.n870 gnd 0.012971f
C2775 vdd.n871 gnd 0.005922f
C2776 vdd.n872 gnd 0.005922f
C2777 vdd.n873 gnd 7.92923f
C2778 vdd.n906 gnd 0.01385f
C2779 vdd.n907 gnd 0.005922f
C2780 vdd.n908 gnd 0.005922f
C2781 vdd.n909 gnd 0.005922f
C2782 vdd.n910 gnd 0.005573f
C2783 vdd.n913 gnd 0.021709f
C2784 vdd.n914 gnd 0.005817f
C2785 vdd.n915 gnd 0.007009f
C2786 vdd.n917 gnd 0.008708f
C2787 vdd.n918 gnd 0.008708f
C2788 vdd.n919 gnd 0.007009f
C2789 vdd.n921 gnd 0.008708f
C2790 vdd.n922 gnd 0.008708f
C2791 vdd.n923 gnd 0.008708f
C2792 vdd.n924 gnd 0.008708f
C2793 vdd.n925 gnd 0.008708f
C2794 vdd.n926 gnd 0.007009f
C2795 vdd.n928 gnd 0.008708f
C2796 vdd.n929 gnd 0.008708f
C2797 vdd.n930 gnd 0.008708f
C2798 vdd.n931 gnd 0.008708f
C2799 vdd.n932 gnd 0.008708f
C2800 vdd.n933 gnd 0.007009f
C2801 vdd.n935 gnd 0.008708f
C2802 vdd.n936 gnd 0.008708f
C2803 vdd.n937 gnd 0.008708f
C2804 vdd.n938 gnd 0.008708f
C2805 vdd.n939 gnd 0.005852f
C2806 vdd.t65 gnd 0.107132f
C2807 vdd.t64 gnd 0.114495f
C2808 vdd.t63 gnd 0.139914f
C2809 vdd.n940 gnd 0.179349f
C2810 vdd.n941 gnd 0.150686f
C2811 vdd.n943 gnd 0.008708f
C2812 vdd.n944 gnd 0.008708f
C2813 vdd.n945 gnd 0.007009f
C2814 vdd.n946 gnd 0.008708f
C2815 vdd.n948 gnd 0.008708f
C2816 vdd.n949 gnd 0.008708f
C2817 vdd.n950 gnd 0.008708f
C2818 vdd.n951 gnd 0.008708f
C2819 vdd.n952 gnd 0.007009f
C2820 vdd.n954 gnd 0.008708f
C2821 vdd.n955 gnd 0.008708f
C2822 vdd.n956 gnd 0.008708f
C2823 vdd.n957 gnd 0.008708f
C2824 vdd.n958 gnd 0.008708f
C2825 vdd.n959 gnd 0.007009f
C2826 vdd.n961 gnd 0.008708f
C2827 vdd.n962 gnd 0.008708f
C2828 vdd.n963 gnd 0.008708f
C2829 vdd.n964 gnd 0.008708f
C2830 vdd.n965 gnd 0.008708f
C2831 vdd.n966 gnd 0.007009f
C2832 vdd.n968 gnd 0.008708f
C2833 vdd.n969 gnd 0.008708f
C2834 vdd.n970 gnd 0.008708f
C2835 vdd.n971 gnd 0.008708f
C2836 vdd.n972 gnd 0.008708f
C2837 vdd.n973 gnd 0.007009f
C2838 vdd.n975 gnd 0.008708f
C2839 vdd.n976 gnd 0.008708f
C2840 vdd.n977 gnd 0.008708f
C2841 vdd.n978 gnd 0.008708f
C2842 vdd.n979 gnd 0.006939f
C2843 vdd.t47 gnd 0.107132f
C2844 vdd.t46 gnd 0.114495f
C2845 vdd.t45 gnd 0.139914f
C2846 vdd.n980 gnd 0.179349f
C2847 vdd.n981 gnd 0.150686f
C2848 vdd.n983 gnd 0.008708f
C2849 vdd.n984 gnd 0.008708f
C2850 vdd.n985 gnd 0.007009f
C2851 vdd.n986 gnd 0.008708f
C2852 vdd.n988 gnd 0.008708f
C2853 vdd.n989 gnd 0.008708f
C2854 vdd.n990 gnd 0.008708f
C2855 vdd.n991 gnd 0.008708f
C2856 vdd.n992 gnd 0.007009f
C2857 vdd.n994 gnd 0.008708f
C2858 vdd.n995 gnd 0.008708f
C2859 vdd.n996 gnd 0.008708f
C2860 vdd.n997 gnd 0.008708f
C2861 vdd.n998 gnd 0.008708f
C2862 vdd.n999 gnd 0.007009f
C2863 vdd.n1001 gnd 0.008708f
C2864 vdd.n1002 gnd 0.008708f
C2865 vdd.n1003 gnd 0.008708f
C2866 vdd.n1004 gnd 0.008708f
C2867 vdd.n1005 gnd 0.008708f
C2868 vdd.n1006 gnd 0.007009f
C2869 vdd.n1008 gnd 0.008708f
C2870 vdd.n1009 gnd 0.008708f
C2871 vdd.n1010 gnd 0.005573f
C2872 vdd.n1011 gnd 0.007009f
C2873 vdd.n1012 gnd 0.005922f
C2874 vdd.n1013 gnd 0.005922f
C2875 vdd.n1014 gnd 0.005922f
C2876 vdd.n1015 gnd 0.005922f
C2877 vdd.n1016 gnd 0.005922f
C2878 vdd.n1017 gnd 0.005922f
C2879 vdd.n1018 gnd 0.005922f
C2880 vdd.n1019 gnd 0.005922f
C2881 vdd.n1020 gnd 0.005922f
C2882 vdd.n1021 gnd 0.005922f
C2883 vdd.n1022 gnd 0.005922f
C2884 vdd.n1023 gnd 0.005922f
C2885 vdd.n1024 gnd 0.005922f
C2886 vdd.n1025 gnd 0.005922f
C2887 vdd.n1026 gnd 0.005922f
C2888 vdd.n1027 gnd 0.005922f
C2889 vdd.n1028 gnd 0.005922f
C2890 vdd.n1029 gnd 0.005922f
C2891 vdd.n1030 gnd 0.005922f
C2892 vdd.n1031 gnd 0.005922f
C2893 vdd.n1032 gnd 0.005922f
C2894 vdd.n1033 gnd 0.005922f
C2895 vdd.n1034 gnd 0.005922f
C2896 vdd.n1035 gnd 0.005922f
C2897 vdd.n1036 gnd 0.005922f
C2898 vdd.n1037 gnd 0.005922f
C2899 vdd.n1038 gnd 0.005922f
C2900 vdd.n1039 gnd 0.005922f
C2901 vdd.n1040 gnd 0.005922f
C2902 vdd.n1041 gnd 0.005922f
C2903 vdd.n1042 gnd 0.005922f
C2904 vdd.t16 gnd 0.239287f
C2905 vdd.t17 gnd 0.24494f
C2906 vdd.t14 gnd 0.156216f
C2907 vdd.n1043 gnd 0.084426f
C2908 vdd.n1044 gnd 0.047889f
C2909 vdd.n1045 gnd 0.008463f
C2910 vdd.n1046 gnd 0.005922f
C2911 vdd.n1047 gnd 0.005922f
C2912 vdd.n1048 gnd 0.005922f
C2913 vdd.n1049 gnd 0.005922f
C2914 vdd.n1050 gnd 0.005922f
C2915 vdd.n1051 gnd 0.005922f
C2916 vdd.n1052 gnd 0.005922f
C2917 vdd.n1053 gnd 0.005922f
C2918 vdd.n1054 gnd 0.005922f
C2919 vdd.n1055 gnd 0.005922f
C2920 vdd.n1056 gnd 0.005922f
C2921 vdd.n1057 gnd 0.005922f
C2922 vdd.n1058 gnd 0.005922f
C2923 vdd.n1059 gnd 0.005922f
C2924 vdd.n1060 gnd 0.005922f
C2925 vdd.n1061 gnd 0.005922f
C2926 vdd.n1062 gnd 0.005922f
C2927 vdd.t30 gnd 0.239287f
C2928 vdd.t31 gnd 0.24494f
C2929 vdd.t29 gnd 0.156216f
C2930 vdd.n1063 gnd 0.084426f
C2931 vdd.n1064 gnd 0.047889f
C2932 vdd.n1065 gnd 0.005922f
C2933 vdd.n1066 gnd 0.005922f
C2934 vdd.n1067 gnd 0.005922f
C2935 vdd.n1068 gnd 0.005922f
C2936 vdd.n1069 gnd 0.005922f
C2937 vdd.n1070 gnd 0.005922f
C2938 vdd.n1071 gnd 0.005922f
C2939 vdd.n1072 gnd 0.005922f
C2940 vdd.n1073 gnd 0.005922f
C2941 vdd.n1074 gnd 0.005922f
C2942 vdd.n1075 gnd 0.005922f
C2943 vdd.n1076 gnd 0.005922f
C2944 vdd.n1077 gnd 0.005922f
C2945 vdd.n1078 gnd 0.005922f
C2946 vdd.n1079 gnd 0.005922f
C2947 vdd.n1080 gnd 0.005922f
C2948 vdd.n1081 gnd 0.005922f
C2949 vdd.n1082 gnd 0.005922f
C2950 vdd.n1083 gnd 0.005922f
C2951 vdd.n1084 gnd 0.005922f
C2952 vdd.n1085 gnd 0.005922f
C2953 vdd.n1086 gnd 0.005922f
C2954 vdd.n1087 gnd 0.005922f
C2955 vdd.n1088 gnd 0.005922f
C2956 vdd.n1089 gnd 0.005922f
C2957 vdd.n1090 gnd 0.005922f
C2958 vdd.n1091 gnd 0.004311f
C2959 vdd.n1092 gnd 0.008463f
C2960 vdd.n1093 gnd 0.004572f
C2961 vdd.n1094 gnd 0.005922f
C2962 vdd.n1095 gnd 0.005922f
C2963 vdd.n1096 gnd 0.005922f
C2964 vdd.n1097 gnd 0.01385f
C2965 vdd.n1098 gnd 0.01385f
C2966 vdd.n1099 gnd 0.012971f
C2967 vdd.n1100 gnd 0.012971f
C2968 vdd.n1101 gnd 0.005922f
C2969 vdd.n1102 gnd 0.005922f
C2970 vdd.n1103 gnd 0.005922f
C2971 vdd.n1104 gnd 0.005922f
C2972 vdd.n1105 gnd 0.005922f
C2973 vdd.n1106 gnd 0.005922f
C2974 vdd.n1107 gnd 0.005922f
C2975 vdd.n1108 gnd 0.005922f
C2976 vdd.n1109 gnd 0.005922f
C2977 vdd.n1110 gnd 0.005922f
C2978 vdd.n1111 gnd 0.005922f
C2979 vdd.n1112 gnd 0.005922f
C2980 vdd.n1113 gnd 0.005922f
C2981 vdd.n1114 gnd 0.005922f
C2982 vdd.n1115 gnd 0.005922f
C2983 vdd.n1116 gnd 0.005922f
C2984 vdd.n1117 gnd 0.005922f
C2985 vdd.n1118 gnd 0.005922f
C2986 vdd.n1119 gnd 0.005922f
C2987 vdd.n1120 gnd 0.005922f
C2988 vdd.n1121 gnd 0.005922f
C2989 vdd.n1122 gnd 0.005922f
C2990 vdd.n1123 gnd 0.005922f
C2991 vdd.n1124 gnd 0.005922f
C2992 vdd.n1125 gnd 0.005922f
C2993 vdd.n1126 gnd 0.005922f
C2994 vdd.n1127 gnd 0.005922f
C2995 vdd.n1128 gnd 0.36042f
C2996 vdd.n1129 gnd 0.005922f
C2997 vdd.n1130 gnd 0.005922f
C2998 vdd.n1131 gnd 0.005922f
C2999 vdd.n1132 gnd 0.005922f
C3000 vdd.n1133 gnd 0.005922f
C3001 vdd.n1134 gnd 0.005922f
C3002 vdd.n1135 gnd 0.005922f
C3003 vdd.n1136 gnd 0.005922f
C3004 vdd.n1137 gnd 0.005922f
C3005 vdd.n1138 gnd 0.005922f
C3006 vdd.n1139 gnd 0.005922f
C3007 vdd.n1140 gnd 0.005922f
C3008 vdd.n1141 gnd 0.005922f
C3009 vdd.n1142 gnd 0.005922f
C3010 vdd.n1143 gnd 0.005922f
C3011 vdd.n1144 gnd 0.005922f
C3012 vdd.n1145 gnd 0.005922f
C3013 vdd.n1146 gnd 0.005922f
C3014 vdd.n1147 gnd 0.005922f
C3015 vdd.n1148 gnd 0.005922f
C3016 vdd.n1149 gnd 0.191334f
C3017 vdd.n1150 gnd 0.005922f
C3018 vdd.n1151 gnd 0.005922f
C3019 vdd.n1152 gnd 0.005922f
C3020 vdd.n1153 gnd 0.005922f
C3021 vdd.n1154 gnd 0.005922f
C3022 vdd.n1155 gnd 0.005922f
C3023 vdd.n1156 gnd 0.005922f
C3024 vdd.n1157 gnd 0.005922f
C3025 vdd.n1158 gnd 0.005922f
C3026 vdd.n1159 gnd 0.005922f
C3027 vdd.n1160 gnd 0.005922f
C3028 vdd.n1161 gnd 0.005922f
C3029 vdd.n1162 gnd 0.005922f
C3030 vdd.n1163 gnd 0.005922f
C3031 vdd.n1164 gnd 0.005922f
C3032 vdd.n1165 gnd 0.005922f
C3033 vdd.n1166 gnd 0.005922f
C3034 vdd.n1167 gnd 0.005922f
C3035 vdd.n1168 gnd 0.005922f
C3036 vdd.n1169 gnd 0.005922f
C3037 vdd.n1170 gnd 0.005922f
C3038 vdd.n1171 gnd 0.005922f
C3039 vdd.n1172 gnd 0.005922f
C3040 vdd.n1173 gnd 0.005922f
C3041 vdd.n1174 gnd 0.005922f
C3042 vdd.n1175 gnd 0.005922f
C3043 vdd.n1176 gnd 0.005922f
C3044 vdd.n1177 gnd 0.012971f
C3045 vdd.n1178 gnd 0.012971f
C3046 vdd.n1179 gnd 0.01385f
C3047 vdd.n1180 gnd 0.005922f
C3048 vdd.n1181 gnd 0.005922f
C3049 vdd.n1182 gnd 0.004572f
C3050 vdd.n1183 gnd 0.005922f
C3051 vdd.n1184 gnd 0.005922f
C3052 vdd.n1185 gnd 0.004311f
C3053 vdd.n1186 gnd 0.005922f
C3054 vdd.n1187 gnd 0.005922f
C3055 vdd.n1188 gnd 0.005922f
C3056 vdd.n1189 gnd 0.005922f
C3057 vdd.n1190 gnd 0.005922f
C3058 vdd.n1191 gnd 0.005922f
C3059 vdd.n1192 gnd 0.005922f
C3060 vdd.n1193 gnd 0.005922f
C3061 vdd.n1194 gnd 0.005922f
C3062 vdd.n1195 gnd 0.005922f
C3063 vdd.n1196 gnd 0.005922f
C3064 vdd.n1197 gnd 0.005922f
C3065 vdd.n1198 gnd 0.005922f
C3066 vdd.n1199 gnd 0.005922f
C3067 vdd.n1200 gnd 0.005922f
C3068 vdd.n1201 gnd 0.005922f
C3069 vdd.n1202 gnd 0.005922f
C3070 vdd.n1203 gnd 0.005922f
C3071 vdd.n1204 gnd 0.005922f
C3072 vdd.n1205 gnd 0.005922f
C3073 vdd.n1206 gnd 0.005922f
C3074 vdd.n1207 gnd 0.005922f
C3075 vdd.n1208 gnd 0.005922f
C3076 vdd.n1209 gnd 0.005922f
C3077 vdd.n1210 gnd 0.005922f
C3078 vdd.n1211 gnd 0.005922f
C3079 vdd.n1212 gnd 0.023733f
C3080 vdd.n1214 gnd 0.021709f
C3081 vdd.n1215 gnd 0.007009f
C3082 vdd.n1217 gnd 0.008708f
C3083 vdd.n1218 gnd 0.007009f
C3084 vdd.n1219 gnd 0.008708f
C3085 vdd.n1221 gnd 0.008708f
C3086 vdd.n1222 gnd 0.008708f
C3087 vdd.n1224 gnd 0.008708f
C3088 vdd.n1225 gnd 0.005817f
C3089 vdd.t23 gnd 0.444963f
C3090 vdd.n1226 gnd 0.008708f
C3091 vdd.n1227 gnd 0.021709f
C3092 vdd.n1228 gnd 0.007009f
C3093 vdd.n1229 gnd 0.008708f
C3094 vdd.n1230 gnd 0.007009f
C3095 vdd.n1231 gnd 0.008708f
C3096 vdd.n1232 gnd 0.889925f
C3097 vdd.n1233 gnd 0.008708f
C3098 vdd.n1234 gnd 0.007009f
C3099 vdd.n1235 gnd 0.007009f
C3100 vdd.n1236 gnd 0.008708f
C3101 vdd.n1237 gnd 0.007009f
C3102 vdd.n1238 gnd 0.008708f
C3103 vdd.t141 gnd 0.444963f
C3104 vdd.n1239 gnd 0.008708f
C3105 vdd.n1240 gnd 0.007009f
C3106 vdd.n1241 gnd 0.008708f
C3107 vdd.n1242 gnd 0.007009f
C3108 vdd.n1243 gnd 0.008708f
C3109 vdd.t86 gnd 0.444963f
C3110 vdd.n1244 gnd 0.008708f
C3111 vdd.n1245 gnd 0.007009f
C3112 vdd.n1246 gnd 0.008708f
C3113 vdd.n1247 gnd 0.007009f
C3114 vdd.n1248 gnd 0.008708f
C3115 vdd.n1249 gnd 0.698591f
C3116 vdd.n1250 gnd 0.738638f
C3117 vdd.t166 gnd 0.444963f
C3118 vdd.n1251 gnd 0.008708f
C3119 vdd.n1252 gnd 0.007009f
C3120 vdd.n1253 gnd 0.004779f
C3121 vdd.n1254 gnd 0.004435f
C3122 vdd.n1255 gnd 0.002453f
C3123 vdd.n1256 gnd 0.005633f
C3124 vdd.n1257 gnd 0.002383f
C3125 vdd.n1258 gnd 0.002523f
C3126 vdd.n1259 gnd 0.004435f
C3127 vdd.n1260 gnd 0.002383f
C3128 vdd.n1261 gnd 0.005633f
C3129 vdd.n1262 gnd 0.002523f
C3130 vdd.n1263 gnd 0.004435f
C3131 vdd.n1264 gnd 0.002383f
C3132 vdd.n1265 gnd 0.004224f
C3133 vdd.n1266 gnd 0.004237f
C3134 vdd.t171 gnd 0.012101f
C3135 vdd.n1267 gnd 0.026925f
C3136 vdd.n1268 gnd 0.140125f
C3137 vdd.n1269 gnd 0.002383f
C3138 vdd.n1270 gnd 0.002523f
C3139 vdd.n1271 gnd 0.005633f
C3140 vdd.n1272 gnd 0.005633f
C3141 vdd.n1273 gnd 0.002523f
C3142 vdd.n1274 gnd 0.002383f
C3143 vdd.n1275 gnd 0.004435f
C3144 vdd.n1276 gnd 0.004435f
C3145 vdd.n1277 gnd 0.002383f
C3146 vdd.n1278 gnd 0.002523f
C3147 vdd.n1279 gnd 0.005633f
C3148 vdd.n1280 gnd 0.005633f
C3149 vdd.n1281 gnd 0.002523f
C3150 vdd.n1282 gnd 0.002383f
C3151 vdd.n1283 gnd 0.004435f
C3152 vdd.n1284 gnd 0.004435f
C3153 vdd.n1285 gnd 0.002383f
C3154 vdd.n1286 gnd 0.002523f
C3155 vdd.n1287 gnd 0.005633f
C3156 vdd.n1288 gnd 0.005633f
C3157 vdd.n1289 gnd 0.013317f
C3158 vdd.n1290 gnd 0.002453f
C3159 vdd.n1291 gnd 0.002383f
C3160 vdd.n1292 gnd 0.011462f
C3161 vdd.n1293 gnd 0.008002f
C3162 vdd.t183 gnd 0.028036f
C3163 vdd.t189 gnd 0.028036f
C3164 vdd.n1294 gnd 0.192681f
C3165 vdd.n1295 gnd 0.151515f
C3166 vdd.t168 gnd 0.028036f
C3167 vdd.t176 gnd 0.028036f
C3168 vdd.n1296 gnd 0.192681f
C3169 vdd.n1297 gnd 0.122271f
C3170 vdd.t92 gnd 0.028036f
C3171 vdd.t195 gnd 0.028036f
C3172 vdd.n1298 gnd 0.192681f
C3173 vdd.n1299 gnd 0.122271f
C3174 vdd.n1300 gnd 0.004779f
C3175 vdd.n1301 gnd 0.004435f
C3176 vdd.n1302 gnd 0.002453f
C3177 vdd.n1303 gnd 0.005633f
C3178 vdd.n1304 gnd 0.002383f
C3179 vdd.n1305 gnd 0.002523f
C3180 vdd.n1306 gnd 0.004435f
C3181 vdd.n1307 gnd 0.002383f
C3182 vdd.n1308 gnd 0.005633f
C3183 vdd.n1309 gnd 0.002523f
C3184 vdd.n1310 gnd 0.004435f
C3185 vdd.n1311 gnd 0.002383f
C3186 vdd.n1312 gnd 0.004224f
C3187 vdd.n1313 gnd 0.004237f
C3188 vdd.t180 gnd 0.012101f
C3189 vdd.n1314 gnd 0.026925f
C3190 vdd.n1315 gnd 0.140125f
C3191 vdd.n1316 gnd 0.002383f
C3192 vdd.n1317 gnd 0.002523f
C3193 vdd.n1318 gnd 0.005633f
C3194 vdd.n1319 gnd 0.005633f
C3195 vdd.n1320 gnd 0.002523f
C3196 vdd.n1321 gnd 0.002383f
C3197 vdd.n1322 gnd 0.004435f
C3198 vdd.n1323 gnd 0.004435f
C3199 vdd.n1324 gnd 0.002383f
C3200 vdd.n1325 gnd 0.002523f
C3201 vdd.n1326 gnd 0.005633f
C3202 vdd.n1327 gnd 0.005633f
C3203 vdd.n1328 gnd 0.002523f
C3204 vdd.n1329 gnd 0.002383f
C3205 vdd.n1330 gnd 0.004435f
C3206 vdd.n1331 gnd 0.004435f
C3207 vdd.n1332 gnd 0.002383f
C3208 vdd.n1333 gnd 0.002523f
C3209 vdd.n1334 gnd 0.005633f
C3210 vdd.n1335 gnd 0.005633f
C3211 vdd.n1336 gnd 0.013317f
C3212 vdd.n1337 gnd 0.002453f
C3213 vdd.n1338 gnd 0.002383f
C3214 vdd.n1339 gnd 0.011462f
C3215 vdd.n1340 gnd 0.007751f
C3216 vdd.n1341 gnd 0.090971f
C3217 vdd.n1342 gnd 0.004779f
C3218 vdd.n1343 gnd 0.004435f
C3219 vdd.n1344 gnd 0.002453f
C3220 vdd.n1345 gnd 0.005633f
C3221 vdd.n1346 gnd 0.002383f
C3222 vdd.n1347 gnd 0.002523f
C3223 vdd.n1348 gnd 0.004435f
C3224 vdd.n1349 gnd 0.002383f
C3225 vdd.n1350 gnd 0.005633f
C3226 vdd.n1351 gnd 0.002523f
C3227 vdd.n1352 gnd 0.004435f
C3228 vdd.n1353 gnd 0.002383f
C3229 vdd.n1354 gnd 0.004224f
C3230 vdd.n1355 gnd 0.004237f
C3231 vdd.t142 gnd 0.012101f
C3232 vdd.n1356 gnd 0.026925f
C3233 vdd.n1357 gnd 0.140125f
C3234 vdd.n1358 gnd 0.002383f
C3235 vdd.n1359 gnd 0.002523f
C3236 vdd.n1360 gnd 0.005633f
C3237 vdd.n1361 gnd 0.005633f
C3238 vdd.n1362 gnd 0.002523f
C3239 vdd.n1363 gnd 0.002383f
C3240 vdd.n1364 gnd 0.004435f
C3241 vdd.n1365 gnd 0.004435f
C3242 vdd.n1366 gnd 0.002383f
C3243 vdd.n1367 gnd 0.002523f
C3244 vdd.n1368 gnd 0.005633f
C3245 vdd.n1369 gnd 0.005633f
C3246 vdd.n1370 gnd 0.002523f
C3247 vdd.n1371 gnd 0.002383f
C3248 vdd.n1372 gnd 0.004435f
C3249 vdd.n1373 gnd 0.004435f
C3250 vdd.n1374 gnd 0.002383f
C3251 vdd.n1375 gnd 0.002523f
C3252 vdd.n1376 gnd 0.005633f
C3253 vdd.n1377 gnd 0.005633f
C3254 vdd.n1378 gnd 0.013317f
C3255 vdd.n1379 gnd 0.002453f
C3256 vdd.n1380 gnd 0.002383f
C3257 vdd.n1381 gnd 0.011462f
C3258 vdd.n1382 gnd 0.008002f
C3259 vdd.t198 gnd 0.028036f
C3260 vdd.t87 gnd 0.028036f
C3261 vdd.n1383 gnd 0.192681f
C3262 vdd.n1384 gnd 0.151515f
C3263 vdd.t199 gnd 0.028036f
C3264 vdd.t149 gnd 0.028036f
C3265 vdd.n1385 gnd 0.192681f
C3266 vdd.n1386 gnd 0.122271f
C3267 vdd.t169 gnd 0.028036f
C3268 vdd.t194 gnd 0.028036f
C3269 vdd.n1387 gnd 0.192681f
C3270 vdd.n1388 gnd 0.122271f
C3271 vdd.n1389 gnd 0.004779f
C3272 vdd.n1390 gnd 0.004435f
C3273 vdd.n1391 gnd 0.002453f
C3274 vdd.n1392 gnd 0.005633f
C3275 vdd.n1393 gnd 0.002383f
C3276 vdd.n1394 gnd 0.002523f
C3277 vdd.n1395 gnd 0.004435f
C3278 vdd.n1396 gnd 0.002383f
C3279 vdd.n1397 gnd 0.005633f
C3280 vdd.n1398 gnd 0.002523f
C3281 vdd.n1399 gnd 0.004435f
C3282 vdd.n1400 gnd 0.002383f
C3283 vdd.n1401 gnd 0.004224f
C3284 vdd.n1402 gnd 0.004237f
C3285 vdd.t150 gnd 0.012101f
C3286 vdd.n1403 gnd 0.026925f
C3287 vdd.n1404 gnd 0.140125f
C3288 vdd.n1405 gnd 0.002383f
C3289 vdd.n1406 gnd 0.002523f
C3290 vdd.n1407 gnd 0.005633f
C3291 vdd.n1408 gnd 0.005633f
C3292 vdd.n1409 gnd 0.002523f
C3293 vdd.n1410 gnd 0.002383f
C3294 vdd.n1411 gnd 0.004435f
C3295 vdd.n1412 gnd 0.004435f
C3296 vdd.n1413 gnd 0.002383f
C3297 vdd.n1414 gnd 0.002523f
C3298 vdd.n1415 gnd 0.005633f
C3299 vdd.n1416 gnd 0.005633f
C3300 vdd.n1417 gnd 0.002523f
C3301 vdd.n1418 gnd 0.002383f
C3302 vdd.n1419 gnd 0.004435f
C3303 vdd.n1420 gnd 0.004435f
C3304 vdd.n1421 gnd 0.002383f
C3305 vdd.n1422 gnd 0.002523f
C3306 vdd.n1423 gnd 0.005633f
C3307 vdd.n1424 gnd 0.005633f
C3308 vdd.n1425 gnd 0.013317f
C3309 vdd.n1426 gnd 0.002453f
C3310 vdd.n1427 gnd 0.002383f
C3311 vdd.n1428 gnd 0.011462f
C3312 vdd.n1429 gnd 0.007751f
C3313 vdd.n1430 gnd 0.054118f
C3314 vdd.n1431 gnd 0.195002f
C3315 vdd.n1432 gnd 0.004779f
C3316 vdd.n1433 gnd 0.004435f
C3317 vdd.n1434 gnd 0.002453f
C3318 vdd.n1435 gnd 0.005633f
C3319 vdd.n1436 gnd 0.002383f
C3320 vdd.n1437 gnd 0.002523f
C3321 vdd.n1438 gnd 0.004435f
C3322 vdd.n1439 gnd 0.002383f
C3323 vdd.n1440 gnd 0.005633f
C3324 vdd.n1441 gnd 0.002523f
C3325 vdd.n1442 gnd 0.004435f
C3326 vdd.n1443 gnd 0.002383f
C3327 vdd.n1444 gnd 0.004224f
C3328 vdd.n1445 gnd 0.004237f
C3329 vdd.t200 gnd 0.012101f
C3330 vdd.n1446 gnd 0.026925f
C3331 vdd.n1447 gnd 0.140125f
C3332 vdd.n1448 gnd 0.002383f
C3333 vdd.n1449 gnd 0.002523f
C3334 vdd.n1450 gnd 0.005633f
C3335 vdd.n1451 gnd 0.005633f
C3336 vdd.n1452 gnd 0.002523f
C3337 vdd.n1453 gnd 0.002383f
C3338 vdd.n1454 gnd 0.004435f
C3339 vdd.n1455 gnd 0.004435f
C3340 vdd.n1456 gnd 0.002383f
C3341 vdd.n1457 gnd 0.002523f
C3342 vdd.n1458 gnd 0.005633f
C3343 vdd.n1459 gnd 0.005633f
C3344 vdd.n1460 gnd 0.002523f
C3345 vdd.n1461 gnd 0.002383f
C3346 vdd.n1462 gnd 0.004435f
C3347 vdd.n1463 gnd 0.004435f
C3348 vdd.n1464 gnd 0.002383f
C3349 vdd.n1465 gnd 0.002523f
C3350 vdd.n1466 gnd 0.005633f
C3351 vdd.n1467 gnd 0.005633f
C3352 vdd.n1468 gnd 0.013317f
C3353 vdd.n1469 gnd 0.002453f
C3354 vdd.n1470 gnd 0.002383f
C3355 vdd.n1471 gnd 0.011462f
C3356 vdd.n1472 gnd 0.008002f
C3357 vdd.t167 gnd 0.028036f
C3358 vdd.t201 gnd 0.028036f
C3359 vdd.n1473 gnd 0.192681f
C3360 vdd.n1474 gnd 0.151515f
C3361 vdd.t159 gnd 0.028036f
C3362 vdd.t144 gnd 0.028036f
C3363 vdd.n1475 gnd 0.192681f
C3364 vdd.n1476 gnd 0.122271f
C3365 vdd.t182 gnd 0.028036f
C3366 vdd.t90 gnd 0.028036f
C3367 vdd.n1477 gnd 0.192681f
C3368 vdd.n1478 gnd 0.122271f
C3369 vdd.n1479 gnd 0.004779f
C3370 vdd.n1480 gnd 0.004435f
C3371 vdd.n1481 gnd 0.002453f
C3372 vdd.n1482 gnd 0.005633f
C3373 vdd.n1483 gnd 0.002383f
C3374 vdd.n1484 gnd 0.002523f
C3375 vdd.n1485 gnd 0.004435f
C3376 vdd.n1486 gnd 0.002383f
C3377 vdd.n1487 gnd 0.005633f
C3378 vdd.n1488 gnd 0.002523f
C3379 vdd.n1489 gnd 0.004435f
C3380 vdd.n1490 gnd 0.002383f
C3381 vdd.n1491 gnd 0.004224f
C3382 vdd.n1492 gnd 0.004237f
C3383 vdd.t146 gnd 0.012101f
C3384 vdd.n1493 gnd 0.026925f
C3385 vdd.n1494 gnd 0.140125f
C3386 vdd.n1495 gnd 0.002383f
C3387 vdd.n1496 gnd 0.002523f
C3388 vdd.n1497 gnd 0.005633f
C3389 vdd.n1498 gnd 0.005633f
C3390 vdd.n1499 gnd 0.002523f
C3391 vdd.n1500 gnd 0.002383f
C3392 vdd.n1501 gnd 0.004435f
C3393 vdd.n1502 gnd 0.004435f
C3394 vdd.n1503 gnd 0.002383f
C3395 vdd.n1504 gnd 0.002523f
C3396 vdd.n1505 gnd 0.005633f
C3397 vdd.n1506 gnd 0.005633f
C3398 vdd.n1507 gnd 0.002523f
C3399 vdd.n1508 gnd 0.002383f
C3400 vdd.n1509 gnd 0.004435f
C3401 vdd.n1510 gnd 0.004435f
C3402 vdd.n1511 gnd 0.002383f
C3403 vdd.n1512 gnd 0.002523f
C3404 vdd.n1513 gnd 0.005633f
C3405 vdd.n1514 gnd 0.005633f
C3406 vdd.n1515 gnd 0.013317f
C3407 vdd.n1516 gnd 0.002453f
C3408 vdd.n1517 gnd 0.002383f
C3409 vdd.n1518 gnd 0.011462f
C3410 vdd.n1519 gnd 0.007751f
C3411 vdd.n1520 gnd 0.054118f
C3412 vdd.n1521 gnd 0.211067f
C3413 vdd.n1522 gnd 1.87887f
C3414 vdd.n1523 gnd 0.513636f
C3415 vdd.n1524 gnd 0.007009f
C3416 vdd.n1525 gnd 0.008708f
C3417 vdd.n1526 gnd 0.547304f
C3418 vdd.n1527 gnd 0.008708f
C3419 vdd.n1528 gnd 0.007009f
C3420 vdd.n1529 gnd 0.008708f
C3421 vdd.n1530 gnd 0.007009f
C3422 vdd.n1531 gnd 0.008708f
C3423 vdd.t89 gnd 0.444963f
C3424 vdd.t158 gnd 0.444963f
C3425 vdd.n1532 gnd 0.008708f
C3426 vdd.n1533 gnd 0.007009f
C3427 vdd.n1534 gnd 0.008708f
C3428 vdd.n1535 gnd 0.007009f
C3429 vdd.n1536 gnd 0.008708f
C3430 vdd.t91 gnd 0.444963f
C3431 vdd.n1537 gnd 0.008708f
C3432 vdd.n1538 gnd 0.007009f
C3433 vdd.n1539 gnd 0.008708f
C3434 vdd.n1540 gnd 0.007009f
C3435 vdd.n1541 gnd 0.008708f
C3436 vdd.t145 gnd 0.444963f
C3437 vdd.n1542 gnd 0.645196f
C3438 vdd.n1543 gnd 0.008708f
C3439 vdd.n1544 gnd 0.007009f
C3440 vdd.n1545 gnd 0.008708f
C3441 vdd.n1546 gnd 0.007009f
C3442 vdd.n1547 gnd 0.008708f
C3443 vdd.n1548 gnd 0.889925f
C3444 vdd.n1549 gnd 0.008708f
C3445 vdd.n1550 gnd 0.007009f
C3446 vdd.n1551 gnd 0.021222f
C3447 vdd.n1552 gnd 0.005817f
C3448 vdd.n1553 gnd 0.021222f
C3449 vdd.t3 gnd 0.444963f
C3450 vdd.n1554 gnd 0.021222f
C3451 vdd.n1555 gnd 0.005817f
C3452 vdd.n1556 gnd 0.008708f
C3453 vdd.n1557 gnd 0.007009f
C3454 vdd.n1558 gnd 0.008708f
C3455 vdd.n1589 gnd 0.021709f
C3456 vdd.n1590 gnd 1.31264f
C3457 vdd.n1591 gnd 0.008708f
C3458 vdd.n1592 gnd 0.007009f
C3459 vdd.n1593 gnd 0.008708f
C3460 vdd.n1594 gnd 0.008708f
C3461 vdd.n1595 gnd 0.008708f
C3462 vdd.n1596 gnd 0.008708f
C3463 vdd.n1597 gnd 0.008708f
C3464 vdd.n1598 gnd 0.007009f
C3465 vdd.n1599 gnd 0.008708f
C3466 vdd.n1600 gnd 0.008708f
C3467 vdd.n1601 gnd 0.008708f
C3468 vdd.n1602 gnd 0.008708f
C3469 vdd.n1603 gnd 0.008708f
C3470 vdd.n1604 gnd 0.007009f
C3471 vdd.n1605 gnd 0.008708f
C3472 vdd.n1606 gnd 0.008708f
C3473 vdd.n1607 gnd 0.008708f
C3474 vdd.n1608 gnd 0.008708f
C3475 vdd.n1609 gnd 0.008708f
C3476 vdd.n1610 gnd 0.007009f
C3477 vdd.n1611 gnd 0.008708f
C3478 vdd.n1612 gnd 0.008708f
C3479 vdd.n1613 gnd 0.008708f
C3480 vdd.n1614 gnd 0.008708f
C3481 vdd.n1615 gnd 0.008708f
C3482 vdd.t43 gnd 0.107132f
C3483 vdd.t44 gnd 0.114495f
C3484 vdd.t42 gnd 0.139914f
C3485 vdd.n1616 gnd 0.179349f
C3486 vdd.n1617 gnd 0.151387f
C3487 vdd.n1618 gnd 0.014999f
C3488 vdd.n1619 gnd 0.008708f
C3489 vdd.n1620 gnd 0.008708f
C3490 vdd.n1621 gnd 0.008708f
C3491 vdd.n1622 gnd 0.008708f
C3492 vdd.n1623 gnd 0.008708f
C3493 vdd.n1624 gnd 0.007009f
C3494 vdd.n1625 gnd 0.008708f
C3495 vdd.n1626 gnd 0.008708f
C3496 vdd.n1627 gnd 0.008708f
C3497 vdd.n1628 gnd 0.008708f
C3498 vdd.n1629 gnd 0.008708f
C3499 vdd.n1630 gnd 0.007009f
C3500 vdd.n1631 gnd 0.008708f
C3501 vdd.n1632 gnd 0.008708f
C3502 vdd.n1633 gnd 0.008708f
C3503 vdd.n1634 gnd 0.008708f
C3504 vdd.n1635 gnd 0.008708f
C3505 vdd.n1636 gnd 0.007009f
C3506 vdd.n1637 gnd 0.008708f
C3507 vdd.n1638 gnd 0.008708f
C3508 vdd.n1639 gnd 0.008708f
C3509 vdd.n1640 gnd 0.008708f
C3510 vdd.n1641 gnd 0.008708f
C3511 vdd.n1642 gnd 0.007009f
C3512 vdd.n1643 gnd 0.008708f
C3513 vdd.n1644 gnd 0.008708f
C3514 vdd.n1645 gnd 0.008708f
C3515 vdd.n1646 gnd 0.008708f
C3516 vdd.n1647 gnd 0.008708f
C3517 vdd.n1648 gnd 0.007009f
C3518 vdd.n1649 gnd 0.008708f
C3519 vdd.n1650 gnd 0.008708f
C3520 vdd.n1651 gnd 0.008708f
C3521 vdd.n1652 gnd 0.008708f
C3522 vdd.n1653 gnd 0.007009f
C3523 vdd.n1654 gnd 0.008708f
C3524 vdd.n1655 gnd 0.008708f
C3525 vdd.n1656 gnd 0.008708f
C3526 vdd.n1657 gnd 0.008708f
C3527 vdd.n1658 gnd 0.008708f
C3528 vdd.n1659 gnd 0.007009f
C3529 vdd.n1660 gnd 0.008708f
C3530 vdd.n1661 gnd 0.008708f
C3531 vdd.n1662 gnd 0.008708f
C3532 vdd.n1663 gnd 0.008708f
C3533 vdd.n1664 gnd 0.008708f
C3534 vdd.n1665 gnd 0.007009f
C3535 vdd.n1666 gnd 0.008708f
C3536 vdd.n1667 gnd 0.008708f
C3537 vdd.n1668 gnd 0.008708f
C3538 vdd.n1669 gnd 0.008708f
C3539 vdd.n1670 gnd 0.008708f
C3540 vdd.n1671 gnd 0.007009f
C3541 vdd.n1672 gnd 0.008708f
C3542 vdd.n1673 gnd 0.008708f
C3543 vdd.n1674 gnd 0.008708f
C3544 vdd.n1675 gnd 0.008708f
C3545 vdd.n1676 gnd 0.008708f
C3546 vdd.n1677 gnd 0.007009f
C3547 vdd.n1678 gnd 0.008708f
C3548 vdd.n1679 gnd 0.008708f
C3549 vdd.n1680 gnd 0.008708f
C3550 vdd.n1681 gnd 0.008708f
C3551 vdd.t4 gnd 0.107132f
C3552 vdd.t5 gnd 0.114495f
C3553 vdd.t2 gnd 0.139914f
C3554 vdd.n1682 gnd 0.179349f
C3555 vdd.n1683 gnd 0.151387f
C3556 vdd.n1684 gnd 0.011495f
C3557 vdd.n1685 gnd 0.003329f
C3558 vdd.n1686 gnd 0.021709f
C3559 vdd.n1687 gnd 0.008708f
C3560 vdd.n1688 gnd 0.00368f
C3561 vdd.n1689 gnd 0.007009f
C3562 vdd.n1690 gnd 0.007009f
C3563 vdd.n1691 gnd 0.008708f
C3564 vdd.n1692 gnd 0.008708f
C3565 vdd.n1693 gnd 0.008708f
C3566 vdd.n1694 gnd 0.007009f
C3567 vdd.n1695 gnd 0.007009f
C3568 vdd.n1696 gnd 0.007009f
C3569 vdd.n1697 gnd 0.008708f
C3570 vdd.n1698 gnd 0.008708f
C3571 vdd.n1699 gnd 0.008708f
C3572 vdd.n1700 gnd 0.007009f
C3573 vdd.n1701 gnd 0.007009f
C3574 vdd.n1702 gnd 0.007009f
C3575 vdd.n1703 gnd 0.008708f
C3576 vdd.n1704 gnd 0.008708f
C3577 vdd.n1705 gnd 0.008708f
C3578 vdd.n1706 gnd 0.007009f
C3579 vdd.n1707 gnd 0.007009f
C3580 vdd.n1708 gnd 0.007009f
C3581 vdd.n1709 gnd 0.008708f
C3582 vdd.n1710 gnd 0.008708f
C3583 vdd.n1711 gnd 0.008708f
C3584 vdd.n1712 gnd 0.007009f
C3585 vdd.n1713 gnd 0.007009f
C3586 vdd.n1714 gnd 0.007009f
C3587 vdd.n1715 gnd 0.008708f
C3588 vdd.n1716 gnd 0.008708f
C3589 vdd.n1717 gnd 0.008708f
C3590 vdd.n1718 gnd 0.006939f
C3591 vdd.n1719 gnd 0.008708f
C3592 vdd.t33 gnd 0.107132f
C3593 vdd.t34 gnd 0.114495f
C3594 vdd.t32 gnd 0.139914f
C3595 vdd.n1720 gnd 0.179349f
C3596 vdd.n1721 gnd 0.151387f
C3597 vdd.n1722 gnd 0.014999f
C3598 vdd.n1723 gnd 0.004766f
C3599 vdd.n1724 gnd 0.008708f
C3600 vdd.n1725 gnd 0.008708f
C3601 vdd.n1726 gnd 0.008708f
C3602 vdd.n1727 gnd 0.007009f
C3603 vdd.n1728 gnd 0.007009f
C3604 vdd.n1729 gnd 0.007009f
C3605 vdd.n1730 gnd 0.008708f
C3606 vdd.n1731 gnd 0.008708f
C3607 vdd.n1732 gnd 0.008708f
C3608 vdd.n1733 gnd 0.007009f
C3609 vdd.n1734 gnd 0.007009f
C3610 vdd.n1735 gnd 0.007009f
C3611 vdd.n1736 gnd 0.008708f
C3612 vdd.n1737 gnd 0.008708f
C3613 vdd.n1738 gnd 0.008708f
C3614 vdd.n1739 gnd 0.007009f
C3615 vdd.n1740 gnd 0.007009f
C3616 vdd.n1741 gnd 0.007009f
C3617 vdd.n1742 gnd 0.008708f
C3618 vdd.n1743 gnd 0.008708f
C3619 vdd.n1744 gnd 0.008708f
C3620 vdd.n1745 gnd 0.007009f
C3621 vdd.n1746 gnd 0.007009f
C3622 vdd.n1747 gnd 0.007009f
C3623 vdd.n1748 gnd 0.008708f
C3624 vdd.n1749 gnd 0.008708f
C3625 vdd.n1750 gnd 0.008708f
C3626 vdd.n1751 gnd 0.007009f
C3627 vdd.n1752 gnd 0.007009f
C3628 vdd.n1753 gnd 0.005852f
C3629 vdd.n1754 gnd 0.008708f
C3630 vdd.n1755 gnd 0.008708f
C3631 vdd.n1756 gnd 0.008708f
C3632 vdd.n1757 gnd 0.005852f
C3633 vdd.n1758 gnd 0.007009f
C3634 vdd.n1759 gnd 0.007009f
C3635 vdd.n1760 gnd 0.008708f
C3636 vdd.n1761 gnd 0.008708f
C3637 vdd.n1762 gnd 0.008708f
C3638 vdd.n1763 gnd 0.007009f
C3639 vdd.n1764 gnd 0.007009f
C3640 vdd.n1765 gnd 0.007009f
C3641 vdd.n1766 gnd 0.008708f
C3642 vdd.n1767 gnd 0.008708f
C3643 vdd.n1768 gnd 0.008708f
C3644 vdd.n1769 gnd 0.007009f
C3645 vdd.n1770 gnd 0.007009f
C3646 vdd.n1771 gnd 0.007009f
C3647 vdd.n1772 gnd 0.008708f
C3648 vdd.n1773 gnd 0.008708f
C3649 vdd.n1774 gnd 0.008708f
C3650 vdd.n1775 gnd 0.007009f
C3651 vdd.n1776 gnd 0.007009f
C3652 vdd.n1777 gnd 0.007009f
C3653 vdd.n1778 gnd 0.008708f
C3654 vdd.n1779 gnd 0.008708f
C3655 vdd.n1780 gnd 0.008708f
C3656 vdd.n1781 gnd 0.007009f
C3657 vdd.n1782 gnd 0.008708f
C3658 vdd.n1783 gnd 2.12692f
C3659 vdd.n1785 gnd 0.021709f
C3660 vdd.n1786 gnd 0.005817f
C3661 vdd.n1787 gnd 0.021709f
C3662 vdd.n1788 gnd 0.021222f
C3663 vdd.n1789 gnd 0.008708f
C3664 vdd.n1790 gnd 0.007009f
C3665 vdd.n1791 gnd 0.008708f
C3666 vdd.n1792 gnd 0.467211f
C3667 vdd.n1793 gnd 0.008708f
C3668 vdd.n1794 gnd 0.007009f
C3669 vdd.n1795 gnd 0.008708f
C3670 vdd.n1796 gnd 0.008708f
C3671 vdd.n1797 gnd 0.008708f
C3672 vdd.n1798 gnd 0.007009f
C3673 vdd.n1799 gnd 0.008708f
C3674 vdd.n1800 gnd 0.796483f
C3675 vdd.n1801 gnd 0.889925f
C3676 vdd.n1802 gnd 0.008708f
C3677 vdd.n1803 gnd 0.007009f
C3678 vdd.n1804 gnd 0.008708f
C3679 vdd.n1805 gnd 0.008708f
C3680 vdd.n1806 gnd 0.008708f
C3681 vdd.n1807 gnd 0.007009f
C3682 vdd.n1808 gnd 0.008708f
C3683 vdd.n1809 gnd 0.538405f
C3684 vdd.n1810 gnd 0.008708f
C3685 vdd.n1811 gnd 0.007009f
C3686 vdd.n1812 gnd 0.008708f
C3687 vdd.n1813 gnd 0.008708f
C3688 vdd.n1814 gnd 0.008708f
C3689 vdd.n1815 gnd 0.007009f
C3690 vdd.n1816 gnd 0.008708f
C3691 vdd.n1817 gnd 0.493909f
C3692 vdd.n1818 gnd 0.689692f
C3693 vdd.n1819 gnd 0.008708f
C3694 vdd.n1820 gnd 0.007009f
C3695 vdd.n1821 gnd 0.008708f
C3696 vdd.n1822 gnd 0.008708f
C3697 vdd.n1823 gnd 0.006693f
C3698 vdd.n1824 gnd 0.008708f
C3699 vdd.n1825 gnd 0.007009f
C3700 vdd.n1826 gnd 0.008708f
C3701 vdd.n1827 gnd 0.738638f
C3702 vdd.n1828 gnd 0.008708f
C3703 vdd.n1829 gnd 0.007009f
C3704 vdd.n1830 gnd 0.008708f
C3705 vdd.n1831 gnd 0.008708f
C3706 vdd.n1832 gnd 0.008708f
C3707 vdd.n1833 gnd 0.007009f
C3708 vdd.n1834 gnd 0.008708f
C3709 vdd.t143 gnd 0.444963f
C3710 vdd.n1835 gnd 0.636297f
C3711 vdd.n1836 gnd 0.008708f
C3712 vdd.n1837 gnd 0.007009f
C3713 vdd.n1838 gnd 0.006693f
C3714 vdd.n1839 gnd 0.008708f
C3715 vdd.n1840 gnd 0.008708f
C3716 vdd.n1841 gnd 0.007009f
C3717 vdd.n1842 gnd 0.008708f
C3718 vdd.n1843 gnd 0.485009f
C3719 vdd.n1844 gnd 0.008708f
C3720 vdd.n1845 gnd 0.007009f
C3721 vdd.n1846 gnd 0.008708f
C3722 vdd.n1847 gnd 0.008708f
C3723 vdd.n1848 gnd 0.008708f
C3724 vdd.n1849 gnd 0.007009f
C3725 vdd.n1850 gnd 0.008708f
C3726 vdd.n1851 gnd 0.627397f
C3727 vdd.n1852 gnd 0.556203f
C3728 vdd.n1853 gnd 0.008708f
C3729 vdd.n1854 gnd 0.007009f
C3730 vdd.n1855 gnd 0.008708f
C3731 vdd.n1856 gnd 0.008708f
C3732 vdd.n1857 gnd 0.008708f
C3733 vdd.n1858 gnd 0.007009f
C3734 vdd.n1859 gnd 0.008708f
C3735 vdd.n1860 gnd 0.707491f
C3736 vdd.n1861 gnd 0.008708f
C3737 vdd.n1862 gnd 0.007009f
C3738 vdd.n1863 gnd 0.008708f
C3739 vdd.n1864 gnd 0.008708f
C3740 vdd.n1865 gnd 0.021222f
C3741 vdd.n1866 gnd 0.008708f
C3742 vdd.n1867 gnd 0.008708f
C3743 vdd.n1868 gnd 0.007009f
C3744 vdd.n1869 gnd 0.008708f
C3745 vdd.n1870 gnd 0.556203f
C3746 vdd.n1871 gnd 0.889925f
C3747 vdd.n1872 gnd 0.008708f
C3748 vdd.n1873 gnd 0.007009f
C3749 vdd.n1874 gnd 0.008708f
C3750 vdd.n1875 gnd 0.008708f
C3751 vdd.n1876 gnd 0.021222f
C3752 vdd.n1877 gnd 0.005817f
C3753 vdd.n1878 gnd 0.021222f
C3754 vdd.n1879 gnd 1.22365f
C3755 vdd.n1880 gnd 0.021222f
C3756 vdd.n1881 gnd 0.021709f
C3757 vdd.n1882 gnd 0.003329f
C3758 vdd.t25 gnd 0.107132f
C3759 vdd.t24 gnd 0.114495f
C3760 vdd.t22 gnd 0.139914f
C3761 vdd.n1883 gnd 0.179349f
C3762 vdd.n1884 gnd 0.150686f
C3763 vdd.n1885 gnd 0.010794f
C3764 vdd.n1886 gnd 0.00368f
C3765 vdd.n1887 gnd 0.007489f
C3766 vdd.n1888 gnd 0.658553f
C3767 vdd.n1890 gnd 0.007009f
C3768 vdd.n1891 gnd 0.007009f
C3769 vdd.n1892 gnd 0.008708f
C3770 vdd.n1894 gnd 0.008708f
C3771 vdd.n1895 gnd 0.008708f
C3772 vdd.n1896 gnd 0.007009f
C3773 vdd.n1897 gnd 0.007009f
C3774 vdd.n1898 gnd 0.007009f
C3775 vdd.n1899 gnd 0.008708f
C3776 vdd.n1901 gnd 0.008708f
C3777 vdd.n1902 gnd 0.008708f
C3778 vdd.n1903 gnd 0.007009f
C3779 vdd.n1904 gnd 0.007009f
C3780 vdd.n1905 gnd 0.007009f
C3781 vdd.n1906 gnd 0.008708f
C3782 vdd.n1908 gnd 0.008708f
C3783 vdd.n1909 gnd 0.008708f
C3784 vdd.n1910 gnd 0.007009f
C3785 vdd.n1911 gnd 0.007009f
C3786 vdd.n1912 gnd 0.007009f
C3787 vdd.n1913 gnd 0.008708f
C3788 vdd.n1915 gnd 0.008708f
C3789 vdd.n1916 gnd 0.008708f
C3790 vdd.n1917 gnd 0.007009f
C3791 vdd.n1918 gnd 0.008708f
C3792 vdd.n1919 gnd 0.008708f
C3793 vdd.n1920 gnd 0.008708f
C3794 vdd.n1921 gnd 0.014298f
C3795 vdd.n1922 gnd 0.004766f
C3796 vdd.n1923 gnd 0.007009f
C3797 vdd.n1924 gnd 0.008708f
C3798 vdd.n1926 gnd 0.008708f
C3799 vdd.n1927 gnd 0.008708f
C3800 vdd.n1928 gnd 0.007009f
C3801 vdd.n1929 gnd 0.007009f
C3802 vdd.n1930 gnd 0.007009f
C3803 vdd.n1931 gnd 0.008708f
C3804 vdd.n1933 gnd 0.008708f
C3805 vdd.n1934 gnd 0.008708f
C3806 vdd.n1935 gnd 0.007009f
C3807 vdd.n1936 gnd 0.007009f
C3808 vdd.n1937 gnd 0.007009f
C3809 vdd.n1938 gnd 0.008708f
C3810 vdd.n1940 gnd 0.008708f
C3811 vdd.n1941 gnd 0.008708f
C3812 vdd.n1942 gnd 0.007009f
C3813 vdd.n1943 gnd 0.007009f
C3814 vdd.n1944 gnd 0.007009f
C3815 vdd.n1945 gnd 0.008708f
C3816 vdd.n1947 gnd 0.008708f
C3817 vdd.n1948 gnd 0.008708f
C3818 vdd.n1949 gnd 0.007009f
C3819 vdd.n1950 gnd 0.007009f
C3820 vdd.n1951 gnd 0.007009f
C3821 vdd.n1952 gnd 0.008708f
C3822 vdd.n1954 gnd 0.008708f
C3823 vdd.n1955 gnd 0.008708f
C3824 vdd.n1956 gnd 0.007009f
C3825 vdd.n1957 gnd 0.008708f
C3826 vdd.n1958 gnd 0.008708f
C3827 vdd.n1959 gnd 0.008708f
C3828 vdd.n1960 gnd 0.014298f
C3829 vdd.n1961 gnd 0.005852f
C3830 vdd.n1962 gnd 0.007009f
C3831 vdd.n1963 gnd 0.008708f
C3832 vdd.n1965 gnd 0.008708f
C3833 vdd.n1966 gnd 0.008708f
C3834 vdd.n1967 gnd 0.007009f
C3835 vdd.n1968 gnd 0.007009f
C3836 vdd.n1969 gnd 0.007009f
C3837 vdd.n1970 gnd 0.008708f
C3838 vdd.n1972 gnd 0.008708f
C3839 vdd.n1973 gnd 0.008708f
C3840 vdd.n1974 gnd 0.007009f
C3841 vdd.n1975 gnd 0.007009f
C3842 vdd.n1976 gnd 0.007009f
C3843 vdd.n1977 gnd 0.008708f
C3844 vdd.n1979 gnd 0.008708f
C3845 vdd.n1980 gnd 0.008708f
C3846 vdd.n1981 gnd 0.007009f
C3847 vdd.n1982 gnd 0.007009f
C3848 vdd.n1983 gnd 0.007009f
C3849 vdd.n1984 gnd 0.008708f
C3850 vdd.n1986 gnd 0.008708f
C3851 vdd.n1987 gnd 0.007009f
C3852 vdd.n1988 gnd 0.007009f
C3853 vdd.n1989 gnd 0.008708f
C3854 vdd.n1991 gnd 0.008708f
C3855 vdd.n1992 gnd 0.008708f
C3856 vdd.n1993 gnd 0.007009f
C3857 vdd.n1994 gnd 0.007489f
C3858 vdd.n1995 gnd 0.658553f
C3859 vdd.n1996 gnd 0.023733f
C3860 vdd.n1997 gnd 0.005922f
C3861 vdd.n1998 gnd 0.005922f
C3862 vdd.n1999 gnd 0.005922f
C3863 vdd.n2000 gnd 0.005922f
C3864 vdd.n2001 gnd 0.005922f
C3865 vdd.n2002 gnd 0.005922f
C3866 vdd.n2003 gnd 0.005922f
C3867 vdd.n2004 gnd 0.005922f
C3868 vdd.n2005 gnd 0.005922f
C3869 vdd.n2006 gnd 0.005922f
C3870 vdd.n2007 gnd 0.005922f
C3871 vdd.n2008 gnd 0.005922f
C3872 vdd.n2009 gnd 0.005922f
C3873 vdd.n2010 gnd 0.005922f
C3874 vdd.n2011 gnd 0.005922f
C3875 vdd.n2012 gnd 0.005922f
C3876 vdd.n2013 gnd 0.005922f
C3877 vdd.n2014 gnd 0.005922f
C3878 vdd.n2015 gnd 0.005922f
C3879 vdd.n2016 gnd 0.005922f
C3880 vdd.n2017 gnd 0.005922f
C3881 vdd.n2018 gnd 0.005922f
C3882 vdd.n2019 gnd 0.005922f
C3883 vdd.n2020 gnd 0.005922f
C3884 vdd.n2021 gnd 0.005922f
C3885 vdd.n2022 gnd 0.005922f
C3886 vdd.n2023 gnd 0.005922f
C3887 vdd.n2024 gnd 0.005922f
C3888 vdd.n2025 gnd 0.005922f
C3889 vdd.n2026 gnd 0.005922f
C3890 vdd.n2027 gnd 0.005922f
C3891 vdd.n2028 gnd 0.01385f
C3892 vdd.n2029 gnd 0.01385f
C3893 vdd.n2031 gnd 7.59106f
C3894 vdd.n2033 gnd 0.01385f
C3895 vdd.n2034 gnd 0.01385f
C3896 vdd.n2035 gnd 0.012971f
C3897 vdd.n2036 gnd 0.005922f
C3898 vdd.n2037 gnd 0.005922f
C3899 vdd.n2038 gnd 0.605149f
C3900 vdd.n2039 gnd 0.005922f
C3901 vdd.n2040 gnd 0.005922f
C3902 vdd.n2041 gnd 0.005922f
C3903 vdd.n2042 gnd 0.005922f
C3904 vdd.n2043 gnd 0.005922f
C3905 vdd.n2044 gnd 0.511707f
C3906 vdd.n2045 gnd 0.005922f
C3907 vdd.n2046 gnd 0.005922f
C3908 vdd.n2047 gnd 0.005922f
C3909 vdd.n2048 gnd 0.005922f
C3910 vdd.n2049 gnd 0.005922f
C3911 vdd.n2050 gnd 0.605149f
C3912 vdd.n2051 gnd 0.005922f
C3913 vdd.n2052 gnd 0.005922f
C3914 vdd.n2053 gnd 0.005922f
C3915 vdd.n2054 gnd 0.005922f
C3916 vdd.n2055 gnd 0.005922f
C3917 vdd.n2056 gnd 0.5918f
C3918 vdd.n2057 gnd 0.005922f
C3919 vdd.n2058 gnd 0.005922f
C3920 vdd.n2059 gnd 0.005922f
C3921 vdd.n2060 gnd 0.005922f
C3922 vdd.n2061 gnd 0.005922f
C3923 vdd.n2062 gnd 0.605149f
C3924 vdd.n2063 gnd 0.005922f
C3925 vdd.n2064 gnd 0.005922f
C3926 vdd.n2065 gnd 0.005922f
C3927 vdd.n2066 gnd 0.005922f
C3928 vdd.n2067 gnd 0.005922f
C3929 vdd.n2068 gnd 0.485009f
C3930 vdd.n2069 gnd 0.005922f
C3931 vdd.n2070 gnd 0.005922f
C3932 vdd.n2071 gnd 0.005051f
C3933 vdd.n2072 gnd 0.017154f
C3934 vdd.n2073 gnd 0.003832f
C3935 vdd.n2074 gnd 0.005922f
C3936 vdd.n2075 gnd 0.35152f
C3937 vdd.n2076 gnd 0.005922f
C3938 vdd.n2077 gnd 0.005922f
C3939 vdd.n2078 gnd 0.005922f
C3940 vdd.n2079 gnd 0.005922f
C3941 vdd.n2080 gnd 0.005922f
C3942 vdd.n2081 gnd 0.387117f
C3943 vdd.n2082 gnd 0.005922f
C3944 vdd.n2083 gnd 0.005922f
C3945 vdd.n2084 gnd 0.005922f
C3946 vdd.n2085 gnd 0.005922f
C3947 vdd.n2086 gnd 0.005922f
C3948 vdd.n2087 gnd 0.520606f
C3949 vdd.n2088 gnd 0.005922f
C3950 vdd.n2089 gnd 0.005922f
C3951 vdd.n2090 gnd 0.005922f
C3952 vdd.n2091 gnd 0.005922f
C3953 vdd.n2092 gnd 0.005922f
C3954 vdd.n2093 gnd 0.498358f
C3955 vdd.n2094 gnd 0.005922f
C3956 vdd.n2095 gnd 0.005922f
C3957 vdd.n2096 gnd 0.005922f
C3958 vdd.n2097 gnd 0.005922f
C3959 vdd.n2098 gnd 0.005922f
C3960 vdd.n2099 gnd 0.364869f
C3961 vdd.n2100 gnd 0.005922f
C3962 vdd.n2101 gnd 0.005922f
C3963 vdd.n2102 gnd 0.005922f
C3964 vdd.n2103 gnd 0.005922f
C3965 vdd.n2104 gnd 0.005922f
C3966 vdd.n2105 gnd 0.191334f
C3967 vdd.n2106 gnd 0.005922f
C3968 vdd.n2107 gnd 0.005922f
C3969 vdd.n2108 gnd 0.005922f
C3970 vdd.n2109 gnd 0.005922f
C3971 vdd.n2110 gnd 0.005922f
C3972 vdd.n2111 gnd 0.315923f
C3973 vdd.n2112 gnd 0.005922f
C3974 vdd.n2113 gnd 0.005922f
C3975 vdd.n2114 gnd 0.005922f
C3976 vdd.n2115 gnd 0.005922f
C3977 vdd.n2116 gnd 0.005922f
C3978 vdd.n2117 gnd 0.605149f
C3979 vdd.n2118 gnd 0.005922f
C3980 vdd.n2119 gnd 0.005922f
C3981 vdd.n2120 gnd 0.005922f
C3982 vdd.n2121 gnd 0.005922f
C3983 vdd.n2122 gnd 0.005922f
C3984 vdd.n2123 gnd 0.005922f
C3985 vdd.n2124 gnd 0.005922f
C3986 vdd.n2125 gnd 0.453862f
C3987 vdd.n2126 gnd 0.005922f
C3988 vdd.n2127 gnd 0.005922f
C3989 vdd.n2128 gnd 0.005922f
C3990 vdd.n2129 gnd 0.005922f
C3991 vdd.n2130 gnd 0.005922f
C3992 vdd.n2131 gnd 0.005922f
C3993 vdd.n2132 gnd 0.378218f
C3994 vdd.n2133 gnd 0.005922f
C3995 vdd.n2134 gnd 0.005922f
C3996 vdd.n2135 gnd 0.005922f
C3997 vdd.n2136 gnd 0.013707f
C3998 vdd.n2137 gnd 0.013114f
C3999 vdd.n2138 gnd 0.005922f
C4000 vdd.n2139 gnd 0.005922f
C4001 vdd.n2140 gnd 0.004572f
C4002 vdd.n2141 gnd 0.005922f
C4003 vdd.n2142 gnd 0.005922f
C4004 vdd.n2143 gnd 0.004311f
C4005 vdd.n2144 gnd 0.005922f
C4006 vdd.n2145 gnd 0.005922f
C4007 vdd.n2146 gnd 0.005922f
C4008 vdd.n2147 gnd 0.005922f
C4009 vdd.n2148 gnd 0.005922f
C4010 vdd.n2149 gnd 0.005922f
C4011 vdd.n2150 gnd 0.005922f
C4012 vdd.n2151 gnd 0.005922f
C4013 vdd.n2152 gnd 0.005922f
C4014 vdd.n2153 gnd 0.005922f
C4015 vdd.n2154 gnd 0.005922f
C4016 vdd.n2155 gnd 0.005922f
C4017 vdd.n2156 gnd 0.005922f
C4018 vdd.n2157 gnd 0.005922f
C4019 vdd.n2158 gnd 0.005922f
C4020 vdd.n2159 gnd 0.005922f
C4021 vdd.n2160 gnd 0.005922f
C4022 vdd.n2161 gnd 0.005922f
C4023 vdd.n2162 gnd 0.005922f
C4024 vdd.n2163 gnd 0.005922f
C4025 vdd.n2164 gnd 0.005922f
C4026 vdd.n2165 gnd 0.005922f
C4027 vdd.n2166 gnd 0.005922f
C4028 vdd.n2167 gnd 0.005922f
C4029 vdd.n2168 gnd 0.005922f
C4030 vdd.n2169 gnd 0.005922f
C4031 vdd.n2170 gnd 0.005922f
C4032 vdd.n2171 gnd 0.005922f
C4033 vdd.n2172 gnd 0.005922f
C4034 vdd.n2173 gnd 0.005922f
C4035 vdd.n2174 gnd 0.005922f
C4036 vdd.n2175 gnd 0.005922f
C4037 vdd.n2176 gnd 0.005922f
C4038 vdd.n2177 gnd 0.005922f
C4039 vdd.n2178 gnd 0.005922f
C4040 vdd.n2179 gnd 0.005922f
C4041 vdd.n2180 gnd 0.005922f
C4042 vdd.n2181 gnd 0.005922f
C4043 vdd.n2182 gnd 0.005922f
C4044 vdd.n2183 gnd 0.005922f
C4045 vdd.n2184 gnd 0.005922f
C4046 vdd.n2185 gnd 0.005922f
C4047 vdd.n2186 gnd 0.005922f
C4048 vdd.n2187 gnd 0.005922f
C4049 vdd.n2188 gnd 0.005922f
C4050 vdd.n2189 gnd 0.005922f
C4051 vdd.n2190 gnd 0.005922f
C4052 vdd.n2191 gnd 0.005922f
C4053 vdd.n2192 gnd 0.005922f
C4054 vdd.n2193 gnd 0.005922f
C4055 vdd.n2194 gnd 0.005922f
C4056 vdd.n2195 gnd 0.005922f
C4057 vdd.n2196 gnd 0.005922f
C4058 vdd.n2197 gnd 0.005922f
C4059 vdd.n2198 gnd 0.005922f
C4060 vdd.n2199 gnd 0.005922f
C4061 vdd.n2200 gnd 0.005922f
C4062 vdd.n2201 gnd 0.005922f
C4063 vdd.n2202 gnd 0.005922f
C4064 vdd.n2203 gnd 0.005922f
C4065 vdd.n2204 gnd 0.01385f
C4066 vdd.n2205 gnd 0.012971f
C4067 vdd.n2206 gnd 0.012971f
C4068 vdd.n2207 gnd 0.720839f
C4069 vdd.n2208 gnd 0.012971f
C4070 vdd.n2209 gnd 0.01385f
C4071 vdd.n2210 gnd 0.013114f
C4072 vdd.n2211 gnd 0.005922f
C4073 vdd.n2212 gnd 0.005922f
C4074 vdd.n2213 gnd 0.005922f
C4075 vdd.n2214 gnd 0.004572f
C4076 vdd.n2215 gnd 0.008463f
C4077 vdd.n2216 gnd 0.004311f
C4078 vdd.n2217 gnd 0.005922f
C4079 vdd.n2218 gnd 0.005922f
C4080 vdd.n2219 gnd 0.005922f
C4081 vdd.n2220 gnd 0.005922f
C4082 vdd.n2221 gnd 0.005922f
C4083 vdd.n2222 gnd 0.005922f
C4084 vdd.n2223 gnd 0.005922f
C4085 vdd.n2224 gnd 0.005922f
C4086 vdd.n2225 gnd 0.005922f
C4087 vdd.n2226 gnd 0.005922f
C4088 vdd.n2227 gnd 0.005922f
C4089 vdd.n2228 gnd 0.005922f
C4090 vdd.n2229 gnd 0.005922f
C4091 vdd.n2230 gnd 0.005922f
C4092 vdd.n2231 gnd 0.005922f
C4093 vdd.n2232 gnd 0.005922f
C4094 vdd.n2233 gnd 0.005922f
C4095 vdd.n2234 gnd 0.005922f
C4096 vdd.n2235 gnd 0.005922f
C4097 vdd.n2236 gnd 0.005922f
C4098 vdd.n2237 gnd 0.005922f
C4099 vdd.n2238 gnd 0.005922f
C4100 vdd.n2239 gnd 0.005922f
C4101 vdd.n2240 gnd 0.005922f
C4102 vdd.n2241 gnd 0.005922f
C4103 vdd.n2242 gnd 0.005922f
C4104 vdd.n2243 gnd 0.005922f
C4105 vdd.n2244 gnd 0.005922f
C4106 vdd.n2245 gnd 0.005922f
C4107 vdd.n2246 gnd 0.005922f
C4108 vdd.n2247 gnd 0.005922f
C4109 vdd.n2248 gnd 0.005922f
C4110 vdd.n2249 gnd 0.005922f
C4111 vdd.n2250 gnd 0.005922f
C4112 vdd.n2251 gnd 0.005922f
C4113 vdd.n2252 gnd 0.005922f
C4114 vdd.n2253 gnd 0.005922f
C4115 vdd.n2254 gnd 0.005922f
C4116 vdd.n2255 gnd 0.005922f
C4117 vdd.n2256 gnd 0.005922f
C4118 vdd.n2257 gnd 0.005922f
C4119 vdd.n2258 gnd 0.005922f
C4120 vdd.n2259 gnd 0.005922f
C4121 vdd.n2260 gnd 0.005922f
C4122 vdd.n2261 gnd 0.005922f
C4123 vdd.n2262 gnd 0.005922f
C4124 vdd.n2263 gnd 0.005922f
C4125 vdd.n2264 gnd 0.005922f
C4126 vdd.n2265 gnd 0.005922f
C4127 vdd.n2266 gnd 0.005922f
C4128 vdd.n2267 gnd 0.005922f
C4129 vdd.n2268 gnd 0.005922f
C4130 vdd.n2269 gnd 0.005922f
C4131 vdd.n2270 gnd 0.005922f
C4132 vdd.n2271 gnd 0.005922f
C4133 vdd.n2272 gnd 0.005922f
C4134 vdd.n2273 gnd 0.005922f
C4135 vdd.n2274 gnd 0.005922f
C4136 vdd.n2275 gnd 0.005922f
C4137 vdd.n2276 gnd 0.005922f
C4138 vdd.n2277 gnd 0.01385f
C4139 vdd.n2278 gnd 0.01385f
C4140 vdd.n2279 gnd 0.738638f
C4141 vdd.t118 gnd 2.62528f
C4142 vdd.t107 gnd 2.62528f
C4143 vdd.n2312 gnd 0.01385f
C4144 vdd.t120 gnd 0.551754f
C4145 vdd.n2313 gnd 0.005922f
C4146 vdd.n2314 gnd 0.005922f
C4147 vdd.t54 gnd 0.239287f
C4148 vdd.t55 gnd 0.24494f
C4149 vdd.t52 gnd 0.156216f
C4150 vdd.n2315 gnd 0.084426f
C4151 vdd.n2316 gnd 0.047889f
C4152 vdd.n2317 gnd 0.005922f
C4153 vdd.t61 gnd 0.239287f
C4154 vdd.t62 gnd 0.24494f
C4155 vdd.t60 gnd 0.156216f
C4156 vdd.n2318 gnd 0.084426f
C4157 vdd.n2319 gnd 0.047889f
C4158 vdd.n2320 gnd 0.008463f
C4159 vdd.n2321 gnd 0.005922f
C4160 vdd.n2322 gnd 0.005922f
C4161 vdd.n2323 gnd 0.005922f
C4162 vdd.n2324 gnd 0.005922f
C4163 vdd.n2325 gnd 0.005922f
C4164 vdd.n2326 gnd 0.005922f
C4165 vdd.n2327 gnd 0.005922f
C4166 vdd.n2328 gnd 0.005922f
C4167 vdd.n2329 gnd 0.005922f
C4168 vdd.n2330 gnd 0.005922f
C4169 vdd.n2331 gnd 0.005922f
C4170 vdd.n2332 gnd 0.005922f
C4171 vdd.n2333 gnd 0.005922f
C4172 vdd.n2334 gnd 0.005922f
C4173 vdd.n2335 gnd 0.005922f
C4174 vdd.n2336 gnd 0.005922f
C4175 vdd.n2337 gnd 0.005922f
C4176 vdd.n2338 gnd 0.005922f
C4177 vdd.n2339 gnd 0.005922f
C4178 vdd.n2340 gnd 0.005922f
C4179 vdd.n2341 gnd 0.005922f
C4180 vdd.n2342 gnd 0.005922f
C4181 vdd.n2343 gnd 0.005922f
C4182 vdd.n2344 gnd 0.005922f
C4183 vdd.n2345 gnd 0.005922f
C4184 vdd.n2346 gnd 0.005922f
C4185 vdd.n2347 gnd 0.005922f
C4186 vdd.n2348 gnd 0.005922f
C4187 vdd.n2349 gnd 0.005922f
C4188 vdd.n2350 gnd 0.005922f
C4189 vdd.n2351 gnd 0.005922f
C4190 vdd.n2352 gnd 0.005922f
C4191 vdd.n2353 gnd 0.005922f
C4192 vdd.n2354 gnd 0.005922f
C4193 vdd.n2355 gnd 0.005922f
C4194 vdd.n2356 gnd 0.005922f
C4195 vdd.n2357 gnd 0.005922f
C4196 vdd.n2358 gnd 0.005922f
C4197 vdd.n2359 gnd 0.005922f
C4198 vdd.n2360 gnd 0.005922f
C4199 vdd.n2361 gnd 0.005922f
C4200 vdd.n2362 gnd 0.005922f
C4201 vdd.n2363 gnd 0.005922f
C4202 vdd.n2364 gnd 0.005922f
C4203 vdd.n2365 gnd 0.005922f
C4204 vdd.n2366 gnd 0.005922f
C4205 vdd.n2367 gnd 0.005922f
C4206 vdd.n2368 gnd 0.005922f
C4207 vdd.n2369 gnd 0.005922f
C4208 vdd.n2370 gnd 0.005922f
C4209 vdd.n2371 gnd 0.005922f
C4210 vdd.n2372 gnd 0.005922f
C4211 vdd.n2373 gnd 0.005922f
C4212 vdd.n2374 gnd 0.005922f
C4213 vdd.n2375 gnd 0.005922f
C4214 vdd.n2376 gnd 0.005922f
C4215 vdd.n2377 gnd 0.005922f
C4216 vdd.n2378 gnd 0.005922f
C4217 vdd.n2379 gnd 0.004311f
C4218 vdd.n2380 gnd 0.005922f
C4219 vdd.n2381 gnd 0.005922f
C4220 vdd.n2382 gnd 0.004572f
C4221 vdd.n2383 gnd 0.005922f
C4222 vdd.n2384 gnd 0.005922f
C4223 vdd.n2385 gnd 0.01385f
C4224 vdd.n2386 gnd 0.012971f
C4225 vdd.n2387 gnd 0.012971f
C4226 vdd.n2388 gnd 0.005922f
C4227 vdd.n2389 gnd 0.005922f
C4228 vdd.n2390 gnd 0.005922f
C4229 vdd.n2391 gnd 0.005922f
C4230 vdd.n2392 gnd 0.005922f
C4231 vdd.n2393 gnd 0.005922f
C4232 vdd.n2394 gnd 0.005922f
C4233 vdd.n2395 gnd 0.005922f
C4234 vdd.n2396 gnd 0.005922f
C4235 vdd.n2397 gnd 0.005922f
C4236 vdd.n2398 gnd 0.005922f
C4237 vdd.n2399 gnd 0.005922f
C4238 vdd.n2400 gnd 0.005922f
C4239 vdd.n2401 gnd 0.005922f
C4240 vdd.n2402 gnd 0.005922f
C4241 vdd.n2403 gnd 0.005922f
C4242 vdd.n2404 gnd 0.005922f
C4243 vdd.n2405 gnd 0.005922f
C4244 vdd.n2406 gnd 0.005922f
C4245 vdd.n2407 gnd 0.005922f
C4246 vdd.n2408 gnd 0.005922f
C4247 vdd.n2409 gnd 0.005922f
C4248 vdd.n2410 gnd 0.005922f
C4249 vdd.n2411 gnd 0.005922f
C4250 vdd.n2412 gnd 0.005922f
C4251 vdd.n2413 gnd 0.005922f
C4252 vdd.n2414 gnd 0.005922f
C4253 vdd.n2415 gnd 0.005922f
C4254 vdd.n2416 gnd 0.005922f
C4255 vdd.n2417 gnd 0.005922f
C4256 vdd.n2418 gnd 0.005922f
C4257 vdd.n2419 gnd 0.005922f
C4258 vdd.n2420 gnd 0.005922f
C4259 vdd.n2421 gnd 0.005922f
C4260 vdd.n2422 gnd 0.005922f
C4261 vdd.n2423 gnd 0.005922f
C4262 vdd.n2424 gnd 0.005922f
C4263 vdd.n2425 gnd 0.005922f
C4264 vdd.n2426 gnd 0.005922f
C4265 vdd.n2427 gnd 0.005922f
C4266 vdd.n2428 gnd 0.005922f
C4267 vdd.n2429 gnd 0.005922f
C4268 vdd.n2430 gnd 0.005922f
C4269 vdd.n2431 gnd 0.005922f
C4270 vdd.n2432 gnd 0.005922f
C4271 vdd.n2433 gnd 0.005922f
C4272 vdd.n2434 gnd 0.005922f
C4273 vdd.n2435 gnd 0.005922f
C4274 vdd.n2436 gnd 0.005922f
C4275 vdd.n2437 gnd 0.005922f
C4276 vdd.n2438 gnd 0.005922f
C4277 vdd.n2439 gnd 0.005922f
C4278 vdd.n2440 gnd 0.005922f
C4279 vdd.n2441 gnd 0.005922f
C4280 vdd.n2442 gnd 0.005922f
C4281 vdd.n2443 gnd 0.005922f
C4282 vdd.n2444 gnd 0.005922f
C4283 vdd.n2445 gnd 0.005922f
C4284 vdd.n2446 gnd 0.005922f
C4285 vdd.n2447 gnd 0.005922f
C4286 vdd.n2448 gnd 0.005922f
C4287 vdd.n2449 gnd 0.005922f
C4288 vdd.n2450 gnd 0.005922f
C4289 vdd.n2451 gnd 0.005922f
C4290 vdd.n2452 gnd 0.005922f
C4291 vdd.n2453 gnd 0.005922f
C4292 vdd.n2454 gnd 0.005922f
C4293 vdd.n2455 gnd 0.005922f
C4294 vdd.n2456 gnd 0.005922f
C4295 vdd.n2457 gnd 0.005922f
C4296 vdd.n2458 gnd 0.005922f
C4297 vdd.n2459 gnd 0.005922f
C4298 vdd.n2460 gnd 0.005922f
C4299 vdd.n2461 gnd 0.191334f
C4300 vdd.n2462 gnd 0.005922f
C4301 vdd.n2463 gnd 0.005922f
C4302 vdd.n2464 gnd 0.005922f
C4303 vdd.n2465 gnd 0.005922f
C4304 vdd.n2466 gnd 0.005922f
C4305 vdd.n2467 gnd 0.005922f
C4306 vdd.n2468 gnd 0.005922f
C4307 vdd.n2469 gnd 0.005922f
C4308 vdd.n2470 gnd 0.005922f
C4309 vdd.n2471 gnd 0.005922f
C4310 vdd.n2472 gnd 0.005922f
C4311 vdd.n2473 gnd 0.005922f
C4312 vdd.n2474 gnd 0.005922f
C4313 vdd.n2475 gnd 0.005922f
C4314 vdd.n2476 gnd 0.378218f
C4315 vdd.n2477 gnd 0.005922f
C4316 vdd.n2478 gnd 0.005922f
C4317 vdd.n2479 gnd 0.005922f
C4318 vdd.n2480 gnd 0.012971f
C4319 vdd.n2481 gnd 0.012971f
C4320 vdd.n2482 gnd 0.01385f
C4321 vdd.n2483 gnd 0.01385f
C4322 vdd.n2484 gnd 0.005922f
C4323 vdd.n2485 gnd 0.005922f
C4324 vdd.n2486 gnd 0.005922f
C4325 vdd.n2487 gnd 0.004572f
C4326 vdd.n2488 gnd 0.008463f
C4327 vdd.n2489 gnd 0.004311f
C4328 vdd.n2490 gnd 0.005922f
C4329 vdd.n2491 gnd 0.005922f
C4330 vdd.n2492 gnd 0.005922f
C4331 vdd.n2493 gnd 0.005922f
C4332 vdd.n2494 gnd 0.005922f
C4333 vdd.n2495 gnd 0.005922f
C4334 vdd.n2496 gnd 0.005922f
C4335 vdd.n2497 gnd 0.005922f
C4336 vdd.n2498 gnd 0.005922f
C4337 vdd.n2499 gnd 0.005922f
C4338 vdd.n2500 gnd 0.005922f
C4339 vdd.n2501 gnd 0.005922f
C4340 vdd.n2502 gnd 0.005922f
C4341 vdd.n2503 gnd 0.005922f
C4342 vdd.n2504 gnd 0.005922f
C4343 vdd.n2505 gnd 0.005922f
C4344 vdd.n2506 gnd 0.005922f
C4345 vdd.n2507 gnd 0.005922f
C4346 vdd.n2508 gnd 0.005922f
C4347 vdd.n2509 gnd 0.005922f
C4348 vdd.n2510 gnd 0.005922f
C4349 vdd.n2511 gnd 0.005922f
C4350 vdd.n2512 gnd 0.005922f
C4351 vdd.n2513 gnd 0.005922f
C4352 vdd.n2514 gnd 0.005922f
C4353 vdd.n2515 gnd 0.005922f
C4354 vdd.n2516 gnd 0.005922f
C4355 vdd.n2517 gnd 0.005922f
C4356 vdd.n2518 gnd 0.005922f
C4357 vdd.n2519 gnd 0.005922f
C4358 vdd.n2520 gnd 0.005922f
C4359 vdd.n2521 gnd 0.005922f
C4360 vdd.n2522 gnd 0.005922f
C4361 vdd.n2523 gnd 0.005922f
C4362 vdd.n2524 gnd 0.005922f
C4363 vdd.n2525 gnd 0.005922f
C4364 vdd.n2526 gnd 0.005922f
C4365 vdd.n2527 gnd 0.005922f
C4366 vdd.n2528 gnd 0.005922f
C4367 vdd.n2529 gnd 0.005922f
C4368 vdd.n2530 gnd 0.005922f
C4369 vdd.n2531 gnd 0.005922f
C4370 vdd.n2532 gnd 0.005922f
C4371 vdd.n2533 gnd 0.005922f
C4372 vdd.n2534 gnd 0.005922f
C4373 vdd.n2535 gnd 0.005922f
C4374 vdd.n2536 gnd 0.005922f
C4375 vdd.n2537 gnd 0.005922f
C4376 vdd.n2538 gnd 0.005922f
C4377 vdd.n2539 gnd 0.005922f
C4378 vdd.n2540 gnd 0.005922f
C4379 vdd.n2541 gnd 0.005922f
C4380 vdd.n2542 gnd 0.005922f
C4381 vdd.n2543 gnd 0.005922f
C4382 vdd.n2544 gnd 0.005922f
C4383 vdd.n2545 gnd 0.005922f
C4384 vdd.n2546 gnd 0.005922f
C4385 vdd.n2547 gnd 0.005922f
C4386 vdd.n2548 gnd 0.005922f
C4387 vdd.n2549 gnd 0.01385f
C4388 vdd.n2550 gnd 0.01385f
C4389 vdd.n2552 gnd 0.738638f
C4390 vdd.n2554 gnd 0.01385f
C4391 vdd.n2555 gnd 0.01385f
C4392 vdd.n2556 gnd 0.012971f
C4393 vdd.n2557 gnd 0.005922f
C4394 vdd.n2558 gnd 0.005922f
C4395 vdd.n2559 gnd 0.320373f
C4396 vdd.n2560 gnd 0.005922f
C4397 vdd.n2561 gnd 0.005922f
C4398 vdd.n2562 gnd 0.005922f
C4399 vdd.n2563 gnd 0.005922f
C4400 vdd.n2564 gnd 0.005922f
C4401 vdd.n2565 gnd 0.36042f
C4402 vdd.n2566 gnd 0.005922f
C4403 vdd.n2567 gnd 0.005922f
C4404 vdd.n2568 gnd 0.005922f
C4405 vdd.n2569 gnd 0.005922f
C4406 vdd.n2570 gnd 0.005922f
C4407 vdd.n2571 gnd 0.605149f
C4408 vdd.n2572 gnd 0.005922f
C4409 vdd.n2573 gnd 0.005922f
C4410 vdd.n2574 gnd 0.005922f
C4411 vdd.n2575 gnd 0.005922f
C4412 vdd.n2576 gnd 0.005922f
C4413 vdd.n2577 gnd 0.400466f
C4414 vdd.n2578 gnd 0.005922f
C4415 vdd.n2579 gnd 0.005922f
C4416 vdd.n2580 gnd 0.005922f
C4417 vdd.n2581 gnd 0.005922f
C4418 vdd.n2582 gnd 0.005922f
C4419 vdd.n2583 gnd 0.533955f
C4420 vdd.n2584 gnd 0.005922f
C4421 vdd.n2585 gnd 0.005922f
C4422 vdd.n2586 gnd 0.005922f
C4423 vdd.n2587 gnd 0.005922f
C4424 vdd.n2588 gnd 0.005922f
C4425 vdd.n2589 gnd 0.485009f
C4426 vdd.n2590 gnd 0.005922f
C4427 vdd.n2591 gnd 0.005922f
C4428 vdd.n2592 gnd 0.005922f
C4429 vdd.n2593 gnd 0.005922f
C4430 vdd.n2594 gnd 0.005922f
C4431 vdd.n2595 gnd 0.35152f
C4432 vdd.n2596 gnd 0.005922f
C4433 vdd.n2597 gnd 0.005922f
C4434 vdd.n2598 gnd 0.005922f
C4435 vdd.n2599 gnd 0.005922f
C4436 vdd.n2600 gnd 0.005922f
C4437 vdd.n2601 gnd 0.191334f
C4438 vdd.n2602 gnd 0.005922f
C4439 vdd.n2603 gnd 0.005922f
C4440 vdd.n2604 gnd 0.005922f
C4441 vdd.n2605 gnd 0.005922f
C4442 vdd.n2606 gnd 0.005922f
C4443 vdd.n2607 gnd 0.520606f
C4444 vdd.n2608 gnd 0.005922f
C4445 vdd.n2609 gnd 0.005922f
C4446 vdd.n2610 gnd 0.005922f
C4447 vdd.n2611 gnd 0.005922f
C4448 vdd.n2612 gnd 0.005922f
C4449 vdd.n2613 gnd 0.605149f
C4450 vdd.n2614 gnd 0.005922f
C4451 vdd.n2615 gnd 0.005922f
C4452 vdd.n2616 gnd 0.003832f
C4453 vdd.n2617 gnd 0.017154f
C4454 vdd.n2618 gnd 0.005051f
C4455 vdd.n2619 gnd 0.005922f
C4456 vdd.n2620 gnd 0.516157f
C4457 vdd.n2621 gnd 0.005922f
C4458 vdd.n2622 gnd 0.005922f
C4459 vdd.n2623 gnd 0.005922f
C4460 vdd.n2624 gnd 0.005922f
C4461 vdd.n2625 gnd 0.005922f
C4462 vdd.n2626 gnd 0.422714f
C4463 vdd.n2627 gnd 0.005922f
C4464 vdd.n2628 gnd 0.005922f
C4465 vdd.n2629 gnd 0.005922f
C4466 vdd.n2630 gnd 0.005922f
C4467 vdd.n2631 gnd 0.005922f
C4468 vdd.n2632 gnd 0.315923f
C4469 vdd.n2633 gnd 0.005922f
C4470 vdd.n2634 gnd 0.005922f
C4471 vdd.n2635 gnd 0.005922f
C4472 vdd.n2636 gnd 0.005922f
C4473 vdd.n2637 gnd 0.005922f
C4474 vdd.n2638 gnd 0.605149f
C4475 vdd.n2639 gnd 0.005922f
C4476 vdd.n2640 gnd 0.005922f
C4477 vdd.n2641 gnd 0.005922f
C4478 vdd.n2642 gnd 0.005922f
C4479 vdd.n2643 gnd 0.005922f
C4480 vdd.n2644 gnd 0.005922f
C4481 vdd.n2646 gnd 0.005922f
C4482 vdd.n2647 gnd 0.005922f
C4483 vdd.n2649 gnd 0.005922f
C4484 vdd.n2650 gnd 0.005922f
C4485 vdd.n2653 gnd 0.005922f
C4486 vdd.n2654 gnd 0.005922f
C4487 vdd.n2655 gnd 0.005922f
C4488 vdd.n2656 gnd 0.005922f
C4489 vdd.n2658 gnd 0.005922f
C4490 vdd.n2659 gnd 0.005922f
C4491 vdd.n2660 gnd 0.005922f
C4492 vdd.n2661 gnd 0.005922f
C4493 vdd.n2662 gnd 0.005922f
C4494 vdd.n2663 gnd 0.005922f
C4495 vdd.n2665 gnd 0.005922f
C4496 vdd.n2666 gnd 0.005922f
C4497 vdd.n2667 gnd 0.005922f
C4498 vdd.n2668 gnd 0.005922f
C4499 vdd.n2669 gnd 0.005922f
C4500 vdd.n2670 gnd 0.005922f
C4501 vdd.n2672 gnd 0.005922f
C4502 vdd.n2673 gnd 0.005922f
C4503 vdd.n2674 gnd 0.005922f
C4504 vdd.n2675 gnd 0.005922f
C4505 vdd.n2676 gnd 0.005922f
C4506 vdd.n2677 gnd 0.005922f
C4507 vdd.n2679 gnd 0.005922f
C4508 vdd.n2680 gnd 0.01385f
C4509 vdd.n2681 gnd 0.01385f
C4510 vdd.n2682 gnd 0.012971f
C4511 vdd.n2683 gnd 0.005922f
C4512 vdd.n2684 gnd 0.005922f
C4513 vdd.n2685 gnd 0.005922f
C4514 vdd.n2686 gnd 0.005922f
C4515 vdd.n2687 gnd 0.005922f
C4516 vdd.n2688 gnd 0.005922f
C4517 vdd.n2689 gnd 0.605149f
C4518 vdd.n2690 gnd 0.005922f
C4519 vdd.n2691 gnd 0.005922f
C4520 vdd.n2692 gnd 0.005922f
C4521 vdd.n2693 gnd 0.005922f
C4522 vdd.n2694 gnd 0.005922f
C4523 vdd.n2695 gnd 0.396017f
C4524 vdd.n2696 gnd 0.005922f
C4525 vdd.n2697 gnd 0.005922f
C4526 vdd.n2698 gnd 0.005922f
C4527 vdd.n2699 gnd 0.013707f
C4528 vdd.n2700 gnd 0.013114f
C4529 vdd.n2701 gnd 0.01385f
C4530 vdd.n2703 gnd 0.005922f
C4531 vdd.n2704 gnd 0.005922f
C4532 vdd.n2705 gnd 0.004572f
C4533 vdd.n2706 gnd 0.008463f
C4534 vdd.n2707 gnd 0.004311f
C4535 vdd.n2708 gnd 0.005922f
C4536 vdd.n2709 gnd 0.005922f
C4537 vdd.n2711 gnd 0.005922f
C4538 vdd.n2712 gnd 0.005922f
C4539 vdd.n2713 gnd 0.005922f
C4540 vdd.n2714 gnd 0.005922f
C4541 vdd.n2715 gnd 0.005922f
C4542 vdd.n2716 gnd 0.005922f
C4543 vdd.n2718 gnd 0.005922f
C4544 vdd.n2719 gnd 0.005922f
C4545 vdd.n2720 gnd 0.005922f
C4546 vdd.n2721 gnd 0.005922f
C4547 vdd.n2722 gnd 0.005922f
C4548 vdd.n2723 gnd 0.005922f
C4549 vdd.n2725 gnd 0.005922f
C4550 vdd.n2726 gnd 0.005922f
C4551 vdd.n2727 gnd 0.005922f
C4552 vdd.n2728 gnd 0.005922f
C4553 vdd.n2729 gnd 0.005922f
C4554 vdd.n2730 gnd 0.005922f
C4555 vdd.n2732 gnd 0.005922f
C4556 vdd.n2733 gnd 0.005922f
C4557 vdd.n2734 gnd 0.005922f
C4558 vdd.n2736 gnd 0.005922f
C4559 vdd.n2737 gnd 0.005922f
C4560 vdd.n2738 gnd 0.005922f
C4561 vdd.n2739 gnd 0.005922f
C4562 vdd.n2740 gnd 0.005922f
C4563 vdd.n2741 gnd 0.005922f
C4564 vdd.n2743 gnd 0.005922f
C4565 vdd.n2744 gnd 0.005922f
C4566 vdd.n2745 gnd 0.005922f
C4567 vdd.n2746 gnd 0.005922f
C4568 vdd.n2747 gnd 0.005922f
C4569 vdd.n2748 gnd 0.005922f
C4570 vdd.n2750 gnd 0.005922f
C4571 vdd.n2751 gnd 0.005922f
C4572 vdd.n2752 gnd 0.005922f
C4573 vdd.n2753 gnd 0.005922f
C4574 vdd.n2754 gnd 0.005922f
C4575 vdd.n2755 gnd 0.005922f
C4576 vdd.n2757 gnd 0.005922f
C4577 vdd.n2758 gnd 0.005922f
C4578 vdd.n2760 gnd 0.005922f
C4579 vdd.n2761 gnd 0.005922f
C4580 vdd.n2762 gnd 0.01385f
C4581 vdd.n2763 gnd 0.012971f
C4582 vdd.n2764 gnd 0.012971f
C4583 vdd.n2765 gnd 0.854328f
C4584 vdd.n2766 gnd 0.012971f
C4585 vdd.n2767 gnd 0.01385f
C4586 vdd.n2768 gnd 0.013114f
C4587 vdd.n2769 gnd 0.005922f
C4588 vdd.n2770 gnd 0.004572f
C4589 vdd.n2771 gnd 0.005922f
C4590 vdd.n2773 gnd 0.005922f
C4591 vdd.n2774 gnd 0.005922f
C4592 vdd.n2775 gnd 0.005922f
C4593 vdd.n2776 gnd 0.005922f
C4594 vdd.n2777 gnd 0.005922f
C4595 vdd.n2778 gnd 0.005922f
C4596 vdd.n2780 gnd 0.005922f
C4597 vdd.n2781 gnd 0.005922f
C4598 vdd.n2782 gnd 0.005922f
C4599 vdd.n2783 gnd 0.005922f
C4600 vdd.n2784 gnd 0.005922f
C4601 vdd.n2785 gnd 0.005922f
C4602 vdd.n2787 gnd 0.005922f
C4603 vdd.n2788 gnd 0.005922f
C4604 vdd.n2789 gnd 0.005922f
C4605 vdd.n2790 gnd 0.005922f
C4606 vdd.n2791 gnd 0.005922f
C4607 vdd.n2792 gnd 0.005922f
C4608 vdd.n2794 gnd 0.005922f
C4609 vdd.n2795 gnd 0.005922f
C4610 vdd.n2797 gnd 0.005922f
C4611 vdd.n2798 gnd 0.020337f
C4612 vdd.n2799 gnd 0.661949f
C4613 vdd.n2800 gnd 0.007489f
C4614 vdd.n2801 gnd 0.021709f
C4615 vdd.n2802 gnd 0.003329f
C4616 vdd.t20 gnd 0.107132f
C4617 vdd.t21 gnd 0.114495f
C4618 vdd.t18 gnd 0.139914f
C4619 vdd.n2803 gnd 0.179349f
C4620 vdd.n2804 gnd 0.150686f
C4621 vdd.n2805 gnd 0.010794f
C4622 vdd.n2806 gnd 0.008708f
C4623 vdd.n2807 gnd 0.00368f
C4624 vdd.n2808 gnd 0.007009f
C4625 vdd.n2809 gnd 0.008708f
C4626 vdd.n2810 gnd 0.008708f
C4627 vdd.n2811 gnd 0.007009f
C4628 vdd.n2812 gnd 0.007009f
C4629 vdd.n2813 gnd 0.008708f
C4630 vdd.n2814 gnd 0.008708f
C4631 vdd.n2815 gnd 0.007009f
C4632 vdd.n2816 gnd 0.007009f
C4633 vdd.n2817 gnd 0.008708f
C4634 vdd.n2818 gnd 0.008708f
C4635 vdd.n2819 gnd 0.007009f
C4636 vdd.n2820 gnd 0.007009f
C4637 vdd.n2821 gnd 0.008708f
C4638 vdd.n2822 gnd 0.008708f
C4639 vdd.n2823 gnd 0.007009f
C4640 vdd.n2824 gnd 0.007009f
C4641 vdd.n2825 gnd 0.008708f
C4642 vdd.n2826 gnd 0.008708f
C4643 vdd.n2827 gnd 0.007009f
C4644 vdd.n2828 gnd 0.007009f
C4645 vdd.n2829 gnd 0.008708f
C4646 vdd.n2830 gnd 0.008708f
C4647 vdd.n2831 gnd 0.007009f
C4648 vdd.n2832 gnd 0.007009f
C4649 vdd.n2833 gnd 0.008708f
C4650 vdd.n2834 gnd 0.008708f
C4651 vdd.n2835 gnd 0.007009f
C4652 vdd.n2836 gnd 0.007009f
C4653 vdd.n2837 gnd 0.008708f
C4654 vdd.n2838 gnd 0.008708f
C4655 vdd.n2839 gnd 0.007009f
C4656 vdd.n2840 gnd 0.007009f
C4657 vdd.n2841 gnd 0.008708f
C4658 vdd.n2842 gnd 0.008708f
C4659 vdd.n2843 gnd 0.007009f
C4660 vdd.n2844 gnd 0.008708f
C4661 vdd.n2845 gnd 0.008708f
C4662 vdd.n2846 gnd 0.007009f
C4663 vdd.n2847 gnd 0.008708f
C4664 vdd.n2848 gnd 0.008708f
C4665 vdd.n2849 gnd 0.008708f
C4666 vdd.n2850 gnd 0.014298f
C4667 vdd.n2851 gnd 0.008708f
C4668 vdd.n2852 gnd 0.008708f
C4669 vdd.n2853 gnd 0.004766f
C4670 vdd.n2854 gnd 0.007009f
C4671 vdd.n2855 gnd 0.008708f
C4672 vdd.n2856 gnd 0.008708f
C4673 vdd.n2857 gnd 0.007009f
C4674 vdd.n2858 gnd 0.007009f
C4675 vdd.n2859 gnd 0.008708f
C4676 vdd.n2860 gnd 0.008708f
C4677 vdd.n2861 gnd 0.007009f
C4678 vdd.n2862 gnd 0.007009f
C4679 vdd.n2863 gnd 0.008708f
C4680 vdd.n2864 gnd 0.008708f
C4681 vdd.n2865 gnd 0.007009f
C4682 vdd.n2866 gnd 0.007009f
C4683 vdd.n2867 gnd 0.008708f
C4684 vdd.n2868 gnd 0.008708f
C4685 vdd.n2869 gnd 0.007009f
C4686 vdd.n2870 gnd 0.007009f
C4687 vdd.n2871 gnd 0.008708f
C4688 vdd.n2872 gnd 0.008708f
C4689 vdd.n2873 gnd 0.007009f
C4690 vdd.n2874 gnd 0.007009f
C4691 vdd.n2875 gnd 0.008708f
C4692 vdd.n2876 gnd 0.008708f
C4693 vdd.n2877 gnd 0.007009f
C4694 vdd.n2878 gnd 0.007009f
C4695 vdd.n2879 gnd 0.008708f
C4696 vdd.n2880 gnd 0.008708f
C4697 vdd.n2881 gnd 0.007009f
C4698 vdd.n2882 gnd 0.007009f
C4699 vdd.n2883 gnd 0.008708f
C4700 vdd.n2884 gnd 0.008708f
C4701 vdd.n2885 gnd 0.007009f
C4702 vdd.n2886 gnd 0.007009f
C4703 vdd.n2887 gnd 0.008708f
C4704 vdd.n2888 gnd 0.008708f
C4705 vdd.n2889 gnd 0.007009f
C4706 vdd.n2890 gnd 0.008708f
C4707 vdd.n2891 gnd 0.008708f
C4708 vdd.n2892 gnd 0.007009f
C4709 vdd.n2893 gnd 0.008708f
C4710 vdd.n2894 gnd 0.008708f
C4711 vdd.n2895 gnd 0.008708f
C4712 vdd.t40 gnd 0.107132f
C4713 vdd.t41 gnd 0.114495f
C4714 vdd.t39 gnd 0.139914f
C4715 vdd.n2896 gnd 0.179349f
C4716 vdd.n2897 gnd 0.150686f
C4717 vdd.n2898 gnd 0.014298f
C4718 vdd.n2899 gnd 0.008708f
C4719 vdd.n2900 gnd 0.008708f
C4720 vdd.n2901 gnd 0.005852f
C4721 vdd.n2902 gnd 0.007009f
C4722 vdd.n2903 gnd 0.008708f
C4723 vdd.n2904 gnd 0.008708f
C4724 vdd.n2905 gnd 0.007009f
C4725 vdd.n2906 gnd 0.007009f
C4726 vdd.n2907 gnd 0.008708f
C4727 vdd.n2908 gnd 0.008708f
C4728 vdd.n2909 gnd 0.007009f
C4729 vdd.n2910 gnd 0.007009f
C4730 vdd.n2911 gnd 0.008708f
C4731 vdd.n2912 gnd 0.008708f
C4732 vdd.n2913 gnd 0.007009f
C4733 vdd.n2914 gnd 0.007009f
C4734 vdd.n2915 gnd 0.008708f
C4735 vdd.n2916 gnd 0.008708f
C4736 vdd.n2917 gnd 0.007009f
C4737 vdd.n2918 gnd 0.007009f
C4738 vdd.n2919 gnd 0.008708f
C4739 vdd.n2920 gnd 0.008708f
C4740 vdd.n2921 gnd 0.007009f
C4741 vdd.n2922 gnd 0.007009f
C4742 vdd.n2923 gnd 0.008708f
C4743 vdd.n2924 gnd 0.008708f
C4744 vdd.n2925 gnd 0.007009f
C4745 vdd.n2926 gnd 0.007009f
C4746 vdd.n2928 gnd 0.661949f
C4747 vdd.n2930 gnd 0.007009f
C4748 vdd.n2931 gnd 0.008708f
C4749 vdd.n2932 gnd 7.92923f
C4750 vdd.n2934 gnd 0.021709f
C4751 vdd.n2935 gnd 0.005817f
C4752 vdd.n2936 gnd 0.021709f
C4753 vdd.n2937 gnd 0.021222f
C4754 vdd.n2938 gnd 0.008708f
C4755 vdd.n2939 gnd 0.007009f
C4756 vdd.n2940 gnd 0.008708f
C4757 vdd.n2941 gnd 0.556203f
C4758 vdd.n2942 gnd 0.008708f
C4759 vdd.n2943 gnd 0.007009f
C4760 vdd.n2944 gnd 0.008708f
C4761 vdd.n2945 gnd 0.008708f
C4762 vdd.n2946 gnd 0.008708f
C4763 vdd.n2947 gnd 0.007009f
C4764 vdd.n2948 gnd 0.008708f
C4765 vdd.n2949 gnd 0.707491f
C4766 vdd.n2950 gnd 0.889925f
C4767 vdd.n2951 gnd 0.008708f
C4768 vdd.n2952 gnd 0.007009f
C4769 vdd.n2953 gnd 0.008708f
C4770 vdd.n2954 gnd 0.008708f
C4771 vdd.n2955 gnd 0.008708f
C4772 vdd.n2956 gnd 0.007009f
C4773 vdd.n2957 gnd 0.008708f
C4774 vdd.n2958 gnd 0.627397f
C4775 vdd.n2959 gnd 0.008708f
C4776 vdd.n2960 gnd 0.007009f
C4777 vdd.n2961 gnd 0.008708f
C4778 vdd.n2962 gnd 0.008708f
C4779 vdd.n2963 gnd 0.008708f
C4780 vdd.n2964 gnd 0.007009f
C4781 vdd.n2965 gnd 0.008708f
C4782 vdd.t78 gnd 0.444963f
C4783 vdd.n2966 gnd 0.738638f
C4784 vdd.n2967 gnd 0.008708f
C4785 vdd.n2968 gnd 0.007009f
C4786 vdd.n2969 gnd 0.008708f
C4787 vdd.n2970 gnd 0.008708f
C4788 vdd.n2971 gnd 0.008708f
C4789 vdd.n2972 gnd 0.007009f
C4790 vdd.n2973 gnd 0.008708f
C4791 vdd.n2974 gnd 0.698591f
C4792 vdd.n2975 gnd 0.008708f
C4793 vdd.n2976 gnd 0.007009f
C4794 vdd.n2977 gnd 0.008708f
C4795 vdd.n2978 gnd 0.008708f
C4796 vdd.n2979 gnd 0.008708f
C4797 vdd.n2980 gnd 0.007009f
C4798 vdd.n2981 gnd 0.007009f
C4799 vdd.n2982 gnd 0.007009f
C4800 vdd.n2983 gnd 0.008708f
C4801 vdd.n2984 gnd 0.008708f
C4802 vdd.n2985 gnd 0.008708f
C4803 vdd.n2986 gnd 0.007009f
C4804 vdd.n2987 gnd 0.007009f
C4805 vdd.n2988 gnd 0.007009f
C4806 vdd.n2989 gnd 0.008708f
C4807 vdd.n2990 gnd 0.008708f
C4808 vdd.n2991 gnd 0.008708f
C4809 vdd.n2992 gnd 0.007009f
C4810 vdd.n2993 gnd 0.007009f
C4811 vdd.n2994 gnd 0.005817f
C4812 vdd.n2995 gnd 0.021222f
C4813 vdd.n2996 gnd 0.021709f
C4814 vdd.n2998 gnd 0.021709f
C4815 vdd.n2999 gnd 0.003329f
C4816 vdd.t77 gnd 0.107132f
C4817 vdd.t76 gnd 0.114495f
C4818 vdd.t75 gnd 0.139914f
C4819 vdd.n3000 gnd 0.179349f
C4820 vdd.n3001 gnd 0.151387f
C4821 vdd.n3002 gnd 0.011495f
C4822 vdd.n3003 gnd 0.00368f
C4823 vdd.n3004 gnd 0.007009f
C4824 vdd.n3005 gnd 0.008708f
C4825 vdd.n3007 gnd 0.008708f
C4826 vdd.n3008 gnd 0.008708f
C4827 vdd.n3009 gnd 0.007009f
C4828 vdd.n3010 gnd 0.007009f
C4829 vdd.n3011 gnd 0.007009f
C4830 vdd.n3012 gnd 0.008708f
C4831 vdd.n3014 gnd 0.008708f
C4832 vdd.n3015 gnd 0.008708f
C4833 vdd.n3016 gnd 0.007009f
C4834 vdd.n3017 gnd 0.007009f
C4835 vdd.n3018 gnd 0.007009f
C4836 vdd.n3019 gnd 0.008708f
C4837 vdd.n3021 gnd 0.008708f
C4838 vdd.n3022 gnd 0.008708f
C4839 vdd.n3023 gnd 0.007009f
C4840 vdd.n3024 gnd 0.007009f
C4841 vdd.n3025 gnd 0.007009f
C4842 vdd.n3026 gnd 0.008708f
C4843 vdd.n3028 gnd 0.008708f
C4844 vdd.n3029 gnd 0.008708f
C4845 vdd.n3030 gnd 0.007009f
C4846 vdd.n3031 gnd 0.007009f
C4847 vdd.n3032 gnd 0.007009f
C4848 vdd.n3033 gnd 0.008708f
C4849 vdd.n3035 gnd 0.008708f
C4850 vdd.n3036 gnd 0.008708f
C4851 vdd.n3037 gnd 0.007009f
C4852 vdd.n3038 gnd 0.008708f
C4853 vdd.n3039 gnd 0.008708f
C4854 vdd.n3040 gnd 0.008708f
C4855 vdd.n3041 gnd 0.014999f
C4856 vdd.n3042 gnd 0.004766f
C4857 vdd.n3043 gnd 0.007009f
C4858 vdd.n3044 gnd 0.008708f
C4859 vdd.n3046 gnd 0.008708f
C4860 vdd.n3047 gnd 0.008708f
C4861 vdd.n3048 gnd 0.007009f
C4862 vdd.n3049 gnd 0.007009f
C4863 vdd.n3050 gnd 0.007009f
C4864 vdd.n3051 gnd 0.008708f
C4865 vdd.n3053 gnd 0.008708f
C4866 vdd.n3054 gnd 0.008708f
C4867 vdd.n3055 gnd 0.007009f
C4868 vdd.n3056 gnd 0.007009f
C4869 vdd.n3057 gnd 0.007009f
C4870 vdd.n3058 gnd 0.008708f
C4871 vdd.n3060 gnd 0.008708f
C4872 vdd.n3061 gnd 0.008708f
C4873 vdd.n3062 gnd 0.007009f
C4874 vdd.n3063 gnd 0.007009f
C4875 vdd.n3064 gnd 0.007009f
C4876 vdd.n3065 gnd 0.008708f
C4877 vdd.n3067 gnd 0.008708f
C4878 vdd.n3068 gnd 0.008708f
C4879 vdd.n3069 gnd 0.007009f
C4880 vdd.n3070 gnd 0.007009f
C4881 vdd.n3071 gnd 0.007009f
C4882 vdd.n3072 gnd 0.008708f
C4883 vdd.n3074 gnd 0.008708f
C4884 vdd.n3075 gnd 0.008708f
C4885 vdd.n3076 gnd 0.007009f
C4886 vdd.n3077 gnd 0.008708f
C4887 vdd.n3078 gnd 0.008708f
C4888 vdd.n3079 gnd 0.008708f
C4889 vdd.n3080 gnd 0.014999f
C4890 vdd.n3081 gnd 0.005852f
C4891 vdd.n3082 gnd 0.007009f
C4892 vdd.n3083 gnd 0.008708f
C4893 vdd.n3085 gnd 0.008708f
C4894 vdd.n3086 gnd 0.008708f
C4895 vdd.n3087 gnd 0.007009f
C4896 vdd.n3088 gnd 0.007009f
C4897 vdd.n3089 gnd 0.007009f
C4898 vdd.n3090 gnd 0.008708f
C4899 vdd.n3092 gnd 0.008708f
C4900 vdd.n3093 gnd 0.008708f
C4901 vdd.n3094 gnd 0.007009f
C4902 vdd.n3095 gnd 0.007009f
C4903 vdd.n3096 gnd 0.007009f
C4904 vdd.n3097 gnd 0.008708f
C4905 vdd.n3099 gnd 0.008708f
C4906 vdd.n3100 gnd 0.008708f
C4907 vdd.n3101 gnd 0.007009f
C4908 vdd.n3102 gnd 0.007009f
C4909 vdd.n3103 gnd 0.007009f
C4910 vdd.n3104 gnd 0.008708f
C4911 vdd.n3106 gnd 0.008708f
C4912 vdd.n3107 gnd 0.008708f
C4913 vdd.n3109 gnd 0.008708f
C4914 vdd.n3110 gnd 0.007009f
C4915 vdd.n3111 gnd 0.007009f
C4916 vdd.n3112 gnd 0.005817f
C4917 vdd.n3113 gnd 0.021709f
C4918 vdd.n3114 gnd 0.021222f
C4919 vdd.n3115 gnd 0.005817f
C4920 vdd.n3116 gnd 0.021222f
C4921 vdd.n3117 gnd 1.31264f
C4922 vdd.t7 gnd 0.444963f
C4923 vdd.n3118 gnd 0.467211f
C4924 vdd.n3119 gnd 0.889925f
C4925 vdd.n3120 gnd 0.008708f
C4926 vdd.n3121 gnd 0.007009f
C4927 vdd.n3122 gnd 0.007009f
C4928 vdd.n3123 gnd 0.007009f
C4929 vdd.n3124 gnd 0.008708f
C4930 vdd.n3125 gnd 0.796483f
C4931 vdd.t84 gnd 0.444963f
C4932 vdd.n3126 gnd 0.538405f
C4933 vdd.n3127 gnd 0.645196f
C4934 vdd.n3128 gnd 0.008708f
C4935 vdd.n3129 gnd 0.007009f
C4936 vdd.n3130 gnd 0.007009f
C4937 vdd.n3131 gnd 0.007009f
C4938 vdd.n3132 gnd 0.008708f
C4939 vdd.n3133 gnd 0.493909f
C4940 vdd.t160 gnd 0.444963f
C4941 vdd.n3134 gnd 0.738638f
C4942 vdd.t164 gnd 0.444963f
C4943 vdd.n3135 gnd 0.547304f
C4944 vdd.n3136 gnd 0.008708f
C4945 vdd.n3137 gnd 0.007009f
C4946 vdd.n3138 gnd 0.006693f
C4947 vdd.n3139 gnd 0.513636f
C4948 vdd.n3140 gnd 1.86896f
C4949 a_n2140_13878.t11 gnd 0.186868f
C4950 a_n2140_13878.t10 gnd 0.186868f
C4951 a_n2140_13878.t5 gnd 0.186868f
C4952 a_n2140_13878.n0 gnd 1.47299f
C4953 a_n2140_13878.t2 gnd 0.186868f
C4954 a_n2140_13878.t4 gnd 0.186868f
C4955 a_n2140_13878.n1 gnd 1.47143f
C4956 a_n2140_13878.n2 gnd 2.05603f
C4957 a_n2140_13878.t12 gnd 0.186868f
C4958 a_n2140_13878.t3 gnd 0.186868f
C4959 a_n2140_13878.n3 gnd 1.47143f
C4960 a_n2140_13878.n4 gnd 1.00289f
C4961 a_n2140_13878.t9 gnd 0.186868f
C4962 a_n2140_13878.t1 gnd 0.186868f
C4963 a_n2140_13878.n5 gnd 1.47143f
C4964 a_n2140_13878.n6 gnd 4.06212f
C4965 a_n2140_13878.t23 gnd 1.74974f
C4966 a_n2140_13878.t16 gnd 0.186868f
C4967 a_n2140_13878.t17 gnd 0.186868f
C4968 a_n2140_13878.n7 gnd 1.3163f
C4969 a_n2140_13878.n8 gnd 1.47077f
C4970 a_n2140_13878.t18 gnd 1.74626f
C4971 a_n2140_13878.n9 gnd 0.740113f
C4972 a_n2140_13878.t19 gnd 1.74626f
C4973 a_n2140_13878.n10 gnd 0.740113f
C4974 a_n2140_13878.t22 gnd 0.186868f
C4975 a_n2140_13878.t21 gnd 0.186868f
C4976 a_n2140_13878.n11 gnd 1.3163f
C4977 a_n2140_13878.n12 gnd 0.74728f
C4978 a_n2140_13878.t20 gnd 1.74626f
C4979 a_n2140_13878.n13 gnd 2.09583f
C4980 a_n2140_13878.n14 gnd 2.85974f
C4981 a_n2140_13878.t6 gnd 0.186868f
C4982 a_n2140_13878.t7 gnd 0.186868f
C4983 a_n2140_13878.n15 gnd 1.47142f
C4984 a_n2140_13878.n16 gnd 2.01665f
C4985 a_n2140_13878.t13 gnd 0.186868f
C4986 a_n2140_13878.t14 gnd 0.186868f
C4987 a_n2140_13878.n17 gnd 1.47143f
C4988 a_n2140_13878.n18 gnd 0.651951f
C4989 a_n2140_13878.t0 gnd 0.186868f
C4990 a_n2140_13878.t8 gnd 0.186868f
C4991 a_n2140_13878.n19 gnd 1.47143f
C4992 a_n2140_13878.n20 gnd 1.32263f
C4993 a_n2140_13878.n21 gnd 1.47386f
C4994 a_n2140_13878.t15 gnd 0.186868f
C4995 a_n2408_n452.n0 gnd 3.95093f
C4996 a_n2408_n452.n1 gnd 2.90522f
C4997 a_n2408_n452.n2 gnd 3.88871f
C4998 a_n2408_n452.n3 gnd 0.820088f
C4999 a_n2408_n452.n4 gnd 0.82009f
C5000 a_n2408_n452.n5 gnd 0.668637f
C5001 a_n2408_n452.n6 gnd 0.204926f
C5002 a_n2408_n452.n7 gnd 0.150932f
C5003 a_n2408_n452.n8 gnd 0.237216f
C5004 a_n2408_n452.n9 gnd 0.183222f
C5005 a_n2408_n452.n10 gnd 0.204926f
C5006 a_n2408_n452.n11 gnd 1.1184f
C5007 a_n2408_n452.n12 gnd 0.150932f
C5008 a_n2408_n452.n13 gnd 0.722632f
C5009 a_n2408_n452.n14 gnd 0.512478f
C5010 a_n2408_n452.n15 gnd 0.215976f
C5011 a_n2408_n452.n16 gnd 0.215976f
C5012 a_n2408_n452.n17 gnd 0.44388f
C5013 a_n2408_n452.n18 gnd 0.215976f
C5014 a_n2408_n452.n19 gnd 0.215976f
C5015 a_n2408_n452.n20 gnd 0.215976f
C5016 a_n2408_n452.n21 gnd 0.747109f
C5017 a_n2408_n452.n22 gnd 0.215976f
C5018 a_n2408_n452.n23 gnd 0.44388f
C5019 a_n2408_n452.n24 gnd 3.3281f
C5020 a_n2408_n452.n25 gnd 0.668661f
C5021 a_n2408_n452.n26 gnd 0.215976f
C5022 a_n2408_n452.n27 gnd 1.7781f
C5023 a_n2408_n452.n28 gnd 2.07945f
C5024 a_n2408_n452.n29 gnd 1.7781f
C5025 a_n2408_n452.n30 gnd 1.89786f
C5026 a_n2408_n452.n31 gnd 0.285304f
C5027 a_n2408_n452.n32 gnd 0.004854f
C5028 a_n2408_n452.n33 gnd 0.010499f
C5029 a_n2408_n452.n34 gnd 0.010499f
C5030 a_n2408_n452.n35 gnd 0.285304f
C5031 a_n2408_n452.n36 gnd 0.285304f
C5032 a_n2408_n452.n37 gnd 0.004854f
C5033 a_n2408_n452.n38 gnd 0.010499f
C5034 a_n2408_n452.n39 gnd 0.010499f
C5035 a_n2408_n452.n40 gnd 0.004854f
C5036 a_n2408_n452.n41 gnd 0.285304f
C5037 a_n2408_n452.n42 gnd 0.285304f
C5038 a_n2408_n452.n43 gnd 0.76008f
C5039 a_n2408_n452.n44 gnd 0.004854f
C5040 a_n2408_n452.n45 gnd 0.010499f
C5041 a_n2408_n452.n46 gnd 0.010499f
C5042 a_n2408_n452.n47 gnd 0.004854f
C5043 a_n2408_n452.n48 gnd 0.285304f
C5044 a_n2408_n452.n49 gnd 0.285304f
C5045 a_n2408_n452.n50 gnd 0.44388f
C5046 a_n2408_n452.n51 gnd 0.004854f
C5047 a_n2408_n452.n52 gnd 0.010499f
C5048 a_n2408_n452.n53 gnd 0.010499f
C5049 a_n2408_n452.n54 gnd 0.004854f
C5050 a_n2408_n452.n55 gnd 0.285304f
C5051 a_n2408_n452.n56 gnd 0.008362f
C5052 a_n2408_n452.n57 gnd 0.285304f
C5053 a_n2408_n452.n58 gnd 0.008362f
C5054 a_n2408_n452.n59 gnd 0.285304f
C5055 a_n2408_n452.n60 gnd 0.008362f
C5056 a_n2408_n452.n61 gnd 0.285304f
C5057 a_n2408_n452.n62 gnd 0.008362f
C5058 a_n2408_n452.n63 gnd 0.285304f
C5059 a_n2408_n452.n64 gnd 0.004854f
C5060 a_n2408_n452.n65 gnd 0.304392f
C5061 a_n2408_n452.t32 gnd 0.149803f
C5062 a_n2408_n452.t11 gnd 0.708488f
C5063 a_n2408_n452.t7 gnd 0.696812f
C5064 a_n2408_n452.t31 gnd 0.696812f
C5065 a_n2408_n452.n66 gnd 0.304392f
C5066 a_n2408_n452.t29 gnd 0.696812f
C5067 a_n2408_n452.t13 gnd 0.696812f
C5068 a_n2408_n452.t9 gnd 0.696812f
C5069 a_n2408_n452.t25 gnd 0.708488f
C5070 a_n2408_n452.t86 gnd 0.708488f
C5071 a_n2408_n452.t67 gnd 0.696812f
C5072 a_n2408_n452.t71 gnd 0.696812f
C5073 a_n2408_n452.n67 gnd 0.304392f
C5074 a_n2408_n452.t61 gnd 0.696812f
C5075 a_n2408_n452.t76 gnd 0.696812f
C5076 a_n2408_n452.t83 gnd 0.696812f
C5077 a_n2408_n452.n68 gnd 0.304392f
C5078 a_n2408_n452.t84 gnd 0.696812f
C5079 a_n2408_n452.t58 gnd 0.708488f
C5080 a_n2408_n452.t18 gnd 1.40268f
C5081 a_n2408_n452.t20 gnd 0.149803f
C5082 a_n2408_n452.t24 gnd 0.149803f
C5083 a_n2408_n452.n69 gnd 1.05521f
C5084 a_n2408_n452.t38 gnd 0.149803f
C5085 a_n2408_n452.t28 gnd 0.149803f
C5086 a_n2408_n452.n70 gnd 1.05521f
C5087 a_n2408_n452.t34 gnd 0.149803f
C5088 a_n2408_n452.t22 gnd 0.149803f
C5089 a_n2408_n452.n71 gnd 1.05521f
C5090 a_n2408_n452.t36 gnd 1.39988f
C5091 a_n2408_n452.t33 gnd 0.696812f
C5092 a_n2408_n452.n72 gnd 0.304392f
C5093 a_n2408_n452.t37 gnd 0.696812f
C5094 a_n2408_n452.t17 gnd 0.708488f
C5095 a_n2408_n452.t19 gnd 0.696812f
C5096 a_n2408_n452.t65 gnd 0.696812f
C5097 a_n2408_n452.n73 gnd 0.304392f
C5098 a_n2408_n452.t79 gnd 0.696812f
C5099 a_n2408_n452.t82 gnd 0.708488f
C5100 a_n2408_n452.t60 gnd 0.696812f
C5101 a_n2408_n452.n74 gnd 0.306874f
C5102 a_n2408_n452.t80 gnd 0.696812f
C5103 a_n2408_n452.n75 gnd 0.304392f
C5104 a_n2408_n452.n76 gnd 0.299809f
C5105 a_n2408_n452.t57 gnd 0.696812f
C5106 a_n2408_n452.n77 gnd 0.299809f
C5107 a_n2408_n452.t74 gnd 0.696812f
C5108 a_n2408_n452.n78 gnd 0.306874f
C5109 a_n2408_n452.t59 gnd 0.708488f
C5110 a_n2408_n452.n79 gnd 0.306874f
C5111 a_n2408_n452.t23 gnd 0.696812f
C5112 a_n2408_n452.n80 gnd 0.304392f
C5113 a_n2408_n452.n81 gnd 0.299809f
C5114 a_n2408_n452.t27 gnd 0.696812f
C5115 a_n2408_n452.n82 gnd 0.299809f
C5116 a_n2408_n452.t21 gnd 0.696812f
C5117 a_n2408_n452.n83 gnd 0.306874f
C5118 a_n2408_n452.t35 gnd 0.708488f
C5119 a_n2408_n452.n84 gnd 1.19872f
C5120 a_n2408_n452.t64 gnd 0.696812f
C5121 a_n2408_n452.n85 gnd 0.302472f
C5122 a_n2408_n452.t70 gnd 0.696812f
C5123 a_n2408_n452.n86 gnd 0.302472f
C5124 a_n2408_n452.t63 gnd 0.696812f
C5125 a_n2408_n452.n87 gnd 0.302472f
C5126 a_n2408_n452.t75 gnd 0.696812f
C5127 a_n2408_n452.n88 gnd 0.302472f
C5128 a_n2408_n452.t66 gnd 0.696812f
C5129 a_n2408_n452.n89 gnd 0.296979f
C5130 a_n2408_n452.t87 gnd 0.696812f
C5131 a_n2408_n452.n90 gnd 0.306363f
C5132 a_n2408_n452.t68 gnd 0.708488f
C5133 a_n2408_n452.t77 gnd 0.696812f
C5134 a_n2408_n452.n91 gnd 0.296979f
C5135 a_n2408_n452.t62 gnd 0.696812f
C5136 a_n2408_n452.n92 gnd 0.306363f
C5137 a_n2408_n452.t72 gnd 0.708488f
C5138 a_n2408_n452.t81 gnd 0.696812f
C5139 a_n2408_n452.n93 gnd 0.296979f
C5140 a_n2408_n452.t69 gnd 0.696812f
C5141 a_n2408_n452.n94 gnd 0.306363f
C5142 a_n2408_n452.t85 gnd 0.708488f
C5143 a_n2408_n452.t73 gnd 0.696812f
C5144 a_n2408_n452.n95 gnd 0.296979f
C5145 a_n2408_n452.t56 gnd 0.696812f
C5146 a_n2408_n452.n96 gnd 0.306363f
C5147 a_n2408_n452.t78 gnd 0.708488f
C5148 a_n2408_n452.n97 gnd 1.45046f
C5149 a_n2408_n452.n98 gnd 0.306874f
C5150 a_n2408_n452.n99 gnd 0.299809f
C5151 a_n2408_n452.n100 gnd 0.299809f
C5152 a_n2408_n452.n101 gnd 0.306874f
C5153 a_n2408_n452.t15 gnd 0.696812f
C5154 a_n2408_n452.n102 gnd 0.306874f
C5155 a_n2408_n452.t53 gnd 0.116514f
C5156 a_n2408_n452.t48 gnd 0.116514f
C5157 a_n2408_n452.n103 gnd 1.03184f
C5158 a_n2408_n452.t6 gnd 0.116514f
C5159 a_n2408_n452.t5 gnd 0.116514f
C5160 a_n2408_n452.n104 gnd 1.02955f
C5161 a_n2408_n452.t4 gnd 0.116514f
C5162 a_n2408_n452.t1 gnd 0.116514f
C5163 a_n2408_n452.n105 gnd 1.02955f
C5164 a_n2408_n452.t49 gnd 0.116514f
C5165 a_n2408_n452.t2 gnd 0.116514f
C5166 a_n2408_n452.n106 gnd 1.03184f
C5167 a_n2408_n452.t45 gnd 0.116514f
C5168 a_n2408_n452.t54 gnd 0.116514f
C5169 a_n2408_n452.n107 gnd 1.02955f
C5170 a_n2408_n452.t41 gnd 0.116514f
C5171 a_n2408_n452.t52 gnd 0.116514f
C5172 a_n2408_n452.n108 gnd 1.02955f
C5173 a_n2408_n452.t42 gnd 0.116514f
C5174 a_n2408_n452.t46 gnd 0.116514f
C5175 a_n2408_n452.n109 gnd 1.02956f
C5176 a_n2408_n452.t40 gnd 0.116514f
C5177 a_n2408_n452.t0 gnd 0.116514f
C5178 a_n2408_n452.n110 gnd 1.02956f
C5179 a_n2408_n452.t55 gnd 0.116514f
C5180 a_n2408_n452.t44 gnd 0.116514f
C5181 a_n2408_n452.n111 gnd 1.02956f
C5182 a_n2408_n452.t51 gnd 0.116514f
C5183 a_n2408_n452.t50 gnd 0.116514f
C5184 a_n2408_n452.n112 gnd 1.03184f
C5185 a_n2408_n452.t3 gnd 0.116514f
C5186 a_n2408_n452.t39 gnd 0.116514f
C5187 a_n2408_n452.n113 gnd 1.02956f
C5188 a_n2408_n452.t43 gnd 0.116514f
C5189 a_n2408_n452.t47 gnd 0.116514f
C5190 a_n2408_n452.n114 gnd 1.02956f
C5191 a_n2408_n452.n115 gnd 0.299809f
C5192 a_n2408_n452.n116 gnd 0.299809f
C5193 a_n2408_n452.n117 gnd 0.306874f
C5194 a_n2408_n452.n118 gnd 0.859759f
C5195 a_n2408_n452.t12 gnd 1.39989f
C5196 a_n2408_n452.t26 gnd 1.40268f
C5197 a_n2408_n452.t10 gnd 0.149803f
C5198 a_n2408_n452.t16 gnd 0.149803f
C5199 a_n2408_n452.n119 gnd 1.05521f
C5200 a_n2408_n452.t30 gnd 0.149803f
C5201 a_n2408_n452.t14 gnd 0.149803f
C5202 a_n2408_n452.n120 gnd 1.05521f
C5203 a_n2408_n452.n121 gnd 1.05522f
C5204 a_n2408_n452.t8 gnd 0.149803f
.ends

