* NGSPICE file created from opamp80.ext - technology: sky130A

.subckt opamp80 gnd CSoutput output vdd plus minus commonsourceibias outputibias diffpairibias
X0 CSoutput.t180 a_n8300_8799.t32 vdd.t293 vdd.t237 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X1 a_n2140_13878.t15 a_n2318_13878.t25 a_n2318_13878.t26 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X2 CSoutput.t183 commonsourceibias.t64 gnd.t228 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X3 a_n2140_13878.t23 a_n2318_13878.t48 vdd.t15 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 CSoutput.t216 a_n2318_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X5 vdd.t292 a_n8300_8799.t33 CSoutput.t179 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X6 gnd.t227 commonsourceibias.t65 CSoutput.t184 gnd.t150 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 a_n8300_8799.t28 plus.t5 a_n2903_n3924.t23 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X8 CSoutput.t35 commonsourceibias.t66 gnd.t226 gnd.t124 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X9 CSoutput.t36 commonsourceibias.t67 gnd.t225 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X10 CSoutput.t178 a_n8300_8799.t34 vdd.t291 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X11 CSoutput.t177 a_n8300_8799.t35 vdd.t290 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X12 minus.t4 gnd.t357 gnd.t359 gnd.t358 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X13 a_n2318_8322.t27 a_n2318_13878.t49 a_n8300_8799.t5 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X14 vdd.t28 CSoutput.t217 output.t16 gnd.t37 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X15 CSoutput.t176 a_n8300_8799.t36 vdd.t289 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X16 CSoutput.t29 commonsourceibias.t68 gnd.t224 gnd.t102 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X17 gnd.t220 commonsourceibias.t69 CSoutput.t30 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X18 CSoutput.t185 commonsourceibias.t70 gnd.t223 gnd.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 gnd.t222 commonsourceibias.t71 CSoutput.t186 gnd.t99 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X20 vdd.t288 a_n8300_8799.t37 CSoutput.t175 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X21 CSoutput.t46 commonsourceibias.t72 gnd.t221 gnd.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X22 CSoutput.t47 commonsourceibias.t73 gnd.t219 gnd.t163 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X23 gnd.t218 commonsourceibias.t74 CSoutput.t206 gnd.t131 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X24 commonsourceibias.t27 commonsourceibias.t26 gnd.t217 gnd.t102 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X25 a_n2318_13878.t0 minus.t5 a_n2903_n3924.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X26 CSoutput.t207 commonsourceibias.t75 gnd.t193 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X27 a_n8300_8799.t14 plus.t6 a_n2903_n3924.t22 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X28 a_n8300_8799.t3 a_n2318_13878.t50 a_n2318_8322.t26 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X29 a_n2318_13878.t42 minus.t6 a_n2903_n3924.t32 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X30 vdd.t287 a_n8300_8799.t38 CSoutput.t174 vdd.t250 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X31 vdd.t286 a_n8300_8799.t39 CSoutput.t173 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X32 CSoutput.t172 a_n8300_8799.t40 vdd.t285 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X33 vdd.t284 a_n8300_8799.t41 CSoutput.t171 vdd.t247 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X34 a_n8300_8799.t24 a_n2318_13878.t51 a_n2318_8322.t25 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X35 CSoutput.t218 a_n2318_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X36 CSoutput.t187 commonsourceibias.t76 gnd.t216 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 gnd.t215 commonsourceibias.t77 CSoutput.t188 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X38 gnd.t356 gnd.t354 gnd.t355 gnd.t281 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X39 CSoutput.t189 commonsourceibias.t78 gnd.t214 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X40 CSoutput.t190 commonsourceibias.t79 gnd.t213 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X41 gnd.t353 gnd.t351 gnd.t352 gnd.t273 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X42 vdd.t129 vdd.t127 vdd.t128 vdd.t55 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X43 CSoutput.t48 commonsourceibias.t80 gnd.t212 gnd.t134 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X44 CSoutput.t170 a_n8300_8799.t42 vdd.t283 vdd.t237 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X45 a_n2903_n3924.t21 plus.t7 a_n8300_8799.t25 gnd.t5 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X46 CSoutput.t169 a_n8300_8799.t43 vdd.t282 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X47 a_n2903_n3924.t7 diffpairibias.t16 gnd.t9 gnd.t8 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X48 a_n2903_n3924.t34 minus.t7 a_n2318_13878.t44 gnd.t59 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X49 CSoutput.t168 a_n8300_8799.t44 vdd.t281 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X50 gnd.t211 commonsourceibias.t81 CSoutput.t49 gnd.t107 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X51 vdd.t280 a_n8300_8799.t45 CSoutput.t167 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X52 CSoutput.t56 commonsourceibias.t82 gnd.t210 gnd.t90 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X53 gnd.t209 commonsourceibias.t24 commonsourceibias.t25 gnd.t104 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X54 CSoutput.t57 commonsourceibias.t83 gnd.t208 gnd.t134 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X55 output.t0 outputibias.t8 gnd.t18 gnd.t17 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X56 CSoutput.t166 a_n8300_8799.t46 vdd.t279 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X57 gnd.t207 commonsourceibias.t84 CSoutput.t201 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X58 a_n2140_13878.t14 a_n2318_13878.t31 a_n2318_13878.t32 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X59 CSoutput.t202 commonsourceibias.t85 gnd.t206 gnd.t118 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X60 gnd.t205 commonsourceibias.t86 CSoutput.t50 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X61 vdd.t29 CSoutput.t219 output.t15 gnd.t36 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X62 a_n2318_13878.t30 a_n2318_13878.t29 a_n2140_13878.t13 vdd.t30 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X63 CSoutput.t51 commonsourceibias.t87 gnd.t204 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X64 gnd.t203 commonsourceibias.t88 CSoutput.t3 gnd.t150 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X65 gnd.t350 gnd.t348 plus.t4 gnd.t349 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X66 CSoutput.t165 a_n8300_8799.t47 vdd.t278 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X67 vdd.t126 vdd.t124 vdd.t125 vdd.t101 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X68 gnd.t202 commonsourceibias.t22 commonsourceibias.t23 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X69 CSoutput.t4 commonsourceibias.t89 gnd.t201 gnd.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X70 gnd.t347 gnd.t344 gnd.t346 gnd.t345 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X71 a_n2903_n3924.t20 plus.t8 a_n8300_8799.t1 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X72 vdd.t263 a_n8300_8799.t48 CSoutput.t164 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X73 gnd.t343 gnd.t341 gnd.t342 gnd.t281 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X74 CSoutput.t31 commonsourceibias.t90 gnd.t200 gnd.t118 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X75 diffpairibias.t15 diffpairibias.t14 gnd.t68 gnd.t67 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X76 CSoutput.t32 commonsourceibias.t91 gnd.t199 gnd.t90 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X77 CSoutput.t208 commonsourceibias.t92 gnd.t198 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X78 gnd.t197 commonsourceibias.t93 CSoutput.t209 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X79 a_n8300_8799.t13 a_n2318_13878.t52 a_n2318_8322.t24 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X80 gnd.t196 commonsourceibias.t94 CSoutput.t191 gnd.t113 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X81 CSoutput.t163 a_n8300_8799.t49 vdd.t277 vdd.t234 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X82 gnd.t195 commonsourceibias.t95 CSoutput.t192 gnd.t82 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X83 vdd.t276 a_n8300_8799.t50 CSoutput.t162 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X84 vdd.t275 a_n8300_8799.t51 CSoutput.t161 vdd.t247 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X85 CSoutput.t37 commonsourceibias.t96 gnd.t194 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X86 diffpairibias.t13 diffpairibias.t12 gnd.t56 gnd.t55 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X87 CSoutput.t160 a_n8300_8799.t52 vdd.t274 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X88 gnd.t192 commonsourceibias.t38 commonsourceibias.t39 gnd.t116 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 gnd.t191 commonsourceibias.t97 CSoutput.t193 gnd.t131 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X90 CSoutput.t54 commonsourceibias.t98 gnd.t190 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 gnd.t189 commonsourceibias.t99 CSoutput.t38 gnd.t116 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X92 gnd.t340 gnd.t338 gnd.t339 gnd.t269 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X93 CSoutput.t24 commonsourceibias.t100 gnd.t188 gnd.t163 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 CSoutput.t210 commonsourceibias.t101 gnd.t187 gnd.t97 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X95 vdd.t273 a_n8300_8799.t53 CSoutput.t159 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X96 CSoutput.t158 a_n8300_8799.t54 vdd.t272 vdd.t256 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X97 gnd.t186 commonsourceibias.t102 CSoutput.t194 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X98 vdd.t123 vdd.t121 vdd.t122 vdd.t91 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X99 CSoutput.t157 a_n8300_8799.t55 vdd.t271 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X100 CSoutput.t156 a_n8300_8799.t56 vdd.t270 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X101 CSoutput.t155 a_n8300_8799.t57 vdd.t269 vdd.t256 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X102 CSoutput.t220 a_n2318_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X103 a_n2903_n3924.t33 minus.t8 a_n2318_13878.t43 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X104 gnd.t185 commonsourceibias.t50 commonsourceibias.t51 gnd.t94 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X105 a_n2903_n3924.t19 plus.t9 a_n8300_8799.t2 gnd.t6 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X106 output.t14 CSoutput.t221 vdd.t296 gnd.t35 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X107 gnd.t184 commonsourceibias.t103 CSoutput.t52 gnd.t116 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 a_n2903_n3924.t36 diffpairibias.t17 gnd.t66 gnd.t65 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X109 vdd.t262 a_n8300_8799.t58 CSoutput.t154 vdd.t226 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X110 gnd.t337 gnd.t335 gnd.t336 gnd.t265 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X111 vdd.t268 a_n8300_8799.t59 CSoutput.t153 vdd.t253 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X112 a_n2318_13878.t18 a_n2318_13878.t17 a_n2140_13878.t12 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X113 vdd.t267 a_n8300_8799.t60 CSoutput.t152 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X114 a_n2903_n3924.t18 plus.t10 a_n8300_8799.t12 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X115 vdd.t266 a_n8300_8799.t61 CSoutput.t151 vdd.t232 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X116 vdd.t265 a_n8300_8799.t62 CSoutput.t150 vdd.t250 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X117 gnd.t183 commonsourceibias.t104 CSoutput.t5 gnd.t107 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X118 a_n8300_8799.t18 a_n2318_13878.t53 a_n2318_8322.t23 vdd.t36 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X119 a_n2318_13878.t16 a_n2318_13878.t15 a_n2140_13878.t11 vdd.t53 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X120 gnd.t334 gnd.t332 gnd.t333 gnd.t265 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X121 CSoutput.t195 commonsourceibias.t105 gnd.t182 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X122 vdd.t264 a_n8300_8799.t63 CSoutput.t149 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X123 CSoutput.t148 a_n8300_8799.t64 vdd.t261 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X124 gnd.t181 commonsourceibias.t106 CSoutput.t39 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X125 vdd.t120 vdd.t118 vdd.t119 vdd.t67 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X126 output.t13 CSoutput.t222 vdd.t297 gnd.t34 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X127 vdd.t117 vdd.t115 vdd.t116 vdd.t105 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X128 gnd.t180 commonsourceibias.t54 commonsourceibias.t55 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X129 gnd.t179 commonsourceibias.t107 CSoutput.t211 gnd.t104 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X130 CSoutput.t147 a_n8300_8799.t65 vdd.t260 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X131 vdd.t114 vdd.t111 vdd.t113 vdd.t112 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X132 output.t18 outputibias.t9 gnd.t64 gnd.t63 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X133 CSoutput.t146 a_n8300_8799.t66 vdd.t259 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X134 CSoutput.t223 a_n2318_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X135 vdd.t258 a_n8300_8799.t67 CSoutput.t145 vdd.t253 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X136 vdd.t299 a_n2318_13878.t54 a_n2318_8322.t11 vdd.t298 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X137 a_n2318_13878.t14 a_n2318_13878.t13 a_n2140_13878.t10 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X138 gnd.t331 gnd.t329 minus.t3 gnd.t330 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X139 vdd.t110 vdd.t108 vdd.t109 vdd.t91 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X140 a_n2318_8322.t10 a_n2318_13878.t55 vdd.t50 vdd.t49 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X141 gnd.t178 commonsourceibias.t108 CSoutput.t196 gnd.t131 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X142 a_n2903_n3924.t37 diffpairibias.t18 gnd.t230 gnd.t229 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X143 output.t12 CSoutput.t224 vdd.t32 gnd.t33 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X144 CSoutput.t144 a_n8300_8799.t68 vdd.t257 vdd.t256 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X145 CSoutput.t143 a_n8300_8799.t69 vdd.t255 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X146 vdd.t33 CSoutput.t225 output.t11 gnd.t32 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X147 gnd.t177 commonsourceibias.t109 CSoutput.t58 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X148 gnd.t176 commonsourceibias.t52 commonsourceibias.t53 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X149 CSoutput.t42 commonsourceibias.t110 gnd.t175 gnd.t163 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X150 gnd.t174 commonsourceibias.t111 CSoutput.t17 gnd.t94 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X151 CSoutput.t33 commonsourceibias.t112 gnd.t173 gnd.t71 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X152 CSoutput.t203 commonsourceibias.t113 gnd.t172 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X153 CSoutput.t226 a_n2318_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X154 gnd.t328 gnd.t326 gnd.t327 gnd.t277 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X155 vdd.t27 a_n2318_13878.t56 a_n2140_13878.t22 vdd.t26 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X156 vdd.t107 vdd.t104 vdd.t106 vdd.t105 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X157 gnd.t325 gnd.t323 gnd.t324 gnd.t265 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X158 vdd.t254 a_n8300_8799.t70 CSoutput.t142 vdd.t253 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X159 vdd.t252 a_n8300_8799.t71 CSoutput.t141 vdd.t232 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X160 vdd.t251 a_n8300_8799.t72 CSoutput.t140 vdd.t250 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X161 a_n8300_8799.t27 plus.t11 a_n2903_n3924.t17 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X162 vdd.t103 vdd.t100 vdd.t102 vdd.t101 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X163 a_n2318_8322.t9 a_n2318_13878.t57 vdd.t6 vdd.t5 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X164 a_n8300_8799.t7 a_n2318_13878.t58 a_n2318_8322.t22 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X165 a_n8300_8799.t15 plus.t12 a_n2903_n3924.t16 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X166 CSoutput.t139 a_n8300_8799.t73 vdd.t249 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X167 diffpairibias.t11 diffpairibias.t10 gnd.t11 gnd.t10 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X168 vdd.t248 a_n8300_8799.t74 CSoutput.t138 vdd.t247 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X169 a_n2318_13878.t28 a_n2318_13878.t27 a_n2140_13878.t9 vdd.t3 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X170 vdd.t246 a_n8300_8799.t75 CSoutput.t137 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X171 CSoutput.t6 commonsourceibias.t114 gnd.t171 gnd.t124 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X172 a_n8300_8799.t0 a_n2318_13878.t59 a_n2318_8322.t21 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X173 CSoutput.t136 a_n8300_8799.t76 vdd.t245 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X174 commonsourceibias.t43 commonsourceibias.t42 gnd.t170 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X175 output.t10 CSoutput.t227 vdd.t34 gnd.t31 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X176 gnd.t169 commonsourceibias.t115 CSoutput.t7 gnd.t150 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X177 a_n2140_13878.t8 a_n2318_13878.t37 a_n2318_13878.t38 vdd.t36 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X178 gnd.t322 gnd.t320 gnd.t321 gnd.t241 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X179 vdd.t99 vdd.t97 vdd.t98 vdd.t67 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X180 gnd.t319 gnd.t316 gnd.t318 gnd.t317 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X181 CSoutput.t197 commonsourceibias.t116 gnd.t168 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X182 output.t9 CSoutput.t228 vdd.t39 gnd.t30 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X183 CSoutput.t135 a_n8300_8799.t77 vdd.t244 vdd.t234 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X184 CSoutput.t198 commonsourceibias.t117 gnd.t167 gnd.t118 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X185 gnd.t315 gnd.t313 gnd.t314 gnd.t273 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X186 vdd.t1 a_n2318_13878.t60 a_n2318_8322.t8 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X187 a_n2140_13878.t7 a_n2318_13878.t23 a_n2318_13878.t24 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X188 outputibias.t7 outputibias.t6 gnd.t51 gnd.t50 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X189 vdd.t243 a_n8300_8799.t78 CSoutput.t134 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X190 a_n2318_13878.t41 minus.t9 a_n2903_n3924.t30 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X191 a_n2903_n3924.t15 plus.t13 a_n8300_8799.t26 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X192 a_n2318_13878.t34 a_n2318_13878.t33 a_n2140_13878.t6 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X193 gnd.t166 commonsourceibias.t118 CSoutput.t40 gnd.t113 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X194 gnd.t165 commonsourceibias.t119 CSoutput.t214 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X195 commonsourceibias.t41 commonsourceibias.t40 gnd.t164 gnd.t163 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 gnd.t162 commonsourceibias.t120 CSoutput.t53 gnd.t99 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X197 outputibias.t5 outputibias.t4 gnd.t53 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X198 plus.t3 gnd.t310 gnd.t312 gnd.t311 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X199 vdd.t242 a_n8300_8799.t79 CSoutput.t133 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X200 CSoutput.t182 commonsourceibias.t121 gnd.t161 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X201 a_n2903_n3924.t28 diffpairibias.t19 gnd.t42 gnd.t41 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X202 gnd.t249 gnd.t247 minus.t2 gnd.t248 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X203 gnd.t309 gnd.t306 gnd.t308 gnd.t307 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X204 a_n2903_n3924.t29 diffpairibias.t20 gnd.t47 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X205 commonsourceibias.t49 commonsourceibias.t48 gnd.t160 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X206 a_n8300_8799.t6 plus.t14 a_n2903_n3924.t14 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X207 vdd.t241 a_n8300_8799.t80 CSoutput.t132 vdd.t226 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X208 vdd.t240 a_n8300_8799.t81 CSoutput.t131 vdd.t188 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X209 gnd.t305 gnd.t303 gnd.t304 gnd.t281 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X210 gnd.t302 gnd.t300 gnd.t301 gnd.t273 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X211 vdd.t40 CSoutput.t229 output.t8 gnd.t29 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X212 CSoutput.t34 commonsourceibias.t122 gnd.t158 gnd.t124 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X213 a_n8300_8799.t22 plus.t15 a_n2903_n3924.t13 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X214 CSoutput.t27 commonsourceibias.t123 gnd.t156 gnd.t97 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 CSoutput.t130 a_n8300_8799.t82 vdd.t239 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X216 CSoutput.t129 a_n8300_8799.t83 vdd.t238 vdd.t237 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X217 commonsourceibias.t47 commonsourceibias.t46 gnd.t157 gnd.t134 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X218 CSoutput.t128 a_n8300_8799.t84 vdd.t236 vdd.t218 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X219 gnd.t155 commonsourceibias.t44 commonsourceibias.t45 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X220 vdd.t41 CSoutput.t230 output.t7 gnd.t28 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X221 diffpairibias.t9 diffpairibias.t8 gnd.t13 gnd.t12 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X222 a_n2140_13878.t21 a_n2318_13878.t61 vdd.t17 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X223 a_n2318_13878.t3 minus.t10 a_n2903_n3924.t3 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X224 vdd.t52 a_n2318_13878.t62 a_n2140_13878.t20 vdd.t51 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X225 CSoutput.t9 commonsourceibias.t124 gnd.t153 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X226 CSoutput.t13 commonsourceibias.t125 gnd.t152 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X227 CSoutput.t127 a_n8300_8799.t85 vdd.t235 vdd.t234 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X228 gnd.t151 commonsourceibias.t10 commonsourceibias.t11 gnd.t150 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X229 a_n2903_n3924.t12 plus.t16 a_n8300_8799.t20 gnd.t59 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X230 vdd.t172 a_n8300_8799.t86 CSoutput.t126 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X231 vdd.t233 a_n8300_8799.t87 CSoutput.t125 vdd.t232 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X232 commonsourceibias.t9 commonsourceibias.t8 gnd.t149 gnd.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X233 outputibias.t3 outputibias.t2 gnd.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X234 CSoutput.t124 a_n8300_8799.t88 vdd.t231 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X235 a_n2140_13878.t5 a_n2318_13878.t19 a_n2318_13878.t20 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X236 gnd.t146 commonsourceibias.t126 CSoutput.t215 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X237 commonsourceibias.t7 commonsourceibias.t6 gnd.t147 gnd.t90 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X238 vdd.t230 a_n8300_8799.t89 CSoutput.t123 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X239 gnd.t145 commonsourceibias.t4 commonsourceibias.t5 gnd.t82 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X240 a_n2903_n3924.t39 minus.t11 a_n2318_13878.t47 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X241 a_n2318_8322.t20 a_n2318_13878.t63 a_n8300_8799.t30 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X242 CSoutput.t20 commonsourceibias.t127 gnd.t144 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X243 CSoutput.t122 a_n8300_8799.t90 vdd.t229 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X244 diffpairibias.t7 diffpairibias.t6 gnd.t49 gnd.t48 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X245 vdd.t174 a_n8300_8799.t91 CSoutput.t121 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X246 commonsourceibias.t21 commonsourceibias.t20 gnd.t143 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X247 vdd.t96 vdd.t94 vdd.t95 vdd.t77 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X248 vdd.t131 a_n2318_13878.t64 a_n2318_8322.t7 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X249 vdd.t228 a_n8300_8799.t92 CSoutput.t120 vdd.t188 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X250 vdd.t227 a_n8300_8799.t93 CSoutput.t119 vdd.t226 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X251 plus.t2 gnd.t297 gnd.t299 gnd.t298 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X252 gnd.t296 gnd.t294 minus.t1 gnd.t295 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X253 gnd.t142 commonsourceibias.t128 CSoutput.t204 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X254 CSoutput.t118 a_n8300_8799.t94 vdd.t225 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X255 gnd.t141 commonsourceibias.t18 commonsourceibias.t19 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X256 CSoutput.t59 commonsourceibias.t129 gnd.t139 gnd.t71 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X257 a_n2140_13878.t19 a_n2318_13878.t65 vdd.t38 vdd.t37 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X258 vdd.t93 vdd.t90 vdd.t92 vdd.t91 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X259 vdd.t89 vdd.t87 vdd.t88 vdd.t77 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X260 output.t6 CSoutput.t231 vdd.t42 gnd.t27 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X261 vdd.t224 a_n8300_8799.t95 CSoutput.t117 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X262 CSoutput.t116 a_n8300_8799.t96 vdd.t223 vdd.t218 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X263 CSoutput.t115 a_n8300_8799.t97 vdd.t222 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X264 CSoutput.t114 a_n8300_8799.t98 vdd.t221 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X265 gnd.t138 commonsourceibias.t130 CSoutput.t8 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X266 gnd.t293 gnd.t290 gnd.t292 gnd.t291 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X267 vdd.t220 a_n8300_8799.t99 CSoutput.t113 vdd.t144 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X268 a_n2903_n3924.t27 diffpairibias.t21 gnd.t39 gnd.t38 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X269 a_n2318_8322.t19 a_n2318_13878.t66 a_n8300_8799.t17 vdd.t3 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X270 vdd.t13 a_n2318_13878.t67 a_n2318_8322.t6 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X271 CSoutput.t112 a_n8300_8799.t100 vdd.t219 vdd.t218 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X272 gnd.t137 commonsourceibias.t16 commonsourceibias.t17 gnd.t107 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X273 a_n8300_8799.t29 plus.t17 a_n2903_n3924.t11 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X274 vdd.t217 a_n8300_8799.t101 CSoutput.t111 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X275 a_n2318_13878.t46 minus.t12 a_n2903_n3924.t38 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X276 CSoutput.t110 a_n8300_8799.t102 vdd.t216 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X277 a_n2903_n3924.t5 minus.t13 a_n2318_13878.t5 gnd.t6 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X278 vdd.t215 a_n8300_8799.t103 CSoutput.t109 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X279 vdd.t214 a_n8300_8799.t104 CSoutput.t108 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X280 vdd.t86 vdd.t84 vdd.t85 vdd.t63 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X281 output.t17 outputibias.t10 gnd.t58 gnd.t57 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X282 gnd.t289 gnd.t287 gnd.t288 gnd.t269 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X283 gnd.t136 commonsourceibias.t14 commonsourceibias.t15 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X284 vdd.t83 vdd.t80 vdd.t82 vdd.t81 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X285 gnd.t286 gnd.t284 gnd.t285 gnd.t269 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X286 CSoutput.t60 commonsourceibias.t131 gnd.t133 gnd.t102 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X287 a_n2903_n3924.t24 minus.t14 a_n2318_13878.t7 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X288 vdd.t213 a_n8300_8799.t105 CSoutput.t107 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X289 vdd.t43 CSoutput.t232 output.t5 gnd.t26 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X290 CSoutput.t106 a_n8300_8799.t106 vdd.t212 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X291 CSoutput.t26 commonsourceibias.t132 gnd.t135 gnd.t134 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X292 output.t19 outputibias.t11 gnd.t237 gnd.t236 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X293 a_n2903_n3924.t4 minus.t15 a_n2318_13878.t4 gnd.t5 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X294 a_n2140_13878.t4 a_n2318_13878.t39 a_n2318_13878.t40 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X295 CSoutput.t105 a_n8300_8799.t107 vdd.t210 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X296 a_n2318_8322.t18 a_n2318_13878.t68 a_n8300_8799.t21 vdd.t30 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X297 vdd.t79 vdd.t76 vdd.t78 vdd.t77 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X298 diffpairibias.t5 diffpairibias.t4 gnd.t232 gnd.t231 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X299 gnd.t283 gnd.t280 gnd.t282 gnd.t281 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X300 CSoutput.t104 a_n8300_8799.t108 vdd.t209 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X301 CSoutput.t103 a_n8300_8799.t109 vdd.t207 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X302 CSoutput.t102 a_n8300_8799.t110 vdd.t205 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X303 gnd.t132 commonsourceibias.t30 commonsourceibias.t31 gnd.t131 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X304 output.t4 CSoutput.t233 vdd.t44 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X305 vdd.t204 a_n8300_8799.t111 CSoutput.t101 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X306 CSoutput.t199 commonsourceibias.t133 gnd.t130 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 vdd.t203 a_n8300_8799.t112 CSoutput.t100 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X308 a_n2318_8322.t5 a_n2318_13878.t69 vdd.t133 vdd.t132 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X309 CSoutput.t99 a_n8300_8799.t113 vdd.t201 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X310 CSoutput.t98 a_n8300_8799.t114 vdd.t199 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X311 vdd.t75 vdd.t73 vdd.t74 vdd.t59 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X312 a_n2903_n3924.t35 minus.t16 a_n2318_13878.t45 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X313 vdd.t145 a_n8300_8799.t115 CSoutput.t97 vdd.t144 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X314 gnd.t128 commonsourceibias.t134 CSoutput.t200 gnd.t104 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X315 CSoutput.t96 a_n8300_8799.t116 vdd.t197 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X316 vdd.t25 a_n2318_13878.t70 a_n2140_13878.t18 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X317 vdd.t196 a_n8300_8799.t117 CSoutput.t95 vdd.t144 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X318 CSoutput.t94 a_n8300_8799.t118 vdd.t195 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X319 CSoutput.t93 a_n8300_8799.t119 vdd.t193 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X320 vdd.t176 a_n8300_8799.t120 CSoutput.t92 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X321 vdd.t192 a_n8300_8799.t121 CSoutput.t91 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X322 gnd.t279 gnd.t276 gnd.t278 gnd.t277 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X323 gnd.t127 commonsourceibias.t135 CSoutput.t43 gnd.t82 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X324 gnd.t246 gnd.t244 plus.t1 gnd.t245 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X325 gnd.t126 commonsourceibias.t136 CSoutput.t212 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X326 vdd.t72 vdd.t70 vdd.t71 vdd.t63 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X327 output.t3 CSoutput.t234 vdd.t45 gnd.t24 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X328 a_n2318_8322.t17 a_n2318_13878.t71 a_n8300_8799.t16 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X329 commonsourceibias.t29 commonsourceibias.t28 gnd.t125 gnd.t124 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 vdd.t46 CSoutput.t235 output.t2 gnd.t23 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X331 CSoutput.t90 a_n8300_8799.t122 vdd.t191 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X332 a_n8300_8799.t8 a_n2318_13878.t72 a_n2318_8322.t16 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X333 vdd.t189 a_n8300_8799.t123 CSoutput.t89 vdd.t188 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X334 a_n2140_13878.t17 a_n2318_13878.t73 vdd.t23 vdd.t22 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X335 gnd.t123 commonsourceibias.t137 CSoutput.t44 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X336 vdd.t187 a_n8300_8799.t124 CSoutput.t88 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X337 CSoutput.t87 a_n8300_8799.t125 vdd.t186 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X338 commonsourceibias.t3 commonsourceibias.t2 gnd.t122 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X339 a_n2903_n3924.t10 plus.t18 a_n8300_8799.t11 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X340 gnd.t275 gnd.t272 gnd.t274 gnd.t273 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X341 a_n2318_13878.t1 minus.t17 a_n2903_n3924.t1 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X342 gnd.t120 commonsourceibias.t138 CSoutput.t45 gnd.t113 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X343 a_n2318_8322.t15 a_n2318_13878.t74 a_n8300_8799.t10 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X344 commonsourceibias.t1 commonsourceibias.t0 gnd.t119 gnd.t118 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X345 gnd.t117 commonsourceibias.t139 CSoutput.t28 gnd.t116 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X346 CSoutput.t55 commonsourceibias.t140 gnd.t115 gnd.t71 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X347 vdd.t184 a_n8300_8799.t126 CSoutput.t86 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X348 gnd.t114 commonsourceibias.t36 commonsourceibias.t37 gnd.t113 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X349 CSoutput.t85 a_n8300_8799.t127 vdd.t182 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X350 CSoutput.t84 a_n8300_8799.t128 vdd.t180 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X351 CSoutput.t83 a_n8300_8799.t129 vdd.t179 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X352 gnd.t271 gnd.t268 gnd.t270 gnd.t269 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X353 a_n2140_13878.t3 a_n2318_13878.t11 a_n2318_13878.t12 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X354 vdd.t178 a_n8300_8799.t130 CSoutput.t82 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X355 gnd.t112 commonsourceibias.t34 commonsourceibias.t35 gnd.t99 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X356 vdd.t69 vdd.t66 vdd.t68 vdd.t67 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X357 vdd.t65 vdd.t62 vdd.t64 vdd.t63 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X358 commonsourceibias.t33 commonsourceibias.t32 gnd.t111 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X359 gnd.t109 commonsourceibias.t141 CSoutput.t181 gnd.t94 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X360 a_n2903_n3924.t26 minus.t18 a_n2318_13878.t8 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X361 a_n2903_n3924.t25 diffpairibias.t22 gnd.t20 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X362 gnd.t108 commonsourceibias.t142 CSoutput.t12 gnd.t107 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X363 vdd.t177 a_n8300_8799.t131 CSoutput.t81 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X364 CSoutput.t25 commonsourceibias.t143 gnd.t106 gnd.t97 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X365 vdd.t170 a_n8300_8799.t132 CSoutput.t80 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X366 gnd.t105 commonsourceibias.t144 CSoutput.t41 gnd.t104 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X367 CSoutput.t79 a_n8300_8799.t133 vdd.t169 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X368 CSoutput.t213 commonsourceibias.t145 gnd.t103 gnd.t102 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X369 a_n2318_13878.t10 a_n2318_13878.t9 a_n2140_13878.t2 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X370 gnd.t267 gnd.t264 gnd.t266 gnd.t265 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X371 a_n8300_8799.t4 a_n2318_13878.t75 a_n2318_8322.t14 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X372 vdd.t19 CSoutput.t236 output.t1 gnd.t22 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X373 vdd.t137 a_n8300_8799.t134 CSoutput.t78 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X374 CSoutput.t77 a_n8300_8799.t135 vdd.t168 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X375 vdd.t166 a_n8300_8799.t136 CSoutput.t76 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X376 CSoutput.t1 commonsourceibias.t146 gnd.t101 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X377 gnd.t100 commonsourceibias.t147 CSoutput.t10 gnd.t99 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X378 commonsourceibias.t57 commonsourceibias.t56 gnd.t98 gnd.t97 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X379 diffpairibias.t3 diffpairibias.t2 gnd.t44 gnd.t43 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X380 vdd.t165 a_n8300_8799.t137 CSoutput.t75 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X381 CSoutput.t74 a_n8300_8799.t138 vdd.t163 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X382 gnd.t263 gnd.t261 plus.t0 gnd.t262 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X383 CSoutput.t237 a_n2318_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X384 minus.t0 gnd.t258 gnd.t260 gnd.t259 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X385 CSoutput.t73 a_n8300_8799.t139 vdd.t162 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X386 a_n2318_8322.t13 a_n2318_13878.t76 a_n8300_8799.t9 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X387 gnd.t96 commonsourceibias.t148 CSoutput.t14 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X388 a_n2318_13878.t2 minus.t19 a_n2903_n3924.t2 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X389 vdd.t158 a_n8300_8799.t140 CSoutput.t72 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X390 gnd.t257 gnd.t254 gnd.t256 gnd.t255 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X391 CSoutput.t71 a_n8300_8799.t141 vdd.t160 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X392 diffpairibias.t1 diffpairibias.t0 gnd.t235 gnd.t234 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X393 gnd.t95 commonsourceibias.t149 CSoutput.t21 gnd.t94 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X394 commonsourceibias.t63 commonsourceibias.t62 gnd.t93 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X395 gnd.t92 commonsourceibias.t150 CSoutput.t0 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X396 CSoutput.t15 commonsourceibias.t151 gnd.t91 gnd.t90 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X397 vdd.t61 vdd.t58 vdd.t60 vdd.t59 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X398 vdd.t295 a_n2318_13878.t77 a_n2140_13878.t16 vdd.t294 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X399 CSoutput.t70 a_n8300_8799.t142 vdd.t156 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X400 vdd.t57 vdd.t54 vdd.t56 vdd.t55 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X401 vdd.t154 a_n8300_8799.t143 CSoutput.t69 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X402 vdd.t152 a_n8300_8799.t144 CSoutput.t68 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X403 gnd.t89 commonsourceibias.t60 commonsourceibias.t61 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X404 CSoutput.t67 a_n8300_8799.t145 vdd.t151 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X405 a_n8300_8799.t19 plus.t19 a_n2903_n3924.t9 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X406 gnd.t74 commonsourceibias.t152 CSoutput.t18 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X407 a_n2318_13878.t6 minus.t20 a_n2903_n3924.t6 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X408 commonsourceibias.t59 commonsourceibias.t58 gnd.t87 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X409 gnd.t85 commonsourceibias.t153 CSoutput.t22 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X410 gnd.t253 gnd.t250 gnd.t252 gnd.t251 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X411 gnd.t83 commonsourceibias.t154 CSoutput.t205 gnd.t82 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X412 a_n2318_8322.t12 a_n2318_13878.t78 a_n8300_8799.t23 vdd.t53 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X413 vdd.t149 a_n8300_8799.t146 CSoutput.t66 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X414 vdd.t147 a_n8300_8799.t147 CSoutput.t65 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X415 vdd.t143 a_n8300_8799.t148 CSoutput.t64 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X416 CSoutput.t63 a_n8300_8799.t149 vdd.t141 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X417 gnd.t81 commonsourceibias.t155 CSoutput.t2 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X418 a_n2318_8322.t4 a_n2318_13878.t79 vdd.t48 vdd.t47 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X419 gnd.t243 gnd.t240 gnd.t242 gnd.t241 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X420 gnd.t80 commonsourceibias.t156 CSoutput.t11 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X421 a_n2140_13878.t1 a_n2318_13878.t21 a_n2318_13878.t22 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X422 gnd.t78 commonsourceibias.t157 CSoutput.t16 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X423 CSoutput.t19 commonsourceibias.t158 gnd.t76 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X424 vdd.t139 a_n8300_8799.t150 CSoutput.t62 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X425 commonsourceibias.t13 commonsourceibias.t12 gnd.t72 gnd.t71 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X426 CSoutput.t23 commonsourceibias.t159 gnd.t70 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X427 outputibias.t1 outputibias.t0 gnd.t239 gnd.t238 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X428 a_n2903_n3924.t8 plus.t20 a_n8300_8799.t31 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X429 a_n2903_n3924.t31 diffpairibias.t23 gnd.t61 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X430 CSoutput.t61 a_n8300_8799.t151 vdd.t135 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X431 a_n2318_13878.t36 a_n2318_13878.t35 a_n2140_13878.t0 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 a_n8300_8799.n221 a_n8300_8799.t141 485.149
R1 a_n8300_8799.n240 a_n8300_8799.t34 485.149
R2 a_n8300_8799.n260 a_n8300_8799.t116 485.149
R3 a_n8300_8799.n160 a_n8300_8799.t99 485.149
R4 a_n8300_8799.n179 a_n8300_8799.t115 485.149
R5 a_n8300_8799.n199 a_n8300_8799.t117 485.149
R6 a_n8300_8799.n53 a_n8300_8799.t81 485.135
R7 a_n8300_8799.n233 a_n8300_8799.t57 464.166
R8 a_n8300_8799.n215 a_n8300_8799.t136 464.166
R9 a_n8300_8799.n232 a_n8300_8799.t98 464.166
R10 a_n8300_8799.n231 a_n8300_8799.t95 464.166
R11 a_n8300_8799.n216 a_n8300_8799.t35 464.166
R12 a_n8300_8799.n230 a_n8300_8799.t103 464.166
R13 a_n8300_8799.n229 a_n8300_8799.t102 464.166
R14 a_n8300_8799.n217 a_n8300_8799.t37 464.166
R15 a_n8300_8799.n228 a_n8300_8799.t36 464.166
R16 a_n8300_8799.n227 a_n8300_8799.t124 464.166
R17 a_n8300_8799.n218 a_n8300_8799.t52 464.166
R18 a_n8300_8799.n226 a_n8300_8799.t41 464.166
R19 a_n8300_8799.n225 a_n8300_8799.t128 464.166
R20 a_n8300_8799.n219 a_n8300_8799.t80 464.166
R21 a_n8300_8799.n224 a_n8300_8799.t56 464.166
R22 a_n8300_8799.n223 a_n8300_8799.t148 464.166
R23 a_n8300_8799.n220 a_n8300_8799.t97 464.166
R24 a_n8300_8799.n222 a_n8300_8799.t59 464.166
R25 a_n8300_8799.n68 a_n8300_8799.t92 485.135
R26 a_n8300_8799.n252 a_n8300_8799.t68 464.166
R27 a_n8300_8799.n234 a_n8300_8799.t150 464.166
R28 a_n8300_8799.n251 a_n8300_8799.t113 464.166
R29 a_n8300_8799.n250 a_n8300_8799.t112 464.166
R30 a_n8300_8799.n235 a_n8300_8799.t46 464.166
R31 a_n8300_8799.n249 a_n8300_8799.t120 464.166
R32 a_n8300_8799.n248 a_n8300_8799.t119 464.166
R33 a_n8300_8799.n236 a_n8300_8799.t48 464.166
R34 a_n8300_8799.n247 a_n8300_8799.t47 464.166
R35 a_n8300_8799.n246 a_n8300_8799.t140 464.166
R36 a_n8300_8799.n237 a_n8300_8799.t65 464.166
R37 a_n8300_8799.n245 a_n8300_8799.t51 464.166
R38 a_n8300_8799.n244 a_n8300_8799.t142 464.166
R39 a_n8300_8799.n238 a_n8300_8799.t93 464.166
R40 a_n8300_8799.n243 a_n8300_8799.t69 464.166
R41 a_n8300_8799.n242 a_n8300_8799.t39 464.166
R42 a_n8300_8799.n239 a_n8300_8799.t114 464.166
R43 a_n8300_8799.n241 a_n8300_8799.t70 464.166
R44 a_n8300_8799.n83 a_n8300_8799.t123 485.135
R45 a_n8300_8799.n272 a_n8300_8799.t54 464.166
R46 a_n8300_8799.n254 a_n8300_8799.t101 464.166
R47 a_n8300_8799.n271 a_n8300_8799.t40 464.166
R48 a_n8300_8799.n270 a_n8300_8799.t60 464.166
R49 a_n8300_8799.n255 a_n8300_8799.t145 464.166
R50 a_n8300_8799.n269 a_n8300_8799.t111 464.166
R51 a_n8300_8799.n268 a_n8300_8799.t139 464.166
R52 a_n8300_8799.n256 a_n8300_8799.t91 464.166
R53 a_n8300_8799.n267 a_n8300_8799.t118 464.166
R54 a_n8300_8799.n266 a_n8300_8799.t50 464.166
R55 a_n8300_8799.n257 a_n8300_8799.t135 464.166
R56 a_n8300_8799.n265 a_n8300_8799.t74 464.166
R57 a_n8300_8799.n264 a_n8300_8799.t129 464.166
R58 a_n8300_8799.n258 a_n8300_8799.t58 464.166
R59 a_n8300_8799.n263 a_n8300_8799.t106 464.166
R60 a_n8300_8799.n262 a_n8300_8799.t45 464.166
R61 a_n8300_8799.n259 a_n8300_8799.t88 464.166
R62 a_n8300_8799.n261 a_n8300_8799.t67 464.166
R63 a_n8300_8799.n161 a_n8300_8799.t138 464.166
R64 a_n8300_8799.n162 a_n8300_8799.t61 464.166
R65 a_n8300_8799.n163 a_n8300_8799.t94 464.166
R66 a_n8300_8799.n164 a_n8300_8799.t132 464.166
R67 a_n8300_8799.n159 a_n8300_8799.t133 464.166
R68 a_n8300_8799.n165 a_n8300_8799.t79 464.166
R69 a_n8300_8799.n166 a_n8300_8799.t110 464.166
R70 a_n8300_8799.n167 a_n8300_8799.t130 464.166
R71 a_n8300_8799.n168 a_n8300_8799.t77 464.166
R72 a_n8300_8799.n158 a_n8300_8799.t78 464.166
R73 a_n8300_8799.n169 a_n8300_8799.t107 464.166
R74 a_n8300_8799.n157 a_n8300_8799.t63 464.166
R75 a_n8300_8799.n170 a_n8300_8799.t64 464.166
R76 a_n8300_8799.n171 a_n8300_8799.t104 464.166
R77 a_n8300_8799.n172 a_n8300_8799.t32 464.166
R78 a_n8300_8799.n173 a_n8300_8799.t62 464.166
R79 a_n8300_8799.n156 a_n8300_8799.t84 464.166
R80 a_n8300_8799.n174 a_n8300_8799.t131 464.166
R81 a_n8300_8799.n180 a_n8300_8799.t151 464.166
R82 a_n8300_8799.n181 a_n8300_8799.t71 464.166
R83 a_n8300_8799.n182 a_n8300_8799.t108 464.166
R84 a_n8300_8799.n183 a_n8300_8799.t146 464.166
R85 a_n8300_8799.n178 a_n8300_8799.t149 464.166
R86 a_n8300_8799.n184 a_n8300_8799.t89 464.166
R87 a_n8300_8799.n185 a_n8300_8799.t127 464.166
R88 a_n8300_8799.n186 a_n8300_8799.t144 464.166
R89 a_n8300_8799.n187 a_n8300_8799.t85 464.166
R90 a_n8300_8799.n177 a_n8300_8799.t86 464.166
R91 a_n8300_8799.n188 a_n8300_8799.t125 464.166
R92 a_n8300_8799.n176 a_n8300_8799.t75 464.166
R93 a_n8300_8799.n189 a_n8300_8799.t76 464.166
R94 a_n8300_8799.n190 a_n8300_8799.t121 464.166
R95 a_n8300_8799.n191 a_n8300_8799.t42 464.166
R96 a_n8300_8799.n192 a_n8300_8799.t72 464.166
R97 a_n8300_8799.n175 a_n8300_8799.t96 464.166
R98 a_n8300_8799.n193 a_n8300_8799.t147 464.166
R99 a_n8300_8799.n200 a_n8300_8799.t66 464.166
R100 a_n8300_8799.n201 a_n8300_8799.t87 464.166
R101 a_n8300_8799.n202 a_n8300_8799.t44 464.166
R102 a_n8300_8799.n203 a_n8300_8799.t105 464.166
R103 a_n8300_8799.n198 a_n8300_8799.t82 464.166
R104 a_n8300_8799.n204 a_n8300_8799.t126 464.166
R105 a_n8300_8799.n205 a_n8300_8799.t73 464.166
R106 a_n8300_8799.n206 a_n8300_8799.t134 464.166
R107 a_n8300_8799.n207 a_n8300_8799.t49 464.166
R108 a_n8300_8799.n197 a_n8300_8799.t33 464.166
R109 a_n8300_8799.n208 a_n8300_8799.t90 464.166
R110 a_n8300_8799.n196 a_n8300_8799.t137 464.166
R111 a_n8300_8799.n209 a_n8300_8799.t109 464.166
R112 a_n8300_8799.n210 a_n8300_8799.t143 464.166
R113 a_n8300_8799.n211 a_n8300_8799.t83 464.166
R114 a_n8300_8799.n212 a_n8300_8799.t38 464.166
R115 a_n8300_8799.n195 a_n8300_8799.t100 464.166
R116 a_n8300_8799.n213 a_n8300_8799.t53 464.166
R117 a_n8300_8799.n44 a_n8300_8799.n67 71.7212
R118 a_n8300_8799.n67 a_n8300_8799.n220 17.8606
R119 a_n8300_8799.n66 a_n8300_8799.n44 76.9909
R120 a_n8300_8799.n223 a_n8300_8799.n66 7.32118
R121 a_n8300_8799.n65 a_n8300_8799.n43 78.3454
R122 a_n8300_8799.n43 a_n8300_8799.n64 72.8951
R123 a_n8300_8799.n63 a_n8300_8799.n45 70.1674
R124 a_n8300_8799.n226 a_n8300_8799.n63 20.9683
R125 a_n8300_8799.n45 a_n8300_8799.n62 72.3034
R126 a_n8300_8799.n62 a_n8300_8799.n218 16.6962
R127 a_n8300_8799.n61 a_n8300_8799.n46 77.6622
R128 a_n8300_8799.n227 a_n8300_8799.n61 5.97853
R129 a_n8300_8799.n60 a_n8300_8799.n46 77.6622
R130 a_n8300_8799.n47 a_n8300_8799.n59 72.3034
R131 a_n8300_8799.n58 a_n8300_8799.n47 70.1674
R132 a_n8300_8799.n230 a_n8300_8799.n58 20.9683
R133 a_n8300_8799.n49 a_n8300_8799.n57 72.8951
R134 a_n8300_8799.n57 a_n8300_8799.n216 15.5127
R135 a_n8300_8799.n56 a_n8300_8799.n49 78.3454
R136 a_n8300_8799.n231 a_n8300_8799.n56 4.61226
R137 a_n8300_8799.n55 a_n8300_8799.n48 76.9909
R138 a_n8300_8799.n48 a_n8300_8799.n54 71.7212
R139 a_n8300_8799.n233 a_n8300_8799.n53 20.9683
R140 a_n8300_8799.n50 a_n8300_8799.n53 70.1674
R141 a_n8300_8799.n36 a_n8300_8799.n82 71.7212
R142 a_n8300_8799.n82 a_n8300_8799.n239 17.8606
R143 a_n8300_8799.n81 a_n8300_8799.n36 76.9909
R144 a_n8300_8799.n242 a_n8300_8799.n81 7.32118
R145 a_n8300_8799.n80 a_n8300_8799.n35 78.3454
R146 a_n8300_8799.n35 a_n8300_8799.n79 72.8951
R147 a_n8300_8799.n78 a_n8300_8799.n37 70.1674
R148 a_n8300_8799.n245 a_n8300_8799.n78 20.9683
R149 a_n8300_8799.n37 a_n8300_8799.n77 72.3034
R150 a_n8300_8799.n77 a_n8300_8799.n237 16.6962
R151 a_n8300_8799.n76 a_n8300_8799.n38 77.6622
R152 a_n8300_8799.n246 a_n8300_8799.n76 5.97853
R153 a_n8300_8799.n75 a_n8300_8799.n38 77.6622
R154 a_n8300_8799.n39 a_n8300_8799.n74 72.3034
R155 a_n8300_8799.n73 a_n8300_8799.n39 70.1674
R156 a_n8300_8799.n249 a_n8300_8799.n73 20.9683
R157 a_n8300_8799.n41 a_n8300_8799.n72 72.8951
R158 a_n8300_8799.n72 a_n8300_8799.n235 15.5127
R159 a_n8300_8799.n71 a_n8300_8799.n41 78.3454
R160 a_n8300_8799.n250 a_n8300_8799.n71 4.61226
R161 a_n8300_8799.n70 a_n8300_8799.n40 76.9909
R162 a_n8300_8799.n40 a_n8300_8799.n69 71.7212
R163 a_n8300_8799.n252 a_n8300_8799.n68 20.9683
R164 a_n8300_8799.n42 a_n8300_8799.n68 70.1674
R165 a_n8300_8799.n28 a_n8300_8799.n97 71.7212
R166 a_n8300_8799.n97 a_n8300_8799.n259 17.8606
R167 a_n8300_8799.n96 a_n8300_8799.n28 76.9909
R168 a_n8300_8799.n262 a_n8300_8799.n96 7.32118
R169 a_n8300_8799.n95 a_n8300_8799.n27 78.3454
R170 a_n8300_8799.n27 a_n8300_8799.n94 72.8951
R171 a_n8300_8799.n93 a_n8300_8799.n29 70.1674
R172 a_n8300_8799.n265 a_n8300_8799.n93 20.9683
R173 a_n8300_8799.n29 a_n8300_8799.n92 72.3034
R174 a_n8300_8799.n92 a_n8300_8799.n257 16.6962
R175 a_n8300_8799.n91 a_n8300_8799.n30 77.6622
R176 a_n8300_8799.n266 a_n8300_8799.n91 5.97853
R177 a_n8300_8799.n90 a_n8300_8799.n30 77.6622
R178 a_n8300_8799.n31 a_n8300_8799.n89 72.3034
R179 a_n8300_8799.n88 a_n8300_8799.n31 70.1674
R180 a_n8300_8799.n269 a_n8300_8799.n88 20.9683
R181 a_n8300_8799.n33 a_n8300_8799.n87 72.8951
R182 a_n8300_8799.n87 a_n8300_8799.n255 15.5127
R183 a_n8300_8799.n86 a_n8300_8799.n33 78.3454
R184 a_n8300_8799.n270 a_n8300_8799.n86 4.61226
R185 a_n8300_8799.n85 a_n8300_8799.n32 76.9909
R186 a_n8300_8799.n32 a_n8300_8799.n84 71.7212
R187 a_n8300_8799.n272 a_n8300_8799.n83 20.9683
R188 a_n8300_8799.n34 a_n8300_8799.n83 70.1674
R189 a_n8300_8799.n20 a_n8300_8799.n112 70.1674
R190 a_n8300_8799.n174 a_n8300_8799.n112 20.9683
R191 a_n8300_8799.n111 a_n8300_8799.n20 71.7212
R192 a_n8300_8799.n111 a_n8300_8799.n156 17.8606
R193 a_n8300_8799.n19 a_n8300_8799.n110 76.9909
R194 a_n8300_8799.n173 a_n8300_8799.n110 7.32118
R195 a_n8300_8799.n109 a_n8300_8799.n19 78.3454
R196 a_n8300_8799.n21 a_n8300_8799.n108 72.8951
R197 a_n8300_8799.n107 a_n8300_8799.n21 70.1674
R198 a_n8300_8799.n107 a_n8300_8799.n157 20.9683
R199 a_n8300_8799.n22 a_n8300_8799.n106 72.3034
R200 a_n8300_8799.n169 a_n8300_8799.n106 16.6962
R201 a_n8300_8799.n105 a_n8300_8799.n22 77.6622
R202 a_n8300_8799.n105 a_n8300_8799.n158 5.97853
R203 a_n8300_8799.n23 a_n8300_8799.n104 77.6622
R204 a_n8300_8799.n103 a_n8300_8799.n23 72.3034
R205 a_n8300_8799.n24 a_n8300_8799.n102 70.1674
R206 a_n8300_8799.n165 a_n8300_8799.n102 20.9683
R207 a_n8300_8799.n101 a_n8300_8799.n24 72.8951
R208 a_n8300_8799.n101 a_n8300_8799.n159 15.5127
R209 a_n8300_8799.n25 a_n8300_8799.n100 78.3454
R210 a_n8300_8799.n164 a_n8300_8799.n100 4.61226
R211 a_n8300_8799.n99 a_n8300_8799.n25 76.9909
R212 a_n8300_8799.n98 a_n8300_8799.n162 17.8606
R213 a_n8300_8799.n98 a_n8300_8799.n26 71.7212
R214 a_n8300_8799.n12 a_n8300_8799.n127 70.1674
R215 a_n8300_8799.n193 a_n8300_8799.n127 20.9683
R216 a_n8300_8799.n126 a_n8300_8799.n12 71.7212
R217 a_n8300_8799.n126 a_n8300_8799.n175 17.8606
R218 a_n8300_8799.n11 a_n8300_8799.n125 76.9909
R219 a_n8300_8799.n192 a_n8300_8799.n125 7.32118
R220 a_n8300_8799.n124 a_n8300_8799.n11 78.3454
R221 a_n8300_8799.n13 a_n8300_8799.n123 72.8951
R222 a_n8300_8799.n122 a_n8300_8799.n13 70.1674
R223 a_n8300_8799.n122 a_n8300_8799.n176 20.9683
R224 a_n8300_8799.n14 a_n8300_8799.n121 72.3034
R225 a_n8300_8799.n188 a_n8300_8799.n121 16.6962
R226 a_n8300_8799.n120 a_n8300_8799.n14 77.6622
R227 a_n8300_8799.n120 a_n8300_8799.n177 5.97853
R228 a_n8300_8799.n15 a_n8300_8799.n119 77.6622
R229 a_n8300_8799.n118 a_n8300_8799.n15 72.3034
R230 a_n8300_8799.n16 a_n8300_8799.n117 70.1674
R231 a_n8300_8799.n184 a_n8300_8799.n117 20.9683
R232 a_n8300_8799.n116 a_n8300_8799.n16 72.8951
R233 a_n8300_8799.n116 a_n8300_8799.n178 15.5127
R234 a_n8300_8799.n17 a_n8300_8799.n115 78.3454
R235 a_n8300_8799.n183 a_n8300_8799.n115 4.61226
R236 a_n8300_8799.n114 a_n8300_8799.n17 76.9909
R237 a_n8300_8799.n113 a_n8300_8799.n181 17.8606
R238 a_n8300_8799.n113 a_n8300_8799.n18 71.7212
R239 a_n8300_8799.n4 a_n8300_8799.n142 70.1674
R240 a_n8300_8799.n213 a_n8300_8799.n142 20.9683
R241 a_n8300_8799.n141 a_n8300_8799.n4 71.7212
R242 a_n8300_8799.n141 a_n8300_8799.n195 17.8606
R243 a_n8300_8799.n3 a_n8300_8799.n140 76.9909
R244 a_n8300_8799.n212 a_n8300_8799.n140 7.32118
R245 a_n8300_8799.n139 a_n8300_8799.n3 78.3454
R246 a_n8300_8799.n5 a_n8300_8799.n138 72.8951
R247 a_n8300_8799.n137 a_n8300_8799.n5 70.1674
R248 a_n8300_8799.n137 a_n8300_8799.n196 20.9683
R249 a_n8300_8799.n6 a_n8300_8799.n136 72.3034
R250 a_n8300_8799.n208 a_n8300_8799.n136 16.6962
R251 a_n8300_8799.n135 a_n8300_8799.n6 77.6622
R252 a_n8300_8799.n135 a_n8300_8799.n197 5.97853
R253 a_n8300_8799.n7 a_n8300_8799.n134 77.6622
R254 a_n8300_8799.n133 a_n8300_8799.n7 72.3034
R255 a_n8300_8799.n8 a_n8300_8799.n132 70.1674
R256 a_n8300_8799.n204 a_n8300_8799.n132 20.9683
R257 a_n8300_8799.n131 a_n8300_8799.n8 72.8951
R258 a_n8300_8799.n131 a_n8300_8799.n198 15.5127
R259 a_n8300_8799.n9 a_n8300_8799.n130 78.3454
R260 a_n8300_8799.n203 a_n8300_8799.n130 4.61226
R261 a_n8300_8799.n129 a_n8300_8799.n9 76.9909
R262 a_n8300_8799.n128 a_n8300_8799.n201 17.8606
R263 a_n8300_8799.n128 a_n8300_8799.n10 71.7212
R264 a_n8300_8799.n281 a_n8300_8799.n280 98.9632
R265 a_n8300_8799.n51 a_n8300_8799.n143 98.9631
R266 a_n8300_8799.n52 a_n8300_8799.n277 98.6055
R267 a_n8300_8799.n52 a_n8300_8799.n278 98.6055
R268 a_n8300_8799.n280 a_n8300_8799.n279 98.6055
R269 a_n8300_8799.n51 a_n8300_8799.n144 98.6055
R270 a_n8300_8799.n51 a_n8300_8799.n145 98.6055
R271 a_n8300_8799.n147 a_n8300_8799.n146 98.6055
R272 a_n8300_8799.n1 a_n8300_8799.n148 81.4626
R273 a_n8300_8799.n2 a_n8300_8799.n152 81.4626
R274 a_n8300_8799.n2 a_n8300_8799.n150 81.4626
R275 a_n8300_8799.n0 a_n8300_8799.n154 80.9324
R276 a_n8300_8799.n1 a_n8300_8799.n155 80.9324
R277 a_n8300_8799.n1 a_n8300_8799.n149 80.9324
R278 a_n8300_8799.n2 a_n8300_8799.n153 80.9324
R279 a_n8300_8799.n2 a_n8300_8799.n151 80.9324
R280 a_n8300_8799.n44 a_n8300_8799.n221 70.4033
R281 a_n8300_8799.n36 a_n8300_8799.n240 70.4033
R282 a_n8300_8799.n28 a_n8300_8799.n260 70.4033
R283 a_n8300_8799.n160 a_n8300_8799.n26 70.4033
R284 a_n8300_8799.n179 a_n8300_8799.n18 70.4033
R285 a_n8300_8799.n199 a_n8300_8799.n10 70.4033
R286 a_n8300_8799.n232 a_n8300_8799.n231 48.2005
R287 a_n8300_8799.n58 a_n8300_8799.n229 20.9683
R288 a_n8300_8799.n228 a_n8300_8799.n227 48.2005
R289 a_n8300_8799.n63 a_n8300_8799.n225 20.9683
R290 a_n8300_8799.n224 a_n8300_8799.n223 48.2005
R291 a_n8300_8799.n251 a_n8300_8799.n250 48.2005
R292 a_n8300_8799.n73 a_n8300_8799.n248 20.9683
R293 a_n8300_8799.n247 a_n8300_8799.n246 48.2005
R294 a_n8300_8799.n78 a_n8300_8799.n244 20.9683
R295 a_n8300_8799.n243 a_n8300_8799.n242 48.2005
R296 a_n8300_8799.n271 a_n8300_8799.n270 48.2005
R297 a_n8300_8799.n88 a_n8300_8799.n268 20.9683
R298 a_n8300_8799.n267 a_n8300_8799.n266 48.2005
R299 a_n8300_8799.n93 a_n8300_8799.n264 20.9683
R300 a_n8300_8799.n263 a_n8300_8799.n262 48.2005
R301 a_n8300_8799.n164 a_n8300_8799.n163 48.2005
R302 a_n8300_8799.n166 a_n8300_8799.n102 20.9683
R303 a_n8300_8799.n168 a_n8300_8799.n158 48.2005
R304 a_n8300_8799.n170 a_n8300_8799.n107 20.9683
R305 a_n8300_8799.n173 a_n8300_8799.n172 48.2005
R306 a_n8300_8799.t43 a_n8300_8799.n112 485.135
R307 a_n8300_8799.n183 a_n8300_8799.n182 48.2005
R308 a_n8300_8799.n185 a_n8300_8799.n117 20.9683
R309 a_n8300_8799.n187 a_n8300_8799.n177 48.2005
R310 a_n8300_8799.n189 a_n8300_8799.n122 20.9683
R311 a_n8300_8799.n192 a_n8300_8799.n191 48.2005
R312 a_n8300_8799.t55 a_n8300_8799.n127 485.135
R313 a_n8300_8799.n203 a_n8300_8799.n202 48.2005
R314 a_n8300_8799.n205 a_n8300_8799.n132 20.9683
R315 a_n8300_8799.n207 a_n8300_8799.n197 48.2005
R316 a_n8300_8799.n209 a_n8300_8799.n137 20.9683
R317 a_n8300_8799.n212 a_n8300_8799.n211 48.2005
R318 a_n8300_8799.t122 a_n8300_8799.n142 485.135
R319 a_n8300_8799.n54 a_n8300_8799.n215 17.8606
R320 a_n8300_8799.n222 a_n8300_8799.n67 25.894
R321 a_n8300_8799.n69 a_n8300_8799.n234 17.8606
R322 a_n8300_8799.n241 a_n8300_8799.n82 25.894
R323 a_n8300_8799.n84 a_n8300_8799.n254 17.8606
R324 a_n8300_8799.n261 a_n8300_8799.n97 25.894
R325 a_n8300_8799.n174 a_n8300_8799.n111 25.894
R326 a_n8300_8799.n193 a_n8300_8799.n126 25.894
R327 a_n8300_8799.n213 a_n8300_8799.n141 25.894
R328 a_n8300_8799.n65 a_n8300_8799.n219 43.3183
R329 a_n8300_8799.n80 a_n8300_8799.n238 43.3183
R330 a_n8300_8799.n95 a_n8300_8799.n258 43.3183
R331 a_n8300_8799.n171 a_n8300_8799.n109 43.3183
R332 a_n8300_8799.n190 a_n8300_8799.n124 43.3183
R333 a_n8300_8799.n210 a_n8300_8799.n139 43.3183
R334 a_n8300_8799.n59 a_n8300_8799.n217 16.6962
R335 a_n8300_8799.n226 a_n8300_8799.n62 27.6507
R336 a_n8300_8799.n74 a_n8300_8799.n236 16.6962
R337 a_n8300_8799.n245 a_n8300_8799.n77 27.6507
R338 a_n8300_8799.n89 a_n8300_8799.n256 16.6962
R339 a_n8300_8799.n265 a_n8300_8799.n92 27.6507
R340 a_n8300_8799.n167 a_n8300_8799.n103 16.6962
R341 a_n8300_8799.n157 a_n8300_8799.n106 27.6507
R342 a_n8300_8799.n186 a_n8300_8799.n118 16.6962
R343 a_n8300_8799.n176 a_n8300_8799.n121 27.6507
R344 a_n8300_8799.n206 a_n8300_8799.n133 16.6962
R345 a_n8300_8799.n196 a_n8300_8799.n136 27.6507
R346 a_n8300_8799.n60 a_n8300_8799.n217 41.7634
R347 a_n8300_8799.n75 a_n8300_8799.n236 41.7634
R348 a_n8300_8799.n90 a_n8300_8799.n256 41.7634
R349 a_n8300_8799.n104 a_n8300_8799.n167 41.7634
R350 a_n8300_8799.n119 a_n8300_8799.n186 41.7634
R351 a_n8300_8799.n134 a_n8300_8799.n206 41.7634
R352 a_n8300_8799.n230 a_n8300_8799.n57 29.3885
R353 a_n8300_8799.n64 a_n8300_8799.n219 15.5127
R354 a_n8300_8799.n249 a_n8300_8799.n72 29.3885
R355 a_n8300_8799.n79 a_n8300_8799.n238 15.5127
R356 a_n8300_8799.n269 a_n8300_8799.n87 29.3885
R357 a_n8300_8799.n94 a_n8300_8799.n258 15.5127
R358 a_n8300_8799.n165 a_n8300_8799.n101 29.3885
R359 a_n8300_8799.n171 a_n8300_8799.n108 15.5127
R360 a_n8300_8799.n184 a_n8300_8799.n116 29.3885
R361 a_n8300_8799.n190 a_n8300_8799.n123 15.5127
R362 a_n8300_8799.n204 a_n8300_8799.n131 29.3885
R363 a_n8300_8799.n210 a_n8300_8799.n138 15.5127
R364 a_n8300_8799.n55 a_n8300_8799.n215 40.1848
R365 a_n8300_8799.n70 a_n8300_8799.n234 40.1848
R366 a_n8300_8799.n85 a_n8300_8799.n254 40.1848
R367 a_n8300_8799.n162 a_n8300_8799.n99 40.1848
R368 a_n8300_8799.n181 a_n8300_8799.n114 40.1848
R369 a_n8300_8799.n201 a_n8300_8799.n129 40.1848
R370 a_n8300_8799.n276 a_n8300_8799.n147 31.7372
R371 a_n8300_8799.n222 a_n8300_8799.n221 20.9576
R372 a_n8300_8799.n241 a_n8300_8799.n240 20.9576
R373 a_n8300_8799.n261 a_n8300_8799.n260 20.9576
R374 a_n8300_8799.n161 a_n8300_8799.n160 20.9576
R375 a_n8300_8799.n180 a_n8300_8799.n179 20.9576
R376 a_n8300_8799.n200 a_n8300_8799.n199 20.9576
R377 a_n8300_8799.n52 a_n8300_8799.n276 18.8589
R378 a_n8300_8799.n55 a_n8300_8799.n232 7.32118
R379 a_n8300_8799.n66 a_n8300_8799.n220 40.1848
R380 a_n8300_8799.n70 a_n8300_8799.n251 7.32118
R381 a_n8300_8799.n81 a_n8300_8799.n239 40.1848
R382 a_n8300_8799.n85 a_n8300_8799.n271 7.32118
R383 a_n8300_8799.n96 a_n8300_8799.n259 40.1848
R384 a_n8300_8799.n163 a_n8300_8799.n99 7.32118
R385 a_n8300_8799.n156 a_n8300_8799.n110 40.1848
R386 a_n8300_8799.n182 a_n8300_8799.n114 7.32118
R387 a_n8300_8799.n175 a_n8300_8799.n125 40.1848
R388 a_n8300_8799.n202 a_n8300_8799.n129 7.32118
R389 a_n8300_8799.n195 a_n8300_8799.n140 40.1848
R390 a_n8300_8799.n225 a_n8300_8799.n64 29.3885
R391 a_n8300_8799.n244 a_n8300_8799.n79 29.3885
R392 a_n8300_8799.n264 a_n8300_8799.n94 29.3885
R393 a_n8300_8799.n108 a_n8300_8799.n170 29.3885
R394 a_n8300_8799.n123 a_n8300_8799.n189 29.3885
R395 a_n8300_8799.n138 a_n8300_8799.n209 29.3885
R396 a_n8300_8799.n60 a_n8300_8799.n228 5.97853
R397 a_n8300_8799.n61 a_n8300_8799.n218 41.7634
R398 a_n8300_8799.n75 a_n8300_8799.n247 5.97853
R399 a_n8300_8799.n76 a_n8300_8799.n237 41.7634
R400 a_n8300_8799.n90 a_n8300_8799.n267 5.97853
R401 a_n8300_8799.n91 a_n8300_8799.n257 41.7634
R402 a_n8300_8799.n168 a_n8300_8799.n104 5.97853
R403 a_n8300_8799.n169 a_n8300_8799.n105 41.7634
R404 a_n8300_8799.n187 a_n8300_8799.n119 5.97853
R405 a_n8300_8799.n188 a_n8300_8799.n120 41.7634
R406 a_n8300_8799.n207 a_n8300_8799.n134 5.97853
R407 a_n8300_8799.n208 a_n8300_8799.n135 41.7634
R408 a_n8300_8799.n275 a_n8300_8799.n1 12.3339
R409 a_n8300_8799.n276 a_n8300_8799.n275 11.4887
R410 a_n8300_8799.n229 a_n8300_8799.n59 27.6507
R411 a_n8300_8799.n248 a_n8300_8799.n74 27.6507
R412 a_n8300_8799.n268 a_n8300_8799.n89 27.6507
R413 a_n8300_8799.n166 a_n8300_8799.n103 27.6507
R414 a_n8300_8799.n185 a_n8300_8799.n118 27.6507
R415 a_n8300_8799.n205 a_n8300_8799.n133 27.6507
R416 a_n8300_8799.n56 a_n8300_8799.n216 43.3183
R417 a_n8300_8799.n65 a_n8300_8799.n224 4.61226
R418 a_n8300_8799.n71 a_n8300_8799.n235 43.3183
R419 a_n8300_8799.n80 a_n8300_8799.n243 4.61226
R420 a_n8300_8799.n86 a_n8300_8799.n255 43.3183
R421 a_n8300_8799.n95 a_n8300_8799.n263 4.61226
R422 a_n8300_8799.n159 a_n8300_8799.n100 43.3183
R423 a_n8300_8799.n172 a_n8300_8799.n109 4.61226
R424 a_n8300_8799.n178 a_n8300_8799.n115 43.3183
R425 a_n8300_8799.n191 a_n8300_8799.n124 4.61226
R426 a_n8300_8799.n198 a_n8300_8799.n130 43.3183
R427 a_n8300_8799.n0 a_n8300_8799.n2 33.2634
R428 a_n8300_8799.n211 a_n8300_8799.n139 4.61226
R429 a_n8300_8799.n253 a_n8300_8799.n50 9.04406
R430 a_n8300_8799.n194 a_n8300_8799.n20 9.04406
R431 a_n8300_8799.n233 a_n8300_8799.n54 25.894
R432 a_n8300_8799.n252 a_n8300_8799.n69 25.894
R433 a_n8300_8799.n272 a_n8300_8799.n84 25.894
R434 a_n8300_8799.n98 a_n8300_8799.n161 25.894
R435 a_n8300_8799.n113 a_n8300_8799.n180 25.894
R436 a_n8300_8799.n128 a_n8300_8799.n200 25.894
R437 a_n8300_8799.n274 a_n8300_8799.n214 6.96667
R438 a_n8300_8799.n274 a_n8300_8799.n273 6.62419
R439 a_n8300_8799.n253 a_n8300_8799.n42 4.93611
R440 a_n8300_8799.n273 a_n8300_8799.n34 4.93611
R441 a_n8300_8799.n194 a_n8300_8799.n12 4.93611
R442 a_n8300_8799.n214 a_n8300_8799.n4 4.93611
R443 a_n8300_8799.n273 a_n8300_8799.n253 4.10845
R444 a_n8300_8799.n214 a_n8300_8799.n194 4.10845
R445 a_n8300_8799.n277 a_n8300_8799.t9 3.61217
R446 a_n8300_8799.n277 a_n8300_8799.t3 3.61217
R447 a_n8300_8799.n278 a_n8300_8799.t21 3.61217
R448 a_n8300_8799.n278 a_n8300_8799.t4 3.61217
R449 a_n8300_8799.n279 a_n8300_8799.t30 3.61217
R450 a_n8300_8799.n279 a_n8300_8799.t18 3.61217
R451 a_n8300_8799.n143 a_n8300_8799.t17 3.61217
R452 a_n8300_8799.n143 a_n8300_8799.t24 3.61217
R453 a_n8300_8799.n144 a_n8300_8799.t5 3.61217
R454 a_n8300_8799.n144 a_n8300_8799.t7 3.61217
R455 a_n8300_8799.n145 a_n8300_8799.t16 3.61217
R456 a_n8300_8799.n145 a_n8300_8799.t8 3.61217
R457 a_n8300_8799.n146 a_n8300_8799.t10 3.61217
R458 a_n8300_8799.n146 a_n8300_8799.t13 3.61217
R459 a_n8300_8799.n281 a_n8300_8799.t23 3.61217
R460 a_n8300_8799.t0 a_n8300_8799.n281 3.61217
R461 a_n8300_8799.n275 a_n8300_8799.n274 3.4105
R462 a_n8300_8799.n154 a_n8300_8799.t12 2.82907
R463 a_n8300_8799.n154 a_n8300_8799.t15 2.82907
R464 a_n8300_8799.n155 a_n8300_8799.t26 2.82907
R465 a_n8300_8799.n155 a_n8300_8799.t6 2.82907
R466 a_n8300_8799.n149 a_n8300_8799.t11 2.82907
R467 a_n8300_8799.n149 a_n8300_8799.t29 2.82907
R468 a_n8300_8799.n148 a_n8300_8799.t2 2.82907
R469 a_n8300_8799.n148 a_n8300_8799.t28 2.82907
R470 a_n8300_8799.n152 a_n8300_8799.t1 2.82907
R471 a_n8300_8799.n152 a_n8300_8799.t27 2.82907
R472 a_n8300_8799.n153 a_n8300_8799.t31 2.82907
R473 a_n8300_8799.n153 a_n8300_8799.t19 2.82907
R474 a_n8300_8799.n151 a_n8300_8799.t20 2.82907
R475 a_n8300_8799.n151 a_n8300_8799.t22 2.82907
R476 a_n8300_8799.n150 a_n8300_8799.t25 2.82907
R477 a_n8300_8799.n150 a_n8300_8799.t14 2.82907
R478 a_n8300_8799.n44 a_n8300_8799.n43 1.13686
R479 a_n8300_8799.n36 a_n8300_8799.n35 1.13686
R480 a_n8300_8799.n28 a_n8300_8799.n27 1.13686
R481 a_n8300_8799.n20 a_n8300_8799.n19 1.13686
R482 a_n8300_8799.n12 a_n8300_8799.n11 1.13686
R483 a_n8300_8799.n4 a_n8300_8799.n3 1.13686
R484 a_n8300_8799.n1 a_n8300_8799.n0 1.06084
R485 a_n8300_8799.n49 a_n8300_8799.n48 0.758076
R486 a_n8300_8799.n49 a_n8300_8799.n47 0.758076
R487 a_n8300_8799.n47 a_n8300_8799.n46 0.758076
R488 a_n8300_8799.n46 a_n8300_8799.n45 0.758076
R489 a_n8300_8799.n43 a_n8300_8799.n45 0.758076
R490 a_n8300_8799.n41 a_n8300_8799.n40 0.758076
R491 a_n8300_8799.n41 a_n8300_8799.n39 0.758076
R492 a_n8300_8799.n39 a_n8300_8799.n38 0.758076
R493 a_n8300_8799.n38 a_n8300_8799.n37 0.758076
R494 a_n8300_8799.n35 a_n8300_8799.n37 0.758076
R495 a_n8300_8799.n33 a_n8300_8799.n32 0.758076
R496 a_n8300_8799.n33 a_n8300_8799.n31 0.758076
R497 a_n8300_8799.n31 a_n8300_8799.n30 0.758076
R498 a_n8300_8799.n30 a_n8300_8799.n29 0.758076
R499 a_n8300_8799.n27 a_n8300_8799.n29 0.758076
R500 a_n8300_8799.n24 a_n8300_8799.n25 0.758076
R501 a_n8300_8799.n23 a_n8300_8799.n24 0.758076
R502 a_n8300_8799.n22 a_n8300_8799.n23 0.758076
R503 a_n8300_8799.n21 a_n8300_8799.n22 0.758076
R504 a_n8300_8799.n19 a_n8300_8799.n21 0.758076
R505 a_n8300_8799.n16 a_n8300_8799.n17 0.758076
R506 a_n8300_8799.n15 a_n8300_8799.n16 0.758076
R507 a_n8300_8799.n14 a_n8300_8799.n15 0.758076
R508 a_n8300_8799.n13 a_n8300_8799.n14 0.758076
R509 a_n8300_8799.n11 a_n8300_8799.n13 0.758076
R510 a_n8300_8799.n8 a_n8300_8799.n9 0.758076
R511 a_n8300_8799.n7 a_n8300_8799.n8 0.758076
R512 a_n8300_8799.n6 a_n8300_8799.n7 0.758076
R513 a_n8300_8799.n5 a_n8300_8799.n6 0.758076
R514 a_n8300_8799.n3 a_n8300_8799.n5 0.758076
R515 a_n8300_8799.n280 a_n8300_8799.n52 0.716017
R516 a_n8300_8799.n147 a_n8300_8799.n51 0.716017
R517 a_n8300_8799.n9 a_n8300_8799.n10 0.568682
R518 a_n8300_8799.n17 a_n8300_8799.n18 0.568682
R519 a_n8300_8799.n25 a_n8300_8799.n26 0.568682
R520 a_n8300_8799.n32 a_n8300_8799.n34 0.568682
R521 a_n8300_8799.n40 a_n8300_8799.n42 0.568682
R522 a_n8300_8799.n48 a_n8300_8799.n50 0.568682
R523 vdd.n327 vdd.n291 756.745
R524 vdd.n268 vdd.n232 756.745
R525 vdd.n225 vdd.n189 756.745
R526 vdd.n166 vdd.n130 756.745
R527 vdd.n124 vdd.n88 756.745
R528 vdd.n65 vdd.n29 756.745
R529 vdd.n2108 vdd.n2072 756.745
R530 vdd.n2167 vdd.n2131 756.745
R531 vdd.n2006 vdd.n1970 756.745
R532 vdd.n2065 vdd.n2029 756.745
R533 vdd.n1905 vdd.n1869 756.745
R534 vdd.n1964 vdd.n1928 756.745
R535 vdd.n1253 vdd.t58 640.208
R536 vdd.n981 vdd.t100 640.208
R537 vdd.n1273 vdd.t73 640.208
R538 vdd.n972 vdd.t124 640.208
R539 vdd.n872 vdd.t80 640.208
R540 vdd.n2704 vdd.t115 640.208
R541 vdd.n832 vdd.t127 640.208
R542 vdd.n2701 vdd.t104 640.208
R543 vdd.n799 vdd.t54 640.208
R544 vdd.n1043 vdd.t111 640.208
R545 vdd.n1679 vdd.t90 592.009
R546 vdd.n1717 vdd.t108 592.009
R547 vdd.n1613 vdd.t121 592.009
R548 vdd.n2269 vdd.t66 592.009
R549 vdd.n1190 vdd.t97 592.009
R550 vdd.n1150 vdd.t118 592.009
R551 vdd.n426 vdd.t87 592.009
R552 vdd.n440 vdd.t76 592.009
R553 vdd.n452 vdd.t94 592.009
R554 vdd.n768 vdd.t70 592.009
R555 vdd.n3276 vdd.t84 592.009
R556 vdd.n688 vdd.t62 592.009
R557 vdd.n328 vdd.n327 585
R558 vdd.n326 vdd.n293 585
R559 vdd.n325 vdd.n324 585
R560 vdd.n296 vdd.n294 585
R561 vdd.n319 vdd.n318 585
R562 vdd.n317 vdd.n316 585
R563 vdd.n300 vdd.n299 585
R564 vdd.n311 vdd.n310 585
R565 vdd.n309 vdd.n308 585
R566 vdd.n304 vdd.n303 585
R567 vdd.n269 vdd.n268 585
R568 vdd.n267 vdd.n234 585
R569 vdd.n266 vdd.n265 585
R570 vdd.n237 vdd.n235 585
R571 vdd.n260 vdd.n259 585
R572 vdd.n258 vdd.n257 585
R573 vdd.n241 vdd.n240 585
R574 vdd.n252 vdd.n251 585
R575 vdd.n250 vdd.n249 585
R576 vdd.n245 vdd.n244 585
R577 vdd.n226 vdd.n225 585
R578 vdd.n224 vdd.n191 585
R579 vdd.n223 vdd.n222 585
R580 vdd.n194 vdd.n192 585
R581 vdd.n217 vdd.n216 585
R582 vdd.n215 vdd.n214 585
R583 vdd.n198 vdd.n197 585
R584 vdd.n209 vdd.n208 585
R585 vdd.n207 vdd.n206 585
R586 vdd.n202 vdd.n201 585
R587 vdd.n167 vdd.n166 585
R588 vdd.n165 vdd.n132 585
R589 vdd.n164 vdd.n163 585
R590 vdd.n135 vdd.n133 585
R591 vdd.n158 vdd.n157 585
R592 vdd.n156 vdd.n155 585
R593 vdd.n139 vdd.n138 585
R594 vdd.n150 vdd.n149 585
R595 vdd.n148 vdd.n147 585
R596 vdd.n143 vdd.n142 585
R597 vdd.n125 vdd.n124 585
R598 vdd.n123 vdd.n90 585
R599 vdd.n122 vdd.n121 585
R600 vdd.n93 vdd.n91 585
R601 vdd.n116 vdd.n115 585
R602 vdd.n114 vdd.n113 585
R603 vdd.n97 vdd.n96 585
R604 vdd.n108 vdd.n107 585
R605 vdd.n106 vdd.n105 585
R606 vdd.n101 vdd.n100 585
R607 vdd.n66 vdd.n65 585
R608 vdd.n64 vdd.n31 585
R609 vdd.n63 vdd.n62 585
R610 vdd.n34 vdd.n32 585
R611 vdd.n57 vdd.n56 585
R612 vdd.n55 vdd.n54 585
R613 vdd.n38 vdd.n37 585
R614 vdd.n49 vdd.n48 585
R615 vdd.n47 vdd.n46 585
R616 vdd.n42 vdd.n41 585
R617 vdd.n2109 vdd.n2108 585
R618 vdd.n2107 vdd.n2074 585
R619 vdd.n2106 vdd.n2105 585
R620 vdd.n2077 vdd.n2075 585
R621 vdd.n2100 vdd.n2099 585
R622 vdd.n2098 vdd.n2097 585
R623 vdd.n2081 vdd.n2080 585
R624 vdd.n2092 vdd.n2091 585
R625 vdd.n2090 vdd.n2089 585
R626 vdd.n2085 vdd.n2084 585
R627 vdd.n2168 vdd.n2167 585
R628 vdd.n2166 vdd.n2133 585
R629 vdd.n2165 vdd.n2164 585
R630 vdd.n2136 vdd.n2134 585
R631 vdd.n2159 vdd.n2158 585
R632 vdd.n2157 vdd.n2156 585
R633 vdd.n2140 vdd.n2139 585
R634 vdd.n2151 vdd.n2150 585
R635 vdd.n2149 vdd.n2148 585
R636 vdd.n2144 vdd.n2143 585
R637 vdd.n2007 vdd.n2006 585
R638 vdd.n2005 vdd.n1972 585
R639 vdd.n2004 vdd.n2003 585
R640 vdd.n1975 vdd.n1973 585
R641 vdd.n1998 vdd.n1997 585
R642 vdd.n1996 vdd.n1995 585
R643 vdd.n1979 vdd.n1978 585
R644 vdd.n1990 vdd.n1989 585
R645 vdd.n1988 vdd.n1987 585
R646 vdd.n1983 vdd.n1982 585
R647 vdd.n2066 vdd.n2065 585
R648 vdd.n2064 vdd.n2031 585
R649 vdd.n2063 vdd.n2062 585
R650 vdd.n2034 vdd.n2032 585
R651 vdd.n2057 vdd.n2056 585
R652 vdd.n2055 vdd.n2054 585
R653 vdd.n2038 vdd.n2037 585
R654 vdd.n2049 vdd.n2048 585
R655 vdd.n2047 vdd.n2046 585
R656 vdd.n2042 vdd.n2041 585
R657 vdd.n1906 vdd.n1905 585
R658 vdd.n1904 vdd.n1871 585
R659 vdd.n1903 vdd.n1902 585
R660 vdd.n1874 vdd.n1872 585
R661 vdd.n1897 vdd.n1896 585
R662 vdd.n1895 vdd.n1894 585
R663 vdd.n1878 vdd.n1877 585
R664 vdd.n1889 vdd.n1888 585
R665 vdd.n1887 vdd.n1886 585
R666 vdd.n1882 vdd.n1881 585
R667 vdd.n1965 vdd.n1964 585
R668 vdd.n1963 vdd.n1930 585
R669 vdd.n1962 vdd.n1961 585
R670 vdd.n1933 vdd.n1931 585
R671 vdd.n1956 vdd.n1955 585
R672 vdd.n1954 vdd.n1953 585
R673 vdd.n1937 vdd.n1936 585
R674 vdd.n1948 vdd.n1947 585
R675 vdd.n1946 vdd.n1945 585
R676 vdd.n1941 vdd.n1940 585
R677 vdd.n3448 vdd.n392 509.269
R678 vdd.n3444 vdd.n393 509.269
R679 vdd.n3316 vdd.n685 509.269
R680 vdd.n3313 vdd.n684 509.269
R681 vdd.n2264 vdd.n1437 509.269
R682 vdd.n2267 vdd.n2266 509.269
R683 vdd.n1586 vdd.n1550 509.269
R684 vdd.n1782 vdd.n1551 509.269
R685 vdd.n305 vdd.t160 329.043
R686 vdd.n246 vdd.t240 329.043
R687 vdd.n203 vdd.t291 329.043
R688 vdd.n144 vdd.t228 329.043
R689 vdd.n102 vdd.t197 329.043
R690 vdd.n43 vdd.t189 329.043
R691 vdd.n2086 vdd.t282 329.043
R692 vdd.n2145 vdd.t220 329.043
R693 vdd.n1984 vdd.t271 329.043
R694 vdd.n2043 vdd.t145 329.043
R695 vdd.n1883 vdd.t191 329.043
R696 vdd.n1942 vdd.t196 329.043
R697 vdd.n1679 vdd.t93 319.788
R698 vdd.n1717 vdd.t110 319.788
R699 vdd.n1613 vdd.t123 319.788
R700 vdd.n2269 vdd.t68 319.788
R701 vdd.n1190 vdd.t98 319.788
R702 vdd.n1150 vdd.t119 319.788
R703 vdd.n426 vdd.t88 319.788
R704 vdd.n440 vdd.t78 319.788
R705 vdd.n452 vdd.t95 319.788
R706 vdd.n768 vdd.t72 319.788
R707 vdd.n3276 vdd.t86 319.788
R708 vdd.n688 vdd.t65 319.788
R709 vdd.n1680 vdd.t92 303.69
R710 vdd.n1718 vdd.t109 303.69
R711 vdd.n1614 vdd.t122 303.69
R712 vdd.n2270 vdd.t69 303.69
R713 vdd.n1191 vdd.t99 303.69
R714 vdd.n1151 vdd.t120 303.69
R715 vdd.n427 vdd.t89 303.69
R716 vdd.n441 vdd.t79 303.69
R717 vdd.n453 vdd.t96 303.69
R718 vdd.n769 vdd.t71 303.69
R719 vdd.n3277 vdd.t85 303.69
R720 vdd.n689 vdd.t64 303.69
R721 vdd.n2936 vdd.n927 291.221
R722 vdd.n3150 vdd.n809 291.221
R723 vdd.n3087 vdd.n806 291.221
R724 vdd.n2868 vdd.n2867 291.221
R725 vdd.n2664 vdd.n969 291.221
R726 vdd.n2595 vdd.n2594 291.221
R727 vdd.n1309 vdd.n1308 291.221
R728 vdd.n2415 vdd.n1075 291.221
R729 vdd.n3066 vdd.n807 291.221
R730 vdd.n3153 vdd.n3152 291.221
R731 vdd.n2772 vdd.n2698 291.221
R732 vdd.n2940 vdd.n931 291.221
R733 vdd.n2592 vdd.n979 291.221
R734 vdd.n977 vdd.n951 291.221
R735 vdd.n1387 vdd.n1116 291.221
R736 vdd.n2419 vdd.n1080 291.221
R737 vdd.n3068 vdd.n807 185
R738 vdd.n3151 vdd.n807 185
R739 vdd.n3070 vdd.n3069 185
R740 vdd.n3069 vdd.n805 185
R741 vdd.n3071 vdd.n839 185
R742 vdd.n3081 vdd.n839 185
R743 vdd.n3072 vdd.n848 185
R744 vdd.n848 vdd.n846 185
R745 vdd.n3074 vdd.n3073 185
R746 vdd.n3075 vdd.n3074 185
R747 vdd.n3027 vdd.n847 185
R748 vdd.n847 vdd.n843 185
R749 vdd.n3026 vdd.n3025 185
R750 vdd.n3025 vdd.n3024 185
R751 vdd.n850 vdd.n849 185
R752 vdd.n851 vdd.n850 185
R753 vdd.n3017 vdd.n3016 185
R754 vdd.n3018 vdd.n3017 185
R755 vdd.n3015 vdd.n860 185
R756 vdd.n860 vdd.n857 185
R757 vdd.n3014 vdd.n3013 185
R758 vdd.n3013 vdd.n3012 185
R759 vdd.n862 vdd.n861 185
R760 vdd.n870 vdd.n862 185
R761 vdd.n3005 vdd.n3004 185
R762 vdd.n3006 vdd.n3005 185
R763 vdd.n3002 vdd.n871 185
R764 vdd.n878 vdd.n871 185
R765 vdd.n3001 vdd.n3000 185
R766 vdd.n3000 vdd.n2999 185
R767 vdd.n874 vdd.n873 185
R768 vdd.n875 vdd.n874 185
R769 vdd.n2992 vdd.n2991 185
R770 vdd.n2993 vdd.n2992 185
R771 vdd.n2990 vdd.n885 185
R772 vdd.n885 vdd.n882 185
R773 vdd.n2989 vdd.n2988 185
R774 vdd.n2988 vdd.n2987 185
R775 vdd.n887 vdd.n886 185
R776 vdd.n895 vdd.n887 185
R777 vdd.n2980 vdd.n2979 185
R778 vdd.n2981 vdd.n2980 185
R779 vdd.n2978 vdd.n896 185
R780 vdd.n901 vdd.n896 185
R781 vdd.n2977 vdd.n2976 185
R782 vdd.n2976 vdd.n2975 185
R783 vdd.n898 vdd.n897 185
R784 vdd.n2847 vdd.n898 185
R785 vdd.n2968 vdd.n2967 185
R786 vdd.n2969 vdd.n2968 185
R787 vdd.n2966 vdd.n908 185
R788 vdd.n908 vdd.n905 185
R789 vdd.n2965 vdd.n2964 185
R790 vdd.n2964 vdd.n2963 185
R791 vdd.n910 vdd.n909 185
R792 vdd.n911 vdd.n910 185
R793 vdd.n2956 vdd.n2955 185
R794 vdd.n2957 vdd.n2956 185
R795 vdd.n2954 vdd.n920 185
R796 vdd.n920 vdd.n917 185
R797 vdd.n2953 vdd.n2952 185
R798 vdd.n2952 vdd.n2951 185
R799 vdd.n922 vdd.n921 185
R800 vdd.n2862 vdd.n922 185
R801 vdd.n2944 vdd.n2943 185
R802 vdd.n2945 vdd.n2944 185
R803 vdd.n2942 vdd.n931 185
R804 vdd.n931 vdd.n928 185
R805 vdd.n2941 vdd.n2940 185
R806 vdd.n933 vdd.n932 185
R807 vdd.n2708 vdd.n2707 185
R808 vdd.n2710 vdd.n2709 185
R809 vdd.n2712 vdd.n2711 185
R810 vdd.n2714 vdd.n2713 185
R811 vdd.n2716 vdd.n2715 185
R812 vdd.n2718 vdd.n2717 185
R813 vdd.n2720 vdd.n2719 185
R814 vdd.n2722 vdd.n2721 185
R815 vdd.n2724 vdd.n2723 185
R816 vdd.n2726 vdd.n2725 185
R817 vdd.n2728 vdd.n2727 185
R818 vdd.n2730 vdd.n2729 185
R819 vdd.n2732 vdd.n2731 185
R820 vdd.n2734 vdd.n2733 185
R821 vdd.n2736 vdd.n2735 185
R822 vdd.n2738 vdd.n2737 185
R823 vdd.n2740 vdd.n2739 185
R824 vdd.n2742 vdd.n2741 185
R825 vdd.n2744 vdd.n2743 185
R826 vdd.n2746 vdd.n2745 185
R827 vdd.n2748 vdd.n2747 185
R828 vdd.n2750 vdd.n2749 185
R829 vdd.n2752 vdd.n2751 185
R830 vdd.n2754 vdd.n2753 185
R831 vdd.n2756 vdd.n2755 185
R832 vdd.n2758 vdd.n2757 185
R833 vdd.n2760 vdd.n2759 185
R834 vdd.n2762 vdd.n2761 185
R835 vdd.n2764 vdd.n2763 185
R836 vdd.n2766 vdd.n2765 185
R837 vdd.n2768 vdd.n2767 185
R838 vdd.n2770 vdd.n2769 185
R839 vdd.n2771 vdd.n2698 185
R840 vdd.n2938 vdd.n2698 185
R841 vdd.n3154 vdd.n3153 185
R842 vdd.n3155 vdd.n798 185
R843 vdd.n3157 vdd.n3156 185
R844 vdd.n3159 vdd.n796 185
R845 vdd.n3161 vdd.n3160 185
R846 vdd.n3162 vdd.n795 185
R847 vdd.n3164 vdd.n3163 185
R848 vdd.n3166 vdd.n793 185
R849 vdd.n3168 vdd.n3167 185
R850 vdd.n3169 vdd.n792 185
R851 vdd.n3171 vdd.n3170 185
R852 vdd.n3173 vdd.n790 185
R853 vdd.n3175 vdd.n3174 185
R854 vdd.n3176 vdd.n789 185
R855 vdd.n3178 vdd.n3177 185
R856 vdd.n3180 vdd.n788 185
R857 vdd.n3181 vdd.n786 185
R858 vdd.n3184 vdd.n3183 185
R859 vdd.n787 vdd.n785 185
R860 vdd.n3040 vdd.n3039 185
R861 vdd.n3042 vdd.n3041 185
R862 vdd.n3044 vdd.n3036 185
R863 vdd.n3046 vdd.n3045 185
R864 vdd.n3047 vdd.n3035 185
R865 vdd.n3049 vdd.n3048 185
R866 vdd.n3051 vdd.n3033 185
R867 vdd.n3053 vdd.n3052 185
R868 vdd.n3054 vdd.n3032 185
R869 vdd.n3056 vdd.n3055 185
R870 vdd.n3058 vdd.n3030 185
R871 vdd.n3060 vdd.n3059 185
R872 vdd.n3061 vdd.n3029 185
R873 vdd.n3063 vdd.n3062 185
R874 vdd.n3065 vdd.n3028 185
R875 vdd.n3067 vdd.n3066 185
R876 vdd.n3066 vdd.n692 185
R877 vdd.n3152 vdd.n802 185
R878 vdd.n3152 vdd.n3151 185
R879 vdd.n2775 vdd.n804 185
R880 vdd.n805 vdd.n804 185
R881 vdd.n2776 vdd.n838 185
R882 vdd.n3081 vdd.n838 185
R883 vdd.n2778 vdd.n2777 185
R884 vdd.n2777 vdd.n846 185
R885 vdd.n2779 vdd.n845 185
R886 vdd.n3075 vdd.n845 185
R887 vdd.n2781 vdd.n2780 185
R888 vdd.n2780 vdd.n843 185
R889 vdd.n2782 vdd.n853 185
R890 vdd.n3024 vdd.n853 185
R891 vdd.n2784 vdd.n2783 185
R892 vdd.n2783 vdd.n851 185
R893 vdd.n2785 vdd.n859 185
R894 vdd.n3018 vdd.n859 185
R895 vdd.n2787 vdd.n2786 185
R896 vdd.n2786 vdd.n857 185
R897 vdd.n2788 vdd.n864 185
R898 vdd.n3012 vdd.n864 185
R899 vdd.n2790 vdd.n2789 185
R900 vdd.n2789 vdd.n870 185
R901 vdd.n2791 vdd.n869 185
R902 vdd.n3006 vdd.n869 185
R903 vdd.n2793 vdd.n2792 185
R904 vdd.n2792 vdd.n878 185
R905 vdd.n2794 vdd.n877 185
R906 vdd.n2999 vdd.n877 185
R907 vdd.n2796 vdd.n2795 185
R908 vdd.n2795 vdd.n875 185
R909 vdd.n2797 vdd.n884 185
R910 vdd.n2993 vdd.n884 185
R911 vdd.n2799 vdd.n2798 185
R912 vdd.n2798 vdd.n882 185
R913 vdd.n2800 vdd.n889 185
R914 vdd.n2987 vdd.n889 185
R915 vdd.n2802 vdd.n2801 185
R916 vdd.n2801 vdd.n895 185
R917 vdd.n2803 vdd.n894 185
R918 vdd.n2981 vdd.n894 185
R919 vdd.n2805 vdd.n2804 185
R920 vdd.n2804 vdd.n901 185
R921 vdd.n2806 vdd.n900 185
R922 vdd.n2975 vdd.n900 185
R923 vdd.n2849 vdd.n2848 185
R924 vdd.n2848 vdd.n2847 185
R925 vdd.n2850 vdd.n907 185
R926 vdd.n2969 vdd.n907 185
R927 vdd.n2852 vdd.n2851 185
R928 vdd.n2851 vdd.n905 185
R929 vdd.n2853 vdd.n913 185
R930 vdd.n2963 vdd.n913 185
R931 vdd.n2855 vdd.n2854 185
R932 vdd.n2854 vdd.n911 185
R933 vdd.n2856 vdd.n919 185
R934 vdd.n2957 vdd.n919 185
R935 vdd.n2858 vdd.n2857 185
R936 vdd.n2857 vdd.n917 185
R937 vdd.n2859 vdd.n924 185
R938 vdd.n2951 vdd.n924 185
R939 vdd.n2861 vdd.n2860 185
R940 vdd.n2862 vdd.n2861 185
R941 vdd.n2774 vdd.n930 185
R942 vdd.n2945 vdd.n930 185
R943 vdd.n2773 vdd.n2772 185
R944 vdd.n2772 vdd.n928 185
R945 vdd.n2264 vdd.n2263 185
R946 vdd.n2265 vdd.n2264 185
R947 vdd.n1438 vdd.n1436 185
R948 vdd.n2256 vdd.n1436 185
R949 vdd.n2259 vdd.n2258 185
R950 vdd.n2258 vdd.n2257 185
R951 vdd.n1441 vdd.n1440 185
R952 vdd.n1442 vdd.n1441 185
R953 vdd.n2245 vdd.n2244 185
R954 vdd.n2246 vdd.n2245 185
R955 vdd.n1450 vdd.n1449 185
R956 vdd.n2237 vdd.n1449 185
R957 vdd.n2240 vdd.n2239 185
R958 vdd.n2239 vdd.n2238 185
R959 vdd.n1453 vdd.n1452 185
R960 vdd.n1460 vdd.n1453 185
R961 vdd.n2228 vdd.n2227 185
R962 vdd.n2229 vdd.n2228 185
R963 vdd.n1462 vdd.n1461 185
R964 vdd.n1461 vdd.n1459 185
R965 vdd.n2223 vdd.n2222 185
R966 vdd.n2222 vdd.n2221 185
R967 vdd.n1465 vdd.n1464 185
R968 vdd.n1466 vdd.n1465 185
R969 vdd.n2212 vdd.n2211 185
R970 vdd.n2213 vdd.n2212 185
R971 vdd.n1473 vdd.n1472 185
R972 vdd.n2204 vdd.n1472 185
R973 vdd.n2207 vdd.n2206 185
R974 vdd.n2206 vdd.n2205 185
R975 vdd.n1476 vdd.n1475 185
R976 vdd.n1482 vdd.n1476 185
R977 vdd.n2195 vdd.n2194 185
R978 vdd.n2196 vdd.n2195 185
R979 vdd.n1484 vdd.n1483 185
R980 vdd.n2187 vdd.n1483 185
R981 vdd.n2190 vdd.n2189 185
R982 vdd.n2189 vdd.n2188 185
R983 vdd.n1487 vdd.n1486 185
R984 vdd.n1488 vdd.n1487 185
R985 vdd.n2178 vdd.n2177 185
R986 vdd.n2179 vdd.n2178 185
R987 vdd.n1496 vdd.n1495 185
R988 vdd.n1495 vdd.n1494 185
R989 vdd.n1866 vdd.n1865 185
R990 vdd.n1865 vdd.n1864 185
R991 vdd.n1499 vdd.n1498 185
R992 vdd.n1505 vdd.n1499 185
R993 vdd.n1855 vdd.n1854 185
R994 vdd.n1856 vdd.n1855 185
R995 vdd.n1507 vdd.n1506 185
R996 vdd.n1847 vdd.n1506 185
R997 vdd.n1850 vdd.n1849 185
R998 vdd.n1849 vdd.n1848 185
R999 vdd.n1510 vdd.n1509 185
R1000 vdd.n1517 vdd.n1510 185
R1001 vdd.n1838 vdd.n1837 185
R1002 vdd.n1839 vdd.n1838 185
R1003 vdd.n1519 vdd.n1518 185
R1004 vdd.n1518 vdd.n1516 185
R1005 vdd.n1833 vdd.n1832 185
R1006 vdd.n1832 vdd.n1831 185
R1007 vdd.n1522 vdd.n1521 185
R1008 vdd.n1523 vdd.n1522 185
R1009 vdd.n1822 vdd.n1821 185
R1010 vdd.n1823 vdd.n1822 185
R1011 vdd.n1530 vdd.n1529 185
R1012 vdd.n1814 vdd.n1529 185
R1013 vdd.n1817 vdd.n1816 185
R1014 vdd.n1816 vdd.n1815 185
R1015 vdd.n1533 vdd.n1532 185
R1016 vdd.n1539 vdd.n1533 185
R1017 vdd.n1805 vdd.n1804 185
R1018 vdd.n1806 vdd.n1805 185
R1019 vdd.n1541 vdd.n1540 185
R1020 vdd.n1797 vdd.n1540 185
R1021 vdd.n1800 vdd.n1799 185
R1022 vdd.n1799 vdd.n1798 185
R1023 vdd.n1544 vdd.n1543 185
R1024 vdd.n1545 vdd.n1544 185
R1025 vdd.n1788 vdd.n1787 185
R1026 vdd.n1789 vdd.n1788 185
R1027 vdd.n1552 vdd.n1551 185
R1028 vdd.n1587 vdd.n1551 185
R1029 vdd.n1783 vdd.n1782 185
R1030 vdd.n1555 vdd.n1554 185
R1031 vdd.n1779 vdd.n1778 185
R1032 vdd.n1780 vdd.n1779 185
R1033 vdd.n1589 vdd.n1588 185
R1034 vdd.n1774 vdd.n1591 185
R1035 vdd.n1773 vdd.n1592 185
R1036 vdd.n1772 vdd.n1593 185
R1037 vdd.n1595 vdd.n1594 185
R1038 vdd.n1768 vdd.n1597 185
R1039 vdd.n1767 vdd.n1598 185
R1040 vdd.n1766 vdd.n1599 185
R1041 vdd.n1601 vdd.n1600 185
R1042 vdd.n1762 vdd.n1603 185
R1043 vdd.n1761 vdd.n1604 185
R1044 vdd.n1760 vdd.n1605 185
R1045 vdd.n1607 vdd.n1606 185
R1046 vdd.n1756 vdd.n1609 185
R1047 vdd.n1755 vdd.n1610 185
R1048 vdd.n1754 vdd.n1611 185
R1049 vdd.n1615 vdd.n1612 185
R1050 vdd.n1750 vdd.n1617 185
R1051 vdd.n1749 vdd.n1618 185
R1052 vdd.n1748 vdd.n1619 185
R1053 vdd.n1621 vdd.n1620 185
R1054 vdd.n1744 vdd.n1623 185
R1055 vdd.n1743 vdd.n1624 185
R1056 vdd.n1742 vdd.n1625 185
R1057 vdd.n1627 vdd.n1626 185
R1058 vdd.n1738 vdd.n1629 185
R1059 vdd.n1737 vdd.n1630 185
R1060 vdd.n1736 vdd.n1631 185
R1061 vdd.n1633 vdd.n1632 185
R1062 vdd.n1732 vdd.n1635 185
R1063 vdd.n1731 vdd.n1636 185
R1064 vdd.n1730 vdd.n1637 185
R1065 vdd.n1639 vdd.n1638 185
R1066 vdd.n1726 vdd.n1641 185
R1067 vdd.n1725 vdd.n1642 185
R1068 vdd.n1724 vdd.n1643 185
R1069 vdd.n1645 vdd.n1644 185
R1070 vdd.n1720 vdd.n1647 185
R1071 vdd.n1719 vdd.n1716 185
R1072 vdd.n1715 vdd.n1648 185
R1073 vdd.n1650 vdd.n1649 185
R1074 vdd.n1711 vdd.n1652 185
R1075 vdd.n1710 vdd.n1653 185
R1076 vdd.n1709 vdd.n1654 185
R1077 vdd.n1656 vdd.n1655 185
R1078 vdd.n1705 vdd.n1658 185
R1079 vdd.n1704 vdd.n1659 185
R1080 vdd.n1703 vdd.n1660 185
R1081 vdd.n1662 vdd.n1661 185
R1082 vdd.n1699 vdd.n1664 185
R1083 vdd.n1698 vdd.n1665 185
R1084 vdd.n1697 vdd.n1666 185
R1085 vdd.n1668 vdd.n1667 185
R1086 vdd.n1693 vdd.n1670 185
R1087 vdd.n1692 vdd.n1671 185
R1088 vdd.n1691 vdd.n1672 185
R1089 vdd.n1674 vdd.n1673 185
R1090 vdd.n1687 vdd.n1676 185
R1091 vdd.n1686 vdd.n1677 185
R1092 vdd.n1685 vdd.n1678 185
R1093 vdd.n1682 vdd.n1586 185
R1094 vdd.n1780 vdd.n1586 185
R1095 vdd.n2268 vdd.n2267 185
R1096 vdd.n2272 vdd.n1432 185
R1097 vdd.n1431 vdd.n1425 185
R1098 vdd.n1429 vdd.n1428 185
R1099 vdd.n1427 vdd.n1221 185
R1100 vdd.n2276 vdd.n1218 185
R1101 vdd.n2278 vdd.n2277 185
R1102 vdd.n2280 vdd.n1216 185
R1103 vdd.n2282 vdd.n2281 185
R1104 vdd.n2283 vdd.n1211 185
R1105 vdd.n2285 vdd.n2284 185
R1106 vdd.n2287 vdd.n1209 185
R1107 vdd.n2289 vdd.n2288 185
R1108 vdd.n2290 vdd.n1204 185
R1109 vdd.n2292 vdd.n2291 185
R1110 vdd.n2294 vdd.n1202 185
R1111 vdd.n2296 vdd.n2295 185
R1112 vdd.n2297 vdd.n1198 185
R1113 vdd.n2299 vdd.n2298 185
R1114 vdd.n2301 vdd.n1195 185
R1115 vdd.n2303 vdd.n2302 185
R1116 vdd.n1196 vdd.n1189 185
R1117 vdd.n2307 vdd.n1193 185
R1118 vdd.n2308 vdd.n1185 185
R1119 vdd.n2310 vdd.n2309 185
R1120 vdd.n2312 vdd.n1183 185
R1121 vdd.n2314 vdd.n2313 185
R1122 vdd.n2315 vdd.n1178 185
R1123 vdd.n2317 vdd.n2316 185
R1124 vdd.n2319 vdd.n1176 185
R1125 vdd.n2321 vdd.n2320 185
R1126 vdd.n2322 vdd.n1171 185
R1127 vdd.n2324 vdd.n2323 185
R1128 vdd.n2326 vdd.n1169 185
R1129 vdd.n2328 vdd.n2327 185
R1130 vdd.n2329 vdd.n1164 185
R1131 vdd.n2331 vdd.n2330 185
R1132 vdd.n2333 vdd.n1162 185
R1133 vdd.n2335 vdd.n2334 185
R1134 vdd.n2336 vdd.n1158 185
R1135 vdd.n2338 vdd.n2337 185
R1136 vdd.n2340 vdd.n1155 185
R1137 vdd.n2342 vdd.n2341 185
R1138 vdd.n1156 vdd.n1149 185
R1139 vdd.n2346 vdd.n1153 185
R1140 vdd.n2347 vdd.n1145 185
R1141 vdd.n2349 vdd.n2348 185
R1142 vdd.n2351 vdd.n1143 185
R1143 vdd.n2353 vdd.n2352 185
R1144 vdd.n2354 vdd.n1138 185
R1145 vdd.n2356 vdd.n2355 185
R1146 vdd.n2358 vdd.n1136 185
R1147 vdd.n2360 vdd.n2359 185
R1148 vdd.n2361 vdd.n1131 185
R1149 vdd.n2363 vdd.n2362 185
R1150 vdd.n2365 vdd.n1129 185
R1151 vdd.n2367 vdd.n2366 185
R1152 vdd.n2368 vdd.n1127 185
R1153 vdd.n2370 vdd.n2369 185
R1154 vdd.n2373 vdd.n2372 185
R1155 vdd.n2375 vdd.n2374 185
R1156 vdd.n2377 vdd.n1125 185
R1157 vdd.n2379 vdd.n2378 185
R1158 vdd.n1437 vdd.n1124 185
R1159 vdd.n2266 vdd.n1435 185
R1160 vdd.n2266 vdd.n2265 185
R1161 vdd.n1445 vdd.n1434 185
R1162 vdd.n2256 vdd.n1434 185
R1163 vdd.n2255 vdd.n2254 185
R1164 vdd.n2257 vdd.n2255 185
R1165 vdd.n1444 vdd.n1443 185
R1166 vdd.n1443 vdd.n1442 185
R1167 vdd.n2248 vdd.n2247 185
R1168 vdd.n2247 vdd.n2246 185
R1169 vdd.n1448 vdd.n1447 185
R1170 vdd.n2237 vdd.n1448 185
R1171 vdd.n2236 vdd.n2235 185
R1172 vdd.n2238 vdd.n2236 185
R1173 vdd.n1455 vdd.n1454 185
R1174 vdd.n1460 vdd.n1454 185
R1175 vdd.n2231 vdd.n2230 185
R1176 vdd.n2230 vdd.n2229 185
R1177 vdd.n1458 vdd.n1457 185
R1178 vdd.n1459 vdd.n1458 185
R1179 vdd.n2220 vdd.n2219 185
R1180 vdd.n2221 vdd.n2220 185
R1181 vdd.n1468 vdd.n1467 185
R1182 vdd.n1467 vdd.n1466 185
R1183 vdd.n2215 vdd.n2214 185
R1184 vdd.n2214 vdd.n2213 185
R1185 vdd.n1471 vdd.n1470 185
R1186 vdd.n2204 vdd.n1471 185
R1187 vdd.n2203 vdd.n2202 185
R1188 vdd.n2205 vdd.n2203 185
R1189 vdd.n1478 vdd.n1477 185
R1190 vdd.n1482 vdd.n1477 185
R1191 vdd.n2198 vdd.n2197 185
R1192 vdd.n2197 vdd.n2196 185
R1193 vdd.n1481 vdd.n1480 185
R1194 vdd.n2187 vdd.n1481 185
R1195 vdd.n2186 vdd.n2185 185
R1196 vdd.n2188 vdd.n2186 185
R1197 vdd.n1490 vdd.n1489 185
R1198 vdd.n1489 vdd.n1488 185
R1199 vdd.n2181 vdd.n2180 185
R1200 vdd.n2180 vdd.n2179 185
R1201 vdd.n1493 vdd.n1492 185
R1202 vdd.n1494 vdd.n1493 185
R1203 vdd.n1863 vdd.n1862 185
R1204 vdd.n1864 vdd.n1863 185
R1205 vdd.n1501 vdd.n1500 185
R1206 vdd.n1505 vdd.n1500 185
R1207 vdd.n1858 vdd.n1857 185
R1208 vdd.n1857 vdd.n1856 185
R1209 vdd.n1504 vdd.n1503 185
R1210 vdd.n1847 vdd.n1504 185
R1211 vdd.n1846 vdd.n1845 185
R1212 vdd.n1848 vdd.n1846 185
R1213 vdd.n1512 vdd.n1511 185
R1214 vdd.n1517 vdd.n1511 185
R1215 vdd.n1841 vdd.n1840 185
R1216 vdd.n1840 vdd.n1839 185
R1217 vdd.n1515 vdd.n1514 185
R1218 vdd.n1516 vdd.n1515 185
R1219 vdd.n1830 vdd.n1829 185
R1220 vdd.n1831 vdd.n1830 185
R1221 vdd.n1525 vdd.n1524 185
R1222 vdd.n1524 vdd.n1523 185
R1223 vdd.n1825 vdd.n1824 185
R1224 vdd.n1824 vdd.n1823 185
R1225 vdd.n1528 vdd.n1527 185
R1226 vdd.n1814 vdd.n1528 185
R1227 vdd.n1813 vdd.n1812 185
R1228 vdd.n1815 vdd.n1813 185
R1229 vdd.n1535 vdd.n1534 185
R1230 vdd.n1539 vdd.n1534 185
R1231 vdd.n1808 vdd.n1807 185
R1232 vdd.n1807 vdd.n1806 185
R1233 vdd.n1538 vdd.n1537 185
R1234 vdd.n1797 vdd.n1538 185
R1235 vdd.n1796 vdd.n1795 185
R1236 vdd.n1798 vdd.n1796 185
R1237 vdd.n1547 vdd.n1546 185
R1238 vdd.n1546 vdd.n1545 185
R1239 vdd.n1791 vdd.n1790 185
R1240 vdd.n1790 vdd.n1789 185
R1241 vdd.n1550 vdd.n1549 185
R1242 vdd.n1587 vdd.n1550 185
R1243 vdd.n971 vdd.n969 185
R1244 vdd.n2593 vdd.n969 185
R1245 vdd.n2515 vdd.n989 185
R1246 vdd.n989 vdd.n976 185
R1247 vdd.n2517 vdd.n2516 185
R1248 vdd.n2518 vdd.n2517 185
R1249 vdd.n2514 vdd.n988 185
R1250 vdd.n1338 vdd.n988 185
R1251 vdd.n2513 vdd.n2512 185
R1252 vdd.n2512 vdd.n2511 185
R1253 vdd.n991 vdd.n990 185
R1254 vdd.n992 vdd.n991 185
R1255 vdd.n2502 vdd.n2501 185
R1256 vdd.n2503 vdd.n2502 185
R1257 vdd.n2500 vdd.n1002 185
R1258 vdd.n1002 vdd.n999 185
R1259 vdd.n2499 vdd.n2498 185
R1260 vdd.n2498 vdd.n2497 185
R1261 vdd.n1004 vdd.n1003 185
R1262 vdd.n1005 vdd.n1004 185
R1263 vdd.n2490 vdd.n2489 185
R1264 vdd.n2491 vdd.n2490 185
R1265 vdd.n2488 vdd.n1013 185
R1266 vdd.n1018 vdd.n1013 185
R1267 vdd.n2487 vdd.n2486 185
R1268 vdd.n2486 vdd.n2485 185
R1269 vdd.n1015 vdd.n1014 185
R1270 vdd.n1024 vdd.n1015 185
R1271 vdd.n2478 vdd.n2477 185
R1272 vdd.n2479 vdd.n2478 185
R1273 vdd.n2476 vdd.n1025 185
R1274 vdd.n1359 vdd.n1025 185
R1275 vdd.n2475 vdd.n2474 185
R1276 vdd.n2474 vdd.n2473 185
R1277 vdd.n1027 vdd.n1026 185
R1278 vdd.n1028 vdd.n1027 185
R1279 vdd.n2466 vdd.n2465 185
R1280 vdd.n2467 vdd.n2466 185
R1281 vdd.n2464 vdd.n1037 185
R1282 vdd.n1037 vdd.n1034 185
R1283 vdd.n2463 vdd.n2462 185
R1284 vdd.n2462 vdd.n2461 185
R1285 vdd.n1039 vdd.n1038 185
R1286 vdd.n1048 vdd.n1039 185
R1287 vdd.n2453 vdd.n2452 185
R1288 vdd.n2454 vdd.n2453 185
R1289 vdd.n2451 vdd.n1049 185
R1290 vdd.n1055 vdd.n1049 185
R1291 vdd.n2450 vdd.n2449 185
R1292 vdd.n2449 vdd.n2448 185
R1293 vdd.n1051 vdd.n1050 185
R1294 vdd.n1052 vdd.n1051 185
R1295 vdd.n2441 vdd.n2440 185
R1296 vdd.n2442 vdd.n2441 185
R1297 vdd.n2439 vdd.n1062 185
R1298 vdd.n1062 vdd.n1059 185
R1299 vdd.n2438 vdd.n2437 185
R1300 vdd.n2437 vdd.n2436 185
R1301 vdd.n1064 vdd.n1063 185
R1302 vdd.n1065 vdd.n1064 185
R1303 vdd.n2429 vdd.n2428 185
R1304 vdd.n2430 vdd.n2429 185
R1305 vdd.n2427 vdd.n1073 185
R1306 vdd.n1079 vdd.n1073 185
R1307 vdd.n2426 vdd.n2425 185
R1308 vdd.n2425 vdd.n2424 185
R1309 vdd.n1075 vdd.n1074 185
R1310 vdd.n1076 vdd.n1075 185
R1311 vdd.n2415 vdd.n2414 185
R1312 vdd.n2413 vdd.n1118 185
R1313 vdd.n2412 vdd.n1117 185
R1314 vdd.n2417 vdd.n1117 185
R1315 vdd.n2411 vdd.n2410 185
R1316 vdd.n2409 vdd.n2408 185
R1317 vdd.n2407 vdd.n2406 185
R1318 vdd.n2405 vdd.n2404 185
R1319 vdd.n2403 vdd.n2402 185
R1320 vdd.n2401 vdd.n2400 185
R1321 vdd.n2399 vdd.n2398 185
R1322 vdd.n2397 vdd.n2396 185
R1323 vdd.n2395 vdd.n2394 185
R1324 vdd.n2393 vdd.n2392 185
R1325 vdd.n2391 vdd.n2390 185
R1326 vdd.n2389 vdd.n2388 185
R1327 vdd.n2387 vdd.n2386 185
R1328 vdd.n2385 vdd.n2384 185
R1329 vdd.n2383 vdd.n2382 185
R1330 vdd.n1275 vdd.n1119 185
R1331 vdd.n1277 vdd.n1276 185
R1332 vdd.n1279 vdd.n1278 185
R1333 vdd.n1281 vdd.n1280 185
R1334 vdd.n1283 vdd.n1282 185
R1335 vdd.n1285 vdd.n1284 185
R1336 vdd.n1287 vdd.n1286 185
R1337 vdd.n1289 vdd.n1288 185
R1338 vdd.n1291 vdd.n1290 185
R1339 vdd.n1293 vdd.n1292 185
R1340 vdd.n1295 vdd.n1294 185
R1341 vdd.n1297 vdd.n1296 185
R1342 vdd.n1299 vdd.n1298 185
R1343 vdd.n1301 vdd.n1300 185
R1344 vdd.n1304 vdd.n1303 185
R1345 vdd.n1306 vdd.n1305 185
R1346 vdd.n1308 vdd.n1307 185
R1347 vdd.n2596 vdd.n2595 185
R1348 vdd.n2598 vdd.n2597 185
R1349 vdd.n2600 vdd.n2599 185
R1350 vdd.n2603 vdd.n2602 185
R1351 vdd.n2605 vdd.n2604 185
R1352 vdd.n2607 vdd.n2606 185
R1353 vdd.n2609 vdd.n2608 185
R1354 vdd.n2611 vdd.n2610 185
R1355 vdd.n2613 vdd.n2612 185
R1356 vdd.n2615 vdd.n2614 185
R1357 vdd.n2617 vdd.n2616 185
R1358 vdd.n2619 vdd.n2618 185
R1359 vdd.n2621 vdd.n2620 185
R1360 vdd.n2623 vdd.n2622 185
R1361 vdd.n2625 vdd.n2624 185
R1362 vdd.n2627 vdd.n2626 185
R1363 vdd.n2629 vdd.n2628 185
R1364 vdd.n2631 vdd.n2630 185
R1365 vdd.n2633 vdd.n2632 185
R1366 vdd.n2635 vdd.n2634 185
R1367 vdd.n2637 vdd.n2636 185
R1368 vdd.n2639 vdd.n2638 185
R1369 vdd.n2641 vdd.n2640 185
R1370 vdd.n2643 vdd.n2642 185
R1371 vdd.n2645 vdd.n2644 185
R1372 vdd.n2647 vdd.n2646 185
R1373 vdd.n2649 vdd.n2648 185
R1374 vdd.n2651 vdd.n2650 185
R1375 vdd.n2653 vdd.n2652 185
R1376 vdd.n2655 vdd.n2654 185
R1377 vdd.n2657 vdd.n2656 185
R1378 vdd.n2659 vdd.n2658 185
R1379 vdd.n2661 vdd.n2660 185
R1380 vdd.n2662 vdd.n970 185
R1381 vdd.n2664 vdd.n2663 185
R1382 vdd.n2665 vdd.n2664 185
R1383 vdd.n2594 vdd.n974 185
R1384 vdd.n2594 vdd.n2593 185
R1385 vdd.n1336 vdd.n975 185
R1386 vdd.n976 vdd.n975 185
R1387 vdd.n1337 vdd.n986 185
R1388 vdd.n2518 vdd.n986 185
R1389 vdd.n1340 vdd.n1339 185
R1390 vdd.n1339 vdd.n1338 185
R1391 vdd.n1341 vdd.n993 185
R1392 vdd.n2511 vdd.n993 185
R1393 vdd.n1343 vdd.n1342 185
R1394 vdd.n1342 vdd.n992 185
R1395 vdd.n1344 vdd.n1000 185
R1396 vdd.n2503 vdd.n1000 185
R1397 vdd.n1346 vdd.n1345 185
R1398 vdd.n1345 vdd.n999 185
R1399 vdd.n1347 vdd.n1006 185
R1400 vdd.n2497 vdd.n1006 185
R1401 vdd.n1349 vdd.n1348 185
R1402 vdd.n1348 vdd.n1005 185
R1403 vdd.n1350 vdd.n1011 185
R1404 vdd.n2491 vdd.n1011 185
R1405 vdd.n1352 vdd.n1351 185
R1406 vdd.n1351 vdd.n1018 185
R1407 vdd.n1353 vdd.n1016 185
R1408 vdd.n2485 vdd.n1016 185
R1409 vdd.n1355 vdd.n1354 185
R1410 vdd.n1354 vdd.n1024 185
R1411 vdd.n1356 vdd.n1022 185
R1412 vdd.n2479 vdd.n1022 185
R1413 vdd.n1358 vdd.n1357 185
R1414 vdd.n1359 vdd.n1358 185
R1415 vdd.n1335 vdd.n1029 185
R1416 vdd.n2473 vdd.n1029 185
R1417 vdd.n1334 vdd.n1333 185
R1418 vdd.n1333 vdd.n1028 185
R1419 vdd.n1332 vdd.n1035 185
R1420 vdd.n2467 vdd.n1035 185
R1421 vdd.n1331 vdd.n1330 185
R1422 vdd.n1330 vdd.n1034 185
R1423 vdd.n1329 vdd.n1040 185
R1424 vdd.n2461 vdd.n1040 185
R1425 vdd.n1328 vdd.n1327 185
R1426 vdd.n1327 vdd.n1048 185
R1427 vdd.n1326 vdd.n1046 185
R1428 vdd.n2454 vdd.n1046 185
R1429 vdd.n1325 vdd.n1324 185
R1430 vdd.n1324 vdd.n1055 185
R1431 vdd.n1323 vdd.n1053 185
R1432 vdd.n2448 vdd.n1053 185
R1433 vdd.n1322 vdd.n1321 185
R1434 vdd.n1321 vdd.n1052 185
R1435 vdd.n1320 vdd.n1060 185
R1436 vdd.n2442 vdd.n1060 185
R1437 vdd.n1319 vdd.n1318 185
R1438 vdd.n1318 vdd.n1059 185
R1439 vdd.n1317 vdd.n1066 185
R1440 vdd.n2436 vdd.n1066 185
R1441 vdd.n1316 vdd.n1315 185
R1442 vdd.n1315 vdd.n1065 185
R1443 vdd.n1314 vdd.n1071 185
R1444 vdd.n2430 vdd.n1071 185
R1445 vdd.n1313 vdd.n1312 185
R1446 vdd.n1312 vdd.n1079 185
R1447 vdd.n1311 vdd.n1077 185
R1448 vdd.n2424 vdd.n1077 185
R1449 vdd.n1310 vdd.n1309 185
R1450 vdd.n1309 vdd.n1076 185
R1451 vdd.n3449 vdd.n3448 185
R1452 vdd.n3448 vdd.n3447 185
R1453 vdd.n3450 vdd.n387 185
R1454 vdd.n387 vdd.n386 185
R1455 vdd.n3452 vdd.n3451 185
R1456 vdd.n3453 vdd.n3452 185
R1457 vdd.n382 vdd.n381 185
R1458 vdd.n3454 vdd.n382 185
R1459 vdd.n3457 vdd.n3456 185
R1460 vdd.n3456 vdd.n3455 185
R1461 vdd.n3458 vdd.n376 185
R1462 vdd.n376 vdd.n375 185
R1463 vdd.n3460 vdd.n3459 185
R1464 vdd.n3461 vdd.n3460 185
R1465 vdd.n371 vdd.n370 185
R1466 vdd.n3462 vdd.n371 185
R1467 vdd.n3465 vdd.n3464 185
R1468 vdd.n3464 vdd.n3463 185
R1469 vdd.n3466 vdd.n365 185
R1470 vdd.n3423 vdd.n365 185
R1471 vdd.n3468 vdd.n3467 185
R1472 vdd.n3469 vdd.n3468 185
R1473 vdd.n360 vdd.n359 185
R1474 vdd.n3470 vdd.n360 185
R1475 vdd.n3473 vdd.n3472 185
R1476 vdd.n3472 vdd.n3471 185
R1477 vdd.n3474 vdd.n354 185
R1478 vdd.n361 vdd.n354 185
R1479 vdd.n3476 vdd.n3475 185
R1480 vdd.n3477 vdd.n3476 185
R1481 vdd.n350 vdd.n349 185
R1482 vdd.n3478 vdd.n350 185
R1483 vdd.n3481 vdd.n3480 185
R1484 vdd.n3480 vdd.n3479 185
R1485 vdd.n3482 vdd.n345 185
R1486 vdd.n345 vdd.n344 185
R1487 vdd.n3484 vdd.n3483 185
R1488 vdd.n3485 vdd.n3484 185
R1489 vdd.n339 vdd.n337 185
R1490 vdd.n3486 vdd.n339 185
R1491 vdd.n3489 vdd.n3488 185
R1492 vdd.n3488 vdd.n3487 185
R1493 vdd.n338 vdd.n336 185
R1494 vdd.n340 vdd.n338 185
R1495 vdd.n3399 vdd.n3398 185
R1496 vdd.n3400 vdd.n3399 185
R1497 vdd.n635 vdd.n634 185
R1498 vdd.n634 vdd.n633 185
R1499 vdd.n3394 vdd.n3393 185
R1500 vdd.n3393 vdd.n3392 185
R1501 vdd.n638 vdd.n637 185
R1502 vdd.n644 vdd.n638 185
R1503 vdd.n3380 vdd.n3379 185
R1504 vdd.n3381 vdd.n3380 185
R1505 vdd.n646 vdd.n645 185
R1506 vdd.n3372 vdd.n645 185
R1507 vdd.n3375 vdd.n3374 185
R1508 vdd.n3374 vdd.n3373 185
R1509 vdd.n649 vdd.n648 185
R1510 vdd.n656 vdd.n649 185
R1511 vdd.n3363 vdd.n3362 185
R1512 vdd.n3364 vdd.n3363 185
R1513 vdd.n658 vdd.n657 185
R1514 vdd.n657 vdd.n655 185
R1515 vdd.n3358 vdd.n3357 185
R1516 vdd.n3357 vdd.n3356 185
R1517 vdd.n661 vdd.n660 185
R1518 vdd.n662 vdd.n661 185
R1519 vdd.n3347 vdd.n3346 185
R1520 vdd.n3348 vdd.n3347 185
R1521 vdd.n669 vdd.n668 185
R1522 vdd.n3339 vdd.n668 185
R1523 vdd.n3342 vdd.n3341 185
R1524 vdd.n3341 vdd.n3340 185
R1525 vdd.n672 vdd.n671 185
R1526 vdd.n679 vdd.n672 185
R1527 vdd.n3330 vdd.n3329 185
R1528 vdd.n3331 vdd.n3330 185
R1529 vdd.n681 vdd.n680 185
R1530 vdd.n680 vdd.n678 185
R1531 vdd.n3325 vdd.n3324 185
R1532 vdd.n3324 vdd.n3323 185
R1533 vdd.n684 vdd.n683 185
R1534 vdd.n723 vdd.n684 185
R1535 vdd.n3313 vdd.n3312 185
R1536 vdd.n3311 vdd.n725 185
R1537 vdd.n3310 vdd.n724 185
R1538 vdd.n3315 vdd.n724 185
R1539 vdd.n729 vdd.n728 185
R1540 vdd.n733 vdd.n732 185
R1541 vdd.n3306 vdd.n734 185
R1542 vdd.n3305 vdd.n3304 185
R1543 vdd.n3303 vdd.n3302 185
R1544 vdd.n3301 vdd.n3300 185
R1545 vdd.n3299 vdd.n3298 185
R1546 vdd.n3297 vdd.n3296 185
R1547 vdd.n3295 vdd.n3294 185
R1548 vdd.n3293 vdd.n3292 185
R1549 vdd.n3291 vdd.n3290 185
R1550 vdd.n3289 vdd.n3288 185
R1551 vdd.n3287 vdd.n3286 185
R1552 vdd.n3285 vdd.n3284 185
R1553 vdd.n3283 vdd.n3282 185
R1554 vdd.n3281 vdd.n3280 185
R1555 vdd.n3279 vdd.n3278 185
R1556 vdd.n3270 vdd.n747 185
R1557 vdd.n3272 vdd.n3271 185
R1558 vdd.n3269 vdd.n3268 185
R1559 vdd.n3267 vdd.n3266 185
R1560 vdd.n3265 vdd.n3264 185
R1561 vdd.n3263 vdd.n3262 185
R1562 vdd.n3261 vdd.n3260 185
R1563 vdd.n3259 vdd.n3258 185
R1564 vdd.n3257 vdd.n3256 185
R1565 vdd.n3255 vdd.n3254 185
R1566 vdd.n3253 vdd.n3252 185
R1567 vdd.n3251 vdd.n3250 185
R1568 vdd.n3249 vdd.n3248 185
R1569 vdd.n3247 vdd.n3246 185
R1570 vdd.n3245 vdd.n3244 185
R1571 vdd.n3243 vdd.n3242 185
R1572 vdd.n3241 vdd.n3240 185
R1573 vdd.n3239 vdd.n3238 185
R1574 vdd.n3237 vdd.n3236 185
R1575 vdd.n3235 vdd.n3234 185
R1576 vdd.n3233 vdd.n3232 185
R1577 vdd.n3231 vdd.n3230 185
R1578 vdd.n3224 vdd.n767 185
R1579 vdd.n3226 vdd.n3225 185
R1580 vdd.n3223 vdd.n3222 185
R1581 vdd.n3221 vdd.n3220 185
R1582 vdd.n3219 vdd.n3218 185
R1583 vdd.n3217 vdd.n3216 185
R1584 vdd.n3215 vdd.n3214 185
R1585 vdd.n3213 vdd.n3212 185
R1586 vdd.n3211 vdd.n3210 185
R1587 vdd.n3209 vdd.n3208 185
R1588 vdd.n3207 vdd.n3206 185
R1589 vdd.n3205 vdd.n3204 185
R1590 vdd.n3203 vdd.n3202 185
R1591 vdd.n3201 vdd.n3200 185
R1592 vdd.n3199 vdd.n3198 185
R1593 vdd.n3197 vdd.n3196 185
R1594 vdd.n3195 vdd.n3194 185
R1595 vdd.n3193 vdd.n3192 185
R1596 vdd.n3191 vdd.n3190 185
R1597 vdd.n3189 vdd.n3188 185
R1598 vdd.n3187 vdd.n691 185
R1599 vdd.n3317 vdd.n3316 185
R1600 vdd.n3316 vdd.n3315 185
R1601 vdd.n3444 vdd.n3443 185
R1602 vdd.n618 vdd.n425 185
R1603 vdd.n617 vdd.n616 185
R1604 vdd.n615 vdd.n614 185
R1605 vdd.n613 vdd.n430 185
R1606 vdd.n609 vdd.n608 185
R1607 vdd.n607 vdd.n606 185
R1608 vdd.n605 vdd.n604 185
R1609 vdd.n603 vdd.n432 185
R1610 vdd.n599 vdd.n598 185
R1611 vdd.n597 vdd.n596 185
R1612 vdd.n595 vdd.n594 185
R1613 vdd.n593 vdd.n434 185
R1614 vdd.n589 vdd.n588 185
R1615 vdd.n587 vdd.n586 185
R1616 vdd.n585 vdd.n584 185
R1617 vdd.n583 vdd.n436 185
R1618 vdd.n579 vdd.n578 185
R1619 vdd.n577 vdd.n576 185
R1620 vdd.n575 vdd.n574 185
R1621 vdd.n573 vdd.n438 185
R1622 vdd.n569 vdd.n568 185
R1623 vdd.n567 vdd.n566 185
R1624 vdd.n565 vdd.n564 185
R1625 vdd.n563 vdd.n442 185
R1626 vdd.n559 vdd.n558 185
R1627 vdd.n557 vdd.n556 185
R1628 vdd.n555 vdd.n554 185
R1629 vdd.n553 vdd.n444 185
R1630 vdd.n549 vdd.n548 185
R1631 vdd.n547 vdd.n546 185
R1632 vdd.n545 vdd.n544 185
R1633 vdd.n543 vdd.n446 185
R1634 vdd.n539 vdd.n538 185
R1635 vdd.n537 vdd.n536 185
R1636 vdd.n535 vdd.n534 185
R1637 vdd.n533 vdd.n448 185
R1638 vdd.n529 vdd.n528 185
R1639 vdd.n527 vdd.n526 185
R1640 vdd.n525 vdd.n524 185
R1641 vdd.n523 vdd.n450 185
R1642 vdd.n519 vdd.n518 185
R1643 vdd.n517 vdd.n516 185
R1644 vdd.n515 vdd.n514 185
R1645 vdd.n513 vdd.n454 185
R1646 vdd.n509 vdd.n508 185
R1647 vdd.n507 vdd.n506 185
R1648 vdd.n505 vdd.n504 185
R1649 vdd.n503 vdd.n456 185
R1650 vdd.n499 vdd.n498 185
R1651 vdd.n497 vdd.n496 185
R1652 vdd.n495 vdd.n494 185
R1653 vdd.n493 vdd.n458 185
R1654 vdd.n489 vdd.n488 185
R1655 vdd.n487 vdd.n486 185
R1656 vdd.n485 vdd.n484 185
R1657 vdd.n483 vdd.n460 185
R1658 vdd.n479 vdd.n478 185
R1659 vdd.n477 vdd.n476 185
R1660 vdd.n475 vdd.n474 185
R1661 vdd.n473 vdd.n462 185
R1662 vdd.n469 vdd.n468 185
R1663 vdd.n467 vdd.n466 185
R1664 vdd.n465 vdd.n392 185
R1665 vdd.n3440 vdd.n393 185
R1666 vdd.n3447 vdd.n393 185
R1667 vdd.n3439 vdd.n3438 185
R1668 vdd.n3438 vdd.n386 185
R1669 vdd.n3437 vdd.n385 185
R1670 vdd.n3453 vdd.n385 185
R1671 vdd.n621 vdd.n384 185
R1672 vdd.n3454 vdd.n384 185
R1673 vdd.n3433 vdd.n383 185
R1674 vdd.n3455 vdd.n383 185
R1675 vdd.n3432 vdd.n3431 185
R1676 vdd.n3431 vdd.n375 185
R1677 vdd.n3430 vdd.n374 185
R1678 vdd.n3461 vdd.n374 185
R1679 vdd.n623 vdd.n373 185
R1680 vdd.n3462 vdd.n373 185
R1681 vdd.n3426 vdd.n372 185
R1682 vdd.n3463 vdd.n372 185
R1683 vdd.n3425 vdd.n3424 185
R1684 vdd.n3424 vdd.n3423 185
R1685 vdd.n3422 vdd.n364 185
R1686 vdd.n3469 vdd.n364 185
R1687 vdd.n625 vdd.n363 185
R1688 vdd.n3470 vdd.n363 185
R1689 vdd.n3418 vdd.n362 185
R1690 vdd.n3471 vdd.n362 185
R1691 vdd.n3417 vdd.n3416 185
R1692 vdd.n3416 vdd.n361 185
R1693 vdd.n3415 vdd.n353 185
R1694 vdd.n3477 vdd.n353 185
R1695 vdd.n627 vdd.n352 185
R1696 vdd.n3478 vdd.n352 185
R1697 vdd.n3411 vdd.n351 185
R1698 vdd.n3479 vdd.n351 185
R1699 vdd.n3410 vdd.n3409 185
R1700 vdd.n3409 vdd.n344 185
R1701 vdd.n3408 vdd.n343 185
R1702 vdd.n3485 vdd.n343 185
R1703 vdd.n629 vdd.n342 185
R1704 vdd.n3486 vdd.n342 185
R1705 vdd.n3404 vdd.n341 185
R1706 vdd.n3487 vdd.n341 185
R1707 vdd.n3403 vdd.n3402 185
R1708 vdd.n3402 vdd.n340 185
R1709 vdd.n3401 vdd.n631 185
R1710 vdd.n3401 vdd.n3400 185
R1711 vdd.n3389 vdd.n632 185
R1712 vdd.n633 vdd.n632 185
R1713 vdd.n3391 vdd.n3390 185
R1714 vdd.n3392 vdd.n3391 185
R1715 vdd.n640 vdd.n639 185
R1716 vdd.n644 vdd.n639 185
R1717 vdd.n3383 vdd.n3382 185
R1718 vdd.n3382 vdd.n3381 185
R1719 vdd.n643 vdd.n642 185
R1720 vdd.n3372 vdd.n643 185
R1721 vdd.n3371 vdd.n3370 185
R1722 vdd.n3373 vdd.n3371 185
R1723 vdd.n651 vdd.n650 185
R1724 vdd.n656 vdd.n650 185
R1725 vdd.n3366 vdd.n3365 185
R1726 vdd.n3365 vdd.n3364 185
R1727 vdd.n654 vdd.n653 185
R1728 vdd.n655 vdd.n654 185
R1729 vdd.n3355 vdd.n3354 185
R1730 vdd.n3356 vdd.n3355 185
R1731 vdd.n664 vdd.n663 185
R1732 vdd.n663 vdd.n662 185
R1733 vdd.n3350 vdd.n3349 185
R1734 vdd.n3349 vdd.n3348 185
R1735 vdd.n667 vdd.n666 185
R1736 vdd.n3339 vdd.n667 185
R1737 vdd.n3338 vdd.n3337 185
R1738 vdd.n3340 vdd.n3338 185
R1739 vdd.n674 vdd.n673 185
R1740 vdd.n679 vdd.n673 185
R1741 vdd.n3333 vdd.n3332 185
R1742 vdd.n3332 vdd.n3331 185
R1743 vdd.n677 vdd.n676 185
R1744 vdd.n678 vdd.n677 185
R1745 vdd.n3322 vdd.n3321 185
R1746 vdd.n3323 vdd.n3322 185
R1747 vdd.n686 vdd.n685 185
R1748 vdd.n723 vdd.n685 185
R1749 vdd.n2936 vdd.n2935 185
R1750 vdd.n2934 vdd.n2700 185
R1751 vdd.n2933 vdd.n2699 185
R1752 vdd.n2938 vdd.n2699 185
R1753 vdd.n2932 vdd.n2931 185
R1754 vdd.n2930 vdd.n2929 185
R1755 vdd.n2928 vdd.n2927 185
R1756 vdd.n2926 vdd.n2925 185
R1757 vdd.n2924 vdd.n2923 185
R1758 vdd.n2922 vdd.n2921 185
R1759 vdd.n2920 vdd.n2919 185
R1760 vdd.n2918 vdd.n2917 185
R1761 vdd.n2916 vdd.n2915 185
R1762 vdd.n2914 vdd.n2913 185
R1763 vdd.n2912 vdd.n2911 185
R1764 vdd.n2910 vdd.n2909 185
R1765 vdd.n2908 vdd.n2907 185
R1766 vdd.n2906 vdd.n2905 185
R1767 vdd.n2904 vdd.n2903 185
R1768 vdd.n2902 vdd.n2901 185
R1769 vdd.n2900 vdd.n2899 185
R1770 vdd.n2898 vdd.n2897 185
R1771 vdd.n2896 vdd.n2895 185
R1772 vdd.n2894 vdd.n2893 185
R1773 vdd.n2892 vdd.n2891 185
R1774 vdd.n2890 vdd.n2889 185
R1775 vdd.n2888 vdd.n2887 185
R1776 vdd.n2886 vdd.n2885 185
R1777 vdd.n2884 vdd.n2883 185
R1778 vdd.n2882 vdd.n2881 185
R1779 vdd.n2880 vdd.n2879 185
R1780 vdd.n2878 vdd.n2877 185
R1781 vdd.n2876 vdd.n2875 185
R1782 vdd.n2873 vdd.n2872 185
R1783 vdd.n2871 vdd.n2870 185
R1784 vdd.n2869 vdd.n2868 185
R1785 vdd.n3087 vdd.n3086 185
R1786 vdd.n3089 vdd.n834 185
R1787 vdd.n3091 vdd.n3090 185
R1788 vdd.n3093 vdd.n831 185
R1789 vdd.n3095 vdd.n3094 185
R1790 vdd.n3097 vdd.n829 185
R1791 vdd.n3099 vdd.n3098 185
R1792 vdd.n3100 vdd.n828 185
R1793 vdd.n3102 vdd.n3101 185
R1794 vdd.n3104 vdd.n826 185
R1795 vdd.n3106 vdd.n3105 185
R1796 vdd.n3107 vdd.n825 185
R1797 vdd.n3109 vdd.n3108 185
R1798 vdd.n3111 vdd.n823 185
R1799 vdd.n3113 vdd.n3112 185
R1800 vdd.n3114 vdd.n822 185
R1801 vdd.n3116 vdd.n3115 185
R1802 vdd.n3118 vdd.n731 185
R1803 vdd.n3120 vdd.n3119 185
R1804 vdd.n3122 vdd.n820 185
R1805 vdd.n3124 vdd.n3123 185
R1806 vdd.n3125 vdd.n819 185
R1807 vdd.n3127 vdd.n3126 185
R1808 vdd.n3129 vdd.n817 185
R1809 vdd.n3131 vdd.n3130 185
R1810 vdd.n3132 vdd.n816 185
R1811 vdd.n3134 vdd.n3133 185
R1812 vdd.n3136 vdd.n814 185
R1813 vdd.n3138 vdd.n3137 185
R1814 vdd.n3139 vdd.n813 185
R1815 vdd.n3141 vdd.n3140 185
R1816 vdd.n3143 vdd.n812 185
R1817 vdd.n3144 vdd.n811 185
R1818 vdd.n3147 vdd.n3146 185
R1819 vdd.n3148 vdd.n809 185
R1820 vdd.n809 vdd.n692 185
R1821 vdd.n3085 vdd.n806 185
R1822 vdd.n3151 vdd.n806 185
R1823 vdd.n3084 vdd.n3083 185
R1824 vdd.n3083 vdd.n805 185
R1825 vdd.n3082 vdd.n836 185
R1826 vdd.n3082 vdd.n3081 185
R1827 vdd.n2816 vdd.n837 185
R1828 vdd.n846 vdd.n837 185
R1829 vdd.n2817 vdd.n844 185
R1830 vdd.n3075 vdd.n844 185
R1831 vdd.n2819 vdd.n2818 185
R1832 vdd.n2818 vdd.n843 185
R1833 vdd.n2820 vdd.n852 185
R1834 vdd.n3024 vdd.n852 185
R1835 vdd.n2822 vdd.n2821 185
R1836 vdd.n2821 vdd.n851 185
R1837 vdd.n2823 vdd.n858 185
R1838 vdd.n3018 vdd.n858 185
R1839 vdd.n2825 vdd.n2824 185
R1840 vdd.n2824 vdd.n857 185
R1841 vdd.n2826 vdd.n863 185
R1842 vdd.n3012 vdd.n863 185
R1843 vdd.n2828 vdd.n2827 185
R1844 vdd.n2827 vdd.n870 185
R1845 vdd.n2829 vdd.n868 185
R1846 vdd.n3006 vdd.n868 185
R1847 vdd.n2831 vdd.n2830 185
R1848 vdd.n2830 vdd.n878 185
R1849 vdd.n2832 vdd.n876 185
R1850 vdd.n2999 vdd.n876 185
R1851 vdd.n2834 vdd.n2833 185
R1852 vdd.n2833 vdd.n875 185
R1853 vdd.n2835 vdd.n883 185
R1854 vdd.n2993 vdd.n883 185
R1855 vdd.n2837 vdd.n2836 185
R1856 vdd.n2836 vdd.n882 185
R1857 vdd.n2838 vdd.n888 185
R1858 vdd.n2987 vdd.n888 185
R1859 vdd.n2840 vdd.n2839 185
R1860 vdd.n2839 vdd.n895 185
R1861 vdd.n2841 vdd.n893 185
R1862 vdd.n2981 vdd.n893 185
R1863 vdd.n2843 vdd.n2842 185
R1864 vdd.n2842 vdd.n901 185
R1865 vdd.n2844 vdd.n899 185
R1866 vdd.n2975 vdd.n899 185
R1867 vdd.n2846 vdd.n2845 185
R1868 vdd.n2847 vdd.n2846 185
R1869 vdd.n2815 vdd.n906 185
R1870 vdd.n2969 vdd.n906 185
R1871 vdd.n2814 vdd.n2813 185
R1872 vdd.n2813 vdd.n905 185
R1873 vdd.n2812 vdd.n912 185
R1874 vdd.n2963 vdd.n912 185
R1875 vdd.n2811 vdd.n2810 185
R1876 vdd.n2810 vdd.n911 185
R1877 vdd.n2809 vdd.n918 185
R1878 vdd.n2957 vdd.n918 185
R1879 vdd.n2808 vdd.n2807 185
R1880 vdd.n2807 vdd.n917 185
R1881 vdd.n2703 vdd.n923 185
R1882 vdd.n2951 vdd.n923 185
R1883 vdd.n2864 vdd.n2863 185
R1884 vdd.n2863 vdd.n2862 185
R1885 vdd.n2865 vdd.n929 185
R1886 vdd.n2945 vdd.n929 185
R1887 vdd.n2867 vdd.n2866 185
R1888 vdd.n2867 vdd.n928 185
R1889 vdd.n927 vdd.n926 185
R1890 vdd.n928 vdd.n927 185
R1891 vdd.n2947 vdd.n2946 185
R1892 vdd.n2946 vdd.n2945 185
R1893 vdd.n2948 vdd.n925 185
R1894 vdd.n2862 vdd.n925 185
R1895 vdd.n2950 vdd.n2949 185
R1896 vdd.n2951 vdd.n2950 185
R1897 vdd.n916 vdd.n915 185
R1898 vdd.n917 vdd.n916 185
R1899 vdd.n2959 vdd.n2958 185
R1900 vdd.n2958 vdd.n2957 185
R1901 vdd.n2960 vdd.n914 185
R1902 vdd.n914 vdd.n911 185
R1903 vdd.n2962 vdd.n2961 185
R1904 vdd.n2963 vdd.n2962 185
R1905 vdd.n904 vdd.n903 185
R1906 vdd.n905 vdd.n904 185
R1907 vdd.n2971 vdd.n2970 185
R1908 vdd.n2970 vdd.n2969 185
R1909 vdd.n2972 vdd.n902 185
R1910 vdd.n2847 vdd.n902 185
R1911 vdd.n2974 vdd.n2973 185
R1912 vdd.n2975 vdd.n2974 185
R1913 vdd.n892 vdd.n891 185
R1914 vdd.n901 vdd.n892 185
R1915 vdd.n2983 vdd.n2982 185
R1916 vdd.n2982 vdd.n2981 185
R1917 vdd.n2984 vdd.n890 185
R1918 vdd.n895 vdd.n890 185
R1919 vdd.n2986 vdd.n2985 185
R1920 vdd.n2987 vdd.n2986 185
R1921 vdd.n881 vdd.n880 185
R1922 vdd.n882 vdd.n881 185
R1923 vdd.n2995 vdd.n2994 185
R1924 vdd.n2994 vdd.n2993 185
R1925 vdd.n2996 vdd.n879 185
R1926 vdd.n879 vdd.n875 185
R1927 vdd.n2998 vdd.n2997 185
R1928 vdd.n2999 vdd.n2998 185
R1929 vdd.n867 vdd.n866 185
R1930 vdd.n878 vdd.n867 185
R1931 vdd.n3008 vdd.n3007 185
R1932 vdd.n3007 vdd.n3006 185
R1933 vdd.n3009 vdd.n865 185
R1934 vdd.n870 vdd.n865 185
R1935 vdd.n3011 vdd.n3010 185
R1936 vdd.n3012 vdd.n3011 185
R1937 vdd.n856 vdd.n855 185
R1938 vdd.n857 vdd.n856 185
R1939 vdd.n3020 vdd.n3019 185
R1940 vdd.n3019 vdd.n3018 185
R1941 vdd.n3021 vdd.n854 185
R1942 vdd.n854 vdd.n851 185
R1943 vdd.n3023 vdd.n3022 185
R1944 vdd.n3024 vdd.n3023 185
R1945 vdd.n842 vdd.n841 185
R1946 vdd.n843 vdd.n842 185
R1947 vdd.n3077 vdd.n3076 185
R1948 vdd.n3076 vdd.n3075 185
R1949 vdd.n3078 vdd.n840 185
R1950 vdd.n846 vdd.n840 185
R1951 vdd.n3080 vdd.n3079 185
R1952 vdd.n3081 vdd.n3080 185
R1953 vdd.n810 vdd.n808 185
R1954 vdd.n808 vdd.n805 185
R1955 vdd.n3150 vdd.n3149 185
R1956 vdd.n3151 vdd.n3150 185
R1957 vdd.n2592 vdd.n2591 185
R1958 vdd.n2593 vdd.n2592 185
R1959 vdd.n980 vdd.n978 185
R1960 vdd.n978 vdd.n976 185
R1961 vdd.n2507 vdd.n987 185
R1962 vdd.n2518 vdd.n987 185
R1963 vdd.n2508 vdd.n996 185
R1964 vdd.n1338 vdd.n996 185
R1965 vdd.n2510 vdd.n2509 185
R1966 vdd.n2511 vdd.n2510 185
R1967 vdd.n2506 vdd.n995 185
R1968 vdd.n995 vdd.n992 185
R1969 vdd.n2505 vdd.n2504 185
R1970 vdd.n2504 vdd.n2503 185
R1971 vdd.n998 vdd.n997 185
R1972 vdd.n999 vdd.n998 185
R1973 vdd.n2496 vdd.n2495 185
R1974 vdd.n2497 vdd.n2496 185
R1975 vdd.n2494 vdd.n1008 185
R1976 vdd.n1008 vdd.n1005 185
R1977 vdd.n2493 vdd.n2492 185
R1978 vdd.n2492 vdd.n2491 185
R1979 vdd.n1010 vdd.n1009 185
R1980 vdd.n1018 vdd.n1010 185
R1981 vdd.n2484 vdd.n2483 185
R1982 vdd.n2485 vdd.n2484 185
R1983 vdd.n2482 vdd.n1019 185
R1984 vdd.n1024 vdd.n1019 185
R1985 vdd.n2481 vdd.n2480 185
R1986 vdd.n2480 vdd.n2479 185
R1987 vdd.n1021 vdd.n1020 185
R1988 vdd.n1359 vdd.n1021 185
R1989 vdd.n2472 vdd.n2471 185
R1990 vdd.n2473 vdd.n2472 185
R1991 vdd.n2470 vdd.n1031 185
R1992 vdd.n1031 vdd.n1028 185
R1993 vdd.n2469 vdd.n2468 185
R1994 vdd.n2468 vdd.n2467 185
R1995 vdd.n1033 vdd.n1032 185
R1996 vdd.n1034 vdd.n1033 185
R1997 vdd.n2460 vdd.n2459 185
R1998 vdd.n2461 vdd.n2460 185
R1999 vdd.n2457 vdd.n1042 185
R2000 vdd.n1048 vdd.n1042 185
R2001 vdd.n2456 vdd.n2455 185
R2002 vdd.n2455 vdd.n2454 185
R2003 vdd.n1045 vdd.n1044 185
R2004 vdd.n1055 vdd.n1045 185
R2005 vdd.n2447 vdd.n2446 185
R2006 vdd.n2448 vdd.n2447 185
R2007 vdd.n2445 vdd.n1056 185
R2008 vdd.n1056 vdd.n1052 185
R2009 vdd.n2444 vdd.n2443 185
R2010 vdd.n2443 vdd.n2442 185
R2011 vdd.n1058 vdd.n1057 185
R2012 vdd.n1059 vdd.n1058 185
R2013 vdd.n2435 vdd.n2434 185
R2014 vdd.n2436 vdd.n2435 185
R2015 vdd.n2433 vdd.n1068 185
R2016 vdd.n1068 vdd.n1065 185
R2017 vdd.n2432 vdd.n2431 185
R2018 vdd.n2431 vdd.n2430 185
R2019 vdd.n1070 vdd.n1069 185
R2020 vdd.n1079 vdd.n1070 185
R2021 vdd.n2423 vdd.n2422 185
R2022 vdd.n2424 vdd.n2423 185
R2023 vdd.n2421 vdd.n1080 185
R2024 vdd.n1080 vdd.n1076 185
R2025 vdd.n2523 vdd.n951 185
R2026 vdd.n2665 vdd.n951 185
R2027 vdd.n2525 vdd.n2524 185
R2028 vdd.n2527 vdd.n2526 185
R2029 vdd.n2529 vdd.n2528 185
R2030 vdd.n2531 vdd.n2530 185
R2031 vdd.n2533 vdd.n2532 185
R2032 vdd.n2535 vdd.n2534 185
R2033 vdd.n2537 vdd.n2536 185
R2034 vdd.n2539 vdd.n2538 185
R2035 vdd.n2541 vdd.n2540 185
R2036 vdd.n2543 vdd.n2542 185
R2037 vdd.n2545 vdd.n2544 185
R2038 vdd.n2547 vdd.n2546 185
R2039 vdd.n2549 vdd.n2548 185
R2040 vdd.n2551 vdd.n2550 185
R2041 vdd.n2553 vdd.n2552 185
R2042 vdd.n2555 vdd.n2554 185
R2043 vdd.n2557 vdd.n2556 185
R2044 vdd.n2559 vdd.n2558 185
R2045 vdd.n2561 vdd.n2560 185
R2046 vdd.n2563 vdd.n2562 185
R2047 vdd.n2565 vdd.n2564 185
R2048 vdd.n2567 vdd.n2566 185
R2049 vdd.n2569 vdd.n2568 185
R2050 vdd.n2571 vdd.n2570 185
R2051 vdd.n2573 vdd.n2572 185
R2052 vdd.n2575 vdd.n2574 185
R2053 vdd.n2577 vdd.n2576 185
R2054 vdd.n2579 vdd.n2578 185
R2055 vdd.n2581 vdd.n2580 185
R2056 vdd.n2583 vdd.n2582 185
R2057 vdd.n2585 vdd.n2584 185
R2058 vdd.n2587 vdd.n2586 185
R2059 vdd.n2589 vdd.n2588 185
R2060 vdd.n2590 vdd.n979 185
R2061 vdd.n2522 vdd.n977 185
R2062 vdd.n2593 vdd.n977 185
R2063 vdd.n2521 vdd.n2520 185
R2064 vdd.n2520 vdd.n976 185
R2065 vdd.n2519 vdd.n984 185
R2066 vdd.n2519 vdd.n2518 185
R2067 vdd.n1256 vdd.n985 185
R2068 vdd.n1338 vdd.n985 185
R2069 vdd.n1257 vdd.n994 185
R2070 vdd.n2511 vdd.n994 185
R2071 vdd.n1259 vdd.n1258 185
R2072 vdd.n1258 vdd.n992 185
R2073 vdd.n1260 vdd.n1001 185
R2074 vdd.n2503 vdd.n1001 185
R2075 vdd.n1262 vdd.n1261 185
R2076 vdd.n1261 vdd.n999 185
R2077 vdd.n1263 vdd.n1007 185
R2078 vdd.n2497 vdd.n1007 185
R2079 vdd.n1265 vdd.n1264 185
R2080 vdd.n1264 vdd.n1005 185
R2081 vdd.n1266 vdd.n1012 185
R2082 vdd.n2491 vdd.n1012 185
R2083 vdd.n1268 vdd.n1267 185
R2084 vdd.n1267 vdd.n1018 185
R2085 vdd.n1269 vdd.n1017 185
R2086 vdd.n2485 vdd.n1017 185
R2087 vdd.n1271 vdd.n1270 185
R2088 vdd.n1270 vdd.n1024 185
R2089 vdd.n1272 vdd.n1023 185
R2090 vdd.n2479 vdd.n1023 185
R2091 vdd.n1361 vdd.n1360 185
R2092 vdd.n1360 vdd.n1359 185
R2093 vdd.n1362 vdd.n1030 185
R2094 vdd.n2473 vdd.n1030 185
R2095 vdd.n1364 vdd.n1363 185
R2096 vdd.n1363 vdd.n1028 185
R2097 vdd.n1365 vdd.n1036 185
R2098 vdd.n2467 vdd.n1036 185
R2099 vdd.n1367 vdd.n1366 185
R2100 vdd.n1366 vdd.n1034 185
R2101 vdd.n1368 vdd.n1041 185
R2102 vdd.n2461 vdd.n1041 185
R2103 vdd.n1370 vdd.n1369 185
R2104 vdd.n1369 vdd.n1048 185
R2105 vdd.n1371 vdd.n1047 185
R2106 vdd.n2454 vdd.n1047 185
R2107 vdd.n1373 vdd.n1372 185
R2108 vdd.n1372 vdd.n1055 185
R2109 vdd.n1374 vdd.n1054 185
R2110 vdd.n2448 vdd.n1054 185
R2111 vdd.n1376 vdd.n1375 185
R2112 vdd.n1375 vdd.n1052 185
R2113 vdd.n1377 vdd.n1061 185
R2114 vdd.n2442 vdd.n1061 185
R2115 vdd.n1379 vdd.n1378 185
R2116 vdd.n1378 vdd.n1059 185
R2117 vdd.n1380 vdd.n1067 185
R2118 vdd.n2436 vdd.n1067 185
R2119 vdd.n1382 vdd.n1381 185
R2120 vdd.n1381 vdd.n1065 185
R2121 vdd.n1383 vdd.n1072 185
R2122 vdd.n2430 vdd.n1072 185
R2123 vdd.n1385 vdd.n1384 185
R2124 vdd.n1384 vdd.n1079 185
R2125 vdd.n1386 vdd.n1078 185
R2126 vdd.n2424 vdd.n1078 185
R2127 vdd.n1388 vdd.n1387 185
R2128 vdd.n1387 vdd.n1076 185
R2129 vdd.n2420 vdd.n2419 185
R2130 vdd.n1082 vdd.n1081 185
R2131 vdd.n1223 vdd.n1222 185
R2132 vdd.n1225 vdd.n1224 185
R2133 vdd.n1227 vdd.n1226 185
R2134 vdd.n1229 vdd.n1228 185
R2135 vdd.n1231 vdd.n1230 185
R2136 vdd.n1233 vdd.n1232 185
R2137 vdd.n1235 vdd.n1234 185
R2138 vdd.n1237 vdd.n1236 185
R2139 vdd.n1239 vdd.n1238 185
R2140 vdd.n1241 vdd.n1240 185
R2141 vdd.n1243 vdd.n1242 185
R2142 vdd.n1245 vdd.n1244 185
R2143 vdd.n1247 vdd.n1246 185
R2144 vdd.n1249 vdd.n1248 185
R2145 vdd.n1251 vdd.n1250 185
R2146 vdd.n1422 vdd.n1252 185
R2147 vdd.n1421 vdd.n1420 185
R2148 vdd.n1419 vdd.n1418 185
R2149 vdd.n1417 vdd.n1416 185
R2150 vdd.n1415 vdd.n1414 185
R2151 vdd.n1413 vdd.n1412 185
R2152 vdd.n1411 vdd.n1410 185
R2153 vdd.n1409 vdd.n1408 185
R2154 vdd.n1407 vdd.n1406 185
R2155 vdd.n1405 vdd.n1404 185
R2156 vdd.n1403 vdd.n1402 185
R2157 vdd.n1401 vdd.n1400 185
R2158 vdd.n1399 vdd.n1398 185
R2159 vdd.n1397 vdd.n1396 185
R2160 vdd.n1395 vdd.n1394 185
R2161 vdd.n1393 vdd.n1392 185
R2162 vdd.n1391 vdd.n1390 185
R2163 vdd.n1389 vdd.n1116 185
R2164 vdd.n2417 vdd.n1116 185
R2165 vdd.n2417 vdd.n1083 179.345
R2166 vdd.n3315 vdd.n692 179.345
R2167 vdd.n327 vdd.n326 171.744
R2168 vdd.n326 vdd.n325 171.744
R2169 vdd.n325 vdd.n294 171.744
R2170 vdd.n318 vdd.n294 171.744
R2171 vdd.n318 vdd.n317 171.744
R2172 vdd.n317 vdd.n299 171.744
R2173 vdd.n310 vdd.n299 171.744
R2174 vdd.n310 vdd.n309 171.744
R2175 vdd.n309 vdd.n303 171.744
R2176 vdd.n268 vdd.n267 171.744
R2177 vdd.n267 vdd.n266 171.744
R2178 vdd.n266 vdd.n235 171.744
R2179 vdd.n259 vdd.n235 171.744
R2180 vdd.n259 vdd.n258 171.744
R2181 vdd.n258 vdd.n240 171.744
R2182 vdd.n251 vdd.n240 171.744
R2183 vdd.n251 vdd.n250 171.744
R2184 vdd.n250 vdd.n244 171.744
R2185 vdd.n225 vdd.n224 171.744
R2186 vdd.n224 vdd.n223 171.744
R2187 vdd.n223 vdd.n192 171.744
R2188 vdd.n216 vdd.n192 171.744
R2189 vdd.n216 vdd.n215 171.744
R2190 vdd.n215 vdd.n197 171.744
R2191 vdd.n208 vdd.n197 171.744
R2192 vdd.n208 vdd.n207 171.744
R2193 vdd.n207 vdd.n201 171.744
R2194 vdd.n166 vdd.n165 171.744
R2195 vdd.n165 vdd.n164 171.744
R2196 vdd.n164 vdd.n133 171.744
R2197 vdd.n157 vdd.n133 171.744
R2198 vdd.n157 vdd.n156 171.744
R2199 vdd.n156 vdd.n138 171.744
R2200 vdd.n149 vdd.n138 171.744
R2201 vdd.n149 vdd.n148 171.744
R2202 vdd.n148 vdd.n142 171.744
R2203 vdd.n124 vdd.n123 171.744
R2204 vdd.n123 vdd.n122 171.744
R2205 vdd.n122 vdd.n91 171.744
R2206 vdd.n115 vdd.n91 171.744
R2207 vdd.n115 vdd.n114 171.744
R2208 vdd.n114 vdd.n96 171.744
R2209 vdd.n107 vdd.n96 171.744
R2210 vdd.n107 vdd.n106 171.744
R2211 vdd.n106 vdd.n100 171.744
R2212 vdd.n65 vdd.n64 171.744
R2213 vdd.n64 vdd.n63 171.744
R2214 vdd.n63 vdd.n32 171.744
R2215 vdd.n56 vdd.n32 171.744
R2216 vdd.n56 vdd.n55 171.744
R2217 vdd.n55 vdd.n37 171.744
R2218 vdd.n48 vdd.n37 171.744
R2219 vdd.n48 vdd.n47 171.744
R2220 vdd.n47 vdd.n41 171.744
R2221 vdd.n2108 vdd.n2107 171.744
R2222 vdd.n2107 vdd.n2106 171.744
R2223 vdd.n2106 vdd.n2075 171.744
R2224 vdd.n2099 vdd.n2075 171.744
R2225 vdd.n2099 vdd.n2098 171.744
R2226 vdd.n2098 vdd.n2080 171.744
R2227 vdd.n2091 vdd.n2080 171.744
R2228 vdd.n2091 vdd.n2090 171.744
R2229 vdd.n2090 vdd.n2084 171.744
R2230 vdd.n2167 vdd.n2166 171.744
R2231 vdd.n2166 vdd.n2165 171.744
R2232 vdd.n2165 vdd.n2134 171.744
R2233 vdd.n2158 vdd.n2134 171.744
R2234 vdd.n2158 vdd.n2157 171.744
R2235 vdd.n2157 vdd.n2139 171.744
R2236 vdd.n2150 vdd.n2139 171.744
R2237 vdd.n2150 vdd.n2149 171.744
R2238 vdd.n2149 vdd.n2143 171.744
R2239 vdd.n2006 vdd.n2005 171.744
R2240 vdd.n2005 vdd.n2004 171.744
R2241 vdd.n2004 vdd.n1973 171.744
R2242 vdd.n1997 vdd.n1973 171.744
R2243 vdd.n1997 vdd.n1996 171.744
R2244 vdd.n1996 vdd.n1978 171.744
R2245 vdd.n1989 vdd.n1978 171.744
R2246 vdd.n1989 vdd.n1988 171.744
R2247 vdd.n1988 vdd.n1982 171.744
R2248 vdd.n2065 vdd.n2064 171.744
R2249 vdd.n2064 vdd.n2063 171.744
R2250 vdd.n2063 vdd.n2032 171.744
R2251 vdd.n2056 vdd.n2032 171.744
R2252 vdd.n2056 vdd.n2055 171.744
R2253 vdd.n2055 vdd.n2037 171.744
R2254 vdd.n2048 vdd.n2037 171.744
R2255 vdd.n2048 vdd.n2047 171.744
R2256 vdd.n2047 vdd.n2041 171.744
R2257 vdd.n1905 vdd.n1904 171.744
R2258 vdd.n1904 vdd.n1903 171.744
R2259 vdd.n1903 vdd.n1872 171.744
R2260 vdd.n1896 vdd.n1872 171.744
R2261 vdd.n1896 vdd.n1895 171.744
R2262 vdd.n1895 vdd.n1877 171.744
R2263 vdd.n1888 vdd.n1877 171.744
R2264 vdd.n1888 vdd.n1887 171.744
R2265 vdd.n1887 vdd.n1881 171.744
R2266 vdd.n1964 vdd.n1963 171.744
R2267 vdd.n1963 vdd.n1962 171.744
R2268 vdd.n1962 vdd.n1931 171.744
R2269 vdd.n1955 vdd.n1931 171.744
R2270 vdd.n1955 vdd.n1954 171.744
R2271 vdd.n1954 vdd.n1936 171.744
R2272 vdd.n1947 vdd.n1936 171.744
R2273 vdd.n1947 vdd.n1946 171.744
R2274 vdd.n1946 vdd.n1940 171.744
R2275 vdd.n468 vdd.n467 146.341
R2276 vdd.n474 vdd.n473 146.341
R2277 vdd.n478 vdd.n477 146.341
R2278 vdd.n484 vdd.n483 146.341
R2279 vdd.n488 vdd.n487 146.341
R2280 vdd.n494 vdd.n493 146.341
R2281 vdd.n498 vdd.n497 146.341
R2282 vdd.n504 vdd.n503 146.341
R2283 vdd.n508 vdd.n507 146.341
R2284 vdd.n514 vdd.n513 146.341
R2285 vdd.n518 vdd.n517 146.341
R2286 vdd.n524 vdd.n523 146.341
R2287 vdd.n528 vdd.n527 146.341
R2288 vdd.n534 vdd.n533 146.341
R2289 vdd.n538 vdd.n537 146.341
R2290 vdd.n544 vdd.n543 146.341
R2291 vdd.n548 vdd.n547 146.341
R2292 vdd.n554 vdd.n553 146.341
R2293 vdd.n558 vdd.n557 146.341
R2294 vdd.n564 vdd.n563 146.341
R2295 vdd.n568 vdd.n567 146.341
R2296 vdd.n574 vdd.n573 146.341
R2297 vdd.n578 vdd.n577 146.341
R2298 vdd.n584 vdd.n583 146.341
R2299 vdd.n588 vdd.n587 146.341
R2300 vdd.n594 vdd.n593 146.341
R2301 vdd.n598 vdd.n597 146.341
R2302 vdd.n604 vdd.n603 146.341
R2303 vdd.n608 vdd.n607 146.341
R2304 vdd.n614 vdd.n613 146.341
R2305 vdd.n616 vdd.n425 146.341
R2306 vdd.n3322 vdd.n685 146.341
R2307 vdd.n3322 vdd.n677 146.341
R2308 vdd.n3332 vdd.n677 146.341
R2309 vdd.n3332 vdd.n673 146.341
R2310 vdd.n3338 vdd.n673 146.341
R2311 vdd.n3338 vdd.n667 146.341
R2312 vdd.n3349 vdd.n667 146.341
R2313 vdd.n3349 vdd.n663 146.341
R2314 vdd.n3355 vdd.n663 146.341
R2315 vdd.n3355 vdd.n654 146.341
R2316 vdd.n3365 vdd.n654 146.341
R2317 vdd.n3365 vdd.n650 146.341
R2318 vdd.n3371 vdd.n650 146.341
R2319 vdd.n3371 vdd.n643 146.341
R2320 vdd.n3382 vdd.n643 146.341
R2321 vdd.n3382 vdd.n639 146.341
R2322 vdd.n3391 vdd.n639 146.341
R2323 vdd.n3391 vdd.n632 146.341
R2324 vdd.n3401 vdd.n632 146.341
R2325 vdd.n3402 vdd.n3401 146.341
R2326 vdd.n3402 vdd.n341 146.341
R2327 vdd.n342 vdd.n341 146.341
R2328 vdd.n343 vdd.n342 146.341
R2329 vdd.n3409 vdd.n343 146.341
R2330 vdd.n3409 vdd.n351 146.341
R2331 vdd.n352 vdd.n351 146.341
R2332 vdd.n353 vdd.n352 146.341
R2333 vdd.n3416 vdd.n353 146.341
R2334 vdd.n3416 vdd.n362 146.341
R2335 vdd.n363 vdd.n362 146.341
R2336 vdd.n364 vdd.n363 146.341
R2337 vdd.n3424 vdd.n364 146.341
R2338 vdd.n3424 vdd.n372 146.341
R2339 vdd.n373 vdd.n372 146.341
R2340 vdd.n374 vdd.n373 146.341
R2341 vdd.n3431 vdd.n374 146.341
R2342 vdd.n3431 vdd.n383 146.341
R2343 vdd.n384 vdd.n383 146.341
R2344 vdd.n385 vdd.n384 146.341
R2345 vdd.n3438 vdd.n385 146.341
R2346 vdd.n3438 vdd.n393 146.341
R2347 vdd.n725 vdd.n724 146.341
R2348 vdd.n728 vdd.n724 146.341
R2349 vdd.n734 vdd.n733 146.341
R2350 vdd.n3304 vdd.n3303 146.341
R2351 vdd.n3300 vdd.n3299 146.341
R2352 vdd.n3296 vdd.n3295 146.341
R2353 vdd.n3292 vdd.n3291 146.341
R2354 vdd.n3288 vdd.n3287 146.341
R2355 vdd.n3284 vdd.n3283 146.341
R2356 vdd.n3280 vdd.n3279 146.341
R2357 vdd.n3271 vdd.n3270 146.341
R2358 vdd.n3268 vdd.n3267 146.341
R2359 vdd.n3264 vdd.n3263 146.341
R2360 vdd.n3260 vdd.n3259 146.341
R2361 vdd.n3256 vdd.n3255 146.341
R2362 vdd.n3252 vdd.n3251 146.341
R2363 vdd.n3248 vdd.n3247 146.341
R2364 vdd.n3244 vdd.n3243 146.341
R2365 vdd.n3240 vdd.n3239 146.341
R2366 vdd.n3236 vdd.n3235 146.341
R2367 vdd.n3232 vdd.n3231 146.341
R2368 vdd.n3225 vdd.n3224 146.341
R2369 vdd.n3222 vdd.n3221 146.341
R2370 vdd.n3218 vdd.n3217 146.341
R2371 vdd.n3214 vdd.n3213 146.341
R2372 vdd.n3210 vdd.n3209 146.341
R2373 vdd.n3206 vdd.n3205 146.341
R2374 vdd.n3202 vdd.n3201 146.341
R2375 vdd.n3198 vdd.n3197 146.341
R2376 vdd.n3194 vdd.n3193 146.341
R2377 vdd.n3190 vdd.n3189 146.341
R2378 vdd.n3316 vdd.n691 146.341
R2379 vdd.n3324 vdd.n684 146.341
R2380 vdd.n3324 vdd.n680 146.341
R2381 vdd.n3330 vdd.n680 146.341
R2382 vdd.n3330 vdd.n672 146.341
R2383 vdd.n3341 vdd.n672 146.341
R2384 vdd.n3341 vdd.n668 146.341
R2385 vdd.n3347 vdd.n668 146.341
R2386 vdd.n3347 vdd.n661 146.341
R2387 vdd.n3357 vdd.n661 146.341
R2388 vdd.n3357 vdd.n657 146.341
R2389 vdd.n3363 vdd.n657 146.341
R2390 vdd.n3363 vdd.n649 146.341
R2391 vdd.n3374 vdd.n649 146.341
R2392 vdd.n3374 vdd.n645 146.341
R2393 vdd.n3380 vdd.n645 146.341
R2394 vdd.n3380 vdd.n638 146.341
R2395 vdd.n3393 vdd.n638 146.341
R2396 vdd.n3393 vdd.n634 146.341
R2397 vdd.n3399 vdd.n634 146.341
R2398 vdd.n3399 vdd.n338 146.341
R2399 vdd.n3488 vdd.n338 146.341
R2400 vdd.n3488 vdd.n339 146.341
R2401 vdd.n3484 vdd.n339 146.341
R2402 vdd.n3484 vdd.n345 146.341
R2403 vdd.n3480 vdd.n345 146.341
R2404 vdd.n3480 vdd.n350 146.341
R2405 vdd.n3476 vdd.n350 146.341
R2406 vdd.n3476 vdd.n354 146.341
R2407 vdd.n3472 vdd.n354 146.341
R2408 vdd.n3472 vdd.n360 146.341
R2409 vdd.n3468 vdd.n360 146.341
R2410 vdd.n3468 vdd.n365 146.341
R2411 vdd.n3464 vdd.n365 146.341
R2412 vdd.n3464 vdd.n371 146.341
R2413 vdd.n3460 vdd.n371 146.341
R2414 vdd.n3460 vdd.n376 146.341
R2415 vdd.n3456 vdd.n376 146.341
R2416 vdd.n3456 vdd.n382 146.341
R2417 vdd.n3452 vdd.n382 146.341
R2418 vdd.n3452 vdd.n387 146.341
R2419 vdd.n3448 vdd.n387 146.341
R2420 vdd.n2378 vdd.n2377 146.341
R2421 vdd.n2375 vdd.n2372 146.341
R2422 vdd.n2370 vdd.n1127 146.341
R2423 vdd.n2366 vdd.n2365 146.341
R2424 vdd.n2363 vdd.n1131 146.341
R2425 vdd.n2359 vdd.n2358 146.341
R2426 vdd.n2356 vdd.n1138 146.341
R2427 vdd.n2352 vdd.n2351 146.341
R2428 vdd.n2349 vdd.n1145 146.341
R2429 vdd.n1156 vdd.n1153 146.341
R2430 vdd.n2341 vdd.n2340 146.341
R2431 vdd.n2338 vdd.n1158 146.341
R2432 vdd.n2334 vdd.n2333 146.341
R2433 vdd.n2331 vdd.n1164 146.341
R2434 vdd.n2327 vdd.n2326 146.341
R2435 vdd.n2324 vdd.n1171 146.341
R2436 vdd.n2320 vdd.n2319 146.341
R2437 vdd.n2317 vdd.n1178 146.341
R2438 vdd.n2313 vdd.n2312 146.341
R2439 vdd.n2310 vdd.n1185 146.341
R2440 vdd.n1196 vdd.n1193 146.341
R2441 vdd.n2302 vdd.n2301 146.341
R2442 vdd.n2299 vdd.n1198 146.341
R2443 vdd.n2295 vdd.n2294 146.341
R2444 vdd.n2292 vdd.n1204 146.341
R2445 vdd.n2288 vdd.n2287 146.341
R2446 vdd.n2285 vdd.n1211 146.341
R2447 vdd.n2281 vdd.n2280 146.341
R2448 vdd.n2278 vdd.n1218 146.341
R2449 vdd.n1429 vdd.n1427 146.341
R2450 vdd.n1432 vdd.n1431 146.341
R2451 vdd.n1790 vdd.n1550 146.341
R2452 vdd.n1790 vdd.n1546 146.341
R2453 vdd.n1796 vdd.n1546 146.341
R2454 vdd.n1796 vdd.n1538 146.341
R2455 vdd.n1807 vdd.n1538 146.341
R2456 vdd.n1807 vdd.n1534 146.341
R2457 vdd.n1813 vdd.n1534 146.341
R2458 vdd.n1813 vdd.n1528 146.341
R2459 vdd.n1824 vdd.n1528 146.341
R2460 vdd.n1824 vdd.n1524 146.341
R2461 vdd.n1830 vdd.n1524 146.341
R2462 vdd.n1830 vdd.n1515 146.341
R2463 vdd.n1840 vdd.n1515 146.341
R2464 vdd.n1840 vdd.n1511 146.341
R2465 vdd.n1846 vdd.n1511 146.341
R2466 vdd.n1846 vdd.n1504 146.341
R2467 vdd.n1857 vdd.n1504 146.341
R2468 vdd.n1857 vdd.n1500 146.341
R2469 vdd.n1863 vdd.n1500 146.341
R2470 vdd.n1863 vdd.n1493 146.341
R2471 vdd.n2180 vdd.n1493 146.341
R2472 vdd.n2180 vdd.n1489 146.341
R2473 vdd.n2186 vdd.n1489 146.341
R2474 vdd.n2186 vdd.n1481 146.341
R2475 vdd.n2197 vdd.n1481 146.341
R2476 vdd.n2197 vdd.n1477 146.341
R2477 vdd.n2203 vdd.n1477 146.341
R2478 vdd.n2203 vdd.n1471 146.341
R2479 vdd.n2214 vdd.n1471 146.341
R2480 vdd.n2214 vdd.n1467 146.341
R2481 vdd.n2220 vdd.n1467 146.341
R2482 vdd.n2220 vdd.n1458 146.341
R2483 vdd.n2230 vdd.n1458 146.341
R2484 vdd.n2230 vdd.n1454 146.341
R2485 vdd.n2236 vdd.n1454 146.341
R2486 vdd.n2236 vdd.n1448 146.341
R2487 vdd.n2247 vdd.n1448 146.341
R2488 vdd.n2247 vdd.n1443 146.341
R2489 vdd.n2255 vdd.n1443 146.341
R2490 vdd.n2255 vdd.n1434 146.341
R2491 vdd.n2266 vdd.n1434 146.341
R2492 vdd.n1779 vdd.n1555 146.341
R2493 vdd.n1779 vdd.n1588 146.341
R2494 vdd.n1592 vdd.n1591 146.341
R2495 vdd.n1594 vdd.n1593 146.341
R2496 vdd.n1598 vdd.n1597 146.341
R2497 vdd.n1600 vdd.n1599 146.341
R2498 vdd.n1604 vdd.n1603 146.341
R2499 vdd.n1606 vdd.n1605 146.341
R2500 vdd.n1610 vdd.n1609 146.341
R2501 vdd.n1612 vdd.n1611 146.341
R2502 vdd.n1618 vdd.n1617 146.341
R2503 vdd.n1620 vdd.n1619 146.341
R2504 vdd.n1624 vdd.n1623 146.341
R2505 vdd.n1626 vdd.n1625 146.341
R2506 vdd.n1630 vdd.n1629 146.341
R2507 vdd.n1632 vdd.n1631 146.341
R2508 vdd.n1636 vdd.n1635 146.341
R2509 vdd.n1638 vdd.n1637 146.341
R2510 vdd.n1642 vdd.n1641 146.341
R2511 vdd.n1644 vdd.n1643 146.341
R2512 vdd.n1716 vdd.n1647 146.341
R2513 vdd.n1649 vdd.n1648 146.341
R2514 vdd.n1653 vdd.n1652 146.341
R2515 vdd.n1655 vdd.n1654 146.341
R2516 vdd.n1659 vdd.n1658 146.341
R2517 vdd.n1661 vdd.n1660 146.341
R2518 vdd.n1665 vdd.n1664 146.341
R2519 vdd.n1667 vdd.n1666 146.341
R2520 vdd.n1671 vdd.n1670 146.341
R2521 vdd.n1673 vdd.n1672 146.341
R2522 vdd.n1677 vdd.n1676 146.341
R2523 vdd.n1678 vdd.n1586 146.341
R2524 vdd.n1788 vdd.n1551 146.341
R2525 vdd.n1788 vdd.n1544 146.341
R2526 vdd.n1799 vdd.n1544 146.341
R2527 vdd.n1799 vdd.n1540 146.341
R2528 vdd.n1805 vdd.n1540 146.341
R2529 vdd.n1805 vdd.n1533 146.341
R2530 vdd.n1816 vdd.n1533 146.341
R2531 vdd.n1816 vdd.n1529 146.341
R2532 vdd.n1822 vdd.n1529 146.341
R2533 vdd.n1822 vdd.n1522 146.341
R2534 vdd.n1832 vdd.n1522 146.341
R2535 vdd.n1832 vdd.n1518 146.341
R2536 vdd.n1838 vdd.n1518 146.341
R2537 vdd.n1838 vdd.n1510 146.341
R2538 vdd.n1849 vdd.n1510 146.341
R2539 vdd.n1849 vdd.n1506 146.341
R2540 vdd.n1855 vdd.n1506 146.341
R2541 vdd.n1855 vdd.n1499 146.341
R2542 vdd.n1865 vdd.n1499 146.341
R2543 vdd.n1865 vdd.n1495 146.341
R2544 vdd.n2178 vdd.n1495 146.341
R2545 vdd.n2178 vdd.n1487 146.341
R2546 vdd.n2189 vdd.n1487 146.341
R2547 vdd.n2189 vdd.n1483 146.341
R2548 vdd.n2195 vdd.n1483 146.341
R2549 vdd.n2195 vdd.n1476 146.341
R2550 vdd.n2206 vdd.n1476 146.341
R2551 vdd.n2206 vdd.n1472 146.341
R2552 vdd.n2212 vdd.n1472 146.341
R2553 vdd.n2212 vdd.n1465 146.341
R2554 vdd.n2222 vdd.n1465 146.341
R2555 vdd.n2222 vdd.n1461 146.341
R2556 vdd.n2228 vdd.n1461 146.341
R2557 vdd.n2228 vdd.n1453 146.341
R2558 vdd.n2239 vdd.n1453 146.341
R2559 vdd.n2239 vdd.n1449 146.341
R2560 vdd.n2245 vdd.n1449 146.341
R2561 vdd.n2245 vdd.n1441 146.341
R2562 vdd.n2258 vdd.n1441 146.341
R2563 vdd.n2258 vdd.n1436 146.341
R2564 vdd.n2264 vdd.n1436 146.341
R2565 vdd.n1253 vdd.t61 127.284
R2566 vdd.n981 vdd.t102 127.284
R2567 vdd.n1273 vdd.t75 127.284
R2568 vdd.n972 vdd.t125 127.284
R2569 vdd.n872 vdd.t82 127.284
R2570 vdd.n872 vdd.t83 127.284
R2571 vdd.n2704 vdd.t117 127.284
R2572 vdd.n832 vdd.t128 127.284
R2573 vdd.n2701 vdd.t107 127.284
R2574 vdd.n799 vdd.t56 127.284
R2575 vdd.n1043 vdd.t113 127.284
R2576 vdd.n1043 vdd.t114 127.284
R2577 vdd.n22 vdd.n20 117.314
R2578 vdd.n17 vdd.n15 117.314
R2579 vdd.n27 vdd.n26 116.927
R2580 vdd.n24 vdd.n23 116.927
R2581 vdd.n22 vdd.n21 116.927
R2582 vdd.n17 vdd.n16 116.927
R2583 vdd.n19 vdd.n18 116.927
R2584 vdd.n27 vdd.n25 116.927
R2585 vdd.n1254 vdd.t60 111.188
R2586 vdd.n982 vdd.t103 111.188
R2587 vdd.n1274 vdd.t74 111.188
R2588 vdd.n973 vdd.t126 111.188
R2589 vdd.n2705 vdd.t116 111.188
R2590 vdd.n833 vdd.t129 111.188
R2591 vdd.n2702 vdd.t106 111.188
R2592 vdd.n800 vdd.t57 111.188
R2593 vdd.n2946 vdd.n927 99.5127
R2594 vdd.n2946 vdd.n925 99.5127
R2595 vdd.n2950 vdd.n925 99.5127
R2596 vdd.n2950 vdd.n916 99.5127
R2597 vdd.n2958 vdd.n916 99.5127
R2598 vdd.n2958 vdd.n914 99.5127
R2599 vdd.n2962 vdd.n914 99.5127
R2600 vdd.n2962 vdd.n904 99.5127
R2601 vdd.n2970 vdd.n904 99.5127
R2602 vdd.n2970 vdd.n902 99.5127
R2603 vdd.n2974 vdd.n902 99.5127
R2604 vdd.n2974 vdd.n892 99.5127
R2605 vdd.n2982 vdd.n892 99.5127
R2606 vdd.n2982 vdd.n890 99.5127
R2607 vdd.n2986 vdd.n890 99.5127
R2608 vdd.n2986 vdd.n881 99.5127
R2609 vdd.n2994 vdd.n881 99.5127
R2610 vdd.n2994 vdd.n879 99.5127
R2611 vdd.n2998 vdd.n879 99.5127
R2612 vdd.n2998 vdd.n867 99.5127
R2613 vdd.n3007 vdd.n867 99.5127
R2614 vdd.n3007 vdd.n865 99.5127
R2615 vdd.n3011 vdd.n865 99.5127
R2616 vdd.n3011 vdd.n856 99.5127
R2617 vdd.n3019 vdd.n856 99.5127
R2618 vdd.n3019 vdd.n854 99.5127
R2619 vdd.n3023 vdd.n854 99.5127
R2620 vdd.n3023 vdd.n842 99.5127
R2621 vdd.n3076 vdd.n842 99.5127
R2622 vdd.n3076 vdd.n840 99.5127
R2623 vdd.n3080 vdd.n840 99.5127
R2624 vdd.n3080 vdd.n808 99.5127
R2625 vdd.n3150 vdd.n808 99.5127
R2626 vdd.n3146 vdd.n809 99.5127
R2627 vdd.n3144 vdd.n3143 99.5127
R2628 vdd.n3141 vdd.n813 99.5127
R2629 vdd.n3137 vdd.n3136 99.5127
R2630 vdd.n3134 vdd.n816 99.5127
R2631 vdd.n3130 vdd.n3129 99.5127
R2632 vdd.n3127 vdd.n819 99.5127
R2633 vdd.n3123 vdd.n3122 99.5127
R2634 vdd.n3120 vdd.n3118 99.5127
R2635 vdd.n3116 vdd.n822 99.5127
R2636 vdd.n3112 vdd.n3111 99.5127
R2637 vdd.n3109 vdd.n825 99.5127
R2638 vdd.n3105 vdd.n3104 99.5127
R2639 vdd.n3102 vdd.n828 99.5127
R2640 vdd.n3098 vdd.n3097 99.5127
R2641 vdd.n3095 vdd.n831 99.5127
R2642 vdd.n3090 vdd.n3089 99.5127
R2643 vdd.n2867 vdd.n929 99.5127
R2644 vdd.n2863 vdd.n929 99.5127
R2645 vdd.n2863 vdd.n923 99.5127
R2646 vdd.n2807 vdd.n923 99.5127
R2647 vdd.n2807 vdd.n918 99.5127
R2648 vdd.n2810 vdd.n918 99.5127
R2649 vdd.n2810 vdd.n912 99.5127
R2650 vdd.n2813 vdd.n912 99.5127
R2651 vdd.n2813 vdd.n906 99.5127
R2652 vdd.n2846 vdd.n906 99.5127
R2653 vdd.n2846 vdd.n899 99.5127
R2654 vdd.n2842 vdd.n899 99.5127
R2655 vdd.n2842 vdd.n893 99.5127
R2656 vdd.n2839 vdd.n893 99.5127
R2657 vdd.n2839 vdd.n888 99.5127
R2658 vdd.n2836 vdd.n888 99.5127
R2659 vdd.n2836 vdd.n883 99.5127
R2660 vdd.n2833 vdd.n883 99.5127
R2661 vdd.n2833 vdd.n876 99.5127
R2662 vdd.n2830 vdd.n876 99.5127
R2663 vdd.n2830 vdd.n868 99.5127
R2664 vdd.n2827 vdd.n868 99.5127
R2665 vdd.n2827 vdd.n863 99.5127
R2666 vdd.n2824 vdd.n863 99.5127
R2667 vdd.n2824 vdd.n858 99.5127
R2668 vdd.n2821 vdd.n858 99.5127
R2669 vdd.n2821 vdd.n852 99.5127
R2670 vdd.n2818 vdd.n852 99.5127
R2671 vdd.n2818 vdd.n844 99.5127
R2672 vdd.n844 vdd.n837 99.5127
R2673 vdd.n3082 vdd.n837 99.5127
R2674 vdd.n3083 vdd.n3082 99.5127
R2675 vdd.n3083 vdd.n806 99.5127
R2676 vdd.n2700 vdd.n2699 99.5127
R2677 vdd.n2931 vdd.n2699 99.5127
R2678 vdd.n2929 vdd.n2928 99.5127
R2679 vdd.n2925 vdd.n2924 99.5127
R2680 vdd.n2921 vdd.n2920 99.5127
R2681 vdd.n2917 vdd.n2916 99.5127
R2682 vdd.n2913 vdd.n2912 99.5127
R2683 vdd.n2909 vdd.n2908 99.5127
R2684 vdd.n2905 vdd.n2904 99.5127
R2685 vdd.n2901 vdd.n2900 99.5127
R2686 vdd.n2897 vdd.n2896 99.5127
R2687 vdd.n2893 vdd.n2892 99.5127
R2688 vdd.n2889 vdd.n2888 99.5127
R2689 vdd.n2885 vdd.n2884 99.5127
R2690 vdd.n2881 vdd.n2880 99.5127
R2691 vdd.n2877 vdd.n2876 99.5127
R2692 vdd.n2872 vdd.n2871 99.5127
R2693 vdd.n2664 vdd.n970 99.5127
R2694 vdd.n2660 vdd.n2659 99.5127
R2695 vdd.n2656 vdd.n2655 99.5127
R2696 vdd.n2652 vdd.n2651 99.5127
R2697 vdd.n2648 vdd.n2647 99.5127
R2698 vdd.n2644 vdd.n2643 99.5127
R2699 vdd.n2640 vdd.n2639 99.5127
R2700 vdd.n2636 vdd.n2635 99.5127
R2701 vdd.n2632 vdd.n2631 99.5127
R2702 vdd.n2628 vdd.n2627 99.5127
R2703 vdd.n2624 vdd.n2623 99.5127
R2704 vdd.n2620 vdd.n2619 99.5127
R2705 vdd.n2616 vdd.n2615 99.5127
R2706 vdd.n2612 vdd.n2611 99.5127
R2707 vdd.n2608 vdd.n2607 99.5127
R2708 vdd.n2604 vdd.n2603 99.5127
R2709 vdd.n2599 vdd.n2598 99.5127
R2710 vdd.n1309 vdd.n1077 99.5127
R2711 vdd.n1312 vdd.n1077 99.5127
R2712 vdd.n1312 vdd.n1071 99.5127
R2713 vdd.n1315 vdd.n1071 99.5127
R2714 vdd.n1315 vdd.n1066 99.5127
R2715 vdd.n1318 vdd.n1066 99.5127
R2716 vdd.n1318 vdd.n1060 99.5127
R2717 vdd.n1321 vdd.n1060 99.5127
R2718 vdd.n1321 vdd.n1053 99.5127
R2719 vdd.n1324 vdd.n1053 99.5127
R2720 vdd.n1324 vdd.n1046 99.5127
R2721 vdd.n1327 vdd.n1046 99.5127
R2722 vdd.n1327 vdd.n1040 99.5127
R2723 vdd.n1330 vdd.n1040 99.5127
R2724 vdd.n1330 vdd.n1035 99.5127
R2725 vdd.n1333 vdd.n1035 99.5127
R2726 vdd.n1333 vdd.n1029 99.5127
R2727 vdd.n1358 vdd.n1029 99.5127
R2728 vdd.n1358 vdd.n1022 99.5127
R2729 vdd.n1354 vdd.n1022 99.5127
R2730 vdd.n1354 vdd.n1016 99.5127
R2731 vdd.n1351 vdd.n1016 99.5127
R2732 vdd.n1351 vdd.n1011 99.5127
R2733 vdd.n1348 vdd.n1011 99.5127
R2734 vdd.n1348 vdd.n1006 99.5127
R2735 vdd.n1345 vdd.n1006 99.5127
R2736 vdd.n1345 vdd.n1000 99.5127
R2737 vdd.n1342 vdd.n1000 99.5127
R2738 vdd.n1342 vdd.n993 99.5127
R2739 vdd.n1339 vdd.n993 99.5127
R2740 vdd.n1339 vdd.n986 99.5127
R2741 vdd.n986 vdd.n975 99.5127
R2742 vdd.n2594 vdd.n975 99.5127
R2743 vdd.n1118 vdd.n1117 99.5127
R2744 vdd.n2410 vdd.n1117 99.5127
R2745 vdd.n2408 vdd.n2407 99.5127
R2746 vdd.n2404 vdd.n2403 99.5127
R2747 vdd.n2400 vdd.n2399 99.5127
R2748 vdd.n2396 vdd.n2395 99.5127
R2749 vdd.n2392 vdd.n2391 99.5127
R2750 vdd.n2388 vdd.n2387 99.5127
R2751 vdd.n2384 vdd.n2383 99.5127
R2752 vdd.n1276 vdd.n1275 99.5127
R2753 vdd.n1280 vdd.n1279 99.5127
R2754 vdd.n1284 vdd.n1283 99.5127
R2755 vdd.n1288 vdd.n1287 99.5127
R2756 vdd.n1292 vdd.n1291 99.5127
R2757 vdd.n1296 vdd.n1295 99.5127
R2758 vdd.n1300 vdd.n1299 99.5127
R2759 vdd.n1305 vdd.n1304 99.5127
R2760 vdd.n2425 vdd.n1075 99.5127
R2761 vdd.n2425 vdd.n1073 99.5127
R2762 vdd.n2429 vdd.n1073 99.5127
R2763 vdd.n2429 vdd.n1064 99.5127
R2764 vdd.n2437 vdd.n1064 99.5127
R2765 vdd.n2437 vdd.n1062 99.5127
R2766 vdd.n2441 vdd.n1062 99.5127
R2767 vdd.n2441 vdd.n1051 99.5127
R2768 vdd.n2449 vdd.n1051 99.5127
R2769 vdd.n2449 vdd.n1049 99.5127
R2770 vdd.n2453 vdd.n1049 99.5127
R2771 vdd.n2453 vdd.n1039 99.5127
R2772 vdd.n2462 vdd.n1039 99.5127
R2773 vdd.n2462 vdd.n1037 99.5127
R2774 vdd.n2466 vdd.n1037 99.5127
R2775 vdd.n2466 vdd.n1027 99.5127
R2776 vdd.n2474 vdd.n1027 99.5127
R2777 vdd.n2474 vdd.n1025 99.5127
R2778 vdd.n2478 vdd.n1025 99.5127
R2779 vdd.n2478 vdd.n1015 99.5127
R2780 vdd.n2486 vdd.n1015 99.5127
R2781 vdd.n2486 vdd.n1013 99.5127
R2782 vdd.n2490 vdd.n1013 99.5127
R2783 vdd.n2490 vdd.n1004 99.5127
R2784 vdd.n2498 vdd.n1004 99.5127
R2785 vdd.n2498 vdd.n1002 99.5127
R2786 vdd.n2502 vdd.n1002 99.5127
R2787 vdd.n2502 vdd.n991 99.5127
R2788 vdd.n2512 vdd.n991 99.5127
R2789 vdd.n2512 vdd.n988 99.5127
R2790 vdd.n2517 vdd.n988 99.5127
R2791 vdd.n2517 vdd.n989 99.5127
R2792 vdd.n989 vdd.n969 99.5127
R2793 vdd.n3066 vdd.n3065 99.5127
R2794 vdd.n3063 vdd.n3029 99.5127
R2795 vdd.n3059 vdd.n3058 99.5127
R2796 vdd.n3056 vdd.n3032 99.5127
R2797 vdd.n3052 vdd.n3051 99.5127
R2798 vdd.n3049 vdd.n3035 99.5127
R2799 vdd.n3045 vdd.n3044 99.5127
R2800 vdd.n3042 vdd.n3039 99.5127
R2801 vdd.n3183 vdd.n787 99.5127
R2802 vdd.n3181 vdd.n3180 99.5127
R2803 vdd.n3178 vdd.n789 99.5127
R2804 vdd.n3174 vdd.n3173 99.5127
R2805 vdd.n3171 vdd.n792 99.5127
R2806 vdd.n3167 vdd.n3166 99.5127
R2807 vdd.n3164 vdd.n795 99.5127
R2808 vdd.n3160 vdd.n3159 99.5127
R2809 vdd.n3157 vdd.n798 99.5127
R2810 vdd.n2772 vdd.n930 99.5127
R2811 vdd.n2861 vdd.n930 99.5127
R2812 vdd.n2861 vdd.n924 99.5127
R2813 vdd.n2857 vdd.n924 99.5127
R2814 vdd.n2857 vdd.n919 99.5127
R2815 vdd.n2854 vdd.n919 99.5127
R2816 vdd.n2854 vdd.n913 99.5127
R2817 vdd.n2851 vdd.n913 99.5127
R2818 vdd.n2851 vdd.n907 99.5127
R2819 vdd.n2848 vdd.n907 99.5127
R2820 vdd.n2848 vdd.n900 99.5127
R2821 vdd.n2804 vdd.n900 99.5127
R2822 vdd.n2804 vdd.n894 99.5127
R2823 vdd.n2801 vdd.n894 99.5127
R2824 vdd.n2801 vdd.n889 99.5127
R2825 vdd.n2798 vdd.n889 99.5127
R2826 vdd.n2798 vdd.n884 99.5127
R2827 vdd.n2795 vdd.n884 99.5127
R2828 vdd.n2795 vdd.n877 99.5127
R2829 vdd.n2792 vdd.n877 99.5127
R2830 vdd.n2792 vdd.n869 99.5127
R2831 vdd.n2789 vdd.n869 99.5127
R2832 vdd.n2789 vdd.n864 99.5127
R2833 vdd.n2786 vdd.n864 99.5127
R2834 vdd.n2786 vdd.n859 99.5127
R2835 vdd.n2783 vdd.n859 99.5127
R2836 vdd.n2783 vdd.n853 99.5127
R2837 vdd.n2780 vdd.n853 99.5127
R2838 vdd.n2780 vdd.n845 99.5127
R2839 vdd.n2777 vdd.n845 99.5127
R2840 vdd.n2777 vdd.n838 99.5127
R2841 vdd.n838 vdd.n804 99.5127
R2842 vdd.n3152 vdd.n804 99.5127
R2843 vdd.n2707 vdd.n933 99.5127
R2844 vdd.n2711 vdd.n2710 99.5127
R2845 vdd.n2715 vdd.n2714 99.5127
R2846 vdd.n2719 vdd.n2718 99.5127
R2847 vdd.n2723 vdd.n2722 99.5127
R2848 vdd.n2727 vdd.n2726 99.5127
R2849 vdd.n2731 vdd.n2730 99.5127
R2850 vdd.n2735 vdd.n2734 99.5127
R2851 vdd.n2739 vdd.n2738 99.5127
R2852 vdd.n2743 vdd.n2742 99.5127
R2853 vdd.n2747 vdd.n2746 99.5127
R2854 vdd.n2751 vdd.n2750 99.5127
R2855 vdd.n2755 vdd.n2754 99.5127
R2856 vdd.n2759 vdd.n2758 99.5127
R2857 vdd.n2763 vdd.n2762 99.5127
R2858 vdd.n2767 vdd.n2766 99.5127
R2859 vdd.n2769 vdd.n2698 99.5127
R2860 vdd.n2944 vdd.n931 99.5127
R2861 vdd.n2944 vdd.n922 99.5127
R2862 vdd.n2952 vdd.n922 99.5127
R2863 vdd.n2952 vdd.n920 99.5127
R2864 vdd.n2956 vdd.n920 99.5127
R2865 vdd.n2956 vdd.n910 99.5127
R2866 vdd.n2964 vdd.n910 99.5127
R2867 vdd.n2964 vdd.n908 99.5127
R2868 vdd.n2968 vdd.n908 99.5127
R2869 vdd.n2968 vdd.n898 99.5127
R2870 vdd.n2976 vdd.n898 99.5127
R2871 vdd.n2976 vdd.n896 99.5127
R2872 vdd.n2980 vdd.n896 99.5127
R2873 vdd.n2980 vdd.n887 99.5127
R2874 vdd.n2988 vdd.n887 99.5127
R2875 vdd.n2988 vdd.n885 99.5127
R2876 vdd.n2992 vdd.n885 99.5127
R2877 vdd.n2992 vdd.n874 99.5127
R2878 vdd.n3000 vdd.n874 99.5127
R2879 vdd.n3000 vdd.n871 99.5127
R2880 vdd.n3005 vdd.n871 99.5127
R2881 vdd.n3005 vdd.n862 99.5127
R2882 vdd.n3013 vdd.n862 99.5127
R2883 vdd.n3013 vdd.n860 99.5127
R2884 vdd.n3017 vdd.n860 99.5127
R2885 vdd.n3017 vdd.n850 99.5127
R2886 vdd.n3025 vdd.n850 99.5127
R2887 vdd.n3025 vdd.n847 99.5127
R2888 vdd.n3074 vdd.n847 99.5127
R2889 vdd.n3074 vdd.n848 99.5127
R2890 vdd.n848 vdd.n839 99.5127
R2891 vdd.n3069 vdd.n839 99.5127
R2892 vdd.n3069 vdd.n807 99.5127
R2893 vdd.n2588 vdd.n2587 99.5127
R2894 vdd.n2584 vdd.n2583 99.5127
R2895 vdd.n2580 vdd.n2579 99.5127
R2896 vdd.n2576 vdd.n2575 99.5127
R2897 vdd.n2572 vdd.n2571 99.5127
R2898 vdd.n2568 vdd.n2567 99.5127
R2899 vdd.n2564 vdd.n2563 99.5127
R2900 vdd.n2560 vdd.n2559 99.5127
R2901 vdd.n2556 vdd.n2555 99.5127
R2902 vdd.n2552 vdd.n2551 99.5127
R2903 vdd.n2548 vdd.n2547 99.5127
R2904 vdd.n2544 vdd.n2543 99.5127
R2905 vdd.n2540 vdd.n2539 99.5127
R2906 vdd.n2536 vdd.n2535 99.5127
R2907 vdd.n2532 vdd.n2531 99.5127
R2908 vdd.n2528 vdd.n2527 99.5127
R2909 vdd.n2524 vdd.n951 99.5127
R2910 vdd.n1387 vdd.n1078 99.5127
R2911 vdd.n1384 vdd.n1078 99.5127
R2912 vdd.n1384 vdd.n1072 99.5127
R2913 vdd.n1381 vdd.n1072 99.5127
R2914 vdd.n1381 vdd.n1067 99.5127
R2915 vdd.n1378 vdd.n1067 99.5127
R2916 vdd.n1378 vdd.n1061 99.5127
R2917 vdd.n1375 vdd.n1061 99.5127
R2918 vdd.n1375 vdd.n1054 99.5127
R2919 vdd.n1372 vdd.n1054 99.5127
R2920 vdd.n1372 vdd.n1047 99.5127
R2921 vdd.n1369 vdd.n1047 99.5127
R2922 vdd.n1369 vdd.n1041 99.5127
R2923 vdd.n1366 vdd.n1041 99.5127
R2924 vdd.n1366 vdd.n1036 99.5127
R2925 vdd.n1363 vdd.n1036 99.5127
R2926 vdd.n1363 vdd.n1030 99.5127
R2927 vdd.n1360 vdd.n1030 99.5127
R2928 vdd.n1360 vdd.n1023 99.5127
R2929 vdd.n1270 vdd.n1023 99.5127
R2930 vdd.n1270 vdd.n1017 99.5127
R2931 vdd.n1267 vdd.n1017 99.5127
R2932 vdd.n1267 vdd.n1012 99.5127
R2933 vdd.n1264 vdd.n1012 99.5127
R2934 vdd.n1264 vdd.n1007 99.5127
R2935 vdd.n1261 vdd.n1007 99.5127
R2936 vdd.n1261 vdd.n1001 99.5127
R2937 vdd.n1258 vdd.n1001 99.5127
R2938 vdd.n1258 vdd.n994 99.5127
R2939 vdd.n994 vdd.n985 99.5127
R2940 vdd.n2519 vdd.n985 99.5127
R2941 vdd.n2520 vdd.n2519 99.5127
R2942 vdd.n2520 vdd.n977 99.5127
R2943 vdd.n1222 vdd.n1082 99.5127
R2944 vdd.n1226 vdd.n1225 99.5127
R2945 vdd.n1230 vdd.n1229 99.5127
R2946 vdd.n1234 vdd.n1233 99.5127
R2947 vdd.n1238 vdd.n1237 99.5127
R2948 vdd.n1242 vdd.n1241 99.5127
R2949 vdd.n1246 vdd.n1245 99.5127
R2950 vdd.n1250 vdd.n1249 99.5127
R2951 vdd.n1420 vdd.n1252 99.5127
R2952 vdd.n1418 vdd.n1417 99.5127
R2953 vdd.n1414 vdd.n1413 99.5127
R2954 vdd.n1410 vdd.n1409 99.5127
R2955 vdd.n1406 vdd.n1405 99.5127
R2956 vdd.n1402 vdd.n1401 99.5127
R2957 vdd.n1398 vdd.n1397 99.5127
R2958 vdd.n1394 vdd.n1393 99.5127
R2959 vdd.n1390 vdd.n1116 99.5127
R2960 vdd.n2423 vdd.n1080 99.5127
R2961 vdd.n2423 vdd.n1070 99.5127
R2962 vdd.n2431 vdd.n1070 99.5127
R2963 vdd.n2431 vdd.n1068 99.5127
R2964 vdd.n2435 vdd.n1068 99.5127
R2965 vdd.n2435 vdd.n1058 99.5127
R2966 vdd.n2443 vdd.n1058 99.5127
R2967 vdd.n2443 vdd.n1056 99.5127
R2968 vdd.n2447 vdd.n1056 99.5127
R2969 vdd.n2447 vdd.n1045 99.5127
R2970 vdd.n2455 vdd.n1045 99.5127
R2971 vdd.n2455 vdd.n1042 99.5127
R2972 vdd.n2460 vdd.n1042 99.5127
R2973 vdd.n2460 vdd.n1033 99.5127
R2974 vdd.n2468 vdd.n1033 99.5127
R2975 vdd.n2468 vdd.n1031 99.5127
R2976 vdd.n2472 vdd.n1031 99.5127
R2977 vdd.n2472 vdd.n1021 99.5127
R2978 vdd.n2480 vdd.n1021 99.5127
R2979 vdd.n2480 vdd.n1019 99.5127
R2980 vdd.n2484 vdd.n1019 99.5127
R2981 vdd.n2484 vdd.n1010 99.5127
R2982 vdd.n2492 vdd.n1010 99.5127
R2983 vdd.n2492 vdd.n1008 99.5127
R2984 vdd.n2496 vdd.n1008 99.5127
R2985 vdd.n2496 vdd.n998 99.5127
R2986 vdd.n2504 vdd.n998 99.5127
R2987 vdd.n2504 vdd.n995 99.5127
R2988 vdd.n2510 vdd.n995 99.5127
R2989 vdd.n2510 vdd.n996 99.5127
R2990 vdd.n996 vdd.n987 99.5127
R2991 vdd.n987 vdd.n978 99.5127
R2992 vdd.n2592 vdd.n978 99.5127
R2993 vdd.n9 vdd.n7 98.9633
R2994 vdd.n2 vdd.n0 98.9633
R2995 vdd.n9 vdd.n8 98.6055
R2996 vdd.n11 vdd.n10 98.6055
R2997 vdd.n13 vdd.n12 98.6055
R2998 vdd.n6 vdd.n5 98.6055
R2999 vdd.n4 vdd.n3 98.6055
R3000 vdd.n2 vdd.n1 98.6055
R3001 vdd.t160 vdd.n303 85.8723
R3002 vdd.t240 vdd.n244 85.8723
R3003 vdd.t291 vdd.n201 85.8723
R3004 vdd.t228 vdd.n142 85.8723
R3005 vdd.t197 vdd.n100 85.8723
R3006 vdd.t189 vdd.n41 85.8723
R3007 vdd.t282 vdd.n2084 85.8723
R3008 vdd.t220 vdd.n2143 85.8723
R3009 vdd.t271 vdd.n1982 85.8723
R3010 vdd.t145 vdd.n2041 85.8723
R3011 vdd.t191 vdd.n1881 85.8723
R3012 vdd.t196 vdd.n1940 85.8723
R3013 vdd.n3003 vdd.n872 78.546
R3014 vdd.n2458 vdd.n1043 78.546
R3015 vdd.n290 vdd.n289 75.1835
R3016 vdd.n288 vdd.n287 75.1835
R3017 vdd.n286 vdd.n285 75.1835
R3018 vdd.n284 vdd.n283 75.1835
R3019 vdd.n282 vdd.n281 75.1835
R3020 vdd.n280 vdd.n279 75.1835
R3021 vdd.n278 vdd.n277 75.1835
R3022 vdd.n276 vdd.n275 75.1835
R3023 vdd.n274 vdd.n273 75.1835
R3024 vdd.n188 vdd.n187 75.1835
R3025 vdd.n186 vdd.n185 75.1835
R3026 vdd.n184 vdd.n183 75.1835
R3027 vdd.n182 vdd.n181 75.1835
R3028 vdd.n180 vdd.n179 75.1835
R3029 vdd.n178 vdd.n177 75.1835
R3030 vdd.n176 vdd.n175 75.1835
R3031 vdd.n174 vdd.n173 75.1835
R3032 vdd.n172 vdd.n171 75.1835
R3033 vdd.n87 vdd.n86 75.1835
R3034 vdd.n85 vdd.n84 75.1835
R3035 vdd.n83 vdd.n82 75.1835
R3036 vdd.n81 vdd.n80 75.1835
R3037 vdd.n79 vdd.n78 75.1835
R3038 vdd.n77 vdd.n76 75.1835
R3039 vdd.n75 vdd.n74 75.1835
R3040 vdd.n73 vdd.n72 75.1835
R3041 vdd.n71 vdd.n70 75.1835
R3042 vdd.n2114 vdd.n2113 75.1835
R3043 vdd.n2116 vdd.n2115 75.1835
R3044 vdd.n2118 vdd.n2117 75.1835
R3045 vdd.n2120 vdd.n2119 75.1835
R3046 vdd.n2122 vdd.n2121 75.1835
R3047 vdd.n2124 vdd.n2123 75.1835
R3048 vdd.n2126 vdd.n2125 75.1835
R3049 vdd.n2128 vdd.n2127 75.1835
R3050 vdd.n2130 vdd.n2129 75.1835
R3051 vdd.n2012 vdd.n2011 75.1835
R3052 vdd.n2014 vdd.n2013 75.1835
R3053 vdd.n2016 vdd.n2015 75.1835
R3054 vdd.n2018 vdd.n2017 75.1835
R3055 vdd.n2020 vdd.n2019 75.1835
R3056 vdd.n2022 vdd.n2021 75.1835
R3057 vdd.n2024 vdd.n2023 75.1835
R3058 vdd.n2026 vdd.n2025 75.1835
R3059 vdd.n2028 vdd.n2027 75.1835
R3060 vdd.n1911 vdd.n1910 75.1835
R3061 vdd.n1913 vdd.n1912 75.1835
R3062 vdd.n1915 vdd.n1914 75.1835
R3063 vdd.n1917 vdd.n1916 75.1835
R3064 vdd.n1919 vdd.n1918 75.1835
R3065 vdd.n1921 vdd.n1920 75.1835
R3066 vdd.n1923 vdd.n1922 75.1835
R3067 vdd.n1925 vdd.n1924 75.1835
R3068 vdd.n1927 vdd.n1926 75.1835
R3069 vdd.n2939 vdd.n2938 72.8958
R3070 vdd.n2938 vdd.n2682 72.8958
R3071 vdd.n2938 vdd.n2683 72.8958
R3072 vdd.n2938 vdd.n2684 72.8958
R3073 vdd.n2938 vdd.n2685 72.8958
R3074 vdd.n2938 vdd.n2686 72.8958
R3075 vdd.n2938 vdd.n2687 72.8958
R3076 vdd.n2938 vdd.n2688 72.8958
R3077 vdd.n2938 vdd.n2689 72.8958
R3078 vdd.n2938 vdd.n2690 72.8958
R3079 vdd.n2938 vdd.n2691 72.8958
R3080 vdd.n2938 vdd.n2692 72.8958
R3081 vdd.n2938 vdd.n2693 72.8958
R3082 vdd.n2938 vdd.n2694 72.8958
R3083 vdd.n2938 vdd.n2695 72.8958
R3084 vdd.n2938 vdd.n2696 72.8958
R3085 vdd.n2938 vdd.n2697 72.8958
R3086 vdd.n803 vdd.n692 72.8958
R3087 vdd.n3158 vdd.n692 72.8958
R3088 vdd.n797 vdd.n692 72.8958
R3089 vdd.n3165 vdd.n692 72.8958
R3090 vdd.n794 vdd.n692 72.8958
R3091 vdd.n3172 vdd.n692 72.8958
R3092 vdd.n791 vdd.n692 72.8958
R3093 vdd.n3179 vdd.n692 72.8958
R3094 vdd.n3182 vdd.n692 72.8958
R3095 vdd.n3038 vdd.n692 72.8958
R3096 vdd.n3043 vdd.n692 72.8958
R3097 vdd.n3037 vdd.n692 72.8958
R3098 vdd.n3050 vdd.n692 72.8958
R3099 vdd.n3034 vdd.n692 72.8958
R3100 vdd.n3057 vdd.n692 72.8958
R3101 vdd.n3031 vdd.n692 72.8958
R3102 vdd.n3064 vdd.n692 72.8958
R3103 vdd.n2417 vdd.n2416 72.8958
R3104 vdd.n2417 vdd.n1084 72.8958
R3105 vdd.n2417 vdd.n1085 72.8958
R3106 vdd.n2417 vdd.n1086 72.8958
R3107 vdd.n2417 vdd.n1087 72.8958
R3108 vdd.n2417 vdd.n1088 72.8958
R3109 vdd.n2417 vdd.n1089 72.8958
R3110 vdd.n2417 vdd.n1090 72.8958
R3111 vdd.n2417 vdd.n1091 72.8958
R3112 vdd.n2417 vdd.n1092 72.8958
R3113 vdd.n2417 vdd.n1093 72.8958
R3114 vdd.n2417 vdd.n1094 72.8958
R3115 vdd.n2417 vdd.n1095 72.8958
R3116 vdd.n2417 vdd.n1096 72.8958
R3117 vdd.n2417 vdd.n1097 72.8958
R3118 vdd.n2417 vdd.n1098 72.8958
R3119 vdd.n2417 vdd.n1099 72.8958
R3120 vdd.n2665 vdd.n952 72.8958
R3121 vdd.n2665 vdd.n953 72.8958
R3122 vdd.n2665 vdd.n954 72.8958
R3123 vdd.n2665 vdd.n955 72.8958
R3124 vdd.n2665 vdd.n956 72.8958
R3125 vdd.n2665 vdd.n957 72.8958
R3126 vdd.n2665 vdd.n958 72.8958
R3127 vdd.n2665 vdd.n959 72.8958
R3128 vdd.n2665 vdd.n960 72.8958
R3129 vdd.n2665 vdd.n961 72.8958
R3130 vdd.n2665 vdd.n962 72.8958
R3131 vdd.n2665 vdd.n963 72.8958
R3132 vdd.n2665 vdd.n964 72.8958
R3133 vdd.n2665 vdd.n965 72.8958
R3134 vdd.n2665 vdd.n966 72.8958
R3135 vdd.n2665 vdd.n967 72.8958
R3136 vdd.n2665 vdd.n968 72.8958
R3137 vdd.n2938 vdd.n2937 72.8958
R3138 vdd.n2938 vdd.n2666 72.8958
R3139 vdd.n2938 vdd.n2667 72.8958
R3140 vdd.n2938 vdd.n2668 72.8958
R3141 vdd.n2938 vdd.n2669 72.8958
R3142 vdd.n2938 vdd.n2670 72.8958
R3143 vdd.n2938 vdd.n2671 72.8958
R3144 vdd.n2938 vdd.n2672 72.8958
R3145 vdd.n2938 vdd.n2673 72.8958
R3146 vdd.n2938 vdd.n2674 72.8958
R3147 vdd.n2938 vdd.n2675 72.8958
R3148 vdd.n2938 vdd.n2676 72.8958
R3149 vdd.n2938 vdd.n2677 72.8958
R3150 vdd.n2938 vdd.n2678 72.8958
R3151 vdd.n2938 vdd.n2679 72.8958
R3152 vdd.n2938 vdd.n2680 72.8958
R3153 vdd.n2938 vdd.n2681 72.8958
R3154 vdd.n3088 vdd.n692 72.8958
R3155 vdd.n835 vdd.n692 72.8958
R3156 vdd.n3096 vdd.n692 72.8958
R3157 vdd.n830 vdd.n692 72.8958
R3158 vdd.n3103 vdd.n692 72.8958
R3159 vdd.n827 vdd.n692 72.8958
R3160 vdd.n3110 vdd.n692 72.8958
R3161 vdd.n824 vdd.n692 72.8958
R3162 vdd.n3117 vdd.n692 72.8958
R3163 vdd.n3121 vdd.n692 72.8958
R3164 vdd.n821 vdd.n692 72.8958
R3165 vdd.n3128 vdd.n692 72.8958
R3166 vdd.n818 vdd.n692 72.8958
R3167 vdd.n3135 vdd.n692 72.8958
R3168 vdd.n815 vdd.n692 72.8958
R3169 vdd.n3142 vdd.n692 72.8958
R3170 vdd.n3145 vdd.n692 72.8958
R3171 vdd.n2665 vdd.n950 72.8958
R3172 vdd.n2665 vdd.n949 72.8958
R3173 vdd.n2665 vdd.n948 72.8958
R3174 vdd.n2665 vdd.n947 72.8958
R3175 vdd.n2665 vdd.n946 72.8958
R3176 vdd.n2665 vdd.n945 72.8958
R3177 vdd.n2665 vdd.n944 72.8958
R3178 vdd.n2665 vdd.n943 72.8958
R3179 vdd.n2665 vdd.n942 72.8958
R3180 vdd.n2665 vdd.n941 72.8958
R3181 vdd.n2665 vdd.n940 72.8958
R3182 vdd.n2665 vdd.n939 72.8958
R3183 vdd.n2665 vdd.n938 72.8958
R3184 vdd.n2665 vdd.n937 72.8958
R3185 vdd.n2665 vdd.n936 72.8958
R3186 vdd.n2665 vdd.n935 72.8958
R3187 vdd.n2665 vdd.n934 72.8958
R3188 vdd.n2418 vdd.n2417 72.8958
R3189 vdd.n2417 vdd.n1100 72.8958
R3190 vdd.n2417 vdd.n1101 72.8958
R3191 vdd.n2417 vdd.n1102 72.8958
R3192 vdd.n2417 vdd.n1103 72.8958
R3193 vdd.n2417 vdd.n1104 72.8958
R3194 vdd.n2417 vdd.n1105 72.8958
R3195 vdd.n2417 vdd.n1106 72.8958
R3196 vdd.n2417 vdd.n1107 72.8958
R3197 vdd.n2417 vdd.n1108 72.8958
R3198 vdd.n2417 vdd.n1109 72.8958
R3199 vdd.n2417 vdd.n1110 72.8958
R3200 vdd.n2417 vdd.n1111 72.8958
R3201 vdd.n2417 vdd.n1112 72.8958
R3202 vdd.n2417 vdd.n1113 72.8958
R3203 vdd.n2417 vdd.n1114 72.8958
R3204 vdd.n2417 vdd.n1115 72.8958
R3205 vdd.n1781 vdd.n1780 66.2847
R3206 vdd.n1780 vdd.n1556 66.2847
R3207 vdd.n1780 vdd.n1557 66.2847
R3208 vdd.n1780 vdd.n1558 66.2847
R3209 vdd.n1780 vdd.n1559 66.2847
R3210 vdd.n1780 vdd.n1560 66.2847
R3211 vdd.n1780 vdd.n1561 66.2847
R3212 vdd.n1780 vdd.n1562 66.2847
R3213 vdd.n1780 vdd.n1563 66.2847
R3214 vdd.n1780 vdd.n1564 66.2847
R3215 vdd.n1780 vdd.n1565 66.2847
R3216 vdd.n1780 vdd.n1566 66.2847
R3217 vdd.n1780 vdd.n1567 66.2847
R3218 vdd.n1780 vdd.n1568 66.2847
R3219 vdd.n1780 vdd.n1569 66.2847
R3220 vdd.n1780 vdd.n1570 66.2847
R3221 vdd.n1780 vdd.n1571 66.2847
R3222 vdd.n1780 vdd.n1572 66.2847
R3223 vdd.n1780 vdd.n1573 66.2847
R3224 vdd.n1780 vdd.n1574 66.2847
R3225 vdd.n1780 vdd.n1575 66.2847
R3226 vdd.n1780 vdd.n1576 66.2847
R3227 vdd.n1780 vdd.n1577 66.2847
R3228 vdd.n1780 vdd.n1578 66.2847
R3229 vdd.n1780 vdd.n1579 66.2847
R3230 vdd.n1780 vdd.n1580 66.2847
R3231 vdd.n1780 vdd.n1581 66.2847
R3232 vdd.n1780 vdd.n1582 66.2847
R3233 vdd.n1780 vdd.n1583 66.2847
R3234 vdd.n1780 vdd.n1584 66.2847
R3235 vdd.n1780 vdd.n1585 66.2847
R3236 vdd.n1433 vdd.n1083 66.2847
R3237 vdd.n1430 vdd.n1083 66.2847
R3238 vdd.n1426 vdd.n1083 66.2847
R3239 vdd.n2279 vdd.n1083 66.2847
R3240 vdd.n1217 vdd.n1083 66.2847
R3241 vdd.n2286 vdd.n1083 66.2847
R3242 vdd.n1210 vdd.n1083 66.2847
R3243 vdd.n2293 vdd.n1083 66.2847
R3244 vdd.n1203 vdd.n1083 66.2847
R3245 vdd.n2300 vdd.n1083 66.2847
R3246 vdd.n1197 vdd.n1083 66.2847
R3247 vdd.n1192 vdd.n1083 66.2847
R3248 vdd.n2311 vdd.n1083 66.2847
R3249 vdd.n1184 vdd.n1083 66.2847
R3250 vdd.n2318 vdd.n1083 66.2847
R3251 vdd.n1177 vdd.n1083 66.2847
R3252 vdd.n2325 vdd.n1083 66.2847
R3253 vdd.n1170 vdd.n1083 66.2847
R3254 vdd.n2332 vdd.n1083 66.2847
R3255 vdd.n1163 vdd.n1083 66.2847
R3256 vdd.n2339 vdd.n1083 66.2847
R3257 vdd.n1157 vdd.n1083 66.2847
R3258 vdd.n1152 vdd.n1083 66.2847
R3259 vdd.n2350 vdd.n1083 66.2847
R3260 vdd.n1144 vdd.n1083 66.2847
R3261 vdd.n2357 vdd.n1083 66.2847
R3262 vdd.n1137 vdd.n1083 66.2847
R3263 vdd.n2364 vdd.n1083 66.2847
R3264 vdd.n1130 vdd.n1083 66.2847
R3265 vdd.n2371 vdd.n1083 66.2847
R3266 vdd.n2376 vdd.n1083 66.2847
R3267 vdd.n1126 vdd.n1083 66.2847
R3268 vdd.n3315 vdd.n3314 66.2847
R3269 vdd.n3315 vdd.n693 66.2847
R3270 vdd.n3315 vdd.n694 66.2847
R3271 vdd.n3315 vdd.n695 66.2847
R3272 vdd.n3315 vdd.n696 66.2847
R3273 vdd.n3315 vdd.n697 66.2847
R3274 vdd.n3315 vdd.n698 66.2847
R3275 vdd.n3315 vdd.n699 66.2847
R3276 vdd.n3315 vdd.n700 66.2847
R3277 vdd.n3315 vdd.n701 66.2847
R3278 vdd.n3315 vdd.n702 66.2847
R3279 vdd.n3315 vdd.n703 66.2847
R3280 vdd.n3315 vdd.n704 66.2847
R3281 vdd.n3315 vdd.n705 66.2847
R3282 vdd.n3315 vdd.n706 66.2847
R3283 vdd.n3315 vdd.n707 66.2847
R3284 vdd.n3315 vdd.n708 66.2847
R3285 vdd.n3315 vdd.n709 66.2847
R3286 vdd.n3315 vdd.n710 66.2847
R3287 vdd.n3315 vdd.n711 66.2847
R3288 vdd.n3315 vdd.n712 66.2847
R3289 vdd.n3315 vdd.n713 66.2847
R3290 vdd.n3315 vdd.n714 66.2847
R3291 vdd.n3315 vdd.n715 66.2847
R3292 vdd.n3315 vdd.n716 66.2847
R3293 vdd.n3315 vdd.n717 66.2847
R3294 vdd.n3315 vdd.n718 66.2847
R3295 vdd.n3315 vdd.n719 66.2847
R3296 vdd.n3315 vdd.n720 66.2847
R3297 vdd.n3315 vdd.n721 66.2847
R3298 vdd.n3315 vdd.n722 66.2847
R3299 vdd.n3446 vdd.n3445 66.2847
R3300 vdd.n3446 vdd.n424 66.2847
R3301 vdd.n3446 vdd.n423 66.2847
R3302 vdd.n3446 vdd.n422 66.2847
R3303 vdd.n3446 vdd.n421 66.2847
R3304 vdd.n3446 vdd.n420 66.2847
R3305 vdd.n3446 vdd.n419 66.2847
R3306 vdd.n3446 vdd.n418 66.2847
R3307 vdd.n3446 vdd.n417 66.2847
R3308 vdd.n3446 vdd.n416 66.2847
R3309 vdd.n3446 vdd.n415 66.2847
R3310 vdd.n3446 vdd.n414 66.2847
R3311 vdd.n3446 vdd.n413 66.2847
R3312 vdd.n3446 vdd.n412 66.2847
R3313 vdd.n3446 vdd.n411 66.2847
R3314 vdd.n3446 vdd.n410 66.2847
R3315 vdd.n3446 vdd.n409 66.2847
R3316 vdd.n3446 vdd.n408 66.2847
R3317 vdd.n3446 vdd.n407 66.2847
R3318 vdd.n3446 vdd.n406 66.2847
R3319 vdd.n3446 vdd.n405 66.2847
R3320 vdd.n3446 vdd.n404 66.2847
R3321 vdd.n3446 vdd.n403 66.2847
R3322 vdd.n3446 vdd.n402 66.2847
R3323 vdd.n3446 vdd.n401 66.2847
R3324 vdd.n3446 vdd.n400 66.2847
R3325 vdd.n3446 vdd.n399 66.2847
R3326 vdd.n3446 vdd.n398 66.2847
R3327 vdd.n3446 vdd.n397 66.2847
R3328 vdd.n3446 vdd.n396 66.2847
R3329 vdd.n3446 vdd.n395 66.2847
R3330 vdd.n3446 vdd.n394 66.2847
R3331 vdd.n467 vdd.n394 52.4337
R3332 vdd.n473 vdd.n395 52.4337
R3333 vdd.n477 vdd.n396 52.4337
R3334 vdd.n483 vdd.n397 52.4337
R3335 vdd.n487 vdd.n398 52.4337
R3336 vdd.n493 vdd.n399 52.4337
R3337 vdd.n497 vdd.n400 52.4337
R3338 vdd.n503 vdd.n401 52.4337
R3339 vdd.n507 vdd.n402 52.4337
R3340 vdd.n513 vdd.n403 52.4337
R3341 vdd.n517 vdd.n404 52.4337
R3342 vdd.n523 vdd.n405 52.4337
R3343 vdd.n527 vdd.n406 52.4337
R3344 vdd.n533 vdd.n407 52.4337
R3345 vdd.n537 vdd.n408 52.4337
R3346 vdd.n543 vdd.n409 52.4337
R3347 vdd.n547 vdd.n410 52.4337
R3348 vdd.n553 vdd.n411 52.4337
R3349 vdd.n557 vdd.n412 52.4337
R3350 vdd.n563 vdd.n413 52.4337
R3351 vdd.n567 vdd.n414 52.4337
R3352 vdd.n573 vdd.n415 52.4337
R3353 vdd.n577 vdd.n416 52.4337
R3354 vdd.n583 vdd.n417 52.4337
R3355 vdd.n587 vdd.n418 52.4337
R3356 vdd.n593 vdd.n419 52.4337
R3357 vdd.n597 vdd.n420 52.4337
R3358 vdd.n603 vdd.n421 52.4337
R3359 vdd.n607 vdd.n422 52.4337
R3360 vdd.n613 vdd.n423 52.4337
R3361 vdd.n616 vdd.n424 52.4337
R3362 vdd.n3445 vdd.n3444 52.4337
R3363 vdd.n3314 vdd.n3313 52.4337
R3364 vdd.n728 vdd.n693 52.4337
R3365 vdd.n734 vdd.n694 52.4337
R3366 vdd.n3303 vdd.n695 52.4337
R3367 vdd.n3299 vdd.n696 52.4337
R3368 vdd.n3295 vdd.n697 52.4337
R3369 vdd.n3291 vdd.n698 52.4337
R3370 vdd.n3287 vdd.n699 52.4337
R3371 vdd.n3283 vdd.n700 52.4337
R3372 vdd.n3279 vdd.n701 52.4337
R3373 vdd.n3271 vdd.n702 52.4337
R3374 vdd.n3267 vdd.n703 52.4337
R3375 vdd.n3263 vdd.n704 52.4337
R3376 vdd.n3259 vdd.n705 52.4337
R3377 vdd.n3255 vdd.n706 52.4337
R3378 vdd.n3251 vdd.n707 52.4337
R3379 vdd.n3247 vdd.n708 52.4337
R3380 vdd.n3243 vdd.n709 52.4337
R3381 vdd.n3239 vdd.n710 52.4337
R3382 vdd.n3235 vdd.n711 52.4337
R3383 vdd.n3231 vdd.n712 52.4337
R3384 vdd.n3225 vdd.n713 52.4337
R3385 vdd.n3221 vdd.n714 52.4337
R3386 vdd.n3217 vdd.n715 52.4337
R3387 vdd.n3213 vdd.n716 52.4337
R3388 vdd.n3209 vdd.n717 52.4337
R3389 vdd.n3205 vdd.n718 52.4337
R3390 vdd.n3201 vdd.n719 52.4337
R3391 vdd.n3197 vdd.n720 52.4337
R3392 vdd.n3193 vdd.n721 52.4337
R3393 vdd.n3189 vdd.n722 52.4337
R3394 vdd.n2378 vdd.n1126 52.4337
R3395 vdd.n2376 vdd.n2375 52.4337
R3396 vdd.n2371 vdd.n2370 52.4337
R3397 vdd.n2366 vdd.n1130 52.4337
R3398 vdd.n2364 vdd.n2363 52.4337
R3399 vdd.n2359 vdd.n1137 52.4337
R3400 vdd.n2357 vdd.n2356 52.4337
R3401 vdd.n2352 vdd.n1144 52.4337
R3402 vdd.n2350 vdd.n2349 52.4337
R3403 vdd.n1153 vdd.n1152 52.4337
R3404 vdd.n2341 vdd.n1157 52.4337
R3405 vdd.n2339 vdd.n2338 52.4337
R3406 vdd.n2334 vdd.n1163 52.4337
R3407 vdd.n2332 vdd.n2331 52.4337
R3408 vdd.n2327 vdd.n1170 52.4337
R3409 vdd.n2325 vdd.n2324 52.4337
R3410 vdd.n2320 vdd.n1177 52.4337
R3411 vdd.n2318 vdd.n2317 52.4337
R3412 vdd.n2313 vdd.n1184 52.4337
R3413 vdd.n2311 vdd.n2310 52.4337
R3414 vdd.n1193 vdd.n1192 52.4337
R3415 vdd.n2302 vdd.n1197 52.4337
R3416 vdd.n2300 vdd.n2299 52.4337
R3417 vdd.n2295 vdd.n1203 52.4337
R3418 vdd.n2293 vdd.n2292 52.4337
R3419 vdd.n2288 vdd.n1210 52.4337
R3420 vdd.n2286 vdd.n2285 52.4337
R3421 vdd.n2281 vdd.n1217 52.4337
R3422 vdd.n2279 vdd.n2278 52.4337
R3423 vdd.n1427 vdd.n1426 52.4337
R3424 vdd.n1431 vdd.n1430 52.4337
R3425 vdd.n2267 vdd.n1433 52.4337
R3426 vdd.n1782 vdd.n1781 52.4337
R3427 vdd.n1588 vdd.n1556 52.4337
R3428 vdd.n1592 vdd.n1557 52.4337
R3429 vdd.n1594 vdd.n1558 52.4337
R3430 vdd.n1598 vdd.n1559 52.4337
R3431 vdd.n1600 vdd.n1560 52.4337
R3432 vdd.n1604 vdd.n1561 52.4337
R3433 vdd.n1606 vdd.n1562 52.4337
R3434 vdd.n1610 vdd.n1563 52.4337
R3435 vdd.n1612 vdd.n1564 52.4337
R3436 vdd.n1618 vdd.n1565 52.4337
R3437 vdd.n1620 vdd.n1566 52.4337
R3438 vdd.n1624 vdd.n1567 52.4337
R3439 vdd.n1626 vdd.n1568 52.4337
R3440 vdd.n1630 vdd.n1569 52.4337
R3441 vdd.n1632 vdd.n1570 52.4337
R3442 vdd.n1636 vdd.n1571 52.4337
R3443 vdd.n1638 vdd.n1572 52.4337
R3444 vdd.n1642 vdd.n1573 52.4337
R3445 vdd.n1644 vdd.n1574 52.4337
R3446 vdd.n1716 vdd.n1575 52.4337
R3447 vdd.n1649 vdd.n1576 52.4337
R3448 vdd.n1653 vdd.n1577 52.4337
R3449 vdd.n1655 vdd.n1578 52.4337
R3450 vdd.n1659 vdd.n1579 52.4337
R3451 vdd.n1661 vdd.n1580 52.4337
R3452 vdd.n1665 vdd.n1581 52.4337
R3453 vdd.n1667 vdd.n1582 52.4337
R3454 vdd.n1671 vdd.n1583 52.4337
R3455 vdd.n1673 vdd.n1584 52.4337
R3456 vdd.n1677 vdd.n1585 52.4337
R3457 vdd.n1781 vdd.n1555 52.4337
R3458 vdd.n1591 vdd.n1556 52.4337
R3459 vdd.n1593 vdd.n1557 52.4337
R3460 vdd.n1597 vdd.n1558 52.4337
R3461 vdd.n1599 vdd.n1559 52.4337
R3462 vdd.n1603 vdd.n1560 52.4337
R3463 vdd.n1605 vdd.n1561 52.4337
R3464 vdd.n1609 vdd.n1562 52.4337
R3465 vdd.n1611 vdd.n1563 52.4337
R3466 vdd.n1617 vdd.n1564 52.4337
R3467 vdd.n1619 vdd.n1565 52.4337
R3468 vdd.n1623 vdd.n1566 52.4337
R3469 vdd.n1625 vdd.n1567 52.4337
R3470 vdd.n1629 vdd.n1568 52.4337
R3471 vdd.n1631 vdd.n1569 52.4337
R3472 vdd.n1635 vdd.n1570 52.4337
R3473 vdd.n1637 vdd.n1571 52.4337
R3474 vdd.n1641 vdd.n1572 52.4337
R3475 vdd.n1643 vdd.n1573 52.4337
R3476 vdd.n1647 vdd.n1574 52.4337
R3477 vdd.n1648 vdd.n1575 52.4337
R3478 vdd.n1652 vdd.n1576 52.4337
R3479 vdd.n1654 vdd.n1577 52.4337
R3480 vdd.n1658 vdd.n1578 52.4337
R3481 vdd.n1660 vdd.n1579 52.4337
R3482 vdd.n1664 vdd.n1580 52.4337
R3483 vdd.n1666 vdd.n1581 52.4337
R3484 vdd.n1670 vdd.n1582 52.4337
R3485 vdd.n1672 vdd.n1583 52.4337
R3486 vdd.n1676 vdd.n1584 52.4337
R3487 vdd.n1678 vdd.n1585 52.4337
R3488 vdd.n1433 vdd.n1432 52.4337
R3489 vdd.n1430 vdd.n1429 52.4337
R3490 vdd.n1426 vdd.n1218 52.4337
R3491 vdd.n2280 vdd.n2279 52.4337
R3492 vdd.n1217 vdd.n1211 52.4337
R3493 vdd.n2287 vdd.n2286 52.4337
R3494 vdd.n1210 vdd.n1204 52.4337
R3495 vdd.n2294 vdd.n2293 52.4337
R3496 vdd.n1203 vdd.n1198 52.4337
R3497 vdd.n2301 vdd.n2300 52.4337
R3498 vdd.n1197 vdd.n1196 52.4337
R3499 vdd.n1192 vdd.n1185 52.4337
R3500 vdd.n2312 vdd.n2311 52.4337
R3501 vdd.n1184 vdd.n1178 52.4337
R3502 vdd.n2319 vdd.n2318 52.4337
R3503 vdd.n1177 vdd.n1171 52.4337
R3504 vdd.n2326 vdd.n2325 52.4337
R3505 vdd.n1170 vdd.n1164 52.4337
R3506 vdd.n2333 vdd.n2332 52.4337
R3507 vdd.n1163 vdd.n1158 52.4337
R3508 vdd.n2340 vdd.n2339 52.4337
R3509 vdd.n1157 vdd.n1156 52.4337
R3510 vdd.n1152 vdd.n1145 52.4337
R3511 vdd.n2351 vdd.n2350 52.4337
R3512 vdd.n1144 vdd.n1138 52.4337
R3513 vdd.n2358 vdd.n2357 52.4337
R3514 vdd.n1137 vdd.n1131 52.4337
R3515 vdd.n2365 vdd.n2364 52.4337
R3516 vdd.n1130 vdd.n1127 52.4337
R3517 vdd.n2372 vdd.n2371 52.4337
R3518 vdd.n2377 vdd.n2376 52.4337
R3519 vdd.n1437 vdd.n1126 52.4337
R3520 vdd.n3314 vdd.n725 52.4337
R3521 vdd.n733 vdd.n693 52.4337
R3522 vdd.n3304 vdd.n694 52.4337
R3523 vdd.n3300 vdd.n695 52.4337
R3524 vdd.n3296 vdd.n696 52.4337
R3525 vdd.n3292 vdd.n697 52.4337
R3526 vdd.n3288 vdd.n698 52.4337
R3527 vdd.n3284 vdd.n699 52.4337
R3528 vdd.n3280 vdd.n700 52.4337
R3529 vdd.n3270 vdd.n701 52.4337
R3530 vdd.n3268 vdd.n702 52.4337
R3531 vdd.n3264 vdd.n703 52.4337
R3532 vdd.n3260 vdd.n704 52.4337
R3533 vdd.n3256 vdd.n705 52.4337
R3534 vdd.n3252 vdd.n706 52.4337
R3535 vdd.n3248 vdd.n707 52.4337
R3536 vdd.n3244 vdd.n708 52.4337
R3537 vdd.n3240 vdd.n709 52.4337
R3538 vdd.n3236 vdd.n710 52.4337
R3539 vdd.n3232 vdd.n711 52.4337
R3540 vdd.n3224 vdd.n712 52.4337
R3541 vdd.n3222 vdd.n713 52.4337
R3542 vdd.n3218 vdd.n714 52.4337
R3543 vdd.n3214 vdd.n715 52.4337
R3544 vdd.n3210 vdd.n716 52.4337
R3545 vdd.n3206 vdd.n717 52.4337
R3546 vdd.n3202 vdd.n718 52.4337
R3547 vdd.n3198 vdd.n719 52.4337
R3548 vdd.n3194 vdd.n720 52.4337
R3549 vdd.n3190 vdd.n721 52.4337
R3550 vdd.n722 vdd.n691 52.4337
R3551 vdd.n3445 vdd.n425 52.4337
R3552 vdd.n614 vdd.n424 52.4337
R3553 vdd.n608 vdd.n423 52.4337
R3554 vdd.n604 vdd.n422 52.4337
R3555 vdd.n598 vdd.n421 52.4337
R3556 vdd.n594 vdd.n420 52.4337
R3557 vdd.n588 vdd.n419 52.4337
R3558 vdd.n584 vdd.n418 52.4337
R3559 vdd.n578 vdd.n417 52.4337
R3560 vdd.n574 vdd.n416 52.4337
R3561 vdd.n568 vdd.n415 52.4337
R3562 vdd.n564 vdd.n414 52.4337
R3563 vdd.n558 vdd.n413 52.4337
R3564 vdd.n554 vdd.n412 52.4337
R3565 vdd.n548 vdd.n411 52.4337
R3566 vdd.n544 vdd.n410 52.4337
R3567 vdd.n538 vdd.n409 52.4337
R3568 vdd.n534 vdd.n408 52.4337
R3569 vdd.n528 vdd.n407 52.4337
R3570 vdd.n524 vdd.n406 52.4337
R3571 vdd.n518 vdd.n405 52.4337
R3572 vdd.n514 vdd.n404 52.4337
R3573 vdd.n508 vdd.n403 52.4337
R3574 vdd.n504 vdd.n402 52.4337
R3575 vdd.n498 vdd.n401 52.4337
R3576 vdd.n494 vdd.n400 52.4337
R3577 vdd.n488 vdd.n399 52.4337
R3578 vdd.n484 vdd.n398 52.4337
R3579 vdd.n478 vdd.n397 52.4337
R3580 vdd.n474 vdd.n396 52.4337
R3581 vdd.n468 vdd.n395 52.4337
R3582 vdd.n394 vdd.n392 52.4337
R3583 vdd.t22 vdd.t130 51.4683
R3584 vdd.n274 vdd.n272 42.0461
R3585 vdd.n172 vdd.n170 42.0461
R3586 vdd.n71 vdd.n69 42.0461
R3587 vdd.n2114 vdd.n2112 42.0461
R3588 vdd.n2012 vdd.n2010 42.0461
R3589 vdd.n1911 vdd.n1909 42.0461
R3590 vdd.n332 vdd.n331 41.6884
R3591 vdd.n230 vdd.n229 41.6884
R3592 vdd.n129 vdd.n128 41.6884
R3593 vdd.n2172 vdd.n2171 41.6884
R3594 vdd.n2070 vdd.n2069 41.6884
R3595 vdd.n1969 vdd.n1968 41.6884
R3596 vdd.n1681 vdd.n1680 41.1157
R3597 vdd.n1719 vdd.n1718 41.1157
R3598 vdd.n1615 vdd.n1614 41.1157
R3599 vdd.n428 vdd.n427 41.1157
R3600 vdd.n566 vdd.n441 41.1157
R3601 vdd.n454 vdd.n453 41.1157
R3602 vdd.n3145 vdd.n3144 39.2114
R3603 vdd.n3142 vdd.n3141 39.2114
R3604 vdd.n3137 vdd.n815 39.2114
R3605 vdd.n3135 vdd.n3134 39.2114
R3606 vdd.n3130 vdd.n818 39.2114
R3607 vdd.n3128 vdd.n3127 39.2114
R3608 vdd.n3123 vdd.n821 39.2114
R3609 vdd.n3121 vdd.n3120 39.2114
R3610 vdd.n3117 vdd.n3116 39.2114
R3611 vdd.n3112 vdd.n824 39.2114
R3612 vdd.n3110 vdd.n3109 39.2114
R3613 vdd.n3105 vdd.n827 39.2114
R3614 vdd.n3103 vdd.n3102 39.2114
R3615 vdd.n3098 vdd.n830 39.2114
R3616 vdd.n3096 vdd.n3095 39.2114
R3617 vdd.n3090 vdd.n835 39.2114
R3618 vdd.n3088 vdd.n3087 39.2114
R3619 vdd.n2937 vdd.n2936 39.2114
R3620 vdd.n2931 vdd.n2666 39.2114
R3621 vdd.n2928 vdd.n2667 39.2114
R3622 vdd.n2924 vdd.n2668 39.2114
R3623 vdd.n2920 vdd.n2669 39.2114
R3624 vdd.n2916 vdd.n2670 39.2114
R3625 vdd.n2912 vdd.n2671 39.2114
R3626 vdd.n2908 vdd.n2672 39.2114
R3627 vdd.n2904 vdd.n2673 39.2114
R3628 vdd.n2900 vdd.n2674 39.2114
R3629 vdd.n2896 vdd.n2675 39.2114
R3630 vdd.n2892 vdd.n2676 39.2114
R3631 vdd.n2888 vdd.n2677 39.2114
R3632 vdd.n2884 vdd.n2678 39.2114
R3633 vdd.n2880 vdd.n2679 39.2114
R3634 vdd.n2876 vdd.n2680 39.2114
R3635 vdd.n2871 vdd.n2681 39.2114
R3636 vdd.n2660 vdd.n968 39.2114
R3637 vdd.n2656 vdd.n967 39.2114
R3638 vdd.n2652 vdd.n966 39.2114
R3639 vdd.n2648 vdd.n965 39.2114
R3640 vdd.n2644 vdd.n964 39.2114
R3641 vdd.n2640 vdd.n963 39.2114
R3642 vdd.n2636 vdd.n962 39.2114
R3643 vdd.n2632 vdd.n961 39.2114
R3644 vdd.n2628 vdd.n960 39.2114
R3645 vdd.n2624 vdd.n959 39.2114
R3646 vdd.n2620 vdd.n958 39.2114
R3647 vdd.n2616 vdd.n957 39.2114
R3648 vdd.n2612 vdd.n956 39.2114
R3649 vdd.n2608 vdd.n955 39.2114
R3650 vdd.n2604 vdd.n954 39.2114
R3651 vdd.n2599 vdd.n953 39.2114
R3652 vdd.n2595 vdd.n952 39.2114
R3653 vdd.n2416 vdd.n2415 39.2114
R3654 vdd.n2410 vdd.n1084 39.2114
R3655 vdd.n2407 vdd.n1085 39.2114
R3656 vdd.n2403 vdd.n1086 39.2114
R3657 vdd.n2399 vdd.n1087 39.2114
R3658 vdd.n2395 vdd.n1088 39.2114
R3659 vdd.n2391 vdd.n1089 39.2114
R3660 vdd.n2387 vdd.n1090 39.2114
R3661 vdd.n2383 vdd.n1091 39.2114
R3662 vdd.n1276 vdd.n1092 39.2114
R3663 vdd.n1280 vdd.n1093 39.2114
R3664 vdd.n1284 vdd.n1094 39.2114
R3665 vdd.n1288 vdd.n1095 39.2114
R3666 vdd.n1292 vdd.n1096 39.2114
R3667 vdd.n1296 vdd.n1097 39.2114
R3668 vdd.n1300 vdd.n1098 39.2114
R3669 vdd.n1305 vdd.n1099 39.2114
R3670 vdd.n3064 vdd.n3063 39.2114
R3671 vdd.n3059 vdd.n3031 39.2114
R3672 vdd.n3057 vdd.n3056 39.2114
R3673 vdd.n3052 vdd.n3034 39.2114
R3674 vdd.n3050 vdd.n3049 39.2114
R3675 vdd.n3045 vdd.n3037 39.2114
R3676 vdd.n3043 vdd.n3042 39.2114
R3677 vdd.n3038 vdd.n787 39.2114
R3678 vdd.n3182 vdd.n3181 39.2114
R3679 vdd.n3179 vdd.n3178 39.2114
R3680 vdd.n3174 vdd.n791 39.2114
R3681 vdd.n3172 vdd.n3171 39.2114
R3682 vdd.n3167 vdd.n794 39.2114
R3683 vdd.n3165 vdd.n3164 39.2114
R3684 vdd.n3160 vdd.n797 39.2114
R3685 vdd.n3158 vdd.n3157 39.2114
R3686 vdd.n3153 vdd.n803 39.2114
R3687 vdd.n2940 vdd.n2939 39.2114
R3688 vdd.n2707 vdd.n2682 39.2114
R3689 vdd.n2711 vdd.n2683 39.2114
R3690 vdd.n2715 vdd.n2684 39.2114
R3691 vdd.n2719 vdd.n2685 39.2114
R3692 vdd.n2723 vdd.n2686 39.2114
R3693 vdd.n2727 vdd.n2687 39.2114
R3694 vdd.n2731 vdd.n2688 39.2114
R3695 vdd.n2735 vdd.n2689 39.2114
R3696 vdd.n2739 vdd.n2690 39.2114
R3697 vdd.n2743 vdd.n2691 39.2114
R3698 vdd.n2747 vdd.n2692 39.2114
R3699 vdd.n2751 vdd.n2693 39.2114
R3700 vdd.n2755 vdd.n2694 39.2114
R3701 vdd.n2759 vdd.n2695 39.2114
R3702 vdd.n2763 vdd.n2696 39.2114
R3703 vdd.n2767 vdd.n2697 39.2114
R3704 vdd.n2939 vdd.n933 39.2114
R3705 vdd.n2710 vdd.n2682 39.2114
R3706 vdd.n2714 vdd.n2683 39.2114
R3707 vdd.n2718 vdd.n2684 39.2114
R3708 vdd.n2722 vdd.n2685 39.2114
R3709 vdd.n2726 vdd.n2686 39.2114
R3710 vdd.n2730 vdd.n2687 39.2114
R3711 vdd.n2734 vdd.n2688 39.2114
R3712 vdd.n2738 vdd.n2689 39.2114
R3713 vdd.n2742 vdd.n2690 39.2114
R3714 vdd.n2746 vdd.n2691 39.2114
R3715 vdd.n2750 vdd.n2692 39.2114
R3716 vdd.n2754 vdd.n2693 39.2114
R3717 vdd.n2758 vdd.n2694 39.2114
R3718 vdd.n2762 vdd.n2695 39.2114
R3719 vdd.n2766 vdd.n2696 39.2114
R3720 vdd.n2769 vdd.n2697 39.2114
R3721 vdd.n803 vdd.n798 39.2114
R3722 vdd.n3159 vdd.n3158 39.2114
R3723 vdd.n797 vdd.n795 39.2114
R3724 vdd.n3166 vdd.n3165 39.2114
R3725 vdd.n794 vdd.n792 39.2114
R3726 vdd.n3173 vdd.n3172 39.2114
R3727 vdd.n791 vdd.n789 39.2114
R3728 vdd.n3180 vdd.n3179 39.2114
R3729 vdd.n3183 vdd.n3182 39.2114
R3730 vdd.n3039 vdd.n3038 39.2114
R3731 vdd.n3044 vdd.n3043 39.2114
R3732 vdd.n3037 vdd.n3035 39.2114
R3733 vdd.n3051 vdd.n3050 39.2114
R3734 vdd.n3034 vdd.n3032 39.2114
R3735 vdd.n3058 vdd.n3057 39.2114
R3736 vdd.n3031 vdd.n3029 39.2114
R3737 vdd.n3065 vdd.n3064 39.2114
R3738 vdd.n2416 vdd.n1118 39.2114
R3739 vdd.n2408 vdd.n1084 39.2114
R3740 vdd.n2404 vdd.n1085 39.2114
R3741 vdd.n2400 vdd.n1086 39.2114
R3742 vdd.n2396 vdd.n1087 39.2114
R3743 vdd.n2392 vdd.n1088 39.2114
R3744 vdd.n2388 vdd.n1089 39.2114
R3745 vdd.n2384 vdd.n1090 39.2114
R3746 vdd.n1275 vdd.n1091 39.2114
R3747 vdd.n1279 vdd.n1092 39.2114
R3748 vdd.n1283 vdd.n1093 39.2114
R3749 vdd.n1287 vdd.n1094 39.2114
R3750 vdd.n1291 vdd.n1095 39.2114
R3751 vdd.n1295 vdd.n1096 39.2114
R3752 vdd.n1299 vdd.n1097 39.2114
R3753 vdd.n1304 vdd.n1098 39.2114
R3754 vdd.n1308 vdd.n1099 39.2114
R3755 vdd.n2598 vdd.n952 39.2114
R3756 vdd.n2603 vdd.n953 39.2114
R3757 vdd.n2607 vdd.n954 39.2114
R3758 vdd.n2611 vdd.n955 39.2114
R3759 vdd.n2615 vdd.n956 39.2114
R3760 vdd.n2619 vdd.n957 39.2114
R3761 vdd.n2623 vdd.n958 39.2114
R3762 vdd.n2627 vdd.n959 39.2114
R3763 vdd.n2631 vdd.n960 39.2114
R3764 vdd.n2635 vdd.n961 39.2114
R3765 vdd.n2639 vdd.n962 39.2114
R3766 vdd.n2643 vdd.n963 39.2114
R3767 vdd.n2647 vdd.n964 39.2114
R3768 vdd.n2651 vdd.n965 39.2114
R3769 vdd.n2655 vdd.n966 39.2114
R3770 vdd.n2659 vdd.n967 39.2114
R3771 vdd.n970 vdd.n968 39.2114
R3772 vdd.n2937 vdd.n2700 39.2114
R3773 vdd.n2929 vdd.n2666 39.2114
R3774 vdd.n2925 vdd.n2667 39.2114
R3775 vdd.n2921 vdd.n2668 39.2114
R3776 vdd.n2917 vdd.n2669 39.2114
R3777 vdd.n2913 vdd.n2670 39.2114
R3778 vdd.n2909 vdd.n2671 39.2114
R3779 vdd.n2905 vdd.n2672 39.2114
R3780 vdd.n2901 vdd.n2673 39.2114
R3781 vdd.n2897 vdd.n2674 39.2114
R3782 vdd.n2893 vdd.n2675 39.2114
R3783 vdd.n2889 vdd.n2676 39.2114
R3784 vdd.n2885 vdd.n2677 39.2114
R3785 vdd.n2881 vdd.n2678 39.2114
R3786 vdd.n2877 vdd.n2679 39.2114
R3787 vdd.n2872 vdd.n2680 39.2114
R3788 vdd.n2868 vdd.n2681 39.2114
R3789 vdd.n3089 vdd.n3088 39.2114
R3790 vdd.n835 vdd.n831 39.2114
R3791 vdd.n3097 vdd.n3096 39.2114
R3792 vdd.n830 vdd.n828 39.2114
R3793 vdd.n3104 vdd.n3103 39.2114
R3794 vdd.n827 vdd.n825 39.2114
R3795 vdd.n3111 vdd.n3110 39.2114
R3796 vdd.n824 vdd.n822 39.2114
R3797 vdd.n3118 vdd.n3117 39.2114
R3798 vdd.n3122 vdd.n3121 39.2114
R3799 vdd.n821 vdd.n819 39.2114
R3800 vdd.n3129 vdd.n3128 39.2114
R3801 vdd.n818 vdd.n816 39.2114
R3802 vdd.n3136 vdd.n3135 39.2114
R3803 vdd.n815 vdd.n813 39.2114
R3804 vdd.n3143 vdd.n3142 39.2114
R3805 vdd.n3146 vdd.n3145 39.2114
R3806 vdd.n979 vdd.n934 39.2114
R3807 vdd.n2587 vdd.n935 39.2114
R3808 vdd.n2583 vdd.n936 39.2114
R3809 vdd.n2579 vdd.n937 39.2114
R3810 vdd.n2575 vdd.n938 39.2114
R3811 vdd.n2571 vdd.n939 39.2114
R3812 vdd.n2567 vdd.n940 39.2114
R3813 vdd.n2563 vdd.n941 39.2114
R3814 vdd.n2559 vdd.n942 39.2114
R3815 vdd.n2555 vdd.n943 39.2114
R3816 vdd.n2551 vdd.n944 39.2114
R3817 vdd.n2547 vdd.n945 39.2114
R3818 vdd.n2543 vdd.n946 39.2114
R3819 vdd.n2539 vdd.n947 39.2114
R3820 vdd.n2535 vdd.n948 39.2114
R3821 vdd.n2531 vdd.n949 39.2114
R3822 vdd.n2527 vdd.n950 39.2114
R3823 vdd.n2419 vdd.n2418 39.2114
R3824 vdd.n1222 vdd.n1100 39.2114
R3825 vdd.n1226 vdd.n1101 39.2114
R3826 vdd.n1230 vdd.n1102 39.2114
R3827 vdd.n1234 vdd.n1103 39.2114
R3828 vdd.n1238 vdd.n1104 39.2114
R3829 vdd.n1242 vdd.n1105 39.2114
R3830 vdd.n1246 vdd.n1106 39.2114
R3831 vdd.n1250 vdd.n1107 39.2114
R3832 vdd.n1420 vdd.n1108 39.2114
R3833 vdd.n1417 vdd.n1109 39.2114
R3834 vdd.n1413 vdd.n1110 39.2114
R3835 vdd.n1409 vdd.n1111 39.2114
R3836 vdd.n1405 vdd.n1112 39.2114
R3837 vdd.n1401 vdd.n1113 39.2114
R3838 vdd.n1397 vdd.n1114 39.2114
R3839 vdd.n1393 vdd.n1115 39.2114
R3840 vdd.n2524 vdd.n950 39.2114
R3841 vdd.n2528 vdd.n949 39.2114
R3842 vdd.n2532 vdd.n948 39.2114
R3843 vdd.n2536 vdd.n947 39.2114
R3844 vdd.n2540 vdd.n946 39.2114
R3845 vdd.n2544 vdd.n945 39.2114
R3846 vdd.n2548 vdd.n944 39.2114
R3847 vdd.n2552 vdd.n943 39.2114
R3848 vdd.n2556 vdd.n942 39.2114
R3849 vdd.n2560 vdd.n941 39.2114
R3850 vdd.n2564 vdd.n940 39.2114
R3851 vdd.n2568 vdd.n939 39.2114
R3852 vdd.n2572 vdd.n938 39.2114
R3853 vdd.n2576 vdd.n937 39.2114
R3854 vdd.n2580 vdd.n936 39.2114
R3855 vdd.n2584 vdd.n935 39.2114
R3856 vdd.n2588 vdd.n934 39.2114
R3857 vdd.n2418 vdd.n1082 39.2114
R3858 vdd.n1225 vdd.n1100 39.2114
R3859 vdd.n1229 vdd.n1101 39.2114
R3860 vdd.n1233 vdd.n1102 39.2114
R3861 vdd.n1237 vdd.n1103 39.2114
R3862 vdd.n1241 vdd.n1104 39.2114
R3863 vdd.n1245 vdd.n1105 39.2114
R3864 vdd.n1249 vdd.n1106 39.2114
R3865 vdd.n1252 vdd.n1107 39.2114
R3866 vdd.n1418 vdd.n1108 39.2114
R3867 vdd.n1414 vdd.n1109 39.2114
R3868 vdd.n1410 vdd.n1110 39.2114
R3869 vdd.n1406 vdd.n1111 39.2114
R3870 vdd.n1402 vdd.n1112 39.2114
R3871 vdd.n1398 vdd.n1113 39.2114
R3872 vdd.n1394 vdd.n1114 39.2114
R3873 vdd.n1390 vdd.n1115 39.2114
R3874 vdd.n2271 vdd.n2270 37.2369
R3875 vdd.n2307 vdd.n1191 37.2369
R3876 vdd.n2346 vdd.n1151 37.2369
R3877 vdd.n3230 vdd.n769 37.2369
R3878 vdd.n3278 vdd.n3277 37.2369
R3879 vdd.n690 vdd.n689 37.2369
R3880 vdd.n2414 vdd.n1074 31.0639
R3881 vdd.n2663 vdd.n971 31.0639
R3882 vdd.n2596 vdd.n974 31.0639
R3883 vdd.n1310 vdd.n1307 31.0639
R3884 vdd.n2869 vdd.n2866 31.0639
R3885 vdd.n3086 vdd.n3085 31.0639
R3886 vdd.n2935 vdd.n926 31.0639
R3887 vdd.n3149 vdd.n3148 31.0639
R3888 vdd.n3068 vdd.n3067 31.0639
R3889 vdd.n3154 vdd.n802 31.0639
R3890 vdd.n2773 vdd.n2771 31.0639
R3891 vdd.n2942 vdd.n2941 31.0639
R3892 vdd.n2421 vdd.n2420 31.0639
R3893 vdd.n2591 vdd.n2590 31.0639
R3894 vdd.n2523 vdd.n2522 31.0639
R3895 vdd.n1389 vdd.n1388 31.0639
R3896 vdd.n1255 vdd.n1254 30.449
R3897 vdd.n983 vdd.n982 30.449
R3898 vdd.n1302 vdd.n1274 30.449
R3899 vdd.n2601 vdd.n973 30.449
R3900 vdd.n2706 vdd.n2705 30.449
R3901 vdd.n3092 vdd.n833 30.449
R3902 vdd.n2874 vdd.n2702 30.449
R3903 vdd.n801 vdd.n800 30.449
R3904 vdd.n1780 vdd.n1587 22.2201
R3905 vdd.n2265 vdd.n1083 22.2201
R3906 vdd.n3315 vdd.n723 22.2201
R3907 vdd.n3447 vdd.n3446 22.2201
R3908 vdd.n1791 vdd.n1549 19.3944
R3909 vdd.n1791 vdd.n1547 19.3944
R3910 vdd.n1795 vdd.n1547 19.3944
R3911 vdd.n1795 vdd.n1537 19.3944
R3912 vdd.n1808 vdd.n1537 19.3944
R3913 vdd.n1808 vdd.n1535 19.3944
R3914 vdd.n1812 vdd.n1535 19.3944
R3915 vdd.n1812 vdd.n1527 19.3944
R3916 vdd.n1825 vdd.n1527 19.3944
R3917 vdd.n1825 vdd.n1525 19.3944
R3918 vdd.n1829 vdd.n1525 19.3944
R3919 vdd.n1829 vdd.n1514 19.3944
R3920 vdd.n1841 vdd.n1514 19.3944
R3921 vdd.n1841 vdd.n1512 19.3944
R3922 vdd.n1845 vdd.n1512 19.3944
R3923 vdd.n1845 vdd.n1503 19.3944
R3924 vdd.n1858 vdd.n1503 19.3944
R3925 vdd.n1858 vdd.n1501 19.3944
R3926 vdd.n1862 vdd.n1501 19.3944
R3927 vdd.n1862 vdd.n1492 19.3944
R3928 vdd.n2181 vdd.n1492 19.3944
R3929 vdd.n2181 vdd.n1490 19.3944
R3930 vdd.n2185 vdd.n1490 19.3944
R3931 vdd.n2185 vdd.n1480 19.3944
R3932 vdd.n2198 vdd.n1480 19.3944
R3933 vdd.n2198 vdd.n1478 19.3944
R3934 vdd.n2202 vdd.n1478 19.3944
R3935 vdd.n2202 vdd.n1470 19.3944
R3936 vdd.n2215 vdd.n1470 19.3944
R3937 vdd.n2215 vdd.n1468 19.3944
R3938 vdd.n2219 vdd.n1468 19.3944
R3939 vdd.n2219 vdd.n1457 19.3944
R3940 vdd.n2231 vdd.n1457 19.3944
R3941 vdd.n2231 vdd.n1455 19.3944
R3942 vdd.n2235 vdd.n1455 19.3944
R3943 vdd.n2235 vdd.n1447 19.3944
R3944 vdd.n2248 vdd.n1447 19.3944
R3945 vdd.n2248 vdd.n1444 19.3944
R3946 vdd.n2254 vdd.n1444 19.3944
R3947 vdd.n2254 vdd.n1445 19.3944
R3948 vdd.n1445 vdd.n1435 19.3944
R3949 vdd.n1715 vdd.n1650 19.3944
R3950 vdd.n1711 vdd.n1650 19.3944
R3951 vdd.n1711 vdd.n1710 19.3944
R3952 vdd.n1710 vdd.n1709 19.3944
R3953 vdd.n1709 vdd.n1656 19.3944
R3954 vdd.n1705 vdd.n1656 19.3944
R3955 vdd.n1705 vdd.n1704 19.3944
R3956 vdd.n1704 vdd.n1703 19.3944
R3957 vdd.n1703 vdd.n1662 19.3944
R3958 vdd.n1699 vdd.n1662 19.3944
R3959 vdd.n1699 vdd.n1698 19.3944
R3960 vdd.n1698 vdd.n1697 19.3944
R3961 vdd.n1697 vdd.n1668 19.3944
R3962 vdd.n1693 vdd.n1668 19.3944
R3963 vdd.n1693 vdd.n1692 19.3944
R3964 vdd.n1692 vdd.n1691 19.3944
R3965 vdd.n1691 vdd.n1674 19.3944
R3966 vdd.n1687 vdd.n1674 19.3944
R3967 vdd.n1687 vdd.n1686 19.3944
R3968 vdd.n1686 vdd.n1685 19.3944
R3969 vdd.n1750 vdd.n1749 19.3944
R3970 vdd.n1749 vdd.n1748 19.3944
R3971 vdd.n1748 vdd.n1621 19.3944
R3972 vdd.n1744 vdd.n1621 19.3944
R3973 vdd.n1744 vdd.n1743 19.3944
R3974 vdd.n1743 vdd.n1742 19.3944
R3975 vdd.n1742 vdd.n1627 19.3944
R3976 vdd.n1738 vdd.n1627 19.3944
R3977 vdd.n1738 vdd.n1737 19.3944
R3978 vdd.n1737 vdd.n1736 19.3944
R3979 vdd.n1736 vdd.n1633 19.3944
R3980 vdd.n1732 vdd.n1633 19.3944
R3981 vdd.n1732 vdd.n1731 19.3944
R3982 vdd.n1731 vdd.n1730 19.3944
R3983 vdd.n1730 vdd.n1639 19.3944
R3984 vdd.n1726 vdd.n1639 19.3944
R3985 vdd.n1726 vdd.n1725 19.3944
R3986 vdd.n1725 vdd.n1724 19.3944
R3987 vdd.n1724 vdd.n1645 19.3944
R3988 vdd.n1720 vdd.n1645 19.3944
R3989 vdd.n1783 vdd.n1554 19.3944
R3990 vdd.n1778 vdd.n1554 19.3944
R3991 vdd.n1778 vdd.n1589 19.3944
R3992 vdd.n1774 vdd.n1589 19.3944
R3993 vdd.n1774 vdd.n1773 19.3944
R3994 vdd.n1773 vdd.n1772 19.3944
R3995 vdd.n1772 vdd.n1595 19.3944
R3996 vdd.n1768 vdd.n1595 19.3944
R3997 vdd.n1768 vdd.n1767 19.3944
R3998 vdd.n1767 vdd.n1766 19.3944
R3999 vdd.n1766 vdd.n1601 19.3944
R4000 vdd.n1762 vdd.n1601 19.3944
R4001 vdd.n1762 vdd.n1761 19.3944
R4002 vdd.n1761 vdd.n1760 19.3944
R4003 vdd.n1760 vdd.n1607 19.3944
R4004 vdd.n1756 vdd.n1607 19.3944
R4005 vdd.n1756 vdd.n1755 19.3944
R4006 vdd.n1755 vdd.n1754 19.3944
R4007 vdd.n2303 vdd.n1189 19.3944
R4008 vdd.n2303 vdd.n1195 19.3944
R4009 vdd.n2298 vdd.n1195 19.3944
R4010 vdd.n2298 vdd.n2297 19.3944
R4011 vdd.n2297 vdd.n2296 19.3944
R4012 vdd.n2296 vdd.n1202 19.3944
R4013 vdd.n2291 vdd.n1202 19.3944
R4014 vdd.n2291 vdd.n2290 19.3944
R4015 vdd.n2290 vdd.n2289 19.3944
R4016 vdd.n2289 vdd.n1209 19.3944
R4017 vdd.n2284 vdd.n1209 19.3944
R4018 vdd.n2284 vdd.n2283 19.3944
R4019 vdd.n2283 vdd.n2282 19.3944
R4020 vdd.n2282 vdd.n1216 19.3944
R4021 vdd.n2277 vdd.n1216 19.3944
R4022 vdd.n2277 vdd.n2276 19.3944
R4023 vdd.n1428 vdd.n1221 19.3944
R4024 vdd.n2272 vdd.n1425 19.3944
R4025 vdd.n2342 vdd.n1149 19.3944
R4026 vdd.n2342 vdd.n1155 19.3944
R4027 vdd.n2337 vdd.n1155 19.3944
R4028 vdd.n2337 vdd.n2336 19.3944
R4029 vdd.n2336 vdd.n2335 19.3944
R4030 vdd.n2335 vdd.n1162 19.3944
R4031 vdd.n2330 vdd.n1162 19.3944
R4032 vdd.n2330 vdd.n2329 19.3944
R4033 vdd.n2329 vdd.n2328 19.3944
R4034 vdd.n2328 vdd.n1169 19.3944
R4035 vdd.n2323 vdd.n1169 19.3944
R4036 vdd.n2323 vdd.n2322 19.3944
R4037 vdd.n2322 vdd.n2321 19.3944
R4038 vdd.n2321 vdd.n1176 19.3944
R4039 vdd.n2316 vdd.n1176 19.3944
R4040 vdd.n2316 vdd.n2315 19.3944
R4041 vdd.n2315 vdd.n2314 19.3944
R4042 vdd.n2314 vdd.n1183 19.3944
R4043 vdd.n2309 vdd.n1183 19.3944
R4044 vdd.n2309 vdd.n2308 19.3944
R4045 vdd.n2379 vdd.n1124 19.3944
R4046 vdd.n2379 vdd.n1125 19.3944
R4047 vdd.n2374 vdd.n2373 19.3944
R4048 vdd.n2369 vdd.n2368 19.3944
R4049 vdd.n2368 vdd.n2367 19.3944
R4050 vdd.n2367 vdd.n1129 19.3944
R4051 vdd.n2362 vdd.n1129 19.3944
R4052 vdd.n2362 vdd.n2361 19.3944
R4053 vdd.n2361 vdd.n2360 19.3944
R4054 vdd.n2360 vdd.n1136 19.3944
R4055 vdd.n2355 vdd.n1136 19.3944
R4056 vdd.n2355 vdd.n2354 19.3944
R4057 vdd.n2354 vdd.n2353 19.3944
R4058 vdd.n2353 vdd.n1143 19.3944
R4059 vdd.n2348 vdd.n1143 19.3944
R4060 vdd.n2348 vdd.n2347 19.3944
R4061 vdd.n1787 vdd.n1552 19.3944
R4062 vdd.n1787 vdd.n1543 19.3944
R4063 vdd.n1800 vdd.n1543 19.3944
R4064 vdd.n1800 vdd.n1541 19.3944
R4065 vdd.n1804 vdd.n1541 19.3944
R4066 vdd.n1804 vdd.n1532 19.3944
R4067 vdd.n1817 vdd.n1532 19.3944
R4068 vdd.n1817 vdd.n1530 19.3944
R4069 vdd.n1821 vdd.n1530 19.3944
R4070 vdd.n1821 vdd.n1521 19.3944
R4071 vdd.n1833 vdd.n1521 19.3944
R4072 vdd.n1833 vdd.n1519 19.3944
R4073 vdd.n1837 vdd.n1519 19.3944
R4074 vdd.n1837 vdd.n1509 19.3944
R4075 vdd.n1850 vdd.n1509 19.3944
R4076 vdd.n1850 vdd.n1507 19.3944
R4077 vdd.n1854 vdd.n1507 19.3944
R4078 vdd.n1854 vdd.n1498 19.3944
R4079 vdd.n1866 vdd.n1498 19.3944
R4080 vdd.n1866 vdd.n1496 19.3944
R4081 vdd.n2177 vdd.n1496 19.3944
R4082 vdd.n2177 vdd.n1486 19.3944
R4083 vdd.n2190 vdd.n1486 19.3944
R4084 vdd.n2190 vdd.n1484 19.3944
R4085 vdd.n2194 vdd.n1484 19.3944
R4086 vdd.n2194 vdd.n1475 19.3944
R4087 vdd.n2207 vdd.n1475 19.3944
R4088 vdd.n2207 vdd.n1473 19.3944
R4089 vdd.n2211 vdd.n1473 19.3944
R4090 vdd.n2211 vdd.n1464 19.3944
R4091 vdd.n2223 vdd.n1464 19.3944
R4092 vdd.n2223 vdd.n1462 19.3944
R4093 vdd.n2227 vdd.n1462 19.3944
R4094 vdd.n2227 vdd.n1452 19.3944
R4095 vdd.n2240 vdd.n1452 19.3944
R4096 vdd.n2240 vdd.n1450 19.3944
R4097 vdd.n2244 vdd.n1450 19.3944
R4098 vdd.n2244 vdd.n1440 19.3944
R4099 vdd.n2259 vdd.n1440 19.3944
R4100 vdd.n2259 vdd.n1438 19.3944
R4101 vdd.n2263 vdd.n1438 19.3944
R4102 vdd.n3321 vdd.n686 19.3944
R4103 vdd.n3321 vdd.n676 19.3944
R4104 vdd.n3333 vdd.n676 19.3944
R4105 vdd.n3333 vdd.n674 19.3944
R4106 vdd.n3337 vdd.n674 19.3944
R4107 vdd.n3337 vdd.n666 19.3944
R4108 vdd.n3350 vdd.n666 19.3944
R4109 vdd.n3350 vdd.n664 19.3944
R4110 vdd.n3354 vdd.n664 19.3944
R4111 vdd.n3354 vdd.n653 19.3944
R4112 vdd.n3366 vdd.n653 19.3944
R4113 vdd.n3366 vdd.n651 19.3944
R4114 vdd.n3370 vdd.n651 19.3944
R4115 vdd.n3370 vdd.n642 19.3944
R4116 vdd.n3383 vdd.n642 19.3944
R4117 vdd.n3383 vdd.n640 19.3944
R4118 vdd.n3390 vdd.n640 19.3944
R4119 vdd.n3390 vdd.n3389 19.3944
R4120 vdd.n3389 vdd.n631 19.3944
R4121 vdd.n3403 vdd.n631 19.3944
R4122 vdd.n3404 vdd.n3403 19.3944
R4123 vdd.n3404 vdd.n629 19.3944
R4124 vdd.n3408 vdd.n629 19.3944
R4125 vdd.n3410 vdd.n3408 19.3944
R4126 vdd.n3411 vdd.n3410 19.3944
R4127 vdd.n3411 vdd.n627 19.3944
R4128 vdd.n3415 vdd.n627 19.3944
R4129 vdd.n3417 vdd.n3415 19.3944
R4130 vdd.n3418 vdd.n3417 19.3944
R4131 vdd.n3418 vdd.n625 19.3944
R4132 vdd.n3422 vdd.n625 19.3944
R4133 vdd.n3425 vdd.n3422 19.3944
R4134 vdd.n3426 vdd.n3425 19.3944
R4135 vdd.n3426 vdd.n623 19.3944
R4136 vdd.n3430 vdd.n623 19.3944
R4137 vdd.n3432 vdd.n3430 19.3944
R4138 vdd.n3433 vdd.n3432 19.3944
R4139 vdd.n3433 vdd.n621 19.3944
R4140 vdd.n3437 vdd.n621 19.3944
R4141 vdd.n3439 vdd.n3437 19.3944
R4142 vdd.n3440 vdd.n3439 19.3944
R4143 vdd.n569 vdd.n438 19.3944
R4144 vdd.n575 vdd.n438 19.3944
R4145 vdd.n576 vdd.n575 19.3944
R4146 vdd.n579 vdd.n576 19.3944
R4147 vdd.n579 vdd.n436 19.3944
R4148 vdd.n585 vdd.n436 19.3944
R4149 vdd.n586 vdd.n585 19.3944
R4150 vdd.n589 vdd.n586 19.3944
R4151 vdd.n589 vdd.n434 19.3944
R4152 vdd.n595 vdd.n434 19.3944
R4153 vdd.n596 vdd.n595 19.3944
R4154 vdd.n599 vdd.n596 19.3944
R4155 vdd.n599 vdd.n432 19.3944
R4156 vdd.n605 vdd.n432 19.3944
R4157 vdd.n606 vdd.n605 19.3944
R4158 vdd.n609 vdd.n606 19.3944
R4159 vdd.n609 vdd.n430 19.3944
R4160 vdd.n615 vdd.n430 19.3944
R4161 vdd.n617 vdd.n615 19.3944
R4162 vdd.n618 vdd.n617 19.3944
R4163 vdd.n516 vdd.n515 19.3944
R4164 vdd.n519 vdd.n516 19.3944
R4165 vdd.n519 vdd.n450 19.3944
R4166 vdd.n525 vdd.n450 19.3944
R4167 vdd.n526 vdd.n525 19.3944
R4168 vdd.n529 vdd.n526 19.3944
R4169 vdd.n529 vdd.n448 19.3944
R4170 vdd.n535 vdd.n448 19.3944
R4171 vdd.n536 vdd.n535 19.3944
R4172 vdd.n539 vdd.n536 19.3944
R4173 vdd.n539 vdd.n446 19.3944
R4174 vdd.n545 vdd.n446 19.3944
R4175 vdd.n546 vdd.n545 19.3944
R4176 vdd.n549 vdd.n546 19.3944
R4177 vdd.n549 vdd.n444 19.3944
R4178 vdd.n555 vdd.n444 19.3944
R4179 vdd.n556 vdd.n555 19.3944
R4180 vdd.n559 vdd.n556 19.3944
R4181 vdd.n559 vdd.n442 19.3944
R4182 vdd.n565 vdd.n442 19.3944
R4183 vdd.n466 vdd.n465 19.3944
R4184 vdd.n469 vdd.n466 19.3944
R4185 vdd.n469 vdd.n462 19.3944
R4186 vdd.n475 vdd.n462 19.3944
R4187 vdd.n476 vdd.n475 19.3944
R4188 vdd.n479 vdd.n476 19.3944
R4189 vdd.n479 vdd.n460 19.3944
R4190 vdd.n485 vdd.n460 19.3944
R4191 vdd.n486 vdd.n485 19.3944
R4192 vdd.n489 vdd.n486 19.3944
R4193 vdd.n489 vdd.n458 19.3944
R4194 vdd.n495 vdd.n458 19.3944
R4195 vdd.n496 vdd.n495 19.3944
R4196 vdd.n499 vdd.n496 19.3944
R4197 vdd.n499 vdd.n456 19.3944
R4198 vdd.n505 vdd.n456 19.3944
R4199 vdd.n506 vdd.n505 19.3944
R4200 vdd.n509 vdd.n506 19.3944
R4201 vdd.n3325 vdd.n683 19.3944
R4202 vdd.n3325 vdd.n681 19.3944
R4203 vdd.n3329 vdd.n681 19.3944
R4204 vdd.n3329 vdd.n671 19.3944
R4205 vdd.n3342 vdd.n671 19.3944
R4206 vdd.n3342 vdd.n669 19.3944
R4207 vdd.n3346 vdd.n669 19.3944
R4208 vdd.n3346 vdd.n660 19.3944
R4209 vdd.n3358 vdd.n660 19.3944
R4210 vdd.n3358 vdd.n658 19.3944
R4211 vdd.n3362 vdd.n658 19.3944
R4212 vdd.n3362 vdd.n648 19.3944
R4213 vdd.n3375 vdd.n648 19.3944
R4214 vdd.n3375 vdd.n646 19.3944
R4215 vdd.n3379 vdd.n646 19.3944
R4216 vdd.n3379 vdd.n637 19.3944
R4217 vdd.n3394 vdd.n637 19.3944
R4218 vdd.n3394 vdd.n635 19.3944
R4219 vdd.n3398 vdd.n635 19.3944
R4220 vdd.n3398 vdd.n336 19.3944
R4221 vdd.n3489 vdd.n336 19.3944
R4222 vdd.n3489 vdd.n337 19.3944
R4223 vdd.n3483 vdd.n337 19.3944
R4224 vdd.n3483 vdd.n3482 19.3944
R4225 vdd.n3482 vdd.n3481 19.3944
R4226 vdd.n3481 vdd.n349 19.3944
R4227 vdd.n3475 vdd.n349 19.3944
R4228 vdd.n3475 vdd.n3474 19.3944
R4229 vdd.n3474 vdd.n3473 19.3944
R4230 vdd.n3473 vdd.n359 19.3944
R4231 vdd.n3467 vdd.n359 19.3944
R4232 vdd.n3467 vdd.n3466 19.3944
R4233 vdd.n3466 vdd.n3465 19.3944
R4234 vdd.n3465 vdd.n370 19.3944
R4235 vdd.n3459 vdd.n370 19.3944
R4236 vdd.n3459 vdd.n3458 19.3944
R4237 vdd.n3458 vdd.n3457 19.3944
R4238 vdd.n3457 vdd.n381 19.3944
R4239 vdd.n3451 vdd.n381 19.3944
R4240 vdd.n3451 vdd.n3450 19.3944
R4241 vdd.n3450 vdd.n3449 19.3944
R4242 vdd.n3272 vdd.n747 19.3944
R4243 vdd.n3272 vdd.n3269 19.3944
R4244 vdd.n3269 vdd.n3266 19.3944
R4245 vdd.n3266 vdd.n3265 19.3944
R4246 vdd.n3265 vdd.n3262 19.3944
R4247 vdd.n3262 vdd.n3261 19.3944
R4248 vdd.n3261 vdd.n3258 19.3944
R4249 vdd.n3258 vdd.n3257 19.3944
R4250 vdd.n3257 vdd.n3254 19.3944
R4251 vdd.n3254 vdd.n3253 19.3944
R4252 vdd.n3253 vdd.n3250 19.3944
R4253 vdd.n3250 vdd.n3249 19.3944
R4254 vdd.n3249 vdd.n3246 19.3944
R4255 vdd.n3246 vdd.n3245 19.3944
R4256 vdd.n3245 vdd.n3242 19.3944
R4257 vdd.n3242 vdd.n3241 19.3944
R4258 vdd.n3241 vdd.n3238 19.3944
R4259 vdd.n3238 vdd.n3237 19.3944
R4260 vdd.n3237 vdd.n3234 19.3944
R4261 vdd.n3234 vdd.n3233 19.3944
R4262 vdd.n3312 vdd.n3311 19.3944
R4263 vdd.n3311 vdd.n3310 19.3944
R4264 vdd.n732 vdd.n729 19.3944
R4265 vdd.n3306 vdd.n3305 19.3944
R4266 vdd.n3305 vdd.n3302 19.3944
R4267 vdd.n3302 vdd.n3301 19.3944
R4268 vdd.n3301 vdd.n3298 19.3944
R4269 vdd.n3298 vdd.n3297 19.3944
R4270 vdd.n3297 vdd.n3294 19.3944
R4271 vdd.n3294 vdd.n3293 19.3944
R4272 vdd.n3293 vdd.n3290 19.3944
R4273 vdd.n3290 vdd.n3289 19.3944
R4274 vdd.n3289 vdd.n3286 19.3944
R4275 vdd.n3286 vdd.n3285 19.3944
R4276 vdd.n3285 vdd.n3282 19.3944
R4277 vdd.n3282 vdd.n3281 19.3944
R4278 vdd.n3226 vdd.n767 19.3944
R4279 vdd.n3226 vdd.n3223 19.3944
R4280 vdd.n3223 vdd.n3220 19.3944
R4281 vdd.n3220 vdd.n3219 19.3944
R4282 vdd.n3219 vdd.n3216 19.3944
R4283 vdd.n3216 vdd.n3215 19.3944
R4284 vdd.n3215 vdd.n3212 19.3944
R4285 vdd.n3212 vdd.n3211 19.3944
R4286 vdd.n3211 vdd.n3208 19.3944
R4287 vdd.n3208 vdd.n3207 19.3944
R4288 vdd.n3207 vdd.n3204 19.3944
R4289 vdd.n3204 vdd.n3203 19.3944
R4290 vdd.n3203 vdd.n3200 19.3944
R4291 vdd.n3200 vdd.n3199 19.3944
R4292 vdd.n3199 vdd.n3196 19.3944
R4293 vdd.n3196 vdd.n3195 19.3944
R4294 vdd.n3192 vdd.n3191 19.3944
R4295 vdd.n3188 vdd.n3187 19.3944
R4296 vdd.n1719 vdd.n1715 19.0066
R4297 vdd.n2307 vdd.n1189 19.0066
R4298 vdd.n569 vdd.n566 19.0066
R4299 vdd.n3230 vdd.n767 19.0066
R4300 vdd.n1254 vdd.n1253 16.0975
R4301 vdd.n982 vdd.n981 16.0975
R4302 vdd.n1680 vdd.n1679 16.0975
R4303 vdd.n1718 vdd.n1717 16.0975
R4304 vdd.n1614 vdd.n1613 16.0975
R4305 vdd.n2270 vdd.n2269 16.0975
R4306 vdd.n1191 vdd.n1190 16.0975
R4307 vdd.n1151 vdd.n1150 16.0975
R4308 vdd.n1274 vdd.n1273 16.0975
R4309 vdd.n973 vdd.n972 16.0975
R4310 vdd.n2705 vdd.n2704 16.0975
R4311 vdd.n427 vdd.n426 16.0975
R4312 vdd.n441 vdd.n440 16.0975
R4313 vdd.n453 vdd.n452 16.0975
R4314 vdd.n769 vdd.n768 16.0975
R4315 vdd.n3277 vdd.n3276 16.0975
R4316 vdd.n833 vdd.n832 16.0975
R4317 vdd.n2702 vdd.n2701 16.0975
R4318 vdd.n689 vdd.n688 16.0975
R4319 vdd.n800 vdd.n799 16.0975
R4320 vdd.t130 vdd.n2665 15.4182
R4321 vdd.n2938 vdd.t22 15.4182
R4322 vdd.n28 vdd.n27 14.5674
R4323 vdd.n2417 vdd.n1076 14.0578
R4324 vdd.n3151 vdd.n692 14.0578
R4325 vdd.n328 vdd.n293 13.1884
R4326 vdd.n269 vdd.n234 13.1884
R4327 vdd.n226 vdd.n191 13.1884
R4328 vdd.n167 vdd.n132 13.1884
R4329 vdd.n125 vdd.n90 13.1884
R4330 vdd.n66 vdd.n31 13.1884
R4331 vdd.n2109 vdd.n2074 13.1884
R4332 vdd.n2168 vdd.n2133 13.1884
R4333 vdd.n2007 vdd.n1972 13.1884
R4334 vdd.n2066 vdd.n2031 13.1884
R4335 vdd.n1906 vdd.n1871 13.1884
R4336 vdd.n1965 vdd.n1930 13.1884
R4337 vdd.n1750 vdd.n1615 12.9944
R4338 vdd.n1754 vdd.n1615 12.9944
R4339 vdd.n2346 vdd.n1149 12.9944
R4340 vdd.n2347 vdd.n2346 12.9944
R4341 vdd.n515 vdd.n454 12.9944
R4342 vdd.n509 vdd.n454 12.9944
R4343 vdd.n3278 vdd.n747 12.9944
R4344 vdd.n3281 vdd.n3278 12.9944
R4345 vdd.n329 vdd.n291 12.8005
R4346 vdd.n324 vdd.n295 12.8005
R4347 vdd.n270 vdd.n232 12.8005
R4348 vdd.n265 vdd.n236 12.8005
R4349 vdd.n227 vdd.n189 12.8005
R4350 vdd.n222 vdd.n193 12.8005
R4351 vdd.n168 vdd.n130 12.8005
R4352 vdd.n163 vdd.n134 12.8005
R4353 vdd.n126 vdd.n88 12.8005
R4354 vdd.n121 vdd.n92 12.8005
R4355 vdd.n67 vdd.n29 12.8005
R4356 vdd.n62 vdd.n33 12.8005
R4357 vdd.n2110 vdd.n2072 12.8005
R4358 vdd.n2105 vdd.n2076 12.8005
R4359 vdd.n2169 vdd.n2131 12.8005
R4360 vdd.n2164 vdd.n2135 12.8005
R4361 vdd.n2008 vdd.n1970 12.8005
R4362 vdd.n2003 vdd.n1974 12.8005
R4363 vdd.n2067 vdd.n2029 12.8005
R4364 vdd.n2062 vdd.n2033 12.8005
R4365 vdd.n1907 vdd.n1869 12.8005
R4366 vdd.n1902 vdd.n1873 12.8005
R4367 vdd.n1966 vdd.n1928 12.8005
R4368 vdd.n1961 vdd.n1932 12.8005
R4369 vdd.n323 vdd.n296 12.0247
R4370 vdd.n264 vdd.n237 12.0247
R4371 vdd.n221 vdd.n194 12.0247
R4372 vdd.n162 vdd.n135 12.0247
R4373 vdd.n120 vdd.n93 12.0247
R4374 vdd.n61 vdd.n34 12.0247
R4375 vdd.n2104 vdd.n2077 12.0247
R4376 vdd.n2163 vdd.n2136 12.0247
R4377 vdd.n2002 vdd.n1975 12.0247
R4378 vdd.n2061 vdd.n2034 12.0247
R4379 vdd.n1901 vdd.n1874 12.0247
R4380 vdd.n1960 vdd.n1933 12.0247
R4381 vdd.n1789 vdd.n1545 11.337
R4382 vdd.n1798 vdd.n1545 11.337
R4383 vdd.n1798 vdd.n1797 11.337
R4384 vdd.n1806 vdd.n1539 11.337
R4385 vdd.n1815 vdd.n1814 11.337
R4386 vdd.n1831 vdd.n1523 11.337
R4387 vdd.n1839 vdd.n1516 11.337
R4388 vdd.n1848 vdd.n1847 11.337
R4389 vdd.n1856 vdd.n1505 11.337
R4390 vdd.n2179 vdd.n1494 11.337
R4391 vdd.n2188 vdd.n1488 11.337
R4392 vdd.n2196 vdd.n1482 11.337
R4393 vdd.n2205 vdd.n2204 11.337
R4394 vdd.n2221 vdd.n1466 11.337
R4395 vdd.n2229 vdd.n1459 11.337
R4396 vdd.n2238 vdd.n2237 11.337
R4397 vdd.n2246 vdd.n1442 11.337
R4398 vdd.n2257 vdd.n1442 11.337
R4399 vdd.n2257 vdd.n2256 11.337
R4400 vdd.n3323 vdd.n678 11.337
R4401 vdd.n3331 vdd.n678 11.337
R4402 vdd.n3331 vdd.n679 11.337
R4403 vdd.n3340 vdd.n3339 11.337
R4404 vdd.n3356 vdd.n662 11.337
R4405 vdd.n3364 vdd.n655 11.337
R4406 vdd.n3373 vdd.n3372 11.337
R4407 vdd.n3381 vdd.n644 11.337
R4408 vdd.n3400 vdd.n633 11.337
R4409 vdd.n3487 vdd.n340 11.337
R4410 vdd.n3485 vdd.n344 11.337
R4411 vdd.n3479 vdd.n3478 11.337
R4412 vdd.n3471 vdd.n361 11.337
R4413 vdd.n3470 vdd.n3469 11.337
R4414 vdd.n3463 vdd.n3462 11.337
R4415 vdd.n3461 vdd.n375 11.337
R4416 vdd.n3455 vdd.n3454 11.337
R4417 vdd.n3454 vdd.n3453 11.337
R4418 vdd.n3453 vdd.n386 11.337
R4419 vdd.n320 vdd.n319 11.249
R4420 vdd.n261 vdd.n260 11.249
R4421 vdd.n218 vdd.n217 11.249
R4422 vdd.n159 vdd.n158 11.249
R4423 vdd.n117 vdd.n116 11.249
R4424 vdd.n58 vdd.n57 11.249
R4425 vdd.n2101 vdd.n2100 11.249
R4426 vdd.n2160 vdd.n2159 11.249
R4427 vdd.n1999 vdd.n1998 11.249
R4428 vdd.n2058 vdd.n2057 11.249
R4429 vdd.n1898 vdd.n1897 11.249
R4430 vdd.n1957 vdd.n1956 11.249
R4431 vdd.n1587 vdd.t91 11.2237
R4432 vdd.n3447 vdd.t77 11.2237
R4433 vdd.t218 vdd.n1460 10.7702
R4434 vdd.n3348 vdd.t138 10.7702
R4435 vdd.n305 vdd.n304 10.7238
R4436 vdd.n246 vdd.n245 10.7238
R4437 vdd.n203 vdd.n202 10.7238
R4438 vdd.n144 vdd.n143 10.7238
R4439 vdd.n102 vdd.n101 10.7238
R4440 vdd.n43 vdd.n42 10.7238
R4441 vdd.n2086 vdd.n2085 10.7238
R4442 vdd.n2145 vdd.n2144 10.7238
R4443 vdd.n1984 vdd.n1983 10.7238
R4444 vdd.n2043 vdd.n2042 10.7238
R4445 vdd.n1883 vdd.n1882 10.7238
R4446 vdd.n1942 vdd.n1941 10.7238
R4447 vdd.n2593 vdd.t49 10.6568
R4448 vdd.t51 vdd.n928 10.6568
R4449 vdd.n2426 vdd.n1074 10.6151
R4450 vdd.n2427 vdd.n2426 10.6151
R4451 vdd.n2428 vdd.n2427 10.6151
R4452 vdd.n2428 vdd.n1063 10.6151
R4453 vdd.n2438 vdd.n1063 10.6151
R4454 vdd.n2439 vdd.n2438 10.6151
R4455 vdd.n2440 vdd.n2439 10.6151
R4456 vdd.n2440 vdd.n1050 10.6151
R4457 vdd.n2450 vdd.n1050 10.6151
R4458 vdd.n2451 vdd.n2450 10.6151
R4459 vdd.n2452 vdd.n2451 10.6151
R4460 vdd.n2452 vdd.n1038 10.6151
R4461 vdd.n2463 vdd.n1038 10.6151
R4462 vdd.n2464 vdd.n2463 10.6151
R4463 vdd.n2465 vdd.n2464 10.6151
R4464 vdd.n2465 vdd.n1026 10.6151
R4465 vdd.n2475 vdd.n1026 10.6151
R4466 vdd.n2476 vdd.n2475 10.6151
R4467 vdd.n2477 vdd.n2476 10.6151
R4468 vdd.n2477 vdd.n1014 10.6151
R4469 vdd.n2487 vdd.n1014 10.6151
R4470 vdd.n2488 vdd.n2487 10.6151
R4471 vdd.n2489 vdd.n2488 10.6151
R4472 vdd.n2489 vdd.n1003 10.6151
R4473 vdd.n2499 vdd.n1003 10.6151
R4474 vdd.n2500 vdd.n2499 10.6151
R4475 vdd.n2501 vdd.n2500 10.6151
R4476 vdd.n2501 vdd.n990 10.6151
R4477 vdd.n2513 vdd.n990 10.6151
R4478 vdd.n2514 vdd.n2513 10.6151
R4479 vdd.n2516 vdd.n2514 10.6151
R4480 vdd.n2516 vdd.n2515 10.6151
R4481 vdd.n2515 vdd.n971 10.6151
R4482 vdd.n2663 vdd.n2662 10.6151
R4483 vdd.n2662 vdd.n2661 10.6151
R4484 vdd.n2661 vdd.n2658 10.6151
R4485 vdd.n2658 vdd.n2657 10.6151
R4486 vdd.n2657 vdd.n2654 10.6151
R4487 vdd.n2654 vdd.n2653 10.6151
R4488 vdd.n2653 vdd.n2650 10.6151
R4489 vdd.n2650 vdd.n2649 10.6151
R4490 vdd.n2649 vdd.n2646 10.6151
R4491 vdd.n2646 vdd.n2645 10.6151
R4492 vdd.n2645 vdd.n2642 10.6151
R4493 vdd.n2642 vdd.n2641 10.6151
R4494 vdd.n2641 vdd.n2638 10.6151
R4495 vdd.n2638 vdd.n2637 10.6151
R4496 vdd.n2637 vdd.n2634 10.6151
R4497 vdd.n2634 vdd.n2633 10.6151
R4498 vdd.n2633 vdd.n2630 10.6151
R4499 vdd.n2630 vdd.n2629 10.6151
R4500 vdd.n2629 vdd.n2626 10.6151
R4501 vdd.n2626 vdd.n2625 10.6151
R4502 vdd.n2625 vdd.n2622 10.6151
R4503 vdd.n2622 vdd.n2621 10.6151
R4504 vdd.n2621 vdd.n2618 10.6151
R4505 vdd.n2618 vdd.n2617 10.6151
R4506 vdd.n2617 vdd.n2614 10.6151
R4507 vdd.n2614 vdd.n2613 10.6151
R4508 vdd.n2613 vdd.n2610 10.6151
R4509 vdd.n2610 vdd.n2609 10.6151
R4510 vdd.n2609 vdd.n2606 10.6151
R4511 vdd.n2606 vdd.n2605 10.6151
R4512 vdd.n2605 vdd.n2602 10.6151
R4513 vdd.n2600 vdd.n2597 10.6151
R4514 vdd.n2597 vdd.n2596 10.6151
R4515 vdd.n1311 vdd.n1310 10.6151
R4516 vdd.n1313 vdd.n1311 10.6151
R4517 vdd.n1314 vdd.n1313 10.6151
R4518 vdd.n1316 vdd.n1314 10.6151
R4519 vdd.n1317 vdd.n1316 10.6151
R4520 vdd.n1319 vdd.n1317 10.6151
R4521 vdd.n1320 vdd.n1319 10.6151
R4522 vdd.n1322 vdd.n1320 10.6151
R4523 vdd.n1323 vdd.n1322 10.6151
R4524 vdd.n1325 vdd.n1323 10.6151
R4525 vdd.n1326 vdd.n1325 10.6151
R4526 vdd.n1328 vdd.n1326 10.6151
R4527 vdd.n1329 vdd.n1328 10.6151
R4528 vdd.n1331 vdd.n1329 10.6151
R4529 vdd.n1332 vdd.n1331 10.6151
R4530 vdd.n1334 vdd.n1332 10.6151
R4531 vdd.n1335 vdd.n1334 10.6151
R4532 vdd.n1357 vdd.n1335 10.6151
R4533 vdd.n1357 vdd.n1356 10.6151
R4534 vdd.n1356 vdd.n1355 10.6151
R4535 vdd.n1355 vdd.n1353 10.6151
R4536 vdd.n1353 vdd.n1352 10.6151
R4537 vdd.n1352 vdd.n1350 10.6151
R4538 vdd.n1350 vdd.n1349 10.6151
R4539 vdd.n1349 vdd.n1347 10.6151
R4540 vdd.n1347 vdd.n1346 10.6151
R4541 vdd.n1346 vdd.n1344 10.6151
R4542 vdd.n1344 vdd.n1343 10.6151
R4543 vdd.n1343 vdd.n1341 10.6151
R4544 vdd.n1341 vdd.n1340 10.6151
R4545 vdd.n1340 vdd.n1337 10.6151
R4546 vdd.n1337 vdd.n1336 10.6151
R4547 vdd.n1336 vdd.n974 10.6151
R4548 vdd.n2414 vdd.n2413 10.6151
R4549 vdd.n2413 vdd.n2412 10.6151
R4550 vdd.n2412 vdd.n2411 10.6151
R4551 vdd.n2411 vdd.n2409 10.6151
R4552 vdd.n2409 vdd.n2406 10.6151
R4553 vdd.n2406 vdd.n2405 10.6151
R4554 vdd.n2405 vdd.n2402 10.6151
R4555 vdd.n2402 vdd.n2401 10.6151
R4556 vdd.n2401 vdd.n2398 10.6151
R4557 vdd.n2398 vdd.n2397 10.6151
R4558 vdd.n2397 vdd.n2394 10.6151
R4559 vdd.n2394 vdd.n2393 10.6151
R4560 vdd.n2393 vdd.n2390 10.6151
R4561 vdd.n2390 vdd.n2389 10.6151
R4562 vdd.n2389 vdd.n2386 10.6151
R4563 vdd.n2386 vdd.n2385 10.6151
R4564 vdd.n2385 vdd.n2382 10.6151
R4565 vdd.n2382 vdd.n1119 10.6151
R4566 vdd.n1277 vdd.n1119 10.6151
R4567 vdd.n1278 vdd.n1277 10.6151
R4568 vdd.n1281 vdd.n1278 10.6151
R4569 vdd.n1282 vdd.n1281 10.6151
R4570 vdd.n1285 vdd.n1282 10.6151
R4571 vdd.n1286 vdd.n1285 10.6151
R4572 vdd.n1289 vdd.n1286 10.6151
R4573 vdd.n1290 vdd.n1289 10.6151
R4574 vdd.n1293 vdd.n1290 10.6151
R4575 vdd.n1294 vdd.n1293 10.6151
R4576 vdd.n1297 vdd.n1294 10.6151
R4577 vdd.n1298 vdd.n1297 10.6151
R4578 vdd.n1301 vdd.n1298 10.6151
R4579 vdd.n1306 vdd.n1303 10.6151
R4580 vdd.n1307 vdd.n1306 10.6151
R4581 vdd.n2866 vdd.n2865 10.6151
R4582 vdd.n2865 vdd.n2864 10.6151
R4583 vdd.n2864 vdd.n2703 10.6151
R4584 vdd.n2808 vdd.n2703 10.6151
R4585 vdd.n2809 vdd.n2808 10.6151
R4586 vdd.n2811 vdd.n2809 10.6151
R4587 vdd.n2812 vdd.n2811 10.6151
R4588 vdd.n2814 vdd.n2812 10.6151
R4589 vdd.n2815 vdd.n2814 10.6151
R4590 vdd.n2845 vdd.n2815 10.6151
R4591 vdd.n2845 vdd.n2844 10.6151
R4592 vdd.n2844 vdd.n2843 10.6151
R4593 vdd.n2843 vdd.n2841 10.6151
R4594 vdd.n2841 vdd.n2840 10.6151
R4595 vdd.n2840 vdd.n2838 10.6151
R4596 vdd.n2838 vdd.n2837 10.6151
R4597 vdd.n2837 vdd.n2835 10.6151
R4598 vdd.n2835 vdd.n2834 10.6151
R4599 vdd.n2834 vdd.n2832 10.6151
R4600 vdd.n2832 vdd.n2831 10.6151
R4601 vdd.n2831 vdd.n2829 10.6151
R4602 vdd.n2829 vdd.n2828 10.6151
R4603 vdd.n2828 vdd.n2826 10.6151
R4604 vdd.n2826 vdd.n2825 10.6151
R4605 vdd.n2825 vdd.n2823 10.6151
R4606 vdd.n2823 vdd.n2822 10.6151
R4607 vdd.n2822 vdd.n2820 10.6151
R4608 vdd.n2820 vdd.n2819 10.6151
R4609 vdd.n2819 vdd.n2817 10.6151
R4610 vdd.n2817 vdd.n2816 10.6151
R4611 vdd.n2816 vdd.n836 10.6151
R4612 vdd.n3084 vdd.n836 10.6151
R4613 vdd.n3085 vdd.n3084 10.6151
R4614 vdd.n2935 vdd.n2934 10.6151
R4615 vdd.n2934 vdd.n2933 10.6151
R4616 vdd.n2933 vdd.n2932 10.6151
R4617 vdd.n2932 vdd.n2930 10.6151
R4618 vdd.n2930 vdd.n2927 10.6151
R4619 vdd.n2927 vdd.n2926 10.6151
R4620 vdd.n2926 vdd.n2923 10.6151
R4621 vdd.n2923 vdd.n2922 10.6151
R4622 vdd.n2922 vdd.n2919 10.6151
R4623 vdd.n2919 vdd.n2918 10.6151
R4624 vdd.n2918 vdd.n2915 10.6151
R4625 vdd.n2915 vdd.n2914 10.6151
R4626 vdd.n2914 vdd.n2911 10.6151
R4627 vdd.n2911 vdd.n2910 10.6151
R4628 vdd.n2910 vdd.n2907 10.6151
R4629 vdd.n2907 vdd.n2906 10.6151
R4630 vdd.n2906 vdd.n2903 10.6151
R4631 vdd.n2903 vdd.n2902 10.6151
R4632 vdd.n2902 vdd.n2899 10.6151
R4633 vdd.n2899 vdd.n2898 10.6151
R4634 vdd.n2898 vdd.n2895 10.6151
R4635 vdd.n2895 vdd.n2894 10.6151
R4636 vdd.n2894 vdd.n2891 10.6151
R4637 vdd.n2891 vdd.n2890 10.6151
R4638 vdd.n2890 vdd.n2887 10.6151
R4639 vdd.n2887 vdd.n2886 10.6151
R4640 vdd.n2886 vdd.n2883 10.6151
R4641 vdd.n2883 vdd.n2882 10.6151
R4642 vdd.n2882 vdd.n2879 10.6151
R4643 vdd.n2879 vdd.n2878 10.6151
R4644 vdd.n2878 vdd.n2875 10.6151
R4645 vdd.n2873 vdd.n2870 10.6151
R4646 vdd.n2870 vdd.n2869 10.6151
R4647 vdd.n2947 vdd.n926 10.6151
R4648 vdd.n2948 vdd.n2947 10.6151
R4649 vdd.n2949 vdd.n2948 10.6151
R4650 vdd.n2949 vdd.n915 10.6151
R4651 vdd.n2959 vdd.n915 10.6151
R4652 vdd.n2960 vdd.n2959 10.6151
R4653 vdd.n2961 vdd.n2960 10.6151
R4654 vdd.n2961 vdd.n903 10.6151
R4655 vdd.n2971 vdd.n903 10.6151
R4656 vdd.n2972 vdd.n2971 10.6151
R4657 vdd.n2973 vdd.n2972 10.6151
R4658 vdd.n2973 vdd.n891 10.6151
R4659 vdd.n2983 vdd.n891 10.6151
R4660 vdd.n2984 vdd.n2983 10.6151
R4661 vdd.n2985 vdd.n2984 10.6151
R4662 vdd.n2985 vdd.n880 10.6151
R4663 vdd.n2995 vdd.n880 10.6151
R4664 vdd.n2996 vdd.n2995 10.6151
R4665 vdd.n2997 vdd.n2996 10.6151
R4666 vdd.n2997 vdd.n866 10.6151
R4667 vdd.n3008 vdd.n866 10.6151
R4668 vdd.n3009 vdd.n3008 10.6151
R4669 vdd.n3010 vdd.n3009 10.6151
R4670 vdd.n3010 vdd.n855 10.6151
R4671 vdd.n3020 vdd.n855 10.6151
R4672 vdd.n3021 vdd.n3020 10.6151
R4673 vdd.n3022 vdd.n3021 10.6151
R4674 vdd.n3022 vdd.n841 10.6151
R4675 vdd.n3077 vdd.n841 10.6151
R4676 vdd.n3078 vdd.n3077 10.6151
R4677 vdd.n3079 vdd.n3078 10.6151
R4678 vdd.n3079 vdd.n810 10.6151
R4679 vdd.n3149 vdd.n810 10.6151
R4680 vdd.n3148 vdd.n3147 10.6151
R4681 vdd.n3147 vdd.n811 10.6151
R4682 vdd.n812 vdd.n811 10.6151
R4683 vdd.n3140 vdd.n812 10.6151
R4684 vdd.n3140 vdd.n3139 10.6151
R4685 vdd.n3139 vdd.n3138 10.6151
R4686 vdd.n3138 vdd.n814 10.6151
R4687 vdd.n3133 vdd.n814 10.6151
R4688 vdd.n3133 vdd.n3132 10.6151
R4689 vdd.n3132 vdd.n3131 10.6151
R4690 vdd.n3131 vdd.n817 10.6151
R4691 vdd.n3126 vdd.n817 10.6151
R4692 vdd.n3126 vdd.n3125 10.6151
R4693 vdd.n3125 vdd.n3124 10.6151
R4694 vdd.n3124 vdd.n820 10.6151
R4695 vdd.n3119 vdd.n820 10.6151
R4696 vdd.n3119 vdd.n731 10.6151
R4697 vdd.n3115 vdd.n731 10.6151
R4698 vdd.n3115 vdd.n3114 10.6151
R4699 vdd.n3114 vdd.n3113 10.6151
R4700 vdd.n3113 vdd.n823 10.6151
R4701 vdd.n3108 vdd.n823 10.6151
R4702 vdd.n3108 vdd.n3107 10.6151
R4703 vdd.n3107 vdd.n3106 10.6151
R4704 vdd.n3106 vdd.n826 10.6151
R4705 vdd.n3101 vdd.n826 10.6151
R4706 vdd.n3101 vdd.n3100 10.6151
R4707 vdd.n3100 vdd.n3099 10.6151
R4708 vdd.n3099 vdd.n829 10.6151
R4709 vdd.n3094 vdd.n829 10.6151
R4710 vdd.n3094 vdd.n3093 10.6151
R4711 vdd.n3091 vdd.n834 10.6151
R4712 vdd.n3086 vdd.n834 10.6151
R4713 vdd.n3067 vdd.n3028 10.6151
R4714 vdd.n3062 vdd.n3028 10.6151
R4715 vdd.n3062 vdd.n3061 10.6151
R4716 vdd.n3061 vdd.n3060 10.6151
R4717 vdd.n3060 vdd.n3030 10.6151
R4718 vdd.n3055 vdd.n3030 10.6151
R4719 vdd.n3055 vdd.n3054 10.6151
R4720 vdd.n3054 vdd.n3053 10.6151
R4721 vdd.n3053 vdd.n3033 10.6151
R4722 vdd.n3048 vdd.n3033 10.6151
R4723 vdd.n3048 vdd.n3047 10.6151
R4724 vdd.n3047 vdd.n3046 10.6151
R4725 vdd.n3046 vdd.n3036 10.6151
R4726 vdd.n3041 vdd.n3036 10.6151
R4727 vdd.n3041 vdd.n3040 10.6151
R4728 vdd.n3040 vdd.n785 10.6151
R4729 vdd.n3184 vdd.n785 10.6151
R4730 vdd.n3184 vdd.n786 10.6151
R4731 vdd.n788 vdd.n786 10.6151
R4732 vdd.n3177 vdd.n788 10.6151
R4733 vdd.n3177 vdd.n3176 10.6151
R4734 vdd.n3176 vdd.n3175 10.6151
R4735 vdd.n3175 vdd.n790 10.6151
R4736 vdd.n3170 vdd.n790 10.6151
R4737 vdd.n3170 vdd.n3169 10.6151
R4738 vdd.n3169 vdd.n3168 10.6151
R4739 vdd.n3168 vdd.n793 10.6151
R4740 vdd.n3163 vdd.n793 10.6151
R4741 vdd.n3163 vdd.n3162 10.6151
R4742 vdd.n3162 vdd.n3161 10.6151
R4743 vdd.n3161 vdd.n796 10.6151
R4744 vdd.n3156 vdd.n3155 10.6151
R4745 vdd.n3155 vdd.n3154 10.6151
R4746 vdd.n2774 vdd.n2773 10.6151
R4747 vdd.n2860 vdd.n2774 10.6151
R4748 vdd.n2860 vdd.n2859 10.6151
R4749 vdd.n2859 vdd.n2858 10.6151
R4750 vdd.n2858 vdd.n2856 10.6151
R4751 vdd.n2856 vdd.n2855 10.6151
R4752 vdd.n2855 vdd.n2853 10.6151
R4753 vdd.n2853 vdd.n2852 10.6151
R4754 vdd.n2852 vdd.n2850 10.6151
R4755 vdd.n2850 vdd.n2849 10.6151
R4756 vdd.n2849 vdd.n2806 10.6151
R4757 vdd.n2806 vdd.n2805 10.6151
R4758 vdd.n2805 vdd.n2803 10.6151
R4759 vdd.n2803 vdd.n2802 10.6151
R4760 vdd.n2802 vdd.n2800 10.6151
R4761 vdd.n2800 vdd.n2799 10.6151
R4762 vdd.n2799 vdd.n2797 10.6151
R4763 vdd.n2797 vdd.n2796 10.6151
R4764 vdd.n2796 vdd.n2794 10.6151
R4765 vdd.n2794 vdd.n2793 10.6151
R4766 vdd.n2793 vdd.n2791 10.6151
R4767 vdd.n2791 vdd.n2790 10.6151
R4768 vdd.n2790 vdd.n2788 10.6151
R4769 vdd.n2788 vdd.n2787 10.6151
R4770 vdd.n2787 vdd.n2785 10.6151
R4771 vdd.n2785 vdd.n2784 10.6151
R4772 vdd.n2784 vdd.n2782 10.6151
R4773 vdd.n2782 vdd.n2781 10.6151
R4774 vdd.n2781 vdd.n2779 10.6151
R4775 vdd.n2779 vdd.n2778 10.6151
R4776 vdd.n2778 vdd.n2776 10.6151
R4777 vdd.n2776 vdd.n2775 10.6151
R4778 vdd.n2775 vdd.n802 10.6151
R4779 vdd.n2941 vdd.n932 10.6151
R4780 vdd.n2708 vdd.n932 10.6151
R4781 vdd.n2709 vdd.n2708 10.6151
R4782 vdd.n2712 vdd.n2709 10.6151
R4783 vdd.n2713 vdd.n2712 10.6151
R4784 vdd.n2716 vdd.n2713 10.6151
R4785 vdd.n2717 vdd.n2716 10.6151
R4786 vdd.n2720 vdd.n2717 10.6151
R4787 vdd.n2721 vdd.n2720 10.6151
R4788 vdd.n2724 vdd.n2721 10.6151
R4789 vdd.n2725 vdd.n2724 10.6151
R4790 vdd.n2728 vdd.n2725 10.6151
R4791 vdd.n2729 vdd.n2728 10.6151
R4792 vdd.n2732 vdd.n2729 10.6151
R4793 vdd.n2733 vdd.n2732 10.6151
R4794 vdd.n2736 vdd.n2733 10.6151
R4795 vdd.n2737 vdd.n2736 10.6151
R4796 vdd.n2740 vdd.n2737 10.6151
R4797 vdd.n2741 vdd.n2740 10.6151
R4798 vdd.n2744 vdd.n2741 10.6151
R4799 vdd.n2745 vdd.n2744 10.6151
R4800 vdd.n2748 vdd.n2745 10.6151
R4801 vdd.n2749 vdd.n2748 10.6151
R4802 vdd.n2752 vdd.n2749 10.6151
R4803 vdd.n2753 vdd.n2752 10.6151
R4804 vdd.n2756 vdd.n2753 10.6151
R4805 vdd.n2757 vdd.n2756 10.6151
R4806 vdd.n2760 vdd.n2757 10.6151
R4807 vdd.n2761 vdd.n2760 10.6151
R4808 vdd.n2764 vdd.n2761 10.6151
R4809 vdd.n2765 vdd.n2764 10.6151
R4810 vdd.n2770 vdd.n2768 10.6151
R4811 vdd.n2771 vdd.n2770 10.6151
R4812 vdd.n2943 vdd.n2942 10.6151
R4813 vdd.n2943 vdd.n921 10.6151
R4814 vdd.n2953 vdd.n921 10.6151
R4815 vdd.n2954 vdd.n2953 10.6151
R4816 vdd.n2955 vdd.n2954 10.6151
R4817 vdd.n2955 vdd.n909 10.6151
R4818 vdd.n2965 vdd.n909 10.6151
R4819 vdd.n2966 vdd.n2965 10.6151
R4820 vdd.n2967 vdd.n2966 10.6151
R4821 vdd.n2967 vdd.n897 10.6151
R4822 vdd.n2977 vdd.n897 10.6151
R4823 vdd.n2978 vdd.n2977 10.6151
R4824 vdd.n2979 vdd.n2978 10.6151
R4825 vdd.n2979 vdd.n886 10.6151
R4826 vdd.n2989 vdd.n886 10.6151
R4827 vdd.n2990 vdd.n2989 10.6151
R4828 vdd.n2991 vdd.n2990 10.6151
R4829 vdd.n2991 vdd.n873 10.6151
R4830 vdd.n3001 vdd.n873 10.6151
R4831 vdd.n3002 vdd.n3001 10.6151
R4832 vdd.n3004 vdd.n861 10.6151
R4833 vdd.n3014 vdd.n861 10.6151
R4834 vdd.n3015 vdd.n3014 10.6151
R4835 vdd.n3016 vdd.n3015 10.6151
R4836 vdd.n3016 vdd.n849 10.6151
R4837 vdd.n3026 vdd.n849 10.6151
R4838 vdd.n3027 vdd.n3026 10.6151
R4839 vdd.n3073 vdd.n3027 10.6151
R4840 vdd.n3073 vdd.n3072 10.6151
R4841 vdd.n3072 vdd.n3071 10.6151
R4842 vdd.n3071 vdd.n3070 10.6151
R4843 vdd.n3070 vdd.n3068 10.6151
R4844 vdd.n2422 vdd.n2421 10.6151
R4845 vdd.n2422 vdd.n1069 10.6151
R4846 vdd.n2432 vdd.n1069 10.6151
R4847 vdd.n2433 vdd.n2432 10.6151
R4848 vdd.n2434 vdd.n2433 10.6151
R4849 vdd.n2434 vdd.n1057 10.6151
R4850 vdd.n2444 vdd.n1057 10.6151
R4851 vdd.n2445 vdd.n2444 10.6151
R4852 vdd.n2446 vdd.n2445 10.6151
R4853 vdd.n2446 vdd.n1044 10.6151
R4854 vdd.n2456 vdd.n1044 10.6151
R4855 vdd.n2457 vdd.n2456 10.6151
R4856 vdd.n2459 vdd.n1032 10.6151
R4857 vdd.n2469 vdd.n1032 10.6151
R4858 vdd.n2470 vdd.n2469 10.6151
R4859 vdd.n2471 vdd.n2470 10.6151
R4860 vdd.n2471 vdd.n1020 10.6151
R4861 vdd.n2481 vdd.n1020 10.6151
R4862 vdd.n2482 vdd.n2481 10.6151
R4863 vdd.n2483 vdd.n2482 10.6151
R4864 vdd.n2483 vdd.n1009 10.6151
R4865 vdd.n2493 vdd.n1009 10.6151
R4866 vdd.n2494 vdd.n2493 10.6151
R4867 vdd.n2495 vdd.n2494 10.6151
R4868 vdd.n2495 vdd.n997 10.6151
R4869 vdd.n2505 vdd.n997 10.6151
R4870 vdd.n2506 vdd.n2505 10.6151
R4871 vdd.n2509 vdd.n2506 10.6151
R4872 vdd.n2509 vdd.n2508 10.6151
R4873 vdd.n2508 vdd.n2507 10.6151
R4874 vdd.n2507 vdd.n980 10.6151
R4875 vdd.n2591 vdd.n980 10.6151
R4876 vdd.n2590 vdd.n2589 10.6151
R4877 vdd.n2589 vdd.n2586 10.6151
R4878 vdd.n2586 vdd.n2585 10.6151
R4879 vdd.n2585 vdd.n2582 10.6151
R4880 vdd.n2582 vdd.n2581 10.6151
R4881 vdd.n2581 vdd.n2578 10.6151
R4882 vdd.n2578 vdd.n2577 10.6151
R4883 vdd.n2577 vdd.n2574 10.6151
R4884 vdd.n2574 vdd.n2573 10.6151
R4885 vdd.n2573 vdd.n2570 10.6151
R4886 vdd.n2570 vdd.n2569 10.6151
R4887 vdd.n2569 vdd.n2566 10.6151
R4888 vdd.n2566 vdd.n2565 10.6151
R4889 vdd.n2565 vdd.n2562 10.6151
R4890 vdd.n2562 vdd.n2561 10.6151
R4891 vdd.n2561 vdd.n2558 10.6151
R4892 vdd.n2558 vdd.n2557 10.6151
R4893 vdd.n2557 vdd.n2554 10.6151
R4894 vdd.n2554 vdd.n2553 10.6151
R4895 vdd.n2553 vdd.n2550 10.6151
R4896 vdd.n2550 vdd.n2549 10.6151
R4897 vdd.n2549 vdd.n2546 10.6151
R4898 vdd.n2546 vdd.n2545 10.6151
R4899 vdd.n2545 vdd.n2542 10.6151
R4900 vdd.n2542 vdd.n2541 10.6151
R4901 vdd.n2541 vdd.n2538 10.6151
R4902 vdd.n2538 vdd.n2537 10.6151
R4903 vdd.n2537 vdd.n2534 10.6151
R4904 vdd.n2534 vdd.n2533 10.6151
R4905 vdd.n2533 vdd.n2530 10.6151
R4906 vdd.n2530 vdd.n2529 10.6151
R4907 vdd.n2526 vdd.n2525 10.6151
R4908 vdd.n2525 vdd.n2523 10.6151
R4909 vdd.n1388 vdd.n1386 10.6151
R4910 vdd.n1386 vdd.n1385 10.6151
R4911 vdd.n1385 vdd.n1383 10.6151
R4912 vdd.n1383 vdd.n1382 10.6151
R4913 vdd.n1382 vdd.n1380 10.6151
R4914 vdd.n1380 vdd.n1379 10.6151
R4915 vdd.n1379 vdd.n1377 10.6151
R4916 vdd.n1377 vdd.n1376 10.6151
R4917 vdd.n1376 vdd.n1374 10.6151
R4918 vdd.n1374 vdd.n1373 10.6151
R4919 vdd.n1373 vdd.n1371 10.6151
R4920 vdd.n1371 vdd.n1370 10.6151
R4921 vdd.n1370 vdd.n1368 10.6151
R4922 vdd.n1368 vdd.n1367 10.6151
R4923 vdd.n1367 vdd.n1365 10.6151
R4924 vdd.n1365 vdd.n1364 10.6151
R4925 vdd.n1364 vdd.n1362 10.6151
R4926 vdd.n1362 vdd.n1361 10.6151
R4927 vdd.n1361 vdd.n1272 10.6151
R4928 vdd.n1272 vdd.n1271 10.6151
R4929 vdd.n1271 vdd.n1269 10.6151
R4930 vdd.n1269 vdd.n1268 10.6151
R4931 vdd.n1268 vdd.n1266 10.6151
R4932 vdd.n1266 vdd.n1265 10.6151
R4933 vdd.n1265 vdd.n1263 10.6151
R4934 vdd.n1263 vdd.n1262 10.6151
R4935 vdd.n1262 vdd.n1260 10.6151
R4936 vdd.n1260 vdd.n1259 10.6151
R4937 vdd.n1259 vdd.n1257 10.6151
R4938 vdd.n1257 vdd.n1256 10.6151
R4939 vdd.n1256 vdd.n984 10.6151
R4940 vdd.n2521 vdd.n984 10.6151
R4941 vdd.n2522 vdd.n2521 10.6151
R4942 vdd.n2420 vdd.n1081 10.6151
R4943 vdd.n1223 vdd.n1081 10.6151
R4944 vdd.n1224 vdd.n1223 10.6151
R4945 vdd.n1227 vdd.n1224 10.6151
R4946 vdd.n1228 vdd.n1227 10.6151
R4947 vdd.n1231 vdd.n1228 10.6151
R4948 vdd.n1232 vdd.n1231 10.6151
R4949 vdd.n1235 vdd.n1232 10.6151
R4950 vdd.n1236 vdd.n1235 10.6151
R4951 vdd.n1239 vdd.n1236 10.6151
R4952 vdd.n1240 vdd.n1239 10.6151
R4953 vdd.n1243 vdd.n1240 10.6151
R4954 vdd.n1244 vdd.n1243 10.6151
R4955 vdd.n1247 vdd.n1244 10.6151
R4956 vdd.n1248 vdd.n1247 10.6151
R4957 vdd.n1251 vdd.n1248 10.6151
R4958 vdd.n1422 vdd.n1251 10.6151
R4959 vdd.n1422 vdd.n1421 10.6151
R4960 vdd.n1421 vdd.n1419 10.6151
R4961 vdd.n1419 vdd.n1416 10.6151
R4962 vdd.n1416 vdd.n1415 10.6151
R4963 vdd.n1415 vdd.n1412 10.6151
R4964 vdd.n1412 vdd.n1411 10.6151
R4965 vdd.n1411 vdd.n1408 10.6151
R4966 vdd.n1408 vdd.n1407 10.6151
R4967 vdd.n1407 vdd.n1404 10.6151
R4968 vdd.n1404 vdd.n1403 10.6151
R4969 vdd.n1403 vdd.n1400 10.6151
R4970 vdd.n1400 vdd.n1399 10.6151
R4971 vdd.n1399 vdd.n1396 10.6151
R4972 vdd.n1396 vdd.n1395 10.6151
R4973 vdd.n1392 vdd.n1391 10.6151
R4974 vdd.n1391 vdd.n1389 10.6151
R4975 vdd.n2213 vdd.t153 10.5435
R4976 vdd.n656 vdd.t150 10.5435
R4977 vdd.n316 vdd.n298 10.4732
R4978 vdd.n257 vdd.n239 10.4732
R4979 vdd.n214 vdd.n196 10.4732
R4980 vdd.n155 vdd.n137 10.4732
R4981 vdd.n113 vdd.n95 10.4732
R4982 vdd.n54 vdd.n36 10.4732
R4983 vdd.n2097 vdd.n2079 10.4732
R4984 vdd.n2156 vdd.n2138 10.4732
R4985 vdd.n1995 vdd.n1977 10.4732
R4986 vdd.n2054 vdd.n2036 10.4732
R4987 vdd.n1894 vdd.n1876 10.4732
R4988 vdd.n1953 vdd.n1935 10.4732
R4989 vdd.t185 vdd.n2187 10.3167
R4990 vdd.n3392 vdd.t173 10.3167
R4991 vdd.n1864 vdd.t136 10.09
R4992 vdd.n3486 vdd.t167 10.09
R4993 vdd.t140 vdd.n1517 9.86327
R4994 vdd.n3477 vdd.t226 9.86327
R4995 vdd.n2382 vdd.n2381 9.78206
R4996 vdd.n3308 vdd.n731 9.78206
R4997 vdd.n3185 vdd.n3184 9.78206
R4998 vdd.n2274 vdd.n1422 9.78206
R4999 vdd.n315 vdd.n300 9.69747
R5000 vdd.n256 vdd.n241 9.69747
R5001 vdd.n213 vdd.n198 9.69747
R5002 vdd.n154 vdd.n139 9.69747
R5003 vdd.n112 vdd.n97 9.69747
R5004 vdd.n53 vdd.n38 9.69747
R5005 vdd.n2096 vdd.n2081 9.69747
R5006 vdd.n2155 vdd.n2140 9.69747
R5007 vdd.n1994 vdd.n1979 9.69747
R5008 vdd.n2053 vdd.n2038 9.69747
R5009 vdd.n1893 vdd.n1878 9.69747
R5010 vdd.n1952 vdd.n1937 9.69747
R5011 vdd.n1823 vdd.t232 9.63654
R5012 vdd.n3423 vdd.t198 9.63654
R5013 vdd.n331 vdd.n330 9.45567
R5014 vdd.n272 vdd.n271 9.45567
R5015 vdd.n229 vdd.n228 9.45567
R5016 vdd.n170 vdd.n169 9.45567
R5017 vdd.n128 vdd.n127 9.45567
R5018 vdd.n69 vdd.n68 9.45567
R5019 vdd.n2112 vdd.n2111 9.45567
R5020 vdd.n2171 vdd.n2170 9.45567
R5021 vdd.n2010 vdd.n2009 9.45567
R5022 vdd.n2069 vdd.n2068 9.45567
R5023 vdd.n1909 vdd.n1908 9.45567
R5024 vdd.n1968 vdd.n1967 9.45567
R5025 vdd.n1797 vdd.t144 9.40981
R5026 vdd.n3455 vdd.t159 9.40981
R5027 vdd.n2344 vdd.n1149 9.3005
R5028 vdd.n2343 vdd.n2342 9.3005
R5029 vdd.n1155 vdd.n1154 9.3005
R5030 vdd.n2337 vdd.n1159 9.3005
R5031 vdd.n2336 vdd.n1160 9.3005
R5032 vdd.n2335 vdd.n1161 9.3005
R5033 vdd.n1165 vdd.n1162 9.3005
R5034 vdd.n2330 vdd.n1166 9.3005
R5035 vdd.n2329 vdd.n1167 9.3005
R5036 vdd.n2328 vdd.n1168 9.3005
R5037 vdd.n1172 vdd.n1169 9.3005
R5038 vdd.n2323 vdd.n1173 9.3005
R5039 vdd.n2322 vdd.n1174 9.3005
R5040 vdd.n2321 vdd.n1175 9.3005
R5041 vdd.n1179 vdd.n1176 9.3005
R5042 vdd.n2316 vdd.n1180 9.3005
R5043 vdd.n2315 vdd.n1181 9.3005
R5044 vdd.n2314 vdd.n1182 9.3005
R5045 vdd.n1186 vdd.n1183 9.3005
R5046 vdd.n2309 vdd.n1187 9.3005
R5047 vdd.n2308 vdd.n1188 9.3005
R5048 vdd.n2307 vdd.n2306 9.3005
R5049 vdd.n2305 vdd.n1189 9.3005
R5050 vdd.n2304 vdd.n2303 9.3005
R5051 vdd.n1195 vdd.n1194 9.3005
R5052 vdd.n2298 vdd.n1199 9.3005
R5053 vdd.n2297 vdd.n1200 9.3005
R5054 vdd.n2296 vdd.n1201 9.3005
R5055 vdd.n1205 vdd.n1202 9.3005
R5056 vdd.n2291 vdd.n1206 9.3005
R5057 vdd.n2290 vdd.n1207 9.3005
R5058 vdd.n2289 vdd.n1208 9.3005
R5059 vdd.n1212 vdd.n1209 9.3005
R5060 vdd.n2284 vdd.n1213 9.3005
R5061 vdd.n2283 vdd.n1214 9.3005
R5062 vdd.n2282 vdd.n1215 9.3005
R5063 vdd.n1219 vdd.n1216 9.3005
R5064 vdd.n2277 vdd.n1220 9.3005
R5065 vdd.n2346 vdd.n2345 9.3005
R5066 vdd.n2368 vdd.n1120 9.3005
R5067 vdd.n2367 vdd.n1128 9.3005
R5068 vdd.n1132 vdd.n1129 9.3005
R5069 vdd.n2362 vdd.n1133 9.3005
R5070 vdd.n2361 vdd.n1134 9.3005
R5071 vdd.n2360 vdd.n1135 9.3005
R5072 vdd.n1139 vdd.n1136 9.3005
R5073 vdd.n2355 vdd.n1140 9.3005
R5074 vdd.n2354 vdd.n1141 9.3005
R5075 vdd.n2353 vdd.n1142 9.3005
R5076 vdd.n1146 vdd.n1143 9.3005
R5077 vdd.n2348 vdd.n1147 9.3005
R5078 vdd.n2347 vdd.n1148 9.3005
R5079 vdd.n2380 vdd.n2379 9.3005
R5080 vdd.n1124 vdd.n1123 9.3005
R5081 vdd.n2177 vdd.n2176 9.3005
R5082 vdd.n1486 vdd.n1485 9.3005
R5083 vdd.n2191 vdd.n2190 9.3005
R5084 vdd.n2192 vdd.n1484 9.3005
R5085 vdd.n2194 vdd.n2193 9.3005
R5086 vdd.n1475 vdd.n1474 9.3005
R5087 vdd.n2208 vdd.n2207 9.3005
R5088 vdd.n2209 vdd.n1473 9.3005
R5089 vdd.n2211 vdd.n2210 9.3005
R5090 vdd.n1464 vdd.n1463 9.3005
R5091 vdd.n2224 vdd.n2223 9.3005
R5092 vdd.n2225 vdd.n1462 9.3005
R5093 vdd.n2227 vdd.n2226 9.3005
R5094 vdd.n1452 vdd.n1451 9.3005
R5095 vdd.n2241 vdd.n2240 9.3005
R5096 vdd.n2242 vdd.n1450 9.3005
R5097 vdd.n2244 vdd.n2243 9.3005
R5098 vdd.n1440 vdd.n1439 9.3005
R5099 vdd.n2260 vdd.n2259 9.3005
R5100 vdd.n2261 vdd.n1438 9.3005
R5101 vdd.n2263 vdd.n2262 9.3005
R5102 vdd.n307 vdd.n306 9.3005
R5103 vdd.n302 vdd.n301 9.3005
R5104 vdd.n313 vdd.n312 9.3005
R5105 vdd.n315 vdd.n314 9.3005
R5106 vdd.n298 vdd.n297 9.3005
R5107 vdd.n321 vdd.n320 9.3005
R5108 vdd.n323 vdd.n322 9.3005
R5109 vdd.n295 vdd.n292 9.3005
R5110 vdd.n330 vdd.n329 9.3005
R5111 vdd.n248 vdd.n247 9.3005
R5112 vdd.n243 vdd.n242 9.3005
R5113 vdd.n254 vdd.n253 9.3005
R5114 vdd.n256 vdd.n255 9.3005
R5115 vdd.n239 vdd.n238 9.3005
R5116 vdd.n262 vdd.n261 9.3005
R5117 vdd.n264 vdd.n263 9.3005
R5118 vdd.n236 vdd.n233 9.3005
R5119 vdd.n271 vdd.n270 9.3005
R5120 vdd.n205 vdd.n204 9.3005
R5121 vdd.n200 vdd.n199 9.3005
R5122 vdd.n211 vdd.n210 9.3005
R5123 vdd.n213 vdd.n212 9.3005
R5124 vdd.n196 vdd.n195 9.3005
R5125 vdd.n219 vdd.n218 9.3005
R5126 vdd.n221 vdd.n220 9.3005
R5127 vdd.n193 vdd.n190 9.3005
R5128 vdd.n228 vdd.n227 9.3005
R5129 vdd.n146 vdd.n145 9.3005
R5130 vdd.n141 vdd.n140 9.3005
R5131 vdd.n152 vdd.n151 9.3005
R5132 vdd.n154 vdd.n153 9.3005
R5133 vdd.n137 vdd.n136 9.3005
R5134 vdd.n160 vdd.n159 9.3005
R5135 vdd.n162 vdd.n161 9.3005
R5136 vdd.n134 vdd.n131 9.3005
R5137 vdd.n169 vdd.n168 9.3005
R5138 vdd.n104 vdd.n103 9.3005
R5139 vdd.n99 vdd.n98 9.3005
R5140 vdd.n110 vdd.n109 9.3005
R5141 vdd.n112 vdd.n111 9.3005
R5142 vdd.n95 vdd.n94 9.3005
R5143 vdd.n118 vdd.n117 9.3005
R5144 vdd.n120 vdd.n119 9.3005
R5145 vdd.n92 vdd.n89 9.3005
R5146 vdd.n127 vdd.n126 9.3005
R5147 vdd.n45 vdd.n44 9.3005
R5148 vdd.n40 vdd.n39 9.3005
R5149 vdd.n51 vdd.n50 9.3005
R5150 vdd.n53 vdd.n52 9.3005
R5151 vdd.n36 vdd.n35 9.3005
R5152 vdd.n59 vdd.n58 9.3005
R5153 vdd.n61 vdd.n60 9.3005
R5154 vdd.n33 vdd.n30 9.3005
R5155 vdd.n68 vdd.n67 9.3005
R5156 vdd.n3230 vdd.n3229 9.3005
R5157 vdd.n3233 vdd.n766 9.3005
R5158 vdd.n3234 vdd.n765 9.3005
R5159 vdd.n3237 vdd.n764 9.3005
R5160 vdd.n3238 vdd.n763 9.3005
R5161 vdd.n3241 vdd.n762 9.3005
R5162 vdd.n3242 vdd.n761 9.3005
R5163 vdd.n3245 vdd.n760 9.3005
R5164 vdd.n3246 vdd.n759 9.3005
R5165 vdd.n3249 vdd.n758 9.3005
R5166 vdd.n3250 vdd.n757 9.3005
R5167 vdd.n3253 vdd.n756 9.3005
R5168 vdd.n3254 vdd.n755 9.3005
R5169 vdd.n3257 vdd.n754 9.3005
R5170 vdd.n3258 vdd.n753 9.3005
R5171 vdd.n3261 vdd.n752 9.3005
R5172 vdd.n3262 vdd.n751 9.3005
R5173 vdd.n3265 vdd.n750 9.3005
R5174 vdd.n3266 vdd.n749 9.3005
R5175 vdd.n3269 vdd.n748 9.3005
R5176 vdd.n3273 vdd.n3272 9.3005
R5177 vdd.n3274 vdd.n747 9.3005
R5178 vdd.n3278 vdd.n3275 9.3005
R5179 vdd.n3281 vdd.n746 9.3005
R5180 vdd.n3282 vdd.n745 9.3005
R5181 vdd.n3285 vdd.n744 9.3005
R5182 vdd.n3286 vdd.n743 9.3005
R5183 vdd.n3289 vdd.n742 9.3005
R5184 vdd.n3290 vdd.n741 9.3005
R5185 vdd.n3293 vdd.n740 9.3005
R5186 vdd.n3294 vdd.n739 9.3005
R5187 vdd.n3297 vdd.n738 9.3005
R5188 vdd.n3298 vdd.n737 9.3005
R5189 vdd.n3301 vdd.n736 9.3005
R5190 vdd.n3302 vdd.n735 9.3005
R5191 vdd.n3305 vdd.n730 9.3005
R5192 vdd.n3311 vdd.n727 9.3005
R5193 vdd.n3312 vdd.n726 9.3005
R5194 vdd.n3326 vdd.n3325 9.3005
R5195 vdd.n3327 vdd.n681 9.3005
R5196 vdd.n3329 vdd.n3328 9.3005
R5197 vdd.n671 vdd.n670 9.3005
R5198 vdd.n3343 vdd.n3342 9.3005
R5199 vdd.n3344 vdd.n669 9.3005
R5200 vdd.n3346 vdd.n3345 9.3005
R5201 vdd.n660 vdd.n659 9.3005
R5202 vdd.n3359 vdd.n3358 9.3005
R5203 vdd.n3360 vdd.n658 9.3005
R5204 vdd.n3362 vdd.n3361 9.3005
R5205 vdd.n648 vdd.n647 9.3005
R5206 vdd.n3376 vdd.n3375 9.3005
R5207 vdd.n3377 vdd.n646 9.3005
R5208 vdd.n3379 vdd.n3378 9.3005
R5209 vdd.n637 vdd.n636 9.3005
R5210 vdd.n3395 vdd.n3394 9.3005
R5211 vdd.n3396 vdd.n635 9.3005
R5212 vdd.n3398 vdd.n3397 9.3005
R5213 vdd.n336 vdd.n334 9.3005
R5214 vdd.n683 vdd.n682 9.3005
R5215 vdd.n3490 vdd.n3489 9.3005
R5216 vdd.n337 vdd.n335 9.3005
R5217 vdd.n3483 vdd.n346 9.3005
R5218 vdd.n3482 vdd.n347 9.3005
R5219 vdd.n3481 vdd.n348 9.3005
R5220 vdd.n355 vdd.n349 9.3005
R5221 vdd.n3475 vdd.n356 9.3005
R5222 vdd.n3474 vdd.n357 9.3005
R5223 vdd.n3473 vdd.n358 9.3005
R5224 vdd.n366 vdd.n359 9.3005
R5225 vdd.n3467 vdd.n367 9.3005
R5226 vdd.n3466 vdd.n368 9.3005
R5227 vdd.n3465 vdd.n369 9.3005
R5228 vdd.n377 vdd.n370 9.3005
R5229 vdd.n3459 vdd.n378 9.3005
R5230 vdd.n3458 vdd.n379 9.3005
R5231 vdd.n3457 vdd.n380 9.3005
R5232 vdd.n388 vdd.n381 9.3005
R5233 vdd.n3451 vdd.n389 9.3005
R5234 vdd.n3450 vdd.n390 9.3005
R5235 vdd.n3449 vdd.n391 9.3005
R5236 vdd.n466 vdd.n463 9.3005
R5237 vdd.n470 vdd.n469 9.3005
R5238 vdd.n471 vdd.n462 9.3005
R5239 vdd.n475 vdd.n472 9.3005
R5240 vdd.n476 vdd.n461 9.3005
R5241 vdd.n480 vdd.n479 9.3005
R5242 vdd.n481 vdd.n460 9.3005
R5243 vdd.n485 vdd.n482 9.3005
R5244 vdd.n486 vdd.n459 9.3005
R5245 vdd.n490 vdd.n489 9.3005
R5246 vdd.n491 vdd.n458 9.3005
R5247 vdd.n495 vdd.n492 9.3005
R5248 vdd.n496 vdd.n457 9.3005
R5249 vdd.n500 vdd.n499 9.3005
R5250 vdd.n501 vdd.n456 9.3005
R5251 vdd.n505 vdd.n502 9.3005
R5252 vdd.n506 vdd.n455 9.3005
R5253 vdd.n510 vdd.n509 9.3005
R5254 vdd.n511 vdd.n454 9.3005
R5255 vdd.n515 vdd.n512 9.3005
R5256 vdd.n516 vdd.n451 9.3005
R5257 vdd.n520 vdd.n519 9.3005
R5258 vdd.n521 vdd.n450 9.3005
R5259 vdd.n525 vdd.n522 9.3005
R5260 vdd.n526 vdd.n449 9.3005
R5261 vdd.n530 vdd.n529 9.3005
R5262 vdd.n531 vdd.n448 9.3005
R5263 vdd.n535 vdd.n532 9.3005
R5264 vdd.n536 vdd.n447 9.3005
R5265 vdd.n540 vdd.n539 9.3005
R5266 vdd.n541 vdd.n446 9.3005
R5267 vdd.n545 vdd.n542 9.3005
R5268 vdd.n546 vdd.n445 9.3005
R5269 vdd.n550 vdd.n549 9.3005
R5270 vdd.n551 vdd.n444 9.3005
R5271 vdd.n555 vdd.n552 9.3005
R5272 vdd.n556 vdd.n443 9.3005
R5273 vdd.n560 vdd.n559 9.3005
R5274 vdd.n561 vdd.n442 9.3005
R5275 vdd.n565 vdd.n562 9.3005
R5276 vdd.n566 vdd.n439 9.3005
R5277 vdd.n570 vdd.n569 9.3005
R5278 vdd.n571 vdd.n438 9.3005
R5279 vdd.n575 vdd.n572 9.3005
R5280 vdd.n576 vdd.n437 9.3005
R5281 vdd.n580 vdd.n579 9.3005
R5282 vdd.n581 vdd.n436 9.3005
R5283 vdd.n585 vdd.n582 9.3005
R5284 vdd.n586 vdd.n435 9.3005
R5285 vdd.n590 vdd.n589 9.3005
R5286 vdd.n591 vdd.n434 9.3005
R5287 vdd.n595 vdd.n592 9.3005
R5288 vdd.n596 vdd.n433 9.3005
R5289 vdd.n600 vdd.n599 9.3005
R5290 vdd.n601 vdd.n432 9.3005
R5291 vdd.n605 vdd.n602 9.3005
R5292 vdd.n606 vdd.n431 9.3005
R5293 vdd.n610 vdd.n609 9.3005
R5294 vdd.n611 vdd.n430 9.3005
R5295 vdd.n615 vdd.n612 9.3005
R5296 vdd.n617 vdd.n429 9.3005
R5297 vdd.n619 vdd.n618 9.3005
R5298 vdd.n3443 vdd.n3442 9.3005
R5299 vdd.n465 vdd.n464 9.3005
R5300 vdd.n3321 vdd.n3320 9.3005
R5301 vdd.n676 vdd.n675 9.3005
R5302 vdd.n3334 vdd.n3333 9.3005
R5303 vdd.n3335 vdd.n674 9.3005
R5304 vdd.n3337 vdd.n3336 9.3005
R5305 vdd.n666 vdd.n665 9.3005
R5306 vdd.n3351 vdd.n3350 9.3005
R5307 vdd.n3352 vdd.n664 9.3005
R5308 vdd.n3354 vdd.n3353 9.3005
R5309 vdd.n653 vdd.n652 9.3005
R5310 vdd.n3367 vdd.n3366 9.3005
R5311 vdd.n3368 vdd.n651 9.3005
R5312 vdd.n3370 vdd.n3369 9.3005
R5313 vdd.n642 vdd.n641 9.3005
R5314 vdd.n3384 vdd.n3383 9.3005
R5315 vdd.n3385 vdd.n640 9.3005
R5316 vdd.n3390 vdd.n3386 9.3005
R5317 vdd.n3389 vdd.n3388 9.3005
R5318 vdd.n3387 vdd.n631 9.3005
R5319 vdd.n3403 vdd.n630 9.3005
R5320 vdd.n3405 vdd.n3404 9.3005
R5321 vdd.n3406 vdd.n629 9.3005
R5322 vdd.n3408 vdd.n3407 9.3005
R5323 vdd.n3410 vdd.n628 9.3005
R5324 vdd.n3412 vdd.n3411 9.3005
R5325 vdd.n3413 vdd.n627 9.3005
R5326 vdd.n3415 vdd.n3414 9.3005
R5327 vdd.n3417 vdd.n626 9.3005
R5328 vdd.n3419 vdd.n3418 9.3005
R5329 vdd.n3420 vdd.n625 9.3005
R5330 vdd.n3422 vdd.n3421 9.3005
R5331 vdd.n3425 vdd.n624 9.3005
R5332 vdd.n3427 vdd.n3426 9.3005
R5333 vdd.n3428 vdd.n623 9.3005
R5334 vdd.n3430 vdd.n3429 9.3005
R5335 vdd.n3432 vdd.n622 9.3005
R5336 vdd.n3434 vdd.n3433 9.3005
R5337 vdd.n3435 vdd.n621 9.3005
R5338 vdd.n3437 vdd.n3436 9.3005
R5339 vdd.n3439 vdd.n620 9.3005
R5340 vdd.n3441 vdd.n3440 9.3005
R5341 vdd.n3319 vdd.n686 9.3005
R5342 vdd.n3318 vdd.n3317 9.3005
R5343 vdd.n3187 vdd.n687 9.3005
R5344 vdd.n3196 vdd.n783 9.3005
R5345 vdd.n3199 vdd.n782 9.3005
R5346 vdd.n3200 vdd.n781 9.3005
R5347 vdd.n3203 vdd.n780 9.3005
R5348 vdd.n3204 vdd.n779 9.3005
R5349 vdd.n3207 vdd.n778 9.3005
R5350 vdd.n3208 vdd.n777 9.3005
R5351 vdd.n3211 vdd.n776 9.3005
R5352 vdd.n3212 vdd.n775 9.3005
R5353 vdd.n3215 vdd.n774 9.3005
R5354 vdd.n3216 vdd.n773 9.3005
R5355 vdd.n3219 vdd.n772 9.3005
R5356 vdd.n3220 vdd.n771 9.3005
R5357 vdd.n3223 vdd.n770 9.3005
R5358 vdd.n3227 vdd.n3226 9.3005
R5359 vdd.n3228 vdd.n767 9.3005
R5360 vdd.n2273 vdd.n2272 9.3005
R5361 vdd.n2268 vdd.n1424 9.3005
R5362 vdd.n1792 vdd.n1791 9.3005
R5363 vdd.n1793 vdd.n1547 9.3005
R5364 vdd.n1795 vdd.n1794 9.3005
R5365 vdd.n1537 vdd.n1536 9.3005
R5366 vdd.n1809 vdd.n1808 9.3005
R5367 vdd.n1810 vdd.n1535 9.3005
R5368 vdd.n1812 vdd.n1811 9.3005
R5369 vdd.n1527 vdd.n1526 9.3005
R5370 vdd.n1826 vdd.n1825 9.3005
R5371 vdd.n1827 vdd.n1525 9.3005
R5372 vdd.n1829 vdd.n1828 9.3005
R5373 vdd.n1514 vdd.n1513 9.3005
R5374 vdd.n1842 vdd.n1841 9.3005
R5375 vdd.n1843 vdd.n1512 9.3005
R5376 vdd.n1845 vdd.n1844 9.3005
R5377 vdd.n1503 vdd.n1502 9.3005
R5378 vdd.n1859 vdd.n1858 9.3005
R5379 vdd.n1860 vdd.n1501 9.3005
R5380 vdd.n1862 vdd.n1861 9.3005
R5381 vdd.n1492 vdd.n1491 9.3005
R5382 vdd.n2182 vdd.n2181 9.3005
R5383 vdd.n2183 vdd.n1490 9.3005
R5384 vdd.n2185 vdd.n2184 9.3005
R5385 vdd.n1480 vdd.n1479 9.3005
R5386 vdd.n2199 vdd.n2198 9.3005
R5387 vdd.n2200 vdd.n1478 9.3005
R5388 vdd.n2202 vdd.n2201 9.3005
R5389 vdd.n1470 vdd.n1469 9.3005
R5390 vdd.n2216 vdd.n2215 9.3005
R5391 vdd.n2217 vdd.n1468 9.3005
R5392 vdd.n2219 vdd.n2218 9.3005
R5393 vdd.n1457 vdd.n1456 9.3005
R5394 vdd.n2232 vdd.n2231 9.3005
R5395 vdd.n2233 vdd.n1455 9.3005
R5396 vdd.n2235 vdd.n2234 9.3005
R5397 vdd.n1447 vdd.n1446 9.3005
R5398 vdd.n2249 vdd.n2248 9.3005
R5399 vdd.n2250 vdd.n1444 9.3005
R5400 vdd.n2254 vdd.n2253 9.3005
R5401 vdd.n2252 vdd.n1445 9.3005
R5402 vdd.n2251 vdd.n1435 9.3005
R5403 vdd.n1549 vdd.n1548 9.3005
R5404 vdd.n1685 vdd.n1684 9.3005
R5405 vdd.n1686 vdd.n1675 9.3005
R5406 vdd.n1688 vdd.n1687 9.3005
R5407 vdd.n1689 vdd.n1674 9.3005
R5408 vdd.n1691 vdd.n1690 9.3005
R5409 vdd.n1692 vdd.n1669 9.3005
R5410 vdd.n1694 vdd.n1693 9.3005
R5411 vdd.n1695 vdd.n1668 9.3005
R5412 vdd.n1697 vdd.n1696 9.3005
R5413 vdd.n1698 vdd.n1663 9.3005
R5414 vdd.n1700 vdd.n1699 9.3005
R5415 vdd.n1701 vdd.n1662 9.3005
R5416 vdd.n1703 vdd.n1702 9.3005
R5417 vdd.n1704 vdd.n1657 9.3005
R5418 vdd.n1706 vdd.n1705 9.3005
R5419 vdd.n1707 vdd.n1656 9.3005
R5420 vdd.n1709 vdd.n1708 9.3005
R5421 vdd.n1710 vdd.n1651 9.3005
R5422 vdd.n1712 vdd.n1711 9.3005
R5423 vdd.n1713 vdd.n1650 9.3005
R5424 vdd.n1715 vdd.n1714 9.3005
R5425 vdd.n1719 vdd.n1646 9.3005
R5426 vdd.n1721 vdd.n1720 9.3005
R5427 vdd.n1722 vdd.n1645 9.3005
R5428 vdd.n1724 vdd.n1723 9.3005
R5429 vdd.n1725 vdd.n1640 9.3005
R5430 vdd.n1727 vdd.n1726 9.3005
R5431 vdd.n1728 vdd.n1639 9.3005
R5432 vdd.n1730 vdd.n1729 9.3005
R5433 vdd.n1731 vdd.n1634 9.3005
R5434 vdd.n1733 vdd.n1732 9.3005
R5435 vdd.n1734 vdd.n1633 9.3005
R5436 vdd.n1736 vdd.n1735 9.3005
R5437 vdd.n1737 vdd.n1628 9.3005
R5438 vdd.n1739 vdd.n1738 9.3005
R5439 vdd.n1740 vdd.n1627 9.3005
R5440 vdd.n1742 vdd.n1741 9.3005
R5441 vdd.n1743 vdd.n1622 9.3005
R5442 vdd.n1745 vdd.n1744 9.3005
R5443 vdd.n1746 vdd.n1621 9.3005
R5444 vdd.n1748 vdd.n1747 9.3005
R5445 vdd.n1749 vdd.n1616 9.3005
R5446 vdd.n1751 vdd.n1750 9.3005
R5447 vdd.n1752 vdd.n1615 9.3005
R5448 vdd.n1754 vdd.n1753 9.3005
R5449 vdd.n1755 vdd.n1608 9.3005
R5450 vdd.n1757 vdd.n1756 9.3005
R5451 vdd.n1758 vdd.n1607 9.3005
R5452 vdd.n1760 vdd.n1759 9.3005
R5453 vdd.n1761 vdd.n1602 9.3005
R5454 vdd.n1763 vdd.n1762 9.3005
R5455 vdd.n1764 vdd.n1601 9.3005
R5456 vdd.n1766 vdd.n1765 9.3005
R5457 vdd.n1767 vdd.n1596 9.3005
R5458 vdd.n1769 vdd.n1768 9.3005
R5459 vdd.n1770 vdd.n1595 9.3005
R5460 vdd.n1772 vdd.n1771 9.3005
R5461 vdd.n1773 vdd.n1590 9.3005
R5462 vdd.n1775 vdd.n1774 9.3005
R5463 vdd.n1776 vdd.n1589 9.3005
R5464 vdd.n1778 vdd.n1777 9.3005
R5465 vdd.n1554 vdd.n1553 9.3005
R5466 vdd.n1784 vdd.n1783 9.3005
R5467 vdd.n1683 vdd.n1682 9.3005
R5468 vdd.n1787 vdd.n1786 9.3005
R5469 vdd.n1543 vdd.n1542 9.3005
R5470 vdd.n1801 vdd.n1800 9.3005
R5471 vdd.n1802 vdd.n1541 9.3005
R5472 vdd.n1804 vdd.n1803 9.3005
R5473 vdd.n1532 vdd.n1531 9.3005
R5474 vdd.n1818 vdd.n1817 9.3005
R5475 vdd.n1819 vdd.n1530 9.3005
R5476 vdd.n1821 vdd.n1820 9.3005
R5477 vdd.n1521 vdd.n1520 9.3005
R5478 vdd.n1834 vdd.n1833 9.3005
R5479 vdd.n1835 vdd.n1519 9.3005
R5480 vdd.n1837 vdd.n1836 9.3005
R5481 vdd.n1509 vdd.n1508 9.3005
R5482 vdd.n1851 vdd.n1850 9.3005
R5483 vdd.n1852 vdd.n1507 9.3005
R5484 vdd.n1854 vdd.n1853 9.3005
R5485 vdd.n1498 vdd.n1497 9.3005
R5486 vdd.n1867 vdd.n1866 9.3005
R5487 vdd.n1868 vdd.n1496 9.3005
R5488 vdd.n1785 vdd.n1552 9.3005
R5489 vdd.n2088 vdd.n2087 9.3005
R5490 vdd.n2083 vdd.n2082 9.3005
R5491 vdd.n2094 vdd.n2093 9.3005
R5492 vdd.n2096 vdd.n2095 9.3005
R5493 vdd.n2079 vdd.n2078 9.3005
R5494 vdd.n2102 vdd.n2101 9.3005
R5495 vdd.n2104 vdd.n2103 9.3005
R5496 vdd.n2076 vdd.n2073 9.3005
R5497 vdd.n2111 vdd.n2110 9.3005
R5498 vdd.n2147 vdd.n2146 9.3005
R5499 vdd.n2142 vdd.n2141 9.3005
R5500 vdd.n2153 vdd.n2152 9.3005
R5501 vdd.n2155 vdd.n2154 9.3005
R5502 vdd.n2138 vdd.n2137 9.3005
R5503 vdd.n2161 vdd.n2160 9.3005
R5504 vdd.n2163 vdd.n2162 9.3005
R5505 vdd.n2135 vdd.n2132 9.3005
R5506 vdd.n2170 vdd.n2169 9.3005
R5507 vdd.n1986 vdd.n1985 9.3005
R5508 vdd.n1981 vdd.n1980 9.3005
R5509 vdd.n1992 vdd.n1991 9.3005
R5510 vdd.n1994 vdd.n1993 9.3005
R5511 vdd.n1977 vdd.n1976 9.3005
R5512 vdd.n2000 vdd.n1999 9.3005
R5513 vdd.n2002 vdd.n2001 9.3005
R5514 vdd.n1974 vdd.n1971 9.3005
R5515 vdd.n2009 vdd.n2008 9.3005
R5516 vdd.n2045 vdd.n2044 9.3005
R5517 vdd.n2040 vdd.n2039 9.3005
R5518 vdd.n2051 vdd.n2050 9.3005
R5519 vdd.n2053 vdd.n2052 9.3005
R5520 vdd.n2036 vdd.n2035 9.3005
R5521 vdd.n2059 vdd.n2058 9.3005
R5522 vdd.n2061 vdd.n2060 9.3005
R5523 vdd.n2033 vdd.n2030 9.3005
R5524 vdd.n2068 vdd.n2067 9.3005
R5525 vdd.n1885 vdd.n1884 9.3005
R5526 vdd.n1880 vdd.n1879 9.3005
R5527 vdd.n1891 vdd.n1890 9.3005
R5528 vdd.n1893 vdd.n1892 9.3005
R5529 vdd.n1876 vdd.n1875 9.3005
R5530 vdd.n1899 vdd.n1898 9.3005
R5531 vdd.n1901 vdd.n1900 9.3005
R5532 vdd.n1873 vdd.n1870 9.3005
R5533 vdd.n1908 vdd.n1907 9.3005
R5534 vdd.n1944 vdd.n1943 9.3005
R5535 vdd.n1939 vdd.n1938 9.3005
R5536 vdd.n1950 vdd.n1949 9.3005
R5537 vdd.n1952 vdd.n1951 9.3005
R5538 vdd.n1935 vdd.n1934 9.3005
R5539 vdd.n1958 vdd.n1957 9.3005
R5540 vdd.n1960 vdd.n1959 9.3005
R5541 vdd.n1932 vdd.n1929 9.3005
R5542 vdd.n1967 vdd.n1966 9.3005
R5543 vdd.n1823 vdd.t208 9.18308
R5544 vdd.n3423 vdd.t142 9.18308
R5545 vdd.n1517 vdd.t183 8.95635
R5546 vdd.n2265 vdd.t67 8.95635
R5547 vdd.n723 vdd.t63 8.95635
R5548 vdd.t155 vdd.n3477 8.95635
R5549 vdd.n312 vdd.n311 8.92171
R5550 vdd.n253 vdd.n252 8.92171
R5551 vdd.n210 vdd.n209 8.92171
R5552 vdd.n151 vdd.n150 8.92171
R5553 vdd.n109 vdd.n108 8.92171
R5554 vdd.n50 vdd.n49 8.92171
R5555 vdd.n2093 vdd.n2092 8.92171
R5556 vdd.n2152 vdd.n2151 8.92171
R5557 vdd.n1991 vdd.n1990 8.92171
R5558 vdd.n2050 vdd.n2049 8.92171
R5559 vdd.n1890 vdd.n1889 8.92171
R5560 vdd.n1949 vdd.n1948 8.92171
R5561 vdd.n231 vdd.n129 8.81535
R5562 vdd.n2071 vdd.n1969 8.81535
R5563 vdd.n1864 vdd.t234 8.72962
R5564 vdd.t157 vdd.n3486 8.72962
R5565 vdd.n2187 vdd.t164 8.50289
R5566 vdd.n3392 vdd.t161 8.50289
R5567 vdd.n28 vdd.n14 8.42249
R5568 vdd.n2213 vdd.t237 8.27616
R5569 vdd.t202 vdd.n656 8.27616
R5570 vdd.n3492 vdd.n3491 8.16225
R5571 vdd.n2175 vdd.n2174 8.16225
R5572 vdd.n308 vdd.n302 8.14595
R5573 vdd.n249 vdd.n243 8.14595
R5574 vdd.n206 vdd.n200 8.14595
R5575 vdd.n147 vdd.n141 8.14595
R5576 vdd.n105 vdd.n99 8.14595
R5577 vdd.n46 vdd.n40 8.14595
R5578 vdd.n2089 vdd.n2083 8.14595
R5579 vdd.n2148 vdd.n2142 8.14595
R5580 vdd.n1987 vdd.n1981 8.14595
R5581 vdd.n2046 vdd.n2040 8.14595
R5582 vdd.n1886 vdd.n1880 8.14595
R5583 vdd.n1945 vdd.n1939 8.14595
R5584 vdd.n1460 vdd.t146 8.04943
R5585 vdd.n3348 vdd.t256 8.04943
R5586 vdd.n2424 vdd.n1076 7.70933
R5587 vdd.n2424 vdd.n1079 7.70933
R5588 vdd.n2430 vdd.n1065 7.70933
R5589 vdd.n2436 vdd.n1065 7.70933
R5590 vdd.n2436 vdd.n1059 7.70933
R5591 vdd.n2442 vdd.n1059 7.70933
R5592 vdd.n2448 vdd.n1052 7.70933
R5593 vdd.n2448 vdd.n1055 7.70933
R5594 vdd.n2454 vdd.n1048 7.70933
R5595 vdd.n2461 vdd.n1034 7.70933
R5596 vdd.n2467 vdd.n1034 7.70933
R5597 vdd.n2473 vdd.n1028 7.70933
R5598 vdd.n2479 vdd.n1024 7.70933
R5599 vdd.n2485 vdd.n1018 7.70933
R5600 vdd.n2497 vdd.n1005 7.70933
R5601 vdd.n2503 vdd.n999 7.70933
R5602 vdd.n2503 vdd.n992 7.70933
R5603 vdd.n2511 vdd.n992 7.70933
R5604 vdd.n2593 vdd.n976 7.70933
R5605 vdd.n2945 vdd.n928 7.70933
R5606 vdd.n2957 vdd.n917 7.70933
R5607 vdd.n2957 vdd.n911 7.70933
R5608 vdd.n2963 vdd.n911 7.70933
R5609 vdd.n2969 vdd.n905 7.70933
R5610 vdd.n2975 vdd.n901 7.70933
R5611 vdd.n2981 vdd.n895 7.70933
R5612 vdd.n2993 vdd.n882 7.70933
R5613 vdd.n2999 vdd.n875 7.70933
R5614 vdd.n2999 vdd.n878 7.70933
R5615 vdd.n3006 vdd.n870 7.70933
R5616 vdd.n3012 vdd.n857 7.70933
R5617 vdd.n3018 vdd.n857 7.70933
R5618 vdd.n3024 vdd.n851 7.70933
R5619 vdd.n3024 vdd.n843 7.70933
R5620 vdd.n3075 vdd.n843 7.70933
R5621 vdd.n3075 vdd.n846 7.70933
R5622 vdd.n3081 vdd.n805 7.70933
R5623 vdd.n3151 vdd.n805 7.70933
R5624 vdd.n3004 vdd.n3003 7.49318
R5625 vdd.n2458 vdd.n2457 7.49318
R5626 vdd.n307 vdd.n304 7.3702
R5627 vdd.n248 vdd.n245 7.3702
R5628 vdd.n205 vdd.n202 7.3702
R5629 vdd.n146 vdd.n143 7.3702
R5630 vdd.n104 vdd.n101 7.3702
R5631 vdd.n45 vdd.n42 7.3702
R5632 vdd.n2088 vdd.n2085 7.3702
R5633 vdd.n2147 vdd.n2144 7.3702
R5634 vdd.n1986 vdd.n1983 7.3702
R5635 vdd.n2045 vdd.n2042 7.3702
R5636 vdd.n1885 vdd.n1882 7.3702
R5637 vdd.n1944 vdd.n1941 7.3702
R5638 vdd.n2442 vdd.t21 7.36923
R5639 vdd.t4 vdd.n851 7.36923
R5640 vdd.n2518 vdd.t298 7.25587
R5641 vdd.n2862 vdd.t16 7.25587
R5642 vdd.n2246 vdd.t190 7.1425
R5643 vdd.n679 vdd.t188 7.1425
R5644 vdd.n1720 vdd.n1719 6.98232
R5645 vdd.n2308 vdd.n2307 6.98232
R5646 vdd.n566 vdd.n565 6.98232
R5647 vdd.n3233 vdd.n3230 6.98232
R5648 vdd.t250 vdd.n1459 6.91577
R5649 vdd.n3356 vdd.t200 6.91577
R5650 vdd.n2205 vdd.t206 6.68904
R5651 vdd.n3372 vdd.t175 6.68904
R5652 vdd.t171 vdd.n1488 6.46231
R5653 vdd.n3400 vdd.t194 6.46231
R5654 vdd.n3492 vdd.n333 6.38151
R5655 vdd.n2174 vdd.n2173 6.38151
R5656 vdd.n1856 vdd.t181 6.23558
R5657 vdd.t247 vdd.n344 6.23558
R5658 vdd.t148 vdd.n1516 6.00885
R5659 vdd.n3471 vdd.t211 6.00885
R5660 vdd.t47 vdd.n1005 5.89549
R5661 vdd.n2969 vdd.t26 5.89549
R5662 vdd.n308 vdd.n307 5.81868
R5663 vdd.n249 vdd.n248 5.81868
R5664 vdd.n206 vdd.n205 5.81868
R5665 vdd.n147 vdd.n146 5.81868
R5666 vdd.n105 vdd.n104 5.81868
R5667 vdd.n46 vdd.n45 5.81868
R5668 vdd.n2089 vdd.n2088 5.81868
R5669 vdd.n2148 vdd.n2147 5.81868
R5670 vdd.n1987 vdd.n1986 5.81868
R5671 vdd.n2046 vdd.n2045 5.81868
R5672 vdd.n1886 vdd.n1885 5.81868
R5673 vdd.n1945 vdd.n1944 5.81868
R5674 vdd.n1815 vdd.t134 5.78212
R5675 vdd.n3462 vdd.t253 5.78212
R5676 vdd.n2601 vdd.n2600 5.77611
R5677 vdd.n1303 vdd.n1302 5.77611
R5678 vdd.n2874 vdd.n2873 5.77611
R5679 vdd.n3092 vdd.n3091 5.77611
R5680 vdd.n3156 vdd.n801 5.77611
R5681 vdd.n2768 vdd.n2706 5.77611
R5682 vdd.n2526 vdd.n983 5.77611
R5683 vdd.n1392 vdd.n1255 5.77611
R5684 vdd.n1682 vdd.n1681 5.62474
R5685 vdd.n2271 vdd.n2268 5.62474
R5686 vdd.n3443 vdd.n428 5.62474
R5687 vdd.n3317 vdd.n690 5.62474
R5688 vdd.n1539 vdd.t134 5.55539
R5689 vdd.t18 vdd.n1028 5.55539
R5690 vdd.n2473 vdd.t9 5.55539
R5691 vdd.t36 vdd.n882 5.55539
R5692 vdd.n2993 vdd.t30 5.55539
R5693 vdd.t253 vdd.n3461 5.55539
R5694 vdd.n1048 vdd.t112 5.44203
R5695 vdd.n3006 vdd.t81 5.44203
R5696 vdd.n1831 vdd.t148 5.32866
R5697 vdd.n2430 vdd.t59 5.32866
R5698 vdd.n1338 vdd.t101 5.32866
R5699 vdd.n2951 vdd.t105 5.32866
R5700 vdd.n846 vdd.t55 5.32866
R5701 vdd.t211 vdd.n3470 5.32866
R5702 vdd.n1847 vdd.t181 5.10193
R5703 vdd.n3479 vdd.t247 5.10193
R5704 vdd.n311 vdd.n302 5.04292
R5705 vdd.n252 vdd.n243 5.04292
R5706 vdd.n209 vdd.n200 5.04292
R5707 vdd.n150 vdd.n141 5.04292
R5708 vdd.n108 vdd.n99 5.04292
R5709 vdd.n49 vdd.n40 5.04292
R5710 vdd.n2092 vdd.n2083 5.04292
R5711 vdd.n2151 vdd.n2142 5.04292
R5712 vdd.n1990 vdd.n1981 5.04292
R5713 vdd.n2049 vdd.n2040 5.04292
R5714 vdd.n1889 vdd.n1880 5.04292
R5715 vdd.n1948 vdd.n1939 5.04292
R5716 vdd.n2479 vdd.t5 4.98857
R5717 vdd.n895 vdd.t24 4.98857
R5718 vdd.n2179 vdd.t171 4.8752
R5719 vdd.t11 vdd.t12 4.8752
R5720 vdd.t10 vdd.t0 4.8752
R5721 vdd.t37 vdd.t53 4.8752
R5722 vdd.t14 vdd.t35 4.8752
R5723 vdd.t194 vdd.n340 4.8752
R5724 vdd.n2602 vdd.n2601 4.83952
R5725 vdd.n1302 vdd.n1301 4.83952
R5726 vdd.n2875 vdd.n2874 4.83952
R5727 vdd.n3093 vdd.n3092 4.83952
R5728 vdd.n801 vdd.n796 4.83952
R5729 vdd.n2765 vdd.n2706 4.83952
R5730 vdd.n2529 vdd.n983 4.83952
R5731 vdd.n1395 vdd.n1255 4.83952
R5732 vdd.n2276 vdd.n2275 4.74817
R5733 vdd.n1428 vdd.n1423 4.74817
R5734 vdd.n1125 vdd.n1122 4.74817
R5735 vdd.n2369 vdd.n1121 4.74817
R5736 vdd.n2374 vdd.n1122 4.74817
R5737 vdd.n2373 vdd.n1121 4.74817
R5738 vdd.n3310 vdd.n3309 4.74817
R5739 vdd.n3307 vdd.n3306 4.74817
R5740 vdd.n3307 vdd.n732 4.74817
R5741 vdd.n3309 vdd.n729 4.74817
R5742 vdd.n3192 vdd.n784 4.74817
R5743 vdd.n3188 vdd.n3186 4.74817
R5744 vdd.n3191 vdd.n3186 4.74817
R5745 vdd.n3195 vdd.n784 4.74817
R5746 vdd.n2275 vdd.n1221 4.74817
R5747 vdd.n1425 vdd.n1423 4.74817
R5748 vdd.n333 vdd.n332 4.7074
R5749 vdd.n231 vdd.n230 4.7074
R5750 vdd.n2173 vdd.n2172 4.7074
R5751 vdd.n2071 vdd.n2070 4.7074
R5752 vdd.n1482 vdd.t206 4.64847
R5753 vdd.n2454 vdd.t8 4.64847
R5754 vdd.n1018 vdd.t3 4.64847
R5755 vdd.n2975 vdd.t2 4.64847
R5756 vdd.n870 vdd.t20 4.64847
R5757 vdd.n3381 vdd.t175 4.64847
R5758 vdd.n2221 vdd.t250 4.42174
R5759 vdd.t200 vdd.n655 4.42174
R5760 vdd.n312 vdd.n300 4.26717
R5761 vdd.n253 vdd.n241 4.26717
R5762 vdd.n210 vdd.n198 4.26717
R5763 vdd.n151 vdd.n139 4.26717
R5764 vdd.n109 vdd.n97 4.26717
R5765 vdd.n50 vdd.n38 4.26717
R5766 vdd.n2093 vdd.n2081 4.26717
R5767 vdd.n2152 vdd.n2140 4.26717
R5768 vdd.n1991 vdd.n1979 4.26717
R5769 vdd.n2050 vdd.n2038 4.26717
R5770 vdd.n1890 vdd.n1878 4.26717
R5771 vdd.n1949 vdd.n1937 4.26717
R5772 vdd.n2237 vdd.t190 4.19501
R5773 vdd.n3340 vdd.t188 4.19501
R5774 vdd.n333 vdd.n231 4.10845
R5775 vdd.n2173 vdd.n2071 4.10845
R5776 vdd.n289 vdd.t222 4.06363
R5777 vdd.n289 vdd.t268 4.06363
R5778 vdd.n287 vdd.t270 4.06363
R5779 vdd.n287 vdd.t143 4.06363
R5780 vdd.n285 vdd.t180 4.06363
R5781 vdd.n285 vdd.t241 4.06363
R5782 vdd.n283 vdd.t274 4.06363
R5783 vdd.n283 vdd.t284 4.06363
R5784 vdd.n281 vdd.t289 4.06363
R5785 vdd.n281 vdd.t187 4.06363
R5786 vdd.n279 vdd.t216 4.06363
R5787 vdd.n279 vdd.t288 4.06363
R5788 vdd.n277 vdd.t290 4.06363
R5789 vdd.n277 vdd.t215 4.06363
R5790 vdd.n275 vdd.t221 4.06363
R5791 vdd.n275 vdd.t224 4.06363
R5792 vdd.n273 vdd.t269 4.06363
R5793 vdd.n273 vdd.t166 4.06363
R5794 vdd.n187 vdd.t199 4.06363
R5795 vdd.n187 vdd.t254 4.06363
R5796 vdd.n185 vdd.t255 4.06363
R5797 vdd.n185 vdd.t286 4.06363
R5798 vdd.n183 vdd.t156 4.06363
R5799 vdd.n183 vdd.t227 4.06363
R5800 vdd.n181 vdd.t260 4.06363
R5801 vdd.n181 vdd.t275 4.06363
R5802 vdd.n179 vdd.t278 4.06363
R5803 vdd.n179 vdd.t158 4.06363
R5804 vdd.n177 vdd.t193 4.06363
R5805 vdd.n177 vdd.t263 4.06363
R5806 vdd.n175 vdd.t279 4.06363
R5807 vdd.n175 vdd.t176 4.06363
R5808 vdd.n173 vdd.t201 4.06363
R5809 vdd.n173 vdd.t203 4.06363
R5810 vdd.n171 vdd.t257 4.06363
R5811 vdd.n171 vdd.t139 4.06363
R5812 vdd.n86 vdd.t231 4.06363
R5813 vdd.n86 vdd.t258 4.06363
R5814 vdd.n84 vdd.t212 4.06363
R5815 vdd.n84 vdd.t280 4.06363
R5816 vdd.n82 vdd.t179 4.06363
R5817 vdd.n82 vdd.t262 4.06363
R5818 vdd.n80 vdd.t168 4.06363
R5819 vdd.n80 vdd.t248 4.06363
R5820 vdd.n78 vdd.t195 4.06363
R5821 vdd.n78 vdd.t276 4.06363
R5822 vdd.n76 vdd.t162 4.06363
R5823 vdd.n76 vdd.t174 4.06363
R5824 vdd.n74 vdd.t151 4.06363
R5825 vdd.n74 vdd.t204 4.06363
R5826 vdd.n72 vdd.t285 4.06363
R5827 vdd.n72 vdd.t267 4.06363
R5828 vdd.n70 vdd.t272 4.06363
R5829 vdd.n70 vdd.t217 4.06363
R5830 vdd.n2113 vdd.t236 4.06363
R5831 vdd.n2113 vdd.t177 4.06363
R5832 vdd.n2115 vdd.t293 4.06363
R5833 vdd.n2115 vdd.t265 4.06363
R5834 vdd.n2117 vdd.t261 4.06363
R5835 vdd.n2117 vdd.t214 4.06363
R5836 vdd.n2119 vdd.t210 4.06363
R5837 vdd.n2119 vdd.t264 4.06363
R5838 vdd.n2121 vdd.t244 4.06363
R5839 vdd.n2121 vdd.t243 4.06363
R5840 vdd.n2123 vdd.t205 4.06363
R5841 vdd.n2123 vdd.t178 4.06363
R5842 vdd.n2125 vdd.t169 4.06363
R5843 vdd.n2125 vdd.t242 4.06363
R5844 vdd.n2127 vdd.t225 4.06363
R5845 vdd.n2127 vdd.t170 4.06363
R5846 vdd.n2129 vdd.t163 4.06363
R5847 vdd.n2129 vdd.t266 4.06363
R5848 vdd.n2011 vdd.t223 4.06363
R5849 vdd.n2011 vdd.t147 4.06363
R5850 vdd.n2013 vdd.t283 4.06363
R5851 vdd.n2013 vdd.t251 4.06363
R5852 vdd.n2015 vdd.t245 4.06363
R5853 vdd.n2015 vdd.t192 4.06363
R5854 vdd.n2017 vdd.t186 4.06363
R5855 vdd.n2017 vdd.t246 4.06363
R5856 vdd.n2019 vdd.t235 4.06363
R5857 vdd.n2019 vdd.t172 4.06363
R5858 vdd.n2021 vdd.t182 4.06363
R5859 vdd.n2021 vdd.t152 4.06363
R5860 vdd.n2023 vdd.t141 4.06363
R5861 vdd.n2023 vdd.t230 4.06363
R5862 vdd.n2025 vdd.t209 4.06363
R5863 vdd.n2025 vdd.t149 4.06363
R5864 vdd.n2027 vdd.t135 4.06363
R5865 vdd.n2027 vdd.t252 4.06363
R5866 vdd.n1910 vdd.t219 4.06363
R5867 vdd.n1910 vdd.t273 4.06363
R5868 vdd.n1912 vdd.t238 4.06363
R5869 vdd.n1912 vdd.t287 4.06363
R5870 vdd.n1914 vdd.t207 4.06363
R5871 vdd.n1914 vdd.t154 4.06363
R5872 vdd.n1916 vdd.t229 4.06363
R5873 vdd.n1916 vdd.t165 4.06363
R5874 vdd.n1918 vdd.t277 4.06363
R5875 vdd.n1918 vdd.t292 4.06363
R5876 vdd.n1920 vdd.t249 4.06363
R5877 vdd.n1920 vdd.t137 4.06363
R5878 vdd.n1922 vdd.t239 4.06363
R5879 vdd.n1922 vdd.t184 4.06363
R5880 vdd.n1924 vdd.t281 4.06363
R5881 vdd.n1924 vdd.t213 4.06363
R5882 vdd.n1926 vdd.t259 4.06363
R5883 vdd.n1926 vdd.t233 4.06363
R5884 vdd.n26 vdd.t45 3.9605
R5885 vdd.n26 vdd.t33 3.9605
R5886 vdd.n23 vdd.t42 3.9605
R5887 vdd.n23 vdd.t43 3.9605
R5888 vdd.n21 vdd.t32 3.9605
R5889 vdd.n21 vdd.t29 3.9605
R5890 vdd.n20 vdd.t44 3.9605
R5891 vdd.n20 vdd.t41 3.9605
R5892 vdd.n15 vdd.t297 3.9605
R5893 vdd.n15 vdd.t46 3.9605
R5894 vdd.n16 vdd.t39 3.9605
R5895 vdd.n16 vdd.t40 3.9605
R5896 vdd.n18 vdd.t34 3.9605
R5897 vdd.n18 vdd.t19 3.9605
R5898 vdd.n25 vdd.t296 3.9605
R5899 vdd.n25 vdd.t28 3.9605
R5900 vdd.n2511 vdd.t132 3.85492
R5901 vdd.n1338 vdd.t132 3.85492
R5902 vdd.n2951 vdd.t294 3.85492
R5903 vdd.t294 vdd.n917 3.85492
R5904 vdd.n7 vdd.t15 3.61217
R5905 vdd.n7 vdd.t25 3.61217
R5906 vdd.n8 vdd.t38 3.61217
R5907 vdd.n8 vdd.t27 3.61217
R5908 vdd.n10 vdd.t17 3.61217
R5909 vdd.n10 vdd.t295 3.61217
R5910 vdd.n12 vdd.t23 3.61217
R5911 vdd.n12 vdd.t52 3.61217
R5912 vdd.n5 vdd.t50 3.61217
R5913 vdd.n5 vdd.t131 3.61217
R5914 vdd.n3 vdd.t133 3.61217
R5915 vdd.n3 vdd.t299 3.61217
R5916 vdd.n1 vdd.t48 3.61217
R5917 vdd.n1 vdd.t1 3.61217
R5918 vdd.n0 vdd.t6 3.61217
R5919 vdd.n0 vdd.t13 3.61217
R5920 vdd.n316 vdd.n315 3.49141
R5921 vdd.n257 vdd.n256 3.49141
R5922 vdd.n214 vdd.n213 3.49141
R5923 vdd.n155 vdd.n154 3.49141
R5924 vdd.n113 vdd.n112 3.49141
R5925 vdd.n54 vdd.n53 3.49141
R5926 vdd.n2097 vdd.n2096 3.49141
R5927 vdd.n2156 vdd.n2155 3.49141
R5928 vdd.n1995 vdd.n1994 3.49141
R5929 vdd.n2054 vdd.n2053 3.49141
R5930 vdd.n1894 vdd.n1893 3.49141
R5931 vdd.n1953 vdd.n1952 3.49141
R5932 vdd.n2665 vdd.t49 3.40145
R5933 vdd.n2938 vdd.t51 3.40145
R5934 vdd.n2238 vdd.t146 3.28809
R5935 vdd.n3339 vdd.t256 3.28809
R5936 vdd.n3003 vdd.n3002 3.12245
R5937 vdd.n2459 vdd.n2458 3.12245
R5938 vdd.t237 vdd.n1466 3.06136
R5939 vdd.n1055 vdd.t8 3.06136
R5940 vdd.n2491 vdd.t3 3.06136
R5941 vdd.n2847 vdd.t2 3.06136
R5942 vdd.n3012 vdd.t20 3.06136
R5943 vdd.n3364 vdd.t202 3.06136
R5944 vdd.n2196 vdd.t164 2.83463
R5945 vdd.n644 vdd.t161 2.83463
R5946 vdd.n1359 vdd.t5 2.72126
R5947 vdd.n2987 vdd.t24 2.72126
R5948 vdd.n319 vdd.n298 2.71565
R5949 vdd.n260 vdd.n239 2.71565
R5950 vdd.n217 vdd.n196 2.71565
R5951 vdd.n158 vdd.n137 2.71565
R5952 vdd.n116 vdd.n95 2.71565
R5953 vdd.n57 vdd.n36 2.71565
R5954 vdd.n2100 vdd.n2079 2.71565
R5955 vdd.n2159 vdd.n2138 2.71565
R5956 vdd.n1998 vdd.n1977 2.71565
R5957 vdd.n2057 vdd.n2036 2.71565
R5958 vdd.n1897 vdd.n1876 2.71565
R5959 vdd.n1956 vdd.n1935 2.71565
R5960 vdd.t234 vdd.n1494 2.6079
R5961 vdd.n3487 vdd.t157 2.6079
R5962 vdd.t0 vdd.n999 2.49453
R5963 vdd.n2963 vdd.t37 2.49453
R5964 vdd.n306 vdd.n305 2.4129
R5965 vdd.n247 vdd.n246 2.4129
R5966 vdd.n204 vdd.n203 2.4129
R5967 vdd.n145 vdd.n144 2.4129
R5968 vdd.n103 vdd.n102 2.4129
R5969 vdd.n44 vdd.n43 2.4129
R5970 vdd.n2087 vdd.n2086 2.4129
R5971 vdd.n2146 vdd.n2145 2.4129
R5972 vdd.n1985 vdd.n1984 2.4129
R5973 vdd.n2044 vdd.n2043 2.4129
R5974 vdd.n1884 vdd.n1883 2.4129
R5975 vdd.n1943 vdd.n1942 2.4129
R5976 vdd.n1848 vdd.t183 2.38117
R5977 vdd.n2256 vdd.t67 2.38117
R5978 vdd.n1079 vdd.t59 2.38117
R5979 vdd.n2518 vdd.t101 2.38117
R5980 vdd.n2862 vdd.t105 2.38117
R5981 vdd.n3081 vdd.t55 2.38117
R5982 vdd.n3323 vdd.t63 2.38117
R5983 vdd.n3478 vdd.t155 2.38117
R5984 vdd.n2381 vdd.n1122 2.27742
R5985 vdd.n2381 vdd.n1121 2.27742
R5986 vdd.n3308 vdd.n3307 2.27742
R5987 vdd.n3309 vdd.n3308 2.27742
R5988 vdd.n3186 vdd.n3185 2.27742
R5989 vdd.n3185 vdd.n784 2.27742
R5990 vdd.n2275 vdd.n2274 2.27742
R5991 vdd.n2274 vdd.n1423 2.27742
R5992 vdd.t208 vdd.n1523 2.15444
R5993 vdd.n2467 vdd.t18 2.15444
R5994 vdd.n1359 vdd.t9 2.15444
R5995 vdd.n2987 vdd.t36 2.15444
R5996 vdd.t30 vdd.n875 2.15444
R5997 vdd.n3469 vdd.t142 2.15444
R5998 vdd.n320 vdd.n296 1.93989
R5999 vdd.n261 vdd.n237 1.93989
R6000 vdd.n218 vdd.n194 1.93989
R6001 vdd.n159 vdd.n135 1.93989
R6002 vdd.n117 vdd.n93 1.93989
R6003 vdd.n58 vdd.n34 1.93989
R6004 vdd.n2101 vdd.n2077 1.93989
R6005 vdd.n2160 vdd.n2136 1.93989
R6006 vdd.n1999 vdd.n1975 1.93989
R6007 vdd.n2058 vdd.n2034 1.93989
R6008 vdd.n1898 vdd.n1874 1.93989
R6009 vdd.n1957 vdd.n1933 1.93989
R6010 vdd.n1806 vdd.t144 1.92771
R6011 vdd.t159 vdd.n375 1.92771
R6012 vdd.n2491 vdd.t47 1.81434
R6013 vdd.n2847 vdd.t26 1.81434
R6014 vdd.n1814 vdd.t232 1.70098
R6015 vdd.n3463 vdd.t198 1.70098
R6016 vdd.n2485 vdd.t12 1.58761
R6017 vdd.n901 vdd.t14 1.58761
R6018 vdd.n1839 vdd.t140 1.47425
R6019 vdd.n361 vdd.t226 1.47425
R6020 vdd.n1505 vdd.t136 1.24752
R6021 vdd.n2461 vdd.t31 1.24752
R6022 vdd.n1024 vdd.t11 1.24752
R6023 vdd.n2981 vdd.t35 1.24752
R6024 vdd.n878 vdd.t7 1.24752
R6025 vdd.t167 vdd.n3485 1.24752
R6026 vdd.n331 vdd.n291 1.16414
R6027 vdd.n324 vdd.n323 1.16414
R6028 vdd.n272 vdd.n232 1.16414
R6029 vdd.n265 vdd.n264 1.16414
R6030 vdd.n229 vdd.n189 1.16414
R6031 vdd.n222 vdd.n221 1.16414
R6032 vdd.n170 vdd.n130 1.16414
R6033 vdd.n163 vdd.n162 1.16414
R6034 vdd.n128 vdd.n88 1.16414
R6035 vdd.n121 vdd.n120 1.16414
R6036 vdd.n69 vdd.n29 1.16414
R6037 vdd.n62 vdd.n61 1.16414
R6038 vdd.n2112 vdd.n2072 1.16414
R6039 vdd.n2105 vdd.n2104 1.16414
R6040 vdd.n2171 vdd.n2131 1.16414
R6041 vdd.n2164 vdd.n2163 1.16414
R6042 vdd.n2010 vdd.n1970 1.16414
R6043 vdd.n2003 vdd.n2002 1.16414
R6044 vdd.n2069 vdd.n2029 1.16414
R6045 vdd.n2062 vdd.n2061 1.16414
R6046 vdd.n1909 vdd.n1869 1.16414
R6047 vdd.n1902 vdd.n1901 1.16414
R6048 vdd.n1968 vdd.n1928 1.16414
R6049 vdd.n1961 vdd.n1960 1.16414
R6050 vdd.n2188 vdd.t185 1.02079
R6051 vdd.t112 vdd.t31 1.02079
R6052 vdd.t7 vdd.t81 1.02079
R6053 vdd.t173 vdd.n633 1.02079
R6054 vdd.n2174 vdd.n28 1.00834
R6055 vdd vdd.n3492 1.0005
R6056 vdd.n1685 vdd.n1681 0.970197
R6057 vdd.n2272 vdd.n2271 0.970197
R6058 vdd.n618 vdd.n428 0.970197
R6059 vdd.n3187 vdd.n690 0.970197
R6060 vdd.n2204 vdd.t153 0.794056
R6061 vdd.n3373 vdd.t150 0.794056
R6062 vdd.n2229 vdd.t218 0.567326
R6063 vdd.t138 vdd.n662 0.567326
R6064 vdd.n2262 vdd.n1123 0.530988
R6065 vdd.n726 vdd.n682 0.530988
R6066 vdd.n464 vdd.n391 0.530988
R6067 vdd.n3442 vdd.n3441 0.530988
R6068 vdd.n3319 vdd.n3318 0.530988
R6069 vdd.n2251 vdd.n1424 0.530988
R6070 vdd.n1683 vdd.n1548 0.530988
R6071 vdd.n1785 vdd.n1784 0.530988
R6072 vdd.n4 vdd.n2 0.459552
R6073 vdd.n11 vdd.n9 0.459552
R6074 vdd.t298 vdd.n976 0.453961
R6075 vdd.n2945 vdd.t16 0.453961
R6076 vdd.n329 vdd.n328 0.388379
R6077 vdd.n295 vdd.n293 0.388379
R6078 vdd.n270 vdd.n269 0.388379
R6079 vdd.n236 vdd.n234 0.388379
R6080 vdd.n227 vdd.n226 0.388379
R6081 vdd.n193 vdd.n191 0.388379
R6082 vdd.n168 vdd.n167 0.388379
R6083 vdd.n134 vdd.n132 0.388379
R6084 vdd.n126 vdd.n125 0.388379
R6085 vdd.n92 vdd.n90 0.388379
R6086 vdd.n67 vdd.n66 0.388379
R6087 vdd.n33 vdd.n31 0.388379
R6088 vdd.n2110 vdd.n2109 0.388379
R6089 vdd.n2076 vdd.n2074 0.388379
R6090 vdd.n2169 vdd.n2168 0.388379
R6091 vdd.n2135 vdd.n2133 0.388379
R6092 vdd.n2008 vdd.n2007 0.388379
R6093 vdd.n1974 vdd.n1972 0.388379
R6094 vdd.n2067 vdd.n2066 0.388379
R6095 vdd.n2033 vdd.n2031 0.388379
R6096 vdd.n1907 vdd.n1906 0.388379
R6097 vdd.n1873 vdd.n1871 0.388379
R6098 vdd.n1966 vdd.n1965 0.388379
R6099 vdd.n1932 vdd.n1930 0.388379
R6100 vdd.n19 vdd.n17 0.387128
R6101 vdd.n24 vdd.n22 0.387128
R6102 vdd.n6 vdd.n4 0.358259
R6103 vdd.n13 vdd.n11 0.358259
R6104 vdd.n276 vdd.n274 0.358259
R6105 vdd.n278 vdd.n276 0.358259
R6106 vdd.n280 vdd.n278 0.358259
R6107 vdd.n282 vdd.n280 0.358259
R6108 vdd.n284 vdd.n282 0.358259
R6109 vdd.n286 vdd.n284 0.358259
R6110 vdd.n288 vdd.n286 0.358259
R6111 vdd.n290 vdd.n288 0.358259
R6112 vdd.n332 vdd.n290 0.358259
R6113 vdd.n174 vdd.n172 0.358259
R6114 vdd.n176 vdd.n174 0.358259
R6115 vdd.n178 vdd.n176 0.358259
R6116 vdd.n180 vdd.n178 0.358259
R6117 vdd.n182 vdd.n180 0.358259
R6118 vdd.n184 vdd.n182 0.358259
R6119 vdd.n186 vdd.n184 0.358259
R6120 vdd.n188 vdd.n186 0.358259
R6121 vdd.n230 vdd.n188 0.358259
R6122 vdd.n73 vdd.n71 0.358259
R6123 vdd.n75 vdd.n73 0.358259
R6124 vdd.n77 vdd.n75 0.358259
R6125 vdd.n79 vdd.n77 0.358259
R6126 vdd.n81 vdd.n79 0.358259
R6127 vdd.n83 vdd.n81 0.358259
R6128 vdd.n85 vdd.n83 0.358259
R6129 vdd.n87 vdd.n85 0.358259
R6130 vdd.n129 vdd.n87 0.358259
R6131 vdd.n2172 vdd.n2130 0.358259
R6132 vdd.n2130 vdd.n2128 0.358259
R6133 vdd.n2128 vdd.n2126 0.358259
R6134 vdd.n2126 vdd.n2124 0.358259
R6135 vdd.n2124 vdd.n2122 0.358259
R6136 vdd.n2122 vdd.n2120 0.358259
R6137 vdd.n2120 vdd.n2118 0.358259
R6138 vdd.n2118 vdd.n2116 0.358259
R6139 vdd.n2116 vdd.n2114 0.358259
R6140 vdd.n2070 vdd.n2028 0.358259
R6141 vdd.n2028 vdd.n2026 0.358259
R6142 vdd.n2026 vdd.n2024 0.358259
R6143 vdd.n2024 vdd.n2022 0.358259
R6144 vdd.n2022 vdd.n2020 0.358259
R6145 vdd.n2020 vdd.n2018 0.358259
R6146 vdd.n2018 vdd.n2016 0.358259
R6147 vdd.n2016 vdd.n2014 0.358259
R6148 vdd.n2014 vdd.n2012 0.358259
R6149 vdd.n1969 vdd.n1927 0.358259
R6150 vdd.n1927 vdd.n1925 0.358259
R6151 vdd.n1925 vdd.n1923 0.358259
R6152 vdd.n1923 vdd.n1921 0.358259
R6153 vdd.n1921 vdd.n1919 0.358259
R6154 vdd.n1919 vdd.n1917 0.358259
R6155 vdd.n1917 vdd.n1915 0.358259
R6156 vdd.n1915 vdd.n1913 0.358259
R6157 vdd.n1913 vdd.n1911 0.358259
R6158 vdd.t21 vdd.n1052 0.340595
R6159 vdd.n2497 vdd.t10 0.340595
R6160 vdd.t53 vdd.n905 0.340595
R6161 vdd.n3018 vdd.t4 0.340595
R6162 vdd.n14 vdd.n6 0.334552
R6163 vdd.n14 vdd.n13 0.334552
R6164 vdd.n27 vdd.n19 0.21707
R6165 vdd.n27 vdd.n24 0.21707
R6166 vdd.n330 vdd.n292 0.155672
R6167 vdd.n322 vdd.n292 0.155672
R6168 vdd.n322 vdd.n321 0.155672
R6169 vdd.n321 vdd.n297 0.155672
R6170 vdd.n314 vdd.n297 0.155672
R6171 vdd.n314 vdd.n313 0.155672
R6172 vdd.n313 vdd.n301 0.155672
R6173 vdd.n306 vdd.n301 0.155672
R6174 vdd.n271 vdd.n233 0.155672
R6175 vdd.n263 vdd.n233 0.155672
R6176 vdd.n263 vdd.n262 0.155672
R6177 vdd.n262 vdd.n238 0.155672
R6178 vdd.n255 vdd.n238 0.155672
R6179 vdd.n255 vdd.n254 0.155672
R6180 vdd.n254 vdd.n242 0.155672
R6181 vdd.n247 vdd.n242 0.155672
R6182 vdd.n228 vdd.n190 0.155672
R6183 vdd.n220 vdd.n190 0.155672
R6184 vdd.n220 vdd.n219 0.155672
R6185 vdd.n219 vdd.n195 0.155672
R6186 vdd.n212 vdd.n195 0.155672
R6187 vdd.n212 vdd.n211 0.155672
R6188 vdd.n211 vdd.n199 0.155672
R6189 vdd.n204 vdd.n199 0.155672
R6190 vdd.n169 vdd.n131 0.155672
R6191 vdd.n161 vdd.n131 0.155672
R6192 vdd.n161 vdd.n160 0.155672
R6193 vdd.n160 vdd.n136 0.155672
R6194 vdd.n153 vdd.n136 0.155672
R6195 vdd.n153 vdd.n152 0.155672
R6196 vdd.n152 vdd.n140 0.155672
R6197 vdd.n145 vdd.n140 0.155672
R6198 vdd.n127 vdd.n89 0.155672
R6199 vdd.n119 vdd.n89 0.155672
R6200 vdd.n119 vdd.n118 0.155672
R6201 vdd.n118 vdd.n94 0.155672
R6202 vdd.n111 vdd.n94 0.155672
R6203 vdd.n111 vdd.n110 0.155672
R6204 vdd.n110 vdd.n98 0.155672
R6205 vdd.n103 vdd.n98 0.155672
R6206 vdd.n68 vdd.n30 0.155672
R6207 vdd.n60 vdd.n30 0.155672
R6208 vdd.n60 vdd.n59 0.155672
R6209 vdd.n59 vdd.n35 0.155672
R6210 vdd.n52 vdd.n35 0.155672
R6211 vdd.n52 vdd.n51 0.155672
R6212 vdd.n51 vdd.n39 0.155672
R6213 vdd.n44 vdd.n39 0.155672
R6214 vdd.n2111 vdd.n2073 0.155672
R6215 vdd.n2103 vdd.n2073 0.155672
R6216 vdd.n2103 vdd.n2102 0.155672
R6217 vdd.n2102 vdd.n2078 0.155672
R6218 vdd.n2095 vdd.n2078 0.155672
R6219 vdd.n2095 vdd.n2094 0.155672
R6220 vdd.n2094 vdd.n2082 0.155672
R6221 vdd.n2087 vdd.n2082 0.155672
R6222 vdd.n2170 vdd.n2132 0.155672
R6223 vdd.n2162 vdd.n2132 0.155672
R6224 vdd.n2162 vdd.n2161 0.155672
R6225 vdd.n2161 vdd.n2137 0.155672
R6226 vdd.n2154 vdd.n2137 0.155672
R6227 vdd.n2154 vdd.n2153 0.155672
R6228 vdd.n2153 vdd.n2141 0.155672
R6229 vdd.n2146 vdd.n2141 0.155672
R6230 vdd.n2009 vdd.n1971 0.155672
R6231 vdd.n2001 vdd.n1971 0.155672
R6232 vdd.n2001 vdd.n2000 0.155672
R6233 vdd.n2000 vdd.n1976 0.155672
R6234 vdd.n1993 vdd.n1976 0.155672
R6235 vdd.n1993 vdd.n1992 0.155672
R6236 vdd.n1992 vdd.n1980 0.155672
R6237 vdd.n1985 vdd.n1980 0.155672
R6238 vdd.n2068 vdd.n2030 0.155672
R6239 vdd.n2060 vdd.n2030 0.155672
R6240 vdd.n2060 vdd.n2059 0.155672
R6241 vdd.n2059 vdd.n2035 0.155672
R6242 vdd.n2052 vdd.n2035 0.155672
R6243 vdd.n2052 vdd.n2051 0.155672
R6244 vdd.n2051 vdd.n2039 0.155672
R6245 vdd.n2044 vdd.n2039 0.155672
R6246 vdd.n1908 vdd.n1870 0.155672
R6247 vdd.n1900 vdd.n1870 0.155672
R6248 vdd.n1900 vdd.n1899 0.155672
R6249 vdd.n1899 vdd.n1875 0.155672
R6250 vdd.n1892 vdd.n1875 0.155672
R6251 vdd.n1892 vdd.n1891 0.155672
R6252 vdd.n1891 vdd.n1879 0.155672
R6253 vdd.n1884 vdd.n1879 0.155672
R6254 vdd.n1967 vdd.n1929 0.155672
R6255 vdd.n1959 vdd.n1929 0.155672
R6256 vdd.n1959 vdd.n1958 0.155672
R6257 vdd.n1958 vdd.n1934 0.155672
R6258 vdd.n1951 vdd.n1934 0.155672
R6259 vdd.n1951 vdd.n1950 0.155672
R6260 vdd.n1950 vdd.n1938 0.155672
R6261 vdd.n1943 vdd.n1938 0.155672
R6262 vdd.n1128 vdd.n1120 0.152939
R6263 vdd.n1132 vdd.n1128 0.152939
R6264 vdd.n1133 vdd.n1132 0.152939
R6265 vdd.n1134 vdd.n1133 0.152939
R6266 vdd.n1135 vdd.n1134 0.152939
R6267 vdd.n1139 vdd.n1135 0.152939
R6268 vdd.n1140 vdd.n1139 0.152939
R6269 vdd.n1141 vdd.n1140 0.152939
R6270 vdd.n1142 vdd.n1141 0.152939
R6271 vdd.n1146 vdd.n1142 0.152939
R6272 vdd.n1147 vdd.n1146 0.152939
R6273 vdd.n1148 vdd.n1147 0.152939
R6274 vdd.n2345 vdd.n1148 0.152939
R6275 vdd.n2345 vdd.n2344 0.152939
R6276 vdd.n2344 vdd.n2343 0.152939
R6277 vdd.n2343 vdd.n1154 0.152939
R6278 vdd.n1159 vdd.n1154 0.152939
R6279 vdd.n1160 vdd.n1159 0.152939
R6280 vdd.n1161 vdd.n1160 0.152939
R6281 vdd.n1165 vdd.n1161 0.152939
R6282 vdd.n1166 vdd.n1165 0.152939
R6283 vdd.n1167 vdd.n1166 0.152939
R6284 vdd.n1168 vdd.n1167 0.152939
R6285 vdd.n1172 vdd.n1168 0.152939
R6286 vdd.n1173 vdd.n1172 0.152939
R6287 vdd.n1174 vdd.n1173 0.152939
R6288 vdd.n1175 vdd.n1174 0.152939
R6289 vdd.n1179 vdd.n1175 0.152939
R6290 vdd.n1180 vdd.n1179 0.152939
R6291 vdd.n1181 vdd.n1180 0.152939
R6292 vdd.n1182 vdd.n1181 0.152939
R6293 vdd.n1186 vdd.n1182 0.152939
R6294 vdd.n1187 vdd.n1186 0.152939
R6295 vdd.n1188 vdd.n1187 0.152939
R6296 vdd.n2306 vdd.n1188 0.152939
R6297 vdd.n2306 vdd.n2305 0.152939
R6298 vdd.n2305 vdd.n2304 0.152939
R6299 vdd.n2304 vdd.n1194 0.152939
R6300 vdd.n1199 vdd.n1194 0.152939
R6301 vdd.n1200 vdd.n1199 0.152939
R6302 vdd.n1201 vdd.n1200 0.152939
R6303 vdd.n1205 vdd.n1201 0.152939
R6304 vdd.n1206 vdd.n1205 0.152939
R6305 vdd.n1207 vdd.n1206 0.152939
R6306 vdd.n1208 vdd.n1207 0.152939
R6307 vdd.n1212 vdd.n1208 0.152939
R6308 vdd.n1213 vdd.n1212 0.152939
R6309 vdd.n1214 vdd.n1213 0.152939
R6310 vdd.n1215 vdd.n1214 0.152939
R6311 vdd.n1219 vdd.n1215 0.152939
R6312 vdd.n1220 vdd.n1219 0.152939
R6313 vdd.n2380 vdd.n1123 0.152939
R6314 vdd.n2176 vdd.n1485 0.152939
R6315 vdd.n2191 vdd.n1485 0.152939
R6316 vdd.n2192 vdd.n2191 0.152939
R6317 vdd.n2193 vdd.n2192 0.152939
R6318 vdd.n2193 vdd.n1474 0.152939
R6319 vdd.n2208 vdd.n1474 0.152939
R6320 vdd.n2209 vdd.n2208 0.152939
R6321 vdd.n2210 vdd.n2209 0.152939
R6322 vdd.n2210 vdd.n1463 0.152939
R6323 vdd.n2224 vdd.n1463 0.152939
R6324 vdd.n2225 vdd.n2224 0.152939
R6325 vdd.n2226 vdd.n2225 0.152939
R6326 vdd.n2226 vdd.n1451 0.152939
R6327 vdd.n2241 vdd.n1451 0.152939
R6328 vdd.n2242 vdd.n2241 0.152939
R6329 vdd.n2243 vdd.n2242 0.152939
R6330 vdd.n2243 vdd.n1439 0.152939
R6331 vdd.n2260 vdd.n1439 0.152939
R6332 vdd.n2261 vdd.n2260 0.152939
R6333 vdd.n2262 vdd.n2261 0.152939
R6334 vdd.n735 vdd.n730 0.152939
R6335 vdd.n736 vdd.n735 0.152939
R6336 vdd.n737 vdd.n736 0.152939
R6337 vdd.n738 vdd.n737 0.152939
R6338 vdd.n739 vdd.n738 0.152939
R6339 vdd.n740 vdd.n739 0.152939
R6340 vdd.n741 vdd.n740 0.152939
R6341 vdd.n742 vdd.n741 0.152939
R6342 vdd.n743 vdd.n742 0.152939
R6343 vdd.n744 vdd.n743 0.152939
R6344 vdd.n745 vdd.n744 0.152939
R6345 vdd.n746 vdd.n745 0.152939
R6346 vdd.n3275 vdd.n746 0.152939
R6347 vdd.n3275 vdd.n3274 0.152939
R6348 vdd.n3274 vdd.n3273 0.152939
R6349 vdd.n3273 vdd.n748 0.152939
R6350 vdd.n749 vdd.n748 0.152939
R6351 vdd.n750 vdd.n749 0.152939
R6352 vdd.n751 vdd.n750 0.152939
R6353 vdd.n752 vdd.n751 0.152939
R6354 vdd.n753 vdd.n752 0.152939
R6355 vdd.n754 vdd.n753 0.152939
R6356 vdd.n755 vdd.n754 0.152939
R6357 vdd.n756 vdd.n755 0.152939
R6358 vdd.n757 vdd.n756 0.152939
R6359 vdd.n758 vdd.n757 0.152939
R6360 vdd.n759 vdd.n758 0.152939
R6361 vdd.n760 vdd.n759 0.152939
R6362 vdd.n761 vdd.n760 0.152939
R6363 vdd.n762 vdd.n761 0.152939
R6364 vdd.n763 vdd.n762 0.152939
R6365 vdd.n764 vdd.n763 0.152939
R6366 vdd.n765 vdd.n764 0.152939
R6367 vdd.n766 vdd.n765 0.152939
R6368 vdd.n3229 vdd.n766 0.152939
R6369 vdd.n3229 vdd.n3228 0.152939
R6370 vdd.n3228 vdd.n3227 0.152939
R6371 vdd.n3227 vdd.n770 0.152939
R6372 vdd.n771 vdd.n770 0.152939
R6373 vdd.n772 vdd.n771 0.152939
R6374 vdd.n773 vdd.n772 0.152939
R6375 vdd.n774 vdd.n773 0.152939
R6376 vdd.n775 vdd.n774 0.152939
R6377 vdd.n776 vdd.n775 0.152939
R6378 vdd.n777 vdd.n776 0.152939
R6379 vdd.n778 vdd.n777 0.152939
R6380 vdd.n779 vdd.n778 0.152939
R6381 vdd.n780 vdd.n779 0.152939
R6382 vdd.n781 vdd.n780 0.152939
R6383 vdd.n782 vdd.n781 0.152939
R6384 vdd.n783 vdd.n782 0.152939
R6385 vdd.n727 vdd.n726 0.152939
R6386 vdd.n3326 vdd.n682 0.152939
R6387 vdd.n3327 vdd.n3326 0.152939
R6388 vdd.n3328 vdd.n3327 0.152939
R6389 vdd.n3328 vdd.n670 0.152939
R6390 vdd.n3343 vdd.n670 0.152939
R6391 vdd.n3344 vdd.n3343 0.152939
R6392 vdd.n3345 vdd.n3344 0.152939
R6393 vdd.n3345 vdd.n659 0.152939
R6394 vdd.n3359 vdd.n659 0.152939
R6395 vdd.n3360 vdd.n3359 0.152939
R6396 vdd.n3361 vdd.n3360 0.152939
R6397 vdd.n3361 vdd.n647 0.152939
R6398 vdd.n3376 vdd.n647 0.152939
R6399 vdd.n3377 vdd.n3376 0.152939
R6400 vdd.n3378 vdd.n3377 0.152939
R6401 vdd.n3378 vdd.n636 0.152939
R6402 vdd.n3395 vdd.n636 0.152939
R6403 vdd.n3396 vdd.n3395 0.152939
R6404 vdd.n3397 vdd.n3396 0.152939
R6405 vdd.n3397 vdd.n334 0.152939
R6406 vdd.n3490 vdd.n335 0.152939
R6407 vdd.n346 vdd.n335 0.152939
R6408 vdd.n347 vdd.n346 0.152939
R6409 vdd.n348 vdd.n347 0.152939
R6410 vdd.n355 vdd.n348 0.152939
R6411 vdd.n356 vdd.n355 0.152939
R6412 vdd.n357 vdd.n356 0.152939
R6413 vdd.n358 vdd.n357 0.152939
R6414 vdd.n366 vdd.n358 0.152939
R6415 vdd.n367 vdd.n366 0.152939
R6416 vdd.n368 vdd.n367 0.152939
R6417 vdd.n369 vdd.n368 0.152939
R6418 vdd.n377 vdd.n369 0.152939
R6419 vdd.n378 vdd.n377 0.152939
R6420 vdd.n379 vdd.n378 0.152939
R6421 vdd.n380 vdd.n379 0.152939
R6422 vdd.n388 vdd.n380 0.152939
R6423 vdd.n389 vdd.n388 0.152939
R6424 vdd.n390 vdd.n389 0.152939
R6425 vdd.n391 vdd.n390 0.152939
R6426 vdd.n464 vdd.n463 0.152939
R6427 vdd.n470 vdd.n463 0.152939
R6428 vdd.n471 vdd.n470 0.152939
R6429 vdd.n472 vdd.n471 0.152939
R6430 vdd.n472 vdd.n461 0.152939
R6431 vdd.n480 vdd.n461 0.152939
R6432 vdd.n481 vdd.n480 0.152939
R6433 vdd.n482 vdd.n481 0.152939
R6434 vdd.n482 vdd.n459 0.152939
R6435 vdd.n490 vdd.n459 0.152939
R6436 vdd.n491 vdd.n490 0.152939
R6437 vdd.n492 vdd.n491 0.152939
R6438 vdd.n492 vdd.n457 0.152939
R6439 vdd.n500 vdd.n457 0.152939
R6440 vdd.n501 vdd.n500 0.152939
R6441 vdd.n502 vdd.n501 0.152939
R6442 vdd.n502 vdd.n455 0.152939
R6443 vdd.n510 vdd.n455 0.152939
R6444 vdd.n511 vdd.n510 0.152939
R6445 vdd.n512 vdd.n511 0.152939
R6446 vdd.n512 vdd.n451 0.152939
R6447 vdd.n520 vdd.n451 0.152939
R6448 vdd.n521 vdd.n520 0.152939
R6449 vdd.n522 vdd.n521 0.152939
R6450 vdd.n522 vdd.n449 0.152939
R6451 vdd.n530 vdd.n449 0.152939
R6452 vdd.n531 vdd.n530 0.152939
R6453 vdd.n532 vdd.n531 0.152939
R6454 vdd.n532 vdd.n447 0.152939
R6455 vdd.n540 vdd.n447 0.152939
R6456 vdd.n541 vdd.n540 0.152939
R6457 vdd.n542 vdd.n541 0.152939
R6458 vdd.n542 vdd.n445 0.152939
R6459 vdd.n550 vdd.n445 0.152939
R6460 vdd.n551 vdd.n550 0.152939
R6461 vdd.n552 vdd.n551 0.152939
R6462 vdd.n552 vdd.n443 0.152939
R6463 vdd.n560 vdd.n443 0.152939
R6464 vdd.n561 vdd.n560 0.152939
R6465 vdd.n562 vdd.n561 0.152939
R6466 vdd.n562 vdd.n439 0.152939
R6467 vdd.n570 vdd.n439 0.152939
R6468 vdd.n571 vdd.n570 0.152939
R6469 vdd.n572 vdd.n571 0.152939
R6470 vdd.n572 vdd.n437 0.152939
R6471 vdd.n580 vdd.n437 0.152939
R6472 vdd.n581 vdd.n580 0.152939
R6473 vdd.n582 vdd.n581 0.152939
R6474 vdd.n582 vdd.n435 0.152939
R6475 vdd.n590 vdd.n435 0.152939
R6476 vdd.n591 vdd.n590 0.152939
R6477 vdd.n592 vdd.n591 0.152939
R6478 vdd.n592 vdd.n433 0.152939
R6479 vdd.n600 vdd.n433 0.152939
R6480 vdd.n601 vdd.n600 0.152939
R6481 vdd.n602 vdd.n601 0.152939
R6482 vdd.n602 vdd.n431 0.152939
R6483 vdd.n610 vdd.n431 0.152939
R6484 vdd.n611 vdd.n610 0.152939
R6485 vdd.n612 vdd.n611 0.152939
R6486 vdd.n612 vdd.n429 0.152939
R6487 vdd.n619 vdd.n429 0.152939
R6488 vdd.n3442 vdd.n619 0.152939
R6489 vdd.n3320 vdd.n3319 0.152939
R6490 vdd.n3320 vdd.n675 0.152939
R6491 vdd.n3334 vdd.n675 0.152939
R6492 vdd.n3335 vdd.n3334 0.152939
R6493 vdd.n3336 vdd.n3335 0.152939
R6494 vdd.n3336 vdd.n665 0.152939
R6495 vdd.n3351 vdd.n665 0.152939
R6496 vdd.n3352 vdd.n3351 0.152939
R6497 vdd.n3353 vdd.n3352 0.152939
R6498 vdd.n3353 vdd.n652 0.152939
R6499 vdd.n3367 vdd.n652 0.152939
R6500 vdd.n3368 vdd.n3367 0.152939
R6501 vdd.n3369 vdd.n3368 0.152939
R6502 vdd.n3369 vdd.n641 0.152939
R6503 vdd.n3384 vdd.n641 0.152939
R6504 vdd.n3385 vdd.n3384 0.152939
R6505 vdd.n3386 vdd.n3385 0.152939
R6506 vdd.n3388 vdd.n3386 0.152939
R6507 vdd.n3388 vdd.n3387 0.152939
R6508 vdd.n3387 vdd.n630 0.152939
R6509 vdd.n3405 vdd.n630 0.152939
R6510 vdd.n3406 vdd.n3405 0.152939
R6511 vdd.n3407 vdd.n3406 0.152939
R6512 vdd.n3407 vdd.n628 0.152939
R6513 vdd.n3412 vdd.n628 0.152939
R6514 vdd.n3413 vdd.n3412 0.152939
R6515 vdd.n3414 vdd.n3413 0.152939
R6516 vdd.n3414 vdd.n626 0.152939
R6517 vdd.n3419 vdd.n626 0.152939
R6518 vdd.n3420 vdd.n3419 0.152939
R6519 vdd.n3421 vdd.n3420 0.152939
R6520 vdd.n3421 vdd.n624 0.152939
R6521 vdd.n3427 vdd.n624 0.152939
R6522 vdd.n3428 vdd.n3427 0.152939
R6523 vdd.n3429 vdd.n3428 0.152939
R6524 vdd.n3429 vdd.n622 0.152939
R6525 vdd.n3434 vdd.n622 0.152939
R6526 vdd.n3435 vdd.n3434 0.152939
R6527 vdd.n3436 vdd.n3435 0.152939
R6528 vdd.n3436 vdd.n620 0.152939
R6529 vdd.n3441 vdd.n620 0.152939
R6530 vdd.n3318 vdd.n687 0.152939
R6531 vdd.n2273 vdd.n1424 0.152939
R6532 vdd.n1792 vdd.n1548 0.152939
R6533 vdd.n1793 vdd.n1792 0.152939
R6534 vdd.n1794 vdd.n1793 0.152939
R6535 vdd.n1794 vdd.n1536 0.152939
R6536 vdd.n1809 vdd.n1536 0.152939
R6537 vdd.n1810 vdd.n1809 0.152939
R6538 vdd.n1811 vdd.n1810 0.152939
R6539 vdd.n1811 vdd.n1526 0.152939
R6540 vdd.n1826 vdd.n1526 0.152939
R6541 vdd.n1827 vdd.n1826 0.152939
R6542 vdd.n1828 vdd.n1827 0.152939
R6543 vdd.n1828 vdd.n1513 0.152939
R6544 vdd.n1842 vdd.n1513 0.152939
R6545 vdd.n1843 vdd.n1842 0.152939
R6546 vdd.n1844 vdd.n1843 0.152939
R6547 vdd.n1844 vdd.n1502 0.152939
R6548 vdd.n1859 vdd.n1502 0.152939
R6549 vdd.n1860 vdd.n1859 0.152939
R6550 vdd.n1861 vdd.n1860 0.152939
R6551 vdd.n1861 vdd.n1491 0.152939
R6552 vdd.n2182 vdd.n1491 0.152939
R6553 vdd.n2183 vdd.n2182 0.152939
R6554 vdd.n2184 vdd.n2183 0.152939
R6555 vdd.n2184 vdd.n1479 0.152939
R6556 vdd.n2199 vdd.n1479 0.152939
R6557 vdd.n2200 vdd.n2199 0.152939
R6558 vdd.n2201 vdd.n2200 0.152939
R6559 vdd.n2201 vdd.n1469 0.152939
R6560 vdd.n2216 vdd.n1469 0.152939
R6561 vdd.n2217 vdd.n2216 0.152939
R6562 vdd.n2218 vdd.n2217 0.152939
R6563 vdd.n2218 vdd.n1456 0.152939
R6564 vdd.n2232 vdd.n1456 0.152939
R6565 vdd.n2233 vdd.n2232 0.152939
R6566 vdd.n2234 vdd.n2233 0.152939
R6567 vdd.n2234 vdd.n1446 0.152939
R6568 vdd.n2249 vdd.n1446 0.152939
R6569 vdd.n2250 vdd.n2249 0.152939
R6570 vdd.n2253 vdd.n2250 0.152939
R6571 vdd.n2253 vdd.n2252 0.152939
R6572 vdd.n2252 vdd.n2251 0.152939
R6573 vdd.n1784 vdd.n1553 0.152939
R6574 vdd.n1777 vdd.n1553 0.152939
R6575 vdd.n1777 vdd.n1776 0.152939
R6576 vdd.n1776 vdd.n1775 0.152939
R6577 vdd.n1775 vdd.n1590 0.152939
R6578 vdd.n1771 vdd.n1590 0.152939
R6579 vdd.n1771 vdd.n1770 0.152939
R6580 vdd.n1770 vdd.n1769 0.152939
R6581 vdd.n1769 vdd.n1596 0.152939
R6582 vdd.n1765 vdd.n1596 0.152939
R6583 vdd.n1765 vdd.n1764 0.152939
R6584 vdd.n1764 vdd.n1763 0.152939
R6585 vdd.n1763 vdd.n1602 0.152939
R6586 vdd.n1759 vdd.n1602 0.152939
R6587 vdd.n1759 vdd.n1758 0.152939
R6588 vdd.n1758 vdd.n1757 0.152939
R6589 vdd.n1757 vdd.n1608 0.152939
R6590 vdd.n1753 vdd.n1608 0.152939
R6591 vdd.n1753 vdd.n1752 0.152939
R6592 vdd.n1752 vdd.n1751 0.152939
R6593 vdd.n1751 vdd.n1616 0.152939
R6594 vdd.n1747 vdd.n1616 0.152939
R6595 vdd.n1747 vdd.n1746 0.152939
R6596 vdd.n1746 vdd.n1745 0.152939
R6597 vdd.n1745 vdd.n1622 0.152939
R6598 vdd.n1741 vdd.n1622 0.152939
R6599 vdd.n1741 vdd.n1740 0.152939
R6600 vdd.n1740 vdd.n1739 0.152939
R6601 vdd.n1739 vdd.n1628 0.152939
R6602 vdd.n1735 vdd.n1628 0.152939
R6603 vdd.n1735 vdd.n1734 0.152939
R6604 vdd.n1734 vdd.n1733 0.152939
R6605 vdd.n1733 vdd.n1634 0.152939
R6606 vdd.n1729 vdd.n1634 0.152939
R6607 vdd.n1729 vdd.n1728 0.152939
R6608 vdd.n1728 vdd.n1727 0.152939
R6609 vdd.n1727 vdd.n1640 0.152939
R6610 vdd.n1723 vdd.n1640 0.152939
R6611 vdd.n1723 vdd.n1722 0.152939
R6612 vdd.n1722 vdd.n1721 0.152939
R6613 vdd.n1721 vdd.n1646 0.152939
R6614 vdd.n1714 vdd.n1646 0.152939
R6615 vdd.n1714 vdd.n1713 0.152939
R6616 vdd.n1713 vdd.n1712 0.152939
R6617 vdd.n1712 vdd.n1651 0.152939
R6618 vdd.n1708 vdd.n1651 0.152939
R6619 vdd.n1708 vdd.n1707 0.152939
R6620 vdd.n1707 vdd.n1706 0.152939
R6621 vdd.n1706 vdd.n1657 0.152939
R6622 vdd.n1702 vdd.n1657 0.152939
R6623 vdd.n1702 vdd.n1701 0.152939
R6624 vdd.n1701 vdd.n1700 0.152939
R6625 vdd.n1700 vdd.n1663 0.152939
R6626 vdd.n1696 vdd.n1663 0.152939
R6627 vdd.n1696 vdd.n1695 0.152939
R6628 vdd.n1695 vdd.n1694 0.152939
R6629 vdd.n1694 vdd.n1669 0.152939
R6630 vdd.n1690 vdd.n1669 0.152939
R6631 vdd.n1690 vdd.n1689 0.152939
R6632 vdd.n1689 vdd.n1688 0.152939
R6633 vdd.n1688 vdd.n1675 0.152939
R6634 vdd.n1684 vdd.n1675 0.152939
R6635 vdd.n1684 vdd.n1683 0.152939
R6636 vdd.n1786 vdd.n1785 0.152939
R6637 vdd.n1786 vdd.n1542 0.152939
R6638 vdd.n1801 vdd.n1542 0.152939
R6639 vdd.n1802 vdd.n1801 0.152939
R6640 vdd.n1803 vdd.n1802 0.152939
R6641 vdd.n1803 vdd.n1531 0.152939
R6642 vdd.n1818 vdd.n1531 0.152939
R6643 vdd.n1819 vdd.n1818 0.152939
R6644 vdd.n1820 vdd.n1819 0.152939
R6645 vdd.n1820 vdd.n1520 0.152939
R6646 vdd.n1834 vdd.n1520 0.152939
R6647 vdd.n1835 vdd.n1834 0.152939
R6648 vdd.n1836 vdd.n1835 0.152939
R6649 vdd.n1836 vdd.n1508 0.152939
R6650 vdd.n1851 vdd.n1508 0.152939
R6651 vdd.n1852 vdd.n1851 0.152939
R6652 vdd.n1853 vdd.n1852 0.152939
R6653 vdd.n1853 vdd.n1497 0.152939
R6654 vdd.n1867 vdd.n1497 0.152939
R6655 vdd.n1868 vdd.n1867 0.152939
R6656 vdd.n1789 vdd.t91 0.113865
R6657 vdd.t77 vdd.n386 0.113865
R6658 vdd.n2381 vdd.n2380 0.110256
R6659 vdd.n3308 vdd.n727 0.110256
R6660 vdd.n3185 vdd.n687 0.110256
R6661 vdd.n2274 vdd.n2273 0.110256
R6662 vdd.n2176 vdd.n2175 0.0695946
R6663 vdd.n3491 vdd.n334 0.0695946
R6664 vdd.n3491 vdd.n3490 0.0695946
R6665 vdd.n2175 vdd.n1868 0.0695946
R6666 vdd.n2381 vdd.n1120 0.0431829
R6667 vdd.n2274 vdd.n1220 0.0431829
R6668 vdd.n3308 vdd.n730 0.0431829
R6669 vdd.n3185 vdd.n783 0.0431829
R6670 vdd vdd.n28 0.00833333
R6671 CSoutput.n19 CSoutput.t233 184.661
R6672 CSoutput.n78 CSoutput.n77 165.8
R6673 CSoutput.n76 CSoutput.n0 165.8
R6674 CSoutput.n75 CSoutput.n74 165.8
R6675 CSoutput.n73 CSoutput.n72 165.8
R6676 CSoutput.n71 CSoutput.n2 165.8
R6677 CSoutput.n69 CSoutput.n68 165.8
R6678 CSoutput.n67 CSoutput.n3 165.8
R6679 CSoutput.n66 CSoutput.n65 165.8
R6680 CSoutput.n63 CSoutput.n4 165.8
R6681 CSoutput.n61 CSoutput.n60 165.8
R6682 CSoutput.n59 CSoutput.n5 165.8
R6683 CSoutput.n58 CSoutput.n57 165.8
R6684 CSoutput.n55 CSoutput.n6 165.8
R6685 CSoutput.n54 CSoutput.n53 165.8
R6686 CSoutput.n52 CSoutput.n51 165.8
R6687 CSoutput.n50 CSoutput.n8 165.8
R6688 CSoutput.n48 CSoutput.n47 165.8
R6689 CSoutput.n46 CSoutput.n9 165.8
R6690 CSoutput.n45 CSoutput.n44 165.8
R6691 CSoutput.n42 CSoutput.n10 165.8
R6692 CSoutput.n41 CSoutput.n40 165.8
R6693 CSoutput.n39 CSoutput.n38 165.8
R6694 CSoutput.n37 CSoutput.n12 165.8
R6695 CSoutput.n35 CSoutput.n34 165.8
R6696 CSoutput.n33 CSoutput.n13 165.8
R6697 CSoutput.n32 CSoutput.n31 165.8
R6698 CSoutput.n29 CSoutput.n14 165.8
R6699 CSoutput.n28 CSoutput.n27 165.8
R6700 CSoutput.n26 CSoutput.n25 165.8
R6701 CSoutput.n24 CSoutput.n16 165.8
R6702 CSoutput.n22 CSoutput.n21 165.8
R6703 CSoutput.n20 CSoutput.n17 165.8
R6704 CSoutput.n77 CSoutput.t235 162.194
R6705 CSoutput.n18 CSoutput.t230 120.501
R6706 CSoutput.n23 CSoutput.t224 120.501
R6707 CSoutput.n15 CSoutput.t219 120.501
R6708 CSoutput.n30 CSoutput.t231 120.501
R6709 CSoutput.n36 CSoutput.t232 120.501
R6710 CSoutput.n11 CSoutput.t221 120.501
R6711 CSoutput.n43 CSoutput.t217 120.501
R6712 CSoutput.n49 CSoutput.t234 120.501
R6713 CSoutput.n7 CSoutput.t225 120.501
R6714 CSoutput.n56 CSoutput.t227 120.501
R6715 CSoutput.n62 CSoutput.t236 120.501
R6716 CSoutput.n64 CSoutput.t228 120.501
R6717 CSoutput.n70 CSoutput.t229 120.501
R6718 CSoutput.n1 CSoutput.t222 120.501
R6719 CSoutput.n330 CSoutput.n328 103.469
R6720 CSoutput.n310 CSoutput.n308 103.469
R6721 CSoutput.n291 CSoutput.n289 103.469
R6722 CSoutput.n120 CSoutput.n118 103.469
R6723 CSoutput.n100 CSoutput.n98 103.469
R6724 CSoutput.n81 CSoutput.n79 103.469
R6725 CSoutput.n344 CSoutput.n343 103.111
R6726 CSoutput.n342 CSoutput.n341 103.111
R6727 CSoutput.n340 CSoutput.n339 103.111
R6728 CSoutput.n338 CSoutput.n337 103.111
R6729 CSoutput.n336 CSoutput.n335 103.111
R6730 CSoutput.n334 CSoutput.n333 103.111
R6731 CSoutput.n332 CSoutput.n331 103.111
R6732 CSoutput.n330 CSoutput.n329 103.111
R6733 CSoutput.n326 CSoutput.n325 103.111
R6734 CSoutput.n324 CSoutput.n323 103.111
R6735 CSoutput.n322 CSoutput.n321 103.111
R6736 CSoutput.n320 CSoutput.n319 103.111
R6737 CSoutput.n318 CSoutput.n317 103.111
R6738 CSoutput.n316 CSoutput.n315 103.111
R6739 CSoutput.n314 CSoutput.n313 103.111
R6740 CSoutput.n312 CSoutput.n311 103.111
R6741 CSoutput.n310 CSoutput.n309 103.111
R6742 CSoutput.n307 CSoutput.n306 103.111
R6743 CSoutput.n305 CSoutput.n304 103.111
R6744 CSoutput.n303 CSoutput.n302 103.111
R6745 CSoutput.n301 CSoutput.n300 103.111
R6746 CSoutput.n299 CSoutput.n298 103.111
R6747 CSoutput.n297 CSoutput.n296 103.111
R6748 CSoutput.n295 CSoutput.n294 103.111
R6749 CSoutput.n293 CSoutput.n292 103.111
R6750 CSoutput.n291 CSoutput.n290 103.111
R6751 CSoutput.n120 CSoutput.n119 103.111
R6752 CSoutput.n122 CSoutput.n121 103.111
R6753 CSoutput.n124 CSoutput.n123 103.111
R6754 CSoutput.n126 CSoutput.n125 103.111
R6755 CSoutput.n128 CSoutput.n127 103.111
R6756 CSoutput.n130 CSoutput.n129 103.111
R6757 CSoutput.n132 CSoutput.n131 103.111
R6758 CSoutput.n134 CSoutput.n133 103.111
R6759 CSoutput.n136 CSoutput.n135 103.111
R6760 CSoutput.n100 CSoutput.n99 103.111
R6761 CSoutput.n102 CSoutput.n101 103.111
R6762 CSoutput.n104 CSoutput.n103 103.111
R6763 CSoutput.n106 CSoutput.n105 103.111
R6764 CSoutput.n108 CSoutput.n107 103.111
R6765 CSoutput.n110 CSoutput.n109 103.111
R6766 CSoutput.n112 CSoutput.n111 103.111
R6767 CSoutput.n114 CSoutput.n113 103.111
R6768 CSoutput.n116 CSoutput.n115 103.111
R6769 CSoutput.n81 CSoutput.n80 103.111
R6770 CSoutput.n83 CSoutput.n82 103.111
R6771 CSoutput.n85 CSoutput.n84 103.111
R6772 CSoutput.n87 CSoutput.n86 103.111
R6773 CSoutput.n89 CSoutput.n88 103.111
R6774 CSoutput.n91 CSoutput.n90 103.111
R6775 CSoutput.n93 CSoutput.n92 103.111
R6776 CSoutput.n95 CSoutput.n94 103.111
R6777 CSoutput.n97 CSoutput.n96 103.111
R6778 CSoutput.n346 CSoutput.n345 103.111
R6779 CSoutput.n382 CSoutput.n380 81.5057
R6780 CSoutput.n366 CSoutput.n364 81.5057
R6781 CSoutput.n351 CSoutput.n349 81.5057
R6782 CSoutput.n430 CSoutput.n428 81.5057
R6783 CSoutput.n414 CSoutput.n412 81.5057
R6784 CSoutput.n399 CSoutput.n397 81.5057
R6785 CSoutput.n394 CSoutput.n393 80.9324
R6786 CSoutput.n392 CSoutput.n391 80.9324
R6787 CSoutput.n390 CSoutput.n389 80.9324
R6788 CSoutput.n388 CSoutput.n387 80.9324
R6789 CSoutput.n386 CSoutput.n385 80.9324
R6790 CSoutput.n384 CSoutput.n383 80.9324
R6791 CSoutput.n382 CSoutput.n381 80.9324
R6792 CSoutput.n378 CSoutput.n377 80.9324
R6793 CSoutput.n376 CSoutput.n375 80.9324
R6794 CSoutput.n374 CSoutput.n373 80.9324
R6795 CSoutput.n372 CSoutput.n371 80.9324
R6796 CSoutput.n370 CSoutput.n369 80.9324
R6797 CSoutput.n368 CSoutput.n367 80.9324
R6798 CSoutput.n366 CSoutput.n365 80.9324
R6799 CSoutput.n363 CSoutput.n362 80.9324
R6800 CSoutput.n361 CSoutput.n360 80.9324
R6801 CSoutput.n359 CSoutput.n358 80.9324
R6802 CSoutput.n357 CSoutput.n356 80.9324
R6803 CSoutput.n355 CSoutput.n354 80.9324
R6804 CSoutput.n353 CSoutput.n352 80.9324
R6805 CSoutput.n351 CSoutput.n350 80.9324
R6806 CSoutput.n430 CSoutput.n429 80.9324
R6807 CSoutput.n432 CSoutput.n431 80.9324
R6808 CSoutput.n434 CSoutput.n433 80.9324
R6809 CSoutput.n436 CSoutput.n435 80.9324
R6810 CSoutput.n438 CSoutput.n437 80.9324
R6811 CSoutput.n440 CSoutput.n439 80.9324
R6812 CSoutput.n442 CSoutput.n441 80.9324
R6813 CSoutput.n414 CSoutput.n413 80.9324
R6814 CSoutput.n416 CSoutput.n415 80.9324
R6815 CSoutput.n418 CSoutput.n417 80.9324
R6816 CSoutput.n420 CSoutput.n419 80.9324
R6817 CSoutput.n422 CSoutput.n421 80.9324
R6818 CSoutput.n424 CSoutput.n423 80.9324
R6819 CSoutput.n426 CSoutput.n425 80.9324
R6820 CSoutput.n399 CSoutput.n398 80.9324
R6821 CSoutput.n401 CSoutput.n400 80.9324
R6822 CSoutput.n403 CSoutput.n402 80.9324
R6823 CSoutput.n405 CSoutput.n404 80.9324
R6824 CSoutput.n407 CSoutput.n406 80.9324
R6825 CSoutput.n409 CSoutput.n408 80.9324
R6826 CSoutput.n411 CSoutput.n410 80.9324
R6827 CSoutput.n25 CSoutput.n24 48.1486
R6828 CSoutput.n69 CSoutput.n3 48.1486
R6829 CSoutput.n38 CSoutput.n37 48.1486
R6830 CSoutput.n42 CSoutput.n41 48.1486
R6831 CSoutput.n51 CSoutput.n50 48.1486
R6832 CSoutput.n55 CSoutput.n54 48.1486
R6833 CSoutput.n22 CSoutput.n17 46.462
R6834 CSoutput.n72 CSoutput.n71 46.462
R6835 CSoutput.n20 CSoutput.n19 44.9055
R6836 CSoutput.n29 CSoutput.n28 43.7635
R6837 CSoutput.n65 CSoutput.n63 43.7635
R6838 CSoutput.n35 CSoutput.n13 41.7396
R6839 CSoutput.n57 CSoutput.n5 41.7396
R6840 CSoutput.n44 CSoutput.n9 37.0171
R6841 CSoutput.n48 CSoutput.n9 37.0171
R6842 CSoutput.n76 CSoutput.n75 34.9932
R6843 CSoutput.n31 CSoutput.n13 32.2947
R6844 CSoutput.n61 CSoutput.n5 32.2947
R6845 CSoutput.n30 CSoutput.n29 29.6014
R6846 CSoutput.n63 CSoutput.n62 29.6014
R6847 CSoutput.n19 CSoutput.n18 28.4085
R6848 CSoutput.n18 CSoutput.n17 25.1176
R6849 CSoutput.n72 CSoutput.n1 25.1176
R6850 CSoutput.n43 CSoutput.n42 22.0922
R6851 CSoutput.n50 CSoutput.n49 22.0922
R6852 CSoutput.n77 CSoutput.n76 21.8586
R6853 CSoutput.n37 CSoutput.n36 18.9681
R6854 CSoutput.n56 CSoutput.n55 18.9681
R6855 CSoutput.n25 CSoutput.n15 17.6292
R6856 CSoutput.n64 CSoutput.n3 17.6292
R6857 CSoutput.n24 CSoutput.n23 15.844
R6858 CSoutput.n70 CSoutput.n69 15.844
R6859 CSoutput.n38 CSoutput.n11 14.5051
R6860 CSoutput.n54 CSoutput.n7 14.5051
R6861 CSoutput.n445 CSoutput.n78 11.4982
R6862 CSoutput.n41 CSoutput.n11 11.3811
R6863 CSoutput.n51 CSoutput.n7 11.3811
R6864 CSoutput.n23 CSoutput.n22 10.0422
R6865 CSoutput.n71 CSoutput.n70 10.0422
R6866 CSoutput.n327 CSoutput.n307 9.25285
R6867 CSoutput.n117 CSoutput.n97 9.25285
R6868 CSoutput.n379 CSoutput.n363 8.98182
R6869 CSoutput.n427 CSoutput.n411 8.98182
R6870 CSoutput.n396 CSoutput.n348 8.67888
R6871 CSoutput.n28 CSoutput.n15 8.25698
R6872 CSoutput.n65 CSoutput.n64 8.25698
R6873 CSoutput.n348 CSoutput.n347 7.12641
R6874 CSoutput.n138 CSoutput.n137 7.12641
R6875 CSoutput.n36 CSoutput.n35 6.91809
R6876 CSoutput.n57 CSoutput.n56 6.91809
R6877 CSoutput.n396 CSoutput.n395 6.02792
R6878 CSoutput.n444 CSoutput.n443 6.02792
R6879 CSoutput.n395 CSoutput.n394 5.25266
R6880 CSoutput.n379 CSoutput.n378 5.25266
R6881 CSoutput.n443 CSoutput.n442 5.25266
R6882 CSoutput.n427 CSoutput.n426 5.25266
R6883 CSoutput.n347 CSoutput.n346 5.1449
R6884 CSoutput.n327 CSoutput.n326 5.1449
R6885 CSoutput.n137 CSoutput.n136 5.1449
R6886 CSoutput.n117 CSoutput.n116 5.1449
R6887 CSoutput.n445 CSoutput.n138 5.08644
R6888 CSoutput.n229 CSoutput.n182 4.5005
R6889 CSoutput.n198 CSoutput.n182 4.5005
R6890 CSoutput.n193 CSoutput.n177 4.5005
R6891 CSoutput.n193 CSoutput.n179 4.5005
R6892 CSoutput.n193 CSoutput.n176 4.5005
R6893 CSoutput.n193 CSoutput.n180 4.5005
R6894 CSoutput.n193 CSoutput.n175 4.5005
R6895 CSoutput.n193 CSoutput.t237 4.5005
R6896 CSoutput.n193 CSoutput.n174 4.5005
R6897 CSoutput.n193 CSoutput.n181 4.5005
R6898 CSoutput.n193 CSoutput.n182 4.5005
R6899 CSoutput.n191 CSoutput.n177 4.5005
R6900 CSoutput.n191 CSoutput.n179 4.5005
R6901 CSoutput.n191 CSoutput.n176 4.5005
R6902 CSoutput.n191 CSoutput.n180 4.5005
R6903 CSoutput.n191 CSoutput.n175 4.5005
R6904 CSoutput.n191 CSoutput.t237 4.5005
R6905 CSoutput.n191 CSoutput.n174 4.5005
R6906 CSoutput.n191 CSoutput.n181 4.5005
R6907 CSoutput.n191 CSoutput.n182 4.5005
R6908 CSoutput.n190 CSoutput.n177 4.5005
R6909 CSoutput.n190 CSoutput.n179 4.5005
R6910 CSoutput.n190 CSoutput.n176 4.5005
R6911 CSoutput.n190 CSoutput.n180 4.5005
R6912 CSoutput.n190 CSoutput.n175 4.5005
R6913 CSoutput.n190 CSoutput.t237 4.5005
R6914 CSoutput.n190 CSoutput.n174 4.5005
R6915 CSoutput.n190 CSoutput.n181 4.5005
R6916 CSoutput.n190 CSoutput.n182 4.5005
R6917 CSoutput.n275 CSoutput.n177 4.5005
R6918 CSoutput.n275 CSoutput.n179 4.5005
R6919 CSoutput.n275 CSoutput.n176 4.5005
R6920 CSoutput.n275 CSoutput.n180 4.5005
R6921 CSoutput.n275 CSoutput.n175 4.5005
R6922 CSoutput.n275 CSoutput.t237 4.5005
R6923 CSoutput.n275 CSoutput.n174 4.5005
R6924 CSoutput.n275 CSoutput.n181 4.5005
R6925 CSoutput.n275 CSoutput.n182 4.5005
R6926 CSoutput.n273 CSoutput.n177 4.5005
R6927 CSoutput.n273 CSoutput.n179 4.5005
R6928 CSoutput.n273 CSoutput.n176 4.5005
R6929 CSoutput.n273 CSoutput.n180 4.5005
R6930 CSoutput.n273 CSoutput.n175 4.5005
R6931 CSoutput.n273 CSoutput.t237 4.5005
R6932 CSoutput.n273 CSoutput.n174 4.5005
R6933 CSoutput.n273 CSoutput.n181 4.5005
R6934 CSoutput.n271 CSoutput.n177 4.5005
R6935 CSoutput.n271 CSoutput.n179 4.5005
R6936 CSoutput.n271 CSoutput.n176 4.5005
R6937 CSoutput.n271 CSoutput.n180 4.5005
R6938 CSoutput.n271 CSoutput.n175 4.5005
R6939 CSoutput.n271 CSoutput.t237 4.5005
R6940 CSoutput.n271 CSoutput.n174 4.5005
R6941 CSoutput.n271 CSoutput.n181 4.5005
R6942 CSoutput.n201 CSoutput.n177 4.5005
R6943 CSoutput.n201 CSoutput.n179 4.5005
R6944 CSoutput.n201 CSoutput.n176 4.5005
R6945 CSoutput.n201 CSoutput.n180 4.5005
R6946 CSoutput.n201 CSoutput.n175 4.5005
R6947 CSoutput.n201 CSoutput.t237 4.5005
R6948 CSoutput.n201 CSoutput.n174 4.5005
R6949 CSoutput.n201 CSoutput.n181 4.5005
R6950 CSoutput.n201 CSoutput.n182 4.5005
R6951 CSoutput.n200 CSoutput.n177 4.5005
R6952 CSoutput.n200 CSoutput.n179 4.5005
R6953 CSoutput.n200 CSoutput.n176 4.5005
R6954 CSoutput.n200 CSoutput.n180 4.5005
R6955 CSoutput.n200 CSoutput.n175 4.5005
R6956 CSoutput.n200 CSoutput.t237 4.5005
R6957 CSoutput.n200 CSoutput.n174 4.5005
R6958 CSoutput.n200 CSoutput.n181 4.5005
R6959 CSoutput.n200 CSoutput.n182 4.5005
R6960 CSoutput.n204 CSoutput.n177 4.5005
R6961 CSoutput.n204 CSoutput.n179 4.5005
R6962 CSoutput.n204 CSoutput.n176 4.5005
R6963 CSoutput.n204 CSoutput.n180 4.5005
R6964 CSoutput.n204 CSoutput.n175 4.5005
R6965 CSoutput.n204 CSoutput.t237 4.5005
R6966 CSoutput.n204 CSoutput.n174 4.5005
R6967 CSoutput.n204 CSoutput.n181 4.5005
R6968 CSoutput.n204 CSoutput.n182 4.5005
R6969 CSoutput.n203 CSoutput.n177 4.5005
R6970 CSoutput.n203 CSoutput.n179 4.5005
R6971 CSoutput.n203 CSoutput.n176 4.5005
R6972 CSoutput.n203 CSoutput.n180 4.5005
R6973 CSoutput.n203 CSoutput.n175 4.5005
R6974 CSoutput.n203 CSoutput.t237 4.5005
R6975 CSoutput.n203 CSoutput.n174 4.5005
R6976 CSoutput.n203 CSoutput.n181 4.5005
R6977 CSoutput.n203 CSoutput.n182 4.5005
R6978 CSoutput.n186 CSoutput.n177 4.5005
R6979 CSoutput.n186 CSoutput.n179 4.5005
R6980 CSoutput.n186 CSoutput.n176 4.5005
R6981 CSoutput.n186 CSoutput.n180 4.5005
R6982 CSoutput.n186 CSoutput.n175 4.5005
R6983 CSoutput.n186 CSoutput.t237 4.5005
R6984 CSoutput.n186 CSoutput.n174 4.5005
R6985 CSoutput.n186 CSoutput.n181 4.5005
R6986 CSoutput.n186 CSoutput.n182 4.5005
R6987 CSoutput.n278 CSoutput.n177 4.5005
R6988 CSoutput.n278 CSoutput.n179 4.5005
R6989 CSoutput.n278 CSoutput.n176 4.5005
R6990 CSoutput.n278 CSoutput.n180 4.5005
R6991 CSoutput.n278 CSoutput.n175 4.5005
R6992 CSoutput.n278 CSoutput.t237 4.5005
R6993 CSoutput.n278 CSoutput.n174 4.5005
R6994 CSoutput.n278 CSoutput.n181 4.5005
R6995 CSoutput.n278 CSoutput.n182 4.5005
R6996 CSoutput.n265 CSoutput.n236 4.5005
R6997 CSoutput.n265 CSoutput.n242 4.5005
R6998 CSoutput.n223 CSoutput.n212 4.5005
R6999 CSoutput.n223 CSoutput.n214 4.5005
R7000 CSoutput.n223 CSoutput.n211 4.5005
R7001 CSoutput.n223 CSoutput.n215 4.5005
R7002 CSoutput.n223 CSoutput.n210 4.5005
R7003 CSoutput.n223 CSoutput.t216 4.5005
R7004 CSoutput.n223 CSoutput.n209 4.5005
R7005 CSoutput.n223 CSoutput.n216 4.5005
R7006 CSoutput.n265 CSoutput.n223 4.5005
R7007 CSoutput.n244 CSoutput.n212 4.5005
R7008 CSoutput.n244 CSoutput.n214 4.5005
R7009 CSoutput.n244 CSoutput.n211 4.5005
R7010 CSoutput.n244 CSoutput.n215 4.5005
R7011 CSoutput.n244 CSoutput.n210 4.5005
R7012 CSoutput.n244 CSoutput.t216 4.5005
R7013 CSoutput.n244 CSoutput.n209 4.5005
R7014 CSoutput.n244 CSoutput.n216 4.5005
R7015 CSoutput.n265 CSoutput.n244 4.5005
R7016 CSoutput.n222 CSoutput.n212 4.5005
R7017 CSoutput.n222 CSoutput.n214 4.5005
R7018 CSoutput.n222 CSoutput.n211 4.5005
R7019 CSoutput.n222 CSoutput.n215 4.5005
R7020 CSoutput.n222 CSoutput.n210 4.5005
R7021 CSoutput.n222 CSoutput.t216 4.5005
R7022 CSoutput.n222 CSoutput.n209 4.5005
R7023 CSoutput.n222 CSoutput.n216 4.5005
R7024 CSoutput.n265 CSoutput.n222 4.5005
R7025 CSoutput.n246 CSoutput.n212 4.5005
R7026 CSoutput.n246 CSoutput.n214 4.5005
R7027 CSoutput.n246 CSoutput.n211 4.5005
R7028 CSoutput.n246 CSoutput.n215 4.5005
R7029 CSoutput.n246 CSoutput.n210 4.5005
R7030 CSoutput.n246 CSoutput.t216 4.5005
R7031 CSoutput.n246 CSoutput.n209 4.5005
R7032 CSoutput.n246 CSoutput.n216 4.5005
R7033 CSoutput.n265 CSoutput.n246 4.5005
R7034 CSoutput.n212 CSoutput.n207 4.5005
R7035 CSoutput.n214 CSoutput.n207 4.5005
R7036 CSoutput.n211 CSoutput.n207 4.5005
R7037 CSoutput.n215 CSoutput.n207 4.5005
R7038 CSoutput.n210 CSoutput.n207 4.5005
R7039 CSoutput.t216 CSoutput.n207 4.5005
R7040 CSoutput.n209 CSoutput.n207 4.5005
R7041 CSoutput.n216 CSoutput.n207 4.5005
R7042 CSoutput.n268 CSoutput.n212 4.5005
R7043 CSoutput.n268 CSoutput.n214 4.5005
R7044 CSoutput.n268 CSoutput.n211 4.5005
R7045 CSoutput.n268 CSoutput.n215 4.5005
R7046 CSoutput.n268 CSoutput.n210 4.5005
R7047 CSoutput.n268 CSoutput.t216 4.5005
R7048 CSoutput.n268 CSoutput.n209 4.5005
R7049 CSoutput.n268 CSoutput.n216 4.5005
R7050 CSoutput.n266 CSoutput.n212 4.5005
R7051 CSoutput.n266 CSoutput.n214 4.5005
R7052 CSoutput.n266 CSoutput.n211 4.5005
R7053 CSoutput.n266 CSoutput.n215 4.5005
R7054 CSoutput.n266 CSoutput.n210 4.5005
R7055 CSoutput.n266 CSoutput.t216 4.5005
R7056 CSoutput.n266 CSoutput.n209 4.5005
R7057 CSoutput.n266 CSoutput.n216 4.5005
R7058 CSoutput.n266 CSoutput.n265 4.5005
R7059 CSoutput.n248 CSoutput.n212 4.5005
R7060 CSoutput.n248 CSoutput.n214 4.5005
R7061 CSoutput.n248 CSoutput.n211 4.5005
R7062 CSoutput.n248 CSoutput.n215 4.5005
R7063 CSoutput.n248 CSoutput.n210 4.5005
R7064 CSoutput.n248 CSoutput.t216 4.5005
R7065 CSoutput.n248 CSoutput.n209 4.5005
R7066 CSoutput.n248 CSoutput.n216 4.5005
R7067 CSoutput.n265 CSoutput.n248 4.5005
R7068 CSoutput.n220 CSoutput.n212 4.5005
R7069 CSoutput.n220 CSoutput.n214 4.5005
R7070 CSoutput.n220 CSoutput.n211 4.5005
R7071 CSoutput.n220 CSoutput.n215 4.5005
R7072 CSoutput.n220 CSoutput.n210 4.5005
R7073 CSoutput.n220 CSoutput.t216 4.5005
R7074 CSoutput.n220 CSoutput.n209 4.5005
R7075 CSoutput.n220 CSoutput.n216 4.5005
R7076 CSoutput.n265 CSoutput.n220 4.5005
R7077 CSoutput.n250 CSoutput.n212 4.5005
R7078 CSoutput.n250 CSoutput.n214 4.5005
R7079 CSoutput.n250 CSoutput.n211 4.5005
R7080 CSoutput.n250 CSoutput.n215 4.5005
R7081 CSoutput.n250 CSoutput.n210 4.5005
R7082 CSoutput.n250 CSoutput.t216 4.5005
R7083 CSoutput.n250 CSoutput.n209 4.5005
R7084 CSoutput.n250 CSoutput.n216 4.5005
R7085 CSoutput.n265 CSoutput.n250 4.5005
R7086 CSoutput.n219 CSoutput.n212 4.5005
R7087 CSoutput.n219 CSoutput.n214 4.5005
R7088 CSoutput.n219 CSoutput.n211 4.5005
R7089 CSoutput.n219 CSoutput.n215 4.5005
R7090 CSoutput.n219 CSoutput.n210 4.5005
R7091 CSoutput.n219 CSoutput.t216 4.5005
R7092 CSoutput.n219 CSoutput.n209 4.5005
R7093 CSoutput.n219 CSoutput.n216 4.5005
R7094 CSoutput.n265 CSoutput.n219 4.5005
R7095 CSoutput.n264 CSoutput.n212 4.5005
R7096 CSoutput.n264 CSoutput.n214 4.5005
R7097 CSoutput.n264 CSoutput.n211 4.5005
R7098 CSoutput.n264 CSoutput.n215 4.5005
R7099 CSoutput.n264 CSoutput.n210 4.5005
R7100 CSoutput.n264 CSoutput.t216 4.5005
R7101 CSoutput.n264 CSoutput.n209 4.5005
R7102 CSoutput.n264 CSoutput.n216 4.5005
R7103 CSoutput.n265 CSoutput.n264 4.5005
R7104 CSoutput.n263 CSoutput.n148 4.5005
R7105 CSoutput.n164 CSoutput.n148 4.5005
R7106 CSoutput.n159 CSoutput.n143 4.5005
R7107 CSoutput.n159 CSoutput.n145 4.5005
R7108 CSoutput.n159 CSoutput.n142 4.5005
R7109 CSoutput.n159 CSoutput.n146 4.5005
R7110 CSoutput.n159 CSoutput.n141 4.5005
R7111 CSoutput.n159 CSoutput.t223 4.5005
R7112 CSoutput.n159 CSoutput.n140 4.5005
R7113 CSoutput.n159 CSoutput.n147 4.5005
R7114 CSoutput.n159 CSoutput.n148 4.5005
R7115 CSoutput.n157 CSoutput.n143 4.5005
R7116 CSoutput.n157 CSoutput.n145 4.5005
R7117 CSoutput.n157 CSoutput.n142 4.5005
R7118 CSoutput.n157 CSoutput.n146 4.5005
R7119 CSoutput.n157 CSoutput.n141 4.5005
R7120 CSoutput.n157 CSoutput.t223 4.5005
R7121 CSoutput.n157 CSoutput.n140 4.5005
R7122 CSoutput.n157 CSoutput.n147 4.5005
R7123 CSoutput.n157 CSoutput.n148 4.5005
R7124 CSoutput.n156 CSoutput.n143 4.5005
R7125 CSoutput.n156 CSoutput.n145 4.5005
R7126 CSoutput.n156 CSoutput.n142 4.5005
R7127 CSoutput.n156 CSoutput.n146 4.5005
R7128 CSoutput.n156 CSoutput.n141 4.5005
R7129 CSoutput.n156 CSoutput.t223 4.5005
R7130 CSoutput.n156 CSoutput.n140 4.5005
R7131 CSoutput.n156 CSoutput.n147 4.5005
R7132 CSoutput.n156 CSoutput.n148 4.5005
R7133 CSoutput.n285 CSoutput.n143 4.5005
R7134 CSoutput.n285 CSoutput.n145 4.5005
R7135 CSoutput.n285 CSoutput.n142 4.5005
R7136 CSoutput.n285 CSoutput.n146 4.5005
R7137 CSoutput.n285 CSoutput.n141 4.5005
R7138 CSoutput.n285 CSoutput.t223 4.5005
R7139 CSoutput.n285 CSoutput.n140 4.5005
R7140 CSoutput.n285 CSoutput.n147 4.5005
R7141 CSoutput.n285 CSoutput.n148 4.5005
R7142 CSoutput.n283 CSoutput.n143 4.5005
R7143 CSoutput.n283 CSoutput.n145 4.5005
R7144 CSoutput.n283 CSoutput.n142 4.5005
R7145 CSoutput.n283 CSoutput.n146 4.5005
R7146 CSoutput.n283 CSoutput.n141 4.5005
R7147 CSoutput.n283 CSoutput.t223 4.5005
R7148 CSoutput.n283 CSoutput.n140 4.5005
R7149 CSoutput.n283 CSoutput.n147 4.5005
R7150 CSoutput.n281 CSoutput.n143 4.5005
R7151 CSoutput.n281 CSoutput.n145 4.5005
R7152 CSoutput.n281 CSoutput.n142 4.5005
R7153 CSoutput.n281 CSoutput.n146 4.5005
R7154 CSoutput.n281 CSoutput.n141 4.5005
R7155 CSoutput.n281 CSoutput.t223 4.5005
R7156 CSoutput.n281 CSoutput.n140 4.5005
R7157 CSoutput.n281 CSoutput.n147 4.5005
R7158 CSoutput.n167 CSoutput.n143 4.5005
R7159 CSoutput.n167 CSoutput.n145 4.5005
R7160 CSoutput.n167 CSoutput.n142 4.5005
R7161 CSoutput.n167 CSoutput.n146 4.5005
R7162 CSoutput.n167 CSoutput.n141 4.5005
R7163 CSoutput.n167 CSoutput.t223 4.5005
R7164 CSoutput.n167 CSoutput.n140 4.5005
R7165 CSoutput.n167 CSoutput.n147 4.5005
R7166 CSoutput.n167 CSoutput.n148 4.5005
R7167 CSoutput.n166 CSoutput.n143 4.5005
R7168 CSoutput.n166 CSoutput.n145 4.5005
R7169 CSoutput.n166 CSoutput.n142 4.5005
R7170 CSoutput.n166 CSoutput.n146 4.5005
R7171 CSoutput.n166 CSoutput.n141 4.5005
R7172 CSoutput.n166 CSoutput.t223 4.5005
R7173 CSoutput.n166 CSoutput.n140 4.5005
R7174 CSoutput.n166 CSoutput.n147 4.5005
R7175 CSoutput.n166 CSoutput.n148 4.5005
R7176 CSoutput.n170 CSoutput.n143 4.5005
R7177 CSoutput.n170 CSoutput.n145 4.5005
R7178 CSoutput.n170 CSoutput.n142 4.5005
R7179 CSoutput.n170 CSoutput.n146 4.5005
R7180 CSoutput.n170 CSoutput.n141 4.5005
R7181 CSoutput.n170 CSoutput.t223 4.5005
R7182 CSoutput.n170 CSoutput.n140 4.5005
R7183 CSoutput.n170 CSoutput.n147 4.5005
R7184 CSoutput.n170 CSoutput.n148 4.5005
R7185 CSoutput.n169 CSoutput.n143 4.5005
R7186 CSoutput.n169 CSoutput.n145 4.5005
R7187 CSoutput.n169 CSoutput.n142 4.5005
R7188 CSoutput.n169 CSoutput.n146 4.5005
R7189 CSoutput.n169 CSoutput.n141 4.5005
R7190 CSoutput.n169 CSoutput.t223 4.5005
R7191 CSoutput.n169 CSoutput.n140 4.5005
R7192 CSoutput.n169 CSoutput.n147 4.5005
R7193 CSoutput.n169 CSoutput.n148 4.5005
R7194 CSoutput.n152 CSoutput.n143 4.5005
R7195 CSoutput.n152 CSoutput.n145 4.5005
R7196 CSoutput.n152 CSoutput.n142 4.5005
R7197 CSoutput.n152 CSoutput.n146 4.5005
R7198 CSoutput.n152 CSoutput.n141 4.5005
R7199 CSoutput.n152 CSoutput.t223 4.5005
R7200 CSoutput.n152 CSoutput.n140 4.5005
R7201 CSoutput.n152 CSoutput.n147 4.5005
R7202 CSoutput.n152 CSoutput.n148 4.5005
R7203 CSoutput.n288 CSoutput.n143 4.5005
R7204 CSoutput.n288 CSoutput.n145 4.5005
R7205 CSoutput.n288 CSoutput.n142 4.5005
R7206 CSoutput.n288 CSoutput.n146 4.5005
R7207 CSoutput.n288 CSoutput.n141 4.5005
R7208 CSoutput.n288 CSoutput.t223 4.5005
R7209 CSoutput.n288 CSoutput.n140 4.5005
R7210 CSoutput.n288 CSoutput.n147 4.5005
R7211 CSoutput.n288 CSoutput.n148 4.5005
R7212 CSoutput.n347 CSoutput.n327 4.10845
R7213 CSoutput.n137 CSoutput.n117 4.10845
R7214 CSoutput.n345 CSoutput.t153 4.06363
R7215 CSoutput.n345 CSoutput.t71 4.06363
R7216 CSoutput.n343 CSoutput.t64 4.06363
R7217 CSoutput.n343 CSoutput.t115 4.06363
R7218 CSoutput.n341 CSoutput.t132 4.06363
R7219 CSoutput.n341 CSoutput.t156 4.06363
R7220 CSoutput.n339 CSoutput.t171 4.06363
R7221 CSoutput.n339 CSoutput.t84 4.06363
R7222 CSoutput.n337 CSoutput.t88 4.06363
R7223 CSoutput.n337 CSoutput.t160 4.06363
R7224 CSoutput.n335 CSoutput.t175 4.06363
R7225 CSoutput.n335 CSoutput.t176 4.06363
R7226 CSoutput.n333 CSoutput.t109 4.06363
R7227 CSoutput.n333 CSoutput.t110 4.06363
R7228 CSoutput.n331 CSoutput.t117 4.06363
R7229 CSoutput.n331 CSoutput.t177 4.06363
R7230 CSoutput.n329 CSoutput.t76 4.06363
R7231 CSoutput.n329 CSoutput.t114 4.06363
R7232 CSoutput.n328 CSoutput.t131 4.06363
R7233 CSoutput.n328 CSoutput.t155 4.06363
R7234 CSoutput.n325 CSoutput.t142 4.06363
R7235 CSoutput.n325 CSoutput.t178 4.06363
R7236 CSoutput.n323 CSoutput.t173 4.06363
R7237 CSoutput.n323 CSoutput.t98 4.06363
R7238 CSoutput.n321 CSoutput.t119 4.06363
R7239 CSoutput.n321 CSoutput.t143 4.06363
R7240 CSoutput.n319 CSoutput.t161 4.06363
R7241 CSoutput.n319 CSoutput.t70 4.06363
R7242 CSoutput.n317 CSoutput.t72 4.06363
R7243 CSoutput.n317 CSoutput.t147 4.06363
R7244 CSoutput.n315 CSoutput.t164 4.06363
R7245 CSoutput.n315 CSoutput.t165 4.06363
R7246 CSoutput.n313 CSoutput.t92 4.06363
R7247 CSoutput.n313 CSoutput.t93 4.06363
R7248 CSoutput.n311 CSoutput.t100 4.06363
R7249 CSoutput.n311 CSoutput.t166 4.06363
R7250 CSoutput.n309 CSoutput.t62 4.06363
R7251 CSoutput.n309 CSoutput.t99 4.06363
R7252 CSoutput.n308 CSoutput.t120 4.06363
R7253 CSoutput.n308 CSoutput.t144 4.06363
R7254 CSoutput.n306 CSoutput.t145 4.06363
R7255 CSoutput.n306 CSoutput.t96 4.06363
R7256 CSoutput.n304 CSoutput.t167 4.06363
R7257 CSoutput.n304 CSoutput.t124 4.06363
R7258 CSoutput.n302 CSoutput.t154 4.06363
R7259 CSoutput.n302 CSoutput.t106 4.06363
R7260 CSoutput.n300 CSoutput.t138 4.06363
R7261 CSoutput.n300 CSoutput.t83 4.06363
R7262 CSoutput.n298 CSoutput.t162 4.06363
R7263 CSoutput.n298 CSoutput.t77 4.06363
R7264 CSoutput.n296 CSoutput.t121 4.06363
R7265 CSoutput.n296 CSoutput.t94 4.06363
R7266 CSoutput.n294 CSoutput.t101 4.06363
R7267 CSoutput.n294 CSoutput.t73 4.06363
R7268 CSoutput.n292 CSoutput.t152 4.06363
R7269 CSoutput.n292 CSoutput.t67 4.06363
R7270 CSoutput.n290 CSoutput.t111 4.06363
R7271 CSoutput.n290 CSoutput.t172 4.06363
R7272 CSoutput.n289 CSoutput.t89 4.06363
R7273 CSoutput.n289 CSoutput.t158 4.06363
R7274 CSoutput.n118 CSoutput.t81 4.06363
R7275 CSoutput.n118 CSoutput.t169 4.06363
R7276 CSoutput.n119 CSoutput.t150 4.06363
R7277 CSoutput.n119 CSoutput.t128 4.06363
R7278 CSoutput.n121 CSoutput.t108 4.06363
R7279 CSoutput.n121 CSoutput.t180 4.06363
R7280 CSoutput.n123 CSoutput.t149 4.06363
R7281 CSoutput.n123 CSoutput.t148 4.06363
R7282 CSoutput.n125 CSoutput.t134 4.06363
R7283 CSoutput.n125 CSoutput.t105 4.06363
R7284 CSoutput.n127 CSoutput.t82 4.06363
R7285 CSoutput.n127 CSoutput.t135 4.06363
R7286 CSoutput.n129 CSoutput.t133 4.06363
R7287 CSoutput.n129 CSoutput.t102 4.06363
R7288 CSoutput.n131 CSoutput.t80 4.06363
R7289 CSoutput.n131 CSoutput.t79 4.06363
R7290 CSoutput.n133 CSoutput.t151 4.06363
R7291 CSoutput.n133 CSoutput.t118 4.06363
R7292 CSoutput.n135 CSoutput.t113 4.06363
R7293 CSoutput.n135 CSoutput.t74 4.06363
R7294 CSoutput.n98 CSoutput.t65 4.06363
R7295 CSoutput.n98 CSoutput.t157 4.06363
R7296 CSoutput.n99 CSoutput.t140 4.06363
R7297 CSoutput.n99 CSoutput.t116 4.06363
R7298 CSoutput.n101 CSoutput.t91 4.06363
R7299 CSoutput.n101 CSoutput.t170 4.06363
R7300 CSoutput.n103 CSoutput.t137 4.06363
R7301 CSoutput.n103 CSoutput.t136 4.06363
R7302 CSoutput.n105 CSoutput.t126 4.06363
R7303 CSoutput.n105 CSoutput.t87 4.06363
R7304 CSoutput.n107 CSoutput.t68 4.06363
R7305 CSoutput.n107 CSoutput.t127 4.06363
R7306 CSoutput.n109 CSoutput.t123 4.06363
R7307 CSoutput.n109 CSoutput.t85 4.06363
R7308 CSoutput.n111 CSoutput.t66 4.06363
R7309 CSoutput.n111 CSoutput.t63 4.06363
R7310 CSoutput.n113 CSoutput.t141 4.06363
R7311 CSoutput.n113 CSoutput.t104 4.06363
R7312 CSoutput.n115 CSoutput.t97 4.06363
R7313 CSoutput.n115 CSoutput.t61 4.06363
R7314 CSoutput.n79 CSoutput.t159 4.06363
R7315 CSoutput.n79 CSoutput.t90 4.06363
R7316 CSoutput.n80 CSoutput.t174 4.06363
R7317 CSoutput.n80 CSoutput.t112 4.06363
R7318 CSoutput.n82 CSoutput.t69 4.06363
R7319 CSoutput.n82 CSoutput.t129 4.06363
R7320 CSoutput.n84 CSoutput.t75 4.06363
R7321 CSoutput.n84 CSoutput.t103 4.06363
R7322 CSoutput.n86 CSoutput.t179 4.06363
R7323 CSoutput.n86 CSoutput.t122 4.06363
R7324 CSoutput.n88 CSoutput.t78 4.06363
R7325 CSoutput.n88 CSoutput.t163 4.06363
R7326 CSoutput.n90 CSoutput.t86 4.06363
R7327 CSoutput.n90 CSoutput.t139 4.06363
R7328 CSoutput.n92 CSoutput.t107 4.06363
R7329 CSoutput.n92 CSoutput.t130 4.06363
R7330 CSoutput.n94 CSoutput.t125 4.06363
R7331 CSoutput.n94 CSoutput.t168 4.06363
R7332 CSoutput.n96 CSoutput.t95 4.06363
R7333 CSoutput.n96 CSoutput.t146 4.06363
R7334 CSoutput.n44 CSoutput.n43 3.79402
R7335 CSoutput.n49 CSoutput.n48 3.79402
R7336 CSoutput.n395 CSoutput.n379 3.72967
R7337 CSoutput.n443 CSoutput.n427 3.72967
R7338 CSoutput.n445 CSoutput.n444 3.57343
R7339 CSoutput.n444 CSoutput.n396 3.08965
R7340 CSoutput.n393 CSoutput.t8 2.82907
R7341 CSoutput.n393 CSoutput.t55 2.82907
R7342 CSoutput.n391 CSoutput.t21 2.82907
R7343 CSoutput.n391 CSoutput.t190 2.82907
R7344 CSoutput.n389 CSoutput.t44 2.82907
R7345 CSoutput.n389 CSoutput.t199 2.82907
R7346 CSoutput.n387 CSoutput.t45 2.82907
R7347 CSoutput.n387 CSoutput.t183 2.82907
R7348 CSoutput.n385 CSoutput.t214 2.82907
R7349 CSoutput.n385 CSoutput.t1 2.82907
R7350 CSoutput.n383 CSoutput.t2 2.82907
R7351 CSoutput.n383 CSoutput.t31 2.82907
R7352 CSoutput.n381 CSoutput.t204 2.82907
R7353 CSoutput.n381 CSoutput.t9 2.82907
R7354 CSoutput.n380 CSoutput.t10 2.82907
R7355 CSoutput.n380 CSoutput.t207 2.82907
R7356 CSoutput.n377 CSoutput.t209 2.82907
R7357 CSoutput.n377 CSoutput.t33 2.82907
R7358 CSoutput.n375 CSoutput.t17 2.82907
R7359 CSoutput.n375 CSoutput.t195 2.82907
R7360 CSoutput.n373 CSoutput.t11 2.82907
R7361 CSoutput.n373 CSoutput.t208 2.82907
R7362 CSoutput.n371 CSoutput.t191 2.82907
R7363 CSoutput.n371 CSoutput.t203 2.82907
R7364 CSoutput.n369 CSoutput.t188 2.82907
R7365 CSoutput.n369 CSoutput.t19 2.82907
R7366 CSoutput.n367 CSoutput.t16 2.82907
R7367 CSoutput.n367 CSoutput.t202 2.82907
R7368 CSoutput.n365 CSoutput.t14 2.82907
R7369 CSoutput.n365 CSoutput.t189 2.82907
R7370 CSoutput.n364 CSoutput.t186 2.82907
R7371 CSoutput.n364 CSoutput.t23 2.82907
R7372 CSoutput.n362 CSoutput.t18 2.82907
R7373 CSoutput.n362 CSoutput.t59 2.82907
R7374 CSoutput.n360 CSoutput.t181 2.82907
R7375 CSoutput.n360 CSoutput.t197 2.82907
R7376 CSoutput.n358 CSoutput.t39 2.82907
R7377 CSoutput.n358 CSoutput.t37 2.82907
R7378 CSoutput.n356 CSoutput.t40 2.82907
R7379 CSoutput.n356 CSoutput.t187 2.82907
R7380 CSoutput.n354 CSoutput.t194 2.82907
R7381 CSoutput.n354 CSoutput.t13 2.82907
R7382 CSoutput.n352 CSoutput.t212 2.82907
R7383 CSoutput.n352 CSoutput.t198 2.82907
R7384 CSoutput.n350 CSoutput.t215 2.82907
R7385 CSoutput.n350 CSoutput.t182 2.82907
R7386 CSoutput.n349 CSoutput.t53 2.82907
R7387 CSoutput.n349 CSoutput.t36 2.82907
R7388 CSoutput.n428 CSoutput.t211 2.82907
R7389 CSoutput.n428 CSoutput.t56 2.82907
R7390 CSoutput.n429 CSoutput.t43 2.82907
R7391 CSoutput.n429 CSoutput.t34 2.82907
R7392 CSoutput.n431 CSoutput.t7 2.82907
R7393 CSoutput.n431 CSoutput.t210 2.82907
R7394 CSoutput.n433 CSoutput.t49 2.82907
R7395 CSoutput.n433 CSoutput.t42 2.82907
R7396 CSoutput.n435 CSoutput.t52 2.82907
R7397 CSoutput.n435 CSoutput.t185 2.82907
R7398 CSoutput.n437 CSoutput.t22 2.82907
R7399 CSoutput.n437 CSoutput.t26 2.82907
R7400 CSoutput.n439 CSoutput.t58 2.82907
R7401 CSoutput.n439 CSoutput.t51 2.82907
R7402 CSoutput.n441 CSoutput.t206 2.82907
R7403 CSoutput.n441 CSoutput.t213 2.82907
R7404 CSoutput.n412 CSoutput.t41 2.82907
R7405 CSoutput.n412 CSoutput.t15 2.82907
R7406 CSoutput.n413 CSoutput.t205 2.82907
R7407 CSoutput.n413 CSoutput.t35 2.82907
R7408 CSoutput.n415 CSoutput.t184 2.82907
R7409 CSoutput.n415 CSoutput.t25 2.82907
R7410 CSoutput.n417 CSoutput.t12 2.82907
R7411 CSoutput.n417 CSoutput.t24 2.82907
R7412 CSoutput.n419 CSoutput.t38 2.82907
R7413 CSoutput.n419 CSoutput.t46 2.82907
R7414 CSoutput.n421 CSoutput.t30 2.82907
R7415 CSoutput.n421 CSoutput.t48 2.82907
R7416 CSoutput.n423 CSoutput.t50 2.82907
R7417 CSoutput.n423 CSoutput.t54 2.82907
R7418 CSoutput.n425 CSoutput.t193 2.82907
R7419 CSoutput.n425 CSoutput.t29 2.82907
R7420 CSoutput.n397 CSoutput.t200 2.82907
R7421 CSoutput.n397 CSoutput.t32 2.82907
R7422 CSoutput.n398 CSoutput.t192 2.82907
R7423 CSoutput.n398 CSoutput.t6 2.82907
R7424 CSoutput.n400 CSoutput.t3 2.82907
R7425 CSoutput.n400 CSoutput.t27 2.82907
R7426 CSoutput.n402 CSoutput.t5 2.82907
R7427 CSoutput.n402 CSoutput.t47 2.82907
R7428 CSoutput.n404 CSoutput.t28 2.82907
R7429 CSoutput.n404 CSoutput.t4 2.82907
R7430 CSoutput.n406 CSoutput.t0 2.82907
R7431 CSoutput.n406 CSoutput.t57 2.82907
R7432 CSoutput.n408 CSoutput.t201 2.82907
R7433 CSoutput.n408 CSoutput.t20 2.82907
R7434 CSoutput.n410 CSoutput.t196 2.82907
R7435 CSoutput.n410 CSoutput.t60 2.82907
R7436 CSoutput.n348 CSoutput.n138 2.78353
R7437 CSoutput.n75 CSoutput.n1 2.45513
R7438 CSoutput.n229 CSoutput.n227 2.251
R7439 CSoutput.n229 CSoutput.n226 2.251
R7440 CSoutput.n229 CSoutput.n225 2.251
R7441 CSoutput.n229 CSoutput.n224 2.251
R7442 CSoutput.n198 CSoutput.n197 2.251
R7443 CSoutput.n198 CSoutput.n196 2.251
R7444 CSoutput.n198 CSoutput.n195 2.251
R7445 CSoutput.n198 CSoutput.n194 2.251
R7446 CSoutput.n271 CSoutput.n270 2.251
R7447 CSoutput.n236 CSoutput.n234 2.251
R7448 CSoutput.n236 CSoutput.n233 2.251
R7449 CSoutput.n236 CSoutput.n232 2.251
R7450 CSoutput.n254 CSoutput.n236 2.251
R7451 CSoutput.n242 CSoutput.n241 2.251
R7452 CSoutput.n242 CSoutput.n240 2.251
R7453 CSoutput.n242 CSoutput.n239 2.251
R7454 CSoutput.n242 CSoutput.n238 2.251
R7455 CSoutput.n268 CSoutput.n208 2.251
R7456 CSoutput.n263 CSoutput.n261 2.251
R7457 CSoutput.n263 CSoutput.n260 2.251
R7458 CSoutput.n263 CSoutput.n259 2.251
R7459 CSoutput.n263 CSoutput.n258 2.251
R7460 CSoutput.n164 CSoutput.n163 2.251
R7461 CSoutput.n164 CSoutput.n162 2.251
R7462 CSoutput.n164 CSoutput.n161 2.251
R7463 CSoutput.n164 CSoutput.n160 2.251
R7464 CSoutput.n281 CSoutput.n280 2.251
R7465 CSoutput.n198 CSoutput.n178 2.2505
R7466 CSoutput.n193 CSoutput.n178 2.2505
R7467 CSoutput.n191 CSoutput.n178 2.2505
R7468 CSoutput.n190 CSoutput.n178 2.2505
R7469 CSoutput.n275 CSoutput.n178 2.2505
R7470 CSoutput.n273 CSoutput.n178 2.2505
R7471 CSoutput.n271 CSoutput.n178 2.2505
R7472 CSoutput.n201 CSoutput.n178 2.2505
R7473 CSoutput.n200 CSoutput.n178 2.2505
R7474 CSoutput.n204 CSoutput.n178 2.2505
R7475 CSoutput.n203 CSoutput.n178 2.2505
R7476 CSoutput.n186 CSoutput.n178 2.2505
R7477 CSoutput.n278 CSoutput.n178 2.2505
R7478 CSoutput.n278 CSoutput.n277 2.2505
R7479 CSoutput.n242 CSoutput.n213 2.2505
R7480 CSoutput.n223 CSoutput.n213 2.2505
R7481 CSoutput.n244 CSoutput.n213 2.2505
R7482 CSoutput.n222 CSoutput.n213 2.2505
R7483 CSoutput.n246 CSoutput.n213 2.2505
R7484 CSoutput.n213 CSoutput.n207 2.2505
R7485 CSoutput.n268 CSoutput.n213 2.2505
R7486 CSoutput.n266 CSoutput.n213 2.2505
R7487 CSoutput.n248 CSoutput.n213 2.2505
R7488 CSoutput.n220 CSoutput.n213 2.2505
R7489 CSoutput.n250 CSoutput.n213 2.2505
R7490 CSoutput.n219 CSoutput.n213 2.2505
R7491 CSoutput.n264 CSoutput.n213 2.2505
R7492 CSoutput.n264 CSoutput.n217 2.2505
R7493 CSoutput.n164 CSoutput.n144 2.2505
R7494 CSoutput.n159 CSoutput.n144 2.2505
R7495 CSoutput.n157 CSoutput.n144 2.2505
R7496 CSoutput.n156 CSoutput.n144 2.2505
R7497 CSoutput.n285 CSoutput.n144 2.2505
R7498 CSoutput.n283 CSoutput.n144 2.2505
R7499 CSoutput.n281 CSoutput.n144 2.2505
R7500 CSoutput.n167 CSoutput.n144 2.2505
R7501 CSoutput.n166 CSoutput.n144 2.2505
R7502 CSoutput.n170 CSoutput.n144 2.2505
R7503 CSoutput.n169 CSoutput.n144 2.2505
R7504 CSoutput.n152 CSoutput.n144 2.2505
R7505 CSoutput.n288 CSoutput.n144 2.2505
R7506 CSoutput.n288 CSoutput.n287 2.2505
R7507 CSoutput.n206 CSoutput.n199 2.25024
R7508 CSoutput.n206 CSoutput.n192 2.25024
R7509 CSoutput.n274 CSoutput.n206 2.25024
R7510 CSoutput.n206 CSoutput.n202 2.25024
R7511 CSoutput.n206 CSoutput.n205 2.25024
R7512 CSoutput.n206 CSoutput.n173 2.25024
R7513 CSoutput.n256 CSoutput.n253 2.25024
R7514 CSoutput.n256 CSoutput.n252 2.25024
R7515 CSoutput.n256 CSoutput.n251 2.25024
R7516 CSoutput.n256 CSoutput.n218 2.25024
R7517 CSoutput.n256 CSoutput.n255 2.25024
R7518 CSoutput.n257 CSoutput.n256 2.25024
R7519 CSoutput.n172 CSoutput.n165 2.25024
R7520 CSoutput.n172 CSoutput.n158 2.25024
R7521 CSoutput.n284 CSoutput.n172 2.25024
R7522 CSoutput.n172 CSoutput.n168 2.25024
R7523 CSoutput.n172 CSoutput.n171 2.25024
R7524 CSoutput.n172 CSoutput.n139 2.25024
R7525 CSoutput.n273 CSoutput.n183 1.50111
R7526 CSoutput.n221 CSoutput.n207 1.50111
R7527 CSoutput.n283 CSoutput.n149 1.50111
R7528 CSoutput.n229 CSoutput.n228 1.501
R7529 CSoutput.n236 CSoutput.n235 1.501
R7530 CSoutput.n263 CSoutput.n262 1.501
R7531 CSoutput.n277 CSoutput.n188 1.12536
R7532 CSoutput.n277 CSoutput.n189 1.12536
R7533 CSoutput.n277 CSoutput.n276 1.12536
R7534 CSoutput.n237 CSoutput.n217 1.12536
R7535 CSoutput.n243 CSoutput.n217 1.12536
R7536 CSoutput.n245 CSoutput.n217 1.12536
R7537 CSoutput.n287 CSoutput.n154 1.12536
R7538 CSoutput.n287 CSoutput.n155 1.12536
R7539 CSoutput.n287 CSoutput.n286 1.12536
R7540 CSoutput.n277 CSoutput.n184 1.12536
R7541 CSoutput.n277 CSoutput.n185 1.12536
R7542 CSoutput.n277 CSoutput.n187 1.12536
R7543 CSoutput.n267 CSoutput.n217 1.12536
R7544 CSoutput.n247 CSoutput.n217 1.12536
R7545 CSoutput.n249 CSoutput.n217 1.12536
R7546 CSoutput.n287 CSoutput.n150 1.12536
R7547 CSoutput.n287 CSoutput.n151 1.12536
R7548 CSoutput.n287 CSoutput.n153 1.12536
R7549 CSoutput.n31 CSoutput.n30 0.669944
R7550 CSoutput.n62 CSoutput.n61 0.669944
R7551 CSoutput.n384 CSoutput.n382 0.573776
R7552 CSoutput.n386 CSoutput.n384 0.573776
R7553 CSoutput.n388 CSoutput.n386 0.573776
R7554 CSoutput.n390 CSoutput.n388 0.573776
R7555 CSoutput.n392 CSoutput.n390 0.573776
R7556 CSoutput.n394 CSoutput.n392 0.573776
R7557 CSoutput.n368 CSoutput.n366 0.573776
R7558 CSoutput.n370 CSoutput.n368 0.573776
R7559 CSoutput.n372 CSoutput.n370 0.573776
R7560 CSoutput.n374 CSoutput.n372 0.573776
R7561 CSoutput.n376 CSoutput.n374 0.573776
R7562 CSoutput.n378 CSoutput.n376 0.573776
R7563 CSoutput.n353 CSoutput.n351 0.573776
R7564 CSoutput.n355 CSoutput.n353 0.573776
R7565 CSoutput.n357 CSoutput.n355 0.573776
R7566 CSoutput.n359 CSoutput.n357 0.573776
R7567 CSoutput.n361 CSoutput.n359 0.573776
R7568 CSoutput.n363 CSoutput.n361 0.573776
R7569 CSoutput.n442 CSoutput.n440 0.573776
R7570 CSoutput.n440 CSoutput.n438 0.573776
R7571 CSoutput.n438 CSoutput.n436 0.573776
R7572 CSoutput.n436 CSoutput.n434 0.573776
R7573 CSoutput.n434 CSoutput.n432 0.573776
R7574 CSoutput.n432 CSoutput.n430 0.573776
R7575 CSoutput.n426 CSoutput.n424 0.573776
R7576 CSoutput.n424 CSoutput.n422 0.573776
R7577 CSoutput.n422 CSoutput.n420 0.573776
R7578 CSoutput.n420 CSoutput.n418 0.573776
R7579 CSoutput.n418 CSoutput.n416 0.573776
R7580 CSoutput.n416 CSoutput.n414 0.573776
R7581 CSoutput.n411 CSoutput.n409 0.573776
R7582 CSoutput.n409 CSoutput.n407 0.573776
R7583 CSoutput.n407 CSoutput.n405 0.573776
R7584 CSoutput.n405 CSoutput.n403 0.573776
R7585 CSoutput.n403 CSoutput.n401 0.573776
R7586 CSoutput.n401 CSoutput.n399 0.573776
R7587 CSoutput.n445 CSoutput.n288 0.53442
R7588 CSoutput.n332 CSoutput.n330 0.358259
R7589 CSoutput.n334 CSoutput.n332 0.358259
R7590 CSoutput.n336 CSoutput.n334 0.358259
R7591 CSoutput.n338 CSoutput.n336 0.358259
R7592 CSoutput.n340 CSoutput.n338 0.358259
R7593 CSoutput.n342 CSoutput.n340 0.358259
R7594 CSoutput.n344 CSoutput.n342 0.358259
R7595 CSoutput.n346 CSoutput.n344 0.358259
R7596 CSoutput.n312 CSoutput.n310 0.358259
R7597 CSoutput.n314 CSoutput.n312 0.358259
R7598 CSoutput.n316 CSoutput.n314 0.358259
R7599 CSoutput.n318 CSoutput.n316 0.358259
R7600 CSoutput.n320 CSoutput.n318 0.358259
R7601 CSoutput.n322 CSoutput.n320 0.358259
R7602 CSoutput.n324 CSoutput.n322 0.358259
R7603 CSoutput.n326 CSoutput.n324 0.358259
R7604 CSoutput.n293 CSoutput.n291 0.358259
R7605 CSoutput.n295 CSoutput.n293 0.358259
R7606 CSoutput.n297 CSoutput.n295 0.358259
R7607 CSoutput.n299 CSoutput.n297 0.358259
R7608 CSoutput.n301 CSoutput.n299 0.358259
R7609 CSoutput.n303 CSoutput.n301 0.358259
R7610 CSoutput.n305 CSoutput.n303 0.358259
R7611 CSoutput.n307 CSoutput.n305 0.358259
R7612 CSoutput.n136 CSoutput.n134 0.358259
R7613 CSoutput.n134 CSoutput.n132 0.358259
R7614 CSoutput.n132 CSoutput.n130 0.358259
R7615 CSoutput.n130 CSoutput.n128 0.358259
R7616 CSoutput.n128 CSoutput.n126 0.358259
R7617 CSoutput.n126 CSoutput.n124 0.358259
R7618 CSoutput.n124 CSoutput.n122 0.358259
R7619 CSoutput.n122 CSoutput.n120 0.358259
R7620 CSoutput.n116 CSoutput.n114 0.358259
R7621 CSoutput.n114 CSoutput.n112 0.358259
R7622 CSoutput.n112 CSoutput.n110 0.358259
R7623 CSoutput.n110 CSoutput.n108 0.358259
R7624 CSoutput.n108 CSoutput.n106 0.358259
R7625 CSoutput.n106 CSoutput.n104 0.358259
R7626 CSoutput.n104 CSoutput.n102 0.358259
R7627 CSoutput.n102 CSoutput.n100 0.358259
R7628 CSoutput.n97 CSoutput.n95 0.358259
R7629 CSoutput.n95 CSoutput.n93 0.358259
R7630 CSoutput.n93 CSoutput.n91 0.358259
R7631 CSoutput.n91 CSoutput.n89 0.358259
R7632 CSoutput.n89 CSoutput.n87 0.358259
R7633 CSoutput.n87 CSoutput.n85 0.358259
R7634 CSoutput.n85 CSoutput.n83 0.358259
R7635 CSoutput.n83 CSoutput.n81 0.358259
R7636 CSoutput.n21 CSoutput.n20 0.169105
R7637 CSoutput.n21 CSoutput.n16 0.169105
R7638 CSoutput.n26 CSoutput.n16 0.169105
R7639 CSoutput.n27 CSoutput.n26 0.169105
R7640 CSoutput.n27 CSoutput.n14 0.169105
R7641 CSoutput.n32 CSoutput.n14 0.169105
R7642 CSoutput.n33 CSoutput.n32 0.169105
R7643 CSoutput.n34 CSoutput.n33 0.169105
R7644 CSoutput.n34 CSoutput.n12 0.169105
R7645 CSoutput.n39 CSoutput.n12 0.169105
R7646 CSoutput.n40 CSoutput.n39 0.169105
R7647 CSoutput.n40 CSoutput.n10 0.169105
R7648 CSoutput.n45 CSoutput.n10 0.169105
R7649 CSoutput.n46 CSoutput.n45 0.169105
R7650 CSoutput.n47 CSoutput.n46 0.169105
R7651 CSoutput.n47 CSoutput.n8 0.169105
R7652 CSoutput.n52 CSoutput.n8 0.169105
R7653 CSoutput.n53 CSoutput.n52 0.169105
R7654 CSoutput.n53 CSoutput.n6 0.169105
R7655 CSoutput.n58 CSoutput.n6 0.169105
R7656 CSoutput.n59 CSoutput.n58 0.169105
R7657 CSoutput.n60 CSoutput.n59 0.169105
R7658 CSoutput.n60 CSoutput.n4 0.169105
R7659 CSoutput.n66 CSoutput.n4 0.169105
R7660 CSoutput.n67 CSoutput.n66 0.169105
R7661 CSoutput.n68 CSoutput.n67 0.169105
R7662 CSoutput.n68 CSoutput.n2 0.169105
R7663 CSoutput.n73 CSoutput.n2 0.169105
R7664 CSoutput.n74 CSoutput.n73 0.169105
R7665 CSoutput.n74 CSoutput.n0 0.169105
R7666 CSoutput.n78 CSoutput.n0 0.169105
R7667 CSoutput.n231 CSoutput.n230 0.0910737
R7668 CSoutput.n282 CSoutput.n279 0.0723685
R7669 CSoutput.n236 CSoutput.n231 0.0522944
R7670 CSoutput.n279 CSoutput.n278 0.0499135
R7671 CSoutput.n230 CSoutput.n229 0.0499135
R7672 CSoutput.n264 CSoutput.n263 0.0464294
R7673 CSoutput.n272 CSoutput.n269 0.0391444
R7674 CSoutput.n231 CSoutput.t226 0.023435
R7675 CSoutput.n279 CSoutput.t218 0.02262
R7676 CSoutput.n230 CSoutput.t220 0.02262
R7677 CSoutput CSoutput.n445 0.0052
R7678 CSoutput.n201 CSoutput.n184 0.00365111
R7679 CSoutput.n204 CSoutput.n185 0.00365111
R7680 CSoutput.n187 CSoutput.n186 0.00365111
R7681 CSoutput.n229 CSoutput.n188 0.00365111
R7682 CSoutput.n193 CSoutput.n189 0.00365111
R7683 CSoutput.n276 CSoutput.n190 0.00365111
R7684 CSoutput.n267 CSoutput.n266 0.00365111
R7685 CSoutput.n247 CSoutput.n220 0.00365111
R7686 CSoutput.n249 CSoutput.n219 0.00365111
R7687 CSoutput.n237 CSoutput.n236 0.00365111
R7688 CSoutput.n243 CSoutput.n223 0.00365111
R7689 CSoutput.n245 CSoutput.n222 0.00365111
R7690 CSoutput.n167 CSoutput.n150 0.00365111
R7691 CSoutput.n170 CSoutput.n151 0.00365111
R7692 CSoutput.n153 CSoutput.n152 0.00365111
R7693 CSoutput.n263 CSoutput.n154 0.00365111
R7694 CSoutput.n159 CSoutput.n155 0.00365111
R7695 CSoutput.n286 CSoutput.n156 0.00365111
R7696 CSoutput.n198 CSoutput.n188 0.00340054
R7697 CSoutput.n191 CSoutput.n189 0.00340054
R7698 CSoutput.n276 CSoutput.n275 0.00340054
R7699 CSoutput.n271 CSoutput.n184 0.00340054
R7700 CSoutput.n200 CSoutput.n185 0.00340054
R7701 CSoutput.n203 CSoutput.n187 0.00340054
R7702 CSoutput.n242 CSoutput.n237 0.00340054
R7703 CSoutput.n244 CSoutput.n243 0.00340054
R7704 CSoutput.n246 CSoutput.n245 0.00340054
R7705 CSoutput.n268 CSoutput.n267 0.00340054
R7706 CSoutput.n248 CSoutput.n247 0.00340054
R7707 CSoutput.n250 CSoutput.n249 0.00340054
R7708 CSoutput.n164 CSoutput.n154 0.00340054
R7709 CSoutput.n157 CSoutput.n155 0.00340054
R7710 CSoutput.n286 CSoutput.n285 0.00340054
R7711 CSoutput.n281 CSoutput.n150 0.00340054
R7712 CSoutput.n166 CSoutput.n151 0.00340054
R7713 CSoutput.n169 CSoutput.n153 0.00340054
R7714 CSoutput.n199 CSoutput.n193 0.00252698
R7715 CSoutput.n192 CSoutput.n190 0.00252698
R7716 CSoutput.n274 CSoutput.n273 0.00252698
R7717 CSoutput.n202 CSoutput.n200 0.00252698
R7718 CSoutput.n205 CSoutput.n203 0.00252698
R7719 CSoutput.n278 CSoutput.n173 0.00252698
R7720 CSoutput.n199 CSoutput.n198 0.00252698
R7721 CSoutput.n192 CSoutput.n191 0.00252698
R7722 CSoutput.n275 CSoutput.n274 0.00252698
R7723 CSoutput.n202 CSoutput.n201 0.00252698
R7724 CSoutput.n205 CSoutput.n204 0.00252698
R7725 CSoutput.n186 CSoutput.n173 0.00252698
R7726 CSoutput.n253 CSoutput.n223 0.00252698
R7727 CSoutput.n252 CSoutput.n222 0.00252698
R7728 CSoutput.n251 CSoutput.n207 0.00252698
R7729 CSoutput.n248 CSoutput.n218 0.00252698
R7730 CSoutput.n255 CSoutput.n250 0.00252698
R7731 CSoutput.n264 CSoutput.n257 0.00252698
R7732 CSoutput.n253 CSoutput.n242 0.00252698
R7733 CSoutput.n252 CSoutput.n244 0.00252698
R7734 CSoutput.n251 CSoutput.n246 0.00252698
R7735 CSoutput.n266 CSoutput.n218 0.00252698
R7736 CSoutput.n255 CSoutput.n220 0.00252698
R7737 CSoutput.n257 CSoutput.n219 0.00252698
R7738 CSoutput.n165 CSoutput.n159 0.00252698
R7739 CSoutput.n158 CSoutput.n156 0.00252698
R7740 CSoutput.n284 CSoutput.n283 0.00252698
R7741 CSoutput.n168 CSoutput.n166 0.00252698
R7742 CSoutput.n171 CSoutput.n169 0.00252698
R7743 CSoutput.n288 CSoutput.n139 0.00252698
R7744 CSoutput.n165 CSoutput.n164 0.00252698
R7745 CSoutput.n158 CSoutput.n157 0.00252698
R7746 CSoutput.n285 CSoutput.n284 0.00252698
R7747 CSoutput.n168 CSoutput.n167 0.00252698
R7748 CSoutput.n171 CSoutput.n170 0.00252698
R7749 CSoutput.n152 CSoutput.n139 0.00252698
R7750 CSoutput.n273 CSoutput.n272 0.0020275
R7751 CSoutput.n272 CSoutput.n271 0.0020275
R7752 CSoutput.n269 CSoutput.n207 0.0020275
R7753 CSoutput.n269 CSoutput.n268 0.0020275
R7754 CSoutput.n283 CSoutput.n282 0.0020275
R7755 CSoutput.n282 CSoutput.n281 0.0020275
R7756 CSoutput.n183 CSoutput.n182 0.00166668
R7757 CSoutput.n265 CSoutput.n221 0.00166668
R7758 CSoutput.n149 CSoutput.n148 0.00166668
R7759 CSoutput.n287 CSoutput.n149 0.00133328
R7760 CSoutput.n221 CSoutput.n217 0.00133328
R7761 CSoutput.n277 CSoutput.n183 0.00133328
R7762 CSoutput.n280 CSoutput.n172 0.001
R7763 CSoutput.n258 CSoutput.n172 0.001
R7764 CSoutput.n160 CSoutput.n140 0.001
R7765 CSoutput.n259 CSoutput.n140 0.001
R7766 CSoutput.n161 CSoutput.n141 0.001
R7767 CSoutput.n260 CSoutput.n141 0.001
R7768 CSoutput.n162 CSoutput.n142 0.001
R7769 CSoutput.n261 CSoutput.n142 0.001
R7770 CSoutput.n163 CSoutput.n143 0.001
R7771 CSoutput.n262 CSoutput.n143 0.001
R7772 CSoutput.n256 CSoutput.n208 0.001
R7773 CSoutput.n256 CSoutput.n254 0.001
R7774 CSoutput.n238 CSoutput.n209 0.001
R7775 CSoutput.n232 CSoutput.n209 0.001
R7776 CSoutput.n239 CSoutput.n210 0.001
R7777 CSoutput.n233 CSoutput.n210 0.001
R7778 CSoutput.n240 CSoutput.n211 0.001
R7779 CSoutput.n234 CSoutput.n211 0.001
R7780 CSoutput.n241 CSoutput.n212 0.001
R7781 CSoutput.n235 CSoutput.n212 0.001
R7782 CSoutput.n270 CSoutput.n206 0.001
R7783 CSoutput.n224 CSoutput.n206 0.001
R7784 CSoutput.n194 CSoutput.n174 0.001
R7785 CSoutput.n225 CSoutput.n174 0.001
R7786 CSoutput.n195 CSoutput.n175 0.001
R7787 CSoutput.n226 CSoutput.n175 0.001
R7788 CSoutput.n196 CSoutput.n176 0.001
R7789 CSoutput.n227 CSoutput.n176 0.001
R7790 CSoutput.n197 CSoutput.n177 0.001
R7791 CSoutput.n228 CSoutput.n177 0.001
R7792 CSoutput.n228 CSoutput.n178 0.001
R7793 CSoutput.n227 CSoutput.n179 0.001
R7794 CSoutput.n226 CSoutput.n180 0.001
R7795 CSoutput.n225 CSoutput.t237 0.001
R7796 CSoutput.n224 CSoutput.n181 0.001
R7797 CSoutput.n197 CSoutput.n179 0.001
R7798 CSoutput.n196 CSoutput.n180 0.001
R7799 CSoutput.n195 CSoutput.t237 0.001
R7800 CSoutput.n194 CSoutput.n181 0.001
R7801 CSoutput.n270 CSoutput.n182 0.001
R7802 CSoutput.n235 CSoutput.n213 0.001
R7803 CSoutput.n234 CSoutput.n214 0.001
R7804 CSoutput.n233 CSoutput.n215 0.001
R7805 CSoutput.n232 CSoutput.t216 0.001
R7806 CSoutput.n254 CSoutput.n216 0.001
R7807 CSoutput.n241 CSoutput.n214 0.001
R7808 CSoutput.n240 CSoutput.n215 0.001
R7809 CSoutput.n239 CSoutput.t216 0.001
R7810 CSoutput.n238 CSoutput.n216 0.001
R7811 CSoutput.n265 CSoutput.n208 0.001
R7812 CSoutput.n262 CSoutput.n144 0.001
R7813 CSoutput.n261 CSoutput.n145 0.001
R7814 CSoutput.n260 CSoutput.n146 0.001
R7815 CSoutput.n259 CSoutput.t223 0.001
R7816 CSoutput.n258 CSoutput.n147 0.001
R7817 CSoutput.n163 CSoutput.n145 0.001
R7818 CSoutput.n162 CSoutput.n146 0.001
R7819 CSoutput.n161 CSoutput.t223 0.001
R7820 CSoutput.n160 CSoutput.n147 0.001
R7821 CSoutput.n280 CSoutput.n148 0.001
R7822 a_n2318_13878.n57 a_n2318_13878.t13 533.335
R7823 a_n2318_13878.n112 a_n2318_13878.t19 512.366
R7824 a_n2318_13878.n64 a_n2318_13878.t9 512.366
R7825 a_n2318_13878.n111 a_n2318_13878.t39 512.366
R7826 a_n2318_13878.n110 a_n2318_13878.t17 512.366
R7827 a_n2318_13878.n65 a_n2318_13878.t11 512.366
R7828 a_n2318_13878.n109 a_n2318_13878.t27 512.366
R7829 a_n2318_13878.n51 a_n2318_13878.t78 533.335
R7830 a_n2318_13878.n108 a_n2318_13878.t59 512.366
R7831 a_n2318_13878.n74 a_n2318_13878.t63 512.366
R7832 a_n2318_13878.n107 a_n2318_13878.t53 512.366
R7833 a_n2318_13878.n106 a_n2318_13878.t68 512.366
R7834 a_n2318_13878.n75 a_n2318_13878.t75 512.366
R7835 a_n2318_13878.n105 a_n2318_13878.t76 512.366
R7836 a_n2318_13878.n36 a_n2318_13878.t15 533.335
R7837 a_n2318_13878.n86 a_n2318_13878.t25 512.366
R7838 a_n2318_13878.n87 a_n2318_13878.t35 512.366
R7839 a_n2318_13878.n88 a_n2318_13878.t37 512.366
R7840 a_n2318_13878.n89 a_n2318_13878.t29 512.366
R7841 a_n2318_13878.n79 a_n2318_13878.t31 512.366
R7842 a_n2318_13878.n90 a_n2318_13878.t33 512.366
R7843 a_n2318_13878.n29 a_n2318_13878.t74 533.335
R7844 a_n2318_13878.n81 a_n2318_13878.t52 512.366
R7845 a_n2318_13878.n82 a_n2318_13878.t71 512.366
R7846 a_n2318_13878.n83 a_n2318_13878.t72 512.366
R7847 a_n2318_13878.n84 a_n2318_13878.t49 512.366
R7848 a_n2318_13878.n80 a_n2318_13878.t58 512.366
R7849 a_n2318_13878.n85 a_n2318_13878.t66 512.366
R7850 a_n2318_13878.n102 a_n2318_13878.t65 512.366
R7851 a_n2318_13878.n92 a_n2318_13878.t56 512.366
R7852 a_n2318_13878.n103 a_n2318_13878.t48 512.366
R7853 a_n2318_13878.n100 a_n2318_13878.t73 512.366
R7854 a_n2318_13878.n93 a_n2318_13878.t62 512.366
R7855 a_n2318_13878.n101 a_n2318_13878.t61 512.366
R7856 a_n2318_13878.n98 a_n2318_13878.t69 512.366
R7857 a_n2318_13878.n94 a_n2318_13878.t54 512.366
R7858 a_n2318_13878.n99 a_n2318_13878.t55 512.366
R7859 a_n2318_13878.n96 a_n2318_13878.t57 512.366
R7860 a_n2318_13878.n95 a_n2318_13878.t67 512.366
R7861 a_n2318_13878.n97 a_n2318_13878.t79 512.366
R7862 a_n2318_13878.n63 a_n2318_13878.n28 70.1674
R7863 a_n2318_13878.n56 a_n2318_13878.n6 70.1674
R7864 a_n2318_13878.n18 a_n2318_13878.n42 70.1674
R7865 a_n2318_13878.n21 a_n2318_13878.n35 70.1674
R7866 a_n2318_13878.n85 a_n2318_13878.n35 20.9683
R7867 a_n2318_13878.n34 a_n2318_13878.n22 72.3034
R7868 a_n2318_13878.n34 a_n2318_13878.n80 16.6962
R7869 a_n2318_13878.n22 a_n2318_13878.n33 77.6622
R7870 a_n2318_13878.n84 a_n2318_13878.n33 5.97853
R7871 a_n2318_13878.n32 a_n2318_13878.n23 77.6622
R7872 a_n2318_13878.n23 a_n2318_13878.n31 72.3034
R7873 a_n2318_13878.n81 a_n2318_13878.n29 20.9683
R7874 a_n2318_13878.n30 a_n2318_13878.n29 70.1674
R7875 a_n2318_13878.n90 a_n2318_13878.n42 20.9683
R7876 a_n2318_13878.n41 a_n2318_13878.n19 72.3034
R7877 a_n2318_13878.n41 a_n2318_13878.n79 16.6962
R7878 a_n2318_13878.n19 a_n2318_13878.n40 77.6622
R7879 a_n2318_13878.n89 a_n2318_13878.n40 5.97853
R7880 a_n2318_13878.n39 a_n2318_13878.n20 77.6622
R7881 a_n2318_13878.n20 a_n2318_13878.n38 72.3034
R7882 a_n2318_13878.n86 a_n2318_13878.n36 20.9683
R7883 a_n2318_13878.n37 a_n2318_13878.n36 70.1674
R7884 a_n2318_13878.n9 a_n2318_13878.n50 70.1674
R7885 a_n2318_13878.n11 a_n2318_13878.n48 70.1674
R7886 a_n2318_13878.n13 a_n2318_13878.n46 70.1674
R7887 a_n2318_13878.n16 a_n2318_13878.n44 70.1674
R7888 a_n2318_13878.n97 a_n2318_13878.n44 20.9683
R7889 a_n2318_13878.n43 a_n2318_13878.n17 75.0448
R7890 a_n2318_13878.n43 a_n2318_13878.n95 11.2134
R7891 a_n2318_13878.n17 a_n2318_13878.n96 161.3
R7892 a_n2318_13878.n99 a_n2318_13878.n46 20.9683
R7893 a_n2318_13878.n45 a_n2318_13878.n14 75.0448
R7894 a_n2318_13878.n45 a_n2318_13878.n94 11.2134
R7895 a_n2318_13878.n14 a_n2318_13878.n98 161.3
R7896 a_n2318_13878.n101 a_n2318_13878.n48 20.9683
R7897 a_n2318_13878.n47 a_n2318_13878.n12 75.0448
R7898 a_n2318_13878.n47 a_n2318_13878.n93 11.2134
R7899 a_n2318_13878.n12 a_n2318_13878.n100 161.3
R7900 a_n2318_13878.n103 a_n2318_13878.n50 20.9683
R7901 a_n2318_13878.n49 a_n2318_13878.n10 75.0448
R7902 a_n2318_13878.n49 a_n2318_13878.n92 11.2134
R7903 a_n2318_13878.n10 a_n2318_13878.n102 161.3
R7904 a_n2318_13878.n105 a_n2318_13878.n56 20.9683
R7905 a_n2318_13878.n7 a_n2318_13878.n55 72.3034
R7906 a_n2318_13878.n55 a_n2318_13878.n75 16.6962
R7907 a_n2318_13878.n54 a_n2318_13878.n7 77.6622
R7908 a_n2318_13878.n106 a_n2318_13878.n54 5.97853
R7909 a_n2318_13878.n53 a_n2318_13878.n5 77.6622
R7910 a_n2318_13878.n5 a_n2318_13878.n52 72.3034
R7911 a_n2318_13878.n108 a_n2318_13878.n51 20.9683
R7912 a_n2318_13878.n8 a_n2318_13878.n51 70.1674
R7913 a_n2318_13878.n109 a_n2318_13878.n63 20.9683
R7914 a_n2318_13878.n28 a_n2318_13878.n62 72.3034
R7915 a_n2318_13878.n62 a_n2318_13878.n65 16.6962
R7916 a_n2318_13878.n61 a_n2318_13878.n60 77.6622
R7917 a_n2318_13878.n110 a_n2318_13878.n61 5.97853
R7918 a_n2318_13878.n59 a_n2318_13878.n4 77.6622
R7919 a_n2318_13878.n4 a_n2318_13878.n58 72.3034
R7920 a_n2318_13878.n112 a_n2318_13878.n57 20.9683
R7921 a_n2318_13878.n3 a_n2318_13878.n57 70.1674
R7922 a_n2318_13878.n1 a_n2318_13878.n72 81.4626
R7923 a_n2318_13878.n2 a_n2318_13878.n68 81.4626
R7924 a_n2318_13878.n2 a_n2318_13878.n66 81.4626
R7925 a_n2318_13878.n1 a_n2318_13878.n73 80.9324
R7926 a_n2318_13878.n1 a_n2318_13878.n71 80.9324
R7927 a_n2318_13878.n0 a_n2318_13878.n70 80.9324
R7928 a_n2318_13878.n2 a_n2318_13878.n69 80.9324
R7929 a_n2318_13878.n2 a_n2318_13878.n67 80.9324
R7930 a_n2318_13878.n26 a_n2318_13878.t22 74.6477
R7931 a_n2318_13878.n24 a_n2318_13878.t16 74.6477
R7932 a_n2318_13878.n27 a_n2318_13878.t14 74.2899
R7933 a_n2318_13878.n25 a_n2318_13878.t24 74.2897
R7934 a_n2318_13878.n26 a_n2318_13878.n114 70.6783
R7935 a_n2318_13878.n26 a_n2318_13878.n115 70.6783
R7936 a_n2318_13878.n25 a_n2318_13878.n78 70.6783
R7937 a_n2318_13878.n24 a_n2318_13878.n77 70.6783
R7938 a_n2318_13878.n24 a_n2318_13878.n76 70.6783
R7939 a_n2318_13878.n116 a_n2318_13878.n27 70.6782
R7940 a_n2318_13878.n111 a_n2318_13878.n110 48.2005
R7941 a_n2318_13878.n63 a_n2318_13878.t21 533.335
R7942 a_n2318_13878.n107 a_n2318_13878.n106 48.2005
R7943 a_n2318_13878.n56 a_n2318_13878.t50 533.335
R7944 a_n2318_13878.n89 a_n2318_13878.n88 48.2005
R7945 a_n2318_13878.t23 a_n2318_13878.n42 533.335
R7946 a_n2318_13878.n84 a_n2318_13878.n83 48.2005
R7947 a_n2318_13878.t51 a_n2318_13878.n35 533.335
R7948 a_n2318_13878.n102 a_n2318_13878.n92 48.2005
R7949 a_n2318_13878.t70 a_n2318_13878.n50 533.335
R7950 a_n2318_13878.n100 a_n2318_13878.n93 48.2005
R7951 a_n2318_13878.t77 a_n2318_13878.n48 533.335
R7952 a_n2318_13878.n98 a_n2318_13878.n94 48.2005
R7953 a_n2318_13878.t64 a_n2318_13878.n46 533.335
R7954 a_n2318_13878.n96 a_n2318_13878.n95 48.2005
R7955 a_n2318_13878.t60 a_n2318_13878.n44 533.335
R7956 a_n2318_13878.n58 a_n2318_13878.n64 16.6962
R7957 a_n2318_13878.n109 a_n2318_13878.n62 27.6507
R7958 a_n2318_13878.n52 a_n2318_13878.n74 16.6962
R7959 a_n2318_13878.n105 a_n2318_13878.n55 27.6507
R7960 a_n2318_13878.n87 a_n2318_13878.n38 16.6962
R7961 a_n2318_13878.n90 a_n2318_13878.n41 27.6507
R7962 a_n2318_13878.n82 a_n2318_13878.n31 16.6962
R7963 a_n2318_13878.n85 a_n2318_13878.n34 27.6507
R7964 a_n2318_13878.n59 a_n2318_13878.n64 41.7634
R7965 a_n2318_13878.n53 a_n2318_13878.n74 41.7634
R7966 a_n2318_13878.n87 a_n2318_13878.n39 41.7634
R7967 a_n2318_13878.n82 a_n2318_13878.n32 41.7634
R7968 a_n2318_13878.n103 a_n2318_13878.n49 35.3134
R7969 a_n2318_13878.n101 a_n2318_13878.n47 35.3134
R7970 a_n2318_13878.n99 a_n2318_13878.n45 35.3134
R7971 a_n2318_13878.n97 a_n2318_13878.n43 35.3134
R7972 a_n2318_13878.n28 a_n2318_13878.n1 23.891
R7973 a_n2318_13878.n30 a_n2318_13878.n15 12.705
R7974 a_n2318_13878.n6 a_n2318_13878.n104 12.5005
R7975 a_n2318_13878.n59 a_n2318_13878.n111 5.97853
R7976 a_n2318_13878.n61 a_n2318_13878.n65 41.7634
R7977 a_n2318_13878.n53 a_n2318_13878.n107 5.97853
R7978 a_n2318_13878.n54 a_n2318_13878.n75 41.7634
R7979 a_n2318_13878.n88 a_n2318_13878.n39 5.97853
R7980 a_n2318_13878.n79 a_n2318_13878.n40 41.7634
R7981 a_n2318_13878.n83 a_n2318_13878.n32 5.97853
R7982 a_n2318_13878.n80 a_n2318_13878.n33 41.7634
R7983 a_n2318_13878.n0 a_n2318_13878.n2 32.5247
R7984 a_n2318_13878.n113 a_n2318_13878.n3 11.1956
R7985 a_n2318_13878.n112 a_n2318_13878.n58 27.6507
R7986 a_n2318_13878.n108 a_n2318_13878.n52 27.6507
R7987 a_n2318_13878.n38 a_n2318_13878.n86 27.6507
R7988 a_n2318_13878.n31 a_n2318_13878.n81 27.6507
R7989 a_n2318_13878.n91 a_n2318_13878.n25 9.85898
R7990 a_n2318_13878.n17 a_n2318_13878.n15 8.73345
R7991 a_n2318_13878.n104 a_n2318_13878.n9 8.73345
R7992 a_n2318_13878.n91 a_n2318_13878.n18 7.36035
R7993 a_n2318_13878.n27 a_n2318_13878.n113 6.01559
R7994 a_n2318_13878.n104 a_n2318_13878.n91 5.3452
R7995 a_n2318_13878.n37 a_n2318_13878.n21 4.01186
R7996 a_n2318_13878.n28 a_n2318_13878.n8 4.0079
R7997 a_n2318_13878.n114 a_n2318_13878.t12 3.61217
R7998 a_n2318_13878.n114 a_n2318_13878.t28 3.61217
R7999 a_n2318_13878.n115 a_n2318_13878.t40 3.61217
R8000 a_n2318_13878.n115 a_n2318_13878.t18 3.61217
R8001 a_n2318_13878.n78 a_n2318_13878.t32 3.61217
R8002 a_n2318_13878.n78 a_n2318_13878.t34 3.61217
R8003 a_n2318_13878.n77 a_n2318_13878.t38 3.61217
R8004 a_n2318_13878.n77 a_n2318_13878.t30 3.61217
R8005 a_n2318_13878.n76 a_n2318_13878.t26 3.61217
R8006 a_n2318_13878.n76 a_n2318_13878.t36 3.61217
R8007 a_n2318_13878.n116 a_n2318_13878.t20 3.61217
R8008 a_n2318_13878.t10 a_n2318_13878.n116 3.61217
R8009 a_n2318_13878.n72 a_n2318_13878.t45 2.82907
R8010 a_n2318_13878.n72 a_n2318_13878.t6 2.82907
R8011 a_n2318_13878.n73 a_n2318_13878.t47 2.82907
R8012 a_n2318_13878.n73 a_n2318_13878.t3 2.82907
R8013 a_n2318_13878.n71 a_n2318_13878.t44 2.82907
R8014 a_n2318_13878.n71 a_n2318_13878.t42 2.82907
R8015 a_n2318_13878.n70 a_n2318_13878.t4 2.82907
R8016 a_n2318_13878.n70 a_n2318_13878.t46 2.82907
R8017 a_n2318_13878.n68 a_n2318_13878.t7 2.82907
R8018 a_n2318_13878.n68 a_n2318_13878.t1 2.82907
R8019 a_n2318_13878.n69 a_n2318_13878.t8 2.82907
R8020 a_n2318_13878.n69 a_n2318_13878.t2 2.82907
R8021 a_n2318_13878.n67 a_n2318_13878.t43 2.82907
R8022 a_n2318_13878.n67 a_n2318_13878.t0 2.82907
R8023 a_n2318_13878.n66 a_n2318_13878.t5 2.82907
R8024 a_n2318_13878.n66 a_n2318_13878.t41 2.82907
R8025 a_n2318_13878.n113 a_n2318_13878.n15 1.30542
R8026 a_n2318_13878.n27 a_n2318_13878.n26 1.07378
R8027 a_n2318_13878.n25 a_n2318_13878.n24 1.07378
R8028 a_n2318_13878.n1 a_n2318_13878.n0 1.06084
R8029 a_n2318_13878.n12 a_n2318_13878.n13 1.04595
R8030 a_n2318_13878.n23 a_n2318_13878.n22 0.758076
R8031 a_n2318_13878.n22 a_n2318_13878.n21 0.758076
R8032 a_n2318_13878.n20 a_n2318_13878.n19 0.758076
R8033 a_n2318_13878.n19 a_n2318_13878.n18 0.758076
R8034 a_n2318_13878.n17 a_n2318_13878.n16 0.758076
R8035 a_n2318_13878.n14 a_n2318_13878.n13 0.758076
R8036 a_n2318_13878.n12 a_n2318_13878.n11 0.758076
R8037 a_n2318_13878.n10 a_n2318_13878.n9 0.758076
R8038 a_n2318_13878.n7 a_n2318_13878.n5 0.758076
R8039 a_n2318_13878.n7 a_n2318_13878.n6 0.758076
R8040 a_n2318_13878.n60 a_n2318_13878.n4 0.758076
R8041 a_n2318_13878.n60 a_n2318_13878.n28 0.724161
R8042 a_n2318_13878.n14 a_n2318_13878.n16 0.67853
R8043 a_n2318_13878.n10 a_n2318_13878.n11 0.67853
R8044 a_n2318_13878.n4 a_n2318_13878.n3 0.568682
R8045 a_n2318_13878.n5 a_n2318_13878.n8 0.568682
R8046 a_n2318_13878.n37 a_n2318_13878.n20 0.568682
R8047 a_n2318_13878.n30 a_n2318_13878.n23 0.568682
R8048 a_n2140_13878.n21 a_n2140_13878.n20 98.9632
R8049 a_n2140_13878.n2 a_n2140_13878.n0 98.7517
R8050 a_n2140_13878.n18 a_n2140_13878.n17 98.6055
R8051 a_n2140_13878.n20 a_n2140_13878.n19 98.6055
R8052 a_n2140_13878.n6 a_n2140_13878.n5 98.6055
R8053 a_n2140_13878.n4 a_n2140_13878.n3 98.6055
R8054 a_n2140_13878.n2 a_n2140_13878.n1 98.6055
R8055 a_n2140_13878.n16 a_n2140_13878.n15 98.6054
R8056 a_n2140_13878.n8 a_n2140_13878.t17 74.6477
R8057 a_n2140_13878.n13 a_n2140_13878.t18 74.2899
R8058 a_n2140_13878.n10 a_n2140_13878.t19 74.2899
R8059 a_n2140_13878.n9 a_n2140_13878.t16 74.2899
R8060 a_n2140_13878.n12 a_n2140_13878.n11 70.6783
R8061 a_n2140_13878.n8 a_n2140_13878.n7 70.6783
R8062 a_n2140_13878.n14 a_n2140_13878.n6 14.2849
R8063 a_n2140_13878.n16 a_n2140_13878.n14 11.9339
R8064 a_n2140_13878.n14 a_n2140_13878.n13 6.95632
R8065 a_n2140_13878.n15 a_n2140_13878.t6 3.61217
R8066 a_n2140_13878.n15 a_n2140_13878.t7 3.61217
R8067 a_n2140_13878.n17 a_n2140_13878.t13 3.61217
R8068 a_n2140_13878.n17 a_n2140_13878.t14 3.61217
R8069 a_n2140_13878.n19 a_n2140_13878.t0 3.61217
R8070 a_n2140_13878.n19 a_n2140_13878.t8 3.61217
R8071 a_n2140_13878.n11 a_n2140_13878.t22 3.61217
R8072 a_n2140_13878.n11 a_n2140_13878.t23 3.61217
R8073 a_n2140_13878.n7 a_n2140_13878.t20 3.61217
R8074 a_n2140_13878.n7 a_n2140_13878.t21 3.61217
R8075 a_n2140_13878.n5 a_n2140_13878.t9 3.61217
R8076 a_n2140_13878.n5 a_n2140_13878.t1 3.61217
R8077 a_n2140_13878.n3 a_n2140_13878.t12 3.61217
R8078 a_n2140_13878.n3 a_n2140_13878.t3 3.61217
R8079 a_n2140_13878.n1 a_n2140_13878.t2 3.61217
R8080 a_n2140_13878.n1 a_n2140_13878.t4 3.61217
R8081 a_n2140_13878.n0 a_n2140_13878.t10 3.61217
R8082 a_n2140_13878.n0 a_n2140_13878.t5 3.61217
R8083 a_n2140_13878.n21 a_n2140_13878.t11 3.61217
R8084 a_n2140_13878.t15 a_n2140_13878.n21 3.61217
R8085 a_n2140_13878.n9 a_n2140_13878.n8 0.358259
R8086 a_n2140_13878.n12 a_n2140_13878.n10 0.358259
R8087 a_n2140_13878.n13 a_n2140_13878.n12 0.358259
R8088 a_n2140_13878.n20 a_n2140_13878.n18 0.358259
R8089 a_n2140_13878.n18 a_n2140_13878.n16 0.358259
R8090 a_n2140_13878.n4 a_n2140_13878.n2 0.146627
R8091 a_n2140_13878.n6 a_n2140_13878.n4 0.146627
R8092 a_n2140_13878.n10 a_n2140_13878.n9 0.101793
R8093 commonsourceibias.n35 commonsourceibias.t12 223.028
R8094 commonsourceibias.n128 commonsourceibias.t129 223.028
R8095 commonsourceibias.n307 commonsourceibias.t140 223.028
R8096 commonsourceibias.n217 commonsourceibias.t112 223.028
R8097 commonsourceibias.n454 commonsourceibias.t30 223.028
R8098 commonsourceibias.n395 commonsourceibias.t108 223.028
R8099 commonsourceibias.n679 commonsourceibias.t74 223.028
R8100 commonsourceibias.n589 commonsourceibias.t97 223.028
R8101 commonsourceibias.n99 commonsourceibias.t34 207.983
R8102 commonsourceibias.n192 commonsourceibias.t120 207.983
R8103 commonsourceibias.n371 commonsourceibias.t147 207.983
R8104 commonsourceibias.n281 commonsourceibias.t71 207.983
R8105 commonsourceibias.n520 commonsourceibias.t6 207.983
R8106 commonsourceibias.n566 commonsourceibias.t91 207.983
R8107 commonsourceibias.n745 commonsourceibias.t82 207.983
R8108 commonsourceibias.n655 commonsourceibias.t151 207.983
R8109 commonsourceibias.n97 commonsourceibias.t42 168.701
R8110 commonsourceibias.n91 commonsourceibias.t60 168.701
R8111 commonsourceibias.n17 commonsourceibias.t32 168.701
R8112 commonsourceibias.n83 commonsourceibias.t22 168.701
R8113 commonsourceibias.n77 commonsourceibias.t0 168.701
R8114 commonsourceibias.n22 commonsourceibias.t18 168.701
R8115 commonsourceibias.n69 commonsourceibias.t62 168.701
R8116 commonsourceibias.n63 commonsourceibias.t36 168.701
R8117 commonsourceibias.n25 commonsourceibias.t48 168.701
R8118 commonsourceibias.n27 commonsourceibias.t14 168.701
R8119 commonsourceibias.n29 commonsourceibias.t20 168.701
R8120 commonsourceibias.n46 commonsourceibias.t50 168.701
R8121 commonsourceibias.n40 commonsourceibias.t2 168.701
R8122 commonsourceibias.n34 commonsourceibias.t52 168.701
R8123 commonsourceibias.n190 commonsourceibias.t67 168.701
R8124 commonsourceibias.n184 commonsourceibias.t126 168.701
R8125 commonsourceibias.n5 commonsourceibias.t121 168.701
R8126 commonsourceibias.n176 commonsourceibias.t136 168.701
R8127 commonsourceibias.n170 commonsourceibias.t117 168.701
R8128 commonsourceibias.n10 commonsourceibias.t102 168.701
R8129 commonsourceibias.n162 commonsourceibias.t125 168.701
R8130 commonsourceibias.n156 commonsourceibias.t118 168.701
R8131 commonsourceibias.n118 commonsourceibias.t76 168.701
R8132 commonsourceibias.n120 commonsourceibias.t106 168.701
R8133 commonsourceibias.n122 commonsourceibias.t96 168.701
R8134 commonsourceibias.n139 commonsourceibias.t141 168.701
R8135 commonsourceibias.n133 commonsourceibias.t116 168.701
R8136 commonsourceibias.n127 commonsourceibias.t152 168.701
R8137 commonsourceibias.n306 commonsourceibias.t130 168.701
R8138 commonsourceibias.n312 commonsourceibias.t79 168.701
R8139 commonsourceibias.n318 commonsourceibias.t149 168.701
R8140 commonsourceibias.n301 commonsourceibias.t133 168.701
R8141 commonsourceibias.n299 commonsourceibias.t137 168.701
R8142 commonsourceibias.n297 commonsourceibias.t64 168.701
R8143 commonsourceibias.n335 commonsourceibias.t138 168.701
R8144 commonsourceibias.n341 commonsourceibias.t146 168.701
R8145 commonsourceibias.n294 commonsourceibias.t119 168.701
R8146 commonsourceibias.n349 commonsourceibias.t90 168.701
R8147 commonsourceibias.n355 commonsourceibias.t155 168.701
R8148 commonsourceibias.n289 commonsourceibias.t124 168.701
R8149 commonsourceibias.n363 commonsourceibias.t128 168.701
R8150 commonsourceibias.n369 commonsourceibias.t75 168.701
R8151 commonsourceibias.n279 commonsourceibias.t159 168.701
R8152 commonsourceibias.n273 commonsourceibias.t148 168.701
R8153 commonsourceibias.n199 commonsourceibias.t78 168.701
R8154 commonsourceibias.n265 commonsourceibias.t157 168.701
R8155 commonsourceibias.n259 commonsourceibias.t85 168.701
R8156 commonsourceibias.n204 commonsourceibias.t77 168.701
R8157 commonsourceibias.n251 commonsourceibias.t158 168.701
R8158 commonsourceibias.n245 commonsourceibias.t94 168.701
R8159 commonsourceibias.n207 commonsourceibias.t113 168.701
R8160 commonsourceibias.n209 commonsourceibias.t156 168.701
R8161 commonsourceibias.n211 commonsourceibias.t92 168.701
R8162 commonsourceibias.n228 commonsourceibias.t111 168.701
R8163 commonsourceibias.n222 commonsourceibias.t105 168.701
R8164 commonsourceibias.n216 commonsourceibias.t93 168.701
R8165 commonsourceibias.n453 commonsourceibias.t26 168.701
R8166 commonsourceibias.n459 commonsourceibias.t44 168.701
R8167 commonsourceibias.n465 commonsourceibias.t58 168.701
R8168 commonsourceibias.n448 commonsourceibias.t54 168.701
R8169 commonsourceibias.n446 commonsourceibias.t46 168.701
R8170 commonsourceibias.n444 commonsourceibias.t38 168.701
R8171 commonsourceibias.n482 commonsourceibias.t8 168.701
R8172 commonsourceibias.n488 commonsourceibias.t16 168.701
R8173 commonsourceibias.n490 commonsourceibias.t40 168.701
R8174 commonsourceibias.n497 commonsourceibias.t10 168.701
R8175 commonsourceibias.n503 commonsourceibias.t56 168.701
R8176 commonsourceibias.n505 commonsourceibias.t4 168.701
R8177 commonsourceibias.n512 commonsourceibias.t28 168.701
R8178 commonsourceibias.n518 commonsourceibias.t24 168.701
R8179 commonsourceibias.n564 commonsourceibias.t134 168.701
R8180 commonsourceibias.n558 commonsourceibias.t114 168.701
R8181 commonsourceibias.n551 commonsourceibias.t95 168.701
R8182 commonsourceibias.n549 commonsourceibias.t123 168.701
R8183 commonsourceibias.n543 commonsourceibias.t88 168.701
R8184 commonsourceibias.n536 commonsourceibias.t73 168.701
R8185 commonsourceibias.n534 commonsourceibias.t104 168.701
R8186 commonsourceibias.n394 commonsourceibias.t131 168.701
R8187 commonsourceibias.n400 commonsourceibias.t84 168.701
R8188 commonsourceibias.n406 commonsourceibias.t127 168.701
R8189 commonsourceibias.n389 commonsourceibias.t150 168.701
R8190 commonsourceibias.n387 commonsourceibias.t83 168.701
R8191 commonsourceibias.n385 commonsourceibias.t139 168.701
R8192 commonsourceibias.n423 commonsourceibias.t89 168.701
R8193 commonsourceibias.n678 commonsourceibias.t145 168.701
R8194 commonsourceibias.n684 commonsourceibias.t109 168.701
R8195 commonsourceibias.n690 commonsourceibias.t87 168.701
R8196 commonsourceibias.n673 commonsourceibias.t153 168.701
R8197 commonsourceibias.n671 commonsourceibias.t132 168.701
R8198 commonsourceibias.n669 commonsourceibias.t103 168.701
R8199 commonsourceibias.n707 commonsourceibias.t70 168.701
R8200 commonsourceibias.n713 commonsourceibias.t81 168.701
R8201 commonsourceibias.n715 commonsourceibias.t110 168.701
R8202 commonsourceibias.n722 commonsourceibias.t115 168.701
R8203 commonsourceibias.n728 commonsourceibias.t101 168.701
R8204 commonsourceibias.n730 commonsourceibias.t135 168.701
R8205 commonsourceibias.n737 commonsourceibias.t122 168.701
R8206 commonsourceibias.n743 commonsourceibias.t107 168.701
R8207 commonsourceibias.n588 commonsourceibias.t68 168.701
R8208 commonsourceibias.n594 commonsourceibias.t86 168.701
R8209 commonsourceibias.n600 commonsourceibias.t98 168.701
R8210 commonsourceibias.n583 commonsourceibias.t69 168.701
R8211 commonsourceibias.n581 commonsourceibias.t80 168.701
R8212 commonsourceibias.n579 commonsourceibias.t99 168.701
R8213 commonsourceibias.n617 commonsourceibias.t72 168.701
R8214 commonsourceibias.n623 commonsourceibias.t142 168.701
R8215 commonsourceibias.n625 commonsourceibias.t100 168.701
R8216 commonsourceibias.n632 commonsourceibias.t65 168.701
R8217 commonsourceibias.n638 commonsourceibias.t143 168.701
R8218 commonsourceibias.n640 commonsourceibias.t154 168.701
R8219 commonsourceibias.n647 commonsourceibias.t66 168.701
R8220 commonsourceibias.n653 commonsourceibias.t144 168.701
R8221 commonsourceibias.n36 commonsourceibias.n33 161.3
R8222 commonsourceibias.n38 commonsourceibias.n37 161.3
R8223 commonsourceibias.n39 commonsourceibias.n32 161.3
R8224 commonsourceibias.n42 commonsourceibias.n41 161.3
R8225 commonsourceibias.n43 commonsourceibias.n31 161.3
R8226 commonsourceibias.n45 commonsourceibias.n44 161.3
R8227 commonsourceibias.n47 commonsourceibias.n30 161.3
R8228 commonsourceibias.n49 commonsourceibias.n48 161.3
R8229 commonsourceibias.n51 commonsourceibias.n50 161.3
R8230 commonsourceibias.n52 commonsourceibias.n28 161.3
R8231 commonsourceibias.n54 commonsourceibias.n53 161.3
R8232 commonsourceibias.n56 commonsourceibias.n55 161.3
R8233 commonsourceibias.n57 commonsourceibias.n26 161.3
R8234 commonsourceibias.n59 commonsourceibias.n58 161.3
R8235 commonsourceibias.n61 commonsourceibias.n60 161.3
R8236 commonsourceibias.n62 commonsourceibias.n24 161.3
R8237 commonsourceibias.n65 commonsourceibias.n64 161.3
R8238 commonsourceibias.n66 commonsourceibias.n23 161.3
R8239 commonsourceibias.n68 commonsourceibias.n67 161.3
R8240 commonsourceibias.n70 commonsourceibias.n21 161.3
R8241 commonsourceibias.n72 commonsourceibias.n71 161.3
R8242 commonsourceibias.n73 commonsourceibias.n20 161.3
R8243 commonsourceibias.n75 commonsourceibias.n74 161.3
R8244 commonsourceibias.n76 commonsourceibias.n19 161.3
R8245 commonsourceibias.n79 commonsourceibias.n78 161.3
R8246 commonsourceibias.n80 commonsourceibias.n18 161.3
R8247 commonsourceibias.n82 commonsourceibias.n81 161.3
R8248 commonsourceibias.n84 commonsourceibias.n16 161.3
R8249 commonsourceibias.n86 commonsourceibias.n85 161.3
R8250 commonsourceibias.n87 commonsourceibias.n15 161.3
R8251 commonsourceibias.n89 commonsourceibias.n88 161.3
R8252 commonsourceibias.n90 commonsourceibias.n14 161.3
R8253 commonsourceibias.n93 commonsourceibias.n92 161.3
R8254 commonsourceibias.n94 commonsourceibias.n13 161.3
R8255 commonsourceibias.n96 commonsourceibias.n95 161.3
R8256 commonsourceibias.n98 commonsourceibias.n12 161.3
R8257 commonsourceibias.n129 commonsourceibias.n126 161.3
R8258 commonsourceibias.n131 commonsourceibias.n130 161.3
R8259 commonsourceibias.n132 commonsourceibias.n125 161.3
R8260 commonsourceibias.n135 commonsourceibias.n134 161.3
R8261 commonsourceibias.n136 commonsourceibias.n124 161.3
R8262 commonsourceibias.n138 commonsourceibias.n137 161.3
R8263 commonsourceibias.n140 commonsourceibias.n123 161.3
R8264 commonsourceibias.n142 commonsourceibias.n141 161.3
R8265 commonsourceibias.n144 commonsourceibias.n143 161.3
R8266 commonsourceibias.n145 commonsourceibias.n121 161.3
R8267 commonsourceibias.n147 commonsourceibias.n146 161.3
R8268 commonsourceibias.n149 commonsourceibias.n148 161.3
R8269 commonsourceibias.n150 commonsourceibias.n119 161.3
R8270 commonsourceibias.n152 commonsourceibias.n151 161.3
R8271 commonsourceibias.n154 commonsourceibias.n153 161.3
R8272 commonsourceibias.n155 commonsourceibias.n117 161.3
R8273 commonsourceibias.n158 commonsourceibias.n157 161.3
R8274 commonsourceibias.n159 commonsourceibias.n11 161.3
R8275 commonsourceibias.n161 commonsourceibias.n160 161.3
R8276 commonsourceibias.n163 commonsourceibias.n9 161.3
R8277 commonsourceibias.n165 commonsourceibias.n164 161.3
R8278 commonsourceibias.n166 commonsourceibias.n8 161.3
R8279 commonsourceibias.n168 commonsourceibias.n167 161.3
R8280 commonsourceibias.n169 commonsourceibias.n7 161.3
R8281 commonsourceibias.n172 commonsourceibias.n171 161.3
R8282 commonsourceibias.n173 commonsourceibias.n6 161.3
R8283 commonsourceibias.n175 commonsourceibias.n174 161.3
R8284 commonsourceibias.n177 commonsourceibias.n4 161.3
R8285 commonsourceibias.n179 commonsourceibias.n178 161.3
R8286 commonsourceibias.n180 commonsourceibias.n3 161.3
R8287 commonsourceibias.n182 commonsourceibias.n181 161.3
R8288 commonsourceibias.n183 commonsourceibias.n2 161.3
R8289 commonsourceibias.n186 commonsourceibias.n185 161.3
R8290 commonsourceibias.n187 commonsourceibias.n1 161.3
R8291 commonsourceibias.n189 commonsourceibias.n188 161.3
R8292 commonsourceibias.n191 commonsourceibias.n0 161.3
R8293 commonsourceibias.n370 commonsourceibias.n284 161.3
R8294 commonsourceibias.n368 commonsourceibias.n367 161.3
R8295 commonsourceibias.n366 commonsourceibias.n285 161.3
R8296 commonsourceibias.n365 commonsourceibias.n364 161.3
R8297 commonsourceibias.n362 commonsourceibias.n286 161.3
R8298 commonsourceibias.n361 commonsourceibias.n360 161.3
R8299 commonsourceibias.n359 commonsourceibias.n287 161.3
R8300 commonsourceibias.n358 commonsourceibias.n357 161.3
R8301 commonsourceibias.n356 commonsourceibias.n288 161.3
R8302 commonsourceibias.n354 commonsourceibias.n353 161.3
R8303 commonsourceibias.n352 commonsourceibias.n290 161.3
R8304 commonsourceibias.n351 commonsourceibias.n350 161.3
R8305 commonsourceibias.n348 commonsourceibias.n291 161.3
R8306 commonsourceibias.n347 commonsourceibias.n346 161.3
R8307 commonsourceibias.n345 commonsourceibias.n292 161.3
R8308 commonsourceibias.n344 commonsourceibias.n343 161.3
R8309 commonsourceibias.n342 commonsourceibias.n293 161.3
R8310 commonsourceibias.n340 commonsourceibias.n339 161.3
R8311 commonsourceibias.n338 commonsourceibias.n295 161.3
R8312 commonsourceibias.n337 commonsourceibias.n336 161.3
R8313 commonsourceibias.n334 commonsourceibias.n296 161.3
R8314 commonsourceibias.n333 commonsourceibias.n332 161.3
R8315 commonsourceibias.n331 commonsourceibias.n330 161.3
R8316 commonsourceibias.n329 commonsourceibias.n298 161.3
R8317 commonsourceibias.n328 commonsourceibias.n327 161.3
R8318 commonsourceibias.n326 commonsourceibias.n325 161.3
R8319 commonsourceibias.n324 commonsourceibias.n300 161.3
R8320 commonsourceibias.n323 commonsourceibias.n322 161.3
R8321 commonsourceibias.n321 commonsourceibias.n320 161.3
R8322 commonsourceibias.n319 commonsourceibias.n302 161.3
R8323 commonsourceibias.n317 commonsourceibias.n316 161.3
R8324 commonsourceibias.n315 commonsourceibias.n303 161.3
R8325 commonsourceibias.n314 commonsourceibias.n313 161.3
R8326 commonsourceibias.n311 commonsourceibias.n304 161.3
R8327 commonsourceibias.n310 commonsourceibias.n309 161.3
R8328 commonsourceibias.n308 commonsourceibias.n305 161.3
R8329 commonsourceibias.n218 commonsourceibias.n215 161.3
R8330 commonsourceibias.n220 commonsourceibias.n219 161.3
R8331 commonsourceibias.n221 commonsourceibias.n214 161.3
R8332 commonsourceibias.n224 commonsourceibias.n223 161.3
R8333 commonsourceibias.n225 commonsourceibias.n213 161.3
R8334 commonsourceibias.n227 commonsourceibias.n226 161.3
R8335 commonsourceibias.n229 commonsourceibias.n212 161.3
R8336 commonsourceibias.n231 commonsourceibias.n230 161.3
R8337 commonsourceibias.n233 commonsourceibias.n232 161.3
R8338 commonsourceibias.n234 commonsourceibias.n210 161.3
R8339 commonsourceibias.n236 commonsourceibias.n235 161.3
R8340 commonsourceibias.n238 commonsourceibias.n237 161.3
R8341 commonsourceibias.n239 commonsourceibias.n208 161.3
R8342 commonsourceibias.n241 commonsourceibias.n240 161.3
R8343 commonsourceibias.n243 commonsourceibias.n242 161.3
R8344 commonsourceibias.n244 commonsourceibias.n206 161.3
R8345 commonsourceibias.n247 commonsourceibias.n246 161.3
R8346 commonsourceibias.n248 commonsourceibias.n205 161.3
R8347 commonsourceibias.n250 commonsourceibias.n249 161.3
R8348 commonsourceibias.n252 commonsourceibias.n203 161.3
R8349 commonsourceibias.n254 commonsourceibias.n253 161.3
R8350 commonsourceibias.n255 commonsourceibias.n202 161.3
R8351 commonsourceibias.n257 commonsourceibias.n256 161.3
R8352 commonsourceibias.n258 commonsourceibias.n201 161.3
R8353 commonsourceibias.n261 commonsourceibias.n260 161.3
R8354 commonsourceibias.n262 commonsourceibias.n200 161.3
R8355 commonsourceibias.n264 commonsourceibias.n263 161.3
R8356 commonsourceibias.n266 commonsourceibias.n198 161.3
R8357 commonsourceibias.n268 commonsourceibias.n267 161.3
R8358 commonsourceibias.n269 commonsourceibias.n197 161.3
R8359 commonsourceibias.n271 commonsourceibias.n270 161.3
R8360 commonsourceibias.n272 commonsourceibias.n196 161.3
R8361 commonsourceibias.n275 commonsourceibias.n274 161.3
R8362 commonsourceibias.n276 commonsourceibias.n195 161.3
R8363 commonsourceibias.n278 commonsourceibias.n277 161.3
R8364 commonsourceibias.n280 commonsourceibias.n194 161.3
R8365 commonsourceibias.n519 commonsourceibias.n433 161.3
R8366 commonsourceibias.n517 commonsourceibias.n516 161.3
R8367 commonsourceibias.n515 commonsourceibias.n434 161.3
R8368 commonsourceibias.n514 commonsourceibias.n513 161.3
R8369 commonsourceibias.n511 commonsourceibias.n435 161.3
R8370 commonsourceibias.n510 commonsourceibias.n509 161.3
R8371 commonsourceibias.n508 commonsourceibias.n436 161.3
R8372 commonsourceibias.n507 commonsourceibias.n506 161.3
R8373 commonsourceibias.n504 commonsourceibias.n437 161.3
R8374 commonsourceibias.n502 commonsourceibias.n501 161.3
R8375 commonsourceibias.n500 commonsourceibias.n438 161.3
R8376 commonsourceibias.n499 commonsourceibias.n498 161.3
R8377 commonsourceibias.n496 commonsourceibias.n439 161.3
R8378 commonsourceibias.n495 commonsourceibias.n494 161.3
R8379 commonsourceibias.n493 commonsourceibias.n440 161.3
R8380 commonsourceibias.n492 commonsourceibias.n491 161.3
R8381 commonsourceibias.n489 commonsourceibias.n441 161.3
R8382 commonsourceibias.n487 commonsourceibias.n486 161.3
R8383 commonsourceibias.n485 commonsourceibias.n442 161.3
R8384 commonsourceibias.n484 commonsourceibias.n483 161.3
R8385 commonsourceibias.n481 commonsourceibias.n443 161.3
R8386 commonsourceibias.n480 commonsourceibias.n479 161.3
R8387 commonsourceibias.n478 commonsourceibias.n477 161.3
R8388 commonsourceibias.n476 commonsourceibias.n445 161.3
R8389 commonsourceibias.n475 commonsourceibias.n474 161.3
R8390 commonsourceibias.n473 commonsourceibias.n472 161.3
R8391 commonsourceibias.n471 commonsourceibias.n447 161.3
R8392 commonsourceibias.n470 commonsourceibias.n469 161.3
R8393 commonsourceibias.n468 commonsourceibias.n467 161.3
R8394 commonsourceibias.n466 commonsourceibias.n449 161.3
R8395 commonsourceibias.n464 commonsourceibias.n463 161.3
R8396 commonsourceibias.n462 commonsourceibias.n450 161.3
R8397 commonsourceibias.n461 commonsourceibias.n460 161.3
R8398 commonsourceibias.n458 commonsourceibias.n451 161.3
R8399 commonsourceibias.n457 commonsourceibias.n456 161.3
R8400 commonsourceibias.n455 commonsourceibias.n452 161.3
R8401 commonsourceibias.n425 commonsourceibias.n424 161.3
R8402 commonsourceibias.n422 commonsourceibias.n384 161.3
R8403 commonsourceibias.n421 commonsourceibias.n420 161.3
R8404 commonsourceibias.n419 commonsourceibias.n418 161.3
R8405 commonsourceibias.n417 commonsourceibias.n386 161.3
R8406 commonsourceibias.n416 commonsourceibias.n415 161.3
R8407 commonsourceibias.n414 commonsourceibias.n413 161.3
R8408 commonsourceibias.n412 commonsourceibias.n388 161.3
R8409 commonsourceibias.n411 commonsourceibias.n410 161.3
R8410 commonsourceibias.n409 commonsourceibias.n408 161.3
R8411 commonsourceibias.n407 commonsourceibias.n390 161.3
R8412 commonsourceibias.n405 commonsourceibias.n404 161.3
R8413 commonsourceibias.n403 commonsourceibias.n391 161.3
R8414 commonsourceibias.n402 commonsourceibias.n401 161.3
R8415 commonsourceibias.n399 commonsourceibias.n392 161.3
R8416 commonsourceibias.n398 commonsourceibias.n397 161.3
R8417 commonsourceibias.n396 commonsourceibias.n393 161.3
R8418 commonsourceibias.n531 commonsourceibias.n383 161.3
R8419 commonsourceibias.n565 commonsourceibias.n374 161.3
R8420 commonsourceibias.n563 commonsourceibias.n562 161.3
R8421 commonsourceibias.n561 commonsourceibias.n375 161.3
R8422 commonsourceibias.n560 commonsourceibias.n559 161.3
R8423 commonsourceibias.n557 commonsourceibias.n376 161.3
R8424 commonsourceibias.n556 commonsourceibias.n555 161.3
R8425 commonsourceibias.n554 commonsourceibias.n377 161.3
R8426 commonsourceibias.n553 commonsourceibias.n552 161.3
R8427 commonsourceibias.n550 commonsourceibias.n378 161.3
R8428 commonsourceibias.n548 commonsourceibias.n547 161.3
R8429 commonsourceibias.n546 commonsourceibias.n379 161.3
R8430 commonsourceibias.n545 commonsourceibias.n544 161.3
R8431 commonsourceibias.n542 commonsourceibias.n380 161.3
R8432 commonsourceibias.n541 commonsourceibias.n540 161.3
R8433 commonsourceibias.n539 commonsourceibias.n381 161.3
R8434 commonsourceibias.n538 commonsourceibias.n537 161.3
R8435 commonsourceibias.n535 commonsourceibias.n382 161.3
R8436 commonsourceibias.n533 commonsourceibias.n532 161.3
R8437 commonsourceibias.n744 commonsourceibias.n658 161.3
R8438 commonsourceibias.n742 commonsourceibias.n741 161.3
R8439 commonsourceibias.n740 commonsourceibias.n659 161.3
R8440 commonsourceibias.n739 commonsourceibias.n738 161.3
R8441 commonsourceibias.n736 commonsourceibias.n660 161.3
R8442 commonsourceibias.n735 commonsourceibias.n734 161.3
R8443 commonsourceibias.n733 commonsourceibias.n661 161.3
R8444 commonsourceibias.n732 commonsourceibias.n731 161.3
R8445 commonsourceibias.n729 commonsourceibias.n662 161.3
R8446 commonsourceibias.n727 commonsourceibias.n726 161.3
R8447 commonsourceibias.n725 commonsourceibias.n663 161.3
R8448 commonsourceibias.n724 commonsourceibias.n723 161.3
R8449 commonsourceibias.n721 commonsourceibias.n664 161.3
R8450 commonsourceibias.n720 commonsourceibias.n719 161.3
R8451 commonsourceibias.n718 commonsourceibias.n665 161.3
R8452 commonsourceibias.n717 commonsourceibias.n716 161.3
R8453 commonsourceibias.n714 commonsourceibias.n666 161.3
R8454 commonsourceibias.n712 commonsourceibias.n711 161.3
R8455 commonsourceibias.n710 commonsourceibias.n667 161.3
R8456 commonsourceibias.n709 commonsourceibias.n708 161.3
R8457 commonsourceibias.n706 commonsourceibias.n668 161.3
R8458 commonsourceibias.n705 commonsourceibias.n704 161.3
R8459 commonsourceibias.n703 commonsourceibias.n702 161.3
R8460 commonsourceibias.n701 commonsourceibias.n670 161.3
R8461 commonsourceibias.n700 commonsourceibias.n699 161.3
R8462 commonsourceibias.n698 commonsourceibias.n697 161.3
R8463 commonsourceibias.n696 commonsourceibias.n672 161.3
R8464 commonsourceibias.n695 commonsourceibias.n694 161.3
R8465 commonsourceibias.n693 commonsourceibias.n692 161.3
R8466 commonsourceibias.n691 commonsourceibias.n674 161.3
R8467 commonsourceibias.n689 commonsourceibias.n688 161.3
R8468 commonsourceibias.n687 commonsourceibias.n675 161.3
R8469 commonsourceibias.n686 commonsourceibias.n685 161.3
R8470 commonsourceibias.n683 commonsourceibias.n676 161.3
R8471 commonsourceibias.n682 commonsourceibias.n681 161.3
R8472 commonsourceibias.n680 commonsourceibias.n677 161.3
R8473 commonsourceibias.n654 commonsourceibias.n568 161.3
R8474 commonsourceibias.n652 commonsourceibias.n651 161.3
R8475 commonsourceibias.n650 commonsourceibias.n569 161.3
R8476 commonsourceibias.n649 commonsourceibias.n648 161.3
R8477 commonsourceibias.n646 commonsourceibias.n570 161.3
R8478 commonsourceibias.n645 commonsourceibias.n644 161.3
R8479 commonsourceibias.n643 commonsourceibias.n571 161.3
R8480 commonsourceibias.n642 commonsourceibias.n641 161.3
R8481 commonsourceibias.n639 commonsourceibias.n572 161.3
R8482 commonsourceibias.n637 commonsourceibias.n636 161.3
R8483 commonsourceibias.n635 commonsourceibias.n573 161.3
R8484 commonsourceibias.n634 commonsourceibias.n633 161.3
R8485 commonsourceibias.n631 commonsourceibias.n574 161.3
R8486 commonsourceibias.n630 commonsourceibias.n629 161.3
R8487 commonsourceibias.n628 commonsourceibias.n575 161.3
R8488 commonsourceibias.n627 commonsourceibias.n626 161.3
R8489 commonsourceibias.n624 commonsourceibias.n576 161.3
R8490 commonsourceibias.n622 commonsourceibias.n621 161.3
R8491 commonsourceibias.n620 commonsourceibias.n577 161.3
R8492 commonsourceibias.n619 commonsourceibias.n618 161.3
R8493 commonsourceibias.n616 commonsourceibias.n578 161.3
R8494 commonsourceibias.n615 commonsourceibias.n614 161.3
R8495 commonsourceibias.n613 commonsourceibias.n612 161.3
R8496 commonsourceibias.n611 commonsourceibias.n580 161.3
R8497 commonsourceibias.n610 commonsourceibias.n609 161.3
R8498 commonsourceibias.n608 commonsourceibias.n607 161.3
R8499 commonsourceibias.n606 commonsourceibias.n582 161.3
R8500 commonsourceibias.n605 commonsourceibias.n604 161.3
R8501 commonsourceibias.n603 commonsourceibias.n602 161.3
R8502 commonsourceibias.n601 commonsourceibias.n584 161.3
R8503 commonsourceibias.n599 commonsourceibias.n598 161.3
R8504 commonsourceibias.n597 commonsourceibias.n585 161.3
R8505 commonsourceibias.n596 commonsourceibias.n595 161.3
R8506 commonsourceibias.n593 commonsourceibias.n586 161.3
R8507 commonsourceibias.n592 commonsourceibias.n591 161.3
R8508 commonsourceibias.n590 commonsourceibias.n587 161.3
R8509 commonsourceibias.n111 commonsourceibias.n109 81.5057
R8510 commonsourceibias.n428 commonsourceibias.n426 81.5057
R8511 commonsourceibias.n111 commonsourceibias.n110 80.9324
R8512 commonsourceibias.n113 commonsourceibias.n112 80.9324
R8513 commonsourceibias.n115 commonsourceibias.n114 80.9324
R8514 commonsourceibias.n108 commonsourceibias.n107 80.9324
R8515 commonsourceibias.n106 commonsourceibias.n105 80.9324
R8516 commonsourceibias.n104 commonsourceibias.n103 80.9324
R8517 commonsourceibias.n102 commonsourceibias.n101 80.9324
R8518 commonsourceibias.n523 commonsourceibias.n522 80.9324
R8519 commonsourceibias.n525 commonsourceibias.n524 80.9324
R8520 commonsourceibias.n527 commonsourceibias.n526 80.9324
R8521 commonsourceibias.n529 commonsourceibias.n528 80.9324
R8522 commonsourceibias.n432 commonsourceibias.n431 80.9324
R8523 commonsourceibias.n430 commonsourceibias.n429 80.9324
R8524 commonsourceibias.n428 commonsourceibias.n427 80.9324
R8525 commonsourceibias.n100 commonsourceibias.n99 80.6037
R8526 commonsourceibias.n193 commonsourceibias.n192 80.6037
R8527 commonsourceibias.n372 commonsourceibias.n371 80.6037
R8528 commonsourceibias.n282 commonsourceibias.n281 80.6037
R8529 commonsourceibias.n521 commonsourceibias.n520 80.6037
R8530 commonsourceibias.n567 commonsourceibias.n566 80.6037
R8531 commonsourceibias.n746 commonsourceibias.n745 80.6037
R8532 commonsourceibias.n656 commonsourceibias.n655 80.6037
R8533 commonsourceibias.n85 commonsourceibias.n84 56.5617
R8534 commonsourceibias.n71 commonsourceibias.n70 56.5617
R8535 commonsourceibias.n62 commonsourceibias.n61 56.5617
R8536 commonsourceibias.n48 commonsourceibias.n47 56.5617
R8537 commonsourceibias.n178 commonsourceibias.n177 56.5617
R8538 commonsourceibias.n164 commonsourceibias.n163 56.5617
R8539 commonsourceibias.n155 commonsourceibias.n154 56.5617
R8540 commonsourceibias.n141 commonsourceibias.n140 56.5617
R8541 commonsourceibias.n320 commonsourceibias.n319 56.5617
R8542 commonsourceibias.n334 commonsourceibias.n333 56.5617
R8543 commonsourceibias.n343 commonsourceibias.n342 56.5617
R8544 commonsourceibias.n357 commonsourceibias.n356 56.5617
R8545 commonsourceibias.n267 commonsourceibias.n266 56.5617
R8546 commonsourceibias.n253 commonsourceibias.n252 56.5617
R8547 commonsourceibias.n244 commonsourceibias.n243 56.5617
R8548 commonsourceibias.n230 commonsourceibias.n229 56.5617
R8549 commonsourceibias.n467 commonsourceibias.n466 56.5617
R8550 commonsourceibias.n481 commonsourceibias.n480 56.5617
R8551 commonsourceibias.n491 commonsourceibias.n489 56.5617
R8552 commonsourceibias.n506 commonsourceibias.n504 56.5617
R8553 commonsourceibias.n552 commonsourceibias.n550 56.5617
R8554 commonsourceibias.n537 commonsourceibias.n535 56.5617
R8555 commonsourceibias.n408 commonsourceibias.n407 56.5617
R8556 commonsourceibias.n422 commonsourceibias.n421 56.5617
R8557 commonsourceibias.n692 commonsourceibias.n691 56.5617
R8558 commonsourceibias.n706 commonsourceibias.n705 56.5617
R8559 commonsourceibias.n716 commonsourceibias.n714 56.5617
R8560 commonsourceibias.n731 commonsourceibias.n729 56.5617
R8561 commonsourceibias.n602 commonsourceibias.n601 56.5617
R8562 commonsourceibias.n616 commonsourceibias.n615 56.5617
R8563 commonsourceibias.n626 commonsourceibias.n624 56.5617
R8564 commonsourceibias.n641 commonsourceibias.n639 56.5617
R8565 commonsourceibias.n76 commonsourceibias.n75 56.0773
R8566 commonsourceibias.n57 commonsourceibias.n56 56.0773
R8567 commonsourceibias.n169 commonsourceibias.n168 56.0773
R8568 commonsourceibias.n150 commonsourceibias.n149 56.0773
R8569 commonsourceibias.n329 commonsourceibias.n328 56.0773
R8570 commonsourceibias.n348 commonsourceibias.n347 56.0773
R8571 commonsourceibias.n258 commonsourceibias.n257 56.0773
R8572 commonsourceibias.n239 commonsourceibias.n238 56.0773
R8573 commonsourceibias.n476 commonsourceibias.n475 56.0773
R8574 commonsourceibias.n496 commonsourceibias.n495 56.0773
R8575 commonsourceibias.n542 commonsourceibias.n541 56.0773
R8576 commonsourceibias.n417 commonsourceibias.n416 56.0773
R8577 commonsourceibias.n701 commonsourceibias.n700 56.0773
R8578 commonsourceibias.n721 commonsourceibias.n720 56.0773
R8579 commonsourceibias.n611 commonsourceibias.n610 56.0773
R8580 commonsourceibias.n631 commonsourceibias.n630 56.0773
R8581 commonsourceibias.n99 commonsourceibias.n98 55.3321
R8582 commonsourceibias.n192 commonsourceibias.n191 55.3321
R8583 commonsourceibias.n371 commonsourceibias.n370 55.3321
R8584 commonsourceibias.n281 commonsourceibias.n280 55.3321
R8585 commonsourceibias.n520 commonsourceibias.n519 55.3321
R8586 commonsourceibias.n566 commonsourceibias.n565 55.3321
R8587 commonsourceibias.n745 commonsourceibias.n744 55.3321
R8588 commonsourceibias.n655 commonsourceibias.n654 55.3321
R8589 commonsourceibias.n90 commonsourceibias.n89 55.1086
R8590 commonsourceibias.n41 commonsourceibias.n31 55.1086
R8591 commonsourceibias.n183 commonsourceibias.n182 55.1086
R8592 commonsourceibias.n134 commonsourceibias.n124 55.1086
R8593 commonsourceibias.n313 commonsourceibias.n303 55.1086
R8594 commonsourceibias.n362 commonsourceibias.n361 55.1086
R8595 commonsourceibias.n272 commonsourceibias.n271 55.1086
R8596 commonsourceibias.n223 commonsourceibias.n213 55.1086
R8597 commonsourceibias.n460 commonsourceibias.n450 55.1086
R8598 commonsourceibias.n511 commonsourceibias.n510 55.1086
R8599 commonsourceibias.n557 commonsourceibias.n556 55.1086
R8600 commonsourceibias.n401 commonsourceibias.n391 55.1086
R8601 commonsourceibias.n685 commonsourceibias.n675 55.1086
R8602 commonsourceibias.n736 commonsourceibias.n735 55.1086
R8603 commonsourceibias.n595 commonsourceibias.n585 55.1086
R8604 commonsourceibias.n646 commonsourceibias.n645 55.1086
R8605 commonsourceibias.n35 commonsourceibias.n34 47.4592
R8606 commonsourceibias.n128 commonsourceibias.n127 47.4592
R8607 commonsourceibias.n307 commonsourceibias.n306 47.4592
R8608 commonsourceibias.n217 commonsourceibias.n216 47.4592
R8609 commonsourceibias.n454 commonsourceibias.n453 47.4592
R8610 commonsourceibias.n395 commonsourceibias.n394 47.4592
R8611 commonsourceibias.n679 commonsourceibias.n678 47.4592
R8612 commonsourceibias.n589 commonsourceibias.n588 47.4592
R8613 commonsourceibias.n308 commonsourceibias.n307 44.0436
R8614 commonsourceibias.n455 commonsourceibias.n454 44.0436
R8615 commonsourceibias.n396 commonsourceibias.n395 44.0436
R8616 commonsourceibias.n680 commonsourceibias.n679 44.0436
R8617 commonsourceibias.n590 commonsourceibias.n589 44.0436
R8618 commonsourceibias.n36 commonsourceibias.n35 44.0436
R8619 commonsourceibias.n129 commonsourceibias.n128 44.0436
R8620 commonsourceibias.n218 commonsourceibias.n217 44.0436
R8621 commonsourceibias.n92 commonsourceibias.n13 42.5146
R8622 commonsourceibias.n39 commonsourceibias.n38 42.5146
R8623 commonsourceibias.n185 commonsourceibias.n1 42.5146
R8624 commonsourceibias.n132 commonsourceibias.n131 42.5146
R8625 commonsourceibias.n311 commonsourceibias.n310 42.5146
R8626 commonsourceibias.n364 commonsourceibias.n285 42.5146
R8627 commonsourceibias.n274 commonsourceibias.n195 42.5146
R8628 commonsourceibias.n221 commonsourceibias.n220 42.5146
R8629 commonsourceibias.n458 commonsourceibias.n457 42.5146
R8630 commonsourceibias.n513 commonsourceibias.n434 42.5146
R8631 commonsourceibias.n559 commonsourceibias.n375 42.5146
R8632 commonsourceibias.n399 commonsourceibias.n398 42.5146
R8633 commonsourceibias.n683 commonsourceibias.n682 42.5146
R8634 commonsourceibias.n738 commonsourceibias.n659 42.5146
R8635 commonsourceibias.n593 commonsourceibias.n592 42.5146
R8636 commonsourceibias.n648 commonsourceibias.n569 42.5146
R8637 commonsourceibias.n78 commonsourceibias.n18 41.5458
R8638 commonsourceibias.n53 commonsourceibias.n52 41.5458
R8639 commonsourceibias.n171 commonsourceibias.n6 41.5458
R8640 commonsourceibias.n146 commonsourceibias.n145 41.5458
R8641 commonsourceibias.n325 commonsourceibias.n324 41.5458
R8642 commonsourceibias.n350 commonsourceibias.n290 41.5458
R8643 commonsourceibias.n260 commonsourceibias.n200 41.5458
R8644 commonsourceibias.n235 commonsourceibias.n234 41.5458
R8645 commonsourceibias.n472 commonsourceibias.n471 41.5458
R8646 commonsourceibias.n498 commonsourceibias.n438 41.5458
R8647 commonsourceibias.n544 commonsourceibias.n379 41.5458
R8648 commonsourceibias.n413 commonsourceibias.n412 41.5458
R8649 commonsourceibias.n697 commonsourceibias.n696 41.5458
R8650 commonsourceibias.n723 commonsourceibias.n663 41.5458
R8651 commonsourceibias.n607 commonsourceibias.n606 41.5458
R8652 commonsourceibias.n633 commonsourceibias.n573 41.5458
R8653 commonsourceibias.n68 commonsourceibias.n23 40.577
R8654 commonsourceibias.n64 commonsourceibias.n23 40.577
R8655 commonsourceibias.n161 commonsourceibias.n11 40.577
R8656 commonsourceibias.n157 commonsourceibias.n11 40.577
R8657 commonsourceibias.n336 commonsourceibias.n295 40.577
R8658 commonsourceibias.n340 commonsourceibias.n295 40.577
R8659 commonsourceibias.n250 commonsourceibias.n205 40.577
R8660 commonsourceibias.n246 commonsourceibias.n205 40.577
R8661 commonsourceibias.n483 commonsourceibias.n442 40.577
R8662 commonsourceibias.n487 commonsourceibias.n442 40.577
R8663 commonsourceibias.n533 commonsourceibias.n383 40.577
R8664 commonsourceibias.n424 commonsourceibias.n383 40.577
R8665 commonsourceibias.n708 commonsourceibias.n667 40.577
R8666 commonsourceibias.n712 commonsourceibias.n667 40.577
R8667 commonsourceibias.n618 commonsourceibias.n577 40.577
R8668 commonsourceibias.n622 commonsourceibias.n577 40.577
R8669 commonsourceibias.n82 commonsourceibias.n18 39.6083
R8670 commonsourceibias.n52 commonsourceibias.n51 39.6083
R8671 commonsourceibias.n175 commonsourceibias.n6 39.6083
R8672 commonsourceibias.n145 commonsourceibias.n144 39.6083
R8673 commonsourceibias.n324 commonsourceibias.n323 39.6083
R8674 commonsourceibias.n354 commonsourceibias.n290 39.6083
R8675 commonsourceibias.n264 commonsourceibias.n200 39.6083
R8676 commonsourceibias.n234 commonsourceibias.n233 39.6083
R8677 commonsourceibias.n471 commonsourceibias.n470 39.6083
R8678 commonsourceibias.n502 commonsourceibias.n438 39.6083
R8679 commonsourceibias.n548 commonsourceibias.n379 39.6083
R8680 commonsourceibias.n412 commonsourceibias.n411 39.6083
R8681 commonsourceibias.n696 commonsourceibias.n695 39.6083
R8682 commonsourceibias.n727 commonsourceibias.n663 39.6083
R8683 commonsourceibias.n606 commonsourceibias.n605 39.6083
R8684 commonsourceibias.n637 commonsourceibias.n573 39.6083
R8685 commonsourceibias.n96 commonsourceibias.n13 38.6395
R8686 commonsourceibias.n38 commonsourceibias.n33 38.6395
R8687 commonsourceibias.n189 commonsourceibias.n1 38.6395
R8688 commonsourceibias.n131 commonsourceibias.n126 38.6395
R8689 commonsourceibias.n310 commonsourceibias.n305 38.6395
R8690 commonsourceibias.n368 commonsourceibias.n285 38.6395
R8691 commonsourceibias.n278 commonsourceibias.n195 38.6395
R8692 commonsourceibias.n220 commonsourceibias.n215 38.6395
R8693 commonsourceibias.n457 commonsourceibias.n452 38.6395
R8694 commonsourceibias.n517 commonsourceibias.n434 38.6395
R8695 commonsourceibias.n563 commonsourceibias.n375 38.6395
R8696 commonsourceibias.n398 commonsourceibias.n393 38.6395
R8697 commonsourceibias.n682 commonsourceibias.n677 38.6395
R8698 commonsourceibias.n742 commonsourceibias.n659 38.6395
R8699 commonsourceibias.n592 commonsourceibias.n587 38.6395
R8700 commonsourceibias.n652 commonsourceibias.n569 38.6395
R8701 commonsourceibias.n89 commonsourceibias.n15 26.0455
R8702 commonsourceibias.n45 commonsourceibias.n31 26.0455
R8703 commonsourceibias.n182 commonsourceibias.n3 26.0455
R8704 commonsourceibias.n138 commonsourceibias.n124 26.0455
R8705 commonsourceibias.n317 commonsourceibias.n303 26.0455
R8706 commonsourceibias.n361 commonsourceibias.n287 26.0455
R8707 commonsourceibias.n271 commonsourceibias.n197 26.0455
R8708 commonsourceibias.n227 commonsourceibias.n213 26.0455
R8709 commonsourceibias.n464 commonsourceibias.n450 26.0455
R8710 commonsourceibias.n510 commonsourceibias.n436 26.0455
R8711 commonsourceibias.n556 commonsourceibias.n377 26.0455
R8712 commonsourceibias.n405 commonsourceibias.n391 26.0455
R8713 commonsourceibias.n689 commonsourceibias.n675 26.0455
R8714 commonsourceibias.n735 commonsourceibias.n661 26.0455
R8715 commonsourceibias.n599 commonsourceibias.n585 26.0455
R8716 commonsourceibias.n645 commonsourceibias.n571 26.0455
R8717 commonsourceibias.n75 commonsourceibias.n20 25.0767
R8718 commonsourceibias.n58 commonsourceibias.n57 25.0767
R8719 commonsourceibias.n168 commonsourceibias.n8 25.0767
R8720 commonsourceibias.n151 commonsourceibias.n150 25.0767
R8721 commonsourceibias.n330 commonsourceibias.n329 25.0767
R8722 commonsourceibias.n347 commonsourceibias.n292 25.0767
R8723 commonsourceibias.n257 commonsourceibias.n202 25.0767
R8724 commonsourceibias.n240 commonsourceibias.n239 25.0767
R8725 commonsourceibias.n477 commonsourceibias.n476 25.0767
R8726 commonsourceibias.n495 commonsourceibias.n440 25.0767
R8727 commonsourceibias.n541 commonsourceibias.n381 25.0767
R8728 commonsourceibias.n418 commonsourceibias.n417 25.0767
R8729 commonsourceibias.n702 commonsourceibias.n701 25.0767
R8730 commonsourceibias.n720 commonsourceibias.n665 25.0767
R8731 commonsourceibias.n612 commonsourceibias.n611 25.0767
R8732 commonsourceibias.n630 commonsourceibias.n575 25.0767
R8733 commonsourceibias.n71 commonsourceibias.n22 24.3464
R8734 commonsourceibias.n61 commonsourceibias.n25 24.3464
R8735 commonsourceibias.n164 commonsourceibias.n10 24.3464
R8736 commonsourceibias.n154 commonsourceibias.n118 24.3464
R8737 commonsourceibias.n333 commonsourceibias.n297 24.3464
R8738 commonsourceibias.n343 commonsourceibias.n294 24.3464
R8739 commonsourceibias.n253 commonsourceibias.n204 24.3464
R8740 commonsourceibias.n243 commonsourceibias.n207 24.3464
R8741 commonsourceibias.n480 commonsourceibias.n444 24.3464
R8742 commonsourceibias.n491 commonsourceibias.n490 24.3464
R8743 commonsourceibias.n537 commonsourceibias.n536 24.3464
R8744 commonsourceibias.n421 commonsourceibias.n385 24.3464
R8745 commonsourceibias.n705 commonsourceibias.n669 24.3464
R8746 commonsourceibias.n716 commonsourceibias.n715 24.3464
R8747 commonsourceibias.n615 commonsourceibias.n579 24.3464
R8748 commonsourceibias.n626 commonsourceibias.n625 24.3464
R8749 commonsourceibias.n85 commonsourceibias.n17 23.8546
R8750 commonsourceibias.n47 commonsourceibias.n46 23.8546
R8751 commonsourceibias.n178 commonsourceibias.n5 23.8546
R8752 commonsourceibias.n140 commonsourceibias.n139 23.8546
R8753 commonsourceibias.n319 commonsourceibias.n318 23.8546
R8754 commonsourceibias.n357 commonsourceibias.n289 23.8546
R8755 commonsourceibias.n267 commonsourceibias.n199 23.8546
R8756 commonsourceibias.n229 commonsourceibias.n228 23.8546
R8757 commonsourceibias.n466 commonsourceibias.n465 23.8546
R8758 commonsourceibias.n506 commonsourceibias.n505 23.8546
R8759 commonsourceibias.n552 commonsourceibias.n551 23.8546
R8760 commonsourceibias.n407 commonsourceibias.n406 23.8546
R8761 commonsourceibias.n691 commonsourceibias.n690 23.8546
R8762 commonsourceibias.n731 commonsourceibias.n730 23.8546
R8763 commonsourceibias.n601 commonsourceibias.n600 23.8546
R8764 commonsourceibias.n641 commonsourceibias.n640 23.8546
R8765 commonsourceibias.n98 commonsourceibias.n97 17.4607
R8766 commonsourceibias.n191 commonsourceibias.n190 17.4607
R8767 commonsourceibias.n370 commonsourceibias.n369 17.4607
R8768 commonsourceibias.n280 commonsourceibias.n279 17.4607
R8769 commonsourceibias.n519 commonsourceibias.n518 17.4607
R8770 commonsourceibias.n565 commonsourceibias.n564 17.4607
R8771 commonsourceibias.n744 commonsourceibias.n743 17.4607
R8772 commonsourceibias.n654 commonsourceibias.n653 17.4607
R8773 commonsourceibias.n84 commonsourceibias.n83 16.9689
R8774 commonsourceibias.n48 commonsourceibias.n29 16.9689
R8775 commonsourceibias.n177 commonsourceibias.n176 16.9689
R8776 commonsourceibias.n141 commonsourceibias.n122 16.9689
R8777 commonsourceibias.n320 commonsourceibias.n301 16.9689
R8778 commonsourceibias.n356 commonsourceibias.n355 16.9689
R8779 commonsourceibias.n266 commonsourceibias.n265 16.9689
R8780 commonsourceibias.n230 commonsourceibias.n211 16.9689
R8781 commonsourceibias.n467 commonsourceibias.n448 16.9689
R8782 commonsourceibias.n504 commonsourceibias.n503 16.9689
R8783 commonsourceibias.n550 commonsourceibias.n549 16.9689
R8784 commonsourceibias.n408 commonsourceibias.n389 16.9689
R8785 commonsourceibias.n692 commonsourceibias.n673 16.9689
R8786 commonsourceibias.n729 commonsourceibias.n728 16.9689
R8787 commonsourceibias.n602 commonsourceibias.n583 16.9689
R8788 commonsourceibias.n639 commonsourceibias.n638 16.9689
R8789 commonsourceibias.n70 commonsourceibias.n69 16.477
R8790 commonsourceibias.n63 commonsourceibias.n62 16.477
R8791 commonsourceibias.n163 commonsourceibias.n162 16.477
R8792 commonsourceibias.n156 commonsourceibias.n155 16.477
R8793 commonsourceibias.n335 commonsourceibias.n334 16.477
R8794 commonsourceibias.n342 commonsourceibias.n341 16.477
R8795 commonsourceibias.n252 commonsourceibias.n251 16.477
R8796 commonsourceibias.n245 commonsourceibias.n244 16.477
R8797 commonsourceibias.n482 commonsourceibias.n481 16.477
R8798 commonsourceibias.n489 commonsourceibias.n488 16.477
R8799 commonsourceibias.n535 commonsourceibias.n534 16.477
R8800 commonsourceibias.n423 commonsourceibias.n422 16.477
R8801 commonsourceibias.n707 commonsourceibias.n706 16.477
R8802 commonsourceibias.n714 commonsourceibias.n713 16.477
R8803 commonsourceibias.n617 commonsourceibias.n616 16.477
R8804 commonsourceibias.n624 commonsourceibias.n623 16.477
R8805 commonsourceibias.n77 commonsourceibias.n76 15.9852
R8806 commonsourceibias.n56 commonsourceibias.n27 15.9852
R8807 commonsourceibias.n170 commonsourceibias.n169 15.9852
R8808 commonsourceibias.n149 commonsourceibias.n120 15.9852
R8809 commonsourceibias.n328 commonsourceibias.n299 15.9852
R8810 commonsourceibias.n349 commonsourceibias.n348 15.9852
R8811 commonsourceibias.n259 commonsourceibias.n258 15.9852
R8812 commonsourceibias.n238 commonsourceibias.n209 15.9852
R8813 commonsourceibias.n475 commonsourceibias.n446 15.9852
R8814 commonsourceibias.n497 commonsourceibias.n496 15.9852
R8815 commonsourceibias.n543 commonsourceibias.n542 15.9852
R8816 commonsourceibias.n416 commonsourceibias.n387 15.9852
R8817 commonsourceibias.n700 commonsourceibias.n671 15.9852
R8818 commonsourceibias.n722 commonsourceibias.n721 15.9852
R8819 commonsourceibias.n610 commonsourceibias.n581 15.9852
R8820 commonsourceibias.n632 commonsourceibias.n631 15.9852
R8821 commonsourceibias.n91 commonsourceibias.n90 15.4934
R8822 commonsourceibias.n41 commonsourceibias.n40 15.4934
R8823 commonsourceibias.n184 commonsourceibias.n183 15.4934
R8824 commonsourceibias.n134 commonsourceibias.n133 15.4934
R8825 commonsourceibias.n313 commonsourceibias.n312 15.4934
R8826 commonsourceibias.n363 commonsourceibias.n362 15.4934
R8827 commonsourceibias.n273 commonsourceibias.n272 15.4934
R8828 commonsourceibias.n223 commonsourceibias.n222 15.4934
R8829 commonsourceibias.n460 commonsourceibias.n459 15.4934
R8830 commonsourceibias.n512 commonsourceibias.n511 15.4934
R8831 commonsourceibias.n558 commonsourceibias.n557 15.4934
R8832 commonsourceibias.n401 commonsourceibias.n400 15.4934
R8833 commonsourceibias.n685 commonsourceibias.n684 15.4934
R8834 commonsourceibias.n737 commonsourceibias.n736 15.4934
R8835 commonsourceibias.n595 commonsourceibias.n594 15.4934
R8836 commonsourceibias.n647 commonsourceibias.n646 15.4934
R8837 commonsourceibias.n102 commonsourceibias.n100 13.2663
R8838 commonsourceibias.n523 commonsourceibias.n521 13.2663
R8839 commonsourceibias.n748 commonsourceibias.n373 10.122
R8840 commonsourceibias.n159 commonsourceibias.n116 9.50363
R8841 commonsourceibias.n531 commonsourceibias.n530 9.50363
R8842 commonsourceibias.n92 commonsourceibias.n91 9.09948
R8843 commonsourceibias.n40 commonsourceibias.n39 9.09948
R8844 commonsourceibias.n185 commonsourceibias.n184 9.09948
R8845 commonsourceibias.n133 commonsourceibias.n132 9.09948
R8846 commonsourceibias.n312 commonsourceibias.n311 9.09948
R8847 commonsourceibias.n364 commonsourceibias.n363 9.09948
R8848 commonsourceibias.n274 commonsourceibias.n273 9.09948
R8849 commonsourceibias.n222 commonsourceibias.n221 9.09948
R8850 commonsourceibias.n459 commonsourceibias.n458 9.09948
R8851 commonsourceibias.n513 commonsourceibias.n512 9.09948
R8852 commonsourceibias.n559 commonsourceibias.n558 9.09948
R8853 commonsourceibias.n400 commonsourceibias.n399 9.09948
R8854 commonsourceibias.n684 commonsourceibias.n683 9.09948
R8855 commonsourceibias.n738 commonsourceibias.n737 9.09948
R8856 commonsourceibias.n594 commonsourceibias.n593 9.09948
R8857 commonsourceibias.n648 commonsourceibias.n647 9.09948
R8858 commonsourceibias.n283 commonsourceibias.n193 8.79451
R8859 commonsourceibias.n657 commonsourceibias.n567 8.79451
R8860 commonsourceibias.n78 commonsourceibias.n77 8.60764
R8861 commonsourceibias.n53 commonsourceibias.n27 8.60764
R8862 commonsourceibias.n171 commonsourceibias.n170 8.60764
R8863 commonsourceibias.n146 commonsourceibias.n120 8.60764
R8864 commonsourceibias.n325 commonsourceibias.n299 8.60764
R8865 commonsourceibias.n350 commonsourceibias.n349 8.60764
R8866 commonsourceibias.n260 commonsourceibias.n259 8.60764
R8867 commonsourceibias.n235 commonsourceibias.n209 8.60764
R8868 commonsourceibias.n472 commonsourceibias.n446 8.60764
R8869 commonsourceibias.n498 commonsourceibias.n497 8.60764
R8870 commonsourceibias.n544 commonsourceibias.n543 8.60764
R8871 commonsourceibias.n413 commonsourceibias.n387 8.60764
R8872 commonsourceibias.n697 commonsourceibias.n671 8.60764
R8873 commonsourceibias.n723 commonsourceibias.n722 8.60764
R8874 commonsourceibias.n607 commonsourceibias.n581 8.60764
R8875 commonsourceibias.n633 commonsourceibias.n632 8.60764
R8876 commonsourceibias.n748 commonsourceibias.n747 8.46921
R8877 commonsourceibias.n69 commonsourceibias.n68 8.11581
R8878 commonsourceibias.n64 commonsourceibias.n63 8.11581
R8879 commonsourceibias.n162 commonsourceibias.n161 8.11581
R8880 commonsourceibias.n157 commonsourceibias.n156 8.11581
R8881 commonsourceibias.n336 commonsourceibias.n335 8.11581
R8882 commonsourceibias.n341 commonsourceibias.n340 8.11581
R8883 commonsourceibias.n251 commonsourceibias.n250 8.11581
R8884 commonsourceibias.n246 commonsourceibias.n245 8.11581
R8885 commonsourceibias.n483 commonsourceibias.n482 8.11581
R8886 commonsourceibias.n488 commonsourceibias.n487 8.11581
R8887 commonsourceibias.n534 commonsourceibias.n533 8.11581
R8888 commonsourceibias.n424 commonsourceibias.n423 8.11581
R8889 commonsourceibias.n708 commonsourceibias.n707 8.11581
R8890 commonsourceibias.n713 commonsourceibias.n712 8.11581
R8891 commonsourceibias.n618 commonsourceibias.n617 8.11581
R8892 commonsourceibias.n623 commonsourceibias.n622 8.11581
R8893 commonsourceibias.n83 commonsourceibias.n82 7.62397
R8894 commonsourceibias.n51 commonsourceibias.n29 7.62397
R8895 commonsourceibias.n176 commonsourceibias.n175 7.62397
R8896 commonsourceibias.n144 commonsourceibias.n122 7.62397
R8897 commonsourceibias.n323 commonsourceibias.n301 7.62397
R8898 commonsourceibias.n355 commonsourceibias.n354 7.62397
R8899 commonsourceibias.n265 commonsourceibias.n264 7.62397
R8900 commonsourceibias.n233 commonsourceibias.n211 7.62397
R8901 commonsourceibias.n470 commonsourceibias.n448 7.62397
R8902 commonsourceibias.n503 commonsourceibias.n502 7.62397
R8903 commonsourceibias.n549 commonsourceibias.n548 7.62397
R8904 commonsourceibias.n411 commonsourceibias.n389 7.62397
R8905 commonsourceibias.n695 commonsourceibias.n673 7.62397
R8906 commonsourceibias.n728 commonsourceibias.n727 7.62397
R8907 commonsourceibias.n605 commonsourceibias.n583 7.62397
R8908 commonsourceibias.n638 commonsourceibias.n637 7.62397
R8909 commonsourceibias.n97 commonsourceibias.n96 7.13213
R8910 commonsourceibias.n34 commonsourceibias.n33 7.13213
R8911 commonsourceibias.n190 commonsourceibias.n189 7.13213
R8912 commonsourceibias.n127 commonsourceibias.n126 7.13213
R8913 commonsourceibias.n306 commonsourceibias.n305 7.13213
R8914 commonsourceibias.n369 commonsourceibias.n368 7.13213
R8915 commonsourceibias.n279 commonsourceibias.n278 7.13213
R8916 commonsourceibias.n216 commonsourceibias.n215 7.13213
R8917 commonsourceibias.n453 commonsourceibias.n452 7.13213
R8918 commonsourceibias.n518 commonsourceibias.n517 7.13213
R8919 commonsourceibias.n564 commonsourceibias.n563 7.13213
R8920 commonsourceibias.n394 commonsourceibias.n393 7.13213
R8921 commonsourceibias.n678 commonsourceibias.n677 7.13213
R8922 commonsourceibias.n743 commonsourceibias.n742 7.13213
R8923 commonsourceibias.n588 commonsourceibias.n587 7.13213
R8924 commonsourceibias.n653 commonsourceibias.n652 7.13213
R8925 commonsourceibias.n373 commonsourceibias.n372 5.06534
R8926 commonsourceibias.n283 commonsourceibias.n282 5.06534
R8927 commonsourceibias.n747 commonsourceibias.n746 5.06534
R8928 commonsourceibias.n657 commonsourceibias.n656 5.06534
R8929 commonsourceibias commonsourceibias.n748 4.04308
R8930 commonsourceibias.n373 commonsourceibias.n283 3.72967
R8931 commonsourceibias.n747 commonsourceibias.n657 3.72967
R8932 commonsourceibias.n109 commonsourceibias.t53 2.82907
R8933 commonsourceibias.n109 commonsourceibias.t13 2.82907
R8934 commonsourceibias.n110 commonsourceibias.t51 2.82907
R8935 commonsourceibias.n110 commonsourceibias.t3 2.82907
R8936 commonsourceibias.n112 commonsourceibias.t15 2.82907
R8937 commonsourceibias.n112 commonsourceibias.t21 2.82907
R8938 commonsourceibias.n114 commonsourceibias.t37 2.82907
R8939 commonsourceibias.n114 commonsourceibias.t49 2.82907
R8940 commonsourceibias.n107 commonsourceibias.t19 2.82907
R8941 commonsourceibias.n107 commonsourceibias.t63 2.82907
R8942 commonsourceibias.n105 commonsourceibias.t23 2.82907
R8943 commonsourceibias.n105 commonsourceibias.t1 2.82907
R8944 commonsourceibias.n103 commonsourceibias.t61 2.82907
R8945 commonsourceibias.n103 commonsourceibias.t33 2.82907
R8946 commonsourceibias.n101 commonsourceibias.t35 2.82907
R8947 commonsourceibias.n101 commonsourceibias.t43 2.82907
R8948 commonsourceibias.n522 commonsourceibias.t25 2.82907
R8949 commonsourceibias.n522 commonsourceibias.t7 2.82907
R8950 commonsourceibias.n524 commonsourceibias.t5 2.82907
R8951 commonsourceibias.n524 commonsourceibias.t29 2.82907
R8952 commonsourceibias.n526 commonsourceibias.t11 2.82907
R8953 commonsourceibias.n526 commonsourceibias.t57 2.82907
R8954 commonsourceibias.n528 commonsourceibias.t17 2.82907
R8955 commonsourceibias.n528 commonsourceibias.t41 2.82907
R8956 commonsourceibias.n431 commonsourceibias.t39 2.82907
R8957 commonsourceibias.n431 commonsourceibias.t9 2.82907
R8958 commonsourceibias.n429 commonsourceibias.t55 2.82907
R8959 commonsourceibias.n429 commonsourceibias.t47 2.82907
R8960 commonsourceibias.n427 commonsourceibias.t45 2.82907
R8961 commonsourceibias.n427 commonsourceibias.t59 2.82907
R8962 commonsourceibias.n426 commonsourceibias.t31 2.82907
R8963 commonsourceibias.n426 commonsourceibias.t27 2.82907
R8964 commonsourceibias.n17 commonsourceibias.n15 0.738255
R8965 commonsourceibias.n46 commonsourceibias.n45 0.738255
R8966 commonsourceibias.n5 commonsourceibias.n3 0.738255
R8967 commonsourceibias.n139 commonsourceibias.n138 0.738255
R8968 commonsourceibias.n318 commonsourceibias.n317 0.738255
R8969 commonsourceibias.n289 commonsourceibias.n287 0.738255
R8970 commonsourceibias.n199 commonsourceibias.n197 0.738255
R8971 commonsourceibias.n228 commonsourceibias.n227 0.738255
R8972 commonsourceibias.n465 commonsourceibias.n464 0.738255
R8973 commonsourceibias.n505 commonsourceibias.n436 0.738255
R8974 commonsourceibias.n551 commonsourceibias.n377 0.738255
R8975 commonsourceibias.n406 commonsourceibias.n405 0.738255
R8976 commonsourceibias.n690 commonsourceibias.n689 0.738255
R8977 commonsourceibias.n730 commonsourceibias.n661 0.738255
R8978 commonsourceibias.n600 commonsourceibias.n599 0.738255
R8979 commonsourceibias.n640 commonsourceibias.n571 0.738255
R8980 commonsourceibias.n104 commonsourceibias.n102 0.573776
R8981 commonsourceibias.n106 commonsourceibias.n104 0.573776
R8982 commonsourceibias.n108 commonsourceibias.n106 0.573776
R8983 commonsourceibias.n115 commonsourceibias.n113 0.573776
R8984 commonsourceibias.n113 commonsourceibias.n111 0.573776
R8985 commonsourceibias.n430 commonsourceibias.n428 0.573776
R8986 commonsourceibias.n432 commonsourceibias.n430 0.573776
R8987 commonsourceibias.n529 commonsourceibias.n527 0.573776
R8988 commonsourceibias.n527 commonsourceibias.n525 0.573776
R8989 commonsourceibias.n525 commonsourceibias.n523 0.573776
R8990 commonsourceibias.n116 commonsourceibias.n108 0.287138
R8991 commonsourceibias.n116 commonsourceibias.n115 0.287138
R8992 commonsourceibias.n530 commonsourceibias.n432 0.287138
R8993 commonsourceibias.n530 commonsourceibias.n529 0.287138
R8994 commonsourceibias.n100 commonsourceibias.n12 0.285035
R8995 commonsourceibias.n193 commonsourceibias.n0 0.285035
R8996 commonsourceibias.n372 commonsourceibias.n284 0.285035
R8997 commonsourceibias.n282 commonsourceibias.n194 0.285035
R8998 commonsourceibias.n521 commonsourceibias.n433 0.285035
R8999 commonsourceibias.n567 commonsourceibias.n374 0.285035
R9000 commonsourceibias.n746 commonsourceibias.n658 0.285035
R9001 commonsourceibias.n656 commonsourceibias.n568 0.285035
R9002 commonsourceibias.n22 commonsourceibias.n20 0.246418
R9003 commonsourceibias.n58 commonsourceibias.n25 0.246418
R9004 commonsourceibias.n10 commonsourceibias.n8 0.246418
R9005 commonsourceibias.n151 commonsourceibias.n118 0.246418
R9006 commonsourceibias.n330 commonsourceibias.n297 0.246418
R9007 commonsourceibias.n294 commonsourceibias.n292 0.246418
R9008 commonsourceibias.n204 commonsourceibias.n202 0.246418
R9009 commonsourceibias.n240 commonsourceibias.n207 0.246418
R9010 commonsourceibias.n477 commonsourceibias.n444 0.246418
R9011 commonsourceibias.n490 commonsourceibias.n440 0.246418
R9012 commonsourceibias.n536 commonsourceibias.n381 0.246418
R9013 commonsourceibias.n418 commonsourceibias.n385 0.246418
R9014 commonsourceibias.n702 commonsourceibias.n669 0.246418
R9015 commonsourceibias.n715 commonsourceibias.n665 0.246418
R9016 commonsourceibias.n612 commonsourceibias.n579 0.246418
R9017 commonsourceibias.n625 commonsourceibias.n575 0.246418
R9018 commonsourceibias.n95 commonsourceibias.n12 0.189894
R9019 commonsourceibias.n95 commonsourceibias.n94 0.189894
R9020 commonsourceibias.n94 commonsourceibias.n93 0.189894
R9021 commonsourceibias.n93 commonsourceibias.n14 0.189894
R9022 commonsourceibias.n88 commonsourceibias.n14 0.189894
R9023 commonsourceibias.n88 commonsourceibias.n87 0.189894
R9024 commonsourceibias.n87 commonsourceibias.n86 0.189894
R9025 commonsourceibias.n86 commonsourceibias.n16 0.189894
R9026 commonsourceibias.n81 commonsourceibias.n16 0.189894
R9027 commonsourceibias.n81 commonsourceibias.n80 0.189894
R9028 commonsourceibias.n80 commonsourceibias.n79 0.189894
R9029 commonsourceibias.n79 commonsourceibias.n19 0.189894
R9030 commonsourceibias.n74 commonsourceibias.n19 0.189894
R9031 commonsourceibias.n74 commonsourceibias.n73 0.189894
R9032 commonsourceibias.n73 commonsourceibias.n72 0.189894
R9033 commonsourceibias.n72 commonsourceibias.n21 0.189894
R9034 commonsourceibias.n67 commonsourceibias.n21 0.189894
R9035 commonsourceibias.n67 commonsourceibias.n66 0.189894
R9036 commonsourceibias.n66 commonsourceibias.n65 0.189894
R9037 commonsourceibias.n65 commonsourceibias.n24 0.189894
R9038 commonsourceibias.n60 commonsourceibias.n24 0.189894
R9039 commonsourceibias.n60 commonsourceibias.n59 0.189894
R9040 commonsourceibias.n59 commonsourceibias.n26 0.189894
R9041 commonsourceibias.n55 commonsourceibias.n26 0.189894
R9042 commonsourceibias.n55 commonsourceibias.n54 0.189894
R9043 commonsourceibias.n54 commonsourceibias.n28 0.189894
R9044 commonsourceibias.n50 commonsourceibias.n28 0.189894
R9045 commonsourceibias.n50 commonsourceibias.n49 0.189894
R9046 commonsourceibias.n49 commonsourceibias.n30 0.189894
R9047 commonsourceibias.n44 commonsourceibias.n30 0.189894
R9048 commonsourceibias.n44 commonsourceibias.n43 0.189894
R9049 commonsourceibias.n43 commonsourceibias.n42 0.189894
R9050 commonsourceibias.n42 commonsourceibias.n32 0.189894
R9051 commonsourceibias.n37 commonsourceibias.n32 0.189894
R9052 commonsourceibias.n37 commonsourceibias.n36 0.189894
R9053 commonsourceibias.n158 commonsourceibias.n117 0.189894
R9054 commonsourceibias.n153 commonsourceibias.n117 0.189894
R9055 commonsourceibias.n153 commonsourceibias.n152 0.189894
R9056 commonsourceibias.n152 commonsourceibias.n119 0.189894
R9057 commonsourceibias.n148 commonsourceibias.n119 0.189894
R9058 commonsourceibias.n148 commonsourceibias.n147 0.189894
R9059 commonsourceibias.n147 commonsourceibias.n121 0.189894
R9060 commonsourceibias.n143 commonsourceibias.n121 0.189894
R9061 commonsourceibias.n143 commonsourceibias.n142 0.189894
R9062 commonsourceibias.n142 commonsourceibias.n123 0.189894
R9063 commonsourceibias.n137 commonsourceibias.n123 0.189894
R9064 commonsourceibias.n137 commonsourceibias.n136 0.189894
R9065 commonsourceibias.n136 commonsourceibias.n135 0.189894
R9066 commonsourceibias.n135 commonsourceibias.n125 0.189894
R9067 commonsourceibias.n130 commonsourceibias.n125 0.189894
R9068 commonsourceibias.n130 commonsourceibias.n129 0.189894
R9069 commonsourceibias.n188 commonsourceibias.n0 0.189894
R9070 commonsourceibias.n188 commonsourceibias.n187 0.189894
R9071 commonsourceibias.n187 commonsourceibias.n186 0.189894
R9072 commonsourceibias.n186 commonsourceibias.n2 0.189894
R9073 commonsourceibias.n181 commonsourceibias.n2 0.189894
R9074 commonsourceibias.n181 commonsourceibias.n180 0.189894
R9075 commonsourceibias.n180 commonsourceibias.n179 0.189894
R9076 commonsourceibias.n179 commonsourceibias.n4 0.189894
R9077 commonsourceibias.n174 commonsourceibias.n4 0.189894
R9078 commonsourceibias.n174 commonsourceibias.n173 0.189894
R9079 commonsourceibias.n173 commonsourceibias.n172 0.189894
R9080 commonsourceibias.n172 commonsourceibias.n7 0.189894
R9081 commonsourceibias.n167 commonsourceibias.n7 0.189894
R9082 commonsourceibias.n167 commonsourceibias.n166 0.189894
R9083 commonsourceibias.n166 commonsourceibias.n165 0.189894
R9084 commonsourceibias.n165 commonsourceibias.n9 0.189894
R9085 commonsourceibias.n160 commonsourceibias.n9 0.189894
R9086 commonsourceibias.n367 commonsourceibias.n284 0.189894
R9087 commonsourceibias.n367 commonsourceibias.n366 0.189894
R9088 commonsourceibias.n366 commonsourceibias.n365 0.189894
R9089 commonsourceibias.n365 commonsourceibias.n286 0.189894
R9090 commonsourceibias.n360 commonsourceibias.n286 0.189894
R9091 commonsourceibias.n360 commonsourceibias.n359 0.189894
R9092 commonsourceibias.n359 commonsourceibias.n358 0.189894
R9093 commonsourceibias.n358 commonsourceibias.n288 0.189894
R9094 commonsourceibias.n353 commonsourceibias.n288 0.189894
R9095 commonsourceibias.n353 commonsourceibias.n352 0.189894
R9096 commonsourceibias.n352 commonsourceibias.n351 0.189894
R9097 commonsourceibias.n351 commonsourceibias.n291 0.189894
R9098 commonsourceibias.n346 commonsourceibias.n291 0.189894
R9099 commonsourceibias.n346 commonsourceibias.n345 0.189894
R9100 commonsourceibias.n345 commonsourceibias.n344 0.189894
R9101 commonsourceibias.n344 commonsourceibias.n293 0.189894
R9102 commonsourceibias.n339 commonsourceibias.n293 0.189894
R9103 commonsourceibias.n339 commonsourceibias.n338 0.189894
R9104 commonsourceibias.n338 commonsourceibias.n337 0.189894
R9105 commonsourceibias.n337 commonsourceibias.n296 0.189894
R9106 commonsourceibias.n332 commonsourceibias.n296 0.189894
R9107 commonsourceibias.n332 commonsourceibias.n331 0.189894
R9108 commonsourceibias.n331 commonsourceibias.n298 0.189894
R9109 commonsourceibias.n327 commonsourceibias.n298 0.189894
R9110 commonsourceibias.n327 commonsourceibias.n326 0.189894
R9111 commonsourceibias.n326 commonsourceibias.n300 0.189894
R9112 commonsourceibias.n322 commonsourceibias.n300 0.189894
R9113 commonsourceibias.n322 commonsourceibias.n321 0.189894
R9114 commonsourceibias.n321 commonsourceibias.n302 0.189894
R9115 commonsourceibias.n316 commonsourceibias.n302 0.189894
R9116 commonsourceibias.n316 commonsourceibias.n315 0.189894
R9117 commonsourceibias.n315 commonsourceibias.n314 0.189894
R9118 commonsourceibias.n314 commonsourceibias.n304 0.189894
R9119 commonsourceibias.n309 commonsourceibias.n304 0.189894
R9120 commonsourceibias.n309 commonsourceibias.n308 0.189894
R9121 commonsourceibias.n277 commonsourceibias.n194 0.189894
R9122 commonsourceibias.n277 commonsourceibias.n276 0.189894
R9123 commonsourceibias.n276 commonsourceibias.n275 0.189894
R9124 commonsourceibias.n275 commonsourceibias.n196 0.189894
R9125 commonsourceibias.n270 commonsourceibias.n196 0.189894
R9126 commonsourceibias.n270 commonsourceibias.n269 0.189894
R9127 commonsourceibias.n269 commonsourceibias.n268 0.189894
R9128 commonsourceibias.n268 commonsourceibias.n198 0.189894
R9129 commonsourceibias.n263 commonsourceibias.n198 0.189894
R9130 commonsourceibias.n263 commonsourceibias.n262 0.189894
R9131 commonsourceibias.n262 commonsourceibias.n261 0.189894
R9132 commonsourceibias.n261 commonsourceibias.n201 0.189894
R9133 commonsourceibias.n256 commonsourceibias.n201 0.189894
R9134 commonsourceibias.n256 commonsourceibias.n255 0.189894
R9135 commonsourceibias.n255 commonsourceibias.n254 0.189894
R9136 commonsourceibias.n254 commonsourceibias.n203 0.189894
R9137 commonsourceibias.n249 commonsourceibias.n203 0.189894
R9138 commonsourceibias.n249 commonsourceibias.n248 0.189894
R9139 commonsourceibias.n248 commonsourceibias.n247 0.189894
R9140 commonsourceibias.n247 commonsourceibias.n206 0.189894
R9141 commonsourceibias.n242 commonsourceibias.n206 0.189894
R9142 commonsourceibias.n242 commonsourceibias.n241 0.189894
R9143 commonsourceibias.n241 commonsourceibias.n208 0.189894
R9144 commonsourceibias.n237 commonsourceibias.n208 0.189894
R9145 commonsourceibias.n237 commonsourceibias.n236 0.189894
R9146 commonsourceibias.n236 commonsourceibias.n210 0.189894
R9147 commonsourceibias.n232 commonsourceibias.n210 0.189894
R9148 commonsourceibias.n232 commonsourceibias.n231 0.189894
R9149 commonsourceibias.n231 commonsourceibias.n212 0.189894
R9150 commonsourceibias.n226 commonsourceibias.n212 0.189894
R9151 commonsourceibias.n226 commonsourceibias.n225 0.189894
R9152 commonsourceibias.n225 commonsourceibias.n224 0.189894
R9153 commonsourceibias.n224 commonsourceibias.n214 0.189894
R9154 commonsourceibias.n219 commonsourceibias.n214 0.189894
R9155 commonsourceibias.n219 commonsourceibias.n218 0.189894
R9156 commonsourceibias.n456 commonsourceibias.n455 0.189894
R9157 commonsourceibias.n456 commonsourceibias.n451 0.189894
R9158 commonsourceibias.n461 commonsourceibias.n451 0.189894
R9159 commonsourceibias.n462 commonsourceibias.n461 0.189894
R9160 commonsourceibias.n463 commonsourceibias.n462 0.189894
R9161 commonsourceibias.n463 commonsourceibias.n449 0.189894
R9162 commonsourceibias.n468 commonsourceibias.n449 0.189894
R9163 commonsourceibias.n469 commonsourceibias.n468 0.189894
R9164 commonsourceibias.n469 commonsourceibias.n447 0.189894
R9165 commonsourceibias.n473 commonsourceibias.n447 0.189894
R9166 commonsourceibias.n474 commonsourceibias.n473 0.189894
R9167 commonsourceibias.n474 commonsourceibias.n445 0.189894
R9168 commonsourceibias.n478 commonsourceibias.n445 0.189894
R9169 commonsourceibias.n479 commonsourceibias.n478 0.189894
R9170 commonsourceibias.n479 commonsourceibias.n443 0.189894
R9171 commonsourceibias.n484 commonsourceibias.n443 0.189894
R9172 commonsourceibias.n485 commonsourceibias.n484 0.189894
R9173 commonsourceibias.n486 commonsourceibias.n485 0.189894
R9174 commonsourceibias.n486 commonsourceibias.n441 0.189894
R9175 commonsourceibias.n492 commonsourceibias.n441 0.189894
R9176 commonsourceibias.n493 commonsourceibias.n492 0.189894
R9177 commonsourceibias.n494 commonsourceibias.n493 0.189894
R9178 commonsourceibias.n494 commonsourceibias.n439 0.189894
R9179 commonsourceibias.n499 commonsourceibias.n439 0.189894
R9180 commonsourceibias.n500 commonsourceibias.n499 0.189894
R9181 commonsourceibias.n501 commonsourceibias.n500 0.189894
R9182 commonsourceibias.n501 commonsourceibias.n437 0.189894
R9183 commonsourceibias.n507 commonsourceibias.n437 0.189894
R9184 commonsourceibias.n508 commonsourceibias.n507 0.189894
R9185 commonsourceibias.n509 commonsourceibias.n508 0.189894
R9186 commonsourceibias.n509 commonsourceibias.n435 0.189894
R9187 commonsourceibias.n514 commonsourceibias.n435 0.189894
R9188 commonsourceibias.n515 commonsourceibias.n514 0.189894
R9189 commonsourceibias.n516 commonsourceibias.n515 0.189894
R9190 commonsourceibias.n516 commonsourceibias.n433 0.189894
R9191 commonsourceibias.n397 commonsourceibias.n396 0.189894
R9192 commonsourceibias.n397 commonsourceibias.n392 0.189894
R9193 commonsourceibias.n402 commonsourceibias.n392 0.189894
R9194 commonsourceibias.n403 commonsourceibias.n402 0.189894
R9195 commonsourceibias.n404 commonsourceibias.n403 0.189894
R9196 commonsourceibias.n404 commonsourceibias.n390 0.189894
R9197 commonsourceibias.n409 commonsourceibias.n390 0.189894
R9198 commonsourceibias.n410 commonsourceibias.n409 0.189894
R9199 commonsourceibias.n410 commonsourceibias.n388 0.189894
R9200 commonsourceibias.n414 commonsourceibias.n388 0.189894
R9201 commonsourceibias.n415 commonsourceibias.n414 0.189894
R9202 commonsourceibias.n415 commonsourceibias.n386 0.189894
R9203 commonsourceibias.n419 commonsourceibias.n386 0.189894
R9204 commonsourceibias.n420 commonsourceibias.n419 0.189894
R9205 commonsourceibias.n420 commonsourceibias.n384 0.189894
R9206 commonsourceibias.n425 commonsourceibias.n384 0.189894
R9207 commonsourceibias.n532 commonsourceibias.n382 0.189894
R9208 commonsourceibias.n538 commonsourceibias.n382 0.189894
R9209 commonsourceibias.n539 commonsourceibias.n538 0.189894
R9210 commonsourceibias.n540 commonsourceibias.n539 0.189894
R9211 commonsourceibias.n540 commonsourceibias.n380 0.189894
R9212 commonsourceibias.n545 commonsourceibias.n380 0.189894
R9213 commonsourceibias.n546 commonsourceibias.n545 0.189894
R9214 commonsourceibias.n547 commonsourceibias.n546 0.189894
R9215 commonsourceibias.n547 commonsourceibias.n378 0.189894
R9216 commonsourceibias.n553 commonsourceibias.n378 0.189894
R9217 commonsourceibias.n554 commonsourceibias.n553 0.189894
R9218 commonsourceibias.n555 commonsourceibias.n554 0.189894
R9219 commonsourceibias.n555 commonsourceibias.n376 0.189894
R9220 commonsourceibias.n560 commonsourceibias.n376 0.189894
R9221 commonsourceibias.n561 commonsourceibias.n560 0.189894
R9222 commonsourceibias.n562 commonsourceibias.n561 0.189894
R9223 commonsourceibias.n562 commonsourceibias.n374 0.189894
R9224 commonsourceibias.n681 commonsourceibias.n680 0.189894
R9225 commonsourceibias.n681 commonsourceibias.n676 0.189894
R9226 commonsourceibias.n686 commonsourceibias.n676 0.189894
R9227 commonsourceibias.n687 commonsourceibias.n686 0.189894
R9228 commonsourceibias.n688 commonsourceibias.n687 0.189894
R9229 commonsourceibias.n688 commonsourceibias.n674 0.189894
R9230 commonsourceibias.n693 commonsourceibias.n674 0.189894
R9231 commonsourceibias.n694 commonsourceibias.n693 0.189894
R9232 commonsourceibias.n694 commonsourceibias.n672 0.189894
R9233 commonsourceibias.n698 commonsourceibias.n672 0.189894
R9234 commonsourceibias.n699 commonsourceibias.n698 0.189894
R9235 commonsourceibias.n699 commonsourceibias.n670 0.189894
R9236 commonsourceibias.n703 commonsourceibias.n670 0.189894
R9237 commonsourceibias.n704 commonsourceibias.n703 0.189894
R9238 commonsourceibias.n704 commonsourceibias.n668 0.189894
R9239 commonsourceibias.n709 commonsourceibias.n668 0.189894
R9240 commonsourceibias.n710 commonsourceibias.n709 0.189894
R9241 commonsourceibias.n711 commonsourceibias.n710 0.189894
R9242 commonsourceibias.n711 commonsourceibias.n666 0.189894
R9243 commonsourceibias.n717 commonsourceibias.n666 0.189894
R9244 commonsourceibias.n718 commonsourceibias.n717 0.189894
R9245 commonsourceibias.n719 commonsourceibias.n718 0.189894
R9246 commonsourceibias.n719 commonsourceibias.n664 0.189894
R9247 commonsourceibias.n724 commonsourceibias.n664 0.189894
R9248 commonsourceibias.n725 commonsourceibias.n724 0.189894
R9249 commonsourceibias.n726 commonsourceibias.n725 0.189894
R9250 commonsourceibias.n726 commonsourceibias.n662 0.189894
R9251 commonsourceibias.n732 commonsourceibias.n662 0.189894
R9252 commonsourceibias.n733 commonsourceibias.n732 0.189894
R9253 commonsourceibias.n734 commonsourceibias.n733 0.189894
R9254 commonsourceibias.n734 commonsourceibias.n660 0.189894
R9255 commonsourceibias.n739 commonsourceibias.n660 0.189894
R9256 commonsourceibias.n740 commonsourceibias.n739 0.189894
R9257 commonsourceibias.n741 commonsourceibias.n740 0.189894
R9258 commonsourceibias.n741 commonsourceibias.n658 0.189894
R9259 commonsourceibias.n591 commonsourceibias.n590 0.189894
R9260 commonsourceibias.n591 commonsourceibias.n586 0.189894
R9261 commonsourceibias.n596 commonsourceibias.n586 0.189894
R9262 commonsourceibias.n597 commonsourceibias.n596 0.189894
R9263 commonsourceibias.n598 commonsourceibias.n597 0.189894
R9264 commonsourceibias.n598 commonsourceibias.n584 0.189894
R9265 commonsourceibias.n603 commonsourceibias.n584 0.189894
R9266 commonsourceibias.n604 commonsourceibias.n603 0.189894
R9267 commonsourceibias.n604 commonsourceibias.n582 0.189894
R9268 commonsourceibias.n608 commonsourceibias.n582 0.189894
R9269 commonsourceibias.n609 commonsourceibias.n608 0.189894
R9270 commonsourceibias.n609 commonsourceibias.n580 0.189894
R9271 commonsourceibias.n613 commonsourceibias.n580 0.189894
R9272 commonsourceibias.n614 commonsourceibias.n613 0.189894
R9273 commonsourceibias.n614 commonsourceibias.n578 0.189894
R9274 commonsourceibias.n619 commonsourceibias.n578 0.189894
R9275 commonsourceibias.n620 commonsourceibias.n619 0.189894
R9276 commonsourceibias.n621 commonsourceibias.n620 0.189894
R9277 commonsourceibias.n621 commonsourceibias.n576 0.189894
R9278 commonsourceibias.n627 commonsourceibias.n576 0.189894
R9279 commonsourceibias.n628 commonsourceibias.n627 0.189894
R9280 commonsourceibias.n629 commonsourceibias.n628 0.189894
R9281 commonsourceibias.n629 commonsourceibias.n574 0.189894
R9282 commonsourceibias.n634 commonsourceibias.n574 0.189894
R9283 commonsourceibias.n635 commonsourceibias.n634 0.189894
R9284 commonsourceibias.n636 commonsourceibias.n635 0.189894
R9285 commonsourceibias.n636 commonsourceibias.n572 0.189894
R9286 commonsourceibias.n642 commonsourceibias.n572 0.189894
R9287 commonsourceibias.n643 commonsourceibias.n642 0.189894
R9288 commonsourceibias.n644 commonsourceibias.n643 0.189894
R9289 commonsourceibias.n644 commonsourceibias.n570 0.189894
R9290 commonsourceibias.n649 commonsourceibias.n570 0.189894
R9291 commonsourceibias.n650 commonsourceibias.n649 0.189894
R9292 commonsourceibias.n651 commonsourceibias.n650 0.189894
R9293 commonsourceibias.n651 commonsourceibias.n568 0.189894
R9294 commonsourceibias.n159 commonsourceibias.n158 0.170955
R9295 commonsourceibias.n160 commonsourceibias.n159 0.170955
R9296 commonsourceibias.n531 commonsourceibias.n425 0.170955
R9297 commonsourceibias.n532 commonsourceibias.n531 0.170955
R9298 gnd.n7129 gnd.n525 1768.67
R9299 gnd.n5093 gnd.n5092 939.716
R9300 gnd.n7604 gnd.n208 795.207
R9301 gnd.n348 gnd.n211 795.207
R9302 gnd.n1787 gnd.n1675 795.207
R9303 gnd.n4398 gnd.n1789 795.207
R9304 gnd.n4835 gnd.n1372 795.207
R9305 gnd.n3161 gnd.n1375 795.207
R9306 gnd.n2807 gnd.n1067 795.207
R9307 gnd.n2763 gnd.n2762 795.207
R9308 gnd.n3223 gnd.n2412 771.183
R9309 gnd.n4123 gnd.n1614 771.183
R9310 gnd.n3154 gnd.n2409 771.183
R9311 gnd.n4180 gnd.n1977 771.183
R9312 gnd.n6475 gnd.n1026 766.379
R9313 gnd.n6391 gnd.n1028 766.379
R9314 gnd.n5603 gnd.n5502 766.379
R9315 gnd.n5601 gnd.n5504 766.379
R9316 gnd.n6472 gnd.n5095 756.769
R9317 gnd.n6441 gnd.n1029 756.769
R9318 gnd.n5735 gnd.n5464 756.769
R9319 gnd.n5721 gnd.n5453 756.769
R9320 gnd.n7602 gnd.n213 739.952
R9321 gnd.n7493 gnd.n210 739.952
R9322 gnd.n4401 gnd.n4400 739.952
R9323 gnd.n4518 gnd.n1721 739.952
R9324 gnd.n4833 gnd.n1377 739.952
R9325 gnd.n2551 gnd.n1374 739.952
R9326 gnd.n4970 gnd.n1140 739.952
R9327 gnd.n5090 gnd.n1071 739.952
R9328 gnd.n6676 gnd.n800 670.282
R9329 gnd.n7130 gnd.n526 670.282
R9330 gnd.n7343 gnd.n399 670.282
R9331 gnd.n2727 gnd.n2726 670.282
R9332 gnd.n6676 gnd.n6675 585
R9333 gnd.n6677 gnd.n6676 585
R9334 gnd.n6674 gnd.n802 585
R9335 gnd.n802 gnd.n801 585
R9336 gnd.n6673 gnd.n6672 585
R9337 gnd.n6672 gnd.n6671 585
R9338 gnd.n807 gnd.n806 585
R9339 gnd.n6670 gnd.n807 585
R9340 gnd.n6668 gnd.n6667 585
R9341 gnd.n6669 gnd.n6668 585
R9342 gnd.n6666 gnd.n809 585
R9343 gnd.n809 gnd.n808 585
R9344 gnd.n6665 gnd.n6664 585
R9345 gnd.n6664 gnd.n6663 585
R9346 gnd.n815 gnd.n814 585
R9347 gnd.n6662 gnd.n815 585
R9348 gnd.n6660 gnd.n6659 585
R9349 gnd.n6661 gnd.n6660 585
R9350 gnd.n6658 gnd.n817 585
R9351 gnd.n817 gnd.n816 585
R9352 gnd.n6657 gnd.n6656 585
R9353 gnd.n6656 gnd.n6655 585
R9354 gnd.n823 gnd.n822 585
R9355 gnd.n6654 gnd.n823 585
R9356 gnd.n6652 gnd.n6651 585
R9357 gnd.n6653 gnd.n6652 585
R9358 gnd.n6650 gnd.n825 585
R9359 gnd.n825 gnd.n824 585
R9360 gnd.n6649 gnd.n6648 585
R9361 gnd.n6648 gnd.n6647 585
R9362 gnd.n831 gnd.n830 585
R9363 gnd.n6646 gnd.n831 585
R9364 gnd.n6644 gnd.n6643 585
R9365 gnd.n6645 gnd.n6644 585
R9366 gnd.n6642 gnd.n833 585
R9367 gnd.n833 gnd.n832 585
R9368 gnd.n6641 gnd.n6640 585
R9369 gnd.n6640 gnd.n6639 585
R9370 gnd.n839 gnd.n838 585
R9371 gnd.n6638 gnd.n839 585
R9372 gnd.n6636 gnd.n6635 585
R9373 gnd.n6637 gnd.n6636 585
R9374 gnd.n6634 gnd.n841 585
R9375 gnd.n841 gnd.n840 585
R9376 gnd.n6633 gnd.n6632 585
R9377 gnd.n6632 gnd.n6631 585
R9378 gnd.n847 gnd.n846 585
R9379 gnd.n6630 gnd.n847 585
R9380 gnd.n6628 gnd.n6627 585
R9381 gnd.n6629 gnd.n6628 585
R9382 gnd.n6626 gnd.n849 585
R9383 gnd.n849 gnd.n848 585
R9384 gnd.n6625 gnd.n6624 585
R9385 gnd.n6624 gnd.n6623 585
R9386 gnd.n855 gnd.n854 585
R9387 gnd.n6622 gnd.n855 585
R9388 gnd.n6620 gnd.n6619 585
R9389 gnd.n6621 gnd.n6620 585
R9390 gnd.n6618 gnd.n857 585
R9391 gnd.n857 gnd.n856 585
R9392 gnd.n6617 gnd.n6616 585
R9393 gnd.n6616 gnd.n6615 585
R9394 gnd.n863 gnd.n862 585
R9395 gnd.n6614 gnd.n863 585
R9396 gnd.n6612 gnd.n6611 585
R9397 gnd.n6613 gnd.n6612 585
R9398 gnd.n6610 gnd.n865 585
R9399 gnd.n865 gnd.n864 585
R9400 gnd.n6609 gnd.n6608 585
R9401 gnd.n6608 gnd.n6607 585
R9402 gnd.n871 gnd.n870 585
R9403 gnd.n6606 gnd.n871 585
R9404 gnd.n6604 gnd.n6603 585
R9405 gnd.n6605 gnd.n6604 585
R9406 gnd.n6602 gnd.n873 585
R9407 gnd.n873 gnd.n872 585
R9408 gnd.n6601 gnd.n6600 585
R9409 gnd.n6600 gnd.n6599 585
R9410 gnd.n879 gnd.n878 585
R9411 gnd.n6598 gnd.n879 585
R9412 gnd.n6596 gnd.n6595 585
R9413 gnd.n6597 gnd.n6596 585
R9414 gnd.n6594 gnd.n881 585
R9415 gnd.n881 gnd.n880 585
R9416 gnd.n6593 gnd.n6592 585
R9417 gnd.n6592 gnd.n6591 585
R9418 gnd.n887 gnd.n886 585
R9419 gnd.n6590 gnd.n887 585
R9420 gnd.n6588 gnd.n6587 585
R9421 gnd.n6589 gnd.n6588 585
R9422 gnd.n6586 gnd.n889 585
R9423 gnd.n889 gnd.n888 585
R9424 gnd.n6585 gnd.n6584 585
R9425 gnd.n6584 gnd.n6583 585
R9426 gnd.n895 gnd.n894 585
R9427 gnd.n6582 gnd.n895 585
R9428 gnd.n6580 gnd.n6579 585
R9429 gnd.n6581 gnd.n6580 585
R9430 gnd.n6578 gnd.n897 585
R9431 gnd.n897 gnd.n896 585
R9432 gnd.n6577 gnd.n6576 585
R9433 gnd.n6576 gnd.n6575 585
R9434 gnd.n903 gnd.n902 585
R9435 gnd.n6574 gnd.n903 585
R9436 gnd.n6572 gnd.n6571 585
R9437 gnd.n6573 gnd.n6572 585
R9438 gnd.n6570 gnd.n905 585
R9439 gnd.n905 gnd.n904 585
R9440 gnd.n6569 gnd.n6568 585
R9441 gnd.n6568 gnd.n6567 585
R9442 gnd.n911 gnd.n910 585
R9443 gnd.n6566 gnd.n911 585
R9444 gnd.n6564 gnd.n6563 585
R9445 gnd.n6565 gnd.n6564 585
R9446 gnd.n6562 gnd.n913 585
R9447 gnd.n913 gnd.n912 585
R9448 gnd.n6561 gnd.n6560 585
R9449 gnd.n6560 gnd.n6559 585
R9450 gnd.n919 gnd.n918 585
R9451 gnd.n6558 gnd.n919 585
R9452 gnd.n6556 gnd.n6555 585
R9453 gnd.n6557 gnd.n6556 585
R9454 gnd.n6554 gnd.n921 585
R9455 gnd.n921 gnd.n920 585
R9456 gnd.n6553 gnd.n6552 585
R9457 gnd.n6552 gnd.n6551 585
R9458 gnd.n927 gnd.n926 585
R9459 gnd.n6550 gnd.n927 585
R9460 gnd.n6548 gnd.n6547 585
R9461 gnd.n6549 gnd.n6548 585
R9462 gnd.n6546 gnd.n929 585
R9463 gnd.n929 gnd.n928 585
R9464 gnd.n6545 gnd.n6544 585
R9465 gnd.n6544 gnd.n6543 585
R9466 gnd.n935 gnd.n934 585
R9467 gnd.n6542 gnd.n935 585
R9468 gnd.n6540 gnd.n6539 585
R9469 gnd.n6541 gnd.n6540 585
R9470 gnd.n6538 gnd.n937 585
R9471 gnd.n937 gnd.n936 585
R9472 gnd.n6537 gnd.n6536 585
R9473 gnd.n6536 gnd.n6535 585
R9474 gnd.n943 gnd.n942 585
R9475 gnd.n6534 gnd.n943 585
R9476 gnd.n6532 gnd.n6531 585
R9477 gnd.n6533 gnd.n6532 585
R9478 gnd.n6530 gnd.n945 585
R9479 gnd.n945 gnd.n944 585
R9480 gnd.n6529 gnd.n6528 585
R9481 gnd.n6528 gnd.n6527 585
R9482 gnd.n951 gnd.n950 585
R9483 gnd.n6526 gnd.n951 585
R9484 gnd.n6524 gnd.n6523 585
R9485 gnd.n6525 gnd.n6524 585
R9486 gnd.n6522 gnd.n953 585
R9487 gnd.n953 gnd.n952 585
R9488 gnd.n6521 gnd.n6520 585
R9489 gnd.n6520 gnd.n6519 585
R9490 gnd.n959 gnd.n958 585
R9491 gnd.n6518 gnd.n959 585
R9492 gnd.n6516 gnd.n6515 585
R9493 gnd.n6517 gnd.n6516 585
R9494 gnd.n6514 gnd.n961 585
R9495 gnd.n961 gnd.n960 585
R9496 gnd.n6513 gnd.n6512 585
R9497 gnd.n6512 gnd.n6511 585
R9498 gnd.n967 gnd.n966 585
R9499 gnd.n6510 gnd.n967 585
R9500 gnd.n800 gnd.n799 585
R9501 gnd.n6678 gnd.n800 585
R9502 gnd.n6681 gnd.n6680 585
R9503 gnd.n6680 gnd.n6679 585
R9504 gnd.n797 gnd.n796 585
R9505 gnd.n796 gnd.n795 585
R9506 gnd.n6686 gnd.n6685 585
R9507 gnd.n6687 gnd.n6686 585
R9508 gnd.n794 gnd.n793 585
R9509 gnd.n6688 gnd.n794 585
R9510 gnd.n6691 gnd.n6690 585
R9511 gnd.n6690 gnd.n6689 585
R9512 gnd.n791 gnd.n790 585
R9513 gnd.n790 gnd.n789 585
R9514 gnd.n6696 gnd.n6695 585
R9515 gnd.n6697 gnd.n6696 585
R9516 gnd.n788 gnd.n787 585
R9517 gnd.n6698 gnd.n788 585
R9518 gnd.n6701 gnd.n6700 585
R9519 gnd.n6700 gnd.n6699 585
R9520 gnd.n785 gnd.n784 585
R9521 gnd.n784 gnd.n783 585
R9522 gnd.n6706 gnd.n6705 585
R9523 gnd.n6707 gnd.n6706 585
R9524 gnd.n782 gnd.n781 585
R9525 gnd.n6708 gnd.n782 585
R9526 gnd.n6711 gnd.n6710 585
R9527 gnd.n6710 gnd.n6709 585
R9528 gnd.n779 gnd.n778 585
R9529 gnd.n778 gnd.n777 585
R9530 gnd.n6716 gnd.n6715 585
R9531 gnd.n6717 gnd.n6716 585
R9532 gnd.n776 gnd.n775 585
R9533 gnd.n6718 gnd.n776 585
R9534 gnd.n6721 gnd.n6720 585
R9535 gnd.n6720 gnd.n6719 585
R9536 gnd.n773 gnd.n772 585
R9537 gnd.n772 gnd.n771 585
R9538 gnd.n6726 gnd.n6725 585
R9539 gnd.n6727 gnd.n6726 585
R9540 gnd.n770 gnd.n769 585
R9541 gnd.n6728 gnd.n770 585
R9542 gnd.n6731 gnd.n6730 585
R9543 gnd.n6730 gnd.n6729 585
R9544 gnd.n767 gnd.n766 585
R9545 gnd.n766 gnd.n765 585
R9546 gnd.n6736 gnd.n6735 585
R9547 gnd.n6737 gnd.n6736 585
R9548 gnd.n764 gnd.n763 585
R9549 gnd.n6738 gnd.n764 585
R9550 gnd.n6741 gnd.n6740 585
R9551 gnd.n6740 gnd.n6739 585
R9552 gnd.n761 gnd.n760 585
R9553 gnd.n760 gnd.n759 585
R9554 gnd.n6746 gnd.n6745 585
R9555 gnd.n6747 gnd.n6746 585
R9556 gnd.n758 gnd.n757 585
R9557 gnd.n6748 gnd.n758 585
R9558 gnd.n6751 gnd.n6750 585
R9559 gnd.n6750 gnd.n6749 585
R9560 gnd.n755 gnd.n754 585
R9561 gnd.n754 gnd.n753 585
R9562 gnd.n6756 gnd.n6755 585
R9563 gnd.n6757 gnd.n6756 585
R9564 gnd.n752 gnd.n751 585
R9565 gnd.n6758 gnd.n752 585
R9566 gnd.n6761 gnd.n6760 585
R9567 gnd.n6760 gnd.n6759 585
R9568 gnd.n749 gnd.n748 585
R9569 gnd.n748 gnd.n747 585
R9570 gnd.n6766 gnd.n6765 585
R9571 gnd.n6767 gnd.n6766 585
R9572 gnd.n746 gnd.n745 585
R9573 gnd.n6768 gnd.n746 585
R9574 gnd.n6771 gnd.n6770 585
R9575 gnd.n6770 gnd.n6769 585
R9576 gnd.n743 gnd.n742 585
R9577 gnd.n742 gnd.n741 585
R9578 gnd.n6776 gnd.n6775 585
R9579 gnd.n6777 gnd.n6776 585
R9580 gnd.n740 gnd.n739 585
R9581 gnd.n6778 gnd.n740 585
R9582 gnd.n6781 gnd.n6780 585
R9583 gnd.n6780 gnd.n6779 585
R9584 gnd.n737 gnd.n736 585
R9585 gnd.n736 gnd.n735 585
R9586 gnd.n6786 gnd.n6785 585
R9587 gnd.n6787 gnd.n6786 585
R9588 gnd.n734 gnd.n733 585
R9589 gnd.n6788 gnd.n734 585
R9590 gnd.n6791 gnd.n6790 585
R9591 gnd.n6790 gnd.n6789 585
R9592 gnd.n731 gnd.n730 585
R9593 gnd.n730 gnd.n729 585
R9594 gnd.n6796 gnd.n6795 585
R9595 gnd.n6797 gnd.n6796 585
R9596 gnd.n728 gnd.n727 585
R9597 gnd.n6798 gnd.n728 585
R9598 gnd.n6801 gnd.n6800 585
R9599 gnd.n6800 gnd.n6799 585
R9600 gnd.n725 gnd.n724 585
R9601 gnd.n724 gnd.n723 585
R9602 gnd.n6806 gnd.n6805 585
R9603 gnd.n6807 gnd.n6806 585
R9604 gnd.n722 gnd.n721 585
R9605 gnd.n6808 gnd.n722 585
R9606 gnd.n6811 gnd.n6810 585
R9607 gnd.n6810 gnd.n6809 585
R9608 gnd.n719 gnd.n718 585
R9609 gnd.n718 gnd.n717 585
R9610 gnd.n6816 gnd.n6815 585
R9611 gnd.n6817 gnd.n6816 585
R9612 gnd.n716 gnd.n715 585
R9613 gnd.n6818 gnd.n716 585
R9614 gnd.n6821 gnd.n6820 585
R9615 gnd.n6820 gnd.n6819 585
R9616 gnd.n713 gnd.n712 585
R9617 gnd.n712 gnd.n711 585
R9618 gnd.n6826 gnd.n6825 585
R9619 gnd.n6827 gnd.n6826 585
R9620 gnd.n710 gnd.n709 585
R9621 gnd.n6828 gnd.n710 585
R9622 gnd.n6831 gnd.n6830 585
R9623 gnd.n6830 gnd.n6829 585
R9624 gnd.n707 gnd.n706 585
R9625 gnd.n706 gnd.n705 585
R9626 gnd.n6836 gnd.n6835 585
R9627 gnd.n6837 gnd.n6836 585
R9628 gnd.n704 gnd.n703 585
R9629 gnd.n6838 gnd.n704 585
R9630 gnd.n6841 gnd.n6840 585
R9631 gnd.n6840 gnd.n6839 585
R9632 gnd.n701 gnd.n700 585
R9633 gnd.n700 gnd.n699 585
R9634 gnd.n6846 gnd.n6845 585
R9635 gnd.n6847 gnd.n6846 585
R9636 gnd.n698 gnd.n697 585
R9637 gnd.n6848 gnd.n698 585
R9638 gnd.n6851 gnd.n6850 585
R9639 gnd.n6850 gnd.n6849 585
R9640 gnd.n695 gnd.n694 585
R9641 gnd.n694 gnd.n693 585
R9642 gnd.n6856 gnd.n6855 585
R9643 gnd.n6857 gnd.n6856 585
R9644 gnd.n692 gnd.n691 585
R9645 gnd.n6858 gnd.n692 585
R9646 gnd.n6861 gnd.n6860 585
R9647 gnd.n6860 gnd.n6859 585
R9648 gnd.n689 gnd.n688 585
R9649 gnd.n688 gnd.n687 585
R9650 gnd.n6866 gnd.n6865 585
R9651 gnd.n6867 gnd.n6866 585
R9652 gnd.n686 gnd.n685 585
R9653 gnd.n6868 gnd.n686 585
R9654 gnd.n6871 gnd.n6870 585
R9655 gnd.n6870 gnd.n6869 585
R9656 gnd.n683 gnd.n682 585
R9657 gnd.n682 gnd.n681 585
R9658 gnd.n6876 gnd.n6875 585
R9659 gnd.n6877 gnd.n6876 585
R9660 gnd.n680 gnd.n679 585
R9661 gnd.n6878 gnd.n680 585
R9662 gnd.n6881 gnd.n6880 585
R9663 gnd.n6880 gnd.n6879 585
R9664 gnd.n677 gnd.n676 585
R9665 gnd.n676 gnd.n675 585
R9666 gnd.n6886 gnd.n6885 585
R9667 gnd.n6887 gnd.n6886 585
R9668 gnd.n674 gnd.n673 585
R9669 gnd.n6888 gnd.n674 585
R9670 gnd.n6891 gnd.n6890 585
R9671 gnd.n6890 gnd.n6889 585
R9672 gnd.n671 gnd.n670 585
R9673 gnd.n670 gnd.n669 585
R9674 gnd.n6896 gnd.n6895 585
R9675 gnd.n6897 gnd.n6896 585
R9676 gnd.n668 gnd.n667 585
R9677 gnd.n6898 gnd.n668 585
R9678 gnd.n6901 gnd.n6900 585
R9679 gnd.n6900 gnd.n6899 585
R9680 gnd.n665 gnd.n664 585
R9681 gnd.n664 gnd.n663 585
R9682 gnd.n6906 gnd.n6905 585
R9683 gnd.n6907 gnd.n6906 585
R9684 gnd.n662 gnd.n661 585
R9685 gnd.n6908 gnd.n662 585
R9686 gnd.n6911 gnd.n6910 585
R9687 gnd.n6910 gnd.n6909 585
R9688 gnd.n659 gnd.n658 585
R9689 gnd.n658 gnd.n657 585
R9690 gnd.n6916 gnd.n6915 585
R9691 gnd.n6917 gnd.n6916 585
R9692 gnd.n656 gnd.n655 585
R9693 gnd.n6918 gnd.n656 585
R9694 gnd.n6921 gnd.n6920 585
R9695 gnd.n6920 gnd.n6919 585
R9696 gnd.n653 gnd.n652 585
R9697 gnd.n652 gnd.n651 585
R9698 gnd.n6926 gnd.n6925 585
R9699 gnd.n6927 gnd.n6926 585
R9700 gnd.n650 gnd.n649 585
R9701 gnd.n6928 gnd.n650 585
R9702 gnd.n6931 gnd.n6930 585
R9703 gnd.n6930 gnd.n6929 585
R9704 gnd.n647 gnd.n646 585
R9705 gnd.n646 gnd.n645 585
R9706 gnd.n6936 gnd.n6935 585
R9707 gnd.n6937 gnd.n6936 585
R9708 gnd.n644 gnd.n643 585
R9709 gnd.n6938 gnd.n644 585
R9710 gnd.n6941 gnd.n6940 585
R9711 gnd.n6940 gnd.n6939 585
R9712 gnd.n641 gnd.n640 585
R9713 gnd.n640 gnd.n639 585
R9714 gnd.n6946 gnd.n6945 585
R9715 gnd.n6947 gnd.n6946 585
R9716 gnd.n638 gnd.n637 585
R9717 gnd.n6948 gnd.n638 585
R9718 gnd.n6951 gnd.n6950 585
R9719 gnd.n6950 gnd.n6949 585
R9720 gnd.n635 gnd.n634 585
R9721 gnd.n634 gnd.n633 585
R9722 gnd.n6956 gnd.n6955 585
R9723 gnd.n6957 gnd.n6956 585
R9724 gnd.n632 gnd.n631 585
R9725 gnd.n6958 gnd.n632 585
R9726 gnd.n6961 gnd.n6960 585
R9727 gnd.n6960 gnd.n6959 585
R9728 gnd.n629 gnd.n628 585
R9729 gnd.n628 gnd.n627 585
R9730 gnd.n6966 gnd.n6965 585
R9731 gnd.n6967 gnd.n6966 585
R9732 gnd.n626 gnd.n625 585
R9733 gnd.n6968 gnd.n626 585
R9734 gnd.n6971 gnd.n6970 585
R9735 gnd.n6970 gnd.n6969 585
R9736 gnd.n623 gnd.n622 585
R9737 gnd.n622 gnd.n621 585
R9738 gnd.n6976 gnd.n6975 585
R9739 gnd.n6977 gnd.n6976 585
R9740 gnd.n620 gnd.n619 585
R9741 gnd.n6978 gnd.n620 585
R9742 gnd.n6981 gnd.n6980 585
R9743 gnd.n6980 gnd.n6979 585
R9744 gnd.n617 gnd.n616 585
R9745 gnd.n616 gnd.n615 585
R9746 gnd.n6986 gnd.n6985 585
R9747 gnd.n6987 gnd.n6986 585
R9748 gnd.n614 gnd.n613 585
R9749 gnd.n6988 gnd.n614 585
R9750 gnd.n6991 gnd.n6990 585
R9751 gnd.n6990 gnd.n6989 585
R9752 gnd.n611 gnd.n610 585
R9753 gnd.n610 gnd.n609 585
R9754 gnd.n6996 gnd.n6995 585
R9755 gnd.n6997 gnd.n6996 585
R9756 gnd.n608 gnd.n607 585
R9757 gnd.n6998 gnd.n608 585
R9758 gnd.n7001 gnd.n7000 585
R9759 gnd.n7000 gnd.n6999 585
R9760 gnd.n605 gnd.n604 585
R9761 gnd.n604 gnd.n603 585
R9762 gnd.n7006 gnd.n7005 585
R9763 gnd.n7007 gnd.n7006 585
R9764 gnd.n602 gnd.n601 585
R9765 gnd.n7008 gnd.n602 585
R9766 gnd.n7011 gnd.n7010 585
R9767 gnd.n7010 gnd.n7009 585
R9768 gnd.n599 gnd.n598 585
R9769 gnd.n598 gnd.n597 585
R9770 gnd.n7016 gnd.n7015 585
R9771 gnd.n7017 gnd.n7016 585
R9772 gnd.n596 gnd.n595 585
R9773 gnd.n7018 gnd.n596 585
R9774 gnd.n7021 gnd.n7020 585
R9775 gnd.n7020 gnd.n7019 585
R9776 gnd.n593 gnd.n592 585
R9777 gnd.n592 gnd.n591 585
R9778 gnd.n7026 gnd.n7025 585
R9779 gnd.n7027 gnd.n7026 585
R9780 gnd.n590 gnd.n589 585
R9781 gnd.n7028 gnd.n590 585
R9782 gnd.n7031 gnd.n7030 585
R9783 gnd.n7030 gnd.n7029 585
R9784 gnd.n587 gnd.n586 585
R9785 gnd.n586 gnd.n585 585
R9786 gnd.n7036 gnd.n7035 585
R9787 gnd.n7037 gnd.n7036 585
R9788 gnd.n584 gnd.n583 585
R9789 gnd.n7038 gnd.n584 585
R9790 gnd.n7041 gnd.n7040 585
R9791 gnd.n7040 gnd.n7039 585
R9792 gnd.n581 gnd.n580 585
R9793 gnd.n580 gnd.n579 585
R9794 gnd.n7046 gnd.n7045 585
R9795 gnd.n7047 gnd.n7046 585
R9796 gnd.n578 gnd.n577 585
R9797 gnd.n7048 gnd.n578 585
R9798 gnd.n7051 gnd.n7050 585
R9799 gnd.n7050 gnd.n7049 585
R9800 gnd.n575 gnd.n574 585
R9801 gnd.n574 gnd.n573 585
R9802 gnd.n7056 gnd.n7055 585
R9803 gnd.n7057 gnd.n7056 585
R9804 gnd.n572 gnd.n571 585
R9805 gnd.n7058 gnd.n572 585
R9806 gnd.n7061 gnd.n7060 585
R9807 gnd.n7060 gnd.n7059 585
R9808 gnd.n569 gnd.n568 585
R9809 gnd.n568 gnd.n567 585
R9810 gnd.n7066 gnd.n7065 585
R9811 gnd.n7067 gnd.n7066 585
R9812 gnd.n566 gnd.n565 585
R9813 gnd.n7068 gnd.n566 585
R9814 gnd.n7071 gnd.n7070 585
R9815 gnd.n7070 gnd.n7069 585
R9816 gnd.n563 gnd.n562 585
R9817 gnd.n562 gnd.n561 585
R9818 gnd.n7076 gnd.n7075 585
R9819 gnd.n7077 gnd.n7076 585
R9820 gnd.n560 gnd.n559 585
R9821 gnd.n7078 gnd.n560 585
R9822 gnd.n7081 gnd.n7080 585
R9823 gnd.n7080 gnd.n7079 585
R9824 gnd.n557 gnd.n556 585
R9825 gnd.n556 gnd.n555 585
R9826 gnd.n7086 gnd.n7085 585
R9827 gnd.n7087 gnd.n7086 585
R9828 gnd.n554 gnd.n553 585
R9829 gnd.n7088 gnd.n554 585
R9830 gnd.n7091 gnd.n7090 585
R9831 gnd.n7090 gnd.n7089 585
R9832 gnd.n551 gnd.n550 585
R9833 gnd.n550 gnd.n549 585
R9834 gnd.n7096 gnd.n7095 585
R9835 gnd.n7097 gnd.n7096 585
R9836 gnd.n548 gnd.n547 585
R9837 gnd.n7098 gnd.n548 585
R9838 gnd.n7101 gnd.n7100 585
R9839 gnd.n7100 gnd.n7099 585
R9840 gnd.n545 gnd.n544 585
R9841 gnd.n544 gnd.n543 585
R9842 gnd.n7106 gnd.n7105 585
R9843 gnd.n7107 gnd.n7106 585
R9844 gnd.n542 gnd.n541 585
R9845 gnd.n7108 gnd.n542 585
R9846 gnd.n7111 gnd.n7110 585
R9847 gnd.n7110 gnd.n7109 585
R9848 gnd.n539 gnd.n538 585
R9849 gnd.n538 gnd.n537 585
R9850 gnd.n7116 gnd.n7115 585
R9851 gnd.n7117 gnd.n7116 585
R9852 gnd.n536 gnd.n535 585
R9853 gnd.n7118 gnd.n536 585
R9854 gnd.n7121 gnd.n7120 585
R9855 gnd.n7120 gnd.n7119 585
R9856 gnd.n533 gnd.n532 585
R9857 gnd.n532 gnd.n531 585
R9858 gnd.n7126 gnd.n7125 585
R9859 gnd.n7127 gnd.n7126 585
R9860 gnd.n530 gnd.n529 585
R9861 gnd.n7128 gnd.n530 585
R9862 gnd.n7131 gnd.n7130 585
R9863 gnd.n7130 gnd.n7129 585
R9864 gnd.n7342 gnd.n403 585
R9865 gnd.n7342 gnd.n7341 585
R9866 gnd.n7336 gnd.n404 585
R9867 gnd.n7340 gnd.n404 585
R9868 gnd.n7338 gnd.n7337 585
R9869 gnd.n7339 gnd.n7338 585
R9870 gnd.n407 gnd.n406 585
R9871 gnd.n406 gnd.n405 585
R9872 gnd.n7331 gnd.n7330 585
R9873 gnd.n7330 gnd.n7329 585
R9874 gnd.n410 gnd.n409 585
R9875 gnd.n7328 gnd.n410 585
R9876 gnd.n7326 gnd.n7325 585
R9877 gnd.n7327 gnd.n7326 585
R9878 gnd.n413 gnd.n412 585
R9879 gnd.n412 gnd.n411 585
R9880 gnd.n7321 gnd.n7320 585
R9881 gnd.n7320 gnd.n7319 585
R9882 gnd.n416 gnd.n415 585
R9883 gnd.n7318 gnd.n416 585
R9884 gnd.n7316 gnd.n7315 585
R9885 gnd.n7317 gnd.n7316 585
R9886 gnd.n419 gnd.n418 585
R9887 gnd.n418 gnd.n417 585
R9888 gnd.n7311 gnd.n7310 585
R9889 gnd.n7310 gnd.n7309 585
R9890 gnd.n422 gnd.n421 585
R9891 gnd.n7308 gnd.n422 585
R9892 gnd.n7306 gnd.n7305 585
R9893 gnd.n7307 gnd.n7306 585
R9894 gnd.n425 gnd.n424 585
R9895 gnd.n424 gnd.n423 585
R9896 gnd.n7301 gnd.n7300 585
R9897 gnd.n7300 gnd.n7299 585
R9898 gnd.n428 gnd.n427 585
R9899 gnd.n7298 gnd.n428 585
R9900 gnd.n7296 gnd.n7295 585
R9901 gnd.n7297 gnd.n7296 585
R9902 gnd.n431 gnd.n430 585
R9903 gnd.n430 gnd.n429 585
R9904 gnd.n7291 gnd.n7290 585
R9905 gnd.n7290 gnd.n7289 585
R9906 gnd.n434 gnd.n433 585
R9907 gnd.n7288 gnd.n434 585
R9908 gnd.n7286 gnd.n7285 585
R9909 gnd.n7287 gnd.n7286 585
R9910 gnd.n437 gnd.n436 585
R9911 gnd.n436 gnd.n435 585
R9912 gnd.n7281 gnd.n7280 585
R9913 gnd.n7280 gnd.n7279 585
R9914 gnd.n440 gnd.n439 585
R9915 gnd.n7278 gnd.n440 585
R9916 gnd.n7276 gnd.n7275 585
R9917 gnd.n7277 gnd.n7276 585
R9918 gnd.n443 gnd.n442 585
R9919 gnd.n442 gnd.n441 585
R9920 gnd.n7271 gnd.n7270 585
R9921 gnd.n7270 gnd.n7269 585
R9922 gnd.n446 gnd.n445 585
R9923 gnd.n7268 gnd.n446 585
R9924 gnd.n7266 gnd.n7265 585
R9925 gnd.n7267 gnd.n7266 585
R9926 gnd.n449 gnd.n448 585
R9927 gnd.n448 gnd.n447 585
R9928 gnd.n7261 gnd.n7260 585
R9929 gnd.n7260 gnd.n7259 585
R9930 gnd.n452 gnd.n451 585
R9931 gnd.n7258 gnd.n452 585
R9932 gnd.n7256 gnd.n7255 585
R9933 gnd.n7257 gnd.n7256 585
R9934 gnd.n455 gnd.n454 585
R9935 gnd.n454 gnd.n453 585
R9936 gnd.n7251 gnd.n7250 585
R9937 gnd.n7250 gnd.n7249 585
R9938 gnd.n458 gnd.n457 585
R9939 gnd.n7248 gnd.n458 585
R9940 gnd.n7246 gnd.n7245 585
R9941 gnd.n7247 gnd.n7246 585
R9942 gnd.n461 gnd.n460 585
R9943 gnd.n460 gnd.n459 585
R9944 gnd.n7241 gnd.n7240 585
R9945 gnd.n7240 gnd.n7239 585
R9946 gnd.n464 gnd.n463 585
R9947 gnd.n7238 gnd.n464 585
R9948 gnd.n7236 gnd.n7235 585
R9949 gnd.n7237 gnd.n7236 585
R9950 gnd.n467 gnd.n466 585
R9951 gnd.n466 gnd.n465 585
R9952 gnd.n7231 gnd.n7230 585
R9953 gnd.n7230 gnd.n7229 585
R9954 gnd.n470 gnd.n469 585
R9955 gnd.n7228 gnd.n470 585
R9956 gnd.n7226 gnd.n7225 585
R9957 gnd.n7227 gnd.n7226 585
R9958 gnd.n473 gnd.n472 585
R9959 gnd.n472 gnd.n471 585
R9960 gnd.n7221 gnd.n7220 585
R9961 gnd.n7220 gnd.n7219 585
R9962 gnd.n476 gnd.n475 585
R9963 gnd.n7218 gnd.n476 585
R9964 gnd.n7216 gnd.n7215 585
R9965 gnd.n7217 gnd.n7216 585
R9966 gnd.n479 gnd.n478 585
R9967 gnd.n478 gnd.n477 585
R9968 gnd.n7211 gnd.n7210 585
R9969 gnd.n7210 gnd.n7209 585
R9970 gnd.n482 gnd.n481 585
R9971 gnd.n7208 gnd.n482 585
R9972 gnd.n7206 gnd.n7205 585
R9973 gnd.n7207 gnd.n7206 585
R9974 gnd.n485 gnd.n484 585
R9975 gnd.n484 gnd.n483 585
R9976 gnd.n7201 gnd.n7200 585
R9977 gnd.n7200 gnd.n7199 585
R9978 gnd.n488 gnd.n487 585
R9979 gnd.n7198 gnd.n488 585
R9980 gnd.n7196 gnd.n7195 585
R9981 gnd.n7197 gnd.n7196 585
R9982 gnd.n491 gnd.n490 585
R9983 gnd.n490 gnd.n489 585
R9984 gnd.n7191 gnd.n7190 585
R9985 gnd.n7190 gnd.n7189 585
R9986 gnd.n494 gnd.n493 585
R9987 gnd.n7188 gnd.n494 585
R9988 gnd.n7186 gnd.n7185 585
R9989 gnd.n7187 gnd.n7186 585
R9990 gnd.n497 gnd.n496 585
R9991 gnd.n496 gnd.n495 585
R9992 gnd.n7181 gnd.n7180 585
R9993 gnd.n7180 gnd.n7179 585
R9994 gnd.n500 gnd.n499 585
R9995 gnd.n7178 gnd.n500 585
R9996 gnd.n7176 gnd.n7175 585
R9997 gnd.n7177 gnd.n7176 585
R9998 gnd.n503 gnd.n502 585
R9999 gnd.n502 gnd.n501 585
R10000 gnd.n7171 gnd.n7170 585
R10001 gnd.n7170 gnd.n7169 585
R10002 gnd.n506 gnd.n505 585
R10003 gnd.n7168 gnd.n506 585
R10004 gnd.n7166 gnd.n7165 585
R10005 gnd.n7167 gnd.n7166 585
R10006 gnd.n509 gnd.n508 585
R10007 gnd.n508 gnd.n507 585
R10008 gnd.n7161 gnd.n7160 585
R10009 gnd.n7160 gnd.n7159 585
R10010 gnd.n512 gnd.n511 585
R10011 gnd.n7158 gnd.n512 585
R10012 gnd.n7156 gnd.n7155 585
R10013 gnd.n7157 gnd.n7156 585
R10014 gnd.n515 gnd.n514 585
R10015 gnd.n514 gnd.n513 585
R10016 gnd.n7151 gnd.n7150 585
R10017 gnd.n7150 gnd.n7149 585
R10018 gnd.n518 gnd.n517 585
R10019 gnd.n7148 gnd.n518 585
R10020 gnd.n7146 gnd.n7145 585
R10021 gnd.n7147 gnd.n7146 585
R10022 gnd.n521 gnd.n520 585
R10023 gnd.n520 gnd.n519 585
R10024 gnd.n7141 gnd.n7140 585
R10025 gnd.n7140 gnd.n7139 585
R10026 gnd.n524 gnd.n523 585
R10027 gnd.n7138 gnd.n524 585
R10028 gnd.n7136 gnd.n7135 585
R10029 gnd.n7137 gnd.n7136 585
R10030 gnd.n527 gnd.n526 585
R10031 gnd.n526 gnd.n525 585
R10032 gnd.n4836 gnd.n4835 585
R10033 gnd.n4835 gnd.n4834 585
R10034 gnd.n4837 gnd.n1368 585
R10035 gnd.n3143 gnd.n1368 585
R10036 gnd.n4839 gnd.n4838 585
R10037 gnd.n4840 gnd.n4839 585
R10038 gnd.n1352 gnd.n1351 585
R10039 gnd.n3136 gnd.n1352 585
R10040 gnd.n4848 gnd.n4847 585
R10041 gnd.n4847 gnd.n4846 585
R10042 gnd.n4849 gnd.n1347 585
R10043 gnd.n3127 gnd.n1347 585
R10044 gnd.n4851 gnd.n4850 585
R10045 gnd.n4852 gnd.n4851 585
R10046 gnd.n1332 gnd.n1331 585
R10047 gnd.n3121 gnd.n1332 585
R10048 gnd.n4860 gnd.n4859 585
R10049 gnd.n4859 gnd.n4858 585
R10050 gnd.n4861 gnd.n1327 585
R10051 gnd.n3038 gnd.n1327 585
R10052 gnd.n4863 gnd.n4862 585
R10053 gnd.n4864 gnd.n4863 585
R10054 gnd.n1312 gnd.n1311 585
R10055 gnd.n3032 gnd.n1312 585
R10056 gnd.n4872 gnd.n4871 585
R10057 gnd.n4871 gnd.n4870 585
R10058 gnd.n4873 gnd.n1307 585
R10059 gnd.n3026 gnd.n1307 585
R10060 gnd.n4875 gnd.n4874 585
R10061 gnd.n4876 gnd.n4875 585
R10062 gnd.n1292 gnd.n1291 585
R10063 gnd.n3055 gnd.n1292 585
R10064 gnd.n4884 gnd.n4883 585
R10065 gnd.n4883 gnd.n4882 585
R10066 gnd.n4885 gnd.n1287 585
R10067 gnd.n3019 gnd.n1287 585
R10068 gnd.n4887 gnd.n4886 585
R10069 gnd.n4888 gnd.n4887 585
R10070 gnd.n1273 gnd.n1272 585
R10071 gnd.n3011 gnd.n1273 585
R10072 gnd.n4896 gnd.n4895 585
R10073 gnd.n4895 gnd.n4894 585
R10074 gnd.n4897 gnd.n1267 585
R10075 gnd.n3004 gnd.n1267 585
R10076 gnd.n4899 gnd.n4898 585
R10077 gnd.n4900 gnd.n4899 585
R10078 gnd.n1268 gnd.n1266 585
R10079 gnd.n2996 gnd.n1266 585
R10080 gnd.n2957 gnd.n2675 585
R10081 gnd.n2967 gnd.n2675 585
R10082 gnd.n2958 gnd.n2684 585
R10083 gnd.n2684 gnd.n2673 585
R10084 gnd.n2960 gnd.n2959 585
R10085 gnd.n2961 gnd.n2960 585
R10086 gnd.n2685 gnd.n2683 585
R10087 gnd.n2948 gnd.n2683 585
R10088 gnd.n2930 gnd.n2929 585
R10089 gnd.n2931 gnd.n2930 585
R10090 gnd.n2704 gnd.n2700 585
R10091 gnd.n2934 gnd.n2700 585
R10092 gnd.n2922 gnd.n2921 585
R10093 gnd.n2923 gnd.n2922 585
R10094 gnd.n1244 gnd.n1243 585
R10095 gnd.n2709 gnd.n1244 585
R10096 gnd.n4910 gnd.n4909 585
R10097 gnd.n4909 gnd.n4908 585
R10098 gnd.n4911 gnd.n1239 585
R10099 gnd.n2872 gnd.n1239 585
R10100 gnd.n4913 gnd.n4912 585
R10101 gnd.n4914 gnd.n4913 585
R10102 gnd.n1223 gnd.n1222 585
R10103 gnd.n2878 gnd.n1223 585
R10104 gnd.n4922 gnd.n4921 585
R10105 gnd.n4921 gnd.n4920 585
R10106 gnd.n4923 gnd.n1218 585
R10107 gnd.n2884 gnd.n1218 585
R10108 gnd.n4925 gnd.n4924 585
R10109 gnd.n4926 gnd.n4925 585
R10110 gnd.n1203 gnd.n1202 585
R10111 gnd.n2890 gnd.n1203 585
R10112 gnd.n4934 gnd.n4933 585
R10113 gnd.n4933 gnd.n4932 585
R10114 gnd.n4935 gnd.n1198 585
R10115 gnd.n2851 gnd.n1198 585
R10116 gnd.n4937 gnd.n4936 585
R10117 gnd.n4938 gnd.n4937 585
R10118 gnd.n1183 gnd.n1182 585
R10119 gnd.n2842 gnd.n1183 585
R10120 gnd.n4946 gnd.n4945 585
R10121 gnd.n4945 gnd.n4944 585
R10122 gnd.n4947 gnd.n1178 585
R10123 gnd.n1178 gnd.n1177 585
R10124 gnd.n4949 gnd.n4948 585
R10125 gnd.n4950 gnd.n4949 585
R10126 gnd.n1164 gnd.n1163 585
R10127 gnd.n1167 gnd.n1164 585
R10128 gnd.n4958 gnd.n4957 585
R10129 gnd.n4957 gnd.n4956 585
R10130 gnd.n4959 gnd.n1157 585
R10131 gnd.n1157 gnd.n1155 585
R10132 gnd.n4961 gnd.n4960 585
R10133 gnd.n4962 gnd.n4961 585
R10134 gnd.n1159 gnd.n1156 585
R10135 gnd.n1156 gnd.n1152 585
R10136 gnd.n1158 gnd.n1143 585
R10137 gnd.n4968 gnd.n1143 585
R10138 gnd.n2762 gnd.n1137 585
R10139 gnd.n2762 gnd.n1068 585
R10140 gnd.n2764 gnd.n2763 585
R10141 gnd.n2766 gnd.n2765 585
R10142 gnd.n2768 gnd.n2767 585
R10143 gnd.n2772 gnd.n2760 585
R10144 gnd.n2774 gnd.n2773 585
R10145 gnd.n2776 gnd.n2775 585
R10146 gnd.n2778 gnd.n2777 585
R10147 gnd.n2782 gnd.n2758 585
R10148 gnd.n2784 gnd.n2783 585
R10149 gnd.n2786 gnd.n2785 585
R10150 gnd.n2788 gnd.n2787 585
R10151 gnd.n2792 gnd.n2756 585
R10152 gnd.n2794 gnd.n2793 585
R10153 gnd.n2796 gnd.n2795 585
R10154 gnd.n2798 gnd.n2797 585
R10155 gnd.n2753 gnd.n2752 585
R10156 gnd.n2802 gnd.n2754 585
R10157 gnd.n2803 gnd.n2749 585
R10158 gnd.n2804 gnd.n1067 585
R10159 gnd.n5092 gnd.n1067 585
R10160 gnd.n3162 gnd.n3161 585
R10161 gnd.n3163 gnd.n2625 585
R10162 gnd.n3164 gnd.n2621 585
R10163 gnd.n2619 gnd.n2610 585
R10164 gnd.n3171 gnd.n2609 585
R10165 gnd.n3172 gnd.n2607 585
R10166 gnd.n2606 gnd.n2599 585
R10167 gnd.n3179 gnd.n2598 585
R10168 gnd.n3180 gnd.n2597 585
R10169 gnd.n2595 gnd.n2587 585
R10170 gnd.n3187 gnd.n2586 585
R10171 gnd.n3188 gnd.n2584 585
R10172 gnd.n2583 gnd.n2576 585
R10173 gnd.n3195 gnd.n2575 585
R10174 gnd.n3196 gnd.n2574 585
R10175 gnd.n2572 gnd.n2564 585
R10176 gnd.n3203 gnd.n2563 585
R10177 gnd.n3204 gnd.n2561 585
R10178 gnd.n2560 gnd.n1372 585
R10179 gnd.n1381 gnd.n1372 585
R10180 gnd.n3146 gnd.n1375 585
R10181 gnd.n4834 gnd.n1375 585
R10182 gnd.n3145 gnd.n3144 585
R10183 gnd.n3144 gnd.n3143 585
R10184 gnd.n2628 gnd.n1366 585
R10185 gnd.n4840 gnd.n1366 585
R10186 gnd.n3135 gnd.n3134 585
R10187 gnd.n3136 gnd.n3135 585
R10188 gnd.n2631 gnd.n1355 585
R10189 gnd.n4846 gnd.n1355 585
R10190 gnd.n3129 gnd.n3128 585
R10191 gnd.n3128 gnd.n3127 585
R10192 gnd.n2633 gnd.n1345 585
R10193 gnd.n4852 gnd.n1345 585
R10194 gnd.n3041 gnd.n2636 585
R10195 gnd.n3121 gnd.n2636 585
R10196 gnd.n3042 gnd.n1335 585
R10197 gnd.n4858 gnd.n1335 585
R10198 gnd.n3043 gnd.n3039 585
R10199 gnd.n3039 gnd.n3038 585
R10200 gnd.n2655 gnd.n1325 585
R10201 gnd.n4864 gnd.n1325 585
R10202 gnd.n3047 gnd.n2654 585
R10203 gnd.n3032 gnd.n2654 585
R10204 gnd.n3048 gnd.n1315 585
R10205 gnd.n4870 gnd.n1315 585
R10206 gnd.n3049 gnd.n2653 585
R10207 gnd.n3026 gnd.n2653 585
R10208 gnd.n2650 gnd.n1305 585
R10209 gnd.n4876 gnd.n1305 585
R10210 gnd.n3054 gnd.n3053 585
R10211 gnd.n3055 gnd.n3054 585
R10212 gnd.n2649 gnd.n1295 585
R10213 gnd.n4882 gnd.n1295 585
R10214 gnd.n3018 gnd.n3017 585
R10215 gnd.n3019 gnd.n3018 585
R10216 gnd.n2658 gnd.n1285 585
R10217 gnd.n4888 gnd.n1285 585
R10218 gnd.n3013 gnd.n3012 585
R10219 gnd.n3012 gnd.n3011 585
R10220 gnd.n2660 gnd.n1276 585
R10221 gnd.n4894 gnd.n1276 585
R10222 gnd.n3003 gnd.n3002 585
R10223 gnd.n3004 gnd.n3003 585
R10224 gnd.n2663 gnd.n1264 585
R10225 gnd.n4900 gnd.n1264 585
R10226 gnd.n2998 gnd.n2997 585
R10227 gnd.n2997 gnd.n2996 585
R10228 gnd.n2666 gnd.n2665 585
R10229 gnd.n2967 gnd.n2666 585
R10230 gnd.n2941 gnd.n2940 585
R10231 gnd.n2940 gnd.n2673 585
R10232 gnd.n2945 gnd.n2681 585
R10233 gnd.n2961 gnd.n2681 585
R10234 gnd.n2947 gnd.n2946 585
R10235 gnd.n2948 gnd.n2947 585
R10236 gnd.n2693 gnd.n2692 585
R10237 gnd.n2931 gnd.n2692 585
R10238 gnd.n2936 gnd.n2935 585
R10239 gnd.n2935 gnd.n2934 585
R10240 gnd.n2696 gnd.n2695 585
R10241 gnd.n2923 gnd.n2696 585
R10242 gnd.n2867 gnd.n2866 585
R10243 gnd.n2866 gnd.n2709 585
R10244 gnd.n2868 gnd.n1247 585
R10245 gnd.n4908 gnd.n1247 585
R10246 gnd.n2874 gnd.n2873 585
R10247 gnd.n2873 gnd.n2872 585
R10248 gnd.n2875 gnd.n1237 585
R10249 gnd.n4914 gnd.n1237 585
R10250 gnd.n2877 gnd.n2876 585
R10251 gnd.n2878 gnd.n2877 585
R10252 gnd.n2740 gnd.n1226 585
R10253 gnd.n4920 gnd.n1226 585
R10254 gnd.n2886 gnd.n2885 585
R10255 gnd.n2885 gnd.n2884 585
R10256 gnd.n2887 gnd.n1216 585
R10257 gnd.n4926 gnd.n1216 585
R10258 gnd.n2889 gnd.n2888 585
R10259 gnd.n2890 gnd.n2889 585
R10260 gnd.n2736 gnd.n1206 585
R10261 gnd.n4932 gnd.n1206 585
R10262 gnd.n2850 gnd.n2849 585
R10263 gnd.n2851 gnd.n2850 585
R10264 gnd.n2742 gnd.n1196 585
R10265 gnd.n4938 gnd.n1196 585
R10266 gnd.n2844 gnd.n2843 585
R10267 gnd.n2843 gnd.n2842 585
R10268 gnd.n2825 gnd.n1186 585
R10269 gnd.n4944 gnd.n1186 585
R10270 gnd.n2824 gnd.n2823 585
R10271 gnd.n2823 gnd.n1177 585
R10272 gnd.n2744 gnd.n1176 585
R10273 gnd.n4950 gnd.n1176 585
R10274 gnd.n2819 gnd.n2818 585
R10275 gnd.n2818 gnd.n1167 585
R10276 gnd.n2817 gnd.n1166 585
R10277 gnd.n4956 gnd.n1166 585
R10278 gnd.n2816 gnd.n2815 585
R10279 gnd.n2815 gnd.n1155 585
R10280 gnd.n2746 gnd.n1154 585
R10281 gnd.n4962 gnd.n1154 585
R10282 gnd.n2811 gnd.n2810 585
R10283 gnd.n2810 gnd.n1152 585
R10284 gnd.n2809 gnd.n1142 585
R10285 gnd.n4968 gnd.n1142 585
R10286 gnd.n2808 gnd.n2807 585
R10287 gnd.n2807 gnd.n1068 585
R10288 gnd.n6476 gnd.n6475 585
R10289 gnd.n6475 gnd.n6474 585
R10290 gnd.n6477 gnd.n1021 585
R10291 gnd.n6384 gnd.n1021 585
R10292 gnd.n6479 gnd.n6478 585
R10293 gnd.n6480 gnd.n6479 585
R10294 gnd.n1022 gnd.n1020 585
R10295 gnd.n1020 gnd.n1016 585
R10296 gnd.n1001 gnd.n1000 585
R10297 gnd.n1005 gnd.n1001 585
R10298 gnd.n6490 gnd.n6489 585
R10299 gnd.n6489 gnd.n6488 585
R10300 gnd.n6491 gnd.n995 585
R10301 gnd.n6373 gnd.n995 585
R10302 gnd.n6493 gnd.n6492 585
R10303 gnd.n6494 gnd.n6493 585
R10304 gnd.n996 gnd.n994 585
R10305 gnd.n994 gnd.n990 585
R10306 gnd.n978 gnd.n977 585
R10307 gnd.n6366 gnd.n978 585
R10308 gnd.n6504 gnd.n6503 585
R10309 gnd.n6503 gnd.n6502 585
R10310 gnd.n6505 gnd.n972 585
R10311 gnd.n6029 gnd.n972 585
R10312 gnd.n6507 gnd.n6506 585
R10313 gnd.n6508 gnd.n6507 585
R10314 gnd.n973 gnd.n971 585
R10315 gnd.n5191 gnd.n971 585
R10316 gnd.n6067 gnd.n6066 585
R10317 gnd.n6066 gnd.n6065 585
R10318 gnd.n5189 gnd.n5188 585
R10319 gnd.n6049 gnd.n5189 585
R10320 gnd.n6041 gnd.n6040 585
R10321 gnd.n6040 gnd.n6039 585
R10322 gnd.n5203 gnd.n5202 585
R10323 gnd.n5211 gnd.n5203 585
R10324 gnd.n6015 gnd.n6014 585
R10325 gnd.n6016 gnd.n6015 585
R10326 gnd.n5214 gnd.n5213 585
R10327 gnd.n5221 gnd.n5213 585
R10328 gnd.n5989 gnd.n5233 585
R10329 gnd.n5233 gnd.n5220 585
R10330 gnd.n5991 gnd.n5990 585
R10331 gnd.n5992 gnd.n5991 585
R10332 gnd.n5234 gnd.n5232 585
R10333 gnd.n5232 gnd.n5228 585
R10334 gnd.n5978 gnd.n5977 585
R10335 gnd.n5977 gnd.n5976 585
R10336 gnd.n5239 gnd.n5238 585
R10337 gnd.n5249 gnd.n5239 585
R10338 gnd.n5967 gnd.n5966 585
R10339 gnd.n5966 gnd.n5965 585
R10340 gnd.n5246 gnd.n5245 585
R10341 gnd.n5953 gnd.n5246 585
R10342 gnd.n5927 gnd.n5331 585
R10343 gnd.n5331 gnd.n5256 585
R10344 gnd.n5929 gnd.n5928 585
R10345 gnd.n5930 gnd.n5929 585
R10346 gnd.n5332 gnd.n5330 585
R10347 gnd.n5340 gnd.n5330 585
R10348 gnd.n5905 gnd.n5352 585
R10349 gnd.n5352 gnd.n5339 585
R10350 gnd.n5907 gnd.n5906 585
R10351 gnd.n5908 gnd.n5907 585
R10352 gnd.n5353 gnd.n5351 585
R10353 gnd.n5351 gnd.n5347 585
R10354 gnd.n5893 gnd.n5892 585
R10355 gnd.n5892 gnd.n5891 585
R10356 gnd.n5358 gnd.n5357 585
R10357 gnd.n5367 gnd.n5358 585
R10358 gnd.n5882 gnd.n5881 585
R10359 gnd.n5881 gnd.n5880 585
R10360 gnd.n5365 gnd.n5364 585
R10361 gnd.n5868 gnd.n5365 585
R10362 gnd.n5840 gnd.n5839 585
R10363 gnd.n5839 gnd.n5374 585
R10364 gnd.n5841 gnd.n5385 585
R10365 gnd.n5832 gnd.n5385 585
R10366 gnd.n5843 gnd.n5842 585
R10367 gnd.n5844 gnd.n5843 585
R10368 gnd.n5386 gnd.n5384 585
R10369 gnd.n5400 gnd.n5384 585
R10370 gnd.n5824 gnd.n5823 585
R10371 gnd.n5823 gnd.n5822 585
R10372 gnd.n5397 gnd.n5396 585
R10373 gnd.n5807 gnd.n5397 585
R10374 gnd.n5794 gnd.n5417 585
R10375 gnd.n5417 gnd.n5407 585
R10376 gnd.n5796 gnd.n5795 585
R10377 gnd.n5797 gnd.n5796 585
R10378 gnd.n5418 gnd.n5416 585
R10379 gnd.n5426 gnd.n5416 585
R10380 gnd.n5770 gnd.n5438 585
R10381 gnd.n5438 gnd.n5425 585
R10382 gnd.n5772 gnd.n5771 585
R10383 gnd.n5773 gnd.n5772 585
R10384 gnd.n5439 gnd.n5437 585
R10385 gnd.n5437 gnd.n5433 585
R10386 gnd.n5758 gnd.n5757 585
R10387 gnd.n5757 gnd.n5756 585
R10388 gnd.n5444 gnd.n5443 585
R10389 gnd.n5448 gnd.n5444 585
R10390 gnd.n5742 gnd.n5741 585
R10391 gnd.n5743 gnd.n5742 585
R10392 gnd.n5459 gnd.n5458 585
R10393 gnd.n5458 gnd.n5454 585
R10394 gnd.n5732 gnd.n5731 585
R10395 gnd.n5733 gnd.n5732 585
R10396 gnd.n5468 gnd.n5467 585
R10397 gnd.n5467 gnd.n5465 585
R10398 gnd.n5726 gnd.n5725 585
R10399 gnd.n5725 gnd.n5724 585
R10400 gnd.n5472 gnd.n5471 585
R10401 gnd.n5480 gnd.n5472 585
R10402 gnd.n5633 gnd.n5632 585
R10403 gnd.n5634 gnd.n5633 585
R10404 gnd.n5482 gnd.n5481 585
R10405 gnd.n5481 gnd.n5479 585
R10406 gnd.n5628 gnd.n5627 585
R10407 gnd.n5627 gnd.n5626 585
R10408 gnd.n5485 gnd.n5484 585
R10409 gnd.n5486 gnd.n5485 585
R10410 gnd.n5617 gnd.n5616 585
R10411 gnd.n5618 gnd.n5617 585
R10412 gnd.n5494 gnd.n5493 585
R10413 gnd.n5493 gnd.n5492 585
R10414 gnd.n5612 gnd.n5611 585
R10415 gnd.n5611 gnd.n5610 585
R10416 gnd.n5497 gnd.n5496 585
R10417 gnd.n5498 gnd.n5497 585
R10418 gnd.n5601 gnd.n5600 585
R10419 gnd.n5602 gnd.n5601 585
R10420 gnd.n5597 gnd.n5504 585
R10421 gnd.n5596 gnd.n5595 585
R10422 gnd.n5593 gnd.n5506 585
R10423 gnd.n5593 gnd.n5503 585
R10424 gnd.n5592 gnd.n5591 585
R10425 gnd.n5590 gnd.n5589 585
R10426 gnd.n5588 gnd.n5511 585
R10427 gnd.n5586 gnd.n5585 585
R10428 gnd.n5584 gnd.n5512 585
R10429 gnd.n5583 gnd.n5582 585
R10430 gnd.n5580 gnd.n5517 585
R10431 gnd.n5578 gnd.n5577 585
R10432 gnd.n5576 gnd.n5518 585
R10433 gnd.n5575 gnd.n5574 585
R10434 gnd.n5572 gnd.n5523 585
R10435 gnd.n5570 gnd.n5569 585
R10436 gnd.n5568 gnd.n5524 585
R10437 gnd.n5567 gnd.n5566 585
R10438 gnd.n5564 gnd.n5529 585
R10439 gnd.n5562 gnd.n5561 585
R10440 gnd.n5560 gnd.n5530 585
R10441 gnd.n5559 gnd.n5558 585
R10442 gnd.n5556 gnd.n5535 585
R10443 gnd.n5554 gnd.n5553 585
R10444 gnd.n5551 gnd.n5536 585
R10445 gnd.n5550 gnd.n5549 585
R10446 gnd.n5547 gnd.n5545 585
R10447 gnd.n5543 gnd.n5502 585
R10448 gnd.n6392 gnd.n6391 585
R10449 gnd.n6393 gnd.n5172 585
R10450 gnd.n6395 gnd.n6394 585
R10451 gnd.n6397 gnd.n5171 585
R10452 gnd.n6399 gnd.n6398 585
R10453 gnd.n6400 gnd.n5162 585
R10454 gnd.n6402 gnd.n6401 585
R10455 gnd.n6404 gnd.n5160 585
R10456 gnd.n6406 gnd.n6405 585
R10457 gnd.n6407 gnd.n5155 585
R10458 gnd.n6409 gnd.n6408 585
R10459 gnd.n6411 gnd.n5153 585
R10460 gnd.n6413 gnd.n6412 585
R10461 gnd.n6414 gnd.n5148 585
R10462 gnd.n6416 gnd.n6415 585
R10463 gnd.n6418 gnd.n5146 585
R10464 gnd.n6420 gnd.n6419 585
R10465 gnd.n6421 gnd.n5141 585
R10466 gnd.n6423 gnd.n6422 585
R10467 gnd.n6425 gnd.n5139 585
R10468 gnd.n6427 gnd.n6426 585
R10469 gnd.n6428 gnd.n5134 585
R10470 gnd.n6430 gnd.n6429 585
R10471 gnd.n6432 gnd.n5132 585
R10472 gnd.n6434 gnd.n6433 585
R10473 gnd.n6435 gnd.n5130 585
R10474 gnd.n6436 gnd.n1026 585
R10475 gnd.n5093 gnd.n1026 585
R10476 gnd.n6387 gnd.n1028 585
R10477 gnd.n6474 gnd.n1028 585
R10478 gnd.n6386 gnd.n6385 585
R10479 gnd.n6385 gnd.n6384 585
R10480 gnd.n6383 gnd.n1018 585
R10481 gnd.n6480 gnd.n1018 585
R10482 gnd.n6377 gnd.n5177 585
R10483 gnd.n6377 gnd.n1016 585
R10484 gnd.n6379 gnd.n6378 585
R10485 gnd.n6378 gnd.n1005 585
R10486 gnd.n6376 gnd.n1003 585
R10487 gnd.n6488 gnd.n1003 585
R10488 gnd.n6375 gnd.n6374 585
R10489 gnd.n6374 gnd.n6373 585
R10490 gnd.n5179 gnd.n992 585
R10491 gnd.n6494 gnd.n992 585
R10492 gnd.n6369 gnd.n6368 585
R10493 gnd.n6368 gnd.n990 585
R10494 gnd.n6367 gnd.n5181 585
R10495 gnd.n6367 gnd.n6366 585
R10496 gnd.n6028 gnd.n980 585
R10497 gnd.n6502 gnd.n980 585
R10498 gnd.n6031 gnd.n6030 585
R10499 gnd.n6030 gnd.n6029 585
R10500 gnd.n6032 gnd.n969 585
R10501 gnd.n6508 gnd.n969 585
R10502 gnd.n6034 gnd.n6033 585
R10503 gnd.n6033 gnd.n5191 585
R10504 gnd.n6035 gnd.n5190 585
R10505 gnd.n6065 gnd.n5190 585
R10506 gnd.n6036 gnd.n5199 585
R10507 gnd.n6049 gnd.n5199 585
R10508 gnd.n6038 gnd.n6037 585
R10509 gnd.n6039 gnd.n6038 585
R10510 gnd.n5206 gnd.n5205 585
R10511 gnd.n5211 gnd.n5205 585
R10512 gnd.n6018 gnd.n6017 585
R10513 gnd.n6017 gnd.n6016 585
R10514 gnd.n5209 gnd.n5208 585
R10515 gnd.n5221 gnd.n5209 585
R10516 gnd.n5943 gnd.n5942 585
R10517 gnd.n5942 gnd.n5220 585
R10518 gnd.n5944 gnd.n5230 585
R10519 gnd.n5992 gnd.n5230 585
R10520 gnd.n5946 gnd.n5945 585
R10521 gnd.n5945 gnd.n5228 585
R10522 gnd.n5947 gnd.n5241 585
R10523 gnd.n5976 gnd.n5241 585
R10524 gnd.n5949 gnd.n5948 585
R10525 gnd.n5948 gnd.n5249 585
R10526 gnd.n5950 gnd.n5248 585
R10527 gnd.n5965 gnd.n5248 585
R10528 gnd.n5952 gnd.n5951 585
R10529 gnd.n5953 gnd.n5952 585
R10530 gnd.n5260 gnd.n5259 585
R10531 gnd.n5259 gnd.n5256 585
R10532 gnd.n5932 gnd.n5931 585
R10533 gnd.n5931 gnd.n5930 585
R10534 gnd.n5327 gnd.n5326 585
R10535 gnd.n5340 gnd.n5327 585
R10536 gnd.n5853 gnd.n5852 585
R10537 gnd.n5852 gnd.n5339 585
R10538 gnd.n5854 gnd.n5349 585
R10539 gnd.n5908 gnd.n5349 585
R10540 gnd.n5857 gnd.n5856 585
R10541 gnd.n5856 gnd.n5347 585
R10542 gnd.n5858 gnd.n5360 585
R10543 gnd.n5891 gnd.n5360 585
R10544 gnd.n5861 gnd.n5860 585
R10545 gnd.n5860 gnd.n5367 585
R10546 gnd.n5862 gnd.n5366 585
R10547 gnd.n5880 gnd.n5366 585
R10548 gnd.n5865 gnd.n5864 585
R10549 gnd.n5868 gnd.n5865 585
R10550 gnd.n5850 gnd.n5376 585
R10551 gnd.n5376 gnd.n5374 585
R10552 gnd.n5381 gnd.n5377 585
R10553 gnd.n5832 gnd.n5381 585
R10554 gnd.n5846 gnd.n5845 585
R10555 gnd.n5845 gnd.n5844 585
R10556 gnd.n5380 gnd.n5379 585
R10557 gnd.n5400 gnd.n5380 585
R10558 gnd.n5804 gnd.n5399 585
R10559 gnd.n5822 gnd.n5399 585
R10560 gnd.n5806 gnd.n5805 585
R10561 gnd.n5807 gnd.n5806 585
R10562 gnd.n5410 gnd.n5409 585
R10563 gnd.n5409 gnd.n5407 585
R10564 gnd.n5799 gnd.n5798 585
R10565 gnd.n5798 gnd.n5797 585
R10566 gnd.n5413 gnd.n5412 585
R10567 gnd.n5426 gnd.n5413 585
R10568 gnd.n5650 gnd.n5649 585
R10569 gnd.n5649 gnd.n5425 585
R10570 gnd.n5651 gnd.n5435 585
R10571 gnd.n5773 gnd.n5435 585
R10572 gnd.n5653 gnd.n5652 585
R10573 gnd.n5652 gnd.n5433 585
R10574 gnd.n5654 gnd.n5445 585
R10575 gnd.n5756 gnd.n5445 585
R10576 gnd.n5656 gnd.n5655 585
R10577 gnd.n5655 gnd.n5448 585
R10578 gnd.n5657 gnd.n5456 585
R10579 gnd.n5743 gnd.n5456 585
R10580 gnd.n5659 gnd.n5658 585
R10581 gnd.n5658 gnd.n5454 585
R10582 gnd.n5660 gnd.n5466 585
R10583 gnd.n5733 gnd.n5466 585
R10584 gnd.n5661 gnd.n5474 585
R10585 gnd.n5474 gnd.n5465 585
R10586 gnd.n5663 gnd.n5662 585
R10587 gnd.n5724 gnd.n5663 585
R10588 gnd.n5475 gnd.n5473 585
R10589 gnd.n5480 gnd.n5473 585
R10590 gnd.n5636 gnd.n5635 585
R10591 gnd.n5635 gnd.n5634 585
R10592 gnd.n5478 gnd.n5477 585
R10593 gnd.n5479 gnd.n5478 585
R10594 gnd.n5625 gnd.n5624 585
R10595 gnd.n5626 gnd.n5625 585
R10596 gnd.n5488 gnd.n5487 585
R10597 gnd.n5487 gnd.n5486 585
R10598 gnd.n5620 gnd.n5619 585
R10599 gnd.n5619 gnd.n5618 585
R10600 gnd.n5491 gnd.n5490 585
R10601 gnd.n5492 gnd.n5491 585
R10602 gnd.n5609 gnd.n5608 585
R10603 gnd.n5610 gnd.n5609 585
R10604 gnd.n5500 gnd.n5499 585
R10605 gnd.n5499 gnd.n5498 585
R10606 gnd.n5604 gnd.n5603 585
R10607 gnd.n5603 gnd.n5602 585
R10608 gnd.n7605 gnd.n7604 585
R10609 gnd.n7604 gnd.n7603 585
R10610 gnd.n7606 gnd.n204 585
R10611 gnd.n209 gnd.n204 585
R10612 gnd.n7608 gnd.n7607 585
R10613 gnd.n7609 gnd.n7608 585
R10614 gnd.n191 gnd.n190 585
R10615 gnd.n194 gnd.n191 585
R10616 gnd.n7617 gnd.n7616 585
R10617 gnd.n7616 gnd.n7615 585
R10618 gnd.n7618 gnd.n186 585
R10619 gnd.n186 gnd.n185 585
R10620 gnd.n7620 gnd.n7619 585
R10621 gnd.n7621 gnd.n7620 585
R10622 gnd.n171 gnd.n170 585
R10623 gnd.n175 gnd.n171 585
R10624 gnd.n7629 gnd.n7628 585
R10625 gnd.n7628 gnd.n7627 585
R10626 gnd.n7630 gnd.n166 585
R10627 gnd.n7438 gnd.n166 585
R10628 gnd.n7632 gnd.n7631 585
R10629 gnd.n7633 gnd.n7632 585
R10630 gnd.n152 gnd.n151 585
R10631 gnd.n7417 gnd.n152 585
R10632 gnd.n7641 gnd.n7640 585
R10633 gnd.n7640 gnd.n7639 585
R10634 gnd.n7642 gnd.n147 585
R10635 gnd.n7408 gnd.n147 585
R10636 gnd.n7644 gnd.n7643 585
R10637 gnd.n7645 gnd.n7644 585
R10638 gnd.n131 gnd.n130 585
R10639 gnd.n7402 gnd.n131 585
R10640 gnd.n7653 gnd.n7652 585
R10641 gnd.n7652 gnd.n7651 585
R10642 gnd.n7654 gnd.n126 585
R10643 gnd.n7394 gnd.n126 585
R10644 gnd.n7656 gnd.n7655 585
R10645 gnd.n7657 gnd.n7656 585
R10646 gnd.n113 gnd.n112 585
R10647 gnd.n7388 gnd.n113 585
R10648 gnd.n7665 gnd.n7664 585
R10649 gnd.n7664 gnd.n7663 585
R10650 gnd.n7666 gnd.n107 585
R10651 gnd.n7380 gnd.n107 585
R10652 gnd.n7668 gnd.n7667 585
R10653 gnd.n7669 gnd.n7668 585
R10654 gnd.n108 gnd.n106 585
R10655 gnd.n7374 gnd.n106 585
R10656 gnd.n4301 gnd.n4300 585
R10657 gnd.n4300 gnd.n381 585
R10658 gnd.n1935 gnd.n88 585
R10659 gnd.n7677 gnd.n88 585
R10660 gnd.n4309 gnd.n4308 585
R10661 gnd.n4308 gnd.n4307 585
R10662 gnd.n4310 gnd.n1925 585
R10663 gnd.n4318 gnd.n1925 585
R10664 gnd.n4312 gnd.n4311 585
R10665 gnd.n4313 gnd.n4312 585
R10666 gnd.n1931 gnd.n1930 585
R10667 gnd.n1930 gnd.n1912 585
R10668 gnd.n1903 gnd.n1902 585
R10669 gnd.n4327 gnd.n1903 585
R10670 gnd.n4333 gnd.n4332 585
R10671 gnd.n4332 gnd.n4331 585
R10672 gnd.n4334 gnd.n1898 585
R10673 gnd.n4289 gnd.n1898 585
R10674 gnd.n4336 gnd.n4335 585
R10675 gnd.n4337 gnd.n4336 585
R10676 gnd.n1883 gnd.n1882 585
R10677 gnd.n4273 gnd.n1883 585
R10678 gnd.n4345 gnd.n4344 585
R10679 gnd.n4344 gnd.n4343 585
R10680 gnd.n4346 gnd.n1878 585
R10681 gnd.n4234 gnd.n1878 585
R10682 gnd.n4348 gnd.n4347 585
R10683 gnd.n4349 gnd.n4348 585
R10684 gnd.n1863 gnd.n1862 585
R10685 gnd.n4225 gnd.n1863 585
R10686 gnd.n4357 gnd.n4356 585
R10687 gnd.n4356 gnd.n4355 585
R10688 gnd.n4358 gnd.n1858 585
R10689 gnd.n4219 gnd.n1858 585
R10690 gnd.n4360 gnd.n4359 585
R10691 gnd.n4361 gnd.n4360 585
R10692 gnd.n1843 gnd.n1842 585
R10693 gnd.n4248 gnd.n1843 585
R10694 gnd.n4369 gnd.n4368 585
R10695 gnd.n4368 gnd.n4367 585
R10696 gnd.n4370 gnd.n1838 585
R10697 gnd.n4212 gnd.n1838 585
R10698 gnd.n4372 gnd.n4371 585
R10699 gnd.n4373 gnd.n4372 585
R10700 gnd.n1823 gnd.n1822 585
R10701 gnd.n4204 gnd.n1823 585
R10702 gnd.n4381 gnd.n4380 585
R10703 gnd.n4380 gnd.n4379 585
R10704 gnd.n4382 gnd.n1816 585
R10705 gnd.n4197 gnd.n1816 585
R10706 gnd.n4384 gnd.n4383 585
R10707 gnd.n4385 gnd.n4384 585
R10708 gnd.n1817 gnd.n1815 585
R10709 gnd.n4189 gnd.n1815 585
R10710 gnd.n1799 gnd.n1792 585
R10711 gnd.n4391 gnd.n1799 585
R10712 gnd.n4396 gnd.n1790 585
R10713 gnd.n1970 gnd.n1790 585
R10714 gnd.n4398 gnd.n4397 585
R10715 gnd.n4399 gnd.n4398 585
R10716 gnd.n1789 gnd.n1629 585
R10717 gnd.n4566 gnd.n1630 585
R10718 gnd.n4565 gnd.n1631 585
R10719 gnd.n1706 gnd.n1632 585
R10720 gnd.n4558 gnd.n1638 585
R10721 gnd.n4557 gnd.n1639 585
R10722 gnd.n1709 gnd.n1640 585
R10723 gnd.n4550 gnd.n1646 585
R10724 gnd.n4549 gnd.n1647 585
R10725 gnd.n1711 gnd.n1648 585
R10726 gnd.n4542 gnd.n1654 585
R10727 gnd.n4541 gnd.n1655 585
R10728 gnd.n1714 gnd.n1656 585
R10729 gnd.n4534 gnd.n1662 585
R10730 gnd.n4533 gnd.n1663 585
R10731 gnd.n1716 gnd.n1664 585
R10732 gnd.n4526 gnd.n1672 585
R10733 gnd.n4525 gnd.n4522 585
R10734 gnd.n1675 gnd.n1673 585
R10735 gnd.n4520 gnd.n1675 585
R10736 gnd.n349 gnd.n348 585
R10737 gnd.n7459 gnd.n344 585
R10738 gnd.n7461 gnd.n7460 585
R10739 gnd.n7463 gnd.n342 585
R10740 gnd.n7465 gnd.n7464 585
R10741 gnd.n7466 gnd.n337 585
R10742 gnd.n7468 gnd.n7467 585
R10743 gnd.n7470 gnd.n335 585
R10744 gnd.n7472 gnd.n7471 585
R10745 gnd.n7473 gnd.n330 585
R10746 gnd.n7475 gnd.n7474 585
R10747 gnd.n7477 gnd.n328 585
R10748 gnd.n7479 gnd.n7478 585
R10749 gnd.n7480 gnd.n323 585
R10750 gnd.n7482 gnd.n7481 585
R10751 gnd.n7484 gnd.n321 585
R10752 gnd.n7486 gnd.n7485 585
R10753 gnd.n7487 gnd.n319 585
R10754 gnd.n7488 gnd.n208 585
R10755 gnd.n212 gnd.n208 585
R10756 gnd.n7455 gnd.n211 585
R10757 gnd.n7603 gnd.n211 585
R10758 gnd.n7454 gnd.n7453 585
R10759 gnd.n7453 gnd.n209 585
R10760 gnd.n7452 gnd.n203 585
R10761 gnd.n7609 gnd.n203 585
R10762 gnd.n354 gnd.n353 585
R10763 gnd.n353 gnd.n194 585
R10764 gnd.n7448 gnd.n193 585
R10765 gnd.n7615 gnd.n193 585
R10766 gnd.n7447 gnd.n7446 585
R10767 gnd.n7446 gnd.n185 585
R10768 gnd.n7445 gnd.n184 585
R10769 gnd.n7621 gnd.n184 585
R10770 gnd.n357 gnd.n356 585
R10771 gnd.n356 gnd.n175 585
R10772 gnd.n7441 gnd.n174 585
R10773 gnd.n7627 gnd.n174 585
R10774 gnd.n7440 gnd.n7439 585
R10775 gnd.n7439 gnd.n7438 585
R10776 gnd.n359 gnd.n165 585
R10777 gnd.n7633 gnd.n165 585
R10778 gnd.n7416 gnd.n7415 585
R10779 gnd.n7417 gnd.n7416 585
R10780 gnd.n363 gnd.n155 585
R10781 gnd.n7639 gnd.n155 585
R10782 gnd.n7410 gnd.n7409 585
R10783 gnd.n7409 gnd.n7408 585
R10784 gnd.n365 gnd.n145 585
R10785 gnd.n7645 gnd.n145 585
R10786 gnd.n7401 gnd.n7400 585
R10787 gnd.n7402 gnd.n7401 585
R10788 gnd.n368 gnd.n134 585
R10789 gnd.n7651 gnd.n134 585
R10790 gnd.n7396 gnd.n7395 585
R10791 gnd.n7395 gnd.n7394 585
R10792 gnd.n370 gnd.n125 585
R10793 gnd.n7657 gnd.n125 585
R10794 gnd.n7387 gnd.n7386 585
R10795 gnd.n7388 gnd.n7387 585
R10796 gnd.n375 gnd.n116 585
R10797 gnd.n7663 gnd.n116 585
R10798 gnd.n7382 gnd.n7381 585
R10799 gnd.n7381 gnd.n7380 585
R10800 gnd.n377 gnd.n104 585
R10801 gnd.n7669 gnd.n104 585
R10802 gnd.n7373 gnd.n7372 585
R10803 gnd.n7374 gnd.n7373 585
R10804 gnd.n84 gnd.n83 585
R10805 gnd.n381 gnd.n84 585
R10806 gnd.n7679 gnd.n7678 585
R10807 gnd.n7678 gnd.n7677 585
R10808 gnd.n7680 gnd.n82 585
R10809 gnd.n4307 gnd.n82 585
R10810 gnd.n1923 gnd.n81 585
R10811 gnd.n4318 gnd.n1923 585
R10812 gnd.n4281 gnd.n1929 585
R10813 gnd.n4313 gnd.n1929 585
R10814 gnd.n4282 gnd.n4279 585
R10815 gnd.n4279 gnd.n1912 585
R10816 gnd.n4283 gnd.n1911 585
R10817 gnd.n4327 gnd.n1911 585
R10818 gnd.n1938 gnd.n1906 585
R10819 gnd.n4331 gnd.n1906 585
R10820 gnd.n4288 gnd.n4287 585
R10821 gnd.n4289 gnd.n4288 585
R10822 gnd.n1937 gnd.n1896 585
R10823 gnd.n4337 gnd.n1896 585
R10824 gnd.n4275 gnd.n4274 585
R10825 gnd.n4274 gnd.n4273 585
R10826 gnd.n1940 gnd.n1886 585
R10827 gnd.n4343 gnd.n1886 585
R10828 gnd.n4236 gnd.n4235 585
R10829 gnd.n4235 gnd.n4234 585
R10830 gnd.n1960 gnd.n1876 585
R10831 gnd.n4349 gnd.n1876 585
R10832 gnd.n4240 gnd.n1959 585
R10833 gnd.n4225 gnd.n1959 585
R10834 gnd.n4241 gnd.n1866 585
R10835 gnd.n4355 gnd.n1866 585
R10836 gnd.n4242 gnd.n1958 585
R10837 gnd.n4219 gnd.n1958 585
R10838 gnd.n1955 gnd.n1856 585
R10839 gnd.n4361 gnd.n1856 585
R10840 gnd.n4247 gnd.n4246 585
R10841 gnd.n4248 gnd.n4247 585
R10842 gnd.n1954 gnd.n1846 585
R10843 gnd.n4367 gnd.n1846 585
R10844 gnd.n4211 gnd.n4210 585
R10845 gnd.n4212 gnd.n4211 585
R10846 gnd.n1962 gnd.n1836 585
R10847 gnd.n4373 gnd.n1836 585
R10848 gnd.n4206 gnd.n4205 585
R10849 gnd.n4205 gnd.n4204 585
R10850 gnd.n1964 gnd.n1826 585
R10851 gnd.n4379 gnd.n1826 585
R10852 gnd.n4196 gnd.n4195 585
R10853 gnd.n4197 gnd.n4196 585
R10854 gnd.n1967 gnd.n1813 585
R10855 gnd.n4385 gnd.n1813 585
R10856 gnd.n4191 gnd.n4190 585
R10857 gnd.n4190 gnd.n4189 585
R10858 gnd.n4188 gnd.n1797 585
R10859 gnd.n4391 gnd.n1797 585
R10860 gnd.n4187 gnd.n1971 585
R10861 gnd.n1971 gnd.n1970 585
R10862 gnd.n1969 gnd.n1787 585
R10863 gnd.n4399 gnd.n1787 585
R10864 gnd.n6472 gnd.n6471 585
R10865 gnd.n6473 gnd.n6472 585
R10866 gnd.n5096 gnd.n5094 585
R10867 gnd.n5094 gnd.n1027 585
R10868 gnd.n1015 gnd.n1014 585
R10869 gnd.n1019 gnd.n1015 585
R10870 gnd.n6483 gnd.n6482 585
R10871 gnd.n6482 gnd.n6481 585
R10872 gnd.n6484 gnd.n1007 585
R10873 gnd.n6354 gnd.n1007 585
R10874 gnd.n6486 gnd.n6485 585
R10875 gnd.n6487 gnd.n6486 585
R10876 gnd.n1008 gnd.n1006 585
R10877 gnd.n1006 gnd.n1002 585
R10878 gnd.n989 gnd.n988 585
R10879 gnd.n993 gnd.n989 585
R10880 gnd.n6497 gnd.n6496 585
R10881 gnd.n6496 gnd.n6495 585
R10882 gnd.n6498 gnd.n983 585
R10883 gnd.n6365 gnd.n983 585
R10884 gnd.n6500 gnd.n6499 585
R10885 gnd.n6501 gnd.n6500 585
R10886 gnd.n984 gnd.n982 585
R10887 gnd.n982 gnd.n979 585
R10888 gnd.n6060 gnd.n6059 585
R10889 gnd.n6059 gnd.n970 585
R10890 gnd.n6061 gnd.n5193 585
R10891 gnd.n5193 gnd.n968 585
R10892 gnd.n6063 gnd.n6062 585
R10893 gnd.n6064 gnd.n6063 585
R10894 gnd.n5194 gnd.n5192 585
R10895 gnd.n6048 gnd.n5192 585
R10896 gnd.n6052 gnd.n6051 585
R10897 gnd.n6051 gnd.n6050 585
R10898 gnd.n5197 gnd.n5196 585
R10899 gnd.n5204 gnd.n5197 585
R10900 gnd.n6002 gnd.n6001 585
R10901 gnd.n6001 gnd.n5212 585
R10902 gnd.n6003 gnd.n5223 585
R10903 gnd.n5223 gnd.n5210 585
R10904 gnd.n6005 gnd.n6004 585
R10905 gnd.n6006 gnd.n6005 585
R10906 gnd.n5224 gnd.n5222 585
R10907 gnd.n5231 gnd.n5222 585
R10908 gnd.n5995 gnd.n5994 585
R10909 gnd.n5994 gnd.n5993 585
R10910 gnd.n5227 gnd.n5226 585
R10911 gnd.n5975 gnd.n5227 585
R10912 gnd.n5961 gnd.n5251 585
R10913 gnd.n5251 gnd.n5240 585
R10914 gnd.n5963 gnd.n5962 585
R10915 gnd.n5964 gnd.n5963 585
R10916 gnd.n5252 gnd.n5250 585
R10917 gnd.n5250 gnd.n5247 585
R10918 gnd.n5956 gnd.n5955 585
R10919 gnd.n5955 gnd.n5954 585
R10920 gnd.n5255 gnd.n5254 585
R10921 gnd.n5329 gnd.n5255 585
R10922 gnd.n5916 gnd.n5342 585
R10923 gnd.n5342 gnd.n5328 585
R10924 gnd.n5918 gnd.n5917 585
R10925 gnd.n5919 gnd.n5918 585
R10926 gnd.n5343 gnd.n5341 585
R10927 gnd.n5350 gnd.n5341 585
R10928 gnd.n5911 gnd.n5910 585
R10929 gnd.n5910 gnd.n5909 585
R10930 gnd.n5346 gnd.n5345 585
R10931 gnd.n5890 gnd.n5346 585
R10932 gnd.n5876 gnd.n5369 585
R10933 gnd.n5369 gnd.n5359 585
R10934 gnd.n5878 gnd.n5877 585
R10935 gnd.n5879 gnd.n5878 585
R10936 gnd.n5370 gnd.n5368 585
R10937 gnd.n5867 gnd.n5368 585
R10938 gnd.n5871 gnd.n5870 585
R10939 gnd.n5870 gnd.n5869 585
R10940 gnd.n5373 gnd.n5372 585
R10941 gnd.n5833 gnd.n5373 585
R10942 gnd.n5817 gnd.n5816 585
R10943 gnd.n5816 gnd.n5383 585
R10944 gnd.n5818 gnd.n5402 585
R10945 gnd.n5402 gnd.n5382 585
R10946 gnd.n5820 gnd.n5819 585
R10947 gnd.n5821 gnd.n5820 585
R10948 gnd.n5403 gnd.n5401 585
R10949 gnd.n5401 gnd.n5398 585
R10950 gnd.n5810 gnd.n5809 585
R10951 gnd.n5809 gnd.n5808 585
R10952 gnd.n5406 gnd.n5405 585
R10953 gnd.n5415 gnd.n5406 585
R10954 gnd.n5781 gnd.n5428 585
R10955 gnd.n5428 gnd.n5414 585
R10956 gnd.n5783 gnd.n5782 585
R10957 gnd.n5784 gnd.n5783 585
R10958 gnd.n5429 gnd.n5427 585
R10959 gnd.n5436 gnd.n5427 585
R10960 gnd.n5776 gnd.n5775 585
R10961 gnd.n5775 gnd.n5774 585
R10962 gnd.n5432 gnd.n5431 585
R10963 gnd.n5755 gnd.n5432 585
R10964 gnd.n5751 gnd.n5750 585
R10965 gnd.n5752 gnd.n5751 585
R10966 gnd.n5450 gnd.n5449 585
R10967 gnd.n5457 gnd.n5449 585
R10968 gnd.n5746 gnd.n5745 585
R10969 gnd.n5745 gnd.n5744 585
R10970 gnd.n5453 gnd.n5452 585
R10971 gnd.n5734 gnd.n5453 585
R10972 gnd.n5721 gnd.n5720 585
R10973 gnd.n5719 gnd.n5672 585
R10974 gnd.n5718 gnd.n5671 585
R10975 gnd.n5723 gnd.n5671 585
R10976 gnd.n5717 gnd.n5716 585
R10977 gnd.n5715 gnd.n5714 585
R10978 gnd.n5713 gnd.n5712 585
R10979 gnd.n5711 gnd.n5710 585
R10980 gnd.n5709 gnd.n5708 585
R10981 gnd.n5707 gnd.n5706 585
R10982 gnd.n5705 gnd.n5704 585
R10983 gnd.n5703 gnd.n5702 585
R10984 gnd.n5701 gnd.n5700 585
R10985 gnd.n5699 gnd.n5698 585
R10986 gnd.n5697 gnd.n5696 585
R10987 gnd.n5695 gnd.n5694 585
R10988 gnd.n5693 gnd.n5692 585
R10989 gnd.n5688 gnd.n5464 585
R10990 gnd.n6441 gnd.n6440 585
R10991 gnd.n6443 gnd.n5125 585
R10992 gnd.n6445 gnd.n6444 585
R10993 gnd.n6446 gnd.n5118 585
R10994 gnd.n6448 gnd.n6447 585
R10995 gnd.n6450 gnd.n5116 585
R10996 gnd.n6452 gnd.n6451 585
R10997 gnd.n6453 gnd.n5111 585
R10998 gnd.n6455 gnd.n6454 585
R10999 gnd.n6457 gnd.n5109 585
R11000 gnd.n6459 gnd.n6458 585
R11001 gnd.n6460 gnd.n5104 585
R11002 gnd.n6462 gnd.n6461 585
R11003 gnd.n6464 gnd.n5102 585
R11004 gnd.n6466 gnd.n6465 585
R11005 gnd.n6467 gnd.n5100 585
R11006 gnd.n6468 gnd.n5095 585
R11007 gnd.n5095 gnd.n5093 585
R11008 gnd.n6348 gnd.n1029 585
R11009 gnd.n6473 gnd.n1029 585
R11010 gnd.n6350 gnd.n6349 585
R11011 gnd.n6350 gnd.n1027 585
R11012 gnd.n6352 gnd.n6351 585
R11013 gnd.n6351 gnd.n1019 585
R11014 gnd.n6353 gnd.n1017 585
R11015 gnd.n6481 gnd.n1017 585
R11016 gnd.n6356 gnd.n6355 585
R11017 gnd.n6355 gnd.n6354 585
R11018 gnd.n6357 gnd.n1004 585
R11019 gnd.n6487 gnd.n1004 585
R11020 gnd.n6359 gnd.n6358 585
R11021 gnd.n6359 gnd.n1002 585
R11022 gnd.n6361 gnd.n6360 585
R11023 gnd.n6360 gnd.n993 585
R11024 gnd.n6362 gnd.n991 585
R11025 gnd.n6495 gnd.n991 585
R11026 gnd.n6364 gnd.n6363 585
R11027 gnd.n6365 gnd.n6364 585
R11028 gnd.n6077 gnd.n981 585
R11029 gnd.n6501 gnd.n981 585
R11030 gnd.n6076 gnd.n6075 585
R11031 gnd.n6075 gnd.n979 585
R11032 gnd.n6074 gnd.n5183 585
R11033 gnd.n6074 gnd.n970 585
R11034 gnd.n6073 gnd.n6072 585
R11035 gnd.n6073 gnd.n968 585
R11036 gnd.n5186 gnd.n5185 585
R11037 gnd.n6064 gnd.n5185 585
R11038 gnd.n6047 gnd.n6046 585
R11039 gnd.n6048 gnd.n6047 585
R11040 gnd.n6045 gnd.n5198 585
R11041 gnd.n6050 gnd.n5198 585
R11042 gnd.n6009 gnd.n5200 585
R11043 gnd.n6009 gnd.n5204 585
R11044 gnd.n6011 gnd.n6010 585
R11045 gnd.n6010 gnd.n5212 585
R11046 gnd.n6008 gnd.n5217 585
R11047 gnd.n6008 gnd.n5210 585
R11048 gnd.n6007 gnd.n5219 585
R11049 gnd.n6007 gnd.n6006 585
R11050 gnd.n5984 gnd.n5218 585
R11051 gnd.n5231 gnd.n5218 585
R11052 gnd.n5983 gnd.n5229 585
R11053 gnd.n5993 gnd.n5229 585
R11054 gnd.n5974 gnd.n5236 585
R11055 gnd.n5975 gnd.n5974 585
R11056 gnd.n5973 gnd.n5972 585
R11057 gnd.n5973 gnd.n5240 585
R11058 gnd.n5971 gnd.n5242 585
R11059 gnd.n5964 gnd.n5242 585
R11060 gnd.n5257 gnd.n5243 585
R11061 gnd.n5257 gnd.n5247 585
R11062 gnd.n5924 gnd.n5258 585
R11063 gnd.n5954 gnd.n5258 585
R11064 gnd.n5923 gnd.n5922 585
R11065 gnd.n5922 gnd.n5329 585
R11066 gnd.n5921 gnd.n5336 585
R11067 gnd.n5921 gnd.n5328 585
R11068 gnd.n5920 gnd.n5338 585
R11069 gnd.n5920 gnd.n5919 585
R11070 gnd.n5899 gnd.n5337 585
R11071 gnd.n5350 gnd.n5337 585
R11072 gnd.n5898 gnd.n5348 585
R11073 gnd.n5909 gnd.n5348 585
R11074 gnd.n5889 gnd.n5355 585
R11075 gnd.n5890 gnd.n5889 585
R11076 gnd.n5888 gnd.n5887 585
R11077 gnd.n5888 gnd.n5359 585
R11078 gnd.n5886 gnd.n5361 585
R11079 gnd.n5879 gnd.n5361 585
R11080 gnd.n5866 gnd.n5362 585
R11081 gnd.n5867 gnd.n5866 585
R11082 gnd.n5836 gnd.n5375 585
R11083 gnd.n5869 gnd.n5375 585
R11084 gnd.n5835 gnd.n5834 585
R11085 gnd.n5834 gnd.n5833 585
R11086 gnd.n5831 gnd.n5392 585
R11087 gnd.n5831 gnd.n5383 585
R11088 gnd.n5830 gnd.n5829 585
R11089 gnd.n5830 gnd.n5382 585
R11090 gnd.n5394 gnd.n5393 585
R11091 gnd.n5821 gnd.n5393 585
R11092 gnd.n5790 gnd.n5789 585
R11093 gnd.n5789 gnd.n5398 585
R11094 gnd.n5791 gnd.n5408 585
R11095 gnd.n5808 gnd.n5408 585
R11096 gnd.n5788 gnd.n5787 585
R11097 gnd.n5787 gnd.n5415 585
R11098 gnd.n5786 gnd.n5422 585
R11099 gnd.n5786 gnd.n5414 585
R11100 gnd.n5785 gnd.n5424 585
R11101 gnd.n5785 gnd.n5784 585
R11102 gnd.n5764 gnd.n5423 585
R11103 gnd.n5436 gnd.n5423 585
R11104 gnd.n5763 gnd.n5434 585
R11105 gnd.n5774 gnd.n5434 585
R11106 gnd.n5754 gnd.n5441 585
R11107 gnd.n5755 gnd.n5754 585
R11108 gnd.n5753 gnd.n5447 585
R11109 gnd.n5753 gnd.n5752 585
R11110 gnd.n5738 gnd.n5446 585
R11111 gnd.n5457 gnd.n5446 585
R11112 gnd.n5737 gnd.n5455 585
R11113 gnd.n5744 gnd.n5455 585
R11114 gnd.n5736 gnd.n5735 585
R11115 gnd.n5735 gnd.n5734 585
R11116 gnd.n3991 gnd.n3990 585
R11117 gnd.n3992 gnd.n3991 585
R11118 gnd.n3902 gnd.n2092 585
R11119 gnd.n2098 gnd.n2092 585
R11120 gnd.n3901 gnd.n3900 585
R11121 gnd.n3900 gnd.n3899 585
R11122 gnd.n2095 gnd.n2094 585
R11123 gnd.n3874 gnd.n2095 585
R11124 gnd.n3888 gnd.n3887 585
R11125 gnd.n3889 gnd.n3888 585
R11126 gnd.n3886 gnd.n2107 585
R11127 gnd.n3880 gnd.n2107 585
R11128 gnd.n3885 gnd.n3884 585
R11129 gnd.n3884 gnd.n3883 585
R11130 gnd.n2109 gnd.n2108 585
R11131 gnd.n3868 gnd.n2109 585
R11132 gnd.n3854 gnd.n3853 585
R11133 gnd.n3853 gnd.n3852 585
R11134 gnd.n3855 gnd.n2123 585
R11135 gnd.n3715 gnd.n2123 585
R11136 gnd.n3857 gnd.n3856 585
R11137 gnd.n3858 gnd.n3857 585
R11138 gnd.n2124 gnd.n2122 585
R11139 gnd.n2122 gnd.n2120 585
R11140 gnd.n3824 gnd.n3823 585
R11141 gnd.n3825 gnd.n3824 585
R11142 gnd.n3822 gnd.n2135 585
R11143 gnd.n2140 gnd.n2135 585
R11144 gnd.n3821 gnd.n3820 585
R11145 gnd.n3820 gnd.n3819 585
R11146 gnd.n2137 gnd.n2136 585
R11147 gnd.n3726 gnd.n2137 585
R11148 gnd.n3808 gnd.n3807 585
R11149 gnd.n3809 gnd.n3808 585
R11150 gnd.n3806 gnd.n2149 585
R11151 gnd.n3801 gnd.n2149 585
R11152 gnd.n3805 gnd.n3804 585
R11153 gnd.n3804 gnd.n3803 585
R11154 gnd.n2151 gnd.n2150 585
R11155 gnd.t2 gnd.n2151 585
R11156 gnd.n3774 gnd.n3773 585
R11157 gnd.n3773 gnd.n2162 585
R11158 gnd.n3775 gnd.n2172 585
R11159 gnd.n3736 gnd.n2172 585
R11160 gnd.n3777 gnd.n3776 585
R11161 gnd.n3778 gnd.n3777 585
R11162 gnd.n3772 gnd.n2171 585
R11163 gnd.n3767 gnd.n2171 585
R11164 gnd.n3771 gnd.n3770 585
R11165 gnd.n3770 gnd.n3769 585
R11166 gnd.n2174 gnd.n2173 585
R11167 gnd.n2184 gnd.n2174 585
R11168 gnd.n3699 gnd.n3698 585
R11169 gnd.n3699 gnd.n2183 585
R11170 gnd.n3703 gnd.n3702 585
R11171 gnd.n3702 gnd.n3701 585
R11172 gnd.n3704 gnd.n2191 585
R11173 gnd.n3749 gnd.n2191 585
R11174 gnd.n3705 gnd.n2202 585
R11175 gnd.n2202 gnd.n2201 585
R11176 gnd.n3707 gnd.n3706 585
R11177 gnd.n3708 gnd.n3707 585
R11178 gnd.n3697 gnd.n2199 585
R11179 gnd.n3692 gnd.n2199 585
R11180 gnd.n3696 gnd.n3695 585
R11181 gnd.n3695 gnd.n3694 585
R11182 gnd.n2204 gnd.n2203 585
R11183 gnd.n3680 gnd.n2204 585
R11184 gnd.n3670 gnd.n2221 585
R11185 gnd.n2221 gnd.n2213 585
R11186 gnd.n3672 gnd.n3671 585
R11187 gnd.n3673 gnd.n3672 585
R11188 gnd.n3669 gnd.n2220 585
R11189 gnd.n2225 gnd.n2220 585
R11190 gnd.n3668 gnd.n3667 585
R11191 gnd.n3667 gnd.n3666 585
R11192 gnd.n2223 gnd.n2222 585
R11193 gnd.n3623 gnd.n2223 585
R11194 gnd.n3653 gnd.n3652 585
R11195 gnd.n3654 gnd.n3653 585
R11196 gnd.n3651 gnd.n2236 585
R11197 gnd.n2236 gnd.n2232 585
R11198 gnd.n3650 gnd.n3649 585
R11199 gnd.n3649 gnd.n3648 585
R11200 gnd.n2238 gnd.n2237 585
R11201 gnd.n3613 gnd.n2238 585
R11202 gnd.n3598 gnd.n3597 585
R11203 gnd.n3597 gnd.n2248 585
R11204 gnd.n3599 gnd.n2259 585
R11205 gnd.n3583 gnd.n2259 585
R11206 gnd.n3601 gnd.n3600 585
R11207 gnd.n3602 gnd.n3601 585
R11208 gnd.n3596 gnd.n2258 585
R11209 gnd.n2258 gnd.n2254 585
R11210 gnd.n3595 gnd.n3594 585
R11211 gnd.n3594 gnd.n3593 585
R11212 gnd.n2261 gnd.n2260 585
R11213 gnd.n3574 gnd.n2261 585
R11214 gnd.n3559 gnd.n3558 585
R11215 gnd.n3558 gnd.n2272 585
R11216 gnd.n3560 gnd.n2283 585
R11217 gnd.n3547 gnd.n2283 585
R11218 gnd.n3562 gnd.n3561 585
R11219 gnd.n3563 gnd.n3562 585
R11220 gnd.n3557 gnd.n2282 585
R11221 gnd.n2282 gnd.n2278 585
R11222 gnd.n3556 gnd.n3555 585
R11223 gnd.n3555 gnd.n3554 585
R11224 gnd.n2285 gnd.n2284 585
R11225 gnd.n3492 gnd.n2285 585
R11226 gnd.n3534 gnd.n3533 585
R11227 gnd.n3535 gnd.n3534 585
R11228 gnd.n3532 gnd.n2300 585
R11229 gnd.n3526 gnd.n2300 585
R11230 gnd.n3531 gnd.n3530 585
R11231 gnd.n3530 gnd.n3529 585
R11232 gnd.n2302 gnd.n2301 585
R11233 gnd.n3519 gnd.n2302 585
R11234 gnd.n3503 gnd.n3502 585
R11235 gnd.n3502 gnd.n3501 585
R11236 gnd.n3504 gnd.n2317 585
R11237 gnd.n3477 gnd.n2317 585
R11238 gnd.n3506 gnd.n3505 585
R11239 gnd.n3507 gnd.n3506 585
R11240 gnd.n2318 gnd.n2316 585
R11241 gnd.t59 gnd.n2316 585
R11242 gnd.n3469 gnd.n3468 585
R11243 gnd.n3470 gnd.n3469 585
R11244 gnd.n3467 gnd.n2322 585
R11245 gnd.n2322 gnd.n1537 585
R11246 gnd.n3466 gnd.n3465 585
R11247 gnd.n3465 gnd.n1535 585
R11248 gnd.n3464 gnd.n2323 585
R11249 gnd.n3464 gnd.n3463 585
R11250 gnd.n1524 gnd.n1523 585
R11251 gnd.n1527 gnd.n1524 585
R11252 gnd.n4683 gnd.n4682 585
R11253 gnd.n4682 gnd.n4681 585
R11254 gnd.n4684 gnd.n1521 585
R11255 gnd.n3383 gnd.n1521 585
R11256 gnd.n4686 gnd.n4685 585
R11257 gnd.n4687 gnd.n4686 585
R11258 gnd.n1522 gnd.n1520 585
R11259 gnd.n1520 gnd.n1517 585
R11260 gnd.n3392 gnd.n3391 585
R11261 gnd.n3393 gnd.n3392 585
R11262 gnd.n1507 gnd.n1506 585
R11263 gnd.n1509 gnd.n1507 585
R11264 gnd.n4697 gnd.n4696 585
R11265 gnd.n4696 gnd.n4695 585
R11266 gnd.n4698 gnd.n1504 585
R11267 gnd.n2341 gnd.n1504 585
R11268 gnd.n4700 gnd.n4699 585
R11269 gnd.n4701 gnd.n4700 585
R11270 gnd.n1505 gnd.n1503 585
R11271 gnd.n2348 gnd.n1503 585
R11272 gnd.n3405 gnd.n3404 585
R11273 gnd.n3406 gnd.n3405 585
R11274 gnd.n1490 gnd.n1489 585
R11275 gnd.n3408 gnd.n1490 585
R11276 gnd.n4711 gnd.n4710 585
R11277 gnd.n4710 gnd.n4709 585
R11278 gnd.n4712 gnd.n1468 585
R11279 gnd.n3415 gnd.n1468 585
R11280 gnd.n4777 gnd.n4776 585
R11281 gnd.n4775 gnd.n1467 585
R11282 gnd.n4774 gnd.n1466 585
R11283 gnd.n4779 gnd.n1466 585
R11284 gnd.n4773 gnd.n4772 585
R11285 gnd.n4771 gnd.n4770 585
R11286 gnd.n4769 gnd.n4768 585
R11287 gnd.n4767 gnd.n4766 585
R11288 gnd.n4765 gnd.n4764 585
R11289 gnd.n4763 gnd.n4762 585
R11290 gnd.n4761 gnd.n4760 585
R11291 gnd.n4759 gnd.n4758 585
R11292 gnd.n4757 gnd.n4756 585
R11293 gnd.n4755 gnd.n4754 585
R11294 gnd.n4753 gnd.n4752 585
R11295 gnd.n4751 gnd.n4750 585
R11296 gnd.n4749 gnd.n4748 585
R11297 gnd.n4747 gnd.n4746 585
R11298 gnd.n4745 gnd.n4744 585
R11299 gnd.n4743 gnd.n4742 585
R11300 gnd.n4741 gnd.n4740 585
R11301 gnd.n4739 gnd.n4738 585
R11302 gnd.n4737 gnd.n4736 585
R11303 gnd.n4735 gnd.n4734 585
R11304 gnd.n4733 gnd.n4732 585
R11305 gnd.n4731 gnd.n4730 585
R11306 gnd.n4729 gnd.n4728 585
R11307 gnd.n4727 gnd.n4726 585
R11308 gnd.n4725 gnd.n4724 585
R11309 gnd.n4723 gnd.n4722 585
R11310 gnd.n4721 gnd.n4720 585
R11311 gnd.n4719 gnd.n4718 585
R11312 gnd.n4717 gnd.n1430 585
R11313 gnd.n4782 gnd.n4781 585
R11314 gnd.n1432 gnd.n1429 585
R11315 gnd.n3311 gnd.n3310 585
R11316 gnd.n3313 gnd.n3312 585
R11317 gnd.n3316 gnd.n3315 585
R11318 gnd.n3318 gnd.n3317 585
R11319 gnd.n3320 gnd.n3319 585
R11320 gnd.n3322 gnd.n3321 585
R11321 gnd.n3324 gnd.n3323 585
R11322 gnd.n3326 gnd.n3325 585
R11323 gnd.n3328 gnd.n3327 585
R11324 gnd.n3330 gnd.n3329 585
R11325 gnd.n3332 gnd.n3331 585
R11326 gnd.n3334 gnd.n3333 585
R11327 gnd.n3336 gnd.n3335 585
R11328 gnd.n3338 gnd.n3337 585
R11329 gnd.n3340 gnd.n3339 585
R11330 gnd.n3342 gnd.n3341 585
R11331 gnd.n3344 gnd.n3343 585
R11332 gnd.n3346 gnd.n3345 585
R11333 gnd.n3348 gnd.n3347 585
R11334 gnd.n3350 gnd.n3349 585
R11335 gnd.n3352 gnd.n3351 585
R11336 gnd.n3354 gnd.n3353 585
R11337 gnd.n3356 gnd.n3355 585
R11338 gnd.n3358 gnd.n3357 585
R11339 gnd.n3360 gnd.n3359 585
R11340 gnd.n3362 gnd.n3361 585
R11341 gnd.n3364 gnd.n3363 585
R11342 gnd.n3366 gnd.n3365 585
R11343 gnd.n3368 gnd.n3367 585
R11344 gnd.n3370 gnd.n3369 585
R11345 gnd.n3371 gnd.n3307 585
R11346 gnd.n3995 gnd.n3994 585
R11347 gnd.n3997 gnd.n3996 585
R11348 gnd.n3999 gnd.n3998 585
R11349 gnd.n4001 gnd.n4000 585
R11350 gnd.n4003 gnd.n4002 585
R11351 gnd.n4005 gnd.n4004 585
R11352 gnd.n4007 gnd.n4006 585
R11353 gnd.n4009 gnd.n4008 585
R11354 gnd.n4011 gnd.n4010 585
R11355 gnd.n4013 gnd.n4012 585
R11356 gnd.n4015 gnd.n4014 585
R11357 gnd.n4017 gnd.n4016 585
R11358 gnd.n4019 gnd.n4018 585
R11359 gnd.n4021 gnd.n4020 585
R11360 gnd.n4023 gnd.n4022 585
R11361 gnd.n4025 gnd.n4024 585
R11362 gnd.n4027 gnd.n4026 585
R11363 gnd.n4029 gnd.n4028 585
R11364 gnd.n4031 gnd.n4030 585
R11365 gnd.n4033 gnd.n4032 585
R11366 gnd.n4035 gnd.n4034 585
R11367 gnd.n4037 gnd.n4036 585
R11368 gnd.n4039 gnd.n4038 585
R11369 gnd.n4041 gnd.n4040 585
R11370 gnd.n4043 gnd.n4042 585
R11371 gnd.n4045 gnd.n4044 585
R11372 gnd.n4047 gnd.n4046 585
R11373 gnd.n4049 gnd.n4048 585
R11374 gnd.n4051 gnd.n4050 585
R11375 gnd.n4054 gnd.n4053 585
R11376 gnd.n4056 gnd.n4055 585
R11377 gnd.n4058 gnd.n4057 585
R11378 gnd.n4060 gnd.n4059 585
R11379 gnd.n3924 gnd.n1750 585
R11380 gnd.n3926 gnd.n3925 585
R11381 gnd.n3928 gnd.n3927 585
R11382 gnd.n3930 gnd.n3929 585
R11383 gnd.n3933 gnd.n3932 585
R11384 gnd.n3935 gnd.n3934 585
R11385 gnd.n3937 gnd.n3936 585
R11386 gnd.n3939 gnd.n3938 585
R11387 gnd.n3941 gnd.n3940 585
R11388 gnd.n3943 gnd.n3942 585
R11389 gnd.n3945 gnd.n3944 585
R11390 gnd.n3947 gnd.n3946 585
R11391 gnd.n3949 gnd.n3948 585
R11392 gnd.n3951 gnd.n3950 585
R11393 gnd.n3953 gnd.n3952 585
R11394 gnd.n3955 gnd.n3954 585
R11395 gnd.n3957 gnd.n3956 585
R11396 gnd.n3959 gnd.n3958 585
R11397 gnd.n3961 gnd.n3960 585
R11398 gnd.n3963 gnd.n3962 585
R11399 gnd.n3965 gnd.n3964 585
R11400 gnd.n3967 gnd.n3966 585
R11401 gnd.n3969 gnd.n3968 585
R11402 gnd.n3971 gnd.n3970 585
R11403 gnd.n3973 gnd.n3972 585
R11404 gnd.n3975 gnd.n3974 585
R11405 gnd.n3977 gnd.n3976 585
R11406 gnd.n3979 gnd.n3978 585
R11407 gnd.n3981 gnd.n3980 585
R11408 gnd.n3983 gnd.n3982 585
R11409 gnd.n3985 gnd.n3984 585
R11410 gnd.n3987 gnd.n3986 585
R11411 gnd.n3988 gnd.n2093 585
R11412 gnd.n3993 gnd.n2089 585
R11413 gnd.n3993 gnd.n3992 585
R11414 gnd.n3872 gnd.n2090 585
R11415 gnd.n2098 gnd.n2090 585
R11416 gnd.n3873 gnd.n2097 585
R11417 gnd.n3899 gnd.n2097 585
R11418 gnd.n3876 gnd.n3875 585
R11419 gnd.n3875 gnd.n3874 585
R11420 gnd.n3877 gnd.n2104 585
R11421 gnd.n3889 gnd.n2104 585
R11422 gnd.n3879 gnd.n3878 585
R11423 gnd.n3880 gnd.n3879 585
R11424 gnd.n3871 gnd.n2111 585
R11425 gnd.n3883 gnd.n2111 585
R11426 gnd.n3870 gnd.n3869 585
R11427 gnd.n3869 gnd.n3868 585
R11428 gnd.n2114 gnd.n2113 585
R11429 gnd.n3852 gnd.n2114 585
R11430 gnd.n3717 gnd.n3716 585
R11431 gnd.n3716 gnd.n3715 585
R11432 gnd.n3718 gnd.n2121 585
R11433 gnd.n3858 gnd.n2121 585
R11434 gnd.n3720 gnd.n3719 585
R11435 gnd.n3719 gnd.n2120 585
R11436 gnd.n3721 gnd.n2134 585
R11437 gnd.n3825 gnd.n2134 585
R11438 gnd.n3723 gnd.n3722 585
R11439 gnd.n3722 gnd.n2140 585
R11440 gnd.n3724 gnd.n2139 585
R11441 gnd.n3819 gnd.n2139 585
R11442 gnd.n3728 gnd.n3727 585
R11443 gnd.n3727 gnd.n3726 585
R11444 gnd.n3729 gnd.n2146 585
R11445 gnd.n3809 gnd.n2146 585
R11446 gnd.n3730 gnd.n2154 585
R11447 gnd.n3801 gnd.n2154 585
R11448 gnd.n3731 gnd.n2153 585
R11449 gnd.n3803 gnd.n2153 585
R11450 gnd.n3733 gnd.n3732 585
R11451 gnd.n3733 gnd.t2 585
R11452 gnd.n3734 gnd.n3712 585
R11453 gnd.n3734 gnd.n2162 585
R11454 gnd.n3738 gnd.n3737 585
R11455 gnd.n3737 gnd.n3736 585
R11456 gnd.n3739 gnd.n2168 585
R11457 gnd.n3778 gnd.n2168 585
R11458 gnd.n3740 gnd.n2177 585
R11459 gnd.n3767 gnd.n2177 585
R11460 gnd.n3741 gnd.n2176 585
R11461 gnd.n3769 gnd.n2176 585
R11462 gnd.n3743 gnd.n3742 585
R11463 gnd.n3743 gnd.n2184 585
R11464 gnd.n3745 gnd.n3744 585
R11465 gnd.n3744 gnd.n2183 585
R11466 gnd.n3746 gnd.n2195 585
R11467 gnd.n3701 gnd.n2195 585
R11468 gnd.n3748 gnd.n3747 585
R11469 gnd.n3749 gnd.n3748 585
R11470 gnd.n3711 gnd.n2194 585
R11471 gnd.n2201 gnd.n2194 585
R11472 gnd.n3710 gnd.n3709 585
R11473 gnd.n3709 gnd.n3708 585
R11474 gnd.n2197 gnd.n2196 585
R11475 gnd.n3692 gnd.n2197 585
R11476 gnd.n3677 gnd.n2206 585
R11477 gnd.n3694 gnd.n2206 585
R11478 gnd.n3679 gnd.n3678 585
R11479 gnd.n3680 gnd.n3679 585
R11480 gnd.n3676 gnd.n2215 585
R11481 gnd.n2215 gnd.n2213 585
R11482 gnd.n3675 gnd.n3674 585
R11483 gnd.n3674 gnd.n3673 585
R11484 gnd.n2217 gnd.n2216 585
R11485 gnd.n2225 gnd.n2217 585
R11486 gnd.n3620 gnd.n2224 585
R11487 gnd.n3666 gnd.n2224 585
R11488 gnd.n3622 gnd.n3621 585
R11489 gnd.n3623 gnd.n3622 585
R11490 gnd.n3619 gnd.n2234 585
R11491 gnd.n3654 gnd.n2234 585
R11492 gnd.n3618 gnd.n3617 585
R11493 gnd.n3617 gnd.n2232 585
R11494 gnd.n3616 gnd.n2240 585
R11495 gnd.n3648 gnd.n2240 585
R11496 gnd.n3615 gnd.n3614 585
R11497 gnd.n3614 gnd.n3613 585
R11498 gnd.n2247 gnd.n2246 585
R11499 gnd.n2248 gnd.n2247 585
R11500 gnd.n3582 gnd.n3581 585
R11501 gnd.n3583 gnd.n3582 585
R11502 gnd.n3580 gnd.n2255 585
R11503 gnd.n3602 gnd.n2255 585
R11504 gnd.n3579 gnd.n3578 585
R11505 gnd.n3578 gnd.n2254 585
R11506 gnd.n3577 gnd.n2263 585
R11507 gnd.n3593 gnd.n2263 585
R11508 gnd.n3576 gnd.n3575 585
R11509 gnd.n3575 gnd.n3574 585
R11510 gnd.n2271 gnd.n2270 585
R11511 gnd.n2272 gnd.n2271 585
R11512 gnd.n3549 gnd.n3548 585
R11513 gnd.n3548 gnd.n3547 585
R11514 gnd.n3550 gnd.n2279 585
R11515 gnd.n3563 gnd.n2279 585
R11516 gnd.n3551 gnd.n2289 585
R11517 gnd.n2289 gnd.n2278 585
R11518 gnd.n3553 gnd.n3552 585
R11519 gnd.n3554 gnd.n3553 585
R11520 gnd.n2290 gnd.n2288 585
R11521 gnd.n3492 gnd.n2288 585
R11522 gnd.n3523 gnd.n2299 585
R11523 gnd.n3535 gnd.n2299 585
R11524 gnd.n3525 gnd.n3524 585
R11525 gnd.n3526 gnd.n3525 585
R11526 gnd.n3522 gnd.n2304 585
R11527 gnd.n3529 gnd.n2304 585
R11528 gnd.n3521 gnd.n3520 585
R11529 gnd.n3520 gnd.n3519 585
R11530 gnd.n2306 gnd.n2305 585
R11531 gnd.n3501 gnd.n2306 585
R11532 gnd.n3476 gnd.n3475 585
R11533 gnd.n3477 gnd.n3476 585
R11534 gnd.n3474 gnd.n2314 585
R11535 gnd.n3507 gnd.n2314 585
R11536 gnd.n3473 gnd.n3472 585
R11537 gnd.n3472 gnd.t59 585
R11538 gnd.n2320 gnd.n2319 585
R11539 gnd.n3470 gnd.n2320 585
R11540 gnd.n3375 gnd.n3374 585
R11541 gnd.n3375 gnd.n1537 585
R11542 gnd.n3377 gnd.n3376 585
R11543 gnd.n3376 gnd.n1535 585
R11544 gnd.n3378 gnd.n2325 585
R11545 gnd.n3463 gnd.n2325 585
R11546 gnd.n3380 gnd.n3379 585
R11547 gnd.n3379 gnd.n1527 585
R11548 gnd.n3381 gnd.n1526 585
R11549 gnd.n4681 gnd.n1526 585
R11550 gnd.n3385 gnd.n3384 585
R11551 gnd.n3384 gnd.n3383 585
R11552 gnd.n3386 gnd.n1518 585
R11553 gnd.n4687 gnd.n1518 585
R11554 gnd.n3388 gnd.n3387 585
R11555 gnd.n3388 gnd.n1517 585
R11556 gnd.n3394 gnd.n3373 585
R11557 gnd.n3394 gnd.n3393 585
R11558 gnd.n3396 gnd.n3395 585
R11559 gnd.n3395 gnd.n1509 585
R11560 gnd.n3397 gnd.n1508 585
R11561 gnd.n4695 gnd.n1508 585
R11562 gnd.n3399 gnd.n3398 585
R11563 gnd.n3398 gnd.n2341 585
R11564 gnd.n3400 gnd.n1501 585
R11565 gnd.n4701 gnd.n1501 585
R11566 gnd.n3402 gnd.n3401 585
R11567 gnd.n3402 gnd.n2348 585
R11568 gnd.n3403 gnd.n3372 585
R11569 gnd.n3406 gnd.n3403 585
R11570 gnd.n3410 gnd.n3409 585
R11571 gnd.n3409 gnd.n3408 585
R11572 gnd.n3411 gnd.n1492 585
R11573 gnd.n4709 gnd.n1492 585
R11574 gnd.n3413 gnd.n3412 585
R11575 gnd.n3415 gnd.n3413 585
R11576 gnd.n4833 gnd.n4832 585
R11577 gnd.n4834 gnd.n4833 585
R11578 gnd.n1363 gnd.n1362 585
R11579 gnd.n3143 gnd.n1363 585
R11580 gnd.n4842 gnd.n4841 585
R11581 gnd.n4841 gnd.n4840 585
R11582 gnd.n4843 gnd.n1357 585
R11583 gnd.n3136 gnd.n1357 585
R11584 gnd.n4845 gnd.n4844 585
R11585 gnd.n4846 gnd.n4845 585
R11586 gnd.n1343 gnd.n1342 585
R11587 gnd.n3127 gnd.n1343 585
R11588 gnd.n4854 gnd.n4853 585
R11589 gnd.n4853 gnd.n4852 585
R11590 gnd.n4855 gnd.n1337 585
R11591 gnd.n3121 gnd.n1337 585
R11592 gnd.n4857 gnd.n4856 585
R11593 gnd.n4858 gnd.n4857 585
R11594 gnd.n1322 gnd.n1321 585
R11595 gnd.n3038 gnd.n1322 585
R11596 gnd.n4866 gnd.n4865 585
R11597 gnd.n4865 gnd.n4864 585
R11598 gnd.n4867 gnd.n1316 585
R11599 gnd.n3032 gnd.n1316 585
R11600 gnd.n4869 gnd.n4868 585
R11601 gnd.n4870 gnd.n4869 585
R11602 gnd.n1303 gnd.n1302 585
R11603 gnd.n3026 gnd.n1303 585
R11604 gnd.n4878 gnd.n4877 585
R11605 gnd.n4877 gnd.n4876 585
R11606 gnd.n4879 gnd.n1297 585
R11607 gnd.n3055 gnd.n1297 585
R11608 gnd.n4881 gnd.n4880 585
R11609 gnd.n4882 gnd.n4881 585
R11610 gnd.n1282 gnd.n1281 585
R11611 gnd.n3019 gnd.n1282 585
R11612 gnd.n4890 gnd.n4889 585
R11613 gnd.n4889 gnd.n4888 585
R11614 gnd.n4891 gnd.n1277 585
R11615 gnd.n3011 gnd.n1277 585
R11616 gnd.n4893 gnd.n4892 585
R11617 gnd.n4894 gnd.n4893 585
R11618 gnd.n1262 gnd.n1260 585
R11619 gnd.n3004 gnd.n1262 585
R11620 gnd.n4902 gnd.n4901 585
R11621 gnd.n4901 gnd.n4900 585
R11622 gnd.n1261 gnd.n1259 585
R11623 gnd.n2996 gnd.n1261 585
R11624 gnd.n2966 gnd.n2965 585
R11625 gnd.n2967 gnd.n2966 585
R11626 gnd.n2964 gnd.n2963 585
R11627 gnd.n2963 gnd.n2673 585
R11628 gnd.n2962 gnd.n2678 585
R11629 gnd.n2962 gnd.n2961 585
R11630 gnd.n2677 gnd.n2676 585
R11631 gnd.n2948 gnd.n2676 585
R11632 gnd.n2932 gnd.n2702 585
R11633 gnd.n2932 gnd.n2931 585
R11634 gnd.n2933 gnd.n1258 585
R11635 gnd.n2934 gnd.n2933 585
R11636 gnd.n2701 gnd.n1252 585
R11637 gnd.n2923 gnd.n2701 585
R11638 gnd.n4905 gnd.n1249 585
R11639 gnd.n2709 gnd.n1249 585
R11640 gnd.n4907 gnd.n4906 585
R11641 gnd.n4908 gnd.n4907 585
R11642 gnd.n1234 gnd.n1233 585
R11643 gnd.n2872 gnd.n1234 585
R11644 gnd.n4916 gnd.n4915 585
R11645 gnd.n4915 gnd.n4914 585
R11646 gnd.n4917 gnd.n1228 585
R11647 gnd.n2878 gnd.n1228 585
R11648 gnd.n4919 gnd.n4918 585
R11649 gnd.n4920 gnd.n4919 585
R11650 gnd.n1214 gnd.n1213 585
R11651 gnd.n2884 gnd.n1214 585
R11652 gnd.n4928 gnd.n4927 585
R11653 gnd.n4927 gnd.n4926 585
R11654 gnd.n4929 gnd.n1208 585
R11655 gnd.n2890 gnd.n1208 585
R11656 gnd.n4931 gnd.n4930 585
R11657 gnd.n4932 gnd.n4931 585
R11658 gnd.n1193 gnd.n1192 585
R11659 gnd.n2851 gnd.n1193 585
R11660 gnd.n4940 gnd.n4939 585
R11661 gnd.n4939 gnd.n4938 585
R11662 gnd.n4941 gnd.n1187 585
R11663 gnd.n2842 gnd.n1187 585
R11664 gnd.n4943 gnd.n4942 585
R11665 gnd.n4944 gnd.n4943 585
R11666 gnd.n1174 gnd.n1173 585
R11667 gnd.n1177 gnd.n1174 585
R11668 gnd.n4952 gnd.n4951 585
R11669 gnd.n4951 gnd.n4950 585
R11670 gnd.n4953 gnd.n1168 585
R11671 gnd.n1168 gnd.n1167 585
R11672 gnd.n4955 gnd.n4954 585
R11673 gnd.n4956 gnd.n4955 585
R11674 gnd.n1151 gnd.n1150 585
R11675 gnd.n1155 gnd.n1151 585
R11676 gnd.n4964 gnd.n4963 585
R11677 gnd.n4963 gnd.n4962 585
R11678 gnd.n4965 gnd.n1144 585
R11679 gnd.n1152 gnd.n1144 585
R11680 gnd.n4967 gnd.n4966 585
R11681 gnd.n4968 gnd.n4967 585
R11682 gnd.n1145 gnd.n1071 585
R11683 gnd.n1071 gnd.n1068 585
R11684 gnd.n5090 gnd.n5089 585
R11685 gnd.n5088 gnd.n1070 585
R11686 gnd.n5087 gnd.n1069 585
R11687 gnd.n5092 gnd.n1069 585
R11688 gnd.n5086 gnd.n5085 585
R11689 gnd.n5084 gnd.n5083 585
R11690 gnd.n5082 gnd.n5081 585
R11691 gnd.n5080 gnd.n5079 585
R11692 gnd.n5078 gnd.n5077 585
R11693 gnd.n5076 gnd.n5075 585
R11694 gnd.n5074 gnd.n5073 585
R11695 gnd.n5072 gnd.n5071 585
R11696 gnd.n5070 gnd.n5069 585
R11697 gnd.n5068 gnd.n5067 585
R11698 gnd.n5066 gnd.n5065 585
R11699 gnd.n5064 gnd.n5063 585
R11700 gnd.n5062 gnd.n5061 585
R11701 gnd.n5060 gnd.n5059 585
R11702 gnd.n5058 gnd.n5057 585
R11703 gnd.n5055 gnd.n5054 585
R11704 gnd.n5053 gnd.n5052 585
R11705 gnd.n5051 gnd.n5050 585
R11706 gnd.n5049 gnd.n5048 585
R11707 gnd.n5047 gnd.n5046 585
R11708 gnd.n5045 gnd.n5044 585
R11709 gnd.n5043 gnd.n5042 585
R11710 gnd.n5041 gnd.n5040 585
R11711 gnd.n5039 gnd.n5038 585
R11712 gnd.n5037 gnd.n5036 585
R11713 gnd.n5035 gnd.n5034 585
R11714 gnd.n5033 gnd.n5032 585
R11715 gnd.n5031 gnd.n5030 585
R11716 gnd.n5029 gnd.n5028 585
R11717 gnd.n5027 gnd.n5026 585
R11718 gnd.n5025 gnd.n5024 585
R11719 gnd.n5023 gnd.n5022 585
R11720 gnd.n5021 gnd.n5020 585
R11721 gnd.n5019 gnd.n5018 585
R11722 gnd.n5017 gnd.n5016 585
R11723 gnd.n5015 gnd.n5014 585
R11724 gnd.n5013 gnd.n5012 585
R11725 gnd.n5011 gnd.n5010 585
R11726 gnd.n5009 gnd.n5008 585
R11727 gnd.n5007 gnd.n5006 585
R11728 gnd.n5005 gnd.n5004 585
R11729 gnd.n5003 gnd.n5002 585
R11730 gnd.n5001 gnd.n5000 585
R11731 gnd.n4999 gnd.n4998 585
R11732 gnd.n4997 gnd.n4996 585
R11733 gnd.n4995 gnd.n4994 585
R11734 gnd.n4993 gnd.n4992 585
R11735 gnd.n4991 gnd.n4990 585
R11736 gnd.n4989 gnd.n4988 585
R11737 gnd.n4987 gnd.n4986 585
R11738 gnd.n4985 gnd.n4984 585
R11739 gnd.n4983 gnd.n4982 585
R11740 gnd.n4981 gnd.n4980 585
R11741 gnd.n4979 gnd.n4978 585
R11742 gnd.n4977 gnd.n4976 585
R11743 gnd.n1140 gnd.n1133 585
R11744 gnd.n2552 gnd.n2551 585
R11745 gnd.n2549 gnd.n2445 585
R11746 gnd.n2548 gnd.n2547 585
R11747 gnd.n2541 gnd.n2447 585
R11748 gnd.n2543 gnd.n2542 585
R11749 gnd.n2539 gnd.n2449 585
R11750 gnd.n2538 gnd.n2537 585
R11751 gnd.n2531 gnd.n2451 585
R11752 gnd.n2533 gnd.n2532 585
R11753 gnd.n2529 gnd.n2453 585
R11754 gnd.n2528 gnd.n2527 585
R11755 gnd.n2521 gnd.n2455 585
R11756 gnd.n2523 gnd.n2522 585
R11757 gnd.n2519 gnd.n2457 585
R11758 gnd.n2518 gnd.n2517 585
R11759 gnd.n2511 gnd.n2459 585
R11760 gnd.n2513 gnd.n2512 585
R11761 gnd.n2509 gnd.n2461 585
R11762 gnd.n2508 gnd.n2507 585
R11763 gnd.n2501 gnd.n2463 585
R11764 gnd.n2503 gnd.n2502 585
R11765 gnd.n2499 gnd.n2467 585
R11766 gnd.n2498 gnd.n2497 585
R11767 gnd.n2491 gnd.n2469 585
R11768 gnd.n2493 gnd.n2492 585
R11769 gnd.n2489 gnd.n2471 585
R11770 gnd.n2488 gnd.n2487 585
R11771 gnd.n2481 gnd.n2473 585
R11772 gnd.n2483 gnd.n2482 585
R11773 gnd.n2479 gnd.n2476 585
R11774 gnd.n2478 gnd.n1425 585
R11775 gnd.n4784 gnd.n1421 585
R11776 gnd.n4786 gnd.n4785 585
R11777 gnd.n4788 gnd.n1419 585
R11778 gnd.n4790 gnd.n4789 585
R11779 gnd.n4791 gnd.n1414 585
R11780 gnd.n4793 gnd.n4792 585
R11781 gnd.n4795 gnd.n1412 585
R11782 gnd.n4797 gnd.n4796 585
R11783 gnd.n4799 gnd.n1405 585
R11784 gnd.n4801 gnd.n4800 585
R11785 gnd.n4803 gnd.n1403 585
R11786 gnd.n4805 gnd.n4804 585
R11787 gnd.n4806 gnd.n1398 585
R11788 gnd.n4808 gnd.n4807 585
R11789 gnd.n4810 gnd.n1396 585
R11790 gnd.n4812 gnd.n4811 585
R11791 gnd.n4813 gnd.n1391 585
R11792 gnd.n4815 gnd.n4814 585
R11793 gnd.n4817 gnd.n1389 585
R11794 gnd.n4819 gnd.n4818 585
R11795 gnd.n4820 gnd.n1383 585
R11796 gnd.n4822 gnd.n4821 585
R11797 gnd.n4824 gnd.n1382 585
R11798 gnd.n4825 gnd.n1380 585
R11799 gnd.n4828 gnd.n4827 585
R11800 gnd.n4829 gnd.n1377 585
R11801 gnd.n1381 gnd.n1377 585
R11802 gnd.n3140 gnd.n1374 585
R11803 gnd.n4834 gnd.n1374 585
R11804 gnd.n3142 gnd.n3141 585
R11805 gnd.n3143 gnd.n3142 585
R11806 gnd.n3139 gnd.n1365 585
R11807 gnd.n4840 gnd.n1365 585
R11808 gnd.n3138 gnd.n3137 585
R11809 gnd.n3137 gnd.n3136 585
R11810 gnd.n2629 gnd.n1354 585
R11811 gnd.n4846 gnd.n1354 585
R11812 gnd.n3126 gnd.n3125 585
R11813 gnd.n3127 gnd.n3126 585
R11814 gnd.n3124 gnd.n1344 585
R11815 gnd.n4852 gnd.n1344 585
R11816 gnd.n3123 gnd.n3122 585
R11817 gnd.n3122 gnd.n3121 585
R11818 gnd.n2634 gnd.n1334 585
R11819 gnd.n4858 gnd.n1334 585
R11820 gnd.n3037 gnd.n3036 585
R11821 gnd.n3038 gnd.n3037 585
R11822 gnd.n3035 gnd.n1324 585
R11823 gnd.n4864 gnd.n1324 585
R11824 gnd.n3034 gnd.n3033 585
R11825 gnd.n3033 gnd.n3032 585
R11826 gnd.n3029 gnd.n1314 585
R11827 gnd.n4870 gnd.n1314 585
R11828 gnd.n3028 gnd.n3027 585
R11829 gnd.n3027 gnd.n3026 585
R11830 gnd.n3025 gnd.n1304 585
R11831 gnd.n4876 gnd.n1304 585
R11832 gnd.n3024 gnd.n2648 585
R11833 gnd.n3055 gnd.n2648 585
R11834 gnd.n3022 gnd.n1294 585
R11835 gnd.n4882 gnd.n1294 585
R11836 gnd.n3021 gnd.n3020 585
R11837 gnd.n3020 gnd.n3019 585
R11838 gnd.n2657 gnd.n1284 585
R11839 gnd.n4888 gnd.n1284 585
R11840 gnd.n3010 gnd.n3009 585
R11841 gnd.n3011 gnd.n3010 585
R11842 gnd.n3007 gnd.n1275 585
R11843 gnd.n4894 gnd.n1275 585
R11844 gnd.n3006 gnd.n3005 585
R11845 gnd.n3005 gnd.n3004 585
R11846 gnd.n2662 gnd.n1263 585
R11847 gnd.n4900 gnd.n1263 585
R11848 gnd.n2954 gnd.n2668 585
R11849 gnd.n2996 gnd.n2668 585
R11850 gnd.n2955 gnd.n2674 585
R11851 gnd.n2967 gnd.n2674 585
R11852 gnd.n2953 gnd.n2952 585
R11853 gnd.n2952 gnd.n2673 585
R11854 gnd.n2951 gnd.n2680 585
R11855 gnd.n2961 gnd.n2680 585
R11856 gnd.n2950 gnd.n2949 585
R11857 gnd.n2949 gnd.n2948 585
R11858 gnd.n2691 gnd.n2689 585
R11859 gnd.n2931 gnd.n2691 585
R11860 gnd.n2926 gnd.n2698 585
R11861 gnd.n2934 gnd.n2698 585
R11862 gnd.n2925 gnd.n2924 585
R11863 gnd.n2924 gnd.n2923 585
R11864 gnd.n2708 gnd.n2707 585
R11865 gnd.n2709 gnd.n2708 585
R11866 gnd.n2869 gnd.n1246 585
R11867 gnd.n4908 gnd.n1246 585
R11868 gnd.n2871 gnd.n2870 585
R11869 gnd.n2872 gnd.n2871 585
R11870 gnd.n2859 gnd.n1236 585
R11871 gnd.n4914 gnd.n1236 585
R11872 gnd.n2880 gnd.n2879 585
R11873 gnd.n2879 gnd.n2878 585
R11874 gnd.n2881 gnd.n1225 585
R11875 gnd.n4920 gnd.n1225 585
R11876 gnd.n2883 gnd.n2882 585
R11877 gnd.n2884 gnd.n2883 585
R11878 gnd.n2857 gnd.n1215 585
R11879 gnd.n4926 gnd.n1215 585
R11880 gnd.n2856 gnd.n2735 585
R11881 gnd.n2890 gnd.n2735 585
R11882 gnd.n2854 gnd.n1205 585
R11883 gnd.n4932 gnd.n1205 585
R11884 gnd.n2853 gnd.n2852 585
R11885 gnd.n2852 gnd.n2851 585
R11886 gnd.n2741 gnd.n1195 585
R11887 gnd.n4938 gnd.n1195 585
R11888 gnd.n2841 gnd.n2840 585
R11889 gnd.n2842 gnd.n2841 585
R11890 gnd.n2838 gnd.n1185 585
R11891 gnd.n4944 gnd.n1185 585
R11892 gnd.n2837 gnd.n2836 585
R11893 gnd.n2836 gnd.n1177 585
R11894 gnd.n2835 gnd.n1175 585
R11895 gnd.n4950 gnd.n1175 585
R11896 gnd.n2834 gnd.n2833 585
R11897 gnd.n2833 gnd.n1167 585
R11898 gnd.n2831 gnd.n1165 585
R11899 gnd.n4956 gnd.n1165 585
R11900 gnd.n2830 gnd.n2829 585
R11901 gnd.n2829 gnd.n1155 585
R11902 gnd.n2828 gnd.n1153 585
R11903 gnd.n4962 gnd.n1153 585
R11904 gnd.n2827 gnd.n1141 585
R11905 gnd.n1152 gnd.n1141 585
R11906 gnd.n4969 gnd.n1139 585
R11907 gnd.n4969 gnd.n4968 585
R11908 gnd.n4971 gnd.n4970 585
R11909 gnd.n4970 gnd.n1068 585
R11910 gnd.n7602 gnd.n7601 585
R11911 gnd.n7603 gnd.n7602 585
R11912 gnd.n201 gnd.n200 585
R11913 gnd.n209 gnd.n201 585
R11914 gnd.n7611 gnd.n7610 585
R11915 gnd.n7610 gnd.n7609 585
R11916 gnd.n7612 gnd.n195 585
R11917 gnd.n195 gnd.n194 585
R11918 gnd.n7614 gnd.n7613 585
R11919 gnd.n7615 gnd.n7614 585
R11920 gnd.n182 gnd.n181 585
R11921 gnd.n185 gnd.n182 585
R11922 gnd.n7623 gnd.n7622 585
R11923 gnd.n7622 gnd.n7621 585
R11924 gnd.n7624 gnd.n176 585
R11925 gnd.n176 gnd.n175 585
R11926 gnd.n7626 gnd.n7625 585
R11927 gnd.n7627 gnd.n7626 585
R11928 gnd.n162 gnd.n161 585
R11929 gnd.n7438 gnd.n162 585
R11930 gnd.n7635 gnd.n7634 585
R11931 gnd.n7634 gnd.n7633 585
R11932 gnd.n7636 gnd.n156 585
R11933 gnd.n7417 gnd.n156 585
R11934 gnd.n7638 gnd.n7637 585
R11935 gnd.n7639 gnd.n7638 585
R11936 gnd.n142 gnd.n141 585
R11937 gnd.n7408 gnd.n142 585
R11938 gnd.n7647 gnd.n7646 585
R11939 gnd.n7646 gnd.n7645 585
R11940 gnd.n7648 gnd.n136 585
R11941 gnd.n7402 gnd.n136 585
R11942 gnd.n7650 gnd.n7649 585
R11943 gnd.n7651 gnd.n7650 585
R11944 gnd.n122 gnd.n121 585
R11945 gnd.n7394 gnd.n122 585
R11946 gnd.n7659 gnd.n7658 585
R11947 gnd.n7658 gnd.n7657 585
R11948 gnd.n7660 gnd.n117 585
R11949 gnd.n7388 gnd.n117 585
R11950 gnd.n7662 gnd.n7661 585
R11951 gnd.n7663 gnd.n7662 585
R11952 gnd.n101 gnd.n99 585
R11953 gnd.n7380 gnd.n101 585
R11954 gnd.n7671 gnd.n7670 585
R11955 gnd.n7670 gnd.n7669 585
R11956 gnd.n100 gnd.n92 585
R11957 gnd.n7374 gnd.n100 585
R11958 gnd.n7674 gnd.n90 585
R11959 gnd.n381 gnd.n90 585
R11960 gnd.n7676 gnd.n7675 585
R11961 gnd.n7677 gnd.n7676 585
R11962 gnd.n4315 gnd.n89 585
R11963 gnd.n4307 gnd.n89 585
R11964 gnd.n4317 gnd.n4316 585
R11965 gnd.n4318 gnd.n4317 585
R11966 gnd.n4314 gnd.n1926 585
R11967 gnd.n4314 gnd.n4313 585
R11968 gnd.n1907 gnd.n97 585
R11969 gnd.n1912 gnd.n1907 585
R11970 gnd.n4328 gnd.n1908 585
R11971 gnd.n4328 gnd.n4327 585
R11972 gnd.n4330 gnd.n4329 585
R11973 gnd.n4331 gnd.n4330 585
R11974 gnd.n1894 gnd.n1893 585
R11975 gnd.n4289 gnd.n1894 585
R11976 gnd.n4339 gnd.n4338 585
R11977 gnd.n4338 gnd.n4337 585
R11978 gnd.n4340 gnd.n1888 585
R11979 gnd.n4273 gnd.n1888 585
R11980 gnd.n4342 gnd.n4341 585
R11981 gnd.n4343 gnd.n4342 585
R11982 gnd.n1873 gnd.n1872 585
R11983 gnd.n4234 gnd.n1873 585
R11984 gnd.n4351 gnd.n4350 585
R11985 gnd.n4350 gnd.n4349 585
R11986 gnd.n4352 gnd.n1867 585
R11987 gnd.n4225 gnd.n1867 585
R11988 gnd.n4354 gnd.n4353 585
R11989 gnd.n4355 gnd.n4354 585
R11990 gnd.n1854 gnd.n1853 585
R11991 gnd.n4219 gnd.n1854 585
R11992 gnd.n4363 gnd.n4362 585
R11993 gnd.n4362 gnd.n4361 585
R11994 gnd.n4364 gnd.n1848 585
R11995 gnd.n4248 gnd.n1848 585
R11996 gnd.n4366 gnd.n4365 585
R11997 gnd.n4367 gnd.n4366 585
R11998 gnd.n1833 gnd.n1832 585
R11999 gnd.n4212 gnd.n1833 585
R12000 gnd.n4375 gnd.n4374 585
R12001 gnd.n4374 gnd.n4373 585
R12002 gnd.n4376 gnd.n1827 585
R12003 gnd.n4204 gnd.n1827 585
R12004 gnd.n4378 gnd.n4377 585
R12005 gnd.n4379 gnd.n4378 585
R12006 gnd.n1810 gnd.n1809 585
R12007 gnd.n4197 gnd.n1810 585
R12008 gnd.n4387 gnd.n4386 585
R12009 gnd.n4386 gnd.n4385 585
R12010 gnd.n4388 gnd.n1801 585
R12011 gnd.n4189 gnd.n1801 585
R12012 gnd.n4390 gnd.n4389 585
R12013 gnd.n4391 gnd.n4390 585
R12014 gnd.n1802 gnd.n1800 585
R12015 gnd.n1970 gnd.n1800 585
R12016 gnd.n1803 gnd.n1721 585
R12017 gnd.n4399 gnd.n1721 585
R12018 gnd.n4518 gnd.n4517 585
R12019 gnd.n4516 gnd.n1720 585
R12020 gnd.n4515 gnd.n1719 585
R12021 gnd.n4520 gnd.n1719 585
R12022 gnd.n4514 gnd.n4513 585
R12023 gnd.n4512 gnd.n4511 585
R12024 gnd.n4510 gnd.n4509 585
R12025 gnd.n4508 gnd.n4507 585
R12026 gnd.n4506 gnd.n4505 585
R12027 gnd.n4504 gnd.n4503 585
R12028 gnd.n4502 gnd.n4501 585
R12029 gnd.n4500 gnd.n4499 585
R12030 gnd.n4498 gnd.n4497 585
R12031 gnd.n4496 gnd.n4495 585
R12032 gnd.n4494 gnd.n4493 585
R12033 gnd.n4492 gnd.n4491 585
R12034 gnd.n4490 gnd.n4489 585
R12035 gnd.n4488 gnd.n4487 585
R12036 gnd.n4486 gnd.n4485 585
R12037 gnd.n4483 gnd.n4482 585
R12038 gnd.n4481 gnd.n4480 585
R12039 gnd.n4479 gnd.n4478 585
R12040 gnd.n4477 gnd.n4476 585
R12041 gnd.n4475 gnd.n4474 585
R12042 gnd.n4473 gnd.n4472 585
R12043 gnd.n4471 gnd.n4470 585
R12044 gnd.n4469 gnd.n4468 585
R12045 gnd.n4466 gnd.n4465 585
R12046 gnd.n4464 gnd.n4463 585
R12047 gnd.n4462 gnd.n4461 585
R12048 gnd.n4460 gnd.n4459 585
R12049 gnd.n4458 gnd.n4457 585
R12050 gnd.n4456 gnd.n4455 585
R12051 gnd.n4454 gnd.n4453 585
R12052 gnd.n4452 gnd.n4451 585
R12053 gnd.n4450 gnd.n4449 585
R12054 gnd.n4448 gnd.n4447 585
R12055 gnd.n4446 gnd.n4445 585
R12056 gnd.n4444 gnd.n4443 585
R12057 gnd.n4442 gnd.n4441 585
R12058 gnd.n4440 gnd.n4439 585
R12059 gnd.n4438 gnd.n4437 585
R12060 gnd.n4436 gnd.n4435 585
R12061 gnd.n4434 gnd.n4433 585
R12062 gnd.n4432 gnd.n4431 585
R12063 gnd.n4430 gnd.n4429 585
R12064 gnd.n4428 gnd.n4427 585
R12065 gnd.n4426 gnd.n4425 585
R12066 gnd.n4424 gnd.n4423 585
R12067 gnd.n4422 gnd.n4421 585
R12068 gnd.n4420 gnd.n4419 585
R12069 gnd.n4418 gnd.n4417 585
R12070 gnd.n4416 gnd.n4415 585
R12071 gnd.n4414 gnd.n4413 585
R12072 gnd.n4412 gnd.n4411 585
R12073 gnd.n4410 gnd.n4409 585
R12074 gnd.n4408 gnd.n4407 585
R12075 gnd.n4402 gnd.n4401 585
R12076 gnd.n7493 gnd.n7492 585
R12077 gnd.n7495 gnd.n315 585
R12078 gnd.n7497 gnd.n7496 585
R12079 gnd.n7498 gnd.n308 585
R12080 gnd.n7500 gnd.n7499 585
R12081 gnd.n7502 gnd.n306 585
R12082 gnd.n7504 gnd.n7503 585
R12083 gnd.n7505 gnd.n301 585
R12084 gnd.n7507 gnd.n7506 585
R12085 gnd.n7509 gnd.n299 585
R12086 gnd.n7511 gnd.n7510 585
R12087 gnd.n7512 gnd.n294 585
R12088 gnd.n7514 gnd.n7513 585
R12089 gnd.n7516 gnd.n292 585
R12090 gnd.n7518 gnd.n7517 585
R12091 gnd.n7519 gnd.n287 585
R12092 gnd.n7521 gnd.n7520 585
R12093 gnd.n7523 gnd.n286 585
R12094 gnd.n7524 gnd.n283 585
R12095 gnd.n7527 gnd.n7526 585
R12096 gnd.n285 gnd.n279 585
R12097 gnd.n7531 gnd.n276 585
R12098 gnd.n7533 gnd.n7532 585
R12099 gnd.n7535 gnd.n274 585
R12100 gnd.n7537 gnd.n7536 585
R12101 gnd.n7538 gnd.n269 585
R12102 gnd.n7540 gnd.n7539 585
R12103 gnd.n7542 gnd.n267 585
R12104 gnd.n7544 gnd.n7543 585
R12105 gnd.n7545 gnd.n262 585
R12106 gnd.n7547 gnd.n7546 585
R12107 gnd.n7549 gnd.n260 585
R12108 gnd.n7551 gnd.n7550 585
R12109 gnd.n7552 gnd.n255 585
R12110 gnd.n7554 gnd.n7553 585
R12111 gnd.n7556 gnd.n253 585
R12112 gnd.n7558 gnd.n7557 585
R12113 gnd.n7559 gnd.n248 585
R12114 gnd.n7561 gnd.n7560 585
R12115 gnd.n7563 gnd.n246 585
R12116 gnd.n7565 gnd.n7564 585
R12117 gnd.n7569 gnd.n241 585
R12118 gnd.n7571 gnd.n7570 585
R12119 gnd.n7573 gnd.n239 585
R12120 gnd.n7575 gnd.n7574 585
R12121 gnd.n7576 gnd.n234 585
R12122 gnd.n7578 gnd.n7577 585
R12123 gnd.n7580 gnd.n232 585
R12124 gnd.n7582 gnd.n7581 585
R12125 gnd.n7583 gnd.n227 585
R12126 gnd.n7585 gnd.n7584 585
R12127 gnd.n7587 gnd.n225 585
R12128 gnd.n7589 gnd.n7588 585
R12129 gnd.n7590 gnd.n220 585
R12130 gnd.n7592 gnd.n7591 585
R12131 gnd.n7594 gnd.n218 585
R12132 gnd.n7596 gnd.n7595 585
R12133 gnd.n7597 gnd.n216 585
R12134 gnd.n7598 gnd.n213 585
R12135 gnd.n213 gnd.n212 585
R12136 gnd.n7423 gnd.n210 585
R12137 gnd.n7603 gnd.n210 585
R12138 gnd.n7425 gnd.n7424 585
R12139 gnd.n7424 gnd.n209 585
R12140 gnd.n7426 gnd.n202 585
R12141 gnd.n7609 gnd.n202 585
R12142 gnd.n7428 gnd.n7427 585
R12143 gnd.n7427 gnd.n194 585
R12144 gnd.n7429 gnd.n192 585
R12145 gnd.n7615 gnd.n192 585
R12146 gnd.n7431 gnd.n7430 585
R12147 gnd.n7430 gnd.n185 585
R12148 gnd.n7432 gnd.n183 585
R12149 gnd.n7621 gnd.n183 585
R12150 gnd.n7434 gnd.n7433 585
R12151 gnd.n7433 gnd.n175 585
R12152 gnd.n7435 gnd.n173 585
R12153 gnd.n7627 gnd.n173 585
R12154 gnd.n7437 gnd.n7436 585
R12155 gnd.n7438 gnd.n7437 585
R12156 gnd.n7420 gnd.n164 585
R12157 gnd.n7633 gnd.n164 585
R12158 gnd.n7419 gnd.n7418 585
R12159 gnd.n7418 gnd.n7417 585
R12160 gnd.n360 gnd.n154 585
R12161 gnd.n7639 gnd.n154 585
R12162 gnd.n7407 gnd.n7406 585
R12163 gnd.n7408 gnd.n7407 585
R12164 gnd.n7405 gnd.n144 585
R12165 gnd.n7645 gnd.n144 585
R12166 gnd.n7404 gnd.n7403 585
R12167 gnd.n7403 gnd.n7402 585
R12168 gnd.n366 gnd.n133 585
R12169 gnd.n7651 gnd.n133 585
R12170 gnd.n7393 gnd.n7392 585
R12171 gnd.n7394 gnd.n7393 585
R12172 gnd.n7391 gnd.n124 585
R12173 gnd.n7657 gnd.n124 585
R12174 gnd.n7390 gnd.n7389 585
R12175 gnd.n7389 gnd.n7388 585
R12176 gnd.n372 gnd.n115 585
R12177 gnd.n7663 gnd.n115 585
R12178 gnd.n7379 gnd.n7378 585
R12179 gnd.n7380 gnd.n7379 585
R12180 gnd.n7377 gnd.n103 585
R12181 gnd.n7669 gnd.n103 585
R12182 gnd.n7376 gnd.n7375 585
R12183 gnd.n7375 gnd.n7374 585
R12184 gnd.n380 gnd.n378 585
R12185 gnd.n381 gnd.n380 585
R12186 gnd.n4304 gnd.n86 585
R12187 gnd.n7677 gnd.n86 585
R12188 gnd.n4306 gnd.n4305 585
R12189 gnd.n4307 gnd.n4306 585
R12190 gnd.n4299 gnd.n1922 585
R12191 gnd.n4318 gnd.n1922 585
R12192 gnd.n4298 gnd.n1928 585
R12193 gnd.n4313 gnd.n1928 585
R12194 gnd.n4297 gnd.n4296 585
R12195 gnd.n4296 gnd.n1912 585
R12196 gnd.n4293 gnd.n1910 585
R12197 gnd.n4327 gnd.n1910 585
R12198 gnd.n4292 gnd.n1905 585
R12199 gnd.n4331 gnd.n1905 585
R12200 gnd.n4291 gnd.n4290 585
R12201 gnd.n4290 gnd.n4289 585
R12202 gnd.n1936 gnd.n1895 585
R12203 gnd.n4337 gnd.n1895 585
R12204 gnd.n4230 gnd.n1941 585
R12205 gnd.n4273 gnd.n1941 585
R12206 gnd.n4231 gnd.n1885 585
R12207 gnd.n4343 gnd.n1885 585
R12208 gnd.n4233 gnd.n4232 585
R12209 gnd.n4234 gnd.n4233 585
R12210 gnd.n4228 gnd.n1875 585
R12211 gnd.n4349 gnd.n1875 585
R12212 gnd.n4227 gnd.n4226 585
R12213 gnd.n4226 gnd.n4225 585
R12214 gnd.n4222 gnd.n1865 585
R12215 gnd.n4355 gnd.n1865 585
R12216 gnd.n4221 gnd.n4220 585
R12217 gnd.n4220 gnd.n4219 585
R12218 gnd.n4218 gnd.n1855 585
R12219 gnd.n4361 gnd.n1855 585
R12220 gnd.n4217 gnd.n1953 585
R12221 gnd.n4248 gnd.n1953 585
R12222 gnd.n4215 gnd.n1845 585
R12223 gnd.n4367 gnd.n1845 585
R12224 gnd.n4214 gnd.n4213 585
R12225 gnd.n4213 gnd.n4212 585
R12226 gnd.n1961 gnd.n1835 585
R12227 gnd.n4373 gnd.n1835 585
R12228 gnd.n4203 gnd.n4202 585
R12229 gnd.n4204 gnd.n4203 585
R12230 gnd.n4200 gnd.n1825 585
R12231 gnd.n4379 gnd.n1825 585
R12232 gnd.n4199 gnd.n4198 585
R12233 gnd.n4198 gnd.n4197 585
R12234 gnd.n1966 gnd.n1812 585
R12235 gnd.n4385 gnd.n1812 585
R12236 gnd.n1795 gnd.n1794 585
R12237 gnd.n4189 gnd.n1795 585
R12238 gnd.n4393 gnd.n4392 585
R12239 gnd.n4392 gnd.n4391 585
R12240 gnd.n4394 gnd.n1784 585
R12241 gnd.n1970 gnd.n1784 585
R12242 gnd.n4400 gnd.n1785 585
R12243 gnd.n4400 gnd.n4399 585
R12244 gnd.n2726 gnd.n2725 585
R12245 gnd.n2726 gnd.n1184 585
R12246 gnd.n7344 gnd.n7343 585
R12247 gnd.n7343 gnd.n172 585
R12248 gnd.n7347 gnd.n399 585
R12249 gnd.n399 gnd.n163 585
R12250 gnd.n7349 gnd.n7348 585
R12251 gnd.n7349 gnd.n362 585
R12252 gnd.n7350 gnd.n398 585
R12253 gnd.n7350 gnd.n153 585
R12254 gnd.n7352 gnd.n7351 585
R12255 gnd.n7351 gnd.n146 585
R12256 gnd.n7353 gnd.n393 585
R12257 gnd.n393 gnd.n143 585
R12258 gnd.n7355 gnd.n7354 585
R12259 gnd.n7355 gnd.n135 585
R12260 gnd.n7356 gnd.n392 585
R12261 gnd.n7356 gnd.n132 585
R12262 gnd.n7358 gnd.n7357 585
R12263 gnd.n7357 gnd.n371 585
R12264 gnd.n7359 gnd.n387 585
R12265 gnd.n387 gnd.n123 585
R12266 gnd.n7361 gnd.n7360 585
R12267 gnd.n7361 gnd.n374 585
R12268 gnd.n7362 gnd.n386 585
R12269 gnd.n7362 gnd.n114 585
R12270 gnd.n7364 gnd.n7363 585
R12271 gnd.n7363 gnd.n105 585
R12272 gnd.n7365 gnd.n383 585
R12273 gnd.n383 gnd.n102 585
R12274 gnd.n7368 gnd.n7367 585
R12275 gnd.n7369 gnd.n7368 585
R12276 gnd.n384 gnd.n382 585
R12277 gnd.n382 gnd.n87 585
R12278 gnd.n1919 gnd.n1917 585
R12279 gnd.n1917 gnd.n85 585
R12280 gnd.n1921 gnd.n1920 585
R12281 gnd.n1924 gnd.n1921 585
R12282 gnd.n4321 gnd.n4320 585
R12283 gnd.n4320 gnd.n4319 585
R12284 gnd.n4322 gnd.n1914 585
R12285 gnd.n1927 gnd.n1914 585
R12286 gnd.n4325 gnd.n4324 585
R12287 gnd.n4326 gnd.n4325 585
R12288 gnd.n1915 gnd.n1913 585
R12289 gnd.n1913 gnd.n1909 585
R12290 gnd.n4268 gnd.n4267 585
R12291 gnd.n4267 gnd.n1904 585
R12292 gnd.n4269 gnd.n1943 585
R12293 gnd.n1943 gnd.n1897 585
R12294 gnd.n4271 gnd.n4270 585
R12295 gnd.n4272 gnd.n4271 585
R12296 gnd.n1944 gnd.n1942 585
R12297 gnd.n1942 gnd.n1887 585
R12298 gnd.n4261 gnd.n4260 585
R12299 gnd.n4260 gnd.n1884 585
R12300 gnd.n4259 gnd.n1946 585
R12301 gnd.n4259 gnd.n1877 585
R12302 gnd.n4258 gnd.n4257 585
R12303 gnd.n4258 gnd.n1874 585
R12304 gnd.n1948 gnd.n1947 585
R12305 gnd.n4224 gnd.n1947 585
R12306 gnd.n4253 gnd.n4252 585
R12307 gnd.n4252 gnd.n1864 585
R12308 gnd.n4251 gnd.n1950 585
R12309 gnd.n4251 gnd.n1857 585
R12310 gnd.n4250 gnd.n1952 585
R12311 gnd.n4250 gnd.n4249 585
R12312 gnd.n4153 gnd.n1951 585
R12313 gnd.n1951 gnd.n1847 585
R12314 gnd.n4155 gnd.n4154 585
R12315 gnd.n4154 gnd.n1844 585
R12316 gnd.n4156 gnd.n4146 585
R12317 gnd.n4146 gnd.n1837 585
R12318 gnd.n4158 gnd.n4157 585
R12319 gnd.n4158 gnd.n1834 585
R12320 gnd.n4159 gnd.n4145 585
R12321 gnd.n4159 gnd.n1965 585
R12322 gnd.n4161 gnd.n4160 585
R12323 gnd.n4160 gnd.n1824 585
R12324 gnd.n4162 gnd.n4140 585
R12325 gnd.n4140 gnd.n1814 585
R12326 gnd.n4164 gnd.n4163 585
R12327 gnd.n4164 gnd.n1811 585
R12328 gnd.n4165 gnd.n4139 585
R12329 gnd.n4165 gnd.n1798 585
R12330 gnd.n4167 gnd.n4166 585
R12331 gnd.n4166 gnd.n1796 585
R12332 gnd.n4168 gnd.n4134 585
R12333 gnd.n4134 gnd.n1788 585
R12334 gnd.n4170 gnd.n4169 585
R12335 gnd.n4170 gnd.n1786 585
R12336 gnd.n4171 gnd.n4133 585
R12337 gnd.n4171 gnd.n1718 585
R12338 gnd.n4173 gnd.n4172 585
R12339 gnd.n4172 gnd.n1676 585
R12340 gnd.n4174 gnd.n2004 585
R12341 gnd.n2004 gnd.n2002 585
R12342 gnd.n4176 gnd.n4175 585
R12343 gnd.n4177 gnd.n4176 585
R12344 gnd.n2005 gnd.n2003 585
R12345 gnd.n2003 gnd.n1978 585
R12346 gnd.n4127 gnd.n4126 585
R12347 gnd.n4126 gnd.n4125 585
R12348 gnd.n2008 gnd.n2007 585
R12349 gnd.n4122 gnd.n2008 585
R12350 gnd.n4108 gnd.n2019 585
R12351 gnd.n2019 gnd.n2009 585
R12352 gnd.n4110 gnd.n4109 585
R12353 gnd.n4111 gnd.n4110 585
R12354 gnd.n2020 gnd.n2018 585
R12355 gnd.n2018 gnd.n2016 585
R12356 gnd.n4103 gnd.n4102 585
R12357 gnd.n4102 gnd.n4101 585
R12358 gnd.n2023 gnd.n2022 585
R12359 gnd.n2024 gnd.n2023 585
R12360 gnd.n4088 gnd.n4087 585
R12361 gnd.n4089 gnd.n4088 585
R12362 gnd.n2033 gnd.n2032 585
R12363 gnd.n2032 gnd.n2030 585
R12364 gnd.n4083 gnd.n4082 585
R12365 gnd.n4082 gnd.n4081 585
R12366 gnd.n2036 gnd.n2035 585
R12367 gnd.n2037 gnd.n2036 585
R12368 gnd.n4068 gnd.n4067 585
R12369 gnd.n4069 gnd.n4068 585
R12370 gnd.n2046 gnd.n2045 585
R12371 gnd.n2045 gnd.n2043 585
R12372 gnd.n4063 gnd.n4062 585
R12373 gnd.n4062 gnd.n4061 585
R12374 gnd.n2049 gnd.n2048 585
R12375 gnd.n2091 gnd.n2049 585
R12376 gnd.n3897 gnd.n3896 585
R12377 gnd.n3898 gnd.n3897 585
R12378 gnd.n2100 gnd.n2099 585
R12379 gnd.n3874 gnd.n2099 585
R12380 gnd.n3892 gnd.n3891 585
R12381 gnd.n3891 gnd.n3890 585
R12382 gnd.n2103 gnd.n2102 585
R12383 gnd.n3882 gnd.n2103 585
R12384 gnd.n3866 gnd.n3865 585
R12385 gnd.n3867 gnd.n3866 585
R12386 gnd.n2116 gnd.n2115 585
R12387 gnd.n2125 gnd.n2115 585
R12388 gnd.n3861 gnd.n3860 585
R12389 gnd.n3860 gnd.n3859 585
R12390 gnd.n2119 gnd.n2118 585
R12391 gnd.n3826 gnd.n2119 585
R12392 gnd.n3817 gnd.n3816 585
R12393 gnd.n3818 gnd.n3817 585
R12394 gnd.n2142 gnd.n2141 585
R12395 gnd.n3725 gnd.n2141 585
R12396 gnd.n3812 gnd.n3811 585
R12397 gnd.n3811 gnd.n3810 585
R12398 gnd.n2145 gnd.n2144 585
R12399 gnd.n3802 gnd.n2145 585
R12400 gnd.n3786 gnd.n3785 585
R12401 gnd.n3787 gnd.n3786 585
R12402 gnd.n2164 gnd.n2163 585
R12403 gnd.n3735 gnd.n2163 585
R12404 gnd.n3781 gnd.n3780 585
R12405 gnd.n3780 gnd.n3779 585
R12406 gnd.n2167 gnd.n2166 585
R12407 gnd.n3768 gnd.n2167 585
R12408 gnd.n3756 gnd.n3755 585
R12409 gnd.n3757 gnd.n3756 585
R12410 gnd.n2186 gnd.n2185 585
R12411 gnd.n3700 gnd.n2185 585
R12412 gnd.n3751 gnd.n3750 585
R12413 gnd.n3750 gnd.n3749 585
R12414 gnd.n2189 gnd.n2188 585
R12415 gnd.n2200 gnd.n2189 585
R12416 gnd.n3690 gnd.n3689 585
R12417 gnd.n3691 gnd.n3690 585
R12418 gnd.n2209 gnd.n2208 585
R12419 gnd.n2208 gnd.n2205 585
R12420 gnd.n3685 gnd.n3684 585
R12421 gnd.n3684 gnd.n3683 585
R12422 gnd.n2212 gnd.n2211 585
R12423 gnd.n2218 gnd.n2212 585
R12424 gnd.n3664 gnd.n3663 585
R12425 gnd.n3665 gnd.n3664 585
R12426 gnd.n2228 gnd.n2227 585
R12427 gnd.n2235 gnd.n2227 585
R12428 gnd.n3659 gnd.n3658 585
R12429 gnd.n3658 gnd.n3657 585
R12430 gnd.n2231 gnd.n2230 585
R12431 gnd.n2239 gnd.n2231 585
R12432 gnd.n3610 gnd.n3609 585
R12433 gnd.n3611 gnd.n3610 585
R12434 gnd.n2250 gnd.n2249 585
R12435 gnd.n2269 gnd.n2249 585
R12436 gnd.n3605 gnd.n3604 585
R12437 gnd.n3604 gnd.n3603 585
R12438 gnd.n2253 gnd.n2252 585
R12439 gnd.n2262 gnd.n2253 585
R12440 gnd.n3571 gnd.n3570 585
R12441 gnd.n3572 gnd.n3571 585
R12442 gnd.n2274 gnd.n2273 585
R12443 gnd.n2291 gnd.n2273 585
R12444 gnd.n3566 gnd.n3565 585
R12445 gnd.n3565 gnd.n3564 585
R12446 gnd.n2277 gnd.n2276 585
R12447 gnd.n3554 gnd.n2277 585
R12448 gnd.n3494 gnd.n3491 585
R12449 gnd.n3494 gnd.n3493 585
R12450 gnd.n3496 gnd.n3495 585
R12451 gnd.n3495 gnd.n2298 585
R12452 gnd.n3497 gnd.n3480 585
R12453 gnd.n3480 gnd.n2303 585
R12454 gnd.n3499 gnd.n3498 585
R12455 gnd.n3500 gnd.n3499 585
R12456 gnd.n3481 gnd.n3479 585
R12457 gnd.n3479 gnd.n2315 585
R12458 gnd.n3484 gnd.n3483 585
R12459 gnd.n3483 gnd.n2313 585
R12460 gnd.n1534 gnd.n1533 585
R12461 gnd.n2321 gnd.n1534 585
R12462 gnd.n4676 gnd.n4675 585
R12463 gnd.n4675 gnd.n4674 585
R12464 gnd.n4677 gnd.n1528 585
R12465 gnd.n2324 gnd.n1528 585
R12466 gnd.n4679 gnd.n4678 585
R12467 gnd.n4680 gnd.n4679 585
R12468 gnd.n1516 gnd.n1515 585
R12469 gnd.n3382 gnd.n1516 585
R12470 gnd.n4690 gnd.n4689 585
R12471 gnd.n4689 gnd.n4688 585
R12472 gnd.n4691 gnd.n1510 585
R12473 gnd.n3390 gnd.n1510 585
R12474 gnd.n4693 gnd.n4692 585
R12475 gnd.n4694 gnd.n4693 585
R12476 gnd.n1500 gnd.n1499 585
R12477 gnd.n2340 gnd.n1500 585
R12478 gnd.n4704 gnd.n4703 585
R12479 gnd.n4703 gnd.n4702 585
R12480 gnd.n4705 gnd.n1494 585
R12481 gnd.n3406 gnd.n1494 585
R12482 gnd.n4707 gnd.n4706 585
R12483 gnd.n4708 gnd.n4707 585
R12484 gnd.n1495 gnd.n1493 585
R12485 gnd.n3414 gnd.n1493 585
R12486 gnd.n3282 gnd.n3281 585
R12487 gnd.n3282 gnd.n1465 585
R12488 gnd.n3284 gnd.n3283 585
R12489 gnd.n3283 gnd.n2361 585
R12490 gnd.n3285 gnd.n2373 585
R12491 gnd.n2373 gnd.n2372 585
R12492 gnd.n3287 gnd.n3286 585
R12493 gnd.n3288 gnd.n3287 585
R12494 gnd.n2374 gnd.n2371 585
R12495 gnd.n2371 gnd.n2368 585
R12496 gnd.n3273 gnd.n3272 585
R12497 gnd.n3272 gnd.n3271 585
R12498 gnd.n2377 gnd.n2376 585
R12499 gnd.n2386 gnd.n2377 585
R12500 gnd.n3248 gnd.n2398 585
R12501 gnd.n2398 gnd.n2385 585
R12502 gnd.n3250 gnd.n3249 585
R12503 gnd.n3251 gnd.n3250 585
R12504 gnd.n2399 gnd.n2397 585
R12505 gnd.n2397 gnd.n2394 585
R12506 gnd.n3243 gnd.n3242 585
R12507 gnd.n3242 gnd.n3241 585
R12508 gnd.n2402 gnd.n2401 585
R12509 gnd.n2411 gnd.n2402 585
R12510 gnd.n3095 gnd.n3094 585
R12511 gnd.n3094 gnd.n2410 585
R12512 gnd.n3096 gnd.n3089 585
R12513 gnd.n3089 gnd.n3088 585
R12514 gnd.n3098 gnd.n3097 585
R12515 gnd.n3098 gnd.n2433 585
R12516 gnd.n3099 gnd.n3086 585
R12517 gnd.n3099 gnd.n2419 585
R12518 gnd.n3103 gnd.n3102 585
R12519 gnd.n3102 gnd.n3101 585
R12520 gnd.n3104 gnd.n3081 585
R12521 gnd.n3100 gnd.n3081 585
R12522 gnd.n3107 gnd.n3105 585
R12523 gnd.n3107 gnd.n3106 585
R12524 gnd.n3108 gnd.n3080 585
R12525 gnd.n3108 gnd.n1376 585
R12526 gnd.n3110 gnd.n3109 585
R12527 gnd.n3109 gnd.n1373 585
R12528 gnd.n3111 gnd.n3075 585
R12529 gnd.n3075 gnd.n1367 585
R12530 gnd.n3113 gnd.n3112 585
R12531 gnd.n3113 gnd.n1364 585
R12532 gnd.n3114 gnd.n3074 585
R12533 gnd.n3114 gnd.n1356 585
R12534 gnd.n3116 gnd.n3115 585
R12535 gnd.n3115 gnd.n1353 585
R12536 gnd.n3117 gnd.n2638 585
R12537 gnd.n2638 gnd.n1346 585
R12538 gnd.n3119 gnd.n3118 585
R12539 gnd.n3120 gnd.n3119 585
R12540 gnd.n2639 gnd.n2637 585
R12541 gnd.n2637 gnd.n1336 585
R12542 gnd.n3068 gnd.n3067 585
R12543 gnd.n3067 gnd.n1333 585
R12544 gnd.n3066 gnd.n2641 585
R12545 gnd.n3066 gnd.n1326 585
R12546 gnd.n3065 gnd.n3064 585
R12547 gnd.n3065 gnd.n1323 585
R12548 gnd.n2643 gnd.n2642 585
R12549 gnd.n3031 gnd.n2642 585
R12550 gnd.n3060 gnd.n3059 585
R12551 gnd.n3059 gnd.n1313 585
R12552 gnd.n3058 gnd.n2645 585
R12553 gnd.n3058 gnd.n1306 585
R12554 gnd.n3057 gnd.n2647 585
R12555 gnd.n3057 gnd.n3056 585
R12556 gnd.n2982 gnd.n2646 585
R12557 gnd.n2646 gnd.n1296 585
R12558 gnd.n2984 gnd.n2983 585
R12559 gnd.n2983 gnd.n1293 585
R12560 gnd.n2985 gnd.n2975 585
R12561 gnd.n2975 gnd.n1286 585
R12562 gnd.n2987 gnd.n2986 585
R12563 gnd.n2987 gnd.n1283 585
R12564 gnd.n2988 gnd.n2974 585
R12565 gnd.n2988 gnd.n2661 585
R12566 gnd.n2990 gnd.n2989 585
R12567 gnd.n2989 gnd.n1274 585
R12568 gnd.n2991 gnd.n2670 585
R12569 gnd.n2670 gnd.n1265 585
R12570 gnd.n2994 gnd.n2993 585
R12571 gnd.n2995 gnd.n2994 585
R12572 gnd.n2972 gnd.n2669 585
R12573 gnd.n2669 gnd.n2667 585
R12574 gnd.n2970 gnd.n2969 585
R12575 gnd.n2969 gnd.n2968 585
R12576 gnd.n2672 gnd.n2671 585
R12577 gnd.n2682 gnd.n2672 585
R12578 gnd.n2911 gnd.n2909 585
R12579 gnd.n2909 gnd.n2679 585
R12580 gnd.n2913 gnd.n2912 585
R12581 gnd.n2913 gnd.n2703 585
R12582 gnd.n2915 gnd.n2914 585
R12583 gnd.n2914 gnd.n2699 585
R12584 gnd.n2916 gnd.n2711 585
R12585 gnd.n2711 gnd.n2697 585
R12586 gnd.n2919 gnd.n2918 585
R12587 gnd.n2920 gnd.n2919 585
R12588 gnd.n2907 gnd.n2710 585
R12589 gnd.n2710 gnd.n1248 585
R12590 gnd.n2901 gnd.n2712 585
R12591 gnd.n2901 gnd.n1245 585
R12592 gnd.n2903 gnd.n2902 585
R12593 gnd.n2902 gnd.n1238 585
R12594 gnd.n2900 gnd.n2714 585
R12595 gnd.n2900 gnd.n1235 585
R12596 gnd.n2899 gnd.n2898 585
R12597 gnd.n2899 gnd.n1227 585
R12598 gnd.n2716 gnd.n2715 585
R12599 gnd.n2715 gnd.n1224 585
R12600 gnd.n2894 gnd.n2893 585
R12601 gnd.n2893 gnd.n1217 585
R12602 gnd.n2892 gnd.n2718 585
R12603 gnd.n2892 gnd.n2891 585
R12604 gnd.n2734 gnd.n2733 585
R12605 gnd.n2734 gnd.n1207 585
R12606 gnd.n2720 gnd.n2719 585
R12607 gnd.n2719 gnd.n1204 585
R12608 gnd.n2729 gnd.n2728 585
R12609 gnd.n2728 gnd.n1197 585
R12610 gnd.n2727 gnd.n2722 585
R12611 gnd.n2727 gnd.n1194 585
R12612 gnd.n4123 gnd.n1612 585
R12613 gnd.n4124 gnd.n4123 585
R12614 gnd.n4587 gnd.n1611 585
R12615 gnd.n4121 gnd.n1611 585
R12616 gnd.n4588 gnd.n1610 585
R12617 gnd.n2017 gnd.n1610 585
R12618 gnd.n4589 gnd.n1609 585
R12619 gnd.n4112 gnd.n1609 585
R12620 gnd.n4099 gnd.n1607 585
R12621 gnd.n4100 gnd.n4099 585
R12622 gnd.n4593 gnd.n1606 585
R12623 gnd.n4098 gnd.n1606 585
R12624 gnd.n4594 gnd.n1605 585
R12625 gnd.n2031 gnd.n1605 585
R12626 gnd.n4595 gnd.n1604 585
R12627 gnd.n4090 gnd.n1604 585
R12628 gnd.n4079 gnd.n1602 585
R12629 gnd.n4080 gnd.n4079 585
R12630 gnd.n4599 gnd.n1601 585
R12631 gnd.n4078 gnd.n1601 585
R12632 gnd.n4600 gnd.n1600 585
R12633 gnd.n2044 gnd.n1600 585
R12634 gnd.n4601 gnd.n1599 585
R12635 gnd.n4070 gnd.n1599 585
R12636 gnd.n2068 gnd.n1597 585
R12637 gnd.n2069 gnd.n2068 585
R12638 gnd.n4605 gnd.n1596 585
R12639 gnd.n2050 gnd.n1596 585
R12640 gnd.n4606 gnd.n1595 585
R12641 gnd.n3836 gnd.n1595 585
R12642 gnd.n4607 gnd.n1594 585
R12643 gnd.n2096 gnd.n1594 585
R12644 gnd.n2105 gnd.n1592 585
R12645 gnd.n2106 gnd.n2105 585
R12646 gnd.n4611 gnd.n1591 585
R12647 gnd.n3881 gnd.n1591 585
R12648 gnd.n4612 gnd.n1590 585
R12649 gnd.n2110 gnd.n1590 585
R12650 gnd.n4613 gnd.n1589 585
R12651 gnd.n3851 gnd.n1589 585
R12652 gnd.n3713 gnd.n1587 585
R12653 gnd.n3714 gnd.n3713 585
R12654 gnd.n4617 gnd.n1586 585
R12655 gnd.n3827 gnd.n1586 585
R12656 gnd.n4618 gnd.n1585 585
R12657 gnd.n2133 gnd.n1585 585
R12658 gnd.n4619 gnd.n1584 585
R12659 gnd.n2138 gnd.n1584 585
R12660 gnd.n2147 gnd.n1582 585
R12661 gnd.n2148 gnd.n2147 585
R12662 gnd.n4623 gnd.n1581 585
R12663 gnd.n3800 gnd.n1581 585
R12664 gnd.n4624 gnd.n1580 585
R12665 gnd.n2152 gnd.n1580 585
R12666 gnd.n4625 gnd.n1579 585
R12667 gnd.n3788 gnd.n1579 585
R12668 gnd.n2169 gnd.n1577 585
R12669 gnd.n2170 gnd.n2169 585
R12670 gnd.n4629 gnd.n1576 585
R12671 gnd.n3766 gnd.n1576 585
R12672 gnd.n4630 gnd.n1575 585
R12673 gnd.n2175 gnd.n1575 585
R12674 gnd.n4631 gnd.n1574 585
R12675 gnd.n3758 gnd.n1574 585
R12676 gnd.n2192 gnd.n1572 585
R12677 gnd.n2193 gnd.n2192 585
R12678 gnd.n4635 gnd.n1571 585
R12679 gnd.n2190 gnd.n1571 585
R12680 gnd.n4636 gnd.n1570 585
R12681 gnd.n2198 gnd.n1570 585
R12682 gnd.n4637 gnd.n1569 585
R12683 gnd.n3693 gnd.n1569 585
R12684 gnd.n3681 gnd.n1567 585
R12685 gnd.n3682 gnd.n3681 585
R12686 gnd.n4641 gnd.n1566 585
R12687 gnd.n2219 gnd.n1566 585
R12688 gnd.n4642 gnd.n1565 585
R12689 gnd.n2226 gnd.n1565 585
R12690 gnd.n4643 gnd.n1564 585
R12691 gnd.n3624 gnd.n1564 585
R12692 gnd.n3655 gnd.n1562 585
R12693 gnd.n3656 gnd.n3655 585
R12694 gnd.n4647 gnd.n1561 585
R12695 gnd.n3647 gnd.n1561 585
R12696 gnd.n4648 gnd.n1560 585
R12697 gnd.n3612 gnd.n1560 585
R12698 gnd.n4649 gnd.n1559 585
R12699 gnd.n3584 gnd.n1559 585
R12700 gnd.n2256 gnd.n1557 585
R12701 gnd.n2257 gnd.n2256 585
R12702 gnd.n4653 gnd.n1556 585
R12703 gnd.n3592 gnd.n1556 585
R12704 gnd.n4654 gnd.n1555 585
R12705 gnd.n3573 gnd.n1555 585
R12706 gnd.n4655 gnd.n1554 585
R12707 gnd.n3546 gnd.n1554 585
R12708 gnd.n2280 gnd.n1552 585
R12709 gnd.n2281 gnd.n2280 585
R12710 gnd.n4659 gnd.n1551 585
R12711 gnd.n2287 gnd.n1551 585
R12712 gnd.n4660 gnd.n1550 585
R12713 gnd.n2286 gnd.n1550 585
R12714 gnd.n4661 gnd.n1549 585
R12715 gnd.n3536 gnd.n1549 585
R12716 gnd.n3527 gnd.n1547 585
R12717 gnd.n3528 gnd.n3527 585
R12718 gnd.n4665 gnd.n1546 585
R12719 gnd.n3518 gnd.n1546 585
R12720 gnd.n4666 gnd.n1545 585
R12721 gnd.n3478 gnd.n1545 585
R12722 gnd.n4667 gnd.n1544 585
R12723 gnd.n3508 gnd.n1544 585
R12724 gnd.n1541 gnd.n1539 585
R12725 gnd.n3471 gnd.n1539 585
R12726 gnd.n4672 gnd.n4671 585
R12727 gnd.n4673 gnd.n4672 585
R12728 gnd.n1540 gnd.n1538 585
R12729 gnd.n3462 gnd.n1538 585
R12730 gnd.n3444 gnd.n3443 585
R12731 gnd.n3443 gnd.n3442 585
R12732 gnd.n3445 gnd.n3441 585
R12733 gnd.n3441 gnd.n1525 585
R12734 gnd.n2336 gnd.n2334 585
R12735 gnd.n2334 gnd.n1519 585
R12736 gnd.n3450 gnd.n3449 585
R12737 gnd.n3451 gnd.n3450 585
R12738 gnd.n2335 gnd.n2333 585
R12739 gnd.n3389 gnd.n2333 585
R12740 gnd.n3437 gnd.n3436 585
R12741 gnd.n3436 gnd.n3435 585
R12742 gnd.n2339 gnd.n2338 585
R12743 gnd.n2339 gnd.n1502 585
R12744 gnd.n3424 gnd.n3423 585
R12745 gnd.n3425 gnd.n3424 585
R12746 gnd.n2350 gnd.n2349 585
R12747 gnd.n3407 gnd.n2349 585
R12748 gnd.n3419 gnd.n3418 585
R12749 gnd.n3418 gnd.n1491 585
R12750 gnd.n3417 gnd.n2352 585
R12751 gnd.n3417 gnd.n3416 585
R12752 gnd.n2364 gnd.n2353 585
R12753 gnd.n2353 gnd.n1433 585
R12754 gnd.n3297 gnd.n3296 585
R12755 gnd.n3298 gnd.n3297 585
R12756 gnd.n2363 gnd.n2362 585
R12757 gnd.n2370 gnd.n2362 585
R12758 gnd.n3291 gnd.n3290 585
R12759 gnd.n3290 gnd.n3289 585
R12760 gnd.n2367 gnd.n2366 585
R12761 gnd.n3270 gnd.n2367 585
R12762 gnd.n2390 gnd.n2388 585
R12763 gnd.n2388 gnd.n2378 585
R12764 gnd.n3260 gnd.n3259 585
R12765 gnd.n3261 gnd.n3260 585
R12766 gnd.n2389 gnd.n2387 585
R12767 gnd.n2396 gnd.n2387 585
R12768 gnd.n3254 gnd.n3253 585
R12769 gnd.n3253 gnd.n3252 585
R12770 gnd.n2393 gnd.n2392 585
R12771 gnd.n3240 gnd.n2393 585
R12772 gnd.n2415 gnd.n2413 585
R12773 gnd.n2413 gnd.n2403 585
R12774 gnd.n3230 gnd.n3229 585
R12775 gnd.n3231 gnd.n3230 585
R12776 gnd.n2414 gnd.n2412 585
R12777 gnd.n3087 gnd.n2412 585
R12778 gnd.n3224 gnd.n3223 585
R12779 gnd.n2418 gnd.n2417 585
R12780 gnd.n3220 gnd.n3219 585
R12781 gnd.n3221 gnd.n3220 585
R12782 gnd.n2435 gnd.n2434 585
R12783 gnd.n3215 gnd.n2437 585
R12784 gnd.n3214 gnd.n2438 585
R12785 gnd.n3213 gnd.n2439 585
R12786 gnd.n2441 gnd.n2440 585
R12787 gnd.n3208 gnd.n2556 585
R12788 gnd.n3207 gnd.n2557 585
R12789 gnd.n2566 gnd.n2558 585
R12790 gnd.n3200 gnd.n2567 585
R12791 gnd.n3199 gnd.n2568 585
R12792 gnd.n2570 gnd.n2569 585
R12793 gnd.n3192 gnd.n2578 585
R12794 gnd.n3191 gnd.n2579 585
R12795 gnd.n2589 gnd.n2580 585
R12796 gnd.n3184 gnd.n2590 585
R12797 gnd.n3183 gnd.n2591 585
R12798 gnd.n2593 gnd.n2592 585
R12799 gnd.n3176 gnd.n2601 585
R12800 gnd.n3175 gnd.n2602 585
R12801 gnd.n2612 gnd.n2603 585
R12802 gnd.n3168 gnd.n2613 585
R12803 gnd.n3167 gnd.n2614 585
R12804 gnd.n3150 gnd.n3149 585
R12805 gnd.n3152 gnd.n3151 585
R12806 gnd.n3157 gnd.n3153 585
R12807 gnd.n3156 gnd.n3154 585
R12808 gnd.n2012 gnd.n1977 585
R12809 gnd.n4124 gnd.n1977 585
R12810 gnd.n4120 gnd.n4119 585
R12811 gnd.n4121 gnd.n4120 585
R12812 gnd.n2011 gnd.n2010 585
R12813 gnd.n2017 gnd.n2010 585
R12814 gnd.n4114 gnd.n4113 585
R12815 gnd.n4113 gnd.n4112 585
R12816 gnd.n2015 gnd.n2014 585
R12817 gnd.n4100 gnd.n2015 585
R12818 gnd.n4097 gnd.n4096 585
R12819 gnd.n4098 gnd.n4097 585
R12820 gnd.n2026 gnd.n2025 585
R12821 gnd.n2031 gnd.n2025 585
R12822 gnd.n4092 gnd.n4091 585
R12823 gnd.n4091 gnd.n4090 585
R12824 gnd.n2029 gnd.n2028 585
R12825 gnd.n4080 gnd.n2029 585
R12826 gnd.n4077 gnd.n4076 585
R12827 gnd.n4078 gnd.n4077 585
R12828 gnd.n2039 gnd.n2038 585
R12829 gnd.n2044 gnd.n2038 585
R12830 gnd.n4072 gnd.n4071 585
R12831 gnd.n4071 gnd.n4070 585
R12832 gnd.n2042 gnd.n2041 585
R12833 gnd.n2069 gnd.n2042 585
R12834 gnd.n3839 gnd.n3838 585
R12835 gnd.n3838 gnd.n2050 585
R12836 gnd.n3837 gnd.n3835 585
R12837 gnd.n3837 gnd.n3836 585
R12838 gnd.n3843 gnd.n3834 585
R12839 gnd.n3834 gnd.n2096 585
R12840 gnd.n3844 gnd.n3833 585
R12841 gnd.n3833 gnd.n2106 585
R12842 gnd.n3845 gnd.n2112 585
R12843 gnd.n3881 gnd.n2112 585
R12844 gnd.n2129 gnd.n2127 585
R12845 gnd.n2127 gnd.n2110 585
R12846 gnd.n3850 gnd.n3849 585
R12847 gnd.n3851 gnd.n3850 585
R12848 gnd.n2128 gnd.n2126 585
R12849 gnd.n3714 gnd.n2126 585
R12850 gnd.n3829 gnd.n3828 585
R12851 gnd.n3828 gnd.n3827 585
R12852 gnd.n2132 gnd.n2131 585
R12853 gnd.n2133 gnd.n2132 585
R12854 gnd.n3794 gnd.n3793 585
R12855 gnd.n3793 gnd.n2138 585
R12856 gnd.n2158 gnd.n2156 585
R12857 gnd.n2156 gnd.n2148 585
R12858 gnd.n3799 gnd.n3798 585
R12859 gnd.n3800 gnd.n3799 585
R12860 gnd.n2157 gnd.n2155 585
R12861 gnd.n2155 gnd.n2152 585
R12862 gnd.n3790 gnd.n3789 585
R12863 gnd.n3789 gnd.n3788 585
R12864 gnd.n2161 gnd.n2160 585
R12865 gnd.n2170 gnd.n2161 585
R12866 gnd.n3765 gnd.n3764 585
R12867 gnd.n3766 gnd.n3765 585
R12868 gnd.n2179 gnd.n2178 585
R12869 gnd.n2178 gnd.n2175 585
R12870 gnd.n3760 gnd.n3759 585
R12871 gnd.n3759 gnd.n3758 585
R12872 gnd.n2182 gnd.n2181 585
R12873 gnd.n2193 gnd.n2182 585
R12874 gnd.n3633 gnd.n3631 585
R12875 gnd.n3631 gnd.n2190 585
R12876 gnd.n3634 gnd.n3630 585
R12877 gnd.n3630 gnd.n2198 585
R12878 gnd.n3635 gnd.n2207 585
R12879 gnd.n3693 gnd.n2207 585
R12880 gnd.n3628 gnd.n2214 585
R12881 gnd.n3682 gnd.n2214 585
R12882 gnd.n3639 gnd.n3627 585
R12883 gnd.n3627 gnd.n2219 585
R12884 gnd.n3640 gnd.n3626 585
R12885 gnd.n3626 gnd.n2226 585
R12886 gnd.n3641 gnd.n3625 585
R12887 gnd.n3625 gnd.n3624 585
R12888 gnd.n2243 gnd.n2233 585
R12889 gnd.n3656 gnd.n2233 585
R12890 gnd.n3646 gnd.n3645 585
R12891 gnd.n3647 gnd.n3646 585
R12892 gnd.n2242 gnd.n2241 585
R12893 gnd.n3612 gnd.n2241 585
R12894 gnd.n3586 gnd.n3585 585
R12895 gnd.n3585 gnd.n3584 585
R12896 gnd.n2267 gnd.n2265 585
R12897 gnd.n2265 gnd.n2257 585
R12898 gnd.n3591 gnd.n3590 585
R12899 gnd.n3592 gnd.n3591 585
R12900 gnd.n2266 gnd.n2264 585
R12901 gnd.n3573 gnd.n2264 585
R12902 gnd.n3545 gnd.n3544 585
R12903 gnd.n3546 gnd.n3545 585
R12904 gnd.n2293 gnd.n2292 585
R12905 gnd.n2292 gnd.n2281 585
R12906 gnd.n3540 gnd.n3539 585
R12907 gnd.n3539 gnd.n2287 585
R12908 gnd.n3538 gnd.n2295 585
R12909 gnd.n3538 gnd.n2286 585
R12910 gnd.n3537 gnd.n2297 585
R12911 gnd.n3537 gnd.n3536 585
R12912 gnd.n2309 gnd.n2296 585
R12913 gnd.n3528 gnd.n2296 585
R12914 gnd.n3517 gnd.n3516 585
R12915 gnd.n3518 gnd.n3517 585
R12916 gnd.n2308 gnd.n2307 585
R12917 gnd.n3478 gnd.n2307 585
R12918 gnd.n3510 gnd.n3509 585
R12919 gnd.n3509 gnd.n3508 585
R12920 gnd.n2312 gnd.n2311 585
R12921 gnd.n3471 gnd.n2312 585
R12922 gnd.n2328 gnd.n1536 585
R12923 gnd.n4673 gnd.n1536 585
R12924 gnd.n3461 gnd.n3460 585
R12925 gnd.n3462 gnd.n3461 585
R12926 gnd.n2327 gnd.n2326 585
R12927 gnd.n3442 gnd.n2326 585
R12928 gnd.n3455 gnd.n3454 585
R12929 gnd.n3454 gnd.n1525 585
R12930 gnd.n3453 gnd.n2330 585
R12931 gnd.n3453 gnd.n1519 585
R12932 gnd.n3452 gnd.n2332 585
R12933 gnd.n3452 gnd.n3451 585
R12934 gnd.n2344 gnd.n2331 585
R12935 gnd.n3389 gnd.n2331 585
R12936 gnd.n3434 gnd.n3433 585
R12937 gnd.n3435 gnd.n3434 585
R12938 gnd.n2343 gnd.n2342 585
R12939 gnd.n2342 gnd.n1502 585
R12940 gnd.n3427 gnd.n3426 585
R12941 gnd.n3426 gnd.n3425 585
R12942 gnd.n2347 gnd.n2346 585
R12943 gnd.n3407 gnd.n2347 585
R12944 gnd.n2357 gnd.n2355 585
R12945 gnd.n2355 gnd.n1491 585
R12946 gnd.n3306 gnd.n3305 585
R12947 gnd.n3416 gnd.n3306 585
R12948 gnd.n2356 gnd.n2354 585
R12949 gnd.n2354 gnd.n1433 585
R12950 gnd.n3300 gnd.n3299 585
R12951 gnd.n3299 gnd.n3298 585
R12952 gnd.n2360 gnd.n2359 585
R12953 gnd.n2370 gnd.n2360 585
R12954 gnd.n2381 gnd.n2369 585
R12955 gnd.n3289 gnd.n2369 585
R12956 gnd.n3269 gnd.n3268 585
R12957 gnd.n3270 gnd.n3269 585
R12958 gnd.n2380 gnd.n2379 585
R12959 gnd.n2379 gnd.n2378 585
R12960 gnd.n3263 gnd.n3262 585
R12961 gnd.n3262 gnd.n3261 585
R12962 gnd.n2384 gnd.n2383 585
R12963 gnd.n2396 gnd.n2384 585
R12964 gnd.n2406 gnd.n2395 585
R12965 gnd.n3252 gnd.n2395 585
R12966 gnd.n3239 gnd.n3238 585
R12967 gnd.n3240 gnd.n3239 585
R12968 gnd.n2405 gnd.n2404 585
R12969 gnd.n2404 gnd.n2403 585
R12970 gnd.n3233 gnd.n3232 585
R12971 gnd.n3232 gnd.n3231 585
R12972 gnd.n2409 gnd.n2408 585
R12973 gnd.n3087 gnd.n2409 585
R12974 gnd.n4529 gnd.n1667 585
R12975 gnd.n4178 gnd.n1667 585
R12976 gnd.n4530 gnd.n1666 585
R12977 gnd.n1996 gnd.n1660 585
R12978 gnd.n4537 gnd.n1659 585
R12979 gnd.n4538 gnd.n1658 585
R12980 gnd.n1993 gnd.n1652 585
R12981 gnd.n4545 gnd.n1651 585
R12982 gnd.n4546 gnd.n1650 585
R12983 gnd.n1991 gnd.n1644 585
R12984 gnd.n4553 gnd.n1643 585
R12985 gnd.n4554 gnd.n1642 585
R12986 gnd.n1988 gnd.n1636 585
R12987 gnd.n4561 gnd.n1635 585
R12988 gnd.n4562 gnd.n1634 585
R12989 gnd.n1986 gnd.n1627 585
R12990 gnd.n4569 gnd.n1626 585
R12991 gnd.n4570 gnd.n1625 585
R12992 gnd.n1983 gnd.n1622 585
R12993 gnd.n4575 gnd.n1621 585
R12994 gnd.n4576 gnd.n1620 585
R12995 gnd.n4577 gnd.n1619 585
R12996 gnd.n1980 gnd.n1617 585
R12997 gnd.n4581 gnd.n1616 585
R12998 gnd.n4582 gnd.n1615 585
R12999 gnd.n4583 gnd.n1614 585
R13000 gnd.n4181 gnd.n4180 585
R13001 gnd.n4182 gnd.n1976 585
R13002 gnd.n2000 gnd.n1975 585
R13003 gnd.n1999 gnd.n1998 585
R13004 gnd.n3991 gnd.n2093 511.721
R13005 gnd.n3994 gnd.n3993 511.721
R13006 gnd.n3413 gnd.n3307 511.721
R13007 gnd.n4777 gnd.n1468 511.721
R13008 gnd.n6678 gnd.n6677 434.747
R13009 gnd.n3308 gnd.t320 389.64
R13010 gnd.n2087 gnd.t276 389.64
R13011 gnd.n4714 gnd.t240 389.64
R13012 gnd.n3922 gnd.t326 389.64
R13013 gnd.n2615 gnd.t306 371.625
R13014 gnd.n4523 gnd.t335 371.625
R13015 gnd.n2622 gnd.t354 371.625
R13016 gnd.n1740 gnd.t332 371.625
R13017 gnd.n1763 gnd.t323 371.625
R13018 gnd.n4403 gnd.t264 371.625
R13019 gnd.n313 gnd.t351 371.625
R13020 gnd.n280 gnd.t272 371.625
R13021 gnd.n7566 gnd.t313 371.625
R13022 gnd.n350 gnd.t300 371.625
R13023 gnd.n1090 gnd.t287 371.625
R13024 gnd.n1112 gnd.t284 371.625
R13025 gnd.n1134 gnd.t268 371.625
R13026 gnd.n2750 gnd.t338 371.625
R13027 gnd.n1409 gnd.t341 371.625
R13028 gnd.n2443 gnd.t280 371.625
R13029 gnd.n2465 gnd.t303 371.625
R13030 gnd.n1668 gnd.t290 371.625
R13031 gnd.n5689 gnd.t316 323.425
R13032 gnd.n5123 gnd.t344 323.425
R13033 gnd.n6334 gnd.n6308 289.615
R13034 gnd.n6302 gnd.n6276 289.615
R13035 gnd.n6270 gnd.n6244 289.615
R13036 gnd.n6239 gnd.n6213 289.615
R13037 gnd.n6207 gnd.n6181 289.615
R13038 gnd.n6175 gnd.n6149 289.615
R13039 gnd.n6143 gnd.n6117 289.615
R13040 gnd.n6112 gnd.n6086 289.615
R13041 gnd.n5539 gnd.t254 279.217
R13042 gnd.n5167 gnd.t250 279.217
R13043 gnd.n1475 gnd.t263 260.649
R13044 gnd.n3914 gnd.t296 260.649
R13045 gnd.n4779 gnd.n4778 256.663
R13046 gnd.n4779 gnd.n1434 256.663
R13047 gnd.n4779 gnd.n1435 256.663
R13048 gnd.n4779 gnd.n1436 256.663
R13049 gnd.n4779 gnd.n1437 256.663
R13050 gnd.n4779 gnd.n1438 256.663
R13051 gnd.n4779 gnd.n1439 256.663
R13052 gnd.n4779 gnd.n1440 256.663
R13053 gnd.n4779 gnd.n1441 256.663
R13054 gnd.n4779 gnd.n1442 256.663
R13055 gnd.n4779 gnd.n1443 256.663
R13056 gnd.n4779 gnd.n1444 256.663
R13057 gnd.n4779 gnd.n1445 256.663
R13058 gnd.n4779 gnd.n1446 256.663
R13059 gnd.n4779 gnd.n1447 256.663
R13060 gnd.n4779 gnd.n1448 256.663
R13061 gnd.n4782 gnd.n1431 256.663
R13062 gnd.n4780 gnd.n4779 256.663
R13063 gnd.n4779 gnd.n1449 256.663
R13064 gnd.n4779 gnd.n1450 256.663
R13065 gnd.n4779 gnd.n1451 256.663
R13066 gnd.n4779 gnd.n1452 256.663
R13067 gnd.n4779 gnd.n1453 256.663
R13068 gnd.n4779 gnd.n1454 256.663
R13069 gnd.n4779 gnd.n1455 256.663
R13070 gnd.n4779 gnd.n1456 256.663
R13071 gnd.n4779 gnd.n1457 256.663
R13072 gnd.n4779 gnd.n1458 256.663
R13073 gnd.n4779 gnd.n1459 256.663
R13074 gnd.n4779 gnd.n1460 256.663
R13075 gnd.n4779 gnd.n1461 256.663
R13076 gnd.n4779 gnd.n1462 256.663
R13077 gnd.n4779 gnd.n1463 256.663
R13078 gnd.n4779 gnd.n1464 256.663
R13079 gnd.n4060 gnd.n2070 256.663
R13080 gnd.n4060 gnd.n2071 256.663
R13081 gnd.n4060 gnd.n2072 256.663
R13082 gnd.n4060 gnd.n2073 256.663
R13083 gnd.n4060 gnd.n2074 256.663
R13084 gnd.n4060 gnd.n2075 256.663
R13085 gnd.n4060 gnd.n2076 256.663
R13086 gnd.n4060 gnd.n2077 256.663
R13087 gnd.n4060 gnd.n2078 256.663
R13088 gnd.n4060 gnd.n2079 256.663
R13089 gnd.n4060 gnd.n2080 256.663
R13090 gnd.n4060 gnd.n2081 256.663
R13091 gnd.n4060 gnd.n2082 256.663
R13092 gnd.n4060 gnd.n2083 256.663
R13093 gnd.n4060 gnd.n2084 256.663
R13094 gnd.n4060 gnd.n2085 256.663
R13095 gnd.n2086 gnd.n1750 256.663
R13096 gnd.n4060 gnd.n2067 256.663
R13097 gnd.n4060 gnd.n2066 256.663
R13098 gnd.n4060 gnd.n2065 256.663
R13099 gnd.n4060 gnd.n2064 256.663
R13100 gnd.n4060 gnd.n2063 256.663
R13101 gnd.n4060 gnd.n2062 256.663
R13102 gnd.n4060 gnd.n2061 256.663
R13103 gnd.n4060 gnd.n2060 256.663
R13104 gnd.n4060 gnd.n2059 256.663
R13105 gnd.n4060 gnd.n2058 256.663
R13106 gnd.n4060 gnd.n2057 256.663
R13107 gnd.n4060 gnd.n2056 256.663
R13108 gnd.n4060 gnd.n2055 256.663
R13109 gnd.n4060 gnd.n2054 256.663
R13110 gnd.n4060 gnd.n2053 256.663
R13111 gnd.n4060 gnd.n2052 256.663
R13112 gnd.n4060 gnd.n2051 256.663
R13113 gnd.n5092 gnd.n1058 242.672
R13114 gnd.n5092 gnd.n1059 242.672
R13115 gnd.n5092 gnd.n1060 242.672
R13116 gnd.n5092 gnd.n1061 242.672
R13117 gnd.n5092 gnd.n1062 242.672
R13118 gnd.n5092 gnd.n1063 242.672
R13119 gnd.n5092 gnd.n1064 242.672
R13120 gnd.n5092 gnd.n1065 242.672
R13121 gnd.n5092 gnd.n1066 242.672
R13122 gnd.n3160 gnd.n1381 242.672
R13123 gnd.n2620 gnd.n1381 242.672
R13124 gnd.n2608 gnd.n1381 242.672
R13125 gnd.n2605 gnd.n1381 242.672
R13126 gnd.n2596 gnd.n1381 242.672
R13127 gnd.n2585 gnd.n1381 242.672
R13128 gnd.n2582 gnd.n1381 242.672
R13129 gnd.n2573 gnd.n1381 242.672
R13130 gnd.n2562 gnd.n1381 242.672
R13131 gnd.n5594 gnd.n5503 242.672
R13132 gnd.n5507 gnd.n5503 242.672
R13133 gnd.n5587 gnd.n5503 242.672
R13134 gnd.n5581 gnd.n5503 242.672
R13135 gnd.n5579 gnd.n5503 242.672
R13136 gnd.n5573 gnd.n5503 242.672
R13137 gnd.n5571 gnd.n5503 242.672
R13138 gnd.n5565 gnd.n5503 242.672
R13139 gnd.n5563 gnd.n5503 242.672
R13140 gnd.n5557 gnd.n5503 242.672
R13141 gnd.n5555 gnd.n5503 242.672
R13142 gnd.n5548 gnd.n5503 242.672
R13143 gnd.n5546 gnd.n5503 242.672
R13144 gnd.n6390 gnd.n5093 242.672
R13145 gnd.n6396 gnd.n5093 242.672
R13146 gnd.n5170 gnd.n5093 242.672
R13147 gnd.n6403 gnd.n5093 242.672
R13148 gnd.n5161 gnd.n5093 242.672
R13149 gnd.n6410 gnd.n5093 242.672
R13150 gnd.n5154 gnd.n5093 242.672
R13151 gnd.n6417 gnd.n5093 242.672
R13152 gnd.n5147 gnd.n5093 242.672
R13153 gnd.n6424 gnd.n5093 242.672
R13154 gnd.n5140 gnd.n5093 242.672
R13155 gnd.n6431 gnd.n5093 242.672
R13156 gnd.n5133 gnd.n5093 242.672
R13157 gnd.n4520 gnd.n1705 242.672
R13158 gnd.n4520 gnd.n1707 242.672
R13159 gnd.n4520 gnd.n1708 242.672
R13160 gnd.n4520 gnd.n1710 242.672
R13161 gnd.n4520 gnd.n1712 242.672
R13162 gnd.n4520 gnd.n1713 242.672
R13163 gnd.n4520 gnd.n1715 242.672
R13164 gnd.n4520 gnd.n1717 242.672
R13165 gnd.n4521 gnd.n4520 242.672
R13166 gnd.n347 gnd.n212 242.672
R13167 gnd.n7462 gnd.n212 242.672
R13168 gnd.n343 gnd.n212 242.672
R13169 gnd.n7469 gnd.n212 242.672
R13170 gnd.n336 gnd.n212 242.672
R13171 gnd.n7476 gnd.n212 242.672
R13172 gnd.n329 gnd.n212 242.672
R13173 gnd.n7483 gnd.n212 242.672
R13174 gnd.n322 gnd.n212 242.672
R13175 gnd.n5723 gnd.n5722 242.672
R13176 gnd.n5723 gnd.n5664 242.672
R13177 gnd.n5723 gnd.n5665 242.672
R13178 gnd.n5723 gnd.n5666 242.672
R13179 gnd.n5723 gnd.n5667 242.672
R13180 gnd.n5723 gnd.n5668 242.672
R13181 gnd.n5723 gnd.n5669 242.672
R13182 gnd.n5723 gnd.n5670 242.672
R13183 gnd.n6442 gnd.n5093 242.672
R13184 gnd.n5126 gnd.n5093 242.672
R13185 gnd.n6449 gnd.n5093 242.672
R13186 gnd.n5117 gnd.n5093 242.672
R13187 gnd.n6456 gnd.n5093 242.672
R13188 gnd.n5110 gnd.n5093 242.672
R13189 gnd.n6463 gnd.n5093 242.672
R13190 gnd.n5103 gnd.n5093 242.672
R13191 gnd.n5092 gnd.n5091 242.672
R13192 gnd.n5092 gnd.n1030 242.672
R13193 gnd.n5092 gnd.n1031 242.672
R13194 gnd.n5092 gnd.n1032 242.672
R13195 gnd.n5092 gnd.n1033 242.672
R13196 gnd.n5092 gnd.n1034 242.672
R13197 gnd.n5092 gnd.n1035 242.672
R13198 gnd.n5092 gnd.n1036 242.672
R13199 gnd.n5092 gnd.n1037 242.672
R13200 gnd.n5092 gnd.n1038 242.672
R13201 gnd.n5092 gnd.n1039 242.672
R13202 gnd.n5092 gnd.n1040 242.672
R13203 gnd.n5092 gnd.n1041 242.672
R13204 gnd.n5092 gnd.n1042 242.672
R13205 gnd.n5092 gnd.n1043 242.672
R13206 gnd.n5092 gnd.n1044 242.672
R13207 gnd.n5092 gnd.n1045 242.672
R13208 gnd.n5092 gnd.n1046 242.672
R13209 gnd.n5092 gnd.n1047 242.672
R13210 gnd.n5092 gnd.n1048 242.672
R13211 gnd.n5092 gnd.n1049 242.672
R13212 gnd.n5092 gnd.n1050 242.672
R13213 gnd.n5092 gnd.n1051 242.672
R13214 gnd.n5092 gnd.n1052 242.672
R13215 gnd.n5092 gnd.n1053 242.672
R13216 gnd.n5092 gnd.n1054 242.672
R13217 gnd.n5092 gnd.n1055 242.672
R13218 gnd.n5092 gnd.n1056 242.672
R13219 gnd.n5092 gnd.n1057 242.672
R13220 gnd.n2550 gnd.n1381 242.672
R13221 gnd.n2446 gnd.n1381 242.672
R13222 gnd.n2540 gnd.n1381 242.672
R13223 gnd.n2450 gnd.n1381 242.672
R13224 gnd.n2530 gnd.n1381 242.672
R13225 gnd.n2454 gnd.n1381 242.672
R13226 gnd.n2520 gnd.n1381 242.672
R13227 gnd.n2458 gnd.n1381 242.672
R13228 gnd.n2510 gnd.n1381 242.672
R13229 gnd.n2462 gnd.n1381 242.672
R13230 gnd.n2500 gnd.n1381 242.672
R13231 gnd.n2468 gnd.n1381 242.672
R13232 gnd.n2490 gnd.n1381 242.672
R13233 gnd.n2472 gnd.n1381 242.672
R13234 gnd.n2480 gnd.n1381 242.672
R13235 gnd.n2477 gnd.n1381 242.672
R13236 gnd.n4783 gnd.n1427 242.672
R13237 gnd.n1426 gnd.n1381 242.672
R13238 gnd.n4787 gnd.n1381 242.672
R13239 gnd.n1420 gnd.n1381 242.672
R13240 gnd.n4794 gnd.n1381 242.672
R13241 gnd.n1413 gnd.n1381 242.672
R13242 gnd.n4802 gnd.n1381 242.672
R13243 gnd.n1404 gnd.n1381 242.672
R13244 gnd.n4809 gnd.n1381 242.672
R13245 gnd.n1397 gnd.n1381 242.672
R13246 gnd.n4816 gnd.n1381 242.672
R13247 gnd.n1390 gnd.n1381 242.672
R13248 gnd.n4823 gnd.n1381 242.672
R13249 gnd.n4826 gnd.n1381 242.672
R13250 gnd.n4520 gnd.n4519 242.672
R13251 gnd.n4520 gnd.n1677 242.672
R13252 gnd.n4520 gnd.n1678 242.672
R13253 gnd.n4520 gnd.n1679 242.672
R13254 gnd.n4520 gnd.n1680 242.672
R13255 gnd.n4520 gnd.n1681 242.672
R13256 gnd.n4520 gnd.n1682 242.672
R13257 gnd.n4520 gnd.n1683 242.672
R13258 gnd.n4520 gnd.n1684 242.672
R13259 gnd.n4520 gnd.n1685 242.672
R13260 gnd.n4520 gnd.n1686 242.672
R13261 gnd.n4520 gnd.n1687 242.672
R13262 gnd.n4520 gnd.n1688 242.672
R13263 gnd.n4467 gnd.n1751 242.672
R13264 gnd.n4520 gnd.n1689 242.672
R13265 gnd.n4520 gnd.n1690 242.672
R13266 gnd.n4520 gnd.n1691 242.672
R13267 gnd.n4520 gnd.n1692 242.672
R13268 gnd.n4520 gnd.n1693 242.672
R13269 gnd.n4520 gnd.n1694 242.672
R13270 gnd.n4520 gnd.n1695 242.672
R13271 gnd.n4520 gnd.n1696 242.672
R13272 gnd.n4520 gnd.n1697 242.672
R13273 gnd.n4520 gnd.n1698 242.672
R13274 gnd.n4520 gnd.n1699 242.672
R13275 gnd.n4520 gnd.n1700 242.672
R13276 gnd.n4520 gnd.n1701 242.672
R13277 gnd.n4520 gnd.n1702 242.672
R13278 gnd.n4520 gnd.n1703 242.672
R13279 gnd.n4520 gnd.n1704 242.672
R13280 gnd.n7494 gnd.n212 242.672
R13281 gnd.n316 gnd.n212 242.672
R13282 gnd.n7501 gnd.n212 242.672
R13283 gnd.n307 gnd.n212 242.672
R13284 gnd.n7508 gnd.n212 242.672
R13285 gnd.n300 gnd.n212 242.672
R13286 gnd.n7515 gnd.n212 242.672
R13287 gnd.n293 gnd.n212 242.672
R13288 gnd.n7522 gnd.n212 242.672
R13289 gnd.n7525 gnd.n212 242.672
R13290 gnd.n284 gnd.n212 242.672
R13291 gnd.n7534 gnd.n212 242.672
R13292 gnd.n275 gnd.n212 242.672
R13293 gnd.n7541 gnd.n212 242.672
R13294 gnd.n268 gnd.n212 242.672
R13295 gnd.n7548 gnd.n212 242.672
R13296 gnd.n261 gnd.n212 242.672
R13297 gnd.n7555 gnd.n212 242.672
R13298 gnd.n254 gnd.n212 242.672
R13299 gnd.n7562 gnd.n212 242.672
R13300 gnd.n247 gnd.n212 242.672
R13301 gnd.n7572 gnd.n212 242.672
R13302 gnd.n240 gnd.n212 242.672
R13303 gnd.n7579 gnd.n212 242.672
R13304 gnd.n233 gnd.n212 242.672
R13305 gnd.n7586 gnd.n212 242.672
R13306 gnd.n226 gnd.n212 242.672
R13307 gnd.n7593 gnd.n212 242.672
R13308 gnd.n219 gnd.n212 242.672
R13309 gnd.n3222 gnd.n3221 242.672
R13310 gnd.n3221 gnd.n2420 242.672
R13311 gnd.n3221 gnd.n2421 242.672
R13312 gnd.n3221 gnd.n2422 242.672
R13313 gnd.n3221 gnd.n2423 242.672
R13314 gnd.n3221 gnd.n2424 242.672
R13315 gnd.n3221 gnd.n2425 242.672
R13316 gnd.n3221 gnd.n2426 242.672
R13317 gnd.n3221 gnd.n2427 242.672
R13318 gnd.n3221 gnd.n2428 242.672
R13319 gnd.n3221 gnd.n2429 242.672
R13320 gnd.n3221 gnd.n2430 242.672
R13321 gnd.n3221 gnd.n2431 242.672
R13322 gnd.n3221 gnd.n2432 242.672
R13323 gnd.n4178 gnd.n1997 242.672
R13324 gnd.n4178 gnd.n1995 242.672
R13325 gnd.n4178 gnd.n1994 242.672
R13326 gnd.n4178 gnd.n1992 242.672
R13327 gnd.n4178 gnd.n1990 242.672
R13328 gnd.n4178 gnd.n1989 242.672
R13329 gnd.n4178 gnd.n1987 242.672
R13330 gnd.n4178 gnd.n1985 242.672
R13331 gnd.n4178 gnd.n1984 242.672
R13332 gnd.n4178 gnd.n1982 242.672
R13333 gnd.n4178 gnd.n1981 242.672
R13334 gnd.n4178 gnd.n1979 242.672
R13335 gnd.n4179 gnd.n4178 242.672
R13336 gnd.n4178 gnd.n2001 242.672
R13337 gnd.n216 gnd.n213 240.244
R13338 gnd.n7595 gnd.n7594 240.244
R13339 gnd.n7592 gnd.n220 240.244
R13340 gnd.n7588 gnd.n7587 240.244
R13341 gnd.n7585 gnd.n227 240.244
R13342 gnd.n7581 gnd.n7580 240.244
R13343 gnd.n7578 gnd.n234 240.244
R13344 gnd.n7574 gnd.n7573 240.244
R13345 gnd.n7571 gnd.n241 240.244
R13346 gnd.n7564 gnd.n7563 240.244
R13347 gnd.n7561 gnd.n248 240.244
R13348 gnd.n7557 gnd.n7556 240.244
R13349 gnd.n7554 gnd.n255 240.244
R13350 gnd.n7550 gnd.n7549 240.244
R13351 gnd.n7547 gnd.n262 240.244
R13352 gnd.n7543 gnd.n7542 240.244
R13353 gnd.n7540 gnd.n269 240.244
R13354 gnd.n7536 gnd.n7535 240.244
R13355 gnd.n7533 gnd.n276 240.244
R13356 gnd.n7526 gnd.n285 240.244
R13357 gnd.n7524 gnd.n7523 240.244
R13358 gnd.n7521 gnd.n287 240.244
R13359 gnd.n7517 gnd.n7516 240.244
R13360 gnd.n7514 gnd.n294 240.244
R13361 gnd.n7510 gnd.n7509 240.244
R13362 gnd.n7507 gnd.n301 240.244
R13363 gnd.n7503 gnd.n7502 240.244
R13364 gnd.n7500 gnd.n308 240.244
R13365 gnd.n7496 gnd.n7495 240.244
R13366 gnd.n4400 gnd.n1784 240.244
R13367 gnd.n4392 gnd.n1784 240.244
R13368 gnd.n4392 gnd.n1795 240.244
R13369 gnd.n1812 gnd.n1795 240.244
R13370 gnd.n4198 gnd.n1812 240.244
R13371 gnd.n4198 gnd.n1825 240.244
R13372 gnd.n4203 gnd.n1825 240.244
R13373 gnd.n4203 gnd.n1835 240.244
R13374 gnd.n4213 gnd.n1835 240.244
R13375 gnd.n4213 gnd.n1845 240.244
R13376 gnd.n1953 gnd.n1845 240.244
R13377 gnd.n1953 gnd.n1855 240.244
R13378 gnd.n4220 gnd.n1855 240.244
R13379 gnd.n4220 gnd.n1865 240.244
R13380 gnd.n4226 gnd.n1865 240.244
R13381 gnd.n4226 gnd.n1875 240.244
R13382 gnd.n4233 gnd.n1875 240.244
R13383 gnd.n4233 gnd.n1885 240.244
R13384 gnd.n1941 gnd.n1885 240.244
R13385 gnd.n1941 gnd.n1895 240.244
R13386 gnd.n4290 gnd.n1895 240.244
R13387 gnd.n4290 gnd.n1905 240.244
R13388 gnd.n1910 gnd.n1905 240.244
R13389 gnd.n4296 gnd.n1910 240.244
R13390 gnd.n4296 gnd.n1928 240.244
R13391 gnd.n1928 gnd.n1922 240.244
R13392 gnd.n4306 gnd.n1922 240.244
R13393 gnd.n4306 gnd.n86 240.244
R13394 gnd.n380 gnd.n86 240.244
R13395 gnd.n7375 gnd.n380 240.244
R13396 gnd.n7375 gnd.n103 240.244
R13397 gnd.n7379 gnd.n103 240.244
R13398 gnd.n7379 gnd.n115 240.244
R13399 gnd.n7389 gnd.n115 240.244
R13400 gnd.n7389 gnd.n124 240.244
R13401 gnd.n7393 gnd.n124 240.244
R13402 gnd.n7393 gnd.n133 240.244
R13403 gnd.n7403 gnd.n133 240.244
R13404 gnd.n7403 gnd.n144 240.244
R13405 gnd.n7407 gnd.n144 240.244
R13406 gnd.n7407 gnd.n154 240.244
R13407 gnd.n7418 gnd.n154 240.244
R13408 gnd.n7418 gnd.n164 240.244
R13409 gnd.n7437 gnd.n164 240.244
R13410 gnd.n7437 gnd.n173 240.244
R13411 gnd.n7433 gnd.n173 240.244
R13412 gnd.n7433 gnd.n183 240.244
R13413 gnd.n7430 gnd.n183 240.244
R13414 gnd.n7430 gnd.n192 240.244
R13415 gnd.n7427 gnd.n192 240.244
R13416 gnd.n7427 gnd.n202 240.244
R13417 gnd.n7424 gnd.n202 240.244
R13418 gnd.n7424 gnd.n210 240.244
R13419 gnd.n1720 gnd.n1719 240.244
R13420 gnd.n4513 gnd.n1719 240.244
R13421 gnd.n4511 gnd.n4510 240.244
R13422 gnd.n4507 gnd.n4506 240.244
R13423 gnd.n4503 gnd.n4502 240.244
R13424 gnd.n4499 gnd.n4498 240.244
R13425 gnd.n4495 gnd.n4494 240.244
R13426 gnd.n4491 gnd.n4490 240.244
R13427 gnd.n4487 gnd.n4486 240.244
R13428 gnd.n4482 gnd.n4481 240.244
R13429 gnd.n4478 gnd.n4477 240.244
R13430 gnd.n4474 gnd.n4473 240.244
R13431 gnd.n4470 gnd.n4469 240.244
R13432 gnd.n4465 gnd.n4464 240.244
R13433 gnd.n4461 gnd.n4460 240.244
R13434 gnd.n4457 gnd.n4456 240.244
R13435 gnd.n4453 gnd.n4452 240.244
R13436 gnd.n4449 gnd.n4448 240.244
R13437 gnd.n4445 gnd.n4444 240.244
R13438 gnd.n4441 gnd.n4440 240.244
R13439 gnd.n4437 gnd.n4436 240.244
R13440 gnd.n4433 gnd.n4432 240.244
R13441 gnd.n4429 gnd.n4428 240.244
R13442 gnd.n4425 gnd.n4424 240.244
R13443 gnd.n4421 gnd.n4420 240.244
R13444 gnd.n4417 gnd.n4416 240.244
R13445 gnd.n4413 gnd.n4412 240.244
R13446 gnd.n4409 gnd.n4408 240.244
R13447 gnd.n1800 gnd.n1721 240.244
R13448 gnd.n4390 gnd.n1800 240.244
R13449 gnd.n4390 gnd.n1801 240.244
R13450 gnd.n4386 gnd.n1801 240.244
R13451 gnd.n4386 gnd.n1810 240.244
R13452 gnd.n4378 gnd.n1810 240.244
R13453 gnd.n4378 gnd.n1827 240.244
R13454 gnd.n4374 gnd.n1827 240.244
R13455 gnd.n4374 gnd.n1833 240.244
R13456 gnd.n4366 gnd.n1833 240.244
R13457 gnd.n4366 gnd.n1848 240.244
R13458 gnd.n4362 gnd.n1848 240.244
R13459 gnd.n4362 gnd.n1854 240.244
R13460 gnd.n4354 gnd.n1854 240.244
R13461 gnd.n4354 gnd.n1867 240.244
R13462 gnd.n4350 gnd.n1867 240.244
R13463 gnd.n4350 gnd.n1873 240.244
R13464 gnd.n4342 gnd.n1873 240.244
R13465 gnd.n4342 gnd.n1888 240.244
R13466 gnd.n4338 gnd.n1888 240.244
R13467 gnd.n4338 gnd.n1894 240.244
R13468 gnd.n4330 gnd.n1894 240.244
R13469 gnd.n4330 gnd.n4328 240.244
R13470 gnd.n4328 gnd.n1907 240.244
R13471 gnd.n4314 gnd.n1907 240.244
R13472 gnd.n4317 gnd.n4314 240.244
R13473 gnd.n4317 gnd.n89 240.244
R13474 gnd.n7676 gnd.n89 240.244
R13475 gnd.n7676 gnd.n90 240.244
R13476 gnd.n100 gnd.n90 240.244
R13477 gnd.n7670 gnd.n100 240.244
R13478 gnd.n7670 gnd.n101 240.244
R13479 gnd.n7662 gnd.n101 240.244
R13480 gnd.n7662 gnd.n117 240.244
R13481 gnd.n7658 gnd.n117 240.244
R13482 gnd.n7658 gnd.n122 240.244
R13483 gnd.n7650 gnd.n122 240.244
R13484 gnd.n7650 gnd.n136 240.244
R13485 gnd.n7646 gnd.n136 240.244
R13486 gnd.n7646 gnd.n142 240.244
R13487 gnd.n7638 gnd.n142 240.244
R13488 gnd.n7638 gnd.n156 240.244
R13489 gnd.n7634 gnd.n156 240.244
R13490 gnd.n7634 gnd.n162 240.244
R13491 gnd.n7626 gnd.n162 240.244
R13492 gnd.n7626 gnd.n176 240.244
R13493 gnd.n7622 gnd.n176 240.244
R13494 gnd.n7622 gnd.n182 240.244
R13495 gnd.n7614 gnd.n182 240.244
R13496 gnd.n7614 gnd.n195 240.244
R13497 gnd.n7610 gnd.n195 240.244
R13498 gnd.n7610 gnd.n201 240.244
R13499 gnd.n7602 gnd.n201 240.244
R13500 gnd.n4827 gnd.n1377 240.244
R13501 gnd.n4825 gnd.n4824 240.244
R13502 gnd.n4822 gnd.n1383 240.244
R13503 gnd.n4818 gnd.n4817 240.244
R13504 gnd.n4815 gnd.n1391 240.244
R13505 gnd.n4811 gnd.n4810 240.244
R13506 gnd.n4808 gnd.n1398 240.244
R13507 gnd.n4804 gnd.n4803 240.244
R13508 gnd.n4801 gnd.n1405 240.244
R13509 gnd.n4796 gnd.n4795 240.244
R13510 gnd.n4793 gnd.n1414 240.244
R13511 gnd.n4789 gnd.n4788 240.244
R13512 gnd.n4786 gnd.n1421 240.244
R13513 gnd.n2479 gnd.n2478 240.244
R13514 gnd.n2482 gnd.n2481 240.244
R13515 gnd.n2489 gnd.n2488 240.244
R13516 gnd.n2492 gnd.n2491 240.244
R13517 gnd.n2499 gnd.n2498 240.244
R13518 gnd.n2502 gnd.n2501 240.244
R13519 gnd.n2509 gnd.n2508 240.244
R13520 gnd.n2512 gnd.n2511 240.244
R13521 gnd.n2519 gnd.n2518 240.244
R13522 gnd.n2522 gnd.n2521 240.244
R13523 gnd.n2529 gnd.n2528 240.244
R13524 gnd.n2532 gnd.n2531 240.244
R13525 gnd.n2539 gnd.n2538 240.244
R13526 gnd.n2542 gnd.n2541 240.244
R13527 gnd.n2549 gnd.n2548 240.244
R13528 gnd.n4970 gnd.n4969 240.244
R13529 gnd.n4969 gnd.n1141 240.244
R13530 gnd.n1153 gnd.n1141 240.244
R13531 gnd.n2829 gnd.n1153 240.244
R13532 gnd.n2829 gnd.n1165 240.244
R13533 gnd.n2833 gnd.n1165 240.244
R13534 gnd.n2833 gnd.n1175 240.244
R13535 gnd.n2836 gnd.n1175 240.244
R13536 gnd.n2836 gnd.n1185 240.244
R13537 gnd.n2841 gnd.n1185 240.244
R13538 gnd.n2841 gnd.n1195 240.244
R13539 gnd.n2852 gnd.n1195 240.244
R13540 gnd.n2852 gnd.n1205 240.244
R13541 gnd.n2735 gnd.n1205 240.244
R13542 gnd.n2735 gnd.n1215 240.244
R13543 gnd.n2883 gnd.n1215 240.244
R13544 gnd.n2883 gnd.n1225 240.244
R13545 gnd.n2879 gnd.n1225 240.244
R13546 gnd.n2879 gnd.n1236 240.244
R13547 gnd.n2871 gnd.n1236 240.244
R13548 gnd.n2871 gnd.n1246 240.244
R13549 gnd.n2708 gnd.n1246 240.244
R13550 gnd.n2924 gnd.n2708 240.244
R13551 gnd.n2924 gnd.n2698 240.244
R13552 gnd.n2698 gnd.n2691 240.244
R13553 gnd.n2949 gnd.n2691 240.244
R13554 gnd.n2949 gnd.n2680 240.244
R13555 gnd.n2952 gnd.n2680 240.244
R13556 gnd.n2952 gnd.n2674 240.244
R13557 gnd.n2674 gnd.n2668 240.244
R13558 gnd.n2668 gnd.n1263 240.244
R13559 gnd.n3005 gnd.n1263 240.244
R13560 gnd.n3005 gnd.n1275 240.244
R13561 gnd.n3010 gnd.n1275 240.244
R13562 gnd.n3010 gnd.n1284 240.244
R13563 gnd.n3020 gnd.n1284 240.244
R13564 gnd.n3020 gnd.n1294 240.244
R13565 gnd.n2648 gnd.n1294 240.244
R13566 gnd.n2648 gnd.n1304 240.244
R13567 gnd.n3027 gnd.n1304 240.244
R13568 gnd.n3027 gnd.n1314 240.244
R13569 gnd.n3033 gnd.n1314 240.244
R13570 gnd.n3033 gnd.n1324 240.244
R13571 gnd.n3037 gnd.n1324 240.244
R13572 gnd.n3037 gnd.n1334 240.244
R13573 gnd.n3122 gnd.n1334 240.244
R13574 gnd.n3122 gnd.n1344 240.244
R13575 gnd.n3126 gnd.n1344 240.244
R13576 gnd.n3126 gnd.n1354 240.244
R13577 gnd.n3137 gnd.n1354 240.244
R13578 gnd.n3137 gnd.n1365 240.244
R13579 gnd.n3142 gnd.n1365 240.244
R13580 gnd.n3142 gnd.n1374 240.244
R13581 gnd.n1070 gnd.n1069 240.244
R13582 gnd.n5085 gnd.n1069 240.244
R13583 gnd.n5083 gnd.n5082 240.244
R13584 gnd.n5079 gnd.n5078 240.244
R13585 gnd.n5075 gnd.n5074 240.244
R13586 gnd.n5071 gnd.n5070 240.244
R13587 gnd.n5067 gnd.n5066 240.244
R13588 gnd.n5063 gnd.n5062 240.244
R13589 gnd.n5059 gnd.n5058 240.244
R13590 gnd.n5054 gnd.n5053 240.244
R13591 gnd.n5050 gnd.n5049 240.244
R13592 gnd.n5046 gnd.n5045 240.244
R13593 gnd.n5042 gnd.n5041 240.244
R13594 gnd.n5038 gnd.n5037 240.244
R13595 gnd.n5034 gnd.n5033 240.244
R13596 gnd.n5030 gnd.n5029 240.244
R13597 gnd.n5026 gnd.n5025 240.244
R13598 gnd.n5022 gnd.n5021 240.244
R13599 gnd.n5018 gnd.n5017 240.244
R13600 gnd.n5014 gnd.n5013 240.244
R13601 gnd.n5010 gnd.n5009 240.244
R13602 gnd.n5006 gnd.n5005 240.244
R13603 gnd.n5002 gnd.n5001 240.244
R13604 gnd.n4998 gnd.n4997 240.244
R13605 gnd.n4994 gnd.n4993 240.244
R13606 gnd.n4990 gnd.n4989 240.244
R13607 gnd.n4986 gnd.n4985 240.244
R13608 gnd.n4982 gnd.n4981 240.244
R13609 gnd.n4978 gnd.n4977 240.244
R13610 gnd.n4967 gnd.n1071 240.244
R13611 gnd.n4967 gnd.n1144 240.244
R13612 gnd.n4963 gnd.n1144 240.244
R13613 gnd.n4963 gnd.n1151 240.244
R13614 gnd.n4955 gnd.n1151 240.244
R13615 gnd.n4955 gnd.n1168 240.244
R13616 gnd.n4951 gnd.n1168 240.244
R13617 gnd.n4951 gnd.n1174 240.244
R13618 gnd.n4943 gnd.n1174 240.244
R13619 gnd.n4943 gnd.n1187 240.244
R13620 gnd.n4939 gnd.n1187 240.244
R13621 gnd.n4939 gnd.n1193 240.244
R13622 gnd.n4931 gnd.n1193 240.244
R13623 gnd.n4931 gnd.n1208 240.244
R13624 gnd.n4927 gnd.n1208 240.244
R13625 gnd.n4927 gnd.n1214 240.244
R13626 gnd.n4919 gnd.n1214 240.244
R13627 gnd.n4919 gnd.n1228 240.244
R13628 gnd.n4915 gnd.n1228 240.244
R13629 gnd.n4915 gnd.n1234 240.244
R13630 gnd.n4907 gnd.n1234 240.244
R13631 gnd.n4907 gnd.n1249 240.244
R13632 gnd.n2701 gnd.n1249 240.244
R13633 gnd.n2933 gnd.n2701 240.244
R13634 gnd.n2933 gnd.n2932 240.244
R13635 gnd.n2932 gnd.n2676 240.244
R13636 gnd.n2962 gnd.n2676 240.244
R13637 gnd.n2963 gnd.n2962 240.244
R13638 gnd.n2966 gnd.n2963 240.244
R13639 gnd.n2966 gnd.n1261 240.244
R13640 gnd.n4901 gnd.n1261 240.244
R13641 gnd.n4901 gnd.n1262 240.244
R13642 gnd.n4893 gnd.n1262 240.244
R13643 gnd.n4893 gnd.n1277 240.244
R13644 gnd.n4889 gnd.n1277 240.244
R13645 gnd.n4889 gnd.n1282 240.244
R13646 gnd.n4881 gnd.n1282 240.244
R13647 gnd.n4881 gnd.n1297 240.244
R13648 gnd.n4877 gnd.n1297 240.244
R13649 gnd.n4877 gnd.n1303 240.244
R13650 gnd.n4869 gnd.n1303 240.244
R13651 gnd.n4869 gnd.n1316 240.244
R13652 gnd.n4865 gnd.n1316 240.244
R13653 gnd.n4865 gnd.n1322 240.244
R13654 gnd.n4857 gnd.n1322 240.244
R13655 gnd.n4857 gnd.n1337 240.244
R13656 gnd.n4853 gnd.n1337 240.244
R13657 gnd.n4853 gnd.n1343 240.244
R13658 gnd.n4845 gnd.n1343 240.244
R13659 gnd.n4845 gnd.n1357 240.244
R13660 gnd.n4841 gnd.n1357 240.244
R13661 gnd.n4841 gnd.n1363 240.244
R13662 gnd.n4833 gnd.n1363 240.244
R13663 gnd.n5100 gnd.n5095 240.244
R13664 gnd.n6465 gnd.n6464 240.244
R13665 gnd.n6462 gnd.n5104 240.244
R13666 gnd.n6458 gnd.n6457 240.244
R13667 gnd.n6455 gnd.n5111 240.244
R13668 gnd.n6451 gnd.n6450 240.244
R13669 gnd.n6448 gnd.n5118 240.244
R13670 gnd.n6444 gnd.n6443 240.244
R13671 gnd.n5735 gnd.n5455 240.244
R13672 gnd.n5455 gnd.n5446 240.244
R13673 gnd.n5753 gnd.n5446 240.244
R13674 gnd.n5754 gnd.n5753 240.244
R13675 gnd.n5754 gnd.n5434 240.244
R13676 gnd.n5434 gnd.n5423 240.244
R13677 gnd.n5785 gnd.n5423 240.244
R13678 gnd.n5786 gnd.n5785 240.244
R13679 gnd.n5787 gnd.n5786 240.244
R13680 gnd.n5787 gnd.n5408 240.244
R13681 gnd.n5789 gnd.n5408 240.244
R13682 gnd.n5789 gnd.n5393 240.244
R13683 gnd.n5830 gnd.n5393 240.244
R13684 gnd.n5831 gnd.n5830 240.244
R13685 gnd.n5834 gnd.n5831 240.244
R13686 gnd.n5834 gnd.n5375 240.244
R13687 gnd.n5866 gnd.n5375 240.244
R13688 gnd.n5866 gnd.n5361 240.244
R13689 gnd.n5888 gnd.n5361 240.244
R13690 gnd.n5889 gnd.n5888 240.244
R13691 gnd.n5889 gnd.n5348 240.244
R13692 gnd.n5348 gnd.n5337 240.244
R13693 gnd.n5920 gnd.n5337 240.244
R13694 gnd.n5921 gnd.n5920 240.244
R13695 gnd.n5922 gnd.n5921 240.244
R13696 gnd.n5922 gnd.n5258 240.244
R13697 gnd.n5258 gnd.n5257 240.244
R13698 gnd.n5257 gnd.n5242 240.244
R13699 gnd.n5973 gnd.n5242 240.244
R13700 gnd.n5974 gnd.n5973 240.244
R13701 gnd.n5974 gnd.n5229 240.244
R13702 gnd.n5229 gnd.n5218 240.244
R13703 gnd.n6007 gnd.n5218 240.244
R13704 gnd.n6008 gnd.n6007 240.244
R13705 gnd.n6010 gnd.n6008 240.244
R13706 gnd.n6010 gnd.n6009 240.244
R13707 gnd.n6009 gnd.n5198 240.244
R13708 gnd.n6047 gnd.n5198 240.244
R13709 gnd.n6047 gnd.n5185 240.244
R13710 gnd.n6073 gnd.n5185 240.244
R13711 gnd.n6074 gnd.n6073 240.244
R13712 gnd.n6075 gnd.n6074 240.244
R13713 gnd.n6075 gnd.n981 240.244
R13714 gnd.n6364 gnd.n981 240.244
R13715 gnd.n6364 gnd.n991 240.244
R13716 gnd.n6360 gnd.n991 240.244
R13717 gnd.n6360 gnd.n6359 240.244
R13718 gnd.n6359 gnd.n1004 240.244
R13719 gnd.n6355 gnd.n1004 240.244
R13720 gnd.n6355 gnd.n1017 240.244
R13721 gnd.n6351 gnd.n1017 240.244
R13722 gnd.n6351 gnd.n6350 240.244
R13723 gnd.n6350 gnd.n1029 240.244
R13724 gnd.n5672 gnd.n5671 240.244
R13725 gnd.n5716 gnd.n5671 240.244
R13726 gnd.n5714 gnd.n5713 240.244
R13727 gnd.n5710 gnd.n5709 240.244
R13728 gnd.n5706 gnd.n5705 240.244
R13729 gnd.n5702 gnd.n5701 240.244
R13730 gnd.n5698 gnd.n5697 240.244
R13731 gnd.n5694 gnd.n5693 240.244
R13732 gnd.n5745 gnd.n5453 240.244
R13733 gnd.n5745 gnd.n5449 240.244
R13734 gnd.n5751 gnd.n5449 240.244
R13735 gnd.n5751 gnd.n5432 240.244
R13736 gnd.n5775 gnd.n5432 240.244
R13737 gnd.n5775 gnd.n5427 240.244
R13738 gnd.n5783 gnd.n5427 240.244
R13739 gnd.n5783 gnd.n5428 240.244
R13740 gnd.n5428 gnd.n5406 240.244
R13741 gnd.n5809 gnd.n5406 240.244
R13742 gnd.n5809 gnd.n5401 240.244
R13743 gnd.n5820 gnd.n5401 240.244
R13744 gnd.n5820 gnd.n5402 240.244
R13745 gnd.n5816 gnd.n5402 240.244
R13746 gnd.n5816 gnd.n5373 240.244
R13747 gnd.n5870 gnd.n5373 240.244
R13748 gnd.n5870 gnd.n5368 240.244
R13749 gnd.n5878 gnd.n5368 240.244
R13750 gnd.n5878 gnd.n5369 240.244
R13751 gnd.n5369 gnd.n5346 240.244
R13752 gnd.n5910 gnd.n5346 240.244
R13753 gnd.n5910 gnd.n5341 240.244
R13754 gnd.n5918 gnd.n5341 240.244
R13755 gnd.n5918 gnd.n5342 240.244
R13756 gnd.n5342 gnd.n5255 240.244
R13757 gnd.n5955 gnd.n5255 240.244
R13758 gnd.n5955 gnd.n5250 240.244
R13759 gnd.n5963 gnd.n5250 240.244
R13760 gnd.n5963 gnd.n5251 240.244
R13761 gnd.n5251 gnd.n5227 240.244
R13762 gnd.n5994 gnd.n5227 240.244
R13763 gnd.n5994 gnd.n5222 240.244
R13764 gnd.n6005 gnd.n5222 240.244
R13765 gnd.n6005 gnd.n5223 240.244
R13766 gnd.n6001 gnd.n5223 240.244
R13767 gnd.n6001 gnd.n5197 240.244
R13768 gnd.n6051 gnd.n5197 240.244
R13769 gnd.n6051 gnd.n5192 240.244
R13770 gnd.n6063 gnd.n5192 240.244
R13771 gnd.n6063 gnd.n5193 240.244
R13772 gnd.n6059 gnd.n5193 240.244
R13773 gnd.n6059 gnd.n982 240.244
R13774 gnd.n6500 gnd.n982 240.244
R13775 gnd.n6500 gnd.n983 240.244
R13776 gnd.n6496 gnd.n983 240.244
R13777 gnd.n6496 gnd.n989 240.244
R13778 gnd.n1006 gnd.n989 240.244
R13779 gnd.n6486 gnd.n1006 240.244
R13780 gnd.n6486 gnd.n1007 240.244
R13781 gnd.n6482 gnd.n1007 240.244
R13782 gnd.n6482 gnd.n1015 240.244
R13783 gnd.n5094 gnd.n1015 240.244
R13784 gnd.n6472 gnd.n5094 240.244
R13785 gnd.n319 gnd.n208 240.244
R13786 gnd.n7485 gnd.n7484 240.244
R13787 gnd.n7482 gnd.n323 240.244
R13788 gnd.n7478 gnd.n7477 240.244
R13789 gnd.n7475 gnd.n330 240.244
R13790 gnd.n7471 gnd.n7470 240.244
R13791 gnd.n7468 gnd.n337 240.244
R13792 gnd.n7464 gnd.n7463 240.244
R13793 gnd.n7461 gnd.n344 240.244
R13794 gnd.n1971 gnd.n1787 240.244
R13795 gnd.n1971 gnd.n1797 240.244
R13796 gnd.n4190 gnd.n1797 240.244
R13797 gnd.n4190 gnd.n1813 240.244
R13798 gnd.n4196 gnd.n1813 240.244
R13799 gnd.n4196 gnd.n1826 240.244
R13800 gnd.n4205 gnd.n1826 240.244
R13801 gnd.n4205 gnd.n1836 240.244
R13802 gnd.n4211 gnd.n1836 240.244
R13803 gnd.n4211 gnd.n1846 240.244
R13804 gnd.n4247 gnd.n1846 240.244
R13805 gnd.n4247 gnd.n1856 240.244
R13806 gnd.n1958 gnd.n1856 240.244
R13807 gnd.n1958 gnd.n1866 240.244
R13808 gnd.n1959 gnd.n1866 240.244
R13809 gnd.n1959 gnd.n1876 240.244
R13810 gnd.n4235 gnd.n1876 240.244
R13811 gnd.n4235 gnd.n1886 240.244
R13812 gnd.n4274 gnd.n1886 240.244
R13813 gnd.n4274 gnd.n1896 240.244
R13814 gnd.n4288 gnd.n1896 240.244
R13815 gnd.n4288 gnd.n1906 240.244
R13816 gnd.n1911 gnd.n1906 240.244
R13817 gnd.n4279 gnd.n1911 240.244
R13818 gnd.n4279 gnd.n1929 240.244
R13819 gnd.n1929 gnd.n1923 240.244
R13820 gnd.n1923 gnd.n82 240.244
R13821 gnd.n7678 gnd.n82 240.244
R13822 gnd.n7678 gnd.n84 240.244
R13823 gnd.n7373 gnd.n84 240.244
R13824 gnd.n7373 gnd.n104 240.244
R13825 gnd.n7381 gnd.n104 240.244
R13826 gnd.n7381 gnd.n116 240.244
R13827 gnd.n7387 gnd.n116 240.244
R13828 gnd.n7387 gnd.n125 240.244
R13829 gnd.n7395 gnd.n125 240.244
R13830 gnd.n7395 gnd.n134 240.244
R13831 gnd.n7401 gnd.n134 240.244
R13832 gnd.n7401 gnd.n145 240.244
R13833 gnd.n7409 gnd.n145 240.244
R13834 gnd.n7409 gnd.n155 240.244
R13835 gnd.n7416 gnd.n155 240.244
R13836 gnd.n7416 gnd.n165 240.244
R13837 gnd.n7439 gnd.n165 240.244
R13838 gnd.n7439 gnd.n174 240.244
R13839 gnd.n356 gnd.n174 240.244
R13840 gnd.n356 gnd.n184 240.244
R13841 gnd.n7446 gnd.n184 240.244
R13842 gnd.n7446 gnd.n193 240.244
R13843 gnd.n353 gnd.n193 240.244
R13844 gnd.n353 gnd.n203 240.244
R13845 gnd.n7453 gnd.n203 240.244
R13846 gnd.n7453 gnd.n211 240.244
R13847 gnd.n1631 gnd.n1630 240.244
R13848 gnd.n1706 gnd.n1638 240.244
R13849 gnd.n1709 gnd.n1639 240.244
R13850 gnd.n1647 gnd.n1646 240.244
R13851 gnd.n1711 gnd.n1654 240.244
R13852 gnd.n1714 gnd.n1655 240.244
R13853 gnd.n1663 gnd.n1662 240.244
R13854 gnd.n1716 gnd.n1672 240.244
R13855 gnd.n4522 gnd.n1675 240.244
R13856 gnd.n4398 gnd.n1790 240.244
R13857 gnd.n1799 gnd.n1790 240.244
R13858 gnd.n1815 gnd.n1799 240.244
R13859 gnd.n4384 gnd.n1815 240.244
R13860 gnd.n4384 gnd.n1816 240.244
R13861 gnd.n4380 gnd.n1816 240.244
R13862 gnd.n4380 gnd.n1823 240.244
R13863 gnd.n4372 gnd.n1823 240.244
R13864 gnd.n4372 gnd.n1838 240.244
R13865 gnd.n4368 gnd.n1838 240.244
R13866 gnd.n4368 gnd.n1843 240.244
R13867 gnd.n4360 gnd.n1843 240.244
R13868 gnd.n4360 gnd.n1858 240.244
R13869 gnd.n4356 gnd.n1858 240.244
R13870 gnd.n4356 gnd.n1863 240.244
R13871 gnd.n4348 gnd.n1863 240.244
R13872 gnd.n4348 gnd.n1878 240.244
R13873 gnd.n4344 gnd.n1878 240.244
R13874 gnd.n4344 gnd.n1883 240.244
R13875 gnd.n4336 gnd.n1883 240.244
R13876 gnd.n4336 gnd.n1898 240.244
R13877 gnd.n4332 gnd.n1898 240.244
R13878 gnd.n4332 gnd.n1903 240.244
R13879 gnd.n1930 gnd.n1903 240.244
R13880 gnd.n4312 gnd.n1930 240.244
R13881 gnd.n4312 gnd.n1925 240.244
R13882 gnd.n4308 gnd.n1925 240.244
R13883 gnd.n4308 gnd.n88 240.244
R13884 gnd.n4300 gnd.n88 240.244
R13885 gnd.n4300 gnd.n106 240.244
R13886 gnd.n7668 gnd.n106 240.244
R13887 gnd.n7668 gnd.n107 240.244
R13888 gnd.n7664 gnd.n107 240.244
R13889 gnd.n7664 gnd.n113 240.244
R13890 gnd.n7656 gnd.n113 240.244
R13891 gnd.n7656 gnd.n126 240.244
R13892 gnd.n7652 gnd.n126 240.244
R13893 gnd.n7652 gnd.n131 240.244
R13894 gnd.n7644 gnd.n131 240.244
R13895 gnd.n7644 gnd.n147 240.244
R13896 gnd.n7640 gnd.n147 240.244
R13897 gnd.n7640 gnd.n152 240.244
R13898 gnd.n7632 gnd.n152 240.244
R13899 gnd.n7632 gnd.n166 240.244
R13900 gnd.n7628 gnd.n166 240.244
R13901 gnd.n7628 gnd.n171 240.244
R13902 gnd.n7620 gnd.n171 240.244
R13903 gnd.n7620 gnd.n186 240.244
R13904 gnd.n7616 gnd.n186 240.244
R13905 gnd.n7616 gnd.n191 240.244
R13906 gnd.n7608 gnd.n191 240.244
R13907 gnd.n7608 gnd.n204 240.244
R13908 gnd.n7604 gnd.n204 240.244
R13909 gnd.n5130 gnd.n1026 240.244
R13910 gnd.n6433 gnd.n6432 240.244
R13911 gnd.n6430 gnd.n5134 240.244
R13912 gnd.n6426 gnd.n6425 240.244
R13913 gnd.n6423 gnd.n5141 240.244
R13914 gnd.n6419 gnd.n6418 240.244
R13915 gnd.n6416 gnd.n5148 240.244
R13916 gnd.n6412 gnd.n6411 240.244
R13917 gnd.n6409 gnd.n5155 240.244
R13918 gnd.n6405 gnd.n6404 240.244
R13919 gnd.n6402 gnd.n5162 240.244
R13920 gnd.n6398 gnd.n6397 240.244
R13921 gnd.n6395 gnd.n5172 240.244
R13922 gnd.n5603 gnd.n5499 240.244
R13923 gnd.n5609 gnd.n5499 240.244
R13924 gnd.n5609 gnd.n5491 240.244
R13925 gnd.n5619 gnd.n5491 240.244
R13926 gnd.n5619 gnd.n5487 240.244
R13927 gnd.n5625 gnd.n5487 240.244
R13928 gnd.n5625 gnd.n5478 240.244
R13929 gnd.n5635 gnd.n5478 240.244
R13930 gnd.n5635 gnd.n5473 240.244
R13931 gnd.n5663 gnd.n5473 240.244
R13932 gnd.n5663 gnd.n5474 240.244
R13933 gnd.n5474 gnd.n5466 240.244
R13934 gnd.n5658 gnd.n5466 240.244
R13935 gnd.n5658 gnd.n5456 240.244
R13936 gnd.n5655 gnd.n5456 240.244
R13937 gnd.n5655 gnd.n5445 240.244
R13938 gnd.n5652 gnd.n5445 240.244
R13939 gnd.n5652 gnd.n5435 240.244
R13940 gnd.n5649 gnd.n5435 240.244
R13941 gnd.n5649 gnd.n5413 240.244
R13942 gnd.n5798 gnd.n5413 240.244
R13943 gnd.n5798 gnd.n5409 240.244
R13944 gnd.n5806 gnd.n5409 240.244
R13945 gnd.n5806 gnd.n5399 240.244
R13946 gnd.n5399 gnd.n5380 240.244
R13947 gnd.n5845 gnd.n5380 240.244
R13948 gnd.n5845 gnd.n5381 240.244
R13949 gnd.n5381 gnd.n5376 240.244
R13950 gnd.n5865 gnd.n5376 240.244
R13951 gnd.n5865 gnd.n5366 240.244
R13952 gnd.n5860 gnd.n5366 240.244
R13953 gnd.n5860 gnd.n5360 240.244
R13954 gnd.n5856 gnd.n5360 240.244
R13955 gnd.n5856 gnd.n5349 240.244
R13956 gnd.n5852 gnd.n5349 240.244
R13957 gnd.n5852 gnd.n5327 240.244
R13958 gnd.n5931 gnd.n5327 240.244
R13959 gnd.n5931 gnd.n5259 240.244
R13960 gnd.n5952 gnd.n5259 240.244
R13961 gnd.n5952 gnd.n5248 240.244
R13962 gnd.n5948 gnd.n5248 240.244
R13963 gnd.n5948 gnd.n5241 240.244
R13964 gnd.n5945 gnd.n5241 240.244
R13965 gnd.n5945 gnd.n5230 240.244
R13966 gnd.n5942 gnd.n5230 240.244
R13967 gnd.n5942 gnd.n5209 240.244
R13968 gnd.n6017 gnd.n5209 240.244
R13969 gnd.n6017 gnd.n5205 240.244
R13970 gnd.n6038 gnd.n5205 240.244
R13971 gnd.n6038 gnd.n5199 240.244
R13972 gnd.n5199 gnd.n5190 240.244
R13973 gnd.n6033 gnd.n5190 240.244
R13974 gnd.n6033 gnd.n969 240.244
R13975 gnd.n6030 gnd.n969 240.244
R13976 gnd.n6030 gnd.n980 240.244
R13977 gnd.n6367 gnd.n980 240.244
R13978 gnd.n6368 gnd.n6367 240.244
R13979 gnd.n6368 gnd.n992 240.244
R13980 gnd.n6374 gnd.n992 240.244
R13981 gnd.n6374 gnd.n1003 240.244
R13982 gnd.n6378 gnd.n1003 240.244
R13983 gnd.n6378 gnd.n6377 240.244
R13984 gnd.n6377 gnd.n1018 240.244
R13985 gnd.n6385 gnd.n1018 240.244
R13986 gnd.n6385 gnd.n1028 240.244
R13987 gnd.n5595 gnd.n5593 240.244
R13988 gnd.n5593 gnd.n5592 240.244
R13989 gnd.n5589 gnd.n5588 240.244
R13990 gnd.n5586 gnd.n5512 240.244
R13991 gnd.n5582 gnd.n5580 240.244
R13992 gnd.n5578 gnd.n5518 240.244
R13993 gnd.n5574 gnd.n5572 240.244
R13994 gnd.n5570 gnd.n5524 240.244
R13995 gnd.n5566 gnd.n5564 240.244
R13996 gnd.n5562 gnd.n5530 240.244
R13997 gnd.n5558 gnd.n5556 240.244
R13998 gnd.n5554 gnd.n5536 240.244
R13999 gnd.n5549 gnd.n5547 240.244
R14000 gnd.n5601 gnd.n5497 240.244
R14001 gnd.n5611 gnd.n5497 240.244
R14002 gnd.n5611 gnd.n5493 240.244
R14003 gnd.n5617 gnd.n5493 240.244
R14004 gnd.n5617 gnd.n5485 240.244
R14005 gnd.n5627 gnd.n5485 240.244
R14006 gnd.n5627 gnd.n5481 240.244
R14007 gnd.n5633 gnd.n5481 240.244
R14008 gnd.n5633 gnd.n5472 240.244
R14009 gnd.n5725 gnd.n5472 240.244
R14010 gnd.n5725 gnd.n5467 240.244
R14011 gnd.n5732 gnd.n5467 240.244
R14012 gnd.n5732 gnd.n5458 240.244
R14013 gnd.n5742 gnd.n5458 240.244
R14014 gnd.n5742 gnd.n5444 240.244
R14015 gnd.n5757 gnd.n5444 240.244
R14016 gnd.n5757 gnd.n5437 240.244
R14017 gnd.n5772 gnd.n5437 240.244
R14018 gnd.n5772 gnd.n5438 240.244
R14019 gnd.n5438 gnd.n5416 240.244
R14020 gnd.n5796 gnd.n5416 240.244
R14021 gnd.n5796 gnd.n5417 240.244
R14022 gnd.n5417 gnd.n5397 240.244
R14023 gnd.n5823 gnd.n5397 240.244
R14024 gnd.n5823 gnd.n5384 240.244
R14025 gnd.n5843 gnd.n5384 240.244
R14026 gnd.n5843 gnd.n5385 240.244
R14027 gnd.n5839 gnd.n5385 240.244
R14028 gnd.n5839 gnd.n5365 240.244
R14029 gnd.n5881 gnd.n5365 240.244
R14030 gnd.n5881 gnd.n5358 240.244
R14031 gnd.n5892 gnd.n5358 240.244
R14032 gnd.n5892 gnd.n5351 240.244
R14033 gnd.n5907 gnd.n5351 240.244
R14034 gnd.n5907 gnd.n5352 240.244
R14035 gnd.n5352 gnd.n5330 240.244
R14036 gnd.n5929 gnd.n5330 240.244
R14037 gnd.n5929 gnd.n5331 240.244
R14038 gnd.n5331 gnd.n5246 240.244
R14039 gnd.n5966 gnd.n5246 240.244
R14040 gnd.n5966 gnd.n5239 240.244
R14041 gnd.n5977 gnd.n5239 240.244
R14042 gnd.n5977 gnd.n5232 240.244
R14043 gnd.n5991 gnd.n5232 240.244
R14044 gnd.n5991 gnd.n5233 240.244
R14045 gnd.n5233 gnd.n5213 240.244
R14046 gnd.n6015 gnd.n5213 240.244
R14047 gnd.n6015 gnd.n5203 240.244
R14048 gnd.n6040 gnd.n5203 240.244
R14049 gnd.n6040 gnd.n5189 240.244
R14050 gnd.n6066 gnd.n5189 240.244
R14051 gnd.n6066 gnd.n971 240.244
R14052 gnd.n6507 gnd.n971 240.244
R14053 gnd.n6507 gnd.n972 240.244
R14054 gnd.n6503 gnd.n972 240.244
R14055 gnd.n6503 gnd.n978 240.244
R14056 gnd.n994 gnd.n978 240.244
R14057 gnd.n6493 gnd.n994 240.244
R14058 gnd.n6493 gnd.n995 240.244
R14059 gnd.n6489 gnd.n995 240.244
R14060 gnd.n6489 gnd.n1001 240.244
R14061 gnd.n1020 gnd.n1001 240.244
R14062 gnd.n6479 gnd.n1020 240.244
R14063 gnd.n6479 gnd.n1021 240.244
R14064 gnd.n6475 gnd.n1021 240.244
R14065 gnd.n2561 gnd.n1372 240.244
R14066 gnd.n2572 gnd.n2563 240.244
R14067 gnd.n2575 gnd.n2574 240.244
R14068 gnd.n2584 gnd.n2583 240.244
R14069 gnd.n2595 gnd.n2586 240.244
R14070 gnd.n2598 gnd.n2597 240.244
R14071 gnd.n2607 gnd.n2606 240.244
R14072 gnd.n2619 gnd.n2609 240.244
R14073 gnd.n2625 gnd.n2621 240.244
R14074 gnd.n2807 gnd.n1142 240.244
R14075 gnd.n2810 gnd.n1142 240.244
R14076 gnd.n2810 gnd.n1154 240.244
R14077 gnd.n2815 gnd.n1154 240.244
R14078 gnd.n2815 gnd.n1166 240.244
R14079 gnd.n2818 gnd.n1166 240.244
R14080 gnd.n2818 gnd.n1176 240.244
R14081 gnd.n2823 gnd.n1176 240.244
R14082 gnd.n2823 gnd.n1186 240.244
R14083 gnd.n2843 gnd.n1186 240.244
R14084 gnd.n2843 gnd.n1196 240.244
R14085 gnd.n2850 gnd.n1196 240.244
R14086 gnd.n2850 gnd.n1206 240.244
R14087 gnd.n2889 gnd.n1206 240.244
R14088 gnd.n2889 gnd.n1216 240.244
R14089 gnd.n2885 gnd.n1216 240.244
R14090 gnd.n2885 gnd.n1226 240.244
R14091 gnd.n2877 gnd.n1226 240.244
R14092 gnd.n2877 gnd.n1237 240.244
R14093 gnd.n2873 gnd.n1237 240.244
R14094 gnd.n2873 gnd.n1247 240.244
R14095 gnd.n2866 gnd.n1247 240.244
R14096 gnd.n2866 gnd.n2696 240.244
R14097 gnd.n2935 gnd.n2696 240.244
R14098 gnd.n2935 gnd.n2692 240.244
R14099 gnd.n2947 gnd.n2692 240.244
R14100 gnd.n2947 gnd.n2681 240.244
R14101 gnd.n2940 gnd.n2681 240.244
R14102 gnd.n2940 gnd.n2666 240.244
R14103 gnd.n2997 gnd.n2666 240.244
R14104 gnd.n2997 gnd.n1264 240.244
R14105 gnd.n3003 gnd.n1264 240.244
R14106 gnd.n3003 gnd.n1276 240.244
R14107 gnd.n3012 gnd.n1276 240.244
R14108 gnd.n3012 gnd.n1285 240.244
R14109 gnd.n3018 gnd.n1285 240.244
R14110 gnd.n3018 gnd.n1295 240.244
R14111 gnd.n3054 gnd.n1295 240.244
R14112 gnd.n3054 gnd.n1305 240.244
R14113 gnd.n2653 gnd.n1305 240.244
R14114 gnd.n2653 gnd.n1315 240.244
R14115 gnd.n2654 gnd.n1315 240.244
R14116 gnd.n2654 gnd.n1325 240.244
R14117 gnd.n3039 gnd.n1325 240.244
R14118 gnd.n3039 gnd.n1335 240.244
R14119 gnd.n2636 gnd.n1335 240.244
R14120 gnd.n2636 gnd.n1345 240.244
R14121 gnd.n3128 gnd.n1345 240.244
R14122 gnd.n3128 gnd.n1355 240.244
R14123 gnd.n3135 gnd.n1355 240.244
R14124 gnd.n3135 gnd.n1366 240.244
R14125 gnd.n3144 gnd.n1366 240.244
R14126 gnd.n3144 gnd.n1375 240.244
R14127 gnd.n2767 gnd.n2766 240.244
R14128 gnd.n2773 gnd.n2772 240.244
R14129 gnd.n2777 gnd.n2776 240.244
R14130 gnd.n2783 gnd.n2782 240.244
R14131 gnd.n2787 gnd.n2786 240.244
R14132 gnd.n2793 gnd.n2792 240.244
R14133 gnd.n2797 gnd.n2796 240.244
R14134 gnd.n2754 gnd.n2753 240.244
R14135 gnd.n2749 gnd.n1067 240.244
R14136 gnd.n2762 gnd.n1143 240.244
R14137 gnd.n1156 gnd.n1143 240.244
R14138 gnd.n4961 gnd.n1156 240.244
R14139 gnd.n4961 gnd.n1157 240.244
R14140 gnd.n4957 gnd.n1157 240.244
R14141 gnd.n4957 gnd.n1164 240.244
R14142 gnd.n4949 gnd.n1164 240.244
R14143 gnd.n4949 gnd.n1178 240.244
R14144 gnd.n4945 gnd.n1178 240.244
R14145 gnd.n4945 gnd.n1183 240.244
R14146 gnd.n4937 gnd.n1183 240.244
R14147 gnd.n4937 gnd.n1198 240.244
R14148 gnd.n4933 gnd.n1198 240.244
R14149 gnd.n4933 gnd.n1203 240.244
R14150 gnd.n4925 gnd.n1203 240.244
R14151 gnd.n4925 gnd.n1218 240.244
R14152 gnd.n4921 gnd.n1218 240.244
R14153 gnd.n4921 gnd.n1223 240.244
R14154 gnd.n4913 gnd.n1223 240.244
R14155 gnd.n4913 gnd.n1239 240.244
R14156 gnd.n4909 gnd.n1239 240.244
R14157 gnd.n4909 gnd.n1244 240.244
R14158 gnd.n2922 gnd.n1244 240.244
R14159 gnd.n2922 gnd.n2700 240.244
R14160 gnd.n2930 gnd.n2700 240.244
R14161 gnd.n2930 gnd.n2683 240.244
R14162 gnd.n2960 gnd.n2683 240.244
R14163 gnd.n2960 gnd.n2684 240.244
R14164 gnd.n2684 gnd.n2675 240.244
R14165 gnd.n2675 gnd.n1266 240.244
R14166 gnd.n4899 gnd.n1266 240.244
R14167 gnd.n4899 gnd.n1267 240.244
R14168 gnd.n4895 gnd.n1267 240.244
R14169 gnd.n4895 gnd.n1273 240.244
R14170 gnd.n4887 gnd.n1273 240.244
R14171 gnd.n4887 gnd.n1287 240.244
R14172 gnd.n4883 gnd.n1287 240.244
R14173 gnd.n4883 gnd.n1292 240.244
R14174 gnd.n4875 gnd.n1292 240.244
R14175 gnd.n4875 gnd.n1307 240.244
R14176 gnd.n4871 gnd.n1307 240.244
R14177 gnd.n4871 gnd.n1312 240.244
R14178 gnd.n4863 gnd.n1312 240.244
R14179 gnd.n4863 gnd.n1327 240.244
R14180 gnd.n4859 gnd.n1327 240.244
R14181 gnd.n4859 gnd.n1332 240.244
R14182 gnd.n4851 gnd.n1332 240.244
R14183 gnd.n4851 gnd.n1347 240.244
R14184 gnd.n4847 gnd.n1347 240.244
R14185 gnd.n4847 gnd.n1352 240.244
R14186 gnd.n4839 gnd.n1352 240.244
R14187 gnd.n4839 gnd.n1368 240.244
R14188 gnd.n4835 gnd.n1368 240.244
R14189 gnd.n6680 gnd.n800 240.244
R14190 gnd.n6680 gnd.n796 240.244
R14191 gnd.n6686 gnd.n796 240.244
R14192 gnd.n6686 gnd.n794 240.244
R14193 gnd.n6690 gnd.n794 240.244
R14194 gnd.n6690 gnd.n790 240.244
R14195 gnd.n6696 gnd.n790 240.244
R14196 gnd.n6696 gnd.n788 240.244
R14197 gnd.n6700 gnd.n788 240.244
R14198 gnd.n6700 gnd.n784 240.244
R14199 gnd.n6706 gnd.n784 240.244
R14200 gnd.n6706 gnd.n782 240.244
R14201 gnd.n6710 gnd.n782 240.244
R14202 gnd.n6710 gnd.n778 240.244
R14203 gnd.n6716 gnd.n778 240.244
R14204 gnd.n6716 gnd.n776 240.244
R14205 gnd.n6720 gnd.n776 240.244
R14206 gnd.n6720 gnd.n772 240.244
R14207 gnd.n6726 gnd.n772 240.244
R14208 gnd.n6726 gnd.n770 240.244
R14209 gnd.n6730 gnd.n770 240.244
R14210 gnd.n6730 gnd.n766 240.244
R14211 gnd.n6736 gnd.n766 240.244
R14212 gnd.n6736 gnd.n764 240.244
R14213 gnd.n6740 gnd.n764 240.244
R14214 gnd.n6740 gnd.n760 240.244
R14215 gnd.n6746 gnd.n760 240.244
R14216 gnd.n6746 gnd.n758 240.244
R14217 gnd.n6750 gnd.n758 240.244
R14218 gnd.n6750 gnd.n754 240.244
R14219 gnd.n6756 gnd.n754 240.244
R14220 gnd.n6756 gnd.n752 240.244
R14221 gnd.n6760 gnd.n752 240.244
R14222 gnd.n6760 gnd.n748 240.244
R14223 gnd.n6766 gnd.n748 240.244
R14224 gnd.n6766 gnd.n746 240.244
R14225 gnd.n6770 gnd.n746 240.244
R14226 gnd.n6770 gnd.n742 240.244
R14227 gnd.n6776 gnd.n742 240.244
R14228 gnd.n6776 gnd.n740 240.244
R14229 gnd.n6780 gnd.n740 240.244
R14230 gnd.n6780 gnd.n736 240.244
R14231 gnd.n6786 gnd.n736 240.244
R14232 gnd.n6786 gnd.n734 240.244
R14233 gnd.n6790 gnd.n734 240.244
R14234 gnd.n6790 gnd.n730 240.244
R14235 gnd.n6796 gnd.n730 240.244
R14236 gnd.n6796 gnd.n728 240.244
R14237 gnd.n6800 gnd.n728 240.244
R14238 gnd.n6800 gnd.n724 240.244
R14239 gnd.n6806 gnd.n724 240.244
R14240 gnd.n6806 gnd.n722 240.244
R14241 gnd.n6810 gnd.n722 240.244
R14242 gnd.n6810 gnd.n718 240.244
R14243 gnd.n6816 gnd.n718 240.244
R14244 gnd.n6816 gnd.n716 240.244
R14245 gnd.n6820 gnd.n716 240.244
R14246 gnd.n6820 gnd.n712 240.244
R14247 gnd.n6826 gnd.n712 240.244
R14248 gnd.n6826 gnd.n710 240.244
R14249 gnd.n6830 gnd.n710 240.244
R14250 gnd.n6830 gnd.n706 240.244
R14251 gnd.n6836 gnd.n706 240.244
R14252 gnd.n6836 gnd.n704 240.244
R14253 gnd.n6840 gnd.n704 240.244
R14254 gnd.n6840 gnd.n700 240.244
R14255 gnd.n6846 gnd.n700 240.244
R14256 gnd.n6846 gnd.n698 240.244
R14257 gnd.n6850 gnd.n698 240.244
R14258 gnd.n6850 gnd.n694 240.244
R14259 gnd.n6856 gnd.n694 240.244
R14260 gnd.n6856 gnd.n692 240.244
R14261 gnd.n6860 gnd.n692 240.244
R14262 gnd.n6860 gnd.n688 240.244
R14263 gnd.n6866 gnd.n688 240.244
R14264 gnd.n6866 gnd.n686 240.244
R14265 gnd.n6870 gnd.n686 240.244
R14266 gnd.n6870 gnd.n682 240.244
R14267 gnd.n6876 gnd.n682 240.244
R14268 gnd.n6876 gnd.n680 240.244
R14269 gnd.n6880 gnd.n680 240.244
R14270 gnd.n6880 gnd.n676 240.244
R14271 gnd.n6886 gnd.n676 240.244
R14272 gnd.n6886 gnd.n674 240.244
R14273 gnd.n6890 gnd.n674 240.244
R14274 gnd.n6890 gnd.n670 240.244
R14275 gnd.n6896 gnd.n670 240.244
R14276 gnd.n6896 gnd.n668 240.244
R14277 gnd.n6900 gnd.n668 240.244
R14278 gnd.n6900 gnd.n664 240.244
R14279 gnd.n6906 gnd.n664 240.244
R14280 gnd.n6906 gnd.n662 240.244
R14281 gnd.n6910 gnd.n662 240.244
R14282 gnd.n6910 gnd.n658 240.244
R14283 gnd.n6916 gnd.n658 240.244
R14284 gnd.n6916 gnd.n656 240.244
R14285 gnd.n6920 gnd.n656 240.244
R14286 gnd.n6920 gnd.n652 240.244
R14287 gnd.n6926 gnd.n652 240.244
R14288 gnd.n6926 gnd.n650 240.244
R14289 gnd.n6930 gnd.n650 240.244
R14290 gnd.n6930 gnd.n646 240.244
R14291 gnd.n6936 gnd.n646 240.244
R14292 gnd.n6936 gnd.n644 240.244
R14293 gnd.n6940 gnd.n644 240.244
R14294 gnd.n6940 gnd.n640 240.244
R14295 gnd.n6946 gnd.n640 240.244
R14296 gnd.n6946 gnd.n638 240.244
R14297 gnd.n6950 gnd.n638 240.244
R14298 gnd.n6950 gnd.n634 240.244
R14299 gnd.n6956 gnd.n634 240.244
R14300 gnd.n6956 gnd.n632 240.244
R14301 gnd.n6960 gnd.n632 240.244
R14302 gnd.n6960 gnd.n628 240.244
R14303 gnd.n6966 gnd.n628 240.244
R14304 gnd.n6966 gnd.n626 240.244
R14305 gnd.n6970 gnd.n626 240.244
R14306 gnd.n6970 gnd.n622 240.244
R14307 gnd.n6976 gnd.n622 240.244
R14308 gnd.n6976 gnd.n620 240.244
R14309 gnd.n6980 gnd.n620 240.244
R14310 gnd.n6980 gnd.n616 240.244
R14311 gnd.n6986 gnd.n616 240.244
R14312 gnd.n6986 gnd.n614 240.244
R14313 gnd.n6990 gnd.n614 240.244
R14314 gnd.n6990 gnd.n610 240.244
R14315 gnd.n6996 gnd.n610 240.244
R14316 gnd.n6996 gnd.n608 240.244
R14317 gnd.n7000 gnd.n608 240.244
R14318 gnd.n7000 gnd.n604 240.244
R14319 gnd.n7006 gnd.n604 240.244
R14320 gnd.n7006 gnd.n602 240.244
R14321 gnd.n7010 gnd.n602 240.244
R14322 gnd.n7010 gnd.n598 240.244
R14323 gnd.n7016 gnd.n598 240.244
R14324 gnd.n7016 gnd.n596 240.244
R14325 gnd.n7020 gnd.n596 240.244
R14326 gnd.n7020 gnd.n592 240.244
R14327 gnd.n7026 gnd.n592 240.244
R14328 gnd.n7026 gnd.n590 240.244
R14329 gnd.n7030 gnd.n590 240.244
R14330 gnd.n7030 gnd.n586 240.244
R14331 gnd.n7036 gnd.n586 240.244
R14332 gnd.n7036 gnd.n584 240.244
R14333 gnd.n7040 gnd.n584 240.244
R14334 gnd.n7040 gnd.n580 240.244
R14335 gnd.n7046 gnd.n580 240.244
R14336 gnd.n7046 gnd.n578 240.244
R14337 gnd.n7050 gnd.n578 240.244
R14338 gnd.n7050 gnd.n574 240.244
R14339 gnd.n7056 gnd.n574 240.244
R14340 gnd.n7056 gnd.n572 240.244
R14341 gnd.n7060 gnd.n572 240.244
R14342 gnd.n7060 gnd.n568 240.244
R14343 gnd.n7066 gnd.n568 240.244
R14344 gnd.n7066 gnd.n566 240.244
R14345 gnd.n7070 gnd.n566 240.244
R14346 gnd.n7070 gnd.n562 240.244
R14347 gnd.n7076 gnd.n562 240.244
R14348 gnd.n7076 gnd.n560 240.244
R14349 gnd.n7080 gnd.n560 240.244
R14350 gnd.n7080 gnd.n556 240.244
R14351 gnd.n7086 gnd.n556 240.244
R14352 gnd.n7086 gnd.n554 240.244
R14353 gnd.n7090 gnd.n554 240.244
R14354 gnd.n7090 gnd.n550 240.244
R14355 gnd.n7096 gnd.n550 240.244
R14356 gnd.n7096 gnd.n548 240.244
R14357 gnd.n7100 gnd.n548 240.244
R14358 gnd.n7100 gnd.n544 240.244
R14359 gnd.n7106 gnd.n544 240.244
R14360 gnd.n7106 gnd.n542 240.244
R14361 gnd.n7110 gnd.n542 240.244
R14362 gnd.n7110 gnd.n538 240.244
R14363 gnd.n7116 gnd.n538 240.244
R14364 gnd.n7116 gnd.n536 240.244
R14365 gnd.n7120 gnd.n536 240.244
R14366 gnd.n7120 gnd.n532 240.244
R14367 gnd.n7126 gnd.n532 240.244
R14368 gnd.n7126 gnd.n530 240.244
R14369 gnd.n7130 gnd.n530 240.244
R14370 gnd.n7136 gnd.n526 240.244
R14371 gnd.n7136 gnd.n524 240.244
R14372 gnd.n7140 gnd.n524 240.244
R14373 gnd.n7140 gnd.n520 240.244
R14374 gnd.n7146 gnd.n520 240.244
R14375 gnd.n7146 gnd.n518 240.244
R14376 gnd.n7150 gnd.n518 240.244
R14377 gnd.n7150 gnd.n514 240.244
R14378 gnd.n7156 gnd.n514 240.244
R14379 gnd.n7156 gnd.n512 240.244
R14380 gnd.n7160 gnd.n512 240.244
R14381 gnd.n7160 gnd.n508 240.244
R14382 gnd.n7166 gnd.n508 240.244
R14383 gnd.n7166 gnd.n506 240.244
R14384 gnd.n7170 gnd.n506 240.244
R14385 gnd.n7170 gnd.n502 240.244
R14386 gnd.n7176 gnd.n502 240.244
R14387 gnd.n7176 gnd.n500 240.244
R14388 gnd.n7180 gnd.n500 240.244
R14389 gnd.n7180 gnd.n496 240.244
R14390 gnd.n7186 gnd.n496 240.244
R14391 gnd.n7186 gnd.n494 240.244
R14392 gnd.n7190 gnd.n494 240.244
R14393 gnd.n7190 gnd.n490 240.244
R14394 gnd.n7196 gnd.n490 240.244
R14395 gnd.n7196 gnd.n488 240.244
R14396 gnd.n7200 gnd.n488 240.244
R14397 gnd.n7200 gnd.n484 240.244
R14398 gnd.n7206 gnd.n484 240.244
R14399 gnd.n7206 gnd.n482 240.244
R14400 gnd.n7210 gnd.n482 240.244
R14401 gnd.n7210 gnd.n478 240.244
R14402 gnd.n7216 gnd.n478 240.244
R14403 gnd.n7216 gnd.n476 240.244
R14404 gnd.n7220 gnd.n476 240.244
R14405 gnd.n7220 gnd.n472 240.244
R14406 gnd.n7226 gnd.n472 240.244
R14407 gnd.n7226 gnd.n470 240.244
R14408 gnd.n7230 gnd.n470 240.244
R14409 gnd.n7230 gnd.n466 240.244
R14410 gnd.n7236 gnd.n466 240.244
R14411 gnd.n7236 gnd.n464 240.244
R14412 gnd.n7240 gnd.n464 240.244
R14413 gnd.n7240 gnd.n460 240.244
R14414 gnd.n7246 gnd.n460 240.244
R14415 gnd.n7246 gnd.n458 240.244
R14416 gnd.n7250 gnd.n458 240.244
R14417 gnd.n7250 gnd.n454 240.244
R14418 gnd.n7256 gnd.n454 240.244
R14419 gnd.n7256 gnd.n452 240.244
R14420 gnd.n7260 gnd.n452 240.244
R14421 gnd.n7260 gnd.n448 240.244
R14422 gnd.n7266 gnd.n448 240.244
R14423 gnd.n7266 gnd.n446 240.244
R14424 gnd.n7270 gnd.n446 240.244
R14425 gnd.n7270 gnd.n442 240.244
R14426 gnd.n7276 gnd.n442 240.244
R14427 gnd.n7276 gnd.n440 240.244
R14428 gnd.n7280 gnd.n440 240.244
R14429 gnd.n7280 gnd.n436 240.244
R14430 gnd.n7286 gnd.n436 240.244
R14431 gnd.n7286 gnd.n434 240.244
R14432 gnd.n7290 gnd.n434 240.244
R14433 gnd.n7290 gnd.n430 240.244
R14434 gnd.n7296 gnd.n430 240.244
R14435 gnd.n7296 gnd.n428 240.244
R14436 gnd.n7300 gnd.n428 240.244
R14437 gnd.n7300 gnd.n424 240.244
R14438 gnd.n7306 gnd.n424 240.244
R14439 gnd.n7306 gnd.n422 240.244
R14440 gnd.n7310 gnd.n422 240.244
R14441 gnd.n7310 gnd.n418 240.244
R14442 gnd.n7316 gnd.n418 240.244
R14443 gnd.n7316 gnd.n416 240.244
R14444 gnd.n7320 gnd.n416 240.244
R14445 gnd.n7320 gnd.n412 240.244
R14446 gnd.n7326 gnd.n412 240.244
R14447 gnd.n7326 gnd.n410 240.244
R14448 gnd.n7330 gnd.n410 240.244
R14449 gnd.n7330 gnd.n406 240.244
R14450 gnd.n7338 gnd.n406 240.244
R14451 gnd.n7338 gnd.n404 240.244
R14452 gnd.n7342 gnd.n404 240.244
R14453 gnd.n7343 gnd.n7342 240.244
R14454 gnd.n2728 gnd.n2727 240.244
R14455 gnd.n2728 gnd.n2719 240.244
R14456 gnd.n2734 gnd.n2719 240.244
R14457 gnd.n2892 gnd.n2734 240.244
R14458 gnd.n2893 gnd.n2892 240.244
R14459 gnd.n2893 gnd.n2715 240.244
R14460 gnd.n2899 gnd.n2715 240.244
R14461 gnd.n2900 gnd.n2899 240.244
R14462 gnd.n2902 gnd.n2900 240.244
R14463 gnd.n2902 gnd.n2901 240.244
R14464 gnd.n2901 gnd.n2710 240.244
R14465 gnd.n2919 gnd.n2710 240.244
R14466 gnd.n2919 gnd.n2711 240.244
R14467 gnd.n2914 gnd.n2711 240.244
R14468 gnd.n2914 gnd.n2913 240.244
R14469 gnd.n2913 gnd.n2909 240.244
R14470 gnd.n2909 gnd.n2672 240.244
R14471 gnd.n2969 gnd.n2672 240.244
R14472 gnd.n2969 gnd.n2669 240.244
R14473 gnd.n2994 gnd.n2669 240.244
R14474 gnd.n2994 gnd.n2670 240.244
R14475 gnd.n2989 gnd.n2670 240.244
R14476 gnd.n2989 gnd.n2988 240.244
R14477 gnd.n2988 gnd.n2987 240.244
R14478 gnd.n2987 gnd.n2975 240.244
R14479 gnd.n2983 gnd.n2975 240.244
R14480 gnd.n2983 gnd.n2646 240.244
R14481 gnd.n3057 gnd.n2646 240.244
R14482 gnd.n3058 gnd.n3057 240.244
R14483 gnd.n3059 gnd.n3058 240.244
R14484 gnd.n3059 gnd.n2642 240.244
R14485 gnd.n3065 gnd.n2642 240.244
R14486 gnd.n3066 gnd.n3065 240.244
R14487 gnd.n3067 gnd.n3066 240.244
R14488 gnd.n3067 gnd.n2637 240.244
R14489 gnd.n3119 gnd.n2637 240.244
R14490 gnd.n3119 gnd.n2638 240.244
R14491 gnd.n3115 gnd.n2638 240.244
R14492 gnd.n3115 gnd.n3114 240.244
R14493 gnd.n3114 gnd.n3113 240.244
R14494 gnd.n3113 gnd.n3075 240.244
R14495 gnd.n3109 gnd.n3075 240.244
R14496 gnd.n3109 gnd.n3108 240.244
R14497 gnd.n3108 gnd.n3107 240.244
R14498 gnd.n3107 gnd.n3081 240.244
R14499 gnd.n3102 gnd.n3081 240.244
R14500 gnd.n3102 gnd.n3099 240.244
R14501 gnd.n3099 gnd.n3098 240.244
R14502 gnd.n3098 gnd.n3089 240.244
R14503 gnd.n3094 gnd.n3089 240.244
R14504 gnd.n3094 gnd.n2402 240.244
R14505 gnd.n3242 gnd.n2402 240.244
R14506 gnd.n3242 gnd.n2397 240.244
R14507 gnd.n3250 gnd.n2397 240.244
R14508 gnd.n3250 gnd.n2398 240.244
R14509 gnd.n2398 gnd.n2377 240.244
R14510 gnd.n3272 gnd.n2377 240.244
R14511 gnd.n3272 gnd.n2371 240.244
R14512 gnd.n3287 gnd.n2371 240.244
R14513 gnd.n3287 gnd.n2373 240.244
R14514 gnd.n3283 gnd.n2373 240.244
R14515 gnd.n3283 gnd.n3282 240.244
R14516 gnd.n3282 gnd.n1493 240.244
R14517 gnd.n4707 gnd.n1493 240.244
R14518 gnd.n4707 gnd.n1494 240.244
R14519 gnd.n4703 gnd.n1494 240.244
R14520 gnd.n4703 gnd.n1500 240.244
R14521 gnd.n4693 gnd.n1500 240.244
R14522 gnd.n4693 gnd.n1510 240.244
R14523 gnd.n4689 gnd.n1510 240.244
R14524 gnd.n4689 gnd.n1516 240.244
R14525 gnd.n4679 gnd.n1516 240.244
R14526 gnd.n4679 gnd.n1528 240.244
R14527 gnd.n4675 gnd.n1528 240.244
R14528 gnd.n4675 gnd.n1534 240.244
R14529 gnd.n3483 gnd.n1534 240.244
R14530 gnd.n3483 gnd.n3479 240.244
R14531 gnd.n3499 gnd.n3479 240.244
R14532 gnd.n3499 gnd.n3480 240.244
R14533 gnd.n3495 gnd.n3480 240.244
R14534 gnd.n3495 gnd.n3494 240.244
R14535 gnd.n3494 gnd.n2277 240.244
R14536 gnd.n3565 gnd.n2277 240.244
R14537 gnd.n3565 gnd.n2273 240.244
R14538 gnd.n3571 gnd.n2273 240.244
R14539 gnd.n3571 gnd.n2253 240.244
R14540 gnd.n3604 gnd.n2253 240.244
R14541 gnd.n3604 gnd.n2249 240.244
R14542 gnd.n3610 gnd.n2249 240.244
R14543 gnd.n3610 gnd.n2231 240.244
R14544 gnd.n3658 gnd.n2231 240.244
R14545 gnd.n3658 gnd.n2227 240.244
R14546 gnd.n3664 gnd.n2227 240.244
R14547 gnd.n3664 gnd.n2212 240.244
R14548 gnd.n3684 gnd.n2212 240.244
R14549 gnd.n3684 gnd.n2208 240.244
R14550 gnd.n3690 gnd.n2208 240.244
R14551 gnd.n3690 gnd.n2189 240.244
R14552 gnd.n3750 gnd.n2189 240.244
R14553 gnd.n3750 gnd.n2185 240.244
R14554 gnd.n3756 gnd.n2185 240.244
R14555 gnd.n3756 gnd.n2167 240.244
R14556 gnd.n3780 gnd.n2167 240.244
R14557 gnd.n3780 gnd.n2163 240.244
R14558 gnd.n3786 gnd.n2163 240.244
R14559 gnd.n3786 gnd.n2145 240.244
R14560 gnd.n3811 gnd.n2145 240.244
R14561 gnd.n3811 gnd.n2141 240.244
R14562 gnd.n3817 gnd.n2141 240.244
R14563 gnd.n3817 gnd.n2119 240.244
R14564 gnd.n3860 gnd.n2119 240.244
R14565 gnd.n3860 gnd.n2115 240.244
R14566 gnd.n3866 gnd.n2115 240.244
R14567 gnd.n3866 gnd.n2103 240.244
R14568 gnd.n3891 gnd.n2103 240.244
R14569 gnd.n3891 gnd.n2099 240.244
R14570 gnd.n3897 gnd.n2099 240.244
R14571 gnd.n3897 gnd.n2049 240.244
R14572 gnd.n4062 gnd.n2049 240.244
R14573 gnd.n4062 gnd.n2045 240.244
R14574 gnd.n4068 gnd.n2045 240.244
R14575 gnd.n4068 gnd.n2036 240.244
R14576 gnd.n4082 gnd.n2036 240.244
R14577 gnd.n4082 gnd.n2032 240.244
R14578 gnd.n4088 gnd.n2032 240.244
R14579 gnd.n4088 gnd.n2023 240.244
R14580 gnd.n4102 gnd.n2023 240.244
R14581 gnd.n4102 gnd.n2018 240.244
R14582 gnd.n4110 gnd.n2018 240.244
R14583 gnd.n4110 gnd.n2019 240.244
R14584 gnd.n2019 gnd.n2008 240.244
R14585 gnd.n4126 gnd.n2008 240.244
R14586 gnd.n4126 gnd.n2003 240.244
R14587 gnd.n4176 gnd.n2003 240.244
R14588 gnd.n4176 gnd.n2004 240.244
R14589 gnd.n4172 gnd.n2004 240.244
R14590 gnd.n4172 gnd.n4171 240.244
R14591 gnd.n4171 gnd.n4170 240.244
R14592 gnd.n4170 gnd.n4134 240.244
R14593 gnd.n4166 gnd.n4134 240.244
R14594 gnd.n4166 gnd.n4165 240.244
R14595 gnd.n4165 gnd.n4164 240.244
R14596 gnd.n4164 gnd.n4140 240.244
R14597 gnd.n4160 gnd.n4140 240.244
R14598 gnd.n4160 gnd.n4159 240.244
R14599 gnd.n4159 gnd.n4158 240.244
R14600 gnd.n4158 gnd.n4146 240.244
R14601 gnd.n4154 gnd.n4146 240.244
R14602 gnd.n4154 gnd.n1951 240.244
R14603 gnd.n4250 gnd.n1951 240.244
R14604 gnd.n4251 gnd.n4250 240.244
R14605 gnd.n4252 gnd.n4251 240.244
R14606 gnd.n4252 gnd.n1947 240.244
R14607 gnd.n4258 gnd.n1947 240.244
R14608 gnd.n4259 gnd.n4258 240.244
R14609 gnd.n4260 gnd.n4259 240.244
R14610 gnd.n4260 gnd.n1942 240.244
R14611 gnd.n4271 gnd.n1942 240.244
R14612 gnd.n4271 gnd.n1943 240.244
R14613 gnd.n4267 gnd.n1943 240.244
R14614 gnd.n4267 gnd.n1913 240.244
R14615 gnd.n4325 gnd.n1913 240.244
R14616 gnd.n4325 gnd.n1914 240.244
R14617 gnd.n4320 gnd.n1914 240.244
R14618 gnd.n4320 gnd.n1921 240.244
R14619 gnd.n1921 gnd.n1917 240.244
R14620 gnd.n1917 gnd.n382 240.244
R14621 gnd.n7368 gnd.n382 240.244
R14622 gnd.n7368 gnd.n383 240.244
R14623 gnd.n7363 gnd.n383 240.244
R14624 gnd.n7363 gnd.n7362 240.244
R14625 gnd.n7362 gnd.n7361 240.244
R14626 gnd.n7361 gnd.n387 240.244
R14627 gnd.n7357 gnd.n387 240.244
R14628 gnd.n7357 gnd.n7356 240.244
R14629 gnd.n7356 gnd.n7355 240.244
R14630 gnd.n7355 gnd.n393 240.244
R14631 gnd.n7351 gnd.n393 240.244
R14632 gnd.n7351 gnd.n7350 240.244
R14633 gnd.n7350 gnd.n7349 240.244
R14634 gnd.n7349 gnd.n399 240.244
R14635 gnd.n6676 gnd.n802 240.244
R14636 gnd.n6672 gnd.n802 240.244
R14637 gnd.n6672 gnd.n807 240.244
R14638 gnd.n6668 gnd.n807 240.244
R14639 gnd.n6668 gnd.n809 240.244
R14640 gnd.n6664 gnd.n809 240.244
R14641 gnd.n6664 gnd.n815 240.244
R14642 gnd.n6660 gnd.n815 240.244
R14643 gnd.n6660 gnd.n817 240.244
R14644 gnd.n6656 gnd.n817 240.244
R14645 gnd.n6656 gnd.n823 240.244
R14646 gnd.n6652 gnd.n823 240.244
R14647 gnd.n6652 gnd.n825 240.244
R14648 gnd.n6648 gnd.n825 240.244
R14649 gnd.n6648 gnd.n831 240.244
R14650 gnd.n6644 gnd.n831 240.244
R14651 gnd.n6644 gnd.n833 240.244
R14652 gnd.n6640 gnd.n833 240.244
R14653 gnd.n6640 gnd.n839 240.244
R14654 gnd.n6636 gnd.n839 240.244
R14655 gnd.n6636 gnd.n841 240.244
R14656 gnd.n6632 gnd.n841 240.244
R14657 gnd.n6632 gnd.n847 240.244
R14658 gnd.n6628 gnd.n847 240.244
R14659 gnd.n6628 gnd.n849 240.244
R14660 gnd.n6624 gnd.n849 240.244
R14661 gnd.n6624 gnd.n855 240.244
R14662 gnd.n6620 gnd.n855 240.244
R14663 gnd.n6620 gnd.n857 240.244
R14664 gnd.n6616 gnd.n857 240.244
R14665 gnd.n6616 gnd.n863 240.244
R14666 gnd.n6612 gnd.n863 240.244
R14667 gnd.n6612 gnd.n865 240.244
R14668 gnd.n6608 gnd.n865 240.244
R14669 gnd.n6608 gnd.n871 240.244
R14670 gnd.n6604 gnd.n871 240.244
R14671 gnd.n6604 gnd.n873 240.244
R14672 gnd.n6600 gnd.n873 240.244
R14673 gnd.n6600 gnd.n879 240.244
R14674 gnd.n6596 gnd.n879 240.244
R14675 gnd.n6596 gnd.n881 240.244
R14676 gnd.n6592 gnd.n881 240.244
R14677 gnd.n6592 gnd.n887 240.244
R14678 gnd.n6588 gnd.n887 240.244
R14679 gnd.n6588 gnd.n889 240.244
R14680 gnd.n6584 gnd.n889 240.244
R14681 gnd.n6584 gnd.n895 240.244
R14682 gnd.n6580 gnd.n895 240.244
R14683 gnd.n6580 gnd.n897 240.244
R14684 gnd.n6576 gnd.n897 240.244
R14685 gnd.n6576 gnd.n903 240.244
R14686 gnd.n6572 gnd.n903 240.244
R14687 gnd.n6572 gnd.n905 240.244
R14688 gnd.n6568 gnd.n905 240.244
R14689 gnd.n6568 gnd.n911 240.244
R14690 gnd.n6564 gnd.n911 240.244
R14691 gnd.n6564 gnd.n913 240.244
R14692 gnd.n6560 gnd.n913 240.244
R14693 gnd.n6560 gnd.n919 240.244
R14694 gnd.n6556 gnd.n919 240.244
R14695 gnd.n6556 gnd.n921 240.244
R14696 gnd.n6552 gnd.n921 240.244
R14697 gnd.n6552 gnd.n927 240.244
R14698 gnd.n6548 gnd.n927 240.244
R14699 gnd.n6548 gnd.n929 240.244
R14700 gnd.n6544 gnd.n929 240.244
R14701 gnd.n6544 gnd.n935 240.244
R14702 gnd.n6540 gnd.n935 240.244
R14703 gnd.n6540 gnd.n937 240.244
R14704 gnd.n6536 gnd.n937 240.244
R14705 gnd.n6536 gnd.n943 240.244
R14706 gnd.n6532 gnd.n943 240.244
R14707 gnd.n6532 gnd.n945 240.244
R14708 gnd.n6528 gnd.n945 240.244
R14709 gnd.n6528 gnd.n951 240.244
R14710 gnd.n6524 gnd.n951 240.244
R14711 gnd.n6524 gnd.n953 240.244
R14712 gnd.n6520 gnd.n953 240.244
R14713 gnd.n6520 gnd.n959 240.244
R14714 gnd.n6516 gnd.n959 240.244
R14715 gnd.n6516 gnd.n961 240.244
R14716 gnd.n6512 gnd.n961 240.244
R14717 gnd.n6512 gnd.n967 240.244
R14718 gnd.n2726 gnd.n967 240.244
R14719 gnd.n3230 gnd.n2412 240.244
R14720 gnd.n3230 gnd.n2413 240.244
R14721 gnd.n2413 gnd.n2393 240.244
R14722 gnd.n3253 gnd.n2393 240.244
R14723 gnd.n3253 gnd.n2387 240.244
R14724 gnd.n3260 gnd.n2387 240.244
R14725 gnd.n3260 gnd.n2388 240.244
R14726 gnd.n2388 gnd.n2367 240.244
R14727 gnd.n3290 gnd.n2367 240.244
R14728 gnd.n3290 gnd.n2362 240.244
R14729 gnd.n3297 gnd.n2362 240.244
R14730 gnd.n3297 gnd.n2353 240.244
R14731 gnd.n3417 gnd.n2353 240.244
R14732 gnd.n3418 gnd.n3417 240.244
R14733 gnd.n3418 gnd.n2349 240.244
R14734 gnd.n3424 gnd.n2349 240.244
R14735 gnd.n3424 gnd.n2339 240.244
R14736 gnd.n3436 gnd.n2339 240.244
R14737 gnd.n3436 gnd.n2333 240.244
R14738 gnd.n3450 gnd.n2333 240.244
R14739 gnd.n3450 gnd.n2334 240.244
R14740 gnd.n3441 gnd.n2334 240.244
R14741 gnd.n3443 gnd.n3441 240.244
R14742 gnd.n3443 gnd.n1538 240.244
R14743 gnd.n4672 gnd.n1538 240.244
R14744 gnd.n4672 gnd.n1539 240.244
R14745 gnd.n1544 gnd.n1539 240.244
R14746 gnd.n1545 gnd.n1544 240.244
R14747 gnd.n1546 gnd.n1545 240.244
R14748 gnd.n3527 gnd.n1546 240.244
R14749 gnd.n3527 gnd.n1549 240.244
R14750 gnd.n1550 gnd.n1549 240.244
R14751 gnd.n1551 gnd.n1550 240.244
R14752 gnd.n2280 gnd.n1551 240.244
R14753 gnd.n2280 gnd.n1554 240.244
R14754 gnd.n1555 gnd.n1554 240.244
R14755 gnd.n1556 gnd.n1555 240.244
R14756 gnd.n2256 gnd.n1556 240.244
R14757 gnd.n2256 gnd.n1559 240.244
R14758 gnd.n1560 gnd.n1559 240.244
R14759 gnd.n1561 gnd.n1560 240.244
R14760 gnd.n3655 gnd.n1561 240.244
R14761 gnd.n3655 gnd.n1564 240.244
R14762 gnd.n1565 gnd.n1564 240.244
R14763 gnd.n1566 gnd.n1565 240.244
R14764 gnd.n3681 gnd.n1566 240.244
R14765 gnd.n3681 gnd.n1569 240.244
R14766 gnd.n1570 gnd.n1569 240.244
R14767 gnd.n1571 gnd.n1570 240.244
R14768 gnd.n2192 gnd.n1571 240.244
R14769 gnd.n2192 gnd.n1574 240.244
R14770 gnd.n1575 gnd.n1574 240.244
R14771 gnd.n1576 gnd.n1575 240.244
R14772 gnd.n2169 gnd.n1576 240.244
R14773 gnd.n2169 gnd.n1579 240.244
R14774 gnd.n1580 gnd.n1579 240.244
R14775 gnd.n1581 gnd.n1580 240.244
R14776 gnd.n2147 gnd.n1581 240.244
R14777 gnd.n2147 gnd.n1584 240.244
R14778 gnd.n1585 gnd.n1584 240.244
R14779 gnd.n1586 gnd.n1585 240.244
R14780 gnd.n3713 gnd.n1586 240.244
R14781 gnd.n3713 gnd.n1589 240.244
R14782 gnd.n1590 gnd.n1589 240.244
R14783 gnd.n1591 gnd.n1590 240.244
R14784 gnd.n2105 gnd.n1591 240.244
R14785 gnd.n2105 gnd.n1594 240.244
R14786 gnd.n1595 gnd.n1594 240.244
R14787 gnd.n1596 gnd.n1595 240.244
R14788 gnd.n2068 gnd.n1596 240.244
R14789 gnd.n2068 gnd.n1599 240.244
R14790 gnd.n1600 gnd.n1599 240.244
R14791 gnd.n1601 gnd.n1600 240.244
R14792 gnd.n4079 gnd.n1601 240.244
R14793 gnd.n4079 gnd.n1604 240.244
R14794 gnd.n1605 gnd.n1604 240.244
R14795 gnd.n1606 gnd.n1605 240.244
R14796 gnd.n4099 gnd.n1606 240.244
R14797 gnd.n4099 gnd.n1609 240.244
R14798 gnd.n1610 gnd.n1609 240.244
R14799 gnd.n1611 gnd.n1610 240.244
R14800 gnd.n4123 gnd.n1611 240.244
R14801 gnd.n3220 gnd.n2418 240.244
R14802 gnd.n3220 gnd.n2434 240.244
R14803 gnd.n2438 gnd.n2437 240.244
R14804 gnd.n2440 gnd.n2439 240.244
R14805 gnd.n2557 gnd.n2556 240.244
R14806 gnd.n2567 gnd.n2566 240.244
R14807 gnd.n2569 gnd.n2568 240.244
R14808 gnd.n2579 gnd.n2578 240.244
R14809 gnd.n2590 gnd.n2589 240.244
R14810 gnd.n2592 gnd.n2591 240.244
R14811 gnd.n2602 gnd.n2601 240.244
R14812 gnd.n2613 gnd.n2612 240.244
R14813 gnd.n3149 gnd.n2614 240.244
R14814 gnd.n3153 gnd.n3152 240.244
R14815 gnd.n3232 gnd.n2409 240.244
R14816 gnd.n3232 gnd.n2404 240.244
R14817 gnd.n3239 gnd.n2404 240.244
R14818 gnd.n3239 gnd.n2395 240.244
R14819 gnd.n2395 gnd.n2384 240.244
R14820 gnd.n3262 gnd.n2384 240.244
R14821 gnd.n3262 gnd.n2379 240.244
R14822 gnd.n3269 gnd.n2379 240.244
R14823 gnd.n3269 gnd.n2369 240.244
R14824 gnd.n2369 gnd.n2360 240.244
R14825 gnd.n3299 gnd.n2360 240.244
R14826 gnd.n3299 gnd.n2354 240.244
R14827 gnd.n3306 gnd.n2354 240.244
R14828 gnd.n3306 gnd.n2355 240.244
R14829 gnd.n2355 gnd.n2347 240.244
R14830 gnd.n3426 gnd.n2347 240.244
R14831 gnd.n3426 gnd.n2342 240.244
R14832 gnd.n3434 gnd.n2342 240.244
R14833 gnd.n3434 gnd.n2331 240.244
R14834 gnd.n3452 gnd.n2331 240.244
R14835 gnd.n3453 gnd.n3452 240.244
R14836 gnd.n3454 gnd.n3453 240.244
R14837 gnd.n3454 gnd.n2326 240.244
R14838 gnd.n3461 gnd.n2326 240.244
R14839 gnd.n3461 gnd.n1536 240.244
R14840 gnd.n2312 gnd.n1536 240.244
R14841 gnd.n3509 gnd.n2312 240.244
R14842 gnd.n3509 gnd.n2307 240.244
R14843 gnd.n3517 gnd.n2307 240.244
R14844 gnd.n3517 gnd.n2296 240.244
R14845 gnd.n3537 gnd.n2296 240.244
R14846 gnd.n3538 gnd.n3537 240.244
R14847 gnd.n3539 gnd.n3538 240.244
R14848 gnd.n3539 gnd.n2292 240.244
R14849 gnd.n3545 gnd.n2292 240.244
R14850 gnd.n3545 gnd.n2264 240.244
R14851 gnd.n3591 gnd.n2264 240.244
R14852 gnd.n3591 gnd.n2265 240.244
R14853 gnd.n3585 gnd.n2265 240.244
R14854 gnd.n3585 gnd.n2241 240.244
R14855 gnd.n3646 gnd.n2241 240.244
R14856 gnd.n3646 gnd.n2233 240.244
R14857 gnd.n3625 gnd.n2233 240.244
R14858 gnd.n3626 gnd.n3625 240.244
R14859 gnd.n3627 gnd.n3626 240.244
R14860 gnd.n3627 gnd.n2214 240.244
R14861 gnd.n2214 gnd.n2207 240.244
R14862 gnd.n3630 gnd.n2207 240.244
R14863 gnd.n3631 gnd.n3630 240.244
R14864 gnd.n3631 gnd.n2182 240.244
R14865 gnd.n3759 gnd.n2182 240.244
R14866 gnd.n3759 gnd.n2178 240.244
R14867 gnd.n3765 gnd.n2178 240.244
R14868 gnd.n3765 gnd.n2161 240.244
R14869 gnd.n3789 gnd.n2161 240.244
R14870 gnd.n3789 gnd.n2155 240.244
R14871 gnd.n3799 gnd.n2155 240.244
R14872 gnd.n3799 gnd.n2156 240.244
R14873 gnd.n3793 gnd.n2156 240.244
R14874 gnd.n3793 gnd.n2132 240.244
R14875 gnd.n3828 gnd.n2132 240.244
R14876 gnd.n3828 gnd.n2126 240.244
R14877 gnd.n3850 gnd.n2126 240.244
R14878 gnd.n3850 gnd.n2127 240.244
R14879 gnd.n2127 gnd.n2112 240.244
R14880 gnd.n3833 gnd.n2112 240.244
R14881 gnd.n3834 gnd.n3833 240.244
R14882 gnd.n3837 gnd.n3834 240.244
R14883 gnd.n3838 gnd.n3837 240.244
R14884 gnd.n3838 gnd.n2042 240.244
R14885 gnd.n4071 gnd.n2042 240.244
R14886 gnd.n4071 gnd.n2038 240.244
R14887 gnd.n4077 gnd.n2038 240.244
R14888 gnd.n4077 gnd.n2029 240.244
R14889 gnd.n4091 gnd.n2029 240.244
R14890 gnd.n4091 gnd.n2025 240.244
R14891 gnd.n4097 gnd.n2025 240.244
R14892 gnd.n4097 gnd.n2015 240.244
R14893 gnd.n4113 gnd.n2015 240.244
R14894 gnd.n4113 gnd.n2010 240.244
R14895 gnd.n4120 gnd.n2010 240.244
R14896 gnd.n4120 gnd.n1977 240.244
R14897 gnd.n1616 gnd.n1615 240.244
R14898 gnd.n1980 gnd.n1619 240.244
R14899 gnd.n1621 gnd.n1620 240.244
R14900 gnd.n1983 gnd.n1625 240.244
R14901 gnd.n1986 gnd.n1626 240.244
R14902 gnd.n1635 gnd.n1634 240.244
R14903 gnd.n1988 gnd.n1642 240.244
R14904 gnd.n1991 gnd.n1643 240.244
R14905 gnd.n1651 gnd.n1650 240.244
R14906 gnd.n1993 gnd.n1658 240.244
R14907 gnd.n1996 gnd.n1659 240.244
R14908 gnd.n1667 gnd.n1666 240.244
R14909 gnd.n1999 gnd.n1667 240.244
R14910 gnd.n2000 gnd.n1976 240.244
R14911 gnd.n1475 gnd.n1474 240.132
R14912 gnd.n3914 gnd.n3913 240.132
R14913 gnd.n6679 gnd.n6678 225.874
R14914 gnd.n6679 gnd.n795 225.874
R14915 gnd.n6687 gnd.n795 225.874
R14916 gnd.n6688 gnd.n6687 225.874
R14917 gnd.n6689 gnd.n6688 225.874
R14918 gnd.n6689 gnd.n789 225.874
R14919 gnd.n6697 gnd.n789 225.874
R14920 gnd.n6698 gnd.n6697 225.874
R14921 gnd.n6699 gnd.n6698 225.874
R14922 gnd.n6699 gnd.n783 225.874
R14923 gnd.n6707 gnd.n783 225.874
R14924 gnd.n6708 gnd.n6707 225.874
R14925 gnd.n6709 gnd.n6708 225.874
R14926 gnd.n6709 gnd.n777 225.874
R14927 gnd.n6717 gnd.n777 225.874
R14928 gnd.n6718 gnd.n6717 225.874
R14929 gnd.n6719 gnd.n6718 225.874
R14930 gnd.n6719 gnd.n771 225.874
R14931 gnd.n6727 gnd.n771 225.874
R14932 gnd.n6728 gnd.n6727 225.874
R14933 gnd.n6729 gnd.n6728 225.874
R14934 gnd.n6729 gnd.n765 225.874
R14935 gnd.n6737 gnd.n765 225.874
R14936 gnd.n6738 gnd.n6737 225.874
R14937 gnd.n6739 gnd.n6738 225.874
R14938 gnd.n6739 gnd.n759 225.874
R14939 gnd.n6747 gnd.n759 225.874
R14940 gnd.n6748 gnd.n6747 225.874
R14941 gnd.n6749 gnd.n6748 225.874
R14942 gnd.n6749 gnd.n753 225.874
R14943 gnd.n6757 gnd.n753 225.874
R14944 gnd.n6758 gnd.n6757 225.874
R14945 gnd.n6759 gnd.n6758 225.874
R14946 gnd.n6759 gnd.n747 225.874
R14947 gnd.n6767 gnd.n747 225.874
R14948 gnd.n6768 gnd.n6767 225.874
R14949 gnd.n6769 gnd.n6768 225.874
R14950 gnd.n6769 gnd.n741 225.874
R14951 gnd.n6777 gnd.n741 225.874
R14952 gnd.n6778 gnd.n6777 225.874
R14953 gnd.n6779 gnd.n6778 225.874
R14954 gnd.n6779 gnd.n735 225.874
R14955 gnd.n6787 gnd.n735 225.874
R14956 gnd.n6788 gnd.n6787 225.874
R14957 gnd.n6789 gnd.n6788 225.874
R14958 gnd.n6789 gnd.n729 225.874
R14959 gnd.n6797 gnd.n729 225.874
R14960 gnd.n6798 gnd.n6797 225.874
R14961 gnd.n6799 gnd.n6798 225.874
R14962 gnd.n6799 gnd.n723 225.874
R14963 gnd.n6807 gnd.n723 225.874
R14964 gnd.n6808 gnd.n6807 225.874
R14965 gnd.n6809 gnd.n6808 225.874
R14966 gnd.n6809 gnd.n717 225.874
R14967 gnd.n6817 gnd.n717 225.874
R14968 gnd.n6818 gnd.n6817 225.874
R14969 gnd.n6819 gnd.n6818 225.874
R14970 gnd.n6819 gnd.n711 225.874
R14971 gnd.n6827 gnd.n711 225.874
R14972 gnd.n6828 gnd.n6827 225.874
R14973 gnd.n6829 gnd.n6828 225.874
R14974 gnd.n6829 gnd.n705 225.874
R14975 gnd.n6837 gnd.n705 225.874
R14976 gnd.n6838 gnd.n6837 225.874
R14977 gnd.n6839 gnd.n6838 225.874
R14978 gnd.n6839 gnd.n699 225.874
R14979 gnd.n6847 gnd.n699 225.874
R14980 gnd.n6848 gnd.n6847 225.874
R14981 gnd.n6849 gnd.n6848 225.874
R14982 gnd.n6849 gnd.n693 225.874
R14983 gnd.n6857 gnd.n693 225.874
R14984 gnd.n6858 gnd.n6857 225.874
R14985 gnd.n6859 gnd.n6858 225.874
R14986 gnd.n6859 gnd.n687 225.874
R14987 gnd.n6867 gnd.n687 225.874
R14988 gnd.n6868 gnd.n6867 225.874
R14989 gnd.n6869 gnd.n6868 225.874
R14990 gnd.n6869 gnd.n681 225.874
R14991 gnd.n6877 gnd.n681 225.874
R14992 gnd.n6878 gnd.n6877 225.874
R14993 gnd.n6879 gnd.n6878 225.874
R14994 gnd.n6879 gnd.n675 225.874
R14995 gnd.n6887 gnd.n675 225.874
R14996 gnd.n6888 gnd.n6887 225.874
R14997 gnd.n6889 gnd.n6888 225.874
R14998 gnd.n6889 gnd.n669 225.874
R14999 gnd.n6897 gnd.n669 225.874
R15000 gnd.n6898 gnd.n6897 225.874
R15001 gnd.n6899 gnd.n6898 225.874
R15002 gnd.n6899 gnd.n663 225.874
R15003 gnd.n6907 gnd.n663 225.874
R15004 gnd.n6908 gnd.n6907 225.874
R15005 gnd.n6909 gnd.n6908 225.874
R15006 gnd.n6909 gnd.n657 225.874
R15007 gnd.n6917 gnd.n657 225.874
R15008 gnd.n6918 gnd.n6917 225.874
R15009 gnd.n6919 gnd.n6918 225.874
R15010 gnd.n6919 gnd.n651 225.874
R15011 gnd.n6927 gnd.n651 225.874
R15012 gnd.n6928 gnd.n6927 225.874
R15013 gnd.n6929 gnd.n6928 225.874
R15014 gnd.n6929 gnd.n645 225.874
R15015 gnd.n6937 gnd.n645 225.874
R15016 gnd.n6938 gnd.n6937 225.874
R15017 gnd.n6939 gnd.n6938 225.874
R15018 gnd.n6939 gnd.n639 225.874
R15019 gnd.n6947 gnd.n639 225.874
R15020 gnd.n6948 gnd.n6947 225.874
R15021 gnd.n6949 gnd.n6948 225.874
R15022 gnd.n6949 gnd.n633 225.874
R15023 gnd.n6957 gnd.n633 225.874
R15024 gnd.n6958 gnd.n6957 225.874
R15025 gnd.n6959 gnd.n6958 225.874
R15026 gnd.n6959 gnd.n627 225.874
R15027 gnd.n6967 gnd.n627 225.874
R15028 gnd.n6968 gnd.n6967 225.874
R15029 gnd.n6969 gnd.n6968 225.874
R15030 gnd.n6969 gnd.n621 225.874
R15031 gnd.n6977 gnd.n621 225.874
R15032 gnd.n6978 gnd.n6977 225.874
R15033 gnd.n6979 gnd.n6978 225.874
R15034 gnd.n6979 gnd.n615 225.874
R15035 gnd.n6987 gnd.n615 225.874
R15036 gnd.n6988 gnd.n6987 225.874
R15037 gnd.n6989 gnd.n6988 225.874
R15038 gnd.n6989 gnd.n609 225.874
R15039 gnd.n6997 gnd.n609 225.874
R15040 gnd.n6998 gnd.n6997 225.874
R15041 gnd.n6999 gnd.n6998 225.874
R15042 gnd.n6999 gnd.n603 225.874
R15043 gnd.n7007 gnd.n603 225.874
R15044 gnd.n7008 gnd.n7007 225.874
R15045 gnd.n7009 gnd.n7008 225.874
R15046 gnd.n7009 gnd.n597 225.874
R15047 gnd.n7017 gnd.n597 225.874
R15048 gnd.n7018 gnd.n7017 225.874
R15049 gnd.n7019 gnd.n7018 225.874
R15050 gnd.n7019 gnd.n591 225.874
R15051 gnd.n7027 gnd.n591 225.874
R15052 gnd.n7028 gnd.n7027 225.874
R15053 gnd.n7029 gnd.n7028 225.874
R15054 gnd.n7029 gnd.n585 225.874
R15055 gnd.n7037 gnd.n585 225.874
R15056 gnd.n7038 gnd.n7037 225.874
R15057 gnd.n7039 gnd.n7038 225.874
R15058 gnd.n7039 gnd.n579 225.874
R15059 gnd.n7047 gnd.n579 225.874
R15060 gnd.n7048 gnd.n7047 225.874
R15061 gnd.n7049 gnd.n7048 225.874
R15062 gnd.n7049 gnd.n573 225.874
R15063 gnd.n7057 gnd.n573 225.874
R15064 gnd.n7058 gnd.n7057 225.874
R15065 gnd.n7059 gnd.n7058 225.874
R15066 gnd.n7059 gnd.n567 225.874
R15067 gnd.n7067 gnd.n567 225.874
R15068 gnd.n7068 gnd.n7067 225.874
R15069 gnd.n7069 gnd.n7068 225.874
R15070 gnd.n7069 gnd.n561 225.874
R15071 gnd.n7077 gnd.n561 225.874
R15072 gnd.n7078 gnd.n7077 225.874
R15073 gnd.n7079 gnd.n7078 225.874
R15074 gnd.n7079 gnd.n555 225.874
R15075 gnd.n7087 gnd.n555 225.874
R15076 gnd.n7088 gnd.n7087 225.874
R15077 gnd.n7089 gnd.n7088 225.874
R15078 gnd.n7089 gnd.n549 225.874
R15079 gnd.n7097 gnd.n549 225.874
R15080 gnd.n7098 gnd.n7097 225.874
R15081 gnd.n7099 gnd.n7098 225.874
R15082 gnd.n7099 gnd.n543 225.874
R15083 gnd.n7107 gnd.n543 225.874
R15084 gnd.n7108 gnd.n7107 225.874
R15085 gnd.n7109 gnd.n7108 225.874
R15086 gnd.n7109 gnd.n537 225.874
R15087 gnd.n7117 gnd.n537 225.874
R15088 gnd.n7118 gnd.n7117 225.874
R15089 gnd.n7119 gnd.n7118 225.874
R15090 gnd.n7119 gnd.n531 225.874
R15091 gnd.n7127 gnd.n531 225.874
R15092 gnd.n7128 gnd.n7127 225.874
R15093 gnd.n7129 gnd.n7128 225.874
R15094 gnd.n5539 gnd.t257 224.174
R15095 gnd.n5167 gnd.t252 224.174
R15096 gnd.n1751 gnd.n1688 199.319
R15097 gnd.n1751 gnd.n1689 199.319
R15098 gnd.n1427 gnd.n1426 199.319
R15099 gnd.n2477 gnd.n1427 199.319
R15100 gnd.n1476 gnd.n1473 186.49
R15101 gnd.n3915 gnd.n3912 186.49
R15102 gnd.n6335 gnd.n6334 185
R15103 gnd.n6333 gnd.n6332 185
R15104 gnd.n6312 gnd.n6311 185
R15105 gnd.n6327 gnd.n6326 185
R15106 gnd.n6325 gnd.n6324 185
R15107 gnd.n6316 gnd.n6315 185
R15108 gnd.n6319 gnd.n6318 185
R15109 gnd.n6303 gnd.n6302 185
R15110 gnd.n6301 gnd.n6300 185
R15111 gnd.n6280 gnd.n6279 185
R15112 gnd.n6295 gnd.n6294 185
R15113 gnd.n6293 gnd.n6292 185
R15114 gnd.n6284 gnd.n6283 185
R15115 gnd.n6287 gnd.n6286 185
R15116 gnd.n6271 gnd.n6270 185
R15117 gnd.n6269 gnd.n6268 185
R15118 gnd.n6248 gnd.n6247 185
R15119 gnd.n6263 gnd.n6262 185
R15120 gnd.n6261 gnd.n6260 185
R15121 gnd.n6252 gnd.n6251 185
R15122 gnd.n6255 gnd.n6254 185
R15123 gnd.n6240 gnd.n6239 185
R15124 gnd.n6238 gnd.n6237 185
R15125 gnd.n6217 gnd.n6216 185
R15126 gnd.n6232 gnd.n6231 185
R15127 gnd.n6230 gnd.n6229 185
R15128 gnd.n6221 gnd.n6220 185
R15129 gnd.n6224 gnd.n6223 185
R15130 gnd.n6208 gnd.n6207 185
R15131 gnd.n6206 gnd.n6205 185
R15132 gnd.n6185 gnd.n6184 185
R15133 gnd.n6200 gnd.n6199 185
R15134 gnd.n6198 gnd.n6197 185
R15135 gnd.n6189 gnd.n6188 185
R15136 gnd.n6192 gnd.n6191 185
R15137 gnd.n6176 gnd.n6175 185
R15138 gnd.n6174 gnd.n6173 185
R15139 gnd.n6153 gnd.n6152 185
R15140 gnd.n6168 gnd.n6167 185
R15141 gnd.n6166 gnd.n6165 185
R15142 gnd.n6157 gnd.n6156 185
R15143 gnd.n6160 gnd.n6159 185
R15144 gnd.n6144 gnd.n6143 185
R15145 gnd.n6142 gnd.n6141 185
R15146 gnd.n6121 gnd.n6120 185
R15147 gnd.n6136 gnd.n6135 185
R15148 gnd.n6134 gnd.n6133 185
R15149 gnd.n6125 gnd.n6124 185
R15150 gnd.n6128 gnd.n6127 185
R15151 gnd.n6113 gnd.n6112 185
R15152 gnd.n6111 gnd.n6110 185
R15153 gnd.n6090 gnd.n6089 185
R15154 gnd.n6105 gnd.n6104 185
R15155 gnd.n6103 gnd.n6102 185
R15156 gnd.n6094 gnd.n6093 185
R15157 gnd.n6097 gnd.n6096 185
R15158 gnd.n5540 gnd.t256 178.987
R15159 gnd.n5168 gnd.t253 178.987
R15160 gnd.n7137 gnd.n525 173.845
R15161 gnd.n7138 gnd.n7137 173.845
R15162 gnd.n7139 gnd.n7138 173.845
R15163 gnd.n7139 gnd.n519 173.845
R15164 gnd.n7147 gnd.n519 173.845
R15165 gnd.n7148 gnd.n7147 173.845
R15166 gnd.n7149 gnd.n7148 173.845
R15167 gnd.n7149 gnd.n513 173.845
R15168 gnd.n7157 gnd.n513 173.845
R15169 gnd.n7158 gnd.n7157 173.845
R15170 gnd.n7159 gnd.n7158 173.845
R15171 gnd.n7159 gnd.n507 173.845
R15172 gnd.n7167 gnd.n507 173.845
R15173 gnd.n7168 gnd.n7167 173.845
R15174 gnd.n7169 gnd.n7168 173.845
R15175 gnd.n7169 gnd.n501 173.845
R15176 gnd.n7177 gnd.n501 173.845
R15177 gnd.n7178 gnd.n7177 173.845
R15178 gnd.n7179 gnd.n7178 173.845
R15179 gnd.n7179 gnd.n495 173.845
R15180 gnd.n7187 gnd.n495 173.845
R15181 gnd.n7188 gnd.n7187 173.845
R15182 gnd.n7189 gnd.n7188 173.845
R15183 gnd.n7189 gnd.n489 173.845
R15184 gnd.n7197 gnd.n489 173.845
R15185 gnd.n7198 gnd.n7197 173.845
R15186 gnd.n7199 gnd.n7198 173.845
R15187 gnd.n7199 gnd.n483 173.845
R15188 gnd.n7207 gnd.n483 173.845
R15189 gnd.n7208 gnd.n7207 173.845
R15190 gnd.n7209 gnd.n7208 173.845
R15191 gnd.n7209 gnd.n477 173.845
R15192 gnd.n7217 gnd.n477 173.845
R15193 gnd.n7218 gnd.n7217 173.845
R15194 gnd.n7219 gnd.n7218 173.845
R15195 gnd.n7219 gnd.n471 173.845
R15196 gnd.n7227 gnd.n471 173.845
R15197 gnd.n7228 gnd.n7227 173.845
R15198 gnd.n7229 gnd.n7228 173.845
R15199 gnd.n7229 gnd.n465 173.845
R15200 gnd.n7237 gnd.n465 173.845
R15201 gnd.n7238 gnd.n7237 173.845
R15202 gnd.n7239 gnd.n7238 173.845
R15203 gnd.n7239 gnd.n459 173.845
R15204 gnd.n7247 gnd.n459 173.845
R15205 gnd.n7248 gnd.n7247 173.845
R15206 gnd.n7249 gnd.n7248 173.845
R15207 gnd.n7249 gnd.n453 173.845
R15208 gnd.n7257 gnd.n453 173.845
R15209 gnd.n7258 gnd.n7257 173.845
R15210 gnd.n7259 gnd.n7258 173.845
R15211 gnd.n7259 gnd.n447 173.845
R15212 gnd.n7267 gnd.n447 173.845
R15213 gnd.n7268 gnd.n7267 173.845
R15214 gnd.n7269 gnd.n7268 173.845
R15215 gnd.n7269 gnd.n441 173.845
R15216 gnd.n7277 gnd.n441 173.845
R15217 gnd.n7278 gnd.n7277 173.845
R15218 gnd.n7279 gnd.n7278 173.845
R15219 gnd.n7279 gnd.n435 173.845
R15220 gnd.n7287 gnd.n435 173.845
R15221 gnd.n7288 gnd.n7287 173.845
R15222 gnd.n7289 gnd.n7288 173.845
R15223 gnd.n7289 gnd.n429 173.845
R15224 gnd.n7297 gnd.n429 173.845
R15225 gnd.n7298 gnd.n7297 173.845
R15226 gnd.n7299 gnd.n7298 173.845
R15227 gnd.n7299 gnd.n423 173.845
R15228 gnd.n7307 gnd.n423 173.845
R15229 gnd.n7308 gnd.n7307 173.845
R15230 gnd.n7309 gnd.n7308 173.845
R15231 gnd.n7309 gnd.n417 173.845
R15232 gnd.n7317 gnd.n417 173.845
R15233 gnd.n7318 gnd.n7317 173.845
R15234 gnd.n7319 gnd.n7318 173.845
R15235 gnd.n7319 gnd.n411 173.845
R15236 gnd.n7327 gnd.n411 173.845
R15237 gnd.n7328 gnd.n7327 173.845
R15238 gnd.n7329 gnd.n7328 173.845
R15239 gnd.n7329 gnd.n405 173.845
R15240 gnd.n7339 gnd.n405 173.845
R15241 gnd.n7340 gnd.n7339 173.845
R15242 gnd.n7341 gnd.n7340 173.845
R15243 gnd.n1 gnd.t39 170.774
R15244 gnd.n7 gnd.t230 170.103
R15245 gnd.n6 gnd.t20 170.103
R15246 gnd.n5 gnd.t47 170.103
R15247 gnd.n4 gnd.t61 170.103
R15248 gnd.n3 gnd.t42 170.103
R15249 gnd.n2 gnd.t9 170.103
R15250 gnd.n1 gnd.t66 170.103
R15251 gnd.n3986 gnd.n3985 163.367
R15252 gnd.n3982 gnd.n3981 163.367
R15253 gnd.n3978 gnd.n3977 163.367
R15254 gnd.n3974 gnd.n3973 163.367
R15255 gnd.n3970 gnd.n3969 163.367
R15256 gnd.n3966 gnd.n3965 163.367
R15257 gnd.n3962 gnd.n3961 163.367
R15258 gnd.n3958 gnd.n3957 163.367
R15259 gnd.n3954 gnd.n3953 163.367
R15260 gnd.n3950 gnd.n3949 163.367
R15261 gnd.n3946 gnd.n3945 163.367
R15262 gnd.n3942 gnd.n3941 163.367
R15263 gnd.n3938 gnd.n3937 163.367
R15264 gnd.n3934 gnd.n3933 163.367
R15265 gnd.n3929 gnd.n3928 163.367
R15266 gnd.n3925 gnd.n3924 163.367
R15267 gnd.n4059 gnd.n4058 163.367
R15268 gnd.n4055 gnd.n4054 163.367
R15269 gnd.n4050 gnd.n4049 163.367
R15270 gnd.n4046 gnd.n4045 163.367
R15271 gnd.n4042 gnd.n4041 163.367
R15272 gnd.n4038 gnd.n4037 163.367
R15273 gnd.n4034 gnd.n4033 163.367
R15274 gnd.n4030 gnd.n4029 163.367
R15275 gnd.n4026 gnd.n4025 163.367
R15276 gnd.n4022 gnd.n4021 163.367
R15277 gnd.n4018 gnd.n4017 163.367
R15278 gnd.n4014 gnd.n4013 163.367
R15279 gnd.n4010 gnd.n4009 163.367
R15280 gnd.n4006 gnd.n4005 163.367
R15281 gnd.n4002 gnd.n4001 163.367
R15282 gnd.n3998 gnd.n3997 163.367
R15283 gnd.n3413 gnd.n1492 163.367
R15284 gnd.n3409 gnd.n1492 163.367
R15285 gnd.n3409 gnd.n3403 163.367
R15286 gnd.n3403 gnd.n3402 163.367
R15287 gnd.n3402 gnd.n1501 163.367
R15288 gnd.n3398 gnd.n1501 163.367
R15289 gnd.n3398 gnd.n1508 163.367
R15290 gnd.n3395 gnd.n1508 163.367
R15291 gnd.n3395 gnd.n3394 163.367
R15292 gnd.n3394 gnd.n3388 163.367
R15293 gnd.n3388 gnd.n1518 163.367
R15294 gnd.n3384 gnd.n1518 163.367
R15295 gnd.n3384 gnd.n1526 163.367
R15296 gnd.n3379 gnd.n1526 163.367
R15297 gnd.n3379 gnd.n2325 163.367
R15298 gnd.n3376 gnd.n2325 163.367
R15299 gnd.n3376 gnd.n3375 163.367
R15300 gnd.n3375 gnd.n2320 163.367
R15301 gnd.n3472 gnd.n2320 163.367
R15302 gnd.n3472 gnd.n2314 163.367
R15303 gnd.n3476 gnd.n2314 163.367
R15304 gnd.n3476 gnd.n2306 163.367
R15305 gnd.n3520 gnd.n2306 163.367
R15306 gnd.n3520 gnd.n2304 163.367
R15307 gnd.n3525 gnd.n2304 163.367
R15308 gnd.n3525 gnd.n2299 163.367
R15309 gnd.n2299 gnd.n2288 163.367
R15310 gnd.n3553 gnd.n2288 163.367
R15311 gnd.n3553 gnd.n2289 163.367
R15312 gnd.n2289 gnd.n2279 163.367
R15313 gnd.n3548 gnd.n2279 163.367
R15314 gnd.n3548 gnd.n2271 163.367
R15315 gnd.n3575 gnd.n2271 163.367
R15316 gnd.n3575 gnd.n2263 163.367
R15317 gnd.n3578 gnd.n2263 163.367
R15318 gnd.n3578 gnd.n2255 163.367
R15319 gnd.n3582 gnd.n2255 163.367
R15320 gnd.n3582 gnd.n2247 163.367
R15321 gnd.n3614 gnd.n2247 163.367
R15322 gnd.n3614 gnd.n2240 163.367
R15323 gnd.n3617 gnd.n2240 163.367
R15324 gnd.n3617 gnd.n2234 163.367
R15325 gnd.n3622 gnd.n2234 163.367
R15326 gnd.n3622 gnd.n2224 163.367
R15327 gnd.n2224 gnd.n2217 163.367
R15328 gnd.n3674 gnd.n2217 163.367
R15329 gnd.n3674 gnd.n2215 163.367
R15330 gnd.n3679 gnd.n2215 163.367
R15331 gnd.n3679 gnd.n2206 163.367
R15332 gnd.n2206 gnd.n2197 163.367
R15333 gnd.n3709 gnd.n2197 163.367
R15334 gnd.n3709 gnd.n2194 163.367
R15335 gnd.n3748 gnd.n2194 163.367
R15336 gnd.n3748 gnd.n2195 163.367
R15337 gnd.n3744 gnd.n2195 163.367
R15338 gnd.n3744 gnd.n3743 163.367
R15339 gnd.n3743 gnd.n2176 163.367
R15340 gnd.n2177 gnd.n2176 163.367
R15341 gnd.n2177 gnd.n2168 163.367
R15342 gnd.n3737 gnd.n2168 163.367
R15343 gnd.n3737 gnd.n3734 163.367
R15344 gnd.n3734 gnd.n3733 163.367
R15345 gnd.n3733 gnd.n2153 163.367
R15346 gnd.n2154 gnd.n2153 163.367
R15347 gnd.n2154 gnd.n2146 163.367
R15348 gnd.n3727 gnd.n2146 163.367
R15349 gnd.n3727 gnd.n2139 163.367
R15350 gnd.n3722 gnd.n2139 163.367
R15351 gnd.n3722 gnd.n2134 163.367
R15352 gnd.n3719 gnd.n2134 163.367
R15353 gnd.n3719 gnd.n2121 163.367
R15354 gnd.n3716 gnd.n2121 163.367
R15355 gnd.n3716 gnd.n2114 163.367
R15356 gnd.n3869 gnd.n2114 163.367
R15357 gnd.n3869 gnd.n2111 163.367
R15358 gnd.n3879 gnd.n2111 163.367
R15359 gnd.n3879 gnd.n2104 163.367
R15360 gnd.n3875 gnd.n2104 163.367
R15361 gnd.n3875 gnd.n2097 163.367
R15362 gnd.n2097 gnd.n2090 163.367
R15363 gnd.n3993 gnd.n2090 163.367
R15364 gnd.n1467 gnd.n1466 163.367
R15365 gnd.n4772 gnd.n1466 163.367
R15366 gnd.n4770 gnd.n4769 163.367
R15367 gnd.n4766 gnd.n4765 163.367
R15368 gnd.n4762 gnd.n4761 163.367
R15369 gnd.n4758 gnd.n4757 163.367
R15370 gnd.n4754 gnd.n4753 163.367
R15371 gnd.n4750 gnd.n4749 163.367
R15372 gnd.n4746 gnd.n4745 163.367
R15373 gnd.n4742 gnd.n4741 163.367
R15374 gnd.n4738 gnd.n4737 163.367
R15375 gnd.n4734 gnd.n4733 163.367
R15376 gnd.n4730 gnd.n4729 163.367
R15377 gnd.n4726 gnd.n4725 163.367
R15378 gnd.n4722 gnd.n4721 163.367
R15379 gnd.n4718 gnd.n4717 163.367
R15380 gnd.n4781 gnd.n1432 163.367
R15381 gnd.n3312 gnd.n3311 163.367
R15382 gnd.n3317 gnd.n3316 163.367
R15383 gnd.n3321 gnd.n3320 163.367
R15384 gnd.n3325 gnd.n3324 163.367
R15385 gnd.n3329 gnd.n3328 163.367
R15386 gnd.n3333 gnd.n3332 163.367
R15387 gnd.n3337 gnd.n3336 163.367
R15388 gnd.n3341 gnd.n3340 163.367
R15389 gnd.n3345 gnd.n3344 163.367
R15390 gnd.n3349 gnd.n3348 163.367
R15391 gnd.n3353 gnd.n3352 163.367
R15392 gnd.n3357 gnd.n3356 163.367
R15393 gnd.n3361 gnd.n3360 163.367
R15394 gnd.n3365 gnd.n3364 163.367
R15395 gnd.n3369 gnd.n3368 163.367
R15396 gnd.n4710 gnd.n1468 163.367
R15397 gnd.n4710 gnd.n1490 163.367
R15398 gnd.n3405 gnd.n1490 163.367
R15399 gnd.n3405 gnd.n1503 163.367
R15400 gnd.n4700 gnd.n1503 163.367
R15401 gnd.n4700 gnd.n1504 163.367
R15402 gnd.n4696 gnd.n1504 163.367
R15403 gnd.n4696 gnd.n1507 163.367
R15404 gnd.n3392 gnd.n1507 163.367
R15405 gnd.n3392 gnd.n1520 163.367
R15406 gnd.n4686 gnd.n1520 163.367
R15407 gnd.n4686 gnd.n1521 163.367
R15408 gnd.n4682 gnd.n1521 163.367
R15409 gnd.n4682 gnd.n1524 163.367
R15410 gnd.n3464 gnd.n1524 163.367
R15411 gnd.n3465 gnd.n3464 163.367
R15412 gnd.n3465 gnd.n2322 163.367
R15413 gnd.n3469 gnd.n2322 163.367
R15414 gnd.n3469 gnd.n2316 163.367
R15415 gnd.n3506 gnd.n2316 163.367
R15416 gnd.n3506 gnd.n2317 163.367
R15417 gnd.n3502 gnd.n2317 163.367
R15418 gnd.n3502 gnd.n2302 163.367
R15419 gnd.n3530 gnd.n2302 163.367
R15420 gnd.n3530 gnd.n2300 163.367
R15421 gnd.n3534 gnd.n2300 163.367
R15422 gnd.n3534 gnd.n2285 163.367
R15423 gnd.n3555 gnd.n2285 163.367
R15424 gnd.n3555 gnd.n2282 163.367
R15425 gnd.n3562 gnd.n2282 163.367
R15426 gnd.n3562 gnd.n2283 163.367
R15427 gnd.n3558 gnd.n2283 163.367
R15428 gnd.n3558 gnd.n2261 163.367
R15429 gnd.n3594 gnd.n2261 163.367
R15430 gnd.n3594 gnd.n2258 163.367
R15431 gnd.n3601 gnd.n2258 163.367
R15432 gnd.n3601 gnd.n2259 163.367
R15433 gnd.n3597 gnd.n2259 163.367
R15434 gnd.n3597 gnd.n2238 163.367
R15435 gnd.n3649 gnd.n2238 163.367
R15436 gnd.n3649 gnd.n2236 163.367
R15437 gnd.n3653 gnd.n2236 163.367
R15438 gnd.n3653 gnd.n2223 163.367
R15439 gnd.n3667 gnd.n2223 163.367
R15440 gnd.n3667 gnd.n2220 163.367
R15441 gnd.n3672 gnd.n2220 163.367
R15442 gnd.n3672 gnd.n2221 163.367
R15443 gnd.n2221 gnd.n2204 163.367
R15444 gnd.n3695 gnd.n2204 163.367
R15445 gnd.n3695 gnd.n2199 163.367
R15446 gnd.n3707 gnd.n2199 163.367
R15447 gnd.n3707 gnd.n2202 163.367
R15448 gnd.n2202 gnd.n2191 163.367
R15449 gnd.n3702 gnd.n2191 163.367
R15450 gnd.n3702 gnd.n3699 163.367
R15451 gnd.n3699 gnd.n2174 163.367
R15452 gnd.n3770 gnd.n2174 163.367
R15453 gnd.n3770 gnd.n2171 163.367
R15454 gnd.n3777 gnd.n2171 163.367
R15455 gnd.n3777 gnd.n2172 163.367
R15456 gnd.n3773 gnd.n2172 163.367
R15457 gnd.n3773 gnd.n2151 163.367
R15458 gnd.n3804 gnd.n2151 163.367
R15459 gnd.n3804 gnd.n2149 163.367
R15460 gnd.n3808 gnd.n2149 163.367
R15461 gnd.n3808 gnd.n2137 163.367
R15462 gnd.n3820 gnd.n2137 163.367
R15463 gnd.n3820 gnd.n2135 163.367
R15464 gnd.n3824 gnd.n2135 163.367
R15465 gnd.n3824 gnd.n2122 163.367
R15466 gnd.n3857 gnd.n2122 163.367
R15467 gnd.n3857 gnd.n2123 163.367
R15468 gnd.n3853 gnd.n2123 163.367
R15469 gnd.n3853 gnd.n2109 163.367
R15470 gnd.n3884 gnd.n2109 163.367
R15471 gnd.n3884 gnd.n2107 163.367
R15472 gnd.n3888 gnd.n2107 163.367
R15473 gnd.n3888 gnd.n2095 163.367
R15474 gnd.n3900 gnd.n2095 163.367
R15475 gnd.n3900 gnd.n2092 163.367
R15476 gnd.n3991 gnd.n2092 163.367
R15477 gnd.n3921 gnd.n3920 156.462
R15478 gnd.n6275 gnd.n6243 153.042
R15479 gnd.n6339 gnd.n6338 152.079
R15480 gnd.n6307 gnd.n6306 152.079
R15481 gnd.n6275 gnd.n6274 152.079
R15482 gnd.n1481 gnd.n1480 152
R15483 gnd.n1482 gnd.n1471 152
R15484 gnd.n1484 gnd.n1483 152
R15485 gnd.n1486 gnd.n1469 152
R15486 gnd.n1488 gnd.n1487 152
R15487 gnd.n3919 gnd.n3903 152
R15488 gnd.n3911 gnd.n3904 152
R15489 gnd.n3910 gnd.n3909 152
R15490 gnd.n3908 gnd.n3905 152
R15491 gnd.n3906 gnd.t294 150.546
R15492 gnd.t58 gnd.n6317 147.661
R15493 gnd.t64 gnd.n6285 147.661
R15494 gnd.t18 gnd.n6253 147.661
R15495 gnd.t237 gnd.n6222 147.661
R15496 gnd.t51 gnd.n6190 147.661
R15497 gnd.t239 gnd.n6158 147.661
R15498 gnd.t16 gnd.n6126 147.661
R15499 gnd.t53 gnd.n6095 147.661
R15500 gnd.n2086 gnd.n2067 143.351
R15501 gnd.n1448 gnd.n1431 143.351
R15502 gnd.n4780 gnd.n1431 143.351
R15503 gnd.n7341 gnd.n212 132.349
R15504 gnd.n1478 gnd.t348 130.484
R15505 gnd.n1487 gnd.t261 126.766
R15506 gnd.n1485 gnd.t310 126.766
R15507 gnd.n1471 gnd.t244 126.766
R15508 gnd.n1479 gnd.t297 126.766
R15509 gnd.n3907 gnd.t357 126.766
R15510 gnd.n3909 gnd.t247 126.766
R15511 gnd.n3918 gnd.t258 126.766
R15512 gnd.n3920 gnd.t329 126.766
R15513 gnd.n4467 gnd.n1750 108.609
R15514 gnd.n4783 gnd.n4782 108.609
R15515 gnd.n6334 gnd.n6333 104.615
R15516 gnd.n6333 gnd.n6311 104.615
R15517 gnd.n6326 gnd.n6311 104.615
R15518 gnd.n6326 gnd.n6325 104.615
R15519 gnd.n6325 gnd.n6315 104.615
R15520 gnd.n6318 gnd.n6315 104.615
R15521 gnd.n6302 gnd.n6301 104.615
R15522 gnd.n6301 gnd.n6279 104.615
R15523 gnd.n6294 gnd.n6279 104.615
R15524 gnd.n6294 gnd.n6293 104.615
R15525 gnd.n6293 gnd.n6283 104.615
R15526 gnd.n6286 gnd.n6283 104.615
R15527 gnd.n6270 gnd.n6269 104.615
R15528 gnd.n6269 gnd.n6247 104.615
R15529 gnd.n6262 gnd.n6247 104.615
R15530 gnd.n6262 gnd.n6261 104.615
R15531 gnd.n6261 gnd.n6251 104.615
R15532 gnd.n6254 gnd.n6251 104.615
R15533 gnd.n6239 gnd.n6238 104.615
R15534 gnd.n6238 gnd.n6216 104.615
R15535 gnd.n6231 gnd.n6216 104.615
R15536 gnd.n6231 gnd.n6230 104.615
R15537 gnd.n6230 gnd.n6220 104.615
R15538 gnd.n6223 gnd.n6220 104.615
R15539 gnd.n6207 gnd.n6206 104.615
R15540 gnd.n6206 gnd.n6184 104.615
R15541 gnd.n6199 gnd.n6184 104.615
R15542 gnd.n6199 gnd.n6198 104.615
R15543 gnd.n6198 gnd.n6188 104.615
R15544 gnd.n6191 gnd.n6188 104.615
R15545 gnd.n6175 gnd.n6174 104.615
R15546 gnd.n6174 gnd.n6152 104.615
R15547 gnd.n6167 gnd.n6152 104.615
R15548 gnd.n6167 gnd.n6166 104.615
R15549 gnd.n6166 gnd.n6156 104.615
R15550 gnd.n6159 gnd.n6156 104.615
R15551 gnd.n6143 gnd.n6142 104.615
R15552 gnd.n6142 gnd.n6120 104.615
R15553 gnd.n6135 gnd.n6120 104.615
R15554 gnd.n6135 gnd.n6134 104.615
R15555 gnd.n6134 gnd.n6124 104.615
R15556 gnd.n6127 gnd.n6124 104.615
R15557 gnd.n6112 gnd.n6111 104.615
R15558 gnd.n6111 gnd.n6089 104.615
R15559 gnd.n6104 gnd.n6089 104.615
R15560 gnd.n6104 gnd.n6103 104.615
R15561 gnd.n6103 gnd.n6093 104.615
R15562 gnd.n6096 gnd.n6093 104.615
R15563 gnd.n5689 gnd.t319 100.632
R15564 gnd.n5123 gnd.t346 100.632
R15565 gnd.n7595 gnd.n219 99.6594
R15566 gnd.n7593 gnd.n7592 99.6594
R15567 gnd.n7588 gnd.n226 99.6594
R15568 gnd.n7586 gnd.n7585 99.6594
R15569 gnd.n7581 gnd.n233 99.6594
R15570 gnd.n7579 gnd.n7578 99.6594
R15571 gnd.n7574 gnd.n240 99.6594
R15572 gnd.n7572 gnd.n7571 99.6594
R15573 gnd.n7564 gnd.n247 99.6594
R15574 gnd.n7562 gnd.n7561 99.6594
R15575 gnd.n7557 gnd.n254 99.6594
R15576 gnd.n7555 gnd.n7554 99.6594
R15577 gnd.n7550 gnd.n261 99.6594
R15578 gnd.n7548 gnd.n7547 99.6594
R15579 gnd.n7543 gnd.n268 99.6594
R15580 gnd.n7541 gnd.n7540 99.6594
R15581 gnd.n7536 gnd.n275 99.6594
R15582 gnd.n7534 gnd.n7533 99.6594
R15583 gnd.n285 gnd.n284 99.6594
R15584 gnd.n7525 gnd.n7524 99.6594
R15585 gnd.n7522 gnd.n7521 99.6594
R15586 gnd.n7517 gnd.n293 99.6594
R15587 gnd.n7515 gnd.n7514 99.6594
R15588 gnd.n7510 gnd.n300 99.6594
R15589 gnd.n7508 gnd.n7507 99.6594
R15590 gnd.n7503 gnd.n307 99.6594
R15591 gnd.n7501 gnd.n7500 99.6594
R15592 gnd.n7496 gnd.n316 99.6594
R15593 gnd.n7494 gnd.n7493 99.6594
R15594 gnd.n4519 gnd.n4518 99.6594
R15595 gnd.n4513 gnd.n1677 99.6594
R15596 gnd.n4510 gnd.n1678 99.6594
R15597 gnd.n4506 gnd.n1679 99.6594
R15598 gnd.n4502 gnd.n1680 99.6594
R15599 gnd.n4498 gnd.n1681 99.6594
R15600 gnd.n4494 gnd.n1682 99.6594
R15601 gnd.n4490 gnd.n1683 99.6594
R15602 gnd.n4486 gnd.n1684 99.6594
R15603 gnd.n4481 gnd.n1685 99.6594
R15604 gnd.n4477 gnd.n1686 99.6594
R15605 gnd.n4473 gnd.n1687 99.6594
R15606 gnd.n4469 gnd.n1688 99.6594
R15607 gnd.n4464 gnd.n1690 99.6594
R15608 gnd.n4460 gnd.n1691 99.6594
R15609 gnd.n4456 gnd.n1692 99.6594
R15610 gnd.n4452 gnd.n1693 99.6594
R15611 gnd.n4448 gnd.n1694 99.6594
R15612 gnd.n4444 gnd.n1695 99.6594
R15613 gnd.n4440 gnd.n1696 99.6594
R15614 gnd.n4436 gnd.n1697 99.6594
R15615 gnd.n4432 gnd.n1698 99.6594
R15616 gnd.n4428 gnd.n1699 99.6594
R15617 gnd.n4424 gnd.n1700 99.6594
R15618 gnd.n4420 gnd.n1701 99.6594
R15619 gnd.n4416 gnd.n1702 99.6594
R15620 gnd.n4412 gnd.n1703 99.6594
R15621 gnd.n4408 gnd.n1704 99.6594
R15622 gnd.n4826 gnd.n4825 99.6594
R15623 gnd.n4823 gnd.n4822 99.6594
R15624 gnd.n4818 gnd.n1390 99.6594
R15625 gnd.n4816 gnd.n4815 99.6594
R15626 gnd.n4811 gnd.n1397 99.6594
R15627 gnd.n4809 gnd.n4808 99.6594
R15628 gnd.n4804 gnd.n1404 99.6594
R15629 gnd.n4802 gnd.n4801 99.6594
R15630 gnd.n4796 gnd.n1413 99.6594
R15631 gnd.n4794 gnd.n4793 99.6594
R15632 gnd.n4789 gnd.n1420 99.6594
R15633 gnd.n4787 gnd.n4786 99.6594
R15634 gnd.n2478 gnd.n2477 99.6594
R15635 gnd.n2482 gnd.n2480 99.6594
R15636 gnd.n2488 gnd.n2472 99.6594
R15637 gnd.n2492 gnd.n2490 99.6594
R15638 gnd.n2498 gnd.n2468 99.6594
R15639 gnd.n2502 gnd.n2500 99.6594
R15640 gnd.n2508 gnd.n2462 99.6594
R15641 gnd.n2512 gnd.n2510 99.6594
R15642 gnd.n2518 gnd.n2458 99.6594
R15643 gnd.n2522 gnd.n2520 99.6594
R15644 gnd.n2528 gnd.n2454 99.6594
R15645 gnd.n2532 gnd.n2530 99.6594
R15646 gnd.n2538 gnd.n2450 99.6594
R15647 gnd.n2542 gnd.n2540 99.6594
R15648 gnd.n2548 gnd.n2446 99.6594
R15649 gnd.n2551 gnd.n2550 99.6594
R15650 gnd.n5091 gnd.n5090 99.6594
R15651 gnd.n5085 gnd.n1030 99.6594
R15652 gnd.n5082 gnd.n1031 99.6594
R15653 gnd.n5078 gnd.n1032 99.6594
R15654 gnd.n5074 gnd.n1033 99.6594
R15655 gnd.n5070 gnd.n1034 99.6594
R15656 gnd.n5066 gnd.n1035 99.6594
R15657 gnd.n5062 gnd.n1036 99.6594
R15658 gnd.n5058 gnd.n1037 99.6594
R15659 gnd.n5053 gnd.n1038 99.6594
R15660 gnd.n5049 gnd.n1039 99.6594
R15661 gnd.n5045 gnd.n1040 99.6594
R15662 gnd.n5041 gnd.n1041 99.6594
R15663 gnd.n5037 gnd.n1042 99.6594
R15664 gnd.n5033 gnd.n1043 99.6594
R15665 gnd.n5029 gnd.n1044 99.6594
R15666 gnd.n5025 gnd.n1045 99.6594
R15667 gnd.n5021 gnd.n1046 99.6594
R15668 gnd.n5017 gnd.n1047 99.6594
R15669 gnd.n5013 gnd.n1048 99.6594
R15670 gnd.n5009 gnd.n1049 99.6594
R15671 gnd.n5005 gnd.n1050 99.6594
R15672 gnd.n5001 gnd.n1051 99.6594
R15673 gnd.n4997 gnd.n1052 99.6594
R15674 gnd.n4993 gnd.n1053 99.6594
R15675 gnd.n4989 gnd.n1054 99.6594
R15676 gnd.n4985 gnd.n1055 99.6594
R15677 gnd.n4981 gnd.n1056 99.6594
R15678 gnd.n4977 gnd.n1057 99.6594
R15679 gnd.n6465 gnd.n5103 99.6594
R15680 gnd.n6463 gnd.n6462 99.6594
R15681 gnd.n6458 gnd.n5110 99.6594
R15682 gnd.n6456 gnd.n6455 99.6594
R15683 gnd.n6451 gnd.n5117 99.6594
R15684 gnd.n6449 gnd.n6448 99.6594
R15685 gnd.n6444 gnd.n5126 99.6594
R15686 gnd.n6442 gnd.n6441 99.6594
R15687 gnd.n5722 gnd.n5721 99.6594
R15688 gnd.n5716 gnd.n5664 99.6594
R15689 gnd.n5713 gnd.n5665 99.6594
R15690 gnd.n5709 gnd.n5666 99.6594
R15691 gnd.n5705 gnd.n5667 99.6594
R15692 gnd.n5701 gnd.n5668 99.6594
R15693 gnd.n5697 gnd.n5669 99.6594
R15694 gnd.n5693 gnd.n5670 99.6594
R15695 gnd.n7485 gnd.n322 99.6594
R15696 gnd.n7483 gnd.n7482 99.6594
R15697 gnd.n7478 gnd.n329 99.6594
R15698 gnd.n7476 gnd.n7475 99.6594
R15699 gnd.n7471 gnd.n336 99.6594
R15700 gnd.n7469 gnd.n7468 99.6594
R15701 gnd.n7464 gnd.n343 99.6594
R15702 gnd.n7462 gnd.n7461 99.6594
R15703 gnd.n348 gnd.n347 99.6594
R15704 gnd.n1789 gnd.n1705 99.6594
R15705 gnd.n1707 gnd.n1631 99.6594
R15706 gnd.n1708 gnd.n1638 99.6594
R15707 gnd.n1710 gnd.n1709 99.6594
R15708 gnd.n1712 gnd.n1647 99.6594
R15709 gnd.n1713 gnd.n1654 99.6594
R15710 gnd.n1715 gnd.n1714 99.6594
R15711 gnd.n1717 gnd.n1663 99.6594
R15712 gnd.n4521 gnd.n1672 99.6594
R15713 gnd.n6433 gnd.n5133 99.6594
R15714 gnd.n6431 gnd.n6430 99.6594
R15715 gnd.n6426 gnd.n5140 99.6594
R15716 gnd.n6424 gnd.n6423 99.6594
R15717 gnd.n6419 gnd.n5147 99.6594
R15718 gnd.n6417 gnd.n6416 99.6594
R15719 gnd.n6412 gnd.n5154 99.6594
R15720 gnd.n6410 gnd.n6409 99.6594
R15721 gnd.n6405 gnd.n5161 99.6594
R15722 gnd.n6403 gnd.n6402 99.6594
R15723 gnd.n6398 gnd.n5170 99.6594
R15724 gnd.n6396 gnd.n6395 99.6594
R15725 gnd.n6391 gnd.n6390 99.6594
R15726 gnd.n5594 gnd.n5504 99.6594
R15727 gnd.n5592 gnd.n5507 99.6594
R15728 gnd.n5588 gnd.n5587 99.6594
R15729 gnd.n5581 gnd.n5512 99.6594
R15730 gnd.n5580 gnd.n5579 99.6594
R15731 gnd.n5573 gnd.n5518 99.6594
R15732 gnd.n5572 gnd.n5571 99.6594
R15733 gnd.n5565 gnd.n5524 99.6594
R15734 gnd.n5564 gnd.n5563 99.6594
R15735 gnd.n5557 gnd.n5530 99.6594
R15736 gnd.n5556 gnd.n5555 99.6594
R15737 gnd.n5548 gnd.n5536 99.6594
R15738 gnd.n5547 gnd.n5546 99.6594
R15739 gnd.n2563 gnd.n2562 99.6594
R15740 gnd.n2574 gnd.n2573 99.6594
R15741 gnd.n2583 gnd.n2582 99.6594
R15742 gnd.n2586 gnd.n2585 99.6594
R15743 gnd.n2597 gnd.n2596 99.6594
R15744 gnd.n2606 gnd.n2605 99.6594
R15745 gnd.n2609 gnd.n2608 99.6594
R15746 gnd.n2621 gnd.n2620 99.6594
R15747 gnd.n3161 gnd.n3160 99.6594
R15748 gnd.n2763 gnd.n1058 99.6594
R15749 gnd.n2767 gnd.n1059 99.6594
R15750 gnd.n2773 gnd.n1060 99.6594
R15751 gnd.n2777 gnd.n1061 99.6594
R15752 gnd.n2783 gnd.n1062 99.6594
R15753 gnd.n2787 gnd.n1063 99.6594
R15754 gnd.n2793 gnd.n1064 99.6594
R15755 gnd.n2797 gnd.n1065 99.6594
R15756 gnd.n2754 gnd.n1066 99.6594
R15757 gnd.n2766 gnd.n1058 99.6594
R15758 gnd.n2772 gnd.n1059 99.6594
R15759 gnd.n2776 gnd.n1060 99.6594
R15760 gnd.n2782 gnd.n1061 99.6594
R15761 gnd.n2786 gnd.n1062 99.6594
R15762 gnd.n2792 gnd.n1063 99.6594
R15763 gnd.n2796 gnd.n1064 99.6594
R15764 gnd.n2753 gnd.n1065 99.6594
R15765 gnd.n2749 gnd.n1066 99.6594
R15766 gnd.n3160 gnd.n2625 99.6594
R15767 gnd.n2620 gnd.n2619 99.6594
R15768 gnd.n2608 gnd.n2607 99.6594
R15769 gnd.n2605 gnd.n2598 99.6594
R15770 gnd.n2596 gnd.n2595 99.6594
R15771 gnd.n2585 gnd.n2584 99.6594
R15772 gnd.n2582 gnd.n2575 99.6594
R15773 gnd.n2573 gnd.n2572 99.6594
R15774 gnd.n2562 gnd.n2561 99.6594
R15775 gnd.n5595 gnd.n5594 99.6594
R15776 gnd.n5589 gnd.n5507 99.6594
R15777 gnd.n5587 gnd.n5586 99.6594
R15778 gnd.n5582 gnd.n5581 99.6594
R15779 gnd.n5579 gnd.n5578 99.6594
R15780 gnd.n5574 gnd.n5573 99.6594
R15781 gnd.n5571 gnd.n5570 99.6594
R15782 gnd.n5566 gnd.n5565 99.6594
R15783 gnd.n5563 gnd.n5562 99.6594
R15784 gnd.n5558 gnd.n5557 99.6594
R15785 gnd.n5555 gnd.n5554 99.6594
R15786 gnd.n5549 gnd.n5548 99.6594
R15787 gnd.n5546 gnd.n5502 99.6594
R15788 gnd.n6390 gnd.n5172 99.6594
R15789 gnd.n6397 gnd.n6396 99.6594
R15790 gnd.n5170 gnd.n5162 99.6594
R15791 gnd.n6404 gnd.n6403 99.6594
R15792 gnd.n5161 gnd.n5155 99.6594
R15793 gnd.n6411 gnd.n6410 99.6594
R15794 gnd.n5154 gnd.n5148 99.6594
R15795 gnd.n6418 gnd.n6417 99.6594
R15796 gnd.n5147 gnd.n5141 99.6594
R15797 gnd.n6425 gnd.n6424 99.6594
R15798 gnd.n5140 gnd.n5134 99.6594
R15799 gnd.n6432 gnd.n6431 99.6594
R15800 gnd.n5133 gnd.n5130 99.6594
R15801 gnd.n1705 gnd.n1630 99.6594
R15802 gnd.n1707 gnd.n1706 99.6594
R15803 gnd.n1708 gnd.n1639 99.6594
R15804 gnd.n1710 gnd.n1646 99.6594
R15805 gnd.n1712 gnd.n1711 99.6594
R15806 gnd.n1713 gnd.n1655 99.6594
R15807 gnd.n1715 gnd.n1662 99.6594
R15808 gnd.n1717 gnd.n1716 99.6594
R15809 gnd.n4522 gnd.n4521 99.6594
R15810 gnd.n347 gnd.n344 99.6594
R15811 gnd.n7463 gnd.n7462 99.6594
R15812 gnd.n343 gnd.n337 99.6594
R15813 gnd.n7470 gnd.n7469 99.6594
R15814 gnd.n336 gnd.n330 99.6594
R15815 gnd.n7477 gnd.n7476 99.6594
R15816 gnd.n329 gnd.n323 99.6594
R15817 gnd.n7484 gnd.n7483 99.6594
R15818 gnd.n322 gnd.n319 99.6594
R15819 gnd.n5722 gnd.n5672 99.6594
R15820 gnd.n5714 gnd.n5664 99.6594
R15821 gnd.n5710 gnd.n5665 99.6594
R15822 gnd.n5706 gnd.n5666 99.6594
R15823 gnd.n5702 gnd.n5667 99.6594
R15824 gnd.n5698 gnd.n5668 99.6594
R15825 gnd.n5694 gnd.n5669 99.6594
R15826 gnd.n5670 gnd.n5464 99.6594
R15827 gnd.n6443 gnd.n6442 99.6594
R15828 gnd.n5126 gnd.n5118 99.6594
R15829 gnd.n6450 gnd.n6449 99.6594
R15830 gnd.n5117 gnd.n5111 99.6594
R15831 gnd.n6457 gnd.n6456 99.6594
R15832 gnd.n5110 gnd.n5104 99.6594
R15833 gnd.n6464 gnd.n6463 99.6594
R15834 gnd.n5103 gnd.n5100 99.6594
R15835 gnd.n5091 gnd.n1070 99.6594
R15836 gnd.n5083 gnd.n1030 99.6594
R15837 gnd.n5079 gnd.n1031 99.6594
R15838 gnd.n5075 gnd.n1032 99.6594
R15839 gnd.n5071 gnd.n1033 99.6594
R15840 gnd.n5067 gnd.n1034 99.6594
R15841 gnd.n5063 gnd.n1035 99.6594
R15842 gnd.n5059 gnd.n1036 99.6594
R15843 gnd.n5054 gnd.n1037 99.6594
R15844 gnd.n5050 gnd.n1038 99.6594
R15845 gnd.n5046 gnd.n1039 99.6594
R15846 gnd.n5042 gnd.n1040 99.6594
R15847 gnd.n5038 gnd.n1041 99.6594
R15848 gnd.n5034 gnd.n1042 99.6594
R15849 gnd.n5030 gnd.n1043 99.6594
R15850 gnd.n5026 gnd.n1044 99.6594
R15851 gnd.n5022 gnd.n1045 99.6594
R15852 gnd.n5018 gnd.n1046 99.6594
R15853 gnd.n5014 gnd.n1047 99.6594
R15854 gnd.n5010 gnd.n1048 99.6594
R15855 gnd.n5006 gnd.n1049 99.6594
R15856 gnd.n5002 gnd.n1050 99.6594
R15857 gnd.n4998 gnd.n1051 99.6594
R15858 gnd.n4994 gnd.n1052 99.6594
R15859 gnd.n4990 gnd.n1053 99.6594
R15860 gnd.n4986 gnd.n1054 99.6594
R15861 gnd.n4982 gnd.n1055 99.6594
R15862 gnd.n4978 gnd.n1056 99.6594
R15863 gnd.n1140 gnd.n1057 99.6594
R15864 gnd.n2550 gnd.n2549 99.6594
R15865 gnd.n2541 gnd.n2446 99.6594
R15866 gnd.n2540 gnd.n2539 99.6594
R15867 gnd.n2531 gnd.n2450 99.6594
R15868 gnd.n2530 gnd.n2529 99.6594
R15869 gnd.n2521 gnd.n2454 99.6594
R15870 gnd.n2520 gnd.n2519 99.6594
R15871 gnd.n2511 gnd.n2458 99.6594
R15872 gnd.n2510 gnd.n2509 99.6594
R15873 gnd.n2501 gnd.n2462 99.6594
R15874 gnd.n2500 gnd.n2499 99.6594
R15875 gnd.n2491 gnd.n2468 99.6594
R15876 gnd.n2490 gnd.n2489 99.6594
R15877 gnd.n2481 gnd.n2472 99.6594
R15878 gnd.n2480 gnd.n2479 99.6594
R15879 gnd.n1426 gnd.n1421 99.6594
R15880 gnd.n4788 gnd.n4787 99.6594
R15881 gnd.n1420 gnd.n1414 99.6594
R15882 gnd.n4795 gnd.n4794 99.6594
R15883 gnd.n1413 gnd.n1405 99.6594
R15884 gnd.n4803 gnd.n4802 99.6594
R15885 gnd.n1404 gnd.n1398 99.6594
R15886 gnd.n4810 gnd.n4809 99.6594
R15887 gnd.n1397 gnd.n1391 99.6594
R15888 gnd.n4817 gnd.n4816 99.6594
R15889 gnd.n1390 gnd.n1383 99.6594
R15890 gnd.n4824 gnd.n4823 99.6594
R15891 gnd.n4827 gnd.n4826 99.6594
R15892 gnd.n4519 gnd.n1720 99.6594
R15893 gnd.n4511 gnd.n1677 99.6594
R15894 gnd.n4507 gnd.n1678 99.6594
R15895 gnd.n4503 gnd.n1679 99.6594
R15896 gnd.n4499 gnd.n1680 99.6594
R15897 gnd.n4495 gnd.n1681 99.6594
R15898 gnd.n4491 gnd.n1682 99.6594
R15899 gnd.n4487 gnd.n1683 99.6594
R15900 gnd.n4482 gnd.n1684 99.6594
R15901 gnd.n4478 gnd.n1685 99.6594
R15902 gnd.n4474 gnd.n1686 99.6594
R15903 gnd.n4470 gnd.n1687 99.6594
R15904 gnd.n4465 gnd.n1689 99.6594
R15905 gnd.n4461 gnd.n1690 99.6594
R15906 gnd.n4457 gnd.n1691 99.6594
R15907 gnd.n4453 gnd.n1692 99.6594
R15908 gnd.n4449 gnd.n1693 99.6594
R15909 gnd.n4445 gnd.n1694 99.6594
R15910 gnd.n4441 gnd.n1695 99.6594
R15911 gnd.n4437 gnd.n1696 99.6594
R15912 gnd.n4433 gnd.n1697 99.6594
R15913 gnd.n4429 gnd.n1698 99.6594
R15914 gnd.n4425 gnd.n1699 99.6594
R15915 gnd.n4421 gnd.n1700 99.6594
R15916 gnd.n4417 gnd.n1701 99.6594
R15917 gnd.n4413 gnd.n1702 99.6594
R15918 gnd.n4409 gnd.n1703 99.6594
R15919 gnd.n4401 gnd.n1704 99.6594
R15920 gnd.n7495 gnd.n7494 99.6594
R15921 gnd.n316 gnd.n308 99.6594
R15922 gnd.n7502 gnd.n7501 99.6594
R15923 gnd.n307 gnd.n301 99.6594
R15924 gnd.n7509 gnd.n7508 99.6594
R15925 gnd.n300 gnd.n294 99.6594
R15926 gnd.n7516 gnd.n7515 99.6594
R15927 gnd.n293 gnd.n287 99.6594
R15928 gnd.n7523 gnd.n7522 99.6594
R15929 gnd.n7526 gnd.n7525 99.6594
R15930 gnd.n284 gnd.n276 99.6594
R15931 gnd.n7535 gnd.n7534 99.6594
R15932 gnd.n275 gnd.n269 99.6594
R15933 gnd.n7542 gnd.n7541 99.6594
R15934 gnd.n268 gnd.n262 99.6594
R15935 gnd.n7549 gnd.n7548 99.6594
R15936 gnd.n261 gnd.n255 99.6594
R15937 gnd.n7556 gnd.n7555 99.6594
R15938 gnd.n254 gnd.n248 99.6594
R15939 gnd.n7563 gnd.n7562 99.6594
R15940 gnd.n247 gnd.n241 99.6594
R15941 gnd.n7573 gnd.n7572 99.6594
R15942 gnd.n240 gnd.n234 99.6594
R15943 gnd.n7580 gnd.n7579 99.6594
R15944 gnd.n233 gnd.n227 99.6594
R15945 gnd.n7587 gnd.n7586 99.6594
R15946 gnd.n226 gnd.n220 99.6594
R15947 gnd.n7594 gnd.n7593 99.6594
R15948 gnd.n219 gnd.n216 99.6594
R15949 gnd.n3223 gnd.n3222 99.6594
R15950 gnd.n2434 gnd.n2420 99.6594
R15951 gnd.n2438 gnd.n2421 99.6594
R15952 gnd.n2440 gnd.n2422 99.6594
R15953 gnd.n2557 gnd.n2423 99.6594
R15954 gnd.n2567 gnd.n2424 99.6594
R15955 gnd.n2569 gnd.n2425 99.6594
R15956 gnd.n2579 gnd.n2426 99.6594
R15957 gnd.n2590 gnd.n2427 99.6594
R15958 gnd.n2592 gnd.n2428 99.6594
R15959 gnd.n2602 gnd.n2429 99.6594
R15960 gnd.n2613 gnd.n2430 99.6594
R15961 gnd.n3149 gnd.n2431 99.6594
R15962 gnd.n3153 gnd.n2432 99.6594
R15963 gnd.n3222 gnd.n2418 99.6594
R15964 gnd.n2437 gnd.n2420 99.6594
R15965 gnd.n2439 gnd.n2421 99.6594
R15966 gnd.n2556 gnd.n2422 99.6594
R15967 gnd.n2566 gnd.n2423 99.6594
R15968 gnd.n2568 gnd.n2424 99.6594
R15969 gnd.n2578 gnd.n2425 99.6594
R15970 gnd.n2589 gnd.n2426 99.6594
R15971 gnd.n2591 gnd.n2427 99.6594
R15972 gnd.n2601 gnd.n2428 99.6594
R15973 gnd.n2612 gnd.n2429 99.6594
R15974 gnd.n2614 gnd.n2430 99.6594
R15975 gnd.n3152 gnd.n2431 99.6594
R15976 gnd.n3154 gnd.n2432 99.6594
R15977 gnd.n1979 gnd.n1615 99.6594
R15978 gnd.n1981 gnd.n1980 99.6594
R15979 gnd.n1982 gnd.n1620 99.6594
R15980 gnd.n1984 gnd.n1983 99.6594
R15981 gnd.n1985 gnd.n1626 99.6594
R15982 gnd.n1987 gnd.n1634 99.6594
R15983 gnd.n1989 gnd.n1988 99.6594
R15984 gnd.n1990 gnd.n1643 99.6594
R15985 gnd.n1992 gnd.n1650 99.6594
R15986 gnd.n1994 gnd.n1993 99.6594
R15987 gnd.n1995 gnd.n1659 99.6594
R15988 gnd.n1997 gnd.n1666 99.6594
R15989 gnd.n2001 gnd.n1999 99.6594
R15990 gnd.n4179 gnd.n1976 99.6594
R15991 gnd.n1997 gnd.n1996 99.6594
R15992 gnd.n1995 gnd.n1658 99.6594
R15993 gnd.n1994 gnd.n1651 99.6594
R15994 gnd.n1992 gnd.n1991 99.6594
R15995 gnd.n1990 gnd.n1642 99.6594
R15996 gnd.n1989 gnd.n1635 99.6594
R15997 gnd.n1987 gnd.n1986 99.6594
R15998 gnd.n1985 gnd.n1625 99.6594
R15999 gnd.n1984 gnd.n1621 99.6594
R16000 gnd.n1982 gnd.n1619 99.6594
R16001 gnd.n1981 gnd.n1616 99.6594
R16002 gnd.n1979 gnd.n1614 99.6594
R16003 gnd.n4180 gnd.n4179 99.6594
R16004 gnd.n2001 gnd.n2000 99.6594
R16005 gnd.n2615 gnd.t309 98.63
R16006 gnd.n4523 gnd.t337 98.63
R16007 gnd.n2622 gnd.t355 98.63
R16008 gnd.n1740 gnd.t334 98.63
R16009 gnd.n1763 gnd.t325 98.63
R16010 gnd.n4403 gnd.t267 98.63
R16011 gnd.n313 gnd.t352 98.63
R16012 gnd.n280 gnd.t274 98.63
R16013 gnd.n7566 gnd.t314 98.63
R16014 gnd.n350 gnd.t301 98.63
R16015 gnd.n1090 gnd.t289 98.63
R16016 gnd.n1112 gnd.t286 98.63
R16017 gnd.n1134 gnd.t271 98.63
R16018 gnd.n2750 gnd.t340 98.63
R16019 gnd.n1409 gnd.t342 98.63
R16020 gnd.n2443 gnd.t282 98.63
R16021 gnd.n2465 gnd.t304 98.63
R16022 gnd.n1668 gnd.t292 98.63
R16023 gnd.n3308 gnd.t322 96.6984
R16024 gnd.n2087 gnd.t278 96.6984
R16025 gnd.n4714 gnd.t243 96.6906
R16026 gnd.n3922 gnd.t327 96.6906
R16027 gnd.n1478 gnd.n1477 81.8399
R16028 gnd.n5690 gnd.t318 74.8376
R16029 gnd.n5124 gnd.t347 74.8376
R16030 gnd.n3309 gnd.t321 72.8438
R16031 gnd.n2088 gnd.t279 72.8438
R16032 gnd.n1479 gnd.n1472 72.8411
R16033 gnd.n1485 gnd.n1470 72.8411
R16034 gnd.n3918 gnd.n3917 72.8411
R16035 gnd.n2616 gnd.t308 72.836
R16036 gnd.n4715 gnd.t242 72.836
R16037 gnd.n3923 gnd.t328 72.836
R16038 gnd.n4524 gnd.t336 72.836
R16039 gnd.n2623 gnd.t356 72.836
R16040 gnd.n1741 gnd.t333 72.836
R16041 gnd.n1764 gnd.t324 72.836
R16042 gnd.n4404 gnd.t266 72.836
R16043 gnd.n314 gnd.t353 72.836
R16044 gnd.n281 gnd.t275 72.836
R16045 gnd.n7567 gnd.t315 72.836
R16046 gnd.n351 gnd.t302 72.836
R16047 gnd.n1091 gnd.t288 72.836
R16048 gnd.n1113 gnd.t285 72.836
R16049 gnd.n1135 gnd.t270 72.836
R16050 gnd.n2751 gnd.t339 72.836
R16051 gnd.n1410 gnd.t343 72.836
R16052 gnd.n2444 gnd.t283 72.836
R16053 gnd.n2466 gnd.t305 72.836
R16054 gnd.n1669 gnd.t293 72.836
R16055 gnd.n3986 gnd.n2051 71.676
R16056 gnd.n3982 gnd.n2052 71.676
R16057 gnd.n3978 gnd.n2053 71.676
R16058 gnd.n3974 gnd.n2054 71.676
R16059 gnd.n3970 gnd.n2055 71.676
R16060 gnd.n3966 gnd.n2056 71.676
R16061 gnd.n3962 gnd.n2057 71.676
R16062 gnd.n3958 gnd.n2058 71.676
R16063 gnd.n3954 gnd.n2059 71.676
R16064 gnd.n3950 gnd.n2060 71.676
R16065 gnd.n3946 gnd.n2061 71.676
R16066 gnd.n3942 gnd.n2062 71.676
R16067 gnd.n3938 gnd.n2063 71.676
R16068 gnd.n3934 gnd.n2064 71.676
R16069 gnd.n3929 gnd.n2065 71.676
R16070 gnd.n3925 gnd.n2066 71.676
R16071 gnd.n4059 gnd.n2086 71.676
R16072 gnd.n4055 gnd.n2085 71.676
R16073 gnd.n4050 gnd.n2084 71.676
R16074 gnd.n4046 gnd.n2083 71.676
R16075 gnd.n4042 gnd.n2082 71.676
R16076 gnd.n4038 gnd.n2081 71.676
R16077 gnd.n4034 gnd.n2080 71.676
R16078 gnd.n4030 gnd.n2079 71.676
R16079 gnd.n4026 gnd.n2078 71.676
R16080 gnd.n4022 gnd.n2077 71.676
R16081 gnd.n4018 gnd.n2076 71.676
R16082 gnd.n4014 gnd.n2075 71.676
R16083 gnd.n4010 gnd.n2074 71.676
R16084 gnd.n4006 gnd.n2073 71.676
R16085 gnd.n4002 gnd.n2072 71.676
R16086 gnd.n3998 gnd.n2071 71.676
R16087 gnd.n3994 gnd.n2070 71.676
R16088 gnd.n4778 gnd.n4777 71.676
R16089 gnd.n4772 gnd.n1434 71.676
R16090 gnd.n4769 gnd.n1435 71.676
R16091 gnd.n4765 gnd.n1436 71.676
R16092 gnd.n4761 gnd.n1437 71.676
R16093 gnd.n4757 gnd.n1438 71.676
R16094 gnd.n4753 gnd.n1439 71.676
R16095 gnd.n4749 gnd.n1440 71.676
R16096 gnd.n4745 gnd.n1441 71.676
R16097 gnd.n4741 gnd.n1442 71.676
R16098 gnd.n4737 gnd.n1443 71.676
R16099 gnd.n4733 gnd.n1444 71.676
R16100 gnd.n4729 gnd.n1445 71.676
R16101 gnd.n4725 gnd.n1446 71.676
R16102 gnd.n4721 gnd.n1447 71.676
R16103 gnd.n4717 gnd.n1448 71.676
R16104 gnd.n1449 gnd.n1432 71.676
R16105 gnd.n3312 gnd.n1450 71.676
R16106 gnd.n3317 gnd.n1451 71.676
R16107 gnd.n3321 gnd.n1452 71.676
R16108 gnd.n3325 gnd.n1453 71.676
R16109 gnd.n3329 gnd.n1454 71.676
R16110 gnd.n3333 gnd.n1455 71.676
R16111 gnd.n3337 gnd.n1456 71.676
R16112 gnd.n3341 gnd.n1457 71.676
R16113 gnd.n3345 gnd.n1458 71.676
R16114 gnd.n3349 gnd.n1459 71.676
R16115 gnd.n3353 gnd.n1460 71.676
R16116 gnd.n3357 gnd.n1461 71.676
R16117 gnd.n3361 gnd.n1462 71.676
R16118 gnd.n3365 gnd.n1463 71.676
R16119 gnd.n3369 gnd.n1464 71.676
R16120 gnd.n4778 gnd.n1467 71.676
R16121 gnd.n4770 gnd.n1434 71.676
R16122 gnd.n4766 gnd.n1435 71.676
R16123 gnd.n4762 gnd.n1436 71.676
R16124 gnd.n4758 gnd.n1437 71.676
R16125 gnd.n4754 gnd.n1438 71.676
R16126 gnd.n4750 gnd.n1439 71.676
R16127 gnd.n4746 gnd.n1440 71.676
R16128 gnd.n4742 gnd.n1441 71.676
R16129 gnd.n4738 gnd.n1442 71.676
R16130 gnd.n4734 gnd.n1443 71.676
R16131 gnd.n4730 gnd.n1444 71.676
R16132 gnd.n4726 gnd.n1445 71.676
R16133 gnd.n4722 gnd.n1446 71.676
R16134 gnd.n4718 gnd.n1447 71.676
R16135 gnd.n4781 gnd.n4780 71.676
R16136 gnd.n3311 gnd.n1449 71.676
R16137 gnd.n3316 gnd.n1450 71.676
R16138 gnd.n3320 gnd.n1451 71.676
R16139 gnd.n3324 gnd.n1452 71.676
R16140 gnd.n3328 gnd.n1453 71.676
R16141 gnd.n3332 gnd.n1454 71.676
R16142 gnd.n3336 gnd.n1455 71.676
R16143 gnd.n3340 gnd.n1456 71.676
R16144 gnd.n3344 gnd.n1457 71.676
R16145 gnd.n3348 gnd.n1458 71.676
R16146 gnd.n3352 gnd.n1459 71.676
R16147 gnd.n3356 gnd.n1460 71.676
R16148 gnd.n3360 gnd.n1461 71.676
R16149 gnd.n3364 gnd.n1462 71.676
R16150 gnd.n3368 gnd.n1463 71.676
R16151 gnd.n3307 gnd.n1464 71.676
R16152 gnd.n3997 gnd.n2070 71.676
R16153 gnd.n4001 gnd.n2071 71.676
R16154 gnd.n4005 gnd.n2072 71.676
R16155 gnd.n4009 gnd.n2073 71.676
R16156 gnd.n4013 gnd.n2074 71.676
R16157 gnd.n4017 gnd.n2075 71.676
R16158 gnd.n4021 gnd.n2076 71.676
R16159 gnd.n4025 gnd.n2077 71.676
R16160 gnd.n4029 gnd.n2078 71.676
R16161 gnd.n4033 gnd.n2079 71.676
R16162 gnd.n4037 gnd.n2080 71.676
R16163 gnd.n4041 gnd.n2081 71.676
R16164 gnd.n4045 gnd.n2082 71.676
R16165 gnd.n4049 gnd.n2083 71.676
R16166 gnd.n4054 gnd.n2084 71.676
R16167 gnd.n4058 gnd.n2085 71.676
R16168 gnd.n3924 gnd.n2067 71.676
R16169 gnd.n3928 gnd.n2066 71.676
R16170 gnd.n3933 gnd.n2065 71.676
R16171 gnd.n3937 gnd.n2064 71.676
R16172 gnd.n3941 gnd.n2063 71.676
R16173 gnd.n3945 gnd.n2062 71.676
R16174 gnd.n3949 gnd.n2061 71.676
R16175 gnd.n3953 gnd.n2060 71.676
R16176 gnd.n3957 gnd.n2059 71.676
R16177 gnd.n3961 gnd.n2058 71.676
R16178 gnd.n3965 gnd.n2057 71.676
R16179 gnd.n3969 gnd.n2056 71.676
R16180 gnd.n3973 gnd.n2055 71.676
R16181 gnd.n3977 gnd.n2054 71.676
R16182 gnd.n3981 gnd.n2053 71.676
R16183 gnd.n3985 gnd.n2052 71.676
R16184 gnd.n2093 gnd.n2051 71.676
R16185 gnd.n8 gnd.t68 69.1507
R16186 gnd.n14 gnd.t235 68.4792
R16187 gnd.n13 gnd.t13 68.4792
R16188 gnd.n12 gnd.t11 68.4792
R16189 gnd.n11 gnd.t49 68.4792
R16190 gnd.n10 gnd.t44 68.4792
R16191 gnd.n9 gnd.t56 68.4792
R16192 gnd.n8 gnd.t232 68.4792
R16193 gnd.n5602 gnd.n5503 64.369
R16194 gnd.n3314 gnd.n3309 59.5399
R16195 gnd.n4052 gnd.n2088 59.5399
R16196 gnd.n4716 gnd.n4715 59.5399
R16197 gnd.n3931 gnd.n3923 59.5399
R16198 gnd.n4713 gnd.n1488 59.1804
R16199 gnd.n6473 gnd.n5093 57.3586
R16200 gnd.n5092 gnd.n1068 57.3586
R16201 gnd.n7603 gnd.n212 57.3586
R16202 gnd.n5309 gnd.t147 56.407
R16203 gnd.n5262 gnd.t210 56.407
R16204 gnd.n5277 gnd.t91 56.407
R16205 gnd.n5293 gnd.t199 56.407
R16206 gnd.n64 gnd.t112 56.407
R16207 gnd.n17 gnd.t100 56.407
R16208 gnd.n32 gnd.t222 56.407
R16209 gnd.n48 gnd.t162 56.407
R16210 gnd.n5322 gnd.t132 55.8337
R16211 gnd.n5275 gnd.t218 55.8337
R16212 gnd.n5290 gnd.t191 55.8337
R16213 gnd.n5306 gnd.t178 55.8337
R16214 gnd.n77 gnd.t72 55.8337
R16215 gnd.n30 gnd.t115 55.8337
R16216 gnd.n45 gnd.t173 55.8337
R16217 gnd.n61 gnd.t139 55.8337
R16218 gnd.n1476 gnd.n1475 54.358
R16219 gnd.n3915 gnd.n3914 54.358
R16220 gnd.n5309 gnd.n5308 53.0052
R16221 gnd.n5311 gnd.n5310 53.0052
R16222 gnd.n5313 gnd.n5312 53.0052
R16223 gnd.n5315 gnd.n5314 53.0052
R16224 gnd.n5317 gnd.n5316 53.0052
R16225 gnd.n5319 gnd.n5318 53.0052
R16226 gnd.n5321 gnd.n5320 53.0052
R16227 gnd.n5262 gnd.n5261 53.0052
R16228 gnd.n5264 gnd.n5263 53.0052
R16229 gnd.n5266 gnd.n5265 53.0052
R16230 gnd.n5268 gnd.n5267 53.0052
R16231 gnd.n5270 gnd.n5269 53.0052
R16232 gnd.n5272 gnd.n5271 53.0052
R16233 gnd.n5274 gnd.n5273 53.0052
R16234 gnd.n5277 gnd.n5276 53.0052
R16235 gnd.n5279 gnd.n5278 53.0052
R16236 gnd.n5281 gnd.n5280 53.0052
R16237 gnd.n5283 gnd.n5282 53.0052
R16238 gnd.n5285 gnd.n5284 53.0052
R16239 gnd.n5287 gnd.n5286 53.0052
R16240 gnd.n5289 gnd.n5288 53.0052
R16241 gnd.n5293 gnd.n5292 53.0052
R16242 gnd.n5295 gnd.n5294 53.0052
R16243 gnd.n5297 gnd.n5296 53.0052
R16244 gnd.n5299 gnd.n5298 53.0052
R16245 gnd.n5301 gnd.n5300 53.0052
R16246 gnd.n5303 gnd.n5302 53.0052
R16247 gnd.n5305 gnd.n5304 53.0052
R16248 gnd.n76 gnd.n75 53.0052
R16249 gnd.n74 gnd.n73 53.0052
R16250 gnd.n72 gnd.n71 53.0052
R16251 gnd.n70 gnd.n69 53.0052
R16252 gnd.n68 gnd.n67 53.0052
R16253 gnd.n66 gnd.n65 53.0052
R16254 gnd.n64 gnd.n63 53.0052
R16255 gnd.n29 gnd.n28 53.0052
R16256 gnd.n27 gnd.n26 53.0052
R16257 gnd.n25 gnd.n24 53.0052
R16258 gnd.n23 gnd.n22 53.0052
R16259 gnd.n21 gnd.n20 53.0052
R16260 gnd.n19 gnd.n18 53.0052
R16261 gnd.n17 gnd.n16 53.0052
R16262 gnd.n44 gnd.n43 53.0052
R16263 gnd.n42 gnd.n41 53.0052
R16264 gnd.n40 gnd.n39 53.0052
R16265 gnd.n38 gnd.n37 53.0052
R16266 gnd.n36 gnd.n35 53.0052
R16267 gnd.n34 gnd.n33 53.0052
R16268 gnd.n32 gnd.n31 53.0052
R16269 gnd.n60 gnd.n59 53.0052
R16270 gnd.n58 gnd.n57 53.0052
R16271 gnd.n56 gnd.n55 53.0052
R16272 gnd.n54 gnd.n53 53.0052
R16273 gnd.n52 gnd.n51 53.0052
R16274 gnd.n50 gnd.n49 53.0052
R16275 gnd.n48 gnd.n47 53.0052
R16276 gnd.n3906 gnd.n3905 52.4801
R16277 gnd.n6318 gnd.t58 52.3082
R16278 gnd.n6286 gnd.t64 52.3082
R16279 gnd.n6254 gnd.t18 52.3082
R16280 gnd.n6223 gnd.t237 52.3082
R16281 gnd.n6191 gnd.t51 52.3082
R16282 gnd.n6159 gnd.t239 52.3082
R16283 gnd.n6127 gnd.t16 52.3082
R16284 gnd.n6096 gnd.t53 52.3082
R16285 gnd.n6148 gnd.n6116 51.4173
R16286 gnd.n6212 gnd.n6211 50.455
R16287 gnd.n6180 gnd.n6179 50.455
R16288 gnd.n6148 gnd.n6147 50.455
R16289 gnd.n5540 gnd.n5539 45.1884
R16290 gnd.n5168 gnd.n5167 45.1884
R16291 gnd.n3989 gnd.n3921 44.3322
R16292 gnd.n1479 gnd.n1478 44.3189
R16293 gnd.n2617 gnd.n2616 42.2793
R16294 gnd.n4525 gnd.n4524 42.2793
R16295 gnd.n5552 gnd.n5540 42.2793
R16296 gnd.n5169 gnd.n5168 42.2793
R16297 gnd.n5692 gnd.n5690 42.2793
R16298 gnd.n5125 gnd.n5124 42.2793
R16299 gnd.n3163 gnd.n2623 42.2793
R16300 gnd.n4484 gnd.n1741 42.2793
R16301 gnd.n4447 gnd.n1764 42.2793
R16302 gnd.n4407 gnd.n4404 42.2793
R16303 gnd.n315 gnd.n314 42.2793
R16304 gnd.n7531 gnd.n281 42.2793
R16305 gnd.n7568 gnd.n7567 42.2793
R16306 gnd.n7459 gnd.n351 42.2793
R16307 gnd.n5056 gnd.n1091 42.2793
R16308 gnd.n5016 gnd.n1113 42.2793
R16309 gnd.n4976 gnd.n1135 42.2793
R16310 gnd.n2803 gnd.n2751 42.2793
R16311 gnd.n4798 gnd.n1410 42.2793
R16312 gnd.n2445 gnd.n2444 42.2793
R16313 gnd.n2467 gnd.n2466 42.2793
R16314 gnd.n1670 gnd.n1669 42.2793
R16315 gnd.n1477 gnd.n1476 41.6274
R16316 gnd.n3916 gnd.n3915 41.6274
R16317 gnd.n1486 gnd.n1485 40.8975
R16318 gnd.n3919 gnd.n3918 40.8975
R16319 gnd.n6677 gnd.n801 39.6473
R16320 gnd.n6671 gnd.n801 39.6473
R16321 gnd.n6671 gnd.n6670 39.6473
R16322 gnd.n6670 gnd.n6669 39.6473
R16323 gnd.n6669 gnd.n808 39.6473
R16324 gnd.n6663 gnd.n808 39.6473
R16325 gnd.n6663 gnd.n6662 39.6473
R16326 gnd.n6662 gnd.n6661 39.6473
R16327 gnd.n6661 gnd.n816 39.6473
R16328 gnd.n6655 gnd.n816 39.6473
R16329 gnd.n6655 gnd.n6654 39.6473
R16330 gnd.n6654 gnd.n6653 39.6473
R16331 gnd.n6653 gnd.n824 39.6473
R16332 gnd.n6647 gnd.n824 39.6473
R16333 gnd.n6647 gnd.n6646 39.6473
R16334 gnd.n6646 gnd.n6645 39.6473
R16335 gnd.n6645 gnd.n832 39.6473
R16336 gnd.n6639 gnd.n832 39.6473
R16337 gnd.n6639 gnd.n6638 39.6473
R16338 gnd.n6638 gnd.n6637 39.6473
R16339 gnd.n6637 gnd.n840 39.6473
R16340 gnd.n6631 gnd.n840 39.6473
R16341 gnd.n6631 gnd.n6630 39.6473
R16342 gnd.n6630 gnd.n6629 39.6473
R16343 gnd.n6629 gnd.n848 39.6473
R16344 gnd.n6623 gnd.n848 39.6473
R16345 gnd.n6623 gnd.n6622 39.6473
R16346 gnd.n6622 gnd.n6621 39.6473
R16347 gnd.n6621 gnd.n856 39.6473
R16348 gnd.n6615 gnd.n856 39.6473
R16349 gnd.n6615 gnd.n6614 39.6473
R16350 gnd.n6614 gnd.n6613 39.6473
R16351 gnd.n6613 gnd.n864 39.6473
R16352 gnd.n6607 gnd.n864 39.6473
R16353 gnd.n6607 gnd.n6606 39.6473
R16354 gnd.n6606 gnd.n6605 39.6473
R16355 gnd.n6605 gnd.n872 39.6473
R16356 gnd.n6599 gnd.n872 39.6473
R16357 gnd.n6599 gnd.n6598 39.6473
R16358 gnd.n6598 gnd.n6597 39.6473
R16359 gnd.n6597 gnd.n880 39.6473
R16360 gnd.n6591 gnd.n880 39.6473
R16361 gnd.n6591 gnd.n6590 39.6473
R16362 gnd.n6590 gnd.n6589 39.6473
R16363 gnd.n6589 gnd.n888 39.6473
R16364 gnd.n6583 gnd.n888 39.6473
R16365 gnd.n6583 gnd.n6582 39.6473
R16366 gnd.n6582 gnd.n6581 39.6473
R16367 gnd.n6581 gnd.n896 39.6473
R16368 gnd.n6575 gnd.n896 39.6473
R16369 gnd.n6575 gnd.n6574 39.6473
R16370 gnd.n6574 gnd.n6573 39.6473
R16371 gnd.n6573 gnd.n904 39.6473
R16372 gnd.n6567 gnd.n904 39.6473
R16373 gnd.n6567 gnd.n6566 39.6473
R16374 gnd.n6566 gnd.n6565 39.6473
R16375 gnd.n6565 gnd.n912 39.6473
R16376 gnd.n6559 gnd.n912 39.6473
R16377 gnd.n6559 gnd.n6558 39.6473
R16378 gnd.n6558 gnd.n6557 39.6473
R16379 gnd.n6557 gnd.n920 39.6473
R16380 gnd.n6551 gnd.n920 39.6473
R16381 gnd.n6551 gnd.n6550 39.6473
R16382 gnd.n6550 gnd.n6549 39.6473
R16383 gnd.n6549 gnd.n928 39.6473
R16384 gnd.n6543 gnd.n928 39.6473
R16385 gnd.n6543 gnd.n6542 39.6473
R16386 gnd.n6542 gnd.n6541 39.6473
R16387 gnd.n6541 gnd.n936 39.6473
R16388 gnd.n6535 gnd.n936 39.6473
R16389 gnd.n6535 gnd.n6534 39.6473
R16390 gnd.n6534 gnd.n6533 39.6473
R16391 gnd.n6533 gnd.n944 39.6473
R16392 gnd.n6527 gnd.n944 39.6473
R16393 gnd.n6527 gnd.n6526 39.6473
R16394 gnd.n6526 gnd.n6525 39.6473
R16395 gnd.n6525 gnd.n952 39.6473
R16396 gnd.n6519 gnd.n952 39.6473
R16397 gnd.n6519 gnd.n6518 39.6473
R16398 gnd.n6518 gnd.n6517 39.6473
R16399 gnd.n6517 gnd.n960 39.6473
R16400 gnd.n6511 gnd.n960 39.6473
R16401 gnd.n6511 gnd.n6510 39.6473
R16402 gnd.n1485 gnd.n1484 35.055
R16403 gnd.n1480 gnd.n1479 35.055
R16404 gnd.n3908 gnd.n3907 35.055
R16405 gnd.n3918 gnd.n3904 35.055
R16406 gnd.n3995 gnd.n2089 33.2493
R16407 gnd.n3412 gnd.n3371 33.2493
R16408 gnd.n5602 gnd.n5498 31.8661
R16409 gnd.n5610 gnd.n5498 31.8661
R16410 gnd.n5618 gnd.n5492 31.8661
R16411 gnd.n5618 gnd.n5486 31.8661
R16412 gnd.n5626 gnd.n5486 31.8661
R16413 gnd.n5626 gnd.n5479 31.8661
R16414 gnd.n5634 gnd.n5479 31.8661
R16415 gnd.n5634 gnd.n5480 31.8661
R16416 gnd.n5733 gnd.n5465 31.8661
R16417 gnd.n4968 gnd.n1068 31.8661
R16418 gnd.n4962 gnd.n1152 31.8661
R16419 gnd.n4962 gnd.n1155 31.8661
R16420 gnd.n4956 gnd.n1155 31.8661
R16421 gnd.n4956 gnd.n1167 31.8661
R16422 gnd.n4950 gnd.n1177 31.8661
R16423 gnd.n3106 gnd.n1376 31.8661
R16424 gnd.n3101 gnd.n3100 31.8661
R16425 gnd.n3101 gnd.n2419 31.8661
R16426 gnd.n3088 gnd.n2433 31.8661
R16427 gnd.n4125 gnd.n1978 31.8661
R16428 gnd.n4177 gnd.n2002 31.8661
R16429 gnd.n2002 gnd.n1676 31.8661
R16430 gnd.n1786 gnd.n1718 31.8661
R16431 gnd.n7627 gnd.n175 31.8661
R16432 gnd.n7621 gnd.n185 31.8661
R16433 gnd.n7615 gnd.n185 31.8661
R16434 gnd.n7615 gnd.n194 31.8661
R16435 gnd.n7609 gnd.n194 31.8661
R16436 gnd.n7603 gnd.n209 31.8661
R16437 gnd.n4938 gnd.n1194 26.7676
R16438 gnd.n4932 gnd.n1204 26.7676
R16439 gnd.n2890 gnd.n1207 26.7676
R16440 gnd.n2884 gnd.n1217 26.7676
R16441 gnd.n4920 gnd.n1224 26.7676
R16442 gnd.n4914 gnd.n1235 26.7676
R16443 gnd.n4908 gnd.n1245 26.7676
R16444 gnd.n2709 gnd.n1248 26.7676
R16445 gnd.n2934 gnd.n2697 26.7676
R16446 gnd.n2931 gnd.n2699 26.7676
R16447 gnd.n2961 gnd.n2679 26.7676
R16448 gnd.n2968 gnd.n2967 26.7676
R16449 gnd.n2996 gnd.n2667 26.7676
R16450 gnd.n3004 gnd.n1265 26.7676
R16451 gnd.n4894 gnd.n1274 26.7676
R16452 gnd.n3011 gnd.n2661 26.7676
R16453 gnd.n4888 gnd.n1283 26.7676
R16454 gnd.n4882 gnd.n1293 26.7676
R16455 gnd.n3055 gnd.n1296 26.7676
R16456 gnd.n3026 gnd.n1306 26.7676
R16457 gnd.n4870 gnd.n1313 26.7676
R16458 gnd.n3032 gnd.n3031 26.7676
R16459 gnd.n4864 gnd.n1323 26.7676
R16460 gnd.n4858 gnd.n1333 26.7676
R16461 gnd.n3121 gnd.n1336 26.7676
R16462 gnd.n3127 gnd.n1346 26.7676
R16463 gnd.n4846 gnd.n1353 26.7676
R16464 gnd.n3136 gnd.n1356 26.7676
R16465 gnd.n4840 gnd.n1364 26.7676
R16466 gnd.n4834 gnd.n1373 26.7676
R16467 gnd.n4399 gnd.n1788 26.7676
R16468 gnd.n4391 gnd.n1798 26.7676
R16469 gnd.n4189 gnd.n1811 26.7676
R16470 gnd.n4385 gnd.n1814 26.7676
R16471 gnd.n4197 gnd.n1824 26.7676
R16472 gnd.n4204 gnd.n1834 26.7676
R16473 gnd.n4373 gnd.n1837 26.7676
R16474 gnd.n4367 gnd.n1847 26.7676
R16475 gnd.n4249 gnd.n4248 26.7676
R16476 gnd.n4361 gnd.n1857 26.7676
R16477 gnd.n4219 gnd.n1864 26.7676
R16478 gnd.n4225 gnd.n1874 26.7676
R16479 gnd.n4349 gnd.n1877 26.7676
R16480 gnd.n4343 gnd.n1887 26.7676
R16481 gnd.n4273 gnd.n4272 26.7676
R16482 gnd.n4337 gnd.n1897 26.7676
R16483 gnd.n4289 gnd.n1904 26.7676
R16484 gnd.n4327 gnd.n4326 26.7676
R16485 gnd.n1927 gnd.n1912 26.7676
R16486 gnd.n4318 gnd.n1924 26.7676
R16487 gnd.n7677 gnd.n87 26.7676
R16488 gnd.n7369 gnd.n381 26.7676
R16489 gnd.n7669 gnd.n105 26.7676
R16490 gnd.n7380 gnd.n114 26.7676
R16491 gnd.n7388 gnd.n123 26.7676
R16492 gnd.n7394 gnd.n132 26.7676
R16493 gnd.n7651 gnd.n135 26.7676
R16494 gnd.n7645 gnd.n146 26.7676
R16495 gnd.n7408 gnd.n153 26.7676
R16496 gnd.n7417 gnd.n163 26.7676
R16497 gnd.n2948 gnd.t148 26.4489
R16498 gnd.n4307 gnd.t113 26.4489
R16499 gnd.n2878 gnd.t84 25.8116
R16500 gnd.n7657 gnd.t129 25.8116
R16501 gnd.n2616 gnd.n2615 25.7944
R16502 gnd.n4524 gnd.n4523 25.7944
R16503 gnd.n5690 gnd.n5689 25.7944
R16504 gnd.n5124 gnd.n5123 25.7944
R16505 gnd.n2623 gnd.n2622 25.7944
R16506 gnd.n1741 gnd.n1740 25.7944
R16507 gnd.n1764 gnd.n1763 25.7944
R16508 gnd.n4404 gnd.n4403 25.7944
R16509 gnd.n314 gnd.n313 25.7944
R16510 gnd.n281 gnd.n280 25.7944
R16511 gnd.n7567 gnd.n7566 25.7944
R16512 gnd.n351 gnd.n350 25.7944
R16513 gnd.n1091 gnd.n1090 25.7944
R16514 gnd.n1113 gnd.n1112 25.7944
R16515 gnd.n1135 gnd.n1134 25.7944
R16516 gnd.n2751 gnd.n2750 25.7944
R16517 gnd.n1410 gnd.n1409 25.7944
R16518 gnd.n2444 gnd.n2443 25.7944
R16519 gnd.n2466 gnd.n2465 25.7944
R16520 gnd.n1669 gnd.n1668 25.7944
R16521 gnd.n2842 gnd.t102 25.1743
R16522 gnd.n7633 gnd.t73 25.1743
R16523 gnd.n5734 gnd.n5454 24.8557
R16524 gnd.n5457 gnd.n5448 24.8557
R16525 gnd.n5755 gnd.n5433 24.8557
R16526 gnd.n5774 gnd.n5773 24.8557
R16527 gnd.n5784 gnd.n5426 24.8557
R16528 gnd.n5797 gnd.n5414 24.8557
R16529 gnd.n5822 gnd.n5398 24.8557
R16530 gnd.n5821 gnd.n5400 24.8557
R16531 gnd.n5844 gnd.n5382 24.8557
R16532 gnd.n5833 gnd.n5374 24.8557
R16533 gnd.n5869 gnd.n5868 24.8557
R16534 gnd.n5879 gnd.n5367 24.8557
R16535 gnd.n5891 gnd.n5359 24.8557
R16536 gnd.n5890 gnd.n5347 24.8557
R16537 gnd.n5909 gnd.n5908 24.8557
R16538 gnd.n5930 gnd.n5328 24.8557
R16539 gnd.n5954 gnd.n5953 24.8557
R16540 gnd.n5965 gnd.n5247 24.8557
R16541 gnd.n5964 gnd.n5249 24.8557
R16542 gnd.n5976 gnd.n5240 24.8557
R16543 gnd.n5993 gnd.n5992 24.8557
R16544 gnd.n5231 gnd.n5220 24.8557
R16545 gnd.n6016 gnd.n5210 24.8557
R16546 gnd.n5212 gnd.n5211 24.8557
R16547 gnd.n6039 gnd.n5204 24.8557
R16548 gnd.n6050 gnd.n6049 24.8557
R16549 gnd.n6064 gnd.n5191 24.8557
R16550 gnd.n6502 gnd.n979 24.8557
R16551 gnd.n6365 gnd.n990 24.8557
R16552 gnd.n6495 gnd.n6494 24.8557
R16553 gnd.n6488 gnd.n1002 24.8557
R16554 gnd.n6487 gnd.n1005 24.8557
R16555 gnd.n6354 gnd.n1016 24.8557
R16556 gnd.n6474 gnd.n1027 24.8557
R16557 gnd.n3309 gnd.n3308 23.855
R16558 gnd.n2088 gnd.n2087 23.855
R16559 gnd.n4715 gnd.n4714 23.855
R16560 gnd.n3923 gnd.n3922 23.855
R16561 gnd.n6510 gnd.n6509 23.7886
R16562 gnd.n5752 gnd.t52 23.2624
R16563 gnd.n5744 gnd.t317 22.6251
R16564 gnd.n4968 gnd.t269 22.6251
R16565 gnd.t154 gnd.n1197 22.6251
R16566 gnd.n3143 gnd.t281 22.6251
R16567 gnd.n1970 gnd.t265 22.6251
R16568 gnd.n362 gnd.t121 22.6251
R16569 gnd.n209 gnd.t273 22.6251
R16570 gnd.t134 gnd.n1238 21.9878
R16571 gnd.n374 gnd.t79 21.9878
R16572 gnd.n5724 gnd.t236 21.3504
R16573 gnd.n2682 gnd.t107 21.3504
R16574 gnd.n4319 gnd.t75 21.3504
R16575 gnd.n4713 gnd.n4712 21.0737
R16576 gnd.n3990 gnd.n3989 21.0737
R16577 gnd.n6029 gnd.t29 20.7131
R16578 gnd.t97 gnd.n1286 20.7131
R16579 gnd.t77 gnd.n1884 20.7131
R16580 gnd.n3106 gnd.n1381 20.3945
R16581 gnd.n4520 gnd.n1718 20.3945
R16582 gnd.t31 gnd.n5221 20.0758
R16583 gnd.t104 gnd.n1326 20.0758
R16584 gnd.t69 gnd.n1844 20.0758
R16585 gnd.n1474 gnd.t312 19.8005
R16586 gnd.n1474 gnd.t246 19.8005
R16587 gnd.n1473 gnd.t299 19.8005
R16588 gnd.n1473 gnd.t350 19.8005
R16589 gnd.n3913 gnd.t359 19.8005
R16590 gnd.n3913 gnd.t249 19.8005
R16591 gnd.n3912 gnd.t260 19.8005
R16592 gnd.n3912 gnd.t331 19.8005
R16593 gnd.n1470 gnd.n1469 19.5087
R16594 gnd.n1483 gnd.n1470 19.5087
R16595 gnd.n1481 gnd.n1472 19.5087
R16596 gnd.n3917 gnd.n3911 19.5087
R16597 gnd.t37 gnd.n5256 19.4385
R16598 gnd.n3233 gnd.n2408 19.3944
R16599 gnd.n3233 gnd.n2405 19.3944
R16600 gnd.n3238 gnd.n2405 19.3944
R16601 gnd.n3238 gnd.n2406 19.3944
R16602 gnd.n2406 gnd.n2383 19.3944
R16603 gnd.n3263 gnd.n2383 19.3944
R16604 gnd.n3263 gnd.n2380 19.3944
R16605 gnd.n3268 gnd.n2380 19.3944
R16606 gnd.n3268 gnd.n2381 19.3944
R16607 gnd.n2381 gnd.n2359 19.3944
R16608 gnd.n3300 gnd.n2359 19.3944
R16609 gnd.n3300 gnd.n2356 19.3944
R16610 gnd.n3305 gnd.n2356 19.3944
R16611 gnd.n3305 gnd.n2357 19.3944
R16612 gnd.n2357 gnd.n2346 19.3944
R16613 gnd.n3427 gnd.n2346 19.3944
R16614 gnd.n3427 gnd.n2343 19.3944
R16615 gnd.n3433 gnd.n2343 19.3944
R16616 gnd.n3433 gnd.n2344 19.3944
R16617 gnd.n2344 gnd.n2332 19.3944
R16618 gnd.n2332 gnd.n2330 19.3944
R16619 gnd.n3455 gnd.n2330 19.3944
R16620 gnd.n3455 gnd.n2327 19.3944
R16621 gnd.n3460 gnd.n2327 19.3944
R16622 gnd.n3460 gnd.n2328 19.3944
R16623 gnd.n2328 gnd.n2311 19.3944
R16624 gnd.n3510 gnd.n2311 19.3944
R16625 gnd.n3510 gnd.n2308 19.3944
R16626 gnd.n3516 gnd.n2308 19.3944
R16627 gnd.n3516 gnd.n2309 19.3944
R16628 gnd.n2309 gnd.n2297 19.3944
R16629 gnd.n2297 gnd.n2295 19.3944
R16630 gnd.n3540 gnd.n2295 19.3944
R16631 gnd.n3540 gnd.n2293 19.3944
R16632 gnd.n3544 gnd.n2293 19.3944
R16633 gnd.n3544 gnd.n2266 19.3944
R16634 gnd.n3590 gnd.n2266 19.3944
R16635 gnd.n3590 gnd.n2267 19.3944
R16636 gnd.n3586 gnd.n2267 19.3944
R16637 gnd.n3586 gnd.n2242 19.3944
R16638 gnd.n3645 gnd.n2242 19.3944
R16639 gnd.n3645 gnd.n2243 19.3944
R16640 gnd.n3641 gnd.n2243 19.3944
R16641 gnd.n3641 gnd.n3640 19.3944
R16642 gnd.n3640 gnd.n3639 19.3944
R16643 gnd.n3639 gnd.n3628 19.3944
R16644 gnd.n3635 gnd.n3628 19.3944
R16645 gnd.n3635 gnd.n3634 19.3944
R16646 gnd.n3634 gnd.n3633 19.3944
R16647 gnd.n3633 gnd.n2181 19.3944
R16648 gnd.n3760 gnd.n2181 19.3944
R16649 gnd.n3760 gnd.n2179 19.3944
R16650 gnd.n3764 gnd.n2179 19.3944
R16651 gnd.n3764 gnd.n2160 19.3944
R16652 gnd.n3790 gnd.n2160 19.3944
R16653 gnd.n3790 gnd.n2157 19.3944
R16654 gnd.n3798 gnd.n2157 19.3944
R16655 gnd.n3798 gnd.n2158 19.3944
R16656 gnd.n3794 gnd.n2158 19.3944
R16657 gnd.n3794 gnd.n2131 19.3944
R16658 gnd.n3829 gnd.n2131 19.3944
R16659 gnd.n3829 gnd.n2128 19.3944
R16660 gnd.n3849 gnd.n2128 19.3944
R16661 gnd.n3849 gnd.n2129 19.3944
R16662 gnd.n3845 gnd.n2129 19.3944
R16663 gnd.n3845 gnd.n3844 19.3944
R16664 gnd.n3844 gnd.n3843 19.3944
R16665 gnd.n3843 gnd.n3835 19.3944
R16666 gnd.n3839 gnd.n3835 19.3944
R16667 gnd.n3839 gnd.n2041 19.3944
R16668 gnd.n4072 gnd.n2041 19.3944
R16669 gnd.n4072 gnd.n2039 19.3944
R16670 gnd.n4076 gnd.n2039 19.3944
R16671 gnd.n4076 gnd.n2028 19.3944
R16672 gnd.n4092 gnd.n2028 19.3944
R16673 gnd.n4092 gnd.n2026 19.3944
R16674 gnd.n4096 gnd.n2026 19.3944
R16675 gnd.n4096 gnd.n2014 19.3944
R16676 gnd.n4114 gnd.n2014 19.3944
R16677 gnd.n4114 gnd.n2011 19.3944
R16678 gnd.n4119 gnd.n2011 19.3944
R16679 gnd.n4119 gnd.n2012 19.3944
R16680 gnd.n3151 gnd.n3150 19.3944
R16681 gnd.n3157 gnd.n3151 19.3944
R16682 gnd.n3157 gnd.n3156 19.3944
R16683 gnd.n3224 gnd.n2417 19.3944
R16684 gnd.n3219 gnd.n2417 19.3944
R16685 gnd.n3219 gnd.n2435 19.3944
R16686 gnd.n3215 gnd.n2435 19.3944
R16687 gnd.n3215 gnd.n3214 19.3944
R16688 gnd.n3214 gnd.n3213 19.3944
R16689 gnd.n3213 gnd.n2441 19.3944
R16690 gnd.n3208 gnd.n2441 19.3944
R16691 gnd.n3208 gnd.n3207 19.3944
R16692 gnd.n3207 gnd.n2558 19.3944
R16693 gnd.n3200 gnd.n2558 19.3944
R16694 gnd.n3200 gnd.n3199 19.3944
R16695 gnd.n3199 gnd.n2570 19.3944
R16696 gnd.n3192 gnd.n2570 19.3944
R16697 gnd.n3192 gnd.n3191 19.3944
R16698 gnd.n3191 gnd.n2580 19.3944
R16699 gnd.n3184 gnd.n2580 19.3944
R16700 gnd.n3184 gnd.n3183 19.3944
R16701 gnd.n3183 gnd.n2593 19.3944
R16702 gnd.n3176 gnd.n2593 19.3944
R16703 gnd.n3176 gnd.n3175 19.3944
R16704 gnd.n3175 gnd.n2603 19.3944
R16705 gnd.n3168 gnd.n2603 19.3944
R16706 gnd.n3168 gnd.n3167 19.3944
R16707 gnd.n4566 gnd.n1629 19.3944
R16708 gnd.n4566 gnd.n4565 19.3944
R16709 gnd.n4565 gnd.n1632 19.3944
R16710 gnd.n4558 gnd.n1632 19.3944
R16711 gnd.n4558 gnd.n4557 19.3944
R16712 gnd.n4557 gnd.n1640 19.3944
R16713 gnd.n4550 gnd.n1640 19.3944
R16714 gnd.n4550 gnd.n4549 19.3944
R16715 gnd.n4549 gnd.n1648 19.3944
R16716 gnd.n4542 gnd.n1648 19.3944
R16717 gnd.n4542 gnd.n4541 19.3944
R16718 gnd.n4541 gnd.n1656 19.3944
R16719 gnd.n4534 gnd.n1656 19.3944
R16720 gnd.n4534 gnd.n4533 19.3944
R16721 gnd.n4533 gnd.n1664 19.3944
R16722 gnd.n4526 gnd.n1664 19.3944
R16723 gnd.n5597 gnd.n5596 19.3944
R16724 gnd.n5596 gnd.n5506 19.3944
R16725 gnd.n5591 gnd.n5506 19.3944
R16726 gnd.n5591 gnd.n5590 19.3944
R16727 gnd.n5590 gnd.n5511 19.3944
R16728 gnd.n5585 gnd.n5511 19.3944
R16729 gnd.n5585 gnd.n5584 19.3944
R16730 gnd.n5584 gnd.n5583 19.3944
R16731 gnd.n5583 gnd.n5517 19.3944
R16732 gnd.n5577 gnd.n5517 19.3944
R16733 gnd.n5577 gnd.n5576 19.3944
R16734 gnd.n5576 gnd.n5575 19.3944
R16735 gnd.n5575 gnd.n5523 19.3944
R16736 gnd.n5569 gnd.n5523 19.3944
R16737 gnd.n5569 gnd.n5568 19.3944
R16738 gnd.n5568 gnd.n5567 19.3944
R16739 gnd.n5567 gnd.n5529 19.3944
R16740 gnd.n5561 gnd.n5529 19.3944
R16741 gnd.n5561 gnd.n5560 19.3944
R16742 gnd.n5560 gnd.n5559 19.3944
R16743 gnd.n5559 gnd.n5535 19.3944
R16744 gnd.n5553 gnd.n5535 19.3944
R16745 gnd.n5551 gnd.n5550 19.3944
R16746 gnd.n5550 gnd.n5545 19.3944
R16747 gnd.n5545 gnd.n5543 19.3944
R16748 gnd.n6394 gnd.n5171 19.3944
R16749 gnd.n6394 gnd.n6393 19.3944
R16750 gnd.n6393 gnd.n6392 19.3944
R16751 gnd.n6436 gnd.n6435 19.3944
R16752 gnd.n6435 gnd.n6434 19.3944
R16753 gnd.n6434 gnd.n5132 19.3944
R16754 gnd.n6429 gnd.n5132 19.3944
R16755 gnd.n6429 gnd.n6428 19.3944
R16756 gnd.n6428 gnd.n6427 19.3944
R16757 gnd.n6427 gnd.n5139 19.3944
R16758 gnd.n6422 gnd.n5139 19.3944
R16759 gnd.n6422 gnd.n6421 19.3944
R16760 gnd.n6421 gnd.n6420 19.3944
R16761 gnd.n6420 gnd.n5146 19.3944
R16762 gnd.n6415 gnd.n5146 19.3944
R16763 gnd.n6415 gnd.n6414 19.3944
R16764 gnd.n6414 gnd.n6413 19.3944
R16765 gnd.n6413 gnd.n5153 19.3944
R16766 gnd.n6408 gnd.n5153 19.3944
R16767 gnd.n6408 gnd.n6407 19.3944
R16768 gnd.n6407 gnd.n6406 19.3944
R16769 gnd.n6406 gnd.n5160 19.3944
R16770 gnd.n6401 gnd.n5160 19.3944
R16771 gnd.n6401 gnd.n6400 19.3944
R16772 gnd.n6400 gnd.n6399 19.3944
R16773 gnd.n5737 gnd.n5736 19.3944
R16774 gnd.n5738 gnd.n5737 19.3944
R16775 gnd.n5738 gnd.n5447 19.3944
R16776 gnd.n5447 gnd.n5441 19.3944
R16777 gnd.n5763 gnd.n5441 19.3944
R16778 gnd.n5764 gnd.n5763 19.3944
R16779 gnd.n5764 gnd.n5424 19.3944
R16780 gnd.n5424 gnd.n5422 19.3944
R16781 gnd.n5788 gnd.n5422 19.3944
R16782 gnd.n5791 gnd.n5788 19.3944
R16783 gnd.n5791 gnd.n5790 19.3944
R16784 gnd.n5790 gnd.n5394 19.3944
R16785 gnd.n5829 gnd.n5394 19.3944
R16786 gnd.n5829 gnd.n5392 19.3944
R16787 gnd.n5835 gnd.n5392 19.3944
R16788 gnd.n5836 gnd.n5835 19.3944
R16789 gnd.n5836 gnd.n5362 19.3944
R16790 gnd.n5886 gnd.n5362 19.3944
R16791 gnd.n5887 gnd.n5886 19.3944
R16792 gnd.n5887 gnd.n5355 19.3944
R16793 gnd.n5898 gnd.n5355 19.3944
R16794 gnd.n5899 gnd.n5898 19.3944
R16795 gnd.n5899 gnd.n5338 19.3944
R16796 gnd.n5338 gnd.n5336 19.3944
R16797 gnd.n5923 gnd.n5336 19.3944
R16798 gnd.n5924 gnd.n5923 19.3944
R16799 gnd.n5924 gnd.n5243 19.3944
R16800 gnd.n5971 gnd.n5243 19.3944
R16801 gnd.n5972 gnd.n5971 19.3944
R16802 gnd.n5972 gnd.n5236 19.3944
R16803 gnd.n5983 gnd.n5236 19.3944
R16804 gnd.n5984 gnd.n5983 19.3944
R16805 gnd.n5984 gnd.n5219 19.3944
R16806 gnd.n5219 gnd.n5217 19.3944
R16807 gnd.n6011 gnd.n5217 19.3944
R16808 gnd.n6011 gnd.n5200 19.3944
R16809 gnd.n6045 gnd.n5200 19.3944
R16810 gnd.n6046 gnd.n6045 19.3944
R16811 gnd.n6046 gnd.n5186 19.3944
R16812 gnd.n6072 gnd.n5186 19.3944
R16813 gnd.n6072 gnd.n5183 19.3944
R16814 gnd.n6076 gnd.n5183 19.3944
R16815 gnd.n6077 gnd.n6076 19.3944
R16816 gnd.n6363 gnd.n6077 19.3944
R16817 gnd.n6363 gnd.n6362 19.3944
R16818 gnd.n6362 gnd.n6361 19.3944
R16819 gnd.n6361 gnd.n6358 19.3944
R16820 gnd.n6358 gnd.n6357 19.3944
R16821 gnd.n6357 gnd.n6356 19.3944
R16822 gnd.n6356 gnd.n6353 19.3944
R16823 gnd.n6353 gnd.n6352 19.3944
R16824 gnd.n6352 gnd.n6349 19.3944
R16825 gnd.n6349 gnd.n6348 19.3944
R16826 gnd.n5720 gnd.n5719 19.3944
R16827 gnd.n5719 gnd.n5718 19.3944
R16828 gnd.n5718 gnd.n5717 19.3944
R16829 gnd.n5717 gnd.n5715 19.3944
R16830 gnd.n5715 gnd.n5712 19.3944
R16831 gnd.n5712 gnd.n5711 19.3944
R16832 gnd.n5711 gnd.n5708 19.3944
R16833 gnd.n5708 gnd.n5707 19.3944
R16834 gnd.n5707 gnd.n5704 19.3944
R16835 gnd.n5704 gnd.n5703 19.3944
R16836 gnd.n5703 gnd.n5700 19.3944
R16837 gnd.n5700 gnd.n5699 19.3944
R16838 gnd.n5699 gnd.n5696 19.3944
R16839 gnd.n5696 gnd.n5695 19.3944
R16840 gnd.n5746 gnd.n5452 19.3944
R16841 gnd.n5746 gnd.n5450 19.3944
R16842 gnd.n5750 gnd.n5450 19.3944
R16843 gnd.n5750 gnd.n5431 19.3944
R16844 gnd.n5776 gnd.n5431 19.3944
R16845 gnd.n5776 gnd.n5429 19.3944
R16846 gnd.n5782 gnd.n5429 19.3944
R16847 gnd.n5782 gnd.n5781 19.3944
R16848 gnd.n5781 gnd.n5405 19.3944
R16849 gnd.n5810 gnd.n5405 19.3944
R16850 gnd.n5810 gnd.n5403 19.3944
R16851 gnd.n5819 gnd.n5403 19.3944
R16852 gnd.n5819 gnd.n5818 19.3944
R16853 gnd.n5818 gnd.n5817 19.3944
R16854 gnd.n5817 gnd.n5372 19.3944
R16855 gnd.n5871 gnd.n5372 19.3944
R16856 gnd.n5871 gnd.n5370 19.3944
R16857 gnd.n5877 gnd.n5370 19.3944
R16858 gnd.n5877 gnd.n5876 19.3944
R16859 gnd.n5876 gnd.n5345 19.3944
R16860 gnd.n5911 gnd.n5345 19.3944
R16861 gnd.n5911 gnd.n5343 19.3944
R16862 gnd.n5917 gnd.n5343 19.3944
R16863 gnd.n5917 gnd.n5916 19.3944
R16864 gnd.n5916 gnd.n5254 19.3944
R16865 gnd.n5956 gnd.n5254 19.3944
R16866 gnd.n5956 gnd.n5252 19.3944
R16867 gnd.n5962 gnd.n5252 19.3944
R16868 gnd.n5962 gnd.n5961 19.3944
R16869 gnd.n5961 gnd.n5226 19.3944
R16870 gnd.n5995 gnd.n5226 19.3944
R16871 gnd.n5995 gnd.n5224 19.3944
R16872 gnd.n6004 gnd.n5224 19.3944
R16873 gnd.n6004 gnd.n6003 19.3944
R16874 gnd.n6003 gnd.n6002 19.3944
R16875 gnd.n6002 gnd.n5196 19.3944
R16876 gnd.n6052 gnd.n5196 19.3944
R16877 gnd.n6052 gnd.n5194 19.3944
R16878 gnd.n6062 gnd.n5194 19.3944
R16879 gnd.n6062 gnd.n6061 19.3944
R16880 gnd.n6061 gnd.n6060 19.3944
R16881 gnd.n6060 gnd.n984 19.3944
R16882 gnd.n6499 gnd.n984 19.3944
R16883 gnd.n6499 gnd.n6498 19.3944
R16884 gnd.n6498 gnd.n6497 19.3944
R16885 gnd.n6497 gnd.n988 19.3944
R16886 gnd.n1008 gnd.n988 19.3944
R16887 gnd.n6485 gnd.n1008 19.3944
R16888 gnd.n6485 gnd.n6484 19.3944
R16889 gnd.n6484 gnd.n6483 19.3944
R16890 gnd.n6483 gnd.n1014 19.3944
R16891 gnd.n5096 gnd.n1014 19.3944
R16892 gnd.n6471 gnd.n5096 19.3944
R16893 gnd.n6468 gnd.n6467 19.3944
R16894 gnd.n6467 gnd.n6466 19.3944
R16895 gnd.n6466 gnd.n5102 19.3944
R16896 gnd.n6461 gnd.n5102 19.3944
R16897 gnd.n6461 gnd.n6460 19.3944
R16898 gnd.n6460 gnd.n6459 19.3944
R16899 gnd.n6459 gnd.n5109 19.3944
R16900 gnd.n6454 gnd.n5109 19.3944
R16901 gnd.n6454 gnd.n6453 19.3944
R16902 gnd.n6453 gnd.n6452 19.3944
R16903 gnd.n6452 gnd.n5116 19.3944
R16904 gnd.n6447 gnd.n5116 19.3944
R16905 gnd.n6447 gnd.n6446 19.3944
R16906 gnd.n6446 gnd.n6445 19.3944
R16907 gnd.n5604 gnd.n5500 19.3944
R16908 gnd.n5608 gnd.n5500 19.3944
R16909 gnd.n5608 gnd.n5490 19.3944
R16910 gnd.n5620 gnd.n5490 19.3944
R16911 gnd.n5620 gnd.n5488 19.3944
R16912 gnd.n5624 gnd.n5488 19.3944
R16913 gnd.n5624 gnd.n5477 19.3944
R16914 gnd.n5636 gnd.n5477 19.3944
R16915 gnd.n5636 gnd.n5475 19.3944
R16916 gnd.n5662 gnd.n5475 19.3944
R16917 gnd.n5662 gnd.n5661 19.3944
R16918 gnd.n5661 gnd.n5660 19.3944
R16919 gnd.n5660 gnd.n5659 19.3944
R16920 gnd.n5659 gnd.n5657 19.3944
R16921 gnd.n5657 gnd.n5656 19.3944
R16922 gnd.n5656 gnd.n5654 19.3944
R16923 gnd.n5654 gnd.n5653 19.3944
R16924 gnd.n5653 gnd.n5651 19.3944
R16925 gnd.n5651 gnd.n5650 19.3944
R16926 gnd.n5650 gnd.n5412 19.3944
R16927 gnd.n5799 gnd.n5412 19.3944
R16928 gnd.n5799 gnd.n5410 19.3944
R16929 gnd.n5805 gnd.n5410 19.3944
R16930 gnd.n5805 gnd.n5804 19.3944
R16931 gnd.n5804 gnd.n5379 19.3944
R16932 gnd.n5846 gnd.n5379 19.3944
R16933 gnd.n5846 gnd.n5377 19.3944
R16934 gnd.n5850 gnd.n5377 19.3944
R16935 gnd.n5864 gnd.n5850 19.3944
R16936 gnd.n5862 gnd.n5861 19.3944
R16937 gnd.n5858 gnd.n5857 19.3944
R16938 gnd.n5854 gnd.n5853 19.3944
R16939 gnd.n5932 gnd.n5326 19.3944
R16940 gnd.n5932 gnd.n5260 19.3944
R16941 gnd.n5951 gnd.n5260 19.3944
R16942 gnd.n5951 gnd.n5950 19.3944
R16943 gnd.n5950 gnd.n5949 19.3944
R16944 gnd.n5949 gnd.n5947 19.3944
R16945 gnd.n5947 gnd.n5946 19.3944
R16946 gnd.n5946 gnd.n5944 19.3944
R16947 gnd.n5944 gnd.n5943 19.3944
R16948 gnd.n5943 gnd.n5208 19.3944
R16949 gnd.n6018 gnd.n5208 19.3944
R16950 gnd.n6018 gnd.n5206 19.3944
R16951 gnd.n6037 gnd.n5206 19.3944
R16952 gnd.n6037 gnd.n6036 19.3944
R16953 gnd.n6036 gnd.n6035 19.3944
R16954 gnd.n6035 gnd.n6034 19.3944
R16955 gnd.n6034 gnd.n6032 19.3944
R16956 gnd.n6032 gnd.n6031 19.3944
R16957 gnd.n6031 gnd.n6028 19.3944
R16958 gnd.n6028 gnd.n5181 19.3944
R16959 gnd.n6369 gnd.n5181 19.3944
R16960 gnd.n6369 gnd.n5179 19.3944
R16961 gnd.n6375 gnd.n5179 19.3944
R16962 gnd.n6376 gnd.n6375 19.3944
R16963 gnd.n6379 gnd.n6376 19.3944
R16964 gnd.n6379 gnd.n5177 19.3944
R16965 gnd.n6383 gnd.n5177 19.3944
R16966 gnd.n6386 gnd.n6383 19.3944
R16967 gnd.n6387 gnd.n6386 19.3944
R16968 gnd.n5600 gnd.n5496 19.3944
R16969 gnd.n5612 gnd.n5496 19.3944
R16970 gnd.n5612 gnd.n5494 19.3944
R16971 gnd.n5616 gnd.n5494 19.3944
R16972 gnd.n5616 gnd.n5484 19.3944
R16973 gnd.n5628 gnd.n5484 19.3944
R16974 gnd.n5628 gnd.n5482 19.3944
R16975 gnd.n5632 gnd.n5482 19.3944
R16976 gnd.n5632 gnd.n5471 19.3944
R16977 gnd.n5726 gnd.n5471 19.3944
R16978 gnd.n5726 gnd.n5468 19.3944
R16979 gnd.n5731 gnd.n5468 19.3944
R16980 gnd.n5731 gnd.n5459 19.3944
R16981 gnd.n5741 gnd.n5459 19.3944
R16982 gnd.n5741 gnd.n5443 19.3944
R16983 gnd.n5758 gnd.n5443 19.3944
R16984 gnd.n5758 gnd.n5439 19.3944
R16985 gnd.n5771 gnd.n5439 19.3944
R16986 gnd.n5771 gnd.n5770 19.3944
R16987 gnd.n5770 gnd.n5418 19.3944
R16988 gnd.n5795 gnd.n5418 19.3944
R16989 gnd.n5795 gnd.n5794 19.3944
R16990 gnd.n5794 gnd.n5396 19.3944
R16991 gnd.n5824 gnd.n5396 19.3944
R16992 gnd.n5824 gnd.n5386 19.3944
R16993 gnd.n5842 gnd.n5386 19.3944
R16994 gnd.n5842 gnd.n5841 19.3944
R16995 gnd.n5841 gnd.n5840 19.3944
R16996 gnd.n5840 gnd.n5364 19.3944
R16997 gnd.n5882 gnd.n5364 19.3944
R16998 gnd.n5882 gnd.n5357 19.3944
R16999 gnd.n5893 gnd.n5357 19.3944
R17000 gnd.n5893 gnd.n5353 19.3944
R17001 gnd.n5906 gnd.n5353 19.3944
R17002 gnd.n5906 gnd.n5905 19.3944
R17003 gnd.n5905 gnd.n5332 19.3944
R17004 gnd.n5928 gnd.n5332 19.3944
R17005 gnd.n5928 gnd.n5927 19.3944
R17006 gnd.n5927 gnd.n5245 19.3944
R17007 gnd.n5967 gnd.n5245 19.3944
R17008 gnd.n5967 gnd.n5238 19.3944
R17009 gnd.n5978 gnd.n5238 19.3944
R17010 gnd.n5978 gnd.n5234 19.3944
R17011 gnd.n5990 gnd.n5234 19.3944
R17012 gnd.n5990 gnd.n5989 19.3944
R17013 gnd.n5989 gnd.n5214 19.3944
R17014 gnd.n6014 gnd.n5214 19.3944
R17015 gnd.n6014 gnd.n5202 19.3944
R17016 gnd.n6041 gnd.n5202 19.3944
R17017 gnd.n6041 gnd.n5188 19.3944
R17018 gnd.n6067 gnd.n5188 19.3944
R17019 gnd.n6067 gnd.n973 19.3944
R17020 gnd.n6506 gnd.n973 19.3944
R17021 gnd.n6506 gnd.n6505 19.3944
R17022 gnd.n6505 gnd.n6504 19.3944
R17023 gnd.n6504 gnd.n977 19.3944
R17024 gnd.n996 gnd.n977 19.3944
R17025 gnd.n6492 gnd.n996 19.3944
R17026 gnd.n6492 gnd.n6491 19.3944
R17027 gnd.n6491 gnd.n6490 19.3944
R17028 gnd.n6490 gnd.n1000 19.3944
R17029 gnd.n1022 gnd.n1000 19.3944
R17030 gnd.n6478 gnd.n1022 19.3944
R17031 gnd.n6478 gnd.n6477 19.3944
R17032 gnd.n6477 gnd.n6476 19.3944
R17033 gnd.n3204 gnd.n2560 19.3944
R17034 gnd.n3204 gnd.n3203 19.3944
R17035 gnd.n3203 gnd.n2564 19.3944
R17036 gnd.n3196 gnd.n2564 19.3944
R17037 gnd.n3196 gnd.n3195 19.3944
R17038 gnd.n3195 gnd.n2576 19.3944
R17039 gnd.n3188 gnd.n2576 19.3944
R17040 gnd.n3188 gnd.n3187 19.3944
R17041 gnd.n3187 gnd.n2587 19.3944
R17042 gnd.n3180 gnd.n2587 19.3944
R17043 gnd.n3180 gnd.n3179 19.3944
R17044 gnd.n3179 gnd.n2599 19.3944
R17045 gnd.n3172 gnd.n2599 19.3944
R17046 gnd.n3172 gnd.n3171 19.3944
R17047 gnd.n3171 gnd.n2610 19.3944
R17048 gnd.n3164 gnd.n2610 19.3944
R17049 gnd.n7135 gnd.n527 19.3944
R17050 gnd.n7135 gnd.n523 19.3944
R17051 gnd.n7141 gnd.n523 19.3944
R17052 gnd.n7141 gnd.n521 19.3944
R17053 gnd.n7145 gnd.n521 19.3944
R17054 gnd.n7145 gnd.n517 19.3944
R17055 gnd.n7151 gnd.n517 19.3944
R17056 gnd.n7151 gnd.n515 19.3944
R17057 gnd.n7155 gnd.n515 19.3944
R17058 gnd.n7155 gnd.n511 19.3944
R17059 gnd.n7161 gnd.n511 19.3944
R17060 gnd.n7161 gnd.n509 19.3944
R17061 gnd.n7165 gnd.n509 19.3944
R17062 gnd.n7165 gnd.n505 19.3944
R17063 gnd.n7171 gnd.n505 19.3944
R17064 gnd.n7171 gnd.n503 19.3944
R17065 gnd.n7175 gnd.n503 19.3944
R17066 gnd.n7175 gnd.n499 19.3944
R17067 gnd.n7181 gnd.n499 19.3944
R17068 gnd.n7181 gnd.n497 19.3944
R17069 gnd.n7185 gnd.n497 19.3944
R17070 gnd.n7185 gnd.n493 19.3944
R17071 gnd.n7191 gnd.n493 19.3944
R17072 gnd.n7191 gnd.n491 19.3944
R17073 gnd.n7195 gnd.n491 19.3944
R17074 gnd.n7195 gnd.n487 19.3944
R17075 gnd.n7201 gnd.n487 19.3944
R17076 gnd.n7201 gnd.n485 19.3944
R17077 gnd.n7205 gnd.n485 19.3944
R17078 gnd.n7205 gnd.n481 19.3944
R17079 gnd.n7211 gnd.n481 19.3944
R17080 gnd.n7211 gnd.n479 19.3944
R17081 gnd.n7215 gnd.n479 19.3944
R17082 gnd.n7215 gnd.n475 19.3944
R17083 gnd.n7221 gnd.n475 19.3944
R17084 gnd.n7221 gnd.n473 19.3944
R17085 gnd.n7225 gnd.n473 19.3944
R17086 gnd.n7225 gnd.n469 19.3944
R17087 gnd.n7231 gnd.n469 19.3944
R17088 gnd.n7231 gnd.n467 19.3944
R17089 gnd.n7235 gnd.n467 19.3944
R17090 gnd.n7235 gnd.n463 19.3944
R17091 gnd.n7241 gnd.n463 19.3944
R17092 gnd.n7241 gnd.n461 19.3944
R17093 gnd.n7245 gnd.n461 19.3944
R17094 gnd.n7245 gnd.n457 19.3944
R17095 gnd.n7251 gnd.n457 19.3944
R17096 gnd.n7251 gnd.n455 19.3944
R17097 gnd.n7255 gnd.n455 19.3944
R17098 gnd.n7255 gnd.n451 19.3944
R17099 gnd.n7261 gnd.n451 19.3944
R17100 gnd.n7261 gnd.n449 19.3944
R17101 gnd.n7265 gnd.n449 19.3944
R17102 gnd.n7265 gnd.n445 19.3944
R17103 gnd.n7271 gnd.n445 19.3944
R17104 gnd.n7271 gnd.n443 19.3944
R17105 gnd.n7275 gnd.n443 19.3944
R17106 gnd.n7275 gnd.n439 19.3944
R17107 gnd.n7281 gnd.n439 19.3944
R17108 gnd.n7281 gnd.n437 19.3944
R17109 gnd.n7285 gnd.n437 19.3944
R17110 gnd.n7285 gnd.n433 19.3944
R17111 gnd.n7291 gnd.n433 19.3944
R17112 gnd.n7291 gnd.n431 19.3944
R17113 gnd.n7295 gnd.n431 19.3944
R17114 gnd.n7295 gnd.n427 19.3944
R17115 gnd.n7301 gnd.n427 19.3944
R17116 gnd.n7301 gnd.n425 19.3944
R17117 gnd.n7305 gnd.n425 19.3944
R17118 gnd.n7305 gnd.n421 19.3944
R17119 gnd.n7311 gnd.n421 19.3944
R17120 gnd.n7311 gnd.n419 19.3944
R17121 gnd.n7315 gnd.n419 19.3944
R17122 gnd.n7315 gnd.n415 19.3944
R17123 gnd.n7321 gnd.n415 19.3944
R17124 gnd.n7321 gnd.n413 19.3944
R17125 gnd.n7325 gnd.n413 19.3944
R17126 gnd.n7325 gnd.n409 19.3944
R17127 gnd.n7331 gnd.n409 19.3944
R17128 gnd.n7331 gnd.n407 19.3944
R17129 gnd.n7337 gnd.n407 19.3944
R17130 gnd.n7337 gnd.n7336 19.3944
R17131 gnd.n7336 gnd.n403 19.3944
R17132 gnd.n7344 gnd.n403 19.3944
R17133 gnd.n6681 gnd.n799 19.3944
R17134 gnd.n6681 gnd.n797 19.3944
R17135 gnd.n6685 gnd.n797 19.3944
R17136 gnd.n6685 gnd.n793 19.3944
R17137 gnd.n6691 gnd.n793 19.3944
R17138 gnd.n6691 gnd.n791 19.3944
R17139 gnd.n6695 gnd.n791 19.3944
R17140 gnd.n6695 gnd.n787 19.3944
R17141 gnd.n6701 gnd.n787 19.3944
R17142 gnd.n6701 gnd.n785 19.3944
R17143 gnd.n6705 gnd.n785 19.3944
R17144 gnd.n6705 gnd.n781 19.3944
R17145 gnd.n6711 gnd.n781 19.3944
R17146 gnd.n6711 gnd.n779 19.3944
R17147 gnd.n6715 gnd.n779 19.3944
R17148 gnd.n6715 gnd.n775 19.3944
R17149 gnd.n6721 gnd.n775 19.3944
R17150 gnd.n6721 gnd.n773 19.3944
R17151 gnd.n6725 gnd.n773 19.3944
R17152 gnd.n6725 gnd.n769 19.3944
R17153 gnd.n6731 gnd.n769 19.3944
R17154 gnd.n6731 gnd.n767 19.3944
R17155 gnd.n6735 gnd.n767 19.3944
R17156 gnd.n6735 gnd.n763 19.3944
R17157 gnd.n6741 gnd.n763 19.3944
R17158 gnd.n6741 gnd.n761 19.3944
R17159 gnd.n6745 gnd.n761 19.3944
R17160 gnd.n6745 gnd.n757 19.3944
R17161 gnd.n6751 gnd.n757 19.3944
R17162 gnd.n6751 gnd.n755 19.3944
R17163 gnd.n6755 gnd.n755 19.3944
R17164 gnd.n6755 gnd.n751 19.3944
R17165 gnd.n6761 gnd.n751 19.3944
R17166 gnd.n6761 gnd.n749 19.3944
R17167 gnd.n6765 gnd.n749 19.3944
R17168 gnd.n6765 gnd.n745 19.3944
R17169 gnd.n6771 gnd.n745 19.3944
R17170 gnd.n6771 gnd.n743 19.3944
R17171 gnd.n6775 gnd.n743 19.3944
R17172 gnd.n6775 gnd.n739 19.3944
R17173 gnd.n6781 gnd.n739 19.3944
R17174 gnd.n6781 gnd.n737 19.3944
R17175 gnd.n6785 gnd.n737 19.3944
R17176 gnd.n6785 gnd.n733 19.3944
R17177 gnd.n6791 gnd.n733 19.3944
R17178 gnd.n6791 gnd.n731 19.3944
R17179 gnd.n6795 gnd.n731 19.3944
R17180 gnd.n6795 gnd.n727 19.3944
R17181 gnd.n6801 gnd.n727 19.3944
R17182 gnd.n6801 gnd.n725 19.3944
R17183 gnd.n6805 gnd.n725 19.3944
R17184 gnd.n6805 gnd.n721 19.3944
R17185 gnd.n6811 gnd.n721 19.3944
R17186 gnd.n6811 gnd.n719 19.3944
R17187 gnd.n6815 gnd.n719 19.3944
R17188 gnd.n6815 gnd.n715 19.3944
R17189 gnd.n6821 gnd.n715 19.3944
R17190 gnd.n6821 gnd.n713 19.3944
R17191 gnd.n6825 gnd.n713 19.3944
R17192 gnd.n6825 gnd.n709 19.3944
R17193 gnd.n6831 gnd.n709 19.3944
R17194 gnd.n6831 gnd.n707 19.3944
R17195 gnd.n6835 gnd.n707 19.3944
R17196 gnd.n6835 gnd.n703 19.3944
R17197 gnd.n6841 gnd.n703 19.3944
R17198 gnd.n6841 gnd.n701 19.3944
R17199 gnd.n6845 gnd.n701 19.3944
R17200 gnd.n6845 gnd.n697 19.3944
R17201 gnd.n6851 gnd.n697 19.3944
R17202 gnd.n6851 gnd.n695 19.3944
R17203 gnd.n6855 gnd.n695 19.3944
R17204 gnd.n6855 gnd.n691 19.3944
R17205 gnd.n6861 gnd.n691 19.3944
R17206 gnd.n6861 gnd.n689 19.3944
R17207 gnd.n6865 gnd.n689 19.3944
R17208 gnd.n6865 gnd.n685 19.3944
R17209 gnd.n6871 gnd.n685 19.3944
R17210 gnd.n6871 gnd.n683 19.3944
R17211 gnd.n6875 gnd.n683 19.3944
R17212 gnd.n6875 gnd.n679 19.3944
R17213 gnd.n6881 gnd.n679 19.3944
R17214 gnd.n6881 gnd.n677 19.3944
R17215 gnd.n6885 gnd.n677 19.3944
R17216 gnd.n6885 gnd.n673 19.3944
R17217 gnd.n6891 gnd.n673 19.3944
R17218 gnd.n6891 gnd.n671 19.3944
R17219 gnd.n6895 gnd.n671 19.3944
R17220 gnd.n6895 gnd.n667 19.3944
R17221 gnd.n6901 gnd.n667 19.3944
R17222 gnd.n6901 gnd.n665 19.3944
R17223 gnd.n6905 gnd.n665 19.3944
R17224 gnd.n6905 gnd.n661 19.3944
R17225 gnd.n6911 gnd.n661 19.3944
R17226 gnd.n6911 gnd.n659 19.3944
R17227 gnd.n6915 gnd.n659 19.3944
R17228 gnd.n6915 gnd.n655 19.3944
R17229 gnd.n6921 gnd.n655 19.3944
R17230 gnd.n6921 gnd.n653 19.3944
R17231 gnd.n6925 gnd.n653 19.3944
R17232 gnd.n6925 gnd.n649 19.3944
R17233 gnd.n6931 gnd.n649 19.3944
R17234 gnd.n6931 gnd.n647 19.3944
R17235 gnd.n6935 gnd.n647 19.3944
R17236 gnd.n6935 gnd.n643 19.3944
R17237 gnd.n6941 gnd.n643 19.3944
R17238 gnd.n6941 gnd.n641 19.3944
R17239 gnd.n6945 gnd.n641 19.3944
R17240 gnd.n6945 gnd.n637 19.3944
R17241 gnd.n6951 gnd.n637 19.3944
R17242 gnd.n6951 gnd.n635 19.3944
R17243 gnd.n6955 gnd.n635 19.3944
R17244 gnd.n6955 gnd.n631 19.3944
R17245 gnd.n6961 gnd.n631 19.3944
R17246 gnd.n6961 gnd.n629 19.3944
R17247 gnd.n6965 gnd.n629 19.3944
R17248 gnd.n6965 gnd.n625 19.3944
R17249 gnd.n6971 gnd.n625 19.3944
R17250 gnd.n6971 gnd.n623 19.3944
R17251 gnd.n6975 gnd.n623 19.3944
R17252 gnd.n6975 gnd.n619 19.3944
R17253 gnd.n6981 gnd.n619 19.3944
R17254 gnd.n6981 gnd.n617 19.3944
R17255 gnd.n6985 gnd.n617 19.3944
R17256 gnd.n6985 gnd.n613 19.3944
R17257 gnd.n6991 gnd.n613 19.3944
R17258 gnd.n6991 gnd.n611 19.3944
R17259 gnd.n6995 gnd.n611 19.3944
R17260 gnd.n6995 gnd.n607 19.3944
R17261 gnd.n7001 gnd.n607 19.3944
R17262 gnd.n7001 gnd.n605 19.3944
R17263 gnd.n7005 gnd.n605 19.3944
R17264 gnd.n7005 gnd.n601 19.3944
R17265 gnd.n7011 gnd.n601 19.3944
R17266 gnd.n7011 gnd.n599 19.3944
R17267 gnd.n7015 gnd.n599 19.3944
R17268 gnd.n7015 gnd.n595 19.3944
R17269 gnd.n7021 gnd.n595 19.3944
R17270 gnd.n7021 gnd.n593 19.3944
R17271 gnd.n7025 gnd.n593 19.3944
R17272 gnd.n7025 gnd.n589 19.3944
R17273 gnd.n7031 gnd.n589 19.3944
R17274 gnd.n7031 gnd.n587 19.3944
R17275 gnd.n7035 gnd.n587 19.3944
R17276 gnd.n7035 gnd.n583 19.3944
R17277 gnd.n7041 gnd.n583 19.3944
R17278 gnd.n7041 gnd.n581 19.3944
R17279 gnd.n7045 gnd.n581 19.3944
R17280 gnd.n7045 gnd.n577 19.3944
R17281 gnd.n7051 gnd.n577 19.3944
R17282 gnd.n7051 gnd.n575 19.3944
R17283 gnd.n7055 gnd.n575 19.3944
R17284 gnd.n7055 gnd.n571 19.3944
R17285 gnd.n7061 gnd.n571 19.3944
R17286 gnd.n7061 gnd.n569 19.3944
R17287 gnd.n7065 gnd.n569 19.3944
R17288 gnd.n7065 gnd.n565 19.3944
R17289 gnd.n7071 gnd.n565 19.3944
R17290 gnd.n7071 gnd.n563 19.3944
R17291 gnd.n7075 gnd.n563 19.3944
R17292 gnd.n7075 gnd.n559 19.3944
R17293 gnd.n7081 gnd.n559 19.3944
R17294 gnd.n7081 gnd.n557 19.3944
R17295 gnd.n7085 gnd.n557 19.3944
R17296 gnd.n7085 gnd.n553 19.3944
R17297 gnd.n7091 gnd.n553 19.3944
R17298 gnd.n7091 gnd.n551 19.3944
R17299 gnd.n7095 gnd.n551 19.3944
R17300 gnd.n7095 gnd.n547 19.3944
R17301 gnd.n7101 gnd.n547 19.3944
R17302 gnd.n7101 gnd.n545 19.3944
R17303 gnd.n7105 gnd.n545 19.3944
R17304 gnd.n7105 gnd.n541 19.3944
R17305 gnd.n7111 gnd.n541 19.3944
R17306 gnd.n7111 gnd.n539 19.3944
R17307 gnd.n7115 gnd.n539 19.3944
R17308 gnd.n7115 gnd.n535 19.3944
R17309 gnd.n7121 gnd.n535 19.3944
R17310 gnd.n7121 gnd.n533 19.3944
R17311 gnd.n7125 gnd.n533 19.3944
R17312 gnd.n7125 gnd.n529 19.3944
R17313 gnd.n7131 gnd.n529 19.3944
R17314 gnd.n4517 gnd.n4516 19.3944
R17315 gnd.n4516 gnd.n4515 19.3944
R17316 gnd.n4515 gnd.n4514 19.3944
R17317 gnd.n4514 gnd.n4512 19.3944
R17318 gnd.n4512 gnd.n4509 19.3944
R17319 gnd.n4509 gnd.n4508 19.3944
R17320 gnd.n4508 gnd.n4505 19.3944
R17321 gnd.n4505 gnd.n4504 19.3944
R17322 gnd.n4504 gnd.n4501 19.3944
R17323 gnd.n4501 gnd.n4500 19.3944
R17324 gnd.n4500 gnd.n4497 19.3944
R17325 gnd.n4497 gnd.n4496 19.3944
R17326 gnd.n4496 gnd.n4493 19.3944
R17327 gnd.n4493 gnd.n4492 19.3944
R17328 gnd.n4492 gnd.n4489 19.3944
R17329 gnd.n4489 gnd.n4488 19.3944
R17330 gnd.n4488 gnd.n4485 19.3944
R17331 gnd.n4483 gnd.n4480 19.3944
R17332 gnd.n4480 gnd.n4479 19.3944
R17333 gnd.n4479 gnd.n4476 19.3944
R17334 gnd.n4476 gnd.n4475 19.3944
R17335 gnd.n4475 gnd.n4472 19.3944
R17336 gnd.n4472 gnd.n4471 19.3944
R17337 gnd.n4471 gnd.n4468 19.3944
R17338 gnd.n4466 gnd.n4463 19.3944
R17339 gnd.n4463 gnd.n4462 19.3944
R17340 gnd.n4462 gnd.n4459 19.3944
R17341 gnd.n4459 gnd.n4458 19.3944
R17342 gnd.n4458 gnd.n4455 19.3944
R17343 gnd.n4455 gnd.n4454 19.3944
R17344 gnd.n4454 gnd.n4451 19.3944
R17345 gnd.n4451 gnd.n4450 19.3944
R17346 gnd.n4446 gnd.n4443 19.3944
R17347 gnd.n4443 gnd.n4442 19.3944
R17348 gnd.n4442 gnd.n4439 19.3944
R17349 gnd.n4439 gnd.n4438 19.3944
R17350 gnd.n4438 gnd.n4435 19.3944
R17351 gnd.n4435 gnd.n4434 19.3944
R17352 gnd.n4434 gnd.n4431 19.3944
R17353 gnd.n4431 gnd.n4430 19.3944
R17354 gnd.n4430 gnd.n4427 19.3944
R17355 gnd.n4427 gnd.n4426 19.3944
R17356 gnd.n4426 gnd.n4423 19.3944
R17357 gnd.n4423 gnd.n4422 19.3944
R17358 gnd.n4422 gnd.n4419 19.3944
R17359 gnd.n4419 gnd.n4418 19.3944
R17360 gnd.n4418 gnd.n4415 19.3944
R17361 gnd.n4415 gnd.n4414 19.3944
R17362 gnd.n4414 gnd.n4411 19.3944
R17363 gnd.n4411 gnd.n4410 19.3944
R17364 gnd.n4394 gnd.n1785 19.3944
R17365 gnd.n4394 gnd.n4393 19.3944
R17366 gnd.n4393 gnd.n1794 19.3944
R17367 gnd.n1966 gnd.n1794 19.3944
R17368 gnd.n4199 gnd.n1966 19.3944
R17369 gnd.n4200 gnd.n4199 19.3944
R17370 gnd.n4202 gnd.n4200 19.3944
R17371 gnd.n4202 gnd.n1961 19.3944
R17372 gnd.n4214 gnd.n1961 19.3944
R17373 gnd.n4215 gnd.n4214 19.3944
R17374 gnd.n4217 gnd.n4215 19.3944
R17375 gnd.n4218 gnd.n4217 19.3944
R17376 gnd.n4221 gnd.n4218 19.3944
R17377 gnd.n4222 gnd.n4221 19.3944
R17378 gnd.n4227 gnd.n4222 19.3944
R17379 gnd.n4228 gnd.n4227 19.3944
R17380 gnd.n4232 gnd.n4228 19.3944
R17381 gnd.n4232 gnd.n4231 19.3944
R17382 gnd.n4231 gnd.n4230 19.3944
R17383 gnd.n4230 gnd.n1936 19.3944
R17384 gnd.n4291 gnd.n1936 19.3944
R17385 gnd.n4292 gnd.n4291 19.3944
R17386 gnd.n4293 gnd.n4292 19.3944
R17387 gnd.n4297 gnd.n4293 19.3944
R17388 gnd.n4298 gnd.n4297 19.3944
R17389 gnd.n4299 gnd.n4298 19.3944
R17390 gnd.n4305 gnd.n4299 19.3944
R17391 gnd.n4305 gnd.n4304 19.3944
R17392 gnd.n4304 gnd.n378 19.3944
R17393 gnd.n7376 gnd.n378 19.3944
R17394 gnd.n7377 gnd.n7376 19.3944
R17395 gnd.n7378 gnd.n7377 19.3944
R17396 gnd.n7378 gnd.n372 19.3944
R17397 gnd.n7390 gnd.n372 19.3944
R17398 gnd.n7391 gnd.n7390 19.3944
R17399 gnd.n7392 gnd.n7391 19.3944
R17400 gnd.n7392 gnd.n366 19.3944
R17401 gnd.n7404 gnd.n366 19.3944
R17402 gnd.n7405 gnd.n7404 19.3944
R17403 gnd.n7406 gnd.n7405 19.3944
R17404 gnd.n7406 gnd.n360 19.3944
R17405 gnd.n7419 gnd.n360 19.3944
R17406 gnd.n7420 gnd.n7419 19.3944
R17407 gnd.n7436 gnd.n7420 19.3944
R17408 gnd.n7436 gnd.n7435 19.3944
R17409 gnd.n7435 gnd.n7434 19.3944
R17410 gnd.n7434 gnd.n7432 19.3944
R17411 gnd.n7432 gnd.n7431 19.3944
R17412 gnd.n7431 gnd.n7429 19.3944
R17413 gnd.n7429 gnd.n7428 19.3944
R17414 gnd.n7428 gnd.n7426 19.3944
R17415 gnd.n7426 gnd.n7425 19.3944
R17416 gnd.n7425 gnd.n7423 19.3944
R17417 gnd.n4397 gnd.n4396 19.3944
R17418 gnd.n4396 gnd.n1792 19.3944
R17419 gnd.n1817 gnd.n1792 19.3944
R17420 gnd.n4383 gnd.n1817 19.3944
R17421 gnd.n4383 gnd.n4382 19.3944
R17422 gnd.n4382 gnd.n4381 19.3944
R17423 gnd.n4381 gnd.n1822 19.3944
R17424 gnd.n4371 gnd.n1822 19.3944
R17425 gnd.n4371 gnd.n4370 19.3944
R17426 gnd.n4370 gnd.n4369 19.3944
R17427 gnd.n4369 gnd.n1842 19.3944
R17428 gnd.n4359 gnd.n1842 19.3944
R17429 gnd.n4359 gnd.n4358 19.3944
R17430 gnd.n4358 gnd.n4357 19.3944
R17431 gnd.n4357 gnd.n1862 19.3944
R17432 gnd.n4347 gnd.n1862 19.3944
R17433 gnd.n4347 gnd.n4346 19.3944
R17434 gnd.n4346 gnd.n4345 19.3944
R17435 gnd.n4345 gnd.n1882 19.3944
R17436 gnd.n4335 gnd.n1882 19.3944
R17437 gnd.n4335 gnd.n4334 19.3944
R17438 gnd.n4334 gnd.n4333 19.3944
R17439 gnd.n4333 gnd.n1902 19.3944
R17440 gnd.n1931 gnd.n1902 19.3944
R17441 gnd.n4311 gnd.n1931 19.3944
R17442 gnd.n4311 gnd.n4310 19.3944
R17443 gnd.n4310 gnd.n4309 19.3944
R17444 gnd.n4309 gnd.n1935 19.3944
R17445 gnd.n4301 gnd.n1935 19.3944
R17446 gnd.n4301 gnd.n108 19.3944
R17447 gnd.n7667 gnd.n108 19.3944
R17448 gnd.n7667 gnd.n7666 19.3944
R17449 gnd.n7666 gnd.n7665 19.3944
R17450 gnd.n7665 gnd.n112 19.3944
R17451 gnd.n7655 gnd.n112 19.3944
R17452 gnd.n7655 gnd.n7654 19.3944
R17453 gnd.n7654 gnd.n7653 19.3944
R17454 gnd.n7653 gnd.n130 19.3944
R17455 gnd.n7643 gnd.n130 19.3944
R17456 gnd.n7643 gnd.n7642 19.3944
R17457 gnd.n7642 gnd.n7641 19.3944
R17458 gnd.n7641 gnd.n151 19.3944
R17459 gnd.n7631 gnd.n151 19.3944
R17460 gnd.n7631 gnd.n7630 19.3944
R17461 gnd.n7630 gnd.n7629 19.3944
R17462 gnd.n7629 gnd.n170 19.3944
R17463 gnd.n7619 gnd.n170 19.3944
R17464 gnd.n7619 gnd.n7618 19.3944
R17465 gnd.n7618 gnd.n7617 19.3944
R17466 gnd.n7617 gnd.n190 19.3944
R17467 gnd.n7607 gnd.n190 19.3944
R17468 gnd.n7607 gnd.n7606 19.3944
R17469 gnd.n7606 gnd.n7605 19.3944
R17470 gnd.n7527 gnd.n279 19.3944
R17471 gnd.n7527 gnd.n283 19.3944
R17472 gnd.n286 gnd.n283 19.3944
R17473 gnd.n7520 gnd.n286 19.3944
R17474 gnd.n7520 gnd.n7519 19.3944
R17475 gnd.n7519 gnd.n7518 19.3944
R17476 gnd.n7518 gnd.n292 19.3944
R17477 gnd.n7513 gnd.n292 19.3944
R17478 gnd.n7513 gnd.n7512 19.3944
R17479 gnd.n7512 gnd.n7511 19.3944
R17480 gnd.n7511 gnd.n299 19.3944
R17481 gnd.n7506 gnd.n299 19.3944
R17482 gnd.n7506 gnd.n7505 19.3944
R17483 gnd.n7505 gnd.n7504 19.3944
R17484 gnd.n7504 gnd.n306 19.3944
R17485 gnd.n7499 gnd.n306 19.3944
R17486 gnd.n7499 gnd.n7498 19.3944
R17487 gnd.n7498 gnd.n7497 19.3944
R17488 gnd.n7565 gnd.n246 19.3944
R17489 gnd.n7560 gnd.n246 19.3944
R17490 gnd.n7560 gnd.n7559 19.3944
R17491 gnd.n7559 gnd.n7558 19.3944
R17492 gnd.n7558 gnd.n253 19.3944
R17493 gnd.n7553 gnd.n253 19.3944
R17494 gnd.n7553 gnd.n7552 19.3944
R17495 gnd.n7552 gnd.n7551 19.3944
R17496 gnd.n7551 gnd.n260 19.3944
R17497 gnd.n7546 gnd.n260 19.3944
R17498 gnd.n7546 gnd.n7545 19.3944
R17499 gnd.n7545 gnd.n7544 19.3944
R17500 gnd.n7544 gnd.n267 19.3944
R17501 gnd.n7539 gnd.n267 19.3944
R17502 gnd.n7539 gnd.n7538 19.3944
R17503 gnd.n7538 gnd.n7537 19.3944
R17504 gnd.n7537 gnd.n274 19.3944
R17505 gnd.n7532 gnd.n274 19.3944
R17506 gnd.n7598 gnd.n7597 19.3944
R17507 gnd.n7597 gnd.n7596 19.3944
R17508 gnd.n7596 gnd.n218 19.3944
R17509 gnd.n7591 gnd.n218 19.3944
R17510 gnd.n7591 gnd.n7590 19.3944
R17511 gnd.n7590 gnd.n7589 19.3944
R17512 gnd.n7589 gnd.n225 19.3944
R17513 gnd.n7584 gnd.n225 19.3944
R17514 gnd.n7584 gnd.n7583 19.3944
R17515 gnd.n7583 gnd.n7582 19.3944
R17516 gnd.n7582 gnd.n232 19.3944
R17517 gnd.n7577 gnd.n232 19.3944
R17518 gnd.n7577 gnd.n7576 19.3944
R17519 gnd.n7576 gnd.n7575 19.3944
R17520 gnd.n7575 gnd.n239 19.3944
R17521 gnd.n7570 gnd.n239 19.3944
R17522 gnd.n7570 gnd.n7569 19.3944
R17523 gnd.n7488 gnd.n7487 19.3944
R17524 gnd.n7487 gnd.n7486 19.3944
R17525 gnd.n7486 gnd.n321 19.3944
R17526 gnd.n7481 gnd.n321 19.3944
R17527 gnd.n7481 gnd.n7480 19.3944
R17528 gnd.n7480 gnd.n7479 19.3944
R17529 gnd.n7479 gnd.n328 19.3944
R17530 gnd.n7474 gnd.n328 19.3944
R17531 gnd.n7474 gnd.n7473 19.3944
R17532 gnd.n7473 gnd.n7472 19.3944
R17533 gnd.n7472 gnd.n335 19.3944
R17534 gnd.n7467 gnd.n335 19.3944
R17535 gnd.n7467 gnd.n7466 19.3944
R17536 gnd.n7466 gnd.n7465 19.3944
R17537 gnd.n7465 gnd.n342 19.3944
R17538 gnd.n7460 gnd.n342 19.3944
R17539 gnd.n4187 gnd.n1969 19.3944
R17540 gnd.n4188 gnd.n4187 19.3944
R17541 gnd.n4191 gnd.n4188 19.3944
R17542 gnd.n4191 gnd.n1967 19.3944
R17543 gnd.n4195 gnd.n1967 19.3944
R17544 gnd.n4195 gnd.n1964 19.3944
R17545 gnd.n4206 gnd.n1964 19.3944
R17546 gnd.n4206 gnd.n1962 19.3944
R17547 gnd.n4210 gnd.n1962 19.3944
R17548 gnd.n4210 gnd.n1954 19.3944
R17549 gnd.n4246 gnd.n1954 19.3944
R17550 gnd.n4246 gnd.n1955 19.3944
R17551 gnd.n4242 gnd.n1955 19.3944
R17552 gnd.n4242 gnd.n4241 19.3944
R17553 gnd.n4241 gnd.n4240 19.3944
R17554 gnd.n4240 gnd.n1960 19.3944
R17555 gnd.n4236 gnd.n1960 19.3944
R17556 gnd.n4236 gnd.n1940 19.3944
R17557 gnd.n4275 gnd.n1940 19.3944
R17558 gnd.n4275 gnd.n1937 19.3944
R17559 gnd.n4287 gnd.n1937 19.3944
R17560 gnd.n4287 gnd.n1938 19.3944
R17561 gnd.n4283 gnd.n1938 19.3944
R17562 gnd.n4283 gnd.n4282 19.3944
R17563 gnd.n4282 gnd.n4281 19.3944
R17564 gnd.n4281 gnd.n81 19.3944
R17565 gnd.n7680 gnd.n81 19.3944
R17566 gnd.n7680 gnd.n7679 19.3944
R17567 gnd.n7679 gnd.n83 19.3944
R17568 gnd.n7372 gnd.n83 19.3944
R17569 gnd.n7372 gnd.n377 19.3944
R17570 gnd.n7382 gnd.n377 19.3944
R17571 gnd.n7382 gnd.n375 19.3944
R17572 gnd.n7386 gnd.n375 19.3944
R17573 gnd.n7386 gnd.n370 19.3944
R17574 gnd.n7396 gnd.n370 19.3944
R17575 gnd.n7396 gnd.n368 19.3944
R17576 gnd.n7400 gnd.n368 19.3944
R17577 gnd.n7400 gnd.n365 19.3944
R17578 gnd.n7410 gnd.n365 19.3944
R17579 gnd.n7410 gnd.n363 19.3944
R17580 gnd.n7415 gnd.n363 19.3944
R17581 gnd.n7415 gnd.n359 19.3944
R17582 gnd.n7440 gnd.n359 19.3944
R17583 gnd.n7441 gnd.n7440 19.3944
R17584 gnd.n7441 gnd.n357 19.3944
R17585 gnd.n7445 gnd.n357 19.3944
R17586 gnd.n7447 gnd.n7445 19.3944
R17587 gnd.n7448 gnd.n7447 19.3944
R17588 gnd.n7448 gnd.n354 19.3944
R17589 gnd.n7452 gnd.n354 19.3944
R17590 gnd.n7454 gnd.n7452 19.3944
R17591 gnd.n7455 gnd.n7454 19.3944
R17592 gnd.n1803 gnd.n1802 19.3944
R17593 gnd.n4389 gnd.n1802 19.3944
R17594 gnd.n4389 gnd.n4388 19.3944
R17595 gnd.n4388 gnd.n4387 19.3944
R17596 gnd.n4387 gnd.n1809 19.3944
R17597 gnd.n4377 gnd.n1809 19.3944
R17598 gnd.n4377 gnd.n4376 19.3944
R17599 gnd.n4376 gnd.n4375 19.3944
R17600 gnd.n4375 gnd.n1832 19.3944
R17601 gnd.n4365 gnd.n1832 19.3944
R17602 gnd.n4365 gnd.n4364 19.3944
R17603 gnd.n4364 gnd.n4363 19.3944
R17604 gnd.n4363 gnd.n1853 19.3944
R17605 gnd.n4353 gnd.n1853 19.3944
R17606 gnd.n4353 gnd.n4352 19.3944
R17607 gnd.n4352 gnd.n4351 19.3944
R17608 gnd.n4351 gnd.n1872 19.3944
R17609 gnd.n4341 gnd.n1872 19.3944
R17610 gnd.n4341 gnd.n4340 19.3944
R17611 gnd.n4340 gnd.n4339 19.3944
R17612 gnd.n4339 gnd.n1893 19.3944
R17613 gnd.n4329 gnd.n1893 19.3944
R17614 gnd.n1908 gnd.n97 19.3944
R17615 gnd.n1926 gnd.n97 19.3944
R17616 gnd.n4316 gnd.n4315 19.3944
R17617 gnd.n7675 gnd.n7674 19.3944
R17618 gnd.n7671 gnd.n92 19.3944
R17619 gnd.n7671 gnd.n99 19.3944
R17620 gnd.n7661 gnd.n99 19.3944
R17621 gnd.n7661 gnd.n7660 19.3944
R17622 gnd.n7660 gnd.n7659 19.3944
R17623 gnd.n7659 gnd.n121 19.3944
R17624 gnd.n7649 gnd.n121 19.3944
R17625 gnd.n7649 gnd.n7648 19.3944
R17626 gnd.n7648 gnd.n7647 19.3944
R17627 gnd.n7647 gnd.n141 19.3944
R17628 gnd.n7637 gnd.n141 19.3944
R17629 gnd.n7637 gnd.n7636 19.3944
R17630 gnd.n7636 gnd.n7635 19.3944
R17631 gnd.n7635 gnd.n161 19.3944
R17632 gnd.n7625 gnd.n161 19.3944
R17633 gnd.n7625 gnd.n7624 19.3944
R17634 gnd.n7624 gnd.n7623 19.3944
R17635 gnd.n7623 gnd.n181 19.3944
R17636 gnd.n7613 gnd.n181 19.3944
R17637 gnd.n7613 gnd.n7612 19.3944
R17638 gnd.n7612 gnd.n7611 19.3944
R17639 gnd.n7611 gnd.n200 19.3944
R17640 gnd.n7601 gnd.n200 19.3944
R17641 gnd.n2729 gnd.n2722 19.3944
R17642 gnd.n2729 gnd.n2720 19.3944
R17643 gnd.n2733 gnd.n2720 19.3944
R17644 gnd.n2733 gnd.n2718 19.3944
R17645 gnd.n2894 gnd.n2718 19.3944
R17646 gnd.n2894 gnd.n2716 19.3944
R17647 gnd.n2898 gnd.n2716 19.3944
R17648 gnd.n2898 gnd.n2714 19.3944
R17649 gnd.n2903 gnd.n2714 19.3944
R17650 gnd.n2903 gnd.n2712 19.3944
R17651 gnd.n2907 gnd.n2712 19.3944
R17652 gnd.n2918 gnd.n2907 19.3944
R17653 gnd.n2916 gnd.n2915 19.3944
R17654 gnd.n2912 gnd.n2911 19.3944
R17655 gnd.n2970 gnd.n2671 19.3944
R17656 gnd.n2993 gnd.n2972 19.3944
R17657 gnd.n2991 gnd.n2990 19.3944
R17658 gnd.n2990 gnd.n2974 19.3944
R17659 gnd.n2986 gnd.n2974 19.3944
R17660 gnd.n2986 gnd.n2985 19.3944
R17661 gnd.n2985 gnd.n2984 19.3944
R17662 gnd.n2984 gnd.n2982 19.3944
R17663 gnd.n2982 gnd.n2647 19.3944
R17664 gnd.n2647 gnd.n2645 19.3944
R17665 gnd.n3060 gnd.n2645 19.3944
R17666 gnd.n3060 gnd.n2643 19.3944
R17667 gnd.n3064 gnd.n2643 19.3944
R17668 gnd.n3064 gnd.n2641 19.3944
R17669 gnd.n3068 gnd.n2641 19.3944
R17670 gnd.n3068 gnd.n2639 19.3944
R17671 gnd.n3118 gnd.n2639 19.3944
R17672 gnd.n3118 gnd.n3117 19.3944
R17673 gnd.n3117 gnd.n3116 19.3944
R17674 gnd.n3116 gnd.n3074 19.3944
R17675 gnd.n3112 gnd.n3074 19.3944
R17676 gnd.n3112 gnd.n3111 19.3944
R17677 gnd.n3111 gnd.n3110 19.3944
R17678 gnd.n3110 gnd.n3080 19.3944
R17679 gnd.n3105 gnd.n3080 19.3944
R17680 gnd.n3105 gnd.n3104 19.3944
R17681 gnd.n3104 gnd.n3103 19.3944
R17682 gnd.n3103 gnd.n3086 19.3944
R17683 gnd.n3097 gnd.n3086 19.3944
R17684 gnd.n3097 gnd.n3096 19.3944
R17685 gnd.n3096 gnd.n3095 19.3944
R17686 gnd.n3095 gnd.n2401 19.3944
R17687 gnd.n3243 gnd.n2401 19.3944
R17688 gnd.n3243 gnd.n2399 19.3944
R17689 gnd.n3249 gnd.n2399 19.3944
R17690 gnd.n3249 gnd.n3248 19.3944
R17691 gnd.n3248 gnd.n2376 19.3944
R17692 gnd.n3273 gnd.n2376 19.3944
R17693 gnd.n3273 gnd.n2374 19.3944
R17694 gnd.n3286 gnd.n2374 19.3944
R17695 gnd.n3286 gnd.n3285 19.3944
R17696 gnd.n3285 gnd.n3284 19.3944
R17697 gnd.n3284 gnd.n3281 19.3944
R17698 gnd.n3281 gnd.n1495 19.3944
R17699 gnd.n4706 gnd.n1495 19.3944
R17700 gnd.n4706 gnd.n4705 19.3944
R17701 gnd.n4705 gnd.n4704 19.3944
R17702 gnd.n4704 gnd.n1499 19.3944
R17703 gnd.n4692 gnd.n1499 19.3944
R17704 gnd.n4692 gnd.n4691 19.3944
R17705 gnd.n4691 gnd.n4690 19.3944
R17706 gnd.n4690 gnd.n1515 19.3944
R17707 gnd.n4678 gnd.n1515 19.3944
R17708 gnd.n4678 gnd.n4677 19.3944
R17709 gnd.n4677 gnd.n4676 19.3944
R17710 gnd.n4676 gnd.n1533 19.3944
R17711 gnd.n3484 gnd.n1533 19.3944
R17712 gnd.n3484 gnd.n3481 19.3944
R17713 gnd.n3498 gnd.n3481 19.3944
R17714 gnd.n3498 gnd.n3497 19.3944
R17715 gnd.n3497 gnd.n3496 19.3944
R17716 gnd.n3496 gnd.n3491 19.3944
R17717 gnd.n3491 gnd.n2276 19.3944
R17718 gnd.n3566 gnd.n2276 19.3944
R17719 gnd.n3566 gnd.n2274 19.3944
R17720 gnd.n3570 gnd.n2274 19.3944
R17721 gnd.n3570 gnd.n2252 19.3944
R17722 gnd.n3605 gnd.n2252 19.3944
R17723 gnd.n3605 gnd.n2250 19.3944
R17724 gnd.n3609 gnd.n2250 19.3944
R17725 gnd.n3609 gnd.n2230 19.3944
R17726 gnd.n3659 gnd.n2230 19.3944
R17727 gnd.n3659 gnd.n2228 19.3944
R17728 gnd.n3663 gnd.n2228 19.3944
R17729 gnd.n3663 gnd.n2211 19.3944
R17730 gnd.n3685 gnd.n2211 19.3944
R17731 gnd.n3685 gnd.n2209 19.3944
R17732 gnd.n3689 gnd.n2209 19.3944
R17733 gnd.n3689 gnd.n2188 19.3944
R17734 gnd.n3751 gnd.n2188 19.3944
R17735 gnd.n3751 gnd.n2186 19.3944
R17736 gnd.n3755 gnd.n2186 19.3944
R17737 gnd.n3755 gnd.n2166 19.3944
R17738 gnd.n3781 gnd.n2166 19.3944
R17739 gnd.n3781 gnd.n2164 19.3944
R17740 gnd.n3785 gnd.n2164 19.3944
R17741 gnd.n3785 gnd.n2144 19.3944
R17742 gnd.n3812 gnd.n2144 19.3944
R17743 gnd.n3812 gnd.n2142 19.3944
R17744 gnd.n3816 gnd.n2142 19.3944
R17745 gnd.n3816 gnd.n2118 19.3944
R17746 gnd.n3861 gnd.n2118 19.3944
R17747 gnd.n3861 gnd.n2116 19.3944
R17748 gnd.n3865 gnd.n2116 19.3944
R17749 gnd.n3865 gnd.n2102 19.3944
R17750 gnd.n3892 gnd.n2102 19.3944
R17751 gnd.n3892 gnd.n2100 19.3944
R17752 gnd.n3896 gnd.n2100 19.3944
R17753 gnd.n3896 gnd.n2048 19.3944
R17754 gnd.n4063 gnd.n2048 19.3944
R17755 gnd.n4063 gnd.n2046 19.3944
R17756 gnd.n4067 gnd.n2046 19.3944
R17757 gnd.n4067 gnd.n2035 19.3944
R17758 gnd.n4083 gnd.n2035 19.3944
R17759 gnd.n4083 gnd.n2033 19.3944
R17760 gnd.n4087 gnd.n2033 19.3944
R17761 gnd.n4087 gnd.n2022 19.3944
R17762 gnd.n4103 gnd.n2022 19.3944
R17763 gnd.n4103 gnd.n2020 19.3944
R17764 gnd.n4109 gnd.n2020 19.3944
R17765 gnd.n4109 gnd.n4108 19.3944
R17766 gnd.n4108 gnd.n2007 19.3944
R17767 gnd.n4127 gnd.n2007 19.3944
R17768 gnd.n4127 gnd.n2005 19.3944
R17769 gnd.n4175 gnd.n2005 19.3944
R17770 gnd.n4175 gnd.n4174 19.3944
R17771 gnd.n4174 gnd.n4173 19.3944
R17772 gnd.n4173 gnd.n4133 19.3944
R17773 gnd.n4169 gnd.n4133 19.3944
R17774 gnd.n4169 gnd.n4168 19.3944
R17775 gnd.n4168 gnd.n4167 19.3944
R17776 gnd.n4167 gnd.n4139 19.3944
R17777 gnd.n4163 gnd.n4139 19.3944
R17778 gnd.n4163 gnd.n4162 19.3944
R17779 gnd.n4162 gnd.n4161 19.3944
R17780 gnd.n4161 gnd.n4145 19.3944
R17781 gnd.n4157 gnd.n4145 19.3944
R17782 gnd.n4157 gnd.n4156 19.3944
R17783 gnd.n4156 gnd.n4155 19.3944
R17784 gnd.n4155 gnd.n4153 19.3944
R17785 gnd.n4153 gnd.n1952 19.3944
R17786 gnd.n1952 gnd.n1950 19.3944
R17787 gnd.n4253 gnd.n1950 19.3944
R17788 gnd.n4253 gnd.n1948 19.3944
R17789 gnd.n4257 gnd.n1948 19.3944
R17790 gnd.n4257 gnd.n1946 19.3944
R17791 gnd.n4261 gnd.n1946 19.3944
R17792 gnd.n4261 gnd.n1944 19.3944
R17793 gnd.n4270 gnd.n1944 19.3944
R17794 gnd.n4270 gnd.n4269 19.3944
R17795 gnd.n4269 gnd.n4268 19.3944
R17796 gnd.n4324 gnd.n1915 19.3944
R17797 gnd.n4322 gnd.n4321 19.3944
R17798 gnd.n1920 gnd.n1919 19.3944
R17799 gnd.n7367 gnd.n384 19.3944
R17800 gnd.n7365 gnd.n7364 19.3944
R17801 gnd.n7364 gnd.n386 19.3944
R17802 gnd.n7360 gnd.n386 19.3944
R17803 gnd.n7360 gnd.n7359 19.3944
R17804 gnd.n7359 gnd.n7358 19.3944
R17805 gnd.n7358 gnd.n392 19.3944
R17806 gnd.n7354 gnd.n392 19.3944
R17807 gnd.n7354 gnd.n7353 19.3944
R17808 gnd.n7353 gnd.n7352 19.3944
R17809 gnd.n7352 gnd.n398 19.3944
R17810 gnd.n7348 gnd.n398 19.3944
R17811 gnd.n7348 gnd.n7347 19.3944
R17812 gnd.n5089 gnd.n5088 19.3944
R17813 gnd.n5088 gnd.n5087 19.3944
R17814 gnd.n5087 gnd.n5086 19.3944
R17815 gnd.n5086 gnd.n5084 19.3944
R17816 gnd.n5084 gnd.n5081 19.3944
R17817 gnd.n5081 gnd.n5080 19.3944
R17818 gnd.n5080 gnd.n5077 19.3944
R17819 gnd.n5077 gnd.n5076 19.3944
R17820 gnd.n5076 gnd.n5073 19.3944
R17821 gnd.n5073 gnd.n5072 19.3944
R17822 gnd.n5072 gnd.n5069 19.3944
R17823 gnd.n5069 gnd.n5068 19.3944
R17824 gnd.n5068 gnd.n5065 19.3944
R17825 gnd.n5065 gnd.n5064 19.3944
R17826 gnd.n5064 gnd.n5061 19.3944
R17827 gnd.n5061 gnd.n5060 19.3944
R17828 gnd.n5060 gnd.n5057 19.3944
R17829 gnd.n5055 gnd.n5052 19.3944
R17830 gnd.n5052 gnd.n5051 19.3944
R17831 gnd.n5051 gnd.n5048 19.3944
R17832 gnd.n5048 gnd.n5047 19.3944
R17833 gnd.n5047 gnd.n5044 19.3944
R17834 gnd.n5044 gnd.n5043 19.3944
R17835 gnd.n5043 gnd.n5040 19.3944
R17836 gnd.n5040 gnd.n5039 19.3944
R17837 gnd.n5039 gnd.n5036 19.3944
R17838 gnd.n5036 gnd.n5035 19.3944
R17839 gnd.n5035 gnd.n5032 19.3944
R17840 gnd.n5032 gnd.n5031 19.3944
R17841 gnd.n5031 gnd.n5028 19.3944
R17842 gnd.n5028 gnd.n5027 19.3944
R17843 gnd.n5027 gnd.n5024 19.3944
R17844 gnd.n5024 gnd.n5023 19.3944
R17845 gnd.n5023 gnd.n5020 19.3944
R17846 gnd.n5020 gnd.n5019 19.3944
R17847 gnd.n5015 gnd.n5012 19.3944
R17848 gnd.n5012 gnd.n5011 19.3944
R17849 gnd.n5011 gnd.n5008 19.3944
R17850 gnd.n5008 gnd.n5007 19.3944
R17851 gnd.n5007 gnd.n5004 19.3944
R17852 gnd.n5004 gnd.n5003 19.3944
R17853 gnd.n5003 gnd.n5000 19.3944
R17854 gnd.n5000 gnd.n4999 19.3944
R17855 gnd.n4999 gnd.n4996 19.3944
R17856 gnd.n4996 gnd.n4995 19.3944
R17857 gnd.n4995 gnd.n4992 19.3944
R17858 gnd.n4992 gnd.n4991 19.3944
R17859 gnd.n4991 gnd.n4988 19.3944
R17860 gnd.n4988 gnd.n4987 19.3944
R17861 gnd.n4987 gnd.n4984 19.3944
R17862 gnd.n4984 gnd.n4983 19.3944
R17863 gnd.n4983 gnd.n4980 19.3944
R17864 gnd.n4980 gnd.n4979 19.3944
R17865 gnd.n2765 gnd.n2764 19.3944
R17866 gnd.n2768 gnd.n2765 19.3944
R17867 gnd.n2768 gnd.n2760 19.3944
R17868 gnd.n2774 gnd.n2760 19.3944
R17869 gnd.n2775 gnd.n2774 19.3944
R17870 gnd.n2778 gnd.n2775 19.3944
R17871 gnd.n2778 gnd.n2758 19.3944
R17872 gnd.n2784 gnd.n2758 19.3944
R17873 gnd.n2785 gnd.n2784 19.3944
R17874 gnd.n2788 gnd.n2785 19.3944
R17875 gnd.n2788 gnd.n2756 19.3944
R17876 gnd.n2794 gnd.n2756 19.3944
R17877 gnd.n2795 gnd.n2794 19.3944
R17878 gnd.n2798 gnd.n2795 19.3944
R17879 gnd.n2798 gnd.n2752 19.3944
R17880 gnd.n2802 gnd.n2752 19.3944
R17881 gnd.n2809 gnd.n2808 19.3944
R17882 gnd.n2811 gnd.n2809 19.3944
R17883 gnd.n2811 gnd.n2746 19.3944
R17884 gnd.n2816 gnd.n2746 19.3944
R17885 gnd.n2817 gnd.n2816 19.3944
R17886 gnd.n2819 gnd.n2817 19.3944
R17887 gnd.n2819 gnd.n2744 19.3944
R17888 gnd.n2824 gnd.n2744 19.3944
R17889 gnd.n2825 gnd.n2824 19.3944
R17890 gnd.n2844 gnd.n2825 19.3944
R17891 gnd.n2844 gnd.n2742 19.3944
R17892 gnd.n2849 gnd.n2742 19.3944
R17893 gnd.n2849 gnd.n2736 19.3944
R17894 gnd.n2888 gnd.n2736 19.3944
R17895 gnd.n2888 gnd.n2887 19.3944
R17896 gnd.n2887 gnd.n2886 19.3944
R17897 gnd.n2886 gnd.n2740 19.3944
R17898 gnd.n2876 gnd.n2740 19.3944
R17899 gnd.n2876 gnd.n2875 19.3944
R17900 gnd.n2875 gnd.n2874 19.3944
R17901 gnd.n2874 gnd.n2868 19.3944
R17902 gnd.n2868 gnd.n2867 19.3944
R17903 gnd.n2867 gnd.n2695 19.3944
R17904 gnd.n2936 gnd.n2695 19.3944
R17905 gnd.n2936 gnd.n2693 19.3944
R17906 gnd.n2946 gnd.n2693 19.3944
R17907 gnd.n2946 gnd.n2945 19.3944
R17908 gnd.n2945 gnd.n2941 19.3944
R17909 gnd.n2941 gnd.n2665 19.3944
R17910 gnd.n2998 gnd.n2665 19.3944
R17911 gnd.n2998 gnd.n2663 19.3944
R17912 gnd.n3002 gnd.n2663 19.3944
R17913 gnd.n3002 gnd.n2660 19.3944
R17914 gnd.n3013 gnd.n2660 19.3944
R17915 gnd.n3013 gnd.n2658 19.3944
R17916 gnd.n3017 gnd.n2658 19.3944
R17917 gnd.n3017 gnd.n2649 19.3944
R17918 gnd.n3053 gnd.n2649 19.3944
R17919 gnd.n3053 gnd.n2650 19.3944
R17920 gnd.n3049 gnd.n2650 19.3944
R17921 gnd.n3049 gnd.n3048 19.3944
R17922 gnd.n3048 gnd.n3047 19.3944
R17923 gnd.n3047 gnd.n2655 19.3944
R17924 gnd.n3043 gnd.n2655 19.3944
R17925 gnd.n3043 gnd.n3042 19.3944
R17926 gnd.n3042 gnd.n3041 19.3944
R17927 gnd.n3041 gnd.n2633 19.3944
R17928 gnd.n3129 gnd.n2633 19.3944
R17929 gnd.n3129 gnd.n2631 19.3944
R17930 gnd.n3134 gnd.n2631 19.3944
R17931 gnd.n3134 gnd.n2628 19.3944
R17932 gnd.n3145 gnd.n2628 19.3944
R17933 gnd.n3146 gnd.n3145 19.3944
R17934 gnd.n4971 gnd.n1139 19.3944
R17935 gnd.n2827 gnd.n1139 19.3944
R17936 gnd.n2828 gnd.n2827 19.3944
R17937 gnd.n2830 gnd.n2828 19.3944
R17938 gnd.n2831 gnd.n2830 19.3944
R17939 gnd.n2834 gnd.n2831 19.3944
R17940 gnd.n2835 gnd.n2834 19.3944
R17941 gnd.n2837 gnd.n2835 19.3944
R17942 gnd.n2838 gnd.n2837 19.3944
R17943 gnd.n2840 gnd.n2838 19.3944
R17944 gnd.n2840 gnd.n2741 19.3944
R17945 gnd.n2853 gnd.n2741 19.3944
R17946 gnd.n2854 gnd.n2853 19.3944
R17947 gnd.n2856 gnd.n2854 19.3944
R17948 gnd.n2857 gnd.n2856 19.3944
R17949 gnd.n2882 gnd.n2857 19.3944
R17950 gnd.n2882 gnd.n2881 19.3944
R17951 gnd.n2881 gnd.n2880 19.3944
R17952 gnd.n2880 gnd.n2859 19.3944
R17953 gnd.n2870 gnd.n2859 19.3944
R17954 gnd.n2870 gnd.n2869 19.3944
R17955 gnd.n2869 gnd.n2707 19.3944
R17956 gnd.n2925 gnd.n2707 19.3944
R17957 gnd.n2926 gnd.n2925 19.3944
R17958 gnd.n2926 gnd.n2689 19.3944
R17959 gnd.n2950 gnd.n2689 19.3944
R17960 gnd.n2951 gnd.n2950 19.3944
R17961 gnd.n2953 gnd.n2951 19.3944
R17962 gnd.n2955 gnd.n2953 19.3944
R17963 gnd.n2955 gnd.n2954 19.3944
R17964 gnd.n2954 gnd.n2662 19.3944
R17965 gnd.n3006 gnd.n2662 19.3944
R17966 gnd.n3007 gnd.n3006 19.3944
R17967 gnd.n3009 gnd.n3007 19.3944
R17968 gnd.n3009 gnd.n2657 19.3944
R17969 gnd.n3021 gnd.n2657 19.3944
R17970 gnd.n3022 gnd.n3021 19.3944
R17971 gnd.n3024 gnd.n3022 19.3944
R17972 gnd.n3025 gnd.n3024 19.3944
R17973 gnd.n3028 gnd.n3025 19.3944
R17974 gnd.n3029 gnd.n3028 19.3944
R17975 gnd.n3034 gnd.n3029 19.3944
R17976 gnd.n3035 gnd.n3034 19.3944
R17977 gnd.n3036 gnd.n3035 19.3944
R17978 gnd.n3036 gnd.n2634 19.3944
R17979 gnd.n3123 gnd.n2634 19.3944
R17980 gnd.n3124 gnd.n3123 19.3944
R17981 gnd.n3125 gnd.n3124 19.3944
R17982 gnd.n3125 gnd.n2629 19.3944
R17983 gnd.n3138 gnd.n2629 19.3944
R17984 gnd.n3139 gnd.n3138 19.3944
R17985 gnd.n3141 gnd.n3139 19.3944
R17986 gnd.n3141 gnd.n3140 19.3944
R17987 gnd.n1158 gnd.n1137 19.3944
R17988 gnd.n1159 gnd.n1158 19.3944
R17989 gnd.n4960 gnd.n1159 19.3944
R17990 gnd.n4960 gnd.n4959 19.3944
R17991 gnd.n4959 gnd.n4958 19.3944
R17992 gnd.n4958 gnd.n1163 19.3944
R17993 gnd.n4948 gnd.n1163 19.3944
R17994 gnd.n4948 gnd.n4947 19.3944
R17995 gnd.n4947 gnd.n4946 19.3944
R17996 gnd.n4946 gnd.n1182 19.3944
R17997 gnd.n4936 gnd.n1182 19.3944
R17998 gnd.n4936 gnd.n4935 19.3944
R17999 gnd.n4935 gnd.n4934 19.3944
R18000 gnd.n4934 gnd.n1202 19.3944
R18001 gnd.n4924 gnd.n1202 19.3944
R18002 gnd.n4924 gnd.n4923 19.3944
R18003 gnd.n4923 gnd.n4922 19.3944
R18004 gnd.n4922 gnd.n1222 19.3944
R18005 gnd.n4912 gnd.n1222 19.3944
R18006 gnd.n4912 gnd.n4911 19.3944
R18007 gnd.n4911 gnd.n4910 19.3944
R18008 gnd.n4910 gnd.n1243 19.3944
R18009 gnd.n2921 gnd.n1243 19.3944
R18010 gnd.n2921 gnd.n2704 19.3944
R18011 gnd.n2929 gnd.n2704 19.3944
R18012 gnd.n2929 gnd.n2685 19.3944
R18013 gnd.n2959 gnd.n2685 19.3944
R18014 gnd.n2959 gnd.n2958 19.3944
R18015 gnd.n2958 gnd.n2957 19.3944
R18016 gnd.n2957 gnd.n1268 19.3944
R18017 gnd.n4898 gnd.n1268 19.3944
R18018 gnd.n4898 gnd.n4897 19.3944
R18019 gnd.n4897 gnd.n4896 19.3944
R18020 gnd.n4896 gnd.n1272 19.3944
R18021 gnd.n4886 gnd.n1272 19.3944
R18022 gnd.n4886 gnd.n4885 19.3944
R18023 gnd.n4885 gnd.n4884 19.3944
R18024 gnd.n4884 gnd.n1291 19.3944
R18025 gnd.n4874 gnd.n1291 19.3944
R18026 gnd.n4874 gnd.n4873 19.3944
R18027 gnd.n4873 gnd.n4872 19.3944
R18028 gnd.n4872 gnd.n1311 19.3944
R18029 gnd.n4862 gnd.n1311 19.3944
R18030 gnd.n4862 gnd.n4861 19.3944
R18031 gnd.n4861 gnd.n4860 19.3944
R18032 gnd.n4860 gnd.n1331 19.3944
R18033 gnd.n4850 gnd.n1331 19.3944
R18034 gnd.n4850 gnd.n4849 19.3944
R18035 gnd.n4849 gnd.n4848 19.3944
R18036 gnd.n4848 gnd.n1351 19.3944
R18037 gnd.n4838 gnd.n1351 19.3944
R18038 gnd.n4838 gnd.n4837 19.3944
R18039 gnd.n4837 gnd.n4836 19.3944
R18040 gnd.n4829 gnd.n4828 19.3944
R18041 gnd.n4828 gnd.n1380 19.3944
R18042 gnd.n1382 gnd.n1380 19.3944
R18043 gnd.n4821 gnd.n1382 19.3944
R18044 gnd.n4821 gnd.n4820 19.3944
R18045 gnd.n4820 gnd.n4819 19.3944
R18046 gnd.n4819 gnd.n1389 19.3944
R18047 gnd.n4814 gnd.n1389 19.3944
R18048 gnd.n4814 gnd.n4813 19.3944
R18049 gnd.n4813 gnd.n4812 19.3944
R18050 gnd.n4812 gnd.n1396 19.3944
R18051 gnd.n4807 gnd.n1396 19.3944
R18052 gnd.n4807 gnd.n4806 19.3944
R18053 gnd.n4806 gnd.n4805 19.3944
R18054 gnd.n4805 gnd.n1403 19.3944
R18055 gnd.n4800 gnd.n1403 19.3944
R18056 gnd.n4800 gnd.n4799 19.3944
R18057 gnd.n2503 gnd.n2463 19.3944
R18058 gnd.n2507 gnd.n2463 19.3944
R18059 gnd.n2507 gnd.n2461 19.3944
R18060 gnd.n2513 gnd.n2461 19.3944
R18061 gnd.n2513 gnd.n2459 19.3944
R18062 gnd.n2517 gnd.n2459 19.3944
R18063 gnd.n2517 gnd.n2457 19.3944
R18064 gnd.n2523 gnd.n2457 19.3944
R18065 gnd.n2523 gnd.n2455 19.3944
R18066 gnd.n2527 gnd.n2455 19.3944
R18067 gnd.n2527 gnd.n2453 19.3944
R18068 gnd.n2533 gnd.n2453 19.3944
R18069 gnd.n2533 gnd.n2451 19.3944
R18070 gnd.n2537 gnd.n2451 19.3944
R18071 gnd.n2537 gnd.n2449 19.3944
R18072 gnd.n2543 gnd.n2449 19.3944
R18073 gnd.n2543 gnd.n2447 19.3944
R18074 gnd.n2547 gnd.n2447 19.3944
R18075 gnd.n2476 gnd.n1425 19.3944
R18076 gnd.n2483 gnd.n2476 19.3944
R18077 gnd.n2483 gnd.n2473 19.3944
R18078 gnd.n2487 gnd.n2473 19.3944
R18079 gnd.n2487 gnd.n2471 19.3944
R18080 gnd.n2493 gnd.n2471 19.3944
R18081 gnd.n2493 gnd.n2469 19.3944
R18082 gnd.n2497 gnd.n2469 19.3944
R18083 gnd.n4797 gnd.n1412 19.3944
R18084 gnd.n4792 gnd.n1412 19.3944
R18085 gnd.n4792 gnd.n4791 19.3944
R18086 gnd.n4791 gnd.n4790 19.3944
R18087 gnd.n4790 gnd.n1419 19.3944
R18088 gnd.n4785 gnd.n1419 19.3944
R18089 gnd.n4785 gnd.n4784 19.3944
R18090 gnd.n4966 gnd.n1145 19.3944
R18091 gnd.n4966 gnd.n4965 19.3944
R18092 gnd.n4965 gnd.n4964 19.3944
R18093 gnd.n4964 gnd.n1150 19.3944
R18094 gnd.n4954 gnd.n1150 19.3944
R18095 gnd.n4954 gnd.n4953 19.3944
R18096 gnd.n4953 gnd.n4952 19.3944
R18097 gnd.n4952 gnd.n1173 19.3944
R18098 gnd.n4942 gnd.n1173 19.3944
R18099 gnd.n4942 gnd.n4941 19.3944
R18100 gnd.n4941 gnd.n4940 19.3944
R18101 gnd.n4940 gnd.n1192 19.3944
R18102 gnd.n4930 gnd.n1192 19.3944
R18103 gnd.n4930 gnd.n4929 19.3944
R18104 gnd.n4929 gnd.n4928 19.3944
R18105 gnd.n4928 gnd.n1213 19.3944
R18106 gnd.n4918 gnd.n1213 19.3944
R18107 gnd.n4918 gnd.n4917 19.3944
R18108 gnd.n4917 gnd.n4916 19.3944
R18109 gnd.n4916 gnd.n1233 19.3944
R18110 gnd.n4906 gnd.n1233 19.3944
R18111 gnd.n4906 gnd.n4905 19.3944
R18112 gnd.n1258 gnd.n1252 19.3944
R18113 gnd.n2702 gnd.n1258 19.3944
R18114 gnd.n2678 gnd.n2677 19.3944
R18115 gnd.n2965 gnd.n2964 19.3944
R18116 gnd.n4902 gnd.n1259 19.3944
R18117 gnd.n4902 gnd.n1260 19.3944
R18118 gnd.n4892 gnd.n1260 19.3944
R18119 gnd.n4892 gnd.n4891 19.3944
R18120 gnd.n4891 gnd.n4890 19.3944
R18121 gnd.n4890 gnd.n1281 19.3944
R18122 gnd.n4880 gnd.n1281 19.3944
R18123 gnd.n4880 gnd.n4879 19.3944
R18124 gnd.n4879 gnd.n4878 19.3944
R18125 gnd.n4878 gnd.n1302 19.3944
R18126 gnd.n4868 gnd.n1302 19.3944
R18127 gnd.n4868 gnd.n4867 19.3944
R18128 gnd.n4867 gnd.n4866 19.3944
R18129 gnd.n4866 gnd.n1321 19.3944
R18130 gnd.n4856 gnd.n1321 19.3944
R18131 gnd.n4856 gnd.n4855 19.3944
R18132 gnd.n4855 gnd.n4854 19.3944
R18133 gnd.n4854 gnd.n1342 19.3944
R18134 gnd.n4844 gnd.n1342 19.3944
R18135 gnd.n4844 gnd.n4843 19.3944
R18136 gnd.n4843 gnd.n4842 19.3944
R18137 gnd.n4842 gnd.n1362 19.3944
R18138 gnd.n4832 gnd.n1362 19.3944
R18139 gnd.n6675 gnd.n6674 19.3944
R18140 gnd.n6674 gnd.n6673 19.3944
R18141 gnd.n6673 gnd.n806 19.3944
R18142 gnd.n6667 gnd.n806 19.3944
R18143 gnd.n6667 gnd.n6666 19.3944
R18144 gnd.n6666 gnd.n6665 19.3944
R18145 gnd.n6665 gnd.n814 19.3944
R18146 gnd.n6659 gnd.n814 19.3944
R18147 gnd.n6659 gnd.n6658 19.3944
R18148 gnd.n6658 gnd.n6657 19.3944
R18149 gnd.n6657 gnd.n822 19.3944
R18150 gnd.n6651 gnd.n822 19.3944
R18151 gnd.n6651 gnd.n6650 19.3944
R18152 gnd.n6650 gnd.n6649 19.3944
R18153 gnd.n6649 gnd.n830 19.3944
R18154 gnd.n6643 gnd.n830 19.3944
R18155 gnd.n6643 gnd.n6642 19.3944
R18156 gnd.n6642 gnd.n6641 19.3944
R18157 gnd.n6641 gnd.n838 19.3944
R18158 gnd.n6635 gnd.n838 19.3944
R18159 gnd.n6635 gnd.n6634 19.3944
R18160 gnd.n6634 gnd.n6633 19.3944
R18161 gnd.n6633 gnd.n846 19.3944
R18162 gnd.n6627 gnd.n846 19.3944
R18163 gnd.n6627 gnd.n6626 19.3944
R18164 gnd.n6626 gnd.n6625 19.3944
R18165 gnd.n6625 gnd.n854 19.3944
R18166 gnd.n6619 gnd.n854 19.3944
R18167 gnd.n6619 gnd.n6618 19.3944
R18168 gnd.n6618 gnd.n6617 19.3944
R18169 gnd.n6617 gnd.n862 19.3944
R18170 gnd.n6611 gnd.n862 19.3944
R18171 gnd.n6611 gnd.n6610 19.3944
R18172 gnd.n6610 gnd.n6609 19.3944
R18173 gnd.n6609 gnd.n870 19.3944
R18174 gnd.n6603 gnd.n870 19.3944
R18175 gnd.n6603 gnd.n6602 19.3944
R18176 gnd.n6602 gnd.n6601 19.3944
R18177 gnd.n6601 gnd.n878 19.3944
R18178 gnd.n6595 gnd.n878 19.3944
R18179 gnd.n6595 gnd.n6594 19.3944
R18180 gnd.n6594 gnd.n6593 19.3944
R18181 gnd.n6593 gnd.n886 19.3944
R18182 gnd.n6587 gnd.n886 19.3944
R18183 gnd.n6587 gnd.n6586 19.3944
R18184 gnd.n6586 gnd.n6585 19.3944
R18185 gnd.n6585 gnd.n894 19.3944
R18186 gnd.n6579 gnd.n894 19.3944
R18187 gnd.n6579 gnd.n6578 19.3944
R18188 gnd.n6578 gnd.n6577 19.3944
R18189 gnd.n6577 gnd.n902 19.3944
R18190 gnd.n6571 gnd.n902 19.3944
R18191 gnd.n6571 gnd.n6570 19.3944
R18192 gnd.n6570 gnd.n6569 19.3944
R18193 gnd.n6569 gnd.n910 19.3944
R18194 gnd.n6563 gnd.n910 19.3944
R18195 gnd.n6563 gnd.n6562 19.3944
R18196 gnd.n6562 gnd.n6561 19.3944
R18197 gnd.n6561 gnd.n918 19.3944
R18198 gnd.n6555 gnd.n918 19.3944
R18199 gnd.n6555 gnd.n6554 19.3944
R18200 gnd.n6554 gnd.n6553 19.3944
R18201 gnd.n6553 gnd.n926 19.3944
R18202 gnd.n6547 gnd.n926 19.3944
R18203 gnd.n6547 gnd.n6546 19.3944
R18204 gnd.n6546 gnd.n6545 19.3944
R18205 gnd.n6545 gnd.n934 19.3944
R18206 gnd.n6539 gnd.n934 19.3944
R18207 gnd.n6539 gnd.n6538 19.3944
R18208 gnd.n6538 gnd.n6537 19.3944
R18209 gnd.n6537 gnd.n942 19.3944
R18210 gnd.n6531 gnd.n942 19.3944
R18211 gnd.n6531 gnd.n6530 19.3944
R18212 gnd.n6530 gnd.n6529 19.3944
R18213 gnd.n6529 gnd.n950 19.3944
R18214 gnd.n6523 gnd.n950 19.3944
R18215 gnd.n6523 gnd.n6522 19.3944
R18216 gnd.n6522 gnd.n6521 19.3944
R18217 gnd.n6521 gnd.n958 19.3944
R18218 gnd.n6515 gnd.n958 19.3944
R18219 gnd.n6515 gnd.n6514 19.3944
R18220 gnd.n6514 gnd.n6513 19.3944
R18221 gnd.n6513 gnd.n966 19.3944
R18222 gnd.n2725 gnd.n966 19.3944
R18223 gnd.n3229 gnd.n2414 19.3944
R18224 gnd.n3229 gnd.n2415 19.3944
R18225 gnd.n2415 gnd.n2392 19.3944
R18226 gnd.n3254 gnd.n2392 19.3944
R18227 gnd.n3254 gnd.n2389 19.3944
R18228 gnd.n3259 gnd.n2389 19.3944
R18229 gnd.n3259 gnd.n2390 19.3944
R18230 gnd.n2390 gnd.n2366 19.3944
R18231 gnd.n3291 gnd.n2366 19.3944
R18232 gnd.n3291 gnd.n2363 19.3944
R18233 gnd.n3296 gnd.n2363 19.3944
R18234 gnd.n3296 gnd.n2364 19.3944
R18235 gnd.n2364 gnd.n2352 19.3944
R18236 gnd.n3419 gnd.n2352 19.3944
R18237 gnd.n3419 gnd.n2350 19.3944
R18238 gnd.n3423 gnd.n2350 19.3944
R18239 gnd.n3423 gnd.n2338 19.3944
R18240 gnd.n3437 gnd.n2338 19.3944
R18241 gnd.n3437 gnd.n2335 19.3944
R18242 gnd.n3449 gnd.n2335 19.3944
R18243 gnd.n3449 gnd.n2336 19.3944
R18244 gnd.n3445 gnd.n2336 19.3944
R18245 gnd.n3445 gnd.n3444 19.3944
R18246 gnd.n3444 gnd.n1540 19.3944
R18247 gnd.n4671 gnd.n1540 19.3944
R18248 gnd.n4671 gnd.n1541 19.3944
R18249 gnd.n4667 gnd.n1541 19.3944
R18250 gnd.n4667 gnd.n4666 19.3944
R18251 gnd.n4666 gnd.n4665 19.3944
R18252 gnd.n4665 gnd.n1547 19.3944
R18253 gnd.n4661 gnd.n1547 19.3944
R18254 gnd.n4661 gnd.n4660 19.3944
R18255 gnd.n4660 gnd.n4659 19.3944
R18256 gnd.n4659 gnd.n1552 19.3944
R18257 gnd.n4655 gnd.n1552 19.3944
R18258 gnd.n4655 gnd.n4654 19.3944
R18259 gnd.n4654 gnd.n4653 19.3944
R18260 gnd.n4653 gnd.n1557 19.3944
R18261 gnd.n4649 gnd.n1557 19.3944
R18262 gnd.n4649 gnd.n4648 19.3944
R18263 gnd.n4648 gnd.n4647 19.3944
R18264 gnd.n4647 gnd.n1562 19.3944
R18265 gnd.n4643 gnd.n1562 19.3944
R18266 gnd.n4643 gnd.n4642 19.3944
R18267 gnd.n4642 gnd.n4641 19.3944
R18268 gnd.n4641 gnd.n1567 19.3944
R18269 gnd.n4637 gnd.n1567 19.3944
R18270 gnd.n4637 gnd.n4636 19.3944
R18271 gnd.n4636 gnd.n4635 19.3944
R18272 gnd.n4635 gnd.n1572 19.3944
R18273 gnd.n4631 gnd.n1572 19.3944
R18274 gnd.n4631 gnd.n4630 19.3944
R18275 gnd.n4630 gnd.n4629 19.3944
R18276 gnd.n4629 gnd.n1577 19.3944
R18277 gnd.n4625 gnd.n1577 19.3944
R18278 gnd.n4625 gnd.n4624 19.3944
R18279 gnd.n4624 gnd.n4623 19.3944
R18280 gnd.n4623 gnd.n1582 19.3944
R18281 gnd.n4619 gnd.n1582 19.3944
R18282 gnd.n4619 gnd.n4618 19.3944
R18283 gnd.n4618 gnd.n4617 19.3944
R18284 gnd.n4617 gnd.n1587 19.3944
R18285 gnd.n4613 gnd.n1587 19.3944
R18286 gnd.n4613 gnd.n4612 19.3944
R18287 gnd.n4612 gnd.n4611 19.3944
R18288 gnd.n4611 gnd.n1592 19.3944
R18289 gnd.n4607 gnd.n1592 19.3944
R18290 gnd.n4607 gnd.n4606 19.3944
R18291 gnd.n4606 gnd.n4605 19.3944
R18292 gnd.n4605 gnd.n1597 19.3944
R18293 gnd.n4601 gnd.n1597 19.3944
R18294 gnd.n4601 gnd.n4600 19.3944
R18295 gnd.n4600 gnd.n4599 19.3944
R18296 gnd.n4599 gnd.n1602 19.3944
R18297 gnd.n4595 gnd.n1602 19.3944
R18298 gnd.n4595 gnd.n4594 19.3944
R18299 gnd.n4594 gnd.n4593 19.3944
R18300 gnd.n4593 gnd.n1607 19.3944
R18301 gnd.n4589 gnd.n1607 19.3944
R18302 gnd.n4589 gnd.n4588 19.3944
R18303 gnd.n4588 gnd.n4587 19.3944
R18304 gnd.n4587 gnd.n1612 19.3944
R18305 gnd.n4583 gnd.n4582 19.3944
R18306 gnd.n4582 gnd.n4581 19.3944
R18307 gnd.n4581 gnd.n1617 19.3944
R18308 gnd.n4577 gnd.n1617 19.3944
R18309 gnd.n4577 gnd.n4576 19.3944
R18310 gnd.n4576 gnd.n4575 19.3944
R18311 gnd.n4575 gnd.n1622 19.3944
R18312 gnd.n4570 gnd.n1622 19.3944
R18313 gnd.n4570 gnd.n4569 19.3944
R18314 gnd.n4569 gnd.n1627 19.3944
R18315 gnd.n4562 gnd.n1627 19.3944
R18316 gnd.n4562 gnd.n4561 19.3944
R18317 gnd.n4561 gnd.n1636 19.3944
R18318 gnd.n4554 gnd.n1636 19.3944
R18319 gnd.n4554 gnd.n4553 19.3944
R18320 gnd.n4553 gnd.n1644 19.3944
R18321 gnd.n4546 gnd.n1644 19.3944
R18322 gnd.n4546 gnd.n4545 19.3944
R18323 gnd.n4545 gnd.n1652 19.3944
R18324 gnd.n4538 gnd.n1652 19.3944
R18325 gnd.n4538 gnd.n4537 19.3944
R18326 gnd.n4537 gnd.n1660 19.3944
R18327 gnd.n4530 gnd.n1660 19.3944
R18328 gnd.n4530 gnd.n4529 19.3944
R18329 gnd.n1998 gnd.n1975 19.3944
R18330 gnd.n4182 gnd.n1975 19.3944
R18331 gnd.n4182 gnd.n4181 19.3944
R18332 gnd.n5880 gnd.t27 18.8012
R18333 gnd.n5919 gnd.t63 18.8012
R18334 gnd.n5723 gnd.n5465 18.4825
R18335 gnd.n6509 gnd.n968 18.4825
R18336 gnd.n4468 gnd.n4467 18.4247
R18337 gnd.n4784 gnd.n4783 18.4247
R18338 gnd.n4526 gnd.n4525 18.2308
R18339 gnd.n3164 gnd.n3163 18.2308
R18340 gnd.n7460 gnd.n7459 18.2308
R18341 gnd.n2803 gnd.n2802 18.2308
R18342 gnd.t28 gnd.n5407 18.1639
R18343 gnd.n1184 gnd.n1177 18.1639
R18344 gnd.n7627 gnd.n172 18.1639
R18345 gnd.n5436 gnd.t25 17.5266
R18346 gnd.t131 gnd.n1167 17.5266
R18347 gnd.n4852 gnd.t90 17.5266
R18348 gnd.n4379 gnd.t99 17.5266
R18349 gnd.n7621 gnd.t71 17.5266
R18350 gnd.t36 gnd.n5383 16.8893
R18351 gnd.n4876 gnd.t82 16.8893
R18352 gnd.n4355 gnd.t110 16.8893
R18353 gnd.n4450 gnd.n4447 16.6793
R18354 gnd.n7532 gnd.n7531 16.6793
R18355 gnd.n5019 gnd.n5016 16.6793
R18356 gnd.n2497 gnd.n2467 16.6793
R18357 gnd.t255 gnd.n5492 16.2519
R18358 gnd.n5350 gnd.t35 16.2519
R18359 gnd.n4900 gnd.t163 16.2519
R18360 gnd.n4331 gnd.t140 16.2519
R18361 gnd.n3221 gnd.n2419 15.9333
R18362 gnd.n3221 gnd.n2433 15.9333
R18363 gnd.n3088 gnd.n3087 15.9333
R18364 gnd.n3087 gnd.n2410 15.9333
R18365 gnd.n3231 gnd.n2410 15.9333
R18366 gnd.n3231 gnd.n2411 15.9333
R18367 gnd.n3241 gnd.n2403 15.9333
R18368 gnd.n3241 gnd.n3240 15.9333
R18369 gnd.n3240 gnd.n2394 15.9333
R18370 gnd.n3252 gnd.n2394 15.9333
R18371 gnd.n3252 gnd.n3251 15.9333
R18372 gnd.n3251 gnd.n2396 15.9333
R18373 gnd.n2396 gnd.n2385 15.9333
R18374 gnd.n3261 gnd.n2385 15.9333
R18375 gnd.n2386 gnd.n2378 15.9333
R18376 gnd.n3271 gnd.n2378 15.9333
R18377 gnd.n3271 gnd.n3270 15.9333
R18378 gnd.n3270 gnd.n2368 15.9333
R18379 gnd.n3289 gnd.n2368 15.9333
R18380 gnd.n3289 gnd.n3288 15.9333
R18381 gnd.n3288 gnd.n2370 15.9333
R18382 gnd.n2372 gnd.n2370 15.9333
R18383 gnd.n3298 gnd.n2361 15.9333
R18384 gnd.n2361 gnd.n1433 15.9333
R18385 gnd.n3416 gnd.n1465 15.9333
R18386 gnd.n3414 gnd.n1491 15.9333
R18387 gnd.n3407 gnd.n3406 15.9333
R18388 gnd.n2340 gnd.n1502 15.9333
R18389 gnd.n3390 gnd.n3389 15.9333
R18390 gnd.n3442 gnd.n2324 15.9333
R18391 gnd.n3508 gnd.n2313 15.9333
R18392 gnd.n3536 gnd.n2298 15.9333
R18393 gnd.n3554 gnd.n2286 15.9333
R18394 gnd.n3554 gnd.n2287 15.9333
R18395 gnd.n2269 gnd.n2257 15.9333
R18396 gnd.n3612 gnd.n2239 15.9333
R18397 gnd.n3657 gnd.n3656 15.9333
R18398 gnd.n3665 gnd.n2226 15.9333
R18399 gnd.n3749 gnd.n2190 15.9333
R18400 gnd.n3749 gnd.n2193 15.9333
R18401 gnd.n3758 gnd.n3757 15.9333
R18402 gnd.n3788 gnd.n3787 15.9333
R18403 gnd.n3725 gnd.n2138 15.9333
R18404 gnd.n3851 gnd.n2125 15.9333
R18405 gnd.n3882 gnd.n3881 15.9333
R18406 gnd.n4061 gnd.n2050 15.9333
R18407 gnd.n4070 gnd.n2043 15.9333
R18408 gnd.n4069 gnd.n2044 15.9333
R18409 gnd.n2044 gnd.n2037 15.9333
R18410 gnd.n4078 gnd.n2037 15.9333
R18411 gnd.n4081 gnd.n4078 15.9333
R18412 gnd.n4081 gnd.n4080 15.9333
R18413 gnd.n4080 gnd.n2030 15.9333
R18414 gnd.n4090 gnd.n2030 15.9333
R18415 gnd.n4090 gnd.n4089 15.9333
R18416 gnd.n2031 gnd.n2024 15.9333
R18417 gnd.n4098 gnd.n2024 15.9333
R18418 gnd.n4101 gnd.n4098 15.9333
R18419 gnd.n4101 gnd.n4100 15.9333
R18420 gnd.n4100 gnd.n2016 15.9333
R18421 gnd.n4112 gnd.n2016 15.9333
R18422 gnd.n4112 gnd.n4111 15.9333
R18423 gnd.n4111 gnd.n2017 15.9333
R18424 gnd.n4121 gnd.n2009 15.9333
R18425 gnd.n4122 gnd.n4121 15.9333
R18426 gnd.n4124 gnd.n4122 15.9333
R18427 gnd.n4125 gnd.n4124 15.9333
R18428 gnd.n4178 gnd.n1978 15.9333
R18429 gnd.n4178 gnd.n4177 15.9333
R18430 gnd.n6319 gnd.n6317 15.6674
R18431 gnd.n6287 gnd.n6285 15.6674
R18432 gnd.n6255 gnd.n6253 15.6674
R18433 gnd.n6224 gnd.n6222 15.6674
R18434 gnd.n6192 gnd.n6190 15.6674
R18435 gnd.n6160 gnd.n6158 15.6674
R18436 gnd.n6128 gnd.n6126 15.6674
R18437 gnd.n6097 gnd.n6095 15.6674
R18438 gnd.n5610 gnd.t255 15.6146
R18439 gnd.t251 gnd.n6480 15.6146
R18440 gnd.n6384 gnd.t345 15.6146
R18441 gnd.n2923 gnd.t116 15.6146
R18442 gnd.t307 gnd.n2403 15.6146
R18443 gnd.n2017 gnd.t291 15.6146
R18444 gnd.n7374 gnd.t159 15.6146
R18445 gnd.n4407 gnd.n4402 15.3217
R18446 gnd.n7492 gnd.n315 15.3217
R18447 gnd.n4976 gnd.n1133 15.3217
R18448 gnd.n2552 gnd.n2445 15.3217
R18449 gnd.n4680 gnd.n1527 15.296
R18450 gnd.n2321 gnd.n1537 15.296
R18451 gnd.n3613 gnd.n3611 15.296
R18452 gnd.n3654 gnd.n2235 15.296
R18453 gnd.n3802 gnd.n3801 15.296
R18454 gnd.n3819 gnd.n3818 15.296
R18455 gnd.n3907 gnd.n3906 15.0827
R18456 gnd.n1477 gnd.n1472 15.0481
R18457 gnd.n3917 gnd.n3916 15.0481
R18458 gnd.n6048 gnd.t30 14.9773
R18459 gnd.n4926 gnd.t86 14.9773
R18460 gnd.n2372 gnd.t67 14.9773
R18461 gnd.t229 gnd.n4069 14.9773
R18462 gnd.n7402 gnd.t94 14.9773
R18463 gnd.n3435 gnd.n2341 14.6587
R18464 gnd.t5 gnd.n1519 14.6587
R18465 gnd.n3528 gnd.n3526 14.6587
R18466 gnd.n3547 gnd.n3546 14.6587
R18467 gnd.n3693 gnd.n3692 14.6587
R18468 gnd.n2184 gnd.n2175 14.6587
R18469 gnd.n3827 gnd.t1 14.6587
R18470 gnd.n3883 gnd.n2110 14.6587
R18471 gnd.n3992 gnd.n2050 14.6587
R18472 gnd.t330 gnd.n2043 14.6587
R18473 gnd.n6501 gnd.t50 14.34
R18474 gnd.t23 gnd.n993 14.34
R18475 gnd.n4950 gnd.t131 14.34
R18476 gnd.t71 gnd.n175 14.34
R18477 gnd.n4688 gnd.n4687 14.0214
R18478 gnd.n3507 gnd.n2315 14.0214
R18479 gnd.n3603 gnd.n3602 14.0214
R18480 gnd.n2225 gnd.n2218 14.0214
R18481 gnd.n3735 gnd.n2162 14.0214
R18482 gnd.n3859 gnd.n2120 14.0214
R18483 gnd.t17 gnd.n5807 13.7027
R18484 gnd.n4944 gnd.n1184 13.7027
R18485 gnd.n2291 gnd.t41 13.7027
R18486 gnd.n3691 gnd.t48 13.7027
R18487 gnd.n7438 gnd.n172 13.7027
R18488 gnd.n5692 gnd.n5688 13.5763
R18489 gnd.n6440 gnd.n5125 13.5763
R18490 gnd.n5724 gnd.n5723 13.384
R18491 gnd.n3501 gnd.n3478 13.384
R18492 gnd.n3593 gnd.n3592 13.384
R18493 gnd.n2219 gnd.n2213 13.384
R18494 gnd.n3778 gnd.n2170 13.384
R18495 gnd.n3715 gnd.n3714 13.384
R18496 gnd.n1488 gnd.n1469 13.1884
R18497 gnd.n1483 gnd.n1482 13.1884
R18498 gnd.n1482 gnd.n1481 13.1884
R18499 gnd.n3910 gnd.n3905 13.1884
R18500 gnd.n3911 gnd.n3910 13.1884
R18501 gnd.n1484 gnd.n1471 13.146
R18502 gnd.n1480 gnd.n1471 13.146
R18503 gnd.n3909 gnd.n3908 13.146
R18504 gnd.n3909 gnd.n3904 13.146
R18505 gnd.n3425 gnd.t65 13.0654
R18506 gnd.t12 gnd.n2106 13.0654
R18507 gnd.n6320 gnd.n6316 12.8005
R18508 gnd.n6288 gnd.n6284 12.8005
R18509 gnd.n6256 gnd.n6252 12.8005
R18510 gnd.n6225 gnd.n6221 12.8005
R18511 gnd.n6193 gnd.n6189 12.8005
R18512 gnd.n6161 gnd.n6157 12.8005
R18513 gnd.n6129 gnd.n6125 12.8005
R18514 gnd.n6098 gnd.n6094 12.8005
R18515 gnd.n4694 gnd.n1509 12.7467
R18516 gnd.n3574 gnd.n3572 12.7467
R18517 gnd.n3680 gnd.n2205 12.7467
R18518 gnd.n4779 gnd.n1465 12.4281
R18519 gnd.n4061 gnd.n4060 12.4281
R18520 gnd.n5695 gnd.n5692 12.4126
R18521 gnd.n6445 gnd.n5125 12.4126
R18522 gnd.n4776 gnd.n4713 12.1761
R18523 gnd.n3989 gnd.n3988 12.1761
R18524 gnd.n3383 gnd.n1525 12.1094
R18525 gnd.t59 gnd.n3471 12.1094
R18526 gnd.t2 gnd.n2152 12.1094
R18527 gnd.n3825 gnd.n2133 12.1094
R18528 gnd.n3836 gnd.t259 12.1094
R18529 gnd.n6324 gnd.n6323 12.0247
R18530 gnd.n6292 gnd.n6291 12.0247
R18531 gnd.n6260 gnd.n6259 12.0247
R18532 gnd.n6229 gnd.n6228 12.0247
R18533 gnd.n6197 gnd.n6196 12.0247
R18534 gnd.n6165 gnd.n6164 12.0247
R18535 gnd.n6133 gnd.n6132 12.0247
R18536 gnd.n6102 gnd.n6101 12.0247
R18537 gnd.n2891 gnd.t86 11.7908
R18538 gnd.t94 gnd.n143 11.7908
R18539 gnd.n3100 gnd.n1381 11.4721
R18540 gnd.t262 gnd.n3415 11.4721
R18541 gnd.n4709 gnd.n4708 11.4721
R18542 gnd.n3898 gnd.n2098 11.4721
R18543 gnd.n4520 gnd.n1676 11.4721
R18544 gnd.n6327 gnd.n6314 11.249
R18545 gnd.n6295 gnd.n6282 11.249
R18546 gnd.n6263 gnd.n6250 11.249
R18547 gnd.n6232 gnd.n6219 11.249
R18548 gnd.n6200 gnd.n6187 11.249
R18549 gnd.n6168 gnd.n6155 11.249
R18550 gnd.n6136 gnd.n6123 11.249
R18551 gnd.n6105 gnd.n6092 11.249
R18552 gnd.n5808 gnd.t17 11.1535
R18553 gnd.t116 gnd.n2920 11.1535
R18554 gnd.n3261 gnd.t38 11.1535
R18555 gnd.n3519 gnd.t55 11.1535
R18556 gnd.t46 gnd.n3767 11.1535
R18557 gnd.t234 gnd.n2031 11.1535
R18558 gnd.t159 gnd.n102 11.1535
R18559 gnd.n3462 gnd.n1535 10.8348
R18560 gnd.n3500 gnd.t62 10.8348
R18561 gnd.n3648 gnd.n3647 10.8348
R18562 gnd.n3647 gnd.n2232 10.8348
R18563 gnd.n3779 gnd.t21 10.8348
R18564 gnd.n3809 gnd.n2148 10.8348
R18565 gnd.n4410 gnd.n4407 10.6672
R18566 gnd.n7497 gnd.n315 10.6672
R18567 gnd.n4979 gnd.n4976 10.6672
R18568 gnd.n2547 gnd.n2445 10.6672
R18569 gnd.n4057 gnd.n4056 10.6151
R18570 gnd.n4056 gnd.n4053 10.6151
R18571 gnd.n4051 gnd.n4048 10.6151
R18572 gnd.n4048 gnd.n4047 10.6151
R18573 gnd.n4047 gnd.n4044 10.6151
R18574 gnd.n4044 gnd.n4043 10.6151
R18575 gnd.n4043 gnd.n4040 10.6151
R18576 gnd.n4040 gnd.n4039 10.6151
R18577 gnd.n4039 gnd.n4036 10.6151
R18578 gnd.n4036 gnd.n4035 10.6151
R18579 gnd.n4035 gnd.n4032 10.6151
R18580 gnd.n4032 gnd.n4031 10.6151
R18581 gnd.n4031 gnd.n4028 10.6151
R18582 gnd.n4028 gnd.n4027 10.6151
R18583 gnd.n4027 gnd.n4024 10.6151
R18584 gnd.n4024 gnd.n4023 10.6151
R18585 gnd.n4023 gnd.n4020 10.6151
R18586 gnd.n4020 gnd.n4019 10.6151
R18587 gnd.n4019 gnd.n4016 10.6151
R18588 gnd.n4016 gnd.n4015 10.6151
R18589 gnd.n4015 gnd.n4012 10.6151
R18590 gnd.n4012 gnd.n4011 10.6151
R18591 gnd.n4011 gnd.n4008 10.6151
R18592 gnd.n4008 gnd.n4007 10.6151
R18593 gnd.n4007 gnd.n4004 10.6151
R18594 gnd.n4004 gnd.n4003 10.6151
R18595 gnd.n4003 gnd.n4000 10.6151
R18596 gnd.n4000 gnd.n3999 10.6151
R18597 gnd.n3999 gnd.n3996 10.6151
R18598 gnd.n3996 gnd.n3995 10.6151
R18599 gnd.n3412 gnd.n3411 10.6151
R18600 gnd.n3411 gnd.n3410 10.6151
R18601 gnd.n3410 gnd.n3372 10.6151
R18602 gnd.n3401 gnd.n3372 10.6151
R18603 gnd.n3401 gnd.n3400 10.6151
R18604 gnd.n3400 gnd.n3399 10.6151
R18605 gnd.n3399 gnd.n3397 10.6151
R18606 gnd.n3397 gnd.n3396 10.6151
R18607 gnd.n3396 gnd.n3373 10.6151
R18608 gnd.n3387 gnd.n3373 10.6151
R18609 gnd.n3387 gnd.n3386 10.6151
R18610 gnd.n3386 gnd.n3385 10.6151
R18611 gnd.n3385 gnd.n3381 10.6151
R18612 gnd.n3381 gnd.n3380 10.6151
R18613 gnd.n3380 gnd.n3378 10.6151
R18614 gnd.n3378 gnd.n3377 10.6151
R18615 gnd.n3377 gnd.n3374 10.6151
R18616 gnd.n3374 gnd.n2319 10.6151
R18617 gnd.n3473 gnd.n2319 10.6151
R18618 gnd.n3474 gnd.n3473 10.6151
R18619 gnd.n3475 gnd.n3474 10.6151
R18620 gnd.n3475 gnd.n2305 10.6151
R18621 gnd.n3521 gnd.n2305 10.6151
R18622 gnd.n3522 gnd.n3521 10.6151
R18623 gnd.n3524 gnd.n3522 10.6151
R18624 gnd.n3524 gnd.n3523 10.6151
R18625 gnd.n3523 gnd.n2290 10.6151
R18626 gnd.n3552 gnd.n2290 10.6151
R18627 gnd.n3552 gnd.n3551 10.6151
R18628 gnd.n3551 gnd.n3550 10.6151
R18629 gnd.n3550 gnd.n3549 10.6151
R18630 gnd.n3549 gnd.n2270 10.6151
R18631 gnd.n3576 gnd.n2270 10.6151
R18632 gnd.n3577 gnd.n3576 10.6151
R18633 gnd.n3579 gnd.n3577 10.6151
R18634 gnd.n3580 gnd.n3579 10.6151
R18635 gnd.n3581 gnd.n3580 10.6151
R18636 gnd.n3581 gnd.n2246 10.6151
R18637 gnd.n3615 gnd.n2246 10.6151
R18638 gnd.n3616 gnd.n3615 10.6151
R18639 gnd.n3618 gnd.n3616 10.6151
R18640 gnd.n3619 gnd.n3618 10.6151
R18641 gnd.n3621 gnd.n3619 10.6151
R18642 gnd.n3621 gnd.n3620 10.6151
R18643 gnd.n3620 gnd.n2216 10.6151
R18644 gnd.n3675 gnd.n2216 10.6151
R18645 gnd.n3676 gnd.n3675 10.6151
R18646 gnd.n3678 gnd.n3676 10.6151
R18647 gnd.n3678 gnd.n3677 10.6151
R18648 gnd.n3677 gnd.n2196 10.6151
R18649 gnd.n3710 gnd.n2196 10.6151
R18650 gnd.n3711 gnd.n3710 10.6151
R18651 gnd.n3747 gnd.n3711 10.6151
R18652 gnd.n3747 gnd.n3746 10.6151
R18653 gnd.n3746 gnd.n3745 10.6151
R18654 gnd.n3745 gnd.n3742 10.6151
R18655 gnd.n3742 gnd.n3741 10.6151
R18656 gnd.n3741 gnd.n3740 10.6151
R18657 gnd.n3740 gnd.n3739 10.6151
R18658 gnd.n3739 gnd.n3738 10.6151
R18659 gnd.n3738 gnd.n3712 10.6151
R18660 gnd.n3732 gnd.n3712 10.6151
R18661 gnd.n3732 gnd.n3731 10.6151
R18662 gnd.n3731 gnd.n3730 10.6151
R18663 gnd.n3730 gnd.n3729 10.6151
R18664 gnd.n3729 gnd.n3728 10.6151
R18665 gnd.n3728 gnd.n3724 10.6151
R18666 gnd.n3724 gnd.n3723 10.6151
R18667 gnd.n3723 gnd.n3721 10.6151
R18668 gnd.n3721 gnd.n3720 10.6151
R18669 gnd.n3720 gnd.n3718 10.6151
R18670 gnd.n3718 gnd.n3717 10.6151
R18671 gnd.n3717 gnd.n2113 10.6151
R18672 gnd.n3870 gnd.n2113 10.6151
R18673 gnd.n3871 gnd.n3870 10.6151
R18674 gnd.n3878 gnd.n3871 10.6151
R18675 gnd.n3878 gnd.n3877 10.6151
R18676 gnd.n3877 gnd.n3876 10.6151
R18677 gnd.n3876 gnd.n3873 10.6151
R18678 gnd.n3873 gnd.n3872 10.6151
R18679 gnd.n3872 gnd.n2089 10.6151
R18680 gnd.n3310 gnd.n1429 10.6151
R18681 gnd.n3313 gnd.n3310 10.6151
R18682 gnd.n3318 gnd.n3315 10.6151
R18683 gnd.n3319 gnd.n3318 10.6151
R18684 gnd.n3322 gnd.n3319 10.6151
R18685 gnd.n3323 gnd.n3322 10.6151
R18686 gnd.n3326 gnd.n3323 10.6151
R18687 gnd.n3327 gnd.n3326 10.6151
R18688 gnd.n3330 gnd.n3327 10.6151
R18689 gnd.n3331 gnd.n3330 10.6151
R18690 gnd.n3334 gnd.n3331 10.6151
R18691 gnd.n3335 gnd.n3334 10.6151
R18692 gnd.n3338 gnd.n3335 10.6151
R18693 gnd.n3339 gnd.n3338 10.6151
R18694 gnd.n3342 gnd.n3339 10.6151
R18695 gnd.n3343 gnd.n3342 10.6151
R18696 gnd.n3346 gnd.n3343 10.6151
R18697 gnd.n3347 gnd.n3346 10.6151
R18698 gnd.n3350 gnd.n3347 10.6151
R18699 gnd.n3351 gnd.n3350 10.6151
R18700 gnd.n3354 gnd.n3351 10.6151
R18701 gnd.n3355 gnd.n3354 10.6151
R18702 gnd.n3358 gnd.n3355 10.6151
R18703 gnd.n3359 gnd.n3358 10.6151
R18704 gnd.n3362 gnd.n3359 10.6151
R18705 gnd.n3363 gnd.n3362 10.6151
R18706 gnd.n3366 gnd.n3363 10.6151
R18707 gnd.n3367 gnd.n3366 10.6151
R18708 gnd.n3370 gnd.n3367 10.6151
R18709 gnd.n3371 gnd.n3370 10.6151
R18710 gnd.n4776 gnd.n4775 10.6151
R18711 gnd.n4775 gnd.n4774 10.6151
R18712 gnd.n4774 gnd.n4773 10.6151
R18713 gnd.n4773 gnd.n4771 10.6151
R18714 gnd.n4771 gnd.n4768 10.6151
R18715 gnd.n4768 gnd.n4767 10.6151
R18716 gnd.n4767 gnd.n4764 10.6151
R18717 gnd.n4764 gnd.n4763 10.6151
R18718 gnd.n4763 gnd.n4760 10.6151
R18719 gnd.n4760 gnd.n4759 10.6151
R18720 gnd.n4759 gnd.n4756 10.6151
R18721 gnd.n4756 gnd.n4755 10.6151
R18722 gnd.n4755 gnd.n4752 10.6151
R18723 gnd.n4752 gnd.n4751 10.6151
R18724 gnd.n4751 gnd.n4748 10.6151
R18725 gnd.n4748 gnd.n4747 10.6151
R18726 gnd.n4747 gnd.n4744 10.6151
R18727 gnd.n4744 gnd.n4743 10.6151
R18728 gnd.n4743 gnd.n4740 10.6151
R18729 gnd.n4740 gnd.n4739 10.6151
R18730 gnd.n4739 gnd.n4736 10.6151
R18731 gnd.n4736 gnd.n4735 10.6151
R18732 gnd.n4735 gnd.n4732 10.6151
R18733 gnd.n4732 gnd.n4731 10.6151
R18734 gnd.n4731 gnd.n4728 10.6151
R18735 gnd.n4728 gnd.n4727 10.6151
R18736 gnd.n4727 gnd.n4724 10.6151
R18737 gnd.n4724 gnd.n4723 10.6151
R18738 gnd.n4720 gnd.n4719 10.6151
R18739 gnd.n4719 gnd.n1430 10.6151
R18740 gnd.n3988 gnd.n3987 10.6151
R18741 gnd.n3987 gnd.n3984 10.6151
R18742 gnd.n3984 gnd.n3983 10.6151
R18743 gnd.n3983 gnd.n3980 10.6151
R18744 gnd.n3980 gnd.n3979 10.6151
R18745 gnd.n3979 gnd.n3976 10.6151
R18746 gnd.n3976 gnd.n3975 10.6151
R18747 gnd.n3975 gnd.n3972 10.6151
R18748 gnd.n3972 gnd.n3971 10.6151
R18749 gnd.n3971 gnd.n3968 10.6151
R18750 gnd.n3968 gnd.n3967 10.6151
R18751 gnd.n3967 gnd.n3964 10.6151
R18752 gnd.n3964 gnd.n3963 10.6151
R18753 gnd.n3963 gnd.n3960 10.6151
R18754 gnd.n3960 gnd.n3959 10.6151
R18755 gnd.n3959 gnd.n3956 10.6151
R18756 gnd.n3956 gnd.n3955 10.6151
R18757 gnd.n3955 gnd.n3952 10.6151
R18758 gnd.n3952 gnd.n3951 10.6151
R18759 gnd.n3951 gnd.n3948 10.6151
R18760 gnd.n3948 gnd.n3947 10.6151
R18761 gnd.n3947 gnd.n3944 10.6151
R18762 gnd.n3944 gnd.n3943 10.6151
R18763 gnd.n3943 gnd.n3940 10.6151
R18764 gnd.n3940 gnd.n3939 10.6151
R18765 gnd.n3939 gnd.n3936 10.6151
R18766 gnd.n3936 gnd.n3935 10.6151
R18767 gnd.n3935 gnd.n3932 10.6151
R18768 gnd.n3930 gnd.n3927 10.6151
R18769 gnd.n3927 gnd.n3926 10.6151
R18770 gnd.n4712 gnd.n4711 10.6151
R18771 gnd.n4711 gnd.n1489 10.6151
R18772 gnd.n3404 gnd.n1489 10.6151
R18773 gnd.n3404 gnd.n1505 10.6151
R18774 gnd.n4699 gnd.n1505 10.6151
R18775 gnd.n4699 gnd.n4698 10.6151
R18776 gnd.n4698 gnd.n4697 10.6151
R18777 gnd.n4697 gnd.n1506 10.6151
R18778 gnd.n3391 gnd.n1506 10.6151
R18779 gnd.n3391 gnd.n1522 10.6151
R18780 gnd.n4685 gnd.n1522 10.6151
R18781 gnd.n4685 gnd.n4684 10.6151
R18782 gnd.n4684 gnd.n4683 10.6151
R18783 gnd.n4683 gnd.n1523 10.6151
R18784 gnd.n2323 gnd.n1523 10.6151
R18785 gnd.n3466 gnd.n2323 10.6151
R18786 gnd.n3467 gnd.n3466 10.6151
R18787 gnd.n3468 gnd.n3467 10.6151
R18788 gnd.n3468 gnd.n2318 10.6151
R18789 gnd.n3505 gnd.n2318 10.6151
R18790 gnd.n3505 gnd.n3504 10.6151
R18791 gnd.n3504 gnd.n3503 10.6151
R18792 gnd.n3503 gnd.n2301 10.6151
R18793 gnd.n3531 gnd.n2301 10.6151
R18794 gnd.n3532 gnd.n3531 10.6151
R18795 gnd.n3533 gnd.n3532 10.6151
R18796 gnd.n3533 gnd.n2284 10.6151
R18797 gnd.n3556 gnd.n2284 10.6151
R18798 gnd.n3557 gnd.n3556 10.6151
R18799 gnd.n3561 gnd.n3557 10.6151
R18800 gnd.n3561 gnd.n3560 10.6151
R18801 gnd.n3560 gnd.n3559 10.6151
R18802 gnd.n3559 gnd.n2260 10.6151
R18803 gnd.n3595 gnd.n2260 10.6151
R18804 gnd.n3596 gnd.n3595 10.6151
R18805 gnd.n3600 gnd.n3596 10.6151
R18806 gnd.n3600 gnd.n3599 10.6151
R18807 gnd.n3599 gnd.n3598 10.6151
R18808 gnd.n3598 gnd.n2237 10.6151
R18809 gnd.n3650 gnd.n2237 10.6151
R18810 gnd.n3651 gnd.n3650 10.6151
R18811 gnd.n3652 gnd.n3651 10.6151
R18812 gnd.n3652 gnd.n2222 10.6151
R18813 gnd.n3668 gnd.n2222 10.6151
R18814 gnd.n3669 gnd.n3668 10.6151
R18815 gnd.n3671 gnd.n3669 10.6151
R18816 gnd.n3671 gnd.n3670 10.6151
R18817 gnd.n3670 gnd.n2203 10.6151
R18818 gnd.n3696 gnd.n2203 10.6151
R18819 gnd.n3697 gnd.n3696 10.6151
R18820 gnd.n3706 gnd.n3697 10.6151
R18821 gnd.n3706 gnd.n3705 10.6151
R18822 gnd.n3705 gnd.n3704 10.6151
R18823 gnd.n3704 gnd.n3703 10.6151
R18824 gnd.n3703 gnd.n3698 10.6151
R18825 gnd.n3698 gnd.n2173 10.6151
R18826 gnd.n3771 gnd.n2173 10.6151
R18827 gnd.n3772 gnd.n3771 10.6151
R18828 gnd.n3776 gnd.n3772 10.6151
R18829 gnd.n3776 gnd.n3775 10.6151
R18830 gnd.n3775 gnd.n3774 10.6151
R18831 gnd.n3774 gnd.n2150 10.6151
R18832 gnd.n3805 gnd.n2150 10.6151
R18833 gnd.n3806 gnd.n3805 10.6151
R18834 gnd.n3807 gnd.n3806 10.6151
R18835 gnd.n3807 gnd.n2136 10.6151
R18836 gnd.n3821 gnd.n2136 10.6151
R18837 gnd.n3822 gnd.n3821 10.6151
R18838 gnd.n3823 gnd.n3822 10.6151
R18839 gnd.n3823 gnd.n2124 10.6151
R18840 gnd.n3856 gnd.n2124 10.6151
R18841 gnd.n3856 gnd.n3855 10.6151
R18842 gnd.n3855 gnd.n3854 10.6151
R18843 gnd.n3854 gnd.n2108 10.6151
R18844 gnd.n3885 gnd.n2108 10.6151
R18845 gnd.n3886 gnd.n3885 10.6151
R18846 gnd.n3887 gnd.n3886 10.6151
R18847 gnd.n3887 gnd.n2094 10.6151
R18848 gnd.n3901 gnd.n2094 10.6151
R18849 gnd.n3902 gnd.n3901 10.6151
R18850 gnd.n3990 gnd.n3902 10.6151
R18851 gnd.n5480 gnd.t236 10.5161
R18852 gnd.n6366 gnd.t50 10.5161
R18853 gnd.n6373 gnd.t23 10.5161
R18854 gnd.n2995 gnd.t163 10.5161
R18855 gnd.n4674 gnd.t8 10.5161
R18856 gnd.n3810 gnd.t10 10.5161
R18857 gnd.n1909 gnd.t140 10.5161
R18858 gnd.n6328 gnd.n6312 10.4732
R18859 gnd.n6296 gnd.n6280 10.4732
R18860 gnd.n6264 gnd.n6248 10.4732
R18861 gnd.n6233 gnd.n6217 10.4732
R18862 gnd.n6201 gnd.n6185 10.4732
R18863 gnd.n6169 gnd.n6153 10.4732
R18864 gnd.n6137 gnd.n6121 10.4732
R18865 gnd.n6106 gnd.n6090 10.4732
R18866 gnd.n4702 gnd.t241 10.1975
R18867 gnd.n3493 gnd.n3492 10.1975
R18868 gnd.n3564 gnd.n2278 10.1975
R18869 gnd.n2201 gnd.n2200 10.1975
R18870 gnd.n3701 gnd.n3700 10.1975
R18871 gnd.n3890 gnd.t277 10.1975
R18872 gnd.n3890 gnd.n3889 10.1975
R18873 gnd.n3899 gnd.n3898 10.1975
R18874 gnd.n6065 gnd.t30 9.87883
R18875 gnd.n3056 gnd.t82 9.87883
R18876 gnd.n3584 gnd.t43 9.87883
R18877 gnd.n3624 gnd.t60 9.87883
R18878 gnd.n4224 gnd.t110 9.87883
R18879 gnd.n6332 gnd.n6331 9.69747
R18880 gnd.n6300 gnd.n6299 9.69747
R18881 gnd.n6268 gnd.n6267 9.69747
R18882 gnd.n6237 gnd.n6236 9.69747
R18883 gnd.n6205 gnd.n6204 9.69747
R18884 gnd.n6173 gnd.n6172 9.69747
R18885 gnd.n6141 gnd.n6140 9.69747
R18886 gnd.n6110 gnd.n6109 9.69747
R18887 gnd.n4681 gnd.n1525 9.56018
R18888 gnd.n3471 gnd.n3470 9.56018
R18889 gnd.n3584 gnd.n2248 9.56018
R18890 gnd.n3624 gnd.n3623 9.56018
R18891 gnd.n3803 gnd.n2152 9.56018
R18892 gnd.n2140 gnd.n2133 9.56018
R18893 gnd.n3852 gnd.t295 9.56018
R18894 gnd.n6338 gnd.n6337 9.45567
R18895 gnd.n6306 gnd.n6305 9.45567
R18896 gnd.n6274 gnd.n6273 9.45567
R18897 gnd.n6243 gnd.n6242 9.45567
R18898 gnd.n6211 gnd.n6210 9.45567
R18899 gnd.n6179 gnd.n6178 9.45567
R18900 gnd.n6147 gnd.n6146 9.45567
R18901 gnd.n6116 gnd.n6115 9.45567
R18902 gnd.n4447 gnd.n4446 9.30959
R18903 gnd.n7531 gnd.n279 9.30959
R18904 gnd.n5016 gnd.n5015 9.30959
R18905 gnd.n2503 gnd.n2467 9.30959
R18906 gnd.n6337 gnd.n6336 9.3005
R18907 gnd.n6310 gnd.n6309 9.3005
R18908 gnd.n6331 gnd.n6330 9.3005
R18909 gnd.n6329 gnd.n6328 9.3005
R18910 gnd.n6314 gnd.n6313 9.3005
R18911 gnd.n6323 gnd.n6322 9.3005
R18912 gnd.n6321 gnd.n6320 9.3005
R18913 gnd.n6305 gnd.n6304 9.3005
R18914 gnd.n6278 gnd.n6277 9.3005
R18915 gnd.n6299 gnd.n6298 9.3005
R18916 gnd.n6297 gnd.n6296 9.3005
R18917 gnd.n6282 gnd.n6281 9.3005
R18918 gnd.n6291 gnd.n6290 9.3005
R18919 gnd.n6289 gnd.n6288 9.3005
R18920 gnd.n6273 gnd.n6272 9.3005
R18921 gnd.n6246 gnd.n6245 9.3005
R18922 gnd.n6267 gnd.n6266 9.3005
R18923 gnd.n6265 gnd.n6264 9.3005
R18924 gnd.n6250 gnd.n6249 9.3005
R18925 gnd.n6259 gnd.n6258 9.3005
R18926 gnd.n6257 gnd.n6256 9.3005
R18927 gnd.n6242 gnd.n6241 9.3005
R18928 gnd.n6215 gnd.n6214 9.3005
R18929 gnd.n6236 gnd.n6235 9.3005
R18930 gnd.n6234 gnd.n6233 9.3005
R18931 gnd.n6219 gnd.n6218 9.3005
R18932 gnd.n6228 gnd.n6227 9.3005
R18933 gnd.n6226 gnd.n6225 9.3005
R18934 gnd.n6210 gnd.n6209 9.3005
R18935 gnd.n6183 gnd.n6182 9.3005
R18936 gnd.n6204 gnd.n6203 9.3005
R18937 gnd.n6202 gnd.n6201 9.3005
R18938 gnd.n6187 gnd.n6186 9.3005
R18939 gnd.n6196 gnd.n6195 9.3005
R18940 gnd.n6194 gnd.n6193 9.3005
R18941 gnd.n6178 gnd.n6177 9.3005
R18942 gnd.n6151 gnd.n6150 9.3005
R18943 gnd.n6172 gnd.n6171 9.3005
R18944 gnd.n6170 gnd.n6169 9.3005
R18945 gnd.n6155 gnd.n6154 9.3005
R18946 gnd.n6164 gnd.n6163 9.3005
R18947 gnd.n6162 gnd.n6161 9.3005
R18948 gnd.n6146 gnd.n6145 9.3005
R18949 gnd.n6119 gnd.n6118 9.3005
R18950 gnd.n6140 gnd.n6139 9.3005
R18951 gnd.n6138 gnd.n6137 9.3005
R18952 gnd.n6123 gnd.n6122 9.3005
R18953 gnd.n6132 gnd.n6131 9.3005
R18954 gnd.n6130 gnd.n6129 9.3005
R18955 gnd.n6115 gnd.n6114 9.3005
R18956 gnd.n6088 gnd.n6087 9.3005
R18957 gnd.n6109 gnd.n6108 9.3005
R18958 gnd.n6107 gnd.n6106 9.3005
R18959 gnd.n6092 gnd.n6091 9.3005
R18960 gnd.n6101 gnd.n6100 9.3005
R18961 gnd.n6099 gnd.n6098 9.3005
R18962 gnd.n6467 gnd.n5099 9.3005
R18963 gnd.n6466 gnd.n5101 9.3005
R18964 gnd.n5105 gnd.n5102 9.3005
R18965 gnd.n6461 gnd.n5106 9.3005
R18966 gnd.n6460 gnd.n5107 9.3005
R18967 gnd.n6459 gnd.n5108 9.3005
R18968 gnd.n5112 gnd.n5109 9.3005
R18969 gnd.n6454 gnd.n5113 9.3005
R18970 gnd.n6453 gnd.n5114 9.3005
R18971 gnd.n6452 gnd.n5115 9.3005
R18972 gnd.n5119 gnd.n5116 9.3005
R18973 gnd.n6447 gnd.n5120 9.3005
R18974 gnd.n6446 gnd.n5121 9.3005
R18975 gnd.n6445 gnd.n5122 9.3005
R18976 gnd.n5127 gnd.n5125 9.3005
R18977 gnd.n6440 gnd.n6439 9.3005
R18978 gnd.n6469 gnd.n6468 9.3005
R18979 gnd.n5747 gnd.n5746 9.3005
R18980 gnd.n5748 gnd.n5450 9.3005
R18981 gnd.n5750 gnd.n5749 9.3005
R18982 gnd.n5431 gnd.n5430 9.3005
R18983 gnd.n5777 gnd.n5776 9.3005
R18984 gnd.n5778 gnd.n5429 9.3005
R18985 gnd.n5782 gnd.n5779 9.3005
R18986 gnd.n5781 gnd.n5780 9.3005
R18987 gnd.n5405 gnd.n5404 9.3005
R18988 gnd.n5811 gnd.n5810 9.3005
R18989 gnd.n5812 gnd.n5403 9.3005
R18990 gnd.n5819 gnd.n5813 9.3005
R18991 gnd.n5818 gnd.n5814 9.3005
R18992 gnd.n5817 gnd.n5815 9.3005
R18993 gnd.n5372 gnd.n5371 9.3005
R18994 gnd.n5872 gnd.n5871 9.3005
R18995 gnd.n5873 gnd.n5370 9.3005
R18996 gnd.n5877 gnd.n5874 9.3005
R18997 gnd.n5876 gnd.n5875 9.3005
R18998 gnd.n5345 gnd.n5344 9.3005
R18999 gnd.n5912 gnd.n5911 9.3005
R19000 gnd.n5913 gnd.n5343 9.3005
R19001 gnd.n5917 gnd.n5914 9.3005
R19002 gnd.n5916 gnd.n5915 9.3005
R19003 gnd.n5254 gnd.n5253 9.3005
R19004 gnd.n5957 gnd.n5956 9.3005
R19005 gnd.n5958 gnd.n5252 9.3005
R19006 gnd.n5962 gnd.n5959 9.3005
R19007 gnd.n5961 gnd.n5960 9.3005
R19008 gnd.n5226 gnd.n5225 9.3005
R19009 gnd.n5996 gnd.n5995 9.3005
R19010 gnd.n5997 gnd.n5224 9.3005
R19011 gnd.n6004 gnd.n5998 9.3005
R19012 gnd.n6003 gnd.n5999 9.3005
R19013 gnd.n6002 gnd.n6000 9.3005
R19014 gnd.n5196 gnd.n5195 9.3005
R19015 gnd.n6053 gnd.n6052 9.3005
R19016 gnd.n6054 gnd.n5194 9.3005
R19017 gnd.n6062 gnd.n6055 9.3005
R19018 gnd.n6061 gnd.n6056 9.3005
R19019 gnd.n6060 gnd.n6058 9.3005
R19020 gnd.n6057 gnd.n984 9.3005
R19021 gnd.n6499 gnd.n985 9.3005
R19022 gnd.n6498 gnd.n986 9.3005
R19023 gnd.n6497 gnd.n987 9.3005
R19024 gnd.n1009 gnd.n988 9.3005
R19025 gnd.n1010 gnd.n1008 9.3005
R19026 gnd.n6485 gnd.n1011 9.3005
R19027 gnd.n6484 gnd.n1012 9.3005
R19028 gnd.n6483 gnd.n1013 9.3005
R19029 gnd.n5097 gnd.n1014 9.3005
R19030 gnd.n5098 gnd.n5096 9.3005
R19031 gnd.n6471 gnd.n6470 9.3005
R19032 gnd.n5452 gnd.n5451 9.3005
R19033 gnd.n5692 gnd.n5691 9.3005
R19034 gnd.n5695 gnd.n5687 9.3005
R19035 gnd.n5696 gnd.n5686 9.3005
R19036 gnd.n5699 gnd.n5685 9.3005
R19037 gnd.n5700 gnd.n5684 9.3005
R19038 gnd.n5703 gnd.n5683 9.3005
R19039 gnd.n5704 gnd.n5682 9.3005
R19040 gnd.n5707 gnd.n5681 9.3005
R19041 gnd.n5708 gnd.n5680 9.3005
R19042 gnd.n5711 gnd.n5679 9.3005
R19043 gnd.n5712 gnd.n5678 9.3005
R19044 gnd.n5715 gnd.n5677 9.3005
R19045 gnd.n5717 gnd.n5676 9.3005
R19046 gnd.n5718 gnd.n5675 9.3005
R19047 gnd.n5719 gnd.n5674 9.3005
R19048 gnd.n5720 gnd.n5673 9.3005
R19049 gnd.n5688 gnd.n5469 9.3005
R19050 gnd.n5737 gnd.n5460 9.3005
R19051 gnd.n5739 gnd.n5738 9.3005
R19052 gnd.n5447 gnd.n5442 9.3005
R19053 gnd.n5760 gnd.n5441 9.3005
R19054 gnd.n5763 gnd.n5762 9.3005
R19055 gnd.n5765 gnd.n5764 9.3005
R19056 gnd.n5768 gnd.n5424 9.3005
R19057 gnd.n5766 gnd.n5422 9.3005
R19058 gnd.n5788 gnd.n5420 9.3005
R19059 gnd.n5792 gnd.n5791 9.3005
R19060 gnd.n5790 gnd.n5395 9.3005
R19061 gnd.n5826 gnd.n5394 9.3005
R19062 gnd.n5829 gnd.n5828 9.3005
R19063 gnd.n5392 gnd.n5391 9.3005
R19064 gnd.n5835 gnd.n5389 9.3005
R19065 gnd.n5837 gnd.n5836 9.3005
R19066 gnd.n5363 gnd.n5362 9.3005
R19067 gnd.n5886 gnd.n5885 9.3005
R19068 gnd.n5887 gnd.n5356 9.3005
R19069 gnd.n5895 gnd.n5355 9.3005
R19070 gnd.n5898 gnd.n5897 9.3005
R19071 gnd.n5900 gnd.n5899 9.3005
R19072 gnd.n5903 gnd.n5338 9.3005
R19073 gnd.n5901 gnd.n5336 9.3005
R19074 gnd.n5923 gnd.n5334 9.3005
R19075 gnd.n5925 gnd.n5924 9.3005
R19076 gnd.n5244 gnd.n5243 9.3005
R19077 gnd.n5971 gnd.n5970 9.3005
R19078 gnd.n5972 gnd.n5237 9.3005
R19079 gnd.n5980 gnd.n5236 9.3005
R19080 gnd.n5983 gnd.n5982 9.3005
R19081 gnd.n5985 gnd.n5984 9.3005
R19082 gnd.n5987 gnd.n5219 9.3005
R19083 gnd.n5217 gnd.n5215 9.3005
R19084 gnd.n6012 gnd.n6011 9.3005
R19085 gnd.n5201 gnd.n5200 9.3005
R19086 gnd.n6045 gnd.n6044 9.3005
R19087 gnd.n6046 gnd.n5187 9.3005
R19088 gnd.n6069 gnd.n5186 9.3005
R19089 gnd.n6072 gnd.n6071 9.3005
R19090 gnd.n5183 gnd.n5182 9.3005
R19091 gnd.n6076 gnd.n5184 9.3005
R19092 gnd.n6078 gnd.n6077 9.3005
R19093 gnd.n6363 gnd.n6080 9.3005
R19094 gnd.n6362 gnd.n6082 9.3005
R19095 gnd.n6361 gnd.n6083 9.3005
R19096 gnd.n6358 gnd.n6084 9.3005
R19097 gnd.n6357 gnd.n6085 9.3005
R19098 gnd.n6356 gnd.n6343 9.3005
R19099 gnd.n6353 gnd.n6345 9.3005
R19100 gnd.n6352 gnd.n6346 9.3005
R19101 gnd.n6349 gnd.n6347 9.3005
R19102 gnd.n6348 gnd.n5128 9.3005
R19103 gnd.n5736 gnd.n5463 9.3005
R19104 gnd.n6435 gnd.n5129 9.3005
R19105 gnd.n6434 gnd.n5131 9.3005
R19106 gnd.n5135 gnd.n5132 9.3005
R19107 gnd.n6429 gnd.n5136 9.3005
R19108 gnd.n6428 gnd.n5137 9.3005
R19109 gnd.n6427 gnd.n5138 9.3005
R19110 gnd.n5142 gnd.n5139 9.3005
R19111 gnd.n6422 gnd.n5143 9.3005
R19112 gnd.n6421 gnd.n5144 9.3005
R19113 gnd.n6420 gnd.n5145 9.3005
R19114 gnd.n5149 gnd.n5146 9.3005
R19115 gnd.n6415 gnd.n5150 9.3005
R19116 gnd.n6414 gnd.n5151 9.3005
R19117 gnd.n6413 gnd.n5152 9.3005
R19118 gnd.n5156 gnd.n5153 9.3005
R19119 gnd.n6408 gnd.n5157 9.3005
R19120 gnd.n6407 gnd.n5158 9.3005
R19121 gnd.n6406 gnd.n5159 9.3005
R19122 gnd.n5163 gnd.n5160 9.3005
R19123 gnd.n6401 gnd.n5164 9.3005
R19124 gnd.n6400 gnd.n5165 9.3005
R19125 gnd.n6399 gnd.n5166 9.3005
R19126 gnd.n5173 gnd.n5171 9.3005
R19127 gnd.n6394 gnd.n5174 9.3005
R19128 gnd.n6393 gnd.n5175 9.3005
R19129 gnd.n6392 gnd.n6389 9.3005
R19130 gnd.n6437 gnd.n6436 9.3005
R19131 gnd.n5933 gnd.n5932 9.3005
R19132 gnd.n5934 gnd.n5260 9.3005
R19133 gnd.n5951 gnd.n5935 9.3005
R19134 gnd.n5950 gnd.n5936 9.3005
R19135 gnd.n5949 gnd.n5937 9.3005
R19136 gnd.n5947 gnd.n5938 9.3005
R19137 gnd.n5946 gnd.n5939 9.3005
R19138 gnd.n5944 gnd.n5940 9.3005
R19139 gnd.n5943 gnd.n5941 9.3005
R19140 gnd.n5208 gnd.n5207 9.3005
R19141 gnd.n6019 gnd.n6018 9.3005
R19142 gnd.n6020 gnd.n5206 9.3005
R19143 gnd.n6037 gnd.n6021 9.3005
R19144 gnd.n6036 gnd.n6022 9.3005
R19145 gnd.n6035 gnd.n6023 9.3005
R19146 gnd.n6034 gnd.n6024 9.3005
R19147 gnd.n6032 gnd.n6025 9.3005
R19148 gnd.n6031 gnd.n6026 9.3005
R19149 gnd.n6028 gnd.n6027 9.3005
R19150 gnd.n5181 gnd.n5180 9.3005
R19151 gnd.n6370 gnd.n6369 9.3005
R19152 gnd.n6371 gnd.n5179 9.3005
R19153 gnd.n6375 gnd.n6372 9.3005
R19154 gnd.n6376 gnd.n5178 9.3005
R19155 gnd.n6380 gnd.n6379 9.3005
R19156 gnd.n6381 gnd.n5177 9.3005
R19157 gnd.n6383 gnd.n6382 9.3005
R19158 gnd.n6386 gnd.n5176 9.3005
R19159 gnd.n6388 gnd.n6387 9.3005
R19160 gnd.n5606 gnd.n5500 9.3005
R19161 gnd.n5608 gnd.n5607 9.3005
R19162 gnd.n5490 gnd.n5489 9.3005
R19163 gnd.n5621 gnd.n5620 9.3005
R19164 gnd.n5622 gnd.n5488 9.3005
R19165 gnd.n5624 gnd.n5623 9.3005
R19166 gnd.n5477 gnd.n5476 9.3005
R19167 gnd.n5637 gnd.n5636 9.3005
R19168 gnd.n5638 gnd.n5475 9.3005
R19169 gnd.n5662 gnd.n5639 9.3005
R19170 gnd.n5661 gnd.n5640 9.3005
R19171 gnd.n5660 gnd.n5641 9.3005
R19172 gnd.n5659 gnd.n5642 9.3005
R19173 gnd.n5657 gnd.n5643 9.3005
R19174 gnd.n5656 gnd.n5644 9.3005
R19175 gnd.n5654 gnd.n5645 9.3005
R19176 gnd.n5653 gnd.n5646 9.3005
R19177 gnd.n5651 gnd.n5647 9.3005
R19178 gnd.n5650 gnd.n5648 9.3005
R19179 gnd.n5412 gnd.n5411 9.3005
R19180 gnd.n5800 gnd.n5799 9.3005
R19181 gnd.n5801 gnd.n5410 9.3005
R19182 gnd.n5805 gnd.n5802 9.3005
R19183 gnd.n5804 gnd.n5803 9.3005
R19184 gnd.n5379 gnd.n5378 9.3005
R19185 gnd.n5847 gnd.n5846 9.3005
R19186 gnd.n5848 gnd.n5377 9.3005
R19187 gnd.n5850 gnd.n5849 9.3005
R19188 gnd.n5605 gnd.n5604 9.3005
R19189 gnd.n5545 gnd.n5544 9.3005
R19190 gnd.n5550 gnd.n5542 9.3005
R19191 gnd.n5551 gnd.n5541 9.3005
R19192 gnd.n5553 gnd.n5538 9.3005
R19193 gnd.n5537 gnd.n5535 9.3005
R19194 gnd.n5559 gnd.n5534 9.3005
R19195 gnd.n5560 gnd.n5533 9.3005
R19196 gnd.n5561 gnd.n5532 9.3005
R19197 gnd.n5531 gnd.n5529 9.3005
R19198 gnd.n5567 gnd.n5528 9.3005
R19199 gnd.n5568 gnd.n5527 9.3005
R19200 gnd.n5569 gnd.n5526 9.3005
R19201 gnd.n5525 gnd.n5523 9.3005
R19202 gnd.n5575 gnd.n5522 9.3005
R19203 gnd.n5576 gnd.n5521 9.3005
R19204 gnd.n5577 gnd.n5520 9.3005
R19205 gnd.n5519 gnd.n5517 9.3005
R19206 gnd.n5583 gnd.n5516 9.3005
R19207 gnd.n5584 gnd.n5515 9.3005
R19208 gnd.n5585 gnd.n5514 9.3005
R19209 gnd.n5513 gnd.n5511 9.3005
R19210 gnd.n5590 gnd.n5510 9.3005
R19211 gnd.n5591 gnd.n5509 9.3005
R19212 gnd.n5508 gnd.n5506 9.3005
R19213 gnd.n5596 gnd.n5505 9.3005
R19214 gnd.n5598 gnd.n5597 9.3005
R19215 gnd.n5543 gnd.n5501 9.3005
R19216 gnd.n5496 gnd.n5495 9.3005
R19217 gnd.n5613 gnd.n5612 9.3005
R19218 gnd.n5614 gnd.n5494 9.3005
R19219 gnd.n5616 gnd.n5615 9.3005
R19220 gnd.n5484 gnd.n5483 9.3005
R19221 gnd.n5629 gnd.n5628 9.3005
R19222 gnd.n5630 gnd.n5482 9.3005
R19223 gnd.n5632 gnd.n5631 9.3005
R19224 gnd.n5471 gnd.n5470 9.3005
R19225 gnd.n5727 gnd.n5726 9.3005
R19226 gnd.n5729 gnd.n5468 9.3005
R19227 gnd.n5731 gnd.n5730 9.3005
R19228 gnd.n5462 gnd.n5459 9.3005
R19229 gnd.n5741 gnd.n5740 9.3005
R19230 gnd.n5461 gnd.n5443 9.3005
R19231 gnd.n5759 gnd.n5758 9.3005
R19232 gnd.n5761 gnd.n5439 9.3005
R19233 gnd.n5771 gnd.n5440 9.3005
R19234 gnd.n5770 gnd.n5769 9.3005
R19235 gnd.n5767 gnd.n5418 9.3005
R19236 gnd.n5795 gnd.n5419 9.3005
R19237 gnd.n5794 gnd.n5793 9.3005
R19238 gnd.n5421 gnd.n5396 9.3005
R19239 gnd.n5825 gnd.n5824 9.3005
R19240 gnd.n5827 gnd.n5386 9.3005
R19241 gnd.n5842 gnd.n5387 9.3005
R19242 gnd.n5841 gnd.n5388 9.3005
R19243 gnd.n5840 gnd.n5838 9.3005
R19244 gnd.n5390 gnd.n5364 9.3005
R19245 gnd.n5883 gnd.n5882 9.3005
R19246 gnd.n5884 gnd.n5357 9.3005
R19247 gnd.n5894 gnd.n5893 9.3005
R19248 gnd.n5896 gnd.n5353 9.3005
R19249 gnd.n5906 gnd.n5354 9.3005
R19250 gnd.n5905 gnd.n5904 9.3005
R19251 gnd.n5902 gnd.n5332 9.3005
R19252 gnd.n5928 gnd.n5333 9.3005
R19253 gnd.n5927 gnd.n5926 9.3005
R19254 gnd.n5335 gnd.n5245 9.3005
R19255 gnd.n5968 gnd.n5967 9.3005
R19256 gnd.n5969 gnd.n5238 9.3005
R19257 gnd.n5979 gnd.n5978 9.3005
R19258 gnd.n5981 gnd.n5234 9.3005
R19259 gnd.n5990 gnd.n5235 9.3005
R19260 gnd.n5989 gnd.n5988 9.3005
R19261 gnd.n5986 gnd.n5214 9.3005
R19262 gnd.n6014 gnd.n6013 9.3005
R19263 gnd.n5216 gnd.n5202 9.3005
R19264 gnd.n6042 gnd.n6041 9.3005
R19265 gnd.n6043 gnd.n5188 9.3005
R19266 gnd.n6068 gnd.n6067 9.3005
R19267 gnd.n6070 gnd.n973 9.3005
R19268 gnd.n6506 gnd.n974 9.3005
R19269 gnd.n6505 gnd.n975 9.3005
R19270 gnd.n6504 gnd.n976 9.3005
R19271 gnd.n6079 gnd.n977 9.3005
R19272 gnd.n6081 gnd.n996 9.3005
R19273 gnd.n6492 gnd.n997 9.3005
R19274 gnd.n6491 gnd.n998 9.3005
R19275 gnd.n6490 gnd.n999 9.3005
R19276 gnd.n6342 gnd.n1000 9.3005
R19277 gnd.n6344 gnd.n1022 9.3005
R19278 gnd.n6478 gnd.n1023 9.3005
R19279 gnd.n6477 gnd.n1024 9.3005
R19280 gnd.n6476 gnd.n1025 9.3005
R19281 gnd.n5600 gnd.n5599 9.3005
R19282 gnd.n799 gnd.n798 9.3005
R19283 gnd.n6682 gnd.n6681 9.3005
R19284 gnd.n6683 gnd.n797 9.3005
R19285 gnd.n6685 gnd.n6684 9.3005
R19286 gnd.n793 gnd.n792 9.3005
R19287 gnd.n6692 gnd.n6691 9.3005
R19288 gnd.n6693 gnd.n791 9.3005
R19289 gnd.n6695 gnd.n6694 9.3005
R19290 gnd.n787 gnd.n786 9.3005
R19291 gnd.n6702 gnd.n6701 9.3005
R19292 gnd.n6703 gnd.n785 9.3005
R19293 gnd.n6705 gnd.n6704 9.3005
R19294 gnd.n781 gnd.n780 9.3005
R19295 gnd.n6712 gnd.n6711 9.3005
R19296 gnd.n6713 gnd.n779 9.3005
R19297 gnd.n6715 gnd.n6714 9.3005
R19298 gnd.n775 gnd.n774 9.3005
R19299 gnd.n6722 gnd.n6721 9.3005
R19300 gnd.n6723 gnd.n773 9.3005
R19301 gnd.n6725 gnd.n6724 9.3005
R19302 gnd.n769 gnd.n768 9.3005
R19303 gnd.n6732 gnd.n6731 9.3005
R19304 gnd.n6733 gnd.n767 9.3005
R19305 gnd.n6735 gnd.n6734 9.3005
R19306 gnd.n763 gnd.n762 9.3005
R19307 gnd.n6742 gnd.n6741 9.3005
R19308 gnd.n6743 gnd.n761 9.3005
R19309 gnd.n6745 gnd.n6744 9.3005
R19310 gnd.n757 gnd.n756 9.3005
R19311 gnd.n6752 gnd.n6751 9.3005
R19312 gnd.n6753 gnd.n755 9.3005
R19313 gnd.n6755 gnd.n6754 9.3005
R19314 gnd.n751 gnd.n750 9.3005
R19315 gnd.n6762 gnd.n6761 9.3005
R19316 gnd.n6763 gnd.n749 9.3005
R19317 gnd.n6765 gnd.n6764 9.3005
R19318 gnd.n745 gnd.n744 9.3005
R19319 gnd.n6772 gnd.n6771 9.3005
R19320 gnd.n6773 gnd.n743 9.3005
R19321 gnd.n6775 gnd.n6774 9.3005
R19322 gnd.n739 gnd.n738 9.3005
R19323 gnd.n6782 gnd.n6781 9.3005
R19324 gnd.n6783 gnd.n737 9.3005
R19325 gnd.n6785 gnd.n6784 9.3005
R19326 gnd.n733 gnd.n732 9.3005
R19327 gnd.n6792 gnd.n6791 9.3005
R19328 gnd.n6793 gnd.n731 9.3005
R19329 gnd.n6795 gnd.n6794 9.3005
R19330 gnd.n727 gnd.n726 9.3005
R19331 gnd.n6802 gnd.n6801 9.3005
R19332 gnd.n6803 gnd.n725 9.3005
R19333 gnd.n6805 gnd.n6804 9.3005
R19334 gnd.n721 gnd.n720 9.3005
R19335 gnd.n6812 gnd.n6811 9.3005
R19336 gnd.n6813 gnd.n719 9.3005
R19337 gnd.n6815 gnd.n6814 9.3005
R19338 gnd.n715 gnd.n714 9.3005
R19339 gnd.n6822 gnd.n6821 9.3005
R19340 gnd.n6823 gnd.n713 9.3005
R19341 gnd.n6825 gnd.n6824 9.3005
R19342 gnd.n709 gnd.n708 9.3005
R19343 gnd.n6832 gnd.n6831 9.3005
R19344 gnd.n6833 gnd.n707 9.3005
R19345 gnd.n6835 gnd.n6834 9.3005
R19346 gnd.n703 gnd.n702 9.3005
R19347 gnd.n6842 gnd.n6841 9.3005
R19348 gnd.n6843 gnd.n701 9.3005
R19349 gnd.n6845 gnd.n6844 9.3005
R19350 gnd.n697 gnd.n696 9.3005
R19351 gnd.n6852 gnd.n6851 9.3005
R19352 gnd.n6853 gnd.n695 9.3005
R19353 gnd.n6855 gnd.n6854 9.3005
R19354 gnd.n691 gnd.n690 9.3005
R19355 gnd.n6862 gnd.n6861 9.3005
R19356 gnd.n6863 gnd.n689 9.3005
R19357 gnd.n6865 gnd.n6864 9.3005
R19358 gnd.n685 gnd.n684 9.3005
R19359 gnd.n6872 gnd.n6871 9.3005
R19360 gnd.n6873 gnd.n683 9.3005
R19361 gnd.n6875 gnd.n6874 9.3005
R19362 gnd.n679 gnd.n678 9.3005
R19363 gnd.n6882 gnd.n6881 9.3005
R19364 gnd.n6883 gnd.n677 9.3005
R19365 gnd.n6885 gnd.n6884 9.3005
R19366 gnd.n673 gnd.n672 9.3005
R19367 gnd.n6892 gnd.n6891 9.3005
R19368 gnd.n6893 gnd.n671 9.3005
R19369 gnd.n6895 gnd.n6894 9.3005
R19370 gnd.n667 gnd.n666 9.3005
R19371 gnd.n6902 gnd.n6901 9.3005
R19372 gnd.n6903 gnd.n665 9.3005
R19373 gnd.n6905 gnd.n6904 9.3005
R19374 gnd.n661 gnd.n660 9.3005
R19375 gnd.n6912 gnd.n6911 9.3005
R19376 gnd.n6913 gnd.n659 9.3005
R19377 gnd.n6915 gnd.n6914 9.3005
R19378 gnd.n655 gnd.n654 9.3005
R19379 gnd.n6922 gnd.n6921 9.3005
R19380 gnd.n6923 gnd.n653 9.3005
R19381 gnd.n6925 gnd.n6924 9.3005
R19382 gnd.n649 gnd.n648 9.3005
R19383 gnd.n6932 gnd.n6931 9.3005
R19384 gnd.n6933 gnd.n647 9.3005
R19385 gnd.n6935 gnd.n6934 9.3005
R19386 gnd.n643 gnd.n642 9.3005
R19387 gnd.n6942 gnd.n6941 9.3005
R19388 gnd.n6943 gnd.n641 9.3005
R19389 gnd.n6945 gnd.n6944 9.3005
R19390 gnd.n637 gnd.n636 9.3005
R19391 gnd.n6952 gnd.n6951 9.3005
R19392 gnd.n6953 gnd.n635 9.3005
R19393 gnd.n6955 gnd.n6954 9.3005
R19394 gnd.n631 gnd.n630 9.3005
R19395 gnd.n6962 gnd.n6961 9.3005
R19396 gnd.n6963 gnd.n629 9.3005
R19397 gnd.n6965 gnd.n6964 9.3005
R19398 gnd.n625 gnd.n624 9.3005
R19399 gnd.n6972 gnd.n6971 9.3005
R19400 gnd.n6973 gnd.n623 9.3005
R19401 gnd.n6975 gnd.n6974 9.3005
R19402 gnd.n619 gnd.n618 9.3005
R19403 gnd.n6982 gnd.n6981 9.3005
R19404 gnd.n6983 gnd.n617 9.3005
R19405 gnd.n6985 gnd.n6984 9.3005
R19406 gnd.n613 gnd.n612 9.3005
R19407 gnd.n6992 gnd.n6991 9.3005
R19408 gnd.n6993 gnd.n611 9.3005
R19409 gnd.n6995 gnd.n6994 9.3005
R19410 gnd.n607 gnd.n606 9.3005
R19411 gnd.n7002 gnd.n7001 9.3005
R19412 gnd.n7003 gnd.n605 9.3005
R19413 gnd.n7005 gnd.n7004 9.3005
R19414 gnd.n601 gnd.n600 9.3005
R19415 gnd.n7012 gnd.n7011 9.3005
R19416 gnd.n7013 gnd.n599 9.3005
R19417 gnd.n7015 gnd.n7014 9.3005
R19418 gnd.n595 gnd.n594 9.3005
R19419 gnd.n7022 gnd.n7021 9.3005
R19420 gnd.n7023 gnd.n593 9.3005
R19421 gnd.n7025 gnd.n7024 9.3005
R19422 gnd.n589 gnd.n588 9.3005
R19423 gnd.n7032 gnd.n7031 9.3005
R19424 gnd.n7033 gnd.n587 9.3005
R19425 gnd.n7035 gnd.n7034 9.3005
R19426 gnd.n583 gnd.n582 9.3005
R19427 gnd.n7042 gnd.n7041 9.3005
R19428 gnd.n7043 gnd.n581 9.3005
R19429 gnd.n7045 gnd.n7044 9.3005
R19430 gnd.n577 gnd.n576 9.3005
R19431 gnd.n7052 gnd.n7051 9.3005
R19432 gnd.n7053 gnd.n575 9.3005
R19433 gnd.n7055 gnd.n7054 9.3005
R19434 gnd.n571 gnd.n570 9.3005
R19435 gnd.n7062 gnd.n7061 9.3005
R19436 gnd.n7063 gnd.n569 9.3005
R19437 gnd.n7065 gnd.n7064 9.3005
R19438 gnd.n565 gnd.n564 9.3005
R19439 gnd.n7072 gnd.n7071 9.3005
R19440 gnd.n7073 gnd.n563 9.3005
R19441 gnd.n7075 gnd.n7074 9.3005
R19442 gnd.n559 gnd.n558 9.3005
R19443 gnd.n7082 gnd.n7081 9.3005
R19444 gnd.n7083 gnd.n557 9.3005
R19445 gnd.n7085 gnd.n7084 9.3005
R19446 gnd.n553 gnd.n552 9.3005
R19447 gnd.n7092 gnd.n7091 9.3005
R19448 gnd.n7093 gnd.n551 9.3005
R19449 gnd.n7095 gnd.n7094 9.3005
R19450 gnd.n547 gnd.n546 9.3005
R19451 gnd.n7102 gnd.n7101 9.3005
R19452 gnd.n7103 gnd.n545 9.3005
R19453 gnd.n7105 gnd.n7104 9.3005
R19454 gnd.n541 gnd.n540 9.3005
R19455 gnd.n7112 gnd.n7111 9.3005
R19456 gnd.n7113 gnd.n539 9.3005
R19457 gnd.n7115 gnd.n7114 9.3005
R19458 gnd.n535 gnd.n534 9.3005
R19459 gnd.n7122 gnd.n7121 9.3005
R19460 gnd.n7123 gnd.n533 9.3005
R19461 gnd.n7125 gnd.n7124 9.3005
R19462 gnd.n529 gnd.n528 9.3005
R19463 gnd.n7132 gnd.n7131 9.3005
R19464 gnd.n7135 gnd.n7134 9.3005
R19465 gnd.n523 gnd.n522 9.3005
R19466 gnd.n7142 gnd.n7141 9.3005
R19467 gnd.n7143 gnd.n521 9.3005
R19468 gnd.n7145 gnd.n7144 9.3005
R19469 gnd.n517 gnd.n516 9.3005
R19470 gnd.n7152 gnd.n7151 9.3005
R19471 gnd.n7153 gnd.n515 9.3005
R19472 gnd.n7155 gnd.n7154 9.3005
R19473 gnd.n511 gnd.n510 9.3005
R19474 gnd.n7162 gnd.n7161 9.3005
R19475 gnd.n7163 gnd.n509 9.3005
R19476 gnd.n7165 gnd.n7164 9.3005
R19477 gnd.n505 gnd.n504 9.3005
R19478 gnd.n7172 gnd.n7171 9.3005
R19479 gnd.n7173 gnd.n503 9.3005
R19480 gnd.n7175 gnd.n7174 9.3005
R19481 gnd.n499 gnd.n498 9.3005
R19482 gnd.n7182 gnd.n7181 9.3005
R19483 gnd.n7183 gnd.n497 9.3005
R19484 gnd.n7185 gnd.n7184 9.3005
R19485 gnd.n493 gnd.n492 9.3005
R19486 gnd.n7192 gnd.n7191 9.3005
R19487 gnd.n7193 gnd.n491 9.3005
R19488 gnd.n7195 gnd.n7194 9.3005
R19489 gnd.n487 gnd.n486 9.3005
R19490 gnd.n7202 gnd.n7201 9.3005
R19491 gnd.n7203 gnd.n485 9.3005
R19492 gnd.n7205 gnd.n7204 9.3005
R19493 gnd.n481 gnd.n480 9.3005
R19494 gnd.n7212 gnd.n7211 9.3005
R19495 gnd.n7213 gnd.n479 9.3005
R19496 gnd.n7215 gnd.n7214 9.3005
R19497 gnd.n475 gnd.n474 9.3005
R19498 gnd.n7222 gnd.n7221 9.3005
R19499 gnd.n7223 gnd.n473 9.3005
R19500 gnd.n7225 gnd.n7224 9.3005
R19501 gnd.n469 gnd.n468 9.3005
R19502 gnd.n7232 gnd.n7231 9.3005
R19503 gnd.n7233 gnd.n467 9.3005
R19504 gnd.n7235 gnd.n7234 9.3005
R19505 gnd.n463 gnd.n462 9.3005
R19506 gnd.n7242 gnd.n7241 9.3005
R19507 gnd.n7243 gnd.n461 9.3005
R19508 gnd.n7245 gnd.n7244 9.3005
R19509 gnd.n457 gnd.n456 9.3005
R19510 gnd.n7252 gnd.n7251 9.3005
R19511 gnd.n7253 gnd.n455 9.3005
R19512 gnd.n7255 gnd.n7254 9.3005
R19513 gnd.n451 gnd.n450 9.3005
R19514 gnd.n7262 gnd.n7261 9.3005
R19515 gnd.n7263 gnd.n449 9.3005
R19516 gnd.n7265 gnd.n7264 9.3005
R19517 gnd.n445 gnd.n444 9.3005
R19518 gnd.n7272 gnd.n7271 9.3005
R19519 gnd.n7273 gnd.n443 9.3005
R19520 gnd.n7275 gnd.n7274 9.3005
R19521 gnd.n439 gnd.n438 9.3005
R19522 gnd.n7282 gnd.n7281 9.3005
R19523 gnd.n7283 gnd.n437 9.3005
R19524 gnd.n7285 gnd.n7284 9.3005
R19525 gnd.n433 gnd.n432 9.3005
R19526 gnd.n7292 gnd.n7291 9.3005
R19527 gnd.n7293 gnd.n431 9.3005
R19528 gnd.n7295 gnd.n7294 9.3005
R19529 gnd.n427 gnd.n426 9.3005
R19530 gnd.n7302 gnd.n7301 9.3005
R19531 gnd.n7303 gnd.n425 9.3005
R19532 gnd.n7305 gnd.n7304 9.3005
R19533 gnd.n421 gnd.n420 9.3005
R19534 gnd.n7312 gnd.n7311 9.3005
R19535 gnd.n7313 gnd.n419 9.3005
R19536 gnd.n7315 gnd.n7314 9.3005
R19537 gnd.n415 gnd.n414 9.3005
R19538 gnd.n7322 gnd.n7321 9.3005
R19539 gnd.n7323 gnd.n413 9.3005
R19540 gnd.n7325 gnd.n7324 9.3005
R19541 gnd.n409 gnd.n408 9.3005
R19542 gnd.n7332 gnd.n7331 9.3005
R19543 gnd.n7333 gnd.n407 9.3005
R19544 gnd.n7337 gnd.n7334 9.3005
R19545 gnd.n7336 gnd.n7335 9.3005
R19546 gnd.n403 gnd.n402 9.3005
R19547 gnd.n7345 gnd.n7344 9.3005
R19548 gnd.n7133 gnd.n527 9.3005
R19549 gnd.n7681 gnd.n7680 9.3005
R19550 gnd.n7679 gnd.n80 9.3005
R19551 gnd.n7370 gnd.n83 9.3005
R19552 gnd.n7372 gnd.n7371 9.3005
R19553 gnd.n377 gnd.n376 9.3005
R19554 gnd.n7383 gnd.n7382 9.3005
R19555 gnd.n7384 gnd.n375 9.3005
R19556 gnd.n7386 gnd.n7385 9.3005
R19557 gnd.n370 gnd.n369 9.3005
R19558 gnd.n7397 gnd.n7396 9.3005
R19559 gnd.n7398 gnd.n368 9.3005
R19560 gnd.n7400 gnd.n7399 9.3005
R19561 gnd.n365 gnd.n364 9.3005
R19562 gnd.n7411 gnd.n7410 9.3005
R19563 gnd.n7412 gnd.n363 9.3005
R19564 gnd.n7415 gnd.n7414 9.3005
R19565 gnd.n7413 gnd.n359 9.3005
R19566 gnd.n7440 gnd.n358 9.3005
R19567 gnd.n7442 gnd.n7441 9.3005
R19568 gnd.n7443 gnd.n357 9.3005
R19569 gnd.n7445 gnd.n7444 9.3005
R19570 gnd.n7447 gnd.n355 9.3005
R19571 gnd.n7449 gnd.n7448 9.3005
R19572 gnd.n7450 gnd.n354 9.3005
R19573 gnd.n7452 gnd.n7451 9.3005
R19574 gnd.n7454 gnd.n352 9.3005
R19575 gnd.n7456 gnd.n7455 9.3005
R19576 gnd.n7487 gnd.n318 9.3005
R19577 gnd.n7486 gnd.n320 9.3005
R19578 gnd.n324 gnd.n321 9.3005
R19579 gnd.n7481 gnd.n325 9.3005
R19580 gnd.n7480 gnd.n326 9.3005
R19581 gnd.n7479 gnd.n327 9.3005
R19582 gnd.n331 gnd.n328 9.3005
R19583 gnd.n7474 gnd.n332 9.3005
R19584 gnd.n7473 gnd.n333 9.3005
R19585 gnd.n7472 gnd.n334 9.3005
R19586 gnd.n338 gnd.n335 9.3005
R19587 gnd.n7467 gnd.n339 9.3005
R19588 gnd.n7466 gnd.n340 9.3005
R19589 gnd.n7465 gnd.n341 9.3005
R19590 gnd.n345 gnd.n342 9.3005
R19591 gnd.n7460 gnd.n346 9.3005
R19592 gnd.n7459 gnd.n7458 9.3005
R19593 gnd.n7457 gnd.n349 9.3005
R19594 gnd.n7489 gnd.n7488 9.3005
R19595 gnd.n7597 gnd.n215 9.3005
R19596 gnd.n7596 gnd.n217 9.3005
R19597 gnd.n221 gnd.n218 9.3005
R19598 gnd.n7591 gnd.n222 9.3005
R19599 gnd.n7590 gnd.n223 9.3005
R19600 gnd.n7589 gnd.n224 9.3005
R19601 gnd.n228 gnd.n225 9.3005
R19602 gnd.n7584 gnd.n229 9.3005
R19603 gnd.n7583 gnd.n230 9.3005
R19604 gnd.n7582 gnd.n231 9.3005
R19605 gnd.n235 gnd.n232 9.3005
R19606 gnd.n7577 gnd.n236 9.3005
R19607 gnd.n7576 gnd.n237 9.3005
R19608 gnd.n7575 gnd.n238 9.3005
R19609 gnd.n242 gnd.n239 9.3005
R19610 gnd.n7570 gnd.n243 9.3005
R19611 gnd.n7569 gnd.n244 9.3005
R19612 gnd.n7565 gnd.n245 9.3005
R19613 gnd.n249 gnd.n246 9.3005
R19614 gnd.n7560 gnd.n250 9.3005
R19615 gnd.n7559 gnd.n251 9.3005
R19616 gnd.n7558 gnd.n252 9.3005
R19617 gnd.n256 gnd.n253 9.3005
R19618 gnd.n7553 gnd.n257 9.3005
R19619 gnd.n7552 gnd.n258 9.3005
R19620 gnd.n7551 gnd.n259 9.3005
R19621 gnd.n263 gnd.n260 9.3005
R19622 gnd.n7546 gnd.n264 9.3005
R19623 gnd.n7545 gnd.n265 9.3005
R19624 gnd.n7544 gnd.n266 9.3005
R19625 gnd.n270 gnd.n267 9.3005
R19626 gnd.n7539 gnd.n271 9.3005
R19627 gnd.n7538 gnd.n272 9.3005
R19628 gnd.n7537 gnd.n273 9.3005
R19629 gnd.n277 gnd.n274 9.3005
R19630 gnd.n7532 gnd.n278 9.3005
R19631 gnd.n7531 gnd.n7530 9.3005
R19632 gnd.n7529 gnd.n279 9.3005
R19633 gnd.n7528 gnd.n7527 9.3005
R19634 gnd.n283 gnd.n282 9.3005
R19635 gnd.n288 gnd.n286 9.3005
R19636 gnd.n7520 gnd.n289 9.3005
R19637 gnd.n7519 gnd.n290 9.3005
R19638 gnd.n7518 gnd.n291 9.3005
R19639 gnd.n295 gnd.n292 9.3005
R19640 gnd.n7513 gnd.n296 9.3005
R19641 gnd.n7512 gnd.n297 9.3005
R19642 gnd.n7511 gnd.n298 9.3005
R19643 gnd.n302 gnd.n299 9.3005
R19644 gnd.n7506 gnd.n303 9.3005
R19645 gnd.n7505 gnd.n304 9.3005
R19646 gnd.n7504 gnd.n305 9.3005
R19647 gnd.n309 gnd.n306 9.3005
R19648 gnd.n7499 gnd.n310 9.3005
R19649 gnd.n7498 gnd.n311 9.3005
R19650 gnd.n7497 gnd.n312 9.3005
R19651 gnd.n317 gnd.n315 9.3005
R19652 gnd.n7492 gnd.n7491 9.3005
R19653 gnd.n7599 gnd.n7598 9.3005
R19654 gnd.n4396 gnd.n4395 9.3005
R19655 gnd.n1793 gnd.n1792 9.3005
R19656 gnd.n1818 gnd.n1817 9.3005
R19657 gnd.n4383 gnd.n1819 9.3005
R19658 gnd.n4382 gnd.n1820 9.3005
R19659 gnd.n4381 gnd.n1821 9.3005
R19660 gnd.n4201 gnd.n1822 9.3005
R19661 gnd.n4371 gnd.n1839 9.3005
R19662 gnd.n4370 gnd.n1840 9.3005
R19663 gnd.n4369 gnd.n1841 9.3005
R19664 gnd.n4216 gnd.n1842 9.3005
R19665 gnd.n4359 gnd.n1859 9.3005
R19666 gnd.n4358 gnd.n1860 9.3005
R19667 gnd.n4357 gnd.n1861 9.3005
R19668 gnd.n4223 gnd.n1862 9.3005
R19669 gnd.n4347 gnd.n1879 9.3005
R19670 gnd.n4346 gnd.n1880 9.3005
R19671 gnd.n4345 gnd.n1881 9.3005
R19672 gnd.n4229 gnd.n1882 9.3005
R19673 gnd.n4335 gnd.n1899 9.3005
R19674 gnd.n4334 gnd.n1900 9.3005
R19675 gnd.n4333 gnd.n1901 9.3005
R19676 gnd.n4294 gnd.n1902 9.3005
R19677 gnd.n4295 gnd.n1931 9.3005
R19678 gnd.n4311 gnd.n1932 9.3005
R19679 gnd.n4310 gnd.n1933 9.3005
R19680 gnd.n4309 gnd.n1934 9.3005
R19681 gnd.n4303 gnd.n1935 9.3005
R19682 gnd.n4302 gnd.n4301 9.3005
R19683 gnd.n379 gnd.n108 9.3005
R19684 gnd.n7667 gnd.n109 9.3005
R19685 gnd.n7666 gnd.n110 9.3005
R19686 gnd.n7665 gnd.n111 9.3005
R19687 gnd.n373 gnd.n112 9.3005
R19688 gnd.n7655 gnd.n127 9.3005
R19689 gnd.n7654 gnd.n128 9.3005
R19690 gnd.n7653 gnd.n129 9.3005
R19691 gnd.n367 gnd.n130 9.3005
R19692 gnd.n7643 gnd.n148 9.3005
R19693 gnd.n7642 gnd.n149 9.3005
R19694 gnd.n7641 gnd.n150 9.3005
R19695 gnd.n361 gnd.n151 9.3005
R19696 gnd.n7631 gnd.n167 9.3005
R19697 gnd.n7630 gnd.n168 9.3005
R19698 gnd.n7629 gnd.n169 9.3005
R19699 gnd.n7421 gnd.n170 9.3005
R19700 gnd.n7619 gnd.n187 9.3005
R19701 gnd.n7618 gnd.n188 9.3005
R19702 gnd.n7617 gnd.n189 9.3005
R19703 gnd.n7422 gnd.n190 9.3005
R19704 gnd.n7607 gnd.n205 9.3005
R19705 gnd.n7606 gnd.n206 9.3005
R19706 gnd.n7605 gnd.n207 9.3005
R19707 gnd.n4397 gnd.n1791 9.3005
R19708 gnd.n4395 gnd.n4394 9.3005
R19709 gnd.n4393 gnd.n1793 9.3005
R19710 gnd.n1818 gnd.n1794 9.3005
R19711 gnd.n1966 gnd.n1819 9.3005
R19712 gnd.n4199 gnd.n1820 9.3005
R19713 gnd.n4200 gnd.n1821 9.3005
R19714 gnd.n4202 gnd.n4201 9.3005
R19715 gnd.n1961 gnd.n1839 9.3005
R19716 gnd.n4214 gnd.n1840 9.3005
R19717 gnd.n4215 gnd.n1841 9.3005
R19718 gnd.n4217 gnd.n4216 9.3005
R19719 gnd.n4218 gnd.n1859 9.3005
R19720 gnd.n4221 gnd.n1860 9.3005
R19721 gnd.n4222 gnd.n1861 9.3005
R19722 gnd.n4227 gnd.n4223 9.3005
R19723 gnd.n4228 gnd.n1879 9.3005
R19724 gnd.n4232 gnd.n1880 9.3005
R19725 gnd.n4231 gnd.n1881 9.3005
R19726 gnd.n4230 gnd.n4229 9.3005
R19727 gnd.n1936 gnd.n1899 9.3005
R19728 gnd.n4291 gnd.n1900 9.3005
R19729 gnd.n4292 gnd.n1901 9.3005
R19730 gnd.n4294 gnd.n4293 9.3005
R19731 gnd.n4297 gnd.n4295 9.3005
R19732 gnd.n4298 gnd.n1932 9.3005
R19733 gnd.n4299 gnd.n1933 9.3005
R19734 gnd.n4305 gnd.n1934 9.3005
R19735 gnd.n4304 gnd.n4303 9.3005
R19736 gnd.n4302 gnd.n378 9.3005
R19737 gnd.n7376 gnd.n379 9.3005
R19738 gnd.n7377 gnd.n109 9.3005
R19739 gnd.n7378 gnd.n110 9.3005
R19740 gnd.n372 gnd.n111 9.3005
R19741 gnd.n7390 gnd.n373 9.3005
R19742 gnd.n7391 gnd.n127 9.3005
R19743 gnd.n7392 gnd.n128 9.3005
R19744 gnd.n366 gnd.n129 9.3005
R19745 gnd.n7404 gnd.n367 9.3005
R19746 gnd.n7405 gnd.n148 9.3005
R19747 gnd.n7406 gnd.n149 9.3005
R19748 gnd.n360 gnd.n150 9.3005
R19749 gnd.n7419 gnd.n361 9.3005
R19750 gnd.n7420 gnd.n167 9.3005
R19751 gnd.n7436 gnd.n168 9.3005
R19752 gnd.n7435 gnd.n169 9.3005
R19753 gnd.n7434 gnd.n7421 9.3005
R19754 gnd.n7432 gnd.n187 9.3005
R19755 gnd.n7431 gnd.n188 9.3005
R19756 gnd.n7429 gnd.n189 9.3005
R19757 gnd.n7428 gnd.n7422 9.3005
R19758 gnd.n7426 gnd.n205 9.3005
R19759 gnd.n7425 gnd.n206 9.3005
R19760 gnd.n7423 gnd.n207 9.3005
R19761 gnd.n1791 gnd.n1785 9.3005
R19762 gnd.n4407 gnd.n4406 9.3005
R19763 gnd.n4410 gnd.n1783 9.3005
R19764 gnd.n4411 gnd.n1782 9.3005
R19765 gnd.n4414 gnd.n1781 9.3005
R19766 gnd.n4415 gnd.n1780 9.3005
R19767 gnd.n4418 gnd.n1779 9.3005
R19768 gnd.n4419 gnd.n1778 9.3005
R19769 gnd.n4422 gnd.n1777 9.3005
R19770 gnd.n4423 gnd.n1776 9.3005
R19771 gnd.n4426 gnd.n1775 9.3005
R19772 gnd.n4427 gnd.n1774 9.3005
R19773 gnd.n4430 gnd.n1773 9.3005
R19774 gnd.n4431 gnd.n1772 9.3005
R19775 gnd.n4434 gnd.n1771 9.3005
R19776 gnd.n4435 gnd.n1770 9.3005
R19777 gnd.n4438 gnd.n1769 9.3005
R19778 gnd.n4439 gnd.n1768 9.3005
R19779 gnd.n4442 gnd.n1767 9.3005
R19780 gnd.n4443 gnd.n1766 9.3005
R19781 gnd.n4446 gnd.n1765 9.3005
R19782 gnd.n4450 gnd.n1761 9.3005
R19783 gnd.n4451 gnd.n1760 9.3005
R19784 gnd.n4454 gnd.n1759 9.3005
R19785 gnd.n4455 gnd.n1758 9.3005
R19786 gnd.n4458 gnd.n1757 9.3005
R19787 gnd.n4459 gnd.n1756 9.3005
R19788 gnd.n4462 gnd.n1755 9.3005
R19789 gnd.n4463 gnd.n1754 9.3005
R19790 gnd.n4466 gnd.n1753 9.3005
R19791 gnd.n4468 gnd.n1749 9.3005
R19792 gnd.n4471 gnd.n1748 9.3005
R19793 gnd.n4472 gnd.n1747 9.3005
R19794 gnd.n4475 gnd.n1746 9.3005
R19795 gnd.n4476 gnd.n1745 9.3005
R19796 gnd.n4479 gnd.n1744 9.3005
R19797 gnd.n4480 gnd.n1743 9.3005
R19798 gnd.n4483 gnd.n1742 9.3005
R19799 gnd.n4485 gnd.n1739 9.3005
R19800 gnd.n4488 gnd.n1738 9.3005
R19801 gnd.n4489 gnd.n1737 9.3005
R19802 gnd.n4492 gnd.n1736 9.3005
R19803 gnd.n4493 gnd.n1735 9.3005
R19804 gnd.n4496 gnd.n1734 9.3005
R19805 gnd.n4497 gnd.n1733 9.3005
R19806 gnd.n4500 gnd.n1732 9.3005
R19807 gnd.n4501 gnd.n1731 9.3005
R19808 gnd.n4504 gnd.n1730 9.3005
R19809 gnd.n4505 gnd.n1729 9.3005
R19810 gnd.n4508 gnd.n1728 9.3005
R19811 gnd.n4509 gnd.n1727 9.3005
R19812 gnd.n4512 gnd.n1726 9.3005
R19813 gnd.n4514 gnd.n1725 9.3005
R19814 gnd.n4515 gnd.n1724 9.3005
R19815 gnd.n4516 gnd.n1723 9.3005
R19816 gnd.n4517 gnd.n1722 9.3005
R19817 gnd.n4447 gnd.n1762 9.3005
R19818 gnd.n4405 gnd.n4402 9.3005
R19819 gnd.n1805 gnd.n1802 9.3005
R19820 gnd.n4389 gnd.n1806 9.3005
R19821 gnd.n4388 gnd.n1807 9.3005
R19822 gnd.n4387 gnd.n1808 9.3005
R19823 gnd.n1828 gnd.n1809 9.3005
R19824 gnd.n4377 gnd.n1829 9.3005
R19825 gnd.n4376 gnd.n1830 9.3005
R19826 gnd.n4375 gnd.n1831 9.3005
R19827 gnd.n1849 gnd.n1832 9.3005
R19828 gnd.n4365 gnd.n1850 9.3005
R19829 gnd.n4364 gnd.n1851 9.3005
R19830 gnd.n4363 gnd.n1852 9.3005
R19831 gnd.n1868 gnd.n1853 9.3005
R19832 gnd.n4353 gnd.n1869 9.3005
R19833 gnd.n4352 gnd.n1870 9.3005
R19834 gnd.n4351 gnd.n1871 9.3005
R19835 gnd.n1889 gnd.n1872 9.3005
R19836 gnd.n4341 gnd.n1890 9.3005
R19837 gnd.n4340 gnd.n1891 9.3005
R19838 gnd.n4339 gnd.n1892 9.3005
R19839 gnd.n1893 gnd.n94 9.3005
R19840 gnd.n99 gnd.n93 9.3005
R19841 gnd.n7661 gnd.n118 9.3005
R19842 gnd.n7660 gnd.n119 9.3005
R19843 gnd.n7659 gnd.n120 9.3005
R19844 gnd.n137 gnd.n121 9.3005
R19845 gnd.n7649 gnd.n138 9.3005
R19846 gnd.n7648 gnd.n139 9.3005
R19847 gnd.n7647 gnd.n140 9.3005
R19848 gnd.n157 gnd.n141 9.3005
R19849 gnd.n7637 gnd.n158 9.3005
R19850 gnd.n7636 gnd.n159 9.3005
R19851 gnd.n7635 gnd.n160 9.3005
R19852 gnd.n177 gnd.n161 9.3005
R19853 gnd.n7625 gnd.n178 9.3005
R19854 gnd.n7624 gnd.n179 9.3005
R19855 gnd.n7623 gnd.n180 9.3005
R19856 gnd.n196 gnd.n181 9.3005
R19857 gnd.n7613 gnd.n197 9.3005
R19858 gnd.n7612 gnd.n198 9.3005
R19859 gnd.n7611 gnd.n199 9.3005
R19860 gnd.n214 gnd.n200 9.3005
R19861 gnd.n7601 gnd.n7600 9.3005
R19862 gnd.n1804 gnd.n1803 9.3005
R19863 gnd.n7672 gnd.n97 9.3005
R19864 gnd.n7672 gnd.n7671 9.3005
R19865 gnd.n2990 gnd.n2973 9.3005
R19866 gnd.n2976 gnd.n2974 9.3005
R19867 gnd.n2986 gnd.n2977 9.3005
R19868 gnd.n2985 gnd.n2978 9.3005
R19869 gnd.n2984 gnd.n2979 9.3005
R19870 gnd.n2982 gnd.n2981 9.3005
R19871 gnd.n2980 gnd.n2647 9.3005
R19872 gnd.n2645 gnd.n2644 9.3005
R19873 gnd.n3061 gnd.n3060 9.3005
R19874 gnd.n3062 gnd.n2643 9.3005
R19875 gnd.n3064 gnd.n3063 9.3005
R19876 gnd.n2641 gnd.n2640 9.3005
R19877 gnd.n3069 gnd.n3068 9.3005
R19878 gnd.n3070 gnd.n2639 9.3005
R19879 gnd.n3118 gnd.n3071 9.3005
R19880 gnd.n3117 gnd.n3072 9.3005
R19881 gnd.n3116 gnd.n3073 9.3005
R19882 gnd.n3076 gnd.n3074 9.3005
R19883 gnd.n3112 gnd.n3077 9.3005
R19884 gnd.n3111 gnd.n3078 9.3005
R19885 gnd.n3110 gnd.n3079 9.3005
R19886 gnd.n3082 gnd.n3080 9.3005
R19887 gnd.n3105 gnd.n3083 9.3005
R19888 gnd.n3104 gnd.n3084 9.3005
R19889 gnd.n3103 gnd.n3085 9.3005
R19890 gnd.n3090 gnd.n3086 9.3005
R19891 gnd.n3097 gnd.n3091 9.3005
R19892 gnd.n3096 gnd.n3092 9.3005
R19893 gnd.n3095 gnd.n3093 9.3005
R19894 gnd.n2401 gnd.n2400 9.3005
R19895 gnd.n3244 gnd.n3243 9.3005
R19896 gnd.n3245 gnd.n2399 9.3005
R19897 gnd.n3249 gnd.n3246 9.3005
R19898 gnd.n3248 gnd.n3247 9.3005
R19899 gnd.n2376 gnd.n2375 9.3005
R19900 gnd.n3274 gnd.n3273 9.3005
R19901 gnd.n3275 gnd.n2374 9.3005
R19902 gnd.n3286 gnd.n3276 9.3005
R19903 gnd.n3285 gnd.n3277 9.3005
R19904 gnd.n3284 gnd.n3278 9.3005
R19905 gnd.n3281 gnd.n3280 9.3005
R19906 gnd.n3279 gnd.n1495 9.3005
R19907 gnd.n4706 gnd.n1496 9.3005
R19908 gnd.n4705 gnd.n1497 9.3005
R19909 gnd.n4704 gnd.n1498 9.3005
R19910 gnd.n1511 gnd.n1499 9.3005
R19911 gnd.n4692 gnd.n1512 9.3005
R19912 gnd.n4691 gnd.n1513 9.3005
R19913 gnd.n4690 gnd.n1514 9.3005
R19914 gnd.n1529 gnd.n1515 9.3005
R19915 gnd.n4678 gnd.n1530 9.3005
R19916 gnd.n4677 gnd.n1531 9.3005
R19917 gnd.n4676 gnd.n1532 9.3005
R19918 gnd.n3482 gnd.n1533 9.3005
R19919 gnd.n3485 gnd.n3484 9.3005
R19920 gnd.n3486 gnd.n3481 9.3005
R19921 gnd.n3498 gnd.n3487 9.3005
R19922 gnd.n3497 gnd.n3488 9.3005
R19923 gnd.n3496 gnd.n3489 9.3005
R19924 gnd.n3491 gnd.n3490 9.3005
R19925 gnd.n2276 gnd.n2275 9.3005
R19926 gnd.n3567 gnd.n3566 9.3005
R19927 gnd.n3568 gnd.n2274 9.3005
R19928 gnd.n3570 gnd.n3569 9.3005
R19929 gnd.n2252 gnd.n2251 9.3005
R19930 gnd.n3606 gnd.n3605 9.3005
R19931 gnd.n3607 gnd.n2250 9.3005
R19932 gnd.n3609 gnd.n3608 9.3005
R19933 gnd.n2230 gnd.n2229 9.3005
R19934 gnd.n3660 gnd.n3659 9.3005
R19935 gnd.n3661 gnd.n2228 9.3005
R19936 gnd.n3663 gnd.n3662 9.3005
R19937 gnd.n2211 gnd.n2210 9.3005
R19938 gnd.n3686 gnd.n3685 9.3005
R19939 gnd.n3687 gnd.n2209 9.3005
R19940 gnd.n3689 gnd.n3688 9.3005
R19941 gnd.n2188 gnd.n2187 9.3005
R19942 gnd.n3752 gnd.n3751 9.3005
R19943 gnd.n3753 gnd.n2186 9.3005
R19944 gnd.n3755 gnd.n3754 9.3005
R19945 gnd.n2166 gnd.n2165 9.3005
R19946 gnd.n3782 gnd.n3781 9.3005
R19947 gnd.n3783 gnd.n2164 9.3005
R19948 gnd.n3785 gnd.n3784 9.3005
R19949 gnd.n2144 gnd.n2143 9.3005
R19950 gnd.n3813 gnd.n3812 9.3005
R19951 gnd.n3814 gnd.n2142 9.3005
R19952 gnd.n3816 gnd.n3815 9.3005
R19953 gnd.n2118 gnd.n2117 9.3005
R19954 gnd.n3862 gnd.n3861 9.3005
R19955 gnd.n3863 gnd.n2116 9.3005
R19956 gnd.n3865 gnd.n3864 9.3005
R19957 gnd.n2102 gnd.n2101 9.3005
R19958 gnd.n3893 gnd.n3892 9.3005
R19959 gnd.n3894 gnd.n2100 9.3005
R19960 gnd.n3896 gnd.n3895 9.3005
R19961 gnd.n2048 gnd.n2047 9.3005
R19962 gnd.n4064 gnd.n4063 9.3005
R19963 gnd.n4065 gnd.n2046 9.3005
R19964 gnd.n4067 gnd.n4066 9.3005
R19965 gnd.n2035 gnd.n2034 9.3005
R19966 gnd.n4084 gnd.n4083 9.3005
R19967 gnd.n4085 gnd.n2033 9.3005
R19968 gnd.n4087 gnd.n4086 9.3005
R19969 gnd.n2022 gnd.n2021 9.3005
R19970 gnd.n4104 gnd.n4103 9.3005
R19971 gnd.n4105 gnd.n2020 9.3005
R19972 gnd.n4109 gnd.n4106 9.3005
R19973 gnd.n4108 gnd.n4107 9.3005
R19974 gnd.n2007 gnd.n2006 9.3005
R19975 gnd.n4128 gnd.n4127 9.3005
R19976 gnd.n4129 gnd.n2005 9.3005
R19977 gnd.n4175 gnd.n4130 9.3005
R19978 gnd.n4174 gnd.n4131 9.3005
R19979 gnd.n4173 gnd.n4132 9.3005
R19980 gnd.n4135 gnd.n4133 9.3005
R19981 gnd.n4169 gnd.n4136 9.3005
R19982 gnd.n4168 gnd.n4137 9.3005
R19983 gnd.n4167 gnd.n4138 9.3005
R19984 gnd.n4141 gnd.n4139 9.3005
R19985 gnd.n4163 gnd.n4142 9.3005
R19986 gnd.n4162 gnd.n4143 9.3005
R19987 gnd.n4161 gnd.n4144 9.3005
R19988 gnd.n4147 gnd.n4145 9.3005
R19989 gnd.n4157 gnd.n4148 9.3005
R19990 gnd.n4156 gnd.n4149 9.3005
R19991 gnd.n4155 gnd.n4150 9.3005
R19992 gnd.n4153 gnd.n4152 9.3005
R19993 gnd.n4151 gnd.n1952 9.3005
R19994 gnd.n1950 gnd.n1949 9.3005
R19995 gnd.n4254 gnd.n4253 9.3005
R19996 gnd.n4255 gnd.n1948 9.3005
R19997 gnd.n4257 gnd.n4256 9.3005
R19998 gnd.n1946 gnd.n1945 9.3005
R19999 gnd.n4262 gnd.n4261 9.3005
R20000 gnd.n4263 gnd.n1944 9.3005
R20001 gnd.n4270 gnd.n4264 9.3005
R20002 gnd.n4269 gnd.n4265 9.3005
R20003 gnd.n7364 gnd.n385 9.3005
R20004 gnd.n388 gnd.n386 9.3005
R20005 gnd.n7360 gnd.n389 9.3005
R20006 gnd.n7359 gnd.n390 9.3005
R20007 gnd.n7358 gnd.n391 9.3005
R20008 gnd.n394 gnd.n392 9.3005
R20009 gnd.n7354 gnd.n395 9.3005
R20010 gnd.n7353 gnd.n396 9.3005
R20011 gnd.n7352 gnd.n397 9.3005
R20012 gnd.n400 gnd.n398 9.3005
R20013 gnd.n7348 gnd.n401 9.3005
R20014 gnd.n7347 gnd.n7346 9.3005
R20015 gnd.n2809 gnd.n2747 9.3005
R20016 gnd.n2812 gnd.n2811 9.3005
R20017 gnd.n2813 gnd.n2746 9.3005
R20018 gnd.n2816 gnd.n2814 9.3005
R20019 gnd.n2817 gnd.n2745 9.3005
R20020 gnd.n2820 gnd.n2819 9.3005
R20021 gnd.n2821 gnd.n2744 9.3005
R20022 gnd.n2824 gnd.n2822 9.3005
R20023 gnd.n2825 gnd.n2743 9.3005
R20024 gnd.n2845 gnd.n2844 9.3005
R20025 gnd.n2846 gnd.n2742 9.3005
R20026 gnd.n2849 gnd.n2848 9.3005
R20027 gnd.n2847 gnd.n2736 9.3005
R20028 gnd.n2888 gnd.n2737 9.3005
R20029 gnd.n2887 gnd.n2738 9.3005
R20030 gnd.n2886 gnd.n2739 9.3005
R20031 gnd.n2860 gnd.n2740 9.3005
R20032 gnd.n2876 gnd.n2861 9.3005
R20033 gnd.n2875 gnd.n2862 9.3005
R20034 gnd.n2874 gnd.n2863 9.3005
R20035 gnd.n2868 gnd.n2864 9.3005
R20036 gnd.n2867 gnd.n2865 9.3005
R20037 gnd.n2695 gnd.n2694 9.3005
R20038 gnd.n2937 gnd.n2936 9.3005
R20039 gnd.n2938 gnd.n2693 9.3005
R20040 gnd.n2946 gnd.n2939 9.3005
R20041 gnd.n2808 gnd.n2806 9.3005
R20042 gnd.n2802 gnd.n2801 9.3005
R20043 gnd.n2800 gnd.n2752 9.3005
R20044 gnd.n2799 gnd.n2798 9.3005
R20045 gnd.n2795 gnd.n2755 9.3005
R20046 gnd.n2794 gnd.n2791 9.3005
R20047 gnd.n2790 gnd.n2756 9.3005
R20048 gnd.n2789 gnd.n2788 9.3005
R20049 gnd.n2785 gnd.n2757 9.3005
R20050 gnd.n2784 gnd.n2781 9.3005
R20051 gnd.n2780 gnd.n2758 9.3005
R20052 gnd.n2779 gnd.n2778 9.3005
R20053 gnd.n2775 gnd.n2759 9.3005
R20054 gnd.n2774 gnd.n2771 9.3005
R20055 gnd.n2770 gnd.n2760 9.3005
R20056 gnd.n2769 gnd.n2768 9.3005
R20057 gnd.n2765 gnd.n2761 9.3005
R20058 gnd.n2764 gnd.n1136 9.3005
R20059 gnd.n2803 gnd.n2748 9.3005
R20060 gnd.n2805 gnd.n2804 9.3005
R20061 gnd.n4784 gnd.n1424 9.3005
R20062 gnd.n4785 gnd.n1423 9.3005
R20063 gnd.n1422 gnd.n1419 9.3005
R20064 gnd.n4790 gnd.n1418 9.3005
R20065 gnd.n4791 gnd.n1417 9.3005
R20066 gnd.n4792 gnd.n1416 9.3005
R20067 gnd.n1415 gnd.n1412 9.3005
R20068 gnd.n4797 gnd.n1411 9.3005
R20069 gnd.n4799 gnd.n1408 9.3005
R20070 gnd.n4800 gnd.n1407 9.3005
R20071 gnd.n1406 gnd.n1403 9.3005
R20072 gnd.n4805 gnd.n1402 9.3005
R20073 gnd.n4806 gnd.n1401 9.3005
R20074 gnd.n4807 gnd.n1400 9.3005
R20075 gnd.n1399 gnd.n1396 9.3005
R20076 gnd.n4812 gnd.n1395 9.3005
R20077 gnd.n4813 gnd.n1394 9.3005
R20078 gnd.n4814 gnd.n1393 9.3005
R20079 gnd.n1392 gnd.n1389 9.3005
R20080 gnd.n4819 gnd.n1388 9.3005
R20081 gnd.n4820 gnd.n1387 9.3005
R20082 gnd.n4821 gnd.n1386 9.3005
R20083 gnd.n1385 gnd.n1382 9.3005
R20084 gnd.n1384 gnd.n1380 9.3005
R20085 gnd.n4828 gnd.n1379 9.3005
R20086 gnd.n4830 gnd.n4829 9.3005
R20087 gnd.n2476 gnd.n2475 9.3005
R20088 gnd.n2484 gnd.n2483 9.3005
R20089 gnd.n2485 gnd.n2473 9.3005
R20090 gnd.n2487 gnd.n2486 9.3005
R20091 gnd.n2471 gnd.n2470 9.3005
R20092 gnd.n2494 gnd.n2493 9.3005
R20093 gnd.n2495 gnd.n2469 9.3005
R20094 gnd.n2497 gnd.n2496 9.3005
R20095 gnd.n2467 gnd.n2464 9.3005
R20096 gnd.n2504 gnd.n2503 9.3005
R20097 gnd.n2505 gnd.n2463 9.3005
R20098 gnd.n2507 gnd.n2506 9.3005
R20099 gnd.n2461 gnd.n2460 9.3005
R20100 gnd.n2514 gnd.n2513 9.3005
R20101 gnd.n2515 gnd.n2459 9.3005
R20102 gnd.n2517 gnd.n2516 9.3005
R20103 gnd.n2457 gnd.n2456 9.3005
R20104 gnd.n2524 gnd.n2523 9.3005
R20105 gnd.n2525 gnd.n2455 9.3005
R20106 gnd.n2527 gnd.n2526 9.3005
R20107 gnd.n2453 gnd.n2452 9.3005
R20108 gnd.n2534 gnd.n2533 9.3005
R20109 gnd.n2535 gnd.n2451 9.3005
R20110 gnd.n2537 gnd.n2536 9.3005
R20111 gnd.n2449 gnd.n2448 9.3005
R20112 gnd.n2544 gnd.n2543 9.3005
R20113 gnd.n2545 gnd.n2447 9.3005
R20114 gnd.n2547 gnd.n2546 9.3005
R20115 gnd.n2445 gnd.n2442 9.3005
R20116 gnd.n2553 gnd.n2552 9.3005
R20117 gnd.n2474 gnd.n1425 9.3005
R20118 gnd.n1158 gnd.n1138 9.3005
R20119 gnd.n2826 gnd.n1159 9.3005
R20120 gnd.n4960 gnd.n1160 9.3005
R20121 gnd.n4959 gnd.n1161 9.3005
R20122 gnd.n4958 gnd.n1162 9.3005
R20123 gnd.n2832 gnd.n1163 9.3005
R20124 gnd.n4948 gnd.n1179 9.3005
R20125 gnd.n4947 gnd.n1180 9.3005
R20126 gnd.n4946 gnd.n1181 9.3005
R20127 gnd.n2839 gnd.n1182 9.3005
R20128 gnd.n4936 gnd.n1199 9.3005
R20129 gnd.n4935 gnd.n1200 9.3005
R20130 gnd.n4934 gnd.n1201 9.3005
R20131 gnd.n2855 gnd.n1202 9.3005
R20132 gnd.n4924 gnd.n1219 9.3005
R20133 gnd.n4923 gnd.n1220 9.3005
R20134 gnd.n4922 gnd.n1221 9.3005
R20135 gnd.n2858 gnd.n1222 9.3005
R20136 gnd.n4912 gnd.n1240 9.3005
R20137 gnd.n4911 gnd.n1241 9.3005
R20138 gnd.n4910 gnd.n1242 9.3005
R20139 gnd.n2706 gnd.n1243 9.3005
R20140 gnd.n2921 gnd.n2705 9.3005
R20141 gnd.n2927 gnd.n2704 9.3005
R20142 gnd.n2929 gnd.n2928 9.3005
R20143 gnd.n2690 gnd.n2685 9.3005
R20144 gnd.n2959 gnd.n2686 9.3005
R20145 gnd.n2958 gnd.n2687 9.3005
R20146 gnd.n2957 gnd.n2956 9.3005
R20147 gnd.n2688 gnd.n1268 9.3005
R20148 gnd.n4898 gnd.n1269 9.3005
R20149 gnd.n4897 gnd.n1270 9.3005
R20150 gnd.n4896 gnd.n1271 9.3005
R20151 gnd.n3008 gnd.n1272 9.3005
R20152 gnd.n4886 gnd.n1288 9.3005
R20153 gnd.n4885 gnd.n1289 9.3005
R20154 gnd.n4884 gnd.n1290 9.3005
R20155 gnd.n3023 gnd.n1291 9.3005
R20156 gnd.n4874 gnd.n1308 9.3005
R20157 gnd.n4873 gnd.n1309 9.3005
R20158 gnd.n4872 gnd.n1310 9.3005
R20159 gnd.n3030 gnd.n1311 9.3005
R20160 gnd.n4862 gnd.n1328 9.3005
R20161 gnd.n4861 gnd.n1329 9.3005
R20162 gnd.n4860 gnd.n1330 9.3005
R20163 gnd.n2635 gnd.n1331 9.3005
R20164 gnd.n4850 gnd.n1348 9.3005
R20165 gnd.n4849 gnd.n1349 9.3005
R20166 gnd.n4848 gnd.n1350 9.3005
R20167 gnd.n2630 gnd.n1351 9.3005
R20168 gnd.n4838 gnd.n1369 9.3005
R20169 gnd.n4837 gnd.n1370 9.3005
R20170 gnd.n4836 gnd.n1371 9.3005
R20171 gnd.n4972 gnd.n1137 9.3005
R20172 gnd.n1139 gnd.n1138 9.3005
R20173 gnd.n2827 gnd.n2826 9.3005
R20174 gnd.n2828 gnd.n1160 9.3005
R20175 gnd.n2830 gnd.n1161 9.3005
R20176 gnd.n2831 gnd.n1162 9.3005
R20177 gnd.n2834 gnd.n2832 9.3005
R20178 gnd.n2835 gnd.n1179 9.3005
R20179 gnd.n2837 gnd.n1180 9.3005
R20180 gnd.n2838 gnd.n1181 9.3005
R20181 gnd.n2840 gnd.n2839 9.3005
R20182 gnd.n2741 gnd.n1199 9.3005
R20183 gnd.n2853 gnd.n1200 9.3005
R20184 gnd.n2854 gnd.n1201 9.3005
R20185 gnd.n2856 gnd.n2855 9.3005
R20186 gnd.n2857 gnd.n1219 9.3005
R20187 gnd.n2882 gnd.n1220 9.3005
R20188 gnd.n2881 gnd.n1221 9.3005
R20189 gnd.n2880 gnd.n2858 9.3005
R20190 gnd.n2859 gnd.n1240 9.3005
R20191 gnd.n2870 gnd.n1241 9.3005
R20192 gnd.n2869 gnd.n1242 9.3005
R20193 gnd.n2707 gnd.n2706 9.3005
R20194 gnd.n2925 gnd.n2705 9.3005
R20195 gnd.n2927 gnd.n2926 9.3005
R20196 gnd.n2928 gnd.n2689 9.3005
R20197 gnd.n2950 gnd.n2690 9.3005
R20198 gnd.n2951 gnd.n2686 9.3005
R20199 gnd.n2953 gnd.n2687 9.3005
R20200 gnd.n2956 gnd.n2955 9.3005
R20201 gnd.n2954 gnd.n2688 9.3005
R20202 gnd.n2662 gnd.n1269 9.3005
R20203 gnd.n3006 gnd.n1270 9.3005
R20204 gnd.n3007 gnd.n1271 9.3005
R20205 gnd.n3009 gnd.n3008 9.3005
R20206 gnd.n2657 gnd.n1288 9.3005
R20207 gnd.n3021 gnd.n1289 9.3005
R20208 gnd.n3022 gnd.n1290 9.3005
R20209 gnd.n3024 gnd.n3023 9.3005
R20210 gnd.n3025 gnd.n1308 9.3005
R20211 gnd.n3028 gnd.n1309 9.3005
R20212 gnd.n3029 gnd.n1310 9.3005
R20213 gnd.n3034 gnd.n3030 9.3005
R20214 gnd.n3035 gnd.n1328 9.3005
R20215 gnd.n3036 gnd.n1329 9.3005
R20216 gnd.n2634 gnd.n1330 9.3005
R20217 gnd.n3123 gnd.n2635 9.3005
R20218 gnd.n3124 gnd.n1348 9.3005
R20219 gnd.n3125 gnd.n1349 9.3005
R20220 gnd.n2629 gnd.n1350 9.3005
R20221 gnd.n3138 gnd.n2630 9.3005
R20222 gnd.n3139 gnd.n1369 9.3005
R20223 gnd.n3141 gnd.n1370 9.3005
R20224 gnd.n3140 gnd.n1371 9.3005
R20225 gnd.n4972 gnd.n4971 9.3005
R20226 gnd.n4976 gnd.n4975 9.3005
R20227 gnd.n4979 gnd.n1132 9.3005
R20228 gnd.n4980 gnd.n1131 9.3005
R20229 gnd.n4983 gnd.n1130 9.3005
R20230 gnd.n4984 gnd.n1129 9.3005
R20231 gnd.n4987 gnd.n1128 9.3005
R20232 gnd.n4988 gnd.n1127 9.3005
R20233 gnd.n4991 gnd.n1126 9.3005
R20234 gnd.n4992 gnd.n1125 9.3005
R20235 gnd.n4995 gnd.n1124 9.3005
R20236 gnd.n4996 gnd.n1123 9.3005
R20237 gnd.n4999 gnd.n1122 9.3005
R20238 gnd.n5000 gnd.n1121 9.3005
R20239 gnd.n5003 gnd.n1120 9.3005
R20240 gnd.n5004 gnd.n1119 9.3005
R20241 gnd.n5007 gnd.n1118 9.3005
R20242 gnd.n5008 gnd.n1117 9.3005
R20243 gnd.n5011 gnd.n1116 9.3005
R20244 gnd.n5012 gnd.n1115 9.3005
R20245 gnd.n5015 gnd.n1114 9.3005
R20246 gnd.n5019 gnd.n1110 9.3005
R20247 gnd.n5020 gnd.n1109 9.3005
R20248 gnd.n5023 gnd.n1108 9.3005
R20249 gnd.n5024 gnd.n1107 9.3005
R20250 gnd.n5027 gnd.n1106 9.3005
R20251 gnd.n5028 gnd.n1105 9.3005
R20252 gnd.n5031 gnd.n1104 9.3005
R20253 gnd.n5032 gnd.n1103 9.3005
R20254 gnd.n5035 gnd.n1102 9.3005
R20255 gnd.n5036 gnd.n1101 9.3005
R20256 gnd.n5039 gnd.n1100 9.3005
R20257 gnd.n5040 gnd.n1099 9.3005
R20258 gnd.n5043 gnd.n1098 9.3005
R20259 gnd.n5044 gnd.n1097 9.3005
R20260 gnd.n5047 gnd.n1096 9.3005
R20261 gnd.n5048 gnd.n1095 9.3005
R20262 gnd.n5051 gnd.n1094 9.3005
R20263 gnd.n5052 gnd.n1093 9.3005
R20264 gnd.n5055 gnd.n1092 9.3005
R20265 gnd.n5057 gnd.n1089 9.3005
R20266 gnd.n5060 gnd.n1088 9.3005
R20267 gnd.n5061 gnd.n1087 9.3005
R20268 gnd.n5064 gnd.n1086 9.3005
R20269 gnd.n5065 gnd.n1085 9.3005
R20270 gnd.n5068 gnd.n1084 9.3005
R20271 gnd.n5069 gnd.n1083 9.3005
R20272 gnd.n5072 gnd.n1082 9.3005
R20273 gnd.n5073 gnd.n1081 9.3005
R20274 gnd.n5076 gnd.n1080 9.3005
R20275 gnd.n5077 gnd.n1079 9.3005
R20276 gnd.n5080 gnd.n1078 9.3005
R20277 gnd.n5081 gnd.n1077 9.3005
R20278 gnd.n5084 gnd.n1076 9.3005
R20279 gnd.n5086 gnd.n1075 9.3005
R20280 gnd.n5087 gnd.n1074 9.3005
R20281 gnd.n5088 gnd.n1073 9.3005
R20282 gnd.n5089 gnd.n1072 9.3005
R20283 gnd.n5016 gnd.n1111 9.3005
R20284 gnd.n4974 gnd.n1133 9.3005
R20285 gnd.n4966 gnd.n1147 9.3005
R20286 gnd.n4965 gnd.n1148 9.3005
R20287 gnd.n4964 gnd.n1149 9.3005
R20288 gnd.n1169 gnd.n1150 9.3005
R20289 gnd.n4954 gnd.n1170 9.3005
R20290 gnd.n4953 gnd.n1171 9.3005
R20291 gnd.n4952 gnd.n1172 9.3005
R20292 gnd.n1188 gnd.n1173 9.3005
R20293 gnd.n4942 gnd.n1189 9.3005
R20294 gnd.n4941 gnd.n1190 9.3005
R20295 gnd.n4940 gnd.n1191 9.3005
R20296 gnd.n1209 gnd.n1192 9.3005
R20297 gnd.n4930 gnd.n1210 9.3005
R20298 gnd.n4929 gnd.n1211 9.3005
R20299 gnd.n4928 gnd.n1212 9.3005
R20300 gnd.n1229 gnd.n1213 9.3005
R20301 gnd.n4918 gnd.n1230 9.3005
R20302 gnd.n4917 gnd.n1231 9.3005
R20303 gnd.n4916 gnd.n1232 9.3005
R20304 gnd.n1250 gnd.n1233 9.3005
R20305 gnd.n4906 gnd.n1251 9.3005
R20306 gnd.n1260 gnd.n1253 9.3005
R20307 gnd.n4892 gnd.n1278 9.3005
R20308 gnd.n4891 gnd.n1279 9.3005
R20309 gnd.n4890 gnd.n1280 9.3005
R20310 gnd.n1298 gnd.n1281 9.3005
R20311 gnd.n4880 gnd.n1299 9.3005
R20312 gnd.n4879 gnd.n1300 9.3005
R20313 gnd.n4878 gnd.n1301 9.3005
R20314 gnd.n1317 gnd.n1302 9.3005
R20315 gnd.n4868 gnd.n1318 9.3005
R20316 gnd.n4867 gnd.n1319 9.3005
R20317 gnd.n4866 gnd.n1320 9.3005
R20318 gnd.n1338 gnd.n1321 9.3005
R20319 gnd.n4856 gnd.n1339 9.3005
R20320 gnd.n4855 gnd.n1340 9.3005
R20321 gnd.n4854 gnd.n1341 9.3005
R20322 gnd.n1358 gnd.n1342 9.3005
R20323 gnd.n4844 gnd.n1359 9.3005
R20324 gnd.n4843 gnd.n1360 9.3005
R20325 gnd.n4842 gnd.n1361 9.3005
R20326 gnd.n1378 gnd.n1362 9.3005
R20327 gnd.n4832 gnd.n4831 9.3005
R20328 gnd.n1146 gnd.n1145 9.3005
R20329 gnd.n4903 gnd.n1258 9.3005
R20330 gnd.n4903 gnd.n4902 9.3005
R20331 gnd.n2730 gnd.n2729 9.3005
R20332 gnd.n2731 gnd.n2720 9.3005
R20333 gnd.n2733 gnd.n2732 9.3005
R20334 gnd.n2718 gnd.n2717 9.3005
R20335 gnd.n2895 gnd.n2894 9.3005
R20336 gnd.n2896 gnd.n2716 9.3005
R20337 gnd.n2898 gnd.n2897 9.3005
R20338 gnd.n2714 gnd.n2713 9.3005
R20339 gnd.n2904 gnd.n2903 9.3005
R20340 gnd.n2905 gnd.n2712 9.3005
R20341 gnd.n2907 gnd.n2906 9.3005
R20342 gnd.n2722 gnd.n2721 9.3005
R20343 gnd.n2723 gnd.n966 9.3005
R20344 gnd.n6513 gnd.n965 9.3005
R20345 gnd.n6514 gnd.n964 9.3005
R20346 gnd.n6515 gnd.n963 9.3005
R20347 gnd.n962 gnd.n958 9.3005
R20348 gnd.n6521 gnd.n957 9.3005
R20349 gnd.n6522 gnd.n956 9.3005
R20350 gnd.n6523 gnd.n955 9.3005
R20351 gnd.n954 gnd.n950 9.3005
R20352 gnd.n6529 gnd.n949 9.3005
R20353 gnd.n6530 gnd.n948 9.3005
R20354 gnd.n6531 gnd.n947 9.3005
R20355 gnd.n946 gnd.n942 9.3005
R20356 gnd.n6537 gnd.n941 9.3005
R20357 gnd.n6538 gnd.n940 9.3005
R20358 gnd.n6539 gnd.n939 9.3005
R20359 gnd.n938 gnd.n934 9.3005
R20360 gnd.n6545 gnd.n933 9.3005
R20361 gnd.n6546 gnd.n932 9.3005
R20362 gnd.n6547 gnd.n931 9.3005
R20363 gnd.n930 gnd.n926 9.3005
R20364 gnd.n6553 gnd.n925 9.3005
R20365 gnd.n6554 gnd.n924 9.3005
R20366 gnd.n6555 gnd.n923 9.3005
R20367 gnd.n922 gnd.n918 9.3005
R20368 gnd.n6561 gnd.n917 9.3005
R20369 gnd.n6562 gnd.n916 9.3005
R20370 gnd.n6563 gnd.n915 9.3005
R20371 gnd.n914 gnd.n910 9.3005
R20372 gnd.n6569 gnd.n909 9.3005
R20373 gnd.n6570 gnd.n908 9.3005
R20374 gnd.n6571 gnd.n907 9.3005
R20375 gnd.n906 gnd.n902 9.3005
R20376 gnd.n6577 gnd.n901 9.3005
R20377 gnd.n6578 gnd.n900 9.3005
R20378 gnd.n6579 gnd.n899 9.3005
R20379 gnd.n898 gnd.n894 9.3005
R20380 gnd.n6585 gnd.n893 9.3005
R20381 gnd.n6586 gnd.n892 9.3005
R20382 gnd.n6587 gnd.n891 9.3005
R20383 gnd.n890 gnd.n886 9.3005
R20384 gnd.n6593 gnd.n885 9.3005
R20385 gnd.n6594 gnd.n884 9.3005
R20386 gnd.n6595 gnd.n883 9.3005
R20387 gnd.n882 gnd.n878 9.3005
R20388 gnd.n6601 gnd.n877 9.3005
R20389 gnd.n6602 gnd.n876 9.3005
R20390 gnd.n6603 gnd.n875 9.3005
R20391 gnd.n874 gnd.n870 9.3005
R20392 gnd.n6609 gnd.n869 9.3005
R20393 gnd.n6610 gnd.n868 9.3005
R20394 gnd.n6611 gnd.n867 9.3005
R20395 gnd.n866 gnd.n862 9.3005
R20396 gnd.n6617 gnd.n861 9.3005
R20397 gnd.n6618 gnd.n860 9.3005
R20398 gnd.n6619 gnd.n859 9.3005
R20399 gnd.n858 gnd.n854 9.3005
R20400 gnd.n6625 gnd.n853 9.3005
R20401 gnd.n6626 gnd.n852 9.3005
R20402 gnd.n6627 gnd.n851 9.3005
R20403 gnd.n850 gnd.n846 9.3005
R20404 gnd.n6633 gnd.n845 9.3005
R20405 gnd.n6634 gnd.n844 9.3005
R20406 gnd.n6635 gnd.n843 9.3005
R20407 gnd.n842 gnd.n838 9.3005
R20408 gnd.n6641 gnd.n837 9.3005
R20409 gnd.n6642 gnd.n836 9.3005
R20410 gnd.n6643 gnd.n835 9.3005
R20411 gnd.n834 gnd.n830 9.3005
R20412 gnd.n6649 gnd.n829 9.3005
R20413 gnd.n6650 gnd.n828 9.3005
R20414 gnd.n6651 gnd.n827 9.3005
R20415 gnd.n826 gnd.n822 9.3005
R20416 gnd.n6657 gnd.n821 9.3005
R20417 gnd.n6658 gnd.n820 9.3005
R20418 gnd.n6659 gnd.n819 9.3005
R20419 gnd.n818 gnd.n814 9.3005
R20420 gnd.n6665 gnd.n813 9.3005
R20421 gnd.n6666 gnd.n812 9.3005
R20422 gnd.n6667 gnd.n811 9.3005
R20423 gnd.n810 gnd.n806 9.3005
R20424 gnd.n6673 gnd.n805 9.3005
R20425 gnd.n6674 gnd.n804 9.3005
R20426 gnd.n6675 gnd.n803 9.3005
R20427 gnd.n2725 gnd.n2724 9.3005
R20428 gnd.n4181 gnd.n1972 9.3005
R20429 gnd.n3234 gnd.n3233 9.3005
R20430 gnd.n3235 gnd.n2405 9.3005
R20431 gnd.n3238 gnd.n3237 9.3005
R20432 gnd.n3236 gnd.n2406 9.3005
R20433 gnd.n2383 gnd.n2382 9.3005
R20434 gnd.n3264 gnd.n3263 9.3005
R20435 gnd.n3265 gnd.n2380 9.3005
R20436 gnd.n3268 gnd.n3267 9.3005
R20437 gnd.n3266 gnd.n2381 9.3005
R20438 gnd.n2359 gnd.n2358 9.3005
R20439 gnd.n3301 gnd.n3300 9.3005
R20440 gnd.n3302 gnd.n2356 9.3005
R20441 gnd.n3305 gnd.n3304 9.3005
R20442 gnd.n3303 gnd.n2357 9.3005
R20443 gnd.n2346 gnd.n2345 9.3005
R20444 gnd.n3428 gnd.n3427 9.3005
R20445 gnd.n3429 gnd.n2343 9.3005
R20446 gnd.n3433 gnd.n3432 9.3005
R20447 gnd.n3431 gnd.n2344 9.3005
R20448 gnd.n3430 gnd.n2332 9.3005
R20449 gnd.n2330 gnd.n2329 9.3005
R20450 gnd.n3456 gnd.n3455 9.3005
R20451 gnd.n3457 gnd.n2327 9.3005
R20452 gnd.n3460 gnd.n3459 9.3005
R20453 gnd.n3458 gnd.n2328 9.3005
R20454 gnd.n2311 gnd.n2310 9.3005
R20455 gnd.n3511 gnd.n3510 9.3005
R20456 gnd.n3512 gnd.n2308 9.3005
R20457 gnd.n3516 gnd.n3515 9.3005
R20458 gnd.n3514 gnd.n2309 9.3005
R20459 gnd.n3513 gnd.n2297 9.3005
R20460 gnd.n2295 gnd.n2294 9.3005
R20461 gnd.n3541 gnd.n3540 9.3005
R20462 gnd.n3542 gnd.n2293 9.3005
R20463 gnd.n3544 gnd.n3543 9.3005
R20464 gnd.n2268 gnd.n2266 9.3005
R20465 gnd.n3590 gnd.n3589 9.3005
R20466 gnd.n3588 gnd.n2267 9.3005
R20467 gnd.n3587 gnd.n3586 9.3005
R20468 gnd.n2244 gnd.n2242 9.3005
R20469 gnd.n3645 gnd.n3644 9.3005
R20470 gnd.n3643 gnd.n2243 9.3005
R20471 gnd.n3642 gnd.n3641 9.3005
R20472 gnd.n3640 gnd.n2245 9.3005
R20473 gnd.n3639 gnd.n3638 9.3005
R20474 gnd.n3637 gnd.n3628 9.3005
R20475 gnd.n3636 gnd.n3635 9.3005
R20476 gnd.n3634 gnd.n3629 9.3005
R20477 gnd.n3633 gnd.n3632 9.3005
R20478 gnd.n2181 gnd.n2180 9.3005
R20479 gnd.n3761 gnd.n3760 9.3005
R20480 gnd.n3762 gnd.n2179 9.3005
R20481 gnd.n3764 gnd.n3763 9.3005
R20482 gnd.n2160 gnd.n2159 9.3005
R20483 gnd.n3791 gnd.n3790 9.3005
R20484 gnd.n3792 gnd.n2157 9.3005
R20485 gnd.n3798 gnd.n3797 9.3005
R20486 gnd.n3796 gnd.n2158 9.3005
R20487 gnd.n3795 gnd.n3794 9.3005
R20488 gnd.n2131 gnd.n2130 9.3005
R20489 gnd.n3830 gnd.n3829 9.3005
R20490 gnd.n3831 gnd.n2128 9.3005
R20491 gnd.n3849 gnd.n3848 9.3005
R20492 gnd.n3847 gnd.n2129 9.3005
R20493 gnd.n3846 gnd.n3845 9.3005
R20494 gnd.n3844 gnd.n3832 9.3005
R20495 gnd.n3843 gnd.n3842 9.3005
R20496 gnd.n3841 gnd.n3835 9.3005
R20497 gnd.n3840 gnd.n3839 9.3005
R20498 gnd.n2041 gnd.n2040 9.3005
R20499 gnd.n4073 gnd.n4072 9.3005
R20500 gnd.n4074 gnd.n2039 9.3005
R20501 gnd.n4076 gnd.n4075 9.3005
R20502 gnd.n2028 gnd.n2027 9.3005
R20503 gnd.n4093 gnd.n4092 9.3005
R20504 gnd.n4094 gnd.n2026 9.3005
R20505 gnd.n4096 gnd.n4095 9.3005
R20506 gnd.n2014 gnd.n2013 9.3005
R20507 gnd.n4115 gnd.n4114 9.3005
R20508 gnd.n4116 gnd.n2011 9.3005
R20509 gnd.n4119 gnd.n4118 9.3005
R20510 gnd.n4117 gnd.n2012 9.3005
R20511 gnd.n2408 gnd.n2407 9.3005
R20512 gnd.n3156 gnd.n3155 9.3005
R20513 gnd.n2945 gnd.n2944 9.3005
R20514 gnd.n2943 gnd.n2941 9.3005
R20515 gnd.n2665 gnd.n2664 9.3005
R20516 gnd.n2999 gnd.n2998 9.3005
R20517 gnd.n3000 gnd.n2663 9.3005
R20518 gnd.n3002 gnd.n3001 9.3005
R20519 gnd.n2660 gnd.n2659 9.3005
R20520 gnd.n3014 gnd.n3013 9.3005
R20521 gnd.n3015 gnd.n2658 9.3005
R20522 gnd.n3017 gnd.n3016 9.3005
R20523 gnd.n2651 gnd.n2649 9.3005
R20524 gnd.n3053 gnd.n3052 9.3005
R20525 gnd.n3051 gnd.n2650 9.3005
R20526 gnd.n3050 gnd.n3049 9.3005
R20527 gnd.n3048 gnd.n2652 9.3005
R20528 gnd.n3047 gnd.n3046 9.3005
R20529 gnd.n3045 gnd.n2655 9.3005
R20530 gnd.n3044 gnd.n3043 9.3005
R20531 gnd.n3042 gnd.n2656 9.3005
R20532 gnd.n3041 gnd.n3040 9.3005
R20533 gnd.n2633 gnd.n2632 9.3005
R20534 gnd.n3130 gnd.n3129 9.3005
R20535 gnd.n3131 gnd.n2631 9.3005
R20536 gnd.n3134 gnd.n3133 9.3005
R20537 gnd.n3132 gnd.n2628 9.3005
R20538 gnd.n3145 gnd.n2627 9.3005
R20539 gnd.n3147 gnd.n3146 9.3005
R20540 gnd.n3205 gnd.n3204 9.3005
R20541 gnd.n3203 gnd.n3202 9.3005
R20542 gnd.n2565 gnd.n2564 9.3005
R20543 gnd.n3197 gnd.n3196 9.3005
R20544 gnd.n3195 gnd.n3194 9.3005
R20545 gnd.n2577 gnd.n2576 9.3005
R20546 gnd.n3189 gnd.n3188 9.3005
R20547 gnd.n3187 gnd.n3186 9.3005
R20548 gnd.n2588 gnd.n2587 9.3005
R20549 gnd.n3181 gnd.n3180 9.3005
R20550 gnd.n3179 gnd.n3178 9.3005
R20551 gnd.n2600 gnd.n2599 9.3005
R20552 gnd.n3173 gnd.n3172 9.3005
R20553 gnd.n3171 gnd.n3170 9.3005
R20554 gnd.n2611 gnd.n2610 9.3005
R20555 gnd.n3165 gnd.n3164 9.3005
R20556 gnd.n3163 gnd.n2624 9.3005
R20557 gnd.n3162 gnd.n3159 9.3005
R20558 gnd.n2560 gnd.n2555 9.3005
R20559 gnd.n3158 gnd.n3157 9.3005
R20560 gnd.n3151 gnd.n2626 9.3005
R20561 gnd.n3150 gnd.n2618 9.3005
R20562 gnd.n3167 gnd.n3166 9.3005
R20563 gnd.n3169 gnd.n3168 9.3005
R20564 gnd.n2604 gnd.n2603 9.3005
R20565 gnd.n3175 gnd.n3174 9.3005
R20566 gnd.n3177 gnd.n3176 9.3005
R20567 gnd.n2594 gnd.n2593 9.3005
R20568 gnd.n3183 gnd.n3182 9.3005
R20569 gnd.n3185 gnd.n3184 9.3005
R20570 gnd.n2581 gnd.n2580 9.3005
R20571 gnd.n3191 gnd.n3190 9.3005
R20572 gnd.n3193 gnd.n3192 9.3005
R20573 gnd.n2571 gnd.n2570 9.3005
R20574 gnd.n3199 gnd.n3198 9.3005
R20575 gnd.n3201 gnd.n3200 9.3005
R20576 gnd.n2559 gnd.n2558 9.3005
R20577 gnd.n3207 gnd.n3206 9.3005
R20578 gnd.n3209 gnd.n3208 9.3005
R20579 gnd.n3210 gnd.n2441 9.3005
R20580 gnd.n3213 gnd.n3212 9.3005
R20581 gnd.n3214 gnd.n2436 9.3005
R20582 gnd.n3216 gnd.n3215 9.3005
R20583 gnd.n3217 gnd.n2435 9.3005
R20584 gnd.n3219 gnd.n3218 9.3005
R20585 gnd.n2417 gnd.n2416 9.3005
R20586 gnd.n3225 gnd.n3224 9.3005
R20587 gnd.n3229 gnd.n3228 9.3005
R20588 gnd.n3227 gnd.n2415 9.3005
R20589 gnd.n2392 gnd.n2391 9.3005
R20590 gnd.n3255 gnd.n3254 9.3005
R20591 gnd.n3256 gnd.n2389 9.3005
R20592 gnd.n3259 gnd.n3258 9.3005
R20593 gnd.n3257 gnd.n2390 9.3005
R20594 gnd.n2366 gnd.n2365 9.3005
R20595 gnd.n3292 gnd.n3291 9.3005
R20596 gnd.n3293 gnd.n2363 9.3005
R20597 gnd.n3296 gnd.n3295 9.3005
R20598 gnd.n3294 gnd.n2364 9.3005
R20599 gnd.n2352 gnd.n2351 9.3005
R20600 gnd.n3420 gnd.n3419 9.3005
R20601 gnd.n3421 gnd.n2350 9.3005
R20602 gnd.n3423 gnd.n3422 9.3005
R20603 gnd.n2338 gnd.n2337 9.3005
R20604 gnd.n3438 gnd.n3437 9.3005
R20605 gnd.n3439 gnd.n2335 9.3005
R20606 gnd.n3449 gnd.n3448 9.3005
R20607 gnd.n3447 gnd.n2336 9.3005
R20608 gnd.n3446 gnd.n3445 9.3005
R20609 gnd.n3444 gnd.n3440 9.3005
R20610 gnd.n1542 gnd.n1540 9.3005
R20611 gnd.n4671 gnd.n4670 9.3005
R20612 gnd.n4669 gnd.n1541 9.3005
R20613 gnd.n4668 gnd.n4667 9.3005
R20614 gnd.n4666 gnd.n1543 9.3005
R20615 gnd.n4665 gnd.n4664 9.3005
R20616 gnd.n4663 gnd.n1547 9.3005
R20617 gnd.n4662 gnd.n4661 9.3005
R20618 gnd.n4660 gnd.n1548 9.3005
R20619 gnd.n4659 gnd.n4658 9.3005
R20620 gnd.n4657 gnd.n1552 9.3005
R20621 gnd.n4656 gnd.n4655 9.3005
R20622 gnd.n4654 gnd.n1553 9.3005
R20623 gnd.n4653 gnd.n4652 9.3005
R20624 gnd.n4651 gnd.n1557 9.3005
R20625 gnd.n4650 gnd.n4649 9.3005
R20626 gnd.n4648 gnd.n1558 9.3005
R20627 gnd.n4647 gnd.n4646 9.3005
R20628 gnd.n4645 gnd.n1562 9.3005
R20629 gnd.n4644 gnd.n4643 9.3005
R20630 gnd.n4642 gnd.n1563 9.3005
R20631 gnd.n4641 gnd.n4640 9.3005
R20632 gnd.n4639 gnd.n1567 9.3005
R20633 gnd.n4638 gnd.n4637 9.3005
R20634 gnd.n4636 gnd.n1568 9.3005
R20635 gnd.n4635 gnd.n4634 9.3005
R20636 gnd.n4633 gnd.n1572 9.3005
R20637 gnd.n4632 gnd.n4631 9.3005
R20638 gnd.n4630 gnd.n1573 9.3005
R20639 gnd.n4629 gnd.n4628 9.3005
R20640 gnd.n4627 gnd.n1577 9.3005
R20641 gnd.n4626 gnd.n4625 9.3005
R20642 gnd.n4624 gnd.n1578 9.3005
R20643 gnd.n4623 gnd.n4622 9.3005
R20644 gnd.n4621 gnd.n1582 9.3005
R20645 gnd.n4620 gnd.n4619 9.3005
R20646 gnd.n4618 gnd.n1583 9.3005
R20647 gnd.n4617 gnd.n4616 9.3005
R20648 gnd.n4615 gnd.n1587 9.3005
R20649 gnd.n4614 gnd.n4613 9.3005
R20650 gnd.n4612 gnd.n1588 9.3005
R20651 gnd.n4611 gnd.n4610 9.3005
R20652 gnd.n4609 gnd.n1592 9.3005
R20653 gnd.n4608 gnd.n4607 9.3005
R20654 gnd.n4606 gnd.n1593 9.3005
R20655 gnd.n4605 gnd.n4604 9.3005
R20656 gnd.n4603 gnd.n1597 9.3005
R20657 gnd.n4602 gnd.n4601 9.3005
R20658 gnd.n4600 gnd.n1598 9.3005
R20659 gnd.n4599 gnd.n4598 9.3005
R20660 gnd.n4597 gnd.n1602 9.3005
R20661 gnd.n4596 gnd.n4595 9.3005
R20662 gnd.n4594 gnd.n1603 9.3005
R20663 gnd.n4593 gnd.n4592 9.3005
R20664 gnd.n4591 gnd.n1607 9.3005
R20665 gnd.n4590 gnd.n4589 9.3005
R20666 gnd.n4588 gnd.n1608 9.3005
R20667 gnd.n4587 gnd.n4586 9.3005
R20668 gnd.n4585 gnd.n1612 9.3005
R20669 gnd.n3226 gnd.n2414 9.3005
R20670 gnd.n4582 gnd.n1613 9.3005
R20671 gnd.n4581 gnd.n4580 9.3005
R20672 gnd.n4579 gnd.n1617 9.3005
R20673 gnd.n4578 gnd.n4577 9.3005
R20674 gnd.n4576 gnd.n1618 9.3005
R20675 gnd.n4575 gnd.n4574 9.3005
R20676 gnd.n4584 gnd.n4583 9.3005
R20677 gnd.n4527 gnd.n4526 9.3005
R20678 gnd.n1665 gnd.n1664 9.3005
R20679 gnd.n4533 gnd.n4532 9.3005
R20680 gnd.n4535 gnd.n4534 9.3005
R20681 gnd.n1657 gnd.n1656 9.3005
R20682 gnd.n4541 gnd.n4540 9.3005
R20683 gnd.n4543 gnd.n4542 9.3005
R20684 gnd.n1649 gnd.n1648 9.3005
R20685 gnd.n4549 gnd.n4548 9.3005
R20686 gnd.n4551 gnd.n4550 9.3005
R20687 gnd.n1641 gnd.n1640 9.3005
R20688 gnd.n4557 gnd.n4556 9.3005
R20689 gnd.n4559 gnd.n4558 9.3005
R20690 gnd.n1633 gnd.n1632 9.3005
R20691 gnd.n4565 gnd.n4564 9.3005
R20692 gnd.n4567 gnd.n4566 9.3005
R20693 gnd.n1629 gnd.n1624 9.3005
R20694 gnd.n4525 gnd.n1674 9.3005
R20695 gnd.n1973 gnd.n1673 9.3005
R20696 gnd.n4572 gnd.n1622 9.3005
R20697 gnd.n4571 gnd.n4570 9.3005
R20698 gnd.n4569 gnd.n4568 9.3005
R20699 gnd.n1628 gnd.n1627 9.3005
R20700 gnd.n4563 gnd.n4562 9.3005
R20701 gnd.n4561 gnd.n4560 9.3005
R20702 gnd.n1637 gnd.n1636 9.3005
R20703 gnd.n4555 gnd.n4554 9.3005
R20704 gnd.n4553 gnd.n4552 9.3005
R20705 gnd.n1645 gnd.n1644 9.3005
R20706 gnd.n4547 gnd.n4546 9.3005
R20707 gnd.n4545 gnd.n4544 9.3005
R20708 gnd.n1653 gnd.n1652 9.3005
R20709 gnd.n4539 gnd.n4538 9.3005
R20710 gnd.n4537 gnd.n4536 9.3005
R20711 gnd.n1661 gnd.n1660 9.3005
R20712 gnd.n4531 gnd.n4530 9.3005
R20713 gnd.n4529 gnd.n4528 9.3005
R20714 gnd.n1998 gnd.n1671 9.3005
R20715 gnd.n1975 gnd.n1974 9.3005
R20716 gnd.n4183 gnd.n4182 9.3005
R20717 gnd.n4187 gnd.n4186 9.3005
R20718 gnd.n4188 gnd.n1968 9.3005
R20719 gnd.n4192 gnd.n4191 9.3005
R20720 gnd.n4193 gnd.n1967 9.3005
R20721 gnd.n4195 gnd.n4194 9.3005
R20722 gnd.n1964 gnd.n1963 9.3005
R20723 gnd.n4207 gnd.n4206 9.3005
R20724 gnd.n4208 gnd.n1962 9.3005
R20725 gnd.n4210 gnd.n4209 9.3005
R20726 gnd.n1956 gnd.n1954 9.3005
R20727 gnd.n4246 gnd.n4245 9.3005
R20728 gnd.n4244 gnd.n1955 9.3005
R20729 gnd.n4243 gnd.n4242 9.3005
R20730 gnd.n4241 gnd.n1957 9.3005
R20731 gnd.n4240 gnd.n4239 9.3005
R20732 gnd.n4238 gnd.n1960 9.3005
R20733 gnd.n4237 gnd.n4236 9.3005
R20734 gnd.n1940 gnd.n1939 9.3005
R20735 gnd.n4276 gnd.n4275 9.3005
R20736 gnd.n4277 gnd.n1937 9.3005
R20737 gnd.n4287 gnd.n4286 9.3005
R20738 gnd.n4285 gnd.n1938 9.3005
R20739 gnd.n4284 gnd.n4283 9.3005
R20740 gnd.n4282 gnd.n4278 9.3005
R20741 gnd.n4281 gnd.n4280 9.3005
R20742 gnd.n81 gnd.n79 9.3005
R20743 gnd.n4185 gnd.n1969 9.3005
R20744 gnd.t32 gnd.n5228 9.24152
R20745 gnd.n6481 gnd.t251 9.24152
R20746 gnd.t345 gnd.n1019 9.24152
R20747 gnd.n1152 gnd.t269 9.24152
R20748 gnd.n3120 gnd.t90 9.24152
R20749 gnd.n1965 gnd.t99 9.24152
R20750 gnd.n7609 gnd.t273 9.24152
R20751 gnd.t238 gnd.t32 8.92286
R20752 gnd.n4695 gnd.n4694 8.92286
R20753 gnd.n3529 gnd.n2303 8.92286
R20754 gnd.n3572 gnd.n2272 8.92286
R20755 gnd.t3 gnd.n2262 8.92286
R20756 gnd.n3683 gnd.t54 8.92286
R20757 gnd.n3694 gnd.n2205 8.92286
R20758 gnd.n3769 gnd.n3768 8.92286
R20759 gnd.n3868 gnd.n3867 8.92286
R20760 gnd.t248 gnd.n2096 8.92286
R20761 gnd.n6335 gnd.n6310 8.92171
R20762 gnd.n6303 gnd.n6278 8.92171
R20763 gnd.n6271 gnd.n6246 8.92171
R20764 gnd.n6240 gnd.n6215 8.92171
R20765 gnd.n6208 gnd.n6183 8.92171
R20766 gnd.n6176 gnd.n6151 8.92171
R20767 gnd.n6144 gnd.n6119 8.92171
R20768 gnd.n6113 gnd.n6088 8.92171
R20769 gnd.n3921 gnd.n3903 8.72777
R20770 gnd.t35 gnd.n5339 8.60421
R20771 gnd.n5291 gnd.n5275 8.43656
R20772 gnd.n46 gnd.n30 8.43656
R20773 gnd.n4708 gnd.t311 8.28555
R20774 gnd.n3451 gnd.t349 8.28555
R20775 gnd.n3463 gnd.t45 8.28555
R20776 gnd.n3478 gnd.n3477 8.28555
R20777 gnd.n3564 gnd.t4 8.28555
R20778 gnd.n3592 gnd.n2254 8.28555
R20779 gnd.n3673 gnd.n2219 8.28555
R20780 gnd.n2200 gnd.t40 8.28555
R20781 gnd.n3736 gnd.n2170 8.28555
R20782 gnd.n3726 gnd.t14 8.28555
R20783 gnd.n6336 gnd.n6308 8.14595
R20784 gnd.n6304 gnd.n6276 8.14595
R20785 gnd.n6272 gnd.n6244 8.14595
R20786 gnd.n6241 gnd.n6213 8.14595
R20787 gnd.n6209 gnd.n6181 8.14595
R20788 gnd.n6177 gnd.n6149 8.14595
R20789 gnd.n6145 gnd.n6117 8.14595
R20790 gnd.n6114 gnd.n6086 8.14595
R20791 gnd.n2942 gnd.n0 8.10675
R20792 gnd.n7683 gnd.n7682 8.10675
R20793 gnd.n6341 gnd.n6340 7.97301
R20794 gnd.n5832 gnd.t36 7.9669
R20795 gnd.n7683 gnd.n78 7.86902
R20796 gnd.n4525 gnd.n1673 7.75808
R20797 gnd.n3163 gnd.n3162 7.75808
R20798 gnd.n7459 gnd.n349 7.75808
R20799 gnd.n2804 gnd.n2803 7.75808
R20800 gnd.n2348 gnd.t245 7.64824
R20801 gnd.n4688 gnd.n1517 7.64824
R20802 gnd.n3477 gnd.n2315 7.64824
R20803 gnd.n3603 gnd.n2254 7.64824
R20804 gnd.n3673 gnd.n2218 7.64824
R20805 gnd.n3736 gnd.n3735 7.64824
R20806 gnd.n3859 gnd.n3858 7.64824
R20807 gnd.n5324 gnd.n5323 7.53171
R20808 gnd.t25 gnd.n5425 7.32958
R20809 gnd.n1487 gnd.n1486 7.30353
R20810 gnd.n3920 gnd.n3919 7.30353
R20811 gnd.n5734 gnd.n5733 7.01093
R20812 gnd.n5744 gnd.n5454 7.01093
R20813 gnd.n5743 gnd.n5457 7.01093
R20814 gnd.n5752 gnd.n5448 7.01093
R20815 gnd.n5756 gnd.n5755 7.01093
R20816 gnd.n5774 gnd.n5433 7.01093
R20817 gnd.n5773 gnd.n5436 7.01093
R20818 gnd.n5784 gnd.n5425 7.01093
R20819 gnd.n5426 gnd.n5414 7.01093
R20820 gnd.n5797 gnd.n5415 7.01093
R20821 gnd.n5808 gnd.n5407 7.01093
R20822 gnd.n5807 gnd.n5398 7.01093
R20823 gnd.n5400 gnd.n5382 7.01093
R20824 gnd.n5844 gnd.n5383 7.01093
R20825 gnd.n5833 gnd.n5832 7.01093
R20826 gnd.n5869 gnd.n5374 7.01093
R20827 gnd.n5880 gnd.n5879 7.01093
R20828 gnd.n5367 gnd.n5359 7.01093
R20829 gnd.n5909 gnd.n5347 7.01093
R20830 gnd.n5908 gnd.n5350 7.01093
R20831 gnd.n5919 gnd.n5339 7.01093
R20832 gnd.n5340 gnd.n5328 7.01093
R20833 gnd.n5930 gnd.n5329 7.01093
R20834 gnd.n5954 gnd.n5256 7.01093
R20835 gnd.n5953 gnd.n5247 7.01093
R20836 gnd.n5249 gnd.n5240 7.01093
R20837 gnd.n5976 gnd.n5975 7.01093
R20838 gnd.n5993 gnd.n5228 7.01093
R20839 gnd.n5992 gnd.n5231 7.01093
R20840 gnd.n6006 gnd.n5220 7.01093
R20841 gnd.n5221 gnd.n5210 7.01093
R20842 gnd.n6016 gnd.n5212 7.01093
R20843 gnd.n6049 gnd.n6048 7.01093
R20844 gnd.n6065 gnd.n6064 7.01093
R20845 gnd.n5191 gnd.n968 7.01093
R20846 gnd.n6508 gnd.n970 7.01093
R20847 gnd.n6029 gnd.n979 7.01093
R20848 gnd.n6502 gnd.n6501 7.01093
R20849 gnd.n6495 gnd.n990 7.01093
R20850 gnd.n6494 gnd.n993 7.01093
R20851 gnd.n6373 gnd.n1002 7.01093
R20852 gnd.n6488 gnd.n6487 7.01093
R20853 gnd.n6354 gnd.n1005 7.01093
R20854 gnd.n6481 gnd.n1016 7.01093
R20855 gnd.n6480 gnd.n1019 7.01093
R20856 gnd.n6384 gnd.n1027 7.01093
R20857 gnd.n6474 gnd.n6473 7.01093
R20858 gnd.n3529 gnd.n3528 7.01093
R20859 gnd.n3546 gnd.n2272 7.01093
R20860 gnd.n3573 gnd.t3 7.01093
R20861 gnd.t54 gnd.n3682 7.01093
R20862 gnd.n3694 gnd.n3693 7.01093
R20863 gnd.n3769 gnd.n2175 7.01093
R20864 gnd.n3868 gnd.n2110 7.01093
R20865 gnd.n3874 gnd.t248 7.01093
R20866 gnd.n5415 gnd.t28 6.69227
R20867 gnd.n5975 gnd.t238 6.69227
R20868 gnd.t34 gnd.n6365 6.69227
R20869 gnd.n4944 gnd.t102 6.69227
R20870 gnd.n3038 gnd.t104 6.69227
R20871 gnd.n3451 gnd.t231 6.69227
R20872 gnd.n3714 gnd.t19 6.69227
R20873 gnd.n4212 gnd.t69 6.69227
R20874 gnd.n7438 gnd.t73 6.69227
R20875 gnd.n4053 gnd.n4052 6.5566
R20876 gnd.n3314 gnd.n3313 6.5566
R20877 gnd.n4720 gnd.n4716 6.5566
R20878 gnd.n3931 gnd.n3930 6.5566
R20879 gnd.n6509 gnd.n6508 6.37362
R20880 gnd.n4681 gnd.n4680 6.37362
R20881 gnd.n3470 gnd.n2321 6.37362
R20882 gnd.n3493 gnd.t233 6.37362
R20883 gnd.n3611 gnd.n2248 6.37362
R20884 gnd.n3623 gnd.n2235 6.37362
R20885 gnd.n3700 gnd.t0 6.37362
R20886 gnd.n3803 gnd.n3802 6.37362
R20887 gnd.n3818 gnd.n2140 6.37362
R20888 gnd.n3150 gnd.n2617 6.20656
R20889 gnd.n1998 gnd.n1670 6.20656
R20890 gnd.n5868 gnd.t15 6.05496
R20891 gnd.n5867 gnd.t27 6.05496
R20892 gnd.t63 gnd.n5340 6.05496
R20893 gnd.t22 gnd.n5204 6.05496
R20894 gnd.n3019 gnd.t97 6.05496
R20895 gnd.n4234 gnd.t77 6.05496
R20896 gnd.n6338 gnd.n6308 5.81868
R20897 gnd.n6306 gnd.n6276 5.81868
R20898 gnd.n6274 gnd.n6244 5.81868
R20899 gnd.n6243 gnd.n6213 5.81868
R20900 gnd.n6211 gnd.n6181 5.81868
R20901 gnd.n6179 gnd.n6149 5.81868
R20902 gnd.n6147 gnd.n6117 5.81868
R20903 gnd.n6116 gnd.n6086 5.81868
R20904 gnd.n3408 gnd.n3407 5.73631
R20905 gnd.n3425 gnd.n2348 5.73631
R20906 gnd.n3492 gnd.n2286 5.73631
R20907 gnd.n2287 gnd.n2278 5.73631
R20908 gnd.n2201 gnd.n2190 5.73631
R20909 gnd.n3701 gnd.n2193 5.73631
R20910 gnd.n3889 gnd.n2106 5.73631
R20911 gnd.n3899 gnd.n2096 5.73631
R20912 gnd.n4057 gnd.n1750 5.62001
R20913 gnd.n4782 gnd.n1429 5.62001
R20914 gnd.n4782 gnd.n1430 5.62001
R20915 gnd.n3926 gnd.n1750 5.62001
R20916 gnd.n5552 gnd.n5551 5.4308
R20917 gnd.n5171 gnd.n5169 5.4308
R20918 gnd.n5329 gnd.t37 5.41765
R20919 gnd.t24 gnd.n5964 5.41765
R20920 gnd.n6050 gnd.t57 5.41765
R20921 gnd.t107 gnd.n2673 5.41765
R20922 gnd.t8 gnd.n4673 5.41765
R20923 gnd.n3800 gnd.t10 5.41765
R20924 gnd.n4313 gnd.t75 5.41765
R20925 gnd.n2842 gnd.n1194 5.09899
R20926 gnd.n4938 gnd.n1197 5.09899
R20927 gnd.n2851 gnd.n1204 5.09899
R20928 gnd.n4932 gnd.n1207 5.09899
R20929 gnd.n2891 gnd.n2890 5.09899
R20930 gnd.n4926 gnd.n1217 5.09899
R20931 gnd.n2884 gnd.n1224 5.09899
R20932 gnd.n4920 gnd.n1227 5.09899
R20933 gnd.n2878 gnd.n1235 5.09899
R20934 gnd.n4914 gnd.n1238 5.09899
R20935 gnd.n2872 gnd.n1245 5.09899
R20936 gnd.n4908 gnd.n1248 5.09899
R20937 gnd.n2920 gnd.n2709 5.09899
R20938 gnd.n2923 gnd.n2697 5.09899
R20939 gnd.n2934 gnd.n2699 5.09899
R20940 gnd.n2931 gnd.n2703 5.09899
R20941 gnd.n2948 gnd.n2679 5.09899
R20942 gnd.n2961 gnd.n2682 5.09899
R20943 gnd.n2968 gnd.n2673 5.09899
R20944 gnd.n2967 gnd.n2667 5.09899
R20945 gnd.n2996 gnd.n2995 5.09899
R20946 gnd.n4900 gnd.n1265 5.09899
R20947 gnd.n3004 gnd.n1274 5.09899
R20948 gnd.n3011 gnd.n1283 5.09899
R20949 gnd.n4888 gnd.n1286 5.09899
R20950 gnd.n3019 gnd.n1293 5.09899
R20951 gnd.n4882 gnd.n1296 5.09899
R20952 gnd.n3056 gnd.n3055 5.09899
R20953 gnd.n4876 gnd.n1306 5.09899
R20954 gnd.n3026 gnd.n1313 5.09899
R20955 gnd.n3032 gnd.n1323 5.09899
R20956 gnd.n4864 gnd.n1326 5.09899
R20957 gnd.n3038 gnd.n1333 5.09899
R20958 gnd.n4858 gnd.n1336 5.09899
R20959 gnd.n3121 gnd.n3120 5.09899
R20960 gnd.n4852 gnd.n1346 5.09899
R20961 gnd.n3127 gnd.n1353 5.09899
R20962 gnd.n4846 gnd.n1356 5.09899
R20963 gnd.n3136 gnd.n1364 5.09899
R20964 gnd.n4840 gnd.n1367 5.09899
R20965 gnd.n3143 gnd.n1373 5.09899
R20966 gnd.n4834 gnd.n1376 5.09899
R20967 gnd.n3393 gnd.t349 5.09899
R20968 gnd.n3463 gnd.n2324 5.09899
R20969 gnd.n4674 gnd.n1535 5.09899
R20970 gnd.n3518 gnd.t62 5.09899
R20971 gnd.n3535 gnd.t233 5.09899
R20972 gnd.n3648 gnd.n2239 5.09899
R20973 gnd.n3657 gnd.n2232 5.09899
R20974 gnd.t0 gnd.n2183 5.09899
R20975 gnd.n3766 gnd.t21 5.09899
R20976 gnd.n3810 gnd.n3809 5.09899
R20977 gnd.n3726 gnd.n3725 5.09899
R20978 gnd.n4399 gnd.n1786 5.09899
R20979 gnd.n1970 gnd.n1788 5.09899
R20980 gnd.n4391 gnd.n1796 5.09899
R20981 gnd.n4189 gnd.n1798 5.09899
R20982 gnd.n4385 gnd.n1811 5.09899
R20983 gnd.n4197 gnd.n1814 5.09899
R20984 gnd.n4379 gnd.n1824 5.09899
R20985 gnd.n4204 gnd.n1965 5.09899
R20986 gnd.n4373 gnd.n1834 5.09899
R20987 gnd.n4212 gnd.n1837 5.09899
R20988 gnd.n4367 gnd.n1844 5.09899
R20989 gnd.n4248 gnd.n1847 5.09899
R20990 gnd.n4219 gnd.n1857 5.09899
R20991 gnd.n4355 gnd.n1864 5.09899
R20992 gnd.n4225 gnd.n4224 5.09899
R20993 gnd.n4349 gnd.n1874 5.09899
R20994 gnd.n4234 gnd.n1877 5.09899
R20995 gnd.n4343 gnd.n1884 5.09899
R20996 gnd.n4273 gnd.n1887 5.09899
R20997 gnd.n4289 gnd.n1897 5.09899
R20998 gnd.n4331 gnd.n1904 5.09899
R20999 gnd.n4327 gnd.n1909 5.09899
R21000 gnd.n4326 gnd.n1912 5.09899
R21001 gnd.n4313 gnd.n1927 5.09899
R21002 gnd.n4319 gnd.n4318 5.09899
R21003 gnd.n4307 gnd.n1924 5.09899
R21004 gnd.n7677 gnd.n85 5.09899
R21005 gnd.n381 gnd.n87 5.09899
R21006 gnd.n7374 gnd.n7369 5.09899
R21007 gnd.n7669 gnd.n102 5.09899
R21008 gnd.n7380 gnd.n105 5.09899
R21009 gnd.n7663 gnd.n114 5.09899
R21010 gnd.n7388 gnd.n374 5.09899
R21011 gnd.n7657 gnd.n123 5.09899
R21012 gnd.n7394 gnd.n371 5.09899
R21013 gnd.n7651 gnd.n132 5.09899
R21014 gnd.n7402 gnd.n135 5.09899
R21015 gnd.n7645 gnd.n143 5.09899
R21016 gnd.n7408 gnd.n146 5.09899
R21017 gnd.n7639 gnd.n153 5.09899
R21018 gnd.n7417 gnd.n362 5.09899
R21019 gnd.n7633 gnd.n163 5.09899
R21020 gnd.n6336 gnd.n6335 5.04292
R21021 gnd.n6304 gnd.n6303 5.04292
R21022 gnd.n6272 gnd.n6271 5.04292
R21023 gnd.n6241 gnd.n6240 5.04292
R21024 gnd.n6209 gnd.n6208 5.04292
R21025 gnd.n6177 gnd.n6176 5.04292
R21026 gnd.n6145 gnd.n6144 5.04292
R21027 gnd.n6114 gnd.n6113 5.04292
R21028 gnd.t26 gnd.n5890 4.78034
R21029 gnd.n6006 gnd.t31 4.78034
R21030 gnd.n2872 gnd.t134 4.78034
R21031 gnd.n4894 gnd.t150 4.78034
R21032 gnd.t38 gnd.n2386 4.78034
R21033 gnd.n4089 gnd.t234 4.78034
R21034 gnd.n4337 gnd.t118 4.78034
R21035 gnd.n7663 gnd.t79 4.78034
R21036 gnd.n5864 gnd.n5863 4.74817
R21037 gnd.n5859 gnd.n5858 4.74817
R21038 gnd.n5855 gnd.n5854 4.74817
R21039 gnd.n5851 gnd.n5326 4.74817
R21040 gnd.n5863 gnd.n5862 4.74817
R21041 gnd.n5861 gnd.n5859 4.74817
R21042 gnd.n5857 gnd.n5855 4.74817
R21043 gnd.n5853 gnd.n5851 4.74817
R21044 gnd.n4329 gnd.n98 4.74817
R21045 gnd.n4316 gnd.n96 4.74817
R21046 gnd.n7675 gnd.n91 4.74817
R21047 gnd.n7673 gnd.n92 4.74817
R21048 gnd.n1908 gnd.n98 4.74817
R21049 gnd.n1926 gnd.n96 4.74817
R21050 gnd.n4315 gnd.n91 4.74817
R21051 gnd.n7674 gnd.n7673 4.74817
R21052 gnd.n2918 gnd.n2917 4.74817
R21053 gnd.n2912 gnd.n2908 4.74817
R21054 gnd.n2910 gnd.n2671 4.74817
R21055 gnd.n2972 gnd.n2971 4.74817
R21056 gnd.n2992 gnd.n2991 4.74817
R21057 gnd.n4266 gnd.n1915 4.74817
R21058 gnd.n4323 gnd.n4322 4.74817
R21059 gnd.n1920 gnd.n1916 4.74817
R21060 gnd.n1918 gnd.n384 4.74817
R21061 gnd.n7366 gnd.n7365 4.74817
R21062 gnd.n4268 gnd.n4266 4.74817
R21063 gnd.n4324 gnd.n4323 4.74817
R21064 gnd.n4321 gnd.n1916 4.74817
R21065 gnd.n1919 gnd.n1918 4.74817
R21066 gnd.n7367 gnd.n7366 4.74817
R21067 gnd.n4905 gnd.n4904 4.74817
R21068 gnd.n2677 gnd.n1257 4.74817
R21069 gnd.n2964 gnd.n1256 4.74817
R21070 gnd.n1259 gnd.n1255 4.74817
R21071 gnd.n4904 gnd.n1252 4.74817
R21072 gnd.n2702 gnd.n1257 4.74817
R21073 gnd.n2678 gnd.n1256 4.74817
R21074 gnd.n2965 gnd.n1255 4.74817
R21075 gnd.n2917 gnd.n2916 4.74817
R21076 gnd.n2915 gnd.n2908 4.74817
R21077 gnd.n2911 gnd.n2910 4.74817
R21078 gnd.n2971 gnd.n2970 4.74817
R21079 gnd.n2993 gnd.n2992 4.74817
R21080 gnd.n5323 gnd.n5322 4.74296
R21081 gnd.n78 gnd.n77 4.74296
R21082 gnd.n5291 gnd.n5290 4.7074
R21083 gnd.n5307 gnd.n5306 4.7074
R21084 gnd.n46 gnd.n45 4.7074
R21085 gnd.n62 gnd.n61 4.7074
R21086 gnd.n5323 gnd.n5307 4.65959
R21087 gnd.n78 gnd.n62 4.65959
R21088 gnd.n4467 gnd.n1752 4.6132
R21089 gnd.n4783 gnd.n1428 4.6132
R21090 gnd.n4709 gnd.n1491 4.46168
R21091 gnd.n4701 gnd.n1502 4.46168
R21092 gnd.n4695 gnd.t298 4.46168
R21093 gnd.n3536 gnd.n3535 4.46168
R21094 gnd.n3563 gnd.n2281 4.46168
R21095 gnd.n3708 gnd.n2198 4.46168
R21096 gnd.n3758 gnd.n2183 4.46168
R21097 gnd.n3836 gnd.n2098 4.46168
R21098 gnd.n3916 gnd.n3903 4.46111
R21099 gnd.n6321 gnd.n6317 4.38594
R21100 gnd.n6289 gnd.n6285 4.38594
R21101 gnd.n6257 gnd.n6253 4.38594
R21102 gnd.n6226 gnd.n6222 4.38594
R21103 gnd.n6194 gnd.n6190 4.38594
R21104 gnd.n6162 gnd.n6158 4.38594
R21105 gnd.n6130 gnd.n6126 4.38594
R21106 gnd.n6099 gnd.n6095 4.38594
R21107 gnd.n6332 gnd.n6310 4.26717
R21108 gnd.n6300 gnd.n6278 4.26717
R21109 gnd.n6268 gnd.n6246 4.26717
R21110 gnd.n6237 gnd.n6215 4.26717
R21111 gnd.n6205 gnd.n6183 4.26717
R21112 gnd.n6173 gnd.n6151 4.26717
R21113 gnd.n6141 gnd.n6119 4.26717
R21114 gnd.n6110 gnd.n6088 4.26717
R21115 gnd.t33 gnd.n5821 4.14303
R21116 gnd.t29 gnd.n970 4.14303
R21117 gnd.n2851 gnd.t154 4.14303
R21118 gnd.n4870 gnd.t124 4.14303
R21119 gnd.t281 gnd.n1367 4.14303
R21120 gnd.t265 gnd.n1796 4.14303
R21121 gnd.n4361 gnd.t88 4.14303
R21122 gnd.n7639 gnd.t121 4.14303
R21123 gnd.n6340 gnd.n6339 4.08274
R21124 gnd.n4052 gnd.n4051 4.05904
R21125 gnd.n3315 gnd.n3314 4.05904
R21126 gnd.n4723 gnd.n4716 4.05904
R21127 gnd.n3932 gnd.n3931 4.05904
R21128 gnd.n15 gnd.n7 3.99943
R21129 gnd.n3383 gnd.n3382 3.82437
R21130 gnd.t59 gnd.n2313 3.82437
R21131 gnd.n3583 gnd.n2269 3.82437
R21132 gnd.n3666 gnd.n3665 3.82437
R21133 gnd.n3787 gnd.t2 3.82437
R21134 gnd.n3826 gnd.n3825 3.82437
R21135 gnd.t259 gnd.n2091 3.82437
R21136 gnd.n5325 gnd.n5324 3.81325
R21137 gnd.n5307 gnd.n5291 3.72967
R21138 gnd.n62 gnd.n46 3.72967
R21139 gnd.n6340 gnd.n6212 3.70378
R21140 gnd.n15 gnd.n14 3.60163
R21141 gnd.n4779 gnd.n1433 3.50571
R21142 gnd.n4060 gnd.n2069 3.50571
R21143 gnd.n6331 gnd.n6312 3.49141
R21144 gnd.n6299 gnd.n6280 3.49141
R21145 gnd.n6267 gnd.n6248 3.49141
R21146 gnd.n6236 gnd.n6217 3.49141
R21147 gnd.n6204 gnd.n6185 3.49141
R21148 gnd.n6172 gnd.n6153 3.49141
R21149 gnd.n6140 gnd.n6121 3.49141
R21150 gnd.n6109 gnd.n6090 3.49141
R21151 gnd.n4485 gnd.n4484 3.29747
R21152 gnd.n4484 gnd.n4483 3.29747
R21153 gnd.n7568 gnd.n7565 3.29747
R21154 gnd.n7569 gnd.n7568 3.29747
R21155 gnd.n5057 gnd.n5056 3.29747
R21156 gnd.n5056 gnd.n5055 3.29747
R21157 gnd.n4799 gnd.n4798 3.29747
R21158 gnd.n4798 gnd.n4797 3.29747
R21159 gnd.n3416 gnd.t262 3.18706
R21160 gnd.n3389 gnd.n1509 3.18706
R21161 gnd.n3519 gnd.n3518 3.18706
R21162 gnd.t4 gnd.n3563 3.18706
R21163 gnd.n3574 gnd.n3573 3.18706
R21164 gnd.n3682 gnd.n3680 3.18706
R21165 gnd.n3708 gnd.t40 3.18706
R21166 gnd.n3767 gnd.n3766 3.18706
R21167 gnd.n3852 gnd.n3851 3.18706
R21168 gnd.n3867 gnd.t295 3.18706
R21169 gnd.n5822 gnd.t33 2.8684
R21170 gnd.n3406 gnd.t65 2.8684
R21171 gnd.n3874 gnd.t12 2.8684
R21172 gnd.n5308 gnd.t125 2.82907
R21173 gnd.n5308 gnd.t209 2.82907
R21174 gnd.n5310 gnd.t98 2.82907
R21175 gnd.n5310 gnd.t145 2.82907
R21176 gnd.n5312 gnd.t164 2.82907
R21177 gnd.n5312 gnd.t151 2.82907
R21178 gnd.n5314 gnd.t149 2.82907
R21179 gnd.n5314 gnd.t137 2.82907
R21180 gnd.n5316 gnd.t157 2.82907
R21181 gnd.n5316 gnd.t192 2.82907
R21182 gnd.n5318 gnd.t87 2.82907
R21183 gnd.n5318 gnd.t180 2.82907
R21184 gnd.n5320 gnd.t217 2.82907
R21185 gnd.n5320 gnd.t155 2.82907
R21186 gnd.n5261 gnd.t158 2.82907
R21187 gnd.n5261 gnd.t179 2.82907
R21188 gnd.n5263 gnd.t187 2.82907
R21189 gnd.n5263 gnd.t127 2.82907
R21190 gnd.n5265 gnd.t175 2.82907
R21191 gnd.n5265 gnd.t169 2.82907
R21192 gnd.n5267 gnd.t223 2.82907
R21193 gnd.n5267 gnd.t211 2.82907
R21194 gnd.n5269 gnd.t135 2.82907
R21195 gnd.n5269 gnd.t184 2.82907
R21196 gnd.n5271 gnd.t204 2.82907
R21197 gnd.n5271 gnd.t85 2.82907
R21198 gnd.n5273 gnd.t103 2.82907
R21199 gnd.n5273 gnd.t177 2.82907
R21200 gnd.n5276 gnd.t226 2.82907
R21201 gnd.n5276 gnd.t105 2.82907
R21202 gnd.n5278 gnd.t106 2.82907
R21203 gnd.n5278 gnd.t83 2.82907
R21204 gnd.n5280 gnd.t188 2.82907
R21205 gnd.n5280 gnd.t227 2.82907
R21206 gnd.n5282 gnd.t221 2.82907
R21207 gnd.n5282 gnd.t108 2.82907
R21208 gnd.n5284 gnd.t212 2.82907
R21209 gnd.n5284 gnd.t189 2.82907
R21210 gnd.n5286 gnd.t190 2.82907
R21211 gnd.n5286 gnd.t220 2.82907
R21212 gnd.n5288 gnd.t224 2.82907
R21213 gnd.n5288 gnd.t205 2.82907
R21214 gnd.n5292 gnd.t171 2.82907
R21215 gnd.n5292 gnd.t128 2.82907
R21216 gnd.n5294 gnd.t156 2.82907
R21217 gnd.n5294 gnd.t195 2.82907
R21218 gnd.n5296 gnd.t219 2.82907
R21219 gnd.n5296 gnd.t203 2.82907
R21220 gnd.n5298 gnd.t201 2.82907
R21221 gnd.n5298 gnd.t183 2.82907
R21222 gnd.n5300 gnd.t208 2.82907
R21223 gnd.n5300 gnd.t117 2.82907
R21224 gnd.n5302 gnd.t144 2.82907
R21225 gnd.n5302 gnd.t92 2.82907
R21226 gnd.n5304 gnd.t133 2.82907
R21227 gnd.n5304 gnd.t207 2.82907
R21228 gnd.n75 gnd.t122 2.82907
R21229 gnd.n75 gnd.t176 2.82907
R21230 gnd.n73 gnd.t143 2.82907
R21231 gnd.n73 gnd.t185 2.82907
R21232 gnd.n71 gnd.t160 2.82907
R21233 gnd.n71 gnd.t136 2.82907
R21234 gnd.n69 gnd.t93 2.82907
R21235 gnd.n69 gnd.t114 2.82907
R21236 gnd.n67 gnd.t119 2.82907
R21237 gnd.n67 gnd.t141 2.82907
R21238 gnd.n65 gnd.t111 2.82907
R21239 gnd.n65 gnd.t202 2.82907
R21240 gnd.n63 gnd.t170 2.82907
R21241 gnd.n63 gnd.t89 2.82907
R21242 gnd.n28 gnd.t213 2.82907
R21243 gnd.n28 gnd.t138 2.82907
R21244 gnd.n26 gnd.t130 2.82907
R21245 gnd.n26 gnd.t95 2.82907
R21246 gnd.n24 gnd.t228 2.82907
R21247 gnd.n24 gnd.t123 2.82907
R21248 gnd.n22 gnd.t101 2.82907
R21249 gnd.n22 gnd.t120 2.82907
R21250 gnd.n20 gnd.t200 2.82907
R21251 gnd.n20 gnd.t165 2.82907
R21252 gnd.n18 gnd.t153 2.82907
R21253 gnd.n18 gnd.t81 2.82907
R21254 gnd.n16 gnd.t193 2.82907
R21255 gnd.n16 gnd.t142 2.82907
R21256 gnd.n43 gnd.t182 2.82907
R21257 gnd.n43 gnd.t197 2.82907
R21258 gnd.n41 gnd.t198 2.82907
R21259 gnd.n41 gnd.t174 2.82907
R21260 gnd.n39 gnd.t172 2.82907
R21261 gnd.n39 gnd.t80 2.82907
R21262 gnd.n37 gnd.t76 2.82907
R21263 gnd.n37 gnd.t196 2.82907
R21264 gnd.n35 gnd.t206 2.82907
R21265 gnd.n35 gnd.t215 2.82907
R21266 gnd.n33 gnd.t214 2.82907
R21267 gnd.n33 gnd.t78 2.82907
R21268 gnd.n31 gnd.t70 2.82907
R21269 gnd.n31 gnd.t96 2.82907
R21270 gnd.n59 gnd.t168 2.82907
R21271 gnd.n59 gnd.t74 2.82907
R21272 gnd.n57 gnd.t194 2.82907
R21273 gnd.n57 gnd.t109 2.82907
R21274 gnd.n55 gnd.t216 2.82907
R21275 gnd.n55 gnd.t181 2.82907
R21276 gnd.n53 gnd.t152 2.82907
R21277 gnd.n53 gnd.t166 2.82907
R21278 gnd.n51 gnd.t167 2.82907
R21279 gnd.n51 gnd.t186 2.82907
R21280 gnd.n49 gnd.t161 2.82907
R21281 gnd.n49 gnd.t126 2.82907
R21282 gnd.n47 gnd.t225 2.82907
R21283 gnd.n47 gnd.t146 2.82907
R21284 gnd.n6328 gnd.n6327 2.71565
R21285 gnd.n6296 gnd.n6295 2.71565
R21286 gnd.n6264 gnd.n6263 2.71565
R21287 gnd.n6233 gnd.n6232 2.71565
R21288 gnd.n6201 gnd.n6200 2.71565
R21289 gnd.n6169 gnd.n6168 2.71565
R21290 gnd.n6137 gnd.n6136 2.71565
R21291 gnd.n6106 gnd.n6105 2.71565
R21292 gnd.n4702 gnd.t245 2.54975
R21293 gnd.n3435 gnd.t298 2.54975
R21294 gnd.n3393 gnd.n3390 2.54975
R21295 gnd.t45 gnd.n3462 2.54975
R21296 gnd.n3501 gnd.n3500 2.54975
R21297 gnd.n3593 gnd.n2262 2.54975
R21298 gnd.n3683 gnd.n2213 2.54975
R21299 gnd.n3779 gnd.n3778 2.54975
R21300 gnd.t14 gnd.n2148 2.54975
R21301 gnd.n3715 gnd.n2125 2.54975
R21302 gnd.t358 gnd.n3880 2.54975
R21303 gnd.n5863 gnd.n5325 2.27742
R21304 gnd.n5859 gnd.n5325 2.27742
R21305 gnd.n5855 gnd.n5325 2.27742
R21306 gnd.n5851 gnd.n5325 2.27742
R21307 gnd.n7672 gnd.n98 2.27742
R21308 gnd.n7672 gnd.n96 2.27742
R21309 gnd.n7672 gnd.n91 2.27742
R21310 gnd.n7673 gnd.n7672 2.27742
R21311 gnd.n4266 gnd.n95 2.27742
R21312 gnd.n4323 gnd.n95 2.27742
R21313 gnd.n1916 gnd.n95 2.27742
R21314 gnd.n1918 gnd.n95 2.27742
R21315 gnd.n7366 gnd.n95 2.27742
R21316 gnd.n4904 gnd.n4903 2.27742
R21317 gnd.n4903 gnd.n1257 2.27742
R21318 gnd.n4903 gnd.n1256 2.27742
R21319 gnd.n4903 gnd.n1255 2.27742
R21320 gnd.n2917 gnd.n1254 2.27742
R21321 gnd.n2908 gnd.n1254 2.27742
R21322 gnd.n2910 gnd.n1254 2.27742
R21323 gnd.n2971 gnd.n1254 2.27742
R21324 gnd.n2992 gnd.n1254 2.27742
R21325 gnd.t317 gnd.n5743 2.23109
R21326 gnd.n5891 gnd.t26 2.23109
R21327 gnd.t41 gnd.n2281 2.23109
R21328 gnd.t48 gnd.n2198 2.23109
R21329 gnd.n6324 gnd.n6314 1.93989
R21330 gnd.n6292 gnd.n6282 1.93989
R21331 gnd.n6260 gnd.n6250 1.93989
R21332 gnd.n6229 gnd.n6219 1.93989
R21333 gnd.n6197 gnd.n6187 1.93989
R21334 gnd.n6165 gnd.n6155 1.93989
R21335 gnd.n6133 gnd.n6123 1.93989
R21336 gnd.n6102 gnd.n6092 1.93989
R21337 gnd.n3408 gnd.t311 1.91244
R21338 gnd.n4687 gnd.n1519 1.91244
R21339 gnd.n3508 gnd.n3507 1.91244
R21340 gnd.n3602 gnd.n2257 1.91244
R21341 gnd.t7 gnd.n3583 1.91244
R21342 gnd.n3666 gnd.t6 1.91244
R21343 gnd.n2226 gnd.n2225 1.91244
R21344 gnd.n3788 gnd.n2162 1.91244
R21345 gnd.n3827 gnd.n2120 1.91244
R21346 gnd.n3881 gnd.t358 1.91244
R21347 gnd.n5756 gnd.t52 1.59378
R21348 gnd.n5965 gnd.t24 1.59378
R21349 gnd.n6039 gnd.t57 1.59378
R21350 gnd.t231 gnd.n1517 1.59378
R21351 gnd.t55 gnd.n2303 1.59378
R21352 gnd.n3768 gnd.t46 1.59378
R21353 gnd.n3858 gnd.t19 1.59378
R21354 gnd.n3415 gnd.n3414 1.27512
R21355 gnd.t241 gnd.n4701 1.27512
R21356 gnd.n2341 gnd.n2340 1.27512
R21357 gnd.n3382 gnd.t5 1.27512
R21358 gnd.n3526 gnd.n2298 1.27512
R21359 gnd.n3547 gnd.n2291 1.27512
R21360 gnd.n3692 gnd.n3691 1.27512
R21361 gnd.n3757 gnd.n2184 1.27512
R21362 gnd.t1 gnd.n3826 1.27512
R21363 gnd.n3883 gnd.n3882 1.27512
R21364 gnd.n3880 gnd.t277 1.27512
R21365 gnd.n3992 gnd.n2091 1.27512
R21366 gnd.n2069 gnd.t330 1.27512
R21367 gnd.n5553 gnd.n5552 1.16414
R21368 gnd.n6399 gnd.n5169 1.16414
R21369 gnd.n6323 gnd.n6316 1.16414
R21370 gnd.n6291 gnd.n6284 1.16414
R21371 gnd.n6259 gnd.n6252 1.16414
R21372 gnd.n6228 gnd.n6221 1.16414
R21373 gnd.n6196 gnd.n6189 1.16414
R21374 gnd.n6164 gnd.n6157 1.16414
R21375 gnd.n6132 gnd.n6125 1.16414
R21376 gnd.n6101 gnd.n6094 1.16414
R21377 gnd.n4467 gnd.n4466 0.970197
R21378 gnd.n4783 gnd.n1425 0.970197
R21379 gnd.n6307 gnd.n6275 0.962709
R21380 gnd.n6339 gnd.n6307 0.962709
R21381 gnd.n6180 gnd.n6148 0.962709
R21382 gnd.n6212 gnd.n6180 0.962709
R21383 gnd.t15 gnd.n5867 0.956468
R21384 gnd.n5211 gnd.t22 0.956468
R21385 gnd.t84 gnd.n1227 0.956468
R21386 gnd.n3031 gnd.t124 0.956468
R21387 gnd.n3298 gnd.t67 0.956468
R21388 gnd.n4070 gnd.t229 0.956468
R21389 gnd.n4249 gnd.t88 0.956468
R21390 gnd.n371 gnd.t129 0.956468
R21391 gnd.n2 gnd.n1 0.672012
R21392 gnd.n3 gnd.n2 0.672012
R21393 gnd.n4 gnd.n3 0.672012
R21394 gnd.n5 gnd.n4 0.672012
R21395 gnd.n6 gnd.n5 0.672012
R21396 gnd.n7 gnd.n6 0.672012
R21397 gnd.n9 gnd.n8 0.672012
R21398 gnd.n10 gnd.n9 0.672012
R21399 gnd.n11 gnd.n10 0.672012
R21400 gnd.n12 gnd.n11 0.672012
R21401 gnd.n13 gnd.n12 0.672012
R21402 gnd.n14 gnd.n13 0.672012
R21403 gnd.n3442 gnd.n1527 0.637812
R21404 gnd.n4673 gnd.n1537 0.637812
R21405 gnd.n3613 gnd.n3612 0.637812
R21406 gnd.n3656 gnd.n3654 0.637812
R21407 gnd.n3801 gnd.n3800 0.637812
R21408 gnd.n3819 gnd.n2138 0.637812
R21409 gnd gnd.n0 0.59317
R21410 gnd.n5322 gnd.n5321 0.573776
R21411 gnd.n5321 gnd.n5319 0.573776
R21412 gnd.n5319 gnd.n5317 0.573776
R21413 gnd.n5317 gnd.n5315 0.573776
R21414 gnd.n5315 gnd.n5313 0.573776
R21415 gnd.n5313 gnd.n5311 0.573776
R21416 gnd.n5311 gnd.n5309 0.573776
R21417 gnd.n5275 gnd.n5274 0.573776
R21418 gnd.n5274 gnd.n5272 0.573776
R21419 gnd.n5272 gnd.n5270 0.573776
R21420 gnd.n5270 gnd.n5268 0.573776
R21421 gnd.n5268 gnd.n5266 0.573776
R21422 gnd.n5266 gnd.n5264 0.573776
R21423 gnd.n5264 gnd.n5262 0.573776
R21424 gnd.n5290 gnd.n5289 0.573776
R21425 gnd.n5289 gnd.n5287 0.573776
R21426 gnd.n5287 gnd.n5285 0.573776
R21427 gnd.n5285 gnd.n5283 0.573776
R21428 gnd.n5283 gnd.n5281 0.573776
R21429 gnd.n5281 gnd.n5279 0.573776
R21430 gnd.n5279 gnd.n5277 0.573776
R21431 gnd.n5306 gnd.n5305 0.573776
R21432 gnd.n5305 gnd.n5303 0.573776
R21433 gnd.n5303 gnd.n5301 0.573776
R21434 gnd.n5301 gnd.n5299 0.573776
R21435 gnd.n5299 gnd.n5297 0.573776
R21436 gnd.n5297 gnd.n5295 0.573776
R21437 gnd.n5295 gnd.n5293 0.573776
R21438 gnd.n66 gnd.n64 0.573776
R21439 gnd.n68 gnd.n66 0.573776
R21440 gnd.n70 gnd.n68 0.573776
R21441 gnd.n72 gnd.n70 0.573776
R21442 gnd.n74 gnd.n72 0.573776
R21443 gnd.n76 gnd.n74 0.573776
R21444 gnd.n77 gnd.n76 0.573776
R21445 gnd.n19 gnd.n17 0.573776
R21446 gnd.n21 gnd.n19 0.573776
R21447 gnd.n23 gnd.n21 0.573776
R21448 gnd.n25 gnd.n23 0.573776
R21449 gnd.n27 gnd.n25 0.573776
R21450 gnd.n29 gnd.n27 0.573776
R21451 gnd.n30 gnd.n29 0.573776
R21452 gnd.n34 gnd.n32 0.573776
R21453 gnd.n36 gnd.n34 0.573776
R21454 gnd.n38 gnd.n36 0.573776
R21455 gnd.n40 gnd.n38 0.573776
R21456 gnd.n42 gnd.n40 0.573776
R21457 gnd.n44 gnd.n42 0.573776
R21458 gnd.n45 gnd.n44 0.573776
R21459 gnd.n50 gnd.n48 0.573776
R21460 gnd.n52 gnd.n50 0.573776
R21461 gnd.n54 gnd.n52 0.573776
R21462 gnd.n56 gnd.n54 0.573776
R21463 gnd.n58 gnd.n56 0.573776
R21464 gnd.n60 gnd.n58 0.573776
R21465 gnd.n61 gnd.n60 0.573776
R21466 gnd.n7684 gnd.n7683 0.553533
R21467 gnd.n7457 gnd.n7456 0.505073
R21468 gnd.n2806 gnd.n2805 0.505073
R21469 gnd.n4117 gnd.n1972 0.489829
R21470 gnd.n3155 gnd.n2407 0.489829
R21471 gnd.n3226 gnd.n3225 0.489829
R21472 gnd.n4585 gnd.n4584 0.489829
R21473 gnd.n6389 gnd.n6388 0.486781
R21474 gnd.n5605 gnd.n5501 0.48678
R21475 gnd.n6470 gnd.n6469 0.480683
R21476 gnd.n5673 gnd.n5451 0.480683
R21477 gnd.n7600 gnd.n7599 0.470012
R21478 gnd.n1804 gnd.n1722 0.470012
R21479 gnd.n4831 gnd.n4830 0.470012
R21480 gnd.n1146 gnd.n1072 0.470012
R21481 gnd.n803 gnd.n798 0.425805
R21482 gnd.n7133 gnd.n7132 0.425805
R21483 gnd.n7346 gnd.n7345 0.425805
R21484 gnd.n2724 gnd.n2721 0.425805
R21485 gnd.n7672 gnd.n95 0.4255
R21486 gnd.n4903 gnd.n1254 0.4255
R21487 gnd.n3167 gnd.n2617 0.388379
R21488 gnd.n6320 gnd.n6319 0.388379
R21489 gnd.n6288 gnd.n6287 0.388379
R21490 gnd.n6256 gnd.n6255 0.388379
R21491 gnd.n6225 gnd.n6224 0.388379
R21492 gnd.n6193 gnd.n6192 0.388379
R21493 gnd.n6161 gnd.n6160 0.388379
R21494 gnd.n6129 gnd.n6128 0.388379
R21495 gnd.n6098 gnd.n6097 0.388379
R21496 gnd.n4529 gnd.n1670 0.388379
R21497 gnd.n7684 gnd.n15 0.374463
R21498 gnd.n6366 gnd.t34 0.319156
R21499 gnd.n2703 gnd.t148 0.319156
R21500 gnd.n2661 gnd.t150 0.319156
R21501 gnd.n2411 gnd.t307 0.319156
R21502 gnd.t43 gnd.t7 0.319156
R21503 gnd.t60 gnd.t6 0.319156
R21504 gnd.t291 gnd.n2009 0.319156
R21505 gnd.n4272 gnd.t118 0.319156
R21506 gnd.t113 gnd.n85 0.319156
R21507 gnd.n5599 gnd.n5598 0.311721
R21508 gnd gnd.n7684 0.295112
R21509 gnd.n7490 gnd.n7489 0.293183
R21510 gnd.n4973 gnd.n1136 0.293183
R21511 gnd.n3148 gnd.n3147 0.27489
R21512 gnd.n4185 gnd.n4184 0.27489
R21513 gnd.n6439 gnd.n6438 0.268793
R21514 gnd.n7491 gnd.n7490 0.258122
R21515 gnd.n4405 gnd.n1623 0.258122
R21516 gnd.n2554 gnd.n2553 0.258122
R21517 gnd.n4974 gnd.n4973 0.258122
R21518 gnd.n6438 gnd.n6437 0.241354
R21519 gnd.n1752 gnd.n1749 0.229039
R21520 gnd.n1753 gnd.n1752 0.229039
R21521 gnd.n1428 gnd.n1424 0.229039
R21522 gnd.n2474 gnd.n1428 0.229039
R21523 gnd.n5728 gnd.n5469 0.206293
R21524 gnd.n5324 gnd.n0 0.169152
R21525 gnd.n6337 gnd.n6309 0.155672
R21526 gnd.n6330 gnd.n6309 0.155672
R21527 gnd.n6330 gnd.n6329 0.155672
R21528 gnd.n6329 gnd.n6313 0.155672
R21529 gnd.n6322 gnd.n6313 0.155672
R21530 gnd.n6322 gnd.n6321 0.155672
R21531 gnd.n6305 gnd.n6277 0.155672
R21532 gnd.n6298 gnd.n6277 0.155672
R21533 gnd.n6298 gnd.n6297 0.155672
R21534 gnd.n6297 gnd.n6281 0.155672
R21535 gnd.n6290 gnd.n6281 0.155672
R21536 gnd.n6290 gnd.n6289 0.155672
R21537 gnd.n6273 gnd.n6245 0.155672
R21538 gnd.n6266 gnd.n6245 0.155672
R21539 gnd.n6266 gnd.n6265 0.155672
R21540 gnd.n6265 gnd.n6249 0.155672
R21541 gnd.n6258 gnd.n6249 0.155672
R21542 gnd.n6258 gnd.n6257 0.155672
R21543 gnd.n6242 gnd.n6214 0.155672
R21544 gnd.n6235 gnd.n6214 0.155672
R21545 gnd.n6235 gnd.n6234 0.155672
R21546 gnd.n6234 gnd.n6218 0.155672
R21547 gnd.n6227 gnd.n6218 0.155672
R21548 gnd.n6227 gnd.n6226 0.155672
R21549 gnd.n6210 gnd.n6182 0.155672
R21550 gnd.n6203 gnd.n6182 0.155672
R21551 gnd.n6203 gnd.n6202 0.155672
R21552 gnd.n6202 gnd.n6186 0.155672
R21553 gnd.n6195 gnd.n6186 0.155672
R21554 gnd.n6195 gnd.n6194 0.155672
R21555 gnd.n6178 gnd.n6150 0.155672
R21556 gnd.n6171 gnd.n6150 0.155672
R21557 gnd.n6171 gnd.n6170 0.155672
R21558 gnd.n6170 gnd.n6154 0.155672
R21559 gnd.n6163 gnd.n6154 0.155672
R21560 gnd.n6163 gnd.n6162 0.155672
R21561 gnd.n6146 gnd.n6118 0.155672
R21562 gnd.n6139 gnd.n6118 0.155672
R21563 gnd.n6139 gnd.n6138 0.155672
R21564 gnd.n6138 gnd.n6122 0.155672
R21565 gnd.n6131 gnd.n6122 0.155672
R21566 gnd.n6131 gnd.n6130 0.155672
R21567 gnd.n6115 gnd.n6087 0.155672
R21568 gnd.n6108 gnd.n6087 0.155672
R21569 gnd.n6108 gnd.n6107 0.155672
R21570 gnd.n6107 gnd.n6091 0.155672
R21571 gnd.n6100 gnd.n6091 0.155672
R21572 gnd.n6100 gnd.n6099 0.155672
R21573 gnd.n6469 gnd.n5099 0.152939
R21574 gnd.n5101 gnd.n5099 0.152939
R21575 gnd.n5105 gnd.n5101 0.152939
R21576 gnd.n5106 gnd.n5105 0.152939
R21577 gnd.n5107 gnd.n5106 0.152939
R21578 gnd.n5108 gnd.n5107 0.152939
R21579 gnd.n5112 gnd.n5108 0.152939
R21580 gnd.n5113 gnd.n5112 0.152939
R21581 gnd.n5114 gnd.n5113 0.152939
R21582 gnd.n5115 gnd.n5114 0.152939
R21583 gnd.n5119 gnd.n5115 0.152939
R21584 gnd.n5120 gnd.n5119 0.152939
R21585 gnd.n5121 gnd.n5120 0.152939
R21586 gnd.n5122 gnd.n5121 0.152939
R21587 gnd.n5127 gnd.n5122 0.152939
R21588 gnd.n6439 gnd.n5127 0.152939
R21589 gnd.n5747 gnd.n5451 0.152939
R21590 gnd.n5748 gnd.n5747 0.152939
R21591 gnd.n5749 gnd.n5748 0.152939
R21592 gnd.n5749 gnd.n5430 0.152939
R21593 gnd.n5777 gnd.n5430 0.152939
R21594 gnd.n5778 gnd.n5777 0.152939
R21595 gnd.n5779 gnd.n5778 0.152939
R21596 gnd.n5780 gnd.n5779 0.152939
R21597 gnd.n5780 gnd.n5404 0.152939
R21598 gnd.n5811 gnd.n5404 0.152939
R21599 gnd.n5812 gnd.n5811 0.152939
R21600 gnd.n5813 gnd.n5812 0.152939
R21601 gnd.n5814 gnd.n5813 0.152939
R21602 gnd.n5815 gnd.n5814 0.152939
R21603 gnd.n5815 gnd.n5371 0.152939
R21604 gnd.n5872 gnd.n5371 0.152939
R21605 gnd.n5873 gnd.n5872 0.152939
R21606 gnd.n5874 gnd.n5873 0.152939
R21607 gnd.n5875 gnd.n5874 0.152939
R21608 gnd.n5875 gnd.n5344 0.152939
R21609 gnd.n5912 gnd.n5344 0.152939
R21610 gnd.n5913 gnd.n5912 0.152939
R21611 gnd.n5914 gnd.n5913 0.152939
R21612 gnd.n5915 gnd.n5914 0.152939
R21613 gnd.n5915 gnd.n5253 0.152939
R21614 gnd.n5957 gnd.n5253 0.152939
R21615 gnd.n5958 gnd.n5957 0.152939
R21616 gnd.n5959 gnd.n5958 0.152939
R21617 gnd.n5960 gnd.n5959 0.152939
R21618 gnd.n5960 gnd.n5225 0.152939
R21619 gnd.n5996 gnd.n5225 0.152939
R21620 gnd.n5997 gnd.n5996 0.152939
R21621 gnd.n5998 gnd.n5997 0.152939
R21622 gnd.n5999 gnd.n5998 0.152939
R21623 gnd.n6000 gnd.n5999 0.152939
R21624 gnd.n6000 gnd.n5195 0.152939
R21625 gnd.n6053 gnd.n5195 0.152939
R21626 gnd.n6054 gnd.n6053 0.152939
R21627 gnd.n6055 gnd.n6054 0.152939
R21628 gnd.n6056 gnd.n6055 0.152939
R21629 gnd.n6058 gnd.n6056 0.152939
R21630 gnd.n6058 gnd.n6057 0.152939
R21631 gnd.n6057 gnd.n985 0.152939
R21632 gnd.n986 gnd.n985 0.152939
R21633 gnd.n987 gnd.n986 0.152939
R21634 gnd.n1009 gnd.n987 0.152939
R21635 gnd.n1010 gnd.n1009 0.152939
R21636 gnd.n1011 gnd.n1010 0.152939
R21637 gnd.n1012 gnd.n1011 0.152939
R21638 gnd.n1013 gnd.n1012 0.152939
R21639 gnd.n5097 gnd.n1013 0.152939
R21640 gnd.n5098 gnd.n5097 0.152939
R21641 gnd.n6470 gnd.n5098 0.152939
R21642 gnd.n5674 gnd.n5673 0.152939
R21643 gnd.n5675 gnd.n5674 0.152939
R21644 gnd.n5676 gnd.n5675 0.152939
R21645 gnd.n5677 gnd.n5676 0.152939
R21646 gnd.n5678 gnd.n5677 0.152939
R21647 gnd.n5679 gnd.n5678 0.152939
R21648 gnd.n5680 gnd.n5679 0.152939
R21649 gnd.n5681 gnd.n5680 0.152939
R21650 gnd.n5682 gnd.n5681 0.152939
R21651 gnd.n5683 gnd.n5682 0.152939
R21652 gnd.n5684 gnd.n5683 0.152939
R21653 gnd.n5685 gnd.n5684 0.152939
R21654 gnd.n5686 gnd.n5685 0.152939
R21655 gnd.n5687 gnd.n5686 0.152939
R21656 gnd.n5691 gnd.n5687 0.152939
R21657 gnd.n5691 gnd.n5469 0.152939
R21658 gnd.n6437 gnd.n5129 0.152939
R21659 gnd.n5131 gnd.n5129 0.152939
R21660 gnd.n5135 gnd.n5131 0.152939
R21661 gnd.n5136 gnd.n5135 0.152939
R21662 gnd.n5137 gnd.n5136 0.152939
R21663 gnd.n5138 gnd.n5137 0.152939
R21664 gnd.n5142 gnd.n5138 0.152939
R21665 gnd.n5143 gnd.n5142 0.152939
R21666 gnd.n5144 gnd.n5143 0.152939
R21667 gnd.n5145 gnd.n5144 0.152939
R21668 gnd.n5149 gnd.n5145 0.152939
R21669 gnd.n5150 gnd.n5149 0.152939
R21670 gnd.n5151 gnd.n5150 0.152939
R21671 gnd.n5152 gnd.n5151 0.152939
R21672 gnd.n5156 gnd.n5152 0.152939
R21673 gnd.n5157 gnd.n5156 0.152939
R21674 gnd.n5158 gnd.n5157 0.152939
R21675 gnd.n5159 gnd.n5158 0.152939
R21676 gnd.n5163 gnd.n5159 0.152939
R21677 gnd.n5164 gnd.n5163 0.152939
R21678 gnd.n5165 gnd.n5164 0.152939
R21679 gnd.n5166 gnd.n5165 0.152939
R21680 gnd.n5173 gnd.n5166 0.152939
R21681 gnd.n5174 gnd.n5173 0.152939
R21682 gnd.n5175 gnd.n5174 0.152939
R21683 gnd.n6389 gnd.n5175 0.152939
R21684 gnd.n5934 gnd.n5933 0.152939
R21685 gnd.n5935 gnd.n5934 0.152939
R21686 gnd.n5936 gnd.n5935 0.152939
R21687 gnd.n5937 gnd.n5936 0.152939
R21688 gnd.n5938 gnd.n5937 0.152939
R21689 gnd.n5939 gnd.n5938 0.152939
R21690 gnd.n5940 gnd.n5939 0.152939
R21691 gnd.n5941 gnd.n5940 0.152939
R21692 gnd.n5941 gnd.n5207 0.152939
R21693 gnd.n6019 gnd.n5207 0.152939
R21694 gnd.n6020 gnd.n6019 0.152939
R21695 gnd.n6021 gnd.n6020 0.152939
R21696 gnd.n6022 gnd.n6021 0.152939
R21697 gnd.n6023 gnd.n6022 0.152939
R21698 gnd.n6024 gnd.n6023 0.152939
R21699 gnd.n6025 gnd.n6024 0.152939
R21700 gnd.n6026 gnd.n6025 0.152939
R21701 gnd.n6027 gnd.n6026 0.152939
R21702 gnd.n6027 gnd.n5180 0.152939
R21703 gnd.n6370 gnd.n5180 0.152939
R21704 gnd.n6371 gnd.n6370 0.152939
R21705 gnd.n6372 gnd.n6371 0.152939
R21706 gnd.n6372 gnd.n5178 0.152939
R21707 gnd.n6380 gnd.n5178 0.152939
R21708 gnd.n6381 gnd.n6380 0.152939
R21709 gnd.n6382 gnd.n6381 0.152939
R21710 gnd.n6382 gnd.n5176 0.152939
R21711 gnd.n6388 gnd.n5176 0.152939
R21712 gnd.n5606 gnd.n5605 0.152939
R21713 gnd.n5607 gnd.n5606 0.152939
R21714 gnd.n5607 gnd.n5489 0.152939
R21715 gnd.n5621 gnd.n5489 0.152939
R21716 gnd.n5622 gnd.n5621 0.152939
R21717 gnd.n5623 gnd.n5622 0.152939
R21718 gnd.n5623 gnd.n5476 0.152939
R21719 gnd.n5637 gnd.n5476 0.152939
R21720 gnd.n5638 gnd.n5637 0.152939
R21721 gnd.n5639 gnd.n5638 0.152939
R21722 gnd.n5640 gnd.n5639 0.152939
R21723 gnd.n5641 gnd.n5640 0.152939
R21724 gnd.n5642 gnd.n5641 0.152939
R21725 gnd.n5643 gnd.n5642 0.152939
R21726 gnd.n5644 gnd.n5643 0.152939
R21727 gnd.n5645 gnd.n5644 0.152939
R21728 gnd.n5646 gnd.n5645 0.152939
R21729 gnd.n5647 gnd.n5646 0.152939
R21730 gnd.n5648 gnd.n5647 0.152939
R21731 gnd.n5648 gnd.n5411 0.152939
R21732 gnd.n5800 gnd.n5411 0.152939
R21733 gnd.n5801 gnd.n5800 0.152939
R21734 gnd.n5802 gnd.n5801 0.152939
R21735 gnd.n5803 gnd.n5802 0.152939
R21736 gnd.n5803 gnd.n5378 0.152939
R21737 gnd.n5847 gnd.n5378 0.152939
R21738 gnd.n5848 gnd.n5847 0.152939
R21739 gnd.n5849 gnd.n5848 0.152939
R21740 gnd.n5598 gnd.n5505 0.152939
R21741 gnd.n5508 gnd.n5505 0.152939
R21742 gnd.n5509 gnd.n5508 0.152939
R21743 gnd.n5510 gnd.n5509 0.152939
R21744 gnd.n5513 gnd.n5510 0.152939
R21745 gnd.n5514 gnd.n5513 0.152939
R21746 gnd.n5515 gnd.n5514 0.152939
R21747 gnd.n5516 gnd.n5515 0.152939
R21748 gnd.n5519 gnd.n5516 0.152939
R21749 gnd.n5520 gnd.n5519 0.152939
R21750 gnd.n5521 gnd.n5520 0.152939
R21751 gnd.n5522 gnd.n5521 0.152939
R21752 gnd.n5525 gnd.n5522 0.152939
R21753 gnd.n5526 gnd.n5525 0.152939
R21754 gnd.n5527 gnd.n5526 0.152939
R21755 gnd.n5528 gnd.n5527 0.152939
R21756 gnd.n5531 gnd.n5528 0.152939
R21757 gnd.n5532 gnd.n5531 0.152939
R21758 gnd.n5533 gnd.n5532 0.152939
R21759 gnd.n5534 gnd.n5533 0.152939
R21760 gnd.n5537 gnd.n5534 0.152939
R21761 gnd.n5538 gnd.n5537 0.152939
R21762 gnd.n5541 gnd.n5538 0.152939
R21763 gnd.n5542 gnd.n5541 0.152939
R21764 gnd.n5544 gnd.n5542 0.152939
R21765 gnd.n5544 gnd.n5501 0.152939
R21766 gnd.n6682 gnd.n798 0.152939
R21767 gnd.n6683 gnd.n6682 0.152939
R21768 gnd.n6684 gnd.n6683 0.152939
R21769 gnd.n6684 gnd.n792 0.152939
R21770 gnd.n6692 gnd.n792 0.152939
R21771 gnd.n6693 gnd.n6692 0.152939
R21772 gnd.n6694 gnd.n6693 0.152939
R21773 gnd.n6694 gnd.n786 0.152939
R21774 gnd.n6702 gnd.n786 0.152939
R21775 gnd.n6703 gnd.n6702 0.152939
R21776 gnd.n6704 gnd.n6703 0.152939
R21777 gnd.n6704 gnd.n780 0.152939
R21778 gnd.n6712 gnd.n780 0.152939
R21779 gnd.n6713 gnd.n6712 0.152939
R21780 gnd.n6714 gnd.n6713 0.152939
R21781 gnd.n6714 gnd.n774 0.152939
R21782 gnd.n6722 gnd.n774 0.152939
R21783 gnd.n6723 gnd.n6722 0.152939
R21784 gnd.n6724 gnd.n6723 0.152939
R21785 gnd.n6724 gnd.n768 0.152939
R21786 gnd.n6732 gnd.n768 0.152939
R21787 gnd.n6733 gnd.n6732 0.152939
R21788 gnd.n6734 gnd.n6733 0.152939
R21789 gnd.n6734 gnd.n762 0.152939
R21790 gnd.n6742 gnd.n762 0.152939
R21791 gnd.n6743 gnd.n6742 0.152939
R21792 gnd.n6744 gnd.n6743 0.152939
R21793 gnd.n6744 gnd.n756 0.152939
R21794 gnd.n6752 gnd.n756 0.152939
R21795 gnd.n6753 gnd.n6752 0.152939
R21796 gnd.n6754 gnd.n6753 0.152939
R21797 gnd.n6754 gnd.n750 0.152939
R21798 gnd.n6762 gnd.n750 0.152939
R21799 gnd.n6763 gnd.n6762 0.152939
R21800 gnd.n6764 gnd.n6763 0.152939
R21801 gnd.n6764 gnd.n744 0.152939
R21802 gnd.n6772 gnd.n744 0.152939
R21803 gnd.n6773 gnd.n6772 0.152939
R21804 gnd.n6774 gnd.n6773 0.152939
R21805 gnd.n6774 gnd.n738 0.152939
R21806 gnd.n6782 gnd.n738 0.152939
R21807 gnd.n6783 gnd.n6782 0.152939
R21808 gnd.n6784 gnd.n6783 0.152939
R21809 gnd.n6784 gnd.n732 0.152939
R21810 gnd.n6792 gnd.n732 0.152939
R21811 gnd.n6793 gnd.n6792 0.152939
R21812 gnd.n6794 gnd.n6793 0.152939
R21813 gnd.n6794 gnd.n726 0.152939
R21814 gnd.n6802 gnd.n726 0.152939
R21815 gnd.n6803 gnd.n6802 0.152939
R21816 gnd.n6804 gnd.n6803 0.152939
R21817 gnd.n6804 gnd.n720 0.152939
R21818 gnd.n6812 gnd.n720 0.152939
R21819 gnd.n6813 gnd.n6812 0.152939
R21820 gnd.n6814 gnd.n6813 0.152939
R21821 gnd.n6814 gnd.n714 0.152939
R21822 gnd.n6822 gnd.n714 0.152939
R21823 gnd.n6823 gnd.n6822 0.152939
R21824 gnd.n6824 gnd.n6823 0.152939
R21825 gnd.n6824 gnd.n708 0.152939
R21826 gnd.n6832 gnd.n708 0.152939
R21827 gnd.n6833 gnd.n6832 0.152939
R21828 gnd.n6834 gnd.n6833 0.152939
R21829 gnd.n6834 gnd.n702 0.152939
R21830 gnd.n6842 gnd.n702 0.152939
R21831 gnd.n6843 gnd.n6842 0.152939
R21832 gnd.n6844 gnd.n6843 0.152939
R21833 gnd.n6844 gnd.n696 0.152939
R21834 gnd.n6852 gnd.n696 0.152939
R21835 gnd.n6853 gnd.n6852 0.152939
R21836 gnd.n6854 gnd.n6853 0.152939
R21837 gnd.n6854 gnd.n690 0.152939
R21838 gnd.n6862 gnd.n690 0.152939
R21839 gnd.n6863 gnd.n6862 0.152939
R21840 gnd.n6864 gnd.n6863 0.152939
R21841 gnd.n6864 gnd.n684 0.152939
R21842 gnd.n6872 gnd.n684 0.152939
R21843 gnd.n6873 gnd.n6872 0.152939
R21844 gnd.n6874 gnd.n6873 0.152939
R21845 gnd.n6874 gnd.n678 0.152939
R21846 gnd.n6882 gnd.n678 0.152939
R21847 gnd.n6883 gnd.n6882 0.152939
R21848 gnd.n6884 gnd.n6883 0.152939
R21849 gnd.n6884 gnd.n672 0.152939
R21850 gnd.n6892 gnd.n672 0.152939
R21851 gnd.n6893 gnd.n6892 0.152939
R21852 gnd.n6894 gnd.n6893 0.152939
R21853 gnd.n6894 gnd.n666 0.152939
R21854 gnd.n6902 gnd.n666 0.152939
R21855 gnd.n6903 gnd.n6902 0.152939
R21856 gnd.n6904 gnd.n6903 0.152939
R21857 gnd.n6904 gnd.n660 0.152939
R21858 gnd.n6912 gnd.n660 0.152939
R21859 gnd.n6913 gnd.n6912 0.152939
R21860 gnd.n6914 gnd.n6913 0.152939
R21861 gnd.n6914 gnd.n654 0.152939
R21862 gnd.n6922 gnd.n654 0.152939
R21863 gnd.n6923 gnd.n6922 0.152939
R21864 gnd.n6924 gnd.n6923 0.152939
R21865 gnd.n6924 gnd.n648 0.152939
R21866 gnd.n6932 gnd.n648 0.152939
R21867 gnd.n6933 gnd.n6932 0.152939
R21868 gnd.n6934 gnd.n6933 0.152939
R21869 gnd.n6934 gnd.n642 0.152939
R21870 gnd.n6942 gnd.n642 0.152939
R21871 gnd.n6943 gnd.n6942 0.152939
R21872 gnd.n6944 gnd.n6943 0.152939
R21873 gnd.n6944 gnd.n636 0.152939
R21874 gnd.n6952 gnd.n636 0.152939
R21875 gnd.n6953 gnd.n6952 0.152939
R21876 gnd.n6954 gnd.n6953 0.152939
R21877 gnd.n6954 gnd.n630 0.152939
R21878 gnd.n6962 gnd.n630 0.152939
R21879 gnd.n6963 gnd.n6962 0.152939
R21880 gnd.n6964 gnd.n6963 0.152939
R21881 gnd.n6964 gnd.n624 0.152939
R21882 gnd.n6972 gnd.n624 0.152939
R21883 gnd.n6973 gnd.n6972 0.152939
R21884 gnd.n6974 gnd.n6973 0.152939
R21885 gnd.n6974 gnd.n618 0.152939
R21886 gnd.n6982 gnd.n618 0.152939
R21887 gnd.n6983 gnd.n6982 0.152939
R21888 gnd.n6984 gnd.n6983 0.152939
R21889 gnd.n6984 gnd.n612 0.152939
R21890 gnd.n6992 gnd.n612 0.152939
R21891 gnd.n6993 gnd.n6992 0.152939
R21892 gnd.n6994 gnd.n6993 0.152939
R21893 gnd.n6994 gnd.n606 0.152939
R21894 gnd.n7002 gnd.n606 0.152939
R21895 gnd.n7003 gnd.n7002 0.152939
R21896 gnd.n7004 gnd.n7003 0.152939
R21897 gnd.n7004 gnd.n600 0.152939
R21898 gnd.n7012 gnd.n600 0.152939
R21899 gnd.n7013 gnd.n7012 0.152939
R21900 gnd.n7014 gnd.n7013 0.152939
R21901 gnd.n7014 gnd.n594 0.152939
R21902 gnd.n7022 gnd.n594 0.152939
R21903 gnd.n7023 gnd.n7022 0.152939
R21904 gnd.n7024 gnd.n7023 0.152939
R21905 gnd.n7024 gnd.n588 0.152939
R21906 gnd.n7032 gnd.n588 0.152939
R21907 gnd.n7033 gnd.n7032 0.152939
R21908 gnd.n7034 gnd.n7033 0.152939
R21909 gnd.n7034 gnd.n582 0.152939
R21910 gnd.n7042 gnd.n582 0.152939
R21911 gnd.n7043 gnd.n7042 0.152939
R21912 gnd.n7044 gnd.n7043 0.152939
R21913 gnd.n7044 gnd.n576 0.152939
R21914 gnd.n7052 gnd.n576 0.152939
R21915 gnd.n7053 gnd.n7052 0.152939
R21916 gnd.n7054 gnd.n7053 0.152939
R21917 gnd.n7054 gnd.n570 0.152939
R21918 gnd.n7062 gnd.n570 0.152939
R21919 gnd.n7063 gnd.n7062 0.152939
R21920 gnd.n7064 gnd.n7063 0.152939
R21921 gnd.n7064 gnd.n564 0.152939
R21922 gnd.n7072 gnd.n564 0.152939
R21923 gnd.n7073 gnd.n7072 0.152939
R21924 gnd.n7074 gnd.n7073 0.152939
R21925 gnd.n7074 gnd.n558 0.152939
R21926 gnd.n7082 gnd.n558 0.152939
R21927 gnd.n7083 gnd.n7082 0.152939
R21928 gnd.n7084 gnd.n7083 0.152939
R21929 gnd.n7084 gnd.n552 0.152939
R21930 gnd.n7092 gnd.n552 0.152939
R21931 gnd.n7093 gnd.n7092 0.152939
R21932 gnd.n7094 gnd.n7093 0.152939
R21933 gnd.n7094 gnd.n546 0.152939
R21934 gnd.n7102 gnd.n546 0.152939
R21935 gnd.n7103 gnd.n7102 0.152939
R21936 gnd.n7104 gnd.n7103 0.152939
R21937 gnd.n7104 gnd.n540 0.152939
R21938 gnd.n7112 gnd.n540 0.152939
R21939 gnd.n7113 gnd.n7112 0.152939
R21940 gnd.n7114 gnd.n7113 0.152939
R21941 gnd.n7114 gnd.n534 0.152939
R21942 gnd.n7122 gnd.n534 0.152939
R21943 gnd.n7123 gnd.n7122 0.152939
R21944 gnd.n7124 gnd.n7123 0.152939
R21945 gnd.n7124 gnd.n528 0.152939
R21946 gnd.n7132 gnd.n528 0.152939
R21947 gnd.n7134 gnd.n7133 0.152939
R21948 gnd.n7134 gnd.n522 0.152939
R21949 gnd.n7142 gnd.n522 0.152939
R21950 gnd.n7143 gnd.n7142 0.152939
R21951 gnd.n7144 gnd.n7143 0.152939
R21952 gnd.n7144 gnd.n516 0.152939
R21953 gnd.n7152 gnd.n516 0.152939
R21954 gnd.n7153 gnd.n7152 0.152939
R21955 gnd.n7154 gnd.n7153 0.152939
R21956 gnd.n7154 gnd.n510 0.152939
R21957 gnd.n7162 gnd.n510 0.152939
R21958 gnd.n7163 gnd.n7162 0.152939
R21959 gnd.n7164 gnd.n7163 0.152939
R21960 gnd.n7164 gnd.n504 0.152939
R21961 gnd.n7172 gnd.n504 0.152939
R21962 gnd.n7173 gnd.n7172 0.152939
R21963 gnd.n7174 gnd.n7173 0.152939
R21964 gnd.n7174 gnd.n498 0.152939
R21965 gnd.n7182 gnd.n498 0.152939
R21966 gnd.n7183 gnd.n7182 0.152939
R21967 gnd.n7184 gnd.n7183 0.152939
R21968 gnd.n7184 gnd.n492 0.152939
R21969 gnd.n7192 gnd.n492 0.152939
R21970 gnd.n7193 gnd.n7192 0.152939
R21971 gnd.n7194 gnd.n7193 0.152939
R21972 gnd.n7194 gnd.n486 0.152939
R21973 gnd.n7202 gnd.n486 0.152939
R21974 gnd.n7203 gnd.n7202 0.152939
R21975 gnd.n7204 gnd.n7203 0.152939
R21976 gnd.n7204 gnd.n480 0.152939
R21977 gnd.n7212 gnd.n480 0.152939
R21978 gnd.n7213 gnd.n7212 0.152939
R21979 gnd.n7214 gnd.n7213 0.152939
R21980 gnd.n7214 gnd.n474 0.152939
R21981 gnd.n7222 gnd.n474 0.152939
R21982 gnd.n7223 gnd.n7222 0.152939
R21983 gnd.n7224 gnd.n7223 0.152939
R21984 gnd.n7224 gnd.n468 0.152939
R21985 gnd.n7232 gnd.n468 0.152939
R21986 gnd.n7233 gnd.n7232 0.152939
R21987 gnd.n7234 gnd.n7233 0.152939
R21988 gnd.n7234 gnd.n462 0.152939
R21989 gnd.n7242 gnd.n462 0.152939
R21990 gnd.n7243 gnd.n7242 0.152939
R21991 gnd.n7244 gnd.n7243 0.152939
R21992 gnd.n7244 gnd.n456 0.152939
R21993 gnd.n7252 gnd.n456 0.152939
R21994 gnd.n7253 gnd.n7252 0.152939
R21995 gnd.n7254 gnd.n7253 0.152939
R21996 gnd.n7254 gnd.n450 0.152939
R21997 gnd.n7262 gnd.n450 0.152939
R21998 gnd.n7263 gnd.n7262 0.152939
R21999 gnd.n7264 gnd.n7263 0.152939
R22000 gnd.n7264 gnd.n444 0.152939
R22001 gnd.n7272 gnd.n444 0.152939
R22002 gnd.n7273 gnd.n7272 0.152939
R22003 gnd.n7274 gnd.n7273 0.152939
R22004 gnd.n7274 gnd.n438 0.152939
R22005 gnd.n7282 gnd.n438 0.152939
R22006 gnd.n7283 gnd.n7282 0.152939
R22007 gnd.n7284 gnd.n7283 0.152939
R22008 gnd.n7284 gnd.n432 0.152939
R22009 gnd.n7292 gnd.n432 0.152939
R22010 gnd.n7293 gnd.n7292 0.152939
R22011 gnd.n7294 gnd.n7293 0.152939
R22012 gnd.n7294 gnd.n426 0.152939
R22013 gnd.n7302 gnd.n426 0.152939
R22014 gnd.n7303 gnd.n7302 0.152939
R22015 gnd.n7304 gnd.n7303 0.152939
R22016 gnd.n7304 gnd.n420 0.152939
R22017 gnd.n7312 gnd.n420 0.152939
R22018 gnd.n7313 gnd.n7312 0.152939
R22019 gnd.n7314 gnd.n7313 0.152939
R22020 gnd.n7314 gnd.n414 0.152939
R22021 gnd.n7322 gnd.n414 0.152939
R22022 gnd.n7323 gnd.n7322 0.152939
R22023 gnd.n7324 gnd.n7323 0.152939
R22024 gnd.n7324 gnd.n408 0.152939
R22025 gnd.n7332 gnd.n408 0.152939
R22026 gnd.n7333 gnd.n7332 0.152939
R22027 gnd.n7334 gnd.n7333 0.152939
R22028 gnd.n7335 gnd.n7334 0.152939
R22029 gnd.n7335 gnd.n402 0.152939
R22030 gnd.n7345 gnd.n402 0.152939
R22031 gnd.n388 gnd.n385 0.152939
R22032 gnd.n389 gnd.n388 0.152939
R22033 gnd.n390 gnd.n389 0.152939
R22034 gnd.n391 gnd.n390 0.152939
R22035 gnd.n394 gnd.n391 0.152939
R22036 gnd.n395 gnd.n394 0.152939
R22037 gnd.n396 gnd.n395 0.152939
R22038 gnd.n397 gnd.n396 0.152939
R22039 gnd.n400 gnd.n397 0.152939
R22040 gnd.n401 gnd.n400 0.152939
R22041 gnd.n7346 gnd.n401 0.152939
R22042 gnd.n118 gnd.n93 0.152939
R22043 gnd.n119 gnd.n118 0.152939
R22044 gnd.n120 gnd.n119 0.152939
R22045 gnd.n137 gnd.n120 0.152939
R22046 gnd.n138 gnd.n137 0.152939
R22047 gnd.n139 gnd.n138 0.152939
R22048 gnd.n140 gnd.n139 0.152939
R22049 gnd.n157 gnd.n140 0.152939
R22050 gnd.n158 gnd.n157 0.152939
R22051 gnd.n159 gnd.n158 0.152939
R22052 gnd.n160 gnd.n159 0.152939
R22053 gnd.n177 gnd.n160 0.152939
R22054 gnd.n178 gnd.n177 0.152939
R22055 gnd.n179 gnd.n178 0.152939
R22056 gnd.n180 gnd.n179 0.152939
R22057 gnd.n196 gnd.n180 0.152939
R22058 gnd.n197 gnd.n196 0.152939
R22059 gnd.n198 gnd.n197 0.152939
R22060 gnd.n199 gnd.n198 0.152939
R22061 gnd.n214 gnd.n199 0.152939
R22062 gnd.n7600 gnd.n214 0.152939
R22063 gnd.n7681 gnd.n80 0.152939
R22064 gnd.n7370 gnd.n80 0.152939
R22065 gnd.n7371 gnd.n7370 0.152939
R22066 gnd.n7371 gnd.n376 0.152939
R22067 gnd.n7383 gnd.n376 0.152939
R22068 gnd.n7384 gnd.n7383 0.152939
R22069 gnd.n7385 gnd.n7384 0.152939
R22070 gnd.n7385 gnd.n369 0.152939
R22071 gnd.n7397 gnd.n369 0.152939
R22072 gnd.n7398 gnd.n7397 0.152939
R22073 gnd.n7399 gnd.n7398 0.152939
R22074 gnd.n7399 gnd.n364 0.152939
R22075 gnd.n7411 gnd.n364 0.152939
R22076 gnd.n7412 gnd.n7411 0.152939
R22077 gnd.n7414 gnd.n7412 0.152939
R22078 gnd.n7414 gnd.n7413 0.152939
R22079 gnd.n7413 gnd.n358 0.152939
R22080 gnd.n7442 gnd.n358 0.152939
R22081 gnd.n7443 gnd.n7442 0.152939
R22082 gnd.n7444 gnd.n7443 0.152939
R22083 gnd.n7444 gnd.n355 0.152939
R22084 gnd.n7449 gnd.n355 0.152939
R22085 gnd.n7450 gnd.n7449 0.152939
R22086 gnd.n7451 gnd.n7450 0.152939
R22087 gnd.n7451 gnd.n352 0.152939
R22088 gnd.n7456 gnd.n352 0.152939
R22089 gnd.n7489 gnd.n318 0.152939
R22090 gnd.n320 gnd.n318 0.152939
R22091 gnd.n324 gnd.n320 0.152939
R22092 gnd.n325 gnd.n324 0.152939
R22093 gnd.n326 gnd.n325 0.152939
R22094 gnd.n327 gnd.n326 0.152939
R22095 gnd.n331 gnd.n327 0.152939
R22096 gnd.n332 gnd.n331 0.152939
R22097 gnd.n333 gnd.n332 0.152939
R22098 gnd.n334 gnd.n333 0.152939
R22099 gnd.n338 gnd.n334 0.152939
R22100 gnd.n339 gnd.n338 0.152939
R22101 gnd.n340 gnd.n339 0.152939
R22102 gnd.n341 gnd.n340 0.152939
R22103 gnd.n345 gnd.n341 0.152939
R22104 gnd.n346 gnd.n345 0.152939
R22105 gnd.n7458 gnd.n346 0.152939
R22106 gnd.n7458 gnd.n7457 0.152939
R22107 gnd.n7599 gnd.n215 0.152939
R22108 gnd.n217 gnd.n215 0.152939
R22109 gnd.n221 gnd.n217 0.152939
R22110 gnd.n222 gnd.n221 0.152939
R22111 gnd.n223 gnd.n222 0.152939
R22112 gnd.n224 gnd.n223 0.152939
R22113 gnd.n228 gnd.n224 0.152939
R22114 gnd.n229 gnd.n228 0.152939
R22115 gnd.n230 gnd.n229 0.152939
R22116 gnd.n231 gnd.n230 0.152939
R22117 gnd.n235 gnd.n231 0.152939
R22118 gnd.n236 gnd.n235 0.152939
R22119 gnd.n237 gnd.n236 0.152939
R22120 gnd.n238 gnd.n237 0.152939
R22121 gnd.n242 gnd.n238 0.152939
R22122 gnd.n243 gnd.n242 0.152939
R22123 gnd.n244 gnd.n243 0.152939
R22124 gnd.n245 gnd.n244 0.152939
R22125 gnd.n249 gnd.n245 0.152939
R22126 gnd.n250 gnd.n249 0.152939
R22127 gnd.n251 gnd.n250 0.152939
R22128 gnd.n252 gnd.n251 0.152939
R22129 gnd.n256 gnd.n252 0.152939
R22130 gnd.n257 gnd.n256 0.152939
R22131 gnd.n258 gnd.n257 0.152939
R22132 gnd.n259 gnd.n258 0.152939
R22133 gnd.n263 gnd.n259 0.152939
R22134 gnd.n264 gnd.n263 0.152939
R22135 gnd.n265 gnd.n264 0.152939
R22136 gnd.n266 gnd.n265 0.152939
R22137 gnd.n270 gnd.n266 0.152939
R22138 gnd.n271 gnd.n270 0.152939
R22139 gnd.n272 gnd.n271 0.152939
R22140 gnd.n273 gnd.n272 0.152939
R22141 gnd.n277 gnd.n273 0.152939
R22142 gnd.n278 gnd.n277 0.152939
R22143 gnd.n7530 gnd.n278 0.152939
R22144 gnd.n7530 gnd.n7529 0.152939
R22145 gnd.n7529 gnd.n7528 0.152939
R22146 gnd.n7528 gnd.n282 0.152939
R22147 gnd.n288 gnd.n282 0.152939
R22148 gnd.n289 gnd.n288 0.152939
R22149 gnd.n290 gnd.n289 0.152939
R22150 gnd.n291 gnd.n290 0.152939
R22151 gnd.n295 gnd.n291 0.152939
R22152 gnd.n296 gnd.n295 0.152939
R22153 gnd.n297 gnd.n296 0.152939
R22154 gnd.n298 gnd.n297 0.152939
R22155 gnd.n302 gnd.n298 0.152939
R22156 gnd.n303 gnd.n302 0.152939
R22157 gnd.n304 gnd.n303 0.152939
R22158 gnd.n305 gnd.n304 0.152939
R22159 gnd.n309 gnd.n305 0.152939
R22160 gnd.n310 gnd.n309 0.152939
R22161 gnd.n311 gnd.n310 0.152939
R22162 gnd.n312 gnd.n311 0.152939
R22163 gnd.n317 gnd.n312 0.152939
R22164 gnd.n7491 gnd.n317 0.152939
R22165 gnd.n1723 gnd.n1722 0.152939
R22166 gnd.n1724 gnd.n1723 0.152939
R22167 gnd.n1725 gnd.n1724 0.152939
R22168 gnd.n1726 gnd.n1725 0.152939
R22169 gnd.n1727 gnd.n1726 0.152939
R22170 gnd.n1728 gnd.n1727 0.152939
R22171 gnd.n1729 gnd.n1728 0.152939
R22172 gnd.n1730 gnd.n1729 0.152939
R22173 gnd.n1731 gnd.n1730 0.152939
R22174 gnd.n1732 gnd.n1731 0.152939
R22175 gnd.n1733 gnd.n1732 0.152939
R22176 gnd.n1734 gnd.n1733 0.152939
R22177 gnd.n1735 gnd.n1734 0.152939
R22178 gnd.n1736 gnd.n1735 0.152939
R22179 gnd.n1737 gnd.n1736 0.152939
R22180 gnd.n1738 gnd.n1737 0.152939
R22181 gnd.n1739 gnd.n1738 0.152939
R22182 gnd.n1742 gnd.n1739 0.152939
R22183 gnd.n1743 gnd.n1742 0.152939
R22184 gnd.n1744 gnd.n1743 0.152939
R22185 gnd.n1745 gnd.n1744 0.152939
R22186 gnd.n1746 gnd.n1745 0.152939
R22187 gnd.n1747 gnd.n1746 0.152939
R22188 gnd.n1748 gnd.n1747 0.152939
R22189 gnd.n1749 gnd.n1748 0.152939
R22190 gnd.n1754 gnd.n1753 0.152939
R22191 gnd.n1755 gnd.n1754 0.152939
R22192 gnd.n1756 gnd.n1755 0.152939
R22193 gnd.n1757 gnd.n1756 0.152939
R22194 gnd.n1758 gnd.n1757 0.152939
R22195 gnd.n1759 gnd.n1758 0.152939
R22196 gnd.n1760 gnd.n1759 0.152939
R22197 gnd.n1761 gnd.n1760 0.152939
R22198 gnd.n1762 gnd.n1761 0.152939
R22199 gnd.n1765 gnd.n1762 0.152939
R22200 gnd.n1766 gnd.n1765 0.152939
R22201 gnd.n1767 gnd.n1766 0.152939
R22202 gnd.n1768 gnd.n1767 0.152939
R22203 gnd.n1769 gnd.n1768 0.152939
R22204 gnd.n1770 gnd.n1769 0.152939
R22205 gnd.n1771 gnd.n1770 0.152939
R22206 gnd.n1772 gnd.n1771 0.152939
R22207 gnd.n1773 gnd.n1772 0.152939
R22208 gnd.n1774 gnd.n1773 0.152939
R22209 gnd.n1775 gnd.n1774 0.152939
R22210 gnd.n1776 gnd.n1775 0.152939
R22211 gnd.n1777 gnd.n1776 0.152939
R22212 gnd.n1778 gnd.n1777 0.152939
R22213 gnd.n1779 gnd.n1778 0.152939
R22214 gnd.n1780 gnd.n1779 0.152939
R22215 gnd.n1781 gnd.n1780 0.152939
R22216 gnd.n1782 gnd.n1781 0.152939
R22217 gnd.n1783 gnd.n1782 0.152939
R22218 gnd.n4406 gnd.n1783 0.152939
R22219 gnd.n4406 gnd.n4405 0.152939
R22220 gnd.n1805 gnd.n1804 0.152939
R22221 gnd.n1806 gnd.n1805 0.152939
R22222 gnd.n1807 gnd.n1806 0.152939
R22223 gnd.n1808 gnd.n1807 0.152939
R22224 gnd.n1828 gnd.n1808 0.152939
R22225 gnd.n1829 gnd.n1828 0.152939
R22226 gnd.n1830 gnd.n1829 0.152939
R22227 gnd.n1831 gnd.n1830 0.152939
R22228 gnd.n1849 gnd.n1831 0.152939
R22229 gnd.n1850 gnd.n1849 0.152939
R22230 gnd.n1851 gnd.n1850 0.152939
R22231 gnd.n1852 gnd.n1851 0.152939
R22232 gnd.n1868 gnd.n1852 0.152939
R22233 gnd.n1869 gnd.n1868 0.152939
R22234 gnd.n1870 gnd.n1869 0.152939
R22235 gnd.n1871 gnd.n1870 0.152939
R22236 gnd.n1889 gnd.n1871 0.152939
R22237 gnd.n1890 gnd.n1889 0.152939
R22238 gnd.n1891 gnd.n1890 0.152939
R22239 gnd.n1892 gnd.n1891 0.152939
R22240 gnd.n1892 gnd.n94 0.152939
R22241 gnd.n2976 gnd.n2973 0.152939
R22242 gnd.n2977 gnd.n2976 0.152939
R22243 gnd.n2978 gnd.n2977 0.152939
R22244 gnd.n2979 gnd.n2978 0.152939
R22245 gnd.n2981 gnd.n2979 0.152939
R22246 gnd.n2981 gnd.n2980 0.152939
R22247 gnd.n2980 gnd.n2644 0.152939
R22248 gnd.n3061 gnd.n2644 0.152939
R22249 gnd.n3062 gnd.n3061 0.152939
R22250 gnd.n3063 gnd.n3062 0.152939
R22251 gnd.n3063 gnd.n2640 0.152939
R22252 gnd.n3069 gnd.n2640 0.152939
R22253 gnd.n3070 gnd.n3069 0.152939
R22254 gnd.n3071 gnd.n3070 0.152939
R22255 gnd.n3072 gnd.n3071 0.152939
R22256 gnd.n3073 gnd.n3072 0.152939
R22257 gnd.n3076 gnd.n3073 0.152939
R22258 gnd.n3077 gnd.n3076 0.152939
R22259 gnd.n3078 gnd.n3077 0.152939
R22260 gnd.n3079 gnd.n3078 0.152939
R22261 gnd.n3082 gnd.n3079 0.152939
R22262 gnd.n3083 gnd.n3082 0.152939
R22263 gnd.n3084 gnd.n3083 0.152939
R22264 gnd.n3085 gnd.n3084 0.152939
R22265 gnd.n3090 gnd.n3085 0.152939
R22266 gnd.n3091 gnd.n3090 0.152939
R22267 gnd.n3092 gnd.n3091 0.152939
R22268 gnd.n3093 gnd.n3092 0.152939
R22269 gnd.n3093 gnd.n2400 0.152939
R22270 gnd.n3244 gnd.n2400 0.152939
R22271 gnd.n3245 gnd.n3244 0.152939
R22272 gnd.n3246 gnd.n3245 0.152939
R22273 gnd.n3247 gnd.n3246 0.152939
R22274 gnd.n3247 gnd.n2375 0.152939
R22275 gnd.n3274 gnd.n2375 0.152939
R22276 gnd.n3275 gnd.n3274 0.152939
R22277 gnd.n3276 gnd.n3275 0.152939
R22278 gnd.n3277 gnd.n3276 0.152939
R22279 gnd.n3278 gnd.n3277 0.152939
R22280 gnd.n3280 gnd.n3278 0.152939
R22281 gnd.n3280 gnd.n3279 0.152939
R22282 gnd.n3279 gnd.n1496 0.152939
R22283 gnd.n1497 gnd.n1496 0.152939
R22284 gnd.n1498 gnd.n1497 0.152939
R22285 gnd.n1511 gnd.n1498 0.152939
R22286 gnd.n1512 gnd.n1511 0.152939
R22287 gnd.n1513 gnd.n1512 0.152939
R22288 gnd.n1514 gnd.n1513 0.152939
R22289 gnd.n1529 gnd.n1514 0.152939
R22290 gnd.n1530 gnd.n1529 0.152939
R22291 gnd.n1531 gnd.n1530 0.152939
R22292 gnd.n1532 gnd.n1531 0.152939
R22293 gnd.n3482 gnd.n1532 0.152939
R22294 gnd.n3485 gnd.n3482 0.152939
R22295 gnd.n3486 gnd.n3485 0.152939
R22296 gnd.n3487 gnd.n3486 0.152939
R22297 gnd.n3488 gnd.n3487 0.152939
R22298 gnd.n3489 gnd.n3488 0.152939
R22299 gnd.n3490 gnd.n3489 0.152939
R22300 gnd.n3490 gnd.n2275 0.152939
R22301 gnd.n3567 gnd.n2275 0.152939
R22302 gnd.n3568 gnd.n3567 0.152939
R22303 gnd.n3569 gnd.n3568 0.152939
R22304 gnd.n3569 gnd.n2251 0.152939
R22305 gnd.n3606 gnd.n2251 0.152939
R22306 gnd.n3607 gnd.n3606 0.152939
R22307 gnd.n3608 gnd.n3607 0.152939
R22308 gnd.n3608 gnd.n2229 0.152939
R22309 gnd.n3660 gnd.n2229 0.152939
R22310 gnd.n3661 gnd.n3660 0.152939
R22311 gnd.n3662 gnd.n3661 0.152939
R22312 gnd.n3662 gnd.n2210 0.152939
R22313 gnd.n3686 gnd.n2210 0.152939
R22314 gnd.n3687 gnd.n3686 0.152939
R22315 gnd.n3688 gnd.n3687 0.152939
R22316 gnd.n3688 gnd.n2187 0.152939
R22317 gnd.n3752 gnd.n2187 0.152939
R22318 gnd.n3753 gnd.n3752 0.152939
R22319 gnd.n3754 gnd.n3753 0.152939
R22320 gnd.n3754 gnd.n2165 0.152939
R22321 gnd.n3782 gnd.n2165 0.152939
R22322 gnd.n3783 gnd.n3782 0.152939
R22323 gnd.n3784 gnd.n3783 0.152939
R22324 gnd.n3784 gnd.n2143 0.152939
R22325 gnd.n3813 gnd.n2143 0.152939
R22326 gnd.n3814 gnd.n3813 0.152939
R22327 gnd.n3815 gnd.n3814 0.152939
R22328 gnd.n3815 gnd.n2117 0.152939
R22329 gnd.n3862 gnd.n2117 0.152939
R22330 gnd.n3863 gnd.n3862 0.152939
R22331 gnd.n3864 gnd.n3863 0.152939
R22332 gnd.n3864 gnd.n2101 0.152939
R22333 gnd.n3893 gnd.n2101 0.152939
R22334 gnd.n3894 gnd.n3893 0.152939
R22335 gnd.n3895 gnd.n3894 0.152939
R22336 gnd.n3895 gnd.n2047 0.152939
R22337 gnd.n4064 gnd.n2047 0.152939
R22338 gnd.n4065 gnd.n4064 0.152939
R22339 gnd.n4066 gnd.n4065 0.152939
R22340 gnd.n4066 gnd.n2034 0.152939
R22341 gnd.n4084 gnd.n2034 0.152939
R22342 gnd.n4085 gnd.n4084 0.152939
R22343 gnd.n4086 gnd.n4085 0.152939
R22344 gnd.n4086 gnd.n2021 0.152939
R22345 gnd.n4104 gnd.n2021 0.152939
R22346 gnd.n4105 gnd.n4104 0.152939
R22347 gnd.n4106 gnd.n4105 0.152939
R22348 gnd.n4107 gnd.n4106 0.152939
R22349 gnd.n4107 gnd.n2006 0.152939
R22350 gnd.n4128 gnd.n2006 0.152939
R22351 gnd.n4129 gnd.n4128 0.152939
R22352 gnd.n4130 gnd.n4129 0.152939
R22353 gnd.n4131 gnd.n4130 0.152939
R22354 gnd.n4132 gnd.n4131 0.152939
R22355 gnd.n4135 gnd.n4132 0.152939
R22356 gnd.n4136 gnd.n4135 0.152939
R22357 gnd.n4137 gnd.n4136 0.152939
R22358 gnd.n4138 gnd.n4137 0.152939
R22359 gnd.n4141 gnd.n4138 0.152939
R22360 gnd.n4142 gnd.n4141 0.152939
R22361 gnd.n4143 gnd.n4142 0.152939
R22362 gnd.n4144 gnd.n4143 0.152939
R22363 gnd.n4147 gnd.n4144 0.152939
R22364 gnd.n4148 gnd.n4147 0.152939
R22365 gnd.n4149 gnd.n4148 0.152939
R22366 gnd.n4150 gnd.n4149 0.152939
R22367 gnd.n4152 gnd.n4150 0.152939
R22368 gnd.n4152 gnd.n4151 0.152939
R22369 gnd.n4151 gnd.n1949 0.152939
R22370 gnd.n4254 gnd.n1949 0.152939
R22371 gnd.n4255 gnd.n4254 0.152939
R22372 gnd.n4256 gnd.n4255 0.152939
R22373 gnd.n4256 gnd.n1945 0.152939
R22374 gnd.n4262 gnd.n1945 0.152939
R22375 gnd.n4263 gnd.n4262 0.152939
R22376 gnd.n4264 gnd.n4263 0.152939
R22377 gnd.n4265 gnd.n4264 0.152939
R22378 gnd.n2806 gnd.n2747 0.152939
R22379 gnd.n2812 gnd.n2747 0.152939
R22380 gnd.n2813 gnd.n2812 0.152939
R22381 gnd.n2814 gnd.n2813 0.152939
R22382 gnd.n2814 gnd.n2745 0.152939
R22383 gnd.n2820 gnd.n2745 0.152939
R22384 gnd.n2821 gnd.n2820 0.152939
R22385 gnd.n2822 gnd.n2821 0.152939
R22386 gnd.n2822 gnd.n2743 0.152939
R22387 gnd.n2845 gnd.n2743 0.152939
R22388 gnd.n2846 gnd.n2845 0.152939
R22389 gnd.n2848 gnd.n2846 0.152939
R22390 gnd.n2848 gnd.n2847 0.152939
R22391 gnd.n2847 gnd.n2737 0.152939
R22392 gnd.n2738 gnd.n2737 0.152939
R22393 gnd.n2739 gnd.n2738 0.152939
R22394 gnd.n2860 gnd.n2739 0.152939
R22395 gnd.n2861 gnd.n2860 0.152939
R22396 gnd.n2862 gnd.n2861 0.152939
R22397 gnd.n2863 gnd.n2862 0.152939
R22398 gnd.n2864 gnd.n2863 0.152939
R22399 gnd.n2865 gnd.n2864 0.152939
R22400 gnd.n2865 gnd.n2694 0.152939
R22401 gnd.n2937 gnd.n2694 0.152939
R22402 gnd.n2938 gnd.n2937 0.152939
R22403 gnd.n2939 gnd.n2938 0.152939
R22404 gnd.n2761 gnd.n1136 0.152939
R22405 gnd.n2769 gnd.n2761 0.152939
R22406 gnd.n2770 gnd.n2769 0.152939
R22407 gnd.n2771 gnd.n2770 0.152939
R22408 gnd.n2771 gnd.n2759 0.152939
R22409 gnd.n2779 gnd.n2759 0.152939
R22410 gnd.n2780 gnd.n2779 0.152939
R22411 gnd.n2781 gnd.n2780 0.152939
R22412 gnd.n2781 gnd.n2757 0.152939
R22413 gnd.n2789 gnd.n2757 0.152939
R22414 gnd.n2790 gnd.n2789 0.152939
R22415 gnd.n2791 gnd.n2790 0.152939
R22416 gnd.n2791 gnd.n2755 0.152939
R22417 gnd.n2799 gnd.n2755 0.152939
R22418 gnd.n2800 gnd.n2799 0.152939
R22419 gnd.n2801 gnd.n2800 0.152939
R22420 gnd.n2801 gnd.n2748 0.152939
R22421 gnd.n2805 gnd.n2748 0.152939
R22422 gnd.n1278 gnd.n1253 0.152939
R22423 gnd.n1279 gnd.n1278 0.152939
R22424 gnd.n1280 gnd.n1279 0.152939
R22425 gnd.n1298 gnd.n1280 0.152939
R22426 gnd.n1299 gnd.n1298 0.152939
R22427 gnd.n1300 gnd.n1299 0.152939
R22428 gnd.n1301 gnd.n1300 0.152939
R22429 gnd.n1317 gnd.n1301 0.152939
R22430 gnd.n1318 gnd.n1317 0.152939
R22431 gnd.n1319 gnd.n1318 0.152939
R22432 gnd.n1320 gnd.n1319 0.152939
R22433 gnd.n1338 gnd.n1320 0.152939
R22434 gnd.n1339 gnd.n1338 0.152939
R22435 gnd.n1340 gnd.n1339 0.152939
R22436 gnd.n1341 gnd.n1340 0.152939
R22437 gnd.n1358 gnd.n1341 0.152939
R22438 gnd.n1359 gnd.n1358 0.152939
R22439 gnd.n1360 gnd.n1359 0.152939
R22440 gnd.n1361 gnd.n1360 0.152939
R22441 gnd.n1378 gnd.n1361 0.152939
R22442 gnd.n4831 gnd.n1378 0.152939
R22443 gnd.n4830 gnd.n1379 0.152939
R22444 gnd.n1384 gnd.n1379 0.152939
R22445 gnd.n1385 gnd.n1384 0.152939
R22446 gnd.n1386 gnd.n1385 0.152939
R22447 gnd.n1387 gnd.n1386 0.152939
R22448 gnd.n1388 gnd.n1387 0.152939
R22449 gnd.n1392 gnd.n1388 0.152939
R22450 gnd.n1393 gnd.n1392 0.152939
R22451 gnd.n1394 gnd.n1393 0.152939
R22452 gnd.n1395 gnd.n1394 0.152939
R22453 gnd.n1399 gnd.n1395 0.152939
R22454 gnd.n1400 gnd.n1399 0.152939
R22455 gnd.n1401 gnd.n1400 0.152939
R22456 gnd.n1402 gnd.n1401 0.152939
R22457 gnd.n1406 gnd.n1402 0.152939
R22458 gnd.n1407 gnd.n1406 0.152939
R22459 gnd.n1408 gnd.n1407 0.152939
R22460 gnd.n1411 gnd.n1408 0.152939
R22461 gnd.n1415 gnd.n1411 0.152939
R22462 gnd.n1416 gnd.n1415 0.152939
R22463 gnd.n1417 gnd.n1416 0.152939
R22464 gnd.n1418 gnd.n1417 0.152939
R22465 gnd.n1422 gnd.n1418 0.152939
R22466 gnd.n1423 gnd.n1422 0.152939
R22467 gnd.n1424 gnd.n1423 0.152939
R22468 gnd.n2475 gnd.n2474 0.152939
R22469 gnd.n2484 gnd.n2475 0.152939
R22470 gnd.n2485 gnd.n2484 0.152939
R22471 gnd.n2486 gnd.n2485 0.152939
R22472 gnd.n2486 gnd.n2470 0.152939
R22473 gnd.n2494 gnd.n2470 0.152939
R22474 gnd.n2495 gnd.n2494 0.152939
R22475 gnd.n2496 gnd.n2495 0.152939
R22476 gnd.n2496 gnd.n2464 0.152939
R22477 gnd.n2504 gnd.n2464 0.152939
R22478 gnd.n2505 gnd.n2504 0.152939
R22479 gnd.n2506 gnd.n2505 0.152939
R22480 gnd.n2506 gnd.n2460 0.152939
R22481 gnd.n2514 gnd.n2460 0.152939
R22482 gnd.n2515 gnd.n2514 0.152939
R22483 gnd.n2516 gnd.n2515 0.152939
R22484 gnd.n2516 gnd.n2456 0.152939
R22485 gnd.n2524 gnd.n2456 0.152939
R22486 gnd.n2525 gnd.n2524 0.152939
R22487 gnd.n2526 gnd.n2525 0.152939
R22488 gnd.n2526 gnd.n2452 0.152939
R22489 gnd.n2534 gnd.n2452 0.152939
R22490 gnd.n2535 gnd.n2534 0.152939
R22491 gnd.n2536 gnd.n2535 0.152939
R22492 gnd.n2536 gnd.n2448 0.152939
R22493 gnd.n2544 gnd.n2448 0.152939
R22494 gnd.n2545 gnd.n2544 0.152939
R22495 gnd.n2546 gnd.n2545 0.152939
R22496 gnd.n2546 gnd.n2442 0.152939
R22497 gnd.n2553 gnd.n2442 0.152939
R22498 gnd.n1073 gnd.n1072 0.152939
R22499 gnd.n1074 gnd.n1073 0.152939
R22500 gnd.n1075 gnd.n1074 0.152939
R22501 gnd.n1076 gnd.n1075 0.152939
R22502 gnd.n1077 gnd.n1076 0.152939
R22503 gnd.n1078 gnd.n1077 0.152939
R22504 gnd.n1079 gnd.n1078 0.152939
R22505 gnd.n1080 gnd.n1079 0.152939
R22506 gnd.n1081 gnd.n1080 0.152939
R22507 gnd.n1082 gnd.n1081 0.152939
R22508 gnd.n1083 gnd.n1082 0.152939
R22509 gnd.n1084 gnd.n1083 0.152939
R22510 gnd.n1085 gnd.n1084 0.152939
R22511 gnd.n1086 gnd.n1085 0.152939
R22512 gnd.n1087 gnd.n1086 0.152939
R22513 gnd.n1088 gnd.n1087 0.152939
R22514 gnd.n1089 gnd.n1088 0.152939
R22515 gnd.n1092 gnd.n1089 0.152939
R22516 gnd.n1093 gnd.n1092 0.152939
R22517 gnd.n1094 gnd.n1093 0.152939
R22518 gnd.n1095 gnd.n1094 0.152939
R22519 gnd.n1096 gnd.n1095 0.152939
R22520 gnd.n1097 gnd.n1096 0.152939
R22521 gnd.n1098 gnd.n1097 0.152939
R22522 gnd.n1099 gnd.n1098 0.152939
R22523 gnd.n1100 gnd.n1099 0.152939
R22524 gnd.n1101 gnd.n1100 0.152939
R22525 gnd.n1102 gnd.n1101 0.152939
R22526 gnd.n1103 gnd.n1102 0.152939
R22527 gnd.n1104 gnd.n1103 0.152939
R22528 gnd.n1105 gnd.n1104 0.152939
R22529 gnd.n1106 gnd.n1105 0.152939
R22530 gnd.n1107 gnd.n1106 0.152939
R22531 gnd.n1108 gnd.n1107 0.152939
R22532 gnd.n1109 gnd.n1108 0.152939
R22533 gnd.n1110 gnd.n1109 0.152939
R22534 gnd.n1111 gnd.n1110 0.152939
R22535 gnd.n1114 gnd.n1111 0.152939
R22536 gnd.n1115 gnd.n1114 0.152939
R22537 gnd.n1116 gnd.n1115 0.152939
R22538 gnd.n1117 gnd.n1116 0.152939
R22539 gnd.n1118 gnd.n1117 0.152939
R22540 gnd.n1119 gnd.n1118 0.152939
R22541 gnd.n1120 gnd.n1119 0.152939
R22542 gnd.n1121 gnd.n1120 0.152939
R22543 gnd.n1122 gnd.n1121 0.152939
R22544 gnd.n1123 gnd.n1122 0.152939
R22545 gnd.n1124 gnd.n1123 0.152939
R22546 gnd.n1125 gnd.n1124 0.152939
R22547 gnd.n1126 gnd.n1125 0.152939
R22548 gnd.n1127 gnd.n1126 0.152939
R22549 gnd.n1128 gnd.n1127 0.152939
R22550 gnd.n1129 gnd.n1128 0.152939
R22551 gnd.n1130 gnd.n1129 0.152939
R22552 gnd.n1131 gnd.n1130 0.152939
R22553 gnd.n1132 gnd.n1131 0.152939
R22554 gnd.n4975 gnd.n1132 0.152939
R22555 gnd.n4975 gnd.n4974 0.152939
R22556 gnd.n1147 gnd.n1146 0.152939
R22557 gnd.n1148 gnd.n1147 0.152939
R22558 gnd.n1149 gnd.n1148 0.152939
R22559 gnd.n1169 gnd.n1149 0.152939
R22560 gnd.n1170 gnd.n1169 0.152939
R22561 gnd.n1171 gnd.n1170 0.152939
R22562 gnd.n1172 gnd.n1171 0.152939
R22563 gnd.n1188 gnd.n1172 0.152939
R22564 gnd.n1189 gnd.n1188 0.152939
R22565 gnd.n1190 gnd.n1189 0.152939
R22566 gnd.n1191 gnd.n1190 0.152939
R22567 gnd.n1209 gnd.n1191 0.152939
R22568 gnd.n1210 gnd.n1209 0.152939
R22569 gnd.n1211 gnd.n1210 0.152939
R22570 gnd.n1212 gnd.n1211 0.152939
R22571 gnd.n1229 gnd.n1212 0.152939
R22572 gnd.n1230 gnd.n1229 0.152939
R22573 gnd.n1231 gnd.n1230 0.152939
R22574 gnd.n1232 gnd.n1231 0.152939
R22575 gnd.n1250 gnd.n1232 0.152939
R22576 gnd.n1251 gnd.n1250 0.152939
R22577 gnd.n2730 gnd.n2721 0.152939
R22578 gnd.n2731 gnd.n2730 0.152939
R22579 gnd.n2732 gnd.n2731 0.152939
R22580 gnd.n2732 gnd.n2717 0.152939
R22581 gnd.n2895 gnd.n2717 0.152939
R22582 gnd.n2896 gnd.n2895 0.152939
R22583 gnd.n2897 gnd.n2896 0.152939
R22584 gnd.n2897 gnd.n2713 0.152939
R22585 gnd.n2904 gnd.n2713 0.152939
R22586 gnd.n2905 gnd.n2904 0.152939
R22587 gnd.n2906 gnd.n2905 0.152939
R22588 gnd.n804 gnd.n803 0.152939
R22589 gnd.n805 gnd.n804 0.152939
R22590 gnd.n810 gnd.n805 0.152939
R22591 gnd.n811 gnd.n810 0.152939
R22592 gnd.n812 gnd.n811 0.152939
R22593 gnd.n813 gnd.n812 0.152939
R22594 gnd.n818 gnd.n813 0.152939
R22595 gnd.n819 gnd.n818 0.152939
R22596 gnd.n820 gnd.n819 0.152939
R22597 gnd.n821 gnd.n820 0.152939
R22598 gnd.n826 gnd.n821 0.152939
R22599 gnd.n827 gnd.n826 0.152939
R22600 gnd.n828 gnd.n827 0.152939
R22601 gnd.n829 gnd.n828 0.152939
R22602 gnd.n834 gnd.n829 0.152939
R22603 gnd.n835 gnd.n834 0.152939
R22604 gnd.n836 gnd.n835 0.152939
R22605 gnd.n837 gnd.n836 0.152939
R22606 gnd.n842 gnd.n837 0.152939
R22607 gnd.n843 gnd.n842 0.152939
R22608 gnd.n844 gnd.n843 0.152939
R22609 gnd.n845 gnd.n844 0.152939
R22610 gnd.n850 gnd.n845 0.152939
R22611 gnd.n851 gnd.n850 0.152939
R22612 gnd.n852 gnd.n851 0.152939
R22613 gnd.n853 gnd.n852 0.152939
R22614 gnd.n858 gnd.n853 0.152939
R22615 gnd.n859 gnd.n858 0.152939
R22616 gnd.n860 gnd.n859 0.152939
R22617 gnd.n861 gnd.n860 0.152939
R22618 gnd.n866 gnd.n861 0.152939
R22619 gnd.n867 gnd.n866 0.152939
R22620 gnd.n868 gnd.n867 0.152939
R22621 gnd.n869 gnd.n868 0.152939
R22622 gnd.n874 gnd.n869 0.152939
R22623 gnd.n875 gnd.n874 0.152939
R22624 gnd.n876 gnd.n875 0.152939
R22625 gnd.n877 gnd.n876 0.152939
R22626 gnd.n882 gnd.n877 0.152939
R22627 gnd.n883 gnd.n882 0.152939
R22628 gnd.n884 gnd.n883 0.152939
R22629 gnd.n885 gnd.n884 0.152939
R22630 gnd.n890 gnd.n885 0.152939
R22631 gnd.n891 gnd.n890 0.152939
R22632 gnd.n892 gnd.n891 0.152939
R22633 gnd.n893 gnd.n892 0.152939
R22634 gnd.n898 gnd.n893 0.152939
R22635 gnd.n899 gnd.n898 0.152939
R22636 gnd.n900 gnd.n899 0.152939
R22637 gnd.n901 gnd.n900 0.152939
R22638 gnd.n906 gnd.n901 0.152939
R22639 gnd.n907 gnd.n906 0.152939
R22640 gnd.n908 gnd.n907 0.152939
R22641 gnd.n909 gnd.n908 0.152939
R22642 gnd.n914 gnd.n909 0.152939
R22643 gnd.n915 gnd.n914 0.152939
R22644 gnd.n916 gnd.n915 0.152939
R22645 gnd.n917 gnd.n916 0.152939
R22646 gnd.n922 gnd.n917 0.152939
R22647 gnd.n923 gnd.n922 0.152939
R22648 gnd.n924 gnd.n923 0.152939
R22649 gnd.n925 gnd.n924 0.152939
R22650 gnd.n930 gnd.n925 0.152939
R22651 gnd.n931 gnd.n930 0.152939
R22652 gnd.n932 gnd.n931 0.152939
R22653 gnd.n933 gnd.n932 0.152939
R22654 gnd.n938 gnd.n933 0.152939
R22655 gnd.n939 gnd.n938 0.152939
R22656 gnd.n940 gnd.n939 0.152939
R22657 gnd.n941 gnd.n940 0.152939
R22658 gnd.n946 gnd.n941 0.152939
R22659 gnd.n947 gnd.n946 0.152939
R22660 gnd.n948 gnd.n947 0.152939
R22661 gnd.n949 gnd.n948 0.152939
R22662 gnd.n954 gnd.n949 0.152939
R22663 gnd.n955 gnd.n954 0.152939
R22664 gnd.n956 gnd.n955 0.152939
R22665 gnd.n957 gnd.n956 0.152939
R22666 gnd.n962 gnd.n957 0.152939
R22667 gnd.n963 gnd.n962 0.152939
R22668 gnd.n964 gnd.n963 0.152939
R22669 gnd.n965 gnd.n964 0.152939
R22670 gnd.n2723 gnd.n965 0.152939
R22671 gnd.n2724 gnd.n2723 0.152939
R22672 gnd.n3234 gnd.n2407 0.152939
R22673 gnd.n3235 gnd.n3234 0.152939
R22674 gnd.n3237 gnd.n3235 0.152939
R22675 gnd.n3237 gnd.n3236 0.152939
R22676 gnd.n3236 gnd.n2382 0.152939
R22677 gnd.n3264 gnd.n2382 0.152939
R22678 gnd.n3265 gnd.n3264 0.152939
R22679 gnd.n3267 gnd.n3265 0.152939
R22680 gnd.n3267 gnd.n3266 0.152939
R22681 gnd.n3266 gnd.n2358 0.152939
R22682 gnd.n3301 gnd.n2358 0.152939
R22683 gnd.n3302 gnd.n3301 0.152939
R22684 gnd.n3304 gnd.n3302 0.152939
R22685 gnd.n3304 gnd.n3303 0.152939
R22686 gnd.n3303 gnd.n2345 0.152939
R22687 gnd.n3428 gnd.n2345 0.152939
R22688 gnd.n3429 gnd.n3428 0.152939
R22689 gnd.n3432 gnd.n3429 0.152939
R22690 gnd.n3432 gnd.n3431 0.152939
R22691 gnd.n3431 gnd.n3430 0.152939
R22692 gnd.n3430 gnd.n2329 0.152939
R22693 gnd.n3456 gnd.n2329 0.152939
R22694 gnd.n3457 gnd.n3456 0.152939
R22695 gnd.n3459 gnd.n3457 0.152939
R22696 gnd.n3459 gnd.n3458 0.152939
R22697 gnd.n3458 gnd.n2310 0.152939
R22698 gnd.n3511 gnd.n2310 0.152939
R22699 gnd.n3512 gnd.n3511 0.152939
R22700 gnd.n3515 gnd.n3512 0.152939
R22701 gnd.n3515 gnd.n3514 0.152939
R22702 gnd.n3514 gnd.n3513 0.152939
R22703 gnd.n3513 gnd.n2294 0.152939
R22704 gnd.n3541 gnd.n2294 0.152939
R22705 gnd.n3542 gnd.n3541 0.152939
R22706 gnd.n3543 gnd.n3542 0.152939
R22707 gnd.n3543 gnd.n2268 0.152939
R22708 gnd.n3589 gnd.n2268 0.152939
R22709 gnd.n3589 gnd.n3588 0.152939
R22710 gnd.n3588 gnd.n3587 0.152939
R22711 gnd.n3587 gnd.n2244 0.152939
R22712 gnd.n3644 gnd.n2244 0.152939
R22713 gnd.n3644 gnd.n3643 0.152939
R22714 gnd.n3643 gnd.n3642 0.152939
R22715 gnd.n3642 gnd.n2245 0.152939
R22716 gnd.n3638 gnd.n2245 0.152939
R22717 gnd.n3638 gnd.n3637 0.152939
R22718 gnd.n3637 gnd.n3636 0.152939
R22719 gnd.n3636 gnd.n3629 0.152939
R22720 gnd.n3632 gnd.n3629 0.152939
R22721 gnd.n3632 gnd.n2180 0.152939
R22722 gnd.n3761 gnd.n2180 0.152939
R22723 gnd.n3762 gnd.n3761 0.152939
R22724 gnd.n3763 gnd.n3762 0.152939
R22725 gnd.n3763 gnd.n2159 0.152939
R22726 gnd.n3791 gnd.n2159 0.152939
R22727 gnd.n3792 gnd.n3791 0.152939
R22728 gnd.n3797 gnd.n3792 0.152939
R22729 gnd.n3797 gnd.n3796 0.152939
R22730 gnd.n3796 gnd.n3795 0.152939
R22731 gnd.n3795 gnd.n2130 0.152939
R22732 gnd.n3830 gnd.n2130 0.152939
R22733 gnd.n3831 gnd.n3830 0.152939
R22734 gnd.n3848 gnd.n3831 0.152939
R22735 gnd.n3848 gnd.n3847 0.152939
R22736 gnd.n3847 gnd.n3846 0.152939
R22737 gnd.n3846 gnd.n3832 0.152939
R22738 gnd.n3842 gnd.n3832 0.152939
R22739 gnd.n3842 gnd.n3841 0.152939
R22740 gnd.n3841 gnd.n3840 0.152939
R22741 gnd.n3840 gnd.n2040 0.152939
R22742 gnd.n4073 gnd.n2040 0.152939
R22743 gnd.n4074 gnd.n4073 0.152939
R22744 gnd.n4075 gnd.n4074 0.152939
R22745 gnd.n4075 gnd.n2027 0.152939
R22746 gnd.n4093 gnd.n2027 0.152939
R22747 gnd.n4094 gnd.n4093 0.152939
R22748 gnd.n4095 gnd.n4094 0.152939
R22749 gnd.n4095 gnd.n2013 0.152939
R22750 gnd.n4115 gnd.n2013 0.152939
R22751 gnd.n4116 gnd.n4115 0.152939
R22752 gnd.n4118 gnd.n4116 0.152939
R22753 gnd.n4118 gnd.n4117 0.152939
R22754 gnd.n2944 gnd.n2943 0.152939
R22755 gnd.n2943 gnd.n2664 0.152939
R22756 gnd.n2999 gnd.n2664 0.152939
R22757 gnd.n3000 gnd.n2999 0.152939
R22758 gnd.n3001 gnd.n3000 0.152939
R22759 gnd.n3001 gnd.n2659 0.152939
R22760 gnd.n3014 gnd.n2659 0.152939
R22761 gnd.n3015 gnd.n3014 0.152939
R22762 gnd.n3016 gnd.n3015 0.152939
R22763 gnd.n3016 gnd.n2651 0.152939
R22764 gnd.n3052 gnd.n2651 0.152939
R22765 gnd.n3052 gnd.n3051 0.152939
R22766 gnd.n3051 gnd.n3050 0.152939
R22767 gnd.n3050 gnd.n2652 0.152939
R22768 gnd.n3046 gnd.n2652 0.152939
R22769 gnd.n3046 gnd.n3045 0.152939
R22770 gnd.n3045 gnd.n3044 0.152939
R22771 gnd.n3044 gnd.n2656 0.152939
R22772 gnd.n3040 gnd.n2656 0.152939
R22773 gnd.n3040 gnd.n2632 0.152939
R22774 gnd.n3130 gnd.n2632 0.152939
R22775 gnd.n3131 gnd.n3130 0.152939
R22776 gnd.n3133 gnd.n3131 0.152939
R22777 gnd.n3133 gnd.n3132 0.152939
R22778 gnd.n3132 gnd.n2627 0.152939
R22779 gnd.n3147 gnd.n2627 0.152939
R22780 gnd.n3225 gnd.n2416 0.152939
R22781 gnd.n3218 gnd.n2416 0.152939
R22782 gnd.n3218 gnd.n3217 0.152939
R22783 gnd.n3217 gnd.n3216 0.152939
R22784 gnd.n3216 gnd.n2436 0.152939
R22785 gnd.n3212 gnd.n2436 0.152939
R22786 gnd.n3228 gnd.n3226 0.152939
R22787 gnd.n3228 gnd.n3227 0.152939
R22788 gnd.n3227 gnd.n2391 0.152939
R22789 gnd.n3255 gnd.n2391 0.152939
R22790 gnd.n3256 gnd.n3255 0.152939
R22791 gnd.n3258 gnd.n3256 0.152939
R22792 gnd.n3258 gnd.n3257 0.152939
R22793 gnd.n3257 gnd.n2365 0.152939
R22794 gnd.n3292 gnd.n2365 0.152939
R22795 gnd.n3293 gnd.n3292 0.152939
R22796 gnd.n3295 gnd.n3293 0.152939
R22797 gnd.n3295 gnd.n3294 0.152939
R22798 gnd.n3294 gnd.n2351 0.152939
R22799 gnd.n3420 gnd.n2351 0.152939
R22800 gnd.n3421 gnd.n3420 0.152939
R22801 gnd.n3422 gnd.n3421 0.152939
R22802 gnd.n3422 gnd.n2337 0.152939
R22803 gnd.n3438 gnd.n2337 0.152939
R22804 gnd.n3439 gnd.n3438 0.152939
R22805 gnd.n3448 gnd.n3439 0.152939
R22806 gnd.n3448 gnd.n3447 0.152939
R22807 gnd.n3447 gnd.n3446 0.152939
R22808 gnd.n3446 gnd.n3440 0.152939
R22809 gnd.n3440 gnd.n1542 0.152939
R22810 gnd.n4670 gnd.n1542 0.152939
R22811 gnd.n4670 gnd.n4669 0.152939
R22812 gnd.n4669 gnd.n4668 0.152939
R22813 gnd.n4668 gnd.n1543 0.152939
R22814 gnd.n4664 gnd.n1543 0.152939
R22815 gnd.n4664 gnd.n4663 0.152939
R22816 gnd.n4663 gnd.n4662 0.152939
R22817 gnd.n4662 gnd.n1548 0.152939
R22818 gnd.n4658 gnd.n1548 0.152939
R22819 gnd.n4658 gnd.n4657 0.152939
R22820 gnd.n4657 gnd.n4656 0.152939
R22821 gnd.n4656 gnd.n1553 0.152939
R22822 gnd.n4652 gnd.n1553 0.152939
R22823 gnd.n4652 gnd.n4651 0.152939
R22824 gnd.n4651 gnd.n4650 0.152939
R22825 gnd.n4650 gnd.n1558 0.152939
R22826 gnd.n4646 gnd.n1558 0.152939
R22827 gnd.n4646 gnd.n4645 0.152939
R22828 gnd.n4645 gnd.n4644 0.152939
R22829 gnd.n4644 gnd.n1563 0.152939
R22830 gnd.n4640 gnd.n1563 0.152939
R22831 gnd.n4640 gnd.n4639 0.152939
R22832 gnd.n4639 gnd.n4638 0.152939
R22833 gnd.n4638 gnd.n1568 0.152939
R22834 gnd.n4634 gnd.n1568 0.152939
R22835 gnd.n4634 gnd.n4633 0.152939
R22836 gnd.n4633 gnd.n4632 0.152939
R22837 gnd.n4632 gnd.n1573 0.152939
R22838 gnd.n4628 gnd.n1573 0.152939
R22839 gnd.n4628 gnd.n4627 0.152939
R22840 gnd.n4627 gnd.n4626 0.152939
R22841 gnd.n4626 gnd.n1578 0.152939
R22842 gnd.n4622 gnd.n1578 0.152939
R22843 gnd.n4622 gnd.n4621 0.152939
R22844 gnd.n4621 gnd.n4620 0.152939
R22845 gnd.n4620 gnd.n1583 0.152939
R22846 gnd.n4616 gnd.n1583 0.152939
R22847 gnd.n4616 gnd.n4615 0.152939
R22848 gnd.n4615 gnd.n4614 0.152939
R22849 gnd.n4614 gnd.n1588 0.152939
R22850 gnd.n4610 gnd.n1588 0.152939
R22851 gnd.n4610 gnd.n4609 0.152939
R22852 gnd.n4609 gnd.n4608 0.152939
R22853 gnd.n4608 gnd.n1593 0.152939
R22854 gnd.n4604 gnd.n1593 0.152939
R22855 gnd.n4604 gnd.n4603 0.152939
R22856 gnd.n4603 gnd.n4602 0.152939
R22857 gnd.n4602 gnd.n1598 0.152939
R22858 gnd.n4598 gnd.n1598 0.152939
R22859 gnd.n4598 gnd.n4597 0.152939
R22860 gnd.n4597 gnd.n4596 0.152939
R22861 gnd.n4596 gnd.n1603 0.152939
R22862 gnd.n4592 gnd.n1603 0.152939
R22863 gnd.n4592 gnd.n4591 0.152939
R22864 gnd.n4591 gnd.n4590 0.152939
R22865 gnd.n4590 gnd.n1608 0.152939
R22866 gnd.n4586 gnd.n1608 0.152939
R22867 gnd.n4586 gnd.n4585 0.152939
R22868 gnd.n4584 gnd.n1613 0.152939
R22869 gnd.n4580 gnd.n1613 0.152939
R22870 gnd.n4580 gnd.n4579 0.152939
R22871 gnd.n4579 gnd.n4578 0.152939
R22872 gnd.n4578 gnd.n1618 0.152939
R22873 gnd.n4574 gnd.n1618 0.152939
R22874 gnd.n4186 gnd.n4185 0.152939
R22875 gnd.n4186 gnd.n1968 0.152939
R22876 gnd.n4192 gnd.n1968 0.152939
R22877 gnd.n4193 gnd.n4192 0.152939
R22878 gnd.n4194 gnd.n4193 0.152939
R22879 gnd.n4194 gnd.n1963 0.152939
R22880 gnd.n4207 gnd.n1963 0.152939
R22881 gnd.n4208 gnd.n4207 0.152939
R22882 gnd.n4209 gnd.n4208 0.152939
R22883 gnd.n4209 gnd.n1956 0.152939
R22884 gnd.n4245 gnd.n1956 0.152939
R22885 gnd.n4245 gnd.n4244 0.152939
R22886 gnd.n4244 gnd.n4243 0.152939
R22887 gnd.n4243 gnd.n1957 0.152939
R22888 gnd.n4239 gnd.n1957 0.152939
R22889 gnd.n4239 gnd.n4238 0.152939
R22890 gnd.n4238 gnd.n4237 0.152939
R22891 gnd.n4237 gnd.n1939 0.152939
R22892 gnd.n4276 gnd.n1939 0.152939
R22893 gnd.n4277 gnd.n4276 0.152939
R22894 gnd.n4286 gnd.n4277 0.152939
R22895 gnd.n4286 gnd.n4285 0.152939
R22896 gnd.n4285 gnd.n4284 0.152939
R22897 gnd.n4284 gnd.n4278 0.152939
R22898 gnd.n4280 gnd.n4278 0.152939
R22899 gnd.n4280 gnd.n79 0.152939
R22900 gnd.n3212 gnd.n3211 0.128549
R22901 gnd.n4574 gnd.n4573 0.128549
R22902 gnd.n2973 gnd.n1254 0.10111
R22903 gnd.n4265 gnd.n95 0.10111
R22904 gnd.n5933 gnd.n5325 0.0767195
R22905 gnd.n5849 gnd.n5325 0.0767195
R22906 gnd.n7672 gnd.n93 0.0767195
R22907 gnd.n7672 gnd.n94 0.0767195
R22908 gnd.n4903 gnd.n1253 0.0767195
R22909 gnd.n4903 gnd.n1251 0.0767195
R22910 gnd.n7682 gnd.n7681 0.0695946
R22911 gnd.n2942 gnd.n2939 0.0695946
R22912 gnd.n2944 gnd.n2942 0.0695946
R22913 gnd.n7682 gnd.n79 0.0695946
R22914 gnd.n3211 gnd.n2554 0.063
R22915 gnd.n4573 gnd.n1623 0.063
R22916 gnd.n385 gnd.n95 0.0523293
R22917 gnd.n2906 gnd.n1254 0.0523293
R22918 gnd.n6438 gnd.n5128 0.0477147
R22919 gnd.n1791 gnd.n1623 0.0477147
R22920 gnd.n7490 gnd.n207 0.0477147
R22921 gnd.n4973 gnd.n4972 0.0477147
R22922 gnd.n2554 gnd.n1371 0.0477147
R22923 gnd.n5599 gnd.n5495 0.0442063
R22924 gnd.n5613 gnd.n5495 0.0442063
R22925 gnd.n5614 gnd.n5613 0.0442063
R22926 gnd.n5615 gnd.n5614 0.0442063
R22927 gnd.n5615 gnd.n5483 0.0442063
R22928 gnd.n5629 gnd.n5483 0.0442063
R22929 gnd.n5630 gnd.n5629 0.0442063
R22930 gnd.n5631 gnd.n5630 0.0442063
R22931 gnd.n5631 gnd.n5470 0.0442063
R22932 gnd.n5727 gnd.n5470 0.0442063
R22933 gnd.n5730 gnd.n5729 0.0344674
R22934 gnd.n4395 gnd.n1791 0.0344674
R22935 gnd.n4395 gnd.n1793 0.0344674
R22936 gnd.n1818 gnd.n1793 0.0344674
R22937 gnd.n1819 gnd.n1818 0.0344674
R22938 gnd.n1820 gnd.n1819 0.0344674
R22939 gnd.n1821 gnd.n1820 0.0344674
R22940 gnd.n4201 gnd.n1821 0.0344674
R22941 gnd.n4201 gnd.n1839 0.0344674
R22942 gnd.n1840 gnd.n1839 0.0344674
R22943 gnd.n1841 gnd.n1840 0.0344674
R22944 gnd.n4216 gnd.n1841 0.0344674
R22945 gnd.n4216 gnd.n1859 0.0344674
R22946 gnd.n1860 gnd.n1859 0.0344674
R22947 gnd.n1861 gnd.n1860 0.0344674
R22948 gnd.n4223 gnd.n1861 0.0344674
R22949 gnd.n4223 gnd.n1879 0.0344674
R22950 gnd.n1880 gnd.n1879 0.0344674
R22951 gnd.n1881 gnd.n1880 0.0344674
R22952 gnd.n4229 gnd.n1881 0.0344674
R22953 gnd.n4229 gnd.n1899 0.0344674
R22954 gnd.n1900 gnd.n1899 0.0344674
R22955 gnd.n1901 gnd.n1900 0.0344674
R22956 gnd.n4294 gnd.n1901 0.0344674
R22957 gnd.n4295 gnd.n4294 0.0344674
R22958 gnd.n4295 gnd.n1932 0.0344674
R22959 gnd.n1933 gnd.n1932 0.0344674
R22960 gnd.n1934 gnd.n1933 0.0344674
R22961 gnd.n4303 gnd.n1934 0.0344674
R22962 gnd.n4303 gnd.n4302 0.0344674
R22963 gnd.n4302 gnd.n379 0.0344674
R22964 gnd.n379 gnd.n109 0.0344674
R22965 gnd.n110 gnd.n109 0.0344674
R22966 gnd.n111 gnd.n110 0.0344674
R22967 gnd.n373 gnd.n111 0.0344674
R22968 gnd.n373 gnd.n127 0.0344674
R22969 gnd.n128 gnd.n127 0.0344674
R22970 gnd.n129 gnd.n128 0.0344674
R22971 gnd.n367 gnd.n129 0.0344674
R22972 gnd.n367 gnd.n148 0.0344674
R22973 gnd.n149 gnd.n148 0.0344674
R22974 gnd.n150 gnd.n149 0.0344674
R22975 gnd.n361 gnd.n150 0.0344674
R22976 gnd.n361 gnd.n167 0.0344674
R22977 gnd.n168 gnd.n167 0.0344674
R22978 gnd.n169 gnd.n168 0.0344674
R22979 gnd.n7421 gnd.n169 0.0344674
R22980 gnd.n7421 gnd.n187 0.0344674
R22981 gnd.n188 gnd.n187 0.0344674
R22982 gnd.n189 gnd.n188 0.0344674
R22983 gnd.n7422 gnd.n189 0.0344674
R22984 gnd.n7422 gnd.n205 0.0344674
R22985 gnd.n206 gnd.n205 0.0344674
R22986 gnd.n207 gnd.n206 0.0344674
R22987 gnd.n4972 gnd.n1138 0.0344674
R22988 gnd.n2826 gnd.n1138 0.0344674
R22989 gnd.n2826 gnd.n1160 0.0344674
R22990 gnd.n1161 gnd.n1160 0.0344674
R22991 gnd.n1162 gnd.n1161 0.0344674
R22992 gnd.n2832 gnd.n1162 0.0344674
R22993 gnd.n2832 gnd.n1179 0.0344674
R22994 gnd.n1180 gnd.n1179 0.0344674
R22995 gnd.n1181 gnd.n1180 0.0344674
R22996 gnd.n2839 gnd.n1181 0.0344674
R22997 gnd.n2839 gnd.n1199 0.0344674
R22998 gnd.n1200 gnd.n1199 0.0344674
R22999 gnd.n1201 gnd.n1200 0.0344674
R23000 gnd.n2855 gnd.n1201 0.0344674
R23001 gnd.n2855 gnd.n1219 0.0344674
R23002 gnd.n1220 gnd.n1219 0.0344674
R23003 gnd.n1221 gnd.n1220 0.0344674
R23004 gnd.n2858 gnd.n1221 0.0344674
R23005 gnd.n2858 gnd.n1240 0.0344674
R23006 gnd.n1241 gnd.n1240 0.0344674
R23007 gnd.n1242 gnd.n1241 0.0344674
R23008 gnd.n2706 gnd.n1242 0.0344674
R23009 gnd.n2706 gnd.n2705 0.0344674
R23010 gnd.n2927 gnd.n2705 0.0344674
R23011 gnd.n2928 gnd.n2927 0.0344674
R23012 gnd.n2928 gnd.n2690 0.0344674
R23013 gnd.n2690 gnd.n2686 0.0344674
R23014 gnd.n2687 gnd.n2686 0.0344674
R23015 gnd.n2956 gnd.n2687 0.0344674
R23016 gnd.n2956 gnd.n2688 0.0344674
R23017 gnd.n2688 gnd.n1269 0.0344674
R23018 gnd.n1270 gnd.n1269 0.0344674
R23019 gnd.n1271 gnd.n1270 0.0344674
R23020 gnd.n3008 gnd.n1271 0.0344674
R23021 gnd.n3008 gnd.n1288 0.0344674
R23022 gnd.n1289 gnd.n1288 0.0344674
R23023 gnd.n1290 gnd.n1289 0.0344674
R23024 gnd.n3023 gnd.n1290 0.0344674
R23025 gnd.n3023 gnd.n1308 0.0344674
R23026 gnd.n1309 gnd.n1308 0.0344674
R23027 gnd.n1310 gnd.n1309 0.0344674
R23028 gnd.n3030 gnd.n1310 0.0344674
R23029 gnd.n3030 gnd.n1328 0.0344674
R23030 gnd.n1329 gnd.n1328 0.0344674
R23031 gnd.n1330 gnd.n1329 0.0344674
R23032 gnd.n2635 gnd.n1330 0.0344674
R23033 gnd.n2635 gnd.n1348 0.0344674
R23034 gnd.n1349 gnd.n1348 0.0344674
R23035 gnd.n1350 gnd.n1349 0.0344674
R23036 gnd.n2630 gnd.n1350 0.0344674
R23037 gnd.n2630 gnd.n1369 0.0344674
R23038 gnd.n1370 gnd.n1369 0.0344674
R23039 gnd.n1371 gnd.n1370 0.0344674
R23040 gnd.n3210 gnd.n3209 0.0344674
R23041 gnd.n4572 gnd.n4571 0.0344674
R23042 gnd.n3158 gnd.n3148 0.029712
R23043 gnd.n4184 gnd.n4183 0.029712
R23044 gnd.n5463 gnd.n5462 0.0269946
R23045 gnd.n5740 gnd.n5460 0.0269946
R23046 gnd.n5739 gnd.n5461 0.0269946
R23047 gnd.n5759 gnd.n5442 0.0269946
R23048 gnd.n5761 gnd.n5760 0.0269946
R23049 gnd.n5762 gnd.n5440 0.0269946
R23050 gnd.n5769 gnd.n5765 0.0269946
R23051 gnd.n5768 gnd.n5767 0.0269946
R23052 gnd.n5766 gnd.n5419 0.0269946
R23053 gnd.n5793 gnd.n5420 0.0269946
R23054 gnd.n5792 gnd.n5421 0.0269946
R23055 gnd.n5825 gnd.n5395 0.0269946
R23056 gnd.n5827 gnd.n5826 0.0269946
R23057 gnd.n5828 gnd.n5387 0.0269946
R23058 gnd.n5391 gnd.n5388 0.0269946
R23059 gnd.n5838 gnd.n5389 0.0269946
R23060 gnd.n5837 gnd.n5390 0.0269946
R23061 gnd.n5883 gnd.n5363 0.0269946
R23062 gnd.n5885 gnd.n5884 0.0269946
R23063 gnd.n5894 gnd.n5356 0.0269946
R23064 gnd.n5896 gnd.n5895 0.0269946
R23065 gnd.n5897 gnd.n5354 0.0269946
R23066 gnd.n5904 gnd.n5900 0.0269946
R23067 gnd.n5903 gnd.n5902 0.0269946
R23068 gnd.n5901 gnd.n5333 0.0269946
R23069 gnd.n5926 gnd.n5334 0.0269946
R23070 gnd.n5925 gnd.n5335 0.0269946
R23071 gnd.n5968 gnd.n5244 0.0269946
R23072 gnd.n5970 gnd.n5969 0.0269946
R23073 gnd.n5979 gnd.n5237 0.0269946
R23074 gnd.n5981 gnd.n5980 0.0269946
R23075 gnd.n5982 gnd.n5235 0.0269946
R23076 gnd.n5988 gnd.n5985 0.0269946
R23077 gnd.n5987 gnd.n5986 0.0269946
R23078 gnd.n6013 gnd.n5215 0.0269946
R23079 gnd.n6012 gnd.n5216 0.0269946
R23080 gnd.n6042 gnd.n5201 0.0269946
R23081 gnd.n6044 gnd.n6043 0.0269946
R23082 gnd.n6068 gnd.n5187 0.0269946
R23083 gnd.n6070 gnd.n6069 0.0269946
R23084 gnd.n6071 gnd.n974 0.0269946
R23085 gnd.n5182 gnd.n975 0.0269946
R23086 gnd.n5184 gnd.n976 0.0269946
R23087 gnd.n6079 gnd.n6078 0.0269946
R23088 gnd.n6081 gnd.n6080 0.0269946
R23089 gnd.n6082 gnd.n997 0.0269946
R23090 gnd.n6083 gnd.n998 0.0269946
R23091 gnd.n6084 gnd.n999 0.0269946
R23092 gnd.n6344 gnd.n6343 0.0269946
R23093 gnd.n6345 gnd.n1023 0.0269946
R23094 gnd.n6346 gnd.n1024 0.0269946
R23095 gnd.n6347 gnd.n1025 0.0269946
R23096 gnd.n3206 gnd.n2555 0.0225788
R23097 gnd.n3205 gnd.n2559 0.0225788
R23098 gnd.n3202 gnd.n3201 0.0225788
R23099 gnd.n3198 gnd.n2565 0.0225788
R23100 gnd.n3197 gnd.n2571 0.0225788
R23101 gnd.n3194 gnd.n3193 0.0225788
R23102 gnd.n3190 gnd.n2577 0.0225788
R23103 gnd.n3189 gnd.n2581 0.0225788
R23104 gnd.n3186 gnd.n3185 0.0225788
R23105 gnd.n3182 gnd.n2588 0.0225788
R23106 gnd.n3181 gnd.n2594 0.0225788
R23107 gnd.n3178 gnd.n3177 0.0225788
R23108 gnd.n3174 gnd.n2600 0.0225788
R23109 gnd.n3173 gnd.n2604 0.0225788
R23110 gnd.n3170 gnd.n3169 0.0225788
R23111 gnd.n3166 gnd.n2611 0.0225788
R23112 gnd.n3165 gnd.n2618 0.0225788
R23113 gnd.n2626 gnd.n2624 0.0225788
R23114 gnd.n3159 gnd.n3158 0.0225788
R23115 gnd.n4568 gnd.n1624 0.0225788
R23116 gnd.n4567 gnd.n1628 0.0225788
R23117 gnd.n4564 gnd.n4563 0.0225788
R23118 gnd.n4560 gnd.n1633 0.0225788
R23119 gnd.n4559 gnd.n1637 0.0225788
R23120 gnd.n4556 gnd.n4555 0.0225788
R23121 gnd.n4552 gnd.n1641 0.0225788
R23122 gnd.n4551 gnd.n1645 0.0225788
R23123 gnd.n4548 gnd.n4547 0.0225788
R23124 gnd.n4544 gnd.n1649 0.0225788
R23125 gnd.n4543 gnd.n1653 0.0225788
R23126 gnd.n4540 gnd.n4539 0.0225788
R23127 gnd.n4536 gnd.n1657 0.0225788
R23128 gnd.n4535 gnd.n1661 0.0225788
R23129 gnd.n4532 gnd.n4531 0.0225788
R23130 gnd.n4528 gnd.n1665 0.0225788
R23131 gnd.n4527 gnd.n1671 0.0225788
R23132 gnd.n1974 gnd.n1674 0.0225788
R23133 gnd.n4183 gnd.n1973 0.0225788
R23134 gnd.n4184 gnd.n1972 0.0218415
R23135 gnd.n3155 gnd.n3148 0.0218415
R23136 gnd.n5729 gnd.n5728 0.0202011
R23137 gnd.n5728 gnd.n5727 0.0148637
R23138 gnd.n6341 gnd.n6085 0.0144266
R23139 gnd.n6342 gnd.n6341 0.0130679
R23140 gnd.n3209 gnd.n2555 0.0123886
R23141 gnd.n3206 gnd.n3205 0.0123886
R23142 gnd.n3202 gnd.n2559 0.0123886
R23143 gnd.n3201 gnd.n2565 0.0123886
R23144 gnd.n3198 gnd.n3197 0.0123886
R23145 gnd.n3194 gnd.n2571 0.0123886
R23146 gnd.n3193 gnd.n2577 0.0123886
R23147 gnd.n3190 gnd.n3189 0.0123886
R23148 gnd.n3186 gnd.n2581 0.0123886
R23149 gnd.n3185 gnd.n2588 0.0123886
R23150 gnd.n3182 gnd.n3181 0.0123886
R23151 gnd.n3178 gnd.n2594 0.0123886
R23152 gnd.n3177 gnd.n2600 0.0123886
R23153 gnd.n3174 gnd.n3173 0.0123886
R23154 gnd.n3170 gnd.n2604 0.0123886
R23155 gnd.n3169 gnd.n2611 0.0123886
R23156 gnd.n3166 gnd.n3165 0.0123886
R23157 gnd.n2624 gnd.n2618 0.0123886
R23158 gnd.n3159 gnd.n2626 0.0123886
R23159 gnd.n4571 gnd.n1624 0.0123886
R23160 gnd.n4568 gnd.n4567 0.0123886
R23161 gnd.n4564 gnd.n1628 0.0123886
R23162 gnd.n4563 gnd.n1633 0.0123886
R23163 gnd.n4560 gnd.n4559 0.0123886
R23164 gnd.n4556 gnd.n1637 0.0123886
R23165 gnd.n4555 gnd.n1641 0.0123886
R23166 gnd.n4552 gnd.n4551 0.0123886
R23167 gnd.n4548 gnd.n1645 0.0123886
R23168 gnd.n4547 gnd.n1649 0.0123886
R23169 gnd.n4544 gnd.n4543 0.0123886
R23170 gnd.n4540 gnd.n1653 0.0123886
R23171 gnd.n4539 gnd.n1657 0.0123886
R23172 gnd.n4536 gnd.n4535 0.0123886
R23173 gnd.n4532 gnd.n1661 0.0123886
R23174 gnd.n4531 gnd.n1665 0.0123886
R23175 gnd.n4528 gnd.n4527 0.0123886
R23176 gnd.n1674 gnd.n1671 0.0123886
R23177 gnd.n1974 gnd.n1973 0.0123886
R23178 gnd.n5730 gnd.n5463 0.00797283
R23179 gnd.n5462 gnd.n5460 0.00797283
R23180 gnd.n5740 gnd.n5739 0.00797283
R23181 gnd.n5461 gnd.n5442 0.00797283
R23182 gnd.n5760 gnd.n5759 0.00797283
R23183 gnd.n5762 gnd.n5761 0.00797283
R23184 gnd.n5765 gnd.n5440 0.00797283
R23185 gnd.n5769 gnd.n5768 0.00797283
R23186 gnd.n5767 gnd.n5766 0.00797283
R23187 gnd.n5420 gnd.n5419 0.00797283
R23188 gnd.n5793 gnd.n5792 0.00797283
R23189 gnd.n5421 gnd.n5395 0.00797283
R23190 gnd.n5826 gnd.n5825 0.00797283
R23191 gnd.n5828 gnd.n5827 0.00797283
R23192 gnd.n5391 gnd.n5387 0.00797283
R23193 gnd.n5389 gnd.n5388 0.00797283
R23194 gnd.n5838 gnd.n5837 0.00797283
R23195 gnd.n5390 gnd.n5363 0.00797283
R23196 gnd.n5885 gnd.n5883 0.00797283
R23197 gnd.n5884 gnd.n5356 0.00797283
R23198 gnd.n5895 gnd.n5894 0.00797283
R23199 gnd.n5897 gnd.n5896 0.00797283
R23200 gnd.n5900 gnd.n5354 0.00797283
R23201 gnd.n5904 gnd.n5903 0.00797283
R23202 gnd.n5902 gnd.n5901 0.00797283
R23203 gnd.n5334 gnd.n5333 0.00797283
R23204 gnd.n5926 gnd.n5925 0.00797283
R23205 gnd.n5335 gnd.n5244 0.00797283
R23206 gnd.n5970 gnd.n5968 0.00797283
R23207 gnd.n5969 gnd.n5237 0.00797283
R23208 gnd.n5980 gnd.n5979 0.00797283
R23209 gnd.n5982 gnd.n5981 0.00797283
R23210 gnd.n5985 gnd.n5235 0.00797283
R23211 gnd.n5988 gnd.n5987 0.00797283
R23212 gnd.n5986 gnd.n5215 0.00797283
R23213 gnd.n6013 gnd.n6012 0.00797283
R23214 gnd.n5216 gnd.n5201 0.00797283
R23215 gnd.n6044 gnd.n6042 0.00797283
R23216 gnd.n6043 gnd.n5187 0.00797283
R23217 gnd.n6069 gnd.n6068 0.00797283
R23218 gnd.n6071 gnd.n6070 0.00797283
R23219 gnd.n5182 gnd.n974 0.00797283
R23220 gnd.n5184 gnd.n975 0.00797283
R23221 gnd.n6078 gnd.n976 0.00797283
R23222 gnd.n6080 gnd.n6079 0.00797283
R23223 gnd.n6082 gnd.n6081 0.00797283
R23224 gnd.n6083 gnd.n997 0.00797283
R23225 gnd.n6084 gnd.n998 0.00797283
R23226 gnd.n6085 gnd.n999 0.00797283
R23227 gnd.n6343 gnd.n6342 0.00797283
R23228 gnd.n6345 gnd.n6344 0.00797283
R23229 gnd.n6346 gnd.n1023 0.00797283
R23230 gnd.n6347 gnd.n1024 0.00797283
R23231 gnd.n5128 gnd.n1025 0.00797283
R23232 gnd.n3211 gnd.n3210 0.00593478
R23233 gnd.n4573 gnd.n4572 0.00593478
R23234 a_n2318_8322.n9 a_n2318_8322.t7 74.6477
R23235 a_n2318_8322.t26 a_n2318_8322.n22 74.6477
R23236 a_n2318_8322.n1 a_n2318_8322.t25 74.6474
R23237 a_n2318_8322.n16 a_n2318_8322.t12 74.2899
R23238 a_n2318_8322.n6 a_n2318_8322.t15 74.2899
R23239 a_n2318_8322.n10 a_n2318_8322.t5 74.2899
R23240 a_n2318_8322.n11 a_n2318_8322.t8 74.2899
R23241 a_n2318_8322.n14 a_n2318_8322.t9 74.2899
R23242 a_n2318_8322.n22 a_n2318_8322.n21 70.6783
R23243 a_n2318_8322.n20 a_n2318_8322.n19 70.6783
R23244 a_n2318_8322.n18 a_n2318_8322.n17 70.6783
R23245 a_n2318_8322.n1 a_n2318_8322.n0 70.6783
R23246 a_n2318_8322.n3 a_n2318_8322.n2 70.6783
R23247 a_n2318_8322.n5 a_n2318_8322.n4 70.6783
R23248 a_n2318_8322.n9 a_n2318_8322.n8 70.6783
R23249 a_n2318_8322.n13 a_n2318_8322.n12 70.6783
R23250 a_n2318_8322.n16 a_n2318_8322.n15 23.4712
R23251 a_n2318_8322.n7 a_n2318_8322.t1 9.85987
R23252 a_n2318_8322.n15 a_n2318_8322.n14 6.95632
R23253 a_n2318_8322.n7 a_n2318_8322.n6 6.19447
R23254 a_n2318_8322.n15 a_n2318_8322.n7 5.3452
R23255 a_n2318_8322.n21 a_n2318_8322.t14 3.61217
R23256 a_n2318_8322.n21 a_n2318_8322.t13 3.61217
R23257 a_n2318_8322.n19 a_n2318_8322.t23 3.61217
R23258 a_n2318_8322.n19 a_n2318_8322.t18 3.61217
R23259 a_n2318_8322.n17 a_n2318_8322.t21 3.61217
R23260 a_n2318_8322.n17 a_n2318_8322.t20 3.61217
R23261 a_n2318_8322.n0 a_n2318_8322.t22 3.61217
R23262 a_n2318_8322.n0 a_n2318_8322.t19 3.61217
R23263 a_n2318_8322.n2 a_n2318_8322.t16 3.61217
R23264 a_n2318_8322.n2 a_n2318_8322.t27 3.61217
R23265 a_n2318_8322.n4 a_n2318_8322.t24 3.61217
R23266 a_n2318_8322.n4 a_n2318_8322.t17 3.61217
R23267 a_n2318_8322.n8 a_n2318_8322.t11 3.61217
R23268 a_n2318_8322.n8 a_n2318_8322.t10 3.61217
R23269 a_n2318_8322.n12 a_n2318_8322.t6 3.61217
R23270 a_n2318_8322.n12 a_n2318_8322.t4 3.61217
R23271 a_n2318_8322.n6 a_n2318_8322.n5 0.358259
R23272 a_n2318_8322.n5 a_n2318_8322.n3 0.358259
R23273 a_n2318_8322.n3 a_n2318_8322.n1 0.358259
R23274 a_n2318_8322.n14 a_n2318_8322.n13 0.358259
R23275 a_n2318_8322.n13 a_n2318_8322.n11 0.358259
R23276 a_n2318_8322.n10 a_n2318_8322.n9 0.358259
R23277 a_n2318_8322.n18 a_n2318_8322.n16 0.358259
R23278 a_n2318_8322.n20 a_n2318_8322.n18 0.358259
R23279 a_n2318_8322.n22 a_n2318_8322.n20 0.358259
R23280 a_n2318_8322.n11 a_n2318_8322.n10 0.101793
R23281 a_n2318_8322.t3 a_n2318_8322.t2 0.0788333
R23282 a_n2318_8322.t0 a_n2318_8322.t3 0.0631667
R23283 a_n2318_8322.t1 a_n2318_8322.t0 0.0471944
R23284 a_n2318_8322.t1 a_n2318_8322.t2 0.0453889
R23285 plus.n46 plus.t9 252.611
R23286 plus.n9 plus.t11 252.611
R23287 plus.n76 plus.t4 243.97
R23288 plus.n72 plus.t12 231.093
R23289 plus.n35 plus.t7 231.093
R23290 plus.n76 plus.n75 223.454
R23291 plus.n78 plus.n77 223.454
R23292 plus.n47 plus.t5 187.445
R23293 plus.n44 plus.t18 187.445
R23294 plus.n42 plus.t17 187.445
R23295 plus.n59 plus.t13 187.445
R23296 plus.n65 plus.t14 187.445
R23297 plus.n38 plus.t10 187.445
R23298 plus.n1 plus.t6 187.445
R23299 plus.n28 plus.t16 187.445
R23300 plus.n22 plus.t15 187.445
R23301 plus.n5 plus.t20 187.445
R23302 plus.n7 plus.t19 187.445
R23303 plus.n10 plus.t8 187.445
R23304 plus.n73 plus.n72 161.3
R23305 plus.n71 plus.n37 161.3
R23306 plus.n70 plus.n69 161.3
R23307 plus.n68 plus.n67 161.3
R23308 plus.n66 plus.n39 161.3
R23309 plus.n64 plus.n63 161.3
R23310 plus.n62 plus.n40 161.3
R23311 plus.n61 plus.n60 161.3
R23312 plus.n58 plus.n41 161.3
R23313 plus.n57 plus.n56 161.3
R23314 plus.n55 plus.n54 161.3
R23315 plus.n53 plus.n43 161.3
R23316 plus.n52 plus.n51 161.3
R23317 plus.n50 plus.n49 161.3
R23318 plus.n48 plus.n45 161.3
R23319 plus.n11 plus.n8 161.3
R23320 plus.n13 plus.n12 161.3
R23321 plus.n15 plus.n14 161.3
R23322 plus.n16 plus.n6 161.3
R23323 plus.n18 plus.n17 161.3
R23324 plus.n20 plus.n19 161.3
R23325 plus.n21 plus.n4 161.3
R23326 plus.n24 plus.n23 161.3
R23327 plus.n25 plus.n3 161.3
R23328 plus.n27 plus.n26 161.3
R23329 plus.n29 plus.n2 161.3
R23330 plus.n31 plus.n30 161.3
R23331 plus.n33 plus.n32 161.3
R23332 plus.n34 plus.n0 161.3
R23333 plus.n36 plus.n35 161.3
R23334 plus.n49 plus.n48 56.5617
R23335 plus.n58 plus.n57 56.5617
R23336 plus.n67 plus.n66 56.5617
R23337 plus.n30 plus.n29 56.5617
R23338 plus.n21 plus.n20 56.5617
R23339 plus.n12 plus.n11 56.5617
R23340 plus.n71 plus.n70 46.3896
R23341 plus.n34 plus.n33 46.3896
R23342 plus.n46 plus.n45 42.8164
R23343 plus.n9 plus.n8 42.8164
R23344 plus.n54 plus.n53 42.5146
R23345 plus.n60 plus.n40 42.5146
R23346 plus.n23 plus.n3 42.5146
R23347 plus.n17 plus.n16 42.5146
R23348 plus.n53 plus.n52 38.6395
R23349 plus.n64 plus.n40 38.6395
R23350 plus.n27 plus.n3 38.6395
R23351 plus.n16 plus.n15 38.6395
R23352 plus.n47 plus.n46 38.2514
R23353 plus.n10 plus.n9 38.2514
R23354 plus.n74 plus.n73 31.491
R23355 plus.n49 plus.n44 19.9199
R23356 plus.n66 plus.n65 19.9199
R23357 plus.n29 plus.n28 19.9199
R23358 plus.n12 plus.n7 19.9199
R23359 plus.n75 plus.t1 19.8005
R23360 plus.n75 plus.t2 19.8005
R23361 plus.n77 plus.t0 19.8005
R23362 plus.n77 plus.t3 19.8005
R23363 plus.n57 plus.n42 17.9525
R23364 plus.n59 plus.n58 17.9525
R23365 plus.n22 plus.n21 17.9525
R23366 plus.n20 plus.n5 17.9525
R23367 plus.n48 plus.n47 15.9852
R23368 plus.n67 plus.n38 15.9852
R23369 plus.n30 plus.n1 15.9852
R23370 plus.n11 plus.n10 15.9852
R23371 plus.n72 plus.n71 15.3369
R23372 plus.n35 plus.n34 15.3369
R23373 plus plus.n79 14.4284
R23374 plus.n74 plus.n36 11.9494
R23375 plus.n70 plus.n38 8.60764
R23376 plus.n33 plus.n1 8.60764
R23377 plus.n54 plus.n42 6.6403
R23378 plus.n60 plus.n59 6.6403
R23379 plus.n23 plus.n22 6.6403
R23380 plus.n17 plus.n5 6.6403
R23381 plus.n79 plus.n78 5.40567
R23382 plus.n52 plus.n44 4.67295
R23383 plus.n65 plus.n64 4.67295
R23384 plus.n28 plus.n27 4.67295
R23385 plus.n15 plus.n7 4.67295
R23386 plus.n79 plus.n74 1.188
R23387 plus.n78 plus.n76 0.716017
R23388 plus.n50 plus.n45 0.189894
R23389 plus.n51 plus.n50 0.189894
R23390 plus.n51 plus.n43 0.189894
R23391 plus.n55 plus.n43 0.189894
R23392 plus.n56 plus.n55 0.189894
R23393 plus.n56 plus.n41 0.189894
R23394 plus.n61 plus.n41 0.189894
R23395 plus.n62 plus.n61 0.189894
R23396 plus.n63 plus.n62 0.189894
R23397 plus.n63 plus.n39 0.189894
R23398 plus.n68 plus.n39 0.189894
R23399 plus.n69 plus.n68 0.189894
R23400 plus.n69 plus.n37 0.189894
R23401 plus.n73 plus.n37 0.189894
R23402 plus.n36 plus.n0 0.189894
R23403 plus.n32 plus.n0 0.189894
R23404 plus.n32 plus.n31 0.189894
R23405 plus.n31 plus.n2 0.189894
R23406 plus.n26 plus.n2 0.189894
R23407 plus.n26 plus.n25 0.189894
R23408 plus.n25 plus.n24 0.189894
R23409 plus.n24 plus.n4 0.189894
R23410 plus.n19 plus.n4 0.189894
R23411 plus.n19 plus.n18 0.189894
R23412 plus.n18 plus.n6 0.189894
R23413 plus.n14 plus.n6 0.189894
R23414 plus.n14 plus.n13 0.189894
R23415 plus.n13 plus.n8 0.189894
R23416 a_n2903_n3924.n0 a_n2903_n3924.t27 214.981
R23417 a_n2903_n3924.n2 a_n2903_n3924.t37 214.452
R23418 a_n2903_n3924.n11 a_n2903_n3924.t25 214.321
R23419 a_n2903_n3924.n12 a_n2903_n3924.t29 214.321
R23420 a_n2903_n3924.n13 a_n2903_n3924.t31 214.321
R23421 a_n2903_n3924.n14 a_n2903_n3924.t28 214.321
R23422 a_n2903_n3924.n15 a_n2903_n3924.t7 214.321
R23423 a_n2903_n3924.n0 a_n2903_n3924.t36 214.321
R23424 a_n2903_n3924.n1 a_n2903_n3924.t19 55.8337
R23425 a_n2903_n3924.n3 a_n2903_n3924.t6 55.8337
R23426 a_n2903_n3924.n10 a_n2903_n3924.t4 55.8337
R23427 a_n2903_n3924.n34 a_n2903_n3924.t16 55.8335
R23428 a_n2903_n3924.n32 a_n2903_n3924.t1 55.8335
R23429 a_n2903_n3924.n25 a_n2903_n3924.t5 55.8335
R23430 a_n2903_n3924.n24 a_n2903_n3924.t17 55.8335
R23431 a_n2903_n3924.n17 a_n2903_n3924.t21 55.8335
R23432 a_n2903_n3924.n36 a_n2903_n3924.n35 53.0052
R23433 a_n2903_n3924.n38 a_n2903_n3924.n37 53.0052
R23434 a_n2903_n3924.n5 a_n2903_n3924.n4 53.0052
R23435 a_n2903_n3924.n7 a_n2903_n3924.n6 53.0052
R23436 a_n2903_n3924.n9 a_n2903_n3924.n8 53.0052
R23437 a_n2903_n3924.n31 a_n2903_n3924.n30 53.0051
R23438 a_n2903_n3924.n29 a_n2903_n3924.n28 53.0051
R23439 a_n2903_n3924.n27 a_n2903_n3924.n26 53.0051
R23440 a_n2903_n3924.n23 a_n2903_n3924.n22 53.0051
R23441 a_n2903_n3924.n21 a_n2903_n3924.n20 53.0051
R23442 a_n2903_n3924.n19 a_n2903_n3924.n18 53.0051
R23443 a_n2903_n3924.n40 a_n2903_n3924.n39 53.0051
R23444 a_n2903_n3924.n16 a_n2903_n3924.n10 12.2417
R23445 a_n2903_n3924.n34 a_n2903_n3924.n33 12.2417
R23446 a_n2903_n3924.n17 a_n2903_n3924.n16 5.16214
R23447 a_n2903_n3924.n33 a_n2903_n3924.n32 5.16214
R23448 a_n2903_n3924.n35 a_n2903_n3924.t14 2.82907
R23449 a_n2903_n3924.n35 a_n2903_n3924.t18 2.82907
R23450 a_n2903_n3924.n37 a_n2903_n3924.t11 2.82907
R23451 a_n2903_n3924.n37 a_n2903_n3924.t15 2.82907
R23452 a_n2903_n3924.n4 a_n2903_n3924.t3 2.82907
R23453 a_n2903_n3924.n4 a_n2903_n3924.t35 2.82907
R23454 a_n2903_n3924.n6 a_n2903_n3924.t32 2.82907
R23455 a_n2903_n3924.n6 a_n2903_n3924.t39 2.82907
R23456 a_n2903_n3924.n8 a_n2903_n3924.t38 2.82907
R23457 a_n2903_n3924.n8 a_n2903_n3924.t34 2.82907
R23458 a_n2903_n3924.n30 a_n2903_n3924.t2 2.82907
R23459 a_n2903_n3924.n30 a_n2903_n3924.t24 2.82907
R23460 a_n2903_n3924.n28 a_n2903_n3924.t0 2.82907
R23461 a_n2903_n3924.n28 a_n2903_n3924.t26 2.82907
R23462 a_n2903_n3924.n26 a_n2903_n3924.t30 2.82907
R23463 a_n2903_n3924.n26 a_n2903_n3924.t33 2.82907
R23464 a_n2903_n3924.n22 a_n2903_n3924.t9 2.82907
R23465 a_n2903_n3924.n22 a_n2903_n3924.t20 2.82907
R23466 a_n2903_n3924.n20 a_n2903_n3924.t13 2.82907
R23467 a_n2903_n3924.n20 a_n2903_n3924.t8 2.82907
R23468 a_n2903_n3924.n18 a_n2903_n3924.t22 2.82907
R23469 a_n2903_n3924.n18 a_n2903_n3924.t12 2.82907
R23470 a_n2903_n3924.t23 a_n2903_n3924.n40 2.82907
R23471 a_n2903_n3924.n40 a_n2903_n3924.t10 2.82907
R23472 a_n2903_n3924.n33 a_n2903_n3924.n2 1.95694
R23473 a_n2903_n3924.n16 a_n2903_n3924.n0 1.95694
R23474 a_n2903_n3924.n0 a_n2903_n3924.n15 0.684366
R23475 a_n2903_n3924.n15 a_n2903_n3924.n14 0.672012
R23476 a_n2903_n3924.n14 a_n2903_n3924.n13 0.672012
R23477 a_n2903_n3924.n13 a_n2903_n3924.n12 0.672012
R23478 a_n2903_n3924.n12 a_n2903_n3924.n11 0.672012
R23479 a_n2903_n3924.n11 a_n2903_n3924.n2 0.541924
R23480 a_n2903_n3924.n19 a_n2903_n3924.n17 0.530672
R23481 a_n2903_n3924.n21 a_n2903_n3924.n19 0.530672
R23482 a_n2903_n3924.n23 a_n2903_n3924.n21 0.530672
R23483 a_n2903_n3924.n24 a_n2903_n3924.n23 0.530672
R23484 a_n2903_n3924.n27 a_n2903_n3924.n25 0.530672
R23485 a_n2903_n3924.n29 a_n2903_n3924.n27 0.530672
R23486 a_n2903_n3924.n31 a_n2903_n3924.n29 0.530672
R23487 a_n2903_n3924.n32 a_n2903_n3924.n31 0.530672
R23488 a_n2903_n3924.n10 a_n2903_n3924.n9 0.530672
R23489 a_n2903_n3924.n9 a_n2903_n3924.n7 0.530672
R23490 a_n2903_n3924.n7 a_n2903_n3924.n5 0.530672
R23491 a_n2903_n3924.n5 a_n2903_n3924.n3 0.530672
R23492 a_n2903_n3924.n39 a_n2903_n3924.n1 0.530672
R23493 a_n2903_n3924.n39 a_n2903_n3924.n38 0.530672
R23494 a_n2903_n3924.n38 a_n2903_n3924.n36 0.530672
R23495 a_n2903_n3924.n36 a_n2903_n3924.n34 0.530672
R23496 a_n2903_n3924.n25 a_n2903_n3924.n24 0.235414
R23497 a_n2903_n3924.n3 a_n2903_n3924.n1 0.235414
R23498 minus.n46 minus.t20 252.611
R23499 minus.n9 minus.t13 252.611
R23500 minus.n78 minus.t3 243.255
R23501 minus.n72 minus.t15 231.093
R23502 minus.n35 minus.t17 231.093
R23503 minus.n77 minus.n75 224.169
R23504 minus.n77 minus.n76 223.454
R23505 minus.n38 minus.t12 187.445
R23506 minus.n65 minus.t7 187.445
R23507 minus.n59 minus.t6 187.445
R23508 minus.n42 minus.t11 187.445
R23509 minus.n44 minus.t10 187.445
R23510 minus.n47 minus.t16 187.445
R23511 minus.n10 minus.t9 187.445
R23512 minus.n7 minus.t8 187.445
R23513 minus.n5 minus.t5 187.445
R23514 minus.n22 minus.t18 187.445
R23515 minus.n28 minus.t19 187.445
R23516 minus.n1 minus.t14 187.445
R23517 minus.n48 minus.n45 161.3
R23518 minus.n50 minus.n49 161.3
R23519 minus.n52 minus.n51 161.3
R23520 minus.n53 minus.n43 161.3
R23521 minus.n55 minus.n54 161.3
R23522 minus.n57 minus.n56 161.3
R23523 minus.n58 minus.n41 161.3
R23524 minus.n61 minus.n60 161.3
R23525 minus.n62 minus.n40 161.3
R23526 minus.n64 minus.n63 161.3
R23527 minus.n66 minus.n39 161.3
R23528 minus.n68 minus.n67 161.3
R23529 minus.n70 minus.n69 161.3
R23530 minus.n71 minus.n37 161.3
R23531 minus.n73 minus.n72 161.3
R23532 minus.n36 minus.n35 161.3
R23533 minus.n34 minus.n0 161.3
R23534 minus.n33 minus.n32 161.3
R23535 minus.n31 minus.n30 161.3
R23536 minus.n29 minus.n2 161.3
R23537 minus.n27 minus.n26 161.3
R23538 minus.n25 minus.n3 161.3
R23539 minus.n24 minus.n23 161.3
R23540 minus.n21 minus.n4 161.3
R23541 minus.n20 minus.n19 161.3
R23542 minus.n18 minus.n17 161.3
R23543 minus.n16 minus.n6 161.3
R23544 minus.n15 minus.n14 161.3
R23545 minus.n13 minus.n12 161.3
R23546 minus.n11 minus.n8 161.3
R23547 minus.n67 minus.n66 56.5617
R23548 minus.n58 minus.n57 56.5617
R23549 minus.n49 minus.n48 56.5617
R23550 minus.n12 minus.n11 56.5617
R23551 minus.n21 minus.n20 56.5617
R23552 minus.n30 minus.n29 56.5617
R23553 minus.n71 minus.n70 46.3896
R23554 minus.n34 minus.n33 46.3896
R23555 minus.n46 minus.n45 42.8164
R23556 minus.n9 minus.n8 42.8164
R23557 minus.n60 minus.n40 42.5146
R23558 minus.n54 minus.n53 42.5146
R23559 minus.n17 minus.n16 42.5146
R23560 minus.n23 minus.n3 42.5146
R23561 minus.n64 minus.n40 38.6395
R23562 minus.n53 minus.n52 38.6395
R23563 minus.n16 minus.n15 38.6395
R23564 minus.n27 minus.n3 38.6395
R23565 minus.n47 minus.n46 38.2514
R23566 minus.n10 minus.n9 38.2514
R23567 minus.n74 minus.n73 31.7069
R23568 minus.n66 minus.n65 19.9199
R23569 minus.n49 minus.n44 19.9199
R23570 minus.n12 minus.n7 19.9199
R23571 minus.n29 minus.n28 19.9199
R23572 minus.n76 minus.t2 19.8005
R23573 minus.n76 minus.t0 19.8005
R23574 minus.n75 minus.t1 19.8005
R23575 minus.n75 minus.t4 19.8005
R23576 minus.n59 minus.n58 17.9525
R23577 minus.n57 minus.n42 17.9525
R23578 minus.n20 minus.n5 17.9525
R23579 minus.n22 minus.n21 17.9525
R23580 minus.n67 minus.n38 15.9852
R23581 minus.n48 minus.n47 15.9852
R23582 minus.n11 minus.n10 15.9852
R23583 minus.n30 minus.n1 15.9852
R23584 minus.n72 minus.n71 15.3369
R23585 minus.n35 minus.n34 15.3369
R23586 minus.n74 minus.n36 12.1653
R23587 minus minus.n79 11.5562
R23588 minus.n70 minus.n38 8.60764
R23589 minus.n33 minus.n1 8.60764
R23590 minus.n60 minus.n59 6.6403
R23591 minus.n54 minus.n42 6.6403
R23592 minus.n17 minus.n5 6.6403
R23593 minus.n23 minus.n22 6.6403
R23594 minus.n79 minus.n78 4.80222
R23595 minus.n65 minus.n64 4.67295
R23596 minus.n52 minus.n44 4.67295
R23597 minus.n15 minus.n7 4.67295
R23598 minus.n28 minus.n27 4.67295
R23599 minus.n79 minus.n74 0.972091
R23600 minus.n78 minus.n77 0.716017
R23601 minus.n73 minus.n37 0.189894
R23602 minus.n69 minus.n37 0.189894
R23603 minus.n69 minus.n68 0.189894
R23604 minus.n68 minus.n39 0.189894
R23605 minus.n63 minus.n39 0.189894
R23606 minus.n63 minus.n62 0.189894
R23607 minus.n62 minus.n61 0.189894
R23608 minus.n61 minus.n41 0.189894
R23609 minus.n56 minus.n41 0.189894
R23610 minus.n56 minus.n55 0.189894
R23611 minus.n55 minus.n43 0.189894
R23612 minus.n51 minus.n43 0.189894
R23613 minus.n51 minus.n50 0.189894
R23614 minus.n50 minus.n45 0.189894
R23615 minus.n13 minus.n8 0.189894
R23616 minus.n14 minus.n13 0.189894
R23617 minus.n14 minus.n6 0.189894
R23618 minus.n18 minus.n6 0.189894
R23619 minus.n19 minus.n18 0.189894
R23620 minus.n19 minus.n4 0.189894
R23621 minus.n24 minus.n4 0.189894
R23622 minus.n25 minus.n24 0.189894
R23623 minus.n26 minus.n25 0.189894
R23624 minus.n26 minus.n2 0.189894
R23625 minus.n31 minus.n2 0.189894
R23626 minus.n32 minus.n31 0.189894
R23627 minus.n32 minus.n0 0.189894
R23628 minus.n36 minus.n0 0.189894
R23629 output.n41 output.n15 289.615
R23630 output.n72 output.n46 289.615
R23631 output.n104 output.n78 289.615
R23632 output.n136 output.n110 289.615
R23633 output.n77 output.n45 197.26
R23634 output.n77 output.n76 196.298
R23635 output.n109 output.n108 196.298
R23636 output.n141 output.n140 196.298
R23637 output.n42 output.n41 185
R23638 output.n40 output.n39 185
R23639 output.n19 output.n18 185
R23640 output.n34 output.n33 185
R23641 output.n32 output.n31 185
R23642 output.n23 output.n22 185
R23643 output.n26 output.n25 185
R23644 output.n73 output.n72 185
R23645 output.n71 output.n70 185
R23646 output.n50 output.n49 185
R23647 output.n65 output.n64 185
R23648 output.n63 output.n62 185
R23649 output.n54 output.n53 185
R23650 output.n57 output.n56 185
R23651 output.n105 output.n104 185
R23652 output.n103 output.n102 185
R23653 output.n82 output.n81 185
R23654 output.n97 output.n96 185
R23655 output.n95 output.n94 185
R23656 output.n86 output.n85 185
R23657 output.n89 output.n88 185
R23658 output.n137 output.n136 185
R23659 output.n135 output.n134 185
R23660 output.n114 output.n113 185
R23661 output.n129 output.n128 185
R23662 output.n127 output.n126 185
R23663 output.n118 output.n117 185
R23664 output.n121 output.n120 185
R23665 output.t17 output.n24 147.661
R23666 output.t18 output.n55 147.661
R23667 output.t0 output.n87 147.661
R23668 output.t19 output.n119 147.661
R23669 output.n41 output.n40 104.615
R23670 output.n40 output.n18 104.615
R23671 output.n33 output.n18 104.615
R23672 output.n33 output.n32 104.615
R23673 output.n32 output.n22 104.615
R23674 output.n25 output.n22 104.615
R23675 output.n72 output.n71 104.615
R23676 output.n71 output.n49 104.615
R23677 output.n64 output.n49 104.615
R23678 output.n64 output.n63 104.615
R23679 output.n63 output.n53 104.615
R23680 output.n56 output.n53 104.615
R23681 output.n104 output.n103 104.615
R23682 output.n103 output.n81 104.615
R23683 output.n96 output.n81 104.615
R23684 output.n96 output.n95 104.615
R23685 output.n95 output.n85 104.615
R23686 output.n88 output.n85 104.615
R23687 output.n136 output.n135 104.615
R23688 output.n135 output.n113 104.615
R23689 output.n128 output.n113 104.615
R23690 output.n128 output.n127 104.615
R23691 output.n127 output.n117 104.615
R23692 output.n120 output.n117 104.615
R23693 output.n1 output.t2 77.056
R23694 output.n14 output.t4 76.6694
R23695 output.n1 output.n0 72.7095
R23696 output.n3 output.n2 72.7095
R23697 output.n5 output.n4 72.7095
R23698 output.n7 output.n6 72.7095
R23699 output.n9 output.n8 72.7095
R23700 output.n11 output.n10 72.7095
R23701 output.n13 output.n12 72.7095
R23702 output.n25 output.t17 52.3082
R23703 output.n56 output.t18 52.3082
R23704 output.n88 output.t0 52.3082
R23705 output.n120 output.t19 52.3082
R23706 output.n26 output.n24 15.6674
R23707 output.n57 output.n55 15.6674
R23708 output.n89 output.n87 15.6674
R23709 output.n121 output.n119 15.6674
R23710 output.n27 output.n23 12.8005
R23711 output.n58 output.n54 12.8005
R23712 output.n90 output.n86 12.8005
R23713 output.n122 output.n118 12.8005
R23714 output.n31 output.n30 12.0247
R23715 output.n62 output.n61 12.0247
R23716 output.n94 output.n93 12.0247
R23717 output.n126 output.n125 12.0247
R23718 output.n34 output.n21 11.249
R23719 output.n65 output.n52 11.249
R23720 output.n97 output.n84 11.249
R23721 output.n129 output.n116 11.249
R23722 output.n35 output.n19 10.4732
R23723 output.n66 output.n50 10.4732
R23724 output.n98 output.n82 10.4732
R23725 output.n130 output.n114 10.4732
R23726 output.n39 output.n38 9.69747
R23727 output.n70 output.n69 9.69747
R23728 output.n102 output.n101 9.69747
R23729 output.n134 output.n133 9.69747
R23730 output.n45 output.n44 9.45567
R23731 output.n76 output.n75 9.45567
R23732 output.n108 output.n107 9.45567
R23733 output.n140 output.n139 9.45567
R23734 output.n44 output.n43 9.3005
R23735 output.n17 output.n16 9.3005
R23736 output.n38 output.n37 9.3005
R23737 output.n36 output.n35 9.3005
R23738 output.n21 output.n20 9.3005
R23739 output.n30 output.n29 9.3005
R23740 output.n28 output.n27 9.3005
R23741 output.n75 output.n74 9.3005
R23742 output.n48 output.n47 9.3005
R23743 output.n69 output.n68 9.3005
R23744 output.n67 output.n66 9.3005
R23745 output.n52 output.n51 9.3005
R23746 output.n61 output.n60 9.3005
R23747 output.n59 output.n58 9.3005
R23748 output.n107 output.n106 9.3005
R23749 output.n80 output.n79 9.3005
R23750 output.n101 output.n100 9.3005
R23751 output.n99 output.n98 9.3005
R23752 output.n84 output.n83 9.3005
R23753 output.n93 output.n92 9.3005
R23754 output.n91 output.n90 9.3005
R23755 output.n139 output.n138 9.3005
R23756 output.n112 output.n111 9.3005
R23757 output.n133 output.n132 9.3005
R23758 output.n131 output.n130 9.3005
R23759 output.n116 output.n115 9.3005
R23760 output.n125 output.n124 9.3005
R23761 output.n123 output.n122 9.3005
R23762 output.n42 output.n17 8.92171
R23763 output.n73 output.n48 8.92171
R23764 output.n105 output.n80 8.92171
R23765 output.n137 output.n112 8.92171
R23766 output output.n141 8.15037
R23767 output.n43 output.n15 8.14595
R23768 output.n74 output.n46 8.14595
R23769 output.n106 output.n78 8.14595
R23770 output.n138 output.n110 8.14595
R23771 output.n45 output.n15 5.81868
R23772 output.n76 output.n46 5.81868
R23773 output.n108 output.n78 5.81868
R23774 output.n140 output.n110 5.81868
R23775 output.n43 output.n42 5.04292
R23776 output.n74 output.n73 5.04292
R23777 output.n106 output.n105 5.04292
R23778 output.n138 output.n137 5.04292
R23779 output.n28 output.n24 4.38594
R23780 output.n59 output.n55 4.38594
R23781 output.n91 output.n87 4.38594
R23782 output.n123 output.n119 4.38594
R23783 output.n39 output.n17 4.26717
R23784 output.n70 output.n48 4.26717
R23785 output.n102 output.n80 4.26717
R23786 output.n134 output.n112 4.26717
R23787 output.n0 output.t8 3.9605
R23788 output.n0 output.t13 3.9605
R23789 output.n2 output.t1 3.9605
R23790 output.n2 output.t9 3.9605
R23791 output.n4 output.t11 3.9605
R23792 output.n4 output.t10 3.9605
R23793 output.n6 output.t16 3.9605
R23794 output.n6 output.t3 3.9605
R23795 output.n8 output.t5 3.9605
R23796 output.n8 output.t14 3.9605
R23797 output.n10 output.t15 3.9605
R23798 output.n10 output.t6 3.9605
R23799 output.n12 output.t7 3.9605
R23800 output.n12 output.t12 3.9605
R23801 output.n38 output.n19 3.49141
R23802 output.n69 output.n50 3.49141
R23803 output.n101 output.n82 3.49141
R23804 output.n133 output.n114 3.49141
R23805 output.n35 output.n34 2.71565
R23806 output.n66 output.n65 2.71565
R23807 output.n98 output.n97 2.71565
R23808 output.n130 output.n129 2.71565
R23809 output.n31 output.n21 1.93989
R23810 output.n62 output.n52 1.93989
R23811 output.n94 output.n84 1.93989
R23812 output.n126 output.n116 1.93989
R23813 output.n30 output.n23 1.16414
R23814 output.n61 output.n54 1.16414
R23815 output.n93 output.n86 1.16414
R23816 output.n125 output.n118 1.16414
R23817 output.n141 output.n109 0.962709
R23818 output.n109 output.n77 0.962709
R23819 output.n27 output.n26 0.388379
R23820 output.n58 output.n57 0.388379
R23821 output.n90 output.n89 0.388379
R23822 output.n122 output.n121 0.388379
R23823 output.n14 output.n13 0.387128
R23824 output.n13 output.n11 0.387128
R23825 output.n11 output.n9 0.387128
R23826 output.n9 output.n7 0.387128
R23827 output.n7 output.n5 0.387128
R23828 output.n5 output.n3 0.387128
R23829 output.n3 output.n1 0.387128
R23830 output.n44 output.n16 0.155672
R23831 output.n37 output.n16 0.155672
R23832 output.n37 output.n36 0.155672
R23833 output.n36 output.n20 0.155672
R23834 output.n29 output.n20 0.155672
R23835 output.n29 output.n28 0.155672
R23836 output.n75 output.n47 0.155672
R23837 output.n68 output.n47 0.155672
R23838 output.n68 output.n67 0.155672
R23839 output.n67 output.n51 0.155672
R23840 output.n60 output.n51 0.155672
R23841 output.n60 output.n59 0.155672
R23842 output.n107 output.n79 0.155672
R23843 output.n100 output.n79 0.155672
R23844 output.n100 output.n99 0.155672
R23845 output.n99 output.n83 0.155672
R23846 output.n92 output.n83 0.155672
R23847 output.n92 output.n91 0.155672
R23848 output.n139 output.n111 0.155672
R23849 output.n132 output.n111 0.155672
R23850 output.n132 output.n131 0.155672
R23851 output.n131 output.n115 0.155672
R23852 output.n124 output.n115 0.155672
R23853 output.n124 output.n123 0.155672
R23854 output output.n14 0.126227
R23855 diffpairibias.n0 diffpairibias.t18 436.822
R23856 diffpairibias.n21 diffpairibias.t19 435.479
R23857 diffpairibias.n20 diffpairibias.t16 435.479
R23858 diffpairibias.n19 diffpairibias.t17 435.479
R23859 diffpairibias.n18 diffpairibias.t21 435.479
R23860 diffpairibias.n0 diffpairibias.t22 435.479
R23861 diffpairibias.n1 diffpairibias.t20 435.479
R23862 diffpairibias.n2 diffpairibias.t23 435.479
R23863 diffpairibias.n10 diffpairibias.t0 377.536
R23864 diffpairibias.n10 diffpairibias.t8 376.193
R23865 diffpairibias.n11 diffpairibias.t10 376.193
R23866 diffpairibias.n12 diffpairibias.t6 376.193
R23867 diffpairibias.n13 diffpairibias.t2 376.193
R23868 diffpairibias.n14 diffpairibias.t12 376.193
R23869 diffpairibias.n15 diffpairibias.t4 376.193
R23870 diffpairibias.n16 diffpairibias.t14 376.193
R23871 diffpairibias.n3 diffpairibias.t1 113.368
R23872 diffpairibias.n3 diffpairibias.t9 112.698
R23873 diffpairibias.n4 diffpairibias.t11 112.698
R23874 diffpairibias.n5 diffpairibias.t7 112.698
R23875 diffpairibias.n6 diffpairibias.t3 112.698
R23876 diffpairibias.n7 diffpairibias.t13 112.698
R23877 diffpairibias.n8 diffpairibias.t5 112.698
R23878 diffpairibias.n9 diffpairibias.t15 112.698
R23879 diffpairibias.n17 diffpairibias.n16 4.77242
R23880 diffpairibias.n17 diffpairibias.n9 4.30807
R23881 diffpairibias.n18 diffpairibias.n17 4.13945
R23882 diffpairibias.n16 diffpairibias.n15 1.34352
R23883 diffpairibias.n15 diffpairibias.n14 1.34352
R23884 diffpairibias.n14 diffpairibias.n13 1.34352
R23885 diffpairibias.n13 diffpairibias.n12 1.34352
R23886 diffpairibias.n12 diffpairibias.n11 1.34352
R23887 diffpairibias.n11 diffpairibias.n10 1.34352
R23888 diffpairibias.n2 diffpairibias.n1 1.34352
R23889 diffpairibias.n1 diffpairibias.n0 1.34352
R23890 diffpairibias.n19 diffpairibias.n18 1.34352
R23891 diffpairibias.n20 diffpairibias.n19 1.34352
R23892 diffpairibias.n21 diffpairibias.n20 1.34352
R23893 diffpairibias.n22 diffpairibias.n21 0.862419
R23894 diffpairibias diffpairibias.n22 0.684875
R23895 diffpairibias.n9 diffpairibias.n8 0.672012
R23896 diffpairibias.n8 diffpairibias.n7 0.672012
R23897 diffpairibias.n7 diffpairibias.n6 0.672012
R23898 diffpairibias.n6 diffpairibias.n5 0.672012
R23899 diffpairibias.n5 diffpairibias.n4 0.672012
R23900 diffpairibias.n4 diffpairibias.n3 0.672012
R23901 diffpairibias.n22 diffpairibias.n2 0.190907
R23902 outputibias.n27 outputibias.n1 289.615
R23903 outputibias.n58 outputibias.n32 289.615
R23904 outputibias.n90 outputibias.n64 289.615
R23905 outputibias.n122 outputibias.n96 289.615
R23906 outputibias.n28 outputibias.n27 185
R23907 outputibias.n26 outputibias.n25 185
R23908 outputibias.n5 outputibias.n4 185
R23909 outputibias.n20 outputibias.n19 185
R23910 outputibias.n18 outputibias.n17 185
R23911 outputibias.n9 outputibias.n8 185
R23912 outputibias.n12 outputibias.n11 185
R23913 outputibias.n59 outputibias.n58 185
R23914 outputibias.n57 outputibias.n56 185
R23915 outputibias.n36 outputibias.n35 185
R23916 outputibias.n51 outputibias.n50 185
R23917 outputibias.n49 outputibias.n48 185
R23918 outputibias.n40 outputibias.n39 185
R23919 outputibias.n43 outputibias.n42 185
R23920 outputibias.n91 outputibias.n90 185
R23921 outputibias.n89 outputibias.n88 185
R23922 outputibias.n68 outputibias.n67 185
R23923 outputibias.n83 outputibias.n82 185
R23924 outputibias.n81 outputibias.n80 185
R23925 outputibias.n72 outputibias.n71 185
R23926 outputibias.n75 outputibias.n74 185
R23927 outputibias.n123 outputibias.n122 185
R23928 outputibias.n121 outputibias.n120 185
R23929 outputibias.n100 outputibias.n99 185
R23930 outputibias.n115 outputibias.n114 185
R23931 outputibias.n113 outputibias.n112 185
R23932 outputibias.n104 outputibias.n103 185
R23933 outputibias.n107 outputibias.n106 185
R23934 outputibias.n0 outputibias.t10 178.945
R23935 outputibias.n133 outputibias.t8 177.018
R23936 outputibias.n132 outputibias.t11 177.018
R23937 outputibias.n0 outputibias.t9 177.018
R23938 outputibias.t7 outputibias.n10 147.661
R23939 outputibias.t1 outputibias.n41 147.661
R23940 outputibias.t3 outputibias.n73 147.661
R23941 outputibias.t5 outputibias.n105 147.661
R23942 outputibias.n128 outputibias.t6 132.363
R23943 outputibias.n128 outputibias.t0 130.436
R23944 outputibias.n129 outputibias.t2 130.436
R23945 outputibias.n130 outputibias.t4 130.436
R23946 outputibias.n27 outputibias.n26 104.615
R23947 outputibias.n26 outputibias.n4 104.615
R23948 outputibias.n19 outputibias.n4 104.615
R23949 outputibias.n19 outputibias.n18 104.615
R23950 outputibias.n18 outputibias.n8 104.615
R23951 outputibias.n11 outputibias.n8 104.615
R23952 outputibias.n58 outputibias.n57 104.615
R23953 outputibias.n57 outputibias.n35 104.615
R23954 outputibias.n50 outputibias.n35 104.615
R23955 outputibias.n50 outputibias.n49 104.615
R23956 outputibias.n49 outputibias.n39 104.615
R23957 outputibias.n42 outputibias.n39 104.615
R23958 outputibias.n90 outputibias.n89 104.615
R23959 outputibias.n89 outputibias.n67 104.615
R23960 outputibias.n82 outputibias.n67 104.615
R23961 outputibias.n82 outputibias.n81 104.615
R23962 outputibias.n81 outputibias.n71 104.615
R23963 outputibias.n74 outputibias.n71 104.615
R23964 outputibias.n122 outputibias.n121 104.615
R23965 outputibias.n121 outputibias.n99 104.615
R23966 outputibias.n114 outputibias.n99 104.615
R23967 outputibias.n114 outputibias.n113 104.615
R23968 outputibias.n113 outputibias.n103 104.615
R23969 outputibias.n106 outputibias.n103 104.615
R23970 outputibias.n63 outputibias.n31 95.6354
R23971 outputibias.n63 outputibias.n62 94.6732
R23972 outputibias.n95 outputibias.n94 94.6732
R23973 outputibias.n127 outputibias.n126 94.6732
R23974 outputibias.n11 outputibias.t7 52.3082
R23975 outputibias.n42 outputibias.t1 52.3082
R23976 outputibias.n74 outputibias.t3 52.3082
R23977 outputibias.n106 outputibias.t5 52.3082
R23978 outputibias.n12 outputibias.n10 15.6674
R23979 outputibias.n43 outputibias.n41 15.6674
R23980 outputibias.n75 outputibias.n73 15.6674
R23981 outputibias.n107 outputibias.n105 15.6674
R23982 outputibias.n13 outputibias.n9 12.8005
R23983 outputibias.n44 outputibias.n40 12.8005
R23984 outputibias.n76 outputibias.n72 12.8005
R23985 outputibias.n108 outputibias.n104 12.8005
R23986 outputibias.n17 outputibias.n16 12.0247
R23987 outputibias.n48 outputibias.n47 12.0247
R23988 outputibias.n80 outputibias.n79 12.0247
R23989 outputibias.n112 outputibias.n111 12.0247
R23990 outputibias.n20 outputibias.n7 11.249
R23991 outputibias.n51 outputibias.n38 11.249
R23992 outputibias.n83 outputibias.n70 11.249
R23993 outputibias.n115 outputibias.n102 11.249
R23994 outputibias.n21 outputibias.n5 10.4732
R23995 outputibias.n52 outputibias.n36 10.4732
R23996 outputibias.n84 outputibias.n68 10.4732
R23997 outputibias.n116 outputibias.n100 10.4732
R23998 outputibias.n25 outputibias.n24 9.69747
R23999 outputibias.n56 outputibias.n55 9.69747
R24000 outputibias.n88 outputibias.n87 9.69747
R24001 outputibias.n120 outputibias.n119 9.69747
R24002 outputibias.n31 outputibias.n30 9.45567
R24003 outputibias.n62 outputibias.n61 9.45567
R24004 outputibias.n94 outputibias.n93 9.45567
R24005 outputibias.n126 outputibias.n125 9.45567
R24006 outputibias.n30 outputibias.n29 9.3005
R24007 outputibias.n3 outputibias.n2 9.3005
R24008 outputibias.n24 outputibias.n23 9.3005
R24009 outputibias.n22 outputibias.n21 9.3005
R24010 outputibias.n7 outputibias.n6 9.3005
R24011 outputibias.n16 outputibias.n15 9.3005
R24012 outputibias.n14 outputibias.n13 9.3005
R24013 outputibias.n61 outputibias.n60 9.3005
R24014 outputibias.n34 outputibias.n33 9.3005
R24015 outputibias.n55 outputibias.n54 9.3005
R24016 outputibias.n53 outputibias.n52 9.3005
R24017 outputibias.n38 outputibias.n37 9.3005
R24018 outputibias.n47 outputibias.n46 9.3005
R24019 outputibias.n45 outputibias.n44 9.3005
R24020 outputibias.n93 outputibias.n92 9.3005
R24021 outputibias.n66 outputibias.n65 9.3005
R24022 outputibias.n87 outputibias.n86 9.3005
R24023 outputibias.n85 outputibias.n84 9.3005
R24024 outputibias.n70 outputibias.n69 9.3005
R24025 outputibias.n79 outputibias.n78 9.3005
R24026 outputibias.n77 outputibias.n76 9.3005
R24027 outputibias.n125 outputibias.n124 9.3005
R24028 outputibias.n98 outputibias.n97 9.3005
R24029 outputibias.n119 outputibias.n118 9.3005
R24030 outputibias.n117 outputibias.n116 9.3005
R24031 outputibias.n102 outputibias.n101 9.3005
R24032 outputibias.n111 outputibias.n110 9.3005
R24033 outputibias.n109 outputibias.n108 9.3005
R24034 outputibias.n28 outputibias.n3 8.92171
R24035 outputibias.n59 outputibias.n34 8.92171
R24036 outputibias.n91 outputibias.n66 8.92171
R24037 outputibias.n123 outputibias.n98 8.92171
R24038 outputibias.n29 outputibias.n1 8.14595
R24039 outputibias.n60 outputibias.n32 8.14595
R24040 outputibias.n92 outputibias.n64 8.14595
R24041 outputibias.n124 outputibias.n96 8.14595
R24042 outputibias.n31 outputibias.n1 5.81868
R24043 outputibias.n62 outputibias.n32 5.81868
R24044 outputibias.n94 outputibias.n64 5.81868
R24045 outputibias.n126 outputibias.n96 5.81868
R24046 outputibias.n131 outputibias.n130 5.20947
R24047 outputibias.n29 outputibias.n28 5.04292
R24048 outputibias.n60 outputibias.n59 5.04292
R24049 outputibias.n92 outputibias.n91 5.04292
R24050 outputibias.n124 outputibias.n123 5.04292
R24051 outputibias.n131 outputibias.n127 4.42209
R24052 outputibias.n14 outputibias.n10 4.38594
R24053 outputibias.n45 outputibias.n41 4.38594
R24054 outputibias.n77 outputibias.n73 4.38594
R24055 outputibias.n109 outputibias.n105 4.38594
R24056 outputibias.n132 outputibias.n131 4.28454
R24057 outputibias.n25 outputibias.n3 4.26717
R24058 outputibias.n56 outputibias.n34 4.26717
R24059 outputibias.n88 outputibias.n66 4.26717
R24060 outputibias.n120 outputibias.n98 4.26717
R24061 outputibias.n24 outputibias.n5 3.49141
R24062 outputibias.n55 outputibias.n36 3.49141
R24063 outputibias.n87 outputibias.n68 3.49141
R24064 outputibias.n119 outputibias.n100 3.49141
R24065 outputibias.n21 outputibias.n20 2.71565
R24066 outputibias.n52 outputibias.n51 2.71565
R24067 outputibias.n84 outputibias.n83 2.71565
R24068 outputibias.n116 outputibias.n115 2.71565
R24069 outputibias.n17 outputibias.n7 1.93989
R24070 outputibias.n48 outputibias.n38 1.93989
R24071 outputibias.n80 outputibias.n70 1.93989
R24072 outputibias.n112 outputibias.n102 1.93989
R24073 outputibias.n130 outputibias.n129 1.9266
R24074 outputibias.n129 outputibias.n128 1.9266
R24075 outputibias.n133 outputibias.n132 1.92658
R24076 outputibias.n134 outputibias.n133 1.29913
R24077 outputibias.n16 outputibias.n9 1.16414
R24078 outputibias.n47 outputibias.n40 1.16414
R24079 outputibias.n79 outputibias.n72 1.16414
R24080 outputibias.n111 outputibias.n104 1.16414
R24081 outputibias.n127 outputibias.n95 0.962709
R24082 outputibias.n95 outputibias.n63 0.962709
R24083 outputibias.n13 outputibias.n12 0.388379
R24084 outputibias.n44 outputibias.n43 0.388379
R24085 outputibias.n76 outputibias.n75 0.388379
R24086 outputibias.n108 outputibias.n107 0.388379
R24087 outputibias.n134 outputibias.n0 0.337251
R24088 outputibias outputibias.n134 0.302375
R24089 outputibias.n30 outputibias.n2 0.155672
R24090 outputibias.n23 outputibias.n2 0.155672
R24091 outputibias.n23 outputibias.n22 0.155672
R24092 outputibias.n22 outputibias.n6 0.155672
R24093 outputibias.n15 outputibias.n6 0.155672
R24094 outputibias.n15 outputibias.n14 0.155672
R24095 outputibias.n61 outputibias.n33 0.155672
R24096 outputibias.n54 outputibias.n33 0.155672
R24097 outputibias.n54 outputibias.n53 0.155672
R24098 outputibias.n53 outputibias.n37 0.155672
R24099 outputibias.n46 outputibias.n37 0.155672
R24100 outputibias.n46 outputibias.n45 0.155672
R24101 outputibias.n93 outputibias.n65 0.155672
R24102 outputibias.n86 outputibias.n65 0.155672
R24103 outputibias.n86 outputibias.n85 0.155672
R24104 outputibias.n85 outputibias.n69 0.155672
R24105 outputibias.n78 outputibias.n69 0.155672
R24106 outputibias.n78 outputibias.n77 0.155672
R24107 outputibias.n125 outputibias.n97 0.155672
R24108 outputibias.n118 outputibias.n97 0.155672
R24109 outputibias.n118 outputibias.n117 0.155672
R24110 outputibias.n117 outputibias.n101 0.155672
R24111 outputibias.n110 outputibias.n101 0.155672
R24112 outputibias.n110 outputibias.n109 0.155672
C0 output outputibias 2.34152f
C1 vdd output 7.23429f
C2 CSoutput output 6.13881f
C3 CSoutput outputibias 0.032386f
C4 vdd CSoutput 0.14092p
C5 commonsourceibias output 0.006808f
C6 minus diffpairibias 3.46e-19
C7 CSoutput minus 2.77524f
C8 vdd plus 0.092938f
C9 plus diffpairibias 2.47e-19
C10 commonsourceibias outputibias 0.003832f
C11 vdd commonsourceibias 0.004218f
C12 CSoutput plus 0.856907f
C13 commonsourceibias diffpairibias 0.06482f
C14 CSoutput commonsourceibias 54.0646f
C15 minus plus 9.171639f
C16 minus commonsourceibias 0.323289f
C17 plus commonsourceibias 0.277692f
C18 diffpairibias gnd 48.980137f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.183542p
C22 plus gnd 32.70674f
C23 minus gnd 26.99455f
C24 CSoutput gnd 0.124832p
C25 vdd gnd 0.473154p
C26 outputibias.t9 gnd 0.11477f
C27 outputibias.t10 gnd 0.115567f
C28 outputibias.n0 gnd 0.130108f
C29 outputibias.n1 gnd 0.001372f
C30 outputibias.n2 gnd 9.76e-19
C31 outputibias.n3 gnd 5.24e-19
C32 outputibias.n4 gnd 0.001239f
C33 outputibias.n5 gnd 5.55e-19
C34 outputibias.n6 gnd 9.76e-19
C35 outputibias.n7 gnd 5.24e-19
C36 outputibias.n8 gnd 0.001239f
C37 outputibias.n9 gnd 5.55e-19
C38 outputibias.n10 gnd 0.004176f
C39 outputibias.t7 gnd 0.00202f
C40 outputibias.n11 gnd 9.3e-19
C41 outputibias.n12 gnd 7.32e-19
C42 outputibias.n13 gnd 5.24e-19
C43 outputibias.n14 gnd 0.02322f
C44 outputibias.n15 gnd 9.76e-19
C45 outputibias.n16 gnd 5.24e-19
C46 outputibias.n17 gnd 5.55e-19
C47 outputibias.n18 gnd 0.001239f
C48 outputibias.n19 gnd 0.001239f
C49 outputibias.n20 gnd 5.55e-19
C50 outputibias.n21 gnd 5.24e-19
C51 outputibias.n22 gnd 9.76e-19
C52 outputibias.n23 gnd 9.76e-19
C53 outputibias.n24 gnd 5.24e-19
C54 outputibias.n25 gnd 5.55e-19
C55 outputibias.n26 gnd 0.001239f
C56 outputibias.n27 gnd 0.002683f
C57 outputibias.n28 gnd 5.55e-19
C58 outputibias.n29 gnd 5.24e-19
C59 outputibias.n30 gnd 0.002256f
C60 outputibias.n31 gnd 0.005781f
C61 outputibias.n32 gnd 0.001372f
C62 outputibias.n33 gnd 9.76e-19
C63 outputibias.n34 gnd 5.24e-19
C64 outputibias.n35 gnd 0.001239f
C65 outputibias.n36 gnd 5.55e-19
C66 outputibias.n37 gnd 9.76e-19
C67 outputibias.n38 gnd 5.24e-19
C68 outputibias.n39 gnd 0.001239f
C69 outputibias.n40 gnd 5.55e-19
C70 outputibias.n41 gnd 0.004176f
C71 outputibias.t1 gnd 0.00202f
C72 outputibias.n42 gnd 9.3e-19
C73 outputibias.n43 gnd 7.32e-19
C74 outputibias.n44 gnd 5.24e-19
C75 outputibias.n45 gnd 0.02322f
C76 outputibias.n46 gnd 9.76e-19
C77 outputibias.n47 gnd 5.24e-19
C78 outputibias.n48 gnd 5.55e-19
C79 outputibias.n49 gnd 0.001239f
C80 outputibias.n50 gnd 0.001239f
C81 outputibias.n51 gnd 5.55e-19
C82 outputibias.n52 gnd 5.24e-19
C83 outputibias.n53 gnd 9.76e-19
C84 outputibias.n54 gnd 9.76e-19
C85 outputibias.n55 gnd 5.24e-19
C86 outputibias.n56 gnd 5.55e-19
C87 outputibias.n57 gnd 0.001239f
C88 outputibias.n58 gnd 0.002683f
C89 outputibias.n59 gnd 5.55e-19
C90 outputibias.n60 gnd 5.24e-19
C91 outputibias.n61 gnd 0.002256f
C92 outputibias.n62 gnd 0.005197f
C93 outputibias.n63 gnd 0.121892f
C94 outputibias.n64 gnd 0.001372f
C95 outputibias.n65 gnd 9.76e-19
C96 outputibias.n66 gnd 5.24e-19
C97 outputibias.n67 gnd 0.001239f
C98 outputibias.n68 gnd 5.55e-19
C99 outputibias.n69 gnd 9.76e-19
C100 outputibias.n70 gnd 5.24e-19
C101 outputibias.n71 gnd 0.001239f
C102 outputibias.n72 gnd 5.55e-19
C103 outputibias.n73 gnd 0.004176f
C104 outputibias.t3 gnd 0.00202f
C105 outputibias.n74 gnd 9.3e-19
C106 outputibias.n75 gnd 7.32e-19
C107 outputibias.n76 gnd 5.24e-19
C108 outputibias.n77 gnd 0.02322f
C109 outputibias.n78 gnd 9.76e-19
C110 outputibias.n79 gnd 5.24e-19
C111 outputibias.n80 gnd 5.55e-19
C112 outputibias.n81 gnd 0.001239f
C113 outputibias.n82 gnd 0.001239f
C114 outputibias.n83 gnd 5.55e-19
C115 outputibias.n84 gnd 5.24e-19
C116 outputibias.n85 gnd 9.76e-19
C117 outputibias.n86 gnd 9.76e-19
C118 outputibias.n87 gnd 5.24e-19
C119 outputibias.n88 gnd 5.55e-19
C120 outputibias.n89 gnd 0.001239f
C121 outputibias.n90 gnd 0.002683f
C122 outputibias.n91 gnd 5.55e-19
C123 outputibias.n92 gnd 5.24e-19
C124 outputibias.n93 gnd 0.002256f
C125 outputibias.n94 gnd 0.005197f
C126 outputibias.n95 gnd 0.064513f
C127 outputibias.n96 gnd 0.001372f
C128 outputibias.n97 gnd 9.76e-19
C129 outputibias.n98 gnd 5.24e-19
C130 outputibias.n99 gnd 0.001239f
C131 outputibias.n100 gnd 5.55e-19
C132 outputibias.n101 gnd 9.76e-19
C133 outputibias.n102 gnd 5.24e-19
C134 outputibias.n103 gnd 0.001239f
C135 outputibias.n104 gnd 5.55e-19
C136 outputibias.n105 gnd 0.004176f
C137 outputibias.t5 gnd 0.00202f
C138 outputibias.n106 gnd 9.3e-19
C139 outputibias.n107 gnd 7.32e-19
C140 outputibias.n108 gnd 5.24e-19
C141 outputibias.n109 gnd 0.02322f
C142 outputibias.n110 gnd 9.76e-19
C143 outputibias.n111 gnd 5.24e-19
C144 outputibias.n112 gnd 5.55e-19
C145 outputibias.n113 gnd 0.001239f
C146 outputibias.n114 gnd 0.001239f
C147 outputibias.n115 gnd 5.55e-19
C148 outputibias.n116 gnd 5.24e-19
C149 outputibias.n117 gnd 9.76e-19
C150 outputibias.n118 gnd 9.76e-19
C151 outputibias.n119 gnd 5.24e-19
C152 outputibias.n120 gnd 5.55e-19
C153 outputibias.n121 gnd 0.001239f
C154 outputibias.n122 gnd 0.002683f
C155 outputibias.n123 gnd 5.55e-19
C156 outputibias.n124 gnd 5.24e-19
C157 outputibias.n125 gnd 0.002256f
C158 outputibias.n126 gnd 0.005197f
C159 outputibias.n127 gnd 0.084814f
C160 outputibias.t4 gnd 0.108319f
C161 outputibias.t2 gnd 0.108319f
C162 outputibias.t0 gnd 0.108319f
C163 outputibias.t6 gnd 0.109238f
C164 outputibias.n128 gnd 0.134674f
C165 outputibias.n129 gnd 0.07244f
C166 outputibias.n130 gnd 0.079818f
C167 outputibias.n131 gnd 0.164901f
C168 outputibias.t11 gnd 0.11477f
C169 outputibias.n132 gnd 0.067481f
C170 outputibias.t8 gnd 0.11477f
C171 outputibias.n133 gnd 0.065115f
C172 outputibias.n134 gnd 0.029159f
C173 diffpairibias.t18 gnd 0.087401f
C174 diffpairibias.t22 gnd 0.087239f
C175 diffpairibias.n0 gnd 0.102784f
C176 diffpairibias.t20 gnd 0.087239f
C177 diffpairibias.n1 gnd 0.050171f
C178 diffpairibias.t23 gnd 0.087239f
C179 diffpairibias.n2 gnd 0.039841f
C180 diffpairibias.t1 gnd 0.083757f
C181 diffpairibias.t9 gnd 0.083392f
C182 diffpairibias.n3 gnd 0.131682f
C183 diffpairibias.t11 gnd 0.083392f
C184 diffpairibias.n4 gnd 0.07027f
C185 diffpairibias.t7 gnd 0.083392f
C186 diffpairibias.n5 gnd 0.07027f
C187 diffpairibias.t3 gnd 0.083392f
C188 diffpairibias.n6 gnd 0.07027f
C189 diffpairibias.t13 gnd 0.083392f
C190 diffpairibias.n7 gnd 0.07027f
C191 diffpairibias.t5 gnd 0.083392f
C192 diffpairibias.n8 gnd 0.07027f
C193 diffpairibias.t15 gnd 0.083392f
C194 diffpairibias.n9 gnd 0.099771f
C195 diffpairibias.t0 gnd 0.08427f
C196 diffpairibias.t8 gnd 0.084123f
C197 diffpairibias.n10 gnd 0.091784f
C198 diffpairibias.t10 gnd 0.084123f
C199 diffpairibias.n11 gnd 0.050681f
C200 diffpairibias.t6 gnd 0.084123f
C201 diffpairibias.n12 gnd 0.050681f
C202 diffpairibias.t2 gnd 0.084123f
C203 diffpairibias.n13 gnd 0.050681f
C204 diffpairibias.t12 gnd 0.084123f
C205 diffpairibias.n14 gnd 0.050681f
C206 diffpairibias.t4 gnd 0.084123f
C207 diffpairibias.n15 gnd 0.050681f
C208 diffpairibias.t14 gnd 0.084123f
C209 diffpairibias.n16 gnd 0.059977f
C210 diffpairibias.n17 gnd 0.226448f
C211 diffpairibias.t21 gnd 0.087239f
C212 diffpairibias.n18 gnd 0.050181f
C213 diffpairibias.t17 gnd 0.087239f
C214 diffpairibias.n19 gnd 0.050171f
C215 diffpairibias.t16 gnd 0.087239f
C216 diffpairibias.n20 gnd 0.050171f
C217 diffpairibias.t19 gnd 0.087239f
C218 diffpairibias.n21 gnd 0.045859f
C219 diffpairibias.n22 gnd 0.046268f
C220 output.t2 gnd 0.464308f
C221 output.t8 gnd 0.044422f
C222 output.t13 gnd 0.044422f
C223 output.n0 gnd 0.364624f
C224 output.n1 gnd 0.614102f
C225 output.t1 gnd 0.044422f
C226 output.t9 gnd 0.044422f
C227 output.n2 gnd 0.364624f
C228 output.n3 gnd 0.350265f
C229 output.t11 gnd 0.044422f
C230 output.t10 gnd 0.044422f
C231 output.n4 gnd 0.364624f
C232 output.n5 gnd 0.350265f
C233 output.t16 gnd 0.044422f
C234 output.t3 gnd 0.044422f
C235 output.n6 gnd 0.364624f
C236 output.n7 gnd 0.350265f
C237 output.t5 gnd 0.044422f
C238 output.t14 gnd 0.044422f
C239 output.n8 gnd 0.364624f
C240 output.n9 gnd 0.350265f
C241 output.t15 gnd 0.044422f
C242 output.t6 gnd 0.044422f
C243 output.n10 gnd 0.364624f
C244 output.n11 gnd 0.350265f
C245 output.t7 gnd 0.044422f
C246 output.t12 gnd 0.044422f
C247 output.n12 gnd 0.364624f
C248 output.n13 gnd 0.350265f
C249 output.t4 gnd 0.462979f
C250 output.n14 gnd 0.28994f
C251 output.n15 gnd 0.015803f
C252 output.n16 gnd 0.011243f
C253 output.n17 gnd 0.006041f
C254 output.n18 gnd 0.01428f
C255 output.n19 gnd 0.006397f
C256 output.n20 gnd 0.011243f
C257 output.n21 gnd 0.006041f
C258 output.n22 gnd 0.01428f
C259 output.n23 gnd 0.006397f
C260 output.n24 gnd 0.048111f
C261 output.t17 gnd 0.023274f
C262 output.n25 gnd 0.01071f
C263 output.n26 gnd 0.008435f
C264 output.n27 gnd 0.006041f
C265 output.n28 gnd 0.267512f
C266 output.n29 gnd 0.011243f
C267 output.n30 gnd 0.006041f
C268 output.n31 gnd 0.006397f
C269 output.n32 gnd 0.01428f
C270 output.n33 gnd 0.01428f
C271 output.n34 gnd 0.006397f
C272 output.n35 gnd 0.006041f
C273 output.n36 gnd 0.011243f
C274 output.n37 gnd 0.011243f
C275 output.n38 gnd 0.006041f
C276 output.n39 gnd 0.006397f
C277 output.n40 gnd 0.01428f
C278 output.n41 gnd 0.030913f
C279 output.n42 gnd 0.006397f
C280 output.n43 gnd 0.006041f
C281 output.n44 gnd 0.025987f
C282 output.n45 gnd 0.097665f
C283 output.n46 gnd 0.015803f
C284 output.n47 gnd 0.011243f
C285 output.n48 gnd 0.006041f
C286 output.n49 gnd 0.01428f
C287 output.n50 gnd 0.006397f
C288 output.n51 gnd 0.011243f
C289 output.n52 gnd 0.006041f
C290 output.n53 gnd 0.01428f
C291 output.n54 gnd 0.006397f
C292 output.n55 gnd 0.048111f
C293 output.t18 gnd 0.023274f
C294 output.n56 gnd 0.01071f
C295 output.n57 gnd 0.008435f
C296 output.n58 gnd 0.006041f
C297 output.n59 gnd 0.267512f
C298 output.n60 gnd 0.011243f
C299 output.n61 gnd 0.006041f
C300 output.n62 gnd 0.006397f
C301 output.n63 gnd 0.01428f
C302 output.n64 gnd 0.01428f
C303 output.n65 gnd 0.006397f
C304 output.n66 gnd 0.006041f
C305 output.n67 gnd 0.011243f
C306 output.n68 gnd 0.011243f
C307 output.n69 gnd 0.006041f
C308 output.n70 gnd 0.006397f
C309 output.n71 gnd 0.01428f
C310 output.n72 gnd 0.030913f
C311 output.n73 gnd 0.006397f
C312 output.n74 gnd 0.006041f
C313 output.n75 gnd 0.025987f
C314 output.n76 gnd 0.09306f
C315 output.n77 gnd 1.65264f
C316 output.n78 gnd 0.015803f
C317 output.n79 gnd 0.011243f
C318 output.n80 gnd 0.006041f
C319 output.n81 gnd 0.01428f
C320 output.n82 gnd 0.006397f
C321 output.n83 gnd 0.011243f
C322 output.n84 gnd 0.006041f
C323 output.n85 gnd 0.01428f
C324 output.n86 gnd 0.006397f
C325 output.n87 gnd 0.048111f
C326 output.t0 gnd 0.023274f
C327 output.n88 gnd 0.01071f
C328 output.n89 gnd 0.008435f
C329 output.n90 gnd 0.006041f
C330 output.n91 gnd 0.267512f
C331 output.n92 gnd 0.011243f
C332 output.n93 gnd 0.006041f
C333 output.n94 gnd 0.006397f
C334 output.n95 gnd 0.01428f
C335 output.n96 gnd 0.01428f
C336 output.n97 gnd 0.006397f
C337 output.n98 gnd 0.006041f
C338 output.n99 gnd 0.011243f
C339 output.n100 gnd 0.011243f
C340 output.n101 gnd 0.006041f
C341 output.n102 gnd 0.006397f
C342 output.n103 gnd 0.01428f
C343 output.n104 gnd 0.030913f
C344 output.n105 gnd 0.006397f
C345 output.n106 gnd 0.006041f
C346 output.n107 gnd 0.025987f
C347 output.n108 gnd 0.09306f
C348 output.n109 gnd 0.713089f
C349 output.n110 gnd 0.015803f
C350 output.n111 gnd 0.011243f
C351 output.n112 gnd 0.006041f
C352 output.n113 gnd 0.01428f
C353 output.n114 gnd 0.006397f
C354 output.n115 gnd 0.011243f
C355 output.n116 gnd 0.006041f
C356 output.n117 gnd 0.01428f
C357 output.n118 gnd 0.006397f
C358 output.n119 gnd 0.048111f
C359 output.t19 gnd 0.023274f
C360 output.n120 gnd 0.01071f
C361 output.n121 gnd 0.008435f
C362 output.n122 gnd 0.006041f
C363 output.n123 gnd 0.267512f
C364 output.n124 gnd 0.011243f
C365 output.n125 gnd 0.006041f
C366 output.n126 gnd 0.006397f
C367 output.n127 gnd 0.01428f
C368 output.n128 gnd 0.01428f
C369 output.n129 gnd 0.006397f
C370 output.n130 gnd 0.006041f
C371 output.n131 gnd 0.011243f
C372 output.n132 gnd 0.011243f
C373 output.n133 gnd 0.006041f
C374 output.n134 gnd 0.006397f
C375 output.n135 gnd 0.01428f
C376 output.n136 gnd 0.030913f
C377 output.n137 gnd 0.006397f
C378 output.n138 gnd 0.006041f
C379 output.n139 gnd 0.025987f
C380 output.n140 gnd 0.09306f
C381 output.n141 gnd 1.67353f
C382 minus.n0 gnd 0.030059f
C383 minus.t14 gnd 0.505432f
C384 minus.n1 gnd 0.204419f
C385 minus.n2 gnd 0.030059f
C386 minus.t19 gnd 0.505432f
C387 minus.n3 gnd 0.024431f
C388 minus.n4 gnd 0.030059f
C389 minus.t18 gnd 0.505432f
C390 minus.t5 gnd 0.505432f
C391 minus.n5 gnd 0.204419f
C392 minus.n6 gnd 0.030059f
C393 minus.t8 gnd 0.505432f
C394 minus.n7 gnd 0.204419f
C395 minus.n8 gnd 0.12903f
C396 minus.t9 gnd 0.505432f
C397 minus.t13 gnd 0.567467f
C398 minus.n9 gnd 0.237182f
C399 minus.n10 gnd 0.236072f
C400 minus.n11 gnd 0.03739f
C401 minus.n12 gnd 0.03514f
C402 minus.n13 gnd 0.030059f
C403 minus.n14 gnd 0.030059f
C404 minus.n15 gnd 0.037653f
C405 minus.n16 gnd 0.024431f
C406 minus.n17 gnd 0.038669f
C407 minus.n18 gnd 0.030059f
C408 minus.n19 gnd 0.030059f
C409 minus.n20 gnd 0.036265f
C410 minus.n21 gnd 0.036265f
C411 minus.n22 gnd 0.204419f
C412 minus.n23 gnd 0.038669f
C413 minus.n24 gnd 0.030059f
C414 minus.n25 gnd 0.030059f
C415 minus.n26 gnd 0.030059f
C416 minus.n27 gnd 0.037653f
C417 minus.n28 gnd 0.204419f
C418 minus.n29 gnd 0.03514f
C419 minus.n30 gnd 0.03739f
C420 minus.n31 gnd 0.030059f
C421 minus.n32 gnd 0.030059f
C422 minus.n33 gnd 0.039147f
C423 minus.n34 gnd 0.01245f
C424 minus.t17 gnd 0.546625f
C425 minus.n35 gnd 0.237424f
C426 minus.n36 gnd 0.353195f
C427 minus.n37 gnd 0.030059f
C428 minus.t15 gnd 0.546625f
C429 minus.t12 gnd 0.505432f
C430 minus.n38 gnd 0.204419f
C431 minus.n39 gnd 0.030059f
C432 minus.t7 gnd 0.505432f
C433 minus.n40 gnd 0.024431f
C434 minus.n41 gnd 0.030059f
C435 minus.t6 gnd 0.505432f
C436 minus.t11 gnd 0.505432f
C437 minus.n42 gnd 0.204419f
C438 minus.n43 gnd 0.030059f
C439 minus.t10 gnd 0.505432f
C440 minus.n44 gnd 0.204419f
C441 minus.n45 gnd 0.12903f
C442 minus.t16 gnd 0.505432f
C443 minus.t20 gnd 0.567467f
C444 minus.n46 gnd 0.237182f
C445 minus.n47 gnd 0.236072f
C446 minus.n48 gnd 0.03739f
C447 minus.n49 gnd 0.03514f
C448 minus.n50 gnd 0.030059f
C449 minus.n51 gnd 0.030059f
C450 minus.n52 gnd 0.037653f
C451 minus.n53 gnd 0.024431f
C452 minus.n54 gnd 0.038669f
C453 minus.n55 gnd 0.030059f
C454 minus.n56 gnd 0.030059f
C455 minus.n57 gnd 0.036265f
C456 minus.n58 gnd 0.036265f
C457 minus.n59 gnd 0.204419f
C458 minus.n60 gnd 0.038669f
C459 minus.n61 gnd 0.030059f
C460 minus.n62 gnd 0.030059f
C461 minus.n63 gnd 0.030059f
C462 minus.n64 gnd 0.037653f
C463 minus.n65 gnd 0.204419f
C464 minus.n66 gnd 0.03514f
C465 minus.n67 gnd 0.03739f
C466 minus.n68 gnd 0.030059f
C467 minus.n69 gnd 0.030059f
C468 minus.n70 gnd 0.039147f
C469 minus.n71 gnd 0.01245f
C470 minus.n72 gnd 0.237424f
C471 minus.n73 gnd 0.936615f
C472 minus.n74 gnd 1.40781f
C473 minus.t1 gnd 0.009266f
C474 minus.t4 gnd 0.009266f
C475 minus.n75 gnd 0.030469f
C476 minus.t2 gnd 0.009266f
C477 minus.t0 gnd 0.009266f
C478 minus.n76 gnd 0.030052f
C479 minus.n77 gnd 0.25648f
C480 minus.t3 gnd 0.051575f
C481 minus.n78 gnd 0.139959f
C482 minus.n79 gnd 1.89864f
C483 a_n2903_n3924.n0 gnd 1.45586f
C484 a_n2903_n3924.t10 gnd 0.088483f
C485 a_n2903_n3924.t19 gnd 0.919619f
C486 a_n2903_n3924.n1 gnd 0.347657f
C487 a_n2903_n3924.t37 gnd 1.14306f
C488 a_n2903_n3924.n2 gnd 1.19083f
C489 a_n2903_n3924.t6 gnd 0.919619f
C490 a_n2903_n3924.n3 gnd 0.347657f
C491 a_n2903_n3924.t3 gnd 0.088483f
C492 a_n2903_n3924.t35 gnd 0.088483f
C493 a_n2903_n3924.n4 gnd 0.722655f
C494 a_n2903_n3924.n5 gnd 0.364177f
C495 a_n2903_n3924.t32 gnd 0.088483f
C496 a_n2903_n3924.t39 gnd 0.088483f
C497 a_n2903_n3924.n6 gnd 0.722655f
C498 a_n2903_n3924.n7 gnd 0.364177f
C499 a_n2903_n3924.t38 gnd 0.088483f
C500 a_n2903_n3924.t34 gnd 0.088483f
C501 a_n2903_n3924.n8 gnd 0.722655f
C502 a_n2903_n3924.n9 gnd 0.364177f
C503 a_n2903_n3924.t4 gnd 0.919619f
C504 a_n2903_n3924.n10 gnd 0.860834f
C505 a_n2903_n3924.t27 gnd 1.14419f
C506 a_n2903_n3924.t25 gnd 1.14261f
C507 a_n2903_n3924.n11 gnd 0.745791f
C508 a_n2903_n3924.t29 gnd 1.14261f
C509 a_n2903_n3924.n12 gnd 0.804756f
C510 a_n2903_n3924.t31 gnd 1.14261f
C511 a_n2903_n3924.n13 gnd 0.804756f
C512 a_n2903_n3924.t28 gnd 1.14261f
C513 a_n2903_n3924.n14 gnd 0.804756f
C514 a_n2903_n3924.t7 gnd 1.14261f
C515 a_n2903_n3924.n15 gnd 0.804756f
C516 a_n2903_n3924.t36 gnd 1.14261f
C517 a_n2903_n3924.n16 gnd 0.834168f
C518 a_n2903_n3924.t21 gnd 0.919616f
C519 a_n2903_n3924.n17 gnd 0.571219f
C520 a_n2903_n3924.t22 gnd 0.088483f
C521 a_n2903_n3924.t12 gnd 0.088483f
C522 a_n2903_n3924.n18 gnd 0.722654f
C523 a_n2903_n3924.n19 gnd 0.364178f
C524 a_n2903_n3924.t13 gnd 0.088483f
C525 a_n2903_n3924.t8 gnd 0.088483f
C526 a_n2903_n3924.n20 gnd 0.722654f
C527 a_n2903_n3924.n21 gnd 0.364178f
C528 a_n2903_n3924.t9 gnd 0.088483f
C529 a_n2903_n3924.t20 gnd 0.088483f
C530 a_n2903_n3924.n22 gnd 0.722654f
C531 a_n2903_n3924.n23 gnd 0.364178f
C532 a_n2903_n3924.t17 gnd 0.919616f
C533 a_n2903_n3924.n24 gnd 0.347661f
C534 a_n2903_n3924.t5 gnd 0.919616f
C535 a_n2903_n3924.n25 gnd 0.347661f
C536 a_n2903_n3924.t30 gnd 0.088483f
C537 a_n2903_n3924.t33 gnd 0.088483f
C538 a_n2903_n3924.n26 gnd 0.722654f
C539 a_n2903_n3924.n27 gnd 0.364178f
C540 a_n2903_n3924.t0 gnd 0.088483f
C541 a_n2903_n3924.t26 gnd 0.088483f
C542 a_n2903_n3924.n28 gnd 0.722654f
C543 a_n2903_n3924.n29 gnd 0.364178f
C544 a_n2903_n3924.t2 gnd 0.088483f
C545 a_n2903_n3924.t24 gnd 0.088483f
C546 a_n2903_n3924.n30 gnd 0.722654f
C547 a_n2903_n3924.n31 gnd 0.364178f
C548 a_n2903_n3924.t1 gnd 0.919616f
C549 a_n2903_n3924.n32 gnd 0.571219f
C550 a_n2903_n3924.n33 gnd 0.834168f
C551 a_n2903_n3924.t16 gnd 0.919616f
C552 a_n2903_n3924.n34 gnd 0.860837f
C553 a_n2903_n3924.t14 gnd 0.088483f
C554 a_n2903_n3924.t18 gnd 0.088483f
C555 a_n2903_n3924.n35 gnd 0.722655f
C556 a_n2903_n3924.n36 gnd 0.364177f
C557 a_n2903_n3924.t11 gnd 0.088483f
C558 a_n2903_n3924.t15 gnd 0.088483f
C559 a_n2903_n3924.n37 gnd 0.722655f
C560 a_n2903_n3924.n38 gnd 0.364177f
C561 a_n2903_n3924.n39 gnd 0.364176f
C562 a_n2903_n3924.n40 gnd 0.722656f
C563 a_n2903_n3924.t23 gnd 0.088483f
C564 plus.n0 gnd 0.022051f
C565 plus.t7 gnd 0.401003f
C566 plus.t6 gnd 0.370784f
C567 plus.n1 gnd 0.149962f
C568 plus.n2 gnd 0.022051f
C569 plus.t16 gnd 0.370784f
C570 plus.n3 gnd 0.017923f
C571 plus.n4 gnd 0.022051f
C572 plus.t15 gnd 0.370784f
C573 plus.t20 gnd 0.370784f
C574 plus.n5 gnd 0.149962f
C575 plus.n6 gnd 0.022051f
C576 plus.t19 gnd 0.370784f
C577 plus.n7 gnd 0.149962f
C578 plus.n8 gnd 0.094656f
C579 plus.t8 gnd 0.370784f
C580 plus.t11 gnd 0.416293f
C581 plus.n9 gnd 0.173997f
C582 plus.n10 gnd 0.173182f
C583 plus.n11 gnd 0.02743f
C584 plus.n12 gnd 0.025779f
C585 plus.n13 gnd 0.022051f
C586 plus.n14 gnd 0.022051f
C587 plus.n15 gnd 0.027622f
C588 plus.n16 gnd 0.017923f
C589 plus.n17 gnd 0.028368f
C590 plus.n18 gnd 0.022051f
C591 plus.n19 gnd 0.022051f
C592 plus.n20 gnd 0.026604f
C593 plus.n21 gnd 0.026604f
C594 plus.n22 gnd 0.149962f
C595 plus.n23 gnd 0.028368f
C596 plus.n24 gnd 0.022051f
C597 plus.n25 gnd 0.022051f
C598 plus.n26 gnd 0.022051f
C599 plus.n27 gnd 0.027622f
C600 plus.n28 gnd 0.149962f
C601 plus.n29 gnd 0.025779f
C602 plus.n30 gnd 0.02743f
C603 plus.n31 gnd 0.022051f
C604 plus.n32 gnd 0.022051f
C605 plus.n33 gnd 0.028719f
C606 plus.n34 gnd 0.009133f
C607 plus.n35 gnd 0.174174f
C608 plus.n36 gnd 0.253432f
C609 plus.n37 gnd 0.022051f
C610 plus.t10 gnd 0.370784f
C611 plus.n38 gnd 0.149962f
C612 plus.n39 gnd 0.022051f
C613 plus.t14 gnd 0.370784f
C614 plus.n40 gnd 0.017923f
C615 plus.n41 gnd 0.022051f
C616 plus.t13 gnd 0.370784f
C617 plus.t17 gnd 0.370784f
C618 plus.n42 gnd 0.149962f
C619 plus.n43 gnd 0.022051f
C620 plus.t18 gnd 0.370784f
C621 plus.n44 gnd 0.149962f
C622 plus.n45 gnd 0.094656f
C623 plus.t5 gnd 0.370784f
C624 plus.t9 gnd 0.416293f
C625 plus.n46 gnd 0.173997f
C626 plus.n47 gnd 0.173182f
C627 plus.n48 gnd 0.02743f
C628 plus.n49 gnd 0.025779f
C629 plus.n50 gnd 0.022051f
C630 plus.n51 gnd 0.022051f
C631 plus.n52 gnd 0.027622f
C632 plus.n53 gnd 0.017923f
C633 plus.n54 gnd 0.028368f
C634 plus.n55 gnd 0.022051f
C635 plus.n56 gnd 0.022051f
C636 plus.n57 gnd 0.026604f
C637 plus.n58 gnd 0.026604f
C638 plus.n59 gnd 0.149962f
C639 plus.n60 gnd 0.028368f
C640 plus.n61 gnd 0.022051f
C641 plus.n62 gnd 0.022051f
C642 plus.n63 gnd 0.022051f
C643 plus.n64 gnd 0.027622f
C644 plus.n65 gnd 0.149962f
C645 plus.n66 gnd 0.025779f
C646 plus.n67 gnd 0.02743f
C647 plus.n68 gnd 0.022051f
C648 plus.n69 gnd 0.022051f
C649 plus.n70 gnd 0.028719f
C650 plus.n71 gnd 0.009133f
C651 plus.t12 gnd 0.401003f
C652 plus.n72 gnd 0.174174f
C653 plus.n73 gnd 0.678265f
C654 plus.n74 gnd 1.02402f
C655 plus.t4 gnd 0.038066f
C656 plus.t1 gnd 0.006798f
C657 plus.t2 gnd 0.006798f
C658 plus.n75 gnd 0.022046f
C659 plus.n76 gnd 0.171146f
C660 plus.t0 gnd 0.006798f
C661 plus.t3 gnd 0.006798f
C662 plus.n77 gnd 0.022046f
C663 plus.n78 gnd 0.128466f
C664 plus.n79 gnd 2.48089f
C665 a_n2318_8322.t2 gnd 39.6105f
C666 a_n2318_8322.t1 gnd 28.4578f
C667 a_n2318_8322.t3 gnd 19.7356f
C668 a_n2318_8322.t0 gnd 39.6105f
C669 a_n2318_8322.t25 gnd 0.897035f
C670 a_n2318_8322.t22 gnd 0.095802f
C671 a_n2318_8322.t19 gnd 0.095802f
C672 a_n2318_8322.n0 gnd 0.674826f
C673 a_n2318_8322.n1 gnd 0.754021f
C674 a_n2318_8322.t16 gnd 0.095802f
C675 a_n2318_8322.t27 gnd 0.095802f
C676 a_n2318_8322.n2 gnd 0.674826f
C677 a_n2318_8322.n3 gnd 0.383107f
C678 a_n2318_8322.t24 gnd 0.095802f
C679 a_n2318_8322.t17 gnd 0.095802f
C680 a_n2318_8322.n4 gnd 0.674826f
C681 a_n2318_8322.n5 gnd 0.383107f
C682 a_n2318_8322.t15 gnd 0.895251f
C683 a_n2318_8322.n6 gnd 0.881306f
C684 a_n2318_8322.n7 gnd 3.41645f
C685 a_n2318_8322.t7 gnd 0.897038f
C686 a_n2318_8322.t11 gnd 0.095802f
C687 a_n2318_8322.t10 gnd 0.095802f
C688 a_n2318_8322.n8 gnd 0.674826f
C689 a_n2318_8322.n9 gnd 0.754019f
C690 a_n2318_8322.t5 gnd 0.895251f
C691 a_n2318_8322.n10 gnd 0.379433f
C692 a_n2318_8322.t8 gnd 0.895251f
C693 a_n2318_8322.n11 gnd 0.379433f
C694 a_n2318_8322.t6 gnd 0.095802f
C695 a_n2318_8322.t4 gnd 0.095802f
C696 a_n2318_8322.n12 gnd 0.674826f
C697 a_n2318_8322.n13 gnd 0.383107f
C698 a_n2318_8322.t9 gnd 0.895251f
C699 a_n2318_8322.n14 gnd 1.07447f
C700 a_n2318_8322.n15 gnd 1.82651f
C701 a_n2318_8322.t12 gnd 0.895251f
C702 a_n2318_8322.n16 gnd 1.5516f
C703 a_n2318_8322.t21 gnd 0.095802f
C704 a_n2318_8322.t20 gnd 0.095802f
C705 a_n2318_8322.n17 gnd 0.674826f
C706 a_n2318_8322.n18 gnd 0.383107f
C707 a_n2318_8322.t23 gnd 0.095802f
C708 a_n2318_8322.t18 gnd 0.095802f
C709 a_n2318_8322.n19 gnd 0.674826f
C710 a_n2318_8322.n20 gnd 0.383107f
C711 a_n2318_8322.t14 gnd 0.095802f
C712 a_n2318_8322.t13 gnd 0.095802f
C713 a_n2318_8322.n21 gnd 0.674826f
C714 a_n2318_8322.n22 gnd 0.754019f
C715 a_n2318_8322.t26 gnd 0.897038f
C716 commonsourceibias.n0 gnd 0.012624f
C717 commonsourceibias.t120 gnd 0.191163f
C718 commonsourceibias.t67 gnd 0.176757f
C719 commonsourceibias.n1 gnd 0.00769f
C720 commonsourceibias.n2 gnd 0.009461f
C721 commonsourceibias.t126 gnd 0.176757f
C722 commonsourceibias.n3 gnd 0.009597f
C723 commonsourceibias.n4 gnd 0.009461f
C724 commonsourceibias.t121 gnd 0.176757f
C725 commonsourceibias.n5 gnd 0.070526f
C726 commonsourceibias.t136 gnd 0.176757f
C727 commonsourceibias.n6 gnd 0.007653f
C728 commonsourceibias.n7 gnd 0.009461f
C729 commonsourceibias.t117 gnd 0.176757f
C730 commonsourceibias.n8 gnd 0.009134f
C731 commonsourceibias.n9 gnd 0.009461f
C732 commonsourceibias.t102 gnd 0.176757f
C733 commonsourceibias.n10 gnd 0.070526f
C734 commonsourceibias.t125 gnd 0.176757f
C735 commonsourceibias.n11 gnd 0.007641f
C736 commonsourceibias.n12 gnd 0.012624f
C737 commonsourceibias.t34 gnd 0.191163f
C738 commonsourceibias.t42 gnd 0.176757f
C739 commonsourceibias.n13 gnd 0.00769f
C740 commonsourceibias.n14 gnd 0.009461f
C741 commonsourceibias.t60 gnd 0.176757f
C742 commonsourceibias.n15 gnd 0.009597f
C743 commonsourceibias.n16 gnd 0.009461f
C744 commonsourceibias.t32 gnd 0.176757f
C745 commonsourceibias.n17 gnd 0.070526f
C746 commonsourceibias.t22 gnd 0.176757f
C747 commonsourceibias.n18 gnd 0.007653f
C748 commonsourceibias.n19 gnd 0.009461f
C749 commonsourceibias.t0 gnd 0.176757f
C750 commonsourceibias.n20 gnd 0.009134f
C751 commonsourceibias.n21 gnd 0.009461f
C752 commonsourceibias.t18 gnd 0.176757f
C753 commonsourceibias.n22 gnd 0.070526f
C754 commonsourceibias.t62 gnd 0.176757f
C755 commonsourceibias.n23 gnd 0.007641f
C756 commonsourceibias.n24 gnd 0.009461f
C757 commonsourceibias.t36 gnd 0.176757f
C758 commonsourceibias.t48 gnd 0.176757f
C759 commonsourceibias.n25 gnd 0.070526f
C760 commonsourceibias.n26 gnd 0.009461f
C761 commonsourceibias.t14 gnd 0.176757f
C762 commonsourceibias.n27 gnd 0.070526f
C763 commonsourceibias.n28 gnd 0.009461f
C764 commonsourceibias.t20 gnd 0.176757f
C765 commonsourceibias.n29 gnd 0.070526f
C766 commonsourceibias.n30 gnd 0.009461f
C767 commonsourceibias.t50 gnd 0.176757f
C768 commonsourceibias.n31 gnd 0.010754f
C769 commonsourceibias.n32 gnd 0.009461f
C770 commonsourceibias.t2 gnd 0.176757f
C771 commonsourceibias.n33 gnd 0.012717f
C772 commonsourceibias.t12 gnd 0.196904f
C773 commonsourceibias.t52 gnd 0.176757f
C774 commonsourceibias.n34 gnd 0.078584f
C775 commonsourceibias.n35 gnd 0.084191f
C776 commonsourceibias.n36 gnd 0.04027f
C777 commonsourceibias.n37 gnd 0.009461f
C778 commonsourceibias.n38 gnd 0.00769f
C779 commonsourceibias.n39 gnd 0.013037f
C780 commonsourceibias.n40 gnd 0.070526f
C781 commonsourceibias.n41 gnd 0.013093f
C782 commonsourceibias.n42 gnd 0.009461f
C783 commonsourceibias.n43 gnd 0.009461f
C784 commonsourceibias.n44 gnd 0.009461f
C785 commonsourceibias.n45 gnd 0.009597f
C786 commonsourceibias.n46 gnd 0.070526f
C787 commonsourceibias.n47 gnd 0.011661f
C788 commonsourceibias.n48 gnd 0.0129f
C789 commonsourceibias.n49 gnd 0.009461f
C790 commonsourceibias.n50 gnd 0.009461f
C791 commonsourceibias.n51 gnd 0.012816f
C792 commonsourceibias.n52 gnd 0.007653f
C793 commonsourceibias.n53 gnd 0.012975f
C794 commonsourceibias.n54 gnd 0.009461f
C795 commonsourceibias.n55 gnd 0.009461f
C796 commonsourceibias.n56 gnd 0.013054f
C797 commonsourceibias.n57 gnd 0.011256f
C798 commonsourceibias.n58 gnd 0.009134f
C799 commonsourceibias.n59 gnd 0.009461f
C800 commonsourceibias.n60 gnd 0.009461f
C801 commonsourceibias.n61 gnd 0.011572f
C802 commonsourceibias.n62 gnd 0.012989f
C803 commonsourceibias.n63 gnd 0.070526f
C804 commonsourceibias.n64 gnd 0.012901f
C805 commonsourceibias.n65 gnd 0.009461f
C806 commonsourceibias.n66 gnd 0.009461f
C807 commonsourceibias.n67 gnd 0.009461f
C808 commonsourceibias.n68 gnd 0.012901f
C809 commonsourceibias.n69 gnd 0.070526f
C810 commonsourceibias.n70 gnd 0.012989f
C811 commonsourceibias.n71 gnd 0.011572f
C812 commonsourceibias.n72 gnd 0.009461f
C813 commonsourceibias.n73 gnd 0.009461f
C814 commonsourceibias.n74 gnd 0.009461f
C815 commonsourceibias.n75 gnd 0.011256f
C816 commonsourceibias.n76 gnd 0.013054f
C817 commonsourceibias.n77 gnd 0.070526f
C818 commonsourceibias.n78 gnd 0.012975f
C819 commonsourceibias.n79 gnd 0.009461f
C820 commonsourceibias.n80 gnd 0.009461f
C821 commonsourceibias.n81 gnd 0.009461f
C822 commonsourceibias.n82 gnd 0.012816f
C823 commonsourceibias.n83 gnd 0.070526f
C824 commonsourceibias.n84 gnd 0.0129f
C825 commonsourceibias.n85 gnd 0.011661f
C826 commonsourceibias.n86 gnd 0.009461f
C827 commonsourceibias.n87 gnd 0.009461f
C828 commonsourceibias.n88 gnd 0.009461f
C829 commonsourceibias.n89 gnd 0.010754f
C830 commonsourceibias.n90 gnd 0.013093f
C831 commonsourceibias.n91 gnd 0.070526f
C832 commonsourceibias.n92 gnd 0.013037f
C833 commonsourceibias.n93 gnd 0.009461f
C834 commonsourceibias.n94 gnd 0.009461f
C835 commonsourceibias.n95 gnd 0.009461f
C836 commonsourceibias.n96 gnd 0.012717f
C837 commonsourceibias.n97 gnd 0.070526f
C838 commonsourceibias.n98 gnd 0.012748f
C839 commonsourceibias.n99 gnd 0.085044f
C840 commonsourceibias.n100 gnd 0.095092f
C841 commonsourceibias.t35 gnd 0.020415f
C842 commonsourceibias.t43 gnd 0.020415f
C843 commonsourceibias.n101 gnd 0.180398f
C844 commonsourceibias.n102 gnd 0.156264f
C845 commonsourceibias.t61 gnd 0.020415f
C846 commonsourceibias.t33 gnd 0.020415f
C847 commonsourceibias.n103 gnd 0.180398f
C848 commonsourceibias.n104 gnd 0.082864f
C849 commonsourceibias.t23 gnd 0.020415f
C850 commonsourceibias.t1 gnd 0.020415f
C851 commonsourceibias.n105 gnd 0.180398f
C852 commonsourceibias.n106 gnd 0.082864f
C853 commonsourceibias.t19 gnd 0.020415f
C854 commonsourceibias.t63 gnd 0.020415f
C855 commonsourceibias.n107 gnd 0.180398f
C856 commonsourceibias.n108 gnd 0.069229f
C857 commonsourceibias.t53 gnd 0.020415f
C858 commonsourceibias.t13 gnd 0.020415f
C859 commonsourceibias.n109 gnd 0.181002f
C860 commonsourceibias.t51 gnd 0.020415f
C861 commonsourceibias.t3 gnd 0.020415f
C862 commonsourceibias.n110 gnd 0.180398f
C863 commonsourceibias.n111 gnd 0.168097f
C864 commonsourceibias.t15 gnd 0.020415f
C865 commonsourceibias.t21 gnd 0.020415f
C866 commonsourceibias.n112 gnd 0.180398f
C867 commonsourceibias.n113 gnd 0.082864f
C868 commonsourceibias.t37 gnd 0.020415f
C869 commonsourceibias.t49 gnd 0.020415f
C870 commonsourceibias.n114 gnd 0.180398f
C871 commonsourceibias.n115 gnd 0.069229f
C872 commonsourceibias.n116 gnd 0.083829f
C873 commonsourceibias.n117 gnd 0.009461f
C874 commonsourceibias.t118 gnd 0.176757f
C875 commonsourceibias.t76 gnd 0.176757f
C876 commonsourceibias.n118 gnd 0.070526f
C877 commonsourceibias.n119 gnd 0.009461f
C878 commonsourceibias.t106 gnd 0.176757f
C879 commonsourceibias.n120 gnd 0.070526f
C880 commonsourceibias.n121 gnd 0.009461f
C881 commonsourceibias.t96 gnd 0.176757f
C882 commonsourceibias.n122 gnd 0.070526f
C883 commonsourceibias.n123 gnd 0.009461f
C884 commonsourceibias.t141 gnd 0.176757f
C885 commonsourceibias.n124 gnd 0.010754f
C886 commonsourceibias.n125 gnd 0.009461f
C887 commonsourceibias.t116 gnd 0.176757f
C888 commonsourceibias.n126 gnd 0.012717f
C889 commonsourceibias.t129 gnd 0.196904f
C890 commonsourceibias.t152 gnd 0.176757f
C891 commonsourceibias.n127 gnd 0.078584f
C892 commonsourceibias.n128 gnd 0.084191f
C893 commonsourceibias.n129 gnd 0.04027f
C894 commonsourceibias.n130 gnd 0.009461f
C895 commonsourceibias.n131 gnd 0.00769f
C896 commonsourceibias.n132 gnd 0.013037f
C897 commonsourceibias.n133 gnd 0.070526f
C898 commonsourceibias.n134 gnd 0.013093f
C899 commonsourceibias.n135 gnd 0.009461f
C900 commonsourceibias.n136 gnd 0.009461f
C901 commonsourceibias.n137 gnd 0.009461f
C902 commonsourceibias.n138 gnd 0.009597f
C903 commonsourceibias.n139 gnd 0.070526f
C904 commonsourceibias.n140 gnd 0.011661f
C905 commonsourceibias.n141 gnd 0.0129f
C906 commonsourceibias.n142 gnd 0.009461f
C907 commonsourceibias.n143 gnd 0.009461f
C908 commonsourceibias.n144 gnd 0.012816f
C909 commonsourceibias.n145 gnd 0.007653f
C910 commonsourceibias.n146 gnd 0.012975f
C911 commonsourceibias.n147 gnd 0.009461f
C912 commonsourceibias.n148 gnd 0.009461f
C913 commonsourceibias.n149 gnd 0.013054f
C914 commonsourceibias.n150 gnd 0.011256f
C915 commonsourceibias.n151 gnd 0.009134f
C916 commonsourceibias.n152 gnd 0.009461f
C917 commonsourceibias.n153 gnd 0.009461f
C918 commonsourceibias.n154 gnd 0.011572f
C919 commonsourceibias.n155 gnd 0.012989f
C920 commonsourceibias.n156 gnd 0.070526f
C921 commonsourceibias.n157 gnd 0.012901f
C922 commonsourceibias.n158 gnd 0.009415f
C923 commonsourceibias.n159 gnd 0.06839f
C924 commonsourceibias.n160 gnd 0.009415f
C925 commonsourceibias.n161 gnd 0.012901f
C926 commonsourceibias.n162 gnd 0.070526f
C927 commonsourceibias.n163 gnd 0.012989f
C928 commonsourceibias.n164 gnd 0.011572f
C929 commonsourceibias.n165 gnd 0.009461f
C930 commonsourceibias.n166 gnd 0.009461f
C931 commonsourceibias.n167 gnd 0.009461f
C932 commonsourceibias.n168 gnd 0.011256f
C933 commonsourceibias.n169 gnd 0.013054f
C934 commonsourceibias.n170 gnd 0.070526f
C935 commonsourceibias.n171 gnd 0.012975f
C936 commonsourceibias.n172 gnd 0.009461f
C937 commonsourceibias.n173 gnd 0.009461f
C938 commonsourceibias.n174 gnd 0.009461f
C939 commonsourceibias.n175 gnd 0.012816f
C940 commonsourceibias.n176 gnd 0.070526f
C941 commonsourceibias.n177 gnd 0.0129f
C942 commonsourceibias.n178 gnd 0.011661f
C943 commonsourceibias.n179 gnd 0.009461f
C944 commonsourceibias.n180 gnd 0.009461f
C945 commonsourceibias.n181 gnd 0.009461f
C946 commonsourceibias.n182 gnd 0.010754f
C947 commonsourceibias.n183 gnd 0.013093f
C948 commonsourceibias.n184 gnd 0.070526f
C949 commonsourceibias.n185 gnd 0.013037f
C950 commonsourceibias.n186 gnd 0.009461f
C951 commonsourceibias.n187 gnd 0.009461f
C952 commonsourceibias.n188 gnd 0.009461f
C953 commonsourceibias.n189 gnd 0.012717f
C954 commonsourceibias.n190 gnd 0.070526f
C955 commonsourceibias.n191 gnd 0.012748f
C956 commonsourceibias.n192 gnd 0.085044f
C957 commonsourceibias.n193 gnd 0.056182f
C958 commonsourceibias.n194 gnd 0.012624f
C959 commonsourceibias.t71 gnd 0.191163f
C960 commonsourceibias.t159 gnd 0.176757f
C961 commonsourceibias.n195 gnd 0.00769f
C962 commonsourceibias.n196 gnd 0.009461f
C963 commonsourceibias.t148 gnd 0.176757f
C964 commonsourceibias.n197 gnd 0.009597f
C965 commonsourceibias.n198 gnd 0.009461f
C966 commonsourceibias.t78 gnd 0.176757f
C967 commonsourceibias.n199 gnd 0.070526f
C968 commonsourceibias.t157 gnd 0.176757f
C969 commonsourceibias.n200 gnd 0.007653f
C970 commonsourceibias.n201 gnd 0.009461f
C971 commonsourceibias.t85 gnd 0.176757f
C972 commonsourceibias.n202 gnd 0.009134f
C973 commonsourceibias.n203 gnd 0.009461f
C974 commonsourceibias.t77 gnd 0.176757f
C975 commonsourceibias.n204 gnd 0.070526f
C976 commonsourceibias.t158 gnd 0.176757f
C977 commonsourceibias.n205 gnd 0.007641f
C978 commonsourceibias.n206 gnd 0.009461f
C979 commonsourceibias.t94 gnd 0.176757f
C980 commonsourceibias.t113 gnd 0.176757f
C981 commonsourceibias.n207 gnd 0.070526f
C982 commonsourceibias.n208 gnd 0.009461f
C983 commonsourceibias.t156 gnd 0.176757f
C984 commonsourceibias.n209 gnd 0.070526f
C985 commonsourceibias.n210 gnd 0.009461f
C986 commonsourceibias.t92 gnd 0.176757f
C987 commonsourceibias.n211 gnd 0.070526f
C988 commonsourceibias.n212 gnd 0.009461f
C989 commonsourceibias.t111 gnd 0.176757f
C990 commonsourceibias.n213 gnd 0.010754f
C991 commonsourceibias.n214 gnd 0.009461f
C992 commonsourceibias.t105 gnd 0.176757f
C993 commonsourceibias.n215 gnd 0.012717f
C994 commonsourceibias.t112 gnd 0.196904f
C995 commonsourceibias.t93 gnd 0.176757f
C996 commonsourceibias.n216 gnd 0.078584f
C997 commonsourceibias.n217 gnd 0.084191f
C998 commonsourceibias.n218 gnd 0.04027f
C999 commonsourceibias.n219 gnd 0.009461f
C1000 commonsourceibias.n220 gnd 0.00769f
C1001 commonsourceibias.n221 gnd 0.013037f
C1002 commonsourceibias.n222 gnd 0.070526f
C1003 commonsourceibias.n223 gnd 0.013093f
C1004 commonsourceibias.n224 gnd 0.009461f
C1005 commonsourceibias.n225 gnd 0.009461f
C1006 commonsourceibias.n226 gnd 0.009461f
C1007 commonsourceibias.n227 gnd 0.009597f
C1008 commonsourceibias.n228 gnd 0.070526f
C1009 commonsourceibias.n229 gnd 0.011661f
C1010 commonsourceibias.n230 gnd 0.0129f
C1011 commonsourceibias.n231 gnd 0.009461f
C1012 commonsourceibias.n232 gnd 0.009461f
C1013 commonsourceibias.n233 gnd 0.012816f
C1014 commonsourceibias.n234 gnd 0.007653f
C1015 commonsourceibias.n235 gnd 0.012975f
C1016 commonsourceibias.n236 gnd 0.009461f
C1017 commonsourceibias.n237 gnd 0.009461f
C1018 commonsourceibias.n238 gnd 0.013054f
C1019 commonsourceibias.n239 gnd 0.011256f
C1020 commonsourceibias.n240 gnd 0.009134f
C1021 commonsourceibias.n241 gnd 0.009461f
C1022 commonsourceibias.n242 gnd 0.009461f
C1023 commonsourceibias.n243 gnd 0.011572f
C1024 commonsourceibias.n244 gnd 0.012989f
C1025 commonsourceibias.n245 gnd 0.070526f
C1026 commonsourceibias.n246 gnd 0.012901f
C1027 commonsourceibias.n247 gnd 0.009461f
C1028 commonsourceibias.n248 gnd 0.009461f
C1029 commonsourceibias.n249 gnd 0.009461f
C1030 commonsourceibias.n250 gnd 0.012901f
C1031 commonsourceibias.n251 gnd 0.070526f
C1032 commonsourceibias.n252 gnd 0.012989f
C1033 commonsourceibias.n253 gnd 0.011572f
C1034 commonsourceibias.n254 gnd 0.009461f
C1035 commonsourceibias.n255 gnd 0.009461f
C1036 commonsourceibias.n256 gnd 0.009461f
C1037 commonsourceibias.n257 gnd 0.011256f
C1038 commonsourceibias.n258 gnd 0.013054f
C1039 commonsourceibias.n259 gnd 0.070526f
C1040 commonsourceibias.n260 gnd 0.012975f
C1041 commonsourceibias.n261 gnd 0.009461f
C1042 commonsourceibias.n262 gnd 0.009461f
C1043 commonsourceibias.n263 gnd 0.009461f
C1044 commonsourceibias.n264 gnd 0.012816f
C1045 commonsourceibias.n265 gnd 0.070526f
C1046 commonsourceibias.n266 gnd 0.0129f
C1047 commonsourceibias.n267 gnd 0.011661f
C1048 commonsourceibias.n268 gnd 0.009461f
C1049 commonsourceibias.n269 gnd 0.009461f
C1050 commonsourceibias.n270 gnd 0.009461f
C1051 commonsourceibias.n271 gnd 0.010754f
C1052 commonsourceibias.n272 gnd 0.013093f
C1053 commonsourceibias.n273 gnd 0.070526f
C1054 commonsourceibias.n274 gnd 0.013037f
C1055 commonsourceibias.n275 gnd 0.009461f
C1056 commonsourceibias.n276 gnd 0.009461f
C1057 commonsourceibias.n277 gnd 0.009461f
C1058 commonsourceibias.n278 gnd 0.012717f
C1059 commonsourceibias.n279 gnd 0.070526f
C1060 commonsourceibias.n280 gnd 0.012748f
C1061 commonsourceibias.n281 gnd 0.085044f
C1062 commonsourceibias.n282 gnd 0.030348f
C1063 commonsourceibias.n283 gnd 0.15151f
C1064 commonsourceibias.n284 gnd 0.012624f
C1065 commonsourceibias.t75 gnd 0.176757f
C1066 commonsourceibias.n285 gnd 0.00769f
C1067 commonsourceibias.n286 gnd 0.009461f
C1068 commonsourceibias.t128 gnd 0.176757f
C1069 commonsourceibias.n287 gnd 0.009597f
C1070 commonsourceibias.n288 gnd 0.009461f
C1071 commonsourceibias.t124 gnd 0.176757f
C1072 commonsourceibias.n289 gnd 0.070526f
C1073 commonsourceibias.t155 gnd 0.176757f
C1074 commonsourceibias.n290 gnd 0.007653f
C1075 commonsourceibias.n291 gnd 0.009461f
C1076 commonsourceibias.t90 gnd 0.176757f
C1077 commonsourceibias.n292 gnd 0.009134f
C1078 commonsourceibias.n293 gnd 0.009461f
C1079 commonsourceibias.t119 gnd 0.176757f
C1080 commonsourceibias.n294 gnd 0.070526f
C1081 commonsourceibias.t146 gnd 0.176757f
C1082 commonsourceibias.n295 gnd 0.007641f
C1083 commonsourceibias.n296 gnd 0.009461f
C1084 commonsourceibias.t138 gnd 0.176757f
C1085 commonsourceibias.t64 gnd 0.176757f
C1086 commonsourceibias.n297 gnd 0.070526f
C1087 commonsourceibias.n298 gnd 0.009461f
C1088 commonsourceibias.t137 gnd 0.176757f
C1089 commonsourceibias.n299 gnd 0.070526f
C1090 commonsourceibias.n300 gnd 0.009461f
C1091 commonsourceibias.t133 gnd 0.176757f
C1092 commonsourceibias.n301 gnd 0.070526f
C1093 commonsourceibias.n302 gnd 0.009461f
C1094 commonsourceibias.t149 gnd 0.176757f
C1095 commonsourceibias.n303 gnd 0.010754f
C1096 commonsourceibias.n304 gnd 0.009461f
C1097 commonsourceibias.t79 gnd 0.176757f
C1098 commonsourceibias.n305 gnd 0.012717f
C1099 commonsourceibias.t140 gnd 0.196904f
C1100 commonsourceibias.t130 gnd 0.176757f
C1101 commonsourceibias.n306 gnd 0.078584f
C1102 commonsourceibias.n307 gnd 0.084191f
C1103 commonsourceibias.n308 gnd 0.04027f
C1104 commonsourceibias.n309 gnd 0.009461f
C1105 commonsourceibias.n310 gnd 0.00769f
C1106 commonsourceibias.n311 gnd 0.013037f
C1107 commonsourceibias.n312 gnd 0.070526f
C1108 commonsourceibias.n313 gnd 0.013093f
C1109 commonsourceibias.n314 gnd 0.009461f
C1110 commonsourceibias.n315 gnd 0.009461f
C1111 commonsourceibias.n316 gnd 0.009461f
C1112 commonsourceibias.n317 gnd 0.009597f
C1113 commonsourceibias.n318 gnd 0.070526f
C1114 commonsourceibias.n319 gnd 0.011661f
C1115 commonsourceibias.n320 gnd 0.0129f
C1116 commonsourceibias.n321 gnd 0.009461f
C1117 commonsourceibias.n322 gnd 0.009461f
C1118 commonsourceibias.n323 gnd 0.012816f
C1119 commonsourceibias.n324 gnd 0.007653f
C1120 commonsourceibias.n325 gnd 0.012975f
C1121 commonsourceibias.n326 gnd 0.009461f
C1122 commonsourceibias.n327 gnd 0.009461f
C1123 commonsourceibias.n328 gnd 0.013054f
C1124 commonsourceibias.n329 gnd 0.011256f
C1125 commonsourceibias.n330 gnd 0.009134f
C1126 commonsourceibias.n331 gnd 0.009461f
C1127 commonsourceibias.n332 gnd 0.009461f
C1128 commonsourceibias.n333 gnd 0.011572f
C1129 commonsourceibias.n334 gnd 0.012989f
C1130 commonsourceibias.n335 gnd 0.070526f
C1131 commonsourceibias.n336 gnd 0.012901f
C1132 commonsourceibias.n337 gnd 0.009461f
C1133 commonsourceibias.n338 gnd 0.009461f
C1134 commonsourceibias.n339 gnd 0.009461f
C1135 commonsourceibias.n340 gnd 0.012901f
C1136 commonsourceibias.n341 gnd 0.070526f
C1137 commonsourceibias.n342 gnd 0.012989f
C1138 commonsourceibias.n343 gnd 0.011572f
C1139 commonsourceibias.n344 gnd 0.009461f
C1140 commonsourceibias.n345 gnd 0.009461f
C1141 commonsourceibias.n346 gnd 0.009461f
C1142 commonsourceibias.n347 gnd 0.011256f
C1143 commonsourceibias.n348 gnd 0.013054f
C1144 commonsourceibias.n349 gnd 0.070526f
C1145 commonsourceibias.n350 gnd 0.012975f
C1146 commonsourceibias.n351 gnd 0.009461f
C1147 commonsourceibias.n352 gnd 0.009461f
C1148 commonsourceibias.n353 gnd 0.009461f
C1149 commonsourceibias.n354 gnd 0.012816f
C1150 commonsourceibias.n355 gnd 0.070526f
C1151 commonsourceibias.n356 gnd 0.0129f
C1152 commonsourceibias.n357 gnd 0.011661f
C1153 commonsourceibias.n358 gnd 0.009461f
C1154 commonsourceibias.n359 gnd 0.009461f
C1155 commonsourceibias.n360 gnd 0.009461f
C1156 commonsourceibias.n361 gnd 0.010754f
C1157 commonsourceibias.n362 gnd 0.013093f
C1158 commonsourceibias.n363 gnd 0.070526f
C1159 commonsourceibias.n364 gnd 0.013037f
C1160 commonsourceibias.n365 gnd 0.009461f
C1161 commonsourceibias.n366 gnd 0.009461f
C1162 commonsourceibias.n367 gnd 0.009461f
C1163 commonsourceibias.n368 gnd 0.012717f
C1164 commonsourceibias.n369 gnd 0.070526f
C1165 commonsourceibias.n370 gnd 0.012748f
C1166 commonsourceibias.t147 gnd 0.191163f
C1167 commonsourceibias.n371 gnd 0.085044f
C1168 commonsourceibias.n372 gnd 0.030348f
C1169 commonsourceibias.n373 gnd 0.449685f
C1170 commonsourceibias.n374 gnd 0.012624f
C1171 commonsourceibias.t91 gnd 0.191163f
C1172 commonsourceibias.t134 gnd 0.176757f
C1173 commonsourceibias.n375 gnd 0.00769f
C1174 commonsourceibias.n376 gnd 0.009461f
C1175 commonsourceibias.t114 gnd 0.176757f
C1176 commonsourceibias.n377 gnd 0.009597f
C1177 commonsourceibias.n378 gnd 0.009461f
C1178 commonsourceibias.t123 gnd 0.176757f
C1179 commonsourceibias.n379 gnd 0.007653f
C1180 commonsourceibias.n380 gnd 0.009461f
C1181 commonsourceibias.t88 gnd 0.176757f
C1182 commonsourceibias.n381 gnd 0.009134f
C1183 commonsourceibias.n382 gnd 0.009461f
C1184 commonsourceibias.t104 gnd 0.176757f
C1185 commonsourceibias.n383 gnd 0.007641f
C1186 commonsourceibias.n384 gnd 0.009461f
C1187 commonsourceibias.t89 gnd 0.176757f
C1188 commonsourceibias.t139 gnd 0.176757f
C1189 commonsourceibias.n385 gnd 0.070526f
C1190 commonsourceibias.n386 gnd 0.009461f
C1191 commonsourceibias.t83 gnd 0.176757f
C1192 commonsourceibias.n387 gnd 0.070526f
C1193 commonsourceibias.n388 gnd 0.009461f
C1194 commonsourceibias.t150 gnd 0.176757f
C1195 commonsourceibias.n389 gnd 0.070526f
C1196 commonsourceibias.n390 gnd 0.009461f
C1197 commonsourceibias.t127 gnd 0.176757f
C1198 commonsourceibias.n391 gnd 0.010754f
C1199 commonsourceibias.n392 gnd 0.009461f
C1200 commonsourceibias.t84 gnd 0.176757f
C1201 commonsourceibias.n393 gnd 0.012717f
C1202 commonsourceibias.t108 gnd 0.196904f
C1203 commonsourceibias.t131 gnd 0.176757f
C1204 commonsourceibias.n394 gnd 0.078584f
C1205 commonsourceibias.n395 gnd 0.084191f
C1206 commonsourceibias.n396 gnd 0.04027f
C1207 commonsourceibias.n397 gnd 0.009461f
C1208 commonsourceibias.n398 gnd 0.00769f
C1209 commonsourceibias.n399 gnd 0.013037f
C1210 commonsourceibias.n400 gnd 0.070526f
C1211 commonsourceibias.n401 gnd 0.013093f
C1212 commonsourceibias.n402 gnd 0.009461f
C1213 commonsourceibias.n403 gnd 0.009461f
C1214 commonsourceibias.n404 gnd 0.009461f
C1215 commonsourceibias.n405 gnd 0.009597f
C1216 commonsourceibias.n406 gnd 0.070526f
C1217 commonsourceibias.n407 gnd 0.011661f
C1218 commonsourceibias.n408 gnd 0.0129f
C1219 commonsourceibias.n409 gnd 0.009461f
C1220 commonsourceibias.n410 gnd 0.009461f
C1221 commonsourceibias.n411 gnd 0.012816f
C1222 commonsourceibias.n412 gnd 0.007653f
C1223 commonsourceibias.n413 gnd 0.012975f
C1224 commonsourceibias.n414 gnd 0.009461f
C1225 commonsourceibias.n415 gnd 0.009461f
C1226 commonsourceibias.n416 gnd 0.013054f
C1227 commonsourceibias.n417 gnd 0.011256f
C1228 commonsourceibias.n418 gnd 0.009134f
C1229 commonsourceibias.n419 gnd 0.009461f
C1230 commonsourceibias.n420 gnd 0.009461f
C1231 commonsourceibias.n421 gnd 0.011572f
C1232 commonsourceibias.n422 gnd 0.012989f
C1233 commonsourceibias.n423 gnd 0.070526f
C1234 commonsourceibias.n424 gnd 0.012901f
C1235 commonsourceibias.n425 gnd 0.009415f
C1236 commonsourceibias.t31 gnd 0.020415f
C1237 commonsourceibias.t27 gnd 0.020415f
C1238 commonsourceibias.n426 gnd 0.181002f
C1239 commonsourceibias.t45 gnd 0.020415f
C1240 commonsourceibias.t59 gnd 0.020415f
C1241 commonsourceibias.n427 gnd 0.180398f
C1242 commonsourceibias.n428 gnd 0.168097f
C1243 commonsourceibias.t55 gnd 0.020415f
C1244 commonsourceibias.t47 gnd 0.020415f
C1245 commonsourceibias.n429 gnd 0.180398f
C1246 commonsourceibias.n430 gnd 0.082864f
C1247 commonsourceibias.t39 gnd 0.020415f
C1248 commonsourceibias.t9 gnd 0.020415f
C1249 commonsourceibias.n431 gnd 0.180398f
C1250 commonsourceibias.n432 gnd 0.069229f
C1251 commonsourceibias.n433 gnd 0.012624f
C1252 commonsourceibias.t24 gnd 0.176757f
C1253 commonsourceibias.n434 gnd 0.00769f
C1254 commonsourceibias.n435 gnd 0.009461f
C1255 commonsourceibias.t28 gnd 0.176757f
C1256 commonsourceibias.n436 gnd 0.009597f
C1257 commonsourceibias.n437 gnd 0.009461f
C1258 commonsourceibias.t56 gnd 0.176757f
C1259 commonsourceibias.n438 gnd 0.007653f
C1260 commonsourceibias.n439 gnd 0.009461f
C1261 commonsourceibias.t10 gnd 0.176757f
C1262 commonsourceibias.n440 gnd 0.009134f
C1263 commonsourceibias.n441 gnd 0.009461f
C1264 commonsourceibias.t16 gnd 0.176757f
C1265 commonsourceibias.n442 gnd 0.007641f
C1266 commonsourceibias.n443 gnd 0.009461f
C1267 commonsourceibias.t8 gnd 0.176757f
C1268 commonsourceibias.t38 gnd 0.176757f
C1269 commonsourceibias.n444 gnd 0.070526f
C1270 commonsourceibias.n445 gnd 0.009461f
C1271 commonsourceibias.t46 gnd 0.176757f
C1272 commonsourceibias.n446 gnd 0.070526f
C1273 commonsourceibias.n447 gnd 0.009461f
C1274 commonsourceibias.t54 gnd 0.176757f
C1275 commonsourceibias.n448 gnd 0.070526f
C1276 commonsourceibias.n449 gnd 0.009461f
C1277 commonsourceibias.t58 gnd 0.176757f
C1278 commonsourceibias.n450 gnd 0.010754f
C1279 commonsourceibias.n451 gnd 0.009461f
C1280 commonsourceibias.t44 gnd 0.176757f
C1281 commonsourceibias.n452 gnd 0.012717f
C1282 commonsourceibias.t30 gnd 0.196904f
C1283 commonsourceibias.t26 gnd 0.176757f
C1284 commonsourceibias.n453 gnd 0.078584f
C1285 commonsourceibias.n454 gnd 0.084191f
C1286 commonsourceibias.n455 gnd 0.04027f
C1287 commonsourceibias.n456 gnd 0.009461f
C1288 commonsourceibias.n457 gnd 0.00769f
C1289 commonsourceibias.n458 gnd 0.013037f
C1290 commonsourceibias.n459 gnd 0.070526f
C1291 commonsourceibias.n460 gnd 0.013093f
C1292 commonsourceibias.n461 gnd 0.009461f
C1293 commonsourceibias.n462 gnd 0.009461f
C1294 commonsourceibias.n463 gnd 0.009461f
C1295 commonsourceibias.n464 gnd 0.009597f
C1296 commonsourceibias.n465 gnd 0.070526f
C1297 commonsourceibias.n466 gnd 0.011661f
C1298 commonsourceibias.n467 gnd 0.0129f
C1299 commonsourceibias.n468 gnd 0.009461f
C1300 commonsourceibias.n469 gnd 0.009461f
C1301 commonsourceibias.n470 gnd 0.012816f
C1302 commonsourceibias.n471 gnd 0.007653f
C1303 commonsourceibias.n472 gnd 0.012975f
C1304 commonsourceibias.n473 gnd 0.009461f
C1305 commonsourceibias.n474 gnd 0.009461f
C1306 commonsourceibias.n475 gnd 0.013054f
C1307 commonsourceibias.n476 gnd 0.011256f
C1308 commonsourceibias.n477 gnd 0.009134f
C1309 commonsourceibias.n478 gnd 0.009461f
C1310 commonsourceibias.n479 gnd 0.009461f
C1311 commonsourceibias.n480 gnd 0.011572f
C1312 commonsourceibias.n481 gnd 0.012989f
C1313 commonsourceibias.n482 gnd 0.070526f
C1314 commonsourceibias.n483 gnd 0.012901f
C1315 commonsourceibias.n484 gnd 0.009461f
C1316 commonsourceibias.n485 gnd 0.009461f
C1317 commonsourceibias.n486 gnd 0.009461f
C1318 commonsourceibias.n487 gnd 0.012901f
C1319 commonsourceibias.n488 gnd 0.070526f
C1320 commonsourceibias.n489 gnd 0.012989f
C1321 commonsourceibias.t40 gnd 0.176757f
C1322 commonsourceibias.n490 gnd 0.070526f
C1323 commonsourceibias.n491 gnd 0.011572f
C1324 commonsourceibias.n492 gnd 0.009461f
C1325 commonsourceibias.n493 gnd 0.009461f
C1326 commonsourceibias.n494 gnd 0.009461f
C1327 commonsourceibias.n495 gnd 0.011256f
C1328 commonsourceibias.n496 gnd 0.013054f
C1329 commonsourceibias.n497 gnd 0.070526f
C1330 commonsourceibias.n498 gnd 0.012975f
C1331 commonsourceibias.n499 gnd 0.009461f
C1332 commonsourceibias.n500 gnd 0.009461f
C1333 commonsourceibias.n501 gnd 0.009461f
C1334 commonsourceibias.n502 gnd 0.012816f
C1335 commonsourceibias.n503 gnd 0.070526f
C1336 commonsourceibias.n504 gnd 0.0129f
C1337 commonsourceibias.t4 gnd 0.176757f
C1338 commonsourceibias.n505 gnd 0.070526f
C1339 commonsourceibias.n506 gnd 0.011661f
C1340 commonsourceibias.n507 gnd 0.009461f
C1341 commonsourceibias.n508 gnd 0.009461f
C1342 commonsourceibias.n509 gnd 0.009461f
C1343 commonsourceibias.n510 gnd 0.010754f
C1344 commonsourceibias.n511 gnd 0.013093f
C1345 commonsourceibias.n512 gnd 0.070526f
C1346 commonsourceibias.n513 gnd 0.013037f
C1347 commonsourceibias.n514 gnd 0.009461f
C1348 commonsourceibias.n515 gnd 0.009461f
C1349 commonsourceibias.n516 gnd 0.009461f
C1350 commonsourceibias.n517 gnd 0.012717f
C1351 commonsourceibias.n518 gnd 0.070526f
C1352 commonsourceibias.n519 gnd 0.012748f
C1353 commonsourceibias.t6 gnd 0.191163f
C1354 commonsourceibias.n520 gnd 0.085044f
C1355 commonsourceibias.n521 gnd 0.095092f
C1356 commonsourceibias.t25 gnd 0.020415f
C1357 commonsourceibias.t7 gnd 0.020415f
C1358 commonsourceibias.n522 gnd 0.180398f
C1359 commonsourceibias.n523 gnd 0.156264f
C1360 commonsourceibias.t5 gnd 0.020415f
C1361 commonsourceibias.t29 gnd 0.020415f
C1362 commonsourceibias.n524 gnd 0.180398f
C1363 commonsourceibias.n525 gnd 0.082864f
C1364 commonsourceibias.t11 gnd 0.020415f
C1365 commonsourceibias.t57 gnd 0.020415f
C1366 commonsourceibias.n526 gnd 0.180398f
C1367 commonsourceibias.n527 gnd 0.082864f
C1368 commonsourceibias.t17 gnd 0.020415f
C1369 commonsourceibias.t41 gnd 0.020415f
C1370 commonsourceibias.n528 gnd 0.180398f
C1371 commonsourceibias.n529 gnd 0.069229f
C1372 commonsourceibias.n530 gnd 0.083829f
C1373 commonsourceibias.n531 gnd 0.06839f
C1374 commonsourceibias.n532 gnd 0.009415f
C1375 commonsourceibias.n533 gnd 0.012901f
C1376 commonsourceibias.n534 gnd 0.070526f
C1377 commonsourceibias.n535 gnd 0.012989f
C1378 commonsourceibias.t73 gnd 0.176757f
C1379 commonsourceibias.n536 gnd 0.070526f
C1380 commonsourceibias.n537 gnd 0.011572f
C1381 commonsourceibias.n538 gnd 0.009461f
C1382 commonsourceibias.n539 gnd 0.009461f
C1383 commonsourceibias.n540 gnd 0.009461f
C1384 commonsourceibias.n541 gnd 0.011256f
C1385 commonsourceibias.n542 gnd 0.013054f
C1386 commonsourceibias.n543 gnd 0.070526f
C1387 commonsourceibias.n544 gnd 0.012975f
C1388 commonsourceibias.n545 gnd 0.009461f
C1389 commonsourceibias.n546 gnd 0.009461f
C1390 commonsourceibias.n547 gnd 0.009461f
C1391 commonsourceibias.n548 gnd 0.012816f
C1392 commonsourceibias.n549 gnd 0.070526f
C1393 commonsourceibias.n550 gnd 0.0129f
C1394 commonsourceibias.t95 gnd 0.176757f
C1395 commonsourceibias.n551 gnd 0.070526f
C1396 commonsourceibias.n552 gnd 0.011661f
C1397 commonsourceibias.n553 gnd 0.009461f
C1398 commonsourceibias.n554 gnd 0.009461f
C1399 commonsourceibias.n555 gnd 0.009461f
C1400 commonsourceibias.n556 gnd 0.010754f
C1401 commonsourceibias.n557 gnd 0.013093f
C1402 commonsourceibias.n558 gnd 0.070526f
C1403 commonsourceibias.n559 gnd 0.013037f
C1404 commonsourceibias.n560 gnd 0.009461f
C1405 commonsourceibias.n561 gnd 0.009461f
C1406 commonsourceibias.n562 gnd 0.009461f
C1407 commonsourceibias.n563 gnd 0.012717f
C1408 commonsourceibias.n564 gnd 0.070526f
C1409 commonsourceibias.n565 gnd 0.012748f
C1410 commonsourceibias.n566 gnd 0.085044f
C1411 commonsourceibias.n567 gnd 0.056182f
C1412 commonsourceibias.n568 gnd 0.012624f
C1413 commonsourceibias.t144 gnd 0.176757f
C1414 commonsourceibias.n569 gnd 0.00769f
C1415 commonsourceibias.n570 gnd 0.009461f
C1416 commonsourceibias.t66 gnd 0.176757f
C1417 commonsourceibias.n571 gnd 0.009597f
C1418 commonsourceibias.n572 gnd 0.009461f
C1419 commonsourceibias.t143 gnd 0.176757f
C1420 commonsourceibias.n573 gnd 0.007653f
C1421 commonsourceibias.n574 gnd 0.009461f
C1422 commonsourceibias.t65 gnd 0.176757f
C1423 commonsourceibias.n575 gnd 0.009134f
C1424 commonsourceibias.n576 gnd 0.009461f
C1425 commonsourceibias.t142 gnd 0.176757f
C1426 commonsourceibias.n577 gnd 0.007641f
C1427 commonsourceibias.n578 gnd 0.009461f
C1428 commonsourceibias.t72 gnd 0.176757f
C1429 commonsourceibias.t99 gnd 0.176757f
C1430 commonsourceibias.n579 gnd 0.070526f
C1431 commonsourceibias.n580 gnd 0.009461f
C1432 commonsourceibias.t80 gnd 0.176757f
C1433 commonsourceibias.n581 gnd 0.070526f
C1434 commonsourceibias.n582 gnd 0.009461f
C1435 commonsourceibias.t69 gnd 0.176757f
C1436 commonsourceibias.n583 gnd 0.070526f
C1437 commonsourceibias.n584 gnd 0.009461f
C1438 commonsourceibias.t98 gnd 0.176757f
C1439 commonsourceibias.n585 gnd 0.010754f
C1440 commonsourceibias.n586 gnd 0.009461f
C1441 commonsourceibias.t86 gnd 0.176757f
C1442 commonsourceibias.n587 gnd 0.012717f
C1443 commonsourceibias.t97 gnd 0.196904f
C1444 commonsourceibias.t68 gnd 0.176757f
C1445 commonsourceibias.n588 gnd 0.078584f
C1446 commonsourceibias.n589 gnd 0.084191f
C1447 commonsourceibias.n590 gnd 0.04027f
C1448 commonsourceibias.n591 gnd 0.009461f
C1449 commonsourceibias.n592 gnd 0.00769f
C1450 commonsourceibias.n593 gnd 0.013037f
C1451 commonsourceibias.n594 gnd 0.070526f
C1452 commonsourceibias.n595 gnd 0.013093f
C1453 commonsourceibias.n596 gnd 0.009461f
C1454 commonsourceibias.n597 gnd 0.009461f
C1455 commonsourceibias.n598 gnd 0.009461f
C1456 commonsourceibias.n599 gnd 0.009597f
C1457 commonsourceibias.n600 gnd 0.070526f
C1458 commonsourceibias.n601 gnd 0.011661f
C1459 commonsourceibias.n602 gnd 0.0129f
C1460 commonsourceibias.n603 gnd 0.009461f
C1461 commonsourceibias.n604 gnd 0.009461f
C1462 commonsourceibias.n605 gnd 0.012816f
C1463 commonsourceibias.n606 gnd 0.007653f
C1464 commonsourceibias.n607 gnd 0.012975f
C1465 commonsourceibias.n608 gnd 0.009461f
C1466 commonsourceibias.n609 gnd 0.009461f
C1467 commonsourceibias.n610 gnd 0.013054f
C1468 commonsourceibias.n611 gnd 0.011256f
C1469 commonsourceibias.n612 gnd 0.009134f
C1470 commonsourceibias.n613 gnd 0.009461f
C1471 commonsourceibias.n614 gnd 0.009461f
C1472 commonsourceibias.n615 gnd 0.011572f
C1473 commonsourceibias.n616 gnd 0.012989f
C1474 commonsourceibias.n617 gnd 0.070526f
C1475 commonsourceibias.n618 gnd 0.012901f
C1476 commonsourceibias.n619 gnd 0.009461f
C1477 commonsourceibias.n620 gnd 0.009461f
C1478 commonsourceibias.n621 gnd 0.009461f
C1479 commonsourceibias.n622 gnd 0.012901f
C1480 commonsourceibias.n623 gnd 0.070526f
C1481 commonsourceibias.n624 gnd 0.012989f
C1482 commonsourceibias.t100 gnd 0.176757f
C1483 commonsourceibias.n625 gnd 0.070526f
C1484 commonsourceibias.n626 gnd 0.011572f
C1485 commonsourceibias.n627 gnd 0.009461f
C1486 commonsourceibias.n628 gnd 0.009461f
C1487 commonsourceibias.n629 gnd 0.009461f
C1488 commonsourceibias.n630 gnd 0.011256f
C1489 commonsourceibias.n631 gnd 0.013054f
C1490 commonsourceibias.n632 gnd 0.070526f
C1491 commonsourceibias.n633 gnd 0.012975f
C1492 commonsourceibias.n634 gnd 0.009461f
C1493 commonsourceibias.n635 gnd 0.009461f
C1494 commonsourceibias.n636 gnd 0.009461f
C1495 commonsourceibias.n637 gnd 0.012816f
C1496 commonsourceibias.n638 gnd 0.070526f
C1497 commonsourceibias.n639 gnd 0.0129f
C1498 commonsourceibias.t154 gnd 0.176757f
C1499 commonsourceibias.n640 gnd 0.070526f
C1500 commonsourceibias.n641 gnd 0.011661f
C1501 commonsourceibias.n642 gnd 0.009461f
C1502 commonsourceibias.n643 gnd 0.009461f
C1503 commonsourceibias.n644 gnd 0.009461f
C1504 commonsourceibias.n645 gnd 0.010754f
C1505 commonsourceibias.n646 gnd 0.013093f
C1506 commonsourceibias.n647 gnd 0.070526f
C1507 commonsourceibias.n648 gnd 0.013037f
C1508 commonsourceibias.n649 gnd 0.009461f
C1509 commonsourceibias.n650 gnd 0.009461f
C1510 commonsourceibias.n651 gnd 0.009461f
C1511 commonsourceibias.n652 gnd 0.012717f
C1512 commonsourceibias.n653 gnd 0.070526f
C1513 commonsourceibias.n654 gnd 0.012748f
C1514 commonsourceibias.t151 gnd 0.191163f
C1515 commonsourceibias.n655 gnd 0.085044f
C1516 commonsourceibias.n656 gnd 0.030348f
C1517 commonsourceibias.n657 gnd 0.15151f
C1518 commonsourceibias.n658 gnd 0.012624f
C1519 commonsourceibias.t107 gnd 0.176757f
C1520 commonsourceibias.n659 gnd 0.00769f
C1521 commonsourceibias.n660 gnd 0.009461f
C1522 commonsourceibias.t122 gnd 0.176757f
C1523 commonsourceibias.n661 gnd 0.009597f
C1524 commonsourceibias.n662 gnd 0.009461f
C1525 commonsourceibias.t101 gnd 0.176757f
C1526 commonsourceibias.n663 gnd 0.007653f
C1527 commonsourceibias.n664 gnd 0.009461f
C1528 commonsourceibias.t115 gnd 0.176757f
C1529 commonsourceibias.n665 gnd 0.009134f
C1530 commonsourceibias.n666 gnd 0.009461f
C1531 commonsourceibias.t81 gnd 0.176757f
C1532 commonsourceibias.n667 gnd 0.007641f
C1533 commonsourceibias.n668 gnd 0.009461f
C1534 commonsourceibias.t70 gnd 0.176757f
C1535 commonsourceibias.t103 gnd 0.176757f
C1536 commonsourceibias.n669 gnd 0.070526f
C1537 commonsourceibias.n670 gnd 0.009461f
C1538 commonsourceibias.t132 gnd 0.176757f
C1539 commonsourceibias.n671 gnd 0.070526f
C1540 commonsourceibias.n672 gnd 0.009461f
C1541 commonsourceibias.t153 gnd 0.176757f
C1542 commonsourceibias.n673 gnd 0.070526f
C1543 commonsourceibias.n674 gnd 0.009461f
C1544 commonsourceibias.t87 gnd 0.176757f
C1545 commonsourceibias.n675 gnd 0.010754f
C1546 commonsourceibias.n676 gnd 0.009461f
C1547 commonsourceibias.t109 gnd 0.176757f
C1548 commonsourceibias.n677 gnd 0.012717f
C1549 commonsourceibias.t74 gnd 0.196904f
C1550 commonsourceibias.t145 gnd 0.176757f
C1551 commonsourceibias.n678 gnd 0.078584f
C1552 commonsourceibias.n679 gnd 0.084191f
C1553 commonsourceibias.n680 gnd 0.04027f
C1554 commonsourceibias.n681 gnd 0.009461f
C1555 commonsourceibias.n682 gnd 0.00769f
C1556 commonsourceibias.n683 gnd 0.013037f
C1557 commonsourceibias.n684 gnd 0.070526f
C1558 commonsourceibias.n685 gnd 0.013093f
C1559 commonsourceibias.n686 gnd 0.009461f
C1560 commonsourceibias.n687 gnd 0.009461f
C1561 commonsourceibias.n688 gnd 0.009461f
C1562 commonsourceibias.n689 gnd 0.009597f
C1563 commonsourceibias.n690 gnd 0.070526f
C1564 commonsourceibias.n691 gnd 0.011661f
C1565 commonsourceibias.n692 gnd 0.0129f
C1566 commonsourceibias.n693 gnd 0.009461f
C1567 commonsourceibias.n694 gnd 0.009461f
C1568 commonsourceibias.n695 gnd 0.012816f
C1569 commonsourceibias.n696 gnd 0.007653f
C1570 commonsourceibias.n697 gnd 0.012975f
C1571 commonsourceibias.n698 gnd 0.009461f
C1572 commonsourceibias.n699 gnd 0.009461f
C1573 commonsourceibias.n700 gnd 0.013054f
C1574 commonsourceibias.n701 gnd 0.011256f
C1575 commonsourceibias.n702 gnd 0.009134f
C1576 commonsourceibias.n703 gnd 0.009461f
C1577 commonsourceibias.n704 gnd 0.009461f
C1578 commonsourceibias.n705 gnd 0.011572f
C1579 commonsourceibias.n706 gnd 0.012989f
C1580 commonsourceibias.n707 gnd 0.070526f
C1581 commonsourceibias.n708 gnd 0.012901f
C1582 commonsourceibias.n709 gnd 0.009461f
C1583 commonsourceibias.n710 gnd 0.009461f
C1584 commonsourceibias.n711 gnd 0.009461f
C1585 commonsourceibias.n712 gnd 0.012901f
C1586 commonsourceibias.n713 gnd 0.070526f
C1587 commonsourceibias.n714 gnd 0.012989f
C1588 commonsourceibias.t110 gnd 0.176757f
C1589 commonsourceibias.n715 gnd 0.070526f
C1590 commonsourceibias.n716 gnd 0.011572f
C1591 commonsourceibias.n717 gnd 0.009461f
C1592 commonsourceibias.n718 gnd 0.009461f
C1593 commonsourceibias.n719 gnd 0.009461f
C1594 commonsourceibias.n720 gnd 0.011256f
C1595 commonsourceibias.n721 gnd 0.013054f
C1596 commonsourceibias.n722 gnd 0.070526f
C1597 commonsourceibias.n723 gnd 0.012975f
C1598 commonsourceibias.n724 gnd 0.009461f
C1599 commonsourceibias.n725 gnd 0.009461f
C1600 commonsourceibias.n726 gnd 0.009461f
C1601 commonsourceibias.n727 gnd 0.012816f
C1602 commonsourceibias.n728 gnd 0.070526f
C1603 commonsourceibias.n729 gnd 0.0129f
C1604 commonsourceibias.t135 gnd 0.176757f
C1605 commonsourceibias.n730 gnd 0.070526f
C1606 commonsourceibias.n731 gnd 0.011661f
C1607 commonsourceibias.n732 gnd 0.009461f
C1608 commonsourceibias.n733 gnd 0.009461f
C1609 commonsourceibias.n734 gnd 0.009461f
C1610 commonsourceibias.n735 gnd 0.010754f
C1611 commonsourceibias.n736 gnd 0.013093f
C1612 commonsourceibias.n737 gnd 0.070526f
C1613 commonsourceibias.n738 gnd 0.013037f
C1614 commonsourceibias.n739 gnd 0.009461f
C1615 commonsourceibias.n740 gnd 0.009461f
C1616 commonsourceibias.n741 gnd 0.009461f
C1617 commonsourceibias.n742 gnd 0.012717f
C1618 commonsourceibias.n743 gnd 0.070526f
C1619 commonsourceibias.n744 gnd 0.012748f
C1620 commonsourceibias.t82 gnd 0.191163f
C1621 commonsourceibias.n745 gnd 0.085044f
C1622 commonsourceibias.n746 gnd 0.030348f
C1623 commonsourceibias.n747 gnd 0.199656f
C1624 commonsourceibias.n748 gnd 5.01419f
C1625 a_n2140_13878.t11 gnd 0.186868f
C1626 a_n2140_13878.t10 gnd 0.186868f
C1627 a_n2140_13878.t5 gnd 0.186868f
C1628 a_n2140_13878.n0 gnd 1.47299f
C1629 a_n2140_13878.t2 gnd 0.186868f
C1630 a_n2140_13878.t4 gnd 0.186868f
C1631 a_n2140_13878.n1 gnd 1.47143f
C1632 a_n2140_13878.n2 gnd 2.05603f
C1633 a_n2140_13878.t12 gnd 0.186868f
C1634 a_n2140_13878.t3 gnd 0.186868f
C1635 a_n2140_13878.n3 gnd 1.47143f
C1636 a_n2140_13878.n4 gnd 1.00289f
C1637 a_n2140_13878.t9 gnd 0.186868f
C1638 a_n2140_13878.t1 gnd 0.186868f
C1639 a_n2140_13878.n5 gnd 1.47143f
C1640 a_n2140_13878.n6 gnd 4.06212f
C1641 a_n2140_13878.t17 gnd 1.74974f
C1642 a_n2140_13878.t20 gnd 0.186868f
C1643 a_n2140_13878.t21 gnd 0.186868f
C1644 a_n2140_13878.n7 gnd 1.3163f
C1645 a_n2140_13878.n8 gnd 1.47077f
C1646 a_n2140_13878.t16 gnd 1.74626f
C1647 a_n2140_13878.n9 gnd 0.740113f
C1648 a_n2140_13878.t19 gnd 1.74626f
C1649 a_n2140_13878.n10 gnd 0.740113f
C1650 a_n2140_13878.t22 gnd 0.186868f
C1651 a_n2140_13878.t23 gnd 0.186868f
C1652 a_n2140_13878.n11 gnd 1.3163f
C1653 a_n2140_13878.n12 gnd 0.74728f
C1654 a_n2140_13878.t18 gnd 1.74626f
C1655 a_n2140_13878.n13 gnd 2.09583f
C1656 a_n2140_13878.n14 gnd 2.85974f
C1657 a_n2140_13878.t6 gnd 0.186868f
C1658 a_n2140_13878.t7 gnd 0.186868f
C1659 a_n2140_13878.n15 gnd 1.47142f
C1660 a_n2140_13878.n16 gnd 2.01665f
C1661 a_n2140_13878.t13 gnd 0.186868f
C1662 a_n2140_13878.t14 gnd 0.186868f
C1663 a_n2140_13878.n17 gnd 1.47143f
C1664 a_n2140_13878.n18 gnd 0.651951f
C1665 a_n2140_13878.t0 gnd 0.186868f
C1666 a_n2140_13878.t8 gnd 0.186868f
C1667 a_n2140_13878.n19 gnd 1.47143f
C1668 a_n2140_13878.n20 gnd 1.32263f
C1669 a_n2140_13878.n21 gnd 1.47386f
C1670 a_n2140_13878.t15 gnd 0.186868f
C1671 a_n2318_13878.n0 gnd 2.73227f
C1672 a_n2318_13878.n1 gnd 3.94723f
C1673 a_n2318_13878.n2 gnd 3.81658f
C1674 a_n2318_13878.n3 gnd 0.652811f
C1675 a_n2318_13878.n4 gnd 0.210856f
C1676 a_n2318_13878.n5 gnd 0.210856f
C1677 a_n2318_13878.n6 gnd 0.729399f
C1678 a_n2318_13878.n7 gnd 0.210856f
C1679 a_n2318_13878.n8 gnd 0.433021f
C1680 a_n2318_13878.n9 gnd 0.652788f
C1681 a_n2318_13878.n10 gnd 0.200068f
C1682 a_n2318_13878.n11 gnd 0.147354f
C1683 a_n2318_13878.n12 gnd 0.231593f
C1684 a_n2318_13878.n13 gnd 0.178879f
C1685 a_n2318_13878.n14 gnd 0.200068f
C1686 a_n2318_13878.n15 gnd 1.09189f
C1687 a_n2318_13878.n16 gnd 0.147354f
C1688 a_n2318_13878.n17 gnd 0.705502f
C1689 a_n2318_13878.n18 gnd 0.50033f
C1690 a_n2318_13878.n19 gnd 0.210856f
C1691 a_n2318_13878.n20 gnd 0.210856f
C1692 a_n2318_13878.n21 gnd 0.433358f
C1693 a_n2318_13878.n22 gnd 0.210856f
C1694 a_n2318_13878.n23 gnd 0.210856f
C1695 a_n2318_13878.n24 gnd 1.73596f
C1696 a_n2318_13878.n25 gnd 2.03016f
C1697 a_n2318_13878.n26 gnd 1.73596f
C1698 a_n2318_13878.n27 gnd 1.85287f
C1699 a_n2318_13878.n28 gnd 3.14412f
C1700 a_n2318_13878.n29 gnd 0.278541f
C1701 a_n2318_13878.n30 gnd 0.742063f
C1702 a_n2318_13878.n31 gnd 0.004739f
C1703 a_n2318_13878.n32 gnd 0.01025f
C1704 a_n2318_13878.n33 gnd 0.01025f
C1705 a_n2318_13878.n34 gnd 0.004739f
C1706 a_n2318_13878.n35 gnd 0.278541f
C1707 a_n2318_13878.n36 gnd 0.278541f
C1708 a_n2318_13878.n37 gnd 0.433358f
C1709 a_n2318_13878.n38 gnd 0.004739f
C1710 a_n2318_13878.n39 gnd 0.01025f
C1711 a_n2318_13878.n40 gnd 0.01025f
C1712 a_n2318_13878.n41 gnd 0.004739f
C1713 a_n2318_13878.n42 gnd 0.278541f
C1714 a_n2318_13878.n43 gnd 0.008164f
C1715 a_n2318_13878.n44 gnd 0.278541f
C1716 a_n2318_13878.n45 gnd 0.008164f
C1717 a_n2318_13878.n46 gnd 0.278541f
C1718 a_n2318_13878.n47 gnd 0.008164f
C1719 a_n2318_13878.n48 gnd 0.278541f
C1720 a_n2318_13878.n49 gnd 0.008164f
C1721 a_n2318_13878.n50 gnd 0.278541f
C1722 a_n2318_13878.n51 gnd 0.278541f
C1723 a_n2318_13878.n52 gnd 0.004739f
C1724 a_n2318_13878.n53 gnd 0.01025f
C1725 a_n2318_13878.n54 gnd 0.01025f
C1726 a_n2318_13878.n55 gnd 0.004739f
C1727 a_n2318_13878.n56 gnd 0.278541f
C1728 a_n2318_13878.n57 gnd 0.278541f
C1729 a_n2318_13878.n58 gnd 0.004739f
C1730 a_n2318_13878.n59 gnd 0.01025f
C1731 a_n2318_13878.n60 gnd 0.105428f
C1732 a_n2318_13878.n61 gnd 0.01025f
C1733 a_n2318_13878.n62 gnd 0.004739f
C1734 a_n2318_13878.n63 gnd 0.278541f
C1735 a_n2318_13878.t20 gnd 0.146252f
C1736 a_n2318_13878.t13 gnd 0.691694f
C1737 a_n2318_13878.t19 gnd 0.680295f
C1738 a_n2318_13878.t9 gnd 0.680295f
C1739 a_n2318_13878.n64 gnd 0.297177f
C1740 a_n2318_13878.t39 gnd 0.680295f
C1741 a_n2318_13878.t17 gnd 0.680295f
C1742 a_n2318_13878.t11 gnd 0.680295f
C1743 a_n2318_13878.n65 gnd 0.297177f
C1744 a_n2318_13878.t27 gnd 0.680295f
C1745 a_n2318_13878.t21 gnd 0.691694f
C1746 a_n2318_13878.t5 gnd 0.113752f
C1747 a_n2318_13878.t41 gnd 0.113752f
C1748 a_n2318_13878.n66 gnd 1.00811f
C1749 a_n2318_13878.t43 gnd 0.113752f
C1750 a_n2318_13878.t0 gnd 0.113752f
C1751 a_n2318_13878.n67 gnd 1.00515f
C1752 a_n2318_13878.t7 gnd 0.113752f
C1753 a_n2318_13878.t1 gnd 0.113752f
C1754 a_n2318_13878.n68 gnd 1.00811f
C1755 a_n2318_13878.t8 gnd 0.113752f
C1756 a_n2318_13878.t2 gnd 0.113752f
C1757 a_n2318_13878.n69 gnd 1.00515f
C1758 a_n2318_13878.t4 gnd 0.113752f
C1759 a_n2318_13878.t46 gnd 0.113752f
C1760 a_n2318_13878.n70 gnd 1.00515f
C1761 a_n2318_13878.t44 gnd 0.113752f
C1762 a_n2318_13878.t42 gnd 0.113752f
C1763 a_n2318_13878.n71 gnd 1.00515f
C1764 a_n2318_13878.t45 gnd 0.113752f
C1765 a_n2318_13878.t6 gnd 0.113752f
C1766 a_n2318_13878.n72 gnd 1.00811f
C1767 a_n2318_13878.t47 gnd 0.113752f
C1768 a_n2318_13878.t3 gnd 0.113752f
C1769 a_n2318_13878.n73 gnd 1.00515f
C1770 a_n2318_13878.t78 gnd 0.691694f
C1771 a_n2318_13878.t59 gnd 0.680295f
C1772 a_n2318_13878.t63 gnd 0.680295f
C1773 a_n2318_13878.n74 gnd 0.297177f
C1774 a_n2318_13878.t53 gnd 0.680295f
C1775 a_n2318_13878.t68 gnd 0.680295f
C1776 a_n2318_13878.t75 gnd 0.680295f
C1777 a_n2318_13878.n75 gnd 0.297177f
C1778 a_n2318_13878.t76 gnd 0.680295f
C1779 a_n2318_13878.t50 gnd 0.691694f
C1780 a_n2318_13878.t16 gnd 1.36943f
C1781 a_n2318_13878.t26 gnd 0.146252f
C1782 a_n2318_13878.t36 gnd 0.146252f
C1783 a_n2318_13878.n76 gnd 1.0302f
C1784 a_n2318_13878.t38 gnd 0.146252f
C1785 a_n2318_13878.t30 gnd 0.146252f
C1786 a_n2318_13878.n77 gnd 1.0302f
C1787 a_n2318_13878.t32 gnd 0.146252f
C1788 a_n2318_13878.t34 gnd 0.146252f
C1789 a_n2318_13878.n78 gnd 1.0302f
C1790 a_n2318_13878.t24 gnd 1.3667f
C1791 a_n2318_13878.t31 gnd 0.680295f
C1792 a_n2318_13878.n79 gnd 0.297177f
C1793 a_n2318_13878.t37 gnd 0.680295f
C1794 a_n2318_13878.t15 gnd 0.691694f
C1795 a_n2318_13878.t25 gnd 0.680295f
C1796 a_n2318_13878.t58 gnd 0.680295f
C1797 a_n2318_13878.n80 gnd 0.297177f
C1798 a_n2318_13878.t72 gnd 0.680295f
C1799 a_n2318_13878.t74 gnd 0.691694f
C1800 a_n2318_13878.t52 gnd 0.680295f
C1801 a_n2318_13878.n81 gnd 0.2996f
C1802 a_n2318_13878.t71 gnd 0.680295f
C1803 a_n2318_13878.n82 gnd 0.297177f
C1804 a_n2318_13878.n83 gnd 0.292702f
C1805 a_n2318_13878.t49 gnd 0.680295f
C1806 a_n2318_13878.n84 gnd 0.292702f
C1807 a_n2318_13878.t66 gnd 0.680295f
C1808 a_n2318_13878.n85 gnd 0.2996f
C1809 a_n2318_13878.t51 gnd 0.691694f
C1810 a_n2318_13878.n86 gnd 0.2996f
C1811 a_n2318_13878.t35 gnd 0.680295f
C1812 a_n2318_13878.n87 gnd 0.297177f
C1813 a_n2318_13878.n88 gnd 0.292702f
C1814 a_n2318_13878.t29 gnd 0.680295f
C1815 a_n2318_13878.n89 gnd 0.292702f
C1816 a_n2318_13878.t33 gnd 0.680295f
C1817 a_n2318_13878.n90 gnd 0.2996f
C1818 a_n2318_13878.t23 gnd 0.691694f
C1819 a_n2318_13878.n91 gnd 1.17031f
C1820 a_n2318_13878.t56 gnd 0.680295f
C1821 a_n2318_13878.n92 gnd 0.295302f
C1822 a_n2318_13878.t62 gnd 0.680295f
C1823 a_n2318_13878.n93 gnd 0.295302f
C1824 a_n2318_13878.t54 gnd 0.680295f
C1825 a_n2318_13878.n94 gnd 0.295302f
C1826 a_n2318_13878.t67 gnd 0.680295f
C1827 a_n2318_13878.n95 gnd 0.295302f
C1828 a_n2318_13878.t57 gnd 0.680295f
C1829 a_n2318_13878.n96 gnd 0.28994f
C1830 a_n2318_13878.t79 gnd 0.680295f
C1831 a_n2318_13878.n97 gnd 0.299101f
C1832 a_n2318_13878.t60 gnd 0.691694f
C1833 a_n2318_13878.t69 gnd 0.680295f
C1834 a_n2318_13878.n98 gnd 0.28994f
C1835 a_n2318_13878.t55 gnd 0.680295f
C1836 a_n2318_13878.n99 gnd 0.299101f
C1837 a_n2318_13878.t64 gnd 0.691694f
C1838 a_n2318_13878.t73 gnd 0.680295f
C1839 a_n2318_13878.n100 gnd 0.28994f
C1840 a_n2318_13878.t61 gnd 0.680295f
C1841 a_n2318_13878.n101 gnd 0.299101f
C1842 a_n2318_13878.t77 gnd 0.691694f
C1843 a_n2318_13878.t65 gnd 0.680295f
C1844 a_n2318_13878.n102 gnd 0.28994f
C1845 a_n2318_13878.t48 gnd 0.680295f
C1846 a_n2318_13878.n103 gnd 0.299101f
C1847 a_n2318_13878.t70 gnd 0.691694f
C1848 a_n2318_13878.n104 gnd 1.41607f
C1849 a_n2318_13878.n105 gnd 0.2996f
C1850 a_n2318_13878.n106 gnd 0.292702f
C1851 a_n2318_13878.n107 gnd 0.292702f
C1852 a_n2318_13878.n108 gnd 0.2996f
C1853 a_n2318_13878.n109 gnd 0.2996f
C1854 a_n2318_13878.n110 gnd 0.292702f
C1855 a_n2318_13878.n111 gnd 0.292702f
C1856 a_n2318_13878.n112 gnd 0.2996f
C1857 a_n2318_13878.n113 gnd 0.839379f
C1858 a_n2318_13878.t14 gnd 1.36671f
C1859 a_n2318_13878.t22 gnd 1.36943f
C1860 a_n2318_13878.t12 gnd 0.146252f
C1861 a_n2318_13878.t28 gnd 0.146252f
C1862 a_n2318_13878.n114 gnd 1.0302f
C1863 a_n2318_13878.t40 gnd 0.146252f
C1864 a_n2318_13878.t18 gnd 0.146252f
C1865 a_n2318_13878.n115 gnd 1.0302f
C1866 a_n2318_13878.n116 gnd 1.0302f
C1867 a_n2318_13878.t10 gnd 0.146252f
C1868 CSoutput.n0 gnd 0.049217f
C1869 CSoutput.t222 gnd 0.325563f
C1870 CSoutput.n1 gnd 0.147008f
C1871 CSoutput.n2 gnd 0.049217f
C1872 CSoutput.t229 gnd 0.325563f
C1873 CSoutput.n3 gnd 0.039009f
C1874 CSoutput.n4 gnd 0.049217f
C1875 CSoutput.t236 gnd 0.325563f
C1876 CSoutput.n5 gnd 0.033638f
C1877 CSoutput.n6 gnd 0.049217f
C1878 CSoutput.t227 gnd 0.325563f
C1879 CSoutput.t225 gnd 0.325563f
C1880 CSoutput.n7 gnd 0.145406f
C1881 CSoutput.n8 gnd 0.049217f
C1882 CSoutput.t234 gnd 0.325563f
C1883 CSoutput.n9 gnd 0.032072f
C1884 CSoutput.n10 gnd 0.049217f
C1885 CSoutput.t217 gnd 0.325563f
C1886 CSoutput.t221 gnd 0.325563f
C1887 CSoutput.n11 gnd 0.145406f
C1888 CSoutput.n12 gnd 0.049217f
C1889 CSoutput.t232 gnd 0.325563f
C1890 CSoutput.n13 gnd 0.033638f
C1891 CSoutput.n14 gnd 0.049217f
C1892 CSoutput.t231 gnd 0.325563f
C1893 CSoutput.t219 gnd 0.325563f
C1894 CSoutput.n15 gnd 0.145406f
C1895 CSoutput.n16 gnd 0.049217f
C1896 CSoutput.t224 gnd 0.325563f
C1897 CSoutput.n17 gnd 0.035927f
C1898 CSoutput.t233 gnd 0.389056f
C1899 CSoutput.t230 gnd 0.325563f
C1900 CSoutput.n18 gnd 0.185627f
C1901 CSoutput.n19 gnd 0.180122f
C1902 CSoutput.n20 gnd 0.208963f
C1903 CSoutput.n21 gnd 0.049217f
C1904 CSoutput.n22 gnd 0.041077f
C1905 CSoutput.n23 gnd 0.145406f
C1906 CSoutput.n24 gnd 0.039597f
C1907 CSoutput.n25 gnd 0.039009f
C1908 CSoutput.n26 gnd 0.049217f
C1909 CSoutput.n27 gnd 0.049217f
C1910 CSoutput.n28 gnd 0.040762f
C1911 CSoutput.n29 gnd 0.034608f
C1912 CSoutput.n30 gnd 0.148643f
C1913 CSoutput.n31 gnd 0.035084f
C1914 CSoutput.n32 gnd 0.049217f
C1915 CSoutput.n33 gnd 0.049217f
C1916 CSoutput.n34 gnd 0.049217f
C1917 CSoutput.n35 gnd 0.040328f
C1918 CSoutput.n36 gnd 0.145406f
C1919 CSoutput.n37 gnd 0.038567f
C1920 CSoutput.n38 gnd 0.040039f
C1921 CSoutput.n39 gnd 0.049217f
C1922 CSoutput.n40 gnd 0.049217f
C1923 CSoutput.n41 gnd 0.041069f
C1924 CSoutput.n42 gnd 0.037537f
C1925 CSoutput.n43 gnd 0.145406f
C1926 CSoutput.n44 gnd 0.038489f
C1927 CSoutput.n45 gnd 0.049217f
C1928 CSoutput.n46 gnd 0.049217f
C1929 CSoutput.n47 gnd 0.049217f
C1930 CSoutput.n48 gnd 0.038489f
C1931 CSoutput.n49 gnd 0.145406f
C1932 CSoutput.n50 gnd 0.037537f
C1933 CSoutput.n51 gnd 0.041069f
C1934 CSoutput.n52 gnd 0.049217f
C1935 CSoutput.n53 gnd 0.049217f
C1936 CSoutput.n54 gnd 0.040039f
C1937 CSoutput.n55 gnd 0.038567f
C1938 CSoutput.n56 gnd 0.145406f
C1939 CSoutput.n57 gnd 0.040328f
C1940 CSoutput.n58 gnd 0.049217f
C1941 CSoutput.n59 gnd 0.049217f
C1942 CSoutput.n60 gnd 0.049217f
C1943 CSoutput.n61 gnd 0.035084f
C1944 CSoutput.n62 gnd 0.148643f
C1945 CSoutput.n63 gnd 0.034608f
C1946 CSoutput.t228 gnd 0.325563f
C1947 CSoutput.n64 gnd 0.145406f
C1948 CSoutput.n65 gnd 0.040762f
C1949 CSoutput.n66 gnd 0.049217f
C1950 CSoutput.n67 gnd 0.049217f
C1951 CSoutput.n68 gnd 0.049217f
C1952 CSoutput.n69 gnd 0.039597f
C1953 CSoutput.n70 gnd 0.145406f
C1954 CSoutput.n71 gnd 0.041077f
C1955 CSoutput.n72 gnd 0.035927f
C1956 CSoutput.n73 gnd 0.049217f
C1957 CSoutput.n74 gnd 0.049217f
C1958 CSoutput.n75 gnd 0.037258f
C1959 CSoutput.n76 gnd 0.022128f
C1960 CSoutput.t235 gnd 0.365793f
C1961 CSoutput.n77 gnd 0.181711f
C1962 CSoutput.n78 gnd 0.743372f
C1963 CSoutput.t159 gnd 0.061392f
C1964 CSoutput.t90 gnd 0.061392f
C1965 CSoutput.n79 gnd 0.475316f
C1966 CSoutput.t174 gnd 0.061392f
C1967 CSoutput.t112 gnd 0.061392f
C1968 CSoutput.n80 gnd 0.474469f
C1969 CSoutput.n81 gnd 0.481585f
C1970 CSoutput.t69 gnd 0.061392f
C1971 CSoutput.t129 gnd 0.061392f
C1972 CSoutput.n82 gnd 0.474469f
C1973 CSoutput.n83 gnd 0.237305f
C1974 CSoutput.t75 gnd 0.061392f
C1975 CSoutput.t103 gnd 0.061392f
C1976 CSoutput.n84 gnd 0.474469f
C1977 CSoutput.n85 gnd 0.237305f
C1978 CSoutput.t179 gnd 0.061392f
C1979 CSoutput.t122 gnd 0.061392f
C1980 CSoutput.n86 gnd 0.474469f
C1981 CSoutput.n87 gnd 0.237305f
C1982 CSoutput.t78 gnd 0.061392f
C1983 CSoutput.t163 gnd 0.061392f
C1984 CSoutput.n88 gnd 0.474469f
C1985 CSoutput.n89 gnd 0.237305f
C1986 CSoutput.t86 gnd 0.061392f
C1987 CSoutput.t139 gnd 0.061392f
C1988 CSoutput.n90 gnd 0.474469f
C1989 CSoutput.n91 gnd 0.237305f
C1990 CSoutput.t107 gnd 0.061392f
C1991 CSoutput.t130 gnd 0.061392f
C1992 CSoutput.n92 gnd 0.474469f
C1993 CSoutput.n93 gnd 0.237305f
C1994 CSoutput.t125 gnd 0.061392f
C1995 CSoutput.t168 gnd 0.061392f
C1996 CSoutput.n94 gnd 0.474469f
C1997 CSoutput.n95 gnd 0.237305f
C1998 CSoutput.t95 gnd 0.061392f
C1999 CSoutput.t146 gnd 0.061392f
C2000 CSoutput.n96 gnd 0.474469f
C2001 CSoutput.n97 gnd 0.435162f
C2002 CSoutput.t65 gnd 0.061392f
C2003 CSoutput.t157 gnd 0.061392f
C2004 CSoutput.n98 gnd 0.475316f
C2005 CSoutput.t140 gnd 0.061392f
C2006 CSoutput.t116 gnd 0.061392f
C2007 CSoutput.n99 gnd 0.474469f
C2008 CSoutput.n100 gnd 0.481585f
C2009 CSoutput.t91 gnd 0.061392f
C2010 CSoutput.t170 gnd 0.061392f
C2011 CSoutput.n101 gnd 0.474469f
C2012 CSoutput.n102 gnd 0.237305f
C2013 CSoutput.t137 gnd 0.061392f
C2014 CSoutput.t136 gnd 0.061392f
C2015 CSoutput.n103 gnd 0.474469f
C2016 CSoutput.n104 gnd 0.237305f
C2017 CSoutput.t126 gnd 0.061392f
C2018 CSoutput.t87 gnd 0.061392f
C2019 CSoutput.n105 gnd 0.474469f
C2020 CSoutput.n106 gnd 0.237305f
C2021 CSoutput.t68 gnd 0.061392f
C2022 CSoutput.t127 gnd 0.061392f
C2023 CSoutput.n107 gnd 0.474469f
C2024 CSoutput.n108 gnd 0.237305f
C2025 CSoutput.t123 gnd 0.061392f
C2026 CSoutput.t85 gnd 0.061392f
C2027 CSoutput.n109 gnd 0.474469f
C2028 CSoutput.n110 gnd 0.237305f
C2029 CSoutput.t66 gnd 0.061392f
C2030 CSoutput.t63 gnd 0.061392f
C2031 CSoutput.n111 gnd 0.474469f
C2032 CSoutput.n112 gnd 0.237305f
C2033 CSoutput.t141 gnd 0.061392f
C2034 CSoutput.t104 gnd 0.061392f
C2035 CSoutput.n113 gnd 0.474469f
C2036 CSoutput.n114 gnd 0.237305f
C2037 CSoutput.t97 gnd 0.061392f
C2038 CSoutput.t61 gnd 0.061392f
C2039 CSoutput.n115 gnd 0.474469f
C2040 CSoutput.n116 gnd 0.353881f
C2041 CSoutput.n117 gnd 0.446242f
C2042 CSoutput.t81 gnd 0.061392f
C2043 CSoutput.t169 gnd 0.061392f
C2044 CSoutput.n118 gnd 0.475316f
C2045 CSoutput.t150 gnd 0.061392f
C2046 CSoutput.t128 gnd 0.061392f
C2047 CSoutput.n119 gnd 0.474469f
C2048 CSoutput.n120 gnd 0.481585f
C2049 CSoutput.t108 gnd 0.061392f
C2050 CSoutput.t180 gnd 0.061392f
C2051 CSoutput.n121 gnd 0.474469f
C2052 CSoutput.n122 gnd 0.237305f
C2053 CSoutput.t149 gnd 0.061392f
C2054 CSoutput.t148 gnd 0.061392f
C2055 CSoutput.n123 gnd 0.474469f
C2056 CSoutput.n124 gnd 0.237305f
C2057 CSoutput.t134 gnd 0.061392f
C2058 CSoutput.t105 gnd 0.061392f
C2059 CSoutput.n125 gnd 0.474469f
C2060 CSoutput.n126 gnd 0.237305f
C2061 CSoutput.t82 gnd 0.061392f
C2062 CSoutput.t135 gnd 0.061392f
C2063 CSoutput.n127 gnd 0.474469f
C2064 CSoutput.n128 gnd 0.237305f
C2065 CSoutput.t133 gnd 0.061392f
C2066 CSoutput.t102 gnd 0.061392f
C2067 CSoutput.n129 gnd 0.474469f
C2068 CSoutput.n130 gnd 0.237305f
C2069 CSoutput.t80 gnd 0.061392f
C2070 CSoutput.t79 gnd 0.061392f
C2071 CSoutput.n131 gnd 0.474469f
C2072 CSoutput.n132 gnd 0.237305f
C2073 CSoutput.t151 gnd 0.061392f
C2074 CSoutput.t118 gnd 0.061392f
C2075 CSoutput.n133 gnd 0.474469f
C2076 CSoutput.n134 gnd 0.237305f
C2077 CSoutput.t113 gnd 0.061392f
C2078 CSoutput.t74 gnd 0.061392f
C2079 CSoutput.n135 gnd 0.474469f
C2080 CSoutput.n136 gnd 0.353881f
C2081 CSoutput.n137 gnd 0.498784f
C2082 CSoutput.n138 gnd 9.29035f
C2083 CSoutput.n140 gnd 0.870649f
C2084 CSoutput.n141 gnd 0.652987f
C2085 CSoutput.n142 gnd 0.870649f
C2086 CSoutput.n143 gnd 0.870649f
C2087 CSoutput.n144 gnd 2.34405f
C2088 CSoutput.n145 gnd 0.870649f
C2089 CSoutput.n146 gnd 0.870649f
C2090 CSoutput.t223 gnd 1.08831f
C2091 CSoutput.n147 gnd 0.870649f
C2092 CSoutput.n148 gnd 0.870649f
C2093 CSoutput.n152 gnd 0.870649f
C2094 CSoutput.n156 gnd 0.870649f
C2095 CSoutput.n157 gnd 0.870649f
C2096 CSoutput.n159 gnd 0.870649f
C2097 CSoutput.n164 gnd 0.870649f
C2098 CSoutput.n166 gnd 0.870649f
C2099 CSoutput.n167 gnd 0.870649f
C2100 CSoutput.n169 gnd 0.870649f
C2101 CSoutput.n170 gnd 0.870649f
C2102 CSoutput.n172 gnd 0.870649f
C2103 CSoutput.t218 gnd 14.548401f
C2104 CSoutput.n174 gnd 0.870649f
C2105 CSoutput.n175 gnd 0.652987f
C2106 CSoutput.n176 gnd 0.870649f
C2107 CSoutput.n177 gnd 0.870649f
C2108 CSoutput.n178 gnd 2.34405f
C2109 CSoutput.n179 gnd 0.870649f
C2110 CSoutput.n180 gnd 0.870649f
C2111 CSoutput.t237 gnd 1.08831f
C2112 CSoutput.n181 gnd 0.870649f
C2113 CSoutput.n182 gnd 0.870649f
C2114 CSoutput.n186 gnd 0.870649f
C2115 CSoutput.n190 gnd 0.870649f
C2116 CSoutput.n191 gnd 0.870649f
C2117 CSoutput.n193 gnd 0.870649f
C2118 CSoutput.n198 gnd 0.870649f
C2119 CSoutput.n200 gnd 0.870649f
C2120 CSoutput.n201 gnd 0.870649f
C2121 CSoutput.n203 gnd 0.870649f
C2122 CSoutput.n204 gnd 0.870649f
C2123 CSoutput.n206 gnd 0.870649f
C2124 CSoutput.n207 gnd 0.652987f
C2125 CSoutput.n209 gnd 0.870649f
C2126 CSoutput.n210 gnd 0.652987f
C2127 CSoutput.n211 gnd 0.870649f
C2128 CSoutput.n212 gnd 0.870649f
C2129 CSoutput.n213 gnd 2.34405f
C2130 CSoutput.n214 gnd 0.870649f
C2131 CSoutput.n215 gnd 0.870649f
C2132 CSoutput.t216 gnd 1.08831f
C2133 CSoutput.n216 gnd 0.870649f
C2134 CSoutput.n217 gnd 2.34405f
C2135 CSoutput.n219 gnd 0.870649f
C2136 CSoutput.n220 gnd 0.870649f
C2137 CSoutput.n222 gnd 0.870649f
C2138 CSoutput.n223 gnd 0.870649f
C2139 CSoutput.t226 gnd 14.311299f
C2140 CSoutput.t220 gnd 14.548401f
C2141 CSoutput.n229 gnd 2.73135f
C2142 CSoutput.n230 gnd 11.1265f
C2143 CSoutput.n231 gnd 11.5921f
C2144 CSoutput.n236 gnd 2.95879f
C2145 CSoutput.n242 gnd 0.870649f
C2146 CSoutput.n244 gnd 0.870649f
C2147 CSoutput.n246 gnd 0.870649f
C2148 CSoutput.n248 gnd 0.870649f
C2149 CSoutput.n250 gnd 0.870649f
C2150 CSoutput.n256 gnd 0.870649f
C2151 CSoutput.n263 gnd 1.59731f
C2152 CSoutput.n264 gnd 1.59731f
C2153 CSoutput.n265 gnd 0.870649f
C2154 CSoutput.n266 gnd 0.870649f
C2155 CSoutput.n268 gnd 0.652987f
C2156 CSoutput.n269 gnd 0.559224f
C2157 CSoutput.n271 gnd 0.652987f
C2158 CSoutput.n272 gnd 0.559224f
C2159 CSoutput.n273 gnd 0.652987f
C2160 CSoutput.n275 gnd 0.870649f
C2161 CSoutput.n277 gnd 2.34405f
C2162 CSoutput.n278 gnd 2.73135f
C2163 CSoutput.n279 gnd 10.2336f
C2164 CSoutput.n281 gnd 0.652987f
C2165 CSoutput.n282 gnd 1.68017f
C2166 CSoutput.n283 gnd 0.652987f
C2167 CSoutput.n285 gnd 0.870649f
C2168 CSoutput.n287 gnd 2.34405f
C2169 CSoutput.n288 gnd 5.10573f
C2170 CSoutput.t89 gnd 0.061392f
C2171 CSoutput.t158 gnd 0.061392f
C2172 CSoutput.n289 gnd 0.475316f
C2173 CSoutput.t111 gnd 0.061392f
C2174 CSoutput.t172 gnd 0.061392f
C2175 CSoutput.n290 gnd 0.474469f
C2176 CSoutput.n291 gnd 0.481585f
C2177 CSoutput.t152 gnd 0.061392f
C2178 CSoutput.t67 gnd 0.061392f
C2179 CSoutput.n292 gnd 0.474469f
C2180 CSoutput.n293 gnd 0.237305f
C2181 CSoutput.t101 gnd 0.061392f
C2182 CSoutput.t73 gnd 0.061392f
C2183 CSoutput.n294 gnd 0.474469f
C2184 CSoutput.n295 gnd 0.237305f
C2185 CSoutput.t121 gnd 0.061392f
C2186 CSoutput.t94 gnd 0.061392f
C2187 CSoutput.n296 gnd 0.474469f
C2188 CSoutput.n297 gnd 0.237305f
C2189 CSoutput.t162 gnd 0.061392f
C2190 CSoutput.t77 gnd 0.061392f
C2191 CSoutput.n298 gnd 0.474469f
C2192 CSoutput.n299 gnd 0.237305f
C2193 CSoutput.t138 gnd 0.061392f
C2194 CSoutput.t83 gnd 0.061392f
C2195 CSoutput.n300 gnd 0.474469f
C2196 CSoutput.n301 gnd 0.237305f
C2197 CSoutput.t154 gnd 0.061392f
C2198 CSoutput.t106 gnd 0.061392f
C2199 CSoutput.n302 gnd 0.474469f
C2200 CSoutput.n303 gnd 0.237305f
C2201 CSoutput.t167 gnd 0.061392f
C2202 CSoutput.t124 gnd 0.061392f
C2203 CSoutput.n304 gnd 0.474469f
C2204 CSoutput.n305 gnd 0.237305f
C2205 CSoutput.t145 gnd 0.061392f
C2206 CSoutput.t96 gnd 0.061392f
C2207 CSoutput.n306 gnd 0.474469f
C2208 CSoutput.n307 gnd 0.435162f
C2209 CSoutput.t120 gnd 0.061392f
C2210 CSoutput.t144 gnd 0.061392f
C2211 CSoutput.n308 gnd 0.475316f
C2212 CSoutput.t62 gnd 0.061392f
C2213 CSoutput.t99 gnd 0.061392f
C2214 CSoutput.n309 gnd 0.474469f
C2215 CSoutput.n310 gnd 0.481585f
C2216 CSoutput.t100 gnd 0.061392f
C2217 CSoutput.t166 gnd 0.061392f
C2218 CSoutput.n311 gnd 0.474469f
C2219 CSoutput.n312 gnd 0.237305f
C2220 CSoutput.t92 gnd 0.061392f
C2221 CSoutput.t93 gnd 0.061392f
C2222 CSoutput.n313 gnd 0.474469f
C2223 CSoutput.n314 gnd 0.237305f
C2224 CSoutput.t164 gnd 0.061392f
C2225 CSoutput.t165 gnd 0.061392f
C2226 CSoutput.n315 gnd 0.474469f
C2227 CSoutput.n316 gnd 0.237305f
C2228 CSoutput.t72 gnd 0.061392f
C2229 CSoutput.t147 gnd 0.061392f
C2230 CSoutput.n317 gnd 0.474469f
C2231 CSoutput.n318 gnd 0.237305f
C2232 CSoutput.t161 gnd 0.061392f
C2233 CSoutput.t70 gnd 0.061392f
C2234 CSoutput.n319 gnd 0.474469f
C2235 CSoutput.n320 gnd 0.237305f
C2236 CSoutput.t119 gnd 0.061392f
C2237 CSoutput.t143 gnd 0.061392f
C2238 CSoutput.n321 gnd 0.474469f
C2239 CSoutput.n322 gnd 0.237305f
C2240 CSoutput.t173 gnd 0.061392f
C2241 CSoutput.t98 gnd 0.061392f
C2242 CSoutput.n323 gnd 0.474469f
C2243 CSoutput.n324 gnd 0.237305f
C2244 CSoutput.t142 gnd 0.061392f
C2245 CSoutput.t178 gnd 0.061392f
C2246 CSoutput.n325 gnd 0.474469f
C2247 CSoutput.n326 gnd 0.353881f
C2248 CSoutput.n327 gnd 0.446242f
C2249 CSoutput.t131 gnd 0.061392f
C2250 CSoutput.t155 gnd 0.061392f
C2251 CSoutput.n328 gnd 0.475316f
C2252 CSoutput.t76 gnd 0.061392f
C2253 CSoutput.t114 gnd 0.061392f
C2254 CSoutput.n329 gnd 0.474469f
C2255 CSoutput.n330 gnd 0.481585f
C2256 CSoutput.t117 gnd 0.061392f
C2257 CSoutput.t177 gnd 0.061392f
C2258 CSoutput.n331 gnd 0.474469f
C2259 CSoutput.n332 gnd 0.237305f
C2260 CSoutput.t109 gnd 0.061392f
C2261 CSoutput.t110 gnd 0.061392f
C2262 CSoutput.n333 gnd 0.474469f
C2263 CSoutput.n334 gnd 0.237305f
C2264 CSoutput.t175 gnd 0.061392f
C2265 CSoutput.t176 gnd 0.061392f
C2266 CSoutput.n335 gnd 0.474469f
C2267 CSoutput.n336 gnd 0.237305f
C2268 CSoutput.t88 gnd 0.061392f
C2269 CSoutput.t160 gnd 0.061392f
C2270 CSoutput.n337 gnd 0.474469f
C2271 CSoutput.n338 gnd 0.237305f
C2272 CSoutput.t171 gnd 0.061392f
C2273 CSoutput.t84 gnd 0.061392f
C2274 CSoutput.n339 gnd 0.474469f
C2275 CSoutput.n340 gnd 0.237305f
C2276 CSoutput.t132 gnd 0.061392f
C2277 CSoutput.t156 gnd 0.061392f
C2278 CSoutput.n341 gnd 0.474469f
C2279 CSoutput.n342 gnd 0.237305f
C2280 CSoutput.t64 gnd 0.061392f
C2281 CSoutput.t115 gnd 0.061392f
C2282 CSoutput.n343 gnd 0.474469f
C2283 CSoutput.n344 gnd 0.237305f
C2284 CSoutput.t153 gnd 0.061392f
C2285 CSoutput.t71 gnd 0.061392f
C2286 CSoutput.n345 gnd 0.474467f
C2287 CSoutput.n346 gnd 0.353883f
C2288 CSoutput.n347 gnd 0.498784f
C2289 CSoutput.n348 gnd 13.267f
C2290 CSoutput.t53 gnd 0.053718f
C2291 CSoutput.t36 gnd 0.053718f
C2292 CSoutput.n349 gnd 0.476259f
C2293 CSoutput.t215 gnd 0.053718f
C2294 CSoutput.t182 gnd 0.053718f
C2295 CSoutput.n350 gnd 0.47467f
C2296 CSoutput.n351 gnd 0.442304f
C2297 CSoutput.t212 gnd 0.053718f
C2298 CSoutput.t198 gnd 0.053718f
C2299 CSoutput.n352 gnd 0.47467f
C2300 CSoutput.n353 gnd 0.218035f
C2301 CSoutput.t194 gnd 0.053718f
C2302 CSoutput.t13 gnd 0.053718f
C2303 CSoutput.n354 gnd 0.47467f
C2304 CSoutput.n355 gnd 0.218035f
C2305 CSoutput.t40 gnd 0.053718f
C2306 CSoutput.t187 gnd 0.053718f
C2307 CSoutput.n356 gnd 0.47467f
C2308 CSoutput.n357 gnd 0.218035f
C2309 CSoutput.t39 gnd 0.053718f
C2310 CSoutput.t37 gnd 0.053718f
C2311 CSoutput.n358 gnd 0.47467f
C2312 CSoutput.n359 gnd 0.218035f
C2313 CSoutput.t181 gnd 0.053718f
C2314 CSoutput.t197 gnd 0.053718f
C2315 CSoutput.n360 gnd 0.47467f
C2316 CSoutput.n361 gnd 0.218035f
C2317 CSoutput.t18 gnd 0.053718f
C2318 CSoutput.t59 gnd 0.053718f
C2319 CSoutput.n362 gnd 0.47467f
C2320 CSoutput.n363 gnd 0.402154f
C2321 CSoutput.t186 gnd 0.053718f
C2322 CSoutput.t23 gnd 0.053718f
C2323 CSoutput.n364 gnd 0.476259f
C2324 CSoutput.t14 gnd 0.053718f
C2325 CSoutput.t189 gnd 0.053718f
C2326 CSoutput.n365 gnd 0.47467f
C2327 CSoutput.n366 gnd 0.442304f
C2328 CSoutput.t16 gnd 0.053718f
C2329 CSoutput.t202 gnd 0.053718f
C2330 CSoutput.n367 gnd 0.47467f
C2331 CSoutput.n368 gnd 0.218035f
C2332 CSoutput.t188 gnd 0.053718f
C2333 CSoutput.t19 gnd 0.053718f
C2334 CSoutput.n369 gnd 0.47467f
C2335 CSoutput.n370 gnd 0.218035f
C2336 CSoutput.t191 gnd 0.053718f
C2337 CSoutput.t203 gnd 0.053718f
C2338 CSoutput.n371 gnd 0.47467f
C2339 CSoutput.n372 gnd 0.218035f
C2340 CSoutput.t11 gnd 0.053718f
C2341 CSoutput.t208 gnd 0.053718f
C2342 CSoutput.n373 gnd 0.47467f
C2343 CSoutput.n374 gnd 0.218035f
C2344 CSoutput.t17 gnd 0.053718f
C2345 CSoutput.t195 gnd 0.053718f
C2346 CSoutput.n375 gnd 0.47467f
C2347 CSoutput.n376 gnd 0.218035f
C2348 CSoutput.t209 gnd 0.053718f
C2349 CSoutput.t33 gnd 0.053718f
C2350 CSoutput.n377 gnd 0.47467f
C2351 CSoutput.n378 gnd 0.331024f
C2352 CSoutput.n379 gnd 0.417524f
C2353 CSoutput.t10 gnd 0.053718f
C2354 CSoutput.t207 gnd 0.053718f
C2355 CSoutput.n380 gnd 0.476259f
C2356 CSoutput.t204 gnd 0.053718f
C2357 CSoutput.t9 gnd 0.053718f
C2358 CSoutput.n381 gnd 0.47467f
C2359 CSoutput.n382 gnd 0.442304f
C2360 CSoutput.t2 gnd 0.053718f
C2361 CSoutput.t31 gnd 0.053718f
C2362 CSoutput.n383 gnd 0.47467f
C2363 CSoutput.n384 gnd 0.218035f
C2364 CSoutput.t214 gnd 0.053718f
C2365 CSoutput.t1 gnd 0.053718f
C2366 CSoutput.n385 gnd 0.47467f
C2367 CSoutput.n386 gnd 0.218035f
C2368 CSoutput.t45 gnd 0.053718f
C2369 CSoutput.t183 gnd 0.053718f
C2370 CSoutput.n387 gnd 0.47467f
C2371 CSoutput.n388 gnd 0.218035f
C2372 CSoutput.t44 gnd 0.053718f
C2373 CSoutput.t199 gnd 0.053718f
C2374 CSoutput.n389 gnd 0.47467f
C2375 CSoutput.n390 gnd 0.218035f
C2376 CSoutput.t21 gnd 0.053718f
C2377 CSoutput.t190 gnd 0.053718f
C2378 CSoutput.n391 gnd 0.47467f
C2379 CSoutput.n392 gnd 0.218035f
C2380 CSoutput.t8 gnd 0.053718f
C2381 CSoutput.t55 gnd 0.053718f
C2382 CSoutput.n393 gnd 0.47467f
C2383 CSoutput.n394 gnd 0.331024f
C2384 CSoutput.n395 gnd 0.448355f
C2385 CSoutput.n396 gnd 13.4517f
C2386 CSoutput.t200 gnd 0.053718f
C2387 CSoutput.t32 gnd 0.053718f
C2388 CSoutput.n397 gnd 0.476259f
C2389 CSoutput.t192 gnd 0.053718f
C2390 CSoutput.t6 gnd 0.053718f
C2391 CSoutput.n398 gnd 0.47467f
C2392 CSoutput.n399 gnd 0.442304f
C2393 CSoutput.t3 gnd 0.053718f
C2394 CSoutput.t27 gnd 0.053718f
C2395 CSoutput.n400 gnd 0.47467f
C2396 CSoutput.n401 gnd 0.218035f
C2397 CSoutput.t5 gnd 0.053718f
C2398 CSoutput.t47 gnd 0.053718f
C2399 CSoutput.n402 gnd 0.47467f
C2400 CSoutput.n403 gnd 0.218035f
C2401 CSoutput.t28 gnd 0.053718f
C2402 CSoutput.t4 gnd 0.053718f
C2403 CSoutput.n404 gnd 0.47467f
C2404 CSoutput.n405 gnd 0.218035f
C2405 CSoutput.t0 gnd 0.053718f
C2406 CSoutput.t57 gnd 0.053718f
C2407 CSoutput.n406 gnd 0.47467f
C2408 CSoutput.n407 gnd 0.218035f
C2409 CSoutput.t201 gnd 0.053718f
C2410 CSoutput.t20 gnd 0.053718f
C2411 CSoutput.n408 gnd 0.47467f
C2412 CSoutput.n409 gnd 0.218035f
C2413 CSoutput.t196 gnd 0.053718f
C2414 CSoutput.t60 gnd 0.053718f
C2415 CSoutput.n410 gnd 0.47467f
C2416 CSoutput.n411 gnd 0.402154f
C2417 CSoutput.t41 gnd 0.053718f
C2418 CSoutput.t15 gnd 0.053718f
C2419 CSoutput.n412 gnd 0.476259f
C2420 CSoutput.t205 gnd 0.053718f
C2421 CSoutput.t35 gnd 0.053718f
C2422 CSoutput.n413 gnd 0.47467f
C2423 CSoutput.n414 gnd 0.442304f
C2424 CSoutput.t184 gnd 0.053718f
C2425 CSoutput.t25 gnd 0.053718f
C2426 CSoutput.n415 gnd 0.47467f
C2427 CSoutput.n416 gnd 0.218035f
C2428 CSoutput.t12 gnd 0.053718f
C2429 CSoutput.t24 gnd 0.053718f
C2430 CSoutput.n417 gnd 0.47467f
C2431 CSoutput.n418 gnd 0.218035f
C2432 CSoutput.t38 gnd 0.053718f
C2433 CSoutput.t46 gnd 0.053718f
C2434 CSoutput.n419 gnd 0.47467f
C2435 CSoutput.n420 gnd 0.218035f
C2436 CSoutput.t30 gnd 0.053718f
C2437 CSoutput.t48 gnd 0.053718f
C2438 CSoutput.n421 gnd 0.47467f
C2439 CSoutput.n422 gnd 0.218035f
C2440 CSoutput.t50 gnd 0.053718f
C2441 CSoutput.t54 gnd 0.053718f
C2442 CSoutput.n423 gnd 0.47467f
C2443 CSoutput.n424 gnd 0.218035f
C2444 CSoutput.t193 gnd 0.053718f
C2445 CSoutput.t29 gnd 0.053718f
C2446 CSoutput.n425 gnd 0.47467f
C2447 CSoutput.n426 gnd 0.331024f
C2448 CSoutput.n427 gnd 0.417524f
C2449 CSoutput.t211 gnd 0.053718f
C2450 CSoutput.t56 gnd 0.053718f
C2451 CSoutput.n428 gnd 0.476259f
C2452 CSoutput.t43 gnd 0.053718f
C2453 CSoutput.t34 gnd 0.053718f
C2454 CSoutput.n429 gnd 0.47467f
C2455 CSoutput.n430 gnd 0.442304f
C2456 CSoutput.t7 gnd 0.053718f
C2457 CSoutput.t210 gnd 0.053718f
C2458 CSoutput.n431 gnd 0.47467f
C2459 CSoutput.n432 gnd 0.218035f
C2460 CSoutput.t49 gnd 0.053718f
C2461 CSoutput.t42 gnd 0.053718f
C2462 CSoutput.n433 gnd 0.47467f
C2463 CSoutput.n434 gnd 0.218035f
C2464 CSoutput.t52 gnd 0.053718f
C2465 CSoutput.t185 gnd 0.053718f
C2466 CSoutput.n435 gnd 0.47467f
C2467 CSoutput.n436 gnd 0.218035f
C2468 CSoutput.t22 gnd 0.053718f
C2469 CSoutput.t26 gnd 0.053718f
C2470 CSoutput.n437 gnd 0.47467f
C2471 CSoutput.n438 gnd 0.218035f
C2472 CSoutput.t58 gnd 0.053718f
C2473 CSoutput.t51 gnd 0.053718f
C2474 CSoutput.n439 gnd 0.47467f
C2475 CSoutput.n440 gnd 0.218035f
C2476 CSoutput.t206 gnd 0.053718f
C2477 CSoutput.t213 gnd 0.053718f
C2478 CSoutput.n441 gnd 0.47467f
C2479 CSoutput.n442 gnd 0.331024f
C2480 CSoutput.n443 gnd 0.448355f
C2481 CSoutput.n444 gnd 7.82108f
C2482 CSoutput.n445 gnd 14.872f
C2483 vdd.t6 gnd 0.039365f
C2484 vdd.t13 gnd 0.039365f
C2485 vdd.n0 gnd 0.310475f
C2486 vdd.t48 gnd 0.039365f
C2487 vdd.t1 gnd 0.039365f
C2488 vdd.n1 gnd 0.309963f
C2489 vdd.n2 gnd 0.285845f
C2490 vdd.t133 gnd 0.039365f
C2491 vdd.t299 gnd 0.039365f
C2492 vdd.n3 gnd 0.309963f
C2493 vdd.n4 gnd 0.144562f
C2494 vdd.t50 gnd 0.039365f
C2495 vdd.t131 gnd 0.039365f
C2496 vdd.n5 gnd 0.309963f
C2497 vdd.n6 gnd 0.135645f
C2498 vdd.t15 gnd 0.039365f
C2499 vdd.t25 gnd 0.039365f
C2500 vdd.n7 gnd 0.310475f
C2501 vdd.t38 gnd 0.039365f
C2502 vdd.t27 gnd 0.039365f
C2503 vdd.n8 gnd 0.309963f
C2504 vdd.n9 gnd 0.285845f
C2505 vdd.t17 gnd 0.039365f
C2506 vdd.t295 gnd 0.039365f
C2507 vdd.n10 gnd 0.309963f
C2508 vdd.n11 gnd 0.144562f
C2509 vdd.t23 gnd 0.039365f
C2510 vdd.t52 gnd 0.039365f
C2511 vdd.n12 gnd 0.309963f
C2512 vdd.n13 gnd 0.135645f
C2513 vdd.n14 gnd 0.095898f
C2514 vdd.t297 gnd 0.021869f
C2515 vdd.t46 gnd 0.021869f
C2516 vdd.n15 gnd 0.201297f
C2517 vdd.t39 gnd 0.021869f
C2518 vdd.t40 gnd 0.021869f
C2519 vdd.n16 gnd 0.200708f
C2520 vdd.n17 gnd 0.349295f
C2521 vdd.t34 gnd 0.021869f
C2522 vdd.t19 gnd 0.021869f
C2523 vdd.n18 gnd 0.200708f
C2524 vdd.n19 gnd 0.144508f
C2525 vdd.t44 gnd 0.021869f
C2526 vdd.t41 gnd 0.021869f
C2527 vdd.n20 gnd 0.201297f
C2528 vdd.t32 gnd 0.021869f
C2529 vdd.t29 gnd 0.021869f
C2530 vdd.n21 gnd 0.200708f
C2531 vdd.n22 gnd 0.349295f
C2532 vdd.t42 gnd 0.021869f
C2533 vdd.t43 gnd 0.021869f
C2534 vdd.n23 gnd 0.200708f
C2535 vdd.n24 gnd 0.144508f
C2536 vdd.t296 gnd 0.021869f
C2537 vdd.t28 gnd 0.021869f
C2538 vdd.n25 gnd 0.200708f
C2539 vdd.t45 gnd 0.021869f
C2540 vdd.t33 gnd 0.021869f
C2541 vdd.n26 gnd 0.200708f
C2542 vdd.n27 gnd 22.0053f
C2543 vdd.n28 gnd 8.55025f
C2544 vdd.n29 gnd 0.005965f
C2545 vdd.n30 gnd 0.005535f
C2546 vdd.n31 gnd 0.003062f
C2547 vdd.n32 gnd 0.00703f
C2548 vdd.n33 gnd 0.002974f
C2549 vdd.n34 gnd 0.003149f
C2550 vdd.n35 gnd 0.005535f
C2551 vdd.n36 gnd 0.002974f
C2552 vdd.n37 gnd 0.00703f
C2553 vdd.n38 gnd 0.003149f
C2554 vdd.n39 gnd 0.005535f
C2555 vdd.n40 gnd 0.002974f
C2556 vdd.n41 gnd 0.005272f
C2557 vdd.n42 gnd 0.005288f
C2558 vdd.t189 gnd 0.015103f
C2559 vdd.n43 gnd 0.033604f
C2560 vdd.n44 gnd 0.174886f
C2561 vdd.n45 gnd 0.002974f
C2562 vdd.n46 gnd 0.003149f
C2563 vdd.n47 gnd 0.00703f
C2564 vdd.n48 gnd 0.00703f
C2565 vdd.n49 gnd 0.003149f
C2566 vdd.n50 gnd 0.002974f
C2567 vdd.n51 gnd 0.005535f
C2568 vdd.n52 gnd 0.005535f
C2569 vdd.n53 gnd 0.002974f
C2570 vdd.n54 gnd 0.003149f
C2571 vdd.n55 gnd 0.00703f
C2572 vdd.n56 gnd 0.00703f
C2573 vdd.n57 gnd 0.003149f
C2574 vdd.n58 gnd 0.002974f
C2575 vdd.n59 gnd 0.005535f
C2576 vdd.n60 gnd 0.005535f
C2577 vdd.n61 gnd 0.002974f
C2578 vdd.n62 gnd 0.003149f
C2579 vdd.n63 gnd 0.00703f
C2580 vdd.n64 gnd 0.00703f
C2581 vdd.n65 gnd 0.01662f
C2582 vdd.n66 gnd 0.003062f
C2583 vdd.n67 gnd 0.002974f
C2584 vdd.n68 gnd 0.014306f
C2585 vdd.n69 gnd 0.009988f
C2586 vdd.t272 gnd 0.034991f
C2587 vdd.t217 gnd 0.034991f
C2588 vdd.n70 gnd 0.240481f
C2589 vdd.n71 gnd 0.189101f
C2590 vdd.t285 gnd 0.034991f
C2591 vdd.t267 gnd 0.034991f
C2592 vdd.n72 gnd 0.240481f
C2593 vdd.n73 gnd 0.152604f
C2594 vdd.t151 gnd 0.034991f
C2595 vdd.t204 gnd 0.034991f
C2596 vdd.n74 gnd 0.240481f
C2597 vdd.n75 gnd 0.152604f
C2598 vdd.t162 gnd 0.034991f
C2599 vdd.t174 gnd 0.034991f
C2600 vdd.n76 gnd 0.240481f
C2601 vdd.n77 gnd 0.152604f
C2602 vdd.t195 gnd 0.034991f
C2603 vdd.t276 gnd 0.034991f
C2604 vdd.n78 gnd 0.240481f
C2605 vdd.n79 gnd 0.152604f
C2606 vdd.t168 gnd 0.034991f
C2607 vdd.t248 gnd 0.034991f
C2608 vdd.n80 gnd 0.240481f
C2609 vdd.n81 gnd 0.152604f
C2610 vdd.t179 gnd 0.034991f
C2611 vdd.t262 gnd 0.034991f
C2612 vdd.n82 gnd 0.240481f
C2613 vdd.n83 gnd 0.152604f
C2614 vdd.t212 gnd 0.034991f
C2615 vdd.t280 gnd 0.034991f
C2616 vdd.n84 gnd 0.240481f
C2617 vdd.n85 gnd 0.152604f
C2618 vdd.t231 gnd 0.034991f
C2619 vdd.t258 gnd 0.034991f
C2620 vdd.n86 gnd 0.240481f
C2621 vdd.n87 gnd 0.152604f
C2622 vdd.n88 gnd 0.005965f
C2623 vdd.n89 gnd 0.005535f
C2624 vdd.n90 gnd 0.003062f
C2625 vdd.n91 gnd 0.00703f
C2626 vdd.n92 gnd 0.002974f
C2627 vdd.n93 gnd 0.003149f
C2628 vdd.n94 gnd 0.005535f
C2629 vdd.n95 gnd 0.002974f
C2630 vdd.n96 gnd 0.00703f
C2631 vdd.n97 gnd 0.003149f
C2632 vdd.n98 gnd 0.005535f
C2633 vdd.n99 gnd 0.002974f
C2634 vdd.n100 gnd 0.005272f
C2635 vdd.n101 gnd 0.005288f
C2636 vdd.t197 gnd 0.015103f
C2637 vdd.n102 gnd 0.033604f
C2638 vdd.n103 gnd 0.174886f
C2639 vdd.n104 gnd 0.002974f
C2640 vdd.n105 gnd 0.003149f
C2641 vdd.n106 gnd 0.00703f
C2642 vdd.n107 gnd 0.00703f
C2643 vdd.n108 gnd 0.003149f
C2644 vdd.n109 gnd 0.002974f
C2645 vdd.n110 gnd 0.005535f
C2646 vdd.n111 gnd 0.005535f
C2647 vdd.n112 gnd 0.002974f
C2648 vdd.n113 gnd 0.003149f
C2649 vdd.n114 gnd 0.00703f
C2650 vdd.n115 gnd 0.00703f
C2651 vdd.n116 gnd 0.003149f
C2652 vdd.n117 gnd 0.002974f
C2653 vdd.n118 gnd 0.005535f
C2654 vdd.n119 gnd 0.005535f
C2655 vdd.n120 gnd 0.002974f
C2656 vdd.n121 gnd 0.003149f
C2657 vdd.n122 gnd 0.00703f
C2658 vdd.n123 gnd 0.00703f
C2659 vdd.n124 gnd 0.01662f
C2660 vdd.n125 gnd 0.003062f
C2661 vdd.n126 gnd 0.002974f
C2662 vdd.n127 gnd 0.014306f
C2663 vdd.n128 gnd 0.009674f
C2664 vdd.n129 gnd 0.113538f
C2665 vdd.n130 gnd 0.005965f
C2666 vdd.n131 gnd 0.005535f
C2667 vdd.n132 gnd 0.003062f
C2668 vdd.n133 gnd 0.00703f
C2669 vdd.n134 gnd 0.002974f
C2670 vdd.n135 gnd 0.003149f
C2671 vdd.n136 gnd 0.005535f
C2672 vdd.n137 gnd 0.002974f
C2673 vdd.n138 gnd 0.00703f
C2674 vdd.n139 gnd 0.003149f
C2675 vdd.n140 gnd 0.005535f
C2676 vdd.n141 gnd 0.002974f
C2677 vdd.n142 gnd 0.005272f
C2678 vdd.n143 gnd 0.005288f
C2679 vdd.t228 gnd 0.015103f
C2680 vdd.n144 gnd 0.033604f
C2681 vdd.n145 gnd 0.174886f
C2682 vdd.n146 gnd 0.002974f
C2683 vdd.n147 gnd 0.003149f
C2684 vdd.n148 gnd 0.00703f
C2685 vdd.n149 gnd 0.00703f
C2686 vdd.n150 gnd 0.003149f
C2687 vdd.n151 gnd 0.002974f
C2688 vdd.n152 gnd 0.005535f
C2689 vdd.n153 gnd 0.005535f
C2690 vdd.n154 gnd 0.002974f
C2691 vdd.n155 gnd 0.003149f
C2692 vdd.n156 gnd 0.00703f
C2693 vdd.n157 gnd 0.00703f
C2694 vdd.n158 gnd 0.003149f
C2695 vdd.n159 gnd 0.002974f
C2696 vdd.n160 gnd 0.005535f
C2697 vdd.n161 gnd 0.005535f
C2698 vdd.n162 gnd 0.002974f
C2699 vdd.n163 gnd 0.003149f
C2700 vdd.n164 gnd 0.00703f
C2701 vdd.n165 gnd 0.00703f
C2702 vdd.n166 gnd 0.01662f
C2703 vdd.n167 gnd 0.003062f
C2704 vdd.n168 gnd 0.002974f
C2705 vdd.n169 gnd 0.014306f
C2706 vdd.n170 gnd 0.009988f
C2707 vdd.t257 gnd 0.034991f
C2708 vdd.t139 gnd 0.034991f
C2709 vdd.n171 gnd 0.240481f
C2710 vdd.n172 gnd 0.189101f
C2711 vdd.t201 gnd 0.034991f
C2712 vdd.t203 gnd 0.034991f
C2713 vdd.n173 gnd 0.240481f
C2714 vdd.n174 gnd 0.152604f
C2715 vdd.t279 gnd 0.034991f
C2716 vdd.t176 gnd 0.034991f
C2717 vdd.n175 gnd 0.240481f
C2718 vdd.n176 gnd 0.152604f
C2719 vdd.t193 gnd 0.034991f
C2720 vdd.t263 gnd 0.034991f
C2721 vdd.n177 gnd 0.240481f
C2722 vdd.n178 gnd 0.152604f
C2723 vdd.t278 gnd 0.034991f
C2724 vdd.t158 gnd 0.034991f
C2725 vdd.n179 gnd 0.240481f
C2726 vdd.n180 gnd 0.152604f
C2727 vdd.t260 gnd 0.034991f
C2728 vdd.t275 gnd 0.034991f
C2729 vdd.n181 gnd 0.240481f
C2730 vdd.n182 gnd 0.152604f
C2731 vdd.t156 gnd 0.034991f
C2732 vdd.t227 gnd 0.034991f
C2733 vdd.n183 gnd 0.240481f
C2734 vdd.n184 gnd 0.152604f
C2735 vdd.t255 gnd 0.034991f
C2736 vdd.t286 gnd 0.034991f
C2737 vdd.n185 gnd 0.240481f
C2738 vdd.n186 gnd 0.152604f
C2739 vdd.t199 gnd 0.034991f
C2740 vdd.t254 gnd 0.034991f
C2741 vdd.n187 gnd 0.240481f
C2742 vdd.n188 gnd 0.152604f
C2743 vdd.n189 gnd 0.005965f
C2744 vdd.n190 gnd 0.005535f
C2745 vdd.n191 gnd 0.003062f
C2746 vdd.n192 gnd 0.00703f
C2747 vdd.n193 gnd 0.002974f
C2748 vdd.n194 gnd 0.003149f
C2749 vdd.n195 gnd 0.005535f
C2750 vdd.n196 gnd 0.002974f
C2751 vdd.n197 gnd 0.00703f
C2752 vdd.n198 gnd 0.003149f
C2753 vdd.n199 gnd 0.005535f
C2754 vdd.n200 gnd 0.002974f
C2755 vdd.n201 gnd 0.005272f
C2756 vdd.n202 gnd 0.005288f
C2757 vdd.t291 gnd 0.015103f
C2758 vdd.n203 gnd 0.033604f
C2759 vdd.n204 gnd 0.174886f
C2760 vdd.n205 gnd 0.002974f
C2761 vdd.n206 gnd 0.003149f
C2762 vdd.n207 gnd 0.00703f
C2763 vdd.n208 gnd 0.00703f
C2764 vdd.n209 gnd 0.003149f
C2765 vdd.n210 gnd 0.002974f
C2766 vdd.n211 gnd 0.005535f
C2767 vdd.n212 gnd 0.005535f
C2768 vdd.n213 gnd 0.002974f
C2769 vdd.n214 gnd 0.003149f
C2770 vdd.n215 gnd 0.00703f
C2771 vdd.n216 gnd 0.00703f
C2772 vdd.n217 gnd 0.003149f
C2773 vdd.n218 gnd 0.002974f
C2774 vdd.n219 gnd 0.005535f
C2775 vdd.n220 gnd 0.005535f
C2776 vdd.n221 gnd 0.002974f
C2777 vdd.n222 gnd 0.003149f
C2778 vdd.n223 gnd 0.00703f
C2779 vdd.n224 gnd 0.00703f
C2780 vdd.n225 gnd 0.01662f
C2781 vdd.n226 gnd 0.003062f
C2782 vdd.n227 gnd 0.002974f
C2783 vdd.n228 gnd 0.014306f
C2784 vdd.n229 gnd 0.009674f
C2785 vdd.n230 gnd 0.067544f
C2786 vdd.n231 gnd 0.243377f
C2787 vdd.n232 gnd 0.005965f
C2788 vdd.n233 gnd 0.005535f
C2789 vdd.n234 gnd 0.003062f
C2790 vdd.n235 gnd 0.00703f
C2791 vdd.n236 gnd 0.002974f
C2792 vdd.n237 gnd 0.003149f
C2793 vdd.n238 gnd 0.005535f
C2794 vdd.n239 gnd 0.002974f
C2795 vdd.n240 gnd 0.00703f
C2796 vdd.n241 gnd 0.003149f
C2797 vdd.n242 gnd 0.005535f
C2798 vdd.n243 gnd 0.002974f
C2799 vdd.n244 gnd 0.005272f
C2800 vdd.n245 gnd 0.005288f
C2801 vdd.t240 gnd 0.015103f
C2802 vdd.n246 gnd 0.033604f
C2803 vdd.n247 gnd 0.174886f
C2804 vdd.n248 gnd 0.002974f
C2805 vdd.n249 gnd 0.003149f
C2806 vdd.n250 gnd 0.00703f
C2807 vdd.n251 gnd 0.00703f
C2808 vdd.n252 gnd 0.003149f
C2809 vdd.n253 gnd 0.002974f
C2810 vdd.n254 gnd 0.005535f
C2811 vdd.n255 gnd 0.005535f
C2812 vdd.n256 gnd 0.002974f
C2813 vdd.n257 gnd 0.003149f
C2814 vdd.n258 gnd 0.00703f
C2815 vdd.n259 gnd 0.00703f
C2816 vdd.n260 gnd 0.003149f
C2817 vdd.n261 gnd 0.002974f
C2818 vdd.n262 gnd 0.005535f
C2819 vdd.n263 gnd 0.005535f
C2820 vdd.n264 gnd 0.002974f
C2821 vdd.n265 gnd 0.003149f
C2822 vdd.n266 gnd 0.00703f
C2823 vdd.n267 gnd 0.00703f
C2824 vdd.n268 gnd 0.01662f
C2825 vdd.n269 gnd 0.003062f
C2826 vdd.n270 gnd 0.002974f
C2827 vdd.n271 gnd 0.014306f
C2828 vdd.n272 gnd 0.009988f
C2829 vdd.t269 gnd 0.034991f
C2830 vdd.t166 gnd 0.034991f
C2831 vdd.n273 gnd 0.240481f
C2832 vdd.n274 gnd 0.189101f
C2833 vdd.t221 gnd 0.034991f
C2834 vdd.t224 gnd 0.034991f
C2835 vdd.n275 gnd 0.240481f
C2836 vdd.n276 gnd 0.152604f
C2837 vdd.t290 gnd 0.034991f
C2838 vdd.t215 gnd 0.034991f
C2839 vdd.n277 gnd 0.240481f
C2840 vdd.n278 gnd 0.152604f
C2841 vdd.t216 gnd 0.034991f
C2842 vdd.t288 gnd 0.034991f
C2843 vdd.n279 gnd 0.240481f
C2844 vdd.n280 gnd 0.152604f
C2845 vdd.t289 gnd 0.034991f
C2846 vdd.t187 gnd 0.034991f
C2847 vdd.n281 gnd 0.240481f
C2848 vdd.n282 gnd 0.152604f
C2849 vdd.t274 gnd 0.034991f
C2850 vdd.t284 gnd 0.034991f
C2851 vdd.n283 gnd 0.240481f
C2852 vdd.n284 gnd 0.152604f
C2853 vdd.t180 gnd 0.034991f
C2854 vdd.t241 gnd 0.034991f
C2855 vdd.n285 gnd 0.240481f
C2856 vdd.n286 gnd 0.152604f
C2857 vdd.t270 gnd 0.034991f
C2858 vdd.t143 gnd 0.034991f
C2859 vdd.n287 gnd 0.240481f
C2860 vdd.n288 gnd 0.152604f
C2861 vdd.t222 gnd 0.034991f
C2862 vdd.t268 gnd 0.034991f
C2863 vdd.n289 gnd 0.240481f
C2864 vdd.n290 gnd 0.152604f
C2865 vdd.n291 gnd 0.005965f
C2866 vdd.n292 gnd 0.005535f
C2867 vdd.n293 gnd 0.003062f
C2868 vdd.n294 gnd 0.00703f
C2869 vdd.n295 gnd 0.002974f
C2870 vdd.n296 gnd 0.003149f
C2871 vdd.n297 gnd 0.005535f
C2872 vdd.n298 gnd 0.002974f
C2873 vdd.n299 gnd 0.00703f
C2874 vdd.n300 gnd 0.003149f
C2875 vdd.n301 gnd 0.005535f
C2876 vdd.n302 gnd 0.002974f
C2877 vdd.n303 gnd 0.005272f
C2878 vdd.n304 gnd 0.005288f
C2879 vdd.t160 gnd 0.015103f
C2880 vdd.n305 gnd 0.033604f
C2881 vdd.n306 gnd 0.174886f
C2882 vdd.n307 gnd 0.002974f
C2883 vdd.n308 gnd 0.003149f
C2884 vdd.n309 gnd 0.00703f
C2885 vdd.n310 gnd 0.00703f
C2886 vdd.n311 gnd 0.003149f
C2887 vdd.n312 gnd 0.002974f
C2888 vdd.n313 gnd 0.005535f
C2889 vdd.n314 gnd 0.005535f
C2890 vdd.n315 gnd 0.002974f
C2891 vdd.n316 gnd 0.003149f
C2892 vdd.n317 gnd 0.00703f
C2893 vdd.n318 gnd 0.00703f
C2894 vdd.n319 gnd 0.003149f
C2895 vdd.n320 gnd 0.002974f
C2896 vdd.n321 gnd 0.005535f
C2897 vdd.n322 gnd 0.005535f
C2898 vdd.n323 gnd 0.002974f
C2899 vdd.n324 gnd 0.003149f
C2900 vdd.n325 gnd 0.00703f
C2901 vdd.n326 gnd 0.00703f
C2902 vdd.n327 gnd 0.01662f
C2903 vdd.n328 gnd 0.003062f
C2904 vdd.n329 gnd 0.002974f
C2905 vdd.n330 gnd 0.014306f
C2906 vdd.n331 gnd 0.009674f
C2907 vdd.n332 gnd 0.067544f
C2908 vdd.n333 gnd 0.278614f
C2909 vdd.n334 gnd 0.008353f
C2910 vdd.n335 gnd 0.010868f
C2911 vdd.n336 gnd 0.008748f
C2912 vdd.n337 gnd 0.008748f
C2913 vdd.n338 gnd 0.010868f
C2914 vdd.n339 gnd 0.010868f
C2915 vdd.n340 gnd 0.794145f
C2916 vdd.n341 gnd 0.010868f
C2917 vdd.n342 gnd 0.010868f
C2918 vdd.n343 gnd 0.010868f
C2919 vdd.n344 gnd 0.860786f
C2920 vdd.n345 gnd 0.010868f
C2921 vdd.n346 gnd 0.010868f
C2922 vdd.n347 gnd 0.010868f
C2923 vdd.n348 gnd 0.010868f
C2924 vdd.n349 gnd 0.008748f
C2925 vdd.n350 gnd 0.010868f
C2926 vdd.t247 gnd 0.555346f
C2927 vdd.n351 gnd 0.010868f
C2928 vdd.n352 gnd 0.010868f
C2929 vdd.n353 gnd 0.010868f
C2930 vdd.t226 gnd 0.555346f
C2931 vdd.n354 gnd 0.010868f
C2932 vdd.n355 gnd 0.010868f
C2933 vdd.n356 gnd 0.010868f
C2934 vdd.n357 gnd 0.010868f
C2935 vdd.n358 gnd 0.010868f
C2936 vdd.n359 gnd 0.008748f
C2937 vdd.n360 gnd 0.010868f
C2938 vdd.n361 gnd 0.627541f
C2939 vdd.n362 gnd 0.010868f
C2940 vdd.n363 gnd 0.010868f
C2941 vdd.n364 gnd 0.010868f
C2942 vdd.t142 gnd 0.555346f
C2943 vdd.n365 gnd 0.010868f
C2944 vdd.n366 gnd 0.010868f
C2945 vdd.n367 gnd 0.010868f
C2946 vdd.n368 gnd 0.010868f
C2947 vdd.n369 gnd 0.010868f
C2948 vdd.n370 gnd 0.008748f
C2949 vdd.n371 gnd 0.010868f
C2950 vdd.t198 gnd 0.555346f
C2951 vdd.n372 gnd 0.010868f
C2952 vdd.n373 gnd 0.010868f
C2953 vdd.n374 gnd 0.010868f
C2954 vdd.n375 gnd 0.649755f
C2955 vdd.n376 gnd 0.010868f
C2956 vdd.n377 gnd 0.010868f
C2957 vdd.n378 gnd 0.010868f
C2958 vdd.n379 gnd 0.010868f
C2959 vdd.n380 gnd 0.010868f
C2960 vdd.n381 gnd 0.008748f
C2961 vdd.n382 gnd 0.010868f
C2962 vdd.t159 gnd 0.555346f
C2963 vdd.n383 gnd 0.010868f
C2964 vdd.n384 gnd 0.010868f
C2965 vdd.n385 gnd 0.010868f
C2966 vdd.n386 gnd 0.560899f
C2967 vdd.n387 gnd 0.010868f
C2968 vdd.n388 gnd 0.010868f
C2969 vdd.n389 gnd 0.010868f
C2970 vdd.n390 gnd 0.010868f
C2971 vdd.n391 gnd 0.026291f
C2972 vdd.n392 gnd 0.026855f
C2973 vdd.t77 gnd 0.555346f
C2974 vdd.n393 gnd 0.026291f
C2975 vdd.n425 gnd 0.010868f
C2976 vdd.t89 gnd 0.133709f
C2977 vdd.t88 gnd 0.142898f
C2978 vdd.t87 gnd 0.174622f
C2979 vdd.n426 gnd 0.223841f
C2980 vdd.n427 gnd 0.188942f
C2981 vdd.n428 gnd 0.014346f
C2982 vdd.n429 gnd 0.010868f
C2983 vdd.n430 gnd 0.008748f
C2984 vdd.n431 gnd 0.010868f
C2985 vdd.n432 gnd 0.008748f
C2986 vdd.n433 gnd 0.010868f
C2987 vdd.n434 gnd 0.008748f
C2988 vdd.n435 gnd 0.010868f
C2989 vdd.n436 gnd 0.008748f
C2990 vdd.n437 gnd 0.010868f
C2991 vdd.n438 gnd 0.008748f
C2992 vdd.n439 gnd 0.010868f
C2993 vdd.t79 gnd 0.133709f
C2994 vdd.t78 gnd 0.142898f
C2995 vdd.t76 gnd 0.174622f
C2996 vdd.n440 gnd 0.223841f
C2997 vdd.n441 gnd 0.188942f
C2998 vdd.n442 gnd 0.008748f
C2999 vdd.n443 gnd 0.010868f
C3000 vdd.n444 gnd 0.008748f
C3001 vdd.n445 gnd 0.010868f
C3002 vdd.n446 gnd 0.008748f
C3003 vdd.n447 gnd 0.010868f
C3004 vdd.n448 gnd 0.008748f
C3005 vdd.n449 gnd 0.010868f
C3006 vdd.n450 gnd 0.008748f
C3007 vdd.n451 gnd 0.010868f
C3008 vdd.t96 gnd 0.133709f
C3009 vdd.t95 gnd 0.142898f
C3010 vdd.t94 gnd 0.174622f
C3011 vdd.n452 gnd 0.223841f
C3012 vdd.n453 gnd 0.188942f
C3013 vdd.n454 gnd 0.01872f
C3014 vdd.n455 gnd 0.010868f
C3015 vdd.n456 gnd 0.008748f
C3016 vdd.n457 gnd 0.010868f
C3017 vdd.n458 gnd 0.008748f
C3018 vdd.n459 gnd 0.010868f
C3019 vdd.n460 gnd 0.008748f
C3020 vdd.n461 gnd 0.010868f
C3021 vdd.n462 gnd 0.008748f
C3022 vdd.n463 gnd 0.010868f
C3023 vdd.n464 gnd 0.026855f
C3024 vdd.n465 gnd 0.007261f
C3025 vdd.n466 gnd 0.008748f
C3026 vdd.n467 gnd 0.010868f
C3027 vdd.n468 gnd 0.010868f
C3028 vdd.n469 gnd 0.008748f
C3029 vdd.n470 gnd 0.010868f
C3030 vdd.n471 gnd 0.010868f
C3031 vdd.n472 gnd 0.010868f
C3032 vdd.n473 gnd 0.010868f
C3033 vdd.n474 gnd 0.010868f
C3034 vdd.n475 gnd 0.008748f
C3035 vdd.n476 gnd 0.008748f
C3036 vdd.n477 gnd 0.010868f
C3037 vdd.n478 gnd 0.010868f
C3038 vdd.n479 gnd 0.008748f
C3039 vdd.n480 gnd 0.010868f
C3040 vdd.n481 gnd 0.010868f
C3041 vdd.n482 gnd 0.010868f
C3042 vdd.n483 gnd 0.010868f
C3043 vdd.n484 gnd 0.010868f
C3044 vdd.n485 gnd 0.008748f
C3045 vdd.n486 gnd 0.008748f
C3046 vdd.n487 gnd 0.010868f
C3047 vdd.n488 gnd 0.010868f
C3048 vdd.n489 gnd 0.008748f
C3049 vdd.n490 gnd 0.010868f
C3050 vdd.n491 gnd 0.010868f
C3051 vdd.n492 gnd 0.010868f
C3052 vdd.n493 gnd 0.010868f
C3053 vdd.n494 gnd 0.010868f
C3054 vdd.n495 gnd 0.008748f
C3055 vdd.n496 gnd 0.008748f
C3056 vdd.n497 gnd 0.010868f
C3057 vdd.n498 gnd 0.010868f
C3058 vdd.n499 gnd 0.008748f
C3059 vdd.n500 gnd 0.010868f
C3060 vdd.n501 gnd 0.010868f
C3061 vdd.n502 gnd 0.010868f
C3062 vdd.n503 gnd 0.010868f
C3063 vdd.n504 gnd 0.010868f
C3064 vdd.n505 gnd 0.008748f
C3065 vdd.n506 gnd 0.008748f
C3066 vdd.n507 gnd 0.010868f
C3067 vdd.n508 gnd 0.010868f
C3068 vdd.n509 gnd 0.007304f
C3069 vdd.n510 gnd 0.010868f
C3070 vdd.n511 gnd 0.010868f
C3071 vdd.n512 gnd 0.010868f
C3072 vdd.n513 gnd 0.010868f
C3073 vdd.n514 gnd 0.010868f
C3074 vdd.n515 gnd 0.007304f
C3075 vdd.n516 gnd 0.008748f
C3076 vdd.n517 gnd 0.010868f
C3077 vdd.n518 gnd 0.010868f
C3078 vdd.n519 gnd 0.008748f
C3079 vdd.n520 gnd 0.010868f
C3080 vdd.n521 gnd 0.010868f
C3081 vdd.n522 gnd 0.010868f
C3082 vdd.n523 gnd 0.010868f
C3083 vdd.n524 gnd 0.010868f
C3084 vdd.n525 gnd 0.008748f
C3085 vdd.n526 gnd 0.008748f
C3086 vdd.n527 gnd 0.010868f
C3087 vdd.n528 gnd 0.010868f
C3088 vdd.n529 gnd 0.008748f
C3089 vdd.n530 gnd 0.010868f
C3090 vdd.n531 gnd 0.010868f
C3091 vdd.n532 gnd 0.010868f
C3092 vdd.n533 gnd 0.010868f
C3093 vdd.n534 gnd 0.010868f
C3094 vdd.n535 gnd 0.008748f
C3095 vdd.n536 gnd 0.008748f
C3096 vdd.n537 gnd 0.010868f
C3097 vdd.n538 gnd 0.010868f
C3098 vdd.n539 gnd 0.008748f
C3099 vdd.n540 gnd 0.010868f
C3100 vdd.n541 gnd 0.010868f
C3101 vdd.n542 gnd 0.010868f
C3102 vdd.n543 gnd 0.010868f
C3103 vdd.n544 gnd 0.010868f
C3104 vdd.n545 gnd 0.008748f
C3105 vdd.n546 gnd 0.008748f
C3106 vdd.n547 gnd 0.010868f
C3107 vdd.n548 gnd 0.010868f
C3108 vdd.n549 gnd 0.008748f
C3109 vdd.n550 gnd 0.010868f
C3110 vdd.n551 gnd 0.010868f
C3111 vdd.n552 gnd 0.010868f
C3112 vdd.n553 gnd 0.010868f
C3113 vdd.n554 gnd 0.010868f
C3114 vdd.n555 gnd 0.008748f
C3115 vdd.n556 gnd 0.008748f
C3116 vdd.n557 gnd 0.010868f
C3117 vdd.n558 gnd 0.010868f
C3118 vdd.n559 gnd 0.008748f
C3119 vdd.n560 gnd 0.010868f
C3120 vdd.n561 gnd 0.010868f
C3121 vdd.n562 gnd 0.010868f
C3122 vdd.n563 gnd 0.010868f
C3123 vdd.n564 gnd 0.010868f
C3124 vdd.n565 gnd 0.005948f
C3125 vdd.n566 gnd 0.01872f
C3126 vdd.n567 gnd 0.010868f
C3127 vdd.n568 gnd 0.010868f
C3128 vdd.n569 gnd 0.00866f
C3129 vdd.n570 gnd 0.010868f
C3130 vdd.n571 gnd 0.010868f
C3131 vdd.n572 gnd 0.010868f
C3132 vdd.n573 gnd 0.010868f
C3133 vdd.n574 gnd 0.010868f
C3134 vdd.n575 gnd 0.008748f
C3135 vdd.n576 gnd 0.008748f
C3136 vdd.n577 gnd 0.010868f
C3137 vdd.n578 gnd 0.010868f
C3138 vdd.n579 gnd 0.008748f
C3139 vdd.n580 gnd 0.010868f
C3140 vdd.n581 gnd 0.010868f
C3141 vdd.n582 gnd 0.010868f
C3142 vdd.n583 gnd 0.010868f
C3143 vdd.n584 gnd 0.010868f
C3144 vdd.n585 gnd 0.008748f
C3145 vdd.n586 gnd 0.008748f
C3146 vdd.n587 gnd 0.010868f
C3147 vdd.n588 gnd 0.010868f
C3148 vdd.n589 gnd 0.008748f
C3149 vdd.n590 gnd 0.010868f
C3150 vdd.n591 gnd 0.010868f
C3151 vdd.n592 gnd 0.010868f
C3152 vdd.n593 gnd 0.010868f
C3153 vdd.n594 gnd 0.010868f
C3154 vdd.n595 gnd 0.008748f
C3155 vdd.n596 gnd 0.008748f
C3156 vdd.n597 gnd 0.010868f
C3157 vdd.n598 gnd 0.010868f
C3158 vdd.n599 gnd 0.008748f
C3159 vdd.n600 gnd 0.010868f
C3160 vdd.n601 gnd 0.010868f
C3161 vdd.n602 gnd 0.010868f
C3162 vdd.n603 gnd 0.010868f
C3163 vdd.n604 gnd 0.010868f
C3164 vdd.n605 gnd 0.008748f
C3165 vdd.n606 gnd 0.008748f
C3166 vdd.n607 gnd 0.010868f
C3167 vdd.n608 gnd 0.010868f
C3168 vdd.n609 gnd 0.008748f
C3169 vdd.n610 gnd 0.010868f
C3170 vdd.n611 gnd 0.010868f
C3171 vdd.n612 gnd 0.010868f
C3172 vdd.n613 gnd 0.010868f
C3173 vdd.n614 gnd 0.010868f
C3174 vdd.n615 gnd 0.008748f
C3175 vdd.n616 gnd 0.010868f
C3176 vdd.n617 gnd 0.008748f
C3177 vdd.n618 gnd 0.004593f
C3178 vdd.n619 gnd 0.010868f
C3179 vdd.n620 gnd 0.010868f
C3180 vdd.n621 gnd 0.008748f
C3181 vdd.n622 gnd 0.010868f
C3182 vdd.n623 gnd 0.008748f
C3183 vdd.n624 gnd 0.010868f
C3184 vdd.n625 gnd 0.008748f
C3185 vdd.n626 gnd 0.010868f
C3186 vdd.n627 gnd 0.008748f
C3187 vdd.n628 gnd 0.010868f
C3188 vdd.n629 gnd 0.008748f
C3189 vdd.n630 gnd 0.010868f
C3190 vdd.n631 gnd 0.008748f
C3191 vdd.n632 gnd 0.010868f
C3192 vdd.n633 gnd 0.605327f
C3193 vdd.t194 gnd 0.555346f
C3194 vdd.n634 gnd 0.010868f
C3195 vdd.n635 gnd 0.008748f
C3196 vdd.n636 gnd 0.010868f
C3197 vdd.n637 gnd 0.008748f
C3198 vdd.n638 gnd 0.010868f
C3199 vdd.t161 gnd 0.555346f
C3200 vdd.n639 gnd 0.010868f
C3201 vdd.n640 gnd 0.008748f
C3202 vdd.n641 gnd 0.010868f
C3203 vdd.n642 gnd 0.008748f
C3204 vdd.n643 gnd 0.010868f
C3205 vdd.t175 gnd 0.555346f
C3206 vdd.n644 gnd 0.694182f
C3207 vdd.n645 gnd 0.010868f
C3208 vdd.n646 gnd 0.008748f
C3209 vdd.n647 gnd 0.010868f
C3210 vdd.n648 gnd 0.008748f
C3211 vdd.n649 gnd 0.010868f
C3212 vdd.t150 gnd 0.555346f
C3213 vdd.n650 gnd 0.010868f
C3214 vdd.n651 gnd 0.008748f
C3215 vdd.n652 gnd 0.010868f
C3216 vdd.n653 gnd 0.008748f
C3217 vdd.n654 gnd 0.010868f
C3218 vdd.n655 gnd 0.771931f
C3219 vdd.n656 gnd 0.921874f
C3220 vdd.t202 gnd 0.555346f
C3221 vdd.n657 gnd 0.010868f
C3222 vdd.n658 gnd 0.008748f
C3223 vdd.n659 gnd 0.010868f
C3224 vdd.n660 gnd 0.008748f
C3225 vdd.n661 gnd 0.010868f
C3226 vdd.n662 gnd 0.583113f
C3227 vdd.n663 gnd 0.010868f
C3228 vdd.n664 gnd 0.008748f
C3229 vdd.n665 gnd 0.010868f
C3230 vdd.n666 gnd 0.008748f
C3231 vdd.n667 gnd 0.010868f
C3232 vdd.t256 gnd 0.555346f
C3233 vdd.t138 gnd 0.555346f
C3234 vdd.n668 gnd 0.010868f
C3235 vdd.n669 gnd 0.008748f
C3236 vdd.n670 gnd 0.010868f
C3237 vdd.n671 gnd 0.008748f
C3238 vdd.n672 gnd 0.010868f
C3239 vdd.t188 gnd 0.555346f
C3240 vdd.n673 gnd 0.010868f
C3241 vdd.n674 gnd 0.008748f
C3242 vdd.n675 gnd 0.010868f
C3243 vdd.n676 gnd 0.008748f
C3244 vdd.n677 gnd 0.010868f
C3245 vdd.n678 gnd 1.11069f
C3246 vdd.n679 gnd 0.905214f
C3247 vdd.n680 gnd 0.010868f
C3248 vdd.n681 gnd 0.008748f
C3249 vdd.n682 gnd 0.026291f
C3250 vdd.n683 gnd 0.007261f
C3251 vdd.n684 gnd 0.026291f
C3252 vdd.t63 gnd 0.555346f
C3253 vdd.n685 gnd 0.026291f
C3254 vdd.n686 gnd 0.007261f
C3255 vdd.n687 gnd 0.009347f
C3256 vdd.t64 gnd 0.133709f
C3257 vdd.t65 gnd 0.142898f
C3258 vdd.t62 gnd 0.174622f
C3259 vdd.n688 gnd 0.223841f
C3260 vdd.n689 gnd 0.188067f
C3261 vdd.n690 gnd 0.013471f
C3262 vdd.n691 gnd 0.010868f
C3263 vdd.n692 gnd 9.4742f
C3264 vdd.n723 gnd 1.5272f
C3265 vdd.n724 gnd 0.010868f
C3266 vdd.n725 gnd 0.010868f
C3267 vdd.n726 gnd 0.026855f
C3268 vdd.n727 gnd 0.009347f
C3269 vdd.n728 gnd 0.010868f
C3270 vdd.n729 gnd 0.008748f
C3271 vdd.n730 gnd 0.006956f
C3272 vdd.n731 gnd 0.025382f
C3273 vdd.n732 gnd 0.008748f
C3274 vdd.n733 gnd 0.010868f
C3275 vdd.n734 gnd 0.010868f
C3276 vdd.n735 gnd 0.010868f
C3277 vdd.n736 gnd 0.010868f
C3278 vdd.n737 gnd 0.010868f
C3279 vdd.n738 gnd 0.010868f
C3280 vdd.n739 gnd 0.010868f
C3281 vdd.n740 gnd 0.010868f
C3282 vdd.n741 gnd 0.010868f
C3283 vdd.n742 gnd 0.010868f
C3284 vdd.n743 gnd 0.010868f
C3285 vdd.n744 gnd 0.010868f
C3286 vdd.n745 gnd 0.010868f
C3287 vdd.n746 gnd 0.010868f
C3288 vdd.n747 gnd 0.007304f
C3289 vdd.n748 gnd 0.010868f
C3290 vdd.n749 gnd 0.010868f
C3291 vdd.n750 gnd 0.010868f
C3292 vdd.n751 gnd 0.010868f
C3293 vdd.n752 gnd 0.010868f
C3294 vdd.n753 gnd 0.010868f
C3295 vdd.n754 gnd 0.010868f
C3296 vdd.n755 gnd 0.010868f
C3297 vdd.n756 gnd 0.010868f
C3298 vdd.n757 gnd 0.010868f
C3299 vdd.n758 gnd 0.010868f
C3300 vdd.n759 gnd 0.010868f
C3301 vdd.n760 gnd 0.010868f
C3302 vdd.n761 gnd 0.010868f
C3303 vdd.n762 gnd 0.010868f
C3304 vdd.n763 gnd 0.010868f
C3305 vdd.n764 gnd 0.010868f
C3306 vdd.n765 gnd 0.010868f
C3307 vdd.n766 gnd 0.010868f
C3308 vdd.n767 gnd 0.00866f
C3309 vdd.t71 gnd 0.133709f
C3310 vdd.t72 gnd 0.142898f
C3311 vdd.t70 gnd 0.174622f
C3312 vdd.n768 gnd 0.223841f
C3313 vdd.n769 gnd 0.188067f
C3314 vdd.n770 gnd 0.010868f
C3315 vdd.n771 gnd 0.010868f
C3316 vdd.n772 gnd 0.010868f
C3317 vdd.n773 gnd 0.010868f
C3318 vdd.n774 gnd 0.010868f
C3319 vdd.n775 gnd 0.010868f
C3320 vdd.n776 gnd 0.010868f
C3321 vdd.n777 gnd 0.010868f
C3322 vdd.n778 gnd 0.010868f
C3323 vdd.n779 gnd 0.010868f
C3324 vdd.n780 gnd 0.010868f
C3325 vdd.n781 gnd 0.010868f
C3326 vdd.n782 gnd 0.010868f
C3327 vdd.n783 gnd 0.006956f
C3328 vdd.n785 gnd 0.00739f
C3329 vdd.n786 gnd 0.00739f
C3330 vdd.n787 gnd 0.00739f
C3331 vdd.n788 gnd 0.00739f
C3332 vdd.n789 gnd 0.00739f
C3333 vdd.n790 gnd 0.00739f
C3334 vdd.n792 gnd 0.00739f
C3335 vdd.n793 gnd 0.00739f
C3336 vdd.n795 gnd 0.00739f
C3337 vdd.n796 gnd 0.00538f
C3338 vdd.n798 gnd 0.00739f
C3339 vdd.t57 gnd 0.298648f
C3340 vdd.t56 gnd 0.305703f
C3341 vdd.t54 gnd 0.194969f
C3342 vdd.n799 gnd 0.10537f
C3343 vdd.n800 gnd 0.059769f
C3344 vdd.n801 gnd 0.010562f
C3345 vdd.n802 gnd 0.017107f
C3346 vdd.n804 gnd 0.00739f
C3347 vdd.n805 gnd 0.755271f
C3348 vdd.n806 gnd 0.016189f
C3349 vdd.n807 gnd 0.016189f
C3350 vdd.n808 gnd 0.00739f
C3351 vdd.n809 gnd 0.017286f
C3352 vdd.n810 gnd 0.00739f
C3353 vdd.n811 gnd 0.00739f
C3354 vdd.n812 gnd 0.00739f
C3355 vdd.n813 gnd 0.00739f
C3356 vdd.n814 gnd 0.00739f
C3357 vdd.n816 gnd 0.00739f
C3358 vdd.n817 gnd 0.00739f
C3359 vdd.n819 gnd 0.00739f
C3360 vdd.n820 gnd 0.00739f
C3361 vdd.n822 gnd 0.00739f
C3362 vdd.n823 gnd 0.00739f
C3363 vdd.n825 gnd 0.00739f
C3364 vdd.n826 gnd 0.00739f
C3365 vdd.n828 gnd 0.00739f
C3366 vdd.n829 gnd 0.00739f
C3367 vdd.n831 gnd 0.00739f
C3368 vdd.t129 gnd 0.298648f
C3369 vdd.t128 gnd 0.305703f
C3370 vdd.t127 gnd 0.194969f
C3371 vdd.n832 gnd 0.10537f
C3372 vdd.n833 gnd 0.059769f
C3373 vdd.n834 gnd 0.00739f
C3374 vdd.n836 gnd 0.00739f
C3375 vdd.n837 gnd 0.00739f
C3376 vdd.t55 gnd 0.377635f
C3377 vdd.n838 gnd 0.00739f
C3378 vdd.n839 gnd 0.00739f
C3379 vdd.n840 gnd 0.00739f
C3380 vdd.n841 gnd 0.00739f
C3381 vdd.n842 gnd 0.00739f
C3382 vdd.n843 gnd 0.755271f
C3383 vdd.n844 gnd 0.00739f
C3384 vdd.n845 gnd 0.00739f
C3385 vdd.n846 gnd 0.638648f
C3386 vdd.n847 gnd 0.00739f
C3387 vdd.n848 gnd 0.00739f
C3388 vdd.n849 gnd 0.00739f
C3389 vdd.n850 gnd 0.00739f
C3390 vdd.n851 gnd 0.73861f
C3391 vdd.n852 gnd 0.00739f
C3392 vdd.n853 gnd 0.00739f
C3393 vdd.n854 gnd 0.00739f
C3394 vdd.n855 gnd 0.00739f
C3395 vdd.n856 gnd 0.00739f
C3396 vdd.n857 gnd 0.755271f
C3397 vdd.n858 gnd 0.00739f
C3398 vdd.n859 gnd 0.00739f
C3399 vdd.t4 gnd 0.377635f
C3400 vdd.n860 gnd 0.00739f
C3401 vdd.n861 gnd 0.00739f
C3402 vdd.n862 gnd 0.00739f
C3403 vdd.t20 gnd 0.377635f
C3404 vdd.n863 gnd 0.00739f
C3405 vdd.n864 gnd 0.00739f
C3406 vdd.n865 gnd 0.00739f
C3407 vdd.n866 gnd 0.00739f
C3408 vdd.n867 gnd 0.00739f
C3409 vdd.t81 gnd 0.316547f
C3410 vdd.n868 gnd 0.00739f
C3411 vdd.n869 gnd 0.00739f
C3412 vdd.n870 gnd 0.605327f
C3413 vdd.n871 gnd 0.00739f
C3414 vdd.t82 gnd 0.305703f
C3415 vdd.t80 gnd 0.194969f
C3416 vdd.t83 gnd 0.305703f
C3417 vdd.n872 gnd 0.171818f
C3418 vdd.n873 gnd 0.00739f
C3419 vdd.n874 gnd 0.00739f
C3420 vdd.n875 gnd 0.483151f
C3421 vdd.n876 gnd 0.00739f
C3422 vdd.n877 gnd 0.00739f
C3423 vdd.t7 gnd 0.111069f
C3424 vdd.n878 gnd 0.438723f
C3425 vdd.n879 gnd 0.00739f
C3426 vdd.n880 gnd 0.00739f
C3427 vdd.n881 gnd 0.00739f
C3428 vdd.n882 gnd 0.649755f
C3429 vdd.n883 gnd 0.00739f
C3430 vdd.n884 gnd 0.00739f
C3431 vdd.t30 gnd 0.377635f
C3432 vdd.n885 gnd 0.00739f
C3433 vdd.n886 gnd 0.00739f
C3434 vdd.n887 gnd 0.00739f
C3435 vdd.t24 gnd 0.377635f
C3436 vdd.n888 gnd 0.00739f
C3437 vdd.n889 gnd 0.00739f
C3438 vdd.t36 gnd 0.377635f
C3439 vdd.n890 gnd 0.00739f
C3440 vdd.n891 gnd 0.00739f
C3441 vdd.n892 gnd 0.00739f
C3442 vdd.t35 gnd 0.299887f
C3443 vdd.n893 gnd 0.00739f
C3444 vdd.n894 gnd 0.00739f
C3445 vdd.n895 gnd 0.621988f
C3446 vdd.n896 gnd 0.00739f
C3447 vdd.n897 gnd 0.00739f
C3448 vdd.n898 gnd 0.00739f
C3449 vdd.t2 gnd 0.377635f
C3450 vdd.n899 gnd 0.00739f
C3451 vdd.n900 gnd 0.00739f
C3452 vdd.t14 gnd 0.316547f
C3453 vdd.n901 gnd 0.455384f
C3454 vdd.n902 gnd 0.00739f
C3455 vdd.n903 gnd 0.00739f
C3456 vdd.n904 gnd 0.00739f
C3457 vdd.n905 gnd 0.394296f
C3458 vdd.n906 gnd 0.00739f
C3459 vdd.n907 gnd 0.00739f
C3460 vdd.t26 gnd 0.377635f
C3461 vdd.n908 gnd 0.00739f
C3462 vdd.n909 gnd 0.00739f
C3463 vdd.n910 gnd 0.00739f
C3464 vdd.n911 gnd 0.755271f
C3465 vdd.n912 gnd 0.00739f
C3466 vdd.n913 gnd 0.00739f
C3467 vdd.t53 gnd 0.255459f
C3468 vdd.t37 gnd 0.360975f
C3469 vdd.n914 gnd 0.00739f
C3470 vdd.n915 gnd 0.00739f
C3471 vdd.n916 gnd 0.00739f
C3472 vdd.n917 gnd 0.566453f
C3473 vdd.n918 gnd 0.00739f
C3474 vdd.n919 gnd 0.00739f
C3475 vdd.n920 gnd 0.00739f
C3476 vdd.n921 gnd 0.00739f
C3477 vdd.n922 gnd 0.00739f
C3478 vdd.t105 gnd 0.377635f
C3479 vdd.n923 gnd 0.00739f
C3480 vdd.n924 gnd 0.00739f
C3481 vdd.t294 gnd 0.377635f
C3482 vdd.n925 gnd 0.00739f
C3483 vdd.n926 gnd 0.016189f
C3484 vdd.n927 gnd 0.016189f
C3485 vdd.n928 gnd 0.899661f
C3486 vdd.n929 gnd 0.00739f
C3487 vdd.n930 gnd 0.00739f
C3488 vdd.t16 gnd 0.377635f
C3489 vdd.n931 gnd 0.016189f
C3490 vdd.n932 gnd 0.00739f
C3491 vdd.n933 gnd 0.00739f
C3492 vdd.t49 gnd 0.688629f
C3493 vdd.n951 gnd 0.017286f
C3494 vdd.n969 gnd 0.016189f
C3495 vdd.n970 gnd 0.00739f
C3496 vdd.n971 gnd 0.016189f
C3497 vdd.t126 gnd 0.298648f
C3498 vdd.t125 gnd 0.305703f
C3499 vdd.t124 gnd 0.194969f
C3500 vdd.n972 gnd 0.10537f
C3501 vdd.n973 gnd 0.059769f
C3502 vdd.n974 gnd 0.017107f
C3503 vdd.n975 gnd 0.00739f
C3504 vdd.n976 gnd 0.399849f
C3505 vdd.n977 gnd 0.016189f
C3506 vdd.n978 gnd 0.00739f
C3507 vdd.n979 gnd 0.017286f
C3508 vdd.n980 gnd 0.00739f
C3509 vdd.t103 gnd 0.298648f
C3510 vdd.t102 gnd 0.305703f
C3511 vdd.t100 gnd 0.194969f
C3512 vdd.n981 gnd 0.10537f
C3513 vdd.n982 gnd 0.059769f
C3514 vdd.n983 gnd 0.010562f
C3515 vdd.n984 gnd 0.00739f
C3516 vdd.n985 gnd 0.00739f
C3517 vdd.t101 gnd 0.377635f
C3518 vdd.n986 gnd 0.00739f
C3519 vdd.t298 gnd 0.377635f
C3520 vdd.n987 gnd 0.00739f
C3521 vdd.n988 gnd 0.00739f
C3522 vdd.n989 gnd 0.00739f
C3523 vdd.n990 gnd 0.00739f
C3524 vdd.n991 gnd 0.00739f
C3525 vdd.n992 gnd 0.755271f
C3526 vdd.n993 gnd 0.00739f
C3527 vdd.n994 gnd 0.00739f
C3528 vdd.t132 gnd 0.377635f
C3529 vdd.n995 gnd 0.00739f
C3530 vdd.n996 gnd 0.00739f
C3531 vdd.n997 gnd 0.00739f
C3532 vdd.n998 gnd 0.00739f
C3533 vdd.n999 gnd 0.499811f
C3534 vdd.n1000 gnd 0.00739f
C3535 vdd.n1001 gnd 0.00739f
C3536 vdd.n1002 gnd 0.00739f
C3537 vdd.n1003 gnd 0.00739f
C3538 vdd.n1004 gnd 0.00739f
C3539 vdd.n1005 gnd 0.666415f
C3540 vdd.n1006 gnd 0.00739f
C3541 vdd.n1007 gnd 0.00739f
C3542 vdd.t0 gnd 0.360975f
C3543 vdd.t10 gnd 0.255459f
C3544 vdd.n1008 gnd 0.00739f
C3545 vdd.n1009 gnd 0.00739f
C3546 vdd.n1010 gnd 0.00739f
C3547 vdd.t3 gnd 0.377635f
C3548 vdd.n1011 gnd 0.00739f
C3549 vdd.n1012 gnd 0.00739f
C3550 vdd.t47 gnd 0.377635f
C3551 vdd.n1013 gnd 0.00739f
C3552 vdd.n1014 gnd 0.00739f
C3553 vdd.n1015 gnd 0.00739f
C3554 vdd.t12 gnd 0.316547f
C3555 vdd.n1016 gnd 0.00739f
C3556 vdd.n1017 gnd 0.00739f
C3557 vdd.n1018 gnd 0.605327f
C3558 vdd.n1019 gnd 0.00739f
C3559 vdd.n1020 gnd 0.00739f
C3560 vdd.n1021 gnd 0.00739f
C3561 vdd.t5 gnd 0.377635f
C3562 vdd.n1022 gnd 0.00739f
C3563 vdd.n1023 gnd 0.00739f
C3564 vdd.t11 gnd 0.299887f
C3565 vdd.n1024 gnd 0.438723f
C3566 vdd.n1025 gnd 0.00739f
C3567 vdd.n1026 gnd 0.00739f
C3568 vdd.n1027 gnd 0.00739f
C3569 vdd.n1028 gnd 0.649755f
C3570 vdd.n1029 gnd 0.00739f
C3571 vdd.n1030 gnd 0.00739f
C3572 vdd.t9 gnd 0.377635f
C3573 vdd.n1031 gnd 0.00739f
C3574 vdd.n1032 gnd 0.00739f
C3575 vdd.n1033 gnd 0.00739f
C3576 vdd.n1034 gnd 0.755271f
C3577 vdd.n1035 gnd 0.00739f
C3578 vdd.n1036 gnd 0.00739f
C3579 vdd.t18 gnd 0.377635f
C3580 vdd.n1037 gnd 0.00739f
C3581 vdd.n1038 gnd 0.00739f
C3582 vdd.n1039 gnd 0.00739f
C3583 vdd.t31 gnd 0.111069f
C3584 vdd.n1040 gnd 0.00739f
C3585 vdd.n1041 gnd 0.00739f
C3586 vdd.n1042 gnd 0.00739f
C3587 vdd.t113 gnd 0.305703f
C3588 vdd.t111 gnd 0.194969f
C3589 vdd.t114 gnd 0.305703f
C3590 vdd.n1043 gnd 0.171818f
C3591 vdd.n1044 gnd 0.00739f
C3592 vdd.n1045 gnd 0.00739f
C3593 vdd.t8 gnd 0.377635f
C3594 vdd.n1046 gnd 0.00739f
C3595 vdd.n1047 gnd 0.00739f
C3596 vdd.t112 gnd 0.316547f
C3597 vdd.n1048 gnd 0.644201f
C3598 vdd.n1049 gnd 0.00739f
C3599 vdd.n1050 gnd 0.00739f
C3600 vdd.n1051 gnd 0.00739f
C3601 vdd.n1052 gnd 0.394296f
C3602 vdd.n1053 gnd 0.00739f
C3603 vdd.n1054 gnd 0.00739f
C3604 vdd.n1055 gnd 0.527579f
C3605 vdd.n1056 gnd 0.00739f
C3606 vdd.n1057 gnd 0.00739f
C3607 vdd.n1058 gnd 0.00739f
C3608 vdd.n1059 gnd 0.755271f
C3609 vdd.n1060 gnd 0.00739f
C3610 vdd.n1061 gnd 0.00739f
C3611 vdd.t21 gnd 0.377635f
C3612 vdd.n1062 gnd 0.00739f
C3613 vdd.n1063 gnd 0.00739f
C3614 vdd.n1064 gnd 0.00739f
C3615 vdd.n1065 gnd 0.755271f
C3616 vdd.n1066 gnd 0.00739f
C3617 vdd.n1067 gnd 0.00739f
C3618 vdd.n1068 gnd 0.00739f
C3619 vdd.n1069 gnd 0.00739f
C3620 vdd.n1070 gnd 0.00739f
C3621 vdd.t59 gnd 0.377635f
C3622 vdd.n1071 gnd 0.00739f
C3623 vdd.n1072 gnd 0.00739f
C3624 vdd.n1073 gnd 0.00739f
C3625 vdd.n1074 gnd 0.016189f
C3626 vdd.n1075 gnd 0.016189f
C3627 vdd.n1076 gnd 1.06626f
C3628 vdd.n1077 gnd 0.00739f
C3629 vdd.n1078 gnd 0.00739f
C3630 vdd.n1079 gnd 0.494258f
C3631 vdd.n1080 gnd 0.016189f
C3632 vdd.n1081 gnd 0.00739f
C3633 vdd.n1082 gnd 0.00739f
C3634 vdd.n1083 gnd 9.874049f
C3635 vdd.n1116 gnd 0.017286f
C3636 vdd.n1117 gnd 0.00739f
C3637 vdd.n1118 gnd 0.00739f
C3638 vdd.n1119 gnd 0.00739f
C3639 vdd.n1120 gnd 0.006956f
C3640 vdd.n1123 gnd 0.026855f
C3641 vdd.n1124 gnd 0.007261f
C3642 vdd.n1125 gnd 0.008748f
C3643 vdd.n1127 gnd 0.010868f
C3644 vdd.n1128 gnd 0.010868f
C3645 vdd.n1129 gnd 0.008748f
C3646 vdd.n1131 gnd 0.010868f
C3647 vdd.n1132 gnd 0.010868f
C3648 vdd.n1133 gnd 0.010868f
C3649 vdd.n1134 gnd 0.010868f
C3650 vdd.n1135 gnd 0.010868f
C3651 vdd.n1136 gnd 0.008748f
C3652 vdd.n1138 gnd 0.010868f
C3653 vdd.n1139 gnd 0.010868f
C3654 vdd.n1140 gnd 0.010868f
C3655 vdd.n1141 gnd 0.010868f
C3656 vdd.n1142 gnd 0.010868f
C3657 vdd.n1143 gnd 0.008748f
C3658 vdd.n1145 gnd 0.010868f
C3659 vdd.n1146 gnd 0.010868f
C3660 vdd.n1147 gnd 0.010868f
C3661 vdd.n1148 gnd 0.010868f
C3662 vdd.n1149 gnd 0.007304f
C3663 vdd.t120 gnd 0.133709f
C3664 vdd.t119 gnd 0.142898f
C3665 vdd.t118 gnd 0.174622f
C3666 vdd.n1150 gnd 0.223841f
C3667 vdd.n1151 gnd 0.188067f
C3668 vdd.n1153 gnd 0.010868f
C3669 vdd.n1154 gnd 0.010868f
C3670 vdd.n1155 gnd 0.008748f
C3671 vdd.n1156 gnd 0.010868f
C3672 vdd.n1158 gnd 0.010868f
C3673 vdd.n1159 gnd 0.010868f
C3674 vdd.n1160 gnd 0.010868f
C3675 vdd.n1161 gnd 0.010868f
C3676 vdd.n1162 gnd 0.008748f
C3677 vdd.n1164 gnd 0.010868f
C3678 vdd.n1165 gnd 0.010868f
C3679 vdd.n1166 gnd 0.010868f
C3680 vdd.n1167 gnd 0.010868f
C3681 vdd.n1168 gnd 0.010868f
C3682 vdd.n1169 gnd 0.008748f
C3683 vdd.n1171 gnd 0.010868f
C3684 vdd.n1172 gnd 0.010868f
C3685 vdd.n1173 gnd 0.010868f
C3686 vdd.n1174 gnd 0.010868f
C3687 vdd.n1175 gnd 0.010868f
C3688 vdd.n1176 gnd 0.008748f
C3689 vdd.n1178 gnd 0.010868f
C3690 vdd.n1179 gnd 0.010868f
C3691 vdd.n1180 gnd 0.010868f
C3692 vdd.n1181 gnd 0.010868f
C3693 vdd.n1182 gnd 0.010868f
C3694 vdd.n1183 gnd 0.008748f
C3695 vdd.n1185 gnd 0.010868f
C3696 vdd.n1186 gnd 0.010868f
C3697 vdd.n1187 gnd 0.010868f
C3698 vdd.n1188 gnd 0.010868f
C3699 vdd.n1189 gnd 0.00866f
C3700 vdd.t99 gnd 0.133709f
C3701 vdd.t98 gnd 0.142898f
C3702 vdd.t97 gnd 0.174622f
C3703 vdd.n1190 gnd 0.223841f
C3704 vdd.n1191 gnd 0.188067f
C3705 vdd.n1193 gnd 0.010868f
C3706 vdd.n1194 gnd 0.010868f
C3707 vdd.n1195 gnd 0.008748f
C3708 vdd.n1196 gnd 0.010868f
C3709 vdd.n1198 gnd 0.010868f
C3710 vdd.n1199 gnd 0.010868f
C3711 vdd.n1200 gnd 0.010868f
C3712 vdd.n1201 gnd 0.010868f
C3713 vdd.n1202 gnd 0.008748f
C3714 vdd.n1204 gnd 0.010868f
C3715 vdd.n1205 gnd 0.010868f
C3716 vdd.n1206 gnd 0.010868f
C3717 vdd.n1207 gnd 0.010868f
C3718 vdd.n1208 gnd 0.010868f
C3719 vdd.n1209 gnd 0.008748f
C3720 vdd.n1211 gnd 0.010868f
C3721 vdd.n1212 gnd 0.010868f
C3722 vdd.n1213 gnd 0.010868f
C3723 vdd.n1214 gnd 0.010868f
C3724 vdd.n1215 gnd 0.010868f
C3725 vdd.n1216 gnd 0.008748f
C3726 vdd.n1218 gnd 0.010868f
C3727 vdd.n1219 gnd 0.010868f
C3728 vdd.n1220 gnd 0.006956f
C3729 vdd.n1221 gnd 0.008748f
C3730 vdd.n1222 gnd 0.00739f
C3731 vdd.n1223 gnd 0.00739f
C3732 vdd.n1224 gnd 0.00739f
C3733 vdd.n1225 gnd 0.00739f
C3734 vdd.n1226 gnd 0.00739f
C3735 vdd.n1227 gnd 0.00739f
C3736 vdd.n1228 gnd 0.00739f
C3737 vdd.n1229 gnd 0.00739f
C3738 vdd.n1230 gnd 0.00739f
C3739 vdd.n1231 gnd 0.00739f
C3740 vdd.n1232 gnd 0.00739f
C3741 vdd.n1233 gnd 0.00739f
C3742 vdd.n1234 gnd 0.00739f
C3743 vdd.n1235 gnd 0.00739f
C3744 vdd.n1236 gnd 0.00739f
C3745 vdd.n1237 gnd 0.00739f
C3746 vdd.n1238 gnd 0.00739f
C3747 vdd.n1239 gnd 0.00739f
C3748 vdd.n1240 gnd 0.00739f
C3749 vdd.n1241 gnd 0.00739f
C3750 vdd.n1242 gnd 0.00739f
C3751 vdd.n1243 gnd 0.00739f
C3752 vdd.n1244 gnd 0.00739f
C3753 vdd.n1245 gnd 0.00739f
C3754 vdd.n1246 gnd 0.00739f
C3755 vdd.n1247 gnd 0.00739f
C3756 vdd.n1248 gnd 0.00739f
C3757 vdd.n1249 gnd 0.00739f
C3758 vdd.n1250 gnd 0.00739f
C3759 vdd.n1251 gnd 0.00739f
C3760 vdd.n1252 gnd 0.00739f
C3761 vdd.t60 gnd 0.298648f
C3762 vdd.t61 gnd 0.305703f
C3763 vdd.t58 gnd 0.194969f
C3764 vdd.n1253 gnd 0.10537f
C3765 vdd.n1254 gnd 0.059769f
C3766 vdd.n1255 gnd 0.010562f
C3767 vdd.n1256 gnd 0.00739f
C3768 vdd.n1257 gnd 0.00739f
C3769 vdd.n1258 gnd 0.00739f
C3770 vdd.n1259 gnd 0.00739f
C3771 vdd.n1260 gnd 0.00739f
C3772 vdd.n1261 gnd 0.00739f
C3773 vdd.n1262 gnd 0.00739f
C3774 vdd.n1263 gnd 0.00739f
C3775 vdd.n1264 gnd 0.00739f
C3776 vdd.n1265 gnd 0.00739f
C3777 vdd.n1266 gnd 0.00739f
C3778 vdd.n1267 gnd 0.00739f
C3779 vdd.n1268 gnd 0.00739f
C3780 vdd.n1269 gnd 0.00739f
C3781 vdd.n1270 gnd 0.00739f
C3782 vdd.n1271 gnd 0.00739f
C3783 vdd.n1272 gnd 0.00739f
C3784 vdd.t74 gnd 0.298648f
C3785 vdd.t75 gnd 0.305703f
C3786 vdd.t73 gnd 0.194969f
C3787 vdd.n1273 gnd 0.10537f
C3788 vdd.n1274 gnd 0.059769f
C3789 vdd.n1275 gnd 0.00739f
C3790 vdd.n1276 gnd 0.00739f
C3791 vdd.n1277 gnd 0.00739f
C3792 vdd.n1278 gnd 0.00739f
C3793 vdd.n1279 gnd 0.00739f
C3794 vdd.n1280 gnd 0.00739f
C3795 vdd.n1281 gnd 0.00739f
C3796 vdd.n1282 gnd 0.00739f
C3797 vdd.n1283 gnd 0.00739f
C3798 vdd.n1284 gnd 0.00739f
C3799 vdd.n1285 gnd 0.00739f
C3800 vdd.n1286 gnd 0.00739f
C3801 vdd.n1287 gnd 0.00739f
C3802 vdd.n1288 gnd 0.00739f
C3803 vdd.n1289 gnd 0.00739f
C3804 vdd.n1290 gnd 0.00739f
C3805 vdd.n1291 gnd 0.00739f
C3806 vdd.n1292 gnd 0.00739f
C3807 vdd.n1293 gnd 0.00739f
C3808 vdd.n1294 gnd 0.00739f
C3809 vdd.n1295 gnd 0.00739f
C3810 vdd.n1296 gnd 0.00739f
C3811 vdd.n1297 gnd 0.00739f
C3812 vdd.n1298 gnd 0.00739f
C3813 vdd.n1299 gnd 0.00739f
C3814 vdd.n1300 gnd 0.00739f
C3815 vdd.n1301 gnd 0.00538f
C3816 vdd.n1302 gnd 0.010562f
C3817 vdd.n1303 gnd 0.005706f
C3818 vdd.n1304 gnd 0.00739f
C3819 vdd.n1305 gnd 0.00739f
C3820 vdd.n1306 gnd 0.00739f
C3821 vdd.n1307 gnd 0.017286f
C3822 vdd.n1308 gnd 0.017286f
C3823 vdd.n1309 gnd 0.016189f
C3824 vdd.n1310 gnd 0.016189f
C3825 vdd.n1311 gnd 0.00739f
C3826 vdd.n1312 gnd 0.00739f
C3827 vdd.n1313 gnd 0.00739f
C3828 vdd.n1314 gnd 0.00739f
C3829 vdd.n1315 gnd 0.00739f
C3830 vdd.n1316 gnd 0.00739f
C3831 vdd.n1317 gnd 0.00739f
C3832 vdd.n1318 gnd 0.00739f
C3833 vdd.n1319 gnd 0.00739f
C3834 vdd.n1320 gnd 0.00739f
C3835 vdd.n1321 gnd 0.00739f
C3836 vdd.n1322 gnd 0.00739f
C3837 vdd.n1323 gnd 0.00739f
C3838 vdd.n1324 gnd 0.00739f
C3839 vdd.n1325 gnd 0.00739f
C3840 vdd.n1326 gnd 0.00739f
C3841 vdd.n1327 gnd 0.00739f
C3842 vdd.n1328 gnd 0.00739f
C3843 vdd.n1329 gnd 0.00739f
C3844 vdd.n1330 gnd 0.00739f
C3845 vdd.n1331 gnd 0.00739f
C3846 vdd.n1332 gnd 0.00739f
C3847 vdd.n1333 gnd 0.00739f
C3848 vdd.n1334 gnd 0.00739f
C3849 vdd.n1335 gnd 0.00739f
C3850 vdd.n1336 gnd 0.00739f
C3851 vdd.n1337 gnd 0.00739f
C3852 vdd.n1338 gnd 0.44983f
C3853 vdd.n1339 gnd 0.00739f
C3854 vdd.n1340 gnd 0.00739f
C3855 vdd.n1341 gnd 0.00739f
C3856 vdd.n1342 gnd 0.00739f
C3857 vdd.n1343 gnd 0.00739f
C3858 vdd.n1344 gnd 0.00739f
C3859 vdd.n1345 gnd 0.00739f
C3860 vdd.n1346 gnd 0.00739f
C3861 vdd.n1347 gnd 0.00739f
C3862 vdd.n1348 gnd 0.00739f
C3863 vdd.n1349 gnd 0.00739f
C3864 vdd.n1350 gnd 0.00739f
C3865 vdd.n1351 gnd 0.00739f
C3866 vdd.n1352 gnd 0.00739f
C3867 vdd.n1353 gnd 0.00739f
C3868 vdd.n1354 gnd 0.00739f
C3869 vdd.n1355 gnd 0.00739f
C3870 vdd.n1356 gnd 0.00739f
C3871 vdd.n1357 gnd 0.00739f
C3872 vdd.n1358 gnd 0.00739f
C3873 vdd.n1359 gnd 0.238799f
C3874 vdd.n1360 gnd 0.00739f
C3875 vdd.n1361 gnd 0.00739f
C3876 vdd.n1362 gnd 0.00739f
C3877 vdd.n1363 gnd 0.00739f
C3878 vdd.n1364 gnd 0.00739f
C3879 vdd.n1365 gnd 0.00739f
C3880 vdd.n1366 gnd 0.00739f
C3881 vdd.n1367 gnd 0.00739f
C3882 vdd.n1368 gnd 0.00739f
C3883 vdd.n1369 gnd 0.00739f
C3884 vdd.n1370 gnd 0.00739f
C3885 vdd.n1371 gnd 0.00739f
C3886 vdd.n1372 gnd 0.00739f
C3887 vdd.n1373 gnd 0.00739f
C3888 vdd.n1374 gnd 0.00739f
C3889 vdd.n1375 gnd 0.00739f
C3890 vdd.n1376 gnd 0.00739f
C3891 vdd.n1377 gnd 0.00739f
C3892 vdd.n1378 gnd 0.00739f
C3893 vdd.n1379 gnd 0.00739f
C3894 vdd.n1380 gnd 0.00739f
C3895 vdd.n1381 gnd 0.00739f
C3896 vdd.n1382 gnd 0.00739f
C3897 vdd.n1383 gnd 0.00739f
C3898 vdd.n1384 gnd 0.00739f
C3899 vdd.n1385 gnd 0.00739f
C3900 vdd.n1386 gnd 0.00739f
C3901 vdd.n1387 gnd 0.016189f
C3902 vdd.n1388 gnd 0.016189f
C3903 vdd.n1389 gnd 0.017286f
C3904 vdd.n1390 gnd 0.00739f
C3905 vdd.n1391 gnd 0.00739f
C3906 vdd.n1392 gnd 0.005706f
C3907 vdd.n1393 gnd 0.00739f
C3908 vdd.n1394 gnd 0.00739f
C3909 vdd.n1395 gnd 0.00538f
C3910 vdd.n1396 gnd 0.00739f
C3911 vdd.n1397 gnd 0.00739f
C3912 vdd.n1398 gnd 0.00739f
C3913 vdd.n1399 gnd 0.00739f
C3914 vdd.n1400 gnd 0.00739f
C3915 vdd.n1401 gnd 0.00739f
C3916 vdd.n1402 gnd 0.00739f
C3917 vdd.n1403 gnd 0.00739f
C3918 vdd.n1404 gnd 0.00739f
C3919 vdd.n1405 gnd 0.00739f
C3920 vdd.n1406 gnd 0.00739f
C3921 vdd.n1407 gnd 0.00739f
C3922 vdd.n1408 gnd 0.00739f
C3923 vdd.n1409 gnd 0.00739f
C3924 vdd.n1410 gnd 0.00739f
C3925 vdd.n1411 gnd 0.00739f
C3926 vdd.n1412 gnd 0.00739f
C3927 vdd.n1413 gnd 0.00739f
C3928 vdd.n1414 gnd 0.00739f
C3929 vdd.n1415 gnd 0.00739f
C3930 vdd.n1416 gnd 0.00739f
C3931 vdd.n1417 gnd 0.00739f
C3932 vdd.n1418 gnd 0.00739f
C3933 vdd.n1419 gnd 0.00739f
C3934 vdd.n1420 gnd 0.00739f
C3935 vdd.n1421 gnd 0.00739f
C3936 vdd.n1422 gnd 0.029621f
C3937 vdd.n1424 gnd 0.026855f
C3938 vdd.n1425 gnd 0.008748f
C3939 vdd.n1427 gnd 0.010868f
C3940 vdd.n1428 gnd 0.008748f
C3941 vdd.n1429 gnd 0.010868f
C3942 vdd.n1431 gnd 0.010868f
C3943 vdd.n1432 gnd 0.010868f
C3944 vdd.n1434 gnd 0.010868f
C3945 vdd.n1435 gnd 0.007261f
C3946 vdd.t67 gnd 0.555346f
C3947 vdd.n1436 gnd 0.010868f
C3948 vdd.n1437 gnd 0.026855f
C3949 vdd.n1438 gnd 0.008748f
C3950 vdd.n1439 gnd 0.010868f
C3951 vdd.n1440 gnd 0.008748f
C3952 vdd.n1441 gnd 0.010868f
C3953 vdd.n1442 gnd 1.11069f
C3954 vdd.n1443 gnd 0.010868f
C3955 vdd.n1444 gnd 0.008748f
C3956 vdd.n1445 gnd 0.008748f
C3957 vdd.n1446 gnd 0.010868f
C3958 vdd.n1447 gnd 0.008748f
C3959 vdd.n1448 gnd 0.010868f
C3960 vdd.t190 gnd 0.555346f
C3961 vdd.n1449 gnd 0.010868f
C3962 vdd.n1450 gnd 0.008748f
C3963 vdd.n1451 gnd 0.010868f
C3964 vdd.n1452 gnd 0.008748f
C3965 vdd.n1453 gnd 0.010868f
C3966 vdd.t146 gnd 0.555346f
C3967 vdd.n1454 gnd 0.010868f
C3968 vdd.n1455 gnd 0.008748f
C3969 vdd.n1456 gnd 0.010868f
C3970 vdd.n1457 gnd 0.008748f
C3971 vdd.n1458 gnd 0.010868f
C3972 vdd.n1459 gnd 0.894107f
C3973 vdd.n1460 gnd 0.921874f
C3974 vdd.t218 gnd 0.555346f
C3975 vdd.n1461 gnd 0.010868f
C3976 vdd.n1462 gnd 0.008748f
C3977 vdd.n1463 gnd 0.010868f
C3978 vdd.n1464 gnd 0.008748f
C3979 vdd.n1465 gnd 0.010868f
C3980 vdd.n1466 gnd 0.705289f
C3981 vdd.n1467 gnd 0.010868f
C3982 vdd.n1468 gnd 0.008748f
C3983 vdd.n1469 gnd 0.010868f
C3984 vdd.n1470 gnd 0.008748f
C3985 vdd.n1471 gnd 0.010868f
C3986 vdd.t153 gnd 0.555346f
C3987 vdd.t237 gnd 0.555346f
C3988 vdd.n1472 gnd 0.010868f
C3989 vdd.n1473 gnd 0.008748f
C3990 vdd.n1474 gnd 0.010868f
C3991 vdd.n1475 gnd 0.008748f
C3992 vdd.n1476 gnd 0.010868f
C3993 vdd.t206 gnd 0.555346f
C3994 vdd.n1477 gnd 0.010868f
C3995 vdd.n1478 gnd 0.008748f
C3996 vdd.n1479 gnd 0.010868f
C3997 vdd.n1480 gnd 0.008748f
C3998 vdd.n1481 gnd 0.010868f
C3999 vdd.t164 gnd 0.555346f
C4000 vdd.n1482 gnd 0.783038f
C4001 vdd.n1483 gnd 0.010868f
C4002 vdd.n1484 gnd 0.008748f
C4003 vdd.n1485 gnd 0.010868f
C4004 vdd.n1486 gnd 0.008748f
C4005 vdd.n1487 gnd 0.010868f
C4006 vdd.n1488 gnd 0.871893f
C4007 vdd.n1489 gnd 0.010868f
C4008 vdd.n1490 gnd 0.008748f
C4009 vdd.n1491 gnd 0.010868f
C4010 vdd.n1492 gnd 0.008748f
C4011 vdd.n1493 gnd 0.010868f
C4012 vdd.n1494 gnd 0.683076f
C4013 vdd.t171 gnd 0.555346f
C4014 vdd.n1495 gnd 0.010868f
C4015 vdd.n1496 gnd 0.008748f
C4016 vdd.n1497 gnd 0.010868f
C4017 vdd.n1498 gnd 0.008748f
C4018 vdd.n1499 gnd 0.010868f
C4019 vdd.t136 gnd 0.555346f
C4020 vdd.n1500 gnd 0.010868f
C4021 vdd.n1501 gnd 0.008748f
C4022 vdd.n1502 gnd 0.010868f
C4023 vdd.n1503 gnd 0.008748f
C4024 vdd.n1504 gnd 0.010868f
C4025 vdd.t181 gnd 0.555346f
C4026 vdd.n1505 gnd 0.616434f
C4027 vdd.n1506 gnd 0.010868f
C4028 vdd.n1507 gnd 0.008748f
C4029 vdd.n1508 gnd 0.010868f
C4030 vdd.n1509 gnd 0.008748f
C4031 vdd.n1510 gnd 0.010868f
C4032 vdd.t183 gnd 0.555346f
C4033 vdd.n1511 gnd 0.010868f
C4034 vdd.n1512 gnd 0.008748f
C4035 vdd.n1513 gnd 0.010868f
C4036 vdd.n1514 gnd 0.008748f
C4037 vdd.n1515 gnd 0.010868f
C4038 vdd.n1516 gnd 0.849679f
C4039 vdd.n1517 gnd 0.921874f
C4040 vdd.t140 gnd 0.555346f
C4041 vdd.n1518 gnd 0.010868f
C4042 vdd.n1519 gnd 0.008748f
C4043 vdd.n1520 gnd 0.010868f
C4044 vdd.n1521 gnd 0.008748f
C4045 vdd.n1522 gnd 0.010868f
C4046 vdd.n1523 gnd 0.660862f
C4047 vdd.n1524 gnd 0.010868f
C4048 vdd.n1525 gnd 0.008748f
C4049 vdd.n1526 gnd 0.010868f
C4050 vdd.n1527 gnd 0.008748f
C4051 vdd.n1528 gnd 0.010868f
C4052 vdd.t232 gnd 0.555346f
C4053 vdd.t208 gnd 0.555346f
C4054 vdd.n1529 gnd 0.010868f
C4055 vdd.n1530 gnd 0.008748f
C4056 vdd.n1531 gnd 0.010868f
C4057 vdd.n1532 gnd 0.008748f
C4058 vdd.n1533 gnd 0.010868f
C4059 vdd.t134 gnd 0.555346f
C4060 vdd.n1534 gnd 0.010868f
C4061 vdd.n1535 gnd 0.008748f
C4062 vdd.n1536 gnd 0.010868f
C4063 vdd.n1537 gnd 0.008748f
C4064 vdd.n1538 gnd 0.010868f
C4065 vdd.t144 gnd 0.555346f
C4066 vdd.n1539 gnd 0.827466f
C4067 vdd.n1540 gnd 0.010868f
C4068 vdd.n1541 gnd 0.008748f
C4069 vdd.n1542 gnd 0.010868f
C4070 vdd.n1543 gnd 0.008748f
C4071 vdd.n1544 gnd 0.010868f
C4072 vdd.n1545 gnd 1.11069f
C4073 vdd.n1546 gnd 0.010868f
C4074 vdd.n1547 gnd 0.008748f
C4075 vdd.n1548 gnd 0.026291f
C4076 vdd.n1549 gnd 0.007261f
C4077 vdd.n1550 gnd 0.026291f
C4078 vdd.t91 gnd 0.555346f
C4079 vdd.n1551 gnd 0.026291f
C4080 vdd.n1552 gnd 0.007261f
C4081 vdd.n1553 gnd 0.010868f
C4082 vdd.n1554 gnd 0.008748f
C4083 vdd.n1555 gnd 0.010868f
C4084 vdd.n1586 gnd 0.026855f
C4085 vdd.n1587 gnd 1.63827f
C4086 vdd.n1588 gnd 0.010868f
C4087 vdd.n1589 gnd 0.008748f
C4088 vdd.n1590 gnd 0.010868f
C4089 vdd.n1591 gnd 0.010868f
C4090 vdd.n1592 gnd 0.010868f
C4091 vdd.n1593 gnd 0.010868f
C4092 vdd.n1594 gnd 0.010868f
C4093 vdd.n1595 gnd 0.008748f
C4094 vdd.n1596 gnd 0.010868f
C4095 vdd.n1597 gnd 0.010868f
C4096 vdd.n1598 gnd 0.010868f
C4097 vdd.n1599 gnd 0.010868f
C4098 vdd.n1600 gnd 0.010868f
C4099 vdd.n1601 gnd 0.008748f
C4100 vdd.n1602 gnd 0.010868f
C4101 vdd.n1603 gnd 0.010868f
C4102 vdd.n1604 gnd 0.010868f
C4103 vdd.n1605 gnd 0.010868f
C4104 vdd.n1606 gnd 0.010868f
C4105 vdd.n1607 gnd 0.008748f
C4106 vdd.n1608 gnd 0.010868f
C4107 vdd.n1609 gnd 0.010868f
C4108 vdd.n1610 gnd 0.010868f
C4109 vdd.n1611 gnd 0.010868f
C4110 vdd.n1612 gnd 0.010868f
C4111 vdd.t122 gnd 0.133709f
C4112 vdd.t123 gnd 0.142898f
C4113 vdd.t121 gnd 0.174622f
C4114 vdd.n1613 gnd 0.223841f
C4115 vdd.n1614 gnd 0.188942f
C4116 vdd.n1615 gnd 0.01872f
C4117 vdd.n1616 gnd 0.010868f
C4118 vdd.n1617 gnd 0.010868f
C4119 vdd.n1618 gnd 0.010868f
C4120 vdd.n1619 gnd 0.010868f
C4121 vdd.n1620 gnd 0.010868f
C4122 vdd.n1621 gnd 0.008748f
C4123 vdd.n1622 gnd 0.010868f
C4124 vdd.n1623 gnd 0.010868f
C4125 vdd.n1624 gnd 0.010868f
C4126 vdd.n1625 gnd 0.010868f
C4127 vdd.n1626 gnd 0.010868f
C4128 vdd.n1627 gnd 0.008748f
C4129 vdd.n1628 gnd 0.010868f
C4130 vdd.n1629 gnd 0.010868f
C4131 vdd.n1630 gnd 0.010868f
C4132 vdd.n1631 gnd 0.010868f
C4133 vdd.n1632 gnd 0.010868f
C4134 vdd.n1633 gnd 0.008748f
C4135 vdd.n1634 gnd 0.010868f
C4136 vdd.n1635 gnd 0.010868f
C4137 vdd.n1636 gnd 0.010868f
C4138 vdd.n1637 gnd 0.010868f
C4139 vdd.n1638 gnd 0.010868f
C4140 vdd.n1639 gnd 0.008748f
C4141 vdd.n1640 gnd 0.010868f
C4142 vdd.n1641 gnd 0.010868f
C4143 vdd.n1642 gnd 0.010868f
C4144 vdd.n1643 gnd 0.010868f
C4145 vdd.n1644 gnd 0.010868f
C4146 vdd.n1645 gnd 0.008748f
C4147 vdd.n1646 gnd 0.010868f
C4148 vdd.n1647 gnd 0.010868f
C4149 vdd.n1648 gnd 0.010868f
C4150 vdd.n1649 gnd 0.010868f
C4151 vdd.n1650 gnd 0.008748f
C4152 vdd.n1651 gnd 0.010868f
C4153 vdd.n1652 gnd 0.010868f
C4154 vdd.n1653 gnd 0.010868f
C4155 vdd.n1654 gnd 0.010868f
C4156 vdd.n1655 gnd 0.010868f
C4157 vdd.n1656 gnd 0.008748f
C4158 vdd.n1657 gnd 0.010868f
C4159 vdd.n1658 gnd 0.010868f
C4160 vdd.n1659 gnd 0.010868f
C4161 vdd.n1660 gnd 0.010868f
C4162 vdd.n1661 gnd 0.010868f
C4163 vdd.n1662 gnd 0.008748f
C4164 vdd.n1663 gnd 0.010868f
C4165 vdd.n1664 gnd 0.010868f
C4166 vdd.n1665 gnd 0.010868f
C4167 vdd.n1666 gnd 0.010868f
C4168 vdd.n1667 gnd 0.010868f
C4169 vdd.n1668 gnd 0.008748f
C4170 vdd.n1669 gnd 0.010868f
C4171 vdd.n1670 gnd 0.010868f
C4172 vdd.n1671 gnd 0.010868f
C4173 vdd.n1672 gnd 0.010868f
C4174 vdd.n1673 gnd 0.010868f
C4175 vdd.n1674 gnd 0.008748f
C4176 vdd.n1675 gnd 0.010868f
C4177 vdd.n1676 gnd 0.010868f
C4178 vdd.n1677 gnd 0.010868f
C4179 vdd.n1678 gnd 0.010868f
C4180 vdd.t92 gnd 0.133709f
C4181 vdd.t93 gnd 0.142898f
C4182 vdd.t90 gnd 0.174622f
C4183 vdd.n1679 gnd 0.223841f
C4184 vdd.n1680 gnd 0.188942f
C4185 vdd.n1681 gnd 0.014346f
C4186 vdd.n1682 gnd 0.004155f
C4187 vdd.n1683 gnd 0.026855f
C4188 vdd.n1684 gnd 0.010868f
C4189 vdd.n1685 gnd 0.004593f
C4190 vdd.n1686 gnd 0.008748f
C4191 vdd.n1687 gnd 0.008748f
C4192 vdd.n1688 gnd 0.010868f
C4193 vdd.n1689 gnd 0.010868f
C4194 vdd.n1690 gnd 0.010868f
C4195 vdd.n1691 gnd 0.008748f
C4196 vdd.n1692 gnd 0.008748f
C4197 vdd.n1693 gnd 0.008748f
C4198 vdd.n1694 gnd 0.010868f
C4199 vdd.n1695 gnd 0.010868f
C4200 vdd.n1696 gnd 0.010868f
C4201 vdd.n1697 gnd 0.008748f
C4202 vdd.n1698 gnd 0.008748f
C4203 vdd.n1699 gnd 0.008748f
C4204 vdd.n1700 gnd 0.010868f
C4205 vdd.n1701 gnd 0.010868f
C4206 vdd.n1702 gnd 0.010868f
C4207 vdd.n1703 gnd 0.008748f
C4208 vdd.n1704 gnd 0.008748f
C4209 vdd.n1705 gnd 0.008748f
C4210 vdd.n1706 gnd 0.010868f
C4211 vdd.n1707 gnd 0.010868f
C4212 vdd.n1708 gnd 0.010868f
C4213 vdd.n1709 gnd 0.008748f
C4214 vdd.n1710 gnd 0.008748f
C4215 vdd.n1711 gnd 0.008748f
C4216 vdd.n1712 gnd 0.010868f
C4217 vdd.n1713 gnd 0.010868f
C4218 vdd.n1714 gnd 0.010868f
C4219 vdd.n1715 gnd 0.00866f
C4220 vdd.n1716 gnd 0.010868f
C4221 vdd.t109 gnd 0.133709f
C4222 vdd.t110 gnd 0.142898f
C4223 vdd.t108 gnd 0.174622f
C4224 vdd.n1717 gnd 0.223841f
C4225 vdd.n1718 gnd 0.188942f
C4226 vdd.n1719 gnd 0.01872f
C4227 vdd.n1720 gnd 0.005948f
C4228 vdd.n1721 gnd 0.010868f
C4229 vdd.n1722 gnd 0.010868f
C4230 vdd.n1723 gnd 0.010868f
C4231 vdd.n1724 gnd 0.008748f
C4232 vdd.n1725 gnd 0.008748f
C4233 vdd.n1726 gnd 0.008748f
C4234 vdd.n1727 gnd 0.010868f
C4235 vdd.n1728 gnd 0.010868f
C4236 vdd.n1729 gnd 0.010868f
C4237 vdd.n1730 gnd 0.008748f
C4238 vdd.n1731 gnd 0.008748f
C4239 vdd.n1732 gnd 0.008748f
C4240 vdd.n1733 gnd 0.010868f
C4241 vdd.n1734 gnd 0.010868f
C4242 vdd.n1735 gnd 0.010868f
C4243 vdd.n1736 gnd 0.008748f
C4244 vdd.n1737 gnd 0.008748f
C4245 vdd.n1738 gnd 0.008748f
C4246 vdd.n1739 gnd 0.010868f
C4247 vdd.n1740 gnd 0.010868f
C4248 vdd.n1741 gnd 0.010868f
C4249 vdd.n1742 gnd 0.008748f
C4250 vdd.n1743 gnd 0.008748f
C4251 vdd.n1744 gnd 0.008748f
C4252 vdd.n1745 gnd 0.010868f
C4253 vdd.n1746 gnd 0.010868f
C4254 vdd.n1747 gnd 0.010868f
C4255 vdd.n1748 gnd 0.008748f
C4256 vdd.n1749 gnd 0.008748f
C4257 vdd.n1750 gnd 0.007304f
C4258 vdd.n1751 gnd 0.010868f
C4259 vdd.n1752 gnd 0.010868f
C4260 vdd.n1753 gnd 0.010868f
C4261 vdd.n1754 gnd 0.007304f
C4262 vdd.n1755 gnd 0.008748f
C4263 vdd.n1756 gnd 0.008748f
C4264 vdd.n1757 gnd 0.010868f
C4265 vdd.n1758 gnd 0.010868f
C4266 vdd.n1759 gnd 0.010868f
C4267 vdd.n1760 gnd 0.008748f
C4268 vdd.n1761 gnd 0.008748f
C4269 vdd.n1762 gnd 0.008748f
C4270 vdd.n1763 gnd 0.010868f
C4271 vdd.n1764 gnd 0.010868f
C4272 vdd.n1765 gnd 0.010868f
C4273 vdd.n1766 gnd 0.008748f
C4274 vdd.n1767 gnd 0.008748f
C4275 vdd.n1768 gnd 0.008748f
C4276 vdd.n1769 gnd 0.010868f
C4277 vdd.n1770 gnd 0.010868f
C4278 vdd.n1771 gnd 0.010868f
C4279 vdd.n1772 gnd 0.008748f
C4280 vdd.n1773 gnd 0.008748f
C4281 vdd.n1774 gnd 0.008748f
C4282 vdd.n1775 gnd 0.010868f
C4283 vdd.n1776 gnd 0.010868f
C4284 vdd.n1777 gnd 0.010868f
C4285 vdd.n1778 gnd 0.008748f
C4286 vdd.n1779 gnd 0.010868f
C4287 vdd.n1780 gnd 2.63234f
C4288 vdd.n1782 gnd 0.026855f
C4289 vdd.n1783 gnd 0.007261f
C4290 vdd.n1784 gnd 0.026855f
C4291 vdd.n1785 gnd 0.026291f
C4292 vdd.n1786 gnd 0.010868f
C4293 vdd.n1787 gnd 0.008748f
C4294 vdd.n1788 gnd 0.010868f
C4295 vdd.n1789 gnd 0.560899f
C4296 vdd.n1790 gnd 0.010868f
C4297 vdd.n1791 gnd 0.008748f
C4298 vdd.n1792 gnd 0.010868f
C4299 vdd.n1793 gnd 0.010868f
C4300 vdd.n1794 gnd 0.010868f
C4301 vdd.n1795 gnd 0.008748f
C4302 vdd.n1796 gnd 0.010868f
C4303 vdd.n1797 gnd 1.01628f
C4304 vdd.n1798 gnd 1.11069f
C4305 vdd.n1799 gnd 0.010868f
C4306 vdd.n1800 gnd 0.008748f
C4307 vdd.n1801 gnd 0.010868f
C4308 vdd.n1802 gnd 0.010868f
C4309 vdd.n1803 gnd 0.010868f
C4310 vdd.n1804 gnd 0.008748f
C4311 vdd.n1805 gnd 0.010868f
C4312 vdd.n1806 gnd 0.649755f
C4313 vdd.n1807 gnd 0.010868f
C4314 vdd.n1808 gnd 0.008748f
C4315 vdd.n1809 gnd 0.010868f
C4316 vdd.n1810 gnd 0.010868f
C4317 vdd.n1811 gnd 0.010868f
C4318 vdd.n1812 gnd 0.008748f
C4319 vdd.n1813 gnd 0.010868f
C4320 vdd.n1814 gnd 0.638648f
C4321 vdd.n1815 gnd 0.838572f
C4322 vdd.n1816 gnd 0.010868f
C4323 vdd.n1817 gnd 0.008748f
C4324 vdd.n1818 gnd 0.010868f
C4325 vdd.n1819 gnd 0.010868f
C4326 vdd.n1820 gnd 0.010868f
C4327 vdd.n1821 gnd 0.008748f
C4328 vdd.n1822 gnd 0.010868f
C4329 vdd.n1823 gnd 0.921874f
C4330 vdd.n1824 gnd 0.010868f
C4331 vdd.n1825 gnd 0.008748f
C4332 vdd.n1826 gnd 0.010868f
C4333 vdd.n1827 gnd 0.010868f
C4334 vdd.n1828 gnd 0.010868f
C4335 vdd.n1829 gnd 0.008748f
C4336 vdd.n1830 gnd 0.010868f
C4337 vdd.t148 gnd 0.555346f
C4338 vdd.n1831 gnd 0.816359f
C4339 vdd.n1832 gnd 0.010868f
C4340 vdd.n1833 gnd 0.008748f
C4341 vdd.n1834 gnd 0.010868f
C4342 vdd.n1835 gnd 0.010868f
C4343 vdd.n1836 gnd 0.010868f
C4344 vdd.n1837 gnd 0.008748f
C4345 vdd.n1838 gnd 0.010868f
C4346 vdd.n1839 gnd 0.627541f
C4347 vdd.n1840 gnd 0.010868f
C4348 vdd.n1841 gnd 0.008748f
C4349 vdd.n1842 gnd 0.010868f
C4350 vdd.n1843 gnd 0.010868f
C4351 vdd.n1844 gnd 0.010868f
C4352 vdd.n1845 gnd 0.008748f
C4353 vdd.n1846 gnd 0.010868f
C4354 vdd.n1847 gnd 0.805252f
C4355 vdd.n1848 gnd 0.671969f
C4356 vdd.n1849 gnd 0.010868f
C4357 vdd.n1850 gnd 0.008748f
C4358 vdd.n1851 gnd 0.010868f
C4359 vdd.n1852 gnd 0.010868f
C4360 vdd.n1853 gnd 0.010868f
C4361 vdd.n1854 gnd 0.008748f
C4362 vdd.n1855 gnd 0.010868f
C4363 vdd.n1856 gnd 0.860786f
C4364 vdd.n1857 gnd 0.010868f
C4365 vdd.n1858 gnd 0.008748f
C4366 vdd.n1859 gnd 0.010868f
C4367 vdd.n1860 gnd 0.010868f
C4368 vdd.n1861 gnd 0.010868f
C4369 vdd.n1862 gnd 0.008748f
C4370 vdd.n1863 gnd 0.010868f
C4371 vdd.t234 gnd 0.555346f
C4372 vdd.n1864 gnd 0.921874f
C4373 vdd.n1865 gnd 0.010868f
C4374 vdd.n1866 gnd 0.008748f
C4375 vdd.n1867 gnd 0.010868f
C4376 vdd.n1868 gnd 0.008353f
C4377 vdd.n1869 gnd 0.005965f
C4378 vdd.n1870 gnd 0.005535f
C4379 vdd.n1871 gnd 0.003062f
C4380 vdd.n1872 gnd 0.00703f
C4381 vdd.n1873 gnd 0.002974f
C4382 vdd.n1874 gnd 0.003149f
C4383 vdd.n1875 gnd 0.005535f
C4384 vdd.n1876 gnd 0.002974f
C4385 vdd.n1877 gnd 0.00703f
C4386 vdd.n1878 gnd 0.003149f
C4387 vdd.n1879 gnd 0.005535f
C4388 vdd.n1880 gnd 0.002974f
C4389 vdd.n1881 gnd 0.005272f
C4390 vdd.n1882 gnd 0.005288f
C4391 vdd.t191 gnd 0.015103f
C4392 vdd.n1883 gnd 0.033604f
C4393 vdd.n1884 gnd 0.174886f
C4394 vdd.n1885 gnd 0.002974f
C4395 vdd.n1886 gnd 0.003149f
C4396 vdd.n1887 gnd 0.00703f
C4397 vdd.n1888 gnd 0.00703f
C4398 vdd.n1889 gnd 0.003149f
C4399 vdd.n1890 gnd 0.002974f
C4400 vdd.n1891 gnd 0.005535f
C4401 vdd.n1892 gnd 0.005535f
C4402 vdd.n1893 gnd 0.002974f
C4403 vdd.n1894 gnd 0.003149f
C4404 vdd.n1895 gnd 0.00703f
C4405 vdd.n1896 gnd 0.00703f
C4406 vdd.n1897 gnd 0.003149f
C4407 vdd.n1898 gnd 0.002974f
C4408 vdd.n1899 gnd 0.005535f
C4409 vdd.n1900 gnd 0.005535f
C4410 vdd.n1901 gnd 0.002974f
C4411 vdd.n1902 gnd 0.003149f
C4412 vdd.n1903 gnd 0.00703f
C4413 vdd.n1904 gnd 0.00703f
C4414 vdd.n1905 gnd 0.01662f
C4415 vdd.n1906 gnd 0.003062f
C4416 vdd.n1907 gnd 0.002974f
C4417 vdd.n1908 gnd 0.014306f
C4418 vdd.n1909 gnd 0.009988f
C4419 vdd.t219 gnd 0.034991f
C4420 vdd.t273 gnd 0.034991f
C4421 vdd.n1910 gnd 0.240481f
C4422 vdd.n1911 gnd 0.189101f
C4423 vdd.t238 gnd 0.034991f
C4424 vdd.t287 gnd 0.034991f
C4425 vdd.n1912 gnd 0.240481f
C4426 vdd.n1913 gnd 0.152604f
C4427 vdd.t207 gnd 0.034991f
C4428 vdd.t154 gnd 0.034991f
C4429 vdd.n1914 gnd 0.240481f
C4430 vdd.n1915 gnd 0.152604f
C4431 vdd.t229 gnd 0.034991f
C4432 vdd.t165 gnd 0.034991f
C4433 vdd.n1916 gnd 0.240481f
C4434 vdd.n1917 gnd 0.152604f
C4435 vdd.t277 gnd 0.034991f
C4436 vdd.t292 gnd 0.034991f
C4437 vdd.n1918 gnd 0.240481f
C4438 vdd.n1919 gnd 0.152604f
C4439 vdd.t249 gnd 0.034991f
C4440 vdd.t137 gnd 0.034991f
C4441 vdd.n1920 gnd 0.240481f
C4442 vdd.n1921 gnd 0.152604f
C4443 vdd.t239 gnd 0.034991f
C4444 vdd.t184 gnd 0.034991f
C4445 vdd.n1922 gnd 0.240481f
C4446 vdd.n1923 gnd 0.152604f
C4447 vdd.t281 gnd 0.034991f
C4448 vdd.t213 gnd 0.034991f
C4449 vdd.n1924 gnd 0.240481f
C4450 vdd.n1925 gnd 0.152604f
C4451 vdd.t259 gnd 0.034991f
C4452 vdd.t233 gnd 0.034991f
C4453 vdd.n1926 gnd 0.240481f
C4454 vdd.n1927 gnd 0.152604f
C4455 vdd.n1928 gnd 0.005965f
C4456 vdd.n1929 gnd 0.005535f
C4457 vdd.n1930 gnd 0.003062f
C4458 vdd.n1931 gnd 0.00703f
C4459 vdd.n1932 gnd 0.002974f
C4460 vdd.n1933 gnd 0.003149f
C4461 vdd.n1934 gnd 0.005535f
C4462 vdd.n1935 gnd 0.002974f
C4463 vdd.n1936 gnd 0.00703f
C4464 vdd.n1937 gnd 0.003149f
C4465 vdd.n1938 gnd 0.005535f
C4466 vdd.n1939 gnd 0.002974f
C4467 vdd.n1940 gnd 0.005272f
C4468 vdd.n1941 gnd 0.005288f
C4469 vdd.t196 gnd 0.015103f
C4470 vdd.n1942 gnd 0.033604f
C4471 vdd.n1943 gnd 0.174886f
C4472 vdd.n1944 gnd 0.002974f
C4473 vdd.n1945 gnd 0.003149f
C4474 vdd.n1946 gnd 0.00703f
C4475 vdd.n1947 gnd 0.00703f
C4476 vdd.n1948 gnd 0.003149f
C4477 vdd.n1949 gnd 0.002974f
C4478 vdd.n1950 gnd 0.005535f
C4479 vdd.n1951 gnd 0.005535f
C4480 vdd.n1952 gnd 0.002974f
C4481 vdd.n1953 gnd 0.003149f
C4482 vdd.n1954 gnd 0.00703f
C4483 vdd.n1955 gnd 0.00703f
C4484 vdd.n1956 gnd 0.003149f
C4485 vdd.n1957 gnd 0.002974f
C4486 vdd.n1958 gnd 0.005535f
C4487 vdd.n1959 gnd 0.005535f
C4488 vdd.n1960 gnd 0.002974f
C4489 vdd.n1961 gnd 0.003149f
C4490 vdd.n1962 gnd 0.00703f
C4491 vdd.n1963 gnd 0.00703f
C4492 vdd.n1964 gnd 0.01662f
C4493 vdd.n1965 gnd 0.003062f
C4494 vdd.n1966 gnd 0.002974f
C4495 vdd.n1967 gnd 0.014306f
C4496 vdd.n1968 gnd 0.009674f
C4497 vdd.n1969 gnd 0.113538f
C4498 vdd.n1970 gnd 0.005965f
C4499 vdd.n1971 gnd 0.005535f
C4500 vdd.n1972 gnd 0.003062f
C4501 vdd.n1973 gnd 0.00703f
C4502 vdd.n1974 gnd 0.002974f
C4503 vdd.n1975 gnd 0.003149f
C4504 vdd.n1976 gnd 0.005535f
C4505 vdd.n1977 gnd 0.002974f
C4506 vdd.n1978 gnd 0.00703f
C4507 vdd.n1979 gnd 0.003149f
C4508 vdd.n1980 gnd 0.005535f
C4509 vdd.n1981 gnd 0.002974f
C4510 vdd.n1982 gnd 0.005272f
C4511 vdd.n1983 gnd 0.005288f
C4512 vdd.t271 gnd 0.015103f
C4513 vdd.n1984 gnd 0.033604f
C4514 vdd.n1985 gnd 0.174886f
C4515 vdd.n1986 gnd 0.002974f
C4516 vdd.n1987 gnd 0.003149f
C4517 vdd.n1988 gnd 0.00703f
C4518 vdd.n1989 gnd 0.00703f
C4519 vdd.n1990 gnd 0.003149f
C4520 vdd.n1991 gnd 0.002974f
C4521 vdd.n1992 gnd 0.005535f
C4522 vdd.n1993 gnd 0.005535f
C4523 vdd.n1994 gnd 0.002974f
C4524 vdd.n1995 gnd 0.003149f
C4525 vdd.n1996 gnd 0.00703f
C4526 vdd.n1997 gnd 0.00703f
C4527 vdd.n1998 gnd 0.003149f
C4528 vdd.n1999 gnd 0.002974f
C4529 vdd.n2000 gnd 0.005535f
C4530 vdd.n2001 gnd 0.005535f
C4531 vdd.n2002 gnd 0.002974f
C4532 vdd.n2003 gnd 0.003149f
C4533 vdd.n2004 gnd 0.00703f
C4534 vdd.n2005 gnd 0.00703f
C4535 vdd.n2006 gnd 0.01662f
C4536 vdd.n2007 gnd 0.003062f
C4537 vdd.n2008 gnd 0.002974f
C4538 vdd.n2009 gnd 0.014306f
C4539 vdd.n2010 gnd 0.009988f
C4540 vdd.t223 gnd 0.034991f
C4541 vdd.t147 gnd 0.034991f
C4542 vdd.n2011 gnd 0.240481f
C4543 vdd.n2012 gnd 0.189101f
C4544 vdd.t283 gnd 0.034991f
C4545 vdd.t251 gnd 0.034991f
C4546 vdd.n2013 gnd 0.240481f
C4547 vdd.n2014 gnd 0.152604f
C4548 vdd.t245 gnd 0.034991f
C4549 vdd.t192 gnd 0.034991f
C4550 vdd.n2015 gnd 0.240481f
C4551 vdd.n2016 gnd 0.152604f
C4552 vdd.t186 gnd 0.034991f
C4553 vdd.t246 gnd 0.034991f
C4554 vdd.n2017 gnd 0.240481f
C4555 vdd.n2018 gnd 0.152604f
C4556 vdd.t235 gnd 0.034991f
C4557 vdd.t172 gnd 0.034991f
C4558 vdd.n2019 gnd 0.240481f
C4559 vdd.n2020 gnd 0.152604f
C4560 vdd.t182 gnd 0.034991f
C4561 vdd.t152 gnd 0.034991f
C4562 vdd.n2021 gnd 0.240481f
C4563 vdd.n2022 gnd 0.152604f
C4564 vdd.t141 gnd 0.034991f
C4565 vdd.t230 gnd 0.034991f
C4566 vdd.n2023 gnd 0.240481f
C4567 vdd.n2024 gnd 0.152604f
C4568 vdd.t209 gnd 0.034991f
C4569 vdd.t149 gnd 0.034991f
C4570 vdd.n2025 gnd 0.240481f
C4571 vdd.n2026 gnd 0.152604f
C4572 vdd.t135 gnd 0.034991f
C4573 vdd.t252 gnd 0.034991f
C4574 vdd.n2027 gnd 0.240481f
C4575 vdd.n2028 gnd 0.152604f
C4576 vdd.n2029 gnd 0.005965f
C4577 vdd.n2030 gnd 0.005535f
C4578 vdd.n2031 gnd 0.003062f
C4579 vdd.n2032 gnd 0.00703f
C4580 vdd.n2033 gnd 0.002974f
C4581 vdd.n2034 gnd 0.003149f
C4582 vdd.n2035 gnd 0.005535f
C4583 vdd.n2036 gnd 0.002974f
C4584 vdd.n2037 gnd 0.00703f
C4585 vdd.n2038 gnd 0.003149f
C4586 vdd.n2039 gnd 0.005535f
C4587 vdd.n2040 gnd 0.002974f
C4588 vdd.n2041 gnd 0.005272f
C4589 vdd.n2042 gnd 0.005288f
C4590 vdd.t145 gnd 0.015103f
C4591 vdd.n2043 gnd 0.033604f
C4592 vdd.n2044 gnd 0.174886f
C4593 vdd.n2045 gnd 0.002974f
C4594 vdd.n2046 gnd 0.003149f
C4595 vdd.n2047 gnd 0.00703f
C4596 vdd.n2048 gnd 0.00703f
C4597 vdd.n2049 gnd 0.003149f
C4598 vdd.n2050 gnd 0.002974f
C4599 vdd.n2051 gnd 0.005535f
C4600 vdd.n2052 gnd 0.005535f
C4601 vdd.n2053 gnd 0.002974f
C4602 vdd.n2054 gnd 0.003149f
C4603 vdd.n2055 gnd 0.00703f
C4604 vdd.n2056 gnd 0.00703f
C4605 vdd.n2057 gnd 0.003149f
C4606 vdd.n2058 gnd 0.002974f
C4607 vdd.n2059 gnd 0.005535f
C4608 vdd.n2060 gnd 0.005535f
C4609 vdd.n2061 gnd 0.002974f
C4610 vdd.n2062 gnd 0.003149f
C4611 vdd.n2063 gnd 0.00703f
C4612 vdd.n2064 gnd 0.00703f
C4613 vdd.n2065 gnd 0.01662f
C4614 vdd.n2066 gnd 0.003062f
C4615 vdd.n2067 gnd 0.002974f
C4616 vdd.n2068 gnd 0.014306f
C4617 vdd.n2069 gnd 0.009674f
C4618 vdd.n2070 gnd 0.067544f
C4619 vdd.n2071 gnd 0.243377f
C4620 vdd.n2072 gnd 0.005965f
C4621 vdd.n2073 gnd 0.005535f
C4622 vdd.n2074 gnd 0.003062f
C4623 vdd.n2075 gnd 0.00703f
C4624 vdd.n2076 gnd 0.002974f
C4625 vdd.n2077 gnd 0.003149f
C4626 vdd.n2078 gnd 0.005535f
C4627 vdd.n2079 gnd 0.002974f
C4628 vdd.n2080 gnd 0.00703f
C4629 vdd.n2081 gnd 0.003149f
C4630 vdd.n2082 gnd 0.005535f
C4631 vdd.n2083 gnd 0.002974f
C4632 vdd.n2084 gnd 0.005272f
C4633 vdd.n2085 gnd 0.005288f
C4634 vdd.t282 gnd 0.015103f
C4635 vdd.n2086 gnd 0.033604f
C4636 vdd.n2087 gnd 0.174886f
C4637 vdd.n2088 gnd 0.002974f
C4638 vdd.n2089 gnd 0.003149f
C4639 vdd.n2090 gnd 0.00703f
C4640 vdd.n2091 gnd 0.00703f
C4641 vdd.n2092 gnd 0.003149f
C4642 vdd.n2093 gnd 0.002974f
C4643 vdd.n2094 gnd 0.005535f
C4644 vdd.n2095 gnd 0.005535f
C4645 vdd.n2096 gnd 0.002974f
C4646 vdd.n2097 gnd 0.003149f
C4647 vdd.n2098 gnd 0.00703f
C4648 vdd.n2099 gnd 0.00703f
C4649 vdd.n2100 gnd 0.003149f
C4650 vdd.n2101 gnd 0.002974f
C4651 vdd.n2102 gnd 0.005535f
C4652 vdd.n2103 gnd 0.005535f
C4653 vdd.n2104 gnd 0.002974f
C4654 vdd.n2105 gnd 0.003149f
C4655 vdd.n2106 gnd 0.00703f
C4656 vdd.n2107 gnd 0.00703f
C4657 vdd.n2108 gnd 0.01662f
C4658 vdd.n2109 gnd 0.003062f
C4659 vdd.n2110 gnd 0.002974f
C4660 vdd.n2111 gnd 0.014306f
C4661 vdd.n2112 gnd 0.009988f
C4662 vdd.t236 gnd 0.034991f
C4663 vdd.t177 gnd 0.034991f
C4664 vdd.n2113 gnd 0.240481f
C4665 vdd.n2114 gnd 0.189101f
C4666 vdd.t293 gnd 0.034991f
C4667 vdd.t265 gnd 0.034991f
C4668 vdd.n2115 gnd 0.240481f
C4669 vdd.n2116 gnd 0.152604f
C4670 vdd.t261 gnd 0.034991f
C4671 vdd.t214 gnd 0.034991f
C4672 vdd.n2117 gnd 0.240481f
C4673 vdd.n2118 gnd 0.152604f
C4674 vdd.t210 gnd 0.034991f
C4675 vdd.t264 gnd 0.034991f
C4676 vdd.n2119 gnd 0.240481f
C4677 vdd.n2120 gnd 0.152604f
C4678 vdd.t244 gnd 0.034991f
C4679 vdd.t243 gnd 0.034991f
C4680 vdd.n2121 gnd 0.240481f
C4681 vdd.n2122 gnd 0.152604f
C4682 vdd.t205 gnd 0.034991f
C4683 vdd.t178 gnd 0.034991f
C4684 vdd.n2123 gnd 0.240481f
C4685 vdd.n2124 gnd 0.152604f
C4686 vdd.t169 gnd 0.034991f
C4687 vdd.t242 gnd 0.034991f
C4688 vdd.n2125 gnd 0.240481f
C4689 vdd.n2126 gnd 0.152604f
C4690 vdd.t225 gnd 0.034991f
C4691 vdd.t170 gnd 0.034991f
C4692 vdd.n2127 gnd 0.240481f
C4693 vdd.n2128 gnd 0.152604f
C4694 vdd.t163 gnd 0.034991f
C4695 vdd.t266 gnd 0.034991f
C4696 vdd.n2129 gnd 0.240481f
C4697 vdd.n2130 gnd 0.152604f
C4698 vdd.n2131 gnd 0.005965f
C4699 vdd.n2132 gnd 0.005535f
C4700 vdd.n2133 gnd 0.003062f
C4701 vdd.n2134 gnd 0.00703f
C4702 vdd.n2135 gnd 0.002974f
C4703 vdd.n2136 gnd 0.003149f
C4704 vdd.n2137 gnd 0.005535f
C4705 vdd.n2138 gnd 0.002974f
C4706 vdd.n2139 gnd 0.00703f
C4707 vdd.n2140 gnd 0.003149f
C4708 vdd.n2141 gnd 0.005535f
C4709 vdd.n2142 gnd 0.002974f
C4710 vdd.n2143 gnd 0.005272f
C4711 vdd.n2144 gnd 0.005288f
C4712 vdd.t220 gnd 0.015103f
C4713 vdd.n2145 gnd 0.033604f
C4714 vdd.n2146 gnd 0.174886f
C4715 vdd.n2147 gnd 0.002974f
C4716 vdd.n2148 gnd 0.003149f
C4717 vdd.n2149 gnd 0.00703f
C4718 vdd.n2150 gnd 0.00703f
C4719 vdd.n2151 gnd 0.003149f
C4720 vdd.n2152 gnd 0.002974f
C4721 vdd.n2153 gnd 0.005535f
C4722 vdd.n2154 gnd 0.005535f
C4723 vdd.n2155 gnd 0.002974f
C4724 vdd.n2156 gnd 0.003149f
C4725 vdd.n2157 gnd 0.00703f
C4726 vdd.n2158 gnd 0.00703f
C4727 vdd.n2159 gnd 0.003149f
C4728 vdd.n2160 gnd 0.002974f
C4729 vdd.n2161 gnd 0.005535f
C4730 vdd.n2162 gnd 0.005535f
C4731 vdd.n2163 gnd 0.002974f
C4732 vdd.n2164 gnd 0.003149f
C4733 vdd.n2165 gnd 0.00703f
C4734 vdd.n2166 gnd 0.00703f
C4735 vdd.n2167 gnd 0.01662f
C4736 vdd.n2168 gnd 0.003062f
C4737 vdd.n2169 gnd 0.002974f
C4738 vdd.n2170 gnd 0.014306f
C4739 vdd.n2171 gnd 0.009674f
C4740 vdd.n2172 gnd 0.067544f
C4741 vdd.n2173 gnd 0.278614f
C4742 vdd.n2174 gnd 2.92276f
C4743 vdd.n2175 gnd 0.641055f
C4744 vdd.n2176 gnd 0.008353f
C4745 vdd.n2177 gnd 0.008748f
C4746 vdd.n2178 gnd 0.010868f
C4747 vdd.n2179 gnd 0.794145f
C4748 vdd.n2180 gnd 0.010868f
C4749 vdd.n2181 gnd 0.008748f
C4750 vdd.n2182 gnd 0.010868f
C4751 vdd.n2183 gnd 0.010868f
C4752 vdd.n2184 gnd 0.010868f
C4753 vdd.n2185 gnd 0.008748f
C4754 vdd.n2186 gnd 0.010868f
C4755 vdd.n2187 gnd 0.921874f
C4756 vdd.t185 gnd 0.555346f
C4757 vdd.n2188 gnd 0.605327f
C4758 vdd.n2189 gnd 0.010868f
C4759 vdd.n2190 gnd 0.008748f
C4760 vdd.n2191 gnd 0.010868f
C4761 vdd.n2192 gnd 0.010868f
C4762 vdd.n2193 gnd 0.010868f
C4763 vdd.n2194 gnd 0.008748f
C4764 vdd.n2195 gnd 0.010868f
C4765 vdd.n2196 gnd 0.694182f
C4766 vdd.n2197 gnd 0.010868f
C4767 vdd.n2198 gnd 0.008748f
C4768 vdd.n2199 gnd 0.010868f
C4769 vdd.n2200 gnd 0.010868f
C4770 vdd.n2201 gnd 0.010868f
C4771 vdd.n2202 gnd 0.008748f
C4772 vdd.n2203 gnd 0.010868f
C4773 vdd.n2204 gnd 0.59422f
C4774 vdd.n2205 gnd 0.883f
C4775 vdd.n2206 gnd 0.010868f
C4776 vdd.n2207 gnd 0.008748f
C4777 vdd.n2208 gnd 0.010868f
C4778 vdd.n2209 gnd 0.010868f
C4779 vdd.n2210 gnd 0.010868f
C4780 vdd.n2211 gnd 0.008748f
C4781 vdd.n2212 gnd 0.010868f
C4782 vdd.n2213 gnd 0.921874f
C4783 vdd.n2214 gnd 0.010868f
C4784 vdd.n2215 gnd 0.008748f
C4785 vdd.n2216 gnd 0.010868f
C4786 vdd.n2217 gnd 0.010868f
C4787 vdd.n2218 gnd 0.010868f
C4788 vdd.n2219 gnd 0.008748f
C4789 vdd.n2220 gnd 0.010868f
C4790 vdd.t250 gnd 0.555346f
C4791 vdd.n2221 gnd 0.771931f
C4792 vdd.n2222 gnd 0.010868f
C4793 vdd.n2223 gnd 0.008748f
C4794 vdd.n2224 gnd 0.010868f
C4795 vdd.n2225 gnd 0.010868f
C4796 vdd.n2226 gnd 0.010868f
C4797 vdd.n2227 gnd 0.008748f
C4798 vdd.n2228 gnd 0.010868f
C4799 vdd.n2229 gnd 0.583113f
C4800 vdd.n2230 gnd 0.010868f
C4801 vdd.n2231 gnd 0.008748f
C4802 vdd.n2232 gnd 0.010868f
C4803 vdd.n2233 gnd 0.010868f
C4804 vdd.n2234 gnd 0.010868f
C4805 vdd.n2235 gnd 0.008748f
C4806 vdd.n2236 gnd 0.010868f
C4807 vdd.n2237 gnd 0.760824f
C4808 vdd.n2238 gnd 0.716396f
C4809 vdd.n2239 gnd 0.010868f
C4810 vdd.n2240 gnd 0.008748f
C4811 vdd.n2241 gnd 0.010868f
C4812 vdd.n2242 gnd 0.010868f
C4813 vdd.n2243 gnd 0.010868f
C4814 vdd.n2244 gnd 0.008748f
C4815 vdd.n2245 gnd 0.010868f
C4816 vdd.n2246 gnd 0.905214f
C4817 vdd.n2247 gnd 0.010868f
C4818 vdd.n2248 gnd 0.008748f
C4819 vdd.n2249 gnd 0.010868f
C4820 vdd.n2250 gnd 0.010868f
C4821 vdd.n2251 gnd 0.026291f
C4822 vdd.n2252 gnd 0.010868f
C4823 vdd.n2253 gnd 0.010868f
C4824 vdd.n2254 gnd 0.008748f
C4825 vdd.n2255 gnd 0.010868f
C4826 vdd.n2256 gnd 0.671969f
C4827 vdd.n2257 gnd 1.11069f
C4828 vdd.n2258 gnd 0.010868f
C4829 vdd.n2259 gnd 0.008748f
C4830 vdd.n2260 gnd 0.010868f
C4831 vdd.n2261 gnd 0.010868f
C4832 vdd.n2262 gnd 0.026291f
C4833 vdd.n2263 gnd 0.007261f
C4834 vdd.n2264 gnd 0.026291f
C4835 vdd.n2265 gnd 1.5272f
C4836 vdd.n2266 gnd 0.026291f
C4837 vdd.n2267 gnd 0.026855f
C4838 vdd.n2268 gnd 0.004155f
C4839 vdd.t69 gnd 0.133709f
C4840 vdd.t68 gnd 0.142898f
C4841 vdd.t66 gnd 0.174622f
C4842 vdd.n2269 gnd 0.223841f
C4843 vdd.n2270 gnd 0.188067f
C4844 vdd.n2271 gnd 0.013471f
C4845 vdd.n2272 gnd 0.004593f
C4846 vdd.n2273 gnd 0.009347f
C4847 vdd.n2274 gnd 0.821922f
C4848 vdd.n2276 gnd 0.008748f
C4849 vdd.n2277 gnd 0.008748f
C4850 vdd.n2278 gnd 0.010868f
C4851 vdd.n2280 gnd 0.010868f
C4852 vdd.n2281 gnd 0.010868f
C4853 vdd.n2282 gnd 0.008748f
C4854 vdd.n2283 gnd 0.008748f
C4855 vdd.n2284 gnd 0.008748f
C4856 vdd.n2285 gnd 0.010868f
C4857 vdd.n2287 gnd 0.010868f
C4858 vdd.n2288 gnd 0.010868f
C4859 vdd.n2289 gnd 0.008748f
C4860 vdd.n2290 gnd 0.008748f
C4861 vdd.n2291 gnd 0.008748f
C4862 vdd.n2292 gnd 0.010868f
C4863 vdd.n2294 gnd 0.010868f
C4864 vdd.n2295 gnd 0.010868f
C4865 vdd.n2296 gnd 0.008748f
C4866 vdd.n2297 gnd 0.008748f
C4867 vdd.n2298 gnd 0.008748f
C4868 vdd.n2299 gnd 0.010868f
C4869 vdd.n2301 gnd 0.010868f
C4870 vdd.n2302 gnd 0.010868f
C4871 vdd.n2303 gnd 0.008748f
C4872 vdd.n2304 gnd 0.010868f
C4873 vdd.n2305 gnd 0.010868f
C4874 vdd.n2306 gnd 0.010868f
C4875 vdd.n2307 gnd 0.017845f
C4876 vdd.n2308 gnd 0.005948f
C4877 vdd.n2309 gnd 0.008748f
C4878 vdd.n2310 gnd 0.010868f
C4879 vdd.n2312 gnd 0.010868f
C4880 vdd.n2313 gnd 0.010868f
C4881 vdd.n2314 gnd 0.008748f
C4882 vdd.n2315 gnd 0.008748f
C4883 vdd.n2316 gnd 0.008748f
C4884 vdd.n2317 gnd 0.010868f
C4885 vdd.n2319 gnd 0.010868f
C4886 vdd.n2320 gnd 0.010868f
C4887 vdd.n2321 gnd 0.008748f
C4888 vdd.n2322 gnd 0.008748f
C4889 vdd.n2323 gnd 0.008748f
C4890 vdd.n2324 gnd 0.010868f
C4891 vdd.n2326 gnd 0.010868f
C4892 vdd.n2327 gnd 0.010868f
C4893 vdd.n2328 gnd 0.008748f
C4894 vdd.n2329 gnd 0.008748f
C4895 vdd.n2330 gnd 0.008748f
C4896 vdd.n2331 gnd 0.010868f
C4897 vdd.n2333 gnd 0.010868f
C4898 vdd.n2334 gnd 0.010868f
C4899 vdd.n2335 gnd 0.008748f
C4900 vdd.n2336 gnd 0.008748f
C4901 vdd.n2337 gnd 0.008748f
C4902 vdd.n2338 gnd 0.010868f
C4903 vdd.n2340 gnd 0.010868f
C4904 vdd.n2341 gnd 0.010868f
C4905 vdd.n2342 gnd 0.008748f
C4906 vdd.n2343 gnd 0.010868f
C4907 vdd.n2344 gnd 0.010868f
C4908 vdd.n2345 gnd 0.010868f
C4909 vdd.n2346 gnd 0.017845f
C4910 vdd.n2347 gnd 0.007304f
C4911 vdd.n2348 gnd 0.008748f
C4912 vdd.n2349 gnd 0.010868f
C4913 vdd.n2351 gnd 0.010868f
C4914 vdd.n2352 gnd 0.010868f
C4915 vdd.n2353 gnd 0.008748f
C4916 vdd.n2354 gnd 0.008748f
C4917 vdd.n2355 gnd 0.008748f
C4918 vdd.n2356 gnd 0.010868f
C4919 vdd.n2358 gnd 0.010868f
C4920 vdd.n2359 gnd 0.010868f
C4921 vdd.n2360 gnd 0.008748f
C4922 vdd.n2361 gnd 0.008748f
C4923 vdd.n2362 gnd 0.008748f
C4924 vdd.n2363 gnd 0.010868f
C4925 vdd.n2365 gnd 0.010868f
C4926 vdd.n2366 gnd 0.010868f
C4927 vdd.n2367 gnd 0.008748f
C4928 vdd.n2368 gnd 0.008748f
C4929 vdd.n2369 gnd 0.008748f
C4930 vdd.n2370 gnd 0.010868f
C4931 vdd.n2372 gnd 0.010868f
C4932 vdd.n2373 gnd 0.008748f
C4933 vdd.n2374 gnd 0.008748f
C4934 vdd.n2375 gnd 0.010868f
C4935 vdd.n2377 gnd 0.010868f
C4936 vdd.n2378 gnd 0.010868f
C4937 vdd.n2379 gnd 0.008748f
C4938 vdd.n2380 gnd 0.009347f
C4939 vdd.n2381 gnd 0.821922f
C4940 vdd.n2382 gnd 0.029621f
C4941 vdd.n2383 gnd 0.00739f
C4942 vdd.n2384 gnd 0.00739f
C4943 vdd.n2385 gnd 0.00739f
C4944 vdd.n2386 gnd 0.00739f
C4945 vdd.n2387 gnd 0.00739f
C4946 vdd.n2388 gnd 0.00739f
C4947 vdd.n2389 gnd 0.00739f
C4948 vdd.n2390 gnd 0.00739f
C4949 vdd.n2391 gnd 0.00739f
C4950 vdd.n2392 gnd 0.00739f
C4951 vdd.n2393 gnd 0.00739f
C4952 vdd.n2394 gnd 0.00739f
C4953 vdd.n2395 gnd 0.00739f
C4954 vdd.n2396 gnd 0.00739f
C4955 vdd.n2397 gnd 0.00739f
C4956 vdd.n2398 gnd 0.00739f
C4957 vdd.n2399 gnd 0.00739f
C4958 vdd.n2400 gnd 0.00739f
C4959 vdd.n2401 gnd 0.00739f
C4960 vdd.n2402 gnd 0.00739f
C4961 vdd.n2403 gnd 0.00739f
C4962 vdd.n2404 gnd 0.00739f
C4963 vdd.n2405 gnd 0.00739f
C4964 vdd.n2406 gnd 0.00739f
C4965 vdd.n2407 gnd 0.00739f
C4966 vdd.n2408 gnd 0.00739f
C4967 vdd.n2409 gnd 0.00739f
C4968 vdd.n2410 gnd 0.00739f
C4969 vdd.n2411 gnd 0.00739f
C4970 vdd.n2412 gnd 0.00739f
C4971 vdd.n2413 gnd 0.00739f
C4972 vdd.n2414 gnd 0.017286f
C4973 vdd.n2415 gnd 0.017286f
C4974 vdd.n2417 gnd 9.4742f
C4975 vdd.n2419 gnd 0.017286f
C4976 vdd.n2420 gnd 0.017286f
C4977 vdd.n2421 gnd 0.016189f
C4978 vdd.n2422 gnd 0.00739f
C4979 vdd.n2423 gnd 0.00739f
C4980 vdd.n2424 gnd 0.755271f
C4981 vdd.n2425 gnd 0.00739f
C4982 vdd.n2426 gnd 0.00739f
C4983 vdd.n2427 gnd 0.00739f
C4984 vdd.n2428 gnd 0.00739f
C4985 vdd.n2429 gnd 0.00739f
C4986 vdd.n2430 gnd 0.638648f
C4987 vdd.n2431 gnd 0.00739f
C4988 vdd.n2432 gnd 0.00739f
C4989 vdd.n2433 gnd 0.00739f
C4990 vdd.n2434 gnd 0.00739f
C4991 vdd.n2435 gnd 0.00739f
C4992 vdd.n2436 gnd 0.755271f
C4993 vdd.n2437 gnd 0.00739f
C4994 vdd.n2438 gnd 0.00739f
C4995 vdd.n2439 gnd 0.00739f
C4996 vdd.n2440 gnd 0.00739f
C4997 vdd.n2441 gnd 0.00739f
C4998 vdd.n2442 gnd 0.73861f
C4999 vdd.n2443 gnd 0.00739f
C5000 vdd.n2444 gnd 0.00739f
C5001 vdd.n2445 gnd 0.00739f
C5002 vdd.n2446 gnd 0.00739f
C5003 vdd.n2447 gnd 0.00739f
C5004 vdd.n2448 gnd 0.755271f
C5005 vdd.n2449 gnd 0.00739f
C5006 vdd.n2450 gnd 0.00739f
C5007 vdd.n2451 gnd 0.00739f
C5008 vdd.n2452 gnd 0.00739f
C5009 vdd.n2453 gnd 0.00739f
C5010 vdd.n2454 gnd 0.605327f
C5011 vdd.n2455 gnd 0.00739f
C5012 vdd.n2456 gnd 0.00739f
C5013 vdd.n2457 gnd 0.006304f
C5014 vdd.n2458 gnd 0.021409f
C5015 vdd.n2459 gnd 0.004782f
C5016 vdd.n2460 gnd 0.00739f
C5017 vdd.n2461 gnd 0.438723f
C5018 vdd.n2462 gnd 0.00739f
C5019 vdd.n2463 gnd 0.00739f
C5020 vdd.n2464 gnd 0.00739f
C5021 vdd.n2465 gnd 0.00739f
C5022 vdd.n2466 gnd 0.00739f
C5023 vdd.n2467 gnd 0.483151f
C5024 vdd.n2468 gnd 0.00739f
C5025 vdd.n2469 gnd 0.00739f
C5026 vdd.n2470 gnd 0.00739f
C5027 vdd.n2471 gnd 0.00739f
C5028 vdd.n2472 gnd 0.00739f
C5029 vdd.n2473 gnd 0.649755f
C5030 vdd.n2474 gnd 0.00739f
C5031 vdd.n2475 gnd 0.00739f
C5032 vdd.n2476 gnd 0.00739f
C5033 vdd.n2477 gnd 0.00739f
C5034 vdd.n2478 gnd 0.00739f
C5035 vdd.n2479 gnd 0.621988f
C5036 vdd.n2480 gnd 0.00739f
C5037 vdd.n2481 gnd 0.00739f
C5038 vdd.n2482 gnd 0.00739f
C5039 vdd.n2483 gnd 0.00739f
C5040 vdd.n2484 gnd 0.00739f
C5041 vdd.n2485 gnd 0.455384f
C5042 vdd.n2486 gnd 0.00739f
C5043 vdd.n2487 gnd 0.00739f
C5044 vdd.n2488 gnd 0.00739f
C5045 vdd.n2489 gnd 0.00739f
C5046 vdd.n2490 gnd 0.00739f
C5047 vdd.n2491 gnd 0.238799f
C5048 vdd.n2492 gnd 0.00739f
C5049 vdd.n2493 gnd 0.00739f
C5050 vdd.n2494 gnd 0.00739f
C5051 vdd.n2495 gnd 0.00739f
C5052 vdd.n2496 gnd 0.00739f
C5053 vdd.n2497 gnd 0.394296f
C5054 vdd.n2498 gnd 0.00739f
C5055 vdd.n2499 gnd 0.00739f
C5056 vdd.n2500 gnd 0.00739f
C5057 vdd.n2501 gnd 0.00739f
C5058 vdd.n2502 gnd 0.00739f
C5059 vdd.n2503 gnd 0.755271f
C5060 vdd.n2504 gnd 0.00739f
C5061 vdd.n2505 gnd 0.00739f
C5062 vdd.n2506 gnd 0.00739f
C5063 vdd.n2507 gnd 0.00739f
C5064 vdd.n2508 gnd 0.00739f
C5065 vdd.n2509 gnd 0.00739f
C5066 vdd.n2510 gnd 0.00739f
C5067 vdd.n2511 gnd 0.566453f
C5068 vdd.n2512 gnd 0.00739f
C5069 vdd.n2513 gnd 0.00739f
C5070 vdd.n2514 gnd 0.00739f
C5071 vdd.n2515 gnd 0.00739f
C5072 vdd.n2516 gnd 0.00739f
C5073 vdd.n2517 gnd 0.00739f
C5074 vdd.n2518 gnd 0.472044f
C5075 vdd.n2519 gnd 0.00739f
C5076 vdd.n2520 gnd 0.00739f
C5077 vdd.n2521 gnd 0.00739f
C5078 vdd.n2522 gnd 0.017107f
C5079 vdd.n2523 gnd 0.016368f
C5080 vdd.n2524 gnd 0.00739f
C5081 vdd.n2525 gnd 0.00739f
C5082 vdd.n2526 gnd 0.005706f
C5083 vdd.n2527 gnd 0.00739f
C5084 vdd.n2528 gnd 0.00739f
C5085 vdd.n2529 gnd 0.00538f
C5086 vdd.n2530 gnd 0.00739f
C5087 vdd.n2531 gnd 0.00739f
C5088 vdd.n2532 gnd 0.00739f
C5089 vdd.n2533 gnd 0.00739f
C5090 vdd.n2534 gnd 0.00739f
C5091 vdd.n2535 gnd 0.00739f
C5092 vdd.n2536 gnd 0.00739f
C5093 vdd.n2537 gnd 0.00739f
C5094 vdd.n2538 gnd 0.00739f
C5095 vdd.n2539 gnd 0.00739f
C5096 vdd.n2540 gnd 0.00739f
C5097 vdd.n2541 gnd 0.00739f
C5098 vdd.n2542 gnd 0.00739f
C5099 vdd.n2543 gnd 0.00739f
C5100 vdd.n2544 gnd 0.00739f
C5101 vdd.n2545 gnd 0.00739f
C5102 vdd.n2546 gnd 0.00739f
C5103 vdd.n2547 gnd 0.00739f
C5104 vdd.n2548 gnd 0.00739f
C5105 vdd.n2549 gnd 0.00739f
C5106 vdd.n2550 gnd 0.00739f
C5107 vdd.n2551 gnd 0.00739f
C5108 vdd.n2552 gnd 0.00739f
C5109 vdd.n2553 gnd 0.00739f
C5110 vdd.n2554 gnd 0.00739f
C5111 vdd.n2555 gnd 0.00739f
C5112 vdd.n2556 gnd 0.00739f
C5113 vdd.n2557 gnd 0.00739f
C5114 vdd.n2558 gnd 0.00739f
C5115 vdd.n2559 gnd 0.00739f
C5116 vdd.n2560 gnd 0.00739f
C5117 vdd.n2561 gnd 0.00739f
C5118 vdd.n2562 gnd 0.00739f
C5119 vdd.n2563 gnd 0.00739f
C5120 vdd.n2564 gnd 0.00739f
C5121 vdd.n2565 gnd 0.00739f
C5122 vdd.n2566 gnd 0.00739f
C5123 vdd.n2567 gnd 0.00739f
C5124 vdd.n2568 gnd 0.00739f
C5125 vdd.n2569 gnd 0.00739f
C5126 vdd.n2570 gnd 0.00739f
C5127 vdd.n2571 gnd 0.00739f
C5128 vdd.n2572 gnd 0.00739f
C5129 vdd.n2573 gnd 0.00739f
C5130 vdd.n2574 gnd 0.00739f
C5131 vdd.n2575 gnd 0.00739f
C5132 vdd.n2576 gnd 0.00739f
C5133 vdd.n2577 gnd 0.00739f
C5134 vdd.n2578 gnd 0.00739f
C5135 vdd.n2579 gnd 0.00739f
C5136 vdd.n2580 gnd 0.00739f
C5137 vdd.n2581 gnd 0.00739f
C5138 vdd.n2582 gnd 0.00739f
C5139 vdd.n2583 gnd 0.00739f
C5140 vdd.n2584 gnd 0.00739f
C5141 vdd.n2585 gnd 0.00739f
C5142 vdd.n2586 gnd 0.00739f
C5143 vdd.n2587 gnd 0.00739f
C5144 vdd.n2588 gnd 0.00739f
C5145 vdd.n2589 gnd 0.00739f
C5146 vdd.n2590 gnd 0.017286f
C5147 vdd.n2591 gnd 0.016189f
C5148 vdd.n2592 gnd 0.016189f
C5149 vdd.n2593 gnd 0.899661f
C5150 vdd.n2594 gnd 0.016189f
C5151 vdd.n2595 gnd 0.017286f
C5152 vdd.n2596 gnd 0.016368f
C5153 vdd.n2597 gnd 0.00739f
C5154 vdd.n2598 gnd 0.00739f
C5155 vdd.n2599 gnd 0.00739f
C5156 vdd.n2600 gnd 0.005706f
C5157 vdd.n2601 gnd 0.010562f
C5158 vdd.n2602 gnd 0.00538f
C5159 vdd.n2603 gnd 0.00739f
C5160 vdd.n2604 gnd 0.00739f
C5161 vdd.n2605 gnd 0.00739f
C5162 vdd.n2606 gnd 0.00739f
C5163 vdd.n2607 gnd 0.00739f
C5164 vdd.n2608 gnd 0.00739f
C5165 vdd.n2609 gnd 0.00739f
C5166 vdd.n2610 gnd 0.00739f
C5167 vdd.n2611 gnd 0.00739f
C5168 vdd.n2612 gnd 0.00739f
C5169 vdd.n2613 gnd 0.00739f
C5170 vdd.n2614 gnd 0.00739f
C5171 vdd.n2615 gnd 0.00739f
C5172 vdd.n2616 gnd 0.00739f
C5173 vdd.n2617 gnd 0.00739f
C5174 vdd.n2618 gnd 0.00739f
C5175 vdd.n2619 gnd 0.00739f
C5176 vdd.n2620 gnd 0.00739f
C5177 vdd.n2621 gnd 0.00739f
C5178 vdd.n2622 gnd 0.00739f
C5179 vdd.n2623 gnd 0.00739f
C5180 vdd.n2624 gnd 0.00739f
C5181 vdd.n2625 gnd 0.00739f
C5182 vdd.n2626 gnd 0.00739f
C5183 vdd.n2627 gnd 0.00739f
C5184 vdd.n2628 gnd 0.00739f
C5185 vdd.n2629 gnd 0.00739f
C5186 vdd.n2630 gnd 0.00739f
C5187 vdd.n2631 gnd 0.00739f
C5188 vdd.n2632 gnd 0.00739f
C5189 vdd.n2633 gnd 0.00739f
C5190 vdd.n2634 gnd 0.00739f
C5191 vdd.n2635 gnd 0.00739f
C5192 vdd.n2636 gnd 0.00739f
C5193 vdd.n2637 gnd 0.00739f
C5194 vdd.n2638 gnd 0.00739f
C5195 vdd.n2639 gnd 0.00739f
C5196 vdd.n2640 gnd 0.00739f
C5197 vdd.n2641 gnd 0.00739f
C5198 vdd.n2642 gnd 0.00739f
C5199 vdd.n2643 gnd 0.00739f
C5200 vdd.n2644 gnd 0.00739f
C5201 vdd.n2645 gnd 0.00739f
C5202 vdd.n2646 gnd 0.00739f
C5203 vdd.n2647 gnd 0.00739f
C5204 vdd.n2648 gnd 0.00739f
C5205 vdd.n2649 gnd 0.00739f
C5206 vdd.n2650 gnd 0.00739f
C5207 vdd.n2651 gnd 0.00739f
C5208 vdd.n2652 gnd 0.00739f
C5209 vdd.n2653 gnd 0.00739f
C5210 vdd.n2654 gnd 0.00739f
C5211 vdd.n2655 gnd 0.00739f
C5212 vdd.n2656 gnd 0.00739f
C5213 vdd.n2657 gnd 0.00739f
C5214 vdd.n2658 gnd 0.00739f
C5215 vdd.n2659 gnd 0.00739f
C5216 vdd.n2660 gnd 0.00739f
C5217 vdd.n2661 gnd 0.00739f
C5218 vdd.n2662 gnd 0.00739f
C5219 vdd.n2663 gnd 0.017286f
C5220 vdd.n2664 gnd 0.017286f
C5221 vdd.n2665 gnd 0.921874f
C5222 vdd.t130 gnd 3.27654f
C5223 vdd.t22 gnd 3.27654f
C5224 vdd.n2698 gnd 0.017286f
C5225 vdd.t51 gnd 0.688629f
C5226 vdd.n2699 gnd 0.00739f
C5227 vdd.n2700 gnd 0.00739f
C5228 vdd.t106 gnd 0.298648f
C5229 vdd.t107 gnd 0.305703f
C5230 vdd.t104 gnd 0.194969f
C5231 vdd.n2701 gnd 0.10537f
C5232 vdd.n2702 gnd 0.059769f
C5233 vdd.n2703 gnd 0.00739f
C5234 vdd.t116 gnd 0.298648f
C5235 vdd.t117 gnd 0.305703f
C5236 vdd.t115 gnd 0.194969f
C5237 vdd.n2704 gnd 0.10537f
C5238 vdd.n2705 gnd 0.059769f
C5239 vdd.n2706 gnd 0.010562f
C5240 vdd.n2707 gnd 0.00739f
C5241 vdd.n2708 gnd 0.00739f
C5242 vdd.n2709 gnd 0.00739f
C5243 vdd.n2710 gnd 0.00739f
C5244 vdd.n2711 gnd 0.00739f
C5245 vdd.n2712 gnd 0.00739f
C5246 vdd.n2713 gnd 0.00739f
C5247 vdd.n2714 gnd 0.00739f
C5248 vdd.n2715 gnd 0.00739f
C5249 vdd.n2716 gnd 0.00739f
C5250 vdd.n2717 gnd 0.00739f
C5251 vdd.n2718 gnd 0.00739f
C5252 vdd.n2719 gnd 0.00739f
C5253 vdd.n2720 gnd 0.00739f
C5254 vdd.n2721 gnd 0.00739f
C5255 vdd.n2722 gnd 0.00739f
C5256 vdd.n2723 gnd 0.00739f
C5257 vdd.n2724 gnd 0.00739f
C5258 vdd.n2725 gnd 0.00739f
C5259 vdd.n2726 gnd 0.00739f
C5260 vdd.n2727 gnd 0.00739f
C5261 vdd.n2728 gnd 0.00739f
C5262 vdd.n2729 gnd 0.00739f
C5263 vdd.n2730 gnd 0.00739f
C5264 vdd.n2731 gnd 0.00739f
C5265 vdd.n2732 gnd 0.00739f
C5266 vdd.n2733 gnd 0.00739f
C5267 vdd.n2734 gnd 0.00739f
C5268 vdd.n2735 gnd 0.00739f
C5269 vdd.n2736 gnd 0.00739f
C5270 vdd.n2737 gnd 0.00739f
C5271 vdd.n2738 gnd 0.00739f
C5272 vdd.n2739 gnd 0.00739f
C5273 vdd.n2740 gnd 0.00739f
C5274 vdd.n2741 gnd 0.00739f
C5275 vdd.n2742 gnd 0.00739f
C5276 vdd.n2743 gnd 0.00739f
C5277 vdd.n2744 gnd 0.00739f
C5278 vdd.n2745 gnd 0.00739f
C5279 vdd.n2746 gnd 0.00739f
C5280 vdd.n2747 gnd 0.00739f
C5281 vdd.n2748 gnd 0.00739f
C5282 vdd.n2749 gnd 0.00739f
C5283 vdd.n2750 gnd 0.00739f
C5284 vdd.n2751 gnd 0.00739f
C5285 vdd.n2752 gnd 0.00739f
C5286 vdd.n2753 gnd 0.00739f
C5287 vdd.n2754 gnd 0.00739f
C5288 vdd.n2755 gnd 0.00739f
C5289 vdd.n2756 gnd 0.00739f
C5290 vdd.n2757 gnd 0.00739f
C5291 vdd.n2758 gnd 0.00739f
C5292 vdd.n2759 gnd 0.00739f
C5293 vdd.n2760 gnd 0.00739f
C5294 vdd.n2761 gnd 0.00739f
C5295 vdd.n2762 gnd 0.00739f
C5296 vdd.n2763 gnd 0.00739f
C5297 vdd.n2764 gnd 0.00739f
C5298 vdd.n2765 gnd 0.00538f
C5299 vdd.n2766 gnd 0.00739f
C5300 vdd.n2767 gnd 0.00739f
C5301 vdd.n2768 gnd 0.005706f
C5302 vdd.n2769 gnd 0.00739f
C5303 vdd.n2770 gnd 0.00739f
C5304 vdd.n2771 gnd 0.017286f
C5305 vdd.n2772 gnd 0.016189f
C5306 vdd.n2773 gnd 0.016189f
C5307 vdd.n2774 gnd 0.00739f
C5308 vdd.n2775 gnd 0.00739f
C5309 vdd.n2776 gnd 0.00739f
C5310 vdd.n2777 gnd 0.00739f
C5311 vdd.n2778 gnd 0.00739f
C5312 vdd.n2779 gnd 0.00739f
C5313 vdd.n2780 gnd 0.00739f
C5314 vdd.n2781 gnd 0.00739f
C5315 vdd.n2782 gnd 0.00739f
C5316 vdd.n2783 gnd 0.00739f
C5317 vdd.n2784 gnd 0.00739f
C5318 vdd.n2785 gnd 0.00739f
C5319 vdd.n2786 gnd 0.00739f
C5320 vdd.n2787 gnd 0.00739f
C5321 vdd.n2788 gnd 0.00739f
C5322 vdd.n2789 gnd 0.00739f
C5323 vdd.n2790 gnd 0.00739f
C5324 vdd.n2791 gnd 0.00739f
C5325 vdd.n2792 gnd 0.00739f
C5326 vdd.n2793 gnd 0.00739f
C5327 vdd.n2794 gnd 0.00739f
C5328 vdd.n2795 gnd 0.00739f
C5329 vdd.n2796 gnd 0.00739f
C5330 vdd.n2797 gnd 0.00739f
C5331 vdd.n2798 gnd 0.00739f
C5332 vdd.n2799 gnd 0.00739f
C5333 vdd.n2800 gnd 0.00739f
C5334 vdd.n2801 gnd 0.00739f
C5335 vdd.n2802 gnd 0.00739f
C5336 vdd.n2803 gnd 0.00739f
C5337 vdd.n2804 gnd 0.00739f
C5338 vdd.n2805 gnd 0.00739f
C5339 vdd.n2806 gnd 0.00739f
C5340 vdd.n2807 gnd 0.00739f
C5341 vdd.n2808 gnd 0.00739f
C5342 vdd.n2809 gnd 0.00739f
C5343 vdd.n2810 gnd 0.00739f
C5344 vdd.n2811 gnd 0.00739f
C5345 vdd.n2812 gnd 0.00739f
C5346 vdd.n2813 gnd 0.00739f
C5347 vdd.n2814 gnd 0.00739f
C5348 vdd.n2815 gnd 0.00739f
C5349 vdd.n2816 gnd 0.00739f
C5350 vdd.n2817 gnd 0.00739f
C5351 vdd.n2818 gnd 0.00739f
C5352 vdd.n2819 gnd 0.00739f
C5353 vdd.n2820 gnd 0.00739f
C5354 vdd.n2821 gnd 0.00739f
C5355 vdd.n2822 gnd 0.00739f
C5356 vdd.n2823 gnd 0.00739f
C5357 vdd.n2824 gnd 0.00739f
C5358 vdd.n2825 gnd 0.00739f
C5359 vdd.n2826 gnd 0.00739f
C5360 vdd.n2827 gnd 0.00739f
C5361 vdd.n2828 gnd 0.00739f
C5362 vdd.n2829 gnd 0.00739f
C5363 vdd.n2830 gnd 0.00739f
C5364 vdd.n2831 gnd 0.00739f
C5365 vdd.n2832 gnd 0.00739f
C5366 vdd.n2833 gnd 0.00739f
C5367 vdd.n2834 gnd 0.00739f
C5368 vdd.n2835 gnd 0.00739f
C5369 vdd.n2836 gnd 0.00739f
C5370 vdd.n2837 gnd 0.00739f
C5371 vdd.n2838 gnd 0.00739f
C5372 vdd.n2839 gnd 0.00739f
C5373 vdd.n2840 gnd 0.00739f
C5374 vdd.n2841 gnd 0.00739f
C5375 vdd.n2842 gnd 0.00739f
C5376 vdd.n2843 gnd 0.00739f
C5377 vdd.n2844 gnd 0.00739f
C5378 vdd.n2845 gnd 0.00739f
C5379 vdd.n2846 gnd 0.00739f
C5380 vdd.n2847 gnd 0.238799f
C5381 vdd.n2848 gnd 0.00739f
C5382 vdd.n2849 gnd 0.00739f
C5383 vdd.n2850 gnd 0.00739f
C5384 vdd.n2851 gnd 0.00739f
C5385 vdd.n2852 gnd 0.00739f
C5386 vdd.n2853 gnd 0.00739f
C5387 vdd.n2854 gnd 0.00739f
C5388 vdd.n2855 gnd 0.00739f
C5389 vdd.n2856 gnd 0.00739f
C5390 vdd.n2857 gnd 0.00739f
C5391 vdd.n2858 gnd 0.00739f
C5392 vdd.n2859 gnd 0.00739f
C5393 vdd.n2860 gnd 0.00739f
C5394 vdd.n2861 gnd 0.00739f
C5395 vdd.n2862 gnd 0.472044f
C5396 vdd.n2863 gnd 0.00739f
C5397 vdd.n2864 gnd 0.00739f
C5398 vdd.n2865 gnd 0.00739f
C5399 vdd.n2866 gnd 0.016189f
C5400 vdd.n2867 gnd 0.016189f
C5401 vdd.n2868 gnd 0.017286f
C5402 vdd.n2869 gnd 0.017286f
C5403 vdd.n2870 gnd 0.00739f
C5404 vdd.n2871 gnd 0.00739f
C5405 vdd.n2872 gnd 0.00739f
C5406 vdd.n2873 gnd 0.005706f
C5407 vdd.n2874 gnd 0.010562f
C5408 vdd.n2875 gnd 0.00538f
C5409 vdd.n2876 gnd 0.00739f
C5410 vdd.n2877 gnd 0.00739f
C5411 vdd.n2878 gnd 0.00739f
C5412 vdd.n2879 gnd 0.00739f
C5413 vdd.n2880 gnd 0.00739f
C5414 vdd.n2881 gnd 0.00739f
C5415 vdd.n2882 gnd 0.00739f
C5416 vdd.n2883 gnd 0.00739f
C5417 vdd.n2884 gnd 0.00739f
C5418 vdd.n2885 gnd 0.00739f
C5419 vdd.n2886 gnd 0.00739f
C5420 vdd.n2887 gnd 0.00739f
C5421 vdd.n2888 gnd 0.00739f
C5422 vdd.n2889 gnd 0.00739f
C5423 vdd.n2890 gnd 0.00739f
C5424 vdd.n2891 gnd 0.00739f
C5425 vdd.n2892 gnd 0.00739f
C5426 vdd.n2893 gnd 0.00739f
C5427 vdd.n2894 gnd 0.00739f
C5428 vdd.n2895 gnd 0.00739f
C5429 vdd.n2896 gnd 0.00739f
C5430 vdd.n2897 gnd 0.00739f
C5431 vdd.n2898 gnd 0.00739f
C5432 vdd.n2899 gnd 0.00739f
C5433 vdd.n2900 gnd 0.00739f
C5434 vdd.n2901 gnd 0.00739f
C5435 vdd.n2902 gnd 0.00739f
C5436 vdd.n2903 gnd 0.00739f
C5437 vdd.n2904 gnd 0.00739f
C5438 vdd.n2905 gnd 0.00739f
C5439 vdd.n2906 gnd 0.00739f
C5440 vdd.n2907 gnd 0.00739f
C5441 vdd.n2908 gnd 0.00739f
C5442 vdd.n2909 gnd 0.00739f
C5443 vdd.n2910 gnd 0.00739f
C5444 vdd.n2911 gnd 0.00739f
C5445 vdd.n2912 gnd 0.00739f
C5446 vdd.n2913 gnd 0.00739f
C5447 vdd.n2914 gnd 0.00739f
C5448 vdd.n2915 gnd 0.00739f
C5449 vdd.n2916 gnd 0.00739f
C5450 vdd.n2917 gnd 0.00739f
C5451 vdd.n2918 gnd 0.00739f
C5452 vdd.n2919 gnd 0.00739f
C5453 vdd.n2920 gnd 0.00739f
C5454 vdd.n2921 gnd 0.00739f
C5455 vdd.n2922 gnd 0.00739f
C5456 vdd.n2923 gnd 0.00739f
C5457 vdd.n2924 gnd 0.00739f
C5458 vdd.n2925 gnd 0.00739f
C5459 vdd.n2926 gnd 0.00739f
C5460 vdd.n2927 gnd 0.00739f
C5461 vdd.n2928 gnd 0.00739f
C5462 vdd.n2929 gnd 0.00739f
C5463 vdd.n2930 gnd 0.00739f
C5464 vdd.n2931 gnd 0.00739f
C5465 vdd.n2932 gnd 0.00739f
C5466 vdd.n2933 gnd 0.00739f
C5467 vdd.n2934 gnd 0.00739f
C5468 vdd.n2935 gnd 0.017286f
C5469 vdd.n2936 gnd 0.017286f
C5470 vdd.n2938 gnd 0.921874f
C5471 vdd.n2940 gnd 0.017286f
C5472 vdd.n2941 gnd 0.017286f
C5473 vdd.n2942 gnd 0.016189f
C5474 vdd.n2943 gnd 0.00739f
C5475 vdd.n2944 gnd 0.00739f
C5476 vdd.n2945 gnd 0.399849f
C5477 vdd.n2946 gnd 0.00739f
C5478 vdd.n2947 gnd 0.00739f
C5479 vdd.n2948 gnd 0.00739f
C5480 vdd.n2949 gnd 0.00739f
C5481 vdd.n2950 gnd 0.00739f
C5482 vdd.n2951 gnd 0.44983f
C5483 vdd.n2952 gnd 0.00739f
C5484 vdd.n2953 gnd 0.00739f
C5485 vdd.n2954 gnd 0.00739f
C5486 vdd.n2955 gnd 0.00739f
C5487 vdd.n2956 gnd 0.00739f
C5488 vdd.n2957 gnd 0.755271f
C5489 vdd.n2958 gnd 0.00739f
C5490 vdd.n2959 gnd 0.00739f
C5491 vdd.n2960 gnd 0.00739f
C5492 vdd.n2961 gnd 0.00739f
C5493 vdd.n2962 gnd 0.00739f
C5494 vdd.n2963 gnd 0.499811f
C5495 vdd.n2964 gnd 0.00739f
C5496 vdd.n2965 gnd 0.00739f
C5497 vdd.n2966 gnd 0.00739f
C5498 vdd.n2967 gnd 0.00739f
C5499 vdd.n2968 gnd 0.00739f
C5500 vdd.n2969 gnd 0.666415f
C5501 vdd.n2970 gnd 0.00739f
C5502 vdd.n2971 gnd 0.00739f
C5503 vdd.n2972 gnd 0.00739f
C5504 vdd.n2973 gnd 0.00739f
C5505 vdd.n2974 gnd 0.00739f
C5506 vdd.n2975 gnd 0.605327f
C5507 vdd.n2976 gnd 0.00739f
C5508 vdd.n2977 gnd 0.00739f
C5509 vdd.n2978 gnd 0.00739f
C5510 vdd.n2979 gnd 0.00739f
C5511 vdd.n2980 gnd 0.00739f
C5512 vdd.n2981 gnd 0.438723f
C5513 vdd.n2982 gnd 0.00739f
C5514 vdd.n2983 gnd 0.00739f
C5515 vdd.n2984 gnd 0.00739f
C5516 vdd.n2985 gnd 0.00739f
C5517 vdd.n2986 gnd 0.00739f
C5518 vdd.n2987 gnd 0.238799f
C5519 vdd.n2988 gnd 0.00739f
C5520 vdd.n2989 gnd 0.00739f
C5521 vdd.n2990 gnd 0.00739f
C5522 vdd.n2991 gnd 0.00739f
C5523 vdd.n2992 gnd 0.00739f
C5524 vdd.n2993 gnd 0.649755f
C5525 vdd.n2994 gnd 0.00739f
C5526 vdd.n2995 gnd 0.00739f
C5527 vdd.n2996 gnd 0.00739f
C5528 vdd.n2997 gnd 0.00739f
C5529 vdd.n2998 gnd 0.00739f
C5530 vdd.n2999 gnd 0.755271f
C5531 vdd.n3000 gnd 0.00739f
C5532 vdd.n3001 gnd 0.00739f
C5533 vdd.n3002 gnd 0.004782f
C5534 vdd.n3003 gnd 0.021409f
C5535 vdd.n3004 gnd 0.006304f
C5536 vdd.n3005 gnd 0.00739f
C5537 vdd.n3006 gnd 0.644201f
C5538 vdd.n3007 gnd 0.00739f
C5539 vdd.n3008 gnd 0.00739f
C5540 vdd.n3009 gnd 0.00739f
C5541 vdd.n3010 gnd 0.00739f
C5542 vdd.n3011 gnd 0.00739f
C5543 vdd.n3012 gnd 0.527579f
C5544 vdd.n3013 gnd 0.00739f
C5545 vdd.n3014 gnd 0.00739f
C5546 vdd.n3015 gnd 0.00739f
C5547 vdd.n3016 gnd 0.00739f
C5548 vdd.n3017 gnd 0.00739f
C5549 vdd.n3018 gnd 0.394296f
C5550 vdd.n3019 gnd 0.00739f
C5551 vdd.n3020 gnd 0.00739f
C5552 vdd.n3021 gnd 0.00739f
C5553 vdd.n3022 gnd 0.00739f
C5554 vdd.n3023 gnd 0.00739f
C5555 vdd.n3024 gnd 0.755271f
C5556 vdd.n3025 gnd 0.00739f
C5557 vdd.n3026 gnd 0.00739f
C5558 vdd.n3027 gnd 0.00739f
C5559 vdd.n3028 gnd 0.00739f
C5560 vdd.n3029 gnd 0.00739f
C5561 vdd.n3030 gnd 0.00739f
C5562 vdd.n3032 gnd 0.00739f
C5563 vdd.n3033 gnd 0.00739f
C5564 vdd.n3035 gnd 0.00739f
C5565 vdd.n3036 gnd 0.00739f
C5566 vdd.n3039 gnd 0.00739f
C5567 vdd.n3040 gnd 0.00739f
C5568 vdd.n3041 gnd 0.00739f
C5569 vdd.n3042 gnd 0.00739f
C5570 vdd.n3044 gnd 0.00739f
C5571 vdd.n3045 gnd 0.00739f
C5572 vdd.n3046 gnd 0.00739f
C5573 vdd.n3047 gnd 0.00739f
C5574 vdd.n3048 gnd 0.00739f
C5575 vdd.n3049 gnd 0.00739f
C5576 vdd.n3051 gnd 0.00739f
C5577 vdd.n3052 gnd 0.00739f
C5578 vdd.n3053 gnd 0.00739f
C5579 vdd.n3054 gnd 0.00739f
C5580 vdd.n3055 gnd 0.00739f
C5581 vdd.n3056 gnd 0.00739f
C5582 vdd.n3058 gnd 0.00739f
C5583 vdd.n3059 gnd 0.00739f
C5584 vdd.n3060 gnd 0.00739f
C5585 vdd.n3061 gnd 0.00739f
C5586 vdd.n3062 gnd 0.00739f
C5587 vdd.n3063 gnd 0.00739f
C5588 vdd.n3065 gnd 0.00739f
C5589 vdd.n3066 gnd 0.017286f
C5590 vdd.n3067 gnd 0.017286f
C5591 vdd.n3068 gnd 0.016189f
C5592 vdd.n3069 gnd 0.00739f
C5593 vdd.n3070 gnd 0.00739f
C5594 vdd.n3071 gnd 0.00739f
C5595 vdd.n3072 gnd 0.00739f
C5596 vdd.n3073 gnd 0.00739f
C5597 vdd.n3074 gnd 0.00739f
C5598 vdd.n3075 gnd 0.755271f
C5599 vdd.n3076 gnd 0.00739f
C5600 vdd.n3077 gnd 0.00739f
C5601 vdd.n3078 gnd 0.00739f
C5602 vdd.n3079 gnd 0.00739f
C5603 vdd.n3080 gnd 0.00739f
C5604 vdd.n3081 gnd 0.494258f
C5605 vdd.n3082 gnd 0.00739f
C5606 vdd.n3083 gnd 0.00739f
C5607 vdd.n3084 gnd 0.00739f
C5608 vdd.n3085 gnd 0.017107f
C5609 vdd.n3086 gnd 0.016368f
C5610 vdd.n3087 gnd 0.017286f
C5611 vdd.n3089 gnd 0.00739f
C5612 vdd.n3090 gnd 0.00739f
C5613 vdd.n3091 gnd 0.005706f
C5614 vdd.n3092 gnd 0.010562f
C5615 vdd.n3093 gnd 0.00538f
C5616 vdd.n3094 gnd 0.00739f
C5617 vdd.n3095 gnd 0.00739f
C5618 vdd.n3097 gnd 0.00739f
C5619 vdd.n3098 gnd 0.00739f
C5620 vdd.n3099 gnd 0.00739f
C5621 vdd.n3100 gnd 0.00739f
C5622 vdd.n3101 gnd 0.00739f
C5623 vdd.n3102 gnd 0.00739f
C5624 vdd.n3104 gnd 0.00739f
C5625 vdd.n3105 gnd 0.00739f
C5626 vdd.n3106 gnd 0.00739f
C5627 vdd.n3107 gnd 0.00739f
C5628 vdd.n3108 gnd 0.00739f
C5629 vdd.n3109 gnd 0.00739f
C5630 vdd.n3111 gnd 0.00739f
C5631 vdd.n3112 gnd 0.00739f
C5632 vdd.n3113 gnd 0.00739f
C5633 vdd.n3114 gnd 0.00739f
C5634 vdd.n3115 gnd 0.00739f
C5635 vdd.n3116 gnd 0.00739f
C5636 vdd.n3118 gnd 0.00739f
C5637 vdd.n3119 gnd 0.00739f
C5638 vdd.n3120 gnd 0.00739f
C5639 vdd.n3122 gnd 0.00739f
C5640 vdd.n3123 gnd 0.00739f
C5641 vdd.n3124 gnd 0.00739f
C5642 vdd.n3125 gnd 0.00739f
C5643 vdd.n3126 gnd 0.00739f
C5644 vdd.n3127 gnd 0.00739f
C5645 vdd.n3129 gnd 0.00739f
C5646 vdd.n3130 gnd 0.00739f
C5647 vdd.n3131 gnd 0.00739f
C5648 vdd.n3132 gnd 0.00739f
C5649 vdd.n3133 gnd 0.00739f
C5650 vdd.n3134 gnd 0.00739f
C5651 vdd.n3136 gnd 0.00739f
C5652 vdd.n3137 gnd 0.00739f
C5653 vdd.n3138 gnd 0.00739f
C5654 vdd.n3139 gnd 0.00739f
C5655 vdd.n3140 gnd 0.00739f
C5656 vdd.n3141 gnd 0.00739f
C5657 vdd.n3143 gnd 0.00739f
C5658 vdd.n3144 gnd 0.00739f
C5659 vdd.n3146 gnd 0.00739f
C5660 vdd.n3147 gnd 0.00739f
C5661 vdd.n3148 gnd 0.017286f
C5662 vdd.n3149 gnd 0.016189f
C5663 vdd.n3150 gnd 0.016189f
C5664 vdd.n3151 gnd 1.06626f
C5665 vdd.n3152 gnd 0.016189f
C5666 vdd.n3153 gnd 0.017286f
C5667 vdd.n3154 gnd 0.016368f
C5668 vdd.n3155 gnd 0.00739f
C5669 vdd.n3156 gnd 0.005706f
C5670 vdd.n3157 gnd 0.00739f
C5671 vdd.n3159 gnd 0.00739f
C5672 vdd.n3160 gnd 0.00739f
C5673 vdd.n3161 gnd 0.00739f
C5674 vdd.n3162 gnd 0.00739f
C5675 vdd.n3163 gnd 0.00739f
C5676 vdd.n3164 gnd 0.00739f
C5677 vdd.n3166 gnd 0.00739f
C5678 vdd.n3167 gnd 0.00739f
C5679 vdd.n3168 gnd 0.00739f
C5680 vdd.n3169 gnd 0.00739f
C5681 vdd.n3170 gnd 0.00739f
C5682 vdd.n3171 gnd 0.00739f
C5683 vdd.n3173 gnd 0.00739f
C5684 vdd.n3174 gnd 0.00739f
C5685 vdd.n3175 gnd 0.00739f
C5686 vdd.n3176 gnd 0.00739f
C5687 vdd.n3177 gnd 0.00739f
C5688 vdd.n3178 gnd 0.00739f
C5689 vdd.n3180 gnd 0.00739f
C5690 vdd.n3181 gnd 0.00739f
C5691 vdd.n3183 gnd 0.00739f
C5692 vdd.n3184 gnd 0.025382f
C5693 vdd.n3185 gnd 0.826161f
C5694 vdd.n3187 gnd 0.004593f
C5695 vdd.n3188 gnd 0.008748f
C5696 vdd.n3189 gnd 0.010868f
C5697 vdd.n3190 gnd 0.010868f
C5698 vdd.n3191 gnd 0.008748f
C5699 vdd.n3192 gnd 0.008748f
C5700 vdd.n3193 gnd 0.010868f
C5701 vdd.n3194 gnd 0.010868f
C5702 vdd.n3195 gnd 0.008748f
C5703 vdd.n3196 gnd 0.008748f
C5704 vdd.n3197 gnd 0.010868f
C5705 vdd.n3198 gnd 0.010868f
C5706 vdd.n3199 gnd 0.008748f
C5707 vdd.n3200 gnd 0.008748f
C5708 vdd.n3201 gnd 0.010868f
C5709 vdd.n3202 gnd 0.010868f
C5710 vdd.n3203 gnd 0.008748f
C5711 vdd.n3204 gnd 0.008748f
C5712 vdd.n3205 gnd 0.010868f
C5713 vdd.n3206 gnd 0.010868f
C5714 vdd.n3207 gnd 0.008748f
C5715 vdd.n3208 gnd 0.008748f
C5716 vdd.n3209 gnd 0.010868f
C5717 vdd.n3210 gnd 0.010868f
C5718 vdd.n3211 gnd 0.008748f
C5719 vdd.n3212 gnd 0.008748f
C5720 vdd.n3213 gnd 0.010868f
C5721 vdd.n3214 gnd 0.010868f
C5722 vdd.n3215 gnd 0.008748f
C5723 vdd.n3216 gnd 0.008748f
C5724 vdd.n3217 gnd 0.010868f
C5725 vdd.n3218 gnd 0.010868f
C5726 vdd.n3219 gnd 0.008748f
C5727 vdd.n3220 gnd 0.008748f
C5728 vdd.n3221 gnd 0.010868f
C5729 vdd.n3222 gnd 0.010868f
C5730 vdd.n3223 gnd 0.008748f
C5731 vdd.n3224 gnd 0.010868f
C5732 vdd.n3225 gnd 0.010868f
C5733 vdd.n3226 gnd 0.008748f
C5734 vdd.n3227 gnd 0.010868f
C5735 vdd.n3228 gnd 0.010868f
C5736 vdd.n3229 gnd 0.010868f
C5737 vdd.n3230 gnd 0.017845f
C5738 vdd.n3231 gnd 0.010868f
C5739 vdd.n3232 gnd 0.010868f
C5740 vdd.n3233 gnd 0.005948f
C5741 vdd.n3234 gnd 0.008748f
C5742 vdd.n3235 gnd 0.010868f
C5743 vdd.n3236 gnd 0.010868f
C5744 vdd.n3237 gnd 0.008748f
C5745 vdd.n3238 gnd 0.008748f
C5746 vdd.n3239 gnd 0.010868f
C5747 vdd.n3240 gnd 0.010868f
C5748 vdd.n3241 gnd 0.008748f
C5749 vdd.n3242 gnd 0.008748f
C5750 vdd.n3243 gnd 0.010868f
C5751 vdd.n3244 gnd 0.010868f
C5752 vdd.n3245 gnd 0.008748f
C5753 vdd.n3246 gnd 0.008748f
C5754 vdd.n3247 gnd 0.010868f
C5755 vdd.n3248 gnd 0.010868f
C5756 vdd.n3249 gnd 0.008748f
C5757 vdd.n3250 gnd 0.008748f
C5758 vdd.n3251 gnd 0.010868f
C5759 vdd.n3252 gnd 0.010868f
C5760 vdd.n3253 gnd 0.008748f
C5761 vdd.n3254 gnd 0.008748f
C5762 vdd.n3255 gnd 0.010868f
C5763 vdd.n3256 gnd 0.010868f
C5764 vdd.n3257 gnd 0.008748f
C5765 vdd.n3258 gnd 0.008748f
C5766 vdd.n3259 gnd 0.010868f
C5767 vdd.n3260 gnd 0.010868f
C5768 vdd.n3261 gnd 0.008748f
C5769 vdd.n3262 gnd 0.008748f
C5770 vdd.n3263 gnd 0.010868f
C5771 vdd.n3264 gnd 0.010868f
C5772 vdd.n3265 gnd 0.008748f
C5773 vdd.n3266 gnd 0.008748f
C5774 vdd.n3267 gnd 0.010868f
C5775 vdd.n3268 gnd 0.010868f
C5776 vdd.n3269 gnd 0.008748f
C5777 vdd.n3270 gnd 0.010868f
C5778 vdd.n3271 gnd 0.010868f
C5779 vdd.n3272 gnd 0.008748f
C5780 vdd.n3273 gnd 0.010868f
C5781 vdd.n3274 gnd 0.010868f
C5782 vdd.n3275 gnd 0.010868f
C5783 vdd.t85 gnd 0.133709f
C5784 vdd.t86 gnd 0.142898f
C5785 vdd.t84 gnd 0.174622f
C5786 vdd.n3276 gnd 0.223841f
C5787 vdd.n3277 gnd 0.188067f
C5788 vdd.n3278 gnd 0.017845f
C5789 vdd.n3279 gnd 0.010868f
C5790 vdd.n3280 gnd 0.010868f
C5791 vdd.n3281 gnd 0.007304f
C5792 vdd.n3282 gnd 0.008748f
C5793 vdd.n3283 gnd 0.010868f
C5794 vdd.n3284 gnd 0.010868f
C5795 vdd.n3285 gnd 0.008748f
C5796 vdd.n3286 gnd 0.008748f
C5797 vdd.n3287 gnd 0.010868f
C5798 vdd.n3288 gnd 0.010868f
C5799 vdd.n3289 gnd 0.008748f
C5800 vdd.n3290 gnd 0.008748f
C5801 vdd.n3291 gnd 0.010868f
C5802 vdd.n3292 gnd 0.010868f
C5803 vdd.n3293 gnd 0.008748f
C5804 vdd.n3294 gnd 0.008748f
C5805 vdd.n3295 gnd 0.010868f
C5806 vdd.n3296 gnd 0.010868f
C5807 vdd.n3297 gnd 0.008748f
C5808 vdd.n3298 gnd 0.008748f
C5809 vdd.n3299 gnd 0.010868f
C5810 vdd.n3300 gnd 0.010868f
C5811 vdd.n3301 gnd 0.008748f
C5812 vdd.n3302 gnd 0.008748f
C5813 vdd.n3303 gnd 0.010868f
C5814 vdd.n3304 gnd 0.010868f
C5815 vdd.n3305 gnd 0.008748f
C5816 vdd.n3306 gnd 0.008748f
C5817 vdd.n3308 gnd 0.826161f
C5818 vdd.n3310 gnd 0.008748f
C5819 vdd.n3311 gnd 0.008748f
C5820 vdd.n3312 gnd 0.007261f
C5821 vdd.n3313 gnd 0.026855f
C5822 vdd.n3315 gnd 9.874049f
C5823 vdd.n3316 gnd 0.026855f
C5824 vdd.n3317 gnd 0.004155f
C5825 vdd.n3318 gnd 0.026855f
C5826 vdd.n3319 gnd 0.026291f
C5827 vdd.n3320 gnd 0.010868f
C5828 vdd.n3321 gnd 0.008748f
C5829 vdd.n3322 gnd 0.010868f
C5830 vdd.n3323 gnd 0.671969f
C5831 vdd.n3324 gnd 0.010868f
C5832 vdd.n3325 gnd 0.008748f
C5833 vdd.n3326 gnd 0.010868f
C5834 vdd.n3327 gnd 0.010868f
C5835 vdd.n3328 gnd 0.010868f
C5836 vdd.n3329 gnd 0.008748f
C5837 vdd.n3330 gnd 0.010868f
C5838 vdd.n3331 gnd 1.11069f
C5839 vdd.n3332 gnd 0.010868f
C5840 vdd.n3333 gnd 0.008748f
C5841 vdd.n3334 gnd 0.010868f
C5842 vdd.n3335 gnd 0.010868f
C5843 vdd.n3336 gnd 0.010868f
C5844 vdd.n3337 gnd 0.008748f
C5845 vdd.n3338 gnd 0.010868f
C5846 vdd.n3339 gnd 0.716396f
C5847 vdd.n3340 gnd 0.760824f
C5848 vdd.n3341 gnd 0.010868f
C5849 vdd.n3342 gnd 0.008748f
C5850 vdd.n3343 gnd 0.010868f
C5851 vdd.n3344 gnd 0.010868f
C5852 vdd.n3345 gnd 0.010868f
C5853 vdd.n3346 gnd 0.008748f
C5854 vdd.n3347 gnd 0.010868f
C5855 vdd.n3348 gnd 0.921874f
C5856 vdd.n3349 gnd 0.010868f
C5857 vdd.n3350 gnd 0.008748f
C5858 vdd.n3351 gnd 0.010868f
C5859 vdd.n3352 gnd 0.010868f
C5860 vdd.n3353 gnd 0.010868f
C5861 vdd.n3354 gnd 0.008748f
C5862 vdd.n3355 gnd 0.010868f
C5863 vdd.t200 gnd 0.555346f
C5864 vdd.n3356 gnd 0.894107f
C5865 vdd.n3357 gnd 0.010868f
C5866 vdd.n3358 gnd 0.008748f
C5867 vdd.n3359 gnd 0.010868f
C5868 vdd.n3360 gnd 0.010868f
C5869 vdd.n3361 gnd 0.010868f
C5870 vdd.n3362 gnd 0.008748f
C5871 vdd.n3363 gnd 0.010868f
C5872 vdd.n3364 gnd 0.705289f
C5873 vdd.n3365 gnd 0.010868f
C5874 vdd.n3366 gnd 0.008748f
C5875 vdd.n3367 gnd 0.010868f
C5876 vdd.n3368 gnd 0.010868f
C5877 vdd.n3369 gnd 0.010868f
C5878 vdd.n3370 gnd 0.008748f
C5879 vdd.n3371 gnd 0.010868f
C5880 vdd.n3372 gnd 0.883f
C5881 vdd.n3373 gnd 0.59422f
C5882 vdd.n3374 gnd 0.010868f
C5883 vdd.n3375 gnd 0.008748f
C5884 vdd.n3376 gnd 0.010868f
C5885 vdd.n3377 gnd 0.010868f
C5886 vdd.n3378 gnd 0.010868f
C5887 vdd.n3379 gnd 0.008748f
C5888 vdd.n3380 gnd 0.010868f
C5889 vdd.n3381 gnd 0.783038f
C5890 vdd.n3382 gnd 0.010868f
C5891 vdd.n3383 gnd 0.008748f
C5892 vdd.n3384 gnd 0.010868f
C5893 vdd.n3385 gnd 0.010868f
C5894 vdd.n3386 gnd 0.010868f
C5895 vdd.n3387 gnd 0.010868f
C5896 vdd.n3388 gnd 0.010868f
C5897 vdd.n3389 gnd 0.008748f
C5898 vdd.n3390 gnd 0.008748f
C5899 vdd.n3391 gnd 0.010868f
C5900 vdd.t173 gnd 0.555346f
C5901 vdd.n3392 gnd 0.921874f
C5902 vdd.n3393 gnd 0.010868f
C5903 vdd.n3394 gnd 0.008748f
C5904 vdd.n3395 gnd 0.010868f
C5905 vdd.n3396 gnd 0.010868f
C5906 vdd.n3397 gnd 0.010868f
C5907 vdd.n3398 gnd 0.008748f
C5908 vdd.n3399 gnd 0.010868f
C5909 vdd.n3400 gnd 0.871893f
C5910 vdd.n3401 gnd 0.010868f
C5911 vdd.n3402 gnd 0.010868f
C5912 vdd.n3403 gnd 0.008748f
C5913 vdd.n3404 gnd 0.008748f
C5914 vdd.n3405 gnd 0.010868f
C5915 vdd.n3406 gnd 0.010868f
C5916 vdd.n3407 gnd 0.010868f
C5917 vdd.n3408 gnd 0.008748f
C5918 vdd.n3409 gnd 0.010868f
C5919 vdd.n3410 gnd 0.008748f
C5920 vdd.n3411 gnd 0.008748f
C5921 vdd.n3412 gnd 0.010868f
C5922 vdd.n3413 gnd 0.010868f
C5923 vdd.n3414 gnd 0.010868f
C5924 vdd.n3415 gnd 0.008748f
C5925 vdd.n3416 gnd 0.010868f
C5926 vdd.n3417 gnd 0.008748f
C5927 vdd.n3418 gnd 0.008748f
C5928 vdd.n3419 gnd 0.010868f
C5929 vdd.n3420 gnd 0.010868f
C5930 vdd.n3421 gnd 0.010868f
C5931 vdd.n3422 gnd 0.008748f
C5932 vdd.n3423 gnd 0.921874f
C5933 vdd.n3424 gnd 0.010868f
C5934 vdd.n3425 gnd 0.008748f
C5935 vdd.n3426 gnd 0.008748f
C5936 vdd.n3427 gnd 0.010868f
C5937 vdd.n3428 gnd 0.010868f
C5938 vdd.n3429 gnd 0.010868f
C5939 vdd.n3430 gnd 0.008748f
C5940 vdd.n3431 gnd 0.010868f
C5941 vdd.n3432 gnd 0.008748f
C5942 vdd.n3433 gnd 0.008748f
C5943 vdd.n3434 gnd 0.010868f
C5944 vdd.n3435 gnd 0.010868f
C5945 vdd.n3436 gnd 0.010868f
C5946 vdd.n3437 gnd 0.008748f
C5947 vdd.n3438 gnd 0.010868f
C5948 vdd.n3439 gnd 0.008748f
C5949 vdd.n3440 gnd 0.007261f
C5950 vdd.n3441 gnd 0.026291f
C5951 vdd.n3442 gnd 0.026855f
C5952 vdd.n3443 gnd 0.004155f
C5953 vdd.n3444 gnd 0.026855f
C5954 vdd.n3446 gnd 2.63234f
C5955 vdd.n3447 gnd 1.63827f
C5956 vdd.n3448 gnd 0.026291f
C5957 vdd.n3449 gnd 0.007261f
C5958 vdd.n3450 gnd 0.008748f
C5959 vdd.n3451 gnd 0.008748f
C5960 vdd.n3452 gnd 0.010868f
C5961 vdd.n3453 gnd 1.11069f
C5962 vdd.n3454 gnd 1.11069f
C5963 vdd.n3455 gnd 1.01628f
C5964 vdd.n3456 gnd 0.010868f
C5965 vdd.n3457 gnd 0.008748f
C5966 vdd.n3458 gnd 0.008748f
C5967 vdd.n3459 gnd 0.008748f
C5968 vdd.n3460 gnd 0.010868f
C5969 vdd.n3461 gnd 0.827466f
C5970 vdd.t253 gnd 0.555346f
C5971 vdd.n3462 gnd 0.838572f
C5972 vdd.n3463 gnd 0.638648f
C5973 vdd.n3464 gnd 0.010868f
C5974 vdd.n3465 gnd 0.008748f
C5975 vdd.n3466 gnd 0.008748f
C5976 vdd.n3467 gnd 0.008748f
C5977 vdd.n3468 gnd 0.010868f
C5978 vdd.n3469 gnd 0.660862f
C5979 vdd.n3470 gnd 0.816359f
C5980 vdd.t211 gnd 0.555346f
C5981 vdd.n3471 gnd 0.849679f
C5982 vdd.n3472 gnd 0.010868f
C5983 vdd.n3473 gnd 0.008748f
C5984 vdd.n3474 gnd 0.008748f
C5985 vdd.n3475 gnd 0.008748f
C5986 vdd.n3476 gnd 0.010868f
C5987 vdd.n3477 gnd 0.921874f
C5988 vdd.t155 gnd 0.555346f
C5989 vdd.n3478 gnd 0.671969f
C5990 vdd.n3479 gnd 0.805252f
C5991 vdd.n3480 gnd 0.010868f
C5992 vdd.n3481 gnd 0.008748f
C5993 vdd.n3482 gnd 0.008748f
C5994 vdd.n3483 gnd 0.008748f
C5995 vdd.n3484 gnd 0.010868f
C5996 vdd.n3485 gnd 0.616434f
C5997 vdd.t167 gnd 0.555346f
C5998 vdd.n3486 gnd 0.921874f
C5999 vdd.t157 gnd 0.555346f
C6000 vdd.n3487 gnd 0.683076f
C6001 vdd.n3488 gnd 0.010868f
C6002 vdd.n3489 gnd 0.008748f
C6003 vdd.n3490 gnd 0.008353f
C6004 vdd.n3491 gnd 0.641055f
C6005 vdd.n3492 gnd 2.91077f
C6006 a_n8300_8799.n0 gnd 2.72381f
C6007 a_n8300_8799.n1 gnd 1.65029f
C6008 a_n8300_8799.n2 gnd 3.77569f
C6009 a_n8300_8799.n3 gnd 0.205925f
C6010 a_n8300_8799.n4 gnd 0.282763f
C6011 a_n8300_8799.n5 gnd 0.205925f
C6012 a_n8300_8799.n6 gnd 0.205925f
C6013 a_n8300_8799.n7 gnd 0.205925f
C6014 a_n8300_8799.n8 gnd 0.205925f
C6015 a_n8300_8799.n9 gnd 0.205925f
C6016 a_n8300_8799.n10 gnd 0.214125f
C6017 a_n8300_8799.n11 gnd 0.205925f
C6018 a_n8300_8799.n12 gnd 0.282763f
C6019 a_n8300_8799.n13 gnd 0.205925f
C6020 a_n8300_8799.n14 gnd 0.205925f
C6021 a_n8300_8799.n15 gnd 0.205925f
C6022 a_n8300_8799.n16 gnd 0.205925f
C6023 a_n8300_8799.n17 gnd 0.205925f
C6024 a_n8300_8799.n18 gnd 0.214125f
C6025 a_n8300_8799.n19 gnd 0.205925f
C6026 a_n8300_8799.n20 gnd 0.44633f
C6027 a_n8300_8799.n21 gnd 0.205925f
C6028 a_n8300_8799.n22 gnd 0.205925f
C6029 a_n8300_8799.n23 gnd 0.205925f
C6030 a_n8300_8799.n24 gnd 0.205925f
C6031 a_n8300_8799.n25 gnd 0.205925f
C6032 a_n8300_8799.n26 gnd 0.214125f
C6033 a_n8300_8799.n27 gnd 0.205925f
C6034 a_n8300_8799.n28 gnd 0.317088f
C6035 a_n8300_8799.n29 gnd 0.205925f
C6036 a_n8300_8799.n30 gnd 0.205925f
C6037 a_n8300_8799.n31 gnd 0.205925f
C6038 a_n8300_8799.n32 gnd 0.205925f
C6039 a_n8300_8799.n33 gnd 0.205925f
C6040 a_n8300_8799.n34 gnd 0.1798f
C6041 a_n8300_8799.n35 gnd 0.205925f
C6042 a_n8300_8799.n36 gnd 0.317088f
C6043 a_n8300_8799.n37 gnd 0.205925f
C6044 a_n8300_8799.n38 gnd 0.205925f
C6045 a_n8300_8799.n39 gnd 0.205925f
C6046 a_n8300_8799.n40 gnd 0.205925f
C6047 a_n8300_8799.n41 gnd 0.205925f
C6048 a_n8300_8799.n42 gnd 0.1798f
C6049 a_n8300_8799.n43 gnd 0.205925f
C6050 a_n8300_8799.n44 gnd 0.317088f
C6051 a_n8300_8799.n45 gnd 0.205925f
C6052 a_n8300_8799.n46 gnd 0.205925f
C6053 a_n8300_8799.n47 gnd 0.205925f
C6054 a_n8300_8799.n48 gnd 0.205925f
C6055 a_n8300_8799.n49 gnd 0.205925f
C6056 a_n8300_8799.n50 gnd 0.343367f
C6057 a_n8300_8799.n51 gnd 1.50927f
C6058 a_n8300_8799.n52 gnd 2.52406f
C6059 a_n8300_8799.n53 gnd 0.247915f
C6060 a_n8300_8799.n54 gnd 0.003624f
C6061 a_n8300_8799.n55 gnd 0.009554f
C6062 a_n8300_8799.n56 gnd 0.010439f
C6063 a_n8300_8799.n57 gnd 0.005516f
C6064 a_n8300_8799.n59 gnd 0.004628f
C6065 a_n8300_8799.n60 gnd 0.01001f
C6066 a_n8300_8799.n61 gnd 0.01001f
C6067 a_n8300_8799.n62 gnd 0.004628f
C6068 a_n8300_8799.n64 gnd 0.005516f
C6069 a_n8300_8799.n65 gnd 0.010439f
C6070 a_n8300_8799.n66 gnd 0.009554f
C6071 a_n8300_8799.n67 gnd 0.003624f
C6072 a_n8300_8799.n68 gnd 0.247915f
C6073 a_n8300_8799.n69 gnd 0.003624f
C6074 a_n8300_8799.n70 gnd 0.009554f
C6075 a_n8300_8799.n71 gnd 0.010439f
C6076 a_n8300_8799.n72 gnd 0.005516f
C6077 a_n8300_8799.n74 gnd 0.004628f
C6078 a_n8300_8799.n75 gnd 0.01001f
C6079 a_n8300_8799.n76 gnd 0.01001f
C6080 a_n8300_8799.n77 gnd 0.004628f
C6081 a_n8300_8799.n79 gnd 0.005516f
C6082 a_n8300_8799.n80 gnd 0.010439f
C6083 a_n8300_8799.n81 gnd 0.009554f
C6084 a_n8300_8799.n82 gnd 0.003624f
C6085 a_n8300_8799.n83 gnd 0.247915f
C6086 a_n8300_8799.n84 gnd 0.003624f
C6087 a_n8300_8799.n85 gnd 0.009554f
C6088 a_n8300_8799.n86 gnd 0.010439f
C6089 a_n8300_8799.n87 gnd 0.005516f
C6090 a_n8300_8799.n89 gnd 0.004628f
C6091 a_n8300_8799.n90 gnd 0.01001f
C6092 a_n8300_8799.n91 gnd 0.01001f
C6093 a_n8300_8799.n92 gnd 0.004628f
C6094 a_n8300_8799.n94 gnd 0.005516f
C6095 a_n8300_8799.n95 gnd 0.010439f
C6096 a_n8300_8799.n96 gnd 0.009554f
C6097 a_n8300_8799.n97 gnd 0.003624f
C6098 a_n8300_8799.n98 gnd 0.003624f
C6099 a_n8300_8799.n99 gnd 0.009554f
C6100 a_n8300_8799.n100 gnd 0.010439f
C6101 a_n8300_8799.n101 gnd 0.005516f
C6102 a_n8300_8799.n103 gnd 0.004628f
C6103 a_n8300_8799.n104 gnd 0.01001f
C6104 a_n8300_8799.n105 gnd 0.01001f
C6105 a_n8300_8799.n106 gnd 0.004628f
C6106 a_n8300_8799.n108 gnd 0.005516f
C6107 a_n8300_8799.n109 gnd 0.010439f
C6108 a_n8300_8799.n110 gnd 0.009554f
C6109 a_n8300_8799.n111 gnd 0.003624f
C6110 a_n8300_8799.n112 gnd 0.247915f
C6111 a_n8300_8799.n113 gnd 0.003624f
C6112 a_n8300_8799.n114 gnd 0.009554f
C6113 a_n8300_8799.n115 gnd 0.010439f
C6114 a_n8300_8799.n116 gnd 0.005516f
C6115 a_n8300_8799.n118 gnd 0.004628f
C6116 a_n8300_8799.n119 gnd 0.01001f
C6117 a_n8300_8799.n120 gnd 0.01001f
C6118 a_n8300_8799.n121 gnd 0.004628f
C6119 a_n8300_8799.n123 gnd 0.005516f
C6120 a_n8300_8799.n124 gnd 0.010439f
C6121 a_n8300_8799.n125 gnd 0.009554f
C6122 a_n8300_8799.n126 gnd 0.003624f
C6123 a_n8300_8799.n127 gnd 0.247915f
C6124 a_n8300_8799.n128 gnd 0.003624f
C6125 a_n8300_8799.n129 gnd 0.009554f
C6126 a_n8300_8799.n130 gnd 0.010439f
C6127 a_n8300_8799.n131 gnd 0.005516f
C6128 a_n8300_8799.n133 gnd 0.004628f
C6129 a_n8300_8799.n134 gnd 0.01001f
C6130 a_n8300_8799.n135 gnd 0.01001f
C6131 a_n8300_8799.n136 gnd 0.004628f
C6132 a_n8300_8799.n138 gnd 0.005516f
C6133 a_n8300_8799.n139 gnd 0.010439f
C6134 a_n8300_8799.n140 gnd 0.009554f
C6135 a_n8300_8799.n141 gnd 0.003624f
C6136 a_n8300_8799.n142 gnd 0.247915f
C6137 a_n8300_8799.t23 gnd 0.142832f
C6138 a_n8300_8799.t17 gnd 0.142832f
C6139 a_n8300_8799.t24 gnd 0.142832f
C6140 a_n8300_8799.n143 gnd 1.12654f
C6141 a_n8300_8799.t5 gnd 0.142832f
C6142 a_n8300_8799.t7 gnd 0.142832f
C6143 a_n8300_8799.n144 gnd 1.12468f
C6144 a_n8300_8799.t16 gnd 0.142832f
C6145 a_n8300_8799.t8 gnd 0.142832f
C6146 a_n8300_8799.n145 gnd 1.12468f
C6147 a_n8300_8799.t10 gnd 0.142832f
C6148 a_n8300_8799.t13 gnd 0.142832f
C6149 a_n8300_8799.n146 gnd 1.12468f
C6150 a_n8300_8799.n147 gnd 3.15899f
C6151 a_n8300_8799.t2 gnd 0.111092f
C6152 a_n8300_8799.t28 gnd 0.111092f
C6153 a_n8300_8799.n148 gnd 0.98454f
C6154 a_n8300_8799.t11 gnd 0.111092f
C6155 a_n8300_8799.t29 gnd 0.111092f
C6156 a_n8300_8799.n149 gnd 0.981645f
C6157 a_n8300_8799.t25 gnd 0.111092f
C6158 a_n8300_8799.t14 gnd 0.111092f
C6159 a_n8300_8799.n150 gnd 0.984539f
C6160 a_n8300_8799.t20 gnd 0.111092f
C6161 a_n8300_8799.t22 gnd 0.111092f
C6162 a_n8300_8799.n151 gnd 0.981644f
C6163 a_n8300_8799.t1 gnd 0.111092f
C6164 a_n8300_8799.t27 gnd 0.111092f
C6165 a_n8300_8799.n152 gnd 0.984539f
C6166 a_n8300_8799.t31 gnd 0.111092f
C6167 a_n8300_8799.t19 gnd 0.111092f
C6168 a_n8300_8799.n153 gnd 0.981644f
C6169 a_n8300_8799.t12 gnd 0.111092f
C6170 a_n8300_8799.t15 gnd 0.111092f
C6171 a_n8300_8799.n154 gnd 0.981645f
C6172 a_n8300_8799.t26 gnd 0.111092f
C6173 a_n8300_8799.t6 gnd 0.111092f
C6174 a_n8300_8799.n155 gnd 0.981645f
C6175 a_n8300_8799.t84 gnd 0.592248f
C6176 a_n8300_8799.n156 gnd 0.266638f
C6177 a_n8300_8799.t32 gnd 0.592248f
C6178 a_n8300_8799.t63 gnd 0.592248f
C6179 a_n8300_8799.n157 gnd 0.268548f
C6180 a_n8300_8799.t64 gnd 0.592248f
C6181 a_n8300_8799.t78 gnd 0.592248f
C6182 a_n8300_8799.n158 gnd 0.261812f
C6183 a_n8300_8799.t130 gnd 0.592248f
C6184 a_n8300_8799.t133 gnd 0.592248f
C6185 a_n8300_8799.n159 gnd 0.265753f
C6186 a_n8300_8799.t94 gnd 0.592248f
C6187 a_n8300_8799.t138 gnd 0.592248f
C6188 a_n8300_8799.t99 gnd 0.603458f
C6189 a_n8300_8799.n160 gnd 0.248275f
C6190 a_n8300_8799.n161 gnd 0.268917f
C6191 a_n8300_8799.t61 gnd 0.592248f
C6192 a_n8300_8799.n162 gnd 0.266638f
C6193 a_n8300_8799.n163 gnd 0.262446f
C6194 a_n8300_8799.t132 gnd 0.592248f
C6195 a_n8300_8799.n164 gnd 0.261177f
C6196 a_n8300_8799.t79 gnd 0.592248f
C6197 a_n8300_8799.n165 gnd 0.268295f
C6198 a_n8300_8799.t110 gnd 0.592248f
C6199 a_n8300_8799.n166 gnd 0.268548f
C6200 a_n8300_8799.n167 gnd 0.266182f
C6201 a_n8300_8799.t77 gnd 0.592248f
C6202 a_n8300_8799.n168 gnd 0.261812f
C6203 a_n8300_8799.t107 gnd 0.592248f
C6204 a_n8300_8799.n169 gnd 0.266182f
C6205 a_n8300_8799.n170 gnd 0.268295f
C6206 a_n8300_8799.t104 gnd 0.592248f
C6207 a_n8300_8799.n171 gnd 0.265753f
C6208 a_n8300_8799.n172 gnd 0.261177f
C6209 a_n8300_8799.t62 gnd 0.592248f
C6210 a_n8300_8799.n173 gnd 0.262446f
C6211 a_n8300_8799.t131 gnd 0.592248f
C6212 a_n8300_8799.n174 gnd 0.268917f
C6213 a_n8300_8799.t43 gnd 0.603448f
C6214 a_n8300_8799.t96 gnd 0.592248f
C6215 a_n8300_8799.n175 gnd 0.266638f
C6216 a_n8300_8799.t42 gnd 0.592248f
C6217 a_n8300_8799.t75 gnd 0.592248f
C6218 a_n8300_8799.n176 gnd 0.268548f
C6219 a_n8300_8799.t76 gnd 0.592248f
C6220 a_n8300_8799.t86 gnd 0.592248f
C6221 a_n8300_8799.n177 gnd 0.261812f
C6222 a_n8300_8799.t144 gnd 0.592248f
C6223 a_n8300_8799.t149 gnd 0.592248f
C6224 a_n8300_8799.n178 gnd 0.265753f
C6225 a_n8300_8799.t108 gnd 0.592248f
C6226 a_n8300_8799.t151 gnd 0.592248f
C6227 a_n8300_8799.t115 gnd 0.603458f
C6228 a_n8300_8799.n179 gnd 0.248275f
C6229 a_n8300_8799.n180 gnd 0.268917f
C6230 a_n8300_8799.t71 gnd 0.592248f
C6231 a_n8300_8799.n181 gnd 0.266638f
C6232 a_n8300_8799.n182 gnd 0.262446f
C6233 a_n8300_8799.t146 gnd 0.592248f
C6234 a_n8300_8799.n183 gnd 0.261177f
C6235 a_n8300_8799.t89 gnd 0.592248f
C6236 a_n8300_8799.n184 gnd 0.268295f
C6237 a_n8300_8799.t127 gnd 0.592248f
C6238 a_n8300_8799.n185 gnd 0.268548f
C6239 a_n8300_8799.n186 gnd 0.266182f
C6240 a_n8300_8799.t85 gnd 0.592248f
C6241 a_n8300_8799.n187 gnd 0.261812f
C6242 a_n8300_8799.t125 gnd 0.592248f
C6243 a_n8300_8799.n188 gnd 0.266182f
C6244 a_n8300_8799.n189 gnd 0.268295f
C6245 a_n8300_8799.t121 gnd 0.592248f
C6246 a_n8300_8799.n190 gnd 0.265753f
C6247 a_n8300_8799.n191 gnd 0.261177f
C6248 a_n8300_8799.t72 gnd 0.592248f
C6249 a_n8300_8799.n192 gnd 0.262446f
C6250 a_n8300_8799.t147 gnd 0.592248f
C6251 a_n8300_8799.n193 gnd 0.268917f
C6252 a_n8300_8799.t55 gnd 0.603448f
C6253 a_n8300_8799.n194 gnd 0.890363f
C6254 a_n8300_8799.t100 gnd 0.592248f
C6255 a_n8300_8799.n195 gnd 0.266638f
C6256 a_n8300_8799.t83 gnd 0.592248f
C6257 a_n8300_8799.t137 gnd 0.592248f
C6258 a_n8300_8799.n196 gnd 0.268548f
C6259 a_n8300_8799.t109 gnd 0.592248f
C6260 a_n8300_8799.t33 gnd 0.592248f
C6261 a_n8300_8799.n197 gnd 0.261812f
C6262 a_n8300_8799.t134 gnd 0.592248f
C6263 a_n8300_8799.t82 gnd 0.592248f
C6264 a_n8300_8799.n198 gnd 0.265753f
C6265 a_n8300_8799.t44 gnd 0.592248f
C6266 a_n8300_8799.t66 gnd 0.592248f
C6267 a_n8300_8799.t117 gnd 0.603458f
C6268 a_n8300_8799.n199 gnd 0.248275f
C6269 a_n8300_8799.n200 gnd 0.268917f
C6270 a_n8300_8799.t87 gnd 0.592248f
C6271 a_n8300_8799.n201 gnd 0.266638f
C6272 a_n8300_8799.n202 gnd 0.262446f
C6273 a_n8300_8799.t105 gnd 0.592248f
C6274 a_n8300_8799.n203 gnd 0.261177f
C6275 a_n8300_8799.t126 gnd 0.592248f
C6276 a_n8300_8799.n204 gnd 0.268295f
C6277 a_n8300_8799.t73 gnd 0.592248f
C6278 a_n8300_8799.n205 gnd 0.268548f
C6279 a_n8300_8799.n206 gnd 0.266182f
C6280 a_n8300_8799.t49 gnd 0.592248f
C6281 a_n8300_8799.n207 gnd 0.261812f
C6282 a_n8300_8799.t90 gnd 0.592248f
C6283 a_n8300_8799.n208 gnd 0.266182f
C6284 a_n8300_8799.n209 gnd 0.268295f
C6285 a_n8300_8799.t143 gnd 0.592248f
C6286 a_n8300_8799.n210 gnd 0.265753f
C6287 a_n8300_8799.n211 gnd 0.261177f
C6288 a_n8300_8799.t38 gnd 0.592248f
C6289 a_n8300_8799.n212 gnd 0.262446f
C6290 a_n8300_8799.t53 gnd 0.592248f
C6291 a_n8300_8799.n213 gnd 0.268917f
C6292 a_n8300_8799.t122 gnd 0.603448f
C6293 a_n8300_8799.n214 gnd 1.55679f
C6294 a_n8300_8799.t81 gnd 0.603448f
C6295 a_n8300_8799.t57 gnd 0.592248f
C6296 a_n8300_8799.t136 gnd 0.592248f
C6297 a_n8300_8799.n215 gnd 0.266638f
C6298 a_n8300_8799.t98 gnd 0.592248f
C6299 a_n8300_8799.t95 gnd 0.592248f
C6300 a_n8300_8799.t35 gnd 0.592248f
C6301 a_n8300_8799.n216 gnd 0.265753f
C6302 a_n8300_8799.t103 gnd 0.592248f
C6303 a_n8300_8799.t102 gnd 0.592248f
C6304 a_n8300_8799.t37 gnd 0.592248f
C6305 a_n8300_8799.n217 gnd 0.266182f
C6306 a_n8300_8799.t36 gnd 0.592248f
C6307 a_n8300_8799.t124 gnd 0.592248f
C6308 a_n8300_8799.t52 gnd 0.592248f
C6309 a_n8300_8799.n218 gnd 0.266182f
C6310 a_n8300_8799.t41 gnd 0.592248f
C6311 a_n8300_8799.t128 gnd 0.592248f
C6312 a_n8300_8799.t80 gnd 0.592248f
C6313 a_n8300_8799.n219 gnd 0.265753f
C6314 a_n8300_8799.t56 gnd 0.592248f
C6315 a_n8300_8799.t148 gnd 0.592248f
C6316 a_n8300_8799.t97 gnd 0.592248f
C6317 a_n8300_8799.n220 gnd 0.266638f
C6318 a_n8300_8799.t141 gnd 0.603458f
C6319 a_n8300_8799.n221 gnd 0.248275f
C6320 a_n8300_8799.t59 gnd 0.592248f
C6321 a_n8300_8799.n222 gnd 0.268917f
C6322 a_n8300_8799.n223 gnd 0.262446f
C6323 a_n8300_8799.n224 gnd 0.261177f
C6324 a_n8300_8799.n225 gnd 0.268295f
C6325 a_n8300_8799.n226 gnd 0.268548f
C6326 a_n8300_8799.n227 gnd 0.261812f
C6327 a_n8300_8799.n228 gnd 0.261812f
C6328 a_n8300_8799.n229 gnd 0.268548f
C6329 a_n8300_8799.n230 gnd 0.268295f
C6330 a_n8300_8799.n231 gnd 0.261177f
C6331 a_n8300_8799.n232 gnd 0.262446f
C6332 a_n8300_8799.n233 gnd 0.268917f
C6333 a_n8300_8799.t92 gnd 0.603448f
C6334 a_n8300_8799.t68 gnd 0.592248f
C6335 a_n8300_8799.t150 gnd 0.592248f
C6336 a_n8300_8799.n234 gnd 0.266638f
C6337 a_n8300_8799.t113 gnd 0.592248f
C6338 a_n8300_8799.t112 gnd 0.592248f
C6339 a_n8300_8799.t46 gnd 0.592248f
C6340 a_n8300_8799.n235 gnd 0.265753f
C6341 a_n8300_8799.t120 gnd 0.592248f
C6342 a_n8300_8799.t119 gnd 0.592248f
C6343 a_n8300_8799.t48 gnd 0.592248f
C6344 a_n8300_8799.n236 gnd 0.266182f
C6345 a_n8300_8799.t47 gnd 0.592248f
C6346 a_n8300_8799.t140 gnd 0.592248f
C6347 a_n8300_8799.t65 gnd 0.592248f
C6348 a_n8300_8799.n237 gnd 0.266182f
C6349 a_n8300_8799.t51 gnd 0.592248f
C6350 a_n8300_8799.t142 gnd 0.592248f
C6351 a_n8300_8799.t93 gnd 0.592248f
C6352 a_n8300_8799.n238 gnd 0.265753f
C6353 a_n8300_8799.t69 gnd 0.592248f
C6354 a_n8300_8799.t39 gnd 0.592248f
C6355 a_n8300_8799.t114 gnd 0.592248f
C6356 a_n8300_8799.n239 gnd 0.266638f
C6357 a_n8300_8799.t34 gnd 0.603458f
C6358 a_n8300_8799.n240 gnd 0.248275f
C6359 a_n8300_8799.t70 gnd 0.592248f
C6360 a_n8300_8799.n241 gnd 0.268917f
C6361 a_n8300_8799.n242 gnd 0.262446f
C6362 a_n8300_8799.n243 gnd 0.261177f
C6363 a_n8300_8799.n244 gnd 0.268295f
C6364 a_n8300_8799.n245 gnd 0.268548f
C6365 a_n8300_8799.n246 gnd 0.261812f
C6366 a_n8300_8799.n247 gnd 0.261812f
C6367 a_n8300_8799.n248 gnd 0.268548f
C6368 a_n8300_8799.n249 gnd 0.268295f
C6369 a_n8300_8799.n250 gnd 0.261177f
C6370 a_n8300_8799.n251 gnd 0.262446f
C6371 a_n8300_8799.n252 gnd 0.268917f
C6372 a_n8300_8799.n253 gnd 0.890363f
C6373 a_n8300_8799.t123 gnd 0.603448f
C6374 a_n8300_8799.t54 gnd 0.592248f
C6375 a_n8300_8799.t101 gnd 0.592248f
C6376 a_n8300_8799.n254 gnd 0.266638f
C6377 a_n8300_8799.t40 gnd 0.592248f
C6378 a_n8300_8799.t60 gnd 0.592248f
C6379 a_n8300_8799.t145 gnd 0.592248f
C6380 a_n8300_8799.n255 gnd 0.265753f
C6381 a_n8300_8799.t111 gnd 0.592248f
C6382 a_n8300_8799.t139 gnd 0.592248f
C6383 a_n8300_8799.t91 gnd 0.592248f
C6384 a_n8300_8799.n256 gnd 0.266182f
C6385 a_n8300_8799.t118 gnd 0.592248f
C6386 a_n8300_8799.t50 gnd 0.592248f
C6387 a_n8300_8799.t135 gnd 0.592248f
C6388 a_n8300_8799.n257 gnd 0.266182f
C6389 a_n8300_8799.t74 gnd 0.592248f
C6390 a_n8300_8799.t129 gnd 0.592248f
C6391 a_n8300_8799.t58 gnd 0.592248f
C6392 a_n8300_8799.n258 gnd 0.265753f
C6393 a_n8300_8799.t106 gnd 0.592248f
C6394 a_n8300_8799.t45 gnd 0.592248f
C6395 a_n8300_8799.t88 gnd 0.592248f
C6396 a_n8300_8799.n259 gnd 0.266638f
C6397 a_n8300_8799.t116 gnd 0.603458f
C6398 a_n8300_8799.n260 gnd 0.248275f
C6399 a_n8300_8799.t67 gnd 0.592248f
C6400 a_n8300_8799.n261 gnd 0.268917f
C6401 a_n8300_8799.n262 gnd 0.262446f
C6402 a_n8300_8799.n263 gnd 0.261177f
C6403 a_n8300_8799.n264 gnd 0.268295f
C6404 a_n8300_8799.n265 gnd 0.268548f
C6405 a_n8300_8799.n266 gnd 0.261812f
C6406 a_n8300_8799.n267 gnd 0.261812f
C6407 a_n8300_8799.n268 gnd 0.268548f
C6408 a_n8300_8799.n269 gnd 0.268295f
C6409 a_n8300_8799.n270 gnd 0.261177f
C6410 a_n8300_8799.n271 gnd 0.262446f
C6411 a_n8300_8799.n272 gnd 0.268917f
C6412 a_n8300_8799.n273 gnd 1.20779f
C6413 a_n8300_8799.n274 gnd 13.8488f
C6414 a_n8300_8799.n275 gnd 4.3344f
C6415 a_n8300_8799.n276 gnd 6.28718f
C6416 a_n8300_8799.t9 gnd 0.142832f
C6417 a_n8300_8799.t3 gnd 0.142832f
C6418 a_n8300_8799.n277 gnd 1.12468f
C6419 a_n8300_8799.t21 gnd 0.142832f
C6420 a_n8300_8799.t4 gnd 0.142832f
C6421 a_n8300_8799.n278 gnd 1.12468f
C6422 a_n8300_8799.t30 gnd 0.142832f
C6423 a_n8300_8799.t18 gnd 0.142832f
C6424 a_n8300_8799.n279 gnd 1.12468f
C6425 a_n8300_8799.n280 gnd 1.01095f
C6426 a_n8300_8799.n281 gnd 1.12654f
C6427 a_n8300_8799.t0 gnd 0.142832f
.ends

