* NGSPICE file created from opamp.ext - technology: sky130A

.subckt opamp CSoutput output vdd plus minus commonsourceibias outputibias diffpairibias
+ gnd
X0 a_n5644_8799.t30 plus.t5 a_n3827_n3924.t26 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X1 gnd.t180 gnd.t177 gnd.t179 gnd.t178 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X2 gnd.t194 commonsourceibias.t46 commonsourceibias.t47 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X3 vdd.t73 a_n5644_8799.t32 CSoutput.t119 vdd.t20 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X4 a_n1986_8322.t19 a_n1996_n452.t44 vdd.t184 vdd.t183 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X5 a_n1808_13878.t11 a_n1996_n452.t19 a_n1996_n452.t20 vdd.t191 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X6 commonsourceibias.t45 commonsourceibias.t44 gnd.t14 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 gnd.t176 gnd.t174 plus.t3 gnd.t175 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X8 a_n3827_n3924.t36 plus.t6 a_n5644_8799.t29 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X9 a_n3827_n3924.t9 diffpairibias.t20 gnd.t193 gnd.t192 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X10 a_n1996_n452.t26 a_n1996_n452.t25 a_n1808_13878.t10 vdd.t77 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X11 a_n1808_13878.t9 a_n1996_n452.t9 a_n1996_n452.t10 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X12 vdd.t156 vdd.t154 vdd.t155 vdd.t129 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X13 a_n1808_13878.t19 a_n1996_n452.t45 vdd.t195 vdd.t194 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X14 CSoutput.t118 a_n5644_8799.t33 vdd.t72 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X15 a_n3827_n3924.t22 minus.t5 a_n1996_n452.t39 gnd.t287 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X16 gnd.t205 commonsourceibias.t42 commonsourceibias.t43 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X17 gnd.t240 commonsourceibias.t48 CSoutput.t71 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X18 commonsourceibias.t41 commonsourceibias.t40 gnd.t208 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 vdd.t153 vdd.t151 vdd.t152 vdd.t104 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X20 a_n1996_n452.t35 minus.t6 a_n3827_n3924.t18 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X21 output.t19 outputibias.t8 gnd.t319 gnd.t318 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X22 gnd.t173 gnd.t171 gnd.t172 gnd.t99 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X23 a_n1986_8322.t11 a_n1996_n452.t46 a_n5644_8799.t5 vdd.t185 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X24 a_n1996_n452.t42 minus.t7 a_n3827_n3924.t46 gnd.t304 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X25 commonsourceibias.t39 commonsourceibias.t38 gnd.t217 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X26 gnd.t302 commonsourceibias.t49 CSoutput.t70 gnd.t254 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X27 CSoutput.t69 commonsourceibias.t50 gnd.t290 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X28 gnd.t170 gnd.t167 gnd.t169 gnd.t168 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X29 a_n3827_n3924.t11 minus.t8 a_n1996_n452.t31 gnd.t204 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X30 CSoutput.t117 a_n5644_8799.t34 vdd.t71 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X31 vdd.t70 a_n5644_8799.t35 CSoutput.t116 vdd.t47 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X32 gnd.t50 commonsourceibias.t36 commonsourceibias.t37 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X33 a_n5644_8799.t8 a_n1996_n452.t47 a_n1986_8322.t10 vdd.t191 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X34 CSoutput.t78 a_n5644_8799.t36 vdd.t69 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X35 vdd.t68 a_n5644_8799.t37 CSoutput.t77 vdd.t63 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X36 a_n3827_n3924.t10 diffpairibias.t21 gnd.t198 gnd.t197 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X37 commonsourceibias.t35 commonsourceibias.t34 gnd.t303 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X38 CSoutput.t76 a_n5644_8799.t38 vdd.t67 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X39 vdd.t150 vdd.t148 vdd.t149 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X40 a_n3827_n3924.t28 plus.t7 a_n5644_8799.t28 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X41 CSoutput.t68 commonsourceibias.t51 gnd.t316 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X42 gnd.t188 commonsourceibias.t32 commonsourceibias.t33 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 output.t15 CSoutput.t120 vdd.t165 gnd.t264 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X44 a_n5644_8799.t27 plus.t8 a_n3827_n3924.t29 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X45 output.t18 outputibias.t9 gnd.t326 gnd.t325 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X46 a_n1808_13878.t8 a_n1996_n452.t23 a_n1996_n452.t24 vdd.t188 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X47 vdd.t66 a_n5644_8799.t39 CSoutput.t94 vdd.t63 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X48 a_n1996_n452.t29 minus.t9 a_n3827_n3924.t6 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X49 diffpairibias.t19 diffpairibias.t18 gnd.t30 gnd.t29 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X50 a_n1996_n452.t14 a_n1996_n452.t13 a_n1808_13878.t7 vdd.t173 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X51 CSoutput.t93 a_n5644_8799.t40 vdd.t65 vdd.t41 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X52 vdd.t147 vdd.t145 vdd.t146 vdd.t114 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X53 CSoutput.t67 commonsourceibias.t52 gnd.t182 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X54 gnd.t166 gnd.t164 gnd.t165 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X55 CSoutput.t66 commonsourceibias.t53 gnd.t220 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X56 plus.t0 gnd.t161 gnd.t163 gnd.t162 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X57 diffpairibias.t17 diffpairibias.t16 gnd.t279 gnd.t278 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X58 gnd.t160 gnd.t158 gnd.t159 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X59 vdd.t144 vdd.t142 vdd.t143 vdd.t93 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X60 gnd.t157 gnd.t155 gnd.t156 gnd.t84 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X61 CSoutput.t121 a_n1986_8322.t23 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X62 vdd.t64 a_n5644_8799.t41 CSoutput.t92 vdd.t63 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X63 CSoutput.t65 commonsourceibias.t54 gnd.t248 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X64 vdd.t62 a_n5644_8799.t42 CSoutput.t108 vdd.t38 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X65 CSoutput.t107 a_n5644_8799.t43 vdd.t61 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X66 gnd.t53 commonsourceibias.t55 CSoutput.t64 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X67 vdd.t60 a_n5644_8799.t44 CSoutput.t99 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X68 gnd.t221 commonsourceibias.t56 CSoutput.t63 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X69 a_n3827_n3924.t27 plus.t9 a_n5644_8799.t26 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X70 CSoutput.t62 commonsourceibias.t57 gnd.t239 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X71 CSoutput.t122 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X72 gnd.t154 gnd.t152 gnd.t153 gnd.t99 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X73 CSoutput.t98 a_n5644_8799.t45 vdd.t59 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 CSoutput.t97 a_n5644_8799.t46 vdd.t58 vdd.t51 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X75 output.t14 CSoutput.t123 vdd.t161 gnd.t273 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X76 a_n3827_n3924.t44 diffpairibias.t22 gnd.t313 gnd.t312 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X77 CSoutput.t91 a_n5644_8799.t47 vdd.t57 vdd.t51 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X78 CSoutput.t61 commonsourceibias.t58 gnd.t329 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X79 vdd.t56 a_n5644_8799.t48 CSoutput.t90 vdd.t49 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X80 outputibias.t7 outputibias.t6 gnd.t228 gnd.t227 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X81 a_n1996_n452.t8 a_n1996_n452.t7 a_n1808_13878.t6 vdd.t185 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X82 CSoutput.t60 commonsourceibias.t59 gnd.t28 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X83 gnd.t16 commonsourceibias.t60 CSoutput.t59 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X84 commonsourceibias.t31 commonsourceibias.t30 gnd.t310 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 a_n1996_n452.t22 a_n1996_n452.t21 a_n1808_13878.t5 vdd.t78 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X86 vdd.t55 a_n5644_8799.t49 CSoutput.t89 vdd.t47 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X87 a_n5644_8799.t4 a_n1996_n452.t48 a_n1986_8322.t9 vdd.t178 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X88 gnd.t151 gnd.t149 gnd.t150 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X89 vdd.t54 a_n5644_8799.t50 CSoutput.t111 vdd.t49 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X90 a_n1996_n452.t34 minus.t10 a_n3827_n3924.t17 gnd.t257 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X91 diffpairibias.t15 diffpairibias.t14 gnd.t281 gnd.t280 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X92 outputibias.t5 outputibias.t4 gnd.t243 gnd.t242 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X93 vdd.t141 vdd.t139 vdd.t140 vdd.t93 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X94 a_n3827_n3924.t21 minus.t11 a_n1996_n452.t38 gnd.t263 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X95 vdd.t53 a_n5644_8799.t51 CSoutput.t110 vdd.t38 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X96 vdd.t138 vdd.t136 vdd.t137 vdd.t122 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X97 CSoutput.t58 commonsourceibias.t61 gnd.t249 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X98 gnd.t12 commonsourceibias.t28 commonsourceibias.t29 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X99 vdd.t135 vdd.t132 vdd.t134 vdd.t133 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X100 gnd.t148 gnd.t146 gnd.t147 gnd.t91 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X101 gnd.t49 commonsourceibias.t62 CSoutput.t57 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X102 output.t13 CSoutput.t124 vdd.t159 gnd.t274 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X103 a_n3827_n3924.t47 diffpairibias.t23 gnd.t322 gnd.t321 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X104 vdd.t131 vdd.t128 vdd.t130 vdd.t129 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X105 a_n3827_n3924.t19 minus.t12 a_n1996_n452.t36 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X106 vdd.t158 CSoutput.t125 output.t12 gnd.t275 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X107 vdd.t3 a_n1996_n452.t49 a_n1986_8322.t18 vdd.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X108 vdd.t127 vdd.t125 vdd.t126 vdd.t118 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X109 a_n1996_n452.t37 minus.t13 a_n3827_n3924.t20 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X110 commonsourceibias.t27 commonsourceibias.t26 gnd.t42 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X111 gnd.t241 commonsourceibias.t63 CSoutput.t56 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X112 CSoutput.t109 a_n5644_8799.t52 vdd.t52 vdd.t51 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X113 a_n1986_8322.t17 a_n1996_n452.t50 vdd.t5 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X114 gnd.t142 gnd.t140 gnd.t141 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X115 a_n3827_n3924.t31 plus.t10 a_n5644_8799.t25 gnd.t307 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X116 a_n3827_n3924.t42 plus.t11 a_n5644_8799.t24 gnd.t306 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X117 gnd.t309 commonsourceibias.t24 commonsourceibias.t25 gnd.t254 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X118 gnd.t145 gnd.t143 gnd.t144 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X119 vdd.t50 a_n5644_8799.t53 CSoutput.t101 vdd.t49 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X120 vdd.t167 CSoutput.t126 output.t11 gnd.t268 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X121 vdd.t180 a_n1996_n452.t51 a_n1808_13878.t18 vdd.t179 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X122 a_n5644_8799.t23 plus.t12 a_n3827_n3924.t38 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X123 CSoutput.t55 commonsourceibias.t64 gnd.t223 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X124 a_n5644_8799.t22 plus.t13 a_n3827_n3924.t23 gnd.t305 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X125 gnd.t43 commonsourceibias.t65 CSoutput.t54 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X126 commonsourceibias.t23 commonsourceibias.t22 gnd.t258 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X127 vdd.t124 vdd.t121 vdd.t123 vdd.t122 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X128 a_n1996_n452.t30 minus.t14 a_n3827_n3924.t7 gnd.t187 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X129 diffpairibias.t13 diffpairibias.t12 gnd.t237 gnd.t236 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X130 vdd.t120 vdd.t117 vdd.t119 vdd.t118 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X131 vdd.t48 a_n5644_8799.t54 CSoutput.t100 vdd.t47 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X132 gnd.t139 gnd.t137 minus.t4 gnd.t138 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X133 a_n5644_8799.t1 a_n1996_n452.t52 a_n1986_8322.t8 vdd.t76 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X134 a_n1986_8322.t16 a_n1996_n452.t53 vdd.t193 vdd.t192 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X135 vdd.t116 vdd.t113 vdd.t115 vdd.t114 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X136 a_n3827_n3924.t5 minus.t15 a_n1996_n452.t28 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X137 a_n1996_n452.t18 a_n1996_n452.t17 a_n1808_13878.t4 vdd.t9 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X138 gnd.t292 commonsourceibias.t66 CSoutput.t53 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X139 gnd.t277 commonsourceibias.t67 CSoutput.t52 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X140 a_n5644_8799.t0 a_n1996_n452.t54 a_n1986_8322.t7 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X141 vdd.t162 CSoutput.t127 output.t10 gnd.t269 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X142 a_n1808_13878.t3 a_n1996_n452.t15 a_n1996_n452.t16 vdd.t178 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X143 output.t9 CSoutput.t128 vdd.t171 gnd.t270 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X144 gnd.t136 gnd.t134 gnd.t135 gnd.t99 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X145 CSoutput.t51 commonsourceibias.t68 gnd.t320 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X146 vdd.t187 a_n1996_n452.t55 a_n1986_8322.t15 vdd.t186 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X147 gnd.t133 gnd.t131 minus.t3 gnd.t132 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X148 gnd.t259 commonsourceibias.t69 CSoutput.t50 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X149 a_n3827_n3924.t37 plus.t14 a_n5644_8799.t21 gnd.t287 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X150 output.t8 CSoutput.t129 vdd.t170 gnd.t288 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X151 gnd.t291 commonsourceibias.t70 CSoutput.t49 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X152 vdd.t112 vdd.t110 vdd.t111 vdd.t104 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X153 a_n3827_n3924.t14 diffpairibias.t24 gnd.t235 gnd.t234 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X154 CSoutput.t96 a_n5644_8799.t55 vdd.t46 vdd.t41 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X155 a_n3827_n3924.t49 diffpairibias.t25 gnd.t328 gnd.t327 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X156 vdd.t45 a_n5644_8799.t56 CSoutput.t95 vdd.t12 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X157 gnd.t130 gnd.t128 gnd.t129 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X158 a_n5644_8799.t20 plus.t15 a_n3827_n3924.t34 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X159 vdd.t44 a_n5644_8799.t57 CSoutput.t104 vdd.t27 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X160 CSoutput.t48 commonsourceibias.t71 gnd.t203 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X161 gnd.t127 gnd.t124 gnd.t126 gnd.t125 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X162 gnd.t123 gnd.t121 gnd.t122 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X163 gnd.t256 commonsourceibias.t72 CSoutput.t47 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X164 diffpairibias.t11 diffpairibias.t10 gnd.t46 gnd.t45 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X165 vdd.t169 CSoutput.t130 output.t7 gnd.t289 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X166 gnd.t48 commonsourceibias.t73 CSoutput.t46 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X167 CSoutput.t45 commonsourceibias.t74 gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X168 CSoutput.t103 a_n5644_8799.t58 vdd.t43 vdd.t31 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X169 vdd.t109 vdd.t107 vdd.t108 vdd.t89 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X170 a_n1808_13878.t17 a_n1996_n452.t56 vdd.t199 vdd.t198 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X171 vdd.t197 a_n1996_n452.t57 a_n1808_13878.t16 vdd.t196 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X172 gnd.t296 commonsourceibias.t75 CSoutput.t44 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X173 diffpairibias.t9 diffpairibias.t8 gnd.t20 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X174 a_n3827_n3924.t2 minus.t16 a_n1996_n452.t1 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X175 CSoutput.t131 a_n1986_8322.t22 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X176 vdd.t106 vdd.t103 vdd.t105 vdd.t104 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X177 gnd.t120 gnd.t118 gnd.t119 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X178 commonsourceibias.t21 commonsourceibias.t20 gnd.t10 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X179 a_n1996_n452.t27 minus.t17 a_n3827_n3924.t4 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X180 diffpairibias.t7 diffpairibias.t6 gnd.t219 gnd.t218 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X181 CSoutput.t102 a_n5644_8799.t59 vdd.t42 vdd.t41 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X182 plus.t4 gnd.t115 gnd.t117 gnd.t116 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X183 a_n1996_n452.t33 minus.t18 a_n3827_n3924.t13 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X184 vdd.t40 a_n5644_8799.t60 CSoutput.t106 vdd.t12 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X185 a_n5644_8799.t19 plus.t16 a_n3827_n3924.t30 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X186 CSoutput.t132 a_n1986_8322.t22 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X187 output.t17 outputibias.t10 gnd.t215 gnd.t214 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X188 CSoutput.t43 commonsourceibias.t76 gnd.t27 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X189 a_n1986_8322.t6 a_n1996_n452.t58 a_n5644_8799.t2 vdd.t77 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X190 gnd.t114 gnd.t112 minus.t2 gnd.t113 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X191 a_n3827_n3924.t3 minus.t19 a_n1996_n452.t2 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X192 gnd.t111 gnd.t109 gnd.t110 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X193 commonsourceibias.t19 commonsourceibias.t18 gnd.t301 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X194 vdd.t39 a_n5644_8799.t61 CSoutput.t105 vdd.t38 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X195 CSoutput.t80 a_n5644_8799.t62 vdd.t37 vdd.t18 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X196 gnd.t108 gnd.t105 gnd.t107 gnd.t106 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X197 vdd.t36 a_n5644_8799.t63 CSoutput.t79 vdd.t27 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X198 vdd.t80 a_n1996_n452.t59 a_n1986_8322.t14 vdd.t79 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X199 CSoutput.t42 commonsourceibias.t77 gnd.t311 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X200 output.t16 outputibias.t11 gnd.t225 gnd.t224 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X201 gnd.t317 commonsourceibias.t78 CSoutput.t41 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X202 CSoutput.t40 commonsourceibias.t79 gnd.t199 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X203 output.t6 CSoutput.t133 vdd.t163 gnd.t293 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X204 gnd.t25 commonsourceibias.t16 commonsourceibias.t17 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X205 gnd.t300 commonsourceibias.t80 CSoutput.t39 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X206 a_n1808_13878.t15 a_n1996_n452.t60 vdd.t190 vdd.t189 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X207 minus.t1 gnd.t102 gnd.t104 gnd.t103 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X208 gnd.t101 gnd.t98 gnd.t100 gnd.t99 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X209 CSoutput.t38 commonsourceibias.t81 gnd.t207 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X210 gnd.t308 commonsourceibias.t82 CSoutput.t37 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X211 CSoutput.t36 commonsourceibias.t83 gnd.t252 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 commonsourceibias.t15 commonsourceibias.t14 gnd.t297 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X213 a_n3827_n3924.t0 diffpairibias.t26 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X214 CSoutput.t86 a_n5644_8799.t64 vdd.t35 vdd.t31 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X215 CSoutput.t35 commonsourceibias.t84 gnd.t238 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X216 gnd.t56 commonsourceibias.t85 CSoutput.t34 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X217 CSoutput.t85 a_n5644_8799.t65 vdd.t34 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X218 vdd.t102 vdd.t100 vdd.t101 vdd.t89 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X219 gnd.t44 commonsourceibias.t86 CSoutput.t33 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X220 CSoutput.t32 commonsourceibias.t87 gnd.t299 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X221 a_n5644_8799.t18 plus.t17 a_n3827_n3924.t33 gnd.t304 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X222 a_n1986_8322.t5 a_n1996_n452.t61 a_n5644_8799.t7 vdd.t9 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X223 vdd.t177 a_n1996_n452.t62 a_n1986_8322.t13 vdd.t176 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X224 vdd.t33 a_n5644_8799.t66 CSoutput.t84 vdd.t20 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X225 CSoutput.t114 a_n5644_8799.t67 vdd.t32 vdd.t31 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X226 CSoutput.t31 commonsourceibias.t88 gnd.t55 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X227 gnd.t331 commonsourceibias.t89 CSoutput.t30 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X228 a_n3827_n3924.t39 plus.t18 a_n5644_8799.t17 gnd.t204 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X229 gnd.t97 gnd.t94 gnd.t96 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X230 diffpairibias.t5 diffpairibias.t4 gnd.t324 gnd.t323 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X231 CSoutput.t29 commonsourceibias.t90 gnd.t230 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X232 gnd.t32 commonsourceibias.t91 CSoutput.t28 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X233 vdd.t99 vdd.t96 vdd.t98 vdd.t97 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X234 CSoutput.t27 commonsourceibias.t92 gnd.t276 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 vdd.t95 vdd.t92 vdd.t94 vdd.t93 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X236 a_n1808_13878.t2 a_n1996_n452.t3 a_n1996_n452.t4 vdd.t175 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X237 gnd.t284 commonsourceibias.t93 CSoutput.t26 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X238 vdd.t160 CSoutput.t134 output.t5 gnd.t294 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X239 a_n3827_n3924.t15 diffpairibias.t27 gnd.t245 gnd.t244 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X240 a_n1986_8322.t4 a_n1996_n452.t63 a_n5644_8799.t6 vdd.t173 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X241 gnd.t59 commonsourceibias.t94 CSoutput.t25 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X242 CSoutput.t24 commonsourceibias.t95 gnd.t232 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X243 gnd.t7 commonsourceibias.t12 commonsourceibias.t13 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X244 outputibias.t3 outputibias.t2 gnd.t211 gnd.t210 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X245 gnd.t37 commonsourceibias.t96 CSoutput.t23 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X246 CSoutput.t113 a_n5644_8799.t68 vdd.t30 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X247 a_n1986_8322.t12 a_n1996_n452.t64 vdd.t75 vdd.t74 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X248 CSoutput.t22 commonsourceibias.t97 gnd.t298 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X249 gnd.t255 commonsourceibias.t98 CSoutput.t21 gnd.t254 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X250 CSoutput.t20 commonsourceibias.t99 gnd.t285 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X251 gnd.t34 commonsourceibias.t100 CSoutput.t19 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X252 gnd.t93 gnd.t90 gnd.t92 gnd.t91 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X253 gnd.t286 commonsourceibias.t101 CSoutput.t18 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X254 commonsourceibias.t11 commonsourceibias.t10 gnd.t295 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X255 minus.t0 gnd.t87 gnd.t89 gnd.t88 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X256 gnd.t184 commonsourceibias.t8 commonsourceibias.t9 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X257 vdd.t1 a_n1996_n452.t65 a_n1808_13878.t14 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X258 a_n3827_n3924.t43 minus.t20 a_n1996_n452.t40 gnd.t307 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X259 output.t4 CSoutput.t135 vdd.t157 gnd.t265 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X260 gnd.t86 gnd.t83 gnd.t85 gnd.t84 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X261 gnd.t51 commonsourceibias.t102 CSoutput.t17 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X262 CSoutput.t16 commonsourceibias.t103 gnd.t189 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X263 vdd.t91 vdd.t88 vdd.t90 vdd.t89 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X264 a_n1996_n452.t0 minus.t21 a_n3827_n3924.t1 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X265 a_n1986_8322.t3 a_n1996_n452.t66 a_n5644_8799.t31 vdd.t174 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X266 gnd.t213 commonsourceibias.t6 commonsourceibias.t7 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X267 vdd.t87 vdd.t85 vdd.t86 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X268 a_n5644_8799.t9 a_n1996_n452.t67 a_n1986_8322.t2 vdd.t175 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X269 a_n1808_13878.t13 a_n1996_n452.t68 vdd.t182 vdd.t181 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X270 vdd.t28 a_n5644_8799.t69 CSoutput.t115 vdd.t27 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X271 CSoutput.t72 a_n5644_8799.t70 vdd.t26 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X272 CSoutput.t15 commonsourceibias.t104 gnd.t216 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X273 a_n5644_8799.t16 plus.t19 a_n3827_n3924.t35 gnd.t187 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X274 vdd.t172 CSoutput.t136 output.t3 gnd.t266 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X275 output.t2 CSoutput.t137 vdd.t166 gnd.t267 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X276 a_n3827_n3924.t12 minus.t22 a_n1996_n452.t32 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X277 gnd.t18 commonsourceibias.t105 CSoutput.t14 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 CSoutput.t13 commonsourceibias.t106 gnd.t231 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X279 a_n3827_n3924.t41 plus.t20 a_n5644_8799.t15 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X280 gnd.t253 commonsourceibias.t4 commonsourceibias.t5 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X281 gnd.t282 commonsourceibias.t2 commonsourceibias.t3 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X282 CSoutput.t88 a_n5644_8799.t71 vdd.t24 vdd.t18 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X283 a_n1808_13878.t1 a_n1996_n452.t11 a_n1996_n452.t12 vdd.t76 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X284 gnd.t201 commonsourceibias.t107 CSoutput.t12 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X285 CSoutput.t11 commonsourceibias.t108 gnd.t41 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X286 a_n3827_n3924.t8 diffpairibias.t28 gnd.t191 gnd.t190 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X287 a_n5644_8799.t14 plus.t21 a_n3827_n3924.t32 gnd.t257 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X288 vdd.t168 CSoutput.t138 output.t1 gnd.t271 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X289 CSoutput.t73 a_n5644_8799.t72 vdd.t23 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X290 gnd.t82 gnd.t80 plus.t2 gnd.t81 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X291 gnd.t75 gnd.t72 gnd.t74 gnd.t73 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X292 vdd.t22 a_n5644_8799.t73 CSoutput.t83 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X293 CSoutput.t10 commonsourceibias.t109 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X294 gnd.t183 commonsourceibias.t110 CSoutput.t9 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X295 diffpairibias.t3 diffpairibias.t2 gnd.t315 gnd.t314 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X296 gnd.t79 gnd.t76 gnd.t78 gnd.t77 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X297 a_n5644_8799.t10 a_n1996_n452.t69 a_n1986_8322.t1 vdd.t188 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X298 a_n1996_n452.t6 a_n1996_n452.t5 a_n1808_13878.t0 vdd.t174 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X299 gnd.t71 gnd.t69 plus.t1 gnd.t70 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X300 a_n3827_n3924.t24 plus.t22 a_n5644_8799.t13 gnd.t263 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X301 vdd.t21 a_n5644_8799.t74 CSoutput.t112 vdd.t20 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X302 gnd.t233 commonsourceibias.t111 CSoutput.t8 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X303 vdd.t164 CSoutput.t139 output.t0 gnd.t272 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X304 CSoutput.t140 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X305 gnd.t68 gnd.t65 gnd.t67 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X306 vdd.t84 vdd.t81 vdd.t83 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X307 CSoutput.t7 commonsourceibias.t112 gnd.t212 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X308 diffpairibias.t1 diffpairibias.t0 gnd.t247 gnd.t246 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X309 a_n3827_n3924.t40 plus.t23 a_n5644_8799.t12 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X310 outputibias.t1 outputibias.t0 gnd.t39 gnd.t38 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X311 a_n5644_8799.t11 plus.t24 a_n3827_n3924.t25 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X312 CSoutput.t141 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X313 a_n3827_n3924.t45 minus.t23 a_n1996_n452.t41 gnd.t306 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X314 gnd.t283 commonsourceibias.t113 CSoutput.t6 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X315 gnd.t64 gnd.t61 gnd.t63 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X316 vdd.t8 a_n1996_n452.t70 a_n1808_13878.t12 vdd.t7 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X317 CSoutput.t82 a_n5644_8799.t75 vdd.t19 vdd.t18 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X318 a_n1996_n452.t43 minus.t24 a_n3827_n3924.t48 gnd.t305 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X319 CSoutput.t5 commonsourceibias.t114 gnd.t60 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X320 gnd.t330 commonsourceibias.t115 CSoutput.t4 gnd.t254 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X321 commonsourceibias.t1 commonsourceibias.t0 gnd.t202 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X322 CSoutput.t75 a_n5644_8799.t76 vdd.t17 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X323 CSoutput.t3 commonsourceibias.t116 gnd.t196 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X324 vdd.t15 a_n5644_8799.t77 CSoutput.t87 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X325 a_n1986_8322.t0 a_n1996_n452.t71 a_n5644_8799.t3 vdd.t78 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X326 vdd.t13 a_n5644_8799.t78 CSoutput.t81 vdd.t12 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X327 CSoutput.t74 a_n5644_8799.t79 vdd.t11 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X328 CSoutput.t2 commonsourceibias.t117 gnd.t22 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X329 gnd.t209 commonsourceibias.t118 CSoutput.t1 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 CSoutput.t0 commonsourceibias.t119 gnd.t58 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X331 a_n3827_n3924.t16 diffpairibias.t29 gnd.t251 gnd.t250 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
R0 plus.n43 plus.t18 322.512
R1 plus.n9 plus.t13 322.512
R2 plus.n42 plus.t17 297.12
R3 plus.n46 plus.t22 297.12
R4 plus.n48 plus.t21 297.12
R5 plus.n52 plus.t23 297.12
R6 plus.n54 plus.t8 297.12
R7 plus.n58 plus.t7 297.12
R8 plus.n60 plus.t12 297.12
R9 plus.n64 plus.t10 297.12
R10 plus.n66 plus.t24 297.12
R11 plus.n32 plus.t14 297.12
R12 plus.n30 plus.t15 297.12
R13 plus.n2 plus.t9 297.12
R14 plus.n24 plus.t5 297.12
R15 plus.n4 plus.t6 297.12
R16 plus.n18 plus.t19 297.12
R17 plus.n6 plus.t20 297.12
R18 plus.n12 plus.t16 297.12
R19 plus.n8 plus.t11 297.12
R20 plus.n70 plus.t1 243.97
R21 plus.n70 plus.n69 223.454
R22 plus.n72 plus.n71 223.454
R23 plus.n67 plus.n66 161.3
R24 plus.n65 plus.n34 161.3
R25 plus.n64 plus.n63 161.3
R26 plus.n62 plus.n35 161.3
R27 plus.n61 plus.n60 161.3
R28 plus.n59 plus.n36 161.3
R29 plus.n58 plus.n57 161.3
R30 plus.n56 plus.n37 161.3
R31 plus.n55 plus.n54 161.3
R32 plus.n53 plus.n38 161.3
R33 plus.n52 plus.n51 161.3
R34 plus.n50 plus.n39 161.3
R35 plus.n49 plus.n48 161.3
R36 plus.n47 plus.n40 161.3
R37 plus.n46 plus.n45 161.3
R38 plus.n44 plus.n41 161.3
R39 plus.n11 plus.n10 161.3
R40 plus.n12 plus.n7 161.3
R41 plus.n14 plus.n13 161.3
R42 plus.n15 plus.n6 161.3
R43 plus.n17 plus.n16 161.3
R44 plus.n18 plus.n5 161.3
R45 plus.n20 plus.n19 161.3
R46 plus.n21 plus.n4 161.3
R47 plus.n23 plus.n22 161.3
R48 plus.n24 plus.n3 161.3
R49 plus.n26 plus.n25 161.3
R50 plus.n27 plus.n2 161.3
R51 plus.n29 plus.n28 161.3
R52 plus.n30 plus.n1 161.3
R53 plus.n31 plus.n0 161.3
R54 plus.n33 plus.n32 161.3
R55 plus.n44 plus.n43 45.0031
R56 plus.n10 plus.n9 45.0031
R57 plus.n66 plus.n65 41.6278
R58 plus.n32 plus.n31 41.6278
R59 plus.n42 plus.n41 37.246
R60 plus.n64 plus.n35 37.246
R61 plus.n30 plus.n29 37.246
R62 plus.n11 plus.n8 37.246
R63 plus.n47 plus.n46 32.8641
R64 plus.n60 plus.n59 32.8641
R65 plus.n25 plus.n2 32.8641
R66 plus.n13 plus.n12 32.8641
R67 plus.n68 plus.n67 31.6047
R68 plus.n48 plus.n39 28.4823
R69 plus.n58 plus.n37 28.4823
R70 plus.n24 plus.n23 28.4823
R71 plus.n17 plus.n6 28.4823
R72 plus.n53 plus.n52 24.1005
R73 plus.n54 plus.n53 24.1005
R74 plus.n19 plus.n4 24.1005
R75 plus.n19 plus.n18 24.1005
R76 plus.n69 plus.t3 19.8005
R77 plus.n69 plus.t4 19.8005
R78 plus.n71 plus.t2 19.8005
R79 plus.n71 plus.t0 19.8005
R80 plus.n52 plus.n39 19.7187
R81 plus.n54 plus.n37 19.7187
R82 plus.n23 plus.n4 19.7187
R83 plus.n18 plus.n17 19.7187
R84 plus.n43 plus.n42 15.6319
R85 plus.n9 plus.n8 15.6319
R86 plus.n48 plus.n47 15.3369
R87 plus.n59 plus.n58 15.3369
R88 plus.n25 plus.n24 15.3369
R89 plus.n13 plus.n6 15.3369
R90 plus plus.n73 14.4015
R91 plus.n68 plus.n33 11.866
R92 plus.n46 plus.n41 10.955
R93 plus.n60 plus.n35 10.955
R94 plus.n29 plus.n2 10.955
R95 plus.n12 plus.n11 10.955
R96 plus.n65 plus.n64 6.57323
R97 plus.n31 plus.n30 6.57323
R98 plus.n73 plus.n72 5.40567
R99 plus.n73 plus.n68 1.188
R100 plus.n72 plus.n70 0.716017
R101 plus.n45 plus.n44 0.189894
R102 plus.n45 plus.n40 0.189894
R103 plus.n49 plus.n40 0.189894
R104 plus.n50 plus.n49 0.189894
R105 plus.n51 plus.n50 0.189894
R106 plus.n51 plus.n38 0.189894
R107 plus.n55 plus.n38 0.189894
R108 plus.n56 plus.n55 0.189894
R109 plus.n57 plus.n56 0.189894
R110 plus.n57 plus.n36 0.189894
R111 plus.n61 plus.n36 0.189894
R112 plus.n62 plus.n61 0.189894
R113 plus.n63 plus.n62 0.189894
R114 plus.n63 plus.n34 0.189894
R115 plus.n67 plus.n34 0.189894
R116 plus.n33 plus.n0 0.189894
R117 plus.n1 plus.n0 0.189894
R118 plus.n28 plus.n1 0.189894
R119 plus.n28 plus.n27 0.189894
R120 plus.n27 plus.n26 0.189894
R121 plus.n26 plus.n3 0.189894
R122 plus.n22 plus.n3 0.189894
R123 plus.n22 plus.n21 0.189894
R124 plus.n21 plus.n20 0.189894
R125 plus.n20 plus.n5 0.189894
R126 plus.n16 plus.n5 0.189894
R127 plus.n16 plus.n15 0.189894
R128 plus.n15 plus.n14 0.189894
R129 plus.n14 plus.n7 0.189894
R130 plus.n10 plus.n7 0.189894
R131 a_n3827_n3924.n10 a_n3827_n3924.t15 214.994
R132 a_n3827_n3924.n7 a_n3827_n3924.t9 214.994
R133 a_n3827_n3924.n10 a_n3827_n3924.t47 214.321
R134 a_n3827_n3924.n10 a_n3827_n3924.t8 214.321
R135 a_n3827_n3924.n9 a_n3827_n3924.t49 214.321
R136 a_n3827_n3924.n9 a_n3827_n3924.t16 214.321
R137 a_n3827_n3924.n8 a_n3827_n3924.t14 214.321
R138 a_n3827_n3924.n8 a_n3827_n3924.t10 214.321
R139 a_n3827_n3924.n7 a_n3827_n3924.t44 214.321
R140 a_n3827_n3924.n7 a_n3827_n3924.t0 214.321
R141 a_n3827_n3924.n4 a_n3827_n3924.t39 55.8337
R142 a_n3827_n3924.n4 a_n3827_n3924.t48 55.8337
R143 a_n3827_n3924.n6 a_n3827_n3924.t22 55.8337
R144 a_n3827_n3924.n3 a_n3827_n3924.t25 55.8335
R145 a_n3827_n3924.n11 a_n3827_n3924.t20 55.8335
R146 a_n3827_n3924.n0 a_n3827_n3924.t11 55.8335
R147 a_n3827_n3924.n0 a_n3827_n3924.t23 55.8335
R148 a_n3827_n3924.n2 a_n3827_n3924.t37 55.8335
R149 a_n3827_n3924.n29 a_n3827_n3924.n11 53.0054
R150 a_n3827_n3924.n3 a_n3827_n3924.n13 53.0052
R151 a_n3827_n3924.n4 a_n3827_n3924.n14 53.0052
R152 a_n3827_n3924.n4 a_n3827_n3924.n15 53.0052
R153 a_n3827_n3924.n4 a_n3827_n3924.n16 53.0052
R154 a_n3827_n3924.n5 a_n3827_n3924.n17 53.0052
R155 a_n3827_n3924.n5 a_n3827_n3924.n18 53.0052
R156 a_n3827_n3924.n6 a_n3827_n3924.n19 53.0052
R157 a_n3827_n3924.n6 a_n3827_n3924.n20 53.0052
R158 a_n3827_n3924.n0 a_n3827_n3924.n12 53.0051
R159 a_n3827_n3924.n0 a_n3827_n3924.n21 53.0051
R160 a_n3827_n3924.n0 a_n3827_n3924.n22 53.0051
R161 a_n3827_n3924.n1 a_n3827_n3924.n23 53.0051
R162 a_n3827_n3924.n1 a_n3827_n3924.n24 53.0051
R163 a_n3827_n3924.n2 a_n3827_n3924.n25 53.0051
R164 a_n3827_n3924.n2 a_n3827_n3924.n26 53.0051
R165 a_n3827_n3924.n27 a_n3827_n3924.n6 12.1986
R166 a_n3827_n3924.n28 a_n3827_n3924.n3 12.1986
R167 a_n3827_n3924.n27 a_n3827_n3924.n2 5.11903
R168 a_n3827_n3924.n11 a_n3827_n3924.n28 5.11903
R169 a_n3827_n3924.n12 a_n3827_n3924.t4 2.82907
R170 a_n3827_n3924.n12 a_n3827_n3924.t2 2.82907
R171 a_n3827_n3924.n21 a_n3827_n3924.t17 2.82907
R172 a_n3827_n3924.n21 a_n3827_n3924.t19 2.82907
R173 a_n3827_n3924.n22 a_n3827_n3924.t46 2.82907
R174 a_n3827_n3924.n22 a_n3827_n3924.t21 2.82907
R175 a_n3827_n3924.n23 a_n3827_n3924.t30 2.82907
R176 a_n3827_n3924.n23 a_n3827_n3924.t42 2.82907
R177 a_n3827_n3924.n24 a_n3827_n3924.t35 2.82907
R178 a_n3827_n3924.n24 a_n3827_n3924.t41 2.82907
R179 a_n3827_n3924.n25 a_n3827_n3924.t26 2.82907
R180 a_n3827_n3924.n25 a_n3827_n3924.t36 2.82907
R181 a_n3827_n3924.n26 a_n3827_n3924.t34 2.82907
R182 a_n3827_n3924.n26 a_n3827_n3924.t27 2.82907
R183 a_n3827_n3924.n13 a_n3827_n3924.t38 2.82907
R184 a_n3827_n3924.n13 a_n3827_n3924.t31 2.82907
R185 a_n3827_n3924.n14 a_n3827_n3924.t29 2.82907
R186 a_n3827_n3924.n14 a_n3827_n3924.t28 2.82907
R187 a_n3827_n3924.n15 a_n3827_n3924.t32 2.82907
R188 a_n3827_n3924.n15 a_n3827_n3924.t40 2.82907
R189 a_n3827_n3924.n16 a_n3827_n3924.t33 2.82907
R190 a_n3827_n3924.n16 a_n3827_n3924.t24 2.82907
R191 a_n3827_n3924.n17 a_n3827_n3924.t6 2.82907
R192 a_n3827_n3924.n17 a_n3827_n3924.t45 2.82907
R193 a_n3827_n3924.n18 a_n3827_n3924.t7 2.82907
R194 a_n3827_n3924.n18 a_n3827_n3924.t5 2.82907
R195 a_n3827_n3924.n19 a_n3827_n3924.t13 2.82907
R196 a_n3827_n3924.n19 a_n3827_n3924.t3 2.82907
R197 a_n3827_n3924.n20 a_n3827_n3924.t18 2.82907
R198 a_n3827_n3924.n20 a_n3827_n3924.t12 2.82907
R199 a_n3827_n3924.t1 a_n3827_n3924.n29 2.82907
R200 a_n3827_n3924.n29 a_n3827_n3924.t43 2.82907
R201 a_n3827_n3924.n8 a_n3827_n3924.n7 2.01503
R202 a_n3827_n3924.n7 a_n3827_n3924.n27 1.95694
R203 a_n3827_n3924.n28 a_n3827_n3924.n10 1.95694
R204 a_n3827_n3924.n6 a_n3827_n3924.n5 1.77636
R205 a_n3827_n3924.n4 a_n3827_n3924.n3 1.77636
R206 a_n3827_n3924.n2 a_n3827_n3924.n1 1.77636
R207 a_n3827_n3924.n11 a_n3827_n3924.n0 1.77636
R208 a_n3827_n3924.n9 a_n3827_n3924.n8 1.34352
R209 a_n3827_n3924.n10 a_n3827_n3924.n9 1.34352
R210 a_n3827_n3924.n1 a_n3827_n3924.n0 1.12334
R211 a_n3827_n3924.n5 a_n3827_n3924.n4 1.12334
R212 a_n5644_8799.n85 a_n5644_8799.t65 485.149
R213 a_n5644_8799.n107 a_n5644_8799.t68 485.149
R214 a_n5644_8799.n130 a_n5644_8799.t34 485.149
R215 a_n5644_8799.n17 a_n5644_8799.t49 485.149
R216 a_n5644_8799.n39 a_n5644_8799.t54 485.149
R217 a_n5644_8799.n62 a_n5644_8799.t35 485.149
R218 a_n5644_8799.n100 a_n5644_8799.t56 464.166
R219 a_n5644_8799.n99 a_n5644_8799.t55 464.166
R220 a_n5644_8799.n81 a_n5644_8799.t42 464.166
R221 a_n5644_8799.n93 a_n5644_8799.t72 464.166
R222 a_n5644_8799.n92 a_n5644_8799.t57 464.166
R223 a_n5644_8799.n84 a_n5644_8799.t47 464.166
R224 a_n5644_8799.n86 a_n5644_8799.t74 464.166
R225 a_n5644_8799.n122 a_n5644_8799.t60 464.166
R226 a_n5644_8799.n121 a_n5644_8799.t59 464.166
R227 a_n5644_8799.n103 a_n5644_8799.t51 464.166
R228 a_n5644_8799.n115 a_n5644_8799.t76 464.166
R229 a_n5644_8799.n114 a_n5644_8799.t63 464.166
R230 a_n5644_8799.n106 a_n5644_8799.t52 464.166
R231 a_n5644_8799.n108 a_n5644_8799.t32 464.166
R232 a_n5644_8799.n145 a_n5644_8799.t78 464.166
R233 a_n5644_8799.n144 a_n5644_8799.t40 464.166
R234 a_n5644_8799.n126 a_n5644_8799.t61 464.166
R235 a_n5644_8799.n138 a_n5644_8799.t33 464.166
R236 a_n5644_8799.n137 a_n5644_8799.t69 464.166
R237 a_n5644_8799.n129 a_n5644_8799.t46 464.166
R238 a_n5644_8799.n131 a_n5644_8799.t66 464.166
R239 a_n5644_8799.n18 a_n5644_8799.t58 464.166
R240 a_n5644_8799.n20 a_n5644_8799.t73 464.166
R241 a_n5644_8799.n24 a_n5644_8799.t38 464.166
R242 a_n5644_8799.n25 a_n5644_8799.t48 464.166
R243 a_n5644_8799.n13 a_n5644_8799.t71 464.166
R244 a_n5644_8799.n31 a_n5644_8799.t37 464.166
R245 a_n5644_8799.n32 a_n5644_8799.t36 464.166
R246 a_n5644_8799.n40 a_n5644_8799.t64 464.166
R247 a_n5644_8799.n42 a_n5644_8799.t77 464.166
R248 a_n5644_8799.n46 a_n5644_8799.t45 464.166
R249 a_n5644_8799.n47 a_n5644_8799.t53 464.166
R250 a_n5644_8799.n35 a_n5644_8799.t75 464.166
R251 a_n5644_8799.n53 a_n5644_8799.t41 464.166
R252 a_n5644_8799.n54 a_n5644_8799.t43 464.166
R253 a_n5644_8799.n63 a_n5644_8799.t67 464.166
R254 a_n5644_8799.n65 a_n5644_8799.t44 464.166
R255 a_n5644_8799.n69 a_n5644_8799.t70 464.166
R256 a_n5644_8799.n70 a_n5644_8799.t50 464.166
R257 a_n5644_8799.n58 a_n5644_8799.t62 464.166
R258 a_n5644_8799.n76 a_n5644_8799.t39 464.166
R259 a_n5644_8799.n77 a_n5644_8799.t79 464.166
R260 a_n5644_8799.n88 a_n5644_8799.n87 161.3
R261 a_n5644_8799.n89 a_n5644_8799.n84 161.3
R262 a_n5644_8799.n91 a_n5644_8799.n90 161.3
R263 a_n5644_8799.n92 a_n5644_8799.n83 161.3
R264 a_n5644_8799.n93 a_n5644_8799.n82 161.3
R265 a_n5644_8799.n95 a_n5644_8799.n94 161.3
R266 a_n5644_8799.n96 a_n5644_8799.n81 161.3
R267 a_n5644_8799.n98 a_n5644_8799.n97 161.3
R268 a_n5644_8799.n99 a_n5644_8799.n80 161.3
R269 a_n5644_8799.n101 a_n5644_8799.n100 161.3
R270 a_n5644_8799.n110 a_n5644_8799.n109 161.3
R271 a_n5644_8799.n111 a_n5644_8799.n106 161.3
R272 a_n5644_8799.n113 a_n5644_8799.n112 161.3
R273 a_n5644_8799.n114 a_n5644_8799.n105 161.3
R274 a_n5644_8799.n115 a_n5644_8799.n104 161.3
R275 a_n5644_8799.n117 a_n5644_8799.n116 161.3
R276 a_n5644_8799.n118 a_n5644_8799.n103 161.3
R277 a_n5644_8799.n120 a_n5644_8799.n119 161.3
R278 a_n5644_8799.n121 a_n5644_8799.n102 161.3
R279 a_n5644_8799.n123 a_n5644_8799.n122 161.3
R280 a_n5644_8799.n133 a_n5644_8799.n132 161.3
R281 a_n5644_8799.n134 a_n5644_8799.n129 161.3
R282 a_n5644_8799.n136 a_n5644_8799.n135 161.3
R283 a_n5644_8799.n137 a_n5644_8799.n128 161.3
R284 a_n5644_8799.n138 a_n5644_8799.n127 161.3
R285 a_n5644_8799.n140 a_n5644_8799.n139 161.3
R286 a_n5644_8799.n141 a_n5644_8799.n126 161.3
R287 a_n5644_8799.n143 a_n5644_8799.n142 161.3
R288 a_n5644_8799.n144 a_n5644_8799.n125 161.3
R289 a_n5644_8799.n146 a_n5644_8799.n145 161.3
R290 a_n5644_8799.n33 a_n5644_8799.n32 161.3
R291 a_n5644_8799.n31 a_n5644_8799.n12 161.3
R292 a_n5644_8799.n30 a_n5644_8799.n29 161.3
R293 a_n5644_8799.n28 a_n5644_8799.n13 161.3
R294 a_n5644_8799.n27 a_n5644_8799.n26 161.3
R295 a_n5644_8799.n25 a_n5644_8799.n14 161.3
R296 a_n5644_8799.n24 a_n5644_8799.n23 161.3
R297 a_n5644_8799.n22 a_n5644_8799.n15 161.3
R298 a_n5644_8799.n21 a_n5644_8799.n20 161.3
R299 a_n5644_8799.n19 a_n5644_8799.n16 161.3
R300 a_n5644_8799.n55 a_n5644_8799.n54 161.3
R301 a_n5644_8799.n53 a_n5644_8799.n34 161.3
R302 a_n5644_8799.n52 a_n5644_8799.n51 161.3
R303 a_n5644_8799.n50 a_n5644_8799.n35 161.3
R304 a_n5644_8799.n49 a_n5644_8799.n48 161.3
R305 a_n5644_8799.n47 a_n5644_8799.n36 161.3
R306 a_n5644_8799.n46 a_n5644_8799.n45 161.3
R307 a_n5644_8799.n44 a_n5644_8799.n37 161.3
R308 a_n5644_8799.n43 a_n5644_8799.n42 161.3
R309 a_n5644_8799.n41 a_n5644_8799.n38 161.3
R310 a_n5644_8799.n78 a_n5644_8799.n77 161.3
R311 a_n5644_8799.n76 a_n5644_8799.n57 161.3
R312 a_n5644_8799.n75 a_n5644_8799.n74 161.3
R313 a_n5644_8799.n73 a_n5644_8799.n58 161.3
R314 a_n5644_8799.n72 a_n5644_8799.n71 161.3
R315 a_n5644_8799.n70 a_n5644_8799.n59 161.3
R316 a_n5644_8799.n69 a_n5644_8799.n68 161.3
R317 a_n5644_8799.n67 a_n5644_8799.n60 161.3
R318 a_n5644_8799.n66 a_n5644_8799.n65 161.3
R319 a_n5644_8799.n64 a_n5644_8799.n61 161.3
R320 a_n5644_8799.n8 a_n5644_8799.n6 98.9633
R321 a_n5644_8799.n3 a_n5644_8799.n1 98.9631
R322 a_n5644_8799.n10 a_n5644_8799.n9 98.6055
R323 a_n5644_8799.n8 a_n5644_8799.n7 98.6055
R324 a_n5644_8799.n3 a_n5644_8799.n2 98.6055
R325 a_n5644_8799.n5 a_n5644_8799.n4 98.6055
R326 a_n5644_8799.n152 a_n5644_8799.n150 81.3764
R327 a_n5644_8799.n161 a_n5644_8799.n159 81.3764
R328 a_n5644_8799.n164 a_n5644_8799.n0 81.3764
R329 a_n5644_8799.n165 a_n5644_8799.n164 80.9326
R330 a_n5644_8799.n158 a_n5644_8799.n157 80.9324
R331 a_n5644_8799.n156 a_n5644_8799.n155 80.9324
R332 a_n5644_8799.n154 a_n5644_8799.n153 80.9324
R333 a_n5644_8799.n152 a_n5644_8799.n151 80.9324
R334 a_n5644_8799.n161 a_n5644_8799.n160 80.9324
R335 a_n5644_8799.n163 a_n5644_8799.n162 80.9324
R336 a_n5644_8799.n88 a_n5644_8799.n85 70.4033
R337 a_n5644_8799.n110 a_n5644_8799.n107 70.4033
R338 a_n5644_8799.n133 a_n5644_8799.n130 70.4033
R339 a_n5644_8799.n17 a_n5644_8799.n16 70.4033
R340 a_n5644_8799.n39 a_n5644_8799.n38 70.4033
R341 a_n5644_8799.n62 a_n5644_8799.n61 70.4033
R342 a_n5644_8799.n100 a_n5644_8799.n99 48.2005
R343 a_n5644_8799.n93 a_n5644_8799.n92 48.2005
R344 a_n5644_8799.n122 a_n5644_8799.n121 48.2005
R345 a_n5644_8799.n115 a_n5644_8799.n114 48.2005
R346 a_n5644_8799.n145 a_n5644_8799.n144 48.2005
R347 a_n5644_8799.n138 a_n5644_8799.n137 48.2005
R348 a_n5644_8799.n25 a_n5644_8799.n24 48.2005
R349 a_n5644_8799.n32 a_n5644_8799.n31 48.2005
R350 a_n5644_8799.n47 a_n5644_8799.n46 48.2005
R351 a_n5644_8799.n54 a_n5644_8799.n53 48.2005
R352 a_n5644_8799.n70 a_n5644_8799.n69 48.2005
R353 a_n5644_8799.n77 a_n5644_8799.n76 48.2005
R354 a_n5644_8799.n98 a_n5644_8799.n81 37.246
R355 a_n5644_8799.n87 a_n5644_8799.n84 37.246
R356 a_n5644_8799.n120 a_n5644_8799.n103 37.246
R357 a_n5644_8799.n109 a_n5644_8799.n106 37.246
R358 a_n5644_8799.n143 a_n5644_8799.n126 37.246
R359 a_n5644_8799.n132 a_n5644_8799.n129 37.246
R360 a_n5644_8799.n20 a_n5644_8799.n19 37.246
R361 a_n5644_8799.n30 a_n5644_8799.n13 37.246
R362 a_n5644_8799.n42 a_n5644_8799.n41 37.246
R363 a_n5644_8799.n52 a_n5644_8799.n35 37.246
R364 a_n5644_8799.n65 a_n5644_8799.n64 37.246
R365 a_n5644_8799.n75 a_n5644_8799.n58 37.246
R366 a_n5644_8799.n94 a_n5644_8799.n81 35.7853
R367 a_n5644_8799.n91 a_n5644_8799.n84 35.7853
R368 a_n5644_8799.n116 a_n5644_8799.n103 35.7853
R369 a_n5644_8799.n113 a_n5644_8799.n106 35.7853
R370 a_n5644_8799.n139 a_n5644_8799.n126 35.7853
R371 a_n5644_8799.n136 a_n5644_8799.n129 35.7853
R372 a_n5644_8799.n20 a_n5644_8799.n15 35.7853
R373 a_n5644_8799.n26 a_n5644_8799.n13 35.7853
R374 a_n5644_8799.n42 a_n5644_8799.n37 35.7853
R375 a_n5644_8799.n48 a_n5644_8799.n35 35.7853
R376 a_n5644_8799.n65 a_n5644_8799.n60 35.7853
R377 a_n5644_8799.n71 a_n5644_8799.n58 35.7853
R378 a_n5644_8799.n163 a_n5644_8799.n158 32.7526
R379 a_n5644_8799.n11 a_n5644_8799.n5 30.7135
R380 a_n5644_8799.n86 a_n5644_8799.n85 20.9576
R381 a_n5644_8799.n108 a_n5644_8799.n107 20.9576
R382 a_n5644_8799.n131 a_n5644_8799.n130 20.9576
R383 a_n5644_8799.n18 a_n5644_8799.n17 20.9576
R384 a_n5644_8799.n40 a_n5644_8799.n39 20.9576
R385 a_n5644_8799.n63 a_n5644_8799.n62 20.9576
R386 a_n5644_8799.n11 a_n5644_8799.n10 17.7361
R387 a_n5644_8799.n94 a_n5644_8799.n93 12.4157
R388 a_n5644_8799.n92 a_n5644_8799.n91 12.4157
R389 a_n5644_8799.n116 a_n5644_8799.n115 12.4157
R390 a_n5644_8799.n114 a_n5644_8799.n113 12.4157
R391 a_n5644_8799.n139 a_n5644_8799.n138 12.4157
R392 a_n5644_8799.n137 a_n5644_8799.n136 12.4157
R393 a_n5644_8799.n24 a_n5644_8799.n15 12.4157
R394 a_n5644_8799.n26 a_n5644_8799.n25 12.4157
R395 a_n5644_8799.n46 a_n5644_8799.n37 12.4157
R396 a_n5644_8799.n48 a_n5644_8799.n47 12.4157
R397 a_n5644_8799.n69 a_n5644_8799.n60 12.4157
R398 a_n5644_8799.n71 a_n5644_8799.n70 12.4157
R399 a_n5644_8799.n154 a_n5644_8799.n149 12.3339
R400 a_n5644_8799.n149 a_n5644_8799.n11 11.4887
R401 a_n5644_8799.n99 a_n5644_8799.n98 10.955
R402 a_n5644_8799.n87 a_n5644_8799.n86 10.955
R403 a_n5644_8799.n121 a_n5644_8799.n120 10.955
R404 a_n5644_8799.n109 a_n5644_8799.n108 10.955
R405 a_n5644_8799.n144 a_n5644_8799.n143 10.955
R406 a_n5644_8799.n132 a_n5644_8799.n131 10.955
R407 a_n5644_8799.n19 a_n5644_8799.n18 10.955
R408 a_n5644_8799.n31 a_n5644_8799.n30 10.955
R409 a_n5644_8799.n41 a_n5644_8799.n40 10.955
R410 a_n5644_8799.n53 a_n5644_8799.n52 10.955
R411 a_n5644_8799.n64 a_n5644_8799.n63 10.955
R412 a_n5644_8799.n76 a_n5644_8799.n75 10.955
R413 a_n5644_8799.n124 a_n5644_8799.n101 9.05164
R414 a_n5644_8799.n56 a_n5644_8799.n33 9.05164
R415 a_n5644_8799.n148 a_n5644_8799.n79 6.86985
R416 a_n5644_8799.n148 a_n5644_8799.n147 6.51296
R417 a_n5644_8799.n124 a_n5644_8799.n123 4.94368
R418 a_n5644_8799.n147 a_n5644_8799.n146 4.94368
R419 a_n5644_8799.n56 a_n5644_8799.n55 4.94368
R420 a_n5644_8799.n79 a_n5644_8799.n78 4.94368
R421 a_n5644_8799.n147 a_n5644_8799.n124 4.10845
R422 a_n5644_8799.n79 a_n5644_8799.n56 4.10845
R423 a_n5644_8799.n9 a_n5644_8799.t6 3.61217
R424 a_n5644_8799.n9 a_n5644_8799.t10 3.61217
R425 a_n5644_8799.n7 a_n5644_8799.t2 3.61217
R426 a_n5644_8799.n7 a_n5644_8799.t4 3.61217
R427 a_n5644_8799.n6 a_n5644_8799.t3 3.61217
R428 a_n5644_8799.n6 a_n5644_8799.t0 3.61217
R429 a_n5644_8799.n1 a_n5644_8799.t7 3.61217
R430 a_n5644_8799.n1 a_n5644_8799.t8 3.61217
R431 a_n5644_8799.n2 a_n5644_8799.t5 3.61217
R432 a_n5644_8799.n2 a_n5644_8799.t1 3.61217
R433 a_n5644_8799.n4 a_n5644_8799.t31 3.61217
R434 a_n5644_8799.n4 a_n5644_8799.t9 3.61217
R435 a_n5644_8799.n149 a_n5644_8799.n148 3.4105
R436 a_n5644_8799.n159 a_n5644_8799.t24 2.82907
R437 a_n5644_8799.n159 a_n5644_8799.t22 2.82907
R438 a_n5644_8799.n160 a_n5644_8799.t15 2.82907
R439 a_n5644_8799.n160 a_n5644_8799.t19 2.82907
R440 a_n5644_8799.n162 a_n5644_8799.t29 2.82907
R441 a_n5644_8799.n162 a_n5644_8799.t16 2.82907
R442 a_n5644_8799.n157 a_n5644_8799.t25 2.82907
R443 a_n5644_8799.n157 a_n5644_8799.t11 2.82907
R444 a_n5644_8799.n155 a_n5644_8799.t28 2.82907
R445 a_n5644_8799.n155 a_n5644_8799.t23 2.82907
R446 a_n5644_8799.n153 a_n5644_8799.t12 2.82907
R447 a_n5644_8799.n153 a_n5644_8799.t27 2.82907
R448 a_n5644_8799.n151 a_n5644_8799.t13 2.82907
R449 a_n5644_8799.n151 a_n5644_8799.t14 2.82907
R450 a_n5644_8799.n150 a_n5644_8799.t17 2.82907
R451 a_n5644_8799.n150 a_n5644_8799.t18 2.82907
R452 a_n5644_8799.n0 a_n5644_8799.t21 2.82907
R453 a_n5644_8799.n0 a_n5644_8799.t20 2.82907
R454 a_n5644_8799.n165 a_n5644_8799.t26 2.82907
R455 a_n5644_8799.t30 a_n5644_8799.n165 2.82907
R456 a_n5644_8799.n154 a_n5644_8799.n152 0.444466
R457 a_n5644_8799.n156 a_n5644_8799.n154 0.444466
R458 a_n5644_8799.n158 a_n5644_8799.n156 0.444466
R459 a_n5644_8799.n164 a_n5644_8799.n163 0.444466
R460 a_n5644_8799.n163 a_n5644_8799.n161 0.444466
R461 a_n5644_8799.n10 a_n5644_8799.n8 0.358259
R462 a_n5644_8799.n5 a_n5644_8799.n3 0.358259
R463 a_n5644_8799.n101 a_n5644_8799.n80 0.189894
R464 a_n5644_8799.n97 a_n5644_8799.n80 0.189894
R465 a_n5644_8799.n97 a_n5644_8799.n96 0.189894
R466 a_n5644_8799.n96 a_n5644_8799.n95 0.189894
R467 a_n5644_8799.n95 a_n5644_8799.n82 0.189894
R468 a_n5644_8799.n83 a_n5644_8799.n82 0.189894
R469 a_n5644_8799.n90 a_n5644_8799.n83 0.189894
R470 a_n5644_8799.n90 a_n5644_8799.n89 0.189894
R471 a_n5644_8799.n89 a_n5644_8799.n88 0.189894
R472 a_n5644_8799.n123 a_n5644_8799.n102 0.189894
R473 a_n5644_8799.n119 a_n5644_8799.n102 0.189894
R474 a_n5644_8799.n119 a_n5644_8799.n118 0.189894
R475 a_n5644_8799.n118 a_n5644_8799.n117 0.189894
R476 a_n5644_8799.n117 a_n5644_8799.n104 0.189894
R477 a_n5644_8799.n105 a_n5644_8799.n104 0.189894
R478 a_n5644_8799.n112 a_n5644_8799.n105 0.189894
R479 a_n5644_8799.n112 a_n5644_8799.n111 0.189894
R480 a_n5644_8799.n111 a_n5644_8799.n110 0.189894
R481 a_n5644_8799.n146 a_n5644_8799.n125 0.189894
R482 a_n5644_8799.n142 a_n5644_8799.n125 0.189894
R483 a_n5644_8799.n142 a_n5644_8799.n141 0.189894
R484 a_n5644_8799.n141 a_n5644_8799.n140 0.189894
R485 a_n5644_8799.n140 a_n5644_8799.n127 0.189894
R486 a_n5644_8799.n128 a_n5644_8799.n127 0.189894
R487 a_n5644_8799.n135 a_n5644_8799.n128 0.189894
R488 a_n5644_8799.n135 a_n5644_8799.n134 0.189894
R489 a_n5644_8799.n134 a_n5644_8799.n133 0.189894
R490 a_n5644_8799.n21 a_n5644_8799.n16 0.189894
R491 a_n5644_8799.n22 a_n5644_8799.n21 0.189894
R492 a_n5644_8799.n23 a_n5644_8799.n22 0.189894
R493 a_n5644_8799.n23 a_n5644_8799.n14 0.189894
R494 a_n5644_8799.n27 a_n5644_8799.n14 0.189894
R495 a_n5644_8799.n28 a_n5644_8799.n27 0.189894
R496 a_n5644_8799.n29 a_n5644_8799.n28 0.189894
R497 a_n5644_8799.n29 a_n5644_8799.n12 0.189894
R498 a_n5644_8799.n33 a_n5644_8799.n12 0.189894
R499 a_n5644_8799.n43 a_n5644_8799.n38 0.189894
R500 a_n5644_8799.n44 a_n5644_8799.n43 0.189894
R501 a_n5644_8799.n45 a_n5644_8799.n44 0.189894
R502 a_n5644_8799.n45 a_n5644_8799.n36 0.189894
R503 a_n5644_8799.n49 a_n5644_8799.n36 0.189894
R504 a_n5644_8799.n50 a_n5644_8799.n49 0.189894
R505 a_n5644_8799.n51 a_n5644_8799.n50 0.189894
R506 a_n5644_8799.n51 a_n5644_8799.n34 0.189894
R507 a_n5644_8799.n55 a_n5644_8799.n34 0.189894
R508 a_n5644_8799.n66 a_n5644_8799.n61 0.189894
R509 a_n5644_8799.n67 a_n5644_8799.n66 0.189894
R510 a_n5644_8799.n68 a_n5644_8799.n67 0.189894
R511 a_n5644_8799.n68 a_n5644_8799.n59 0.189894
R512 a_n5644_8799.n72 a_n5644_8799.n59 0.189894
R513 a_n5644_8799.n73 a_n5644_8799.n72 0.189894
R514 a_n5644_8799.n74 a_n5644_8799.n73 0.189894
R515 a_n5644_8799.n74 a_n5644_8799.n57 0.189894
R516 a_n5644_8799.n78 a_n5644_8799.n57 0.189894
R517 gnd.n5620 gnd.n4173 939.716
R518 gnd.n6110 gnd.n643 893.337
R519 gnd.n6740 gnd.n165 838.452
R520 gnd.n6851 gnd.n6750 838.452
R521 gnd.n322 gnd.n273 838.452
R522 gnd.n6344 gnd.n502 838.452
R523 gnd.n1340 gnd.n1329 838.452
R524 gnd.n2569 gnd.n2568 838.452
R525 gnd.n2365 gnd.n1060 838.452
R526 gnd.n4051 gnd.n1133 838.452
R527 gnd.n7057 gnd.n161 783.196
R528 gnd.n7061 gnd.n7060 783.196
R529 gnd.n501 gnd.n500 783.196
R530 gnd.n6548 gnd.n277 783.196
R531 gnd.n3920 gnd.n1333 783.196
R532 gnd.n2248 gnd.n2247 783.196
R533 gnd.n1136 gnd.n1135 783.196
R534 gnd.n4171 gnd.n1064 783.196
R535 gnd.n5528 gnd.n1009 766.379
R536 gnd.n5531 gnd.n5530 766.379
R537 gnd.n4770 gnd.n4673 766.379
R538 gnd.n4766 gnd.n4671 766.379
R539 gnd.n5619 gnd.n4182 756.769
R540 gnd.n5522 gnd.n5521 756.769
R541 gnd.n4863 gnd.n4580 756.769
R542 gnd.n4861 gnd.n4583 756.769
R543 gnd.n2634 gnd.n2079 711.122
R544 gnd.n6370 gnd.n460 711.122
R545 gnd.n2636 gnd.n2076 711.122
R546 gnd.n6372 gnd.n456 711.122
R547 gnd.n5791 gnd.n839 655.866
R548 gnd.n6111 gnd.n644 655.866
R549 gnd.n6325 gnd.n517 655.866
R550 gnd.n2518 gnd.n1007 655.866
R551 gnd.n842 gnd.n839 585
R552 gnd.n5789 gnd.n839 585
R553 gnd.n5787 gnd.n5786 585
R554 gnd.n5788 gnd.n5787 585
R555 gnd.n5785 gnd.n841 585
R556 gnd.n841 gnd.n840 585
R557 gnd.n5784 gnd.n5783 585
R558 gnd.n5783 gnd.n5782 585
R559 gnd.n847 gnd.n846 585
R560 gnd.n5781 gnd.n847 585
R561 gnd.n5779 gnd.n5778 585
R562 gnd.n5780 gnd.n5779 585
R563 gnd.n5777 gnd.n849 585
R564 gnd.n849 gnd.n848 585
R565 gnd.n5776 gnd.n5775 585
R566 gnd.n5775 gnd.n5774 585
R567 gnd.n855 gnd.n854 585
R568 gnd.n5773 gnd.n855 585
R569 gnd.n5771 gnd.n5770 585
R570 gnd.n5772 gnd.n5771 585
R571 gnd.n5769 gnd.n857 585
R572 gnd.n857 gnd.n856 585
R573 gnd.n5768 gnd.n5767 585
R574 gnd.n5767 gnd.n5766 585
R575 gnd.n863 gnd.n862 585
R576 gnd.n5765 gnd.n863 585
R577 gnd.n5763 gnd.n5762 585
R578 gnd.n5764 gnd.n5763 585
R579 gnd.n5761 gnd.n865 585
R580 gnd.n865 gnd.n864 585
R581 gnd.n5760 gnd.n5759 585
R582 gnd.n5759 gnd.n5758 585
R583 gnd.n871 gnd.n870 585
R584 gnd.n5757 gnd.n871 585
R585 gnd.n5755 gnd.n5754 585
R586 gnd.n5756 gnd.n5755 585
R587 gnd.n5753 gnd.n873 585
R588 gnd.n873 gnd.n872 585
R589 gnd.n5752 gnd.n5751 585
R590 gnd.n5751 gnd.n5750 585
R591 gnd.n879 gnd.n878 585
R592 gnd.n5749 gnd.n879 585
R593 gnd.n5747 gnd.n5746 585
R594 gnd.n5748 gnd.n5747 585
R595 gnd.n5745 gnd.n881 585
R596 gnd.n881 gnd.n880 585
R597 gnd.n5744 gnd.n5743 585
R598 gnd.n5743 gnd.n5742 585
R599 gnd.n887 gnd.n886 585
R600 gnd.n5741 gnd.n887 585
R601 gnd.n5739 gnd.n5738 585
R602 gnd.n5740 gnd.n5739 585
R603 gnd.n5737 gnd.n889 585
R604 gnd.n889 gnd.n888 585
R605 gnd.n5736 gnd.n5735 585
R606 gnd.n5735 gnd.n5734 585
R607 gnd.n895 gnd.n894 585
R608 gnd.n5733 gnd.n895 585
R609 gnd.n5731 gnd.n5730 585
R610 gnd.n5732 gnd.n5731 585
R611 gnd.n5729 gnd.n897 585
R612 gnd.n897 gnd.n896 585
R613 gnd.n5728 gnd.n5727 585
R614 gnd.n5727 gnd.n5726 585
R615 gnd.n903 gnd.n902 585
R616 gnd.n5725 gnd.n903 585
R617 gnd.n5723 gnd.n5722 585
R618 gnd.n5724 gnd.n5723 585
R619 gnd.n5721 gnd.n905 585
R620 gnd.n905 gnd.n904 585
R621 gnd.n5720 gnd.n5719 585
R622 gnd.n5719 gnd.n5718 585
R623 gnd.n911 gnd.n910 585
R624 gnd.n5717 gnd.n911 585
R625 gnd.n5715 gnd.n5714 585
R626 gnd.n5716 gnd.n5715 585
R627 gnd.n5713 gnd.n913 585
R628 gnd.n913 gnd.n912 585
R629 gnd.n5712 gnd.n5711 585
R630 gnd.n5711 gnd.n5710 585
R631 gnd.n919 gnd.n918 585
R632 gnd.n5709 gnd.n919 585
R633 gnd.n5707 gnd.n5706 585
R634 gnd.n5708 gnd.n5707 585
R635 gnd.n5705 gnd.n921 585
R636 gnd.n921 gnd.n920 585
R637 gnd.n5704 gnd.n5703 585
R638 gnd.n5703 gnd.n5702 585
R639 gnd.n927 gnd.n926 585
R640 gnd.n5701 gnd.n927 585
R641 gnd.n5699 gnd.n5698 585
R642 gnd.n5700 gnd.n5699 585
R643 gnd.n5697 gnd.n929 585
R644 gnd.n929 gnd.n928 585
R645 gnd.n5696 gnd.n5695 585
R646 gnd.n5695 gnd.n5694 585
R647 gnd.n935 gnd.n934 585
R648 gnd.n5693 gnd.n935 585
R649 gnd.n5691 gnd.n5690 585
R650 gnd.n5692 gnd.n5691 585
R651 gnd.n5689 gnd.n937 585
R652 gnd.n937 gnd.n936 585
R653 gnd.n5688 gnd.n5687 585
R654 gnd.n5687 gnd.n5686 585
R655 gnd.n943 gnd.n942 585
R656 gnd.n5685 gnd.n943 585
R657 gnd.n5683 gnd.n5682 585
R658 gnd.n5684 gnd.n5683 585
R659 gnd.n5681 gnd.n945 585
R660 gnd.n945 gnd.n944 585
R661 gnd.n5680 gnd.n5679 585
R662 gnd.n5679 gnd.n5678 585
R663 gnd.n951 gnd.n950 585
R664 gnd.n5677 gnd.n951 585
R665 gnd.n5675 gnd.n5674 585
R666 gnd.n5676 gnd.n5675 585
R667 gnd.n5673 gnd.n953 585
R668 gnd.n953 gnd.n952 585
R669 gnd.n5672 gnd.n5671 585
R670 gnd.n5671 gnd.n5670 585
R671 gnd.n959 gnd.n958 585
R672 gnd.n5669 gnd.n959 585
R673 gnd.n5667 gnd.n5666 585
R674 gnd.n5668 gnd.n5667 585
R675 gnd.n5665 gnd.n961 585
R676 gnd.n961 gnd.n960 585
R677 gnd.n5664 gnd.n5663 585
R678 gnd.n5663 gnd.n5662 585
R679 gnd.n967 gnd.n966 585
R680 gnd.n5661 gnd.n967 585
R681 gnd.n5659 gnd.n5658 585
R682 gnd.n5660 gnd.n5659 585
R683 gnd.n5657 gnd.n969 585
R684 gnd.n969 gnd.n968 585
R685 gnd.n5656 gnd.n5655 585
R686 gnd.n5655 gnd.n5654 585
R687 gnd.n975 gnd.n974 585
R688 gnd.n5653 gnd.n975 585
R689 gnd.n5651 gnd.n5650 585
R690 gnd.n5652 gnd.n5651 585
R691 gnd.n5649 gnd.n977 585
R692 gnd.n977 gnd.n976 585
R693 gnd.n5648 gnd.n5647 585
R694 gnd.n5647 gnd.n5646 585
R695 gnd.n983 gnd.n982 585
R696 gnd.n5645 gnd.n983 585
R697 gnd.n5643 gnd.n5642 585
R698 gnd.n5644 gnd.n5643 585
R699 gnd.n5641 gnd.n985 585
R700 gnd.n985 gnd.n984 585
R701 gnd.n5640 gnd.n5639 585
R702 gnd.n5639 gnd.n5638 585
R703 gnd.n991 gnd.n990 585
R704 gnd.n5637 gnd.n991 585
R705 gnd.n5635 gnd.n5634 585
R706 gnd.n5636 gnd.n5635 585
R707 gnd.n5633 gnd.n993 585
R708 gnd.n993 gnd.n992 585
R709 gnd.n5632 gnd.n5631 585
R710 gnd.n5631 gnd.n5630 585
R711 gnd.n999 gnd.n998 585
R712 gnd.n5629 gnd.n999 585
R713 gnd.n5627 gnd.n5626 585
R714 gnd.n5628 gnd.n5627 585
R715 gnd.n5625 gnd.n1001 585
R716 gnd.n1001 gnd.n1000 585
R717 gnd.n5624 gnd.n5623 585
R718 gnd.n5623 gnd.n5622 585
R719 gnd.n5792 gnd.n5791 585
R720 gnd.n5791 gnd.n5790 585
R721 gnd.n837 gnd.n836 585
R722 gnd.n836 gnd.n835 585
R723 gnd.n5797 gnd.n5796 585
R724 gnd.n5798 gnd.n5797 585
R725 gnd.n834 gnd.n833 585
R726 gnd.n5799 gnd.n834 585
R727 gnd.n5802 gnd.n5801 585
R728 gnd.n5801 gnd.n5800 585
R729 gnd.n831 gnd.n830 585
R730 gnd.n830 gnd.n829 585
R731 gnd.n5807 gnd.n5806 585
R732 gnd.n5808 gnd.n5807 585
R733 gnd.n828 gnd.n827 585
R734 gnd.n5809 gnd.n828 585
R735 gnd.n5812 gnd.n5811 585
R736 gnd.n5811 gnd.n5810 585
R737 gnd.n825 gnd.n824 585
R738 gnd.n824 gnd.n823 585
R739 gnd.n5817 gnd.n5816 585
R740 gnd.n5818 gnd.n5817 585
R741 gnd.n822 gnd.n821 585
R742 gnd.n5819 gnd.n822 585
R743 gnd.n5822 gnd.n5821 585
R744 gnd.n5821 gnd.n5820 585
R745 gnd.n819 gnd.n818 585
R746 gnd.n818 gnd.n817 585
R747 gnd.n5827 gnd.n5826 585
R748 gnd.n5828 gnd.n5827 585
R749 gnd.n816 gnd.n815 585
R750 gnd.n5829 gnd.n816 585
R751 gnd.n5832 gnd.n5831 585
R752 gnd.n5831 gnd.n5830 585
R753 gnd.n813 gnd.n812 585
R754 gnd.n812 gnd.n811 585
R755 gnd.n5837 gnd.n5836 585
R756 gnd.n5838 gnd.n5837 585
R757 gnd.n810 gnd.n809 585
R758 gnd.n5839 gnd.n810 585
R759 gnd.n5842 gnd.n5841 585
R760 gnd.n5841 gnd.n5840 585
R761 gnd.n807 gnd.n806 585
R762 gnd.n806 gnd.n805 585
R763 gnd.n5847 gnd.n5846 585
R764 gnd.n5848 gnd.n5847 585
R765 gnd.n804 gnd.n803 585
R766 gnd.n5849 gnd.n804 585
R767 gnd.n5852 gnd.n5851 585
R768 gnd.n5851 gnd.n5850 585
R769 gnd.n801 gnd.n800 585
R770 gnd.n800 gnd.n799 585
R771 gnd.n5857 gnd.n5856 585
R772 gnd.n5858 gnd.n5857 585
R773 gnd.n798 gnd.n797 585
R774 gnd.n5859 gnd.n798 585
R775 gnd.n5862 gnd.n5861 585
R776 gnd.n5861 gnd.n5860 585
R777 gnd.n795 gnd.n794 585
R778 gnd.n794 gnd.n793 585
R779 gnd.n5867 gnd.n5866 585
R780 gnd.n5868 gnd.n5867 585
R781 gnd.n792 gnd.n791 585
R782 gnd.n5869 gnd.n792 585
R783 gnd.n5872 gnd.n5871 585
R784 gnd.n5871 gnd.n5870 585
R785 gnd.n789 gnd.n788 585
R786 gnd.n788 gnd.n787 585
R787 gnd.n5877 gnd.n5876 585
R788 gnd.n5878 gnd.n5877 585
R789 gnd.n786 gnd.n785 585
R790 gnd.n5879 gnd.n786 585
R791 gnd.n5882 gnd.n5881 585
R792 gnd.n5881 gnd.n5880 585
R793 gnd.n783 gnd.n782 585
R794 gnd.n782 gnd.n781 585
R795 gnd.n5887 gnd.n5886 585
R796 gnd.n5888 gnd.n5887 585
R797 gnd.n780 gnd.n779 585
R798 gnd.n5889 gnd.n780 585
R799 gnd.n5892 gnd.n5891 585
R800 gnd.n5891 gnd.n5890 585
R801 gnd.n777 gnd.n776 585
R802 gnd.n776 gnd.n775 585
R803 gnd.n5897 gnd.n5896 585
R804 gnd.n5898 gnd.n5897 585
R805 gnd.n774 gnd.n773 585
R806 gnd.n5899 gnd.n774 585
R807 gnd.n5902 gnd.n5901 585
R808 gnd.n5901 gnd.n5900 585
R809 gnd.n771 gnd.n770 585
R810 gnd.n770 gnd.n769 585
R811 gnd.n5907 gnd.n5906 585
R812 gnd.n5908 gnd.n5907 585
R813 gnd.n768 gnd.n767 585
R814 gnd.n5909 gnd.n768 585
R815 gnd.n5912 gnd.n5911 585
R816 gnd.n5911 gnd.n5910 585
R817 gnd.n765 gnd.n764 585
R818 gnd.n764 gnd.n763 585
R819 gnd.n5917 gnd.n5916 585
R820 gnd.n5918 gnd.n5917 585
R821 gnd.n762 gnd.n761 585
R822 gnd.n5919 gnd.n762 585
R823 gnd.n5922 gnd.n5921 585
R824 gnd.n5921 gnd.n5920 585
R825 gnd.n759 gnd.n758 585
R826 gnd.n758 gnd.n757 585
R827 gnd.n5927 gnd.n5926 585
R828 gnd.n5928 gnd.n5927 585
R829 gnd.n756 gnd.n755 585
R830 gnd.n5929 gnd.n756 585
R831 gnd.n5932 gnd.n5931 585
R832 gnd.n5931 gnd.n5930 585
R833 gnd.n753 gnd.n752 585
R834 gnd.n752 gnd.n751 585
R835 gnd.n5937 gnd.n5936 585
R836 gnd.n5938 gnd.n5937 585
R837 gnd.n750 gnd.n749 585
R838 gnd.n5939 gnd.n750 585
R839 gnd.n5942 gnd.n5941 585
R840 gnd.n5941 gnd.n5940 585
R841 gnd.n747 gnd.n746 585
R842 gnd.n746 gnd.n745 585
R843 gnd.n5947 gnd.n5946 585
R844 gnd.n5948 gnd.n5947 585
R845 gnd.n744 gnd.n743 585
R846 gnd.n5949 gnd.n744 585
R847 gnd.n5952 gnd.n5951 585
R848 gnd.n5951 gnd.n5950 585
R849 gnd.n741 gnd.n740 585
R850 gnd.n740 gnd.n739 585
R851 gnd.n5957 gnd.n5956 585
R852 gnd.n5958 gnd.n5957 585
R853 gnd.n738 gnd.n737 585
R854 gnd.n5959 gnd.n738 585
R855 gnd.n5962 gnd.n5961 585
R856 gnd.n5961 gnd.n5960 585
R857 gnd.n735 gnd.n734 585
R858 gnd.n734 gnd.n733 585
R859 gnd.n5967 gnd.n5966 585
R860 gnd.n5968 gnd.n5967 585
R861 gnd.n732 gnd.n731 585
R862 gnd.n5969 gnd.n732 585
R863 gnd.n5972 gnd.n5971 585
R864 gnd.n5971 gnd.n5970 585
R865 gnd.n729 gnd.n728 585
R866 gnd.n728 gnd.n727 585
R867 gnd.n5977 gnd.n5976 585
R868 gnd.n5978 gnd.n5977 585
R869 gnd.n726 gnd.n725 585
R870 gnd.n5979 gnd.n726 585
R871 gnd.n5982 gnd.n5981 585
R872 gnd.n5981 gnd.n5980 585
R873 gnd.n723 gnd.n722 585
R874 gnd.n722 gnd.n721 585
R875 gnd.n5987 gnd.n5986 585
R876 gnd.n5988 gnd.n5987 585
R877 gnd.n720 gnd.n719 585
R878 gnd.n5989 gnd.n720 585
R879 gnd.n5992 gnd.n5991 585
R880 gnd.n5991 gnd.n5990 585
R881 gnd.n717 gnd.n716 585
R882 gnd.n716 gnd.n715 585
R883 gnd.n5997 gnd.n5996 585
R884 gnd.n5998 gnd.n5997 585
R885 gnd.n714 gnd.n713 585
R886 gnd.n5999 gnd.n714 585
R887 gnd.n6002 gnd.n6001 585
R888 gnd.n6001 gnd.n6000 585
R889 gnd.n711 gnd.n710 585
R890 gnd.n710 gnd.n709 585
R891 gnd.n6007 gnd.n6006 585
R892 gnd.n6008 gnd.n6007 585
R893 gnd.n708 gnd.n707 585
R894 gnd.n6009 gnd.n708 585
R895 gnd.n6012 gnd.n6011 585
R896 gnd.n6011 gnd.n6010 585
R897 gnd.n705 gnd.n704 585
R898 gnd.n704 gnd.n703 585
R899 gnd.n6017 gnd.n6016 585
R900 gnd.n6018 gnd.n6017 585
R901 gnd.n702 gnd.n701 585
R902 gnd.n6019 gnd.n702 585
R903 gnd.n6022 gnd.n6021 585
R904 gnd.n6021 gnd.n6020 585
R905 gnd.n699 gnd.n698 585
R906 gnd.n698 gnd.n697 585
R907 gnd.n6027 gnd.n6026 585
R908 gnd.n6028 gnd.n6027 585
R909 gnd.n696 gnd.n695 585
R910 gnd.n6029 gnd.n696 585
R911 gnd.n6032 gnd.n6031 585
R912 gnd.n6031 gnd.n6030 585
R913 gnd.n693 gnd.n692 585
R914 gnd.n692 gnd.n691 585
R915 gnd.n6037 gnd.n6036 585
R916 gnd.n6038 gnd.n6037 585
R917 gnd.n690 gnd.n689 585
R918 gnd.n6039 gnd.n690 585
R919 gnd.n6042 gnd.n6041 585
R920 gnd.n6041 gnd.n6040 585
R921 gnd.n687 gnd.n686 585
R922 gnd.n686 gnd.n685 585
R923 gnd.n6047 gnd.n6046 585
R924 gnd.n6048 gnd.n6047 585
R925 gnd.n684 gnd.n683 585
R926 gnd.n6049 gnd.n684 585
R927 gnd.n6052 gnd.n6051 585
R928 gnd.n6051 gnd.n6050 585
R929 gnd.n681 gnd.n680 585
R930 gnd.n680 gnd.n679 585
R931 gnd.n6057 gnd.n6056 585
R932 gnd.n6058 gnd.n6057 585
R933 gnd.n678 gnd.n677 585
R934 gnd.n6059 gnd.n678 585
R935 gnd.n6062 gnd.n6061 585
R936 gnd.n6061 gnd.n6060 585
R937 gnd.n675 gnd.n674 585
R938 gnd.n674 gnd.n673 585
R939 gnd.n6067 gnd.n6066 585
R940 gnd.n6068 gnd.n6067 585
R941 gnd.n672 gnd.n671 585
R942 gnd.n6069 gnd.n672 585
R943 gnd.n6072 gnd.n6071 585
R944 gnd.n6071 gnd.n6070 585
R945 gnd.n669 gnd.n668 585
R946 gnd.n668 gnd.n667 585
R947 gnd.n6077 gnd.n6076 585
R948 gnd.n6078 gnd.n6077 585
R949 gnd.n666 gnd.n665 585
R950 gnd.n6079 gnd.n666 585
R951 gnd.n6082 gnd.n6081 585
R952 gnd.n6081 gnd.n6080 585
R953 gnd.n663 gnd.n662 585
R954 gnd.n662 gnd.n661 585
R955 gnd.n6087 gnd.n6086 585
R956 gnd.n6088 gnd.n6087 585
R957 gnd.n660 gnd.n659 585
R958 gnd.n6089 gnd.n660 585
R959 gnd.n6092 gnd.n6091 585
R960 gnd.n6091 gnd.n6090 585
R961 gnd.n657 gnd.n656 585
R962 gnd.n656 gnd.n655 585
R963 gnd.n6097 gnd.n6096 585
R964 gnd.n6098 gnd.n6097 585
R965 gnd.n654 gnd.n653 585
R966 gnd.n6099 gnd.n654 585
R967 gnd.n6102 gnd.n6101 585
R968 gnd.n6101 gnd.n6100 585
R969 gnd.n651 gnd.n650 585
R970 gnd.n650 gnd.n649 585
R971 gnd.n6107 gnd.n6106 585
R972 gnd.n6108 gnd.n6107 585
R973 gnd.n648 gnd.n647 585
R974 gnd.n6109 gnd.n648 585
R975 gnd.n6112 gnd.n6111 585
R976 gnd.n6111 gnd.n6110 585
R977 gnd.n6324 gnd.n521 585
R978 gnd.n6324 gnd.n6323 585
R979 gnd.n6317 gnd.n522 585
R980 gnd.n6321 gnd.n522 585
R981 gnd.n6319 gnd.n6318 585
R982 gnd.n6320 gnd.n6319 585
R983 gnd.n525 gnd.n524 585
R984 gnd.n524 gnd.n523 585
R985 gnd.n6312 gnd.n6311 585
R986 gnd.n6311 gnd.n6310 585
R987 gnd.n528 gnd.n527 585
R988 gnd.n6309 gnd.n528 585
R989 gnd.n6307 gnd.n6306 585
R990 gnd.n6308 gnd.n6307 585
R991 gnd.n531 gnd.n530 585
R992 gnd.n530 gnd.n529 585
R993 gnd.n6302 gnd.n6301 585
R994 gnd.n6301 gnd.n6300 585
R995 gnd.n534 gnd.n533 585
R996 gnd.n6299 gnd.n534 585
R997 gnd.n6297 gnd.n6296 585
R998 gnd.n6298 gnd.n6297 585
R999 gnd.n537 gnd.n536 585
R1000 gnd.n536 gnd.n535 585
R1001 gnd.n6292 gnd.n6291 585
R1002 gnd.n6291 gnd.n6290 585
R1003 gnd.n540 gnd.n539 585
R1004 gnd.n6289 gnd.n540 585
R1005 gnd.n6287 gnd.n6286 585
R1006 gnd.n6288 gnd.n6287 585
R1007 gnd.n543 gnd.n542 585
R1008 gnd.n542 gnd.n541 585
R1009 gnd.n6282 gnd.n6281 585
R1010 gnd.n6281 gnd.n6280 585
R1011 gnd.n546 gnd.n545 585
R1012 gnd.n6279 gnd.n546 585
R1013 gnd.n6277 gnd.n6276 585
R1014 gnd.n6278 gnd.n6277 585
R1015 gnd.n549 gnd.n548 585
R1016 gnd.n548 gnd.n547 585
R1017 gnd.n6272 gnd.n6271 585
R1018 gnd.n6271 gnd.n6270 585
R1019 gnd.n552 gnd.n551 585
R1020 gnd.n6269 gnd.n552 585
R1021 gnd.n6267 gnd.n6266 585
R1022 gnd.n6268 gnd.n6267 585
R1023 gnd.n555 gnd.n554 585
R1024 gnd.n554 gnd.n553 585
R1025 gnd.n6262 gnd.n6261 585
R1026 gnd.n6261 gnd.n6260 585
R1027 gnd.n558 gnd.n557 585
R1028 gnd.n6259 gnd.n558 585
R1029 gnd.n6257 gnd.n6256 585
R1030 gnd.n6258 gnd.n6257 585
R1031 gnd.n561 gnd.n560 585
R1032 gnd.n560 gnd.n559 585
R1033 gnd.n6252 gnd.n6251 585
R1034 gnd.n6251 gnd.n6250 585
R1035 gnd.n564 gnd.n563 585
R1036 gnd.n6249 gnd.n564 585
R1037 gnd.n6247 gnd.n6246 585
R1038 gnd.n6248 gnd.n6247 585
R1039 gnd.n567 gnd.n566 585
R1040 gnd.n566 gnd.n565 585
R1041 gnd.n6242 gnd.n6241 585
R1042 gnd.n6241 gnd.n6240 585
R1043 gnd.n570 gnd.n569 585
R1044 gnd.n6239 gnd.n570 585
R1045 gnd.n6237 gnd.n6236 585
R1046 gnd.n6238 gnd.n6237 585
R1047 gnd.n573 gnd.n572 585
R1048 gnd.n572 gnd.n571 585
R1049 gnd.n6232 gnd.n6231 585
R1050 gnd.n6231 gnd.n6230 585
R1051 gnd.n576 gnd.n575 585
R1052 gnd.n6229 gnd.n576 585
R1053 gnd.n6227 gnd.n6226 585
R1054 gnd.n6228 gnd.n6227 585
R1055 gnd.n579 gnd.n578 585
R1056 gnd.n578 gnd.n577 585
R1057 gnd.n6222 gnd.n6221 585
R1058 gnd.n6221 gnd.n6220 585
R1059 gnd.n582 gnd.n581 585
R1060 gnd.n6219 gnd.n582 585
R1061 gnd.n6217 gnd.n6216 585
R1062 gnd.n6218 gnd.n6217 585
R1063 gnd.n585 gnd.n584 585
R1064 gnd.n584 gnd.n583 585
R1065 gnd.n6212 gnd.n6211 585
R1066 gnd.n6211 gnd.n6210 585
R1067 gnd.n588 gnd.n587 585
R1068 gnd.n6209 gnd.n588 585
R1069 gnd.n6207 gnd.n6206 585
R1070 gnd.n6208 gnd.n6207 585
R1071 gnd.n591 gnd.n590 585
R1072 gnd.n590 gnd.n589 585
R1073 gnd.n6202 gnd.n6201 585
R1074 gnd.n6201 gnd.n6200 585
R1075 gnd.n594 gnd.n593 585
R1076 gnd.n6199 gnd.n594 585
R1077 gnd.n6197 gnd.n6196 585
R1078 gnd.n6198 gnd.n6197 585
R1079 gnd.n597 gnd.n596 585
R1080 gnd.n596 gnd.n595 585
R1081 gnd.n6192 gnd.n6191 585
R1082 gnd.n6191 gnd.n6190 585
R1083 gnd.n600 gnd.n599 585
R1084 gnd.n6189 gnd.n600 585
R1085 gnd.n6187 gnd.n6186 585
R1086 gnd.n6188 gnd.n6187 585
R1087 gnd.n603 gnd.n602 585
R1088 gnd.n602 gnd.n601 585
R1089 gnd.n6182 gnd.n6181 585
R1090 gnd.n6181 gnd.n6180 585
R1091 gnd.n606 gnd.n605 585
R1092 gnd.n6179 gnd.n606 585
R1093 gnd.n6177 gnd.n6176 585
R1094 gnd.n6178 gnd.n6177 585
R1095 gnd.n609 gnd.n608 585
R1096 gnd.n608 gnd.n607 585
R1097 gnd.n6172 gnd.n6171 585
R1098 gnd.n6171 gnd.n6170 585
R1099 gnd.n612 gnd.n611 585
R1100 gnd.n6169 gnd.n612 585
R1101 gnd.n6167 gnd.n6166 585
R1102 gnd.n6168 gnd.n6167 585
R1103 gnd.n615 gnd.n614 585
R1104 gnd.n614 gnd.n613 585
R1105 gnd.n6162 gnd.n6161 585
R1106 gnd.n6161 gnd.n6160 585
R1107 gnd.n618 gnd.n617 585
R1108 gnd.n6159 gnd.n618 585
R1109 gnd.n6157 gnd.n6156 585
R1110 gnd.n6158 gnd.n6157 585
R1111 gnd.n621 gnd.n620 585
R1112 gnd.n620 gnd.n619 585
R1113 gnd.n6152 gnd.n6151 585
R1114 gnd.n6151 gnd.n6150 585
R1115 gnd.n624 gnd.n623 585
R1116 gnd.n6149 gnd.n624 585
R1117 gnd.n6147 gnd.n6146 585
R1118 gnd.n6148 gnd.n6147 585
R1119 gnd.n627 gnd.n626 585
R1120 gnd.n626 gnd.n625 585
R1121 gnd.n6142 gnd.n6141 585
R1122 gnd.n6141 gnd.n6140 585
R1123 gnd.n630 gnd.n629 585
R1124 gnd.n6139 gnd.n630 585
R1125 gnd.n6137 gnd.n6136 585
R1126 gnd.n6138 gnd.n6137 585
R1127 gnd.n633 gnd.n632 585
R1128 gnd.n632 gnd.n631 585
R1129 gnd.n6132 gnd.n6131 585
R1130 gnd.n6131 gnd.n6130 585
R1131 gnd.n636 gnd.n635 585
R1132 gnd.n6129 gnd.n636 585
R1133 gnd.n6127 gnd.n6126 585
R1134 gnd.n6128 gnd.n6127 585
R1135 gnd.n639 gnd.n638 585
R1136 gnd.n638 gnd.n637 585
R1137 gnd.n6122 gnd.n6121 585
R1138 gnd.n6121 gnd.n6120 585
R1139 gnd.n642 gnd.n641 585
R1140 gnd.n6119 gnd.n642 585
R1141 gnd.n6117 gnd.n6116 585
R1142 gnd.n6118 gnd.n6117 585
R1143 gnd.n645 gnd.n644 585
R1144 gnd.n644 gnd.n643 585
R1145 gnd.n1329 gnd.n1328 585
R1146 gnd.n2567 gnd.n1329 585
R1147 gnd.n3929 gnd.n3928 585
R1148 gnd.n3928 gnd.n3927 585
R1149 gnd.n3930 gnd.n1324 585
R1150 gnd.n2535 gnd.n1324 585
R1151 gnd.n3932 gnd.n3931 585
R1152 gnd.n3933 gnd.n3932 585
R1153 gnd.n1308 gnd.n1307 585
R1154 gnd.n2505 gnd.n1308 585
R1155 gnd.n3941 gnd.n3940 585
R1156 gnd.n3940 gnd.n3939 585
R1157 gnd.n3942 gnd.n1303 585
R1158 gnd.n2496 gnd.n1303 585
R1159 gnd.n3944 gnd.n3943 585
R1160 gnd.n3945 gnd.n3944 585
R1161 gnd.n1288 gnd.n1287 585
R1162 gnd.n1299 gnd.n1288 585
R1163 gnd.n3953 gnd.n3952 585
R1164 gnd.n3952 gnd.n3951 585
R1165 gnd.n3954 gnd.n1283 585
R1166 gnd.n1283 gnd.n1282 585
R1167 gnd.n3956 gnd.n3955 585
R1168 gnd.n3957 gnd.n3956 585
R1169 gnd.n1268 gnd.n1267 585
R1170 gnd.n1272 gnd.n1268 585
R1171 gnd.n3965 gnd.n3964 585
R1172 gnd.n3964 gnd.n3963 585
R1173 gnd.n3966 gnd.n1263 585
R1174 gnd.n1269 gnd.n1263 585
R1175 gnd.n3968 gnd.n3967 585
R1176 gnd.n3969 gnd.n3968 585
R1177 gnd.n1250 gnd.n1249 585
R1178 gnd.n1253 gnd.n1250 585
R1179 gnd.n3977 gnd.n3976 585
R1180 gnd.n3976 gnd.n3975 585
R1181 gnd.n3978 gnd.n1245 585
R1182 gnd.n1245 gnd.n1244 585
R1183 gnd.n3980 gnd.n3979 585
R1184 gnd.n3981 gnd.n3980 585
R1185 gnd.n1230 gnd.n1229 585
R1186 gnd.n1234 gnd.n1230 585
R1187 gnd.n3989 gnd.n3988 585
R1188 gnd.n3988 gnd.n3987 585
R1189 gnd.n3990 gnd.n1225 585
R1190 gnd.n1231 gnd.n1225 585
R1191 gnd.n3992 gnd.n3991 585
R1192 gnd.n3993 gnd.n3992 585
R1193 gnd.n1212 gnd.n1211 585
R1194 gnd.n1222 gnd.n1212 585
R1195 gnd.n4001 gnd.n4000 585
R1196 gnd.n4000 gnd.n3999 585
R1197 gnd.n4002 gnd.n1207 585
R1198 gnd.n1207 gnd.n1206 585
R1199 gnd.n4004 gnd.n4003 585
R1200 gnd.n4005 gnd.n4004 585
R1201 gnd.n1192 gnd.n1191 585
R1202 gnd.n1196 gnd.n1192 585
R1203 gnd.n4013 gnd.n4012 585
R1204 gnd.n4012 gnd.n4011 585
R1205 gnd.n4014 gnd.n1187 585
R1206 gnd.n1193 gnd.n1187 585
R1207 gnd.n4016 gnd.n4015 585
R1208 gnd.n4017 gnd.n4016 585
R1209 gnd.n1174 gnd.n1173 585
R1210 gnd.n1184 gnd.n1174 585
R1211 gnd.n4025 gnd.n4024 585
R1212 gnd.n4024 gnd.n4023 585
R1213 gnd.n4026 gnd.n1169 585
R1214 gnd.n1169 gnd.n1168 585
R1215 gnd.n4028 gnd.n4027 585
R1216 gnd.n4029 gnd.n4028 585
R1217 gnd.n1156 gnd.n1155 585
R1218 gnd.n1159 gnd.n1156 585
R1219 gnd.n4037 gnd.n4036 585
R1220 gnd.n4036 gnd.n4035 585
R1221 gnd.n4038 gnd.n1150 585
R1222 gnd.n1150 gnd.n1149 585
R1223 gnd.n4040 gnd.n4039 585
R1224 gnd.n4041 gnd.n4040 585
R1225 gnd.n1151 gnd.n1134 585
R1226 gnd.n1146 gnd.n1134 585
R1227 gnd.n4050 gnd.n1132 585
R1228 gnd.n4050 gnd.n4049 585
R1229 gnd.n4052 gnd.n4051 585
R1230 gnd.n4051 gnd.n1061 585
R1231 gnd.n2323 gnd.n1133 585
R1232 gnd.n2325 gnd.n2324 585
R1233 gnd.n2327 gnd.n2326 585
R1234 gnd.n2331 gnd.n2321 585
R1235 gnd.n2333 gnd.n2332 585
R1236 gnd.n2335 gnd.n2334 585
R1237 gnd.n2337 gnd.n2336 585
R1238 gnd.n2341 gnd.n2319 585
R1239 gnd.n2343 gnd.n2342 585
R1240 gnd.n2345 gnd.n2344 585
R1241 gnd.n2347 gnd.n2346 585
R1242 gnd.n2351 gnd.n2317 585
R1243 gnd.n2353 gnd.n2352 585
R1244 gnd.n2355 gnd.n2354 585
R1245 gnd.n2357 gnd.n2356 585
R1246 gnd.n2314 gnd.n2313 585
R1247 gnd.n2361 gnd.n2315 585
R1248 gnd.n2362 gnd.n2310 585
R1249 gnd.n2363 gnd.n1060 585
R1250 gnd.n4173 gnd.n1060 585
R1251 gnd.n2570 gnd.n2569 585
R1252 gnd.n2571 gnd.n2149 585
R1253 gnd.n2572 gnd.n2145 585
R1254 gnd.n2137 gnd.n2136 585
R1255 gnd.n2579 gnd.n2135 585
R1256 gnd.n2580 gnd.n2134 585
R1257 gnd.n2133 gnd.n2127 585
R1258 gnd.n2587 gnd.n2126 585
R1259 gnd.n2588 gnd.n2125 585
R1260 gnd.n2119 gnd.n2118 585
R1261 gnd.n2595 gnd.n2117 585
R1262 gnd.n2596 gnd.n2116 585
R1263 gnd.n2115 gnd.n2109 585
R1264 gnd.n2603 gnd.n2108 585
R1265 gnd.n2604 gnd.n2107 585
R1266 gnd.n2101 gnd.n2100 585
R1267 gnd.n2611 gnd.n2099 585
R1268 gnd.n2612 gnd.n2098 585
R1269 gnd.n2097 gnd.n1340 585
R1270 gnd.n3919 gnd.n1340 585
R1271 gnd.n2568 gnd.n2151 585
R1272 gnd.n2568 gnd.n2567 585
R1273 gnd.n2538 gnd.n1331 585
R1274 gnd.n3927 gnd.n1331 585
R1275 gnd.n2537 gnd.n2536 585
R1276 gnd.n2536 gnd.n2535 585
R1277 gnd.n2283 gnd.n1322 585
R1278 gnd.n3933 gnd.n1322 585
R1279 gnd.n2504 gnd.n2503 585
R1280 gnd.n2505 gnd.n2504 585
R1281 gnd.n2286 gnd.n1311 585
R1282 gnd.n3939 gnd.n1311 585
R1283 gnd.n2498 gnd.n2497 585
R1284 gnd.n2497 gnd.n2496 585
R1285 gnd.n2432 gnd.n1301 585
R1286 gnd.n3945 gnd.n1301 585
R1287 gnd.n2431 gnd.n2289 585
R1288 gnd.n2289 gnd.n1299 585
R1289 gnd.n2288 gnd.n1290 585
R1290 gnd.n3951 gnd.n1290 585
R1291 gnd.n2427 gnd.n2426 585
R1292 gnd.n2426 gnd.n1282 585
R1293 gnd.n2425 gnd.n1281 585
R1294 gnd.n3957 gnd.n1281 585
R1295 gnd.n2424 gnd.n2292 585
R1296 gnd.n2292 gnd.n1272 585
R1297 gnd.n2291 gnd.n1271 585
R1298 gnd.n3963 gnd.n1271 585
R1299 gnd.n2420 gnd.n2419 585
R1300 gnd.n2419 gnd.n1269 585
R1301 gnd.n2418 gnd.n1262 585
R1302 gnd.n3969 gnd.n1262 585
R1303 gnd.n2417 gnd.n2295 585
R1304 gnd.n2295 gnd.n1253 585
R1305 gnd.n2294 gnd.n1252 585
R1306 gnd.n3975 gnd.n1252 585
R1307 gnd.n2413 gnd.n2412 585
R1308 gnd.n2412 gnd.n1244 585
R1309 gnd.n2411 gnd.n1243 585
R1310 gnd.n3981 gnd.n1243 585
R1311 gnd.n2410 gnd.n2298 585
R1312 gnd.n2298 gnd.n1234 585
R1313 gnd.n2297 gnd.n1233 585
R1314 gnd.n3987 gnd.n1233 585
R1315 gnd.n2406 gnd.n2405 585
R1316 gnd.n2405 gnd.n1231 585
R1317 gnd.n2404 gnd.n1224 585
R1318 gnd.n3993 gnd.n1224 585
R1319 gnd.n2403 gnd.n2402 585
R1320 gnd.n2402 gnd.n1222 585
R1321 gnd.n2300 gnd.n1214 585
R1322 gnd.n3999 gnd.n1214 585
R1323 gnd.n2398 gnd.n2397 585
R1324 gnd.n2397 gnd.n1206 585
R1325 gnd.n2396 gnd.n1205 585
R1326 gnd.n4005 gnd.n1205 585
R1327 gnd.n2395 gnd.n2394 585
R1328 gnd.n2394 gnd.n1196 585
R1329 gnd.n2302 gnd.n1195 585
R1330 gnd.n4011 gnd.n1195 585
R1331 gnd.n2390 gnd.n2389 585
R1332 gnd.n2389 gnd.n1193 585
R1333 gnd.n2388 gnd.n1186 585
R1334 gnd.n4017 gnd.n1186 585
R1335 gnd.n2387 gnd.n2386 585
R1336 gnd.n2386 gnd.n1184 585
R1337 gnd.n2304 gnd.n1176 585
R1338 gnd.n4023 gnd.n1176 585
R1339 gnd.n2382 gnd.n2381 585
R1340 gnd.n2381 gnd.n1168 585
R1341 gnd.n2380 gnd.n1167 585
R1342 gnd.n4029 gnd.n1167 585
R1343 gnd.n2379 gnd.n2378 585
R1344 gnd.n2378 gnd.n1159 585
R1345 gnd.n2306 gnd.n1158 585
R1346 gnd.n4035 gnd.n1158 585
R1347 gnd.n2374 gnd.n2373 585
R1348 gnd.n2373 gnd.n1149 585
R1349 gnd.n2372 gnd.n1148 585
R1350 gnd.n4041 gnd.n1148 585
R1351 gnd.n2371 gnd.n2370 585
R1352 gnd.n2370 gnd.n1146 585
R1353 gnd.n2308 gnd.n1138 585
R1354 gnd.n4049 gnd.n1138 585
R1355 gnd.n2366 gnd.n2365 585
R1356 gnd.n2365 gnd.n1061 585
R1357 gnd.n5528 gnd.n5527 585
R1358 gnd.n5529 gnd.n5528 585
R1359 gnd.n4235 gnd.n4234 585
R1360 gnd.n4241 gnd.n4234 585
R1361 gnd.n5503 gnd.n4253 585
R1362 gnd.n4253 gnd.n4240 585
R1363 gnd.n5505 gnd.n5504 585
R1364 gnd.n5506 gnd.n5505 585
R1365 gnd.n4254 gnd.n4252 585
R1366 gnd.n4252 gnd.n4248 585
R1367 gnd.n5237 gnd.n5236 585
R1368 gnd.n5236 gnd.n5235 585
R1369 gnd.n4259 gnd.n4258 585
R1370 gnd.n5206 gnd.n4259 585
R1371 gnd.n5226 gnd.n5225 585
R1372 gnd.n5225 gnd.n5224 585
R1373 gnd.n4266 gnd.n4265 585
R1374 gnd.n5212 gnd.n4266 585
R1375 gnd.n5182 gnd.n4286 585
R1376 gnd.n4286 gnd.n4285 585
R1377 gnd.n5184 gnd.n5183 585
R1378 gnd.n5185 gnd.n5184 585
R1379 gnd.n4287 gnd.n4284 585
R1380 gnd.n4295 gnd.n4284 585
R1381 gnd.n5160 gnd.n4307 585
R1382 gnd.n4307 gnd.n4294 585
R1383 gnd.n5162 gnd.n5161 585
R1384 gnd.n5163 gnd.n5162 585
R1385 gnd.n4308 gnd.n4306 585
R1386 gnd.n4306 gnd.n4302 585
R1387 gnd.n5148 gnd.n5147 585
R1388 gnd.n5147 gnd.n5146 585
R1389 gnd.n4313 gnd.n4312 585
R1390 gnd.n4323 gnd.n4313 585
R1391 gnd.n5137 gnd.n5136 585
R1392 gnd.n5136 gnd.n5135 585
R1393 gnd.n4320 gnd.n4319 585
R1394 gnd.n5123 gnd.n4320 585
R1395 gnd.n5097 gnd.n4341 585
R1396 gnd.n4341 gnd.n4330 585
R1397 gnd.n5099 gnd.n5098 585
R1398 gnd.n5100 gnd.n5099 585
R1399 gnd.n4342 gnd.n4340 585
R1400 gnd.n4350 gnd.n4340 585
R1401 gnd.n5075 gnd.n4362 585
R1402 gnd.n4362 gnd.n4349 585
R1403 gnd.n5077 gnd.n5076 585
R1404 gnd.n5078 gnd.n5077 585
R1405 gnd.n4363 gnd.n4361 585
R1406 gnd.n4361 gnd.n4357 585
R1407 gnd.n5063 gnd.n5062 585
R1408 gnd.n5062 gnd.n5061 585
R1409 gnd.n4368 gnd.n4367 585
R1410 gnd.n4377 gnd.n4368 585
R1411 gnd.n5052 gnd.n5051 585
R1412 gnd.n5051 gnd.n5050 585
R1413 gnd.n4375 gnd.n4374 585
R1414 gnd.n5038 gnd.n4375 585
R1415 gnd.n4476 gnd.n4475 585
R1416 gnd.n4476 gnd.n4384 585
R1417 gnd.n4995 gnd.n4994 585
R1418 gnd.n4994 gnd.n4993 585
R1419 gnd.n4996 gnd.n4470 585
R1420 gnd.n4481 gnd.n4470 585
R1421 gnd.n4998 gnd.n4997 585
R1422 gnd.n4999 gnd.n4998 585
R1423 gnd.n4471 gnd.n4469 585
R1424 gnd.n4494 gnd.n4469 585
R1425 gnd.n4454 gnd.n4453 585
R1426 gnd.n4457 gnd.n4454 585
R1427 gnd.n5009 gnd.n5008 585
R1428 gnd.n5008 gnd.n5007 585
R1429 gnd.n5010 gnd.n4448 585
R1430 gnd.n4969 gnd.n4448 585
R1431 gnd.n5012 gnd.n5011 585
R1432 gnd.n5013 gnd.n5012 585
R1433 gnd.n4449 gnd.n4447 585
R1434 gnd.n4508 gnd.n4447 585
R1435 gnd.n4961 gnd.n4960 585
R1436 gnd.n4960 gnd.n4959 585
R1437 gnd.n4505 gnd.n4504 585
R1438 gnd.n4943 gnd.n4505 585
R1439 gnd.n4930 gnd.n4524 585
R1440 gnd.n4524 gnd.n4523 585
R1441 gnd.n4932 gnd.n4931 585
R1442 gnd.n4933 gnd.n4932 585
R1443 gnd.n4525 gnd.n4522 585
R1444 gnd.n4531 gnd.n4522 585
R1445 gnd.n4911 gnd.n4910 585
R1446 gnd.n4912 gnd.n4911 585
R1447 gnd.n4542 gnd.n4541 585
R1448 gnd.n4541 gnd.n4537 585
R1449 gnd.n4901 gnd.n4900 585
R1450 gnd.n4902 gnd.n4901 585
R1451 gnd.n4552 gnd.n4551 585
R1452 gnd.n4557 gnd.n4551 585
R1453 gnd.n4879 gnd.n4570 585
R1454 gnd.n4570 gnd.n4556 585
R1455 gnd.n4881 gnd.n4880 585
R1456 gnd.n4882 gnd.n4881 585
R1457 gnd.n4571 gnd.n4569 585
R1458 gnd.n4569 gnd.n4565 585
R1459 gnd.n4870 gnd.n4869 585
R1460 gnd.n4871 gnd.n4870 585
R1461 gnd.n4578 gnd.n4577 585
R1462 gnd.n4582 gnd.n4577 585
R1463 gnd.n4847 gnd.n4599 585
R1464 gnd.n4599 gnd.n4581 585
R1465 gnd.n4849 gnd.n4848 585
R1466 gnd.n4850 gnd.n4849 585
R1467 gnd.n4600 gnd.n4598 585
R1468 gnd.n4598 gnd.n4589 585
R1469 gnd.n4842 gnd.n4841 585
R1470 gnd.n4841 gnd.n4840 585
R1471 gnd.n4647 gnd.n4646 585
R1472 gnd.n4648 gnd.n4647 585
R1473 gnd.n4801 gnd.n4800 585
R1474 gnd.n4802 gnd.n4801 585
R1475 gnd.n4657 gnd.n4656 585
R1476 gnd.n4656 gnd.n4655 585
R1477 gnd.n4796 gnd.n4795 585
R1478 gnd.n4795 gnd.n4794 585
R1479 gnd.n4660 gnd.n4659 585
R1480 gnd.n4661 gnd.n4660 585
R1481 gnd.n4785 gnd.n4784 585
R1482 gnd.n4786 gnd.n4785 585
R1483 gnd.n4668 gnd.n4667 585
R1484 gnd.n4777 gnd.n4667 585
R1485 gnd.n4780 gnd.n4779 585
R1486 gnd.n4779 gnd.n4778 585
R1487 gnd.n4671 gnd.n4670 585
R1488 gnd.n4672 gnd.n4671 585
R1489 gnd.n4766 gnd.n4765 585
R1490 gnd.n4764 gnd.n4690 585
R1491 gnd.n4763 gnd.n4689 585
R1492 gnd.n4768 gnd.n4689 585
R1493 gnd.n4762 gnd.n4761 585
R1494 gnd.n4760 gnd.n4759 585
R1495 gnd.n4758 gnd.n4757 585
R1496 gnd.n4756 gnd.n4755 585
R1497 gnd.n4754 gnd.n4753 585
R1498 gnd.n4752 gnd.n4751 585
R1499 gnd.n4750 gnd.n4749 585
R1500 gnd.n4748 gnd.n4747 585
R1501 gnd.n4746 gnd.n4745 585
R1502 gnd.n4744 gnd.n4743 585
R1503 gnd.n4742 gnd.n4741 585
R1504 gnd.n4740 gnd.n4739 585
R1505 gnd.n4738 gnd.n4737 585
R1506 gnd.n4736 gnd.n4735 585
R1507 gnd.n4734 gnd.n4733 585
R1508 gnd.n4732 gnd.n4731 585
R1509 gnd.n4730 gnd.n4729 585
R1510 gnd.n4728 gnd.n4727 585
R1511 gnd.n4726 gnd.n4725 585
R1512 gnd.n4724 gnd.n4723 585
R1513 gnd.n4722 gnd.n4721 585
R1514 gnd.n4720 gnd.n4719 585
R1515 gnd.n4677 gnd.n4676 585
R1516 gnd.n4771 gnd.n4770 585
R1517 gnd.n5532 gnd.n5531 585
R1518 gnd.n5534 gnd.n5533 585
R1519 gnd.n5536 gnd.n5535 585
R1520 gnd.n5538 gnd.n5537 585
R1521 gnd.n5540 gnd.n5539 585
R1522 gnd.n5542 gnd.n5541 585
R1523 gnd.n5544 gnd.n5543 585
R1524 gnd.n5546 gnd.n5545 585
R1525 gnd.n5548 gnd.n5547 585
R1526 gnd.n5550 gnd.n5549 585
R1527 gnd.n5552 gnd.n5551 585
R1528 gnd.n5554 gnd.n5553 585
R1529 gnd.n5556 gnd.n5555 585
R1530 gnd.n5558 gnd.n5557 585
R1531 gnd.n5560 gnd.n5559 585
R1532 gnd.n5562 gnd.n5561 585
R1533 gnd.n5564 gnd.n5563 585
R1534 gnd.n5566 gnd.n5565 585
R1535 gnd.n5568 gnd.n5567 585
R1536 gnd.n5570 gnd.n5569 585
R1537 gnd.n5572 gnd.n5571 585
R1538 gnd.n5574 gnd.n5573 585
R1539 gnd.n5576 gnd.n5575 585
R1540 gnd.n5578 gnd.n5577 585
R1541 gnd.n5580 gnd.n5579 585
R1542 gnd.n5581 gnd.n4202 585
R1543 gnd.n5582 gnd.n1009 585
R1544 gnd.n5620 gnd.n1009 585
R1545 gnd.n5530 gnd.n4232 585
R1546 gnd.n5530 gnd.n5529 585
R1547 gnd.n5199 gnd.n4231 585
R1548 gnd.n4241 gnd.n4231 585
R1549 gnd.n5201 gnd.n5200 585
R1550 gnd.n5200 gnd.n4240 585
R1551 gnd.n5202 gnd.n4250 585
R1552 gnd.n5506 gnd.n4250 585
R1553 gnd.n5204 gnd.n5203 585
R1554 gnd.n5203 gnd.n4248 585
R1555 gnd.n5205 gnd.n4261 585
R1556 gnd.n5235 gnd.n4261 585
R1557 gnd.n5208 gnd.n5207 585
R1558 gnd.n5207 gnd.n5206 585
R1559 gnd.n5209 gnd.n4268 585
R1560 gnd.n5224 gnd.n4268 585
R1561 gnd.n5211 gnd.n5210 585
R1562 gnd.n5212 gnd.n5211 585
R1563 gnd.n4278 gnd.n4277 585
R1564 gnd.n4285 gnd.n4277 585
R1565 gnd.n5187 gnd.n5186 585
R1566 gnd.n5186 gnd.n5185 585
R1567 gnd.n4281 gnd.n4280 585
R1568 gnd.n4295 gnd.n4281 585
R1569 gnd.n5113 gnd.n5112 585
R1570 gnd.n5112 gnd.n4294 585
R1571 gnd.n5114 gnd.n4304 585
R1572 gnd.n5163 gnd.n4304 585
R1573 gnd.n5116 gnd.n5115 585
R1574 gnd.n5115 gnd.n4302 585
R1575 gnd.n5117 gnd.n4315 585
R1576 gnd.n5146 gnd.n4315 585
R1577 gnd.n5119 gnd.n5118 585
R1578 gnd.n5118 gnd.n4323 585
R1579 gnd.n5120 gnd.n4322 585
R1580 gnd.n5135 gnd.n4322 585
R1581 gnd.n5122 gnd.n5121 585
R1582 gnd.n5123 gnd.n5122 585
R1583 gnd.n4334 gnd.n4333 585
R1584 gnd.n4333 gnd.n4330 585
R1585 gnd.n5102 gnd.n5101 585
R1586 gnd.n5101 gnd.n5100 585
R1587 gnd.n4337 gnd.n4336 585
R1588 gnd.n4350 gnd.n4337 585
R1589 gnd.n5026 gnd.n5025 585
R1590 gnd.n5025 gnd.n4349 585
R1591 gnd.n5027 gnd.n4359 585
R1592 gnd.n5078 gnd.n4359 585
R1593 gnd.n5029 gnd.n5028 585
R1594 gnd.n5028 gnd.n4357 585
R1595 gnd.n5030 gnd.n4370 585
R1596 gnd.n5061 gnd.n4370 585
R1597 gnd.n5032 gnd.n5031 585
R1598 gnd.n5031 gnd.n4377 585
R1599 gnd.n5033 gnd.n4376 585
R1600 gnd.n5050 gnd.n4376 585
R1601 gnd.n5035 gnd.n5034 585
R1602 gnd.n5038 gnd.n5035 585
R1603 gnd.n4387 gnd.n4386 585
R1604 gnd.n4386 gnd.n4384 585
R1605 gnd.n4478 gnd.n4477 585
R1606 gnd.n4993 gnd.n4477 585
R1607 gnd.n4480 gnd.n4479 585
R1608 gnd.n4481 gnd.n4480 585
R1609 gnd.n4491 gnd.n4467 585
R1610 gnd.n4999 gnd.n4467 585
R1611 gnd.n4493 gnd.n4492 585
R1612 gnd.n4494 gnd.n4493 585
R1613 gnd.n4490 gnd.n4489 585
R1614 gnd.n4490 gnd.n4457 585
R1615 gnd.n4488 gnd.n4455 585
R1616 gnd.n5007 gnd.n4455 585
R1617 gnd.n4444 gnd.n4442 585
R1618 gnd.n4969 gnd.n4444 585
R1619 gnd.n5015 gnd.n5014 585
R1620 gnd.n5014 gnd.n5013 585
R1621 gnd.n4443 gnd.n4441 585
R1622 gnd.n4508 gnd.n4443 585
R1623 gnd.n4940 gnd.n4507 585
R1624 gnd.n4959 gnd.n4507 585
R1625 gnd.n4942 gnd.n4941 585
R1626 gnd.n4943 gnd.n4942 585
R1627 gnd.n4517 gnd.n4516 585
R1628 gnd.n4523 gnd.n4516 585
R1629 gnd.n4935 gnd.n4934 585
R1630 gnd.n4934 gnd.n4933 585
R1631 gnd.n4520 gnd.n4519 585
R1632 gnd.n4531 gnd.n4520 585
R1633 gnd.n4820 gnd.n4539 585
R1634 gnd.n4912 gnd.n4539 585
R1635 gnd.n4822 gnd.n4821 585
R1636 gnd.n4821 gnd.n4537 585
R1637 gnd.n4823 gnd.n4550 585
R1638 gnd.n4902 gnd.n4550 585
R1639 gnd.n4825 gnd.n4824 585
R1640 gnd.n4825 gnd.n4557 585
R1641 gnd.n4827 gnd.n4826 585
R1642 gnd.n4826 gnd.n4556 585
R1643 gnd.n4828 gnd.n4567 585
R1644 gnd.n4882 gnd.n4567 585
R1645 gnd.n4830 gnd.n4829 585
R1646 gnd.n4829 gnd.n4565 585
R1647 gnd.n4831 gnd.n4576 585
R1648 gnd.n4871 gnd.n4576 585
R1649 gnd.n4833 gnd.n4832 585
R1650 gnd.n4833 gnd.n4582 585
R1651 gnd.n4835 gnd.n4834 585
R1652 gnd.n4834 gnd.n4581 585
R1653 gnd.n4836 gnd.n4597 585
R1654 gnd.n4850 gnd.n4597 585
R1655 gnd.n4837 gnd.n4650 585
R1656 gnd.n4650 gnd.n4589 585
R1657 gnd.n4839 gnd.n4838 585
R1658 gnd.n4840 gnd.n4839 585
R1659 gnd.n4651 gnd.n4649 585
R1660 gnd.n4649 gnd.n4648 585
R1661 gnd.n4804 gnd.n4803 585
R1662 gnd.n4803 gnd.n4802 585
R1663 gnd.n4654 gnd.n4653 585
R1664 gnd.n4655 gnd.n4654 585
R1665 gnd.n4793 gnd.n4792 585
R1666 gnd.n4794 gnd.n4793 585
R1667 gnd.n4663 gnd.n4662 585
R1668 gnd.n4662 gnd.n4661 585
R1669 gnd.n4788 gnd.n4787 585
R1670 gnd.n4787 gnd.n4786 585
R1671 gnd.n4666 gnd.n4665 585
R1672 gnd.n4777 gnd.n4666 585
R1673 gnd.n4776 gnd.n4775 585
R1674 gnd.n4778 gnd.n4776 585
R1675 gnd.n4674 gnd.n4673 585
R1676 gnd.n4673 gnd.n4672 585
R1677 gnd.n7066 gnd.n165 585
R1678 gnd.n165 gnd.n164 585
R1679 gnd.n7068 gnd.n7067 585
R1680 gnd.n7069 gnd.n7068 585
R1681 gnd.n151 gnd.n150 585
R1682 gnd.n154 gnd.n151 585
R1683 gnd.n7077 gnd.n7076 585
R1684 gnd.n7076 gnd.n7075 585
R1685 gnd.n7078 gnd.n146 585
R1686 gnd.n146 gnd.n145 585
R1687 gnd.n7080 gnd.n7079 585
R1688 gnd.n7081 gnd.n7080 585
R1689 gnd.n132 gnd.n131 585
R1690 gnd.n142 gnd.n132 585
R1691 gnd.n7089 gnd.n7088 585
R1692 gnd.n7088 gnd.n7087 585
R1693 gnd.n7090 gnd.n127 585
R1694 gnd.n127 gnd.n126 585
R1695 gnd.n7092 gnd.n7091 585
R1696 gnd.n7093 gnd.n7092 585
R1697 gnd.n113 gnd.n112 585
R1698 gnd.n116 gnd.n113 585
R1699 gnd.n7101 gnd.n7100 585
R1700 gnd.n7100 gnd.n7099 585
R1701 gnd.n7102 gnd.n108 585
R1702 gnd.n108 gnd.n107 585
R1703 gnd.n7104 gnd.n7103 585
R1704 gnd.n7105 gnd.n7104 585
R1705 gnd.n94 gnd.n93 585
R1706 gnd.n104 gnd.n94 585
R1707 gnd.n7113 gnd.n7112 585
R1708 gnd.n7112 gnd.n7111 585
R1709 gnd.n7114 gnd.n88 585
R1710 gnd.n88 gnd.n86 585
R1711 gnd.n7116 gnd.n7115 585
R1712 gnd.n7117 gnd.n7116 585
R1713 gnd.n89 gnd.n87 585
R1714 gnd.n87 gnd.n74 585
R1715 gnd.n6699 gnd.n75 585
R1716 gnd.n7123 gnd.n75 585
R1717 gnd.n6698 gnd.n6697 585
R1718 gnd.n6697 gnd.n6696 585
R1719 gnd.n170 gnd.n169 585
R1720 gnd.n171 gnd.n170 585
R1721 gnd.n6690 gnd.n6689 585
R1722 gnd.n6689 gnd.n6688 585
R1723 gnd.n176 gnd.n175 585
R1724 gnd.n188 gnd.n176 585
R1725 gnd.n6676 gnd.n6675 585
R1726 gnd.n6677 gnd.n6676 585
R1727 gnd.n190 gnd.n189 585
R1728 gnd.n6668 gnd.n189 585
R1729 gnd.n6640 gnd.n6639 585
R1730 gnd.n6639 gnd.n194 585
R1731 gnd.n6641 gnd.n202 585
R1732 gnd.n6655 gnd.n202 585
R1733 gnd.n6642 gnd.n214 585
R1734 gnd.n214 gnd.n212 585
R1735 gnd.n6644 gnd.n6643 585
R1736 gnd.n6645 gnd.n6644 585
R1737 gnd.n215 gnd.n213 585
R1738 gnd.n213 gnd.n209 585
R1739 gnd.n6617 gnd.n223 585
R1740 gnd.n6629 gnd.n223 585
R1741 gnd.n6618 gnd.n233 585
R1742 gnd.n233 gnd.n221 585
R1743 gnd.n6620 gnd.n6619 585
R1744 gnd.n6621 gnd.n6620 585
R1745 gnd.n234 gnd.n232 585
R1746 gnd.n6610 gnd.n232 585
R1747 gnd.n6576 gnd.n6575 585
R1748 gnd.n6575 gnd.n239 585
R1749 gnd.n6577 gnd.n248 585
R1750 gnd.n6591 gnd.n248 585
R1751 gnd.n6578 gnd.n260 585
R1752 gnd.n6569 gnd.n260 585
R1753 gnd.n6580 gnd.n6579 585
R1754 gnd.n6581 gnd.n6580 585
R1755 gnd.n261 gnd.n259 585
R1756 gnd.n6565 gnd.n259 585
R1757 gnd.n6341 gnd.n6340 585
R1758 gnd.n6340 gnd.n6339 585
R1759 gnd.n6342 gnd.n276 585
R1760 gnd.n6556 gnd.n276 585
R1761 gnd.n6344 gnd.n6343 585
R1762 gnd.n6345 gnd.n6344 585
R1763 gnd.n502 gnd.n398 585
R1764 gnd.n6426 gnd.n399 585
R1765 gnd.n6425 gnd.n400 585
R1766 gnd.n407 gnd.n401 585
R1767 gnd.n6418 gnd.n408 585
R1768 gnd.n6417 gnd.n409 585
R1769 gnd.n411 gnd.n410 585
R1770 gnd.n6410 gnd.n417 585
R1771 gnd.n6409 gnd.n418 585
R1772 gnd.n425 gnd.n419 585
R1773 gnd.n6402 gnd.n426 585
R1774 gnd.n6401 gnd.n427 585
R1775 gnd.n429 gnd.n428 585
R1776 gnd.n6394 gnd.n435 585
R1777 gnd.n6393 gnd.n436 585
R1778 gnd.n445 gnd.n437 585
R1779 gnd.n6386 gnd.n446 585
R1780 gnd.n6385 gnd.n6382 585
R1781 gnd.n447 gnd.n322 585
R1782 gnd.n6546 gnd.n322 585
R1783 gnd.n6851 gnd.n6850 585
R1784 gnd.n6753 gnd.n6749 585
R1785 gnd.n6801 gnd.n6800 585
R1786 gnd.n6799 gnd.n6798 585
R1787 gnd.n6797 gnd.n6796 585
R1788 gnd.n6790 gnd.n6755 585
R1789 gnd.n6792 gnd.n6791 585
R1790 gnd.n6789 gnd.n6788 585
R1791 gnd.n6787 gnd.n6786 585
R1792 gnd.n6780 gnd.n6757 585
R1793 gnd.n6782 gnd.n6781 585
R1794 gnd.n6779 gnd.n6778 585
R1795 gnd.n6777 gnd.n6776 585
R1796 gnd.n6770 gnd.n6759 585
R1797 gnd.n6772 gnd.n6771 585
R1798 gnd.n6769 gnd.n6768 585
R1799 gnd.n6767 gnd.n6766 585
R1800 gnd.n6763 gnd.n6762 585
R1801 gnd.n6761 gnd.n6740 585
R1802 gnd.n7058 gnd.n6740 585
R1803 gnd.n6847 gnd.n6750 585
R1804 gnd.n6750 gnd.n164 585
R1805 gnd.n6846 gnd.n163 585
R1806 gnd.n7069 gnd.n163 585
R1807 gnd.n6845 gnd.n6844 585
R1808 gnd.n6844 gnd.n154 585
R1809 gnd.n6805 gnd.n153 585
R1810 gnd.n7075 gnd.n153 585
R1811 gnd.n6840 gnd.n6839 585
R1812 gnd.n6839 gnd.n145 585
R1813 gnd.n6838 gnd.n144 585
R1814 gnd.n7081 gnd.n144 585
R1815 gnd.n6837 gnd.n6836 585
R1816 gnd.n6836 gnd.n142 585
R1817 gnd.n6807 gnd.n134 585
R1818 gnd.n7087 gnd.n134 585
R1819 gnd.n6832 gnd.n6831 585
R1820 gnd.n6831 gnd.n126 585
R1821 gnd.n6830 gnd.n125 585
R1822 gnd.n7093 gnd.n125 585
R1823 gnd.n6829 gnd.n6828 585
R1824 gnd.n6828 gnd.n116 585
R1825 gnd.n6809 gnd.n115 585
R1826 gnd.n7099 gnd.n115 585
R1827 gnd.n6824 gnd.n6823 585
R1828 gnd.n6823 gnd.n107 585
R1829 gnd.n6822 gnd.n106 585
R1830 gnd.n7105 gnd.n106 585
R1831 gnd.n6821 gnd.n6820 585
R1832 gnd.n6820 gnd.n104 585
R1833 gnd.n6811 gnd.n96 585
R1834 gnd.n7111 gnd.n96 585
R1835 gnd.n6816 gnd.n6815 585
R1836 gnd.n6815 gnd.n86 585
R1837 gnd.n6814 gnd.n85 585
R1838 gnd.n7117 gnd.n85 585
R1839 gnd.n72 gnd.n71 585
R1840 gnd.n74 gnd.n72 585
R1841 gnd.n7125 gnd.n7124 585
R1842 gnd.n7124 gnd.n7123 585
R1843 gnd.n7126 gnd.n70 585
R1844 gnd.n6696 gnd.n70 585
R1845 gnd.n178 gnd.n68 585
R1846 gnd.n178 gnd.n171 585
R1847 gnd.n6661 gnd.n179 585
R1848 gnd.n6688 gnd.n179 585
R1849 gnd.n6662 gnd.n6660 585
R1850 gnd.n6660 gnd.n188 585
R1851 gnd.n197 gnd.n187 585
R1852 gnd.n6677 gnd.n187 585
R1853 gnd.n6667 gnd.n6666 585
R1854 gnd.n6668 gnd.n6667 585
R1855 gnd.n196 gnd.n195 585
R1856 gnd.n195 gnd.n194 585
R1857 gnd.n6657 gnd.n6656 585
R1858 gnd.n6656 gnd.n6655 585
R1859 gnd.n200 gnd.n199 585
R1860 gnd.n212 gnd.n200 585
R1861 gnd.n6599 gnd.n211 585
R1862 gnd.n6645 gnd.n211 585
R1863 gnd.n6602 gnd.n6598 585
R1864 gnd.n6598 gnd.n209 585
R1865 gnd.n6603 gnd.n222 585
R1866 gnd.n6629 gnd.n222 585
R1867 gnd.n6604 gnd.n6597 585
R1868 gnd.n6597 gnd.n221 585
R1869 gnd.n242 gnd.n231 585
R1870 gnd.n6621 gnd.n231 585
R1871 gnd.n6609 gnd.n6608 585
R1872 gnd.n6610 gnd.n6609 585
R1873 gnd.n241 gnd.n240 585
R1874 gnd.n240 gnd.n239 585
R1875 gnd.n6593 gnd.n6592 585
R1876 gnd.n6592 gnd.n6591 585
R1877 gnd.n245 gnd.n244 585
R1878 gnd.n6569 gnd.n245 585
R1879 gnd.n270 gnd.n257 585
R1880 gnd.n6581 gnd.n257 585
R1881 gnd.n6564 gnd.n6563 585
R1882 gnd.n6565 gnd.n6564 585
R1883 gnd.n269 gnd.n268 585
R1884 gnd.n6339 gnd.n268 585
R1885 gnd.n6558 gnd.n6557 585
R1886 gnd.n6557 gnd.n6556 585
R1887 gnd.n273 gnd.n272 585
R1888 gnd.n6345 gnd.n273 585
R1889 gnd.n5515 gnd.n4182 585
R1890 gnd.n4182 gnd.n1008 585
R1891 gnd.n5516 gnd.n4243 585
R1892 gnd.n4243 gnd.n4233 585
R1893 gnd.n5518 gnd.n5517 585
R1894 gnd.n5519 gnd.n5518 585
R1895 gnd.n4244 gnd.n4242 585
R1896 gnd.n4251 gnd.n4242 585
R1897 gnd.n5509 gnd.n5508 585
R1898 gnd.n5508 gnd.n5507 585
R1899 gnd.n4247 gnd.n4246 585
R1900 gnd.n5234 gnd.n4247 585
R1901 gnd.n5220 gnd.n4270 585
R1902 gnd.n4270 gnd.n4260 585
R1903 gnd.n5222 gnd.n5221 585
R1904 gnd.n5223 gnd.n5222 585
R1905 gnd.n4271 gnd.n4269 585
R1906 gnd.n4269 gnd.n4267 585
R1907 gnd.n5215 gnd.n5214 585
R1908 gnd.n5214 gnd.n5213 585
R1909 gnd.n4274 gnd.n4273 585
R1910 gnd.n4283 gnd.n4274 585
R1911 gnd.n5171 gnd.n4297 585
R1912 gnd.n4297 gnd.n4282 585
R1913 gnd.n5173 gnd.n5172 585
R1914 gnd.n5174 gnd.n5173 585
R1915 gnd.n4298 gnd.n4296 585
R1916 gnd.n4305 gnd.n4296 585
R1917 gnd.n5166 gnd.n5165 585
R1918 gnd.n5165 gnd.n5164 585
R1919 gnd.n4301 gnd.n4300 585
R1920 gnd.n5145 gnd.n4301 585
R1921 gnd.n5131 gnd.n4325 585
R1922 gnd.n4325 gnd.n4314 585
R1923 gnd.n5133 gnd.n5132 585
R1924 gnd.n5134 gnd.n5133 585
R1925 gnd.n4326 gnd.n4324 585
R1926 gnd.n4324 gnd.n4321 585
R1927 gnd.n5126 gnd.n5125 585
R1928 gnd.n5125 gnd.n5124 585
R1929 gnd.n4329 gnd.n4328 585
R1930 gnd.n4339 gnd.n4329 585
R1931 gnd.n5086 gnd.n4352 585
R1932 gnd.n4352 gnd.n4338 585
R1933 gnd.n5088 gnd.n5087 585
R1934 gnd.n5089 gnd.n5088 585
R1935 gnd.n4353 gnd.n4351 585
R1936 gnd.n4360 gnd.n4351 585
R1937 gnd.n5081 gnd.n5080 585
R1938 gnd.n5080 gnd.n5079 585
R1939 gnd.n4356 gnd.n4355 585
R1940 gnd.n5060 gnd.n4356 585
R1941 gnd.n5046 gnd.n4379 585
R1942 gnd.n4379 gnd.n4369 585
R1943 gnd.n5048 gnd.n5047 585
R1944 gnd.n5049 gnd.n5048 585
R1945 gnd.n4380 gnd.n4378 585
R1946 gnd.n5037 gnd.n4378 585
R1947 gnd.n5041 gnd.n5040 585
R1948 gnd.n5040 gnd.n5039 585
R1949 gnd.n4383 gnd.n4382 585
R1950 gnd.n4992 gnd.n4383 585
R1951 gnd.n4485 gnd.n4484 585
R1952 gnd.n4486 gnd.n4485 585
R1953 gnd.n4465 gnd.n4464 585
R1954 gnd.n4468 gnd.n4465 585
R1955 gnd.n5002 gnd.n5001 585
R1956 gnd.n5001 gnd.n5000 585
R1957 gnd.n5003 gnd.n4459 585
R1958 gnd.n4495 gnd.n4459 585
R1959 gnd.n5005 gnd.n5004 585
R1960 gnd.n5006 gnd.n5005 585
R1961 gnd.n4460 gnd.n4458 585
R1962 gnd.n4970 gnd.n4458 585
R1963 gnd.n4954 gnd.n4953 585
R1964 gnd.n4953 gnd.n4446 585
R1965 gnd.n4955 gnd.n4510 585
R1966 gnd.n4510 gnd.n4445 585
R1967 gnd.n4957 gnd.n4956 585
R1968 gnd.n4958 gnd.n4957 585
R1969 gnd.n4511 gnd.n4509 585
R1970 gnd.n4509 gnd.n4506 585
R1971 gnd.n4946 gnd.n4945 585
R1972 gnd.n4945 gnd.n4944 585
R1973 gnd.n4514 gnd.n4513 585
R1974 gnd.n4521 gnd.n4514 585
R1975 gnd.n4920 gnd.n4919 585
R1976 gnd.n4921 gnd.n4920 585
R1977 gnd.n4533 gnd.n4532 585
R1978 gnd.n4540 gnd.n4532 585
R1979 gnd.n4915 gnd.n4914 585
R1980 gnd.n4914 gnd.n4913 585
R1981 gnd.n4536 gnd.n4535 585
R1982 gnd.n4903 gnd.n4536 585
R1983 gnd.n4890 gnd.n4560 585
R1984 gnd.n4560 gnd.n4559 585
R1985 gnd.n4892 gnd.n4891 585
R1986 gnd.n4893 gnd.n4892 585
R1987 gnd.n4561 gnd.n4558 585
R1988 gnd.n4568 gnd.n4558 585
R1989 gnd.n4885 gnd.n4884 585
R1990 gnd.n4884 gnd.n4883 585
R1991 gnd.n4564 gnd.n4563 585
R1992 gnd.n4872 gnd.n4564 585
R1993 gnd.n4859 gnd.n4585 585
R1994 gnd.n4585 gnd.n4584 585
R1995 gnd.n4861 gnd.n4860 585
R1996 gnd.n4862 gnd.n4861 585
R1997 gnd.n4855 gnd.n4583 585
R1998 gnd.n4854 gnd.n4853 585
R1999 gnd.n4588 gnd.n4587 585
R2000 gnd.n4851 gnd.n4588 585
R2001 gnd.n4610 gnd.n4609 585
R2002 gnd.n4613 gnd.n4612 585
R2003 gnd.n4611 gnd.n4606 585
R2004 gnd.n4618 gnd.n4617 585
R2005 gnd.n4620 gnd.n4619 585
R2006 gnd.n4623 gnd.n4622 585
R2007 gnd.n4621 gnd.n4604 585
R2008 gnd.n4628 gnd.n4627 585
R2009 gnd.n4630 gnd.n4629 585
R2010 gnd.n4633 gnd.n4632 585
R2011 gnd.n4631 gnd.n4602 585
R2012 gnd.n4638 gnd.n4637 585
R2013 gnd.n4642 gnd.n4639 585
R2014 gnd.n4643 gnd.n4580 585
R2015 gnd.n5521 gnd.n4197 585
R2016 gnd.n5588 gnd.n5587 585
R2017 gnd.n5590 gnd.n5589 585
R2018 gnd.n5592 gnd.n5591 585
R2019 gnd.n5594 gnd.n5593 585
R2020 gnd.n5596 gnd.n5595 585
R2021 gnd.n5598 gnd.n5597 585
R2022 gnd.n5600 gnd.n5599 585
R2023 gnd.n5602 gnd.n5601 585
R2024 gnd.n5604 gnd.n5603 585
R2025 gnd.n5606 gnd.n5605 585
R2026 gnd.n5608 gnd.n5607 585
R2027 gnd.n5610 gnd.n5609 585
R2028 gnd.n5613 gnd.n5612 585
R2029 gnd.n5611 gnd.n4185 585
R2030 gnd.n5617 gnd.n4183 585
R2031 gnd.n5619 gnd.n5618 585
R2032 gnd.n5620 gnd.n5619 585
R2033 gnd.n5522 gnd.n4238 585
R2034 gnd.n5522 gnd.n1008 585
R2035 gnd.n5524 gnd.n5523 585
R2036 gnd.n5523 gnd.n4233 585
R2037 gnd.n5520 gnd.n4237 585
R2038 gnd.n5520 gnd.n5519 585
R2039 gnd.n5499 gnd.n4239 585
R2040 gnd.n4251 gnd.n4239 585
R2041 gnd.n5498 gnd.n4249 585
R2042 gnd.n5507 gnd.n4249 585
R2043 gnd.n5233 gnd.n4256 585
R2044 gnd.n5234 gnd.n5233 585
R2045 gnd.n5232 gnd.n5231 585
R2046 gnd.n5232 gnd.n4260 585
R2047 gnd.n5230 gnd.n4262 585
R2048 gnd.n5223 gnd.n4262 585
R2049 gnd.n4275 gnd.n4263 585
R2050 gnd.n4275 gnd.n4267 585
R2051 gnd.n5179 gnd.n4276 585
R2052 gnd.n5213 gnd.n4276 585
R2053 gnd.n5178 gnd.n5177 585
R2054 gnd.n5177 gnd.n4283 585
R2055 gnd.n5176 gnd.n4291 585
R2056 gnd.n5176 gnd.n4282 585
R2057 gnd.n5175 gnd.n4293 585
R2058 gnd.n5175 gnd.n5174 585
R2059 gnd.n5154 gnd.n4292 585
R2060 gnd.n4305 gnd.n4292 585
R2061 gnd.n5153 gnd.n4303 585
R2062 gnd.n5164 gnd.n4303 585
R2063 gnd.n5144 gnd.n4310 585
R2064 gnd.n5145 gnd.n5144 585
R2065 gnd.n5143 gnd.n5142 585
R2066 gnd.n5143 gnd.n4314 585
R2067 gnd.n5141 gnd.n4316 585
R2068 gnd.n5134 gnd.n4316 585
R2069 gnd.n4331 gnd.n4317 585
R2070 gnd.n4331 gnd.n4321 585
R2071 gnd.n5094 gnd.n4332 585
R2072 gnd.n5124 gnd.n4332 585
R2073 gnd.n5093 gnd.n5092 585
R2074 gnd.n5092 gnd.n4339 585
R2075 gnd.n5091 gnd.n4346 585
R2076 gnd.n5091 gnd.n4338 585
R2077 gnd.n5090 gnd.n4348 585
R2078 gnd.n5090 gnd.n5089 585
R2079 gnd.n5069 gnd.n4347 585
R2080 gnd.n4360 gnd.n4347 585
R2081 gnd.n5068 gnd.n4358 585
R2082 gnd.n5079 gnd.n4358 585
R2083 gnd.n5059 gnd.n4365 585
R2084 gnd.n5060 gnd.n5059 585
R2085 gnd.n5058 gnd.n5057 585
R2086 gnd.n5058 gnd.n4369 585
R2087 gnd.n5056 gnd.n4371 585
R2088 gnd.n5049 gnd.n4371 585
R2089 gnd.n5036 gnd.n4372 585
R2090 gnd.n5037 gnd.n5036 585
R2091 gnd.n4989 gnd.n4385 585
R2092 gnd.n5039 gnd.n4385 585
R2093 gnd.n4991 gnd.n4990 585
R2094 gnd.n4992 gnd.n4991 585
R2095 gnd.n4984 gnd.n4487 585
R2096 gnd.n4487 gnd.n4486 585
R2097 gnd.n4982 gnd.n4981 585
R2098 gnd.n4981 gnd.n4468 585
R2099 gnd.n4979 gnd.n4466 585
R2100 gnd.n5000 gnd.n4466 585
R2101 gnd.n4497 gnd.n4496 585
R2102 gnd.n4496 gnd.n4495 585
R2103 gnd.n4973 gnd.n4456 585
R2104 gnd.n5006 gnd.n4456 585
R2105 gnd.n4972 gnd.n4971 585
R2106 gnd.n4971 gnd.n4970 585
R2107 gnd.n4968 gnd.n4499 585
R2108 gnd.n4968 gnd.n4446 585
R2109 gnd.n4967 gnd.n4966 585
R2110 gnd.n4967 gnd.n4445 585
R2111 gnd.n4502 gnd.n4501 585
R2112 gnd.n4958 gnd.n4501 585
R2113 gnd.n4926 gnd.n4925 585
R2114 gnd.n4925 gnd.n4506 585
R2115 gnd.n4927 gnd.n4515 585
R2116 gnd.n4944 gnd.n4515 585
R2117 gnd.n4924 gnd.n4923 585
R2118 gnd.n4923 gnd.n4521 585
R2119 gnd.n4922 gnd.n4529 585
R2120 gnd.n4922 gnd.n4921 585
R2121 gnd.n4907 gnd.n4530 585
R2122 gnd.n4540 gnd.n4530 585
R2123 gnd.n4906 gnd.n4538 585
R2124 gnd.n4913 gnd.n4538 585
R2125 gnd.n4905 gnd.n4904 585
R2126 gnd.n4904 gnd.n4903 585
R2127 gnd.n4549 gnd.n4546 585
R2128 gnd.n4559 gnd.n4549 585
R2129 gnd.n4895 gnd.n4894 585
R2130 gnd.n4894 gnd.n4893 585
R2131 gnd.n4555 gnd.n4554 585
R2132 gnd.n4568 gnd.n4555 585
R2133 gnd.n4875 gnd.n4566 585
R2134 gnd.n4883 gnd.n4566 585
R2135 gnd.n4874 gnd.n4873 585
R2136 gnd.n4873 gnd.n4872 585
R2137 gnd.n4575 gnd.n4573 585
R2138 gnd.n4584 gnd.n4575 585
R2139 gnd.n4864 gnd.n4863 585
R2140 gnd.n4863 gnd.n4862 585
R2141 gnd.n3493 gnd.n3492 585
R2142 gnd.n3494 gnd.n3493 585
R2143 gnd.n3404 gnd.n1677 585
R2144 gnd.n1683 gnd.n1677 585
R2145 gnd.n3403 gnd.n3402 585
R2146 gnd.n3402 gnd.n3401 585
R2147 gnd.n1680 gnd.n1679 585
R2148 gnd.n3372 gnd.n1680 585
R2149 gnd.n3385 gnd.n3384 585
R2150 gnd.n3386 gnd.n3385 585
R2151 gnd.n3383 gnd.n1695 585
R2152 gnd.n3378 gnd.n1695 585
R2153 gnd.n3382 gnd.n3381 585
R2154 gnd.n3381 gnd.n3380 585
R2155 gnd.n1697 gnd.n1696 585
R2156 gnd.n3366 gnd.n1697 585
R2157 gnd.n3328 gnd.n3325 585
R2158 gnd.n3328 gnd.n3327 585
R2159 gnd.n3329 gnd.n3324 585
R2160 gnd.n3329 gnd.n1711 585
R2161 gnd.n3331 gnd.n3330 585
R2162 gnd.n3330 gnd.n1710 585
R2163 gnd.n3332 gnd.n1722 585
R2164 gnd.n3312 gnd.n1722 585
R2165 gnd.n3334 gnd.n3333 585
R2166 gnd.n3335 gnd.n3334 585
R2167 gnd.n3323 gnd.n1721 585
R2168 gnd.n3318 gnd.n1721 585
R2169 gnd.n3322 gnd.n3321 585
R2170 gnd.n3321 gnd.n3320 585
R2171 gnd.n1724 gnd.n1723 585
R2172 gnd.n3303 gnd.n1724 585
R2173 gnd.n3289 gnd.n1742 585
R2174 gnd.n1742 gnd.n1741 585
R2175 gnd.n3291 gnd.n3290 585
R2176 gnd.n3292 gnd.n3291 585
R2177 gnd.n3288 gnd.n1738 585
R2178 gnd.n3283 gnd.n1738 585
R2179 gnd.n3287 gnd.n3286 585
R2180 gnd.n3286 gnd.n3285 585
R2181 gnd.n1744 gnd.n1743 585
R2182 gnd.n3267 gnd.n1744 585
R2183 gnd.n3255 gnd.n1763 585
R2184 gnd.n1763 gnd.n1754 585
R2185 gnd.n3257 gnd.n3256 585
R2186 gnd.n3258 gnd.n3257 585
R2187 gnd.n3254 gnd.n1762 585
R2188 gnd.n3217 gnd.n1762 585
R2189 gnd.n3253 gnd.n3252 585
R2190 gnd.n3252 gnd.n3251 585
R2191 gnd.n1765 gnd.n1764 585
R2192 gnd.n3214 gnd.n1765 585
R2193 gnd.n3239 gnd.n3238 585
R2194 gnd.n3240 gnd.n3239 585
R2195 gnd.n3237 gnd.n1776 585
R2196 gnd.n1776 gnd.n1772 585
R2197 gnd.n3236 gnd.n3235 585
R2198 gnd.n3235 gnd.n3234 585
R2199 gnd.n1778 gnd.n1777 585
R2200 gnd.n3204 gnd.n1778 585
R2201 gnd.n3190 gnd.n3189 585
R2202 gnd.n3189 gnd.n1788 585
R2203 gnd.n3191 gnd.n1798 585
R2204 gnd.n3174 gnd.n1798 585
R2205 gnd.n3193 gnd.n3192 585
R2206 gnd.n3194 gnd.n3193 585
R2207 gnd.n3188 gnd.n1797 585
R2208 gnd.n1797 gnd.n1794 585
R2209 gnd.n3187 gnd.n3186 585
R2210 gnd.n3186 gnd.n3185 585
R2211 gnd.n1800 gnd.n1799 585
R2212 gnd.n3165 gnd.n1800 585
R2213 gnd.n3150 gnd.n3149 585
R2214 gnd.n3149 gnd.n1811 585
R2215 gnd.n3151 gnd.n1821 585
R2216 gnd.n3134 gnd.n1821 585
R2217 gnd.n3153 gnd.n3152 585
R2218 gnd.n3154 gnd.n3153 585
R2219 gnd.n3148 gnd.n1820 585
R2220 gnd.n1820 gnd.n1817 585
R2221 gnd.n3147 gnd.n3146 585
R2222 gnd.n3146 gnd.n3145 585
R2223 gnd.n1823 gnd.n1822 585
R2224 gnd.n3125 gnd.n1823 585
R2225 gnd.n3110 gnd.n3109 585
R2226 gnd.n3109 gnd.n1834 585
R2227 gnd.n3111 gnd.n1843 585
R2228 gnd.n3095 gnd.n1843 585
R2229 gnd.n3113 gnd.n3112 585
R2230 gnd.n3114 gnd.n3113 585
R2231 gnd.n3108 gnd.n1842 585
R2232 gnd.n3101 gnd.n1842 585
R2233 gnd.n3107 gnd.n3106 585
R2234 gnd.n3106 gnd.n3105 585
R2235 gnd.n1845 gnd.n1844 585
R2236 gnd.n3068 gnd.n1845 585
R2237 gnd.n3081 gnd.n3080 585
R2238 gnd.n3082 gnd.n3081 585
R2239 gnd.n3079 gnd.n1857 585
R2240 gnd.n3074 gnd.n1857 585
R2241 gnd.n3078 gnd.n3077 585
R2242 gnd.n3077 gnd.n3076 585
R2243 gnd.n1859 gnd.n1858 585
R2244 gnd.n3055 gnd.n1859 585
R2245 gnd.n3046 gnd.n1876 585
R2246 gnd.n1876 gnd.n1868 585
R2247 gnd.n3048 gnd.n3047 585
R2248 gnd.n3049 gnd.n3048 585
R2249 gnd.n3045 gnd.n1875 585
R2250 gnd.n1881 gnd.n1875 585
R2251 gnd.n3044 gnd.n3043 585
R2252 gnd.n3043 gnd.n3042 585
R2253 gnd.n1878 gnd.n1877 585
R2254 gnd.n2842 gnd.n1878 585
R2255 gnd.n3029 gnd.n3028 585
R2256 gnd.n3030 gnd.n3029 585
R2257 gnd.n3027 gnd.n1891 585
R2258 gnd.n1891 gnd.n1887 585
R2259 gnd.n3026 gnd.n3025 585
R2260 gnd.n3025 gnd.n3024 585
R2261 gnd.n1893 gnd.n1892 585
R2262 gnd.n2850 gnd.n1893 585
R2263 gnd.n2998 gnd.n2997 585
R2264 gnd.n2999 gnd.n2998 585
R2265 gnd.n2996 gnd.n1906 585
R2266 gnd.n1906 gnd.n1903 585
R2267 gnd.n2995 gnd.n2994 585
R2268 gnd.n2994 gnd.n2993 585
R2269 gnd.n1908 gnd.n1907 585
R2270 gnd.n2857 gnd.n1908 585
R2271 gnd.n2978 gnd.n2977 585
R2272 gnd.n2979 gnd.n2978 585
R2273 gnd.n2976 gnd.n1919 585
R2274 gnd.n2971 gnd.n1919 585
R2275 gnd.n2975 gnd.n2974 585
R2276 gnd.n2974 gnd.n2973 585
R2277 gnd.n1921 gnd.n1920 585
R2278 gnd.n2959 gnd.n1921 585
R2279 gnd.n2945 gnd.n1942 585
R2280 gnd.n2864 gnd.n1942 585
R2281 gnd.n2947 gnd.n2946 585
R2282 gnd.n2948 gnd.n2947 585
R2283 gnd.n2944 gnd.n1941 585
R2284 gnd.n1941 gnd.n1938 585
R2285 gnd.n2943 gnd.n2942 585
R2286 gnd.n2942 gnd.n2941 585
R2287 gnd.n1944 gnd.n1943 585
R2288 gnd.n2873 gnd.n1944 585
R2289 gnd.n2929 gnd.n2928 585
R2290 gnd.n2930 gnd.n2929 585
R2291 gnd.n2927 gnd.n1954 585
R2292 gnd.n1954 gnd.n1951 585
R2293 gnd.n2926 gnd.n2925 585
R2294 gnd.n2925 gnd.n2924 585
R2295 gnd.n1956 gnd.n1955 585
R2296 gnd.n2881 gnd.n1956 585
R2297 gnd.n2911 gnd.n2910 585
R2298 gnd.n2912 gnd.n2911 585
R2299 gnd.n2909 gnd.n1967 585
R2300 gnd.n2904 gnd.n1967 585
R2301 gnd.n2908 gnd.n2907 585
R2302 gnd.n2907 gnd.n2906 585
R2303 gnd.n1470 gnd.n1469 585
R2304 gnd.n2887 gnd.n1470 585
R2305 gnd.n3797 gnd.n3796 585
R2306 gnd.n3796 gnd.n3795 585
R2307 gnd.n3798 gnd.n1448 585
R2308 gnd.n2893 gnd.n1448 585
R2309 gnd.n3863 gnd.n3862 585
R2310 gnd.n3861 gnd.n1447 585
R2311 gnd.n3860 gnd.n1446 585
R2312 gnd.n3865 gnd.n1446 585
R2313 gnd.n3859 gnd.n3858 585
R2314 gnd.n3857 gnd.n3856 585
R2315 gnd.n3855 gnd.n3854 585
R2316 gnd.n3853 gnd.n3852 585
R2317 gnd.n3851 gnd.n3850 585
R2318 gnd.n3849 gnd.n3848 585
R2319 gnd.n3847 gnd.n3846 585
R2320 gnd.n3845 gnd.n3844 585
R2321 gnd.n3843 gnd.n3842 585
R2322 gnd.n3841 gnd.n3840 585
R2323 gnd.n3839 gnd.n3838 585
R2324 gnd.n3837 gnd.n3836 585
R2325 gnd.n3835 gnd.n3834 585
R2326 gnd.n3833 gnd.n3832 585
R2327 gnd.n3831 gnd.n3830 585
R2328 gnd.n3829 gnd.n3828 585
R2329 gnd.n3827 gnd.n3826 585
R2330 gnd.n3825 gnd.n3824 585
R2331 gnd.n3823 gnd.n3822 585
R2332 gnd.n3821 gnd.n3820 585
R2333 gnd.n3819 gnd.n3818 585
R2334 gnd.n3817 gnd.n3816 585
R2335 gnd.n3815 gnd.n3814 585
R2336 gnd.n3813 gnd.n3812 585
R2337 gnd.n3811 gnd.n3810 585
R2338 gnd.n3809 gnd.n3808 585
R2339 gnd.n3807 gnd.n3806 585
R2340 gnd.n3805 gnd.n3804 585
R2341 gnd.n3803 gnd.n1410 585
R2342 gnd.n3868 gnd.n3867 585
R2343 gnd.n1412 gnd.n1409 585
R2344 gnd.n2779 gnd.n2778 585
R2345 gnd.n2781 gnd.n2780 585
R2346 gnd.n2784 gnd.n2783 585
R2347 gnd.n2786 gnd.n2785 585
R2348 gnd.n2788 gnd.n2787 585
R2349 gnd.n2790 gnd.n2789 585
R2350 gnd.n2792 gnd.n2791 585
R2351 gnd.n2794 gnd.n2793 585
R2352 gnd.n2796 gnd.n2795 585
R2353 gnd.n2798 gnd.n2797 585
R2354 gnd.n2800 gnd.n2799 585
R2355 gnd.n2802 gnd.n2801 585
R2356 gnd.n2804 gnd.n2803 585
R2357 gnd.n2806 gnd.n2805 585
R2358 gnd.n2808 gnd.n2807 585
R2359 gnd.n2810 gnd.n2809 585
R2360 gnd.n2812 gnd.n2811 585
R2361 gnd.n2814 gnd.n2813 585
R2362 gnd.n2816 gnd.n2815 585
R2363 gnd.n2818 gnd.n2817 585
R2364 gnd.n2820 gnd.n2819 585
R2365 gnd.n2822 gnd.n2821 585
R2366 gnd.n2824 gnd.n2823 585
R2367 gnd.n2826 gnd.n2825 585
R2368 gnd.n2828 gnd.n2827 585
R2369 gnd.n2830 gnd.n2829 585
R2370 gnd.n2832 gnd.n2831 585
R2371 gnd.n2834 gnd.n2833 585
R2372 gnd.n2836 gnd.n2835 585
R2373 gnd.n2838 gnd.n2837 585
R2374 gnd.n2839 gnd.n2775 585
R2375 gnd.n3497 gnd.n3496 585
R2376 gnd.n3499 gnd.n3498 585
R2377 gnd.n3501 gnd.n3500 585
R2378 gnd.n3503 gnd.n3502 585
R2379 gnd.n3505 gnd.n3504 585
R2380 gnd.n3507 gnd.n3506 585
R2381 gnd.n3509 gnd.n3508 585
R2382 gnd.n3511 gnd.n3510 585
R2383 gnd.n3513 gnd.n3512 585
R2384 gnd.n3515 gnd.n3514 585
R2385 gnd.n3517 gnd.n3516 585
R2386 gnd.n3519 gnd.n3518 585
R2387 gnd.n3521 gnd.n3520 585
R2388 gnd.n3523 gnd.n3522 585
R2389 gnd.n3525 gnd.n3524 585
R2390 gnd.n3527 gnd.n3526 585
R2391 gnd.n3529 gnd.n3528 585
R2392 gnd.n3531 gnd.n3530 585
R2393 gnd.n3533 gnd.n3532 585
R2394 gnd.n3535 gnd.n3534 585
R2395 gnd.n3537 gnd.n3536 585
R2396 gnd.n3539 gnd.n3538 585
R2397 gnd.n3541 gnd.n3540 585
R2398 gnd.n3543 gnd.n3542 585
R2399 gnd.n3545 gnd.n3544 585
R2400 gnd.n3547 gnd.n3546 585
R2401 gnd.n3549 gnd.n3548 585
R2402 gnd.n3551 gnd.n3550 585
R2403 gnd.n3553 gnd.n3552 585
R2404 gnd.n3556 gnd.n3555 585
R2405 gnd.n3558 gnd.n3557 585
R2406 gnd.n3560 gnd.n3559 585
R2407 gnd.n3562 gnd.n3561 585
R2408 gnd.n3426 gnd.n351 585
R2409 gnd.n3428 gnd.n3427 585
R2410 gnd.n3430 gnd.n3429 585
R2411 gnd.n3432 gnd.n3431 585
R2412 gnd.n3435 gnd.n3434 585
R2413 gnd.n3437 gnd.n3436 585
R2414 gnd.n3439 gnd.n3438 585
R2415 gnd.n3441 gnd.n3440 585
R2416 gnd.n3443 gnd.n3442 585
R2417 gnd.n3445 gnd.n3444 585
R2418 gnd.n3447 gnd.n3446 585
R2419 gnd.n3449 gnd.n3448 585
R2420 gnd.n3451 gnd.n3450 585
R2421 gnd.n3453 gnd.n3452 585
R2422 gnd.n3455 gnd.n3454 585
R2423 gnd.n3457 gnd.n3456 585
R2424 gnd.n3459 gnd.n3458 585
R2425 gnd.n3461 gnd.n3460 585
R2426 gnd.n3463 gnd.n3462 585
R2427 gnd.n3465 gnd.n3464 585
R2428 gnd.n3467 gnd.n3466 585
R2429 gnd.n3469 gnd.n3468 585
R2430 gnd.n3471 gnd.n3470 585
R2431 gnd.n3473 gnd.n3472 585
R2432 gnd.n3475 gnd.n3474 585
R2433 gnd.n3477 gnd.n3476 585
R2434 gnd.n3479 gnd.n3478 585
R2435 gnd.n3481 gnd.n3480 585
R2436 gnd.n3483 gnd.n3482 585
R2437 gnd.n3485 gnd.n3484 585
R2438 gnd.n3487 gnd.n3486 585
R2439 gnd.n3489 gnd.n3488 585
R2440 gnd.n3490 gnd.n1678 585
R2441 gnd.n3495 gnd.n1673 585
R2442 gnd.n3495 gnd.n3494 585
R2443 gnd.n3370 gnd.n1674 585
R2444 gnd.n1683 gnd.n1674 585
R2445 gnd.n3371 gnd.n1682 585
R2446 gnd.n3401 gnd.n1682 585
R2447 gnd.n3374 gnd.n3373 585
R2448 gnd.n3373 gnd.n3372 585
R2449 gnd.n3375 gnd.n1691 585
R2450 gnd.n3386 gnd.n1691 585
R2451 gnd.n3377 gnd.n3376 585
R2452 gnd.n3378 gnd.n3377 585
R2453 gnd.n3369 gnd.n1699 585
R2454 gnd.n3380 gnd.n1699 585
R2455 gnd.n3368 gnd.n3367 585
R2456 gnd.n3367 gnd.n3366 585
R2457 gnd.n1702 gnd.n1701 585
R2458 gnd.n3327 gnd.n1702 585
R2459 gnd.n3309 gnd.n3308 585
R2460 gnd.n3309 gnd.n1711 585
R2461 gnd.n3310 gnd.n3307 585
R2462 gnd.n3310 gnd.n1710 585
R2463 gnd.n3314 gnd.n3313 585
R2464 gnd.n3313 gnd.n3312 585
R2465 gnd.n3315 gnd.n1719 585
R2466 gnd.n3335 gnd.n1719 585
R2467 gnd.n3317 gnd.n3316 585
R2468 gnd.n3318 gnd.n3317 585
R2469 gnd.n3306 gnd.n1725 585
R2470 gnd.n3320 gnd.n1725 585
R2471 gnd.n3305 gnd.n3304 585
R2472 gnd.n3304 gnd.n3303 585
R2473 gnd.n1727 gnd.n1726 585
R2474 gnd.n1741 gnd.n1727 585
R2475 gnd.n3262 gnd.n1736 585
R2476 gnd.n3292 gnd.n1736 585
R2477 gnd.n3263 gnd.n1747 585
R2478 gnd.n3283 gnd.n1747 585
R2479 gnd.n3264 gnd.n1746 585
R2480 gnd.n3285 gnd.n1746 585
R2481 gnd.n3266 gnd.n3265 585
R2482 gnd.n3267 gnd.n3266 585
R2483 gnd.n3261 gnd.n1756 585
R2484 gnd.n1756 gnd.n1754 585
R2485 gnd.n3260 gnd.n3259 585
R2486 gnd.n3259 gnd.n3258 585
R2487 gnd.n1758 gnd.n1757 585
R2488 gnd.n3217 gnd.n1758 585
R2489 gnd.n3211 gnd.n1766 585
R2490 gnd.n3251 gnd.n1766 585
R2491 gnd.n3213 gnd.n3212 585
R2492 gnd.n3214 gnd.n3213 585
R2493 gnd.n3210 gnd.n1774 585
R2494 gnd.n3240 gnd.n1774 585
R2495 gnd.n3209 gnd.n3208 585
R2496 gnd.n3208 gnd.n1772 585
R2497 gnd.n3207 gnd.n1780 585
R2498 gnd.n3234 gnd.n1780 585
R2499 gnd.n3206 gnd.n3205 585
R2500 gnd.n3205 gnd.n3204 585
R2501 gnd.n1787 gnd.n1786 585
R2502 gnd.n1788 gnd.n1787 585
R2503 gnd.n3173 gnd.n3172 585
R2504 gnd.n3174 gnd.n3173 585
R2505 gnd.n3171 gnd.n1795 585
R2506 gnd.n3194 gnd.n1795 585
R2507 gnd.n3170 gnd.n3169 585
R2508 gnd.n3169 gnd.n1794 585
R2509 gnd.n3168 gnd.n1802 585
R2510 gnd.n3185 gnd.n1802 585
R2511 gnd.n3167 gnd.n3166 585
R2512 gnd.n3166 gnd.n3165 585
R2513 gnd.n1810 gnd.n1809 585
R2514 gnd.n1811 gnd.n1810 585
R2515 gnd.n3133 gnd.n3132 585
R2516 gnd.n3134 gnd.n3133 585
R2517 gnd.n3131 gnd.n1818 585
R2518 gnd.n3154 gnd.n1818 585
R2519 gnd.n3130 gnd.n3129 585
R2520 gnd.n3129 gnd.n1817 585
R2521 gnd.n3128 gnd.n1825 585
R2522 gnd.n3145 gnd.n1825 585
R2523 gnd.n3127 gnd.n3126 585
R2524 gnd.n3126 gnd.n3125 585
R2525 gnd.n1833 gnd.n1832 585
R2526 gnd.n1834 gnd.n1833 585
R2527 gnd.n3097 gnd.n3096 585
R2528 gnd.n3096 gnd.n3095 585
R2529 gnd.n3098 gnd.n1840 585
R2530 gnd.n3114 gnd.n1840 585
R2531 gnd.n3100 gnd.n3099 585
R2532 gnd.n3101 gnd.n3100 585
R2533 gnd.n1849 gnd.n1847 585
R2534 gnd.n3105 gnd.n1847 585
R2535 gnd.n3070 gnd.n3069 585
R2536 gnd.n3069 gnd.n3068 585
R2537 gnd.n3071 gnd.n1856 585
R2538 gnd.n3082 gnd.n1856 585
R2539 gnd.n3073 gnd.n3072 585
R2540 gnd.n3074 gnd.n3073 585
R2541 gnd.n1862 gnd.n1861 585
R2542 gnd.n3076 gnd.n1861 585
R2543 gnd.n3054 gnd.n3053 585
R2544 gnd.n3055 gnd.n3054 585
R2545 gnd.n3052 gnd.n1870 585
R2546 gnd.n1870 gnd.n1868 585
R2547 gnd.n3051 gnd.n3050 585
R2548 gnd.n3050 gnd.n3049 585
R2549 gnd.n1872 gnd.n1871 585
R2550 gnd.n1881 gnd.n1872 585
R2551 gnd.n2840 gnd.n1880 585
R2552 gnd.n3042 gnd.n1880 585
R2553 gnd.n2844 gnd.n2843 585
R2554 gnd.n2843 gnd.n2842 585
R2555 gnd.n2845 gnd.n1888 585
R2556 gnd.n3030 gnd.n1888 585
R2557 gnd.n2847 gnd.n2846 585
R2558 gnd.n2846 gnd.n1887 585
R2559 gnd.n2848 gnd.n1895 585
R2560 gnd.n3024 gnd.n1895 585
R2561 gnd.n2852 gnd.n2851 585
R2562 gnd.n2851 gnd.n2850 585
R2563 gnd.n2853 gnd.n1904 585
R2564 gnd.n2999 gnd.n1904 585
R2565 gnd.n2855 gnd.n2854 585
R2566 gnd.n2854 gnd.n1903 585
R2567 gnd.n2856 gnd.n1910 585
R2568 gnd.n2993 gnd.n1910 585
R2569 gnd.n2859 gnd.n2858 585
R2570 gnd.n2858 gnd.n2857 585
R2571 gnd.n2860 gnd.n1917 585
R2572 gnd.n2979 gnd.n1917 585
R2573 gnd.n2861 gnd.n1924 585
R2574 gnd.n2971 gnd.n1924 585
R2575 gnd.n2862 gnd.n1923 585
R2576 gnd.n2973 gnd.n1923 585
R2577 gnd.n2863 gnd.n1932 585
R2578 gnd.n2959 gnd.n1932 585
R2579 gnd.n2866 gnd.n2865 585
R2580 gnd.n2865 gnd.n2864 585
R2581 gnd.n2867 gnd.n1939 585
R2582 gnd.n2948 gnd.n1939 585
R2583 gnd.n2869 gnd.n2868 585
R2584 gnd.n2868 gnd.n1938 585
R2585 gnd.n2870 gnd.n1945 585
R2586 gnd.n2941 gnd.n1945 585
R2587 gnd.n2875 gnd.n2874 585
R2588 gnd.n2874 gnd.n2873 585
R2589 gnd.n2876 gnd.n1952 585
R2590 gnd.n2930 gnd.n1952 585
R2591 gnd.n2878 gnd.n2877 585
R2592 gnd.n2877 gnd.n1951 585
R2593 gnd.n2879 gnd.n1958 585
R2594 gnd.n2924 gnd.n1958 585
R2595 gnd.n2883 gnd.n2882 585
R2596 gnd.n2882 gnd.n2881 585
R2597 gnd.n2884 gnd.n1965 585
R2598 gnd.n2912 gnd.n1965 585
R2599 gnd.n2885 gnd.n1970 585
R2600 gnd.n2904 gnd.n1970 585
R2601 gnd.n2886 gnd.n1969 585
R2602 gnd.n2906 gnd.n1969 585
R2603 gnd.n2889 gnd.n2888 585
R2604 gnd.n2888 gnd.n2887 585
R2605 gnd.n2890 gnd.n1472 585
R2606 gnd.n3795 gnd.n1472 585
R2607 gnd.n2892 gnd.n2891 585
R2608 gnd.n2893 gnd.n2892 585
R2609 gnd.n3924 gnd.n1333 585
R2610 gnd.n2567 gnd.n1333 585
R2611 gnd.n3926 gnd.n3925 585
R2612 gnd.n3927 gnd.n3926 585
R2613 gnd.n1319 gnd.n1318 585
R2614 gnd.n2535 gnd.n1319 585
R2615 gnd.n3935 gnd.n3934 585
R2616 gnd.n3934 gnd.n3933 585
R2617 gnd.n3936 gnd.n1313 585
R2618 gnd.n2505 gnd.n1313 585
R2619 gnd.n3938 gnd.n3937 585
R2620 gnd.n3939 gnd.n3938 585
R2621 gnd.n1298 gnd.n1297 585
R2622 gnd.n2496 gnd.n1298 585
R2623 gnd.n3947 gnd.n3946 585
R2624 gnd.n3946 gnd.n3945 585
R2625 gnd.n3948 gnd.n1292 585
R2626 gnd.n1299 gnd.n1292 585
R2627 gnd.n3950 gnd.n3949 585
R2628 gnd.n3951 gnd.n3950 585
R2629 gnd.n1279 gnd.n1278 585
R2630 gnd.n1282 gnd.n1279 585
R2631 gnd.n3959 gnd.n3958 585
R2632 gnd.n3958 gnd.n3957 585
R2633 gnd.n3960 gnd.n1273 585
R2634 gnd.n1273 gnd.n1272 585
R2635 gnd.n3962 gnd.n3961 585
R2636 gnd.n3963 gnd.n3962 585
R2637 gnd.n1260 gnd.n1259 585
R2638 gnd.n1269 gnd.n1260 585
R2639 gnd.n3971 gnd.n3970 585
R2640 gnd.n3970 gnd.n3969 585
R2641 gnd.n3972 gnd.n1254 585
R2642 gnd.n1254 gnd.n1253 585
R2643 gnd.n3974 gnd.n3973 585
R2644 gnd.n3975 gnd.n3974 585
R2645 gnd.n1241 gnd.n1240 585
R2646 gnd.n1244 gnd.n1241 585
R2647 gnd.n3983 gnd.n3982 585
R2648 gnd.n3982 gnd.n3981 585
R2649 gnd.n3984 gnd.n1235 585
R2650 gnd.n1235 gnd.n1234 585
R2651 gnd.n3986 gnd.n3985 585
R2652 gnd.n3987 gnd.n3986 585
R2653 gnd.n1221 gnd.n1220 585
R2654 gnd.n1231 gnd.n1221 585
R2655 gnd.n3995 gnd.n3994 585
R2656 gnd.n3994 gnd.n3993 585
R2657 gnd.n3996 gnd.n1215 585
R2658 gnd.n1222 gnd.n1215 585
R2659 gnd.n3998 gnd.n3997 585
R2660 gnd.n3999 gnd.n3998 585
R2661 gnd.n1203 gnd.n1202 585
R2662 gnd.n1206 gnd.n1203 585
R2663 gnd.n4007 gnd.n4006 585
R2664 gnd.n4006 gnd.n4005 585
R2665 gnd.n4008 gnd.n1197 585
R2666 gnd.n1197 gnd.n1196 585
R2667 gnd.n4010 gnd.n4009 585
R2668 gnd.n4011 gnd.n4010 585
R2669 gnd.n1183 gnd.n1182 585
R2670 gnd.n1193 gnd.n1183 585
R2671 gnd.n4019 gnd.n4018 585
R2672 gnd.n4018 gnd.n4017 585
R2673 gnd.n4020 gnd.n1177 585
R2674 gnd.n1184 gnd.n1177 585
R2675 gnd.n4022 gnd.n4021 585
R2676 gnd.n4023 gnd.n4022 585
R2677 gnd.n1165 gnd.n1164 585
R2678 gnd.n1168 gnd.n1165 585
R2679 gnd.n4031 gnd.n4030 585
R2680 gnd.n4030 gnd.n4029 585
R2681 gnd.n4032 gnd.n1160 585
R2682 gnd.n1160 gnd.n1159 585
R2683 gnd.n4034 gnd.n4033 585
R2684 gnd.n4035 gnd.n4034 585
R2685 gnd.n1145 gnd.n1144 585
R2686 gnd.n1149 gnd.n1145 585
R2687 gnd.n4043 gnd.n4042 585
R2688 gnd.n4042 gnd.n4041 585
R2689 gnd.n1141 gnd.n1139 585
R2690 gnd.n1146 gnd.n1139 585
R2691 gnd.n4048 gnd.n4047 585
R2692 gnd.n4049 gnd.n4048 585
R2693 gnd.n1140 gnd.n1064 585
R2694 gnd.n1064 gnd.n1061 585
R2695 gnd.n4171 gnd.n4170 585
R2696 gnd.n4169 gnd.n1063 585
R2697 gnd.n4168 gnd.n1062 585
R2698 gnd.n4173 gnd.n1062 585
R2699 gnd.n4167 gnd.n4166 585
R2700 gnd.n4165 gnd.n4164 585
R2701 gnd.n4163 gnd.n4162 585
R2702 gnd.n4161 gnd.n4160 585
R2703 gnd.n4159 gnd.n4158 585
R2704 gnd.n4157 gnd.n4156 585
R2705 gnd.n4155 gnd.n4154 585
R2706 gnd.n4153 gnd.n4152 585
R2707 gnd.n4151 gnd.n4150 585
R2708 gnd.n4149 gnd.n4148 585
R2709 gnd.n4147 gnd.n4146 585
R2710 gnd.n4145 gnd.n4144 585
R2711 gnd.n4143 gnd.n4142 585
R2712 gnd.n4141 gnd.n4140 585
R2713 gnd.n4139 gnd.n4138 585
R2714 gnd.n4136 gnd.n4135 585
R2715 gnd.n4134 gnd.n4133 585
R2716 gnd.n4132 gnd.n4131 585
R2717 gnd.n4130 gnd.n4129 585
R2718 gnd.n4128 gnd.n4127 585
R2719 gnd.n4126 gnd.n4125 585
R2720 gnd.n4124 gnd.n4123 585
R2721 gnd.n4122 gnd.n4121 585
R2722 gnd.n4120 gnd.n4119 585
R2723 gnd.n4118 gnd.n4117 585
R2724 gnd.n4116 gnd.n4115 585
R2725 gnd.n4114 gnd.n4113 585
R2726 gnd.n4112 gnd.n4111 585
R2727 gnd.n4110 gnd.n4109 585
R2728 gnd.n4108 gnd.n4107 585
R2729 gnd.n4106 gnd.n4105 585
R2730 gnd.n4104 gnd.n4103 585
R2731 gnd.n4102 gnd.n4101 585
R2732 gnd.n4100 gnd.n4099 585
R2733 gnd.n4098 gnd.n4097 585
R2734 gnd.n4096 gnd.n4095 585
R2735 gnd.n4094 gnd.n4093 585
R2736 gnd.n4092 gnd.n4091 585
R2737 gnd.n4090 gnd.n4089 585
R2738 gnd.n4088 gnd.n4087 585
R2739 gnd.n4086 gnd.n4085 585
R2740 gnd.n4084 gnd.n4083 585
R2741 gnd.n4082 gnd.n4081 585
R2742 gnd.n4080 gnd.n4079 585
R2743 gnd.n4078 gnd.n4077 585
R2744 gnd.n4076 gnd.n4075 585
R2745 gnd.n4074 gnd.n4073 585
R2746 gnd.n4072 gnd.n4071 585
R2747 gnd.n4070 gnd.n4069 585
R2748 gnd.n4068 gnd.n4067 585
R2749 gnd.n4066 gnd.n4065 585
R2750 gnd.n4064 gnd.n4063 585
R2751 gnd.n4062 gnd.n4061 585
R2752 gnd.n4060 gnd.n4059 585
R2753 gnd.n4058 gnd.n4057 585
R2754 gnd.n1135 gnd.n1126 585
R2755 gnd.n2247 gnd.n2246 585
R2756 gnd.n2240 gnd.n2154 585
R2757 gnd.n2242 gnd.n2241 585
R2758 gnd.n2239 gnd.n2238 585
R2759 gnd.n2237 gnd.n2236 585
R2760 gnd.n2230 gnd.n2156 585
R2761 gnd.n2232 gnd.n2231 585
R2762 gnd.n2229 gnd.n2228 585
R2763 gnd.n2227 gnd.n2226 585
R2764 gnd.n2220 gnd.n2158 585
R2765 gnd.n2222 gnd.n2221 585
R2766 gnd.n2219 gnd.n2218 585
R2767 gnd.n2217 gnd.n2216 585
R2768 gnd.n2210 gnd.n2160 585
R2769 gnd.n2212 gnd.n2211 585
R2770 gnd.n2209 gnd.n2208 585
R2771 gnd.n2207 gnd.n2206 585
R2772 gnd.n2200 gnd.n2162 585
R2773 gnd.n2202 gnd.n2201 585
R2774 gnd.n2199 gnd.n2198 585
R2775 gnd.n2197 gnd.n2196 585
R2776 gnd.n2190 gnd.n2166 585
R2777 gnd.n2192 gnd.n2191 585
R2778 gnd.n2189 gnd.n2188 585
R2779 gnd.n2187 gnd.n2186 585
R2780 gnd.n2180 gnd.n2168 585
R2781 gnd.n2182 gnd.n2181 585
R2782 gnd.n2179 gnd.n2178 585
R2783 gnd.n2177 gnd.n2176 585
R2784 gnd.n2172 gnd.n2171 585
R2785 gnd.n2170 gnd.n1406 585
R2786 gnd.n3871 gnd.n3870 585
R2787 gnd.n3873 gnd.n3872 585
R2788 gnd.n3875 gnd.n3874 585
R2789 gnd.n3877 gnd.n3876 585
R2790 gnd.n3879 gnd.n3878 585
R2791 gnd.n3881 gnd.n3880 585
R2792 gnd.n3883 gnd.n3882 585
R2793 gnd.n3885 gnd.n3884 585
R2794 gnd.n3888 gnd.n3887 585
R2795 gnd.n3890 gnd.n3889 585
R2796 gnd.n3892 gnd.n3891 585
R2797 gnd.n3894 gnd.n3893 585
R2798 gnd.n3896 gnd.n3895 585
R2799 gnd.n3898 gnd.n3897 585
R2800 gnd.n3900 gnd.n3899 585
R2801 gnd.n3902 gnd.n3901 585
R2802 gnd.n3904 gnd.n3903 585
R2803 gnd.n3906 gnd.n3905 585
R2804 gnd.n3908 gnd.n3907 585
R2805 gnd.n3910 gnd.n3909 585
R2806 gnd.n3912 gnd.n3911 585
R2807 gnd.n3914 gnd.n3913 585
R2808 gnd.n3915 gnd.n1379 585
R2809 gnd.n3917 gnd.n3916 585
R2810 gnd.n1338 gnd.n1337 585
R2811 gnd.n3921 gnd.n3920 585
R2812 gnd.n3920 gnd.n3919 585
R2813 gnd.n2510 gnd.n2248 585
R2814 gnd.n2567 gnd.n2248 585
R2815 gnd.n2511 gnd.n1330 585
R2816 gnd.n3927 gnd.n1330 585
R2817 gnd.n2513 gnd.n2512 585
R2818 gnd.n2535 gnd.n2513 585
R2819 gnd.n2508 gnd.n1321 585
R2820 gnd.n3933 gnd.n1321 585
R2821 gnd.n2507 gnd.n2506 585
R2822 gnd.n2506 gnd.n2505 585
R2823 gnd.n2284 gnd.n1310 585
R2824 gnd.n3939 gnd.n1310 585
R2825 gnd.n2495 gnd.n2494 585
R2826 gnd.n2496 gnd.n2495 585
R2827 gnd.n2493 gnd.n1300 585
R2828 gnd.n3945 gnd.n1300 585
R2829 gnd.n2492 gnd.n2491 585
R2830 gnd.n2491 gnd.n1299 585
R2831 gnd.n2489 gnd.n1289 585
R2832 gnd.n3951 gnd.n1289 585
R2833 gnd.n2488 gnd.n2487 585
R2834 gnd.n2487 gnd.n1282 585
R2835 gnd.n2486 gnd.n1280 585
R2836 gnd.n3957 gnd.n1280 585
R2837 gnd.n2485 gnd.n2484 585
R2838 gnd.n2484 gnd.n1272 585
R2839 gnd.n2482 gnd.n1270 585
R2840 gnd.n3963 gnd.n1270 585
R2841 gnd.n2481 gnd.n2480 585
R2842 gnd.n2480 gnd.n1269 585
R2843 gnd.n2479 gnd.n1261 585
R2844 gnd.n3969 gnd.n1261 585
R2845 gnd.n2478 gnd.n2477 585
R2846 gnd.n2477 gnd.n1253 585
R2847 gnd.n2475 gnd.n1251 585
R2848 gnd.n3975 gnd.n1251 585
R2849 gnd.n2474 gnd.n2473 585
R2850 gnd.n2473 gnd.n1244 585
R2851 gnd.n2472 gnd.n1242 585
R2852 gnd.n3981 gnd.n1242 585
R2853 gnd.n2471 gnd.n2470 585
R2854 gnd.n2470 gnd.n1234 585
R2855 gnd.n2468 gnd.n1232 585
R2856 gnd.n3987 gnd.n1232 585
R2857 gnd.n2467 gnd.n2466 585
R2858 gnd.n2466 gnd.n1231 585
R2859 gnd.n2465 gnd.n1223 585
R2860 gnd.n3993 gnd.n1223 585
R2861 gnd.n2464 gnd.n2463 585
R2862 gnd.n2463 gnd.n1222 585
R2863 gnd.n2461 gnd.n1213 585
R2864 gnd.n3999 gnd.n1213 585
R2865 gnd.n2460 gnd.n2459 585
R2866 gnd.n2459 gnd.n1206 585
R2867 gnd.n2458 gnd.n1204 585
R2868 gnd.n4005 gnd.n1204 585
R2869 gnd.n2457 gnd.n2456 585
R2870 gnd.n2456 gnd.n1196 585
R2871 gnd.n2454 gnd.n1194 585
R2872 gnd.n4011 gnd.n1194 585
R2873 gnd.n2453 gnd.n2452 585
R2874 gnd.n2452 gnd.n1193 585
R2875 gnd.n2451 gnd.n1185 585
R2876 gnd.n4017 gnd.n1185 585
R2877 gnd.n2450 gnd.n2449 585
R2878 gnd.n2449 gnd.n1184 585
R2879 gnd.n2447 gnd.n1175 585
R2880 gnd.n4023 gnd.n1175 585
R2881 gnd.n2446 gnd.n2445 585
R2882 gnd.n2445 gnd.n1168 585
R2883 gnd.n2444 gnd.n1166 585
R2884 gnd.n4029 gnd.n1166 585
R2885 gnd.n2443 gnd.n2442 585
R2886 gnd.n2442 gnd.n1159 585
R2887 gnd.n2440 gnd.n1157 585
R2888 gnd.n4035 gnd.n1157 585
R2889 gnd.n2439 gnd.n2438 585
R2890 gnd.n2438 gnd.n1149 585
R2891 gnd.n2437 gnd.n1147 585
R2892 gnd.n4041 gnd.n1147 585
R2893 gnd.n2436 gnd.n2435 585
R2894 gnd.n2435 gnd.n1146 585
R2895 gnd.n2433 gnd.n1137 585
R2896 gnd.n4049 gnd.n1137 585
R2897 gnd.n1136 gnd.n1130 585
R2898 gnd.n1136 gnd.n1061 585
R2899 gnd.n161 gnd.n160 585
R2900 gnd.n164 gnd.n161 585
R2901 gnd.n7071 gnd.n7070 585
R2902 gnd.n7070 gnd.n7069 585
R2903 gnd.n7072 gnd.n155 585
R2904 gnd.n155 gnd.n154 585
R2905 gnd.n7074 gnd.n7073 585
R2906 gnd.n7075 gnd.n7074 585
R2907 gnd.n141 gnd.n140 585
R2908 gnd.n145 gnd.n141 585
R2909 gnd.n7083 gnd.n7082 585
R2910 gnd.n7082 gnd.n7081 585
R2911 gnd.n7084 gnd.n135 585
R2912 gnd.n142 gnd.n135 585
R2913 gnd.n7086 gnd.n7085 585
R2914 gnd.n7087 gnd.n7086 585
R2915 gnd.n123 gnd.n122 585
R2916 gnd.n126 gnd.n123 585
R2917 gnd.n7095 gnd.n7094 585
R2918 gnd.n7094 gnd.n7093 585
R2919 gnd.n7096 gnd.n117 585
R2920 gnd.n117 gnd.n116 585
R2921 gnd.n7098 gnd.n7097 585
R2922 gnd.n7099 gnd.n7098 585
R2923 gnd.n103 gnd.n102 585
R2924 gnd.n107 gnd.n103 585
R2925 gnd.n7107 gnd.n7106 585
R2926 gnd.n7106 gnd.n7105 585
R2927 gnd.n7108 gnd.n97 585
R2928 gnd.n104 gnd.n97 585
R2929 gnd.n7110 gnd.n7109 585
R2930 gnd.n7111 gnd.n7110 585
R2931 gnd.n83 gnd.n82 585
R2932 gnd.n86 gnd.n83 585
R2933 gnd.n7119 gnd.n7118 585
R2934 gnd.n7118 gnd.n7117 585
R2935 gnd.n7120 gnd.n77 585
R2936 gnd.n77 gnd.n74 585
R2937 gnd.n7122 gnd.n7121 585
R2938 gnd.n7123 gnd.n7122 585
R2939 gnd.n78 gnd.n76 585
R2940 gnd.n6696 gnd.n76 585
R2941 gnd.n6685 gnd.n181 585
R2942 gnd.n181 gnd.n171 585
R2943 gnd.n6687 gnd.n6686 585
R2944 gnd.n6688 gnd.n6687 585
R2945 gnd.n182 gnd.n180 585
R2946 gnd.n188 gnd.n180 585
R2947 gnd.n6679 gnd.n6678 585
R2948 gnd.n6678 gnd.n6677 585
R2949 gnd.n185 gnd.n184 585
R2950 gnd.n6668 gnd.n185 585
R2951 gnd.n6652 gnd.n204 585
R2952 gnd.n204 gnd.n194 585
R2953 gnd.n6654 gnd.n6653 585
R2954 gnd.n6655 gnd.n6654 585
R2955 gnd.n205 gnd.n203 585
R2956 gnd.n212 gnd.n203 585
R2957 gnd.n6647 gnd.n6646 585
R2958 gnd.n6646 gnd.n6645 585
R2959 gnd.n208 gnd.n207 585
R2960 gnd.n209 gnd.n208 585
R2961 gnd.n6628 gnd.n6627 585
R2962 gnd.n6629 gnd.n6628 585
R2963 gnd.n225 gnd.n224 585
R2964 gnd.n224 gnd.n221 585
R2965 gnd.n6623 gnd.n6622 585
R2966 gnd.n6622 gnd.n6621 585
R2967 gnd.n228 gnd.n227 585
R2968 gnd.n6610 gnd.n228 585
R2969 gnd.n6588 gnd.n250 585
R2970 gnd.n250 gnd.n239 585
R2971 gnd.n6590 gnd.n6589 585
R2972 gnd.n6591 gnd.n6590 585
R2973 gnd.n251 gnd.n249 585
R2974 gnd.n6569 gnd.n249 585
R2975 gnd.n6583 gnd.n6582 585
R2976 gnd.n6582 gnd.n6581 585
R2977 gnd.n254 gnd.n253 585
R2978 gnd.n6565 gnd.n254 585
R2979 gnd.n280 gnd.n278 585
R2980 gnd.n6339 gnd.n278 585
R2981 gnd.n6555 gnd.n6554 585
R2982 gnd.n6556 gnd.n6555 585
R2983 gnd.n279 gnd.n277 585
R2984 gnd.n6345 gnd.n277 585
R2985 gnd.n6549 gnd.n6548 585
R2986 gnd.n283 gnd.n282 585
R2987 gnd.n6545 gnd.n6544 585
R2988 gnd.n6546 gnd.n6545 585
R2989 gnd.n6543 gnd.n324 585
R2990 gnd.n6542 gnd.n6541 585
R2991 gnd.n6540 gnd.n6539 585
R2992 gnd.n6538 gnd.n6537 585
R2993 gnd.n6536 gnd.n6535 585
R2994 gnd.n6534 gnd.n6533 585
R2995 gnd.n6532 gnd.n6531 585
R2996 gnd.n6530 gnd.n6529 585
R2997 gnd.n6528 gnd.n6527 585
R2998 gnd.n6526 gnd.n6525 585
R2999 gnd.n6524 gnd.n6523 585
R3000 gnd.n6522 gnd.n6521 585
R3001 gnd.n6520 gnd.n6519 585
R3002 gnd.n6518 gnd.n6517 585
R3003 gnd.n6516 gnd.n6515 585
R3004 gnd.n6513 gnd.n6512 585
R3005 gnd.n6511 gnd.n6510 585
R3006 gnd.n6509 gnd.n6508 585
R3007 gnd.n6507 gnd.n6506 585
R3008 gnd.n6505 gnd.n6504 585
R3009 gnd.n6503 gnd.n6502 585
R3010 gnd.n6501 gnd.n6500 585
R3011 gnd.n6499 gnd.n6498 585
R3012 gnd.n6496 gnd.n6495 585
R3013 gnd.n6494 gnd.n6493 585
R3014 gnd.n6492 gnd.n6491 585
R3015 gnd.n6490 gnd.n6489 585
R3016 gnd.n6488 gnd.n6487 585
R3017 gnd.n6486 gnd.n6485 585
R3018 gnd.n6484 gnd.n6483 585
R3019 gnd.n6482 gnd.n6481 585
R3020 gnd.n6480 gnd.n6479 585
R3021 gnd.n6478 gnd.n6477 585
R3022 gnd.n6476 gnd.n6475 585
R3023 gnd.n6474 gnd.n6473 585
R3024 gnd.n6472 gnd.n6471 585
R3025 gnd.n6470 gnd.n6469 585
R3026 gnd.n6468 gnd.n6467 585
R3027 gnd.n6466 gnd.n6465 585
R3028 gnd.n6464 gnd.n6463 585
R3029 gnd.n6462 gnd.n6461 585
R3030 gnd.n6460 gnd.n6459 585
R3031 gnd.n6458 gnd.n6457 585
R3032 gnd.n6456 gnd.n6455 585
R3033 gnd.n6454 gnd.n6453 585
R3034 gnd.n6452 gnd.n6451 585
R3035 gnd.n6450 gnd.n6449 585
R3036 gnd.n6448 gnd.n6447 585
R3037 gnd.n6446 gnd.n6445 585
R3038 gnd.n6444 gnd.n6443 585
R3039 gnd.n6442 gnd.n6441 585
R3040 gnd.n6440 gnd.n6439 585
R3041 gnd.n6438 gnd.n6437 585
R3042 gnd.n500 gnd.n385 585
R3043 gnd.n7062 gnd.n7061 585
R3044 gnd.n6739 gnd.n6738 585
R3045 gnd.n6939 gnd.n6938 585
R3046 gnd.n6941 gnd.n6940 585
R3047 gnd.n6943 gnd.n6942 585
R3048 gnd.n6945 gnd.n6944 585
R3049 gnd.n6947 gnd.n6946 585
R3050 gnd.n6949 gnd.n6948 585
R3051 gnd.n6951 gnd.n6950 585
R3052 gnd.n6953 gnd.n6952 585
R3053 gnd.n6955 gnd.n6954 585
R3054 gnd.n6957 gnd.n6956 585
R3055 gnd.n6959 gnd.n6958 585
R3056 gnd.n6961 gnd.n6960 585
R3057 gnd.n6963 gnd.n6962 585
R3058 gnd.n6965 gnd.n6964 585
R3059 gnd.n6967 gnd.n6966 585
R3060 gnd.n6969 gnd.n6968 585
R3061 gnd.n6971 gnd.n6970 585
R3062 gnd.n6974 gnd.n6973 585
R3063 gnd.n6972 gnd.n6918 585
R3064 gnd.n6979 gnd.n6978 585
R3065 gnd.n6981 gnd.n6980 585
R3066 gnd.n6983 gnd.n6982 585
R3067 gnd.n6985 gnd.n6984 585
R3068 gnd.n6987 gnd.n6986 585
R3069 gnd.n6989 gnd.n6988 585
R3070 gnd.n6991 gnd.n6990 585
R3071 gnd.n6993 gnd.n6992 585
R3072 gnd.n6995 gnd.n6994 585
R3073 gnd.n6997 gnd.n6996 585
R3074 gnd.n6999 gnd.n6998 585
R3075 gnd.n7001 gnd.n7000 585
R3076 gnd.n7003 gnd.n7002 585
R3077 gnd.n7005 gnd.n7004 585
R3078 gnd.n7007 gnd.n7006 585
R3079 gnd.n7009 gnd.n7008 585
R3080 gnd.n7011 gnd.n7010 585
R3081 gnd.n7013 gnd.n7012 585
R3082 gnd.n7015 gnd.n7014 585
R3083 gnd.n7017 gnd.n7016 585
R3084 gnd.n7022 gnd.n7021 585
R3085 gnd.n7024 gnd.n7023 585
R3086 gnd.n7026 gnd.n7025 585
R3087 gnd.n7028 gnd.n7027 585
R3088 gnd.n7030 gnd.n7029 585
R3089 gnd.n7032 gnd.n7031 585
R3090 gnd.n7034 gnd.n7033 585
R3091 gnd.n7036 gnd.n7035 585
R3092 gnd.n7038 gnd.n7037 585
R3093 gnd.n7040 gnd.n7039 585
R3094 gnd.n7042 gnd.n7041 585
R3095 gnd.n7044 gnd.n7043 585
R3096 gnd.n7046 gnd.n7045 585
R3097 gnd.n7048 gnd.n7047 585
R3098 gnd.n7051 gnd.n7050 585
R3099 gnd.n7049 gnd.n6884 585
R3100 gnd.n7055 gnd.n6881 585
R3101 gnd.n7057 gnd.n7056 585
R3102 gnd.n7058 gnd.n7057 585
R3103 gnd.n7060 gnd.n6733 585
R3104 gnd.n7060 gnd.n164 585
R3105 gnd.n6732 gnd.n162 585
R3106 gnd.n7069 gnd.n162 585
R3107 gnd.n6731 gnd.n6730 585
R3108 gnd.n6730 gnd.n154 585
R3109 gnd.n6728 gnd.n152 585
R3110 gnd.n7075 gnd.n152 585
R3111 gnd.n6727 gnd.n6726 585
R3112 gnd.n6726 gnd.n145 585
R3113 gnd.n6725 gnd.n143 585
R3114 gnd.n7081 gnd.n143 585
R3115 gnd.n6724 gnd.n6723 585
R3116 gnd.n6723 gnd.n142 585
R3117 gnd.n6721 gnd.n133 585
R3118 gnd.n7087 gnd.n133 585
R3119 gnd.n6720 gnd.n6719 585
R3120 gnd.n6719 gnd.n126 585
R3121 gnd.n6718 gnd.n124 585
R3122 gnd.n7093 gnd.n124 585
R3123 gnd.n6717 gnd.n6716 585
R3124 gnd.n6716 gnd.n116 585
R3125 gnd.n6714 gnd.n114 585
R3126 gnd.n7099 gnd.n114 585
R3127 gnd.n6713 gnd.n6712 585
R3128 gnd.n6712 gnd.n107 585
R3129 gnd.n6711 gnd.n105 585
R3130 gnd.n7105 gnd.n105 585
R3131 gnd.n6710 gnd.n6709 585
R3132 gnd.n6709 gnd.n104 585
R3133 gnd.n6707 gnd.n95 585
R3134 gnd.n7111 gnd.n95 585
R3135 gnd.n6706 gnd.n6705 585
R3136 gnd.n6705 gnd.n86 585
R3137 gnd.n6704 gnd.n84 585
R3138 gnd.n7117 gnd.n84 585
R3139 gnd.n6703 gnd.n6702 585
R3140 gnd.n6702 gnd.n74 585
R3141 gnd.n167 gnd.n73 585
R3142 gnd.n7123 gnd.n73 585
R3143 gnd.n6695 gnd.n6694 585
R3144 gnd.n6696 gnd.n6695 585
R3145 gnd.n6693 gnd.n172 585
R3146 gnd.n172 gnd.n171 585
R3147 gnd.n177 gnd.n173 585
R3148 gnd.n6688 gnd.n177 585
R3149 gnd.n6672 gnd.n6671 585
R3150 gnd.n6671 gnd.n188 585
R3151 gnd.n6673 gnd.n186 585
R3152 gnd.n6677 gnd.n186 585
R3153 gnd.n6670 gnd.n6669 585
R3154 gnd.n6669 gnd.n6668 585
R3155 gnd.n193 gnd.n192 585
R3156 gnd.n194 gnd.n193 585
R3157 gnd.n6636 gnd.n201 585
R3158 gnd.n6655 gnd.n201 585
R3159 gnd.n6635 gnd.n6634 585
R3160 gnd.n6634 gnd.n212 585
R3161 gnd.n6633 gnd.n210 585
R3162 gnd.n6645 gnd.n210 585
R3163 gnd.n6632 gnd.n6631 585
R3164 gnd.n6631 gnd.n209 585
R3165 gnd.n6630 gnd.n218 585
R3166 gnd.n6630 gnd.n6629 585
R3167 gnd.n6614 gnd.n220 585
R3168 gnd.n221 gnd.n220 585
R3169 gnd.n6613 gnd.n230 585
R3170 gnd.n6621 gnd.n230 585
R3171 gnd.n6612 gnd.n6611 585
R3172 gnd.n6611 gnd.n6610 585
R3173 gnd.n238 gnd.n236 585
R3174 gnd.n239 gnd.n238 585
R3175 gnd.n6572 gnd.n247 585
R3176 gnd.n6591 gnd.n247 585
R3177 gnd.n6571 gnd.n6570 585
R3178 gnd.n6570 gnd.n6569 585
R3179 gnd.n6568 gnd.n256 585
R3180 gnd.n6581 gnd.n256 585
R3181 gnd.n6567 gnd.n6566 585
R3182 gnd.n6566 gnd.n6565 585
R3183 gnd.n266 gnd.n264 585
R3184 gnd.n6339 gnd.n266 585
R3185 gnd.n504 gnd.n275 585
R3186 gnd.n6556 gnd.n275 585
R3187 gnd.n503 gnd.n501 585
R3188 gnd.n6345 gnd.n501 585
R3189 gnd.n1007 gnd.n1006 585
R3190 gnd.n1291 gnd.n1007 585
R3191 gnd.n6326 gnd.n6325 585
R3192 gnd.n6325 gnd.n229 585
R3193 gnd.n6329 gnd.n517 585
R3194 gnd.n517 gnd.n516 585
R3195 gnd.n6331 gnd.n6330 585
R3196 gnd.n6331 gnd.n246 585
R3197 gnd.n6332 gnd.n515 585
R3198 gnd.n6332 gnd.n258 585
R3199 gnd.n6334 gnd.n6333 585
R3200 gnd.n6333 gnd.n255 585
R3201 gnd.n6335 gnd.n507 585
R3202 gnd.n507 gnd.n267 585
R3203 gnd.n6337 gnd.n6336 585
R3204 gnd.n6338 gnd.n6337 585
R3205 gnd.n508 gnd.n498 585
R3206 gnd.n498 gnd.n274 585
R3207 gnd.n6347 gnd.n499 585
R3208 gnd.n6347 gnd.n6346 585
R3209 gnd.n6348 gnd.n497 585
R3210 gnd.n6348 gnd.n323 585
R3211 gnd.n6350 gnd.n6349 585
R3212 gnd.n6349 gnd.n284 585
R3213 gnd.n6351 gnd.n492 585
R3214 gnd.n492 gnd.n490 585
R3215 gnd.n6353 gnd.n6352 585
R3216 gnd.n6354 gnd.n6353 585
R3217 gnd.n493 gnd.n491 585
R3218 gnd.n491 gnd.n470 585
R3219 gnd.n3670 gnd.n3669 585
R3220 gnd.n3669 gnd.n458 585
R3221 gnd.n3671 gnd.n1577 585
R3222 gnd.n1577 gnd.n457 585
R3223 gnd.n3673 gnd.n3672 585
R3224 gnd.n3674 gnd.n3673 585
R3225 gnd.n1578 gnd.n1576 585
R3226 gnd.n1576 gnd.n1573 585
R3227 gnd.n3662 gnd.n3661 585
R3228 gnd.n3661 gnd.n3660 585
R3229 gnd.n1581 gnd.n1580 585
R3230 gnd.n3648 gnd.n1581 585
R3231 gnd.n3646 gnd.n3645 585
R3232 gnd.n3647 gnd.n3646 585
R3233 gnd.n1591 gnd.n1590 585
R3234 gnd.n3637 gnd.n1590 585
R3235 gnd.n3641 gnd.n3640 585
R3236 gnd.n3640 gnd.n3639 585
R3237 gnd.n1594 gnd.n1593 585
R3238 gnd.n3627 gnd.n1594 585
R3239 gnd.n3625 gnd.n3624 585
R3240 gnd.n3626 gnd.n3625 585
R3241 gnd.n1603 gnd.n1602 585
R3242 gnd.n3616 gnd.n1602 585
R3243 gnd.n3620 gnd.n3619 585
R3244 gnd.n3619 gnd.n3618 585
R3245 gnd.n1606 gnd.n1605 585
R3246 gnd.n3606 gnd.n1606 585
R3247 gnd.n3604 gnd.n3603 585
R3248 gnd.n3605 gnd.n3604 585
R3249 gnd.n1615 gnd.n1614 585
R3250 gnd.n3595 gnd.n1614 585
R3251 gnd.n3599 gnd.n3598 585
R3252 gnd.n3598 gnd.n3597 585
R3253 gnd.n1618 gnd.n1617 585
R3254 gnd.n3585 gnd.n1618 585
R3255 gnd.n3582 gnd.n3581 585
R3256 gnd.n3583 gnd.n3582 585
R3257 gnd.n1626 gnd.n1625 585
R3258 gnd.n3573 gnd.n1625 585
R3259 gnd.n3577 gnd.n3576 585
R3260 gnd.n3576 gnd.n3575 585
R3261 gnd.n1629 gnd.n1628 585
R3262 gnd.n3563 gnd.n1629 585
R3263 gnd.n3396 gnd.n3395 585
R3264 gnd.n3395 gnd.n1636 585
R3265 gnd.n3397 gnd.n1686 585
R3266 gnd.n1686 gnd.n1675 585
R3267 gnd.n3399 gnd.n3398 585
R3268 gnd.n3400 gnd.n3399 585
R3269 gnd.n1687 gnd.n1685 585
R3270 gnd.n1693 gnd.n1685 585
R3271 gnd.n3389 gnd.n3388 585
R3272 gnd.n3388 gnd.n3387 585
R3273 gnd.n1690 gnd.n1689 585
R3274 gnd.n1698 gnd.n1690 585
R3275 gnd.n3343 gnd.n1713 585
R3276 gnd.n1713 gnd.n1703 585
R3277 gnd.n3345 gnd.n3344 585
R3278 gnd.n3346 gnd.n3345 585
R3279 gnd.n1714 gnd.n1712 585
R3280 gnd.n3311 gnd.n1712 585
R3281 gnd.n3338 gnd.n3337 585
R3282 gnd.n3337 gnd.n3336 585
R3283 gnd.n1717 gnd.n1716 585
R3284 gnd.n3319 gnd.n1717 585
R3285 gnd.n3278 gnd.n3277 585
R3286 gnd.n3277 gnd.n1728 585
R3287 gnd.n3279 gnd.n1749 585
R3288 gnd.n1749 gnd.n1737 585
R3289 gnd.n3281 gnd.n3280 585
R3290 gnd.n3282 gnd.n3281 585
R3291 gnd.n1750 gnd.n1748 585
R3292 gnd.n1748 gnd.n1745 585
R3293 gnd.n3271 gnd.n3270 585
R3294 gnd.n3270 gnd.n3269 585
R3295 gnd.n1753 gnd.n1752 585
R3296 gnd.n1759 gnd.n1753 585
R3297 gnd.n3249 gnd.n3248 585
R3298 gnd.n3250 gnd.n3249 585
R3299 gnd.n1768 gnd.n1767 585
R3300 gnd.n1775 gnd.n1767 585
R3301 gnd.n3244 gnd.n3243 585
R3302 gnd.n3243 gnd.n3242 585
R3303 gnd.n1771 gnd.n1770 585
R3304 gnd.n1779 gnd.n1771 585
R3305 gnd.n3202 gnd.n3201 585
R3306 gnd.n3203 gnd.n3202 585
R3307 gnd.n1790 gnd.n1789 585
R3308 gnd.n1808 gnd.n1789 585
R3309 gnd.n3197 gnd.n3196 585
R3310 gnd.n3196 gnd.n3195 585
R3311 gnd.n1793 gnd.n1792 585
R3312 gnd.n1801 gnd.n1793 585
R3313 gnd.n3162 gnd.n3161 585
R3314 gnd.n3163 gnd.n3162 585
R3315 gnd.n1813 gnd.n1812 585
R3316 gnd.n1831 gnd.n1812 585
R3317 gnd.n3157 gnd.n3156 585
R3318 gnd.n3156 gnd.n3155 585
R3319 gnd.n1816 gnd.n1815 585
R3320 gnd.n1824 gnd.n1816 585
R3321 gnd.n3122 gnd.n3121 585
R3322 gnd.n3123 gnd.n3122 585
R3323 gnd.n1836 gnd.n1835 585
R3324 gnd.n3094 gnd.n1835 585
R3325 gnd.n3117 gnd.n3116 585
R3326 gnd.n3116 gnd.n3115 585
R3327 gnd.n1839 gnd.n1838 585
R3328 gnd.n3104 gnd.n1839 585
R3329 gnd.n3066 gnd.n3065 585
R3330 gnd.n3067 gnd.n3066 585
R3331 gnd.n1864 gnd.n1863 585
R3332 gnd.n1863 gnd.n1855 585
R3333 gnd.n3061 gnd.n3060 585
R3334 gnd.n3060 gnd.n1860 585
R3335 gnd.n3059 gnd.n1866 585
R3336 gnd.n3059 gnd.n3058 585
R3337 gnd.n3038 gnd.n1867 585
R3338 gnd.n1873 gnd.n1867 585
R3339 gnd.n3040 gnd.n3039 585
R3340 gnd.n3041 gnd.n3040 585
R3341 gnd.n1883 gnd.n1882 585
R3342 gnd.n2841 gnd.n1882 585
R3343 gnd.n3033 gnd.n3032 585
R3344 gnd.n3032 gnd.n3031 585
R3345 gnd.n1886 gnd.n1885 585
R3346 gnd.n1894 gnd.n1886 585
R3347 gnd.n2987 gnd.n1912 585
R3348 gnd.n1912 gnd.n1905 585
R3349 gnd.n2989 gnd.n2988 585
R3350 gnd.n2990 gnd.n2989 585
R3351 gnd.n1913 gnd.n1911 585
R3352 gnd.n1911 gnd.n1909 585
R3353 gnd.n2982 gnd.n2981 585
R3354 gnd.n2981 gnd.n2980 585
R3355 gnd.n1916 gnd.n1915 585
R3356 gnd.n2972 gnd.n1916 585
R3357 gnd.n2957 gnd.n2956 585
R3358 gnd.n2958 gnd.n2957 585
R3359 gnd.n1934 gnd.n1933 585
R3360 gnd.n1940 gnd.n1933 585
R3361 gnd.n2952 gnd.n2951 585
R3362 gnd.n2951 gnd.n2950 585
R3363 gnd.n1937 gnd.n1936 585
R3364 gnd.n2872 gnd.n1937 585
R3365 gnd.n2920 gnd.n1960 585
R3366 gnd.n1960 gnd.n1953 585
R3367 gnd.n2922 gnd.n2921 585
R3368 gnd.n2923 gnd.n2922 585
R3369 gnd.n1961 gnd.n1959 585
R3370 gnd.n2880 gnd.n1959 585
R3371 gnd.n2915 gnd.n2914 585
R3372 gnd.n2914 gnd.n2913 585
R3373 gnd.n1964 gnd.n1963 585
R3374 gnd.n2905 gnd.n1964 585
R3375 gnd.n2752 gnd.n2748 585
R3376 gnd.n2748 gnd.n1474 585
R3377 gnd.n2754 gnd.n2753 585
R3378 gnd.n2754 gnd.n1471 585
R3379 gnd.n2755 gnd.n2747 585
R3380 gnd.n2755 gnd.n1445 585
R3381 gnd.n2758 gnd.n2757 585
R3382 gnd.n2757 gnd.n2756 585
R3383 gnd.n2759 gnd.n1991 585
R3384 gnd.n1991 gnd.n1979 585
R3385 gnd.n2761 gnd.n2760 585
R3386 gnd.n2762 gnd.n2761 585
R3387 gnd.n1992 gnd.n1990 585
R3388 gnd.n1990 gnd.n1987 585
R3389 gnd.n2741 gnd.n2740 585
R3390 gnd.n2740 gnd.n2739 585
R3391 gnd.n1995 gnd.n1994 585
R3392 gnd.n2004 gnd.n1995 585
R3393 gnd.n2712 gnd.n2016 585
R3394 gnd.n2016 gnd.n2003 585
R3395 gnd.n2714 gnd.n2713 585
R3396 gnd.n2715 gnd.n2714 585
R3397 gnd.n2017 gnd.n2015 585
R3398 gnd.n2015 gnd.n2012 585
R3399 gnd.n2707 gnd.n2706 585
R3400 gnd.n2706 gnd.n2705 585
R3401 gnd.n2020 gnd.n2019 585
R3402 gnd.n2028 gnd.n2020 585
R3403 gnd.n2682 gnd.n2041 585
R3404 gnd.n2041 gnd.n2027 585
R3405 gnd.n2684 gnd.n2683 585
R3406 gnd.n2685 gnd.n2684 585
R3407 gnd.n2042 gnd.n2040 585
R3408 gnd.n2040 gnd.n2037 585
R3409 gnd.n2677 gnd.n2676 585
R3410 gnd.n2676 gnd.n2675 585
R3411 gnd.n2045 gnd.n2044 585
R3412 gnd.n2054 gnd.n2045 585
R3413 gnd.n2652 gnd.n2066 585
R3414 gnd.n2066 gnd.n2053 585
R3415 gnd.n2654 gnd.n2653 585
R3416 gnd.n2655 gnd.n2654 585
R3417 gnd.n2067 gnd.n2065 585
R3418 gnd.n2065 gnd.n2062 585
R3419 gnd.n2647 gnd.n2646 585
R3420 gnd.n2646 gnd.n2645 585
R3421 gnd.n2070 gnd.n2069 585
R3422 gnd.n2078 gnd.n2070 585
R3423 gnd.n2552 gnd.n2546 585
R3424 gnd.n2546 gnd.n2077 585
R3425 gnd.n2554 gnd.n2553 585
R3426 gnd.n2555 gnd.n2554 585
R3427 gnd.n2547 gnd.n2256 585
R3428 gnd.n2558 gnd.n2256 585
R3429 gnd.n2560 gnd.n2255 585
R3430 gnd.n2560 gnd.n2559 585
R3431 gnd.n2562 gnd.n2561 585
R3432 gnd.n2561 gnd.n1350 585
R3433 gnd.n2563 gnd.n2250 585
R3434 gnd.n2250 gnd.n1339 585
R3435 gnd.n2565 gnd.n2564 585
R3436 gnd.n2566 gnd.n2565 585
R3437 gnd.n2251 gnd.n2249 585
R3438 gnd.n2249 gnd.n1332 585
R3439 gnd.n2533 gnd.n2532 585
R3440 gnd.n2534 gnd.n2533 585
R3441 gnd.n2515 gnd.n2514 585
R3442 gnd.n2514 gnd.n1323 585
R3443 gnd.n2527 gnd.n2526 585
R3444 gnd.n2526 gnd.n1320 585
R3445 gnd.n2525 gnd.n2517 585
R3446 gnd.n2525 gnd.n1312 585
R3447 gnd.n2524 gnd.n2523 585
R3448 gnd.n2524 gnd.n1309 585
R3449 gnd.n2519 gnd.n2518 585
R3450 gnd.n2518 gnd.n1302 585
R3451 gnd.n6370 gnd.n6369 585
R3452 gnd.n6371 gnd.n6370 585
R3453 gnd.n461 gnd.n459 585
R3454 gnd.n1575 gnd.n459 585
R3455 gnd.n3678 gnd.n3676 585
R3456 gnd.n3676 gnd.n3675 585
R3457 gnd.n3679 gnd.n1572 585
R3458 gnd.n3659 gnd.n1572 585
R3459 gnd.n3680 gnd.n1571 585
R3460 gnd.n1582 gnd.n1571 585
R3461 gnd.n3649 gnd.n1569 585
R3462 gnd.n3650 gnd.n3649 585
R3463 gnd.n3684 gnd.n1568 585
R3464 gnd.n1589 gnd.n1568 585
R3465 gnd.n3685 gnd.n1567 585
R3466 gnd.n3638 gnd.n1567 585
R3467 gnd.n3686 gnd.n1566 585
R3468 gnd.n1595 gnd.n1566 585
R3469 gnd.n3628 gnd.n1564 585
R3470 gnd.n3629 gnd.n3628 585
R3471 gnd.n3690 gnd.n1563 585
R3472 gnd.n1601 gnd.n1563 585
R3473 gnd.n3691 gnd.n1562 585
R3474 gnd.n3617 gnd.n1562 585
R3475 gnd.n3692 gnd.n1561 585
R3476 gnd.n1607 gnd.n1561 585
R3477 gnd.n3607 gnd.n1559 585
R3478 gnd.n3608 gnd.n3607 585
R3479 gnd.n3696 gnd.n1558 585
R3480 gnd.n1613 gnd.n1558 585
R3481 gnd.n3697 gnd.n1557 585
R3482 gnd.n3596 gnd.n1557 585
R3483 gnd.n3698 gnd.n1556 585
R3484 gnd.n3584 gnd.n1556 585
R3485 gnd.n3586 gnd.n1554 585
R3486 gnd.n3587 gnd.n3586 585
R3487 gnd.n3702 gnd.n1553 585
R3488 gnd.n1624 gnd.n1553 585
R3489 gnd.n3703 gnd.n1552 585
R3490 gnd.n3574 gnd.n1552 585
R3491 gnd.n3704 gnd.n1551 585
R3492 gnd.n1630 gnd.n1551 585
R3493 gnd.n3564 gnd.n1549 585
R3494 gnd.n3565 gnd.n3564 585
R3495 gnd.n3708 gnd.n1548 585
R3496 gnd.n1676 gnd.n1548 585
R3497 gnd.n3709 gnd.n1547 585
R3498 gnd.n1684 gnd.n1547 585
R3499 gnd.n3710 gnd.n1546 585
R3500 gnd.n1681 gnd.n1546 585
R3501 gnd.n1694 gnd.n1544 585
R3502 gnd.n3386 gnd.n1694 585
R3503 gnd.n3714 gnd.n1543 585
R3504 gnd.n3379 gnd.n1543 585
R3505 gnd.n3715 gnd.n1542 585
R3506 gnd.n3365 gnd.n1542 585
R3507 gnd.n3716 gnd.n1541 585
R3508 gnd.n3326 gnd.n1541 585
R3509 gnd.n3347 gnd.n1539 585
R3510 gnd.n3348 gnd.n3347 585
R3511 gnd.n3720 gnd.n1538 585
R3512 gnd.n1720 gnd.n1538 585
R3513 gnd.n3721 gnd.n1537 585
R3514 gnd.n1718 gnd.n1537 585
R3515 gnd.n3722 gnd.n1536 585
R3516 gnd.n3302 gnd.n1536 585
R3517 gnd.n1739 gnd.n1534 585
R3518 gnd.n1740 gnd.n1739 585
R3519 gnd.n3726 gnd.n1533 585
R3520 gnd.n3293 gnd.n1533 585
R3521 gnd.n3727 gnd.n1532 585
R3522 gnd.n3284 gnd.n1532 585
R3523 gnd.n3728 gnd.n1531 585
R3524 gnd.n3268 gnd.n1531 585
R3525 gnd.n1760 gnd.n1529 585
R3526 gnd.n1761 gnd.n1760 585
R3527 gnd.n3732 gnd.n1528 585
R3528 gnd.n3218 gnd.n1528 585
R3529 gnd.n3733 gnd.n1527 585
R3530 gnd.n3215 gnd.n1527 585
R3531 gnd.n3734 gnd.n1526 585
R3532 gnd.n3241 gnd.n1526 585
R3533 gnd.n3232 gnd.n1524 585
R3534 gnd.n3233 gnd.n3232 585
R3535 gnd.n3738 gnd.n1523 585
R3536 gnd.n3204 gnd.n1523 585
R3537 gnd.n3739 gnd.n1522 585
R3538 gnd.n3175 gnd.n1522 585
R3539 gnd.n3740 gnd.n1521 585
R3540 gnd.n1796 gnd.n1521 585
R3541 gnd.n3183 gnd.n1519 585
R3542 gnd.n3184 gnd.n3183 585
R3543 gnd.n3744 gnd.n1518 585
R3544 gnd.n3164 gnd.n1518 585
R3545 gnd.n3745 gnd.n1517 585
R3546 gnd.n3135 gnd.n1517 585
R3547 gnd.n3746 gnd.n1516 585
R3548 gnd.n1819 gnd.n1516 585
R3549 gnd.n3143 gnd.n1514 585
R3550 gnd.n3144 gnd.n3143 585
R3551 gnd.n3750 gnd.n1513 585
R3552 gnd.n3124 gnd.n1513 585
R3553 gnd.n3751 gnd.n1512 585
R3554 gnd.n3093 gnd.n1512 585
R3555 gnd.n3752 gnd.n1511 585
R3556 gnd.n1841 gnd.n1511 585
R3557 gnd.n3102 gnd.n1509 585
R3558 gnd.n3103 gnd.n3102 585
R3559 gnd.n3756 gnd.n1508 585
R3560 gnd.n1846 gnd.n1508 585
R3561 gnd.n3757 gnd.n1507 585
R3562 gnd.n3083 gnd.n1507 585
R3563 gnd.n3758 gnd.n1506 585
R3564 gnd.n3075 gnd.n1506 585
R3565 gnd.n3056 gnd.n1504 585
R3566 gnd.n3057 gnd.n3056 585
R3567 gnd.n3762 gnd.n1503 585
R3568 gnd.n1874 gnd.n1503 585
R3569 gnd.n3763 gnd.n1502 585
R3570 gnd.n1881 gnd.n1502 585
R3571 gnd.n3764 gnd.n1501 585
R3572 gnd.n1879 gnd.n1501 585
R3573 gnd.n1889 gnd.n1499 585
R3574 gnd.n1890 gnd.n1889 585
R3575 gnd.n3768 gnd.n1498 585
R3576 gnd.n3023 gnd.n1498 585
R3577 gnd.n3769 gnd.n1497 585
R3578 gnd.n2849 gnd.n1497 585
R3579 gnd.n3770 gnd.n1496 585
R3580 gnd.n3000 gnd.n1496 585
R3581 gnd.n2991 gnd.n1494 585
R3582 gnd.n2992 gnd.n2991 585
R3583 gnd.n3774 gnd.n1493 585
R3584 gnd.n1918 gnd.n1493 585
R3585 gnd.n3775 gnd.n1492 585
R3586 gnd.n2970 gnd.n1492 585
R3587 gnd.n3776 gnd.n1491 585
R3588 gnd.n1922 gnd.n1491 585
R3589 gnd.n2960 gnd.n1489 585
R3590 gnd.n2961 gnd.n2960 585
R3591 gnd.n3780 gnd.n1488 585
R3592 gnd.n2949 gnd.n1488 585
R3593 gnd.n3781 gnd.n1487 585
R3594 gnd.n2940 gnd.n1487 585
R3595 gnd.n3782 gnd.n1486 585
R3596 gnd.n2871 gnd.n1486 585
R3597 gnd.n2931 gnd.n1484 585
R3598 gnd.n2932 gnd.n2931 585
R3599 gnd.n3786 gnd.n1483 585
R3600 gnd.n1957 gnd.n1483 585
R3601 gnd.n3787 gnd.n1482 585
R3602 gnd.n1966 gnd.n1482 585
R3603 gnd.n3788 gnd.n1481 585
R3604 gnd.n2904 gnd.n1481 585
R3605 gnd.n1478 gnd.n1476 585
R3606 gnd.n1968 gnd.n1476 585
R3607 gnd.n3793 gnd.n3792 585
R3608 gnd.n3794 gnd.n3793 585
R3609 gnd.n1477 gnd.n1475 585
R3610 gnd.n2894 gnd.n1475 585
R3611 gnd.n1983 gnd.n1981 585
R3612 gnd.n1981 gnd.n1413 585
R3613 gnd.n2771 gnd.n2770 585
R3614 gnd.n2772 gnd.n2771 585
R3615 gnd.n1982 gnd.n1980 585
R3616 gnd.n1989 gnd.n1980 585
R3617 gnd.n2765 gnd.n2764 585
R3618 gnd.n2764 gnd.n2763 585
R3619 gnd.n1986 gnd.n1985 585
R3620 gnd.n2738 gnd.n1986 585
R3621 gnd.n2008 gnd.n2006 585
R3622 gnd.n2006 gnd.n1996 585
R3623 gnd.n2724 gnd.n2723 585
R3624 gnd.n2725 gnd.n2724 585
R3625 gnd.n2007 gnd.n2005 585
R3626 gnd.n2014 gnd.n2005 585
R3627 gnd.n2718 gnd.n2717 585
R3628 gnd.n2717 gnd.n2716 585
R3629 gnd.n2011 gnd.n2010 585
R3630 gnd.n2704 gnd.n2011 585
R3631 gnd.n2033 gnd.n2031 585
R3632 gnd.n2031 gnd.n2030 585
R3633 gnd.n2694 gnd.n2693 585
R3634 gnd.n2695 gnd.n2694 585
R3635 gnd.n2032 gnd.n2029 585
R3636 gnd.n2039 gnd.n2029 585
R3637 gnd.n2688 gnd.n2687 585
R3638 gnd.n2687 gnd.n2686 585
R3639 gnd.n2036 gnd.n2035 585
R3640 gnd.n2674 gnd.n2036 585
R3641 gnd.n2058 gnd.n2056 585
R3642 gnd.n2056 gnd.n2046 585
R3643 gnd.n2664 gnd.n2663 585
R3644 gnd.n2665 gnd.n2664 585
R3645 gnd.n2057 gnd.n2055 585
R3646 gnd.n2064 gnd.n2055 585
R3647 gnd.n2658 gnd.n2657 585
R3648 gnd.n2657 gnd.n2656 585
R3649 gnd.n2061 gnd.n2060 585
R3650 gnd.n2644 gnd.n2061 585
R3651 gnd.n2081 gnd.n2080 585
R3652 gnd.n2080 gnd.n2071 585
R3653 gnd.n2634 gnd.n2633 585
R3654 gnd.n2635 gnd.n2634 585
R3655 gnd.n2629 gnd.n2079 585
R3656 gnd.n2628 gnd.n2083 585
R3657 gnd.n2627 gnd.n2084 585
R3658 gnd.n2557 gnd.n2084 585
R3659 gnd.n2257 gnd.n2085 585
R3660 gnd.n2623 gnd.n2087 585
R3661 gnd.n2622 gnd.n2088 585
R3662 gnd.n2621 gnd.n2089 585
R3663 gnd.n2260 gnd.n2090 585
R3664 gnd.n2616 gnd.n2093 585
R3665 gnd.n2615 gnd.n2094 585
R3666 gnd.n2262 gnd.n2095 585
R3667 gnd.n2608 gnd.n2103 585
R3668 gnd.n2607 gnd.n2104 585
R3669 gnd.n2265 gnd.n2105 585
R3670 gnd.n2600 gnd.n2111 585
R3671 gnd.n2599 gnd.n2112 585
R3672 gnd.n2267 gnd.n2113 585
R3673 gnd.n2592 gnd.n2121 585
R3674 gnd.n2591 gnd.n2122 585
R3675 gnd.n2270 gnd.n2123 585
R3676 gnd.n2584 gnd.n2129 585
R3677 gnd.n2583 gnd.n2130 585
R3678 gnd.n2272 gnd.n2131 585
R3679 gnd.n2576 gnd.n2139 585
R3680 gnd.n2575 gnd.n2140 585
R3681 gnd.n2278 gnd.n2277 585
R3682 gnd.n2280 gnd.n2276 585
R3683 gnd.n2544 gnd.n2543 585
R3684 gnd.n2281 gnd.n2076 585
R3685 gnd.n6373 gnd.n6372 585
R3686 gnd.n6372 gnd.n6371 585
R3687 gnd.n455 gnd.n454 585
R3688 gnd.n1575 gnd.n455 585
R3689 gnd.n1585 gnd.n1574 585
R3690 gnd.n3675 gnd.n1574 585
R3691 gnd.n3658 gnd.n3657 585
R3692 gnd.n3659 gnd.n3658 585
R3693 gnd.n1584 gnd.n1583 585
R3694 gnd.n1583 gnd.n1582 585
R3695 gnd.n3652 gnd.n3651 585
R3696 gnd.n3651 gnd.n3650 585
R3697 gnd.n1588 gnd.n1587 585
R3698 gnd.n1589 gnd.n1588 585
R3699 gnd.n3636 gnd.n3635 585
R3700 gnd.n3638 gnd.n3636 585
R3701 gnd.n1597 gnd.n1596 585
R3702 gnd.n1596 gnd.n1595 585
R3703 gnd.n3631 gnd.n3630 585
R3704 gnd.n3630 gnd.n3629 585
R3705 gnd.n1600 gnd.n1599 585
R3706 gnd.n1601 gnd.n1600 585
R3707 gnd.n3615 gnd.n3614 585
R3708 gnd.n3617 gnd.n3615 585
R3709 gnd.n1609 gnd.n1608 585
R3710 gnd.n1608 gnd.n1607 585
R3711 gnd.n3610 gnd.n3609 585
R3712 gnd.n3609 gnd.n3608 585
R3713 gnd.n1612 gnd.n1611 585
R3714 gnd.n1613 gnd.n1612 585
R3715 gnd.n3594 gnd.n3593 585
R3716 gnd.n3596 gnd.n3594 585
R3717 gnd.n1620 gnd.n1619 585
R3718 gnd.n3584 gnd.n1619 585
R3719 gnd.n3589 gnd.n3588 585
R3720 gnd.n3588 gnd.n3587 585
R3721 gnd.n1623 gnd.n1622 585
R3722 gnd.n1624 gnd.n1623 585
R3723 gnd.n3572 gnd.n3571 585
R3724 gnd.n3574 gnd.n3572 585
R3725 gnd.n1632 gnd.n1631 585
R3726 gnd.n1631 gnd.n1630 585
R3727 gnd.n3567 gnd.n3566 585
R3728 gnd.n3566 gnd.n3565 585
R3729 gnd.n1635 gnd.n1634 585
R3730 gnd.n1676 gnd.n1635 585
R3731 gnd.n3357 gnd.n3355 585
R3732 gnd.n3355 gnd.n1684 585
R3733 gnd.n3358 gnd.n3354 585
R3734 gnd.n3354 gnd.n1681 585
R3735 gnd.n3359 gnd.n1692 585
R3736 gnd.n3386 gnd.n1692 585
R3737 gnd.n1706 gnd.n1700 585
R3738 gnd.n3379 gnd.n1700 585
R3739 gnd.n3364 gnd.n3363 585
R3740 gnd.n3365 gnd.n3364 585
R3741 gnd.n1705 gnd.n1704 585
R3742 gnd.n3326 gnd.n1704 585
R3743 gnd.n3350 gnd.n3349 585
R3744 gnd.n3349 gnd.n3348 585
R3745 gnd.n1709 gnd.n1708 585
R3746 gnd.n1720 gnd.n1709 585
R3747 gnd.n1732 gnd.n1730 585
R3748 gnd.n1730 gnd.n1718 585
R3749 gnd.n3301 gnd.n3300 585
R3750 gnd.n3302 gnd.n3301 585
R3751 gnd.n1731 gnd.n1729 585
R3752 gnd.n1740 gnd.n1729 585
R3753 gnd.n3295 gnd.n3294 585
R3754 gnd.n3294 gnd.n3293 585
R3755 gnd.n1735 gnd.n1734 585
R3756 gnd.n3284 gnd.n1735 585
R3757 gnd.n3221 gnd.n1755 585
R3758 gnd.n3268 gnd.n1755 585
R3759 gnd.n3224 gnd.n3220 585
R3760 gnd.n3220 gnd.n1761 585
R3761 gnd.n3225 gnd.n3219 585
R3762 gnd.n3219 gnd.n3218 585
R3763 gnd.n3226 gnd.n3216 585
R3764 gnd.n3216 gnd.n3215 585
R3765 gnd.n1783 gnd.n1773 585
R3766 gnd.n3241 gnd.n1773 585
R3767 gnd.n3231 gnd.n3230 585
R3768 gnd.n3233 gnd.n3231 585
R3769 gnd.n1782 gnd.n1781 585
R3770 gnd.n3204 gnd.n1781 585
R3771 gnd.n3177 gnd.n3176 585
R3772 gnd.n3176 gnd.n3175 585
R3773 gnd.n1806 gnd.n1804 585
R3774 gnd.n1804 gnd.n1796 585
R3775 gnd.n3182 gnd.n3181 585
R3776 gnd.n3184 gnd.n3182 585
R3777 gnd.n1805 gnd.n1803 585
R3778 gnd.n3164 gnd.n1803 585
R3779 gnd.n3137 gnd.n3136 585
R3780 gnd.n3136 gnd.n3135 585
R3781 gnd.n1829 gnd.n1827 585
R3782 gnd.n1827 gnd.n1819 585
R3783 gnd.n3142 gnd.n3141 585
R3784 gnd.n3144 gnd.n3142 585
R3785 gnd.n1828 gnd.n1826 585
R3786 gnd.n3124 gnd.n1826 585
R3787 gnd.n3092 gnd.n3091 585
R3788 gnd.n3093 gnd.n3092 585
R3789 gnd.n1851 gnd.n1850 585
R3790 gnd.n1850 gnd.n1841 585
R3791 gnd.n3087 gnd.n1848 585
R3792 gnd.n3103 gnd.n1848 585
R3793 gnd.n3086 gnd.n3085 585
R3794 gnd.n3085 gnd.n1846 585
R3795 gnd.n3084 gnd.n1853 585
R3796 gnd.n3084 gnd.n3083 585
R3797 gnd.n3011 gnd.n1854 585
R3798 gnd.n3075 gnd.n1854 585
R3799 gnd.n3009 gnd.n1869 585
R3800 gnd.n3057 gnd.n1869 585
R3801 gnd.n3015 gnd.n3008 585
R3802 gnd.n3008 gnd.n1874 585
R3803 gnd.n3016 gnd.n3007 585
R3804 gnd.n3007 gnd.n1881 585
R3805 gnd.n3017 gnd.n3006 585
R3806 gnd.n3006 gnd.n1879 585
R3807 gnd.n1899 gnd.n1897 585
R3808 gnd.n1897 gnd.n1890 585
R3809 gnd.n3022 gnd.n3021 585
R3810 gnd.n3023 gnd.n3022 585
R3811 gnd.n1898 gnd.n1896 585
R3812 gnd.n2849 gnd.n1896 585
R3813 gnd.n3002 gnd.n3001 585
R3814 gnd.n3001 gnd.n3000 585
R3815 gnd.n1902 gnd.n1901 585
R3816 gnd.n2992 gnd.n1902 585
R3817 gnd.n1928 gnd.n1926 585
R3818 gnd.n1926 gnd.n1918 585
R3819 gnd.n2969 gnd.n2968 585
R3820 gnd.n2970 gnd.n2969 585
R3821 gnd.n1927 gnd.n1925 585
R3822 gnd.n1925 gnd.n1922 585
R3823 gnd.n2963 gnd.n2962 585
R3824 gnd.n2962 gnd.n2961 585
R3825 gnd.n1931 gnd.n1930 585
R3826 gnd.n2949 gnd.n1931 585
R3827 gnd.n2939 gnd.n2938 585
R3828 gnd.n2940 gnd.n2939 585
R3829 gnd.n1947 gnd.n1946 585
R3830 gnd.n2871 gnd.n1946 585
R3831 gnd.n2934 gnd.n2933 585
R3832 gnd.n2933 gnd.n2932 585
R3833 gnd.n1950 gnd.n1949 585
R3834 gnd.n1957 gnd.n1950 585
R3835 gnd.n1974 gnd.n1972 585
R3836 gnd.n1972 gnd.n1966 585
R3837 gnd.n2903 gnd.n2902 585
R3838 gnd.n2904 gnd.n2903 585
R3839 gnd.n1973 gnd.n1971 585
R3840 gnd.n1971 gnd.n1968 585
R3841 gnd.n2897 gnd.n1473 585
R3842 gnd.n3794 gnd.n1473 585
R3843 gnd.n2896 gnd.n2895 585
R3844 gnd.n2895 gnd.n2894 585
R3845 gnd.n2774 gnd.n1976 585
R3846 gnd.n2774 gnd.n1413 585
R3847 gnd.n2773 gnd.n1978 585
R3848 gnd.n2773 gnd.n2772 585
R3849 gnd.n2732 gnd.n1977 585
R3850 gnd.n1989 gnd.n1977 585
R3851 gnd.n1999 gnd.n1988 585
R3852 gnd.n2763 gnd.n1988 585
R3853 gnd.n2737 gnd.n2736 585
R3854 gnd.n2738 gnd.n2737 585
R3855 gnd.n1998 gnd.n1997 585
R3856 gnd.n1997 gnd.n1996 585
R3857 gnd.n2727 gnd.n2726 585
R3858 gnd.n2726 gnd.n2725 585
R3859 gnd.n2002 gnd.n2001 585
R3860 gnd.n2014 gnd.n2002 585
R3861 gnd.n2023 gnd.n2013 585
R3862 gnd.n2716 gnd.n2013 585
R3863 gnd.n2703 gnd.n2702 585
R3864 gnd.n2704 gnd.n2703 585
R3865 gnd.n2022 gnd.n2021 585
R3866 gnd.n2030 gnd.n2021 585
R3867 gnd.n2697 gnd.n2696 585
R3868 gnd.n2696 gnd.n2695 585
R3869 gnd.n2026 gnd.n2025 585
R3870 gnd.n2039 gnd.n2026 585
R3871 gnd.n2049 gnd.n2038 585
R3872 gnd.n2686 gnd.n2038 585
R3873 gnd.n2673 gnd.n2672 585
R3874 gnd.n2674 gnd.n2673 585
R3875 gnd.n2048 gnd.n2047 585
R3876 gnd.n2047 gnd.n2046 585
R3877 gnd.n2667 gnd.n2666 585
R3878 gnd.n2666 gnd.n2665 585
R3879 gnd.n2052 gnd.n2051 585
R3880 gnd.n2064 gnd.n2052 585
R3881 gnd.n2074 gnd.n2063 585
R3882 gnd.n2656 gnd.n2063 585
R3883 gnd.n2643 gnd.n2642 585
R3884 gnd.n2644 gnd.n2643 585
R3885 gnd.n2073 gnd.n2072 585
R3886 gnd.n2072 gnd.n2071 585
R3887 gnd.n2637 gnd.n2636 585
R3888 gnd.n2636 gnd.n2635 585
R3889 gnd.n6389 gnd.n440 585
R3890 gnd.n6355 gnd.n440 585
R3891 gnd.n6390 gnd.n439 585
R3892 gnd.n485 gnd.n433 585
R3893 gnd.n6397 gnd.n432 585
R3894 gnd.n6398 gnd.n431 585
R3895 gnd.n482 gnd.n423 585
R3896 gnd.n6405 gnd.n422 585
R3897 gnd.n6406 gnd.n421 585
R3898 gnd.n480 gnd.n415 585
R3899 gnd.n6413 gnd.n414 585
R3900 gnd.n6414 gnd.n413 585
R3901 gnd.n477 gnd.n405 585
R3902 gnd.n6421 gnd.n404 585
R3903 gnd.n6422 gnd.n403 585
R3904 gnd.n475 gnd.n395 585
R3905 gnd.n6429 gnd.n394 585
R3906 gnd.n6430 gnd.n393 585
R3907 gnd.n6431 gnd.n392 585
R3908 gnd.n6357 gnd.n391 585
R3909 gnd.n6359 gnd.n6358 585
R3910 gnd.n6360 gnd.n468 585
R3911 gnd.n472 gnd.n466 585
R3912 gnd.n6364 gnd.n465 585
R3913 gnd.n6365 gnd.n464 585
R3914 gnd.n6366 gnd.n460 585
R3915 gnd.n456 gnd.n452 585
R3916 gnd.n6378 gnd.n451 585
R3917 gnd.n6379 gnd.n450 585
R3918 gnd.n487 gnd.n449 585
R3919 gnd.n3493 gnd.n1678 473.281
R3920 gnd.n3496 gnd.n3495 473.281
R3921 gnd.n2892 gnd.n2775 473.281
R3922 gnd.n3863 gnd.n1448 473.281
R3923 gnd.n2776 gnd.t155 443.966
R3924 gnd.n1671 gnd.t90 443.966
R3925 gnd.n3800 gnd.t83 443.966
R3926 gnd.n3424 gnd.t146 443.966
R3927 gnd.n2141 gnd.t105 371.625
R3928 gnd.n6383 gnd.t65 371.625
R3929 gnd.n6736 gnd.t118 371.625
R3930 gnd.n6919 gnd.t128 371.625
R3931 gnd.n7018 gnd.t140 371.625
R3932 gnd.n341 gnd.t158 371.625
R3933 gnd.n364 gnd.t164 371.625
R3934 gnd.n386 gnd.t121 371.625
R3935 gnd.n6751 gnd.t61 371.625
R3936 gnd.n2146 gnd.t98 371.625
R3937 gnd.n2311 gnd.t94 371.625
R3938 gnd.n1083 gnd.t109 371.625
R3939 gnd.n1105 gnd.t143 371.625
R3940 gnd.n1127 gnd.t149 371.625
R3941 gnd.n1396 gnd.t134 371.625
R3942 gnd.n2152 gnd.t152 371.625
R3943 gnd.n2164 gnd.t171 371.625
R3944 gnd.n441 gnd.t72 371.625
R3945 gnd.n5790 gnd.n5789 348.315
R3946 gnd.n4640 gnd.t124 323.425
R3947 gnd.n4198 gnd.t177 323.425
R3948 gnd.n5488 gnd.n5462 289.615
R3949 gnd.n5456 gnd.n5430 289.615
R3950 gnd.n5424 gnd.n5398 289.615
R3951 gnd.n5393 gnd.n5367 289.615
R3952 gnd.n5361 gnd.n5335 289.615
R3953 gnd.n5329 gnd.n5303 289.615
R3954 gnd.n5297 gnd.n5271 289.615
R3955 gnd.n5266 gnd.n5240 289.615
R3956 gnd.n4714 gnd.t167 279.217
R3957 gnd.n4224 gnd.t76 279.217
R3958 gnd.n1455 gnd.t82 260.649
R3959 gnd.n3416 gnd.t114 260.649
R3960 gnd.n3865 gnd.n3864 256.663
R3961 gnd.n3865 gnd.n1414 256.663
R3962 gnd.n3865 gnd.n1415 256.663
R3963 gnd.n3865 gnd.n1416 256.663
R3964 gnd.n3865 gnd.n1417 256.663
R3965 gnd.n3865 gnd.n1418 256.663
R3966 gnd.n3865 gnd.n1419 256.663
R3967 gnd.n3865 gnd.n1420 256.663
R3968 gnd.n3865 gnd.n1421 256.663
R3969 gnd.n3865 gnd.n1422 256.663
R3970 gnd.n3865 gnd.n1423 256.663
R3971 gnd.n3865 gnd.n1424 256.663
R3972 gnd.n3865 gnd.n1425 256.663
R3973 gnd.n3865 gnd.n1426 256.663
R3974 gnd.n3865 gnd.n1427 256.663
R3975 gnd.n3865 gnd.n1428 256.663
R3976 gnd.n3868 gnd.n1411 256.663
R3977 gnd.n3866 gnd.n3865 256.663
R3978 gnd.n3865 gnd.n1429 256.663
R3979 gnd.n3865 gnd.n1430 256.663
R3980 gnd.n3865 gnd.n1431 256.663
R3981 gnd.n3865 gnd.n1432 256.663
R3982 gnd.n3865 gnd.n1433 256.663
R3983 gnd.n3865 gnd.n1434 256.663
R3984 gnd.n3865 gnd.n1435 256.663
R3985 gnd.n3865 gnd.n1436 256.663
R3986 gnd.n3865 gnd.n1437 256.663
R3987 gnd.n3865 gnd.n1438 256.663
R3988 gnd.n3865 gnd.n1439 256.663
R3989 gnd.n3865 gnd.n1440 256.663
R3990 gnd.n3865 gnd.n1441 256.663
R3991 gnd.n3865 gnd.n1442 256.663
R3992 gnd.n3865 gnd.n1443 256.663
R3993 gnd.n3865 gnd.n1444 256.663
R3994 gnd.n3562 gnd.n1654 256.663
R3995 gnd.n3562 gnd.n1655 256.663
R3996 gnd.n3562 gnd.n1656 256.663
R3997 gnd.n3562 gnd.n1657 256.663
R3998 gnd.n3562 gnd.n1658 256.663
R3999 gnd.n3562 gnd.n1659 256.663
R4000 gnd.n3562 gnd.n1660 256.663
R4001 gnd.n3562 gnd.n1661 256.663
R4002 gnd.n3562 gnd.n1662 256.663
R4003 gnd.n3562 gnd.n1663 256.663
R4004 gnd.n3562 gnd.n1664 256.663
R4005 gnd.n3562 gnd.n1665 256.663
R4006 gnd.n3562 gnd.n1666 256.663
R4007 gnd.n3562 gnd.n1667 256.663
R4008 gnd.n3562 gnd.n1668 256.663
R4009 gnd.n3562 gnd.n1669 256.663
R4010 gnd.n1670 gnd.n351 256.663
R4011 gnd.n3562 gnd.n1653 256.663
R4012 gnd.n3562 gnd.n1652 256.663
R4013 gnd.n3562 gnd.n1651 256.663
R4014 gnd.n3562 gnd.n1650 256.663
R4015 gnd.n3562 gnd.n1649 256.663
R4016 gnd.n3562 gnd.n1648 256.663
R4017 gnd.n3562 gnd.n1647 256.663
R4018 gnd.n3562 gnd.n1646 256.663
R4019 gnd.n3562 gnd.n1645 256.663
R4020 gnd.n3562 gnd.n1644 256.663
R4021 gnd.n3562 gnd.n1643 256.663
R4022 gnd.n3562 gnd.n1642 256.663
R4023 gnd.n3562 gnd.n1641 256.663
R4024 gnd.n3562 gnd.n1640 256.663
R4025 gnd.n3562 gnd.n1639 256.663
R4026 gnd.n3562 gnd.n1638 256.663
R4027 gnd.n3562 gnd.n1637 256.663
R4028 gnd.n4173 gnd.n1051 242.672
R4029 gnd.n4173 gnd.n1052 242.672
R4030 gnd.n4173 gnd.n1053 242.672
R4031 gnd.n4173 gnd.n1054 242.672
R4032 gnd.n4173 gnd.n1055 242.672
R4033 gnd.n4173 gnd.n1056 242.672
R4034 gnd.n4173 gnd.n1057 242.672
R4035 gnd.n4173 gnd.n1058 242.672
R4036 gnd.n4173 gnd.n1059 242.672
R4037 gnd.n3919 gnd.n1349 242.672
R4038 gnd.n3919 gnd.n1348 242.672
R4039 gnd.n3919 gnd.n1347 242.672
R4040 gnd.n3919 gnd.n1346 242.672
R4041 gnd.n3919 gnd.n1345 242.672
R4042 gnd.n3919 gnd.n1344 242.672
R4043 gnd.n3919 gnd.n1343 242.672
R4044 gnd.n3919 gnd.n1342 242.672
R4045 gnd.n3919 gnd.n1341 242.672
R4046 gnd.n4768 gnd.n4767 242.672
R4047 gnd.n4768 gnd.n4678 242.672
R4048 gnd.n4768 gnd.n4679 242.672
R4049 gnd.n4768 gnd.n4680 242.672
R4050 gnd.n4768 gnd.n4681 242.672
R4051 gnd.n4768 gnd.n4682 242.672
R4052 gnd.n4768 gnd.n4683 242.672
R4053 gnd.n4768 gnd.n4684 242.672
R4054 gnd.n4768 gnd.n4685 242.672
R4055 gnd.n4768 gnd.n4686 242.672
R4056 gnd.n4768 gnd.n4687 242.672
R4057 gnd.n4768 gnd.n4688 242.672
R4058 gnd.n4769 gnd.n4768 242.672
R4059 gnd.n5620 gnd.n1022 242.672
R4060 gnd.n5620 gnd.n1021 242.672
R4061 gnd.n5620 gnd.n1020 242.672
R4062 gnd.n5620 gnd.n1019 242.672
R4063 gnd.n5620 gnd.n1018 242.672
R4064 gnd.n5620 gnd.n1017 242.672
R4065 gnd.n5620 gnd.n1016 242.672
R4066 gnd.n5620 gnd.n1015 242.672
R4067 gnd.n5620 gnd.n1014 242.672
R4068 gnd.n5620 gnd.n1013 242.672
R4069 gnd.n5620 gnd.n1012 242.672
R4070 gnd.n5620 gnd.n1011 242.672
R4071 gnd.n5620 gnd.n1010 242.672
R4072 gnd.n6546 gnd.n313 242.672
R4073 gnd.n6546 gnd.n314 242.672
R4074 gnd.n6546 gnd.n315 242.672
R4075 gnd.n6546 gnd.n316 242.672
R4076 gnd.n6546 gnd.n317 242.672
R4077 gnd.n6546 gnd.n318 242.672
R4078 gnd.n6546 gnd.n319 242.672
R4079 gnd.n6546 gnd.n320 242.672
R4080 gnd.n6546 gnd.n321 242.672
R4081 gnd.n7058 gnd.n6852 242.672
R4082 gnd.n7058 gnd.n6748 242.672
R4083 gnd.n7058 gnd.n6747 242.672
R4084 gnd.n7058 gnd.n6746 242.672
R4085 gnd.n7058 gnd.n6745 242.672
R4086 gnd.n7058 gnd.n6744 242.672
R4087 gnd.n7058 gnd.n6743 242.672
R4088 gnd.n7058 gnd.n6742 242.672
R4089 gnd.n7058 gnd.n6741 242.672
R4090 gnd.n4852 gnd.n4851 242.672
R4091 gnd.n4851 gnd.n4590 242.672
R4092 gnd.n4851 gnd.n4591 242.672
R4093 gnd.n4851 gnd.n4592 242.672
R4094 gnd.n4851 gnd.n4593 242.672
R4095 gnd.n4851 gnd.n4594 242.672
R4096 gnd.n4851 gnd.n4595 242.672
R4097 gnd.n4851 gnd.n4596 242.672
R4098 gnd.n5620 gnd.n4174 242.672
R4099 gnd.n5620 gnd.n4175 242.672
R4100 gnd.n5620 gnd.n4176 242.672
R4101 gnd.n5620 gnd.n4177 242.672
R4102 gnd.n5620 gnd.n4178 242.672
R4103 gnd.n5620 gnd.n4179 242.672
R4104 gnd.n5620 gnd.n4180 242.672
R4105 gnd.n5620 gnd.n4181 242.672
R4106 gnd.n4173 gnd.n4172 242.672
R4107 gnd.n4173 gnd.n1023 242.672
R4108 gnd.n4173 gnd.n1024 242.672
R4109 gnd.n4173 gnd.n1025 242.672
R4110 gnd.n4173 gnd.n1026 242.672
R4111 gnd.n4173 gnd.n1027 242.672
R4112 gnd.n4173 gnd.n1028 242.672
R4113 gnd.n4173 gnd.n1029 242.672
R4114 gnd.n4173 gnd.n1030 242.672
R4115 gnd.n4173 gnd.n1031 242.672
R4116 gnd.n4173 gnd.n1032 242.672
R4117 gnd.n4173 gnd.n1033 242.672
R4118 gnd.n4173 gnd.n1034 242.672
R4119 gnd.n4173 gnd.n1035 242.672
R4120 gnd.n4173 gnd.n1036 242.672
R4121 gnd.n4173 gnd.n1037 242.672
R4122 gnd.n4173 gnd.n1038 242.672
R4123 gnd.n4173 gnd.n1039 242.672
R4124 gnd.n4173 gnd.n1040 242.672
R4125 gnd.n4173 gnd.n1041 242.672
R4126 gnd.n4173 gnd.n1042 242.672
R4127 gnd.n4173 gnd.n1043 242.672
R4128 gnd.n4173 gnd.n1044 242.672
R4129 gnd.n4173 gnd.n1045 242.672
R4130 gnd.n4173 gnd.n1046 242.672
R4131 gnd.n4173 gnd.n1047 242.672
R4132 gnd.n4173 gnd.n1048 242.672
R4133 gnd.n4173 gnd.n1049 242.672
R4134 gnd.n4173 gnd.n1050 242.672
R4135 gnd.n3919 gnd.n1351 242.672
R4136 gnd.n3919 gnd.n1352 242.672
R4137 gnd.n3919 gnd.n1353 242.672
R4138 gnd.n3919 gnd.n1354 242.672
R4139 gnd.n3919 gnd.n1355 242.672
R4140 gnd.n3919 gnd.n1356 242.672
R4141 gnd.n3919 gnd.n1357 242.672
R4142 gnd.n3919 gnd.n1358 242.672
R4143 gnd.n3919 gnd.n1359 242.672
R4144 gnd.n3919 gnd.n1360 242.672
R4145 gnd.n3919 gnd.n1361 242.672
R4146 gnd.n3919 gnd.n1362 242.672
R4147 gnd.n3919 gnd.n1363 242.672
R4148 gnd.n3919 gnd.n1364 242.672
R4149 gnd.n3919 gnd.n1365 242.672
R4150 gnd.n3919 gnd.n1366 242.672
R4151 gnd.n3869 gnd.n1407 242.672
R4152 gnd.n3919 gnd.n1367 242.672
R4153 gnd.n3919 gnd.n1368 242.672
R4154 gnd.n3919 gnd.n1369 242.672
R4155 gnd.n3919 gnd.n1370 242.672
R4156 gnd.n3919 gnd.n1371 242.672
R4157 gnd.n3919 gnd.n1372 242.672
R4158 gnd.n3919 gnd.n1373 242.672
R4159 gnd.n3919 gnd.n1374 242.672
R4160 gnd.n3919 gnd.n1375 242.672
R4161 gnd.n3919 gnd.n1376 242.672
R4162 gnd.n3919 gnd.n1377 242.672
R4163 gnd.n3919 gnd.n1378 242.672
R4164 gnd.n3919 gnd.n3918 242.672
R4165 gnd.n6547 gnd.n6546 242.672
R4166 gnd.n6546 gnd.n285 242.672
R4167 gnd.n6546 gnd.n286 242.672
R4168 gnd.n6546 gnd.n287 242.672
R4169 gnd.n6546 gnd.n288 242.672
R4170 gnd.n6546 gnd.n289 242.672
R4171 gnd.n6546 gnd.n290 242.672
R4172 gnd.n6546 gnd.n291 242.672
R4173 gnd.n6546 gnd.n292 242.672
R4174 gnd.n6546 gnd.n293 242.672
R4175 gnd.n6546 gnd.n294 242.672
R4176 gnd.n6546 gnd.n295 242.672
R4177 gnd.n6546 gnd.n296 242.672
R4178 gnd.n6497 gnd.n352 242.672
R4179 gnd.n6546 gnd.n297 242.672
R4180 gnd.n6546 gnd.n298 242.672
R4181 gnd.n6546 gnd.n299 242.672
R4182 gnd.n6546 gnd.n300 242.672
R4183 gnd.n6546 gnd.n301 242.672
R4184 gnd.n6546 gnd.n302 242.672
R4185 gnd.n6546 gnd.n303 242.672
R4186 gnd.n6546 gnd.n304 242.672
R4187 gnd.n6546 gnd.n305 242.672
R4188 gnd.n6546 gnd.n306 242.672
R4189 gnd.n6546 gnd.n307 242.672
R4190 gnd.n6546 gnd.n308 242.672
R4191 gnd.n6546 gnd.n309 242.672
R4192 gnd.n6546 gnd.n310 242.672
R4193 gnd.n6546 gnd.n311 242.672
R4194 gnd.n6546 gnd.n312 242.672
R4195 gnd.n7059 gnd.n7058 242.672
R4196 gnd.n7058 gnd.n6853 242.672
R4197 gnd.n7058 gnd.n6854 242.672
R4198 gnd.n7058 gnd.n6855 242.672
R4199 gnd.n7058 gnd.n6856 242.672
R4200 gnd.n7058 gnd.n6857 242.672
R4201 gnd.n7058 gnd.n6858 242.672
R4202 gnd.n7058 gnd.n6859 242.672
R4203 gnd.n7058 gnd.n6860 242.672
R4204 gnd.n7058 gnd.n6861 242.672
R4205 gnd.n7058 gnd.n6862 242.672
R4206 gnd.n7058 gnd.n6863 242.672
R4207 gnd.n7058 gnd.n6864 242.672
R4208 gnd.n7058 gnd.n6865 242.672
R4209 gnd.n7058 gnd.n6866 242.672
R4210 gnd.n7058 gnd.n6867 242.672
R4211 gnd.n7058 gnd.n6868 242.672
R4212 gnd.n7058 gnd.n6869 242.672
R4213 gnd.n7058 gnd.n6870 242.672
R4214 gnd.n7058 gnd.n6871 242.672
R4215 gnd.n7058 gnd.n6872 242.672
R4216 gnd.n7058 gnd.n6873 242.672
R4217 gnd.n7058 gnd.n6874 242.672
R4218 gnd.n7058 gnd.n6875 242.672
R4219 gnd.n7058 gnd.n6876 242.672
R4220 gnd.n7058 gnd.n6877 242.672
R4221 gnd.n7058 gnd.n6878 242.672
R4222 gnd.n7058 gnd.n6879 242.672
R4223 gnd.n7058 gnd.n6880 242.672
R4224 gnd.n2557 gnd.n2556 242.672
R4225 gnd.n2557 gnd.n2258 242.672
R4226 gnd.n2557 gnd.n2259 242.672
R4227 gnd.n2557 gnd.n2261 242.672
R4228 gnd.n2557 gnd.n2263 242.672
R4229 gnd.n2557 gnd.n2264 242.672
R4230 gnd.n2557 gnd.n2266 242.672
R4231 gnd.n2557 gnd.n2268 242.672
R4232 gnd.n2557 gnd.n2269 242.672
R4233 gnd.n2557 gnd.n2271 242.672
R4234 gnd.n2557 gnd.n2273 242.672
R4235 gnd.n2557 gnd.n2274 242.672
R4236 gnd.n2557 gnd.n2275 242.672
R4237 gnd.n2557 gnd.n2545 242.672
R4238 gnd.n6355 gnd.n486 242.672
R4239 gnd.n6355 gnd.n484 242.672
R4240 gnd.n6355 gnd.n483 242.672
R4241 gnd.n6355 gnd.n481 242.672
R4242 gnd.n6355 gnd.n479 242.672
R4243 gnd.n6355 gnd.n478 242.672
R4244 gnd.n6355 gnd.n476 242.672
R4245 gnd.n6355 gnd.n474 242.672
R4246 gnd.n6356 gnd.n6355 242.672
R4247 gnd.n6355 gnd.n469 242.672
R4248 gnd.n6355 gnd.n473 242.672
R4249 gnd.n6355 gnd.n471 242.672
R4250 gnd.n6355 gnd.n489 242.672
R4251 gnd.n6355 gnd.n488 242.672
R4252 gnd.n7057 gnd.n6881 240.244
R4253 gnd.n7050 gnd.n7049 240.244
R4254 gnd.n7047 gnd.n7046 240.244
R4255 gnd.n7043 gnd.n7042 240.244
R4256 gnd.n7039 gnd.n7038 240.244
R4257 gnd.n7035 gnd.n7034 240.244
R4258 gnd.n7031 gnd.n7030 240.244
R4259 gnd.n7027 gnd.n7026 240.244
R4260 gnd.n7023 gnd.n7022 240.244
R4261 gnd.n7016 gnd.n7015 240.244
R4262 gnd.n7012 gnd.n7011 240.244
R4263 gnd.n7008 gnd.n7007 240.244
R4264 gnd.n7004 gnd.n7003 240.244
R4265 gnd.n7000 gnd.n6999 240.244
R4266 gnd.n6996 gnd.n6995 240.244
R4267 gnd.n6992 gnd.n6991 240.244
R4268 gnd.n6988 gnd.n6987 240.244
R4269 gnd.n6984 gnd.n6983 240.244
R4270 gnd.n6980 gnd.n6979 240.244
R4271 gnd.n6973 gnd.n6972 240.244
R4272 gnd.n6970 gnd.n6969 240.244
R4273 gnd.n6966 gnd.n6965 240.244
R4274 gnd.n6962 gnd.n6961 240.244
R4275 gnd.n6958 gnd.n6957 240.244
R4276 gnd.n6954 gnd.n6953 240.244
R4277 gnd.n6950 gnd.n6949 240.244
R4278 gnd.n6946 gnd.n6945 240.244
R4279 gnd.n6942 gnd.n6941 240.244
R4280 gnd.n6938 gnd.n6739 240.244
R4281 gnd.n501 gnd.n275 240.244
R4282 gnd.n275 gnd.n266 240.244
R4283 gnd.n6566 gnd.n266 240.244
R4284 gnd.n6566 gnd.n256 240.244
R4285 gnd.n6570 gnd.n256 240.244
R4286 gnd.n6570 gnd.n247 240.244
R4287 gnd.n247 gnd.n238 240.244
R4288 gnd.n6611 gnd.n238 240.244
R4289 gnd.n6611 gnd.n230 240.244
R4290 gnd.n230 gnd.n220 240.244
R4291 gnd.n6630 gnd.n220 240.244
R4292 gnd.n6631 gnd.n6630 240.244
R4293 gnd.n6631 gnd.n210 240.244
R4294 gnd.n6634 gnd.n210 240.244
R4295 gnd.n6634 gnd.n201 240.244
R4296 gnd.n201 gnd.n193 240.244
R4297 gnd.n6669 gnd.n193 240.244
R4298 gnd.n6669 gnd.n186 240.244
R4299 gnd.n6671 gnd.n186 240.244
R4300 gnd.n6671 gnd.n177 240.244
R4301 gnd.n177 gnd.n172 240.244
R4302 gnd.n6695 gnd.n172 240.244
R4303 gnd.n6695 gnd.n73 240.244
R4304 gnd.n6702 gnd.n73 240.244
R4305 gnd.n6702 gnd.n84 240.244
R4306 gnd.n6705 gnd.n84 240.244
R4307 gnd.n6705 gnd.n95 240.244
R4308 gnd.n6709 gnd.n95 240.244
R4309 gnd.n6709 gnd.n105 240.244
R4310 gnd.n6712 gnd.n105 240.244
R4311 gnd.n6712 gnd.n114 240.244
R4312 gnd.n6716 gnd.n114 240.244
R4313 gnd.n6716 gnd.n124 240.244
R4314 gnd.n6719 gnd.n124 240.244
R4315 gnd.n6719 gnd.n133 240.244
R4316 gnd.n6723 gnd.n133 240.244
R4317 gnd.n6723 gnd.n143 240.244
R4318 gnd.n6726 gnd.n143 240.244
R4319 gnd.n6726 gnd.n152 240.244
R4320 gnd.n6730 gnd.n152 240.244
R4321 gnd.n6730 gnd.n162 240.244
R4322 gnd.n7060 gnd.n162 240.244
R4323 gnd.n6545 gnd.n283 240.244
R4324 gnd.n6545 gnd.n324 240.244
R4325 gnd.n6541 gnd.n6540 240.244
R4326 gnd.n6537 gnd.n6536 240.244
R4327 gnd.n6533 gnd.n6532 240.244
R4328 gnd.n6529 gnd.n6528 240.244
R4329 gnd.n6525 gnd.n6524 240.244
R4330 gnd.n6521 gnd.n6520 240.244
R4331 gnd.n6517 gnd.n6516 240.244
R4332 gnd.n6512 gnd.n6511 240.244
R4333 gnd.n6508 gnd.n6507 240.244
R4334 gnd.n6504 gnd.n6503 240.244
R4335 gnd.n6500 gnd.n6499 240.244
R4336 gnd.n6495 gnd.n6494 240.244
R4337 gnd.n6491 gnd.n6490 240.244
R4338 gnd.n6487 gnd.n6486 240.244
R4339 gnd.n6483 gnd.n6482 240.244
R4340 gnd.n6479 gnd.n6478 240.244
R4341 gnd.n6475 gnd.n6474 240.244
R4342 gnd.n6471 gnd.n6470 240.244
R4343 gnd.n6467 gnd.n6466 240.244
R4344 gnd.n6463 gnd.n6462 240.244
R4345 gnd.n6459 gnd.n6458 240.244
R4346 gnd.n6455 gnd.n6454 240.244
R4347 gnd.n6451 gnd.n6450 240.244
R4348 gnd.n6447 gnd.n6446 240.244
R4349 gnd.n6443 gnd.n6442 240.244
R4350 gnd.n6439 gnd.n6438 240.244
R4351 gnd.n6555 gnd.n277 240.244
R4352 gnd.n6555 gnd.n278 240.244
R4353 gnd.n278 gnd.n254 240.244
R4354 gnd.n6582 gnd.n254 240.244
R4355 gnd.n6582 gnd.n249 240.244
R4356 gnd.n6590 gnd.n249 240.244
R4357 gnd.n6590 gnd.n250 240.244
R4358 gnd.n250 gnd.n228 240.244
R4359 gnd.n6622 gnd.n228 240.244
R4360 gnd.n6622 gnd.n224 240.244
R4361 gnd.n6628 gnd.n224 240.244
R4362 gnd.n6628 gnd.n208 240.244
R4363 gnd.n6646 gnd.n208 240.244
R4364 gnd.n6646 gnd.n203 240.244
R4365 gnd.n6654 gnd.n203 240.244
R4366 gnd.n6654 gnd.n204 240.244
R4367 gnd.n204 gnd.n185 240.244
R4368 gnd.n6678 gnd.n185 240.244
R4369 gnd.n6678 gnd.n180 240.244
R4370 gnd.n6687 gnd.n180 240.244
R4371 gnd.n6687 gnd.n181 240.244
R4372 gnd.n181 gnd.n76 240.244
R4373 gnd.n7122 gnd.n76 240.244
R4374 gnd.n7122 gnd.n77 240.244
R4375 gnd.n7118 gnd.n77 240.244
R4376 gnd.n7118 gnd.n83 240.244
R4377 gnd.n7110 gnd.n83 240.244
R4378 gnd.n7110 gnd.n97 240.244
R4379 gnd.n7106 gnd.n97 240.244
R4380 gnd.n7106 gnd.n103 240.244
R4381 gnd.n7098 gnd.n103 240.244
R4382 gnd.n7098 gnd.n117 240.244
R4383 gnd.n7094 gnd.n117 240.244
R4384 gnd.n7094 gnd.n123 240.244
R4385 gnd.n7086 gnd.n123 240.244
R4386 gnd.n7086 gnd.n135 240.244
R4387 gnd.n7082 gnd.n135 240.244
R4388 gnd.n7082 gnd.n141 240.244
R4389 gnd.n7074 gnd.n141 240.244
R4390 gnd.n7074 gnd.n155 240.244
R4391 gnd.n7070 gnd.n155 240.244
R4392 gnd.n7070 gnd.n161 240.244
R4393 gnd.n3920 gnd.n1338 240.244
R4394 gnd.n3917 gnd.n1379 240.244
R4395 gnd.n3913 gnd.n3912 240.244
R4396 gnd.n3909 gnd.n3908 240.244
R4397 gnd.n3905 gnd.n3904 240.244
R4398 gnd.n3901 gnd.n3900 240.244
R4399 gnd.n3897 gnd.n3896 240.244
R4400 gnd.n3893 gnd.n3892 240.244
R4401 gnd.n3889 gnd.n3888 240.244
R4402 gnd.n3884 gnd.n3883 240.244
R4403 gnd.n3880 gnd.n3879 240.244
R4404 gnd.n3876 gnd.n3875 240.244
R4405 gnd.n3872 gnd.n3871 240.244
R4406 gnd.n2171 gnd.n2170 240.244
R4407 gnd.n2178 gnd.n2177 240.244
R4408 gnd.n2181 gnd.n2180 240.244
R4409 gnd.n2188 gnd.n2187 240.244
R4410 gnd.n2191 gnd.n2190 240.244
R4411 gnd.n2198 gnd.n2197 240.244
R4412 gnd.n2201 gnd.n2200 240.244
R4413 gnd.n2208 gnd.n2207 240.244
R4414 gnd.n2211 gnd.n2210 240.244
R4415 gnd.n2218 gnd.n2217 240.244
R4416 gnd.n2221 gnd.n2220 240.244
R4417 gnd.n2228 gnd.n2227 240.244
R4418 gnd.n2231 gnd.n2230 240.244
R4419 gnd.n2238 gnd.n2237 240.244
R4420 gnd.n2241 gnd.n2240 240.244
R4421 gnd.n1137 gnd.n1136 240.244
R4422 gnd.n2435 gnd.n1137 240.244
R4423 gnd.n2435 gnd.n1147 240.244
R4424 gnd.n2438 gnd.n1147 240.244
R4425 gnd.n2438 gnd.n1157 240.244
R4426 gnd.n2442 gnd.n1157 240.244
R4427 gnd.n2442 gnd.n1166 240.244
R4428 gnd.n2445 gnd.n1166 240.244
R4429 gnd.n2445 gnd.n1175 240.244
R4430 gnd.n2449 gnd.n1175 240.244
R4431 gnd.n2449 gnd.n1185 240.244
R4432 gnd.n2452 gnd.n1185 240.244
R4433 gnd.n2452 gnd.n1194 240.244
R4434 gnd.n2456 gnd.n1194 240.244
R4435 gnd.n2456 gnd.n1204 240.244
R4436 gnd.n2459 gnd.n1204 240.244
R4437 gnd.n2459 gnd.n1213 240.244
R4438 gnd.n2463 gnd.n1213 240.244
R4439 gnd.n2463 gnd.n1223 240.244
R4440 gnd.n2466 gnd.n1223 240.244
R4441 gnd.n2466 gnd.n1232 240.244
R4442 gnd.n2470 gnd.n1232 240.244
R4443 gnd.n2470 gnd.n1242 240.244
R4444 gnd.n2473 gnd.n1242 240.244
R4445 gnd.n2473 gnd.n1251 240.244
R4446 gnd.n2477 gnd.n1251 240.244
R4447 gnd.n2477 gnd.n1261 240.244
R4448 gnd.n2480 gnd.n1261 240.244
R4449 gnd.n2480 gnd.n1270 240.244
R4450 gnd.n2484 gnd.n1270 240.244
R4451 gnd.n2484 gnd.n1280 240.244
R4452 gnd.n2487 gnd.n1280 240.244
R4453 gnd.n2487 gnd.n1289 240.244
R4454 gnd.n2491 gnd.n1289 240.244
R4455 gnd.n2491 gnd.n1300 240.244
R4456 gnd.n2495 gnd.n1300 240.244
R4457 gnd.n2495 gnd.n1310 240.244
R4458 gnd.n2506 gnd.n1310 240.244
R4459 gnd.n2506 gnd.n1321 240.244
R4460 gnd.n2513 gnd.n1321 240.244
R4461 gnd.n2513 gnd.n1330 240.244
R4462 gnd.n2248 gnd.n1330 240.244
R4463 gnd.n1063 gnd.n1062 240.244
R4464 gnd.n4166 gnd.n1062 240.244
R4465 gnd.n4164 gnd.n4163 240.244
R4466 gnd.n4160 gnd.n4159 240.244
R4467 gnd.n4156 gnd.n4155 240.244
R4468 gnd.n4152 gnd.n4151 240.244
R4469 gnd.n4148 gnd.n4147 240.244
R4470 gnd.n4144 gnd.n4143 240.244
R4471 gnd.n4140 gnd.n4139 240.244
R4472 gnd.n4135 gnd.n4134 240.244
R4473 gnd.n4131 gnd.n4130 240.244
R4474 gnd.n4127 gnd.n4126 240.244
R4475 gnd.n4123 gnd.n4122 240.244
R4476 gnd.n4119 gnd.n4118 240.244
R4477 gnd.n4115 gnd.n4114 240.244
R4478 gnd.n4111 gnd.n4110 240.244
R4479 gnd.n4107 gnd.n4106 240.244
R4480 gnd.n4103 gnd.n4102 240.244
R4481 gnd.n4099 gnd.n4098 240.244
R4482 gnd.n4095 gnd.n4094 240.244
R4483 gnd.n4091 gnd.n4090 240.244
R4484 gnd.n4087 gnd.n4086 240.244
R4485 gnd.n4083 gnd.n4082 240.244
R4486 gnd.n4079 gnd.n4078 240.244
R4487 gnd.n4075 gnd.n4074 240.244
R4488 gnd.n4071 gnd.n4070 240.244
R4489 gnd.n4067 gnd.n4066 240.244
R4490 gnd.n4063 gnd.n4062 240.244
R4491 gnd.n4059 gnd.n4058 240.244
R4492 gnd.n4048 gnd.n1064 240.244
R4493 gnd.n4048 gnd.n1139 240.244
R4494 gnd.n4042 gnd.n1139 240.244
R4495 gnd.n4042 gnd.n1145 240.244
R4496 gnd.n4034 gnd.n1145 240.244
R4497 gnd.n4034 gnd.n1160 240.244
R4498 gnd.n4030 gnd.n1160 240.244
R4499 gnd.n4030 gnd.n1165 240.244
R4500 gnd.n4022 gnd.n1165 240.244
R4501 gnd.n4022 gnd.n1177 240.244
R4502 gnd.n4018 gnd.n1177 240.244
R4503 gnd.n4018 gnd.n1183 240.244
R4504 gnd.n4010 gnd.n1183 240.244
R4505 gnd.n4010 gnd.n1197 240.244
R4506 gnd.n4006 gnd.n1197 240.244
R4507 gnd.n4006 gnd.n1203 240.244
R4508 gnd.n3998 gnd.n1203 240.244
R4509 gnd.n3998 gnd.n1215 240.244
R4510 gnd.n3994 gnd.n1215 240.244
R4511 gnd.n3994 gnd.n1221 240.244
R4512 gnd.n3986 gnd.n1221 240.244
R4513 gnd.n3986 gnd.n1235 240.244
R4514 gnd.n3982 gnd.n1235 240.244
R4515 gnd.n3982 gnd.n1241 240.244
R4516 gnd.n3974 gnd.n1241 240.244
R4517 gnd.n3974 gnd.n1254 240.244
R4518 gnd.n3970 gnd.n1254 240.244
R4519 gnd.n3970 gnd.n1260 240.244
R4520 gnd.n3962 gnd.n1260 240.244
R4521 gnd.n3962 gnd.n1273 240.244
R4522 gnd.n3958 gnd.n1273 240.244
R4523 gnd.n3958 gnd.n1279 240.244
R4524 gnd.n3950 gnd.n1279 240.244
R4525 gnd.n3950 gnd.n1292 240.244
R4526 gnd.n3946 gnd.n1292 240.244
R4527 gnd.n3946 gnd.n1298 240.244
R4528 gnd.n3938 gnd.n1298 240.244
R4529 gnd.n3938 gnd.n1313 240.244
R4530 gnd.n3934 gnd.n1313 240.244
R4531 gnd.n3934 gnd.n1319 240.244
R4532 gnd.n3926 gnd.n1319 240.244
R4533 gnd.n3926 gnd.n1333 240.244
R4534 gnd.n5619 gnd.n4183 240.244
R4535 gnd.n5612 gnd.n5611 240.244
R4536 gnd.n5609 gnd.n5608 240.244
R4537 gnd.n5605 gnd.n5604 240.244
R4538 gnd.n5601 gnd.n5600 240.244
R4539 gnd.n5597 gnd.n5596 240.244
R4540 gnd.n5593 gnd.n5592 240.244
R4541 gnd.n5589 gnd.n5588 240.244
R4542 gnd.n4863 gnd.n4575 240.244
R4543 gnd.n4873 gnd.n4575 240.244
R4544 gnd.n4873 gnd.n4566 240.244
R4545 gnd.n4566 gnd.n4555 240.244
R4546 gnd.n4894 gnd.n4555 240.244
R4547 gnd.n4894 gnd.n4549 240.244
R4548 gnd.n4904 gnd.n4549 240.244
R4549 gnd.n4904 gnd.n4538 240.244
R4550 gnd.n4538 gnd.n4530 240.244
R4551 gnd.n4922 gnd.n4530 240.244
R4552 gnd.n4923 gnd.n4922 240.244
R4553 gnd.n4923 gnd.n4515 240.244
R4554 gnd.n4925 gnd.n4515 240.244
R4555 gnd.n4925 gnd.n4501 240.244
R4556 gnd.n4967 gnd.n4501 240.244
R4557 gnd.n4968 gnd.n4967 240.244
R4558 gnd.n4971 gnd.n4968 240.244
R4559 gnd.n4971 gnd.n4456 240.244
R4560 gnd.n4496 gnd.n4456 240.244
R4561 gnd.n4496 gnd.n4466 240.244
R4562 gnd.n4981 gnd.n4466 240.244
R4563 gnd.n4981 gnd.n4487 240.244
R4564 gnd.n4991 gnd.n4487 240.244
R4565 gnd.n4991 gnd.n4385 240.244
R4566 gnd.n5036 gnd.n4385 240.244
R4567 gnd.n5036 gnd.n4371 240.244
R4568 gnd.n5058 gnd.n4371 240.244
R4569 gnd.n5059 gnd.n5058 240.244
R4570 gnd.n5059 gnd.n4358 240.244
R4571 gnd.n4358 gnd.n4347 240.244
R4572 gnd.n5090 gnd.n4347 240.244
R4573 gnd.n5091 gnd.n5090 240.244
R4574 gnd.n5092 gnd.n5091 240.244
R4575 gnd.n5092 gnd.n4332 240.244
R4576 gnd.n4332 gnd.n4331 240.244
R4577 gnd.n4331 gnd.n4316 240.244
R4578 gnd.n5143 gnd.n4316 240.244
R4579 gnd.n5144 gnd.n5143 240.244
R4580 gnd.n5144 gnd.n4303 240.244
R4581 gnd.n4303 gnd.n4292 240.244
R4582 gnd.n5175 gnd.n4292 240.244
R4583 gnd.n5176 gnd.n5175 240.244
R4584 gnd.n5177 gnd.n5176 240.244
R4585 gnd.n5177 gnd.n4276 240.244
R4586 gnd.n4276 gnd.n4275 240.244
R4587 gnd.n4275 gnd.n4262 240.244
R4588 gnd.n5232 gnd.n4262 240.244
R4589 gnd.n5233 gnd.n5232 240.244
R4590 gnd.n5233 gnd.n4249 240.244
R4591 gnd.n4249 gnd.n4239 240.244
R4592 gnd.n5520 gnd.n4239 240.244
R4593 gnd.n5523 gnd.n5520 240.244
R4594 gnd.n5523 gnd.n5522 240.244
R4595 gnd.n4853 gnd.n4588 240.244
R4596 gnd.n4609 gnd.n4588 240.244
R4597 gnd.n4612 gnd.n4611 240.244
R4598 gnd.n4619 gnd.n4618 240.244
R4599 gnd.n4622 gnd.n4621 240.244
R4600 gnd.n4629 gnd.n4628 240.244
R4601 gnd.n4632 gnd.n4631 240.244
R4602 gnd.n4639 gnd.n4638 240.244
R4603 gnd.n4861 gnd.n4585 240.244
R4604 gnd.n4585 gnd.n4564 240.244
R4605 gnd.n4884 gnd.n4564 240.244
R4606 gnd.n4884 gnd.n4558 240.244
R4607 gnd.n4892 gnd.n4558 240.244
R4608 gnd.n4892 gnd.n4560 240.244
R4609 gnd.n4560 gnd.n4536 240.244
R4610 gnd.n4914 gnd.n4536 240.244
R4611 gnd.n4914 gnd.n4532 240.244
R4612 gnd.n4920 gnd.n4532 240.244
R4613 gnd.n4920 gnd.n4514 240.244
R4614 gnd.n4945 gnd.n4514 240.244
R4615 gnd.n4945 gnd.n4509 240.244
R4616 gnd.n4957 gnd.n4509 240.244
R4617 gnd.n4957 gnd.n4510 240.244
R4618 gnd.n4953 gnd.n4510 240.244
R4619 gnd.n4953 gnd.n4458 240.244
R4620 gnd.n5005 gnd.n4458 240.244
R4621 gnd.n5005 gnd.n4459 240.244
R4622 gnd.n5001 gnd.n4459 240.244
R4623 gnd.n5001 gnd.n4465 240.244
R4624 gnd.n4485 gnd.n4465 240.244
R4625 gnd.n4485 gnd.n4383 240.244
R4626 gnd.n5040 gnd.n4383 240.244
R4627 gnd.n5040 gnd.n4378 240.244
R4628 gnd.n5048 gnd.n4378 240.244
R4629 gnd.n5048 gnd.n4379 240.244
R4630 gnd.n4379 gnd.n4356 240.244
R4631 gnd.n5080 gnd.n4356 240.244
R4632 gnd.n5080 gnd.n4351 240.244
R4633 gnd.n5088 gnd.n4351 240.244
R4634 gnd.n5088 gnd.n4352 240.244
R4635 gnd.n4352 gnd.n4329 240.244
R4636 gnd.n5125 gnd.n4329 240.244
R4637 gnd.n5125 gnd.n4324 240.244
R4638 gnd.n5133 gnd.n4324 240.244
R4639 gnd.n5133 gnd.n4325 240.244
R4640 gnd.n4325 gnd.n4301 240.244
R4641 gnd.n5165 gnd.n4301 240.244
R4642 gnd.n5165 gnd.n4296 240.244
R4643 gnd.n5173 gnd.n4296 240.244
R4644 gnd.n5173 gnd.n4297 240.244
R4645 gnd.n4297 gnd.n4274 240.244
R4646 gnd.n5214 gnd.n4274 240.244
R4647 gnd.n5214 gnd.n4269 240.244
R4648 gnd.n5222 gnd.n4269 240.244
R4649 gnd.n5222 gnd.n4270 240.244
R4650 gnd.n4270 gnd.n4247 240.244
R4651 gnd.n5508 gnd.n4247 240.244
R4652 gnd.n5508 gnd.n4242 240.244
R4653 gnd.n5518 gnd.n4242 240.244
R4654 gnd.n5518 gnd.n4243 240.244
R4655 gnd.n4243 gnd.n4182 240.244
R4656 gnd.n6762 gnd.n6740 240.244
R4657 gnd.n6768 gnd.n6767 240.244
R4658 gnd.n6771 gnd.n6770 240.244
R4659 gnd.n6778 gnd.n6777 240.244
R4660 gnd.n6781 gnd.n6780 240.244
R4661 gnd.n6788 gnd.n6787 240.244
R4662 gnd.n6791 gnd.n6790 240.244
R4663 gnd.n6798 gnd.n6797 240.244
R4664 gnd.n6800 gnd.n6749 240.244
R4665 gnd.n6557 gnd.n273 240.244
R4666 gnd.n6557 gnd.n268 240.244
R4667 gnd.n6564 gnd.n268 240.244
R4668 gnd.n6564 gnd.n257 240.244
R4669 gnd.n257 gnd.n245 240.244
R4670 gnd.n6592 gnd.n245 240.244
R4671 gnd.n6592 gnd.n240 240.244
R4672 gnd.n6609 gnd.n240 240.244
R4673 gnd.n6609 gnd.n231 240.244
R4674 gnd.n6597 gnd.n231 240.244
R4675 gnd.n6597 gnd.n222 240.244
R4676 gnd.n6598 gnd.n222 240.244
R4677 gnd.n6598 gnd.n211 240.244
R4678 gnd.n211 gnd.n200 240.244
R4679 gnd.n6656 gnd.n200 240.244
R4680 gnd.n6656 gnd.n195 240.244
R4681 gnd.n6667 gnd.n195 240.244
R4682 gnd.n6667 gnd.n187 240.244
R4683 gnd.n6660 gnd.n187 240.244
R4684 gnd.n6660 gnd.n179 240.244
R4685 gnd.n179 gnd.n178 240.244
R4686 gnd.n178 gnd.n70 240.244
R4687 gnd.n7124 gnd.n70 240.244
R4688 gnd.n7124 gnd.n72 240.244
R4689 gnd.n85 gnd.n72 240.244
R4690 gnd.n6815 gnd.n85 240.244
R4691 gnd.n6815 gnd.n96 240.244
R4692 gnd.n6820 gnd.n96 240.244
R4693 gnd.n6820 gnd.n106 240.244
R4694 gnd.n6823 gnd.n106 240.244
R4695 gnd.n6823 gnd.n115 240.244
R4696 gnd.n6828 gnd.n115 240.244
R4697 gnd.n6828 gnd.n125 240.244
R4698 gnd.n6831 gnd.n125 240.244
R4699 gnd.n6831 gnd.n134 240.244
R4700 gnd.n6836 gnd.n134 240.244
R4701 gnd.n6836 gnd.n144 240.244
R4702 gnd.n6839 gnd.n144 240.244
R4703 gnd.n6839 gnd.n153 240.244
R4704 gnd.n6844 gnd.n153 240.244
R4705 gnd.n6844 gnd.n163 240.244
R4706 gnd.n6750 gnd.n163 240.244
R4707 gnd.n400 gnd.n399 240.244
R4708 gnd.n408 gnd.n407 240.244
R4709 gnd.n410 gnd.n409 240.244
R4710 gnd.n418 gnd.n417 240.244
R4711 gnd.n426 gnd.n425 240.244
R4712 gnd.n428 gnd.n427 240.244
R4713 gnd.n436 gnd.n435 240.244
R4714 gnd.n446 gnd.n445 240.244
R4715 gnd.n6382 gnd.n322 240.244
R4716 gnd.n6344 gnd.n276 240.244
R4717 gnd.n6340 gnd.n276 240.244
R4718 gnd.n6340 gnd.n259 240.244
R4719 gnd.n6580 gnd.n259 240.244
R4720 gnd.n6580 gnd.n260 240.244
R4721 gnd.n260 gnd.n248 240.244
R4722 gnd.n6575 gnd.n248 240.244
R4723 gnd.n6575 gnd.n232 240.244
R4724 gnd.n6620 gnd.n232 240.244
R4725 gnd.n6620 gnd.n233 240.244
R4726 gnd.n233 gnd.n223 240.244
R4727 gnd.n223 gnd.n213 240.244
R4728 gnd.n6644 gnd.n213 240.244
R4729 gnd.n6644 gnd.n214 240.244
R4730 gnd.n214 gnd.n202 240.244
R4731 gnd.n6639 gnd.n202 240.244
R4732 gnd.n6639 gnd.n189 240.244
R4733 gnd.n6676 gnd.n189 240.244
R4734 gnd.n6676 gnd.n176 240.244
R4735 gnd.n6689 gnd.n176 240.244
R4736 gnd.n6689 gnd.n170 240.244
R4737 gnd.n6697 gnd.n170 240.244
R4738 gnd.n6697 gnd.n75 240.244
R4739 gnd.n87 gnd.n75 240.244
R4740 gnd.n7116 gnd.n87 240.244
R4741 gnd.n7116 gnd.n88 240.244
R4742 gnd.n7112 gnd.n88 240.244
R4743 gnd.n7112 gnd.n94 240.244
R4744 gnd.n7104 gnd.n94 240.244
R4745 gnd.n7104 gnd.n108 240.244
R4746 gnd.n7100 gnd.n108 240.244
R4747 gnd.n7100 gnd.n113 240.244
R4748 gnd.n7092 gnd.n113 240.244
R4749 gnd.n7092 gnd.n127 240.244
R4750 gnd.n7088 gnd.n127 240.244
R4751 gnd.n7088 gnd.n132 240.244
R4752 gnd.n7080 gnd.n132 240.244
R4753 gnd.n7080 gnd.n146 240.244
R4754 gnd.n7076 gnd.n146 240.244
R4755 gnd.n7076 gnd.n151 240.244
R4756 gnd.n7068 gnd.n151 240.244
R4757 gnd.n7068 gnd.n165 240.244
R4758 gnd.n4202 gnd.n1009 240.244
R4759 gnd.n5579 gnd.n5578 240.244
R4760 gnd.n5575 gnd.n5574 240.244
R4761 gnd.n5571 gnd.n5570 240.244
R4762 gnd.n5567 gnd.n5566 240.244
R4763 gnd.n5563 gnd.n5562 240.244
R4764 gnd.n5559 gnd.n5558 240.244
R4765 gnd.n5555 gnd.n5554 240.244
R4766 gnd.n5551 gnd.n5550 240.244
R4767 gnd.n5547 gnd.n5546 240.244
R4768 gnd.n5543 gnd.n5542 240.244
R4769 gnd.n5539 gnd.n5538 240.244
R4770 gnd.n5535 gnd.n5534 240.244
R4771 gnd.n4776 gnd.n4673 240.244
R4772 gnd.n4776 gnd.n4666 240.244
R4773 gnd.n4787 gnd.n4666 240.244
R4774 gnd.n4787 gnd.n4662 240.244
R4775 gnd.n4793 gnd.n4662 240.244
R4776 gnd.n4793 gnd.n4654 240.244
R4777 gnd.n4803 gnd.n4654 240.244
R4778 gnd.n4803 gnd.n4649 240.244
R4779 gnd.n4839 gnd.n4649 240.244
R4780 gnd.n4839 gnd.n4650 240.244
R4781 gnd.n4650 gnd.n4597 240.244
R4782 gnd.n4834 gnd.n4597 240.244
R4783 gnd.n4834 gnd.n4833 240.244
R4784 gnd.n4833 gnd.n4576 240.244
R4785 gnd.n4829 gnd.n4576 240.244
R4786 gnd.n4829 gnd.n4567 240.244
R4787 gnd.n4826 gnd.n4567 240.244
R4788 gnd.n4826 gnd.n4825 240.244
R4789 gnd.n4825 gnd.n4550 240.244
R4790 gnd.n4821 gnd.n4550 240.244
R4791 gnd.n4821 gnd.n4539 240.244
R4792 gnd.n4539 gnd.n4520 240.244
R4793 gnd.n4934 gnd.n4520 240.244
R4794 gnd.n4934 gnd.n4516 240.244
R4795 gnd.n4942 gnd.n4516 240.244
R4796 gnd.n4942 gnd.n4507 240.244
R4797 gnd.n4507 gnd.n4443 240.244
R4798 gnd.n5014 gnd.n4443 240.244
R4799 gnd.n5014 gnd.n4444 240.244
R4800 gnd.n4455 gnd.n4444 240.244
R4801 gnd.n4490 gnd.n4455 240.244
R4802 gnd.n4493 gnd.n4490 240.244
R4803 gnd.n4493 gnd.n4467 240.244
R4804 gnd.n4480 gnd.n4467 240.244
R4805 gnd.n4480 gnd.n4477 240.244
R4806 gnd.n4477 gnd.n4386 240.244
R4807 gnd.n5035 gnd.n4386 240.244
R4808 gnd.n5035 gnd.n4376 240.244
R4809 gnd.n5031 gnd.n4376 240.244
R4810 gnd.n5031 gnd.n4370 240.244
R4811 gnd.n5028 gnd.n4370 240.244
R4812 gnd.n5028 gnd.n4359 240.244
R4813 gnd.n5025 gnd.n4359 240.244
R4814 gnd.n5025 gnd.n4337 240.244
R4815 gnd.n5101 gnd.n4337 240.244
R4816 gnd.n5101 gnd.n4333 240.244
R4817 gnd.n5122 gnd.n4333 240.244
R4818 gnd.n5122 gnd.n4322 240.244
R4819 gnd.n5118 gnd.n4322 240.244
R4820 gnd.n5118 gnd.n4315 240.244
R4821 gnd.n5115 gnd.n4315 240.244
R4822 gnd.n5115 gnd.n4304 240.244
R4823 gnd.n5112 gnd.n4304 240.244
R4824 gnd.n5112 gnd.n4281 240.244
R4825 gnd.n5186 gnd.n4281 240.244
R4826 gnd.n5186 gnd.n4277 240.244
R4827 gnd.n5211 gnd.n4277 240.244
R4828 gnd.n5211 gnd.n4268 240.244
R4829 gnd.n5207 gnd.n4268 240.244
R4830 gnd.n5207 gnd.n4261 240.244
R4831 gnd.n5203 gnd.n4261 240.244
R4832 gnd.n5203 gnd.n4250 240.244
R4833 gnd.n5200 gnd.n4250 240.244
R4834 gnd.n5200 gnd.n4231 240.244
R4835 gnd.n5530 gnd.n4231 240.244
R4836 gnd.n4690 gnd.n4689 240.244
R4837 gnd.n4761 gnd.n4689 240.244
R4838 gnd.n4759 gnd.n4758 240.244
R4839 gnd.n4755 gnd.n4754 240.244
R4840 gnd.n4751 gnd.n4750 240.244
R4841 gnd.n4747 gnd.n4746 240.244
R4842 gnd.n4743 gnd.n4742 240.244
R4843 gnd.n4739 gnd.n4738 240.244
R4844 gnd.n4735 gnd.n4734 240.244
R4845 gnd.n4731 gnd.n4730 240.244
R4846 gnd.n4727 gnd.n4726 240.244
R4847 gnd.n4723 gnd.n4722 240.244
R4848 gnd.n4719 gnd.n4677 240.244
R4849 gnd.n4779 gnd.n4671 240.244
R4850 gnd.n4779 gnd.n4667 240.244
R4851 gnd.n4785 gnd.n4667 240.244
R4852 gnd.n4785 gnd.n4660 240.244
R4853 gnd.n4795 gnd.n4660 240.244
R4854 gnd.n4795 gnd.n4656 240.244
R4855 gnd.n4801 gnd.n4656 240.244
R4856 gnd.n4801 gnd.n4647 240.244
R4857 gnd.n4841 gnd.n4647 240.244
R4858 gnd.n4841 gnd.n4598 240.244
R4859 gnd.n4849 gnd.n4598 240.244
R4860 gnd.n4849 gnd.n4599 240.244
R4861 gnd.n4599 gnd.n4577 240.244
R4862 gnd.n4870 gnd.n4577 240.244
R4863 gnd.n4870 gnd.n4569 240.244
R4864 gnd.n4881 gnd.n4569 240.244
R4865 gnd.n4881 gnd.n4570 240.244
R4866 gnd.n4570 gnd.n4551 240.244
R4867 gnd.n4901 gnd.n4551 240.244
R4868 gnd.n4901 gnd.n4541 240.244
R4869 gnd.n4911 gnd.n4541 240.244
R4870 gnd.n4911 gnd.n4522 240.244
R4871 gnd.n4932 gnd.n4522 240.244
R4872 gnd.n4932 gnd.n4524 240.244
R4873 gnd.n4524 gnd.n4505 240.244
R4874 gnd.n4960 gnd.n4505 240.244
R4875 gnd.n4960 gnd.n4447 240.244
R4876 gnd.n5012 gnd.n4447 240.244
R4877 gnd.n5012 gnd.n4448 240.244
R4878 gnd.n5008 gnd.n4448 240.244
R4879 gnd.n5008 gnd.n4454 240.244
R4880 gnd.n4469 gnd.n4454 240.244
R4881 gnd.n4998 gnd.n4469 240.244
R4882 gnd.n4998 gnd.n4470 240.244
R4883 gnd.n4994 gnd.n4470 240.244
R4884 gnd.n4994 gnd.n4476 240.244
R4885 gnd.n4476 gnd.n4375 240.244
R4886 gnd.n5051 gnd.n4375 240.244
R4887 gnd.n5051 gnd.n4368 240.244
R4888 gnd.n5062 gnd.n4368 240.244
R4889 gnd.n5062 gnd.n4361 240.244
R4890 gnd.n5077 gnd.n4361 240.244
R4891 gnd.n5077 gnd.n4362 240.244
R4892 gnd.n4362 gnd.n4340 240.244
R4893 gnd.n5099 gnd.n4340 240.244
R4894 gnd.n5099 gnd.n4341 240.244
R4895 gnd.n4341 gnd.n4320 240.244
R4896 gnd.n5136 gnd.n4320 240.244
R4897 gnd.n5136 gnd.n4313 240.244
R4898 gnd.n5147 gnd.n4313 240.244
R4899 gnd.n5147 gnd.n4306 240.244
R4900 gnd.n5162 gnd.n4306 240.244
R4901 gnd.n5162 gnd.n4307 240.244
R4902 gnd.n4307 gnd.n4284 240.244
R4903 gnd.n5184 gnd.n4284 240.244
R4904 gnd.n5184 gnd.n4286 240.244
R4905 gnd.n4286 gnd.n4266 240.244
R4906 gnd.n5225 gnd.n4266 240.244
R4907 gnd.n5225 gnd.n4259 240.244
R4908 gnd.n5236 gnd.n4259 240.244
R4909 gnd.n5236 gnd.n4252 240.244
R4910 gnd.n5505 gnd.n4252 240.244
R4911 gnd.n5505 gnd.n4253 240.244
R4912 gnd.n4253 gnd.n4234 240.244
R4913 gnd.n5528 gnd.n4234 240.244
R4914 gnd.n2098 gnd.n1340 240.244
R4915 gnd.n2100 gnd.n2099 240.244
R4916 gnd.n2108 gnd.n2107 240.244
R4917 gnd.n2116 gnd.n2115 240.244
R4918 gnd.n2118 gnd.n2117 240.244
R4919 gnd.n2126 gnd.n2125 240.244
R4920 gnd.n2134 gnd.n2133 240.244
R4921 gnd.n2136 gnd.n2135 240.244
R4922 gnd.n2149 gnd.n2145 240.244
R4923 gnd.n2365 gnd.n1138 240.244
R4924 gnd.n2370 gnd.n1138 240.244
R4925 gnd.n2370 gnd.n1148 240.244
R4926 gnd.n2373 gnd.n1148 240.244
R4927 gnd.n2373 gnd.n1158 240.244
R4928 gnd.n2378 gnd.n1158 240.244
R4929 gnd.n2378 gnd.n1167 240.244
R4930 gnd.n2381 gnd.n1167 240.244
R4931 gnd.n2381 gnd.n1176 240.244
R4932 gnd.n2386 gnd.n1176 240.244
R4933 gnd.n2386 gnd.n1186 240.244
R4934 gnd.n2389 gnd.n1186 240.244
R4935 gnd.n2389 gnd.n1195 240.244
R4936 gnd.n2394 gnd.n1195 240.244
R4937 gnd.n2394 gnd.n1205 240.244
R4938 gnd.n2397 gnd.n1205 240.244
R4939 gnd.n2397 gnd.n1214 240.244
R4940 gnd.n2402 gnd.n1214 240.244
R4941 gnd.n2402 gnd.n1224 240.244
R4942 gnd.n2405 gnd.n1224 240.244
R4943 gnd.n2405 gnd.n1233 240.244
R4944 gnd.n2298 gnd.n1233 240.244
R4945 gnd.n2298 gnd.n1243 240.244
R4946 gnd.n2412 gnd.n1243 240.244
R4947 gnd.n2412 gnd.n1252 240.244
R4948 gnd.n2295 gnd.n1252 240.244
R4949 gnd.n2295 gnd.n1262 240.244
R4950 gnd.n2419 gnd.n1262 240.244
R4951 gnd.n2419 gnd.n1271 240.244
R4952 gnd.n2292 gnd.n1271 240.244
R4953 gnd.n2292 gnd.n1281 240.244
R4954 gnd.n2426 gnd.n1281 240.244
R4955 gnd.n2426 gnd.n1290 240.244
R4956 gnd.n2289 gnd.n1290 240.244
R4957 gnd.n2289 gnd.n1301 240.244
R4958 gnd.n2497 gnd.n1301 240.244
R4959 gnd.n2497 gnd.n1311 240.244
R4960 gnd.n2504 gnd.n1311 240.244
R4961 gnd.n2504 gnd.n1322 240.244
R4962 gnd.n2536 gnd.n1322 240.244
R4963 gnd.n2536 gnd.n1331 240.244
R4964 gnd.n2568 gnd.n1331 240.244
R4965 gnd.n2326 gnd.n2325 240.244
R4966 gnd.n2332 gnd.n2331 240.244
R4967 gnd.n2336 gnd.n2335 240.244
R4968 gnd.n2342 gnd.n2341 240.244
R4969 gnd.n2346 gnd.n2345 240.244
R4970 gnd.n2352 gnd.n2351 240.244
R4971 gnd.n2356 gnd.n2355 240.244
R4972 gnd.n2315 gnd.n2314 240.244
R4973 gnd.n2310 gnd.n1060 240.244
R4974 gnd.n4051 gnd.n4050 240.244
R4975 gnd.n4050 gnd.n1134 240.244
R4976 gnd.n4040 gnd.n1134 240.244
R4977 gnd.n4040 gnd.n1150 240.244
R4978 gnd.n4036 gnd.n1150 240.244
R4979 gnd.n4036 gnd.n1156 240.244
R4980 gnd.n4028 gnd.n1156 240.244
R4981 gnd.n4028 gnd.n1169 240.244
R4982 gnd.n4024 gnd.n1169 240.244
R4983 gnd.n4024 gnd.n1174 240.244
R4984 gnd.n4016 gnd.n1174 240.244
R4985 gnd.n4016 gnd.n1187 240.244
R4986 gnd.n4012 gnd.n1187 240.244
R4987 gnd.n4012 gnd.n1192 240.244
R4988 gnd.n4004 gnd.n1192 240.244
R4989 gnd.n4004 gnd.n1207 240.244
R4990 gnd.n4000 gnd.n1207 240.244
R4991 gnd.n4000 gnd.n1212 240.244
R4992 gnd.n3992 gnd.n1212 240.244
R4993 gnd.n3992 gnd.n1225 240.244
R4994 gnd.n3988 gnd.n1225 240.244
R4995 gnd.n3988 gnd.n1230 240.244
R4996 gnd.n3980 gnd.n1230 240.244
R4997 gnd.n3980 gnd.n1245 240.244
R4998 gnd.n3976 gnd.n1245 240.244
R4999 gnd.n3976 gnd.n1250 240.244
R5000 gnd.n3968 gnd.n1250 240.244
R5001 gnd.n3968 gnd.n1263 240.244
R5002 gnd.n3964 gnd.n1263 240.244
R5003 gnd.n3964 gnd.n1268 240.244
R5004 gnd.n3956 gnd.n1268 240.244
R5005 gnd.n3956 gnd.n1283 240.244
R5006 gnd.n3952 gnd.n1283 240.244
R5007 gnd.n3952 gnd.n1288 240.244
R5008 gnd.n3944 gnd.n1288 240.244
R5009 gnd.n3944 gnd.n1303 240.244
R5010 gnd.n3940 gnd.n1303 240.244
R5011 gnd.n3940 gnd.n1308 240.244
R5012 gnd.n3932 gnd.n1308 240.244
R5013 gnd.n3932 gnd.n1324 240.244
R5014 gnd.n3928 gnd.n1324 240.244
R5015 gnd.n3928 gnd.n1329 240.244
R5016 gnd.n5791 gnd.n836 240.244
R5017 gnd.n5797 gnd.n836 240.244
R5018 gnd.n5797 gnd.n834 240.244
R5019 gnd.n5801 gnd.n834 240.244
R5020 gnd.n5801 gnd.n830 240.244
R5021 gnd.n5807 gnd.n830 240.244
R5022 gnd.n5807 gnd.n828 240.244
R5023 gnd.n5811 gnd.n828 240.244
R5024 gnd.n5811 gnd.n824 240.244
R5025 gnd.n5817 gnd.n824 240.244
R5026 gnd.n5817 gnd.n822 240.244
R5027 gnd.n5821 gnd.n822 240.244
R5028 gnd.n5821 gnd.n818 240.244
R5029 gnd.n5827 gnd.n818 240.244
R5030 gnd.n5827 gnd.n816 240.244
R5031 gnd.n5831 gnd.n816 240.244
R5032 gnd.n5831 gnd.n812 240.244
R5033 gnd.n5837 gnd.n812 240.244
R5034 gnd.n5837 gnd.n810 240.244
R5035 gnd.n5841 gnd.n810 240.244
R5036 gnd.n5841 gnd.n806 240.244
R5037 gnd.n5847 gnd.n806 240.244
R5038 gnd.n5847 gnd.n804 240.244
R5039 gnd.n5851 gnd.n804 240.244
R5040 gnd.n5851 gnd.n800 240.244
R5041 gnd.n5857 gnd.n800 240.244
R5042 gnd.n5857 gnd.n798 240.244
R5043 gnd.n5861 gnd.n798 240.244
R5044 gnd.n5861 gnd.n794 240.244
R5045 gnd.n5867 gnd.n794 240.244
R5046 gnd.n5867 gnd.n792 240.244
R5047 gnd.n5871 gnd.n792 240.244
R5048 gnd.n5871 gnd.n788 240.244
R5049 gnd.n5877 gnd.n788 240.244
R5050 gnd.n5877 gnd.n786 240.244
R5051 gnd.n5881 gnd.n786 240.244
R5052 gnd.n5881 gnd.n782 240.244
R5053 gnd.n5887 gnd.n782 240.244
R5054 gnd.n5887 gnd.n780 240.244
R5055 gnd.n5891 gnd.n780 240.244
R5056 gnd.n5891 gnd.n776 240.244
R5057 gnd.n5897 gnd.n776 240.244
R5058 gnd.n5897 gnd.n774 240.244
R5059 gnd.n5901 gnd.n774 240.244
R5060 gnd.n5901 gnd.n770 240.244
R5061 gnd.n5907 gnd.n770 240.244
R5062 gnd.n5907 gnd.n768 240.244
R5063 gnd.n5911 gnd.n768 240.244
R5064 gnd.n5911 gnd.n764 240.244
R5065 gnd.n5917 gnd.n764 240.244
R5066 gnd.n5917 gnd.n762 240.244
R5067 gnd.n5921 gnd.n762 240.244
R5068 gnd.n5921 gnd.n758 240.244
R5069 gnd.n5927 gnd.n758 240.244
R5070 gnd.n5927 gnd.n756 240.244
R5071 gnd.n5931 gnd.n756 240.244
R5072 gnd.n5931 gnd.n752 240.244
R5073 gnd.n5937 gnd.n752 240.244
R5074 gnd.n5937 gnd.n750 240.244
R5075 gnd.n5941 gnd.n750 240.244
R5076 gnd.n5941 gnd.n746 240.244
R5077 gnd.n5947 gnd.n746 240.244
R5078 gnd.n5947 gnd.n744 240.244
R5079 gnd.n5951 gnd.n744 240.244
R5080 gnd.n5951 gnd.n740 240.244
R5081 gnd.n5957 gnd.n740 240.244
R5082 gnd.n5957 gnd.n738 240.244
R5083 gnd.n5961 gnd.n738 240.244
R5084 gnd.n5961 gnd.n734 240.244
R5085 gnd.n5967 gnd.n734 240.244
R5086 gnd.n5967 gnd.n732 240.244
R5087 gnd.n5971 gnd.n732 240.244
R5088 gnd.n5971 gnd.n728 240.244
R5089 gnd.n5977 gnd.n728 240.244
R5090 gnd.n5977 gnd.n726 240.244
R5091 gnd.n5981 gnd.n726 240.244
R5092 gnd.n5981 gnd.n722 240.244
R5093 gnd.n5987 gnd.n722 240.244
R5094 gnd.n5987 gnd.n720 240.244
R5095 gnd.n5991 gnd.n720 240.244
R5096 gnd.n5991 gnd.n716 240.244
R5097 gnd.n5997 gnd.n716 240.244
R5098 gnd.n5997 gnd.n714 240.244
R5099 gnd.n6001 gnd.n714 240.244
R5100 gnd.n6001 gnd.n710 240.244
R5101 gnd.n6007 gnd.n710 240.244
R5102 gnd.n6007 gnd.n708 240.244
R5103 gnd.n6011 gnd.n708 240.244
R5104 gnd.n6011 gnd.n704 240.244
R5105 gnd.n6017 gnd.n704 240.244
R5106 gnd.n6017 gnd.n702 240.244
R5107 gnd.n6021 gnd.n702 240.244
R5108 gnd.n6021 gnd.n698 240.244
R5109 gnd.n6027 gnd.n698 240.244
R5110 gnd.n6027 gnd.n696 240.244
R5111 gnd.n6031 gnd.n696 240.244
R5112 gnd.n6031 gnd.n692 240.244
R5113 gnd.n6037 gnd.n692 240.244
R5114 gnd.n6037 gnd.n690 240.244
R5115 gnd.n6041 gnd.n690 240.244
R5116 gnd.n6041 gnd.n686 240.244
R5117 gnd.n6047 gnd.n686 240.244
R5118 gnd.n6047 gnd.n684 240.244
R5119 gnd.n6051 gnd.n684 240.244
R5120 gnd.n6051 gnd.n680 240.244
R5121 gnd.n6057 gnd.n680 240.244
R5122 gnd.n6057 gnd.n678 240.244
R5123 gnd.n6061 gnd.n678 240.244
R5124 gnd.n6061 gnd.n674 240.244
R5125 gnd.n6067 gnd.n674 240.244
R5126 gnd.n6067 gnd.n672 240.244
R5127 gnd.n6071 gnd.n672 240.244
R5128 gnd.n6071 gnd.n668 240.244
R5129 gnd.n6077 gnd.n668 240.244
R5130 gnd.n6077 gnd.n666 240.244
R5131 gnd.n6081 gnd.n666 240.244
R5132 gnd.n6081 gnd.n662 240.244
R5133 gnd.n6087 gnd.n662 240.244
R5134 gnd.n6087 gnd.n660 240.244
R5135 gnd.n6091 gnd.n660 240.244
R5136 gnd.n6091 gnd.n656 240.244
R5137 gnd.n6097 gnd.n656 240.244
R5138 gnd.n6097 gnd.n654 240.244
R5139 gnd.n6101 gnd.n654 240.244
R5140 gnd.n6101 gnd.n650 240.244
R5141 gnd.n6107 gnd.n650 240.244
R5142 gnd.n6107 gnd.n648 240.244
R5143 gnd.n6111 gnd.n648 240.244
R5144 gnd.n6117 gnd.n644 240.244
R5145 gnd.n6117 gnd.n642 240.244
R5146 gnd.n6121 gnd.n642 240.244
R5147 gnd.n6121 gnd.n638 240.244
R5148 gnd.n6127 gnd.n638 240.244
R5149 gnd.n6127 gnd.n636 240.244
R5150 gnd.n6131 gnd.n636 240.244
R5151 gnd.n6131 gnd.n632 240.244
R5152 gnd.n6137 gnd.n632 240.244
R5153 gnd.n6137 gnd.n630 240.244
R5154 gnd.n6141 gnd.n630 240.244
R5155 gnd.n6141 gnd.n626 240.244
R5156 gnd.n6147 gnd.n626 240.244
R5157 gnd.n6147 gnd.n624 240.244
R5158 gnd.n6151 gnd.n624 240.244
R5159 gnd.n6151 gnd.n620 240.244
R5160 gnd.n6157 gnd.n620 240.244
R5161 gnd.n6157 gnd.n618 240.244
R5162 gnd.n6161 gnd.n618 240.244
R5163 gnd.n6161 gnd.n614 240.244
R5164 gnd.n6167 gnd.n614 240.244
R5165 gnd.n6167 gnd.n612 240.244
R5166 gnd.n6171 gnd.n612 240.244
R5167 gnd.n6171 gnd.n608 240.244
R5168 gnd.n6177 gnd.n608 240.244
R5169 gnd.n6177 gnd.n606 240.244
R5170 gnd.n6181 gnd.n606 240.244
R5171 gnd.n6181 gnd.n602 240.244
R5172 gnd.n6187 gnd.n602 240.244
R5173 gnd.n6187 gnd.n600 240.244
R5174 gnd.n6191 gnd.n600 240.244
R5175 gnd.n6191 gnd.n596 240.244
R5176 gnd.n6197 gnd.n596 240.244
R5177 gnd.n6197 gnd.n594 240.244
R5178 gnd.n6201 gnd.n594 240.244
R5179 gnd.n6201 gnd.n590 240.244
R5180 gnd.n6207 gnd.n590 240.244
R5181 gnd.n6207 gnd.n588 240.244
R5182 gnd.n6211 gnd.n588 240.244
R5183 gnd.n6211 gnd.n584 240.244
R5184 gnd.n6217 gnd.n584 240.244
R5185 gnd.n6217 gnd.n582 240.244
R5186 gnd.n6221 gnd.n582 240.244
R5187 gnd.n6221 gnd.n578 240.244
R5188 gnd.n6227 gnd.n578 240.244
R5189 gnd.n6227 gnd.n576 240.244
R5190 gnd.n6231 gnd.n576 240.244
R5191 gnd.n6231 gnd.n572 240.244
R5192 gnd.n6237 gnd.n572 240.244
R5193 gnd.n6237 gnd.n570 240.244
R5194 gnd.n6241 gnd.n570 240.244
R5195 gnd.n6241 gnd.n566 240.244
R5196 gnd.n6247 gnd.n566 240.244
R5197 gnd.n6247 gnd.n564 240.244
R5198 gnd.n6251 gnd.n564 240.244
R5199 gnd.n6251 gnd.n560 240.244
R5200 gnd.n6257 gnd.n560 240.244
R5201 gnd.n6257 gnd.n558 240.244
R5202 gnd.n6261 gnd.n558 240.244
R5203 gnd.n6261 gnd.n554 240.244
R5204 gnd.n6267 gnd.n554 240.244
R5205 gnd.n6267 gnd.n552 240.244
R5206 gnd.n6271 gnd.n552 240.244
R5207 gnd.n6271 gnd.n548 240.244
R5208 gnd.n6277 gnd.n548 240.244
R5209 gnd.n6277 gnd.n546 240.244
R5210 gnd.n6281 gnd.n546 240.244
R5211 gnd.n6281 gnd.n542 240.244
R5212 gnd.n6287 gnd.n542 240.244
R5213 gnd.n6287 gnd.n540 240.244
R5214 gnd.n6291 gnd.n540 240.244
R5215 gnd.n6291 gnd.n536 240.244
R5216 gnd.n6297 gnd.n536 240.244
R5217 gnd.n6297 gnd.n534 240.244
R5218 gnd.n6301 gnd.n534 240.244
R5219 gnd.n6301 gnd.n530 240.244
R5220 gnd.n6307 gnd.n530 240.244
R5221 gnd.n6307 gnd.n528 240.244
R5222 gnd.n6311 gnd.n528 240.244
R5223 gnd.n6311 gnd.n524 240.244
R5224 gnd.n6319 gnd.n524 240.244
R5225 gnd.n6319 gnd.n522 240.244
R5226 gnd.n6324 gnd.n522 240.244
R5227 gnd.n6325 gnd.n6324 240.244
R5228 gnd.n2524 gnd.n2518 240.244
R5229 gnd.n2525 gnd.n2524 240.244
R5230 gnd.n2526 gnd.n2525 240.244
R5231 gnd.n2526 gnd.n2514 240.244
R5232 gnd.n2533 gnd.n2514 240.244
R5233 gnd.n2533 gnd.n2249 240.244
R5234 gnd.n2565 gnd.n2249 240.244
R5235 gnd.n2565 gnd.n2250 240.244
R5236 gnd.n2561 gnd.n2250 240.244
R5237 gnd.n2561 gnd.n2560 240.244
R5238 gnd.n2560 gnd.n2256 240.244
R5239 gnd.n2554 gnd.n2256 240.244
R5240 gnd.n2554 gnd.n2546 240.244
R5241 gnd.n2546 gnd.n2070 240.244
R5242 gnd.n2646 gnd.n2070 240.244
R5243 gnd.n2646 gnd.n2065 240.244
R5244 gnd.n2654 gnd.n2065 240.244
R5245 gnd.n2654 gnd.n2066 240.244
R5246 gnd.n2066 gnd.n2045 240.244
R5247 gnd.n2676 gnd.n2045 240.244
R5248 gnd.n2676 gnd.n2040 240.244
R5249 gnd.n2684 gnd.n2040 240.244
R5250 gnd.n2684 gnd.n2041 240.244
R5251 gnd.n2041 gnd.n2020 240.244
R5252 gnd.n2706 gnd.n2020 240.244
R5253 gnd.n2706 gnd.n2015 240.244
R5254 gnd.n2714 gnd.n2015 240.244
R5255 gnd.n2714 gnd.n2016 240.244
R5256 gnd.n2016 gnd.n1995 240.244
R5257 gnd.n2740 gnd.n1995 240.244
R5258 gnd.n2740 gnd.n1990 240.244
R5259 gnd.n2761 gnd.n1990 240.244
R5260 gnd.n2761 gnd.n1991 240.244
R5261 gnd.n2757 gnd.n1991 240.244
R5262 gnd.n2757 gnd.n2755 240.244
R5263 gnd.n2755 gnd.n2754 240.244
R5264 gnd.n2754 gnd.n2748 240.244
R5265 gnd.n2748 gnd.n1964 240.244
R5266 gnd.n2914 gnd.n1964 240.244
R5267 gnd.n2914 gnd.n1959 240.244
R5268 gnd.n2922 gnd.n1959 240.244
R5269 gnd.n2922 gnd.n1960 240.244
R5270 gnd.n1960 gnd.n1937 240.244
R5271 gnd.n2951 gnd.n1937 240.244
R5272 gnd.n2951 gnd.n1933 240.244
R5273 gnd.n2957 gnd.n1933 240.244
R5274 gnd.n2957 gnd.n1916 240.244
R5275 gnd.n2981 gnd.n1916 240.244
R5276 gnd.n2981 gnd.n1911 240.244
R5277 gnd.n2989 gnd.n1911 240.244
R5278 gnd.n2989 gnd.n1912 240.244
R5279 gnd.n1912 gnd.n1886 240.244
R5280 gnd.n3032 gnd.n1886 240.244
R5281 gnd.n3032 gnd.n1882 240.244
R5282 gnd.n3040 gnd.n1882 240.244
R5283 gnd.n3040 gnd.n1867 240.244
R5284 gnd.n3059 gnd.n1867 240.244
R5285 gnd.n3060 gnd.n3059 240.244
R5286 gnd.n3060 gnd.n1863 240.244
R5287 gnd.n3066 gnd.n1863 240.244
R5288 gnd.n3066 gnd.n1839 240.244
R5289 gnd.n3116 gnd.n1839 240.244
R5290 gnd.n3116 gnd.n1835 240.244
R5291 gnd.n3122 gnd.n1835 240.244
R5292 gnd.n3122 gnd.n1816 240.244
R5293 gnd.n3156 gnd.n1816 240.244
R5294 gnd.n3156 gnd.n1812 240.244
R5295 gnd.n3162 gnd.n1812 240.244
R5296 gnd.n3162 gnd.n1793 240.244
R5297 gnd.n3196 gnd.n1793 240.244
R5298 gnd.n3196 gnd.n1789 240.244
R5299 gnd.n3202 gnd.n1789 240.244
R5300 gnd.n3202 gnd.n1771 240.244
R5301 gnd.n3243 gnd.n1771 240.244
R5302 gnd.n3243 gnd.n1767 240.244
R5303 gnd.n3249 gnd.n1767 240.244
R5304 gnd.n3249 gnd.n1753 240.244
R5305 gnd.n3270 gnd.n1753 240.244
R5306 gnd.n3270 gnd.n1748 240.244
R5307 gnd.n3281 gnd.n1748 240.244
R5308 gnd.n3281 gnd.n1749 240.244
R5309 gnd.n3277 gnd.n1749 240.244
R5310 gnd.n3277 gnd.n1717 240.244
R5311 gnd.n3337 gnd.n1717 240.244
R5312 gnd.n3337 gnd.n1712 240.244
R5313 gnd.n3345 gnd.n1712 240.244
R5314 gnd.n3345 gnd.n1713 240.244
R5315 gnd.n1713 gnd.n1690 240.244
R5316 gnd.n3388 gnd.n1690 240.244
R5317 gnd.n3388 gnd.n1685 240.244
R5318 gnd.n3399 gnd.n1685 240.244
R5319 gnd.n3399 gnd.n1686 240.244
R5320 gnd.n3395 gnd.n1686 240.244
R5321 gnd.n3395 gnd.n1629 240.244
R5322 gnd.n3576 gnd.n1629 240.244
R5323 gnd.n3576 gnd.n1625 240.244
R5324 gnd.n3582 gnd.n1625 240.244
R5325 gnd.n3582 gnd.n1618 240.244
R5326 gnd.n3598 gnd.n1618 240.244
R5327 gnd.n3598 gnd.n1614 240.244
R5328 gnd.n3604 gnd.n1614 240.244
R5329 gnd.n3604 gnd.n1606 240.244
R5330 gnd.n3619 gnd.n1606 240.244
R5331 gnd.n3619 gnd.n1602 240.244
R5332 gnd.n3625 gnd.n1602 240.244
R5333 gnd.n3625 gnd.n1594 240.244
R5334 gnd.n3640 gnd.n1594 240.244
R5335 gnd.n3640 gnd.n1590 240.244
R5336 gnd.n3646 gnd.n1590 240.244
R5337 gnd.n3646 gnd.n1581 240.244
R5338 gnd.n3661 gnd.n1581 240.244
R5339 gnd.n3661 gnd.n1576 240.244
R5340 gnd.n3673 gnd.n1576 240.244
R5341 gnd.n3673 gnd.n1577 240.244
R5342 gnd.n3669 gnd.n1577 240.244
R5343 gnd.n3669 gnd.n491 240.244
R5344 gnd.n6353 gnd.n491 240.244
R5345 gnd.n6353 gnd.n492 240.244
R5346 gnd.n6349 gnd.n492 240.244
R5347 gnd.n6349 gnd.n6348 240.244
R5348 gnd.n6348 gnd.n6347 240.244
R5349 gnd.n6347 gnd.n498 240.244
R5350 gnd.n6337 gnd.n498 240.244
R5351 gnd.n6337 gnd.n507 240.244
R5352 gnd.n6333 gnd.n507 240.244
R5353 gnd.n6333 gnd.n6332 240.244
R5354 gnd.n6332 gnd.n6331 240.244
R5355 gnd.n6331 gnd.n517 240.244
R5356 gnd.n5787 gnd.n839 240.244
R5357 gnd.n5787 gnd.n841 240.244
R5358 gnd.n5783 gnd.n841 240.244
R5359 gnd.n5783 gnd.n847 240.244
R5360 gnd.n5779 gnd.n847 240.244
R5361 gnd.n5779 gnd.n849 240.244
R5362 gnd.n5775 gnd.n849 240.244
R5363 gnd.n5775 gnd.n855 240.244
R5364 gnd.n5771 gnd.n855 240.244
R5365 gnd.n5771 gnd.n857 240.244
R5366 gnd.n5767 gnd.n857 240.244
R5367 gnd.n5767 gnd.n863 240.244
R5368 gnd.n5763 gnd.n863 240.244
R5369 gnd.n5763 gnd.n865 240.244
R5370 gnd.n5759 gnd.n865 240.244
R5371 gnd.n5759 gnd.n871 240.244
R5372 gnd.n5755 gnd.n871 240.244
R5373 gnd.n5755 gnd.n873 240.244
R5374 gnd.n5751 gnd.n873 240.244
R5375 gnd.n5751 gnd.n879 240.244
R5376 gnd.n5747 gnd.n879 240.244
R5377 gnd.n5747 gnd.n881 240.244
R5378 gnd.n5743 gnd.n881 240.244
R5379 gnd.n5743 gnd.n887 240.244
R5380 gnd.n5739 gnd.n887 240.244
R5381 gnd.n5739 gnd.n889 240.244
R5382 gnd.n5735 gnd.n889 240.244
R5383 gnd.n5735 gnd.n895 240.244
R5384 gnd.n5731 gnd.n895 240.244
R5385 gnd.n5731 gnd.n897 240.244
R5386 gnd.n5727 gnd.n897 240.244
R5387 gnd.n5727 gnd.n903 240.244
R5388 gnd.n5723 gnd.n903 240.244
R5389 gnd.n5723 gnd.n905 240.244
R5390 gnd.n5719 gnd.n905 240.244
R5391 gnd.n5719 gnd.n911 240.244
R5392 gnd.n5715 gnd.n911 240.244
R5393 gnd.n5715 gnd.n913 240.244
R5394 gnd.n5711 gnd.n913 240.244
R5395 gnd.n5711 gnd.n919 240.244
R5396 gnd.n5707 gnd.n919 240.244
R5397 gnd.n5707 gnd.n921 240.244
R5398 gnd.n5703 gnd.n921 240.244
R5399 gnd.n5703 gnd.n927 240.244
R5400 gnd.n5699 gnd.n927 240.244
R5401 gnd.n5699 gnd.n929 240.244
R5402 gnd.n5695 gnd.n929 240.244
R5403 gnd.n5695 gnd.n935 240.244
R5404 gnd.n5691 gnd.n935 240.244
R5405 gnd.n5691 gnd.n937 240.244
R5406 gnd.n5687 gnd.n937 240.244
R5407 gnd.n5687 gnd.n943 240.244
R5408 gnd.n5683 gnd.n943 240.244
R5409 gnd.n5683 gnd.n945 240.244
R5410 gnd.n5679 gnd.n945 240.244
R5411 gnd.n5679 gnd.n951 240.244
R5412 gnd.n5675 gnd.n951 240.244
R5413 gnd.n5675 gnd.n953 240.244
R5414 gnd.n5671 gnd.n953 240.244
R5415 gnd.n5671 gnd.n959 240.244
R5416 gnd.n5667 gnd.n959 240.244
R5417 gnd.n5667 gnd.n961 240.244
R5418 gnd.n5663 gnd.n961 240.244
R5419 gnd.n5663 gnd.n967 240.244
R5420 gnd.n5659 gnd.n967 240.244
R5421 gnd.n5659 gnd.n969 240.244
R5422 gnd.n5655 gnd.n969 240.244
R5423 gnd.n5655 gnd.n975 240.244
R5424 gnd.n5651 gnd.n975 240.244
R5425 gnd.n5651 gnd.n977 240.244
R5426 gnd.n5647 gnd.n977 240.244
R5427 gnd.n5647 gnd.n983 240.244
R5428 gnd.n5643 gnd.n983 240.244
R5429 gnd.n5643 gnd.n985 240.244
R5430 gnd.n5639 gnd.n985 240.244
R5431 gnd.n5639 gnd.n991 240.244
R5432 gnd.n5635 gnd.n991 240.244
R5433 gnd.n5635 gnd.n993 240.244
R5434 gnd.n5631 gnd.n993 240.244
R5435 gnd.n5631 gnd.n999 240.244
R5436 gnd.n5627 gnd.n999 240.244
R5437 gnd.n5627 gnd.n1001 240.244
R5438 gnd.n5623 gnd.n1001 240.244
R5439 gnd.n5623 gnd.n1007 240.244
R5440 gnd.n2634 gnd.n2080 240.244
R5441 gnd.n2080 gnd.n2061 240.244
R5442 gnd.n2657 gnd.n2061 240.244
R5443 gnd.n2657 gnd.n2055 240.244
R5444 gnd.n2664 gnd.n2055 240.244
R5445 gnd.n2664 gnd.n2056 240.244
R5446 gnd.n2056 gnd.n2036 240.244
R5447 gnd.n2687 gnd.n2036 240.244
R5448 gnd.n2687 gnd.n2029 240.244
R5449 gnd.n2694 gnd.n2029 240.244
R5450 gnd.n2694 gnd.n2031 240.244
R5451 gnd.n2031 gnd.n2011 240.244
R5452 gnd.n2717 gnd.n2011 240.244
R5453 gnd.n2717 gnd.n2005 240.244
R5454 gnd.n2724 gnd.n2005 240.244
R5455 gnd.n2724 gnd.n2006 240.244
R5456 gnd.n2006 gnd.n1986 240.244
R5457 gnd.n2764 gnd.n1986 240.244
R5458 gnd.n2764 gnd.n1980 240.244
R5459 gnd.n2771 gnd.n1980 240.244
R5460 gnd.n2771 gnd.n1981 240.244
R5461 gnd.n1981 gnd.n1475 240.244
R5462 gnd.n3793 gnd.n1475 240.244
R5463 gnd.n3793 gnd.n1476 240.244
R5464 gnd.n1481 gnd.n1476 240.244
R5465 gnd.n1482 gnd.n1481 240.244
R5466 gnd.n1483 gnd.n1482 240.244
R5467 gnd.n2931 gnd.n1483 240.244
R5468 gnd.n2931 gnd.n1486 240.244
R5469 gnd.n1487 gnd.n1486 240.244
R5470 gnd.n1488 gnd.n1487 240.244
R5471 gnd.n2960 gnd.n1488 240.244
R5472 gnd.n2960 gnd.n1491 240.244
R5473 gnd.n1492 gnd.n1491 240.244
R5474 gnd.n1493 gnd.n1492 240.244
R5475 gnd.n2991 gnd.n1493 240.244
R5476 gnd.n2991 gnd.n1496 240.244
R5477 gnd.n1497 gnd.n1496 240.244
R5478 gnd.n1498 gnd.n1497 240.244
R5479 gnd.n1889 gnd.n1498 240.244
R5480 gnd.n1889 gnd.n1501 240.244
R5481 gnd.n1502 gnd.n1501 240.244
R5482 gnd.n1503 gnd.n1502 240.244
R5483 gnd.n3056 gnd.n1503 240.244
R5484 gnd.n3056 gnd.n1506 240.244
R5485 gnd.n1507 gnd.n1506 240.244
R5486 gnd.n1508 gnd.n1507 240.244
R5487 gnd.n3102 gnd.n1508 240.244
R5488 gnd.n3102 gnd.n1511 240.244
R5489 gnd.n1512 gnd.n1511 240.244
R5490 gnd.n1513 gnd.n1512 240.244
R5491 gnd.n3143 gnd.n1513 240.244
R5492 gnd.n3143 gnd.n1516 240.244
R5493 gnd.n1517 gnd.n1516 240.244
R5494 gnd.n1518 gnd.n1517 240.244
R5495 gnd.n3183 gnd.n1518 240.244
R5496 gnd.n3183 gnd.n1521 240.244
R5497 gnd.n1522 gnd.n1521 240.244
R5498 gnd.n1523 gnd.n1522 240.244
R5499 gnd.n3232 gnd.n1523 240.244
R5500 gnd.n3232 gnd.n1526 240.244
R5501 gnd.n1527 gnd.n1526 240.244
R5502 gnd.n1528 gnd.n1527 240.244
R5503 gnd.n1760 gnd.n1528 240.244
R5504 gnd.n1760 gnd.n1531 240.244
R5505 gnd.n1532 gnd.n1531 240.244
R5506 gnd.n1533 gnd.n1532 240.244
R5507 gnd.n1739 gnd.n1533 240.244
R5508 gnd.n1739 gnd.n1536 240.244
R5509 gnd.n1537 gnd.n1536 240.244
R5510 gnd.n1538 gnd.n1537 240.244
R5511 gnd.n3347 gnd.n1538 240.244
R5512 gnd.n3347 gnd.n1541 240.244
R5513 gnd.n1542 gnd.n1541 240.244
R5514 gnd.n1543 gnd.n1542 240.244
R5515 gnd.n1694 gnd.n1543 240.244
R5516 gnd.n1694 gnd.n1546 240.244
R5517 gnd.n1547 gnd.n1546 240.244
R5518 gnd.n1548 gnd.n1547 240.244
R5519 gnd.n3564 gnd.n1548 240.244
R5520 gnd.n3564 gnd.n1551 240.244
R5521 gnd.n1552 gnd.n1551 240.244
R5522 gnd.n1553 gnd.n1552 240.244
R5523 gnd.n3586 gnd.n1553 240.244
R5524 gnd.n3586 gnd.n1556 240.244
R5525 gnd.n1557 gnd.n1556 240.244
R5526 gnd.n1558 gnd.n1557 240.244
R5527 gnd.n3607 gnd.n1558 240.244
R5528 gnd.n3607 gnd.n1561 240.244
R5529 gnd.n1562 gnd.n1561 240.244
R5530 gnd.n1563 gnd.n1562 240.244
R5531 gnd.n3628 gnd.n1563 240.244
R5532 gnd.n3628 gnd.n1566 240.244
R5533 gnd.n1567 gnd.n1566 240.244
R5534 gnd.n1568 gnd.n1567 240.244
R5535 gnd.n3649 gnd.n1568 240.244
R5536 gnd.n3649 gnd.n1571 240.244
R5537 gnd.n1572 gnd.n1571 240.244
R5538 gnd.n3676 gnd.n1572 240.244
R5539 gnd.n3676 gnd.n459 240.244
R5540 gnd.n6370 gnd.n459 240.244
R5541 gnd.n2084 gnd.n2083 240.244
R5542 gnd.n2257 gnd.n2084 240.244
R5543 gnd.n2088 gnd.n2087 240.244
R5544 gnd.n2260 gnd.n2089 240.244
R5545 gnd.n2094 gnd.n2093 240.244
R5546 gnd.n2262 gnd.n2103 240.244
R5547 gnd.n2265 gnd.n2104 240.244
R5548 gnd.n2112 gnd.n2111 240.244
R5549 gnd.n2267 gnd.n2121 240.244
R5550 gnd.n2270 gnd.n2122 240.244
R5551 gnd.n2130 gnd.n2129 240.244
R5552 gnd.n2272 gnd.n2139 240.244
R5553 gnd.n2277 gnd.n2140 240.244
R5554 gnd.n2544 gnd.n2276 240.244
R5555 gnd.n2636 gnd.n2072 240.244
R5556 gnd.n2643 gnd.n2072 240.244
R5557 gnd.n2643 gnd.n2063 240.244
R5558 gnd.n2063 gnd.n2052 240.244
R5559 gnd.n2666 gnd.n2052 240.244
R5560 gnd.n2666 gnd.n2047 240.244
R5561 gnd.n2673 gnd.n2047 240.244
R5562 gnd.n2673 gnd.n2038 240.244
R5563 gnd.n2038 gnd.n2026 240.244
R5564 gnd.n2696 gnd.n2026 240.244
R5565 gnd.n2696 gnd.n2021 240.244
R5566 gnd.n2703 gnd.n2021 240.244
R5567 gnd.n2703 gnd.n2013 240.244
R5568 gnd.n2013 gnd.n2002 240.244
R5569 gnd.n2726 gnd.n2002 240.244
R5570 gnd.n2726 gnd.n1997 240.244
R5571 gnd.n2737 gnd.n1997 240.244
R5572 gnd.n2737 gnd.n1988 240.244
R5573 gnd.n1988 gnd.n1977 240.244
R5574 gnd.n2773 gnd.n1977 240.244
R5575 gnd.n2774 gnd.n2773 240.244
R5576 gnd.n2895 gnd.n2774 240.244
R5577 gnd.n2895 gnd.n1473 240.244
R5578 gnd.n1971 gnd.n1473 240.244
R5579 gnd.n2903 gnd.n1971 240.244
R5580 gnd.n2903 gnd.n1972 240.244
R5581 gnd.n1972 gnd.n1950 240.244
R5582 gnd.n2933 gnd.n1950 240.244
R5583 gnd.n2933 gnd.n1946 240.244
R5584 gnd.n2939 gnd.n1946 240.244
R5585 gnd.n2939 gnd.n1931 240.244
R5586 gnd.n2962 gnd.n1931 240.244
R5587 gnd.n2962 gnd.n1925 240.244
R5588 gnd.n2969 gnd.n1925 240.244
R5589 gnd.n2969 gnd.n1926 240.244
R5590 gnd.n1926 gnd.n1902 240.244
R5591 gnd.n3001 gnd.n1902 240.244
R5592 gnd.n3001 gnd.n1896 240.244
R5593 gnd.n3022 gnd.n1896 240.244
R5594 gnd.n3022 gnd.n1897 240.244
R5595 gnd.n3006 gnd.n1897 240.244
R5596 gnd.n3007 gnd.n3006 240.244
R5597 gnd.n3008 gnd.n3007 240.244
R5598 gnd.n3008 gnd.n1869 240.244
R5599 gnd.n1869 gnd.n1854 240.244
R5600 gnd.n3084 gnd.n1854 240.244
R5601 gnd.n3085 gnd.n3084 240.244
R5602 gnd.n3085 gnd.n1848 240.244
R5603 gnd.n1850 gnd.n1848 240.244
R5604 gnd.n3092 gnd.n1850 240.244
R5605 gnd.n3092 gnd.n1826 240.244
R5606 gnd.n3142 gnd.n1826 240.244
R5607 gnd.n3142 gnd.n1827 240.244
R5608 gnd.n3136 gnd.n1827 240.244
R5609 gnd.n3136 gnd.n1803 240.244
R5610 gnd.n3182 gnd.n1803 240.244
R5611 gnd.n3182 gnd.n1804 240.244
R5612 gnd.n3176 gnd.n1804 240.244
R5613 gnd.n3176 gnd.n1781 240.244
R5614 gnd.n3231 gnd.n1781 240.244
R5615 gnd.n3231 gnd.n1773 240.244
R5616 gnd.n3216 gnd.n1773 240.244
R5617 gnd.n3219 gnd.n3216 240.244
R5618 gnd.n3220 gnd.n3219 240.244
R5619 gnd.n3220 gnd.n1755 240.244
R5620 gnd.n1755 gnd.n1735 240.244
R5621 gnd.n3294 gnd.n1735 240.244
R5622 gnd.n3294 gnd.n1729 240.244
R5623 gnd.n3301 gnd.n1729 240.244
R5624 gnd.n3301 gnd.n1730 240.244
R5625 gnd.n1730 gnd.n1709 240.244
R5626 gnd.n3349 gnd.n1709 240.244
R5627 gnd.n3349 gnd.n1704 240.244
R5628 gnd.n3364 gnd.n1704 240.244
R5629 gnd.n3364 gnd.n1700 240.244
R5630 gnd.n1700 gnd.n1692 240.244
R5631 gnd.n3354 gnd.n1692 240.244
R5632 gnd.n3355 gnd.n3354 240.244
R5633 gnd.n3355 gnd.n1635 240.244
R5634 gnd.n3566 gnd.n1635 240.244
R5635 gnd.n3566 gnd.n1631 240.244
R5636 gnd.n3572 gnd.n1631 240.244
R5637 gnd.n3572 gnd.n1623 240.244
R5638 gnd.n3588 gnd.n1623 240.244
R5639 gnd.n3588 gnd.n1619 240.244
R5640 gnd.n3594 gnd.n1619 240.244
R5641 gnd.n3594 gnd.n1612 240.244
R5642 gnd.n3609 gnd.n1612 240.244
R5643 gnd.n3609 gnd.n1608 240.244
R5644 gnd.n3615 gnd.n1608 240.244
R5645 gnd.n3615 gnd.n1600 240.244
R5646 gnd.n3630 gnd.n1600 240.244
R5647 gnd.n3630 gnd.n1596 240.244
R5648 gnd.n3636 gnd.n1596 240.244
R5649 gnd.n3636 gnd.n1588 240.244
R5650 gnd.n3651 gnd.n1588 240.244
R5651 gnd.n3651 gnd.n1583 240.244
R5652 gnd.n3658 gnd.n1583 240.244
R5653 gnd.n3658 gnd.n1574 240.244
R5654 gnd.n1574 gnd.n455 240.244
R5655 gnd.n6372 gnd.n455 240.244
R5656 gnd.n465 gnd.n464 240.244
R5657 gnd.n472 gnd.n468 240.244
R5658 gnd.n6358 gnd.n6357 240.244
R5659 gnd.n393 gnd.n392 240.244
R5660 gnd.n475 gnd.n394 240.244
R5661 gnd.n404 gnd.n403 240.244
R5662 gnd.n477 gnd.n413 240.244
R5663 gnd.n480 gnd.n414 240.244
R5664 gnd.n422 gnd.n421 240.244
R5665 gnd.n482 gnd.n431 240.244
R5666 gnd.n485 gnd.n432 240.244
R5667 gnd.n440 gnd.n439 240.244
R5668 gnd.n487 gnd.n440 240.244
R5669 gnd.n451 gnd.n450 240.244
R5670 gnd.n1455 gnd.n1454 240.132
R5671 gnd.n3416 gnd.n3415 240.132
R5672 gnd.n5790 gnd.n835 225.874
R5673 gnd.n5798 gnd.n835 225.874
R5674 gnd.n5799 gnd.n5798 225.874
R5675 gnd.n5800 gnd.n5799 225.874
R5676 gnd.n5800 gnd.n829 225.874
R5677 gnd.n5808 gnd.n829 225.874
R5678 gnd.n5809 gnd.n5808 225.874
R5679 gnd.n5810 gnd.n5809 225.874
R5680 gnd.n5810 gnd.n823 225.874
R5681 gnd.n5818 gnd.n823 225.874
R5682 gnd.n5819 gnd.n5818 225.874
R5683 gnd.n5820 gnd.n5819 225.874
R5684 gnd.n5820 gnd.n817 225.874
R5685 gnd.n5828 gnd.n817 225.874
R5686 gnd.n5829 gnd.n5828 225.874
R5687 gnd.n5830 gnd.n5829 225.874
R5688 gnd.n5830 gnd.n811 225.874
R5689 gnd.n5838 gnd.n811 225.874
R5690 gnd.n5839 gnd.n5838 225.874
R5691 gnd.n5840 gnd.n5839 225.874
R5692 gnd.n5840 gnd.n805 225.874
R5693 gnd.n5848 gnd.n805 225.874
R5694 gnd.n5849 gnd.n5848 225.874
R5695 gnd.n5850 gnd.n5849 225.874
R5696 gnd.n5850 gnd.n799 225.874
R5697 gnd.n5858 gnd.n799 225.874
R5698 gnd.n5859 gnd.n5858 225.874
R5699 gnd.n5860 gnd.n5859 225.874
R5700 gnd.n5860 gnd.n793 225.874
R5701 gnd.n5868 gnd.n793 225.874
R5702 gnd.n5869 gnd.n5868 225.874
R5703 gnd.n5870 gnd.n5869 225.874
R5704 gnd.n5870 gnd.n787 225.874
R5705 gnd.n5878 gnd.n787 225.874
R5706 gnd.n5879 gnd.n5878 225.874
R5707 gnd.n5880 gnd.n5879 225.874
R5708 gnd.n5880 gnd.n781 225.874
R5709 gnd.n5888 gnd.n781 225.874
R5710 gnd.n5889 gnd.n5888 225.874
R5711 gnd.n5890 gnd.n5889 225.874
R5712 gnd.n5890 gnd.n775 225.874
R5713 gnd.n5898 gnd.n775 225.874
R5714 gnd.n5899 gnd.n5898 225.874
R5715 gnd.n5900 gnd.n5899 225.874
R5716 gnd.n5900 gnd.n769 225.874
R5717 gnd.n5908 gnd.n769 225.874
R5718 gnd.n5909 gnd.n5908 225.874
R5719 gnd.n5910 gnd.n5909 225.874
R5720 gnd.n5910 gnd.n763 225.874
R5721 gnd.n5918 gnd.n763 225.874
R5722 gnd.n5919 gnd.n5918 225.874
R5723 gnd.n5920 gnd.n5919 225.874
R5724 gnd.n5920 gnd.n757 225.874
R5725 gnd.n5928 gnd.n757 225.874
R5726 gnd.n5929 gnd.n5928 225.874
R5727 gnd.n5930 gnd.n5929 225.874
R5728 gnd.n5930 gnd.n751 225.874
R5729 gnd.n5938 gnd.n751 225.874
R5730 gnd.n5939 gnd.n5938 225.874
R5731 gnd.n5940 gnd.n5939 225.874
R5732 gnd.n5940 gnd.n745 225.874
R5733 gnd.n5948 gnd.n745 225.874
R5734 gnd.n5949 gnd.n5948 225.874
R5735 gnd.n5950 gnd.n5949 225.874
R5736 gnd.n5950 gnd.n739 225.874
R5737 gnd.n5958 gnd.n739 225.874
R5738 gnd.n5959 gnd.n5958 225.874
R5739 gnd.n5960 gnd.n5959 225.874
R5740 gnd.n5960 gnd.n733 225.874
R5741 gnd.n5968 gnd.n733 225.874
R5742 gnd.n5969 gnd.n5968 225.874
R5743 gnd.n5970 gnd.n5969 225.874
R5744 gnd.n5970 gnd.n727 225.874
R5745 gnd.n5978 gnd.n727 225.874
R5746 gnd.n5979 gnd.n5978 225.874
R5747 gnd.n5980 gnd.n5979 225.874
R5748 gnd.n5980 gnd.n721 225.874
R5749 gnd.n5988 gnd.n721 225.874
R5750 gnd.n5989 gnd.n5988 225.874
R5751 gnd.n5990 gnd.n5989 225.874
R5752 gnd.n5990 gnd.n715 225.874
R5753 gnd.n5998 gnd.n715 225.874
R5754 gnd.n5999 gnd.n5998 225.874
R5755 gnd.n6000 gnd.n5999 225.874
R5756 gnd.n6000 gnd.n709 225.874
R5757 gnd.n6008 gnd.n709 225.874
R5758 gnd.n6009 gnd.n6008 225.874
R5759 gnd.n6010 gnd.n6009 225.874
R5760 gnd.n6010 gnd.n703 225.874
R5761 gnd.n6018 gnd.n703 225.874
R5762 gnd.n6019 gnd.n6018 225.874
R5763 gnd.n6020 gnd.n6019 225.874
R5764 gnd.n6020 gnd.n697 225.874
R5765 gnd.n6028 gnd.n697 225.874
R5766 gnd.n6029 gnd.n6028 225.874
R5767 gnd.n6030 gnd.n6029 225.874
R5768 gnd.n6030 gnd.n691 225.874
R5769 gnd.n6038 gnd.n691 225.874
R5770 gnd.n6039 gnd.n6038 225.874
R5771 gnd.n6040 gnd.n6039 225.874
R5772 gnd.n6040 gnd.n685 225.874
R5773 gnd.n6048 gnd.n685 225.874
R5774 gnd.n6049 gnd.n6048 225.874
R5775 gnd.n6050 gnd.n6049 225.874
R5776 gnd.n6050 gnd.n679 225.874
R5777 gnd.n6058 gnd.n679 225.874
R5778 gnd.n6059 gnd.n6058 225.874
R5779 gnd.n6060 gnd.n6059 225.874
R5780 gnd.n6060 gnd.n673 225.874
R5781 gnd.n6068 gnd.n673 225.874
R5782 gnd.n6069 gnd.n6068 225.874
R5783 gnd.n6070 gnd.n6069 225.874
R5784 gnd.n6070 gnd.n667 225.874
R5785 gnd.n6078 gnd.n667 225.874
R5786 gnd.n6079 gnd.n6078 225.874
R5787 gnd.n6080 gnd.n6079 225.874
R5788 gnd.n6080 gnd.n661 225.874
R5789 gnd.n6088 gnd.n661 225.874
R5790 gnd.n6089 gnd.n6088 225.874
R5791 gnd.n6090 gnd.n6089 225.874
R5792 gnd.n6090 gnd.n655 225.874
R5793 gnd.n6098 gnd.n655 225.874
R5794 gnd.n6099 gnd.n6098 225.874
R5795 gnd.n6100 gnd.n6099 225.874
R5796 gnd.n6100 gnd.n649 225.874
R5797 gnd.n6108 gnd.n649 225.874
R5798 gnd.n6109 gnd.n6108 225.874
R5799 gnd.n6110 gnd.n6109 225.874
R5800 gnd.n4714 gnd.t170 224.174
R5801 gnd.n4224 gnd.t78 224.174
R5802 gnd.n352 gnd.n296 199.319
R5803 gnd.n352 gnd.n297 199.319
R5804 gnd.n1407 gnd.n1367 199.319
R5805 gnd.n1407 gnd.n1366 199.319
R5806 gnd.n1456 gnd.n1453 186.49
R5807 gnd.n3417 gnd.n3414 186.49
R5808 gnd.n5489 gnd.n5488 185
R5809 gnd.n5487 gnd.n5486 185
R5810 gnd.n5466 gnd.n5465 185
R5811 gnd.n5481 gnd.n5480 185
R5812 gnd.n5479 gnd.n5478 185
R5813 gnd.n5470 gnd.n5469 185
R5814 gnd.n5473 gnd.n5472 185
R5815 gnd.n5457 gnd.n5456 185
R5816 gnd.n5455 gnd.n5454 185
R5817 gnd.n5434 gnd.n5433 185
R5818 gnd.n5449 gnd.n5448 185
R5819 gnd.n5447 gnd.n5446 185
R5820 gnd.n5438 gnd.n5437 185
R5821 gnd.n5441 gnd.n5440 185
R5822 gnd.n5425 gnd.n5424 185
R5823 gnd.n5423 gnd.n5422 185
R5824 gnd.n5402 gnd.n5401 185
R5825 gnd.n5417 gnd.n5416 185
R5826 gnd.n5415 gnd.n5414 185
R5827 gnd.n5406 gnd.n5405 185
R5828 gnd.n5409 gnd.n5408 185
R5829 gnd.n5394 gnd.n5393 185
R5830 gnd.n5392 gnd.n5391 185
R5831 gnd.n5371 gnd.n5370 185
R5832 gnd.n5386 gnd.n5385 185
R5833 gnd.n5384 gnd.n5383 185
R5834 gnd.n5375 gnd.n5374 185
R5835 gnd.n5378 gnd.n5377 185
R5836 gnd.n5362 gnd.n5361 185
R5837 gnd.n5360 gnd.n5359 185
R5838 gnd.n5339 gnd.n5338 185
R5839 gnd.n5354 gnd.n5353 185
R5840 gnd.n5352 gnd.n5351 185
R5841 gnd.n5343 gnd.n5342 185
R5842 gnd.n5346 gnd.n5345 185
R5843 gnd.n5330 gnd.n5329 185
R5844 gnd.n5328 gnd.n5327 185
R5845 gnd.n5307 gnd.n5306 185
R5846 gnd.n5322 gnd.n5321 185
R5847 gnd.n5320 gnd.n5319 185
R5848 gnd.n5311 gnd.n5310 185
R5849 gnd.n5314 gnd.n5313 185
R5850 gnd.n5298 gnd.n5297 185
R5851 gnd.n5296 gnd.n5295 185
R5852 gnd.n5275 gnd.n5274 185
R5853 gnd.n5290 gnd.n5289 185
R5854 gnd.n5288 gnd.n5287 185
R5855 gnd.n5279 gnd.n5278 185
R5856 gnd.n5282 gnd.n5281 185
R5857 gnd.n5267 gnd.n5266 185
R5858 gnd.n5265 gnd.n5264 185
R5859 gnd.n5244 gnd.n5243 185
R5860 gnd.n5259 gnd.n5258 185
R5861 gnd.n5257 gnd.n5256 185
R5862 gnd.n5248 gnd.n5247 185
R5863 gnd.n5251 gnd.n5250 185
R5864 gnd.n4715 gnd.t169 178.987
R5865 gnd.n4225 gnd.t79 178.987
R5866 gnd.n1 gnd.t193 170.774
R5867 gnd.n9 gnd.t245 170.103
R5868 gnd.n8 gnd.t322 170.103
R5869 gnd.n7 gnd.t191 170.103
R5870 gnd.n6 gnd.t328 170.103
R5871 gnd.n5 gnd.t251 170.103
R5872 gnd.n4 gnd.t235 170.103
R5873 gnd.n3 gnd.t198 170.103
R5874 gnd.n2 gnd.t313 170.103
R5875 gnd.n1 gnd.t1 170.103
R5876 gnd.n6497 gnd.n351 164.544
R5877 gnd.n3869 gnd.n3868 164.544
R5878 gnd.n3488 gnd.n3487 163.367
R5879 gnd.n3484 gnd.n3483 163.367
R5880 gnd.n3480 gnd.n3479 163.367
R5881 gnd.n3476 gnd.n3475 163.367
R5882 gnd.n3472 gnd.n3471 163.367
R5883 gnd.n3468 gnd.n3467 163.367
R5884 gnd.n3464 gnd.n3463 163.367
R5885 gnd.n3460 gnd.n3459 163.367
R5886 gnd.n3456 gnd.n3455 163.367
R5887 gnd.n3452 gnd.n3451 163.367
R5888 gnd.n3448 gnd.n3447 163.367
R5889 gnd.n3444 gnd.n3443 163.367
R5890 gnd.n3440 gnd.n3439 163.367
R5891 gnd.n3436 gnd.n3435 163.367
R5892 gnd.n3431 gnd.n3430 163.367
R5893 gnd.n3427 gnd.n3426 163.367
R5894 gnd.n3561 gnd.n3560 163.367
R5895 gnd.n3557 gnd.n3556 163.367
R5896 gnd.n3552 gnd.n3551 163.367
R5897 gnd.n3548 gnd.n3547 163.367
R5898 gnd.n3544 gnd.n3543 163.367
R5899 gnd.n3540 gnd.n3539 163.367
R5900 gnd.n3536 gnd.n3535 163.367
R5901 gnd.n3532 gnd.n3531 163.367
R5902 gnd.n3528 gnd.n3527 163.367
R5903 gnd.n3524 gnd.n3523 163.367
R5904 gnd.n3520 gnd.n3519 163.367
R5905 gnd.n3516 gnd.n3515 163.367
R5906 gnd.n3512 gnd.n3511 163.367
R5907 gnd.n3508 gnd.n3507 163.367
R5908 gnd.n3504 gnd.n3503 163.367
R5909 gnd.n3500 gnd.n3499 163.367
R5910 gnd.n2892 gnd.n1472 163.367
R5911 gnd.n2888 gnd.n1472 163.367
R5912 gnd.n2888 gnd.n1969 163.367
R5913 gnd.n1970 gnd.n1969 163.367
R5914 gnd.n1970 gnd.n1965 163.367
R5915 gnd.n2882 gnd.n1965 163.367
R5916 gnd.n2882 gnd.n1958 163.367
R5917 gnd.n2877 gnd.n1958 163.367
R5918 gnd.n2877 gnd.n1952 163.367
R5919 gnd.n2874 gnd.n1952 163.367
R5920 gnd.n2874 gnd.n1945 163.367
R5921 gnd.n2868 gnd.n1945 163.367
R5922 gnd.n2868 gnd.n1939 163.367
R5923 gnd.n2865 gnd.n1939 163.367
R5924 gnd.n2865 gnd.n1932 163.367
R5925 gnd.n1932 gnd.n1923 163.367
R5926 gnd.n1924 gnd.n1923 163.367
R5927 gnd.n1924 gnd.n1917 163.367
R5928 gnd.n2858 gnd.n1917 163.367
R5929 gnd.n2858 gnd.n1910 163.367
R5930 gnd.n2854 gnd.n1910 163.367
R5931 gnd.n2854 gnd.n1904 163.367
R5932 gnd.n2851 gnd.n1904 163.367
R5933 gnd.n2851 gnd.n1895 163.367
R5934 gnd.n2846 gnd.n1895 163.367
R5935 gnd.n2846 gnd.n1888 163.367
R5936 gnd.n2843 gnd.n1888 163.367
R5937 gnd.n2843 gnd.n1880 163.367
R5938 gnd.n1880 gnd.n1872 163.367
R5939 gnd.n3050 gnd.n1872 163.367
R5940 gnd.n3050 gnd.n1870 163.367
R5941 gnd.n3054 gnd.n1870 163.367
R5942 gnd.n3054 gnd.n1861 163.367
R5943 gnd.n3073 gnd.n1861 163.367
R5944 gnd.n3073 gnd.n1856 163.367
R5945 gnd.n3069 gnd.n1856 163.367
R5946 gnd.n3069 gnd.n1847 163.367
R5947 gnd.n3100 gnd.n1847 163.367
R5948 gnd.n3100 gnd.n1840 163.367
R5949 gnd.n3096 gnd.n1840 163.367
R5950 gnd.n3096 gnd.n1833 163.367
R5951 gnd.n3126 gnd.n1833 163.367
R5952 gnd.n3126 gnd.n1825 163.367
R5953 gnd.n3129 gnd.n1825 163.367
R5954 gnd.n3129 gnd.n1818 163.367
R5955 gnd.n3133 gnd.n1818 163.367
R5956 gnd.n3133 gnd.n1810 163.367
R5957 gnd.n3166 gnd.n1810 163.367
R5958 gnd.n3166 gnd.n1802 163.367
R5959 gnd.n3169 gnd.n1802 163.367
R5960 gnd.n3169 gnd.n1795 163.367
R5961 gnd.n3173 gnd.n1795 163.367
R5962 gnd.n3173 gnd.n1787 163.367
R5963 gnd.n3205 gnd.n1787 163.367
R5964 gnd.n3205 gnd.n1780 163.367
R5965 gnd.n3208 gnd.n1780 163.367
R5966 gnd.n3208 gnd.n1774 163.367
R5967 gnd.n3213 gnd.n1774 163.367
R5968 gnd.n3213 gnd.n1766 163.367
R5969 gnd.n1766 gnd.n1758 163.367
R5970 gnd.n3259 gnd.n1758 163.367
R5971 gnd.n3259 gnd.n1756 163.367
R5972 gnd.n3266 gnd.n1756 163.367
R5973 gnd.n3266 gnd.n1746 163.367
R5974 gnd.n1747 gnd.n1746 163.367
R5975 gnd.n1747 gnd.n1736 163.367
R5976 gnd.n1736 gnd.n1727 163.367
R5977 gnd.n3304 gnd.n1727 163.367
R5978 gnd.n3304 gnd.n1725 163.367
R5979 gnd.n3317 gnd.n1725 163.367
R5980 gnd.n3317 gnd.n1719 163.367
R5981 gnd.n3313 gnd.n1719 163.367
R5982 gnd.n3313 gnd.n3310 163.367
R5983 gnd.n3310 gnd.n3309 163.367
R5984 gnd.n3309 gnd.n1702 163.367
R5985 gnd.n3367 gnd.n1702 163.367
R5986 gnd.n3367 gnd.n1699 163.367
R5987 gnd.n3377 gnd.n1699 163.367
R5988 gnd.n3377 gnd.n1691 163.367
R5989 gnd.n3373 gnd.n1691 163.367
R5990 gnd.n3373 gnd.n1682 163.367
R5991 gnd.n1682 gnd.n1674 163.367
R5992 gnd.n3495 gnd.n1674 163.367
R5993 gnd.n1447 gnd.n1446 163.367
R5994 gnd.n3858 gnd.n1446 163.367
R5995 gnd.n3856 gnd.n3855 163.367
R5996 gnd.n3852 gnd.n3851 163.367
R5997 gnd.n3848 gnd.n3847 163.367
R5998 gnd.n3844 gnd.n3843 163.367
R5999 gnd.n3840 gnd.n3839 163.367
R6000 gnd.n3836 gnd.n3835 163.367
R6001 gnd.n3832 gnd.n3831 163.367
R6002 gnd.n3828 gnd.n3827 163.367
R6003 gnd.n3824 gnd.n3823 163.367
R6004 gnd.n3820 gnd.n3819 163.367
R6005 gnd.n3816 gnd.n3815 163.367
R6006 gnd.n3812 gnd.n3811 163.367
R6007 gnd.n3808 gnd.n3807 163.367
R6008 gnd.n3804 gnd.n3803 163.367
R6009 gnd.n3867 gnd.n1412 163.367
R6010 gnd.n2780 gnd.n2779 163.367
R6011 gnd.n2785 gnd.n2784 163.367
R6012 gnd.n2789 gnd.n2788 163.367
R6013 gnd.n2793 gnd.n2792 163.367
R6014 gnd.n2797 gnd.n2796 163.367
R6015 gnd.n2801 gnd.n2800 163.367
R6016 gnd.n2805 gnd.n2804 163.367
R6017 gnd.n2809 gnd.n2808 163.367
R6018 gnd.n2813 gnd.n2812 163.367
R6019 gnd.n2817 gnd.n2816 163.367
R6020 gnd.n2821 gnd.n2820 163.367
R6021 gnd.n2825 gnd.n2824 163.367
R6022 gnd.n2829 gnd.n2828 163.367
R6023 gnd.n2833 gnd.n2832 163.367
R6024 gnd.n2837 gnd.n2836 163.367
R6025 gnd.n3796 gnd.n1448 163.367
R6026 gnd.n3796 gnd.n1470 163.367
R6027 gnd.n2907 gnd.n1470 163.367
R6028 gnd.n2907 gnd.n1967 163.367
R6029 gnd.n2911 gnd.n1967 163.367
R6030 gnd.n2911 gnd.n1956 163.367
R6031 gnd.n2925 gnd.n1956 163.367
R6032 gnd.n2925 gnd.n1954 163.367
R6033 gnd.n2929 gnd.n1954 163.367
R6034 gnd.n2929 gnd.n1944 163.367
R6035 gnd.n2942 gnd.n1944 163.367
R6036 gnd.n2942 gnd.n1941 163.367
R6037 gnd.n2947 gnd.n1941 163.367
R6038 gnd.n2947 gnd.n1942 163.367
R6039 gnd.n1942 gnd.n1921 163.367
R6040 gnd.n2974 gnd.n1921 163.367
R6041 gnd.n2974 gnd.n1919 163.367
R6042 gnd.n2978 gnd.n1919 163.367
R6043 gnd.n2978 gnd.n1908 163.367
R6044 gnd.n2994 gnd.n1908 163.367
R6045 gnd.n2994 gnd.n1906 163.367
R6046 gnd.n2998 gnd.n1906 163.367
R6047 gnd.n2998 gnd.n1893 163.367
R6048 gnd.n3025 gnd.n1893 163.367
R6049 gnd.n3025 gnd.n1891 163.367
R6050 gnd.n3029 gnd.n1891 163.367
R6051 gnd.n3029 gnd.n1878 163.367
R6052 gnd.n3043 gnd.n1878 163.367
R6053 gnd.n3043 gnd.n1875 163.367
R6054 gnd.n3048 gnd.n1875 163.367
R6055 gnd.n3048 gnd.n1876 163.367
R6056 gnd.n1876 gnd.n1859 163.367
R6057 gnd.n3077 gnd.n1859 163.367
R6058 gnd.n3077 gnd.n1857 163.367
R6059 gnd.n3081 gnd.n1857 163.367
R6060 gnd.n3081 gnd.n1845 163.367
R6061 gnd.n3106 gnd.n1845 163.367
R6062 gnd.n3106 gnd.n1842 163.367
R6063 gnd.n3113 gnd.n1842 163.367
R6064 gnd.n3113 gnd.n1843 163.367
R6065 gnd.n3109 gnd.n1843 163.367
R6066 gnd.n3109 gnd.n1823 163.367
R6067 gnd.n3146 gnd.n1823 163.367
R6068 gnd.n3146 gnd.n1820 163.367
R6069 gnd.n3153 gnd.n1820 163.367
R6070 gnd.n3153 gnd.n1821 163.367
R6071 gnd.n3149 gnd.n1821 163.367
R6072 gnd.n3149 gnd.n1800 163.367
R6073 gnd.n3186 gnd.n1800 163.367
R6074 gnd.n3186 gnd.n1797 163.367
R6075 gnd.n3193 gnd.n1797 163.367
R6076 gnd.n3193 gnd.n1798 163.367
R6077 gnd.n3189 gnd.n1798 163.367
R6078 gnd.n3189 gnd.n1778 163.367
R6079 gnd.n3235 gnd.n1778 163.367
R6080 gnd.n3235 gnd.n1776 163.367
R6081 gnd.n3239 gnd.n1776 163.367
R6082 gnd.n3239 gnd.n1765 163.367
R6083 gnd.n3252 gnd.n1765 163.367
R6084 gnd.n3252 gnd.n1762 163.367
R6085 gnd.n3257 gnd.n1762 163.367
R6086 gnd.n3257 gnd.n1763 163.367
R6087 gnd.n1763 gnd.n1744 163.367
R6088 gnd.n3286 gnd.n1744 163.367
R6089 gnd.n3286 gnd.n1738 163.367
R6090 gnd.n3291 gnd.n1738 163.367
R6091 gnd.n3291 gnd.n1742 163.367
R6092 gnd.n1742 gnd.n1724 163.367
R6093 gnd.n3321 gnd.n1724 163.367
R6094 gnd.n3321 gnd.n1721 163.367
R6095 gnd.n3334 gnd.n1721 163.367
R6096 gnd.n3334 gnd.n1722 163.367
R6097 gnd.n3330 gnd.n1722 163.367
R6098 gnd.n3330 gnd.n3329 163.367
R6099 gnd.n3329 gnd.n3328 163.367
R6100 gnd.n3328 gnd.n1697 163.367
R6101 gnd.n3381 gnd.n1697 163.367
R6102 gnd.n3381 gnd.n1695 163.367
R6103 gnd.n3385 gnd.n1695 163.367
R6104 gnd.n3385 gnd.n1680 163.367
R6105 gnd.n3402 gnd.n1680 163.367
R6106 gnd.n3402 gnd.n1677 163.367
R6107 gnd.n3493 gnd.n1677 163.367
R6108 gnd.n3423 gnd.n3422 156.462
R6109 gnd.n5429 gnd.n5397 153.042
R6110 gnd.n5493 gnd.n5492 152.079
R6111 gnd.n5461 gnd.n5460 152.079
R6112 gnd.n5429 gnd.n5428 152.079
R6113 gnd.n1461 gnd.n1460 152
R6114 gnd.n1462 gnd.n1451 152
R6115 gnd.n1464 gnd.n1463 152
R6116 gnd.n1466 gnd.n1449 152
R6117 gnd.n1468 gnd.n1467 152
R6118 gnd.n3421 gnd.n3405 152
R6119 gnd.n3413 gnd.n3406 152
R6120 gnd.n3412 gnd.n3411 152
R6121 gnd.n3410 gnd.n3407 152
R6122 gnd.n3408 gnd.t112 150.546
R6123 gnd.t215 gnd.n5471 147.661
R6124 gnd.t326 gnd.n5439 147.661
R6125 gnd.t319 gnd.n5407 147.661
R6126 gnd.t225 gnd.n5376 147.661
R6127 gnd.t228 gnd.n5344 147.661
R6128 gnd.t39 gnd.n5312 147.661
R6129 gnd.t211 gnd.n5280 147.661
R6130 gnd.t243 gnd.n5249 147.661
R6131 gnd.n1670 gnd.n1653 143.351
R6132 gnd.n1428 gnd.n1411 143.351
R6133 gnd.n3866 gnd.n1411 143.351
R6134 gnd.n1458 gnd.t69 130.484
R6135 gnd.n1467 gnd.t80 126.766
R6136 gnd.n1465 gnd.t161 126.766
R6137 gnd.n1451 gnd.t174 126.766
R6138 gnd.n1459 gnd.t115 126.766
R6139 gnd.n3409 gnd.t87 126.766
R6140 gnd.n3411 gnd.t131 126.766
R6141 gnd.n3420 gnd.t102 126.766
R6142 gnd.n3422 gnd.t137 126.766
R6143 gnd.n5488 gnd.n5487 104.615
R6144 gnd.n5487 gnd.n5465 104.615
R6145 gnd.n5480 gnd.n5465 104.615
R6146 gnd.n5480 gnd.n5479 104.615
R6147 gnd.n5479 gnd.n5469 104.615
R6148 gnd.n5472 gnd.n5469 104.615
R6149 gnd.n5456 gnd.n5455 104.615
R6150 gnd.n5455 gnd.n5433 104.615
R6151 gnd.n5448 gnd.n5433 104.615
R6152 gnd.n5448 gnd.n5447 104.615
R6153 gnd.n5447 gnd.n5437 104.615
R6154 gnd.n5440 gnd.n5437 104.615
R6155 gnd.n5424 gnd.n5423 104.615
R6156 gnd.n5423 gnd.n5401 104.615
R6157 gnd.n5416 gnd.n5401 104.615
R6158 gnd.n5416 gnd.n5415 104.615
R6159 gnd.n5415 gnd.n5405 104.615
R6160 gnd.n5408 gnd.n5405 104.615
R6161 gnd.n5393 gnd.n5392 104.615
R6162 gnd.n5392 gnd.n5370 104.615
R6163 gnd.n5385 gnd.n5370 104.615
R6164 gnd.n5385 gnd.n5384 104.615
R6165 gnd.n5384 gnd.n5374 104.615
R6166 gnd.n5377 gnd.n5374 104.615
R6167 gnd.n5361 gnd.n5360 104.615
R6168 gnd.n5360 gnd.n5338 104.615
R6169 gnd.n5353 gnd.n5338 104.615
R6170 gnd.n5353 gnd.n5352 104.615
R6171 gnd.n5352 gnd.n5342 104.615
R6172 gnd.n5345 gnd.n5342 104.615
R6173 gnd.n5329 gnd.n5328 104.615
R6174 gnd.n5328 gnd.n5306 104.615
R6175 gnd.n5321 gnd.n5306 104.615
R6176 gnd.n5321 gnd.n5320 104.615
R6177 gnd.n5320 gnd.n5310 104.615
R6178 gnd.n5313 gnd.n5310 104.615
R6179 gnd.n5297 gnd.n5296 104.615
R6180 gnd.n5296 gnd.n5274 104.615
R6181 gnd.n5289 gnd.n5274 104.615
R6182 gnd.n5289 gnd.n5288 104.615
R6183 gnd.n5288 gnd.n5278 104.615
R6184 gnd.n5281 gnd.n5278 104.615
R6185 gnd.n5266 gnd.n5265 104.615
R6186 gnd.n5265 gnd.n5243 104.615
R6187 gnd.n5258 gnd.n5243 104.615
R6188 gnd.n5258 gnd.n5257 104.615
R6189 gnd.n5257 gnd.n5247 104.615
R6190 gnd.n5250 gnd.n5247 104.615
R6191 gnd.n4640 gnd.t127 100.632
R6192 gnd.n4198 gnd.t179 100.632
R6193 gnd.n7049 gnd.n6880 99.6594
R6194 gnd.n7047 gnd.n6879 99.6594
R6195 gnd.n7043 gnd.n6878 99.6594
R6196 gnd.n7039 gnd.n6877 99.6594
R6197 gnd.n7035 gnd.n6876 99.6594
R6198 gnd.n7031 gnd.n6875 99.6594
R6199 gnd.n7027 gnd.n6874 99.6594
R6200 gnd.n7023 gnd.n6873 99.6594
R6201 gnd.n7016 gnd.n6872 99.6594
R6202 gnd.n7012 gnd.n6871 99.6594
R6203 gnd.n7008 gnd.n6870 99.6594
R6204 gnd.n7004 gnd.n6869 99.6594
R6205 gnd.n7000 gnd.n6868 99.6594
R6206 gnd.n6996 gnd.n6867 99.6594
R6207 gnd.n6992 gnd.n6866 99.6594
R6208 gnd.n6988 gnd.n6865 99.6594
R6209 gnd.n6984 gnd.n6864 99.6594
R6210 gnd.n6980 gnd.n6863 99.6594
R6211 gnd.n6972 gnd.n6862 99.6594
R6212 gnd.n6970 gnd.n6861 99.6594
R6213 gnd.n6966 gnd.n6860 99.6594
R6214 gnd.n6962 gnd.n6859 99.6594
R6215 gnd.n6958 gnd.n6858 99.6594
R6216 gnd.n6954 gnd.n6857 99.6594
R6217 gnd.n6950 gnd.n6856 99.6594
R6218 gnd.n6946 gnd.n6855 99.6594
R6219 gnd.n6942 gnd.n6854 99.6594
R6220 gnd.n6938 gnd.n6853 99.6594
R6221 gnd.n7061 gnd.n7059 99.6594
R6222 gnd.n6548 gnd.n6547 99.6594
R6223 gnd.n324 gnd.n285 99.6594
R6224 gnd.n6540 gnd.n286 99.6594
R6225 gnd.n6536 gnd.n287 99.6594
R6226 gnd.n6532 gnd.n288 99.6594
R6227 gnd.n6528 gnd.n289 99.6594
R6228 gnd.n6524 gnd.n290 99.6594
R6229 gnd.n6520 gnd.n291 99.6594
R6230 gnd.n6516 gnd.n292 99.6594
R6231 gnd.n6511 gnd.n293 99.6594
R6232 gnd.n6507 gnd.n294 99.6594
R6233 gnd.n6503 gnd.n295 99.6594
R6234 gnd.n6499 gnd.n296 99.6594
R6235 gnd.n6494 gnd.n298 99.6594
R6236 gnd.n6490 gnd.n299 99.6594
R6237 gnd.n6486 gnd.n300 99.6594
R6238 gnd.n6482 gnd.n301 99.6594
R6239 gnd.n6478 gnd.n302 99.6594
R6240 gnd.n6474 gnd.n303 99.6594
R6241 gnd.n6470 gnd.n304 99.6594
R6242 gnd.n6466 gnd.n305 99.6594
R6243 gnd.n6462 gnd.n306 99.6594
R6244 gnd.n6458 gnd.n307 99.6594
R6245 gnd.n6454 gnd.n308 99.6594
R6246 gnd.n6450 gnd.n309 99.6594
R6247 gnd.n6446 gnd.n310 99.6594
R6248 gnd.n6442 gnd.n311 99.6594
R6249 gnd.n6438 gnd.n312 99.6594
R6250 gnd.n3918 gnd.n3917 99.6594
R6251 gnd.n3913 gnd.n1378 99.6594
R6252 gnd.n3909 gnd.n1377 99.6594
R6253 gnd.n3905 gnd.n1376 99.6594
R6254 gnd.n3901 gnd.n1375 99.6594
R6255 gnd.n3897 gnd.n1374 99.6594
R6256 gnd.n3893 gnd.n1373 99.6594
R6257 gnd.n3889 gnd.n1372 99.6594
R6258 gnd.n3884 gnd.n1371 99.6594
R6259 gnd.n3880 gnd.n1370 99.6594
R6260 gnd.n3876 gnd.n1369 99.6594
R6261 gnd.n3872 gnd.n1368 99.6594
R6262 gnd.n2170 gnd.n1366 99.6594
R6263 gnd.n2177 gnd.n1365 99.6594
R6264 gnd.n2181 gnd.n1364 99.6594
R6265 gnd.n2187 gnd.n1363 99.6594
R6266 gnd.n2191 gnd.n1362 99.6594
R6267 gnd.n2197 gnd.n1361 99.6594
R6268 gnd.n2201 gnd.n1360 99.6594
R6269 gnd.n2207 gnd.n1359 99.6594
R6270 gnd.n2211 gnd.n1358 99.6594
R6271 gnd.n2217 gnd.n1357 99.6594
R6272 gnd.n2221 gnd.n1356 99.6594
R6273 gnd.n2227 gnd.n1355 99.6594
R6274 gnd.n2231 gnd.n1354 99.6594
R6275 gnd.n2237 gnd.n1353 99.6594
R6276 gnd.n2241 gnd.n1352 99.6594
R6277 gnd.n2247 gnd.n1351 99.6594
R6278 gnd.n4172 gnd.n4171 99.6594
R6279 gnd.n4166 gnd.n1023 99.6594
R6280 gnd.n4163 gnd.n1024 99.6594
R6281 gnd.n4159 gnd.n1025 99.6594
R6282 gnd.n4155 gnd.n1026 99.6594
R6283 gnd.n4151 gnd.n1027 99.6594
R6284 gnd.n4147 gnd.n1028 99.6594
R6285 gnd.n4143 gnd.n1029 99.6594
R6286 gnd.n4139 gnd.n1030 99.6594
R6287 gnd.n4134 gnd.n1031 99.6594
R6288 gnd.n4130 gnd.n1032 99.6594
R6289 gnd.n4126 gnd.n1033 99.6594
R6290 gnd.n4122 gnd.n1034 99.6594
R6291 gnd.n4118 gnd.n1035 99.6594
R6292 gnd.n4114 gnd.n1036 99.6594
R6293 gnd.n4110 gnd.n1037 99.6594
R6294 gnd.n4106 gnd.n1038 99.6594
R6295 gnd.n4102 gnd.n1039 99.6594
R6296 gnd.n4098 gnd.n1040 99.6594
R6297 gnd.n4094 gnd.n1041 99.6594
R6298 gnd.n4090 gnd.n1042 99.6594
R6299 gnd.n4086 gnd.n1043 99.6594
R6300 gnd.n4082 gnd.n1044 99.6594
R6301 gnd.n4078 gnd.n1045 99.6594
R6302 gnd.n4074 gnd.n1046 99.6594
R6303 gnd.n4070 gnd.n1047 99.6594
R6304 gnd.n4066 gnd.n1048 99.6594
R6305 gnd.n4062 gnd.n1049 99.6594
R6306 gnd.n4058 gnd.n1050 99.6594
R6307 gnd.n5611 gnd.n4181 99.6594
R6308 gnd.n5609 gnd.n4180 99.6594
R6309 gnd.n5605 gnd.n4179 99.6594
R6310 gnd.n5601 gnd.n4178 99.6594
R6311 gnd.n5597 gnd.n4177 99.6594
R6312 gnd.n5593 gnd.n4176 99.6594
R6313 gnd.n5589 gnd.n4175 99.6594
R6314 gnd.n5521 gnd.n4174 99.6594
R6315 gnd.n4852 gnd.n4583 99.6594
R6316 gnd.n4609 gnd.n4590 99.6594
R6317 gnd.n4611 gnd.n4591 99.6594
R6318 gnd.n4619 gnd.n4592 99.6594
R6319 gnd.n4621 gnd.n4593 99.6594
R6320 gnd.n4629 gnd.n4594 99.6594
R6321 gnd.n4631 gnd.n4595 99.6594
R6322 gnd.n4639 gnd.n4596 99.6594
R6323 gnd.n6767 gnd.n6741 99.6594
R6324 gnd.n6771 gnd.n6742 99.6594
R6325 gnd.n6777 gnd.n6743 99.6594
R6326 gnd.n6781 gnd.n6744 99.6594
R6327 gnd.n6787 gnd.n6745 99.6594
R6328 gnd.n6791 gnd.n6746 99.6594
R6329 gnd.n6797 gnd.n6747 99.6594
R6330 gnd.n6800 gnd.n6748 99.6594
R6331 gnd.n6852 gnd.n6851 99.6594
R6332 gnd.n502 gnd.n313 99.6594
R6333 gnd.n400 gnd.n314 99.6594
R6334 gnd.n408 gnd.n315 99.6594
R6335 gnd.n410 gnd.n316 99.6594
R6336 gnd.n418 gnd.n317 99.6594
R6337 gnd.n426 gnd.n318 99.6594
R6338 gnd.n428 gnd.n319 99.6594
R6339 gnd.n436 gnd.n320 99.6594
R6340 gnd.n446 gnd.n321 99.6594
R6341 gnd.n5579 gnd.n1010 99.6594
R6342 gnd.n5575 gnd.n1011 99.6594
R6343 gnd.n5571 gnd.n1012 99.6594
R6344 gnd.n5567 gnd.n1013 99.6594
R6345 gnd.n5563 gnd.n1014 99.6594
R6346 gnd.n5559 gnd.n1015 99.6594
R6347 gnd.n5555 gnd.n1016 99.6594
R6348 gnd.n5551 gnd.n1017 99.6594
R6349 gnd.n5547 gnd.n1018 99.6594
R6350 gnd.n5543 gnd.n1019 99.6594
R6351 gnd.n5539 gnd.n1020 99.6594
R6352 gnd.n5535 gnd.n1021 99.6594
R6353 gnd.n5531 gnd.n1022 99.6594
R6354 gnd.n4767 gnd.n4766 99.6594
R6355 gnd.n4761 gnd.n4678 99.6594
R6356 gnd.n4758 gnd.n4679 99.6594
R6357 gnd.n4754 gnd.n4680 99.6594
R6358 gnd.n4750 gnd.n4681 99.6594
R6359 gnd.n4746 gnd.n4682 99.6594
R6360 gnd.n4742 gnd.n4683 99.6594
R6361 gnd.n4738 gnd.n4684 99.6594
R6362 gnd.n4734 gnd.n4685 99.6594
R6363 gnd.n4730 gnd.n4686 99.6594
R6364 gnd.n4726 gnd.n4687 99.6594
R6365 gnd.n4722 gnd.n4688 99.6594
R6366 gnd.n4769 gnd.n4677 99.6594
R6367 gnd.n2099 gnd.n1341 99.6594
R6368 gnd.n2107 gnd.n1342 99.6594
R6369 gnd.n2115 gnd.n1343 99.6594
R6370 gnd.n2117 gnd.n1344 99.6594
R6371 gnd.n2125 gnd.n1345 99.6594
R6372 gnd.n2133 gnd.n1346 99.6594
R6373 gnd.n2135 gnd.n1347 99.6594
R6374 gnd.n2145 gnd.n1348 99.6594
R6375 gnd.n2569 gnd.n1349 99.6594
R6376 gnd.n1133 gnd.n1051 99.6594
R6377 gnd.n2326 gnd.n1052 99.6594
R6378 gnd.n2332 gnd.n1053 99.6594
R6379 gnd.n2336 gnd.n1054 99.6594
R6380 gnd.n2342 gnd.n1055 99.6594
R6381 gnd.n2346 gnd.n1056 99.6594
R6382 gnd.n2352 gnd.n1057 99.6594
R6383 gnd.n2356 gnd.n1058 99.6594
R6384 gnd.n2315 gnd.n1059 99.6594
R6385 gnd.n2325 gnd.n1051 99.6594
R6386 gnd.n2331 gnd.n1052 99.6594
R6387 gnd.n2335 gnd.n1053 99.6594
R6388 gnd.n2341 gnd.n1054 99.6594
R6389 gnd.n2345 gnd.n1055 99.6594
R6390 gnd.n2351 gnd.n1056 99.6594
R6391 gnd.n2355 gnd.n1057 99.6594
R6392 gnd.n2314 gnd.n1058 99.6594
R6393 gnd.n2310 gnd.n1059 99.6594
R6394 gnd.n2149 gnd.n1349 99.6594
R6395 gnd.n2136 gnd.n1348 99.6594
R6396 gnd.n2134 gnd.n1347 99.6594
R6397 gnd.n2126 gnd.n1346 99.6594
R6398 gnd.n2118 gnd.n1345 99.6594
R6399 gnd.n2116 gnd.n1344 99.6594
R6400 gnd.n2108 gnd.n1343 99.6594
R6401 gnd.n2100 gnd.n1342 99.6594
R6402 gnd.n2098 gnd.n1341 99.6594
R6403 gnd.n4767 gnd.n4690 99.6594
R6404 gnd.n4759 gnd.n4678 99.6594
R6405 gnd.n4755 gnd.n4679 99.6594
R6406 gnd.n4751 gnd.n4680 99.6594
R6407 gnd.n4747 gnd.n4681 99.6594
R6408 gnd.n4743 gnd.n4682 99.6594
R6409 gnd.n4739 gnd.n4683 99.6594
R6410 gnd.n4735 gnd.n4684 99.6594
R6411 gnd.n4731 gnd.n4685 99.6594
R6412 gnd.n4727 gnd.n4686 99.6594
R6413 gnd.n4723 gnd.n4687 99.6594
R6414 gnd.n4719 gnd.n4688 99.6594
R6415 gnd.n4770 gnd.n4769 99.6594
R6416 gnd.n5534 gnd.n1022 99.6594
R6417 gnd.n5538 gnd.n1021 99.6594
R6418 gnd.n5542 gnd.n1020 99.6594
R6419 gnd.n5546 gnd.n1019 99.6594
R6420 gnd.n5550 gnd.n1018 99.6594
R6421 gnd.n5554 gnd.n1017 99.6594
R6422 gnd.n5558 gnd.n1016 99.6594
R6423 gnd.n5562 gnd.n1015 99.6594
R6424 gnd.n5566 gnd.n1014 99.6594
R6425 gnd.n5570 gnd.n1013 99.6594
R6426 gnd.n5574 gnd.n1012 99.6594
R6427 gnd.n5578 gnd.n1011 99.6594
R6428 gnd.n4202 gnd.n1010 99.6594
R6429 gnd.n399 gnd.n313 99.6594
R6430 gnd.n407 gnd.n314 99.6594
R6431 gnd.n409 gnd.n315 99.6594
R6432 gnd.n417 gnd.n316 99.6594
R6433 gnd.n425 gnd.n317 99.6594
R6434 gnd.n427 gnd.n318 99.6594
R6435 gnd.n435 gnd.n319 99.6594
R6436 gnd.n445 gnd.n320 99.6594
R6437 gnd.n6382 gnd.n321 99.6594
R6438 gnd.n6852 gnd.n6749 99.6594
R6439 gnd.n6798 gnd.n6748 99.6594
R6440 gnd.n6790 gnd.n6747 99.6594
R6441 gnd.n6788 gnd.n6746 99.6594
R6442 gnd.n6780 gnd.n6745 99.6594
R6443 gnd.n6778 gnd.n6744 99.6594
R6444 gnd.n6770 gnd.n6743 99.6594
R6445 gnd.n6768 gnd.n6742 99.6594
R6446 gnd.n6762 gnd.n6741 99.6594
R6447 gnd.n4853 gnd.n4852 99.6594
R6448 gnd.n4612 gnd.n4590 99.6594
R6449 gnd.n4618 gnd.n4591 99.6594
R6450 gnd.n4622 gnd.n4592 99.6594
R6451 gnd.n4628 gnd.n4593 99.6594
R6452 gnd.n4632 gnd.n4594 99.6594
R6453 gnd.n4638 gnd.n4595 99.6594
R6454 gnd.n4596 gnd.n4580 99.6594
R6455 gnd.n5588 gnd.n4174 99.6594
R6456 gnd.n5592 gnd.n4175 99.6594
R6457 gnd.n5596 gnd.n4176 99.6594
R6458 gnd.n5600 gnd.n4177 99.6594
R6459 gnd.n5604 gnd.n4178 99.6594
R6460 gnd.n5608 gnd.n4179 99.6594
R6461 gnd.n5612 gnd.n4180 99.6594
R6462 gnd.n4183 gnd.n4181 99.6594
R6463 gnd.n4172 gnd.n1063 99.6594
R6464 gnd.n4164 gnd.n1023 99.6594
R6465 gnd.n4160 gnd.n1024 99.6594
R6466 gnd.n4156 gnd.n1025 99.6594
R6467 gnd.n4152 gnd.n1026 99.6594
R6468 gnd.n4148 gnd.n1027 99.6594
R6469 gnd.n4144 gnd.n1028 99.6594
R6470 gnd.n4140 gnd.n1029 99.6594
R6471 gnd.n4135 gnd.n1030 99.6594
R6472 gnd.n4131 gnd.n1031 99.6594
R6473 gnd.n4127 gnd.n1032 99.6594
R6474 gnd.n4123 gnd.n1033 99.6594
R6475 gnd.n4119 gnd.n1034 99.6594
R6476 gnd.n4115 gnd.n1035 99.6594
R6477 gnd.n4111 gnd.n1036 99.6594
R6478 gnd.n4107 gnd.n1037 99.6594
R6479 gnd.n4103 gnd.n1038 99.6594
R6480 gnd.n4099 gnd.n1039 99.6594
R6481 gnd.n4095 gnd.n1040 99.6594
R6482 gnd.n4091 gnd.n1041 99.6594
R6483 gnd.n4087 gnd.n1042 99.6594
R6484 gnd.n4083 gnd.n1043 99.6594
R6485 gnd.n4079 gnd.n1044 99.6594
R6486 gnd.n4075 gnd.n1045 99.6594
R6487 gnd.n4071 gnd.n1046 99.6594
R6488 gnd.n4067 gnd.n1047 99.6594
R6489 gnd.n4063 gnd.n1048 99.6594
R6490 gnd.n4059 gnd.n1049 99.6594
R6491 gnd.n1135 gnd.n1050 99.6594
R6492 gnd.n2240 gnd.n1351 99.6594
R6493 gnd.n2238 gnd.n1352 99.6594
R6494 gnd.n2230 gnd.n1353 99.6594
R6495 gnd.n2228 gnd.n1354 99.6594
R6496 gnd.n2220 gnd.n1355 99.6594
R6497 gnd.n2218 gnd.n1356 99.6594
R6498 gnd.n2210 gnd.n1357 99.6594
R6499 gnd.n2208 gnd.n1358 99.6594
R6500 gnd.n2200 gnd.n1359 99.6594
R6501 gnd.n2198 gnd.n1360 99.6594
R6502 gnd.n2190 gnd.n1361 99.6594
R6503 gnd.n2188 gnd.n1362 99.6594
R6504 gnd.n2180 gnd.n1363 99.6594
R6505 gnd.n2178 gnd.n1364 99.6594
R6506 gnd.n2171 gnd.n1365 99.6594
R6507 gnd.n3871 gnd.n1367 99.6594
R6508 gnd.n3875 gnd.n1368 99.6594
R6509 gnd.n3879 gnd.n1369 99.6594
R6510 gnd.n3883 gnd.n1370 99.6594
R6511 gnd.n3888 gnd.n1371 99.6594
R6512 gnd.n3892 gnd.n1372 99.6594
R6513 gnd.n3896 gnd.n1373 99.6594
R6514 gnd.n3900 gnd.n1374 99.6594
R6515 gnd.n3904 gnd.n1375 99.6594
R6516 gnd.n3908 gnd.n1376 99.6594
R6517 gnd.n3912 gnd.n1377 99.6594
R6518 gnd.n1379 gnd.n1378 99.6594
R6519 gnd.n3918 gnd.n1338 99.6594
R6520 gnd.n6547 gnd.n283 99.6594
R6521 gnd.n6541 gnd.n285 99.6594
R6522 gnd.n6537 gnd.n286 99.6594
R6523 gnd.n6533 gnd.n287 99.6594
R6524 gnd.n6529 gnd.n288 99.6594
R6525 gnd.n6525 gnd.n289 99.6594
R6526 gnd.n6521 gnd.n290 99.6594
R6527 gnd.n6517 gnd.n291 99.6594
R6528 gnd.n6512 gnd.n292 99.6594
R6529 gnd.n6508 gnd.n293 99.6594
R6530 gnd.n6504 gnd.n294 99.6594
R6531 gnd.n6500 gnd.n295 99.6594
R6532 gnd.n6495 gnd.n297 99.6594
R6533 gnd.n6491 gnd.n298 99.6594
R6534 gnd.n6487 gnd.n299 99.6594
R6535 gnd.n6483 gnd.n300 99.6594
R6536 gnd.n6479 gnd.n301 99.6594
R6537 gnd.n6475 gnd.n302 99.6594
R6538 gnd.n6471 gnd.n303 99.6594
R6539 gnd.n6467 gnd.n304 99.6594
R6540 gnd.n6463 gnd.n305 99.6594
R6541 gnd.n6459 gnd.n306 99.6594
R6542 gnd.n6455 gnd.n307 99.6594
R6543 gnd.n6451 gnd.n308 99.6594
R6544 gnd.n6447 gnd.n309 99.6594
R6545 gnd.n6443 gnd.n310 99.6594
R6546 gnd.n6439 gnd.n311 99.6594
R6547 gnd.n500 gnd.n312 99.6594
R6548 gnd.n7059 gnd.n6739 99.6594
R6549 gnd.n6941 gnd.n6853 99.6594
R6550 gnd.n6945 gnd.n6854 99.6594
R6551 gnd.n6949 gnd.n6855 99.6594
R6552 gnd.n6953 gnd.n6856 99.6594
R6553 gnd.n6957 gnd.n6857 99.6594
R6554 gnd.n6961 gnd.n6858 99.6594
R6555 gnd.n6965 gnd.n6859 99.6594
R6556 gnd.n6969 gnd.n6860 99.6594
R6557 gnd.n6973 gnd.n6861 99.6594
R6558 gnd.n6979 gnd.n6862 99.6594
R6559 gnd.n6983 gnd.n6863 99.6594
R6560 gnd.n6987 gnd.n6864 99.6594
R6561 gnd.n6991 gnd.n6865 99.6594
R6562 gnd.n6995 gnd.n6866 99.6594
R6563 gnd.n6999 gnd.n6867 99.6594
R6564 gnd.n7003 gnd.n6868 99.6594
R6565 gnd.n7007 gnd.n6869 99.6594
R6566 gnd.n7011 gnd.n6870 99.6594
R6567 gnd.n7015 gnd.n6871 99.6594
R6568 gnd.n7022 gnd.n6872 99.6594
R6569 gnd.n7026 gnd.n6873 99.6594
R6570 gnd.n7030 gnd.n6874 99.6594
R6571 gnd.n7034 gnd.n6875 99.6594
R6572 gnd.n7038 gnd.n6876 99.6594
R6573 gnd.n7042 gnd.n6877 99.6594
R6574 gnd.n7046 gnd.n6878 99.6594
R6575 gnd.n7050 gnd.n6879 99.6594
R6576 gnd.n6881 gnd.n6880 99.6594
R6577 gnd.n2556 gnd.n2079 99.6594
R6578 gnd.n2258 gnd.n2257 99.6594
R6579 gnd.n2259 gnd.n2088 99.6594
R6580 gnd.n2261 gnd.n2260 99.6594
R6581 gnd.n2263 gnd.n2094 99.6594
R6582 gnd.n2264 gnd.n2103 99.6594
R6583 gnd.n2266 gnd.n2265 99.6594
R6584 gnd.n2268 gnd.n2112 99.6594
R6585 gnd.n2269 gnd.n2121 99.6594
R6586 gnd.n2271 gnd.n2270 99.6594
R6587 gnd.n2273 gnd.n2130 99.6594
R6588 gnd.n2274 gnd.n2139 99.6594
R6589 gnd.n2277 gnd.n2275 99.6594
R6590 gnd.n2545 gnd.n2544 99.6594
R6591 gnd.n2556 gnd.n2083 99.6594
R6592 gnd.n2258 gnd.n2087 99.6594
R6593 gnd.n2259 gnd.n2089 99.6594
R6594 gnd.n2261 gnd.n2093 99.6594
R6595 gnd.n2263 gnd.n2262 99.6594
R6596 gnd.n2264 gnd.n2104 99.6594
R6597 gnd.n2266 gnd.n2111 99.6594
R6598 gnd.n2268 gnd.n2267 99.6594
R6599 gnd.n2269 gnd.n2122 99.6594
R6600 gnd.n2271 gnd.n2129 99.6594
R6601 gnd.n2273 gnd.n2272 99.6594
R6602 gnd.n2274 gnd.n2140 99.6594
R6603 gnd.n2276 gnd.n2275 99.6594
R6604 gnd.n2545 gnd.n2076 99.6594
R6605 gnd.n471 gnd.n464 99.6594
R6606 gnd.n473 gnd.n472 99.6594
R6607 gnd.n6358 gnd.n469 99.6594
R6608 gnd.n6356 gnd.n392 99.6594
R6609 gnd.n474 gnd.n394 99.6594
R6610 gnd.n476 gnd.n403 99.6594
R6611 gnd.n478 gnd.n477 99.6594
R6612 gnd.n479 gnd.n414 99.6594
R6613 gnd.n481 gnd.n421 99.6594
R6614 gnd.n483 gnd.n482 99.6594
R6615 gnd.n484 gnd.n432 99.6594
R6616 gnd.n486 gnd.n439 99.6594
R6617 gnd.n488 gnd.n487 99.6594
R6618 gnd.n489 gnd.n451 99.6594
R6619 gnd.n486 gnd.n485 99.6594
R6620 gnd.n484 gnd.n431 99.6594
R6621 gnd.n483 gnd.n422 99.6594
R6622 gnd.n481 gnd.n480 99.6594
R6623 gnd.n479 gnd.n413 99.6594
R6624 gnd.n478 gnd.n404 99.6594
R6625 gnd.n476 gnd.n475 99.6594
R6626 gnd.n474 gnd.n393 99.6594
R6627 gnd.n6357 gnd.n6356 99.6594
R6628 gnd.n469 gnd.n468 99.6594
R6629 gnd.n473 gnd.n465 99.6594
R6630 gnd.n471 gnd.n460 99.6594
R6631 gnd.n489 gnd.n456 99.6594
R6632 gnd.n488 gnd.n450 99.6594
R6633 gnd.n2141 gnd.t108 98.63
R6634 gnd.n6383 gnd.t68 98.63
R6635 gnd.n6736 gnd.t119 98.63
R6636 gnd.n6919 gnd.t129 98.63
R6637 gnd.n7018 gnd.t141 98.63
R6638 gnd.n341 gnd.t160 98.63
R6639 gnd.n364 gnd.t166 98.63
R6640 gnd.n386 gnd.t123 98.63
R6641 gnd.n6751 gnd.t63 98.63
R6642 gnd.n2146 gnd.t100 98.63
R6643 gnd.n2311 gnd.t97 98.63
R6644 gnd.n1083 gnd.t111 98.63
R6645 gnd.n1105 gnd.t145 98.63
R6646 gnd.n1127 gnd.t151 98.63
R6647 gnd.n1396 gnd.t135 98.63
R6648 gnd.n2152 gnd.t153 98.63
R6649 gnd.n2164 gnd.t172 98.63
R6650 gnd.n441 gnd.t74 98.63
R6651 gnd.n2776 gnd.t157 92.8196
R6652 gnd.n1671 gnd.t92 92.8196
R6653 gnd.n3800 gnd.t86 92.8118
R6654 gnd.n3424 gnd.t147 92.8118
R6655 gnd.n6118 gnd.n643 87.1465
R6656 gnd.n6119 gnd.n6118 87.1465
R6657 gnd.n6120 gnd.n6119 87.1465
R6658 gnd.n6120 gnd.n637 87.1465
R6659 gnd.n6128 gnd.n637 87.1465
R6660 gnd.n6129 gnd.n6128 87.1465
R6661 gnd.n6130 gnd.n6129 87.1465
R6662 gnd.n6130 gnd.n631 87.1465
R6663 gnd.n6138 gnd.n631 87.1465
R6664 gnd.n6139 gnd.n6138 87.1465
R6665 gnd.n6140 gnd.n6139 87.1465
R6666 gnd.n6140 gnd.n625 87.1465
R6667 gnd.n6148 gnd.n625 87.1465
R6668 gnd.n6149 gnd.n6148 87.1465
R6669 gnd.n6150 gnd.n6149 87.1465
R6670 gnd.n6150 gnd.n619 87.1465
R6671 gnd.n6158 gnd.n619 87.1465
R6672 gnd.n6159 gnd.n6158 87.1465
R6673 gnd.n6160 gnd.n6159 87.1465
R6674 gnd.n6160 gnd.n613 87.1465
R6675 gnd.n6168 gnd.n613 87.1465
R6676 gnd.n6169 gnd.n6168 87.1465
R6677 gnd.n6170 gnd.n6169 87.1465
R6678 gnd.n6170 gnd.n607 87.1465
R6679 gnd.n6178 gnd.n607 87.1465
R6680 gnd.n6179 gnd.n6178 87.1465
R6681 gnd.n6180 gnd.n6179 87.1465
R6682 gnd.n6180 gnd.n601 87.1465
R6683 gnd.n6188 gnd.n601 87.1465
R6684 gnd.n6189 gnd.n6188 87.1465
R6685 gnd.n6190 gnd.n6189 87.1465
R6686 gnd.n6190 gnd.n595 87.1465
R6687 gnd.n6198 gnd.n595 87.1465
R6688 gnd.n6199 gnd.n6198 87.1465
R6689 gnd.n6200 gnd.n6199 87.1465
R6690 gnd.n6200 gnd.n589 87.1465
R6691 gnd.n6208 gnd.n589 87.1465
R6692 gnd.n6209 gnd.n6208 87.1465
R6693 gnd.n6210 gnd.n6209 87.1465
R6694 gnd.n6210 gnd.n583 87.1465
R6695 gnd.n6218 gnd.n583 87.1465
R6696 gnd.n6219 gnd.n6218 87.1465
R6697 gnd.n6220 gnd.n6219 87.1465
R6698 gnd.n6220 gnd.n577 87.1465
R6699 gnd.n6228 gnd.n577 87.1465
R6700 gnd.n6229 gnd.n6228 87.1465
R6701 gnd.n6230 gnd.n6229 87.1465
R6702 gnd.n6230 gnd.n571 87.1465
R6703 gnd.n6238 gnd.n571 87.1465
R6704 gnd.n6239 gnd.n6238 87.1465
R6705 gnd.n6240 gnd.n6239 87.1465
R6706 gnd.n6240 gnd.n565 87.1465
R6707 gnd.n6248 gnd.n565 87.1465
R6708 gnd.n6249 gnd.n6248 87.1465
R6709 gnd.n6250 gnd.n6249 87.1465
R6710 gnd.n6250 gnd.n559 87.1465
R6711 gnd.n6258 gnd.n559 87.1465
R6712 gnd.n6259 gnd.n6258 87.1465
R6713 gnd.n6260 gnd.n6259 87.1465
R6714 gnd.n6260 gnd.n553 87.1465
R6715 gnd.n6268 gnd.n553 87.1465
R6716 gnd.n6269 gnd.n6268 87.1465
R6717 gnd.n6270 gnd.n6269 87.1465
R6718 gnd.n6270 gnd.n547 87.1465
R6719 gnd.n6278 gnd.n547 87.1465
R6720 gnd.n6279 gnd.n6278 87.1465
R6721 gnd.n6280 gnd.n6279 87.1465
R6722 gnd.n6280 gnd.n541 87.1465
R6723 gnd.n6288 gnd.n541 87.1465
R6724 gnd.n6289 gnd.n6288 87.1465
R6725 gnd.n6290 gnd.n6289 87.1465
R6726 gnd.n6290 gnd.n535 87.1465
R6727 gnd.n6298 gnd.n535 87.1465
R6728 gnd.n6299 gnd.n6298 87.1465
R6729 gnd.n6300 gnd.n6299 87.1465
R6730 gnd.n6300 gnd.n529 87.1465
R6731 gnd.n6308 gnd.n529 87.1465
R6732 gnd.n6309 gnd.n6308 87.1465
R6733 gnd.n6310 gnd.n6309 87.1465
R6734 gnd.n6310 gnd.n523 87.1465
R6735 gnd.n6320 gnd.n523 87.1465
R6736 gnd.n6321 gnd.n6320 87.1465
R6737 gnd.n6323 gnd.n6321 87.1465
R6738 gnd.n1458 gnd.n1457 81.8399
R6739 gnd.n4641 gnd.t126 74.8376
R6740 gnd.n4199 gnd.t180 74.8376
R6741 gnd.n2777 gnd.t156 72.8438
R6742 gnd.n1672 gnd.t93 72.8438
R6743 gnd.n1459 gnd.n1452 72.8411
R6744 gnd.n1465 gnd.n1450 72.8411
R6745 gnd.n3420 gnd.n3419 72.8411
R6746 gnd.n2142 gnd.t107 72.836
R6747 gnd.n3801 gnd.t85 72.836
R6748 gnd.n3425 gnd.t148 72.836
R6749 gnd.n6384 gnd.t67 72.836
R6750 gnd.n6737 gnd.t120 72.836
R6751 gnd.n6920 gnd.t130 72.836
R6752 gnd.n7019 gnd.t142 72.836
R6753 gnd.n342 gnd.t159 72.836
R6754 gnd.n365 gnd.t165 72.836
R6755 gnd.n387 gnd.t122 72.836
R6756 gnd.n6752 gnd.t64 72.836
R6757 gnd.n2147 gnd.t101 72.836
R6758 gnd.n2312 gnd.t96 72.836
R6759 gnd.n1084 gnd.t110 72.836
R6760 gnd.n1106 gnd.t144 72.836
R6761 gnd.n1128 gnd.t150 72.836
R6762 gnd.n1397 gnd.t136 72.836
R6763 gnd.n2153 gnd.t154 72.836
R6764 gnd.n2165 gnd.t173 72.836
R6765 gnd.n442 gnd.t75 72.836
R6766 gnd.n3488 gnd.n1637 71.676
R6767 gnd.n3484 gnd.n1638 71.676
R6768 gnd.n3480 gnd.n1639 71.676
R6769 gnd.n3476 gnd.n1640 71.676
R6770 gnd.n3472 gnd.n1641 71.676
R6771 gnd.n3468 gnd.n1642 71.676
R6772 gnd.n3464 gnd.n1643 71.676
R6773 gnd.n3460 gnd.n1644 71.676
R6774 gnd.n3456 gnd.n1645 71.676
R6775 gnd.n3452 gnd.n1646 71.676
R6776 gnd.n3448 gnd.n1647 71.676
R6777 gnd.n3444 gnd.n1648 71.676
R6778 gnd.n3440 gnd.n1649 71.676
R6779 gnd.n3436 gnd.n1650 71.676
R6780 gnd.n3431 gnd.n1651 71.676
R6781 gnd.n3427 gnd.n1652 71.676
R6782 gnd.n3561 gnd.n1670 71.676
R6783 gnd.n3557 gnd.n1669 71.676
R6784 gnd.n3552 gnd.n1668 71.676
R6785 gnd.n3548 gnd.n1667 71.676
R6786 gnd.n3544 gnd.n1666 71.676
R6787 gnd.n3540 gnd.n1665 71.676
R6788 gnd.n3536 gnd.n1664 71.676
R6789 gnd.n3532 gnd.n1663 71.676
R6790 gnd.n3528 gnd.n1662 71.676
R6791 gnd.n3524 gnd.n1661 71.676
R6792 gnd.n3520 gnd.n1660 71.676
R6793 gnd.n3516 gnd.n1659 71.676
R6794 gnd.n3512 gnd.n1658 71.676
R6795 gnd.n3508 gnd.n1657 71.676
R6796 gnd.n3504 gnd.n1656 71.676
R6797 gnd.n3500 gnd.n1655 71.676
R6798 gnd.n3496 gnd.n1654 71.676
R6799 gnd.n3864 gnd.n3863 71.676
R6800 gnd.n3858 gnd.n1414 71.676
R6801 gnd.n3855 gnd.n1415 71.676
R6802 gnd.n3851 gnd.n1416 71.676
R6803 gnd.n3847 gnd.n1417 71.676
R6804 gnd.n3843 gnd.n1418 71.676
R6805 gnd.n3839 gnd.n1419 71.676
R6806 gnd.n3835 gnd.n1420 71.676
R6807 gnd.n3831 gnd.n1421 71.676
R6808 gnd.n3827 gnd.n1422 71.676
R6809 gnd.n3823 gnd.n1423 71.676
R6810 gnd.n3819 gnd.n1424 71.676
R6811 gnd.n3815 gnd.n1425 71.676
R6812 gnd.n3811 gnd.n1426 71.676
R6813 gnd.n3807 gnd.n1427 71.676
R6814 gnd.n3803 gnd.n1428 71.676
R6815 gnd.n1429 gnd.n1412 71.676
R6816 gnd.n2780 gnd.n1430 71.676
R6817 gnd.n2785 gnd.n1431 71.676
R6818 gnd.n2789 gnd.n1432 71.676
R6819 gnd.n2793 gnd.n1433 71.676
R6820 gnd.n2797 gnd.n1434 71.676
R6821 gnd.n2801 gnd.n1435 71.676
R6822 gnd.n2805 gnd.n1436 71.676
R6823 gnd.n2809 gnd.n1437 71.676
R6824 gnd.n2813 gnd.n1438 71.676
R6825 gnd.n2817 gnd.n1439 71.676
R6826 gnd.n2821 gnd.n1440 71.676
R6827 gnd.n2825 gnd.n1441 71.676
R6828 gnd.n2829 gnd.n1442 71.676
R6829 gnd.n2833 gnd.n1443 71.676
R6830 gnd.n2837 gnd.n1444 71.676
R6831 gnd.n3864 gnd.n1447 71.676
R6832 gnd.n3856 gnd.n1414 71.676
R6833 gnd.n3852 gnd.n1415 71.676
R6834 gnd.n3848 gnd.n1416 71.676
R6835 gnd.n3844 gnd.n1417 71.676
R6836 gnd.n3840 gnd.n1418 71.676
R6837 gnd.n3836 gnd.n1419 71.676
R6838 gnd.n3832 gnd.n1420 71.676
R6839 gnd.n3828 gnd.n1421 71.676
R6840 gnd.n3824 gnd.n1422 71.676
R6841 gnd.n3820 gnd.n1423 71.676
R6842 gnd.n3816 gnd.n1424 71.676
R6843 gnd.n3812 gnd.n1425 71.676
R6844 gnd.n3808 gnd.n1426 71.676
R6845 gnd.n3804 gnd.n1427 71.676
R6846 gnd.n3867 gnd.n3866 71.676
R6847 gnd.n2779 gnd.n1429 71.676
R6848 gnd.n2784 gnd.n1430 71.676
R6849 gnd.n2788 gnd.n1431 71.676
R6850 gnd.n2792 gnd.n1432 71.676
R6851 gnd.n2796 gnd.n1433 71.676
R6852 gnd.n2800 gnd.n1434 71.676
R6853 gnd.n2804 gnd.n1435 71.676
R6854 gnd.n2808 gnd.n1436 71.676
R6855 gnd.n2812 gnd.n1437 71.676
R6856 gnd.n2816 gnd.n1438 71.676
R6857 gnd.n2820 gnd.n1439 71.676
R6858 gnd.n2824 gnd.n1440 71.676
R6859 gnd.n2828 gnd.n1441 71.676
R6860 gnd.n2832 gnd.n1442 71.676
R6861 gnd.n2836 gnd.n1443 71.676
R6862 gnd.n2775 gnd.n1444 71.676
R6863 gnd.n3499 gnd.n1654 71.676
R6864 gnd.n3503 gnd.n1655 71.676
R6865 gnd.n3507 gnd.n1656 71.676
R6866 gnd.n3511 gnd.n1657 71.676
R6867 gnd.n3515 gnd.n1658 71.676
R6868 gnd.n3519 gnd.n1659 71.676
R6869 gnd.n3523 gnd.n1660 71.676
R6870 gnd.n3527 gnd.n1661 71.676
R6871 gnd.n3531 gnd.n1662 71.676
R6872 gnd.n3535 gnd.n1663 71.676
R6873 gnd.n3539 gnd.n1664 71.676
R6874 gnd.n3543 gnd.n1665 71.676
R6875 gnd.n3547 gnd.n1666 71.676
R6876 gnd.n3551 gnd.n1667 71.676
R6877 gnd.n3556 gnd.n1668 71.676
R6878 gnd.n3560 gnd.n1669 71.676
R6879 gnd.n3426 gnd.n1653 71.676
R6880 gnd.n3430 gnd.n1652 71.676
R6881 gnd.n3435 gnd.n1651 71.676
R6882 gnd.n3439 gnd.n1650 71.676
R6883 gnd.n3443 gnd.n1649 71.676
R6884 gnd.n3447 gnd.n1648 71.676
R6885 gnd.n3451 gnd.n1647 71.676
R6886 gnd.n3455 gnd.n1646 71.676
R6887 gnd.n3459 gnd.n1645 71.676
R6888 gnd.n3463 gnd.n1644 71.676
R6889 gnd.n3467 gnd.n1643 71.676
R6890 gnd.n3471 gnd.n1642 71.676
R6891 gnd.n3475 gnd.n1641 71.676
R6892 gnd.n3479 gnd.n1640 71.676
R6893 gnd.n3483 gnd.n1639 71.676
R6894 gnd.n3487 gnd.n1638 71.676
R6895 gnd.n1678 gnd.n1637 71.676
R6896 gnd.n10 gnd.t20 69.1507
R6897 gnd.n18 gnd.t281 68.4792
R6898 gnd.n17 gnd.t247 68.4792
R6899 gnd.n16 gnd.t46 68.4792
R6900 gnd.n15 gnd.t237 68.4792
R6901 gnd.n14 gnd.t219 68.4792
R6902 gnd.n13 gnd.t315 68.4792
R6903 gnd.n12 gnd.t279 68.4792
R6904 gnd.n11 gnd.t324 68.4792
R6905 gnd.n10 gnd.t30 68.4792
R6906 gnd.n4768 gnd.n4672 64.369
R6907 gnd.n4173 gnd.n1061 63.0944
R6908 gnd.n7058 gnd.n164 63.0944
R6909 gnd.n2782 gnd.n2777 59.5399
R6910 gnd.n3554 gnd.n1672 59.5399
R6911 gnd.n3802 gnd.n3801 59.5399
R6912 gnd.n3433 gnd.n3425 59.5399
R6913 gnd.n3799 gnd.n1468 59.1804
R6914 gnd.n4427 gnd.t42 56.407
R6915 gnd.n4392 gnd.t316 56.407
R6916 gnd.n4403 gnd.t5 56.407
R6917 gnd.n4415 gnd.t60 56.407
R6918 gnd.n56 gnd.t25 56.407
R6919 gnd.n21 gnd.t233 56.407
R6920 gnd.n32 gnd.t331 56.407
R6921 gnd.n44 gnd.t221 56.407
R6922 gnd.n4436 gnd.t253 55.8337
R6923 gnd.n4401 gnd.t53 55.8337
R6924 gnd.n4412 gnd.t300 55.8337
R6925 gnd.n4424 gnd.t291 55.8337
R6926 gnd.n65 gnd.t303 55.8337
R6927 gnd.n30 gnd.t22 55.8337
R6928 gnd.n41 gnd.t298 55.8337
R6929 gnd.n53 gnd.t232 55.8337
R6930 gnd.n1456 gnd.n1455 54.358
R6931 gnd.n3417 gnd.n3416 54.358
R6932 gnd.n4427 gnd.n4426 53.0052
R6933 gnd.n4429 gnd.n4428 53.0052
R6934 gnd.n4431 gnd.n4430 53.0052
R6935 gnd.n4433 gnd.n4432 53.0052
R6936 gnd.n4435 gnd.n4434 53.0052
R6937 gnd.n4392 gnd.n4391 53.0052
R6938 gnd.n4394 gnd.n4393 53.0052
R6939 gnd.n4396 gnd.n4395 53.0052
R6940 gnd.n4398 gnd.n4397 53.0052
R6941 gnd.n4400 gnd.n4399 53.0052
R6942 gnd.n4403 gnd.n4402 53.0052
R6943 gnd.n4405 gnd.n4404 53.0052
R6944 gnd.n4407 gnd.n4406 53.0052
R6945 gnd.n4409 gnd.n4408 53.0052
R6946 gnd.n4411 gnd.n4410 53.0052
R6947 gnd.n4415 gnd.n4414 53.0052
R6948 gnd.n4417 gnd.n4416 53.0052
R6949 gnd.n4419 gnd.n4418 53.0052
R6950 gnd.n4421 gnd.n4420 53.0052
R6951 gnd.n4423 gnd.n4422 53.0052
R6952 gnd.n64 gnd.n63 53.0052
R6953 gnd.n62 gnd.n61 53.0052
R6954 gnd.n60 gnd.n59 53.0052
R6955 gnd.n58 gnd.n57 53.0052
R6956 gnd.n56 gnd.n55 53.0052
R6957 gnd.n29 gnd.n28 53.0052
R6958 gnd.n27 gnd.n26 53.0052
R6959 gnd.n25 gnd.n24 53.0052
R6960 gnd.n23 gnd.n22 53.0052
R6961 gnd.n21 gnd.n20 53.0052
R6962 gnd.n40 gnd.n39 53.0052
R6963 gnd.n38 gnd.n37 53.0052
R6964 gnd.n36 gnd.n35 53.0052
R6965 gnd.n34 gnd.n33 53.0052
R6966 gnd.n32 gnd.n31 53.0052
R6967 gnd.n52 gnd.n51 53.0052
R6968 gnd.n50 gnd.n49 53.0052
R6969 gnd.n48 gnd.n47 53.0052
R6970 gnd.n46 gnd.n45 53.0052
R6971 gnd.n44 gnd.n43 53.0052
R6972 gnd.n3408 gnd.n3407 52.4801
R6973 gnd.n5472 gnd.t215 52.3082
R6974 gnd.n5440 gnd.t326 52.3082
R6975 gnd.n5408 gnd.t319 52.3082
R6976 gnd.n5377 gnd.t225 52.3082
R6977 gnd.n5345 gnd.t228 52.3082
R6978 gnd.n5313 gnd.t39 52.3082
R6979 gnd.n5281 gnd.t211 52.3082
R6980 gnd.n5250 gnd.t243 52.3082
R6981 gnd.n6323 gnd.n6322 52.2881
R6982 gnd.n5621 gnd.n5620 51.9414
R6983 gnd.n5302 gnd.n5270 51.4173
R6984 gnd.n5366 gnd.n5365 50.455
R6985 gnd.n5334 gnd.n5333 50.455
R6986 gnd.n5302 gnd.n5301 50.455
R6987 gnd.n4715 gnd.n4714 45.1884
R6988 gnd.n4225 gnd.n4224 45.1884
R6989 gnd.n3491 gnd.n3423 44.3322
R6990 gnd.n1459 gnd.n1458 44.3189
R6991 gnd.n2143 gnd.n2142 42.4732
R6992 gnd.n443 gnd.n442 42.4732
R6993 gnd.n6385 gnd.n6384 42.2793
R6994 gnd.n6738 gnd.n6737 42.2793
R6995 gnd.n6978 gnd.n6920 42.2793
R6996 gnd.n7020 gnd.n7019 42.2793
R6997 gnd.n6514 gnd.n342 42.2793
R6998 gnd.n6477 gnd.n365 42.2793
R6999 gnd.n6437 gnd.n387 42.2793
R7000 gnd.n6753 gnd.n6752 42.2793
R7001 gnd.n4716 gnd.n4715 42.2793
R7002 gnd.n4226 gnd.n4225 42.2793
R7003 gnd.n4642 gnd.n4641 42.2793
R7004 gnd.n5587 gnd.n4199 42.2793
R7005 gnd.n2571 gnd.n2147 42.2793
R7006 gnd.n2362 gnd.n2312 42.2793
R7007 gnd.n4137 gnd.n1084 42.2793
R7008 gnd.n4097 gnd.n1106 42.2793
R7009 gnd.n4057 gnd.n1128 42.2793
R7010 gnd.n3886 gnd.n1397 42.2793
R7011 gnd.n2154 gnd.n2153 42.2793
R7012 gnd.n2166 gnd.n2165 42.2793
R7013 gnd.n1457 gnd.n1456 41.6274
R7014 gnd.n3418 gnd.n3417 41.6274
R7015 gnd.n1466 gnd.n1465 40.8975
R7016 gnd.n3421 gnd.n3420 40.8975
R7017 gnd.n1465 gnd.n1464 35.055
R7018 gnd.n1460 gnd.n1459 35.055
R7019 gnd.n3410 gnd.n3409 35.055
R7020 gnd.n3420 gnd.n3406 35.055
R7021 gnd.n5789 gnd.n5788 32.3154
R7022 gnd.n5788 gnd.n840 32.3154
R7023 gnd.n5782 gnd.n840 32.3154
R7024 gnd.n5782 gnd.n5781 32.3154
R7025 gnd.n5781 gnd.n5780 32.3154
R7026 gnd.n5780 gnd.n848 32.3154
R7027 gnd.n5774 gnd.n848 32.3154
R7028 gnd.n5774 gnd.n5773 32.3154
R7029 gnd.n5773 gnd.n5772 32.3154
R7030 gnd.n5772 gnd.n856 32.3154
R7031 gnd.n5766 gnd.n856 32.3154
R7032 gnd.n5766 gnd.n5765 32.3154
R7033 gnd.n5765 gnd.n5764 32.3154
R7034 gnd.n5764 gnd.n864 32.3154
R7035 gnd.n5758 gnd.n864 32.3154
R7036 gnd.n5758 gnd.n5757 32.3154
R7037 gnd.n5757 gnd.n5756 32.3154
R7038 gnd.n5756 gnd.n872 32.3154
R7039 gnd.n5750 gnd.n872 32.3154
R7040 gnd.n5750 gnd.n5749 32.3154
R7041 gnd.n5749 gnd.n5748 32.3154
R7042 gnd.n5748 gnd.n880 32.3154
R7043 gnd.n5742 gnd.n880 32.3154
R7044 gnd.n5742 gnd.n5741 32.3154
R7045 gnd.n5741 gnd.n5740 32.3154
R7046 gnd.n5740 gnd.n888 32.3154
R7047 gnd.n5734 gnd.n888 32.3154
R7048 gnd.n5734 gnd.n5733 32.3154
R7049 gnd.n5733 gnd.n5732 32.3154
R7050 gnd.n5732 gnd.n896 32.3154
R7051 gnd.n5726 gnd.n896 32.3154
R7052 gnd.n5726 gnd.n5725 32.3154
R7053 gnd.n5725 gnd.n5724 32.3154
R7054 gnd.n5724 gnd.n904 32.3154
R7055 gnd.n5718 gnd.n904 32.3154
R7056 gnd.n5718 gnd.n5717 32.3154
R7057 gnd.n5717 gnd.n5716 32.3154
R7058 gnd.n5716 gnd.n912 32.3154
R7059 gnd.n5710 gnd.n912 32.3154
R7060 gnd.n5710 gnd.n5709 32.3154
R7061 gnd.n5709 gnd.n5708 32.3154
R7062 gnd.n5708 gnd.n920 32.3154
R7063 gnd.n5702 gnd.n920 32.3154
R7064 gnd.n5702 gnd.n5701 32.3154
R7065 gnd.n5701 gnd.n5700 32.3154
R7066 gnd.n5700 gnd.n928 32.3154
R7067 gnd.n5694 gnd.n928 32.3154
R7068 gnd.n5694 gnd.n5693 32.3154
R7069 gnd.n5693 gnd.n5692 32.3154
R7070 gnd.n5692 gnd.n936 32.3154
R7071 gnd.n5686 gnd.n936 32.3154
R7072 gnd.n5686 gnd.n5685 32.3154
R7073 gnd.n5685 gnd.n5684 32.3154
R7074 gnd.n5684 gnd.n944 32.3154
R7075 gnd.n5678 gnd.n944 32.3154
R7076 gnd.n5678 gnd.n5677 32.3154
R7077 gnd.n5677 gnd.n5676 32.3154
R7078 gnd.n5676 gnd.n952 32.3154
R7079 gnd.n5670 gnd.n952 32.3154
R7080 gnd.n5670 gnd.n5669 32.3154
R7081 gnd.n5669 gnd.n5668 32.3154
R7082 gnd.n5668 gnd.n960 32.3154
R7083 gnd.n5662 gnd.n960 32.3154
R7084 gnd.n5662 gnd.n5661 32.3154
R7085 gnd.n5661 gnd.n5660 32.3154
R7086 gnd.n5660 gnd.n968 32.3154
R7087 gnd.n5654 gnd.n968 32.3154
R7088 gnd.n5654 gnd.n5653 32.3154
R7089 gnd.n5653 gnd.n5652 32.3154
R7090 gnd.n5652 gnd.n976 32.3154
R7091 gnd.n5646 gnd.n976 32.3154
R7092 gnd.n5646 gnd.n5645 32.3154
R7093 gnd.n5645 gnd.n5644 32.3154
R7094 gnd.n5644 gnd.n984 32.3154
R7095 gnd.n5638 gnd.n984 32.3154
R7096 gnd.n5638 gnd.n5637 32.3154
R7097 gnd.n5637 gnd.n5636 32.3154
R7098 gnd.n5636 gnd.n992 32.3154
R7099 gnd.n5630 gnd.n992 32.3154
R7100 gnd.n5630 gnd.n5629 32.3154
R7101 gnd.n5629 gnd.n5628 32.3154
R7102 gnd.n5628 gnd.n1000 32.3154
R7103 gnd.n5622 gnd.n1000 32.3154
R7104 gnd.n4778 gnd.n4672 31.8661
R7105 gnd.n4778 gnd.n4777 31.8661
R7106 gnd.n4786 gnd.n4661 31.8661
R7107 gnd.n4794 gnd.n4661 31.8661
R7108 gnd.n4794 gnd.n4655 31.8661
R7109 gnd.n4802 gnd.n4655 31.8661
R7110 gnd.n4802 gnd.n4648 31.8661
R7111 gnd.n4840 gnd.n4648 31.8661
R7112 gnd.n4850 gnd.n4581 31.8661
R7113 gnd.n4049 gnd.n1061 31.8661
R7114 gnd.n4041 gnd.n1146 31.8661
R7115 gnd.n4041 gnd.n1149 31.8661
R7116 gnd.n4035 gnd.n1149 31.8661
R7117 gnd.n4035 gnd.n1159 31.8661
R7118 gnd.n4029 gnd.n1168 31.8661
R7119 gnd.n4023 gnd.n1168 31.8661
R7120 gnd.n4017 gnd.n1184 31.8661
R7121 gnd.n4011 gnd.n1193 31.8661
R7122 gnd.n4011 gnd.n1196 31.8661
R7123 gnd.n4005 gnd.n1206 31.8661
R7124 gnd.n3999 gnd.n1206 31.8661
R7125 gnd.n3993 gnd.n1222 31.8661
R7126 gnd.n3987 gnd.n1231 31.8661
R7127 gnd.n3987 gnd.n1234 31.8661
R7128 gnd.n3981 gnd.n1244 31.8661
R7129 gnd.n3975 gnd.n1253 31.8661
R7130 gnd.n3969 gnd.n1253 31.8661
R7131 gnd.n3963 gnd.n1269 31.8661
R7132 gnd.n3963 gnd.n1272 31.8661
R7133 gnd.n3957 gnd.n1282 31.8661
R7134 gnd.n3945 gnd.n1299 31.8661
R7135 gnd.n2566 gnd.n1339 31.8661
R7136 gnd.n2559 gnd.n1350 31.8661
R7137 gnd.n2559 gnd.n2558 31.8661
R7138 gnd.n2555 gnd.n2077 31.8661
R7139 gnd.n470 gnd.n458 31.8661
R7140 gnd.n6354 gnd.n490 31.8661
R7141 gnd.n490 gnd.n284 31.8661
R7142 gnd.n6346 gnd.n323 31.8661
R7143 gnd.n6610 gnd.n239 31.8661
R7144 gnd.n6629 gnd.n221 31.8661
R7145 gnd.n6645 gnd.n209 31.8661
R7146 gnd.n6645 gnd.n212 31.8661
R7147 gnd.n6655 gnd.n194 31.8661
R7148 gnd.n6668 gnd.n194 31.8661
R7149 gnd.n6677 gnd.n188 31.8661
R7150 gnd.n6688 gnd.n171 31.8661
R7151 gnd.n6696 gnd.n171 31.8661
R7152 gnd.n7123 gnd.n74 31.8661
R7153 gnd.n7117 gnd.n86 31.8661
R7154 gnd.n7111 gnd.n86 31.8661
R7155 gnd.n7105 gnd.n104 31.8661
R7156 gnd.n7105 gnd.n107 31.8661
R7157 gnd.n7099 gnd.n116 31.8661
R7158 gnd.n7093 gnd.n126 31.8661
R7159 gnd.n7087 gnd.n126 31.8661
R7160 gnd.n7081 gnd.n142 31.8661
R7161 gnd.n7081 gnd.n145 31.8661
R7162 gnd.n7075 gnd.n145 31.8661
R7163 gnd.n7075 gnd.n154 31.8661
R7164 gnd.n7069 gnd.n164 31.8661
R7165 gnd.n1222 gnd.t36 31.5474
R7166 gnd.t222 gnd.n1244 31.5474
R7167 gnd.n6677 gnd.t17 31.5474
R7168 gnd.t40 gnd.n74 31.5474
R7169 gnd.n1184 gnd.t195 30.9101
R7170 gnd.t31 gnd.n1282 30.9101
R7171 gnd.t2 gnd.n221 30.9101
R7172 gnd.n3497 gnd.n1673 30.7517
R7173 gnd.n2891 gnd.n2839 30.7517
R7174 gnd.n3939 gnd.n1309 28.6795
R7175 gnd.n2505 gnd.n1312 28.6795
R7176 gnd.n3933 gnd.n1320 28.6795
R7177 gnd.n2535 gnd.n1323 28.6795
R7178 gnd.n2567 gnd.n1332 28.6795
R7179 gnd.n6345 gnd.n274 28.6795
R7180 gnd.n6339 gnd.n267 28.6795
R7181 gnd.n6565 gnd.n255 28.6795
R7182 gnd.n6581 gnd.n258 28.6795
R7183 gnd.n6569 gnd.n246 28.6795
R7184 gnd.n3919 gnd.n1339 28.0422
R7185 gnd.n6546 gnd.n323 28.0422
R7186 gnd.n2142 gnd.n2141 25.7944
R7187 gnd.n6384 gnd.n6383 25.7944
R7188 gnd.n6737 gnd.n6736 25.7944
R7189 gnd.n6920 gnd.n6919 25.7944
R7190 gnd.n7019 gnd.n7018 25.7944
R7191 gnd.n342 gnd.n341 25.7944
R7192 gnd.n365 gnd.n364 25.7944
R7193 gnd.n387 gnd.n386 25.7944
R7194 gnd.n6752 gnd.n6751 25.7944
R7195 gnd.n4641 gnd.n4640 25.7944
R7196 gnd.n4199 gnd.n4198 25.7944
R7197 gnd.n2147 gnd.n2146 25.7944
R7198 gnd.n2312 gnd.n2311 25.7944
R7199 gnd.n1084 gnd.n1083 25.7944
R7200 gnd.n1106 gnd.n1105 25.7944
R7201 gnd.n1128 gnd.n1127 25.7944
R7202 gnd.n1397 gnd.n1396 25.7944
R7203 gnd.n2153 gnd.n2152 25.7944
R7204 gnd.n2165 gnd.n2164 25.7944
R7205 gnd.n442 gnd.n441 25.7944
R7206 gnd.n4862 gnd.n4582 24.8557
R7207 gnd.n4872 gnd.n4565 24.8557
R7208 gnd.n4568 gnd.n4556 24.8557
R7209 gnd.n4893 gnd.n4557 24.8557
R7210 gnd.n4903 gnd.n4537 24.8557
R7211 gnd.n4913 gnd.n4912 24.8557
R7212 gnd.n4523 gnd.n4521 24.8557
R7213 gnd.n4944 gnd.n4943 24.8557
R7214 gnd.n4959 gnd.n4506 24.8557
R7215 gnd.n5013 gnd.n4445 24.8557
R7216 gnd.n4969 gnd.n4446 24.8557
R7217 gnd.n5006 gnd.n4457 24.8557
R7218 gnd.n4495 gnd.n4494 24.8557
R7219 gnd.n5000 gnd.n4999 24.8557
R7220 gnd.n4481 gnd.n4468 24.8557
R7221 gnd.n5039 gnd.n5038 24.8557
R7222 gnd.n5049 gnd.n4377 24.8557
R7223 gnd.n5061 gnd.n4369 24.8557
R7224 gnd.n5060 gnd.n4357 24.8557
R7225 gnd.n5079 gnd.n5078 24.8557
R7226 gnd.n5089 gnd.n4350 24.8557
R7227 gnd.n5100 gnd.n4338 24.8557
R7228 gnd.n5124 gnd.n5123 24.8557
R7229 gnd.n5135 gnd.n4321 24.8557
R7230 gnd.n5134 gnd.n4323 24.8557
R7231 gnd.n5146 gnd.n4314 24.8557
R7232 gnd.n5164 gnd.n5163 24.8557
R7233 gnd.n4305 gnd.n4294 24.8557
R7234 gnd.n5185 gnd.n4282 24.8557
R7235 gnd.n5213 gnd.n5212 24.8557
R7236 gnd.n5224 gnd.n4267 24.8557
R7237 gnd.n5235 gnd.n4260 24.8557
R7238 gnd.n5234 gnd.n4248 24.8557
R7239 gnd.n5507 gnd.n5506 24.8557
R7240 gnd.n5529 gnd.n4233 24.8557
R7241 gnd.n2558 gnd.n2557 23.8997
R7242 gnd.n6355 gnd.n6354 23.8997
R7243 gnd.n4883 gnd.t242 23.2624
R7244 gnd.n4584 gnd.t125 22.6251
R7245 gnd.n6322 gnd.t200 22.3064
R7246 gnd.n4017 gnd.t6 21.9878
R7247 gnd.n3957 gnd.t9 21.9878
R7248 gnd.n6629 gnd.t15 21.9878
R7249 gnd.n7099 gnd.t13 21.9878
R7250 gnd.t224 gnd.n4589 21.3504
R7251 gnd.n3993 gnd.t26 21.3504
R7252 gnd.n3981 gnd.t11 21.3504
R7253 gnd.n188 gnd.t181 21.3504
R7254 gnd.n7123 gnd.t33 21.3504
R7255 gnd.t275 gnd.n4295 20.7131
R7256 gnd.n4005 gnd.t206 20.7131
R7257 gnd.n3969 gnd.t47 20.7131
R7258 gnd.n6655 gnd.t54 20.7131
R7259 gnd.n7111 gnd.t254 20.7131
R7260 gnd.t273 gnd.n4330 20.0758
R7261 gnd.n4029 gnd.t52 20.0758
R7262 gnd.n7087 gnd.t21 20.0758
R7263 gnd.n2777 gnd.n2776 19.9763
R7264 gnd.n1672 gnd.n1671 19.9763
R7265 gnd.n3801 gnd.n3800 19.9763
R7266 gnd.n3425 gnd.n3424 19.9763
R7267 gnd.n1454 gnd.t163 19.8005
R7268 gnd.n1454 gnd.t176 19.8005
R7269 gnd.n1453 gnd.t117 19.8005
R7270 gnd.n1453 gnd.t71 19.8005
R7271 gnd.n3415 gnd.t89 19.8005
R7272 gnd.n3415 gnd.t133 19.8005
R7273 gnd.n3414 gnd.t104 19.8005
R7274 gnd.n3414 gnd.t139 19.8005
R7275 gnd.n1450 gnd.n1449 19.5087
R7276 gnd.n1463 gnd.n1450 19.5087
R7277 gnd.n1461 gnd.n1452 19.5087
R7278 gnd.n3419 gnd.n3413 19.5087
R7279 gnd.n5050 gnd.t266 19.4385
R7280 gnd.n2637 gnd.n2073 19.3944
R7281 gnd.n2642 gnd.n2073 19.3944
R7282 gnd.n2642 gnd.n2074 19.3944
R7283 gnd.n2074 gnd.n2051 19.3944
R7284 gnd.n2667 gnd.n2051 19.3944
R7285 gnd.n2667 gnd.n2048 19.3944
R7286 gnd.n2672 gnd.n2048 19.3944
R7287 gnd.n2672 gnd.n2049 19.3944
R7288 gnd.n2049 gnd.n2025 19.3944
R7289 gnd.n2697 gnd.n2025 19.3944
R7290 gnd.n2697 gnd.n2022 19.3944
R7291 gnd.n2702 gnd.n2022 19.3944
R7292 gnd.n2702 gnd.n2023 19.3944
R7293 gnd.n2023 gnd.n2001 19.3944
R7294 gnd.n2727 gnd.n2001 19.3944
R7295 gnd.n2727 gnd.n1998 19.3944
R7296 gnd.n2736 gnd.n1998 19.3944
R7297 gnd.n2736 gnd.n1999 19.3944
R7298 gnd.n2732 gnd.n1999 19.3944
R7299 gnd.n2732 gnd.n1978 19.3944
R7300 gnd.n1978 gnd.n1976 19.3944
R7301 gnd.n2896 gnd.n1976 19.3944
R7302 gnd.n2897 gnd.n2896 19.3944
R7303 gnd.n2897 gnd.n1973 19.3944
R7304 gnd.n2902 gnd.n1973 19.3944
R7305 gnd.n2902 gnd.n1974 19.3944
R7306 gnd.n1974 gnd.n1949 19.3944
R7307 gnd.n2934 gnd.n1949 19.3944
R7308 gnd.n2934 gnd.n1947 19.3944
R7309 gnd.n2938 gnd.n1947 19.3944
R7310 gnd.n2938 gnd.n1930 19.3944
R7311 gnd.n2963 gnd.n1930 19.3944
R7312 gnd.n2963 gnd.n1927 19.3944
R7313 gnd.n2968 gnd.n1927 19.3944
R7314 gnd.n2968 gnd.n1928 19.3944
R7315 gnd.n1928 gnd.n1901 19.3944
R7316 gnd.n3002 gnd.n1901 19.3944
R7317 gnd.n3002 gnd.n1898 19.3944
R7318 gnd.n3021 gnd.n1898 19.3944
R7319 gnd.n3021 gnd.n1899 19.3944
R7320 gnd.n3017 gnd.n1899 19.3944
R7321 gnd.n3017 gnd.n3016 19.3944
R7322 gnd.n3016 gnd.n3015 19.3944
R7323 gnd.n3015 gnd.n3009 19.3944
R7324 gnd.n3011 gnd.n3009 19.3944
R7325 gnd.n3011 gnd.n1853 19.3944
R7326 gnd.n3086 gnd.n1853 19.3944
R7327 gnd.n3087 gnd.n3086 19.3944
R7328 gnd.n3087 gnd.n1851 19.3944
R7329 gnd.n3091 gnd.n1851 19.3944
R7330 gnd.n3091 gnd.n1828 19.3944
R7331 gnd.n3141 gnd.n1828 19.3944
R7332 gnd.n3141 gnd.n1829 19.3944
R7333 gnd.n3137 gnd.n1829 19.3944
R7334 gnd.n3137 gnd.n1805 19.3944
R7335 gnd.n3181 gnd.n1805 19.3944
R7336 gnd.n3181 gnd.n1806 19.3944
R7337 gnd.n3177 gnd.n1806 19.3944
R7338 gnd.n3177 gnd.n1782 19.3944
R7339 gnd.n3230 gnd.n1782 19.3944
R7340 gnd.n3230 gnd.n1783 19.3944
R7341 gnd.n3226 gnd.n1783 19.3944
R7342 gnd.n3226 gnd.n3225 19.3944
R7343 gnd.n3225 gnd.n3224 19.3944
R7344 gnd.n3224 gnd.n3221 19.3944
R7345 gnd.n3221 gnd.n1734 19.3944
R7346 gnd.n3295 gnd.n1734 19.3944
R7347 gnd.n3295 gnd.n1731 19.3944
R7348 gnd.n3300 gnd.n1731 19.3944
R7349 gnd.n3300 gnd.n1732 19.3944
R7350 gnd.n1732 gnd.n1708 19.3944
R7351 gnd.n3350 gnd.n1708 19.3944
R7352 gnd.n3350 gnd.n1705 19.3944
R7353 gnd.n3363 gnd.n1705 19.3944
R7354 gnd.n3363 gnd.n1706 19.3944
R7355 gnd.n3359 gnd.n1706 19.3944
R7356 gnd.n3359 gnd.n3358 19.3944
R7357 gnd.n3358 gnd.n3357 19.3944
R7358 gnd.n3357 gnd.n1634 19.3944
R7359 gnd.n3567 gnd.n1634 19.3944
R7360 gnd.n3567 gnd.n1632 19.3944
R7361 gnd.n3571 gnd.n1632 19.3944
R7362 gnd.n3571 gnd.n1622 19.3944
R7363 gnd.n3589 gnd.n1622 19.3944
R7364 gnd.n3589 gnd.n1620 19.3944
R7365 gnd.n3593 gnd.n1620 19.3944
R7366 gnd.n3593 gnd.n1611 19.3944
R7367 gnd.n3610 gnd.n1611 19.3944
R7368 gnd.n3610 gnd.n1609 19.3944
R7369 gnd.n3614 gnd.n1609 19.3944
R7370 gnd.n3614 gnd.n1599 19.3944
R7371 gnd.n3631 gnd.n1599 19.3944
R7372 gnd.n3631 gnd.n1597 19.3944
R7373 gnd.n3635 gnd.n1597 19.3944
R7374 gnd.n3635 gnd.n1587 19.3944
R7375 gnd.n3652 gnd.n1587 19.3944
R7376 gnd.n3652 gnd.n1584 19.3944
R7377 gnd.n3657 gnd.n1584 19.3944
R7378 gnd.n3657 gnd.n1585 19.3944
R7379 gnd.n1585 gnd.n454 19.3944
R7380 gnd.n6373 gnd.n454 19.3944
R7381 gnd.n2280 gnd.n2278 19.3944
R7382 gnd.n2543 gnd.n2280 19.3944
R7383 gnd.n2543 gnd.n2281 19.3944
R7384 gnd.n2629 gnd.n2628 19.3944
R7385 gnd.n2628 gnd.n2627 19.3944
R7386 gnd.n2627 gnd.n2085 19.3944
R7387 gnd.n2623 gnd.n2085 19.3944
R7388 gnd.n2623 gnd.n2622 19.3944
R7389 gnd.n2622 gnd.n2621 19.3944
R7390 gnd.n2621 gnd.n2090 19.3944
R7391 gnd.n2616 gnd.n2090 19.3944
R7392 gnd.n2616 gnd.n2615 19.3944
R7393 gnd.n2615 gnd.n2095 19.3944
R7394 gnd.n2608 gnd.n2095 19.3944
R7395 gnd.n2608 gnd.n2607 19.3944
R7396 gnd.n2607 gnd.n2105 19.3944
R7397 gnd.n2600 gnd.n2105 19.3944
R7398 gnd.n2600 gnd.n2599 19.3944
R7399 gnd.n2599 gnd.n2113 19.3944
R7400 gnd.n2592 gnd.n2113 19.3944
R7401 gnd.n2592 gnd.n2591 19.3944
R7402 gnd.n2591 gnd.n2123 19.3944
R7403 gnd.n2584 gnd.n2123 19.3944
R7404 gnd.n2584 gnd.n2583 19.3944
R7405 gnd.n2583 gnd.n2131 19.3944
R7406 gnd.n2576 gnd.n2131 19.3944
R7407 gnd.n2576 gnd.n2575 19.3944
R7408 gnd.n6426 gnd.n398 19.3944
R7409 gnd.n6426 gnd.n6425 19.3944
R7410 gnd.n6425 gnd.n401 19.3944
R7411 gnd.n6418 gnd.n401 19.3944
R7412 gnd.n6418 gnd.n6417 19.3944
R7413 gnd.n6417 gnd.n411 19.3944
R7414 gnd.n6410 gnd.n411 19.3944
R7415 gnd.n6410 gnd.n6409 19.3944
R7416 gnd.n6409 gnd.n419 19.3944
R7417 gnd.n6402 gnd.n419 19.3944
R7418 gnd.n6402 gnd.n6401 19.3944
R7419 gnd.n6401 gnd.n429 19.3944
R7420 gnd.n6394 gnd.n429 19.3944
R7421 gnd.n6394 gnd.n6393 19.3944
R7422 gnd.n6393 gnd.n437 19.3944
R7423 gnd.n6386 gnd.n437 19.3944
R7424 gnd.n504 gnd.n503 19.3944
R7425 gnd.n504 gnd.n264 19.3944
R7426 gnd.n6567 gnd.n264 19.3944
R7427 gnd.n6568 gnd.n6567 19.3944
R7428 gnd.n6571 gnd.n6568 19.3944
R7429 gnd.n6572 gnd.n6571 19.3944
R7430 gnd.n6572 gnd.n236 19.3944
R7431 gnd.n6612 gnd.n236 19.3944
R7432 gnd.n6613 gnd.n6612 19.3944
R7433 gnd.n6614 gnd.n6613 19.3944
R7434 gnd.n6614 gnd.n218 19.3944
R7435 gnd.n6632 gnd.n218 19.3944
R7436 gnd.n6633 gnd.n6632 19.3944
R7437 gnd.n6635 gnd.n6633 19.3944
R7438 gnd.n6636 gnd.n6635 19.3944
R7439 gnd.n6636 gnd.n192 19.3944
R7440 gnd.n6670 gnd.n192 19.3944
R7441 gnd.n6673 gnd.n6670 19.3944
R7442 gnd.n6673 gnd.n6672 19.3944
R7443 gnd.n6672 gnd.n173 19.3944
R7444 gnd.n6693 gnd.n173 19.3944
R7445 gnd.n6694 gnd.n6693 19.3944
R7446 gnd.n6694 gnd.n167 19.3944
R7447 gnd.n6703 gnd.n167 19.3944
R7448 gnd.n6704 gnd.n6703 19.3944
R7449 gnd.n6706 gnd.n6704 19.3944
R7450 gnd.n6707 gnd.n6706 19.3944
R7451 gnd.n6710 gnd.n6707 19.3944
R7452 gnd.n6711 gnd.n6710 19.3944
R7453 gnd.n6713 gnd.n6711 19.3944
R7454 gnd.n6714 gnd.n6713 19.3944
R7455 gnd.n6717 gnd.n6714 19.3944
R7456 gnd.n6718 gnd.n6717 19.3944
R7457 gnd.n6720 gnd.n6718 19.3944
R7458 gnd.n6721 gnd.n6720 19.3944
R7459 gnd.n6724 gnd.n6721 19.3944
R7460 gnd.n6725 gnd.n6724 19.3944
R7461 gnd.n6727 gnd.n6725 19.3944
R7462 gnd.n6728 gnd.n6727 19.3944
R7463 gnd.n6731 gnd.n6728 19.3944
R7464 gnd.n6732 gnd.n6731 19.3944
R7465 gnd.n6733 gnd.n6732 19.3944
R7466 gnd.n6974 gnd.n6918 19.3944
R7467 gnd.n6974 gnd.n6971 19.3944
R7468 gnd.n6971 gnd.n6968 19.3944
R7469 gnd.n6968 gnd.n6967 19.3944
R7470 gnd.n6967 gnd.n6964 19.3944
R7471 gnd.n6964 gnd.n6963 19.3944
R7472 gnd.n6963 gnd.n6960 19.3944
R7473 gnd.n6960 gnd.n6959 19.3944
R7474 gnd.n6959 gnd.n6956 19.3944
R7475 gnd.n6956 gnd.n6955 19.3944
R7476 gnd.n6955 gnd.n6952 19.3944
R7477 gnd.n6952 gnd.n6951 19.3944
R7478 gnd.n6951 gnd.n6948 19.3944
R7479 gnd.n6948 gnd.n6947 19.3944
R7480 gnd.n6947 gnd.n6944 19.3944
R7481 gnd.n6944 gnd.n6943 19.3944
R7482 gnd.n6943 gnd.n6940 19.3944
R7483 gnd.n6940 gnd.n6939 19.3944
R7484 gnd.n7017 gnd.n7014 19.3944
R7485 gnd.n7014 gnd.n7013 19.3944
R7486 gnd.n7013 gnd.n7010 19.3944
R7487 gnd.n7010 gnd.n7009 19.3944
R7488 gnd.n7009 gnd.n7006 19.3944
R7489 gnd.n7006 gnd.n7005 19.3944
R7490 gnd.n7005 gnd.n7002 19.3944
R7491 gnd.n7002 gnd.n7001 19.3944
R7492 gnd.n7001 gnd.n6998 19.3944
R7493 gnd.n6998 gnd.n6997 19.3944
R7494 gnd.n6997 gnd.n6994 19.3944
R7495 gnd.n6994 gnd.n6993 19.3944
R7496 gnd.n6993 gnd.n6990 19.3944
R7497 gnd.n6990 gnd.n6989 19.3944
R7498 gnd.n6989 gnd.n6986 19.3944
R7499 gnd.n6986 gnd.n6985 19.3944
R7500 gnd.n6985 gnd.n6982 19.3944
R7501 gnd.n6982 gnd.n6981 19.3944
R7502 gnd.n7056 gnd.n7055 19.3944
R7503 gnd.n7055 gnd.n6884 19.3944
R7504 gnd.n7051 gnd.n6884 19.3944
R7505 gnd.n7051 gnd.n7048 19.3944
R7506 gnd.n7048 gnd.n7045 19.3944
R7507 gnd.n7045 gnd.n7044 19.3944
R7508 gnd.n7044 gnd.n7041 19.3944
R7509 gnd.n7041 gnd.n7040 19.3944
R7510 gnd.n7040 gnd.n7037 19.3944
R7511 gnd.n7037 gnd.n7036 19.3944
R7512 gnd.n7036 gnd.n7033 19.3944
R7513 gnd.n7033 gnd.n7032 19.3944
R7514 gnd.n7032 gnd.n7029 19.3944
R7515 gnd.n7029 gnd.n7028 19.3944
R7516 gnd.n7028 gnd.n7025 19.3944
R7517 gnd.n7025 gnd.n7024 19.3944
R7518 gnd.n7024 gnd.n7021 19.3944
R7519 gnd.n6554 gnd.n279 19.3944
R7520 gnd.n6554 gnd.n280 19.3944
R7521 gnd.n280 gnd.n253 19.3944
R7522 gnd.n6583 gnd.n253 19.3944
R7523 gnd.n6583 gnd.n251 19.3944
R7524 gnd.n6589 gnd.n251 19.3944
R7525 gnd.n6589 gnd.n6588 19.3944
R7526 gnd.n6588 gnd.n227 19.3944
R7527 gnd.n6623 gnd.n227 19.3944
R7528 gnd.n6623 gnd.n225 19.3944
R7529 gnd.n6627 gnd.n225 19.3944
R7530 gnd.n6627 gnd.n207 19.3944
R7531 gnd.n6647 gnd.n207 19.3944
R7532 gnd.n6647 gnd.n205 19.3944
R7533 gnd.n6653 gnd.n205 19.3944
R7534 gnd.n6653 gnd.n6652 19.3944
R7535 gnd.n6652 gnd.n184 19.3944
R7536 gnd.n6679 gnd.n184 19.3944
R7537 gnd.n6679 gnd.n182 19.3944
R7538 gnd.n6686 gnd.n182 19.3944
R7539 gnd.n6686 gnd.n6685 19.3944
R7540 gnd.n6685 gnd.n78 19.3944
R7541 gnd.n7121 gnd.n78 19.3944
R7542 gnd.n7121 gnd.n7120 19.3944
R7543 gnd.n7120 gnd.n7119 19.3944
R7544 gnd.n7119 gnd.n82 19.3944
R7545 gnd.n7109 gnd.n82 19.3944
R7546 gnd.n7109 gnd.n7108 19.3944
R7547 gnd.n7108 gnd.n7107 19.3944
R7548 gnd.n7107 gnd.n102 19.3944
R7549 gnd.n7097 gnd.n102 19.3944
R7550 gnd.n7097 gnd.n7096 19.3944
R7551 gnd.n7096 gnd.n7095 19.3944
R7552 gnd.n7095 gnd.n122 19.3944
R7553 gnd.n7085 gnd.n122 19.3944
R7554 gnd.n7085 gnd.n7084 19.3944
R7555 gnd.n7084 gnd.n7083 19.3944
R7556 gnd.n7083 gnd.n140 19.3944
R7557 gnd.n7073 gnd.n140 19.3944
R7558 gnd.n7073 gnd.n7072 19.3944
R7559 gnd.n7072 gnd.n7071 19.3944
R7560 gnd.n7071 gnd.n160 19.3944
R7561 gnd.n6549 gnd.n282 19.3944
R7562 gnd.n6544 gnd.n282 19.3944
R7563 gnd.n6544 gnd.n6543 19.3944
R7564 gnd.n6543 gnd.n6542 19.3944
R7565 gnd.n6542 gnd.n6539 19.3944
R7566 gnd.n6539 gnd.n6538 19.3944
R7567 gnd.n6538 gnd.n6535 19.3944
R7568 gnd.n6535 gnd.n6534 19.3944
R7569 gnd.n6534 gnd.n6531 19.3944
R7570 gnd.n6531 gnd.n6530 19.3944
R7571 gnd.n6530 gnd.n6527 19.3944
R7572 gnd.n6527 gnd.n6526 19.3944
R7573 gnd.n6526 gnd.n6523 19.3944
R7574 gnd.n6523 gnd.n6522 19.3944
R7575 gnd.n6522 gnd.n6519 19.3944
R7576 gnd.n6519 gnd.n6518 19.3944
R7577 gnd.n6518 gnd.n6515 19.3944
R7578 gnd.n6513 gnd.n6510 19.3944
R7579 gnd.n6510 gnd.n6509 19.3944
R7580 gnd.n6509 gnd.n6506 19.3944
R7581 gnd.n6506 gnd.n6505 19.3944
R7582 gnd.n6505 gnd.n6502 19.3944
R7583 gnd.n6502 gnd.n6501 19.3944
R7584 gnd.n6501 gnd.n6498 19.3944
R7585 gnd.n6496 gnd.n6493 19.3944
R7586 gnd.n6493 gnd.n6492 19.3944
R7587 gnd.n6492 gnd.n6489 19.3944
R7588 gnd.n6489 gnd.n6488 19.3944
R7589 gnd.n6488 gnd.n6485 19.3944
R7590 gnd.n6485 gnd.n6484 19.3944
R7591 gnd.n6484 gnd.n6481 19.3944
R7592 gnd.n6481 gnd.n6480 19.3944
R7593 gnd.n6476 gnd.n6473 19.3944
R7594 gnd.n6473 gnd.n6472 19.3944
R7595 gnd.n6472 gnd.n6469 19.3944
R7596 gnd.n6469 gnd.n6468 19.3944
R7597 gnd.n6468 gnd.n6465 19.3944
R7598 gnd.n6465 gnd.n6464 19.3944
R7599 gnd.n6464 gnd.n6461 19.3944
R7600 gnd.n6461 gnd.n6460 19.3944
R7601 gnd.n6460 gnd.n6457 19.3944
R7602 gnd.n6457 gnd.n6456 19.3944
R7603 gnd.n6456 gnd.n6453 19.3944
R7604 gnd.n6453 gnd.n6452 19.3944
R7605 gnd.n6452 gnd.n6449 19.3944
R7606 gnd.n6449 gnd.n6448 19.3944
R7607 gnd.n6448 gnd.n6445 19.3944
R7608 gnd.n6445 gnd.n6444 19.3944
R7609 gnd.n6444 gnd.n6441 19.3944
R7610 gnd.n6441 gnd.n6440 19.3944
R7611 gnd.n6763 gnd.n6761 19.3944
R7612 gnd.n6766 gnd.n6763 19.3944
R7613 gnd.n6769 gnd.n6766 19.3944
R7614 gnd.n6772 gnd.n6769 19.3944
R7615 gnd.n6772 gnd.n6759 19.3944
R7616 gnd.n6776 gnd.n6759 19.3944
R7617 gnd.n6779 gnd.n6776 19.3944
R7618 gnd.n6782 gnd.n6779 19.3944
R7619 gnd.n6782 gnd.n6757 19.3944
R7620 gnd.n6786 gnd.n6757 19.3944
R7621 gnd.n6789 gnd.n6786 19.3944
R7622 gnd.n6792 gnd.n6789 19.3944
R7623 gnd.n6792 gnd.n6755 19.3944
R7624 gnd.n6796 gnd.n6755 19.3944
R7625 gnd.n6799 gnd.n6796 19.3944
R7626 gnd.n6801 gnd.n6799 19.3944
R7627 gnd.n6558 gnd.n272 19.3944
R7628 gnd.n6558 gnd.n269 19.3944
R7629 gnd.n6563 gnd.n269 19.3944
R7630 gnd.n6563 gnd.n270 19.3944
R7631 gnd.n270 gnd.n244 19.3944
R7632 gnd.n6593 gnd.n244 19.3944
R7633 gnd.n6593 gnd.n241 19.3944
R7634 gnd.n6608 gnd.n241 19.3944
R7635 gnd.n6608 gnd.n242 19.3944
R7636 gnd.n6604 gnd.n242 19.3944
R7637 gnd.n6604 gnd.n6603 19.3944
R7638 gnd.n6603 gnd.n6602 19.3944
R7639 gnd.n6602 gnd.n6599 19.3944
R7640 gnd.n6599 gnd.n199 19.3944
R7641 gnd.n6657 gnd.n199 19.3944
R7642 gnd.n6657 gnd.n196 19.3944
R7643 gnd.n6666 gnd.n196 19.3944
R7644 gnd.n6666 gnd.n197 19.3944
R7645 gnd.n6662 gnd.n197 19.3944
R7646 gnd.n6662 gnd.n6661 19.3944
R7647 gnd.n6661 gnd.n68 19.3944
R7648 gnd.n7126 gnd.n68 19.3944
R7649 gnd.n7126 gnd.n7125 19.3944
R7650 gnd.n7125 gnd.n71 19.3944
R7651 gnd.n6814 gnd.n71 19.3944
R7652 gnd.n6816 gnd.n6814 19.3944
R7653 gnd.n6816 gnd.n6811 19.3944
R7654 gnd.n6821 gnd.n6811 19.3944
R7655 gnd.n6822 gnd.n6821 19.3944
R7656 gnd.n6824 gnd.n6822 19.3944
R7657 gnd.n6824 gnd.n6809 19.3944
R7658 gnd.n6829 gnd.n6809 19.3944
R7659 gnd.n6830 gnd.n6829 19.3944
R7660 gnd.n6832 gnd.n6830 19.3944
R7661 gnd.n6832 gnd.n6807 19.3944
R7662 gnd.n6837 gnd.n6807 19.3944
R7663 gnd.n6838 gnd.n6837 19.3944
R7664 gnd.n6840 gnd.n6838 19.3944
R7665 gnd.n6840 gnd.n6805 19.3944
R7666 gnd.n6845 gnd.n6805 19.3944
R7667 gnd.n6846 gnd.n6845 19.3944
R7668 gnd.n6847 gnd.n6846 19.3944
R7669 gnd.n6343 gnd.n6342 19.3944
R7670 gnd.n6342 gnd.n6341 19.3944
R7671 gnd.n6341 gnd.n261 19.3944
R7672 gnd.n6579 gnd.n261 19.3944
R7673 gnd.n6579 gnd.n6578 19.3944
R7674 gnd.n6578 gnd.n6577 19.3944
R7675 gnd.n6577 gnd.n6576 19.3944
R7676 gnd.n6576 gnd.n234 19.3944
R7677 gnd.n6619 gnd.n234 19.3944
R7678 gnd.n6619 gnd.n6618 19.3944
R7679 gnd.n6618 gnd.n6617 19.3944
R7680 gnd.n6617 gnd.n215 19.3944
R7681 gnd.n6643 gnd.n215 19.3944
R7682 gnd.n6643 gnd.n6642 19.3944
R7683 gnd.n6642 gnd.n6641 19.3944
R7684 gnd.n6641 gnd.n6640 19.3944
R7685 gnd.n6640 gnd.n190 19.3944
R7686 gnd.n6675 gnd.n190 19.3944
R7687 gnd.n6675 gnd.n175 19.3944
R7688 gnd.n6690 gnd.n175 19.3944
R7689 gnd.n6690 gnd.n169 19.3944
R7690 gnd.n6698 gnd.n169 19.3944
R7691 gnd.n6699 gnd.n6698 19.3944
R7692 gnd.n6699 gnd.n89 19.3944
R7693 gnd.n7115 gnd.n89 19.3944
R7694 gnd.n7115 gnd.n7114 19.3944
R7695 gnd.n7114 gnd.n7113 19.3944
R7696 gnd.n7113 gnd.n93 19.3944
R7697 gnd.n7103 gnd.n93 19.3944
R7698 gnd.n7103 gnd.n7102 19.3944
R7699 gnd.n7102 gnd.n7101 19.3944
R7700 gnd.n7101 gnd.n112 19.3944
R7701 gnd.n7091 gnd.n112 19.3944
R7702 gnd.n7091 gnd.n7090 19.3944
R7703 gnd.n7090 gnd.n7089 19.3944
R7704 gnd.n7089 gnd.n131 19.3944
R7705 gnd.n7079 gnd.n131 19.3944
R7706 gnd.n7079 gnd.n7078 19.3944
R7707 gnd.n7078 gnd.n7077 19.3944
R7708 gnd.n7077 gnd.n150 19.3944
R7709 gnd.n7067 gnd.n150 19.3944
R7710 gnd.n7067 gnd.n7066 19.3944
R7711 gnd.n4765 gnd.n4764 19.3944
R7712 gnd.n4764 gnd.n4763 19.3944
R7713 gnd.n4763 gnd.n4762 19.3944
R7714 gnd.n4762 gnd.n4760 19.3944
R7715 gnd.n4760 gnd.n4757 19.3944
R7716 gnd.n4757 gnd.n4756 19.3944
R7717 gnd.n4756 gnd.n4753 19.3944
R7718 gnd.n4753 gnd.n4752 19.3944
R7719 gnd.n4752 gnd.n4749 19.3944
R7720 gnd.n4749 gnd.n4748 19.3944
R7721 gnd.n4748 gnd.n4745 19.3944
R7722 gnd.n4745 gnd.n4744 19.3944
R7723 gnd.n4744 gnd.n4741 19.3944
R7724 gnd.n4741 gnd.n4740 19.3944
R7725 gnd.n4740 gnd.n4737 19.3944
R7726 gnd.n4737 gnd.n4736 19.3944
R7727 gnd.n4736 gnd.n4733 19.3944
R7728 gnd.n4733 gnd.n4732 19.3944
R7729 gnd.n4732 gnd.n4729 19.3944
R7730 gnd.n4729 gnd.n4728 19.3944
R7731 gnd.n4728 gnd.n4725 19.3944
R7732 gnd.n4725 gnd.n4724 19.3944
R7733 gnd.n4721 gnd.n4720 19.3944
R7734 gnd.n4720 gnd.n4676 19.3944
R7735 gnd.n4771 gnd.n4676 19.3944
R7736 gnd.n5537 gnd.n5536 19.3944
R7737 gnd.n5536 gnd.n5533 19.3944
R7738 gnd.n5533 gnd.n5532 19.3944
R7739 gnd.n5582 gnd.n5581 19.3944
R7740 gnd.n5581 gnd.n5580 19.3944
R7741 gnd.n5580 gnd.n5577 19.3944
R7742 gnd.n5577 gnd.n5576 19.3944
R7743 gnd.n5576 gnd.n5573 19.3944
R7744 gnd.n5573 gnd.n5572 19.3944
R7745 gnd.n5572 gnd.n5569 19.3944
R7746 gnd.n5569 gnd.n5568 19.3944
R7747 gnd.n5568 gnd.n5565 19.3944
R7748 gnd.n5565 gnd.n5564 19.3944
R7749 gnd.n5564 gnd.n5561 19.3944
R7750 gnd.n5561 gnd.n5560 19.3944
R7751 gnd.n5560 gnd.n5557 19.3944
R7752 gnd.n5557 gnd.n5556 19.3944
R7753 gnd.n5556 gnd.n5553 19.3944
R7754 gnd.n5553 gnd.n5552 19.3944
R7755 gnd.n5552 gnd.n5549 19.3944
R7756 gnd.n5549 gnd.n5548 19.3944
R7757 gnd.n5548 gnd.n5545 19.3944
R7758 gnd.n5545 gnd.n5544 19.3944
R7759 gnd.n5544 gnd.n5541 19.3944
R7760 gnd.n5541 gnd.n5540 19.3944
R7761 gnd.n4864 gnd.n4573 19.3944
R7762 gnd.n4874 gnd.n4573 19.3944
R7763 gnd.n4875 gnd.n4874 19.3944
R7764 gnd.n4875 gnd.n4554 19.3944
R7765 gnd.n4895 gnd.n4554 19.3944
R7766 gnd.n4895 gnd.n4546 19.3944
R7767 gnd.n4905 gnd.n4546 19.3944
R7768 gnd.n4906 gnd.n4905 19.3944
R7769 gnd.n4907 gnd.n4906 19.3944
R7770 gnd.n4907 gnd.n4529 19.3944
R7771 gnd.n4924 gnd.n4529 19.3944
R7772 gnd.n4927 gnd.n4924 19.3944
R7773 gnd.n4927 gnd.n4926 19.3944
R7774 gnd.n4926 gnd.n4502 19.3944
R7775 gnd.n4966 gnd.n4502 19.3944
R7776 gnd.n4966 gnd.n4499 19.3944
R7777 gnd.n4972 gnd.n4499 19.3944
R7778 gnd.n4973 gnd.n4972 19.3944
R7779 gnd.n4973 gnd.n4497 19.3944
R7780 gnd.n4979 gnd.n4497 19.3944
R7781 gnd.n4982 gnd.n4979 19.3944
R7782 gnd.n4984 gnd.n4982 19.3944
R7783 gnd.n4990 gnd.n4984 19.3944
R7784 gnd.n4990 gnd.n4989 19.3944
R7785 gnd.n4989 gnd.n4372 19.3944
R7786 gnd.n5056 gnd.n4372 19.3944
R7787 gnd.n5057 gnd.n5056 19.3944
R7788 gnd.n5057 gnd.n4365 19.3944
R7789 gnd.n5068 gnd.n4365 19.3944
R7790 gnd.n5069 gnd.n5068 19.3944
R7791 gnd.n5069 gnd.n4348 19.3944
R7792 gnd.n4348 gnd.n4346 19.3944
R7793 gnd.n5093 gnd.n4346 19.3944
R7794 gnd.n5094 gnd.n5093 19.3944
R7795 gnd.n5094 gnd.n4317 19.3944
R7796 gnd.n5141 gnd.n4317 19.3944
R7797 gnd.n5142 gnd.n5141 19.3944
R7798 gnd.n5142 gnd.n4310 19.3944
R7799 gnd.n5153 gnd.n4310 19.3944
R7800 gnd.n5154 gnd.n5153 19.3944
R7801 gnd.n5154 gnd.n4293 19.3944
R7802 gnd.n4293 gnd.n4291 19.3944
R7803 gnd.n5178 gnd.n4291 19.3944
R7804 gnd.n5179 gnd.n5178 19.3944
R7805 gnd.n5179 gnd.n4263 19.3944
R7806 gnd.n5230 gnd.n4263 19.3944
R7807 gnd.n5231 gnd.n5230 19.3944
R7808 gnd.n5231 gnd.n4256 19.3944
R7809 gnd.n5498 gnd.n4256 19.3944
R7810 gnd.n5499 gnd.n5498 19.3944
R7811 gnd.n5499 gnd.n4237 19.3944
R7812 gnd.n5524 gnd.n4237 19.3944
R7813 gnd.n5524 gnd.n4238 19.3944
R7814 gnd.n4855 gnd.n4854 19.3944
R7815 gnd.n4854 gnd.n4587 19.3944
R7816 gnd.n4610 gnd.n4587 19.3944
R7817 gnd.n4613 gnd.n4610 19.3944
R7818 gnd.n4613 gnd.n4606 19.3944
R7819 gnd.n4617 gnd.n4606 19.3944
R7820 gnd.n4620 gnd.n4617 19.3944
R7821 gnd.n4623 gnd.n4620 19.3944
R7822 gnd.n4623 gnd.n4604 19.3944
R7823 gnd.n4627 gnd.n4604 19.3944
R7824 gnd.n4630 gnd.n4627 19.3944
R7825 gnd.n4633 gnd.n4630 19.3944
R7826 gnd.n4633 gnd.n4602 19.3944
R7827 gnd.n4637 gnd.n4602 19.3944
R7828 gnd.n4860 gnd.n4859 19.3944
R7829 gnd.n4859 gnd.n4563 19.3944
R7830 gnd.n4885 gnd.n4563 19.3944
R7831 gnd.n4885 gnd.n4561 19.3944
R7832 gnd.n4891 gnd.n4561 19.3944
R7833 gnd.n4891 gnd.n4890 19.3944
R7834 gnd.n4890 gnd.n4535 19.3944
R7835 gnd.n4915 gnd.n4535 19.3944
R7836 gnd.n4915 gnd.n4533 19.3944
R7837 gnd.n4919 gnd.n4533 19.3944
R7838 gnd.n4919 gnd.n4513 19.3944
R7839 gnd.n4946 gnd.n4513 19.3944
R7840 gnd.n4946 gnd.n4511 19.3944
R7841 gnd.n4956 gnd.n4511 19.3944
R7842 gnd.n4956 gnd.n4955 19.3944
R7843 gnd.n4955 gnd.n4954 19.3944
R7844 gnd.n4954 gnd.n4460 19.3944
R7845 gnd.n5004 gnd.n4460 19.3944
R7846 gnd.n5004 gnd.n5003 19.3944
R7847 gnd.n5003 gnd.n5002 19.3944
R7848 gnd.n5002 gnd.n4464 19.3944
R7849 gnd.n4484 gnd.n4464 19.3944
R7850 gnd.n4484 gnd.n4382 19.3944
R7851 gnd.n5041 gnd.n4382 19.3944
R7852 gnd.n5041 gnd.n4380 19.3944
R7853 gnd.n5047 gnd.n4380 19.3944
R7854 gnd.n5047 gnd.n5046 19.3944
R7855 gnd.n5046 gnd.n4355 19.3944
R7856 gnd.n5081 gnd.n4355 19.3944
R7857 gnd.n5081 gnd.n4353 19.3944
R7858 gnd.n5087 gnd.n4353 19.3944
R7859 gnd.n5087 gnd.n5086 19.3944
R7860 gnd.n5086 gnd.n4328 19.3944
R7861 gnd.n5126 gnd.n4328 19.3944
R7862 gnd.n5126 gnd.n4326 19.3944
R7863 gnd.n5132 gnd.n4326 19.3944
R7864 gnd.n5132 gnd.n5131 19.3944
R7865 gnd.n5131 gnd.n4300 19.3944
R7866 gnd.n5166 gnd.n4300 19.3944
R7867 gnd.n5166 gnd.n4298 19.3944
R7868 gnd.n5172 gnd.n4298 19.3944
R7869 gnd.n5172 gnd.n5171 19.3944
R7870 gnd.n5171 gnd.n4273 19.3944
R7871 gnd.n5215 gnd.n4273 19.3944
R7872 gnd.n5215 gnd.n4271 19.3944
R7873 gnd.n5221 gnd.n4271 19.3944
R7874 gnd.n5221 gnd.n5220 19.3944
R7875 gnd.n5220 gnd.n4246 19.3944
R7876 gnd.n5509 gnd.n4246 19.3944
R7877 gnd.n5509 gnd.n4244 19.3944
R7878 gnd.n5517 gnd.n4244 19.3944
R7879 gnd.n5517 gnd.n5516 19.3944
R7880 gnd.n5516 gnd.n5515 19.3944
R7881 gnd.n5618 gnd.n5617 19.3944
R7882 gnd.n5617 gnd.n4185 19.3944
R7883 gnd.n5613 gnd.n4185 19.3944
R7884 gnd.n5613 gnd.n5610 19.3944
R7885 gnd.n5610 gnd.n5607 19.3944
R7886 gnd.n5607 gnd.n5606 19.3944
R7887 gnd.n5606 gnd.n5603 19.3944
R7888 gnd.n5603 gnd.n5602 19.3944
R7889 gnd.n5602 gnd.n5599 19.3944
R7890 gnd.n5599 gnd.n5598 19.3944
R7891 gnd.n5598 gnd.n5595 19.3944
R7892 gnd.n5595 gnd.n5594 19.3944
R7893 gnd.n5594 gnd.n5591 19.3944
R7894 gnd.n5591 gnd.n5590 19.3944
R7895 gnd.n4775 gnd.n4674 19.3944
R7896 gnd.n4775 gnd.n4665 19.3944
R7897 gnd.n4788 gnd.n4665 19.3944
R7898 gnd.n4788 gnd.n4663 19.3944
R7899 gnd.n4792 gnd.n4663 19.3944
R7900 gnd.n4792 gnd.n4653 19.3944
R7901 gnd.n4804 gnd.n4653 19.3944
R7902 gnd.n4804 gnd.n4651 19.3944
R7903 gnd.n4838 gnd.n4651 19.3944
R7904 gnd.n4838 gnd.n4837 19.3944
R7905 gnd.n4837 gnd.n4836 19.3944
R7906 gnd.n4836 gnd.n4835 19.3944
R7907 gnd.n4835 gnd.n4832 19.3944
R7908 gnd.n4832 gnd.n4831 19.3944
R7909 gnd.n4831 gnd.n4830 19.3944
R7910 gnd.n4830 gnd.n4828 19.3944
R7911 gnd.n4828 gnd.n4827 19.3944
R7912 gnd.n4827 gnd.n4824 19.3944
R7913 gnd.n4824 gnd.n4823 19.3944
R7914 gnd.n4823 gnd.n4822 19.3944
R7915 gnd.n4822 gnd.n4820 19.3944
R7916 gnd.n4820 gnd.n4519 19.3944
R7917 gnd.n4935 gnd.n4519 19.3944
R7918 gnd.n4935 gnd.n4517 19.3944
R7919 gnd.n4941 gnd.n4517 19.3944
R7920 gnd.n4941 gnd.n4940 19.3944
R7921 gnd.n4940 gnd.n4441 19.3944
R7922 gnd.n5015 gnd.n4441 19.3944
R7923 gnd.n5015 gnd.n4442 19.3944
R7924 gnd.n4489 gnd.n4488 19.3944
R7925 gnd.n4492 gnd.n4491 19.3944
R7926 gnd.n4479 gnd.n4478 19.3944
R7927 gnd.n5034 gnd.n4387 19.3944
R7928 gnd.n5034 gnd.n5033 19.3944
R7929 gnd.n5033 gnd.n5032 19.3944
R7930 gnd.n5032 gnd.n5030 19.3944
R7931 gnd.n5030 gnd.n5029 19.3944
R7932 gnd.n5029 gnd.n5027 19.3944
R7933 gnd.n5027 gnd.n5026 19.3944
R7934 gnd.n5026 gnd.n4336 19.3944
R7935 gnd.n5102 gnd.n4336 19.3944
R7936 gnd.n5102 gnd.n4334 19.3944
R7937 gnd.n5121 gnd.n4334 19.3944
R7938 gnd.n5121 gnd.n5120 19.3944
R7939 gnd.n5120 gnd.n5119 19.3944
R7940 gnd.n5119 gnd.n5117 19.3944
R7941 gnd.n5117 gnd.n5116 19.3944
R7942 gnd.n5116 gnd.n5114 19.3944
R7943 gnd.n5114 gnd.n5113 19.3944
R7944 gnd.n5113 gnd.n4280 19.3944
R7945 gnd.n5187 gnd.n4280 19.3944
R7946 gnd.n5187 gnd.n4278 19.3944
R7947 gnd.n5210 gnd.n4278 19.3944
R7948 gnd.n5210 gnd.n5209 19.3944
R7949 gnd.n5209 gnd.n5208 19.3944
R7950 gnd.n5208 gnd.n5205 19.3944
R7951 gnd.n5205 gnd.n5204 19.3944
R7952 gnd.n5204 gnd.n5202 19.3944
R7953 gnd.n5202 gnd.n5201 19.3944
R7954 gnd.n5201 gnd.n5199 19.3944
R7955 gnd.n5199 gnd.n4232 19.3944
R7956 gnd.n4780 gnd.n4670 19.3944
R7957 gnd.n4780 gnd.n4668 19.3944
R7958 gnd.n4784 gnd.n4668 19.3944
R7959 gnd.n4784 gnd.n4659 19.3944
R7960 gnd.n4796 gnd.n4659 19.3944
R7961 gnd.n4796 gnd.n4657 19.3944
R7962 gnd.n4800 gnd.n4657 19.3944
R7963 gnd.n4800 gnd.n4646 19.3944
R7964 gnd.n4842 gnd.n4646 19.3944
R7965 gnd.n4842 gnd.n4600 19.3944
R7966 gnd.n4848 gnd.n4600 19.3944
R7967 gnd.n4848 gnd.n4847 19.3944
R7968 gnd.n4847 gnd.n4578 19.3944
R7969 gnd.n4869 gnd.n4578 19.3944
R7970 gnd.n4869 gnd.n4571 19.3944
R7971 gnd.n4880 gnd.n4571 19.3944
R7972 gnd.n4880 gnd.n4879 19.3944
R7973 gnd.n4879 gnd.n4552 19.3944
R7974 gnd.n4900 gnd.n4552 19.3944
R7975 gnd.n4900 gnd.n4542 19.3944
R7976 gnd.n4910 gnd.n4542 19.3944
R7977 gnd.n4910 gnd.n4525 19.3944
R7978 gnd.n4931 gnd.n4525 19.3944
R7979 gnd.n4931 gnd.n4930 19.3944
R7980 gnd.n4930 gnd.n4504 19.3944
R7981 gnd.n4961 gnd.n4504 19.3944
R7982 gnd.n4961 gnd.n4449 19.3944
R7983 gnd.n5011 gnd.n4449 19.3944
R7984 gnd.n5011 gnd.n5010 19.3944
R7985 gnd.n5010 gnd.n5009 19.3944
R7986 gnd.n5009 gnd.n4453 19.3944
R7987 gnd.n4471 gnd.n4453 19.3944
R7988 gnd.n4997 gnd.n4471 19.3944
R7989 gnd.n4997 gnd.n4996 19.3944
R7990 gnd.n4996 gnd.n4995 19.3944
R7991 gnd.n4995 gnd.n4475 19.3944
R7992 gnd.n4475 gnd.n4374 19.3944
R7993 gnd.n5052 gnd.n4374 19.3944
R7994 gnd.n5052 gnd.n4367 19.3944
R7995 gnd.n5063 gnd.n4367 19.3944
R7996 gnd.n5063 gnd.n4363 19.3944
R7997 gnd.n5076 gnd.n4363 19.3944
R7998 gnd.n5076 gnd.n5075 19.3944
R7999 gnd.n5075 gnd.n4342 19.3944
R8000 gnd.n5098 gnd.n4342 19.3944
R8001 gnd.n5098 gnd.n5097 19.3944
R8002 gnd.n5097 gnd.n4319 19.3944
R8003 gnd.n5137 gnd.n4319 19.3944
R8004 gnd.n5137 gnd.n4312 19.3944
R8005 gnd.n5148 gnd.n4312 19.3944
R8006 gnd.n5148 gnd.n4308 19.3944
R8007 gnd.n5161 gnd.n4308 19.3944
R8008 gnd.n5161 gnd.n5160 19.3944
R8009 gnd.n5160 gnd.n4287 19.3944
R8010 gnd.n5183 gnd.n4287 19.3944
R8011 gnd.n5183 gnd.n5182 19.3944
R8012 gnd.n5182 gnd.n4265 19.3944
R8013 gnd.n5226 gnd.n4265 19.3944
R8014 gnd.n5226 gnd.n4258 19.3944
R8015 gnd.n5237 gnd.n4258 19.3944
R8016 gnd.n5237 gnd.n4254 19.3944
R8017 gnd.n5504 gnd.n4254 19.3944
R8018 gnd.n5504 gnd.n5503 19.3944
R8019 gnd.n5503 gnd.n4235 19.3944
R8020 gnd.n5527 gnd.n4235 19.3944
R8021 gnd.n2612 gnd.n2097 19.3944
R8022 gnd.n2612 gnd.n2611 19.3944
R8023 gnd.n2611 gnd.n2101 19.3944
R8024 gnd.n2604 gnd.n2101 19.3944
R8025 gnd.n2604 gnd.n2603 19.3944
R8026 gnd.n2603 gnd.n2109 19.3944
R8027 gnd.n2596 gnd.n2109 19.3944
R8028 gnd.n2596 gnd.n2595 19.3944
R8029 gnd.n2595 gnd.n2119 19.3944
R8030 gnd.n2588 gnd.n2119 19.3944
R8031 gnd.n2588 gnd.n2587 19.3944
R8032 gnd.n2587 gnd.n2127 19.3944
R8033 gnd.n2580 gnd.n2127 19.3944
R8034 gnd.n2580 gnd.n2579 19.3944
R8035 gnd.n2579 gnd.n2137 19.3944
R8036 gnd.n2572 gnd.n2137 19.3944
R8037 gnd.n2433 gnd.n1130 19.3944
R8038 gnd.n2436 gnd.n2433 19.3944
R8039 gnd.n2437 gnd.n2436 19.3944
R8040 gnd.n2439 gnd.n2437 19.3944
R8041 gnd.n2440 gnd.n2439 19.3944
R8042 gnd.n2443 gnd.n2440 19.3944
R8043 gnd.n2444 gnd.n2443 19.3944
R8044 gnd.n2446 gnd.n2444 19.3944
R8045 gnd.n2447 gnd.n2446 19.3944
R8046 gnd.n2450 gnd.n2447 19.3944
R8047 gnd.n2451 gnd.n2450 19.3944
R8048 gnd.n2453 gnd.n2451 19.3944
R8049 gnd.n2454 gnd.n2453 19.3944
R8050 gnd.n2457 gnd.n2454 19.3944
R8051 gnd.n2458 gnd.n2457 19.3944
R8052 gnd.n2460 gnd.n2458 19.3944
R8053 gnd.n2461 gnd.n2460 19.3944
R8054 gnd.n2464 gnd.n2461 19.3944
R8055 gnd.n2465 gnd.n2464 19.3944
R8056 gnd.n2467 gnd.n2465 19.3944
R8057 gnd.n2468 gnd.n2467 19.3944
R8058 gnd.n2471 gnd.n2468 19.3944
R8059 gnd.n2472 gnd.n2471 19.3944
R8060 gnd.n2474 gnd.n2472 19.3944
R8061 gnd.n2475 gnd.n2474 19.3944
R8062 gnd.n2478 gnd.n2475 19.3944
R8063 gnd.n2479 gnd.n2478 19.3944
R8064 gnd.n2481 gnd.n2479 19.3944
R8065 gnd.n2482 gnd.n2481 19.3944
R8066 gnd.n2485 gnd.n2482 19.3944
R8067 gnd.n2486 gnd.n2485 19.3944
R8068 gnd.n2488 gnd.n2486 19.3944
R8069 gnd.n2489 gnd.n2488 19.3944
R8070 gnd.n2492 gnd.n2489 19.3944
R8071 gnd.n2493 gnd.n2492 19.3944
R8072 gnd.n2494 gnd.n2493 19.3944
R8073 gnd.n2494 gnd.n2284 19.3944
R8074 gnd.n2507 gnd.n2284 19.3944
R8075 gnd.n2508 gnd.n2507 19.3944
R8076 gnd.n2512 gnd.n2508 19.3944
R8077 gnd.n2512 gnd.n2511 19.3944
R8078 gnd.n2511 gnd.n2510 19.3944
R8079 gnd.n2324 gnd.n2323 19.3944
R8080 gnd.n2327 gnd.n2324 19.3944
R8081 gnd.n2327 gnd.n2321 19.3944
R8082 gnd.n2333 gnd.n2321 19.3944
R8083 gnd.n2334 gnd.n2333 19.3944
R8084 gnd.n2337 gnd.n2334 19.3944
R8085 gnd.n2337 gnd.n2319 19.3944
R8086 gnd.n2343 gnd.n2319 19.3944
R8087 gnd.n2344 gnd.n2343 19.3944
R8088 gnd.n2347 gnd.n2344 19.3944
R8089 gnd.n2347 gnd.n2317 19.3944
R8090 gnd.n2353 gnd.n2317 19.3944
R8091 gnd.n2354 gnd.n2353 19.3944
R8092 gnd.n2357 gnd.n2354 19.3944
R8093 gnd.n2357 gnd.n2313 19.3944
R8094 gnd.n2361 gnd.n2313 19.3944
R8095 gnd.n2366 gnd.n2308 19.3944
R8096 gnd.n2371 gnd.n2308 19.3944
R8097 gnd.n2372 gnd.n2371 19.3944
R8098 gnd.n2374 gnd.n2372 19.3944
R8099 gnd.n2374 gnd.n2306 19.3944
R8100 gnd.n2379 gnd.n2306 19.3944
R8101 gnd.n2380 gnd.n2379 19.3944
R8102 gnd.n2382 gnd.n2380 19.3944
R8103 gnd.n2382 gnd.n2304 19.3944
R8104 gnd.n2387 gnd.n2304 19.3944
R8105 gnd.n2388 gnd.n2387 19.3944
R8106 gnd.n2390 gnd.n2388 19.3944
R8107 gnd.n2390 gnd.n2302 19.3944
R8108 gnd.n2395 gnd.n2302 19.3944
R8109 gnd.n2396 gnd.n2395 19.3944
R8110 gnd.n2398 gnd.n2396 19.3944
R8111 gnd.n2398 gnd.n2300 19.3944
R8112 gnd.n2403 gnd.n2300 19.3944
R8113 gnd.n2404 gnd.n2403 19.3944
R8114 gnd.n2406 gnd.n2404 19.3944
R8115 gnd.n2406 gnd.n2297 19.3944
R8116 gnd.n2410 gnd.n2297 19.3944
R8117 gnd.n2411 gnd.n2410 19.3944
R8118 gnd.n2413 gnd.n2411 19.3944
R8119 gnd.n2413 gnd.n2294 19.3944
R8120 gnd.n2417 gnd.n2294 19.3944
R8121 gnd.n2418 gnd.n2417 19.3944
R8122 gnd.n2420 gnd.n2418 19.3944
R8123 gnd.n2420 gnd.n2291 19.3944
R8124 gnd.n2424 gnd.n2291 19.3944
R8125 gnd.n2425 gnd.n2424 19.3944
R8126 gnd.n2427 gnd.n2425 19.3944
R8127 gnd.n2427 gnd.n2288 19.3944
R8128 gnd.n2431 gnd.n2288 19.3944
R8129 gnd.n2432 gnd.n2431 19.3944
R8130 gnd.n2498 gnd.n2432 19.3944
R8131 gnd.n2498 gnd.n2286 19.3944
R8132 gnd.n2503 gnd.n2286 19.3944
R8133 gnd.n2503 gnd.n2283 19.3944
R8134 gnd.n2537 gnd.n2283 19.3944
R8135 gnd.n2538 gnd.n2537 19.3944
R8136 gnd.n2538 gnd.n2151 19.3944
R8137 gnd.n4170 gnd.n4169 19.3944
R8138 gnd.n4169 gnd.n4168 19.3944
R8139 gnd.n4168 gnd.n4167 19.3944
R8140 gnd.n4167 gnd.n4165 19.3944
R8141 gnd.n4165 gnd.n4162 19.3944
R8142 gnd.n4162 gnd.n4161 19.3944
R8143 gnd.n4161 gnd.n4158 19.3944
R8144 gnd.n4158 gnd.n4157 19.3944
R8145 gnd.n4157 gnd.n4154 19.3944
R8146 gnd.n4154 gnd.n4153 19.3944
R8147 gnd.n4153 gnd.n4150 19.3944
R8148 gnd.n4150 gnd.n4149 19.3944
R8149 gnd.n4149 gnd.n4146 19.3944
R8150 gnd.n4146 gnd.n4145 19.3944
R8151 gnd.n4145 gnd.n4142 19.3944
R8152 gnd.n4142 gnd.n4141 19.3944
R8153 gnd.n4141 gnd.n4138 19.3944
R8154 gnd.n4136 gnd.n4133 19.3944
R8155 gnd.n4133 gnd.n4132 19.3944
R8156 gnd.n4132 gnd.n4129 19.3944
R8157 gnd.n4129 gnd.n4128 19.3944
R8158 gnd.n4128 gnd.n4125 19.3944
R8159 gnd.n4125 gnd.n4124 19.3944
R8160 gnd.n4124 gnd.n4121 19.3944
R8161 gnd.n4121 gnd.n4120 19.3944
R8162 gnd.n4120 gnd.n4117 19.3944
R8163 gnd.n4117 gnd.n4116 19.3944
R8164 gnd.n4116 gnd.n4113 19.3944
R8165 gnd.n4113 gnd.n4112 19.3944
R8166 gnd.n4112 gnd.n4109 19.3944
R8167 gnd.n4109 gnd.n4108 19.3944
R8168 gnd.n4108 gnd.n4105 19.3944
R8169 gnd.n4105 gnd.n4104 19.3944
R8170 gnd.n4104 gnd.n4101 19.3944
R8171 gnd.n4101 gnd.n4100 19.3944
R8172 gnd.n4096 gnd.n4093 19.3944
R8173 gnd.n4093 gnd.n4092 19.3944
R8174 gnd.n4092 gnd.n4089 19.3944
R8175 gnd.n4089 gnd.n4088 19.3944
R8176 gnd.n4088 gnd.n4085 19.3944
R8177 gnd.n4085 gnd.n4084 19.3944
R8178 gnd.n4084 gnd.n4081 19.3944
R8179 gnd.n4081 gnd.n4080 19.3944
R8180 gnd.n4080 gnd.n4077 19.3944
R8181 gnd.n4077 gnd.n4076 19.3944
R8182 gnd.n4076 gnd.n4073 19.3944
R8183 gnd.n4073 gnd.n4072 19.3944
R8184 gnd.n4072 gnd.n4069 19.3944
R8185 gnd.n4069 gnd.n4068 19.3944
R8186 gnd.n4068 gnd.n4065 19.3944
R8187 gnd.n4065 gnd.n4064 19.3944
R8188 gnd.n4064 gnd.n4061 19.3944
R8189 gnd.n4061 gnd.n4060 19.3944
R8190 gnd.n3921 gnd.n1337 19.3944
R8191 gnd.n3916 gnd.n1337 19.3944
R8192 gnd.n3916 gnd.n3915 19.3944
R8193 gnd.n3915 gnd.n3914 19.3944
R8194 gnd.n3914 gnd.n3911 19.3944
R8195 gnd.n3911 gnd.n3910 19.3944
R8196 gnd.n3910 gnd.n3907 19.3944
R8197 gnd.n3907 gnd.n3906 19.3944
R8198 gnd.n3906 gnd.n3903 19.3944
R8199 gnd.n3903 gnd.n3902 19.3944
R8200 gnd.n3902 gnd.n3899 19.3944
R8201 gnd.n3899 gnd.n3898 19.3944
R8202 gnd.n3898 gnd.n3895 19.3944
R8203 gnd.n3895 gnd.n3894 19.3944
R8204 gnd.n3894 gnd.n3891 19.3944
R8205 gnd.n3891 gnd.n3890 19.3944
R8206 gnd.n3890 gnd.n3887 19.3944
R8207 gnd.n2199 gnd.n2196 19.3944
R8208 gnd.n2202 gnd.n2199 19.3944
R8209 gnd.n2202 gnd.n2162 19.3944
R8210 gnd.n2206 gnd.n2162 19.3944
R8211 gnd.n2209 gnd.n2206 19.3944
R8212 gnd.n2212 gnd.n2209 19.3944
R8213 gnd.n2212 gnd.n2160 19.3944
R8214 gnd.n2216 gnd.n2160 19.3944
R8215 gnd.n2219 gnd.n2216 19.3944
R8216 gnd.n2222 gnd.n2219 19.3944
R8217 gnd.n2222 gnd.n2158 19.3944
R8218 gnd.n2226 gnd.n2158 19.3944
R8219 gnd.n2229 gnd.n2226 19.3944
R8220 gnd.n2232 gnd.n2229 19.3944
R8221 gnd.n2232 gnd.n2156 19.3944
R8222 gnd.n2236 gnd.n2156 19.3944
R8223 gnd.n2239 gnd.n2236 19.3944
R8224 gnd.n2242 gnd.n2239 19.3944
R8225 gnd.n2172 gnd.n1406 19.3944
R8226 gnd.n2176 gnd.n2172 19.3944
R8227 gnd.n2179 gnd.n2176 19.3944
R8228 gnd.n2182 gnd.n2179 19.3944
R8229 gnd.n2182 gnd.n2168 19.3944
R8230 gnd.n2186 gnd.n2168 19.3944
R8231 gnd.n2189 gnd.n2186 19.3944
R8232 gnd.n2192 gnd.n2189 19.3944
R8233 gnd.n3885 gnd.n3882 19.3944
R8234 gnd.n3882 gnd.n3881 19.3944
R8235 gnd.n3881 gnd.n3878 19.3944
R8236 gnd.n3878 gnd.n3877 19.3944
R8237 gnd.n3877 gnd.n3874 19.3944
R8238 gnd.n3874 gnd.n3873 19.3944
R8239 gnd.n3873 gnd.n3870 19.3944
R8240 gnd.n4047 gnd.n1140 19.3944
R8241 gnd.n4047 gnd.n1141 19.3944
R8242 gnd.n4043 gnd.n1141 19.3944
R8243 gnd.n4043 gnd.n1144 19.3944
R8244 gnd.n4033 gnd.n1144 19.3944
R8245 gnd.n4033 gnd.n4032 19.3944
R8246 gnd.n4032 gnd.n4031 19.3944
R8247 gnd.n4031 gnd.n1164 19.3944
R8248 gnd.n4021 gnd.n1164 19.3944
R8249 gnd.n4021 gnd.n4020 19.3944
R8250 gnd.n4020 gnd.n4019 19.3944
R8251 gnd.n4019 gnd.n1182 19.3944
R8252 gnd.n4009 gnd.n1182 19.3944
R8253 gnd.n4009 gnd.n4008 19.3944
R8254 gnd.n4008 gnd.n4007 19.3944
R8255 gnd.n4007 gnd.n1202 19.3944
R8256 gnd.n3997 gnd.n1202 19.3944
R8257 gnd.n3997 gnd.n3996 19.3944
R8258 gnd.n3996 gnd.n3995 19.3944
R8259 gnd.n3995 gnd.n1220 19.3944
R8260 gnd.n3985 gnd.n1220 19.3944
R8261 gnd.n3985 gnd.n3984 19.3944
R8262 gnd.n3984 gnd.n3983 19.3944
R8263 gnd.n3983 gnd.n1240 19.3944
R8264 gnd.n3973 gnd.n1240 19.3944
R8265 gnd.n3973 gnd.n3972 19.3944
R8266 gnd.n3972 gnd.n3971 19.3944
R8267 gnd.n3971 gnd.n1259 19.3944
R8268 gnd.n3961 gnd.n1259 19.3944
R8269 gnd.n3961 gnd.n3960 19.3944
R8270 gnd.n3960 gnd.n3959 19.3944
R8271 gnd.n3959 gnd.n1278 19.3944
R8272 gnd.n3949 gnd.n1278 19.3944
R8273 gnd.n3949 gnd.n3948 19.3944
R8274 gnd.n3948 gnd.n3947 19.3944
R8275 gnd.n3947 gnd.n1297 19.3944
R8276 gnd.n3937 gnd.n1297 19.3944
R8277 gnd.n3937 gnd.n3936 19.3944
R8278 gnd.n3936 gnd.n3935 19.3944
R8279 gnd.n3935 gnd.n1318 19.3944
R8280 gnd.n3925 gnd.n1318 19.3944
R8281 gnd.n3925 gnd.n3924 19.3944
R8282 gnd.n4052 gnd.n1132 19.3944
R8283 gnd.n1151 gnd.n1132 19.3944
R8284 gnd.n4039 gnd.n1151 19.3944
R8285 gnd.n4039 gnd.n4038 19.3944
R8286 gnd.n4038 gnd.n4037 19.3944
R8287 gnd.n4037 gnd.n1155 19.3944
R8288 gnd.n4027 gnd.n1155 19.3944
R8289 gnd.n4027 gnd.n4026 19.3944
R8290 gnd.n4026 gnd.n4025 19.3944
R8291 gnd.n4025 gnd.n1173 19.3944
R8292 gnd.n4015 gnd.n1173 19.3944
R8293 gnd.n4015 gnd.n4014 19.3944
R8294 gnd.n4014 gnd.n4013 19.3944
R8295 gnd.n4013 gnd.n1191 19.3944
R8296 gnd.n4003 gnd.n1191 19.3944
R8297 gnd.n4003 gnd.n4002 19.3944
R8298 gnd.n4002 gnd.n4001 19.3944
R8299 gnd.n4001 gnd.n1211 19.3944
R8300 gnd.n3991 gnd.n1211 19.3944
R8301 gnd.n3991 gnd.n3990 19.3944
R8302 gnd.n3990 gnd.n3989 19.3944
R8303 gnd.n3989 gnd.n1229 19.3944
R8304 gnd.n3979 gnd.n1229 19.3944
R8305 gnd.n3979 gnd.n3978 19.3944
R8306 gnd.n3978 gnd.n3977 19.3944
R8307 gnd.n3977 gnd.n1249 19.3944
R8308 gnd.n3967 gnd.n1249 19.3944
R8309 gnd.n3967 gnd.n3966 19.3944
R8310 gnd.n3966 gnd.n3965 19.3944
R8311 gnd.n3965 gnd.n1267 19.3944
R8312 gnd.n3955 gnd.n1267 19.3944
R8313 gnd.n3955 gnd.n3954 19.3944
R8314 gnd.n3954 gnd.n3953 19.3944
R8315 gnd.n3953 gnd.n1287 19.3944
R8316 gnd.n3943 gnd.n1287 19.3944
R8317 gnd.n3943 gnd.n3942 19.3944
R8318 gnd.n3942 gnd.n3941 19.3944
R8319 gnd.n3941 gnd.n1307 19.3944
R8320 gnd.n3931 gnd.n1307 19.3944
R8321 gnd.n3931 gnd.n3930 19.3944
R8322 gnd.n3930 gnd.n3929 19.3944
R8323 gnd.n3929 gnd.n1328 19.3944
R8324 gnd.n2523 gnd.n2519 19.3944
R8325 gnd.n2523 gnd.n2517 19.3944
R8326 gnd.n2527 gnd.n2517 19.3944
R8327 gnd.n2527 gnd.n2515 19.3944
R8328 gnd.n2532 gnd.n2515 19.3944
R8329 gnd.n2532 gnd.n2251 19.3944
R8330 gnd.n2564 gnd.n2251 19.3944
R8331 gnd.n2564 gnd.n2563 19.3944
R8332 gnd.n2563 gnd.n2562 19.3944
R8333 gnd.n2562 gnd.n2255 19.3944
R8334 gnd.n2547 gnd.n2255 19.3944
R8335 gnd.n2553 gnd.n2547 19.3944
R8336 gnd.n2553 gnd.n2552 19.3944
R8337 gnd.n2552 gnd.n2069 19.3944
R8338 gnd.n2647 gnd.n2069 19.3944
R8339 gnd.n2647 gnd.n2067 19.3944
R8340 gnd.n2653 gnd.n2067 19.3944
R8341 gnd.n2653 gnd.n2652 19.3944
R8342 gnd.n2652 gnd.n2044 19.3944
R8343 gnd.n2677 gnd.n2044 19.3944
R8344 gnd.n2677 gnd.n2042 19.3944
R8345 gnd.n2683 gnd.n2042 19.3944
R8346 gnd.n2683 gnd.n2682 19.3944
R8347 gnd.n2682 gnd.n2019 19.3944
R8348 gnd.n2707 gnd.n2019 19.3944
R8349 gnd.n2707 gnd.n2017 19.3944
R8350 gnd.n2713 gnd.n2017 19.3944
R8351 gnd.n2713 gnd.n2712 19.3944
R8352 gnd.n2712 gnd.n1994 19.3944
R8353 gnd.n2741 gnd.n1994 19.3944
R8354 gnd.n2741 gnd.n1992 19.3944
R8355 gnd.n2760 gnd.n1992 19.3944
R8356 gnd.n2760 gnd.n2759 19.3944
R8357 gnd.n2759 gnd.n2758 19.3944
R8358 gnd.n2758 gnd.n2747 19.3944
R8359 gnd.n2753 gnd.n2747 19.3944
R8360 gnd.n2753 gnd.n2752 19.3944
R8361 gnd.n2752 gnd.n1963 19.3944
R8362 gnd.n2915 gnd.n1963 19.3944
R8363 gnd.n2915 gnd.n1961 19.3944
R8364 gnd.n2921 gnd.n1961 19.3944
R8365 gnd.n2921 gnd.n2920 19.3944
R8366 gnd.n2920 gnd.n1936 19.3944
R8367 gnd.n2952 gnd.n1936 19.3944
R8368 gnd.n2952 gnd.n1934 19.3944
R8369 gnd.n2956 gnd.n1934 19.3944
R8370 gnd.n2956 gnd.n1915 19.3944
R8371 gnd.n2982 gnd.n1915 19.3944
R8372 gnd.n2982 gnd.n1913 19.3944
R8373 gnd.n2988 gnd.n1913 19.3944
R8374 gnd.n2988 gnd.n2987 19.3944
R8375 gnd.n2987 gnd.n1885 19.3944
R8376 gnd.n3033 gnd.n1885 19.3944
R8377 gnd.n3033 gnd.n1883 19.3944
R8378 gnd.n3039 gnd.n1883 19.3944
R8379 gnd.n3039 gnd.n3038 19.3944
R8380 gnd.n3038 gnd.n1866 19.3944
R8381 gnd.n3061 gnd.n1866 19.3944
R8382 gnd.n3061 gnd.n1864 19.3944
R8383 gnd.n3065 gnd.n1864 19.3944
R8384 gnd.n3065 gnd.n1838 19.3944
R8385 gnd.n3117 gnd.n1838 19.3944
R8386 gnd.n3117 gnd.n1836 19.3944
R8387 gnd.n3121 gnd.n1836 19.3944
R8388 gnd.n3121 gnd.n1815 19.3944
R8389 gnd.n3157 gnd.n1815 19.3944
R8390 gnd.n3157 gnd.n1813 19.3944
R8391 gnd.n3161 gnd.n1813 19.3944
R8392 gnd.n3161 gnd.n1792 19.3944
R8393 gnd.n3197 gnd.n1792 19.3944
R8394 gnd.n3197 gnd.n1790 19.3944
R8395 gnd.n3201 gnd.n1790 19.3944
R8396 gnd.n3201 gnd.n1770 19.3944
R8397 gnd.n3244 gnd.n1770 19.3944
R8398 gnd.n3244 gnd.n1768 19.3944
R8399 gnd.n3248 gnd.n1768 19.3944
R8400 gnd.n3248 gnd.n1752 19.3944
R8401 gnd.n3271 gnd.n1752 19.3944
R8402 gnd.n3271 gnd.n1750 19.3944
R8403 gnd.n3280 gnd.n1750 19.3944
R8404 gnd.n3280 gnd.n3279 19.3944
R8405 gnd.n3279 gnd.n3278 19.3944
R8406 gnd.n3278 gnd.n1716 19.3944
R8407 gnd.n3338 gnd.n1716 19.3944
R8408 gnd.n3338 gnd.n1714 19.3944
R8409 gnd.n3344 gnd.n1714 19.3944
R8410 gnd.n3344 gnd.n3343 19.3944
R8411 gnd.n3343 gnd.n1689 19.3944
R8412 gnd.n3389 gnd.n1689 19.3944
R8413 gnd.n3389 gnd.n1687 19.3944
R8414 gnd.n3398 gnd.n1687 19.3944
R8415 gnd.n3398 gnd.n3397 19.3944
R8416 gnd.n3397 gnd.n3396 19.3944
R8417 gnd.n3396 gnd.n1628 19.3944
R8418 gnd.n3577 gnd.n1628 19.3944
R8419 gnd.n3577 gnd.n1626 19.3944
R8420 gnd.n3581 gnd.n1626 19.3944
R8421 gnd.n3581 gnd.n1617 19.3944
R8422 gnd.n3599 gnd.n1617 19.3944
R8423 gnd.n3599 gnd.n1615 19.3944
R8424 gnd.n3603 gnd.n1615 19.3944
R8425 gnd.n3603 gnd.n1605 19.3944
R8426 gnd.n3620 gnd.n1605 19.3944
R8427 gnd.n3620 gnd.n1603 19.3944
R8428 gnd.n3624 gnd.n1603 19.3944
R8429 gnd.n3624 gnd.n1593 19.3944
R8430 gnd.n3641 gnd.n1593 19.3944
R8431 gnd.n3641 gnd.n1591 19.3944
R8432 gnd.n3645 gnd.n1591 19.3944
R8433 gnd.n3645 gnd.n1580 19.3944
R8434 gnd.n3662 gnd.n1580 19.3944
R8435 gnd.n3662 gnd.n1578 19.3944
R8436 gnd.n3672 gnd.n1578 19.3944
R8437 gnd.n3672 gnd.n3671 19.3944
R8438 gnd.n3671 gnd.n3670 19.3944
R8439 gnd.n3670 gnd.n493 19.3944
R8440 gnd.n6352 gnd.n493 19.3944
R8441 gnd.n6352 gnd.n6351 19.3944
R8442 gnd.n6351 gnd.n6350 19.3944
R8443 gnd.n6350 gnd.n497 19.3944
R8444 gnd.n499 gnd.n497 19.3944
R8445 gnd.n508 gnd.n499 19.3944
R8446 gnd.n6336 gnd.n508 19.3944
R8447 gnd.n6336 gnd.n6335 19.3944
R8448 gnd.n6335 gnd.n6334 19.3944
R8449 gnd.n6334 gnd.n515 19.3944
R8450 gnd.n6330 gnd.n515 19.3944
R8451 gnd.n6330 gnd.n6329 19.3944
R8452 gnd.n6116 gnd.n645 19.3944
R8453 gnd.n6116 gnd.n641 19.3944
R8454 gnd.n6122 gnd.n641 19.3944
R8455 gnd.n6122 gnd.n639 19.3944
R8456 gnd.n6126 gnd.n639 19.3944
R8457 gnd.n6126 gnd.n635 19.3944
R8458 gnd.n6132 gnd.n635 19.3944
R8459 gnd.n6132 gnd.n633 19.3944
R8460 gnd.n6136 gnd.n633 19.3944
R8461 gnd.n6136 gnd.n629 19.3944
R8462 gnd.n6142 gnd.n629 19.3944
R8463 gnd.n6142 gnd.n627 19.3944
R8464 gnd.n6146 gnd.n627 19.3944
R8465 gnd.n6146 gnd.n623 19.3944
R8466 gnd.n6152 gnd.n623 19.3944
R8467 gnd.n6152 gnd.n621 19.3944
R8468 gnd.n6156 gnd.n621 19.3944
R8469 gnd.n6156 gnd.n617 19.3944
R8470 gnd.n6162 gnd.n617 19.3944
R8471 gnd.n6162 gnd.n615 19.3944
R8472 gnd.n6166 gnd.n615 19.3944
R8473 gnd.n6166 gnd.n611 19.3944
R8474 gnd.n6172 gnd.n611 19.3944
R8475 gnd.n6172 gnd.n609 19.3944
R8476 gnd.n6176 gnd.n609 19.3944
R8477 gnd.n6176 gnd.n605 19.3944
R8478 gnd.n6182 gnd.n605 19.3944
R8479 gnd.n6182 gnd.n603 19.3944
R8480 gnd.n6186 gnd.n603 19.3944
R8481 gnd.n6186 gnd.n599 19.3944
R8482 gnd.n6192 gnd.n599 19.3944
R8483 gnd.n6192 gnd.n597 19.3944
R8484 gnd.n6196 gnd.n597 19.3944
R8485 gnd.n6196 gnd.n593 19.3944
R8486 gnd.n6202 gnd.n593 19.3944
R8487 gnd.n6202 gnd.n591 19.3944
R8488 gnd.n6206 gnd.n591 19.3944
R8489 gnd.n6206 gnd.n587 19.3944
R8490 gnd.n6212 gnd.n587 19.3944
R8491 gnd.n6212 gnd.n585 19.3944
R8492 gnd.n6216 gnd.n585 19.3944
R8493 gnd.n6216 gnd.n581 19.3944
R8494 gnd.n6222 gnd.n581 19.3944
R8495 gnd.n6222 gnd.n579 19.3944
R8496 gnd.n6226 gnd.n579 19.3944
R8497 gnd.n6226 gnd.n575 19.3944
R8498 gnd.n6232 gnd.n575 19.3944
R8499 gnd.n6232 gnd.n573 19.3944
R8500 gnd.n6236 gnd.n573 19.3944
R8501 gnd.n6236 gnd.n569 19.3944
R8502 gnd.n6242 gnd.n569 19.3944
R8503 gnd.n6242 gnd.n567 19.3944
R8504 gnd.n6246 gnd.n567 19.3944
R8505 gnd.n6246 gnd.n563 19.3944
R8506 gnd.n6252 gnd.n563 19.3944
R8507 gnd.n6252 gnd.n561 19.3944
R8508 gnd.n6256 gnd.n561 19.3944
R8509 gnd.n6256 gnd.n557 19.3944
R8510 gnd.n6262 gnd.n557 19.3944
R8511 gnd.n6262 gnd.n555 19.3944
R8512 gnd.n6266 gnd.n555 19.3944
R8513 gnd.n6266 gnd.n551 19.3944
R8514 gnd.n6272 gnd.n551 19.3944
R8515 gnd.n6272 gnd.n549 19.3944
R8516 gnd.n6276 gnd.n549 19.3944
R8517 gnd.n6276 gnd.n545 19.3944
R8518 gnd.n6282 gnd.n545 19.3944
R8519 gnd.n6282 gnd.n543 19.3944
R8520 gnd.n6286 gnd.n543 19.3944
R8521 gnd.n6286 gnd.n539 19.3944
R8522 gnd.n6292 gnd.n539 19.3944
R8523 gnd.n6292 gnd.n537 19.3944
R8524 gnd.n6296 gnd.n537 19.3944
R8525 gnd.n6296 gnd.n533 19.3944
R8526 gnd.n6302 gnd.n533 19.3944
R8527 gnd.n6302 gnd.n531 19.3944
R8528 gnd.n6306 gnd.n531 19.3944
R8529 gnd.n6306 gnd.n527 19.3944
R8530 gnd.n6312 gnd.n527 19.3944
R8531 gnd.n6312 gnd.n525 19.3944
R8532 gnd.n6318 gnd.n525 19.3944
R8533 gnd.n6318 gnd.n6317 19.3944
R8534 gnd.n6317 gnd.n521 19.3944
R8535 gnd.n6326 gnd.n521 19.3944
R8536 gnd.n5792 gnd.n837 19.3944
R8537 gnd.n5796 gnd.n837 19.3944
R8538 gnd.n5796 gnd.n833 19.3944
R8539 gnd.n5802 gnd.n833 19.3944
R8540 gnd.n5802 gnd.n831 19.3944
R8541 gnd.n5806 gnd.n831 19.3944
R8542 gnd.n5806 gnd.n827 19.3944
R8543 gnd.n5812 gnd.n827 19.3944
R8544 gnd.n5812 gnd.n825 19.3944
R8545 gnd.n5816 gnd.n825 19.3944
R8546 gnd.n5816 gnd.n821 19.3944
R8547 gnd.n5822 gnd.n821 19.3944
R8548 gnd.n5822 gnd.n819 19.3944
R8549 gnd.n5826 gnd.n819 19.3944
R8550 gnd.n5826 gnd.n815 19.3944
R8551 gnd.n5832 gnd.n815 19.3944
R8552 gnd.n5832 gnd.n813 19.3944
R8553 gnd.n5836 gnd.n813 19.3944
R8554 gnd.n5836 gnd.n809 19.3944
R8555 gnd.n5842 gnd.n809 19.3944
R8556 gnd.n5842 gnd.n807 19.3944
R8557 gnd.n5846 gnd.n807 19.3944
R8558 gnd.n5846 gnd.n803 19.3944
R8559 gnd.n5852 gnd.n803 19.3944
R8560 gnd.n5852 gnd.n801 19.3944
R8561 gnd.n5856 gnd.n801 19.3944
R8562 gnd.n5856 gnd.n797 19.3944
R8563 gnd.n5862 gnd.n797 19.3944
R8564 gnd.n5862 gnd.n795 19.3944
R8565 gnd.n5866 gnd.n795 19.3944
R8566 gnd.n5866 gnd.n791 19.3944
R8567 gnd.n5872 gnd.n791 19.3944
R8568 gnd.n5872 gnd.n789 19.3944
R8569 gnd.n5876 gnd.n789 19.3944
R8570 gnd.n5876 gnd.n785 19.3944
R8571 gnd.n5882 gnd.n785 19.3944
R8572 gnd.n5882 gnd.n783 19.3944
R8573 gnd.n5886 gnd.n783 19.3944
R8574 gnd.n5886 gnd.n779 19.3944
R8575 gnd.n5892 gnd.n779 19.3944
R8576 gnd.n5892 gnd.n777 19.3944
R8577 gnd.n5896 gnd.n777 19.3944
R8578 gnd.n5896 gnd.n773 19.3944
R8579 gnd.n5902 gnd.n773 19.3944
R8580 gnd.n5902 gnd.n771 19.3944
R8581 gnd.n5906 gnd.n771 19.3944
R8582 gnd.n5906 gnd.n767 19.3944
R8583 gnd.n5912 gnd.n767 19.3944
R8584 gnd.n5912 gnd.n765 19.3944
R8585 gnd.n5916 gnd.n765 19.3944
R8586 gnd.n5916 gnd.n761 19.3944
R8587 gnd.n5922 gnd.n761 19.3944
R8588 gnd.n5922 gnd.n759 19.3944
R8589 gnd.n5926 gnd.n759 19.3944
R8590 gnd.n5926 gnd.n755 19.3944
R8591 gnd.n5932 gnd.n755 19.3944
R8592 gnd.n5932 gnd.n753 19.3944
R8593 gnd.n5936 gnd.n753 19.3944
R8594 gnd.n5936 gnd.n749 19.3944
R8595 gnd.n5942 gnd.n749 19.3944
R8596 gnd.n5942 gnd.n747 19.3944
R8597 gnd.n5946 gnd.n747 19.3944
R8598 gnd.n5946 gnd.n743 19.3944
R8599 gnd.n5952 gnd.n743 19.3944
R8600 gnd.n5952 gnd.n741 19.3944
R8601 gnd.n5956 gnd.n741 19.3944
R8602 gnd.n5956 gnd.n737 19.3944
R8603 gnd.n5962 gnd.n737 19.3944
R8604 gnd.n5962 gnd.n735 19.3944
R8605 gnd.n5966 gnd.n735 19.3944
R8606 gnd.n5966 gnd.n731 19.3944
R8607 gnd.n5972 gnd.n731 19.3944
R8608 gnd.n5972 gnd.n729 19.3944
R8609 gnd.n5976 gnd.n729 19.3944
R8610 gnd.n5976 gnd.n725 19.3944
R8611 gnd.n5982 gnd.n725 19.3944
R8612 gnd.n5982 gnd.n723 19.3944
R8613 gnd.n5986 gnd.n723 19.3944
R8614 gnd.n5986 gnd.n719 19.3944
R8615 gnd.n5992 gnd.n719 19.3944
R8616 gnd.n5992 gnd.n717 19.3944
R8617 gnd.n5996 gnd.n717 19.3944
R8618 gnd.n5996 gnd.n713 19.3944
R8619 gnd.n6002 gnd.n713 19.3944
R8620 gnd.n6002 gnd.n711 19.3944
R8621 gnd.n6006 gnd.n711 19.3944
R8622 gnd.n6006 gnd.n707 19.3944
R8623 gnd.n6012 gnd.n707 19.3944
R8624 gnd.n6012 gnd.n705 19.3944
R8625 gnd.n6016 gnd.n705 19.3944
R8626 gnd.n6016 gnd.n701 19.3944
R8627 gnd.n6022 gnd.n701 19.3944
R8628 gnd.n6022 gnd.n699 19.3944
R8629 gnd.n6026 gnd.n699 19.3944
R8630 gnd.n6026 gnd.n695 19.3944
R8631 gnd.n6032 gnd.n695 19.3944
R8632 gnd.n6032 gnd.n693 19.3944
R8633 gnd.n6036 gnd.n693 19.3944
R8634 gnd.n6036 gnd.n689 19.3944
R8635 gnd.n6042 gnd.n689 19.3944
R8636 gnd.n6042 gnd.n687 19.3944
R8637 gnd.n6046 gnd.n687 19.3944
R8638 gnd.n6046 gnd.n683 19.3944
R8639 gnd.n6052 gnd.n683 19.3944
R8640 gnd.n6052 gnd.n681 19.3944
R8641 gnd.n6056 gnd.n681 19.3944
R8642 gnd.n6056 gnd.n677 19.3944
R8643 gnd.n6062 gnd.n677 19.3944
R8644 gnd.n6062 gnd.n675 19.3944
R8645 gnd.n6066 gnd.n675 19.3944
R8646 gnd.n6066 gnd.n671 19.3944
R8647 gnd.n6072 gnd.n671 19.3944
R8648 gnd.n6072 gnd.n669 19.3944
R8649 gnd.n6076 gnd.n669 19.3944
R8650 gnd.n6076 gnd.n665 19.3944
R8651 gnd.n6082 gnd.n665 19.3944
R8652 gnd.n6082 gnd.n663 19.3944
R8653 gnd.n6086 gnd.n663 19.3944
R8654 gnd.n6086 gnd.n659 19.3944
R8655 gnd.n6092 gnd.n659 19.3944
R8656 gnd.n6092 gnd.n657 19.3944
R8657 gnd.n6096 gnd.n657 19.3944
R8658 gnd.n6096 gnd.n653 19.3944
R8659 gnd.n6102 gnd.n653 19.3944
R8660 gnd.n6102 gnd.n651 19.3944
R8661 gnd.n6106 gnd.n651 19.3944
R8662 gnd.n6106 gnd.n647 19.3944
R8663 gnd.n6112 gnd.n647 19.3944
R8664 gnd.n5786 gnd.n842 19.3944
R8665 gnd.n5786 gnd.n5785 19.3944
R8666 gnd.n5785 gnd.n5784 19.3944
R8667 gnd.n5784 gnd.n846 19.3944
R8668 gnd.n5778 gnd.n846 19.3944
R8669 gnd.n5778 gnd.n5777 19.3944
R8670 gnd.n5777 gnd.n5776 19.3944
R8671 gnd.n5776 gnd.n854 19.3944
R8672 gnd.n5770 gnd.n854 19.3944
R8673 gnd.n5770 gnd.n5769 19.3944
R8674 gnd.n5769 gnd.n5768 19.3944
R8675 gnd.n5768 gnd.n862 19.3944
R8676 gnd.n5762 gnd.n862 19.3944
R8677 gnd.n5762 gnd.n5761 19.3944
R8678 gnd.n5761 gnd.n5760 19.3944
R8679 gnd.n5760 gnd.n870 19.3944
R8680 gnd.n5754 gnd.n870 19.3944
R8681 gnd.n5754 gnd.n5753 19.3944
R8682 gnd.n5753 gnd.n5752 19.3944
R8683 gnd.n5752 gnd.n878 19.3944
R8684 gnd.n5746 gnd.n878 19.3944
R8685 gnd.n5746 gnd.n5745 19.3944
R8686 gnd.n5745 gnd.n5744 19.3944
R8687 gnd.n5744 gnd.n886 19.3944
R8688 gnd.n5738 gnd.n886 19.3944
R8689 gnd.n5738 gnd.n5737 19.3944
R8690 gnd.n5737 gnd.n5736 19.3944
R8691 gnd.n5736 gnd.n894 19.3944
R8692 gnd.n5730 gnd.n894 19.3944
R8693 gnd.n5730 gnd.n5729 19.3944
R8694 gnd.n5729 gnd.n5728 19.3944
R8695 gnd.n5728 gnd.n902 19.3944
R8696 gnd.n5722 gnd.n902 19.3944
R8697 gnd.n5722 gnd.n5721 19.3944
R8698 gnd.n5721 gnd.n5720 19.3944
R8699 gnd.n5720 gnd.n910 19.3944
R8700 gnd.n5714 gnd.n910 19.3944
R8701 gnd.n5714 gnd.n5713 19.3944
R8702 gnd.n5713 gnd.n5712 19.3944
R8703 gnd.n5712 gnd.n918 19.3944
R8704 gnd.n5706 gnd.n918 19.3944
R8705 gnd.n5706 gnd.n5705 19.3944
R8706 gnd.n5705 gnd.n5704 19.3944
R8707 gnd.n5704 gnd.n926 19.3944
R8708 gnd.n5698 gnd.n926 19.3944
R8709 gnd.n5698 gnd.n5697 19.3944
R8710 gnd.n5697 gnd.n5696 19.3944
R8711 gnd.n5696 gnd.n934 19.3944
R8712 gnd.n5690 gnd.n934 19.3944
R8713 gnd.n5690 gnd.n5689 19.3944
R8714 gnd.n5689 gnd.n5688 19.3944
R8715 gnd.n5688 gnd.n942 19.3944
R8716 gnd.n5682 gnd.n942 19.3944
R8717 gnd.n5682 gnd.n5681 19.3944
R8718 gnd.n5681 gnd.n5680 19.3944
R8719 gnd.n5680 gnd.n950 19.3944
R8720 gnd.n5674 gnd.n950 19.3944
R8721 gnd.n5674 gnd.n5673 19.3944
R8722 gnd.n5673 gnd.n5672 19.3944
R8723 gnd.n5672 gnd.n958 19.3944
R8724 gnd.n5666 gnd.n958 19.3944
R8725 gnd.n5666 gnd.n5665 19.3944
R8726 gnd.n5665 gnd.n5664 19.3944
R8727 gnd.n5664 gnd.n966 19.3944
R8728 gnd.n5658 gnd.n966 19.3944
R8729 gnd.n5658 gnd.n5657 19.3944
R8730 gnd.n5657 gnd.n5656 19.3944
R8731 gnd.n5656 gnd.n974 19.3944
R8732 gnd.n5650 gnd.n974 19.3944
R8733 gnd.n5650 gnd.n5649 19.3944
R8734 gnd.n5649 gnd.n5648 19.3944
R8735 gnd.n5648 gnd.n982 19.3944
R8736 gnd.n5642 gnd.n982 19.3944
R8737 gnd.n5642 gnd.n5641 19.3944
R8738 gnd.n5641 gnd.n5640 19.3944
R8739 gnd.n5640 gnd.n990 19.3944
R8740 gnd.n5634 gnd.n990 19.3944
R8741 gnd.n5634 gnd.n5633 19.3944
R8742 gnd.n5633 gnd.n5632 19.3944
R8743 gnd.n5632 gnd.n998 19.3944
R8744 gnd.n5626 gnd.n998 19.3944
R8745 gnd.n5626 gnd.n5625 19.3944
R8746 gnd.n5625 gnd.n5624 19.3944
R8747 gnd.n5624 gnd.n1006 19.3944
R8748 gnd.n2633 gnd.n2081 19.3944
R8749 gnd.n2081 gnd.n2060 19.3944
R8750 gnd.n2658 gnd.n2060 19.3944
R8751 gnd.n2658 gnd.n2057 19.3944
R8752 gnd.n2663 gnd.n2057 19.3944
R8753 gnd.n2663 gnd.n2058 19.3944
R8754 gnd.n2058 gnd.n2035 19.3944
R8755 gnd.n2688 gnd.n2035 19.3944
R8756 gnd.n2688 gnd.n2032 19.3944
R8757 gnd.n2693 gnd.n2032 19.3944
R8758 gnd.n2693 gnd.n2033 19.3944
R8759 gnd.n2033 gnd.n2010 19.3944
R8760 gnd.n2718 gnd.n2010 19.3944
R8761 gnd.n2718 gnd.n2007 19.3944
R8762 gnd.n2723 gnd.n2007 19.3944
R8763 gnd.n2723 gnd.n2008 19.3944
R8764 gnd.n2008 gnd.n1985 19.3944
R8765 gnd.n2765 gnd.n1985 19.3944
R8766 gnd.n2765 gnd.n1982 19.3944
R8767 gnd.n2770 gnd.n1982 19.3944
R8768 gnd.n2770 gnd.n1983 19.3944
R8769 gnd.n1983 gnd.n1477 19.3944
R8770 gnd.n3792 gnd.n1477 19.3944
R8771 gnd.n3792 gnd.n1478 19.3944
R8772 gnd.n3788 gnd.n1478 19.3944
R8773 gnd.n3788 gnd.n3787 19.3944
R8774 gnd.n3787 gnd.n3786 19.3944
R8775 gnd.n3786 gnd.n1484 19.3944
R8776 gnd.n3782 gnd.n1484 19.3944
R8777 gnd.n3782 gnd.n3781 19.3944
R8778 gnd.n3781 gnd.n3780 19.3944
R8779 gnd.n3780 gnd.n1489 19.3944
R8780 gnd.n3776 gnd.n1489 19.3944
R8781 gnd.n3776 gnd.n3775 19.3944
R8782 gnd.n3775 gnd.n3774 19.3944
R8783 gnd.n3774 gnd.n1494 19.3944
R8784 gnd.n3770 gnd.n1494 19.3944
R8785 gnd.n3770 gnd.n3769 19.3944
R8786 gnd.n3769 gnd.n3768 19.3944
R8787 gnd.n3768 gnd.n1499 19.3944
R8788 gnd.n3764 gnd.n1499 19.3944
R8789 gnd.n3764 gnd.n3763 19.3944
R8790 gnd.n3763 gnd.n3762 19.3944
R8791 gnd.n3762 gnd.n1504 19.3944
R8792 gnd.n3758 gnd.n1504 19.3944
R8793 gnd.n3758 gnd.n3757 19.3944
R8794 gnd.n3757 gnd.n3756 19.3944
R8795 gnd.n3756 gnd.n1509 19.3944
R8796 gnd.n3752 gnd.n1509 19.3944
R8797 gnd.n3752 gnd.n3751 19.3944
R8798 gnd.n3751 gnd.n3750 19.3944
R8799 gnd.n3750 gnd.n1514 19.3944
R8800 gnd.n3746 gnd.n1514 19.3944
R8801 gnd.n3746 gnd.n3745 19.3944
R8802 gnd.n3745 gnd.n3744 19.3944
R8803 gnd.n3744 gnd.n1519 19.3944
R8804 gnd.n3740 gnd.n1519 19.3944
R8805 gnd.n3740 gnd.n3739 19.3944
R8806 gnd.n3739 gnd.n3738 19.3944
R8807 gnd.n3738 gnd.n1524 19.3944
R8808 gnd.n3734 gnd.n1524 19.3944
R8809 gnd.n3734 gnd.n3733 19.3944
R8810 gnd.n3733 gnd.n3732 19.3944
R8811 gnd.n3732 gnd.n1529 19.3944
R8812 gnd.n3728 gnd.n1529 19.3944
R8813 gnd.n3728 gnd.n3727 19.3944
R8814 gnd.n3727 gnd.n3726 19.3944
R8815 gnd.n3726 gnd.n1534 19.3944
R8816 gnd.n3722 gnd.n1534 19.3944
R8817 gnd.n3722 gnd.n3721 19.3944
R8818 gnd.n3721 gnd.n3720 19.3944
R8819 gnd.n3720 gnd.n1539 19.3944
R8820 gnd.n3716 gnd.n1539 19.3944
R8821 gnd.n3716 gnd.n3715 19.3944
R8822 gnd.n3715 gnd.n3714 19.3944
R8823 gnd.n3714 gnd.n1544 19.3944
R8824 gnd.n3710 gnd.n1544 19.3944
R8825 gnd.n3710 gnd.n3709 19.3944
R8826 gnd.n3709 gnd.n3708 19.3944
R8827 gnd.n3708 gnd.n1549 19.3944
R8828 gnd.n3704 gnd.n1549 19.3944
R8829 gnd.n3704 gnd.n3703 19.3944
R8830 gnd.n3703 gnd.n3702 19.3944
R8831 gnd.n3702 gnd.n1554 19.3944
R8832 gnd.n3698 gnd.n1554 19.3944
R8833 gnd.n3698 gnd.n3697 19.3944
R8834 gnd.n3697 gnd.n3696 19.3944
R8835 gnd.n3696 gnd.n1559 19.3944
R8836 gnd.n3692 gnd.n1559 19.3944
R8837 gnd.n3692 gnd.n3691 19.3944
R8838 gnd.n3691 gnd.n3690 19.3944
R8839 gnd.n3690 gnd.n1564 19.3944
R8840 gnd.n3686 gnd.n1564 19.3944
R8841 gnd.n3686 gnd.n3685 19.3944
R8842 gnd.n3685 gnd.n3684 19.3944
R8843 gnd.n3684 gnd.n1569 19.3944
R8844 gnd.n3680 gnd.n1569 19.3944
R8845 gnd.n3680 gnd.n3679 19.3944
R8846 gnd.n3679 gnd.n3678 19.3944
R8847 gnd.n3678 gnd.n461 19.3944
R8848 gnd.n6369 gnd.n461 19.3944
R8849 gnd.n6366 gnd.n6365 19.3944
R8850 gnd.n6365 gnd.n6364 19.3944
R8851 gnd.n6364 gnd.n466 19.3944
R8852 gnd.n6360 gnd.n466 19.3944
R8853 gnd.n6360 gnd.n6359 19.3944
R8854 gnd.n6359 gnd.n391 19.3944
R8855 gnd.n6431 gnd.n391 19.3944
R8856 gnd.n6431 gnd.n6430 19.3944
R8857 gnd.n6430 gnd.n6429 19.3944
R8858 gnd.n6429 gnd.n395 19.3944
R8859 gnd.n6422 gnd.n395 19.3944
R8860 gnd.n6422 gnd.n6421 19.3944
R8861 gnd.n6421 gnd.n405 19.3944
R8862 gnd.n6414 gnd.n405 19.3944
R8863 gnd.n6414 gnd.n6413 19.3944
R8864 gnd.n6413 gnd.n415 19.3944
R8865 gnd.n6406 gnd.n415 19.3944
R8866 gnd.n6406 gnd.n6405 19.3944
R8867 gnd.n6405 gnd.n423 19.3944
R8868 gnd.n6398 gnd.n423 19.3944
R8869 gnd.n6398 gnd.n6397 19.3944
R8870 gnd.n6397 gnd.n433 19.3944
R8871 gnd.n6390 gnd.n433 19.3944
R8872 gnd.n6390 gnd.n6389 19.3944
R8873 gnd.n6379 gnd.n449 19.3944
R8874 gnd.n6379 gnd.n6378 19.3944
R8875 gnd.n6378 gnd.n452 19.3944
R8876 gnd.n5622 gnd.n5621 19.3895
R8877 gnd.n5007 gnd.t288 18.8012
R8878 gnd.n4992 gnd.t325 18.8012
R8879 gnd.n3799 gnd.n3798 18.5761
R8880 gnd.n3492 gnd.n3491 18.5761
R8881 gnd.n4851 gnd.n4850 18.4825
R8882 gnd.n6498 gnd.n6497 18.4247
R8883 gnd.n3870 gnd.n3869 18.4247
R8884 gnd.n6386 gnd.n6385 18.2308
R8885 gnd.n6801 gnd.n6753 18.2308
R8886 gnd.n2572 gnd.n2571 18.2308
R8887 gnd.n2362 gnd.n2361 18.2308
R8888 gnd.t268 gnd.n4531 18.1639
R8889 gnd.n3951 gnd.n1291 18.1639
R8890 gnd.n6621 gnd.n229 18.1639
R8891 gnd.n4559 gnd.t267 17.5266
R8892 gnd.n4958 gnd.t272 16.8893
R8893 gnd.n4049 gnd.t95 16.8893
R8894 gnd.t4 gnd.n1302 16.8893
R8895 gnd.n3927 gnd.t99 16.8893
R8896 gnd.n6556 gnd.t66 16.8893
R8897 gnd.n516 gnd.t24 16.8893
R8898 gnd.n7069 gnd.t62 16.8893
R8899 gnd.n6981 gnd.n6978 16.6793
R8900 gnd.n6480 gnd.n6477 16.6793
R8901 gnd.n4100 gnd.n4097 16.6793
R8902 gnd.n2192 gnd.n2166 16.6793
R8903 gnd.n4786 gnd.t168 16.2519
R8904 gnd.n4486 gnd.t274 16.2519
R8905 gnd.n2635 gnd.n2077 15.9333
R8906 gnd.n2635 gnd.n2078 15.9333
R8907 gnd.n2078 gnd.n2071 15.9333
R8908 gnd.n2645 gnd.n2071 15.9333
R8909 gnd.n2644 gnd.n2062 15.9333
R8910 gnd.n2656 gnd.n2062 15.9333
R8911 gnd.n2656 gnd.n2655 15.9333
R8912 gnd.n2655 gnd.n2064 15.9333
R8913 gnd.n2064 gnd.n2053 15.9333
R8914 gnd.n2665 gnd.n2053 15.9333
R8915 gnd.n2665 gnd.n2054 15.9333
R8916 gnd.n2054 gnd.n2046 15.9333
R8917 gnd.n2675 gnd.n2046 15.9333
R8918 gnd.n2674 gnd.n2037 15.9333
R8919 gnd.n2686 gnd.n2037 15.9333
R8920 gnd.n2686 gnd.n2685 15.9333
R8921 gnd.n2685 gnd.n2039 15.9333
R8922 gnd.n2039 gnd.n2027 15.9333
R8923 gnd.n2695 gnd.n2027 15.9333
R8924 gnd.n2695 gnd.n2028 15.9333
R8925 gnd.n2030 gnd.n2028 15.9333
R8926 gnd.n2705 gnd.n2704 15.9333
R8927 gnd.n2704 gnd.n2012 15.9333
R8928 gnd.n2716 gnd.n2012 15.9333
R8929 gnd.n2716 gnd.n2715 15.9333
R8930 gnd.n2715 gnd.n2014 15.9333
R8931 gnd.n2014 gnd.n2003 15.9333
R8932 gnd.n2725 gnd.n2003 15.9333
R8933 gnd.n2725 gnd.n2004 15.9333
R8934 gnd.n2739 gnd.n1996 15.9333
R8935 gnd.n2739 gnd.n2738 15.9333
R8936 gnd.n2738 gnd.n1987 15.9333
R8937 gnd.n2763 gnd.n1987 15.9333
R8938 gnd.n2763 gnd.n2762 15.9333
R8939 gnd.n2762 gnd.n1989 15.9333
R8940 gnd.n1989 gnd.n1979 15.9333
R8941 gnd.n2772 gnd.n1979 15.9333
R8942 gnd.n2756 gnd.n1413 15.9333
R8943 gnd.n2894 gnd.n1445 15.9333
R8944 gnd.n3794 gnd.n1474 15.9333
R8945 gnd.n2905 gnd.n2904 15.9333
R8946 gnd.n2880 gnd.n1957 15.9333
R8947 gnd.n2950 gnd.n2949 15.9333
R8948 gnd.n2958 gnd.n1922 15.9333
R8949 gnd.n3041 gnd.n1881 15.9333
R8950 gnd.n3083 gnd.n1855 15.9333
R8951 gnd.n3104 gnd.n3103 15.9333
R8952 gnd.n3094 gnd.n3093 15.9333
R8953 gnd.n3124 gnd.n1824 15.9333
R8954 gnd.n1831 gnd.n1819 15.9333
R8955 gnd.n3164 gnd.n1801 15.9333
R8956 gnd.n3204 gnd.n1779 15.9333
R8957 gnd.n1740 gnd.n1728 15.9333
R8958 gnd.n3336 gnd.n1718 15.9333
R8959 gnd.n3348 gnd.n3346 15.9333
R8960 gnd.n3365 gnd.n1698 15.9333
R8961 gnd.n3386 gnd.n1693 15.9333
R8962 gnd.n3400 gnd.n1684 15.9333
R8963 gnd.n1676 gnd.n1636 15.9333
R8964 gnd.n3575 gnd.n1630 15.9333
R8965 gnd.n3575 gnd.n3574 15.9333
R8966 gnd.n3574 gnd.n3573 15.9333
R8967 gnd.n3573 gnd.n1624 15.9333
R8968 gnd.n3583 gnd.n1624 15.9333
R8969 gnd.n3587 gnd.n3583 15.9333
R8970 gnd.n3587 gnd.n3585 15.9333
R8971 gnd.n3585 gnd.n3584 15.9333
R8972 gnd.n3597 gnd.n3596 15.9333
R8973 gnd.n3596 gnd.n3595 15.9333
R8974 gnd.n3595 gnd.n1613 15.9333
R8975 gnd.n3605 gnd.n1613 15.9333
R8976 gnd.n3608 gnd.n3605 15.9333
R8977 gnd.n3608 gnd.n3606 15.9333
R8978 gnd.n3606 gnd.n1607 15.9333
R8979 gnd.n3618 gnd.n1607 15.9333
R8980 gnd.n3617 gnd.n3616 15.9333
R8981 gnd.n3616 gnd.n1601 15.9333
R8982 gnd.n3626 gnd.n1601 15.9333
R8983 gnd.n3629 gnd.n3626 15.9333
R8984 gnd.n3629 gnd.n3627 15.9333
R8985 gnd.n3627 gnd.n1595 15.9333
R8986 gnd.n3639 gnd.n1595 15.9333
R8987 gnd.n3639 gnd.n3638 15.9333
R8988 gnd.n3637 gnd.n1589 15.9333
R8989 gnd.n3647 gnd.n1589 15.9333
R8990 gnd.n3650 gnd.n3647 15.9333
R8991 gnd.n3650 gnd.n3648 15.9333
R8992 gnd.n3648 gnd.n1582 15.9333
R8993 gnd.n3660 gnd.n1582 15.9333
R8994 gnd.n3660 gnd.n3659 15.9333
R8995 gnd.n3659 gnd.n1573 15.9333
R8996 gnd.n3675 gnd.n1573 15.9333
R8997 gnd.n3674 gnd.n1575 15.9333
R8998 gnd.n1575 gnd.n457 15.9333
R8999 gnd.n6371 gnd.n457 15.9333
R9000 gnd.n6371 gnd.n458 15.9333
R9001 gnd.n5473 gnd.n5471 15.6674
R9002 gnd.n5441 gnd.n5439 15.6674
R9003 gnd.n5409 gnd.n5407 15.6674
R9004 gnd.n5378 gnd.n5376 15.6674
R9005 gnd.n5346 gnd.n5344 15.6674
R9006 gnd.n5314 gnd.n5312 15.6674
R9007 gnd.n5282 gnd.n5280 15.6674
R9008 gnd.n5251 gnd.n5249 15.6674
R9009 gnd.n4777 gnd.t168 15.6146
R9010 gnd.t77 gnd.n4240 15.6146
R9011 gnd.t178 gnd.n4241 15.6146
R9012 gnd.n7062 gnd.n6738 15.3217
R9013 gnd.n6437 gnd.n385 15.3217
R9014 gnd.n4057 gnd.n1126 15.3217
R9015 gnd.n2246 gnd.n2154 15.3217
R9016 gnd.n2961 gnd.n2959 15.296
R9017 gnd.n2979 gnd.n1918 15.296
R9018 gnd.t229 gnd.n2990 15.296
R9019 gnd.n3095 gnd.n1841 15.296
R9020 gnd.n3145 gnd.n3144 15.296
R9021 gnd.n3269 gnd.t23 15.296
R9022 gnd.n3284 gnd.n3283 15.296
R9023 gnd.n3303 gnd.n3302 15.296
R9024 gnd.n3409 gnd.n3408 15.0827
R9025 gnd.n1457 gnd.n1452 15.0481
R9026 gnd.n3419 gnd.n3418 15.0481
R9027 gnd.n5145 gnd.t265 14.9773
R9028 gnd.n1146 gnd.t95 14.9773
R9029 gnd.n2772 gnd.t29 14.9773
R9030 gnd.t321 gnd.n1630 14.9773
R9031 gnd.t62 gnd.n154 14.9773
R9032 gnd.n3795 gnd.n1471 14.6587
R9033 gnd.n3031 gnd.n3030 14.6587
R9034 gnd.n3240 gnd.n1775 14.6587
R9035 gnd.n3366 gnd.n1703 14.6587
R9036 gnd.t227 gnd.n4283 14.34
R9037 gnd.n5223 gnd.t271 14.34
R9038 gnd.t116 gnd.n2923 14.0214
R9039 gnd.n2940 gnd.n1938 14.0214
R9040 gnd.n3000 gnd.n1903 14.0214
R9041 gnd.n3105 gnd.n1846 14.0214
R9042 gnd.n3135 gnd.n3134 14.0214
R9043 gnd.n1761 gnd.n1754 14.0214
R9044 gnd.n3335 gnd.n1720 14.0214
R9045 gnd.t138 gnd.n3563 14.0214
R9046 gnd.n4933 gnd.t318 13.7027
R9047 gnd.n1299 gnd.n1291 13.7027
R9048 gnd.t234 gnd.n3057 13.7027
R9049 gnd.t218 gnd.n1796 13.7027
R9050 gnd.n6610 gnd.n229 13.7027
R9051 gnd.n4643 gnd.n4642 13.5763
R9052 gnd.n5587 gnd.n4197 13.5763
R9053 gnd.n4851 gnd.n4589 13.384
R9054 gnd.n2873 gnd.n2872 13.384
R9055 gnd.n2850 gnd.n1905 13.384
R9056 gnd.t35 gnd.n1894 13.384
R9057 gnd.n3250 gnd.t57 13.384
R9058 gnd.n3217 gnd.n1759 13.384
R9059 gnd.n3311 gnd.n1710 13.384
R9060 gnd.n1468 gnd.n1449 13.1884
R9061 gnd.n1463 gnd.n1462 13.1884
R9062 gnd.n1462 gnd.n1461 13.1884
R9063 gnd.n3412 gnd.n3407 13.1884
R9064 gnd.n3413 gnd.n3412 13.1884
R9065 gnd.n1464 gnd.n1451 13.146
R9066 gnd.n1460 gnd.n1451 13.146
R9067 gnd.n3411 gnd.n3410 13.146
R9068 gnd.n3411 gnd.n3406 13.146
R9069 gnd.n3865 gnd.n1445 13.0654
R9070 gnd.n3387 gnd.t45 13.0654
R9071 gnd.n3562 gnd.n1636 13.0654
R9072 gnd.n5474 gnd.n5470 12.8005
R9073 gnd.n5442 gnd.n5438 12.8005
R9074 gnd.n5410 gnd.n5406 12.8005
R9075 gnd.n5379 gnd.n5375 12.8005
R9076 gnd.n5347 gnd.n5343 12.8005
R9077 gnd.n5315 gnd.n5311 12.8005
R9078 gnd.n5283 gnd.n5279 12.8005
R9079 gnd.n5252 gnd.n5248 12.8005
R9080 gnd.n2932 gnd.n2930 12.7467
R9081 gnd.n3075 gnd.n3074 12.7467
R9082 gnd.n3185 gnd.n3184 12.7467
R9083 gnd.n3326 gnd.n1711 12.7467
R9084 gnd.t192 gnd.n2674 12.4281
R9085 gnd.n3638 gnd.t280 12.4281
R9086 gnd.n4642 gnd.n4637 12.4126
R9087 gnd.n5590 gnd.n5587 12.4126
R9088 gnd.n3862 gnd.n3799 12.1761
R9089 gnd.n3491 gnd.n3490 12.1761
R9090 gnd.n2948 gnd.n1940 12.1094
R9091 gnd.n2993 gnd.n1909 12.1094
R9092 gnd.n3267 gnd.n1745 12.1094
R9093 gnd.n3319 gnd.n3318 12.1094
R9094 gnd.n5478 gnd.n5477 12.0247
R9095 gnd.n5446 gnd.n5445 12.0247
R9096 gnd.n5414 gnd.n5413 12.0247
R9097 gnd.n5383 gnd.n5382 12.0247
R9098 gnd.n5351 gnd.n5350 12.0247
R9099 gnd.n5319 gnd.n5318 12.0247
R9100 gnd.n5287 gnd.n5286 12.0247
R9101 gnd.n5256 gnd.n5255 12.0247
R9102 gnd.t52 gnd.n1159 11.7908
R9103 gnd.n2496 gnd.t4 11.7908
R9104 gnd.n2534 gnd.t99 11.7908
R9105 gnd.n6338 gnd.t66 11.7908
R9106 gnd.n6591 gnd.t24 11.7908
R9107 gnd.n142 gnd.t21 11.7908
R9108 gnd.n2881 gnd.n1966 11.4721
R9109 gnd.n2841 gnd.t187 11.4721
R9110 gnd.n2842 gnd.n1879 11.4721
R9111 gnd.n1874 gnd.n1868 11.4721
R9112 gnd.n3175 gnd.n3174 11.4721
R9113 gnd.n3233 gnd.n1772 11.4721
R9114 gnd.n3242 gnd.t261 11.4721
R9115 gnd.n3380 gnd.n3379 11.4721
R9116 gnd.n3401 gnd.n1681 11.4721
R9117 gnd.n1683 gnd.t103 11.4721
R9118 gnd.n5481 gnd.n5468 11.249
R9119 gnd.n5449 gnd.n5436 11.249
R9120 gnd.n5417 gnd.n5404 11.249
R9121 gnd.n5386 gnd.n5373 11.249
R9122 gnd.n5354 gnd.n5341 11.249
R9123 gnd.n5322 gnd.n5309 11.249
R9124 gnd.n5290 gnd.n5277 11.249
R9125 gnd.n5259 gnd.n5246 11.249
R9126 gnd.n4921 gnd.t318 11.1535
R9127 gnd.t206 gnd.n1196 11.1535
R9128 gnd.n1269 gnd.t47 11.1535
R9129 gnd.n2004 gnd.t0 11.1535
R9130 gnd.n3024 gnd.t278 11.1535
R9131 gnd.n3251 gnd.t327 11.1535
R9132 gnd.n3597 gnd.t246 11.1535
R9133 gnd.n212 gnd.t54 11.1535
R9134 gnd.n104 gnd.t254 11.1535
R9135 gnd.n2973 gnd.n2972 10.8348
R9136 gnd.n2972 gnd.n2971 10.8348
R9137 gnd.n3123 gnd.n1834 10.8348
R9138 gnd.n3125 gnd.n3123 10.8348
R9139 gnd.n3292 gnd.n1737 10.8348
R9140 gnd.n1741 gnd.n1737 10.8348
R9141 gnd.n6939 gnd.n6738 10.6672
R9142 gnd.n6440 gnd.n6437 10.6672
R9143 gnd.n4060 gnd.n4057 10.6672
R9144 gnd.n2242 gnd.n2154 10.6672
R9145 gnd.n3559 gnd.n3558 10.6151
R9146 gnd.n3558 gnd.n3555 10.6151
R9147 gnd.n3553 gnd.n3550 10.6151
R9148 gnd.n3550 gnd.n3549 10.6151
R9149 gnd.n3549 gnd.n3546 10.6151
R9150 gnd.n3546 gnd.n3545 10.6151
R9151 gnd.n3545 gnd.n3542 10.6151
R9152 gnd.n3542 gnd.n3541 10.6151
R9153 gnd.n3541 gnd.n3538 10.6151
R9154 gnd.n3538 gnd.n3537 10.6151
R9155 gnd.n3537 gnd.n3534 10.6151
R9156 gnd.n3534 gnd.n3533 10.6151
R9157 gnd.n3533 gnd.n3530 10.6151
R9158 gnd.n3530 gnd.n3529 10.6151
R9159 gnd.n3529 gnd.n3526 10.6151
R9160 gnd.n3526 gnd.n3525 10.6151
R9161 gnd.n3525 gnd.n3522 10.6151
R9162 gnd.n3522 gnd.n3521 10.6151
R9163 gnd.n3521 gnd.n3518 10.6151
R9164 gnd.n3518 gnd.n3517 10.6151
R9165 gnd.n3517 gnd.n3514 10.6151
R9166 gnd.n3514 gnd.n3513 10.6151
R9167 gnd.n3513 gnd.n3510 10.6151
R9168 gnd.n3510 gnd.n3509 10.6151
R9169 gnd.n3509 gnd.n3506 10.6151
R9170 gnd.n3506 gnd.n3505 10.6151
R9171 gnd.n3505 gnd.n3502 10.6151
R9172 gnd.n3502 gnd.n3501 10.6151
R9173 gnd.n3501 gnd.n3498 10.6151
R9174 gnd.n3498 gnd.n3497 10.6151
R9175 gnd.n2891 gnd.n2890 10.6151
R9176 gnd.n2890 gnd.n2889 10.6151
R9177 gnd.n2889 gnd.n2886 10.6151
R9178 gnd.n2886 gnd.n2885 10.6151
R9179 gnd.n2885 gnd.n2884 10.6151
R9180 gnd.n2884 gnd.n2883 10.6151
R9181 gnd.n2883 gnd.n2879 10.6151
R9182 gnd.n2879 gnd.n2878 10.6151
R9183 gnd.n2878 gnd.n2876 10.6151
R9184 gnd.n2876 gnd.n2875 10.6151
R9185 gnd.n2875 gnd.n2870 10.6151
R9186 gnd.n2870 gnd.n2869 10.6151
R9187 gnd.n2869 gnd.n2867 10.6151
R9188 gnd.n2867 gnd.n2866 10.6151
R9189 gnd.n2866 gnd.n2863 10.6151
R9190 gnd.n2863 gnd.n2862 10.6151
R9191 gnd.n2862 gnd.n2861 10.6151
R9192 gnd.n2861 gnd.n2860 10.6151
R9193 gnd.n2860 gnd.n2859 10.6151
R9194 gnd.n2859 gnd.n2856 10.6151
R9195 gnd.n2856 gnd.n2855 10.6151
R9196 gnd.n2855 gnd.n2853 10.6151
R9197 gnd.n2853 gnd.n2852 10.6151
R9198 gnd.n2852 gnd.n2848 10.6151
R9199 gnd.n2848 gnd.n2847 10.6151
R9200 gnd.n2847 gnd.n2845 10.6151
R9201 gnd.n2845 gnd.n2844 10.6151
R9202 gnd.n2844 gnd.n2840 10.6151
R9203 gnd.n2840 gnd.n1871 10.6151
R9204 gnd.n3051 gnd.n1871 10.6151
R9205 gnd.n3052 gnd.n3051 10.6151
R9206 gnd.n3053 gnd.n3052 10.6151
R9207 gnd.n3053 gnd.n1862 10.6151
R9208 gnd.n3072 gnd.n1862 10.6151
R9209 gnd.n3072 gnd.n3071 10.6151
R9210 gnd.n3071 gnd.n3070 10.6151
R9211 gnd.n3070 gnd.n1849 10.6151
R9212 gnd.n3099 gnd.n1849 10.6151
R9213 gnd.n3099 gnd.n3098 10.6151
R9214 gnd.n3098 gnd.n3097 10.6151
R9215 gnd.n3097 gnd.n1832 10.6151
R9216 gnd.n3127 gnd.n1832 10.6151
R9217 gnd.n3128 gnd.n3127 10.6151
R9218 gnd.n3130 gnd.n3128 10.6151
R9219 gnd.n3131 gnd.n3130 10.6151
R9220 gnd.n3132 gnd.n3131 10.6151
R9221 gnd.n3132 gnd.n1809 10.6151
R9222 gnd.n3167 gnd.n1809 10.6151
R9223 gnd.n3168 gnd.n3167 10.6151
R9224 gnd.n3170 gnd.n3168 10.6151
R9225 gnd.n3171 gnd.n3170 10.6151
R9226 gnd.n3172 gnd.n3171 10.6151
R9227 gnd.n3172 gnd.n1786 10.6151
R9228 gnd.n3206 gnd.n1786 10.6151
R9229 gnd.n3207 gnd.n3206 10.6151
R9230 gnd.n3209 gnd.n3207 10.6151
R9231 gnd.n3210 gnd.n3209 10.6151
R9232 gnd.n3212 gnd.n3210 10.6151
R9233 gnd.n3212 gnd.n3211 10.6151
R9234 gnd.n3211 gnd.n1757 10.6151
R9235 gnd.n3260 gnd.n1757 10.6151
R9236 gnd.n3261 gnd.n3260 10.6151
R9237 gnd.n3265 gnd.n3261 10.6151
R9238 gnd.n3265 gnd.n3264 10.6151
R9239 gnd.n3264 gnd.n3263 10.6151
R9240 gnd.n3263 gnd.n3262 10.6151
R9241 gnd.n3262 gnd.n1726 10.6151
R9242 gnd.n3305 gnd.n1726 10.6151
R9243 gnd.n3306 gnd.n3305 10.6151
R9244 gnd.n3316 gnd.n3306 10.6151
R9245 gnd.n3316 gnd.n3315 10.6151
R9246 gnd.n3315 gnd.n3314 10.6151
R9247 gnd.n3314 gnd.n3307 10.6151
R9248 gnd.n3308 gnd.n3307 10.6151
R9249 gnd.n3308 gnd.n1701 10.6151
R9250 gnd.n3368 gnd.n1701 10.6151
R9251 gnd.n3369 gnd.n3368 10.6151
R9252 gnd.n3376 gnd.n3369 10.6151
R9253 gnd.n3376 gnd.n3375 10.6151
R9254 gnd.n3375 gnd.n3374 10.6151
R9255 gnd.n3374 gnd.n3371 10.6151
R9256 gnd.n3371 gnd.n3370 10.6151
R9257 gnd.n3370 gnd.n1673 10.6151
R9258 gnd.n2778 gnd.n1409 10.6151
R9259 gnd.n2781 gnd.n2778 10.6151
R9260 gnd.n2786 gnd.n2783 10.6151
R9261 gnd.n2787 gnd.n2786 10.6151
R9262 gnd.n2790 gnd.n2787 10.6151
R9263 gnd.n2791 gnd.n2790 10.6151
R9264 gnd.n2794 gnd.n2791 10.6151
R9265 gnd.n2795 gnd.n2794 10.6151
R9266 gnd.n2798 gnd.n2795 10.6151
R9267 gnd.n2799 gnd.n2798 10.6151
R9268 gnd.n2802 gnd.n2799 10.6151
R9269 gnd.n2803 gnd.n2802 10.6151
R9270 gnd.n2806 gnd.n2803 10.6151
R9271 gnd.n2807 gnd.n2806 10.6151
R9272 gnd.n2810 gnd.n2807 10.6151
R9273 gnd.n2811 gnd.n2810 10.6151
R9274 gnd.n2814 gnd.n2811 10.6151
R9275 gnd.n2815 gnd.n2814 10.6151
R9276 gnd.n2818 gnd.n2815 10.6151
R9277 gnd.n2819 gnd.n2818 10.6151
R9278 gnd.n2822 gnd.n2819 10.6151
R9279 gnd.n2823 gnd.n2822 10.6151
R9280 gnd.n2826 gnd.n2823 10.6151
R9281 gnd.n2827 gnd.n2826 10.6151
R9282 gnd.n2830 gnd.n2827 10.6151
R9283 gnd.n2831 gnd.n2830 10.6151
R9284 gnd.n2834 gnd.n2831 10.6151
R9285 gnd.n2835 gnd.n2834 10.6151
R9286 gnd.n2838 gnd.n2835 10.6151
R9287 gnd.n2839 gnd.n2838 10.6151
R9288 gnd.n3862 gnd.n3861 10.6151
R9289 gnd.n3861 gnd.n3860 10.6151
R9290 gnd.n3860 gnd.n3859 10.6151
R9291 gnd.n3859 gnd.n3857 10.6151
R9292 gnd.n3857 gnd.n3854 10.6151
R9293 gnd.n3854 gnd.n3853 10.6151
R9294 gnd.n3853 gnd.n3850 10.6151
R9295 gnd.n3850 gnd.n3849 10.6151
R9296 gnd.n3849 gnd.n3846 10.6151
R9297 gnd.n3846 gnd.n3845 10.6151
R9298 gnd.n3845 gnd.n3842 10.6151
R9299 gnd.n3842 gnd.n3841 10.6151
R9300 gnd.n3841 gnd.n3838 10.6151
R9301 gnd.n3838 gnd.n3837 10.6151
R9302 gnd.n3837 gnd.n3834 10.6151
R9303 gnd.n3834 gnd.n3833 10.6151
R9304 gnd.n3833 gnd.n3830 10.6151
R9305 gnd.n3830 gnd.n3829 10.6151
R9306 gnd.n3829 gnd.n3826 10.6151
R9307 gnd.n3826 gnd.n3825 10.6151
R9308 gnd.n3825 gnd.n3822 10.6151
R9309 gnd.n3822 gnd.n3821 10.6151
R9310 gnd.n3821 gnd.n3818 10.6151
R9311 gnd.n3818 gnd.n3817 10.6151
R9312 gnd.n3817 gnd.n3814 10.6151
R9313 gnd.n3814 gnd.n3813 10.6151
R9314 gnd.n3813 gnd.n3810 10.6151
R9315 gnd.n3810 gnd.n3809 10.6151
R9316 gnd.n3806 gnd.n3805 10.6151
R9317 gnd.n3805 gnd.n1410 10.6151
R9318 gnd.n3490 gnd.n3489 10.6151
R9319 gnd.n3489 gnd.n3486 10.6151
R9320 gnd.n3486 gnd.n3485 10.6151
R9321 gnd.n3485 gnd.n3482 10.6151
R9322 gnd.n3482 gnd.n3481 10.6151
R9323 gnd.n3481 gnd.n3478 10.6151
R9324 gnd.n3478 gnd.n3477 10.6151
R9325 gnd.n3477 gnd.n3474 10.6151
R9326 gnd.n3474 gnd.n3473 10.6151
R9327 gnd.n3473 gnd.n3470 10.6151
R9328 gnd.n3470 gnd.n3469 10.6151
R9329 gnd.n3469 gnd.n3466 10.6151
R9330 gnd.n3466 gnd.n3465 10.6151
R9331 gnd.n3465 gnd.n3462 10.6151
R9332 gnd.n3462 gnd.n3461 10.6151
R9333 gnd.n3461 gnd.n3458 10.6151
R9334 gnd.n3458 gnd.n3457 10.6151
R9335 gnd.n3457 gnd.n3454 10.6151
R9336 gnd.n3454 gnd.n3453 10.6151
R9337 gnd.n3453 gnd.n3450 10.6151
R9338 gnd.n3450 gnd.n3449 10.6151
R9339 gnd.n3449 gnd.n3446 10.6151
R9340 gnd.n3446 gnd.n3445 10.6151
R9341 gnd.n3445 gnd.n3442 10.6151
R9342 gnd.n3442 gnd.n3441 10.6151
R9343 gnd.n3441 gnd.n3438 10.6151
R9344 gnd.n3438 gnd.n3437 10.6151
R9345 gnd.n3437 gnd.n3434 10.6151
R9346 gnd.n3432 gnd.n3429 10.6151
R9347 gnd.n3429 gnd.n3428 10.6151
R9348 gnd.n3798 gnd.n3797 10.6151
R9349 gnd.n3797 gnd.n1469 10.6151
R9350 gnd.n2908 gnd.n1469 10.6151
R9351 gnd.n2909 gnd.n2908 10.6151
R9352 gnd.n2910 gnd.n2909 10.6151
R9353 gnd.n2910 gnd.n1955 10.6151
R9354 gnd.n2926 gnd.n1955 10.6151
R9355 gnd.n2927 gnd.n2926 10.6151
R9356 gnd.n2928 gnd.n2927 10.6151
R9357 gnd.n2928 gnd.n1943 10.6151
R9358 gnd.n2943 gnd.n1943 10.6151
R9359 gnd.n2944 gnd.n2943 10.6151
R9360 gnd.n2946 gnd.n2944 10.6151
R9361 gnd.n2946 gnd.n2945 10.6151
R9362 gnd.n2945 gnd.n1920 10.6151
R9363 gnd.n2975 gnd.n1920 10.6151
R9364 gnd.n2976 gnd.n2975 10.6151
R9365 gnd.n2977 gnd.n2976 10.6151
R9366 gnd.n2977 gnd.n1907 10.6151
R9367 gnd.n2995 gnd.n1907 10.6151
R9368 gnd.n2996 gnd.n2995 10.6151
R9369 gnd.n2997 gnd.n2996 10.6151
R9370 gnd.n2997 gnd.n1892 10.6151
R9371 gnd.n3026 gnd.n1892 10.6151
R9372 gnd.n3027 gnd.n3026 10.6151
R9373 gnd.n3028 gnd.n3027 10.6151
R9374 gnd.n3028 gnd.n1877 10.6151
R9375 gnd.n3044 gnd.n1877 10.6151
R9376 gnd.n3045 gnd.n3044 10.6151
R9377 gnd.n3047 gnd.n3045 10.6151
R9378 gnd.n3047 gnd.n3046 10.6151
R9379 gnd.n3046 gnd.n1858 10.6151
R9380 gnd.n3078 gnd.n1858 10.6151
R9381 gnd.n3079 gnd.n3078 10.6151
R9382 gnd.n3080 gnd.n3079 10.6151
R9383 gnd.n3080 gnd.n1844 10.6151
R9384 gnd.n3107 gnd.n1844 10.6151
R9385 gnd.n3108 gnd.n3107 10.6151
R9386 gnd.n3112 gnd.n3108 10.6151
R9387 gnd.n3112 gnd.n3111 10.6151
R9388 gnd.n3111 gnd.n3110 10.6151
R9389 gnd.n3110 gnd.n1822 10.6151
R9390 gnd.n3147 gnd.n1822 10.6151
R9391 gnd.n3148 gnd.n3147 10.6151
R9392 gnd.n3152 gnd.n3148 10.6151
R9393 gnd.n3152 gnd.n3151 10.6151
R9394 gnd.n3151 gnd.n3150 10.6151
R9395 gnd.n3150 gnd.n1799 10.6151
R9396 gnd.n3187 gnd.n1799 10.6151
R9397 gnd.n3188 gnd.n3187 10.6151
R9398 gnd.n3192 gnd.n3188 10.6151
R9399 gnd.n3192 gnd.n3191 10.6151
R9400 gnd.n3191 gnd.n3190 10.6151
R9401 gnd.n3190 gnd.n1777 10.6151
R9402 gnd.n3236 gnd.n1777 10.6151
R9403 gnd.n3237 gnd.n3236 10.6151
R9404 gnd.n3238 gnd.n3237 10.6151
R9405 gnd.n3238 gnd.n1764 10.6151
R9406 gnd.n3253 gnd.n1764 10.6151
R9407 gnd.n3254 gnd.n3253 10.6151
R9408 gnd.n3256 gnd.n3254 10.6151
R9409 gnd.n3256 gnd.n3255 10.6151
R9410 gnd.n3255 gnd.n1743 10.6151
R9411 gnd.n3287 gnd.n1743 10.6151
R9412 gnd.n3288 gnd.n3287 10.6151
R9413 gnd.n3290 gnd.n3288 10.6151
R9414 gnd.n3290 gnd.n3289 10.6151
R9415 gnd.n3289 gnd.n1723 10.6151
R9416 gnd.n3322 gnd.n1723 10.6151
R9417 gnd.n3323 gnd.n3322 10.6151
R9418 gnd.n3333 gnd.n3323 10.6151
R9419 gnd.n3333 gnd.n3332 10.6151
R9420 gnd.n3332 gnd.n3331 10.6151
R9421 gnd.n3331 gnd.n3324 10.6151
R9422 gnd.n3325 gnd.n3324 10.6151
R9423 gnd.n3325 gnd.n1696 10.6151
R9424 gnd.n3382 gnd.n1696 10.6151
R9425 gnd.n3383 gnd.n3382 10.6151
R9426 gnd.n3384 gnd.n3383 10.6151
R9427 gnd.n3384 gnd.n1679 10.6151
R9428 gnd.n3403 gnd.n1679 10.6151
R9429 gnd.n3404 gnd.n3403 10.6151
R9430 gnd.n3492 gnd.n3404 10.6151
R9431 gnd.n4840 gnd.t224 10.5161
R9432 gnd.n4285 gnd.t227 10.5161
R9433 gnd.n5206 gnd.t271 10.5161
R9434 gnd.n1231 gnd.t26 10.5161
R9435 gnd.t11 gnd.n1234 10.5161
R9436 gnd.n2970 gnd.t197 10.5161
R9437 gnd.n3293 gnd.t236 10.5161
R9438 gnd.n6688 gnd.t181 10.5161
R9439 gnd.n6696 gnd.t33 10.5161
R9440 gnd.n5482 gnd.n5466 10.4732
R9441 gnd.n5450 gnd.n5434 10.4732
R9442 gnd.n5418 gnd.n5402 10.4732
R9443 gnd.n5387 gnd.n5371 10.4732
R9444 gnd.n5355 gnd.n5339 10.4732
R9445 gnd.n5323 gnd.n5307 10.4732
R9446 gnd.n5291 gnd.n5275 10.4732
R9447 gnd.n5260 gnd.n5244 10.4732
R9448 gnd.n2906 gnd.n1968 10.1975
R9449 gnd.n2912 gnd.n1966 10.1975
R9450 gnd.n3042 gnd.n1879 10.1975
R9451 gnd.n3049 gnd.n1874 10.1975
R9452 gnd.n3175 gnd.n1788 10.1975
R9453 gnd.n3234 gnd.n3233 10.1975
R9454 gnd.t265 gnd.n4302 9.87883
R9455 gnd.n1193 gnd.t6 9.87883
R9456 gnd.t9 gnd.n1272 9.87883
R9457 gnd.t312 gnd.t175 9.87883
R9458 gnd.t15 gnd.n209 9.87883
R9459 gnd.t13 gnd.n107 9.87883
R9460 gnd.n5486 gnd.n5485 9.69747
R9461 gnd.n5454 gnd.n5453 9.69747
R9462 gnd.n5422 gnd.n5421 9.69747
R9463 gnd.n5391 gnd.n5390 9.69747
R9464 gnd.n5359 gnd.n5358 9.69747
R9465 gnd.n5327 gnd.n5326 9.69747
R9466 gnd.n5295 gnd.n5294 9.69747
R9467 gnd.n5264 gnd.n5263 9.69747
R9468 gnd.n2864 gnd.n1940 9.56018
R9469 gnd.n2857 gnd.n1909 9.56018
R9470 gnd.t185 gnd.n1873 9.56018
R9471 gnd.n3115 gnd.n3114 9.56018
R9472 gnd.n3155 gnd.n1817 9.56018
R9473 gnd.t257 gnd.n3203 9.56018
R9474 gnd.n3285 gnd.n1745 9.56018
R9475 gnd.n3320 gnd.n3319 9.56018
R9476 gnd.n5492 gnd.n5491 9.45567
R9477 gnd.n5460 gnd.n5459 9.45567
R9478 gnd.n5428 gnd.n5427 9.45567
R9479 gnd.n5397 gnd.n5396 9.45567
R9480 gnd.n5365 gnd.n5364 9.45567
R9481 gnd.n5333 gnd.n5332 9.45567
R9482 gnd.n5301 gnd.n5300 9.45567
R9483 gnd.n5270 gnd.n5269 9.45567
R9484 gnd.n6978 gnd.n6918 9.30959
R9485 gnd.n6477 gnd.n6476 9.30959
R9486 gnd.n4097 gnd.n4096 9.30959
R9487 gnd.n2196 gnd.n2166 9.30959
R9488 gnd.n6437 gnd.n6436 9.3005
R9489 gnd.n6440 gnd.n384 9.3005
R9490 gnd.n6441 gnd.n383 9.3005
R9491 gnd.n6444 gnd.n382 9.3005
R9492 gnd.n6445 gnd.n381 9.3005
R9493 gnd.n6448 gnd.n380 9.3005
R9494 gnd.n6449 gnd.n379 9.3005
R9495 gnd.n6452 gnd.n378 9.3005
R9496 gnd.n6453 gnd.n377 9.3005
R9497 gnd.n6456 gnd.n376 9.3005
R9498 gnd.n6457 gnd.n375 9.3005
R9499 gnd.n6460 gnd.n374 9.3005
R9500 gnd.n6461 gnd.n373 9.3005
R9501 gnd.n6464 gnd.n372 9.3005
R9502 gnd.n6465 gnd.n371 9.3005
R9503 gnd.n6468 gnd.n370 9.3005
R9504 gnd.n6469 gnd.n369 9.3005
R9505 gnd.n6472 gnd.n368 9.3005
R9506 gnd.n6473 gnd.n367 9.3005
R9507 gnd.n6476 gnd.n366 9.3005
R9508 gnd.n6480 gnd.n362 9.3005
R9509 gnd.n6481 gnd.n361 9.3005
R9510 gnd.n6484 gnd.n360 9.3005
R9511 gnd.n6485 gnd.n359 9.3005
R9512 gnd.n6488 gnd.n358 9.3005
R9513 gnd.n6489 gnd.n357 9.3005
R9514 gnd.n6492 gnd.n356 9.3005
R9515 gnd.n6493 gnd.n355 9.3005
R9516 gnd.n6496 gnd.n354 9.3005
R9517 gnd.n6498 gnd.n350 9.3005
R9518 gnd.n6501 gnd.n349 9.3005
R9519 gnd.n6502 gnd.n348 9.3005
R9520 gnd.n6505 gnd.n347 9.3005
R9521 gnd.n6506 gnd.n346 9.3005
R9522 gnd.n6509 gnd.n345 9.3005
R9523 gnd.n6510 gnd.n344 9.3005
R9524 gnd.n6513 gnd.n343 9.3005
R9525 gnd.n6515 gnd.n340 9.3005
R9526 gnd.n6518 gnd.n339 9.3005
R9527 gnd.n6519 gnd.n338 9.3005
R9528 gnd.n6522 gnd.n337 9.3005
R9529 gnd.n6523 gnd.n336 9.3005
R9530 gnd.n6526 gnd.n335 9.3005
R9531 gnd.n6527 gnd.n334 9.3005
R9532 gnd.n6530 gnd.n333 9.3005
R9533 gnd.n6531 gnd.n332 9.3005
R9534 gnd.n6534 gnd.n331 9.3005
R9535 gnd.n6535 gnd.n330 9.3005
R9536 gnd.n6538 gnd.n329 9.3005
R9537 gnd.n6539 gnd.n328 9.3005
R9538 gnd.n6542 gnd.n327 9.3005
R9539 gnd.n6543 gnd.n326 9.3005
R9540 gnd.n6544 gnd.n325 9.3005
R9541 gnd.n282 gnd.n281 9.3005
R9542 gnd.n6550 gnd.n6549 9.3005
R9543 gnd.n6477 gnd.n363 9.3005
R9544 gnd.n6435 gnd.n385 9.3005
R9545 gnd.n6554 gnd.n6553 9.3005
R9546 gnd.n6552 gnd.n280 9.3005
R9547 gnd.n253 gnd.n252 9.3005
R9548 gnd.n6584 gnd.n6583 9.3005
R9549 gnd.n6585 gnd.n251 9.3005
R9550 gnd.n6589 gnd.n6586 9.3005
R9551 gnd.n6588 gnd.n6587 9.3005
R9552 gnd.n227 gnd.n226 9.3005
R9553 gnd.n6624 gnd.n6623 9.3005
R9554 gnd.n6625 gnd.n225 9.3005
R9555 gnd.n6627 gnd.n6626 9.3005
R9556 gnd.n207 gnd.n206 9.3005
R9557 gnd.n6648 gnd.n6647 9.3005
R9558 gnd.n6649 gnd.n205 9.3005
R9559 gnd.n6653 gnd.n6650 9.3005
R9560 gnd.n6652 gnd.n6651 9.3005
R9561 gnd.n6551 gnd.n279 9.3005
R9562 gnd.n184 gnd.n183 9.3005
R9563 gnd.n6680 gnd.n6679 9.3005
R9564 gnd.n6681 gnd.n182 9.3005
R9565 gnd.n6686 gnd.n6682 9.3005
R9566 gnd.n6685 gnd.n6684 9.3005
R9567 gnd.n6683 gnd.n78 9.3005
R9568 gnd.n7121 gnd.n79 9.3005
R9569 gnd.n7120 gnd.n80 9.3005
R9570 gnd.n7119 gnd.n81 9.3005
R9571 gnd.n98 gnd.n82 9.3005
R9572 gnd.n7109 gnd.n99 9.3005
R9573 gnd.n7108 gnd.n100 9.3005
R9574 gnd.n7107 gnd.n101 9.3005
R9575 gnd.n118 gnd.n102 9.3005
R9576 gnd.n7097 gnd.n119 9.3005
R9577 gnd.n7096 gnd.n120 9.3005
R9578 gnd.n7095 gnd.n121 9.3005
R9579 gnd.n136 gnd.n122 9.3005
R9580 gnd.n7085 gnd.n137 9.3005
R9581 gnd.n7084 gnd.n138 9.3005
R9582 gnd.n7083 gnd.n139 9.3005
R9583 gnd.n156 gnd.n140 9.3005
R9584 gnd.n7073 gnd.n157 9.3005
R9585 gnd.n7072 gnd.n158 9.3005
R9586 gnd.n7071 gnd.n159 9.3005
R9587 gnd.n6882 gnd.n160 9.3005
R9588 gnd.n7127 gnd.n7126 9.3005
R9589 gnd.n7125 gnd.n69 9.3005
R9590 gnd.n6812 gnd.n71 9.3005
R9591 gnd.n6814 gnd.n6813 9.3005
R9592 gnd.n6817 gnd.n6816 9.3005
R9593 gnd.n6818 gnd.n6811 9.3005
R9594 gnd.n6821 gnd.n6819 9.3005
R9595 gnd.n6822 gnd.n6810 9.3005
R9596 gnd.n6825 gnd.n6824 9.3005
R9597 gnd.n6826 gnd.n6809 9.3005
R9598 gnd.n6829 gnd.n6827 9.3005
R9599 gnd.n6830 gnd.n6808 9.3005
R9600 gnd.n6833 gnd.n6832 9.3005
R9601 gnd.n6834 gnd.n6807 9.3005
R9602 gnd.n6837 gnd.n6835 9.3005
R9603 gnd.n6838 gnd.n6806 9.3005
R9604 gnd.n6841 gnd.n6840 9.3005
R9605 gnd.n6842 gnd.n6805 9.3005
R9606 gnd.n6845 gnd.n6843 9.3005
R9607 gnd.n6846 gnd.n6804 9.3005
R9608 gnd.n6848 gnd.n6847 9.3005
R9609 gnd.n6764 gnd.n6763 9.3005
R9610 gnd.n6766 gnd.n6765 9.3005
R9611 gnd.n6769 gnd.n6760 9.3005
R9612 gnd.n6773 gnd.n6772 9.3005
R9613 gnd.n6774 gnd.n6759 9.3005
R9614 gnd.n6776 gnd.n6775 9.3005
R9615 gnd.n6779 gnd.n6758 9.3005
R9616 gnd.n6783 gnd.n6782 9.3005
R9617 gnd.n6784 gnd.n6757 9.3005
R9618 gnd.n6786 gnd.n6785 9.3005
R9619 gnd.n6789 gnd.n6756 9.3005
R9620 gnd.n6793 gnd.n6792 9.3005
R9621 gnd.n6794 gnd.n6755 9.3005
R9622 gnd.n6796 gnd.n6795 9.3005
R9623 gnd.n6799 gnd.n6754 9.3005
R9624 gnd.n6802 gnd.n6801 9.3005
R9625 gnd.n6803 gnd.n6753 9.3005
R9626 gnd.n6850 gnd.n6849 9.3005
R9627 gnd.n6761 gnd.n6734 9.3005
R9628 gnd.n7055 gnd.n7054 9.3005
R9629 gnd.n7053 gnd.n6884 9.3005
R9630 gnd.n7052 gnd.n7051 9.3005
R9631 gnd.n7048 gnd.n6885 9.3005
R9632 gnd.n7045 gnd.n6886 9.3005
R9633 gnd.n7044 gnd.n6887 9.3005
R9634 gnd.n7041 gnd.n6888 9.3005
R9635 gnd.n7040 gnd.n6889 9.3005
R9636 gnd.n7037 gnd.n6890 9.3005
R9637 gnd.n7036 gnd.n6891 9.3005
R9638 gnd.n7033 gnd.n6892 9.3005
R9639 gnd.n7032 gnd.n6893 9.3005
R9640 gnd.n7029 gnd.n6894 9.3005
R9641 gnd.n7028 gnd.n6895 9.3005
R9642 gnd.n7025 gnd.n6896 9.3005
R9643 gnd.n7024 gnd.n6897 9.3005
R9644 gnd.n7021 gnd.n6898 9.3005
R9645 gnd.n7017 gnd.n6899 9.3005
R9646 gnd.n7014 gnd.n6900 9.3005
R9647 gnd.n7013 gnd.n6901 9.3005
R9648 gnd.n7010 gnd.n6902 9.3005
R9649 gnd.n7009 gnd.n6903 9.3005
R9650 gnd.n7006 gnd.n6904 9.3005
R9651 gnd.n7005 gnd.n6905 9.3005
R9652 gnd.n7002 gnd.n6906 9.3005
R9653 gnd.n7001 gnd.n6907 9.3005
R9654 gnd.n6998 gnd.n6908 9.3005
R9655 gnd.n6997 gnd.n6909 9.3005
R9656 gnd.n6994 gnd.n6910 9.3005
R9657 gnd.n6993 gnd.n6911 9.3005
R9658 gnd.n6990 gnd.n6912 9.3005
R9659 gnd.n6989 gnd.n6913 9.3005
R9660 gnd.n6986 gnd.n6914 9.3005
R9661 gnd.n6985 gnd.n6915 9.3005
R9662 gnd.n6982 gnd.n6916 9.3005
R9663 gnd.n6981 gnd.n6917 9.3005
R9664 gnd.n6978 gnd.n6977 9.3005
R9665 gnd.n6976 gnd.n6918 9.3005
R9666 gnd.n6975 gnd.n6974 9.3005
R9667 gnd.n6971 gnd.n6921 9.3005
R9668 gnd.n6968 gnd.n6922 9.3005
R9669 gnd.n6967 gnd.n6923 9.3005
R9670 gnd.n6964 gnd.n6924 9.3005
R9671 gnd.n6963 gnd.n6925 9.3005
R9672 gnd.n6960 gnd.n6926 9.3005
R9673 gnd.n6959 gnd.n6927 9.3005
R9674 gnd.n6956 gnd.n6928 9.3005
R9675 gnd.n6955 gnd.n6929 9.3005
R9676 gnd.n6952 gnd.n6930 9.3005
R9677 gnd.n6951 gnd.n6931 9.3005
R9678 gnd.n6948 gnd.n6932 9.3005
R9679 gnd.n6947 gnd.n6933 9.3005
R9680 gnd.n6944 gnd.n6934 9.3005
R9681 gnd.n6943 gnd.n6935 9.3005
R9682 gnd.n6940 gnd.n6936 9.3005
R9683 gnd.n6939 gnd.n6937 9.3005
R9684 gnd.n6738 gnd.n6735 9.3005
R9685 gnd.n7063 gnd.n7062 9.3005
R9686 gnd.n7056 gnd.n6883 9.3005
R9687 gnd.n505 gnd.n504 9.3005
R9688 gnd.n506 gnd.n264 9.3005
R9689 gnd.n6567 gnd.n265 9.3005
R9690 gnd.n6568 gnd.n262 9.3005
R9691 gnd.n6571 gnd.n263 9.3005
R9692 gnd.n6573 gnd.n6572 9.3005
R9693 gnd.n6574 gnd.n236 9.3005
R9694 gnd.n6612 gnd.n237 9.3005
R9695 gnd.n6613 gnd.n235 9.3005
R9696 gnd.n6615 gnd.n6614 9.3005
R9697 gnd.n6616 gnd.n218 9.3005
R9698 gnd.n6632 gnd.n219 9.3005
R9699 gnd.n6633 gnd.n216 9.3005
R9700 gnd.n6635 gnd.n217 9.3005
R9701 gnd.n6637 gnd.n6636 9.3005
R9702 gnd.n6638 gnd.n192 9.3005
R9703 gnd.n6670 gnd.n191 9.3005
R9704 gnd.n6674 gnd.n6673 9.3005
R9705 gnd.n6672 gnd.n174 9.3005
R9706 gnd.n6691 gnd.n173 9.3005
R9707 gnd.n6693 gnd.n6692 9.3005
R9708 gnd.n6694 gnd.n168 9.3005
R9709 gnd.n6700 gnd.n167 9.3005
R9710 gnd.n6703 gnd.n6701 9.3005
R9711 gnd.n6704 gnd.n90 9.3005
R9712 gnd.n6706 gnd.n91 9.3005
R9713 gnd.n6707 gnd.n92 9.3005
R9714 gnd.n6710 gnd.n6708 9.3005
R9715 gnd.n6711 gnd.n109 9.3005
R9716 gnd.n6713 gnd.n110 9.3005
R9717 gnd.n6714 gnd.n111 9.3005
R9718 gnd.n6717 gnd.n6715 9.3005
R9719 gnd.n6718 gnd.n128 9.3005
R9720 gnd.n6720 gnd.n129 9.3005
R9721 gnd.n6721 gnd.n130 9.3005
R9722 gnd.n6724 gnd.n6722 9.3005
R9723 gnd.n6725 gnd.n147 9.3005
R9724 gnd.n6727 gnd.n148 9.3005
R9725 gnd.n6728 gnd.n149 9.3005
R9726 gnd.n6731 gnd.n6729 9.3005
R9727 gnd.n6732 gnd.n166 9.3005
R9728 gnd.n7065 gnd.n6733 9.3005
R9729 gnd.n503 gnd.n388 9.3005
R9730 gnd.n6342 gnd.n505 9.3005
R9731 gnd.n6341 gnd.n506 9.3005
R9732 gnd.n265 gnd.n261 9.3005
R9733 gnd.n6579 gnd.n262 9.3005
R9734 gnd.n6578 gnd.n263 9.3005
R9735 gnd.n6577 gnd.n6573 9.3005
R9736 gnd.n6576 gnd.n6574 9.3005
R9737 gnd.n237 gnd.n234 9.3005
R9738 gnd.n6619 gnd.n235 9.3005
R9739 gnd.n6618 gnd.n6615 9.3005
R9740 gnd.n6617 gnd.n6616 9.3005
R9741 gnd.n219 gnd.n215 9.3005
R9742 gnd.n6643 gnd.n216 9.3005
R9743 gnd.n6642 gnd.n217 9.3005
R9744 gnd.n6641 gnd.n6637 9.3005
R9745 gnd.n6640 gnd.n6638 9.3005
R9746 gnd.n191 gnd.n190 9.3005
R9747 gnd.n6675 gnd.n6674 9.3005
R9748 gnd.n175 gnd.n174 9.3005
R9749 gnd.n6691 gnd.n6690 9.3005
R9750 gnd.n6692 gnd.n169 9.3005
R9751 gnd.n6698 gnd.n168 9.3005
R9752 gnd.n6700 gnd.n6699 9.3005
R9753 gnd.n6701 gnd.n89 9.3005
R9754 gnd.n7115 gnd.n90 9.3005
R9755 gnd.n7114 gnd.n91 9.3005
R9756 gnd.n7113 gnd.n92 9.3005
R9757 gnd.n6708 gnd.n93 9.3005
R9758 gnd.n7103 gnd.n109 9.3005
R9759 gnd.n7102 gnd.n110 9.3005
R9760 gnd.n7101 gnd.n111 9.3005
R9761 gnd.n6715 gnd.n112 9.3005
R9762 gnd.n7091 gnd.n128 9.3005
R9763 gnd.n7090 gnd.n129 9.3005
R9764 gnd.n7089 gnd.n130 9.3005
R9765 gnd.n6722 gnd.n131 9.3005
R9766 gnd.n7079 gnd.n147 9.3005
R9767 gnd.n7078 gnd.n148 9.3005
R9768 gnd.n7077 gnd.n149 9.3005
R9769 gnd.n6729 gnd.n150 9.3005
R9770 gnd.n7067 gnd.n166 9.3005
R9771 gnd.n7066 gnd.n7065 9.3005
R9772 gnd.n6343 gnd.n388 9.3005
R9773 gnd.n5491 gnd.n5490 9.3005
R9774 gnd.n5464 gnd.n5463 9.3005
R9775 gnd.n5485 gnd.n5484 9.3005
R9776 gnd.n5483 gnd.n5482 9.3005
R9777 gnd.n5468 gnd.n5467 9.3005
R9778 gnd.n5477 gnd.n5476 9.3005
R9779 gnd.n5475 gnd.n5474 9.3005
R9780 gnd.n5459 gnd.n5458 9.3005
R9781 gnd.n5432 gnd.n5431 9.3005
R9782 gnd.n5453 gnd.n5452 9.3005
R9783 gnd.n5451 gnd.n5450 9.3005
R9784 gnd.n5436 gnd.n5435 9.3005
R9785 gnd.n5445 gnd.n5444 9.3005
R9786 gnd.n5443 gnd.n5442 9.3005
R9787 gnd.n5427 gnd.n5426 9.3005
R9788 gnd.n5400 gnd.n5399 9.3005
R9789 gnd.n5421 gnd.n5420 9.3005
R9790 gnd.n5419 gnd.n5418 9.3005
R9791 gnd.n5404 gnd.n5403 9.3005
R9792 gnd.n5413 gnd.n5412 9.3005
R9793 gnd.n5411 gnd.n5410 9.3005
R9794 gnd.n5396 gnd.n5395 9.3005
R9795 gnd.n5369 gnd.n5368 9.3005
R9796 gnd.n5390 gnd.n5389 9.3005
R9797 gnd.n5388 gnd.n5387 9.3005
R9798 gnd.n5373 gnd.n5372 9.3005
R9799 gnd.n5382 gnd.n5381 9.3005
R9800 gnd.n5380 gnd.n5379 9.3005
R9801 gnd.n5364 gnd.n5363 9.3005
R9802 gnd.n5337 gnd.n5336 9.3005
R9803 gnd.n5358 gnd.n5357 9.3005
R9804 gnd.n5356 gnd.n5355 9.3005
R9805 gnd.n5341 gnd.n5340 9.3005
R9806 gnd.n5350 gnd.n5349 9.3005
R9807 gnd.n5348 gnd.n5347 9.3005
R9808 gnd.n5332 gnd.n5331 9.3005
R9809 gnd.n5305 gnd.n5304 9.3005
R9810 gnd.n5326 gnd.n5325 9.3005
R9811 gnd.n5324 gnd.n5323 9.3005
R9812 gnd.n5309 gnd.n5308 9.3005
R9813 gnd.n5318 gnd.n5317 9.3005
R9814 gnd.n5316 gnd.n5315 9.3005
R9815 gnd.n5300 gnd.n5299 9.3005
R9816 gnd.n5273 gnd.n5272 9.3005
R9817 gnd.n5294 gnd.n5293 9.3005
R9818 gnd.n5292 gnd.n5291 9.3005
R9819 gnd.n5277 gnd.n5276 9.3005
R9820 gnd.n5286 gnd.n5285 9.3005
R9821 gnd.n5284 gnd.n5283 9.3005
R9822 gnd.n5269 gnd.n5268 9.3005
R9823 gnd.n5242 gnd.n5241 9.3005
R9824 gnd.n5263 gnd.n5262 9.3005
R9825 gnd.n5261 gnd.n5260 9.3005
R9826 gnd.n5246 gnd.n5245 9.3005
R9827 gnd.n5255 gnd.n5254 9.3005
R9828 gnd.n5253 gnd.n5252 9.3005
R9829 gnd.n5617 gnd.n5616 9.3005
R9830 gnd.n5615 gnd.n4185 9.3005
R9831 gnd.n5614 gnd.n5613 9.3005
R9832 gnd.n5610 gnd.n4186 9.3005
R9833 gnd.n5607 gnd.n4187 9.3005
R9834 gnd.n5606 gnd.n4188 9.3005
R9835 gnd.n5603 gnd.n4189 9.3005
R9836 gnd.n5602 gnd.n4190 9.3005
R9837 gnd.n5599 gnd.n4191 9.3005
R9838 gnd.n5598 gnd.n4192 9.3005
R9839 gnd.n5595 gnd.n4193 9.3005
R9840 gnd.n5594 gnd.n4194 9.3005
R9841 gnd.n5591 gnd.n4195 9.3005
R9842 gnd.n5590 gnd.n4196 9.3005
R9843 gnd.n5587 gnd.n5586 9.3005
R9844 gnd.n5585 gnd.n4197 9.3005
R9845 gnd.n5618 gnd.n4184 9.3005
R9846 gnd.n4859 gnd.n4858 9.3005
R9847 gnd.n4563 gnd.n4562 9.3005
R9848 gnd.n4886 gnd.n4885 9.3005
R9849 gnd.n4887 gnd.n4561 9.3005
R9850 gnd.n4891 gnd.n4888 9.3005
R9851 gnd.n4890 gnd.n4889 9.3005
R9852 gnd.n4535 gnd.n4534 9.3005
R9853 gnd.n4916 gnd.n4915 9.3005
R9854 gnd.n4917 gnd.n4533 9.3005
R9855 gnd.n4919 gnd.n4918 9.3005
R9856 gnd.n4513 gnd.n4512 9.3005
R9857 gnd.n4947 gnd.n4946 9.3005
R9858 gnd.n4948 gnd.n4511 9.3005
R9859 gnd.n4956 gnd.n4949 9.3005
R9860 gnd.n4955 gnd.n4950 9.3005
R9861 gnd.n4954 gnd.n4952 9.3005
R9862 gnd.n4951 gnd.n4460 9.3005
R9863 gnd.n5004 gnd.n4461 9.3005
R9864 gnd.n5003 gnd.n4462 9.3005
R9865 gnd.n5002 gnd.n4463 9.3005
R9866 gnd.n4482 gnd.n4464 9.3005
R9867 gnd.n4484 gnd.n4483 9.3005
R9868 gnd.n4382 gnd.n4381 9.3005
R9869 gnd.n5042 gnd.n5041 9.3005
R9870 gnd.n5043 gnd.n4380 9.3005
R9871 gnd.n5047 gnd.n5044 9.3005
R9872 gnd.n5046 gnd.n5045 9.3005
R9873 gnd.n4355 gnd.n4354 9.3005
R9874 gnd.n5082 gnd.n5081 9.3005
R9875 gnd.n5083 gnd.n4353 9.3005
R9876 gnd.n5087 gnd.n5084 9.3005
R9877 gnd.n5086 gnd.n5085 9.3005
R9878 gnd.n4328 gnd.n4327 9.3005
R9879 gnd.n5127 gnd.n5126 9.3005
R9880 gnd.n5128 gnd.n4326 9.3005
R9881 gnd.n5132 gnd.n5129 9.3005
R9882 gnd.n5131 gnd.n5130 9.3005
R9883 gnd.n4300 gnd.n4299 9.3005
R9884 gnd.n5167 gnd.n5166 9.3005
R9885 gnd.n5168 gnd.n4298 9.3005
R9886 gnd.n5172 gnd.n5169 9.3005
R9887 gnd.n5171 gnd.n5170 9.3005
R9888 gnd.n4273 gnd.n4272 9.3005
R9889 gnd.n5216 gnd.n5215 9.3005
R9890 gnd.n5217 gnd.n4271 9.3005
R9891 gnd.n5221 gnd.n5218 9.3005
R9892 gnd.n5220 gnd.n5219 9.3005
R9893 gnd.n4246 gnd.n4245 9.3005
R9894 gnd.n5510 gnd.n5509 9.3005
R9895 gnd.n5511 gnd.n4244 9.3005
R9896 gnd.n5517 gnd.n5512 9.3005
R9897 gnd.n5516 gnd.n5513 9.3005
R9898 gnd.n5515 gnd.n5514 9.3005
R9899 gnd.n4860 gnd.n4857 9.3005
R9900 gnd.n4642 gnd.n4601 9.3005
R9901 gnd.n4637 gnd.n4636 9.3005
R9902 gnd.n4635 gnd.n4602 9.3005
R9903 gnd.n4634 gnd.n4633 9.3005
R9904 gnd.n4630 gnd.n4603 9.3005
R9905 gnd.n4627 gnd.n4626 9.3005
R9906 gnd.n4625 gnd.n4604 9.3005
R9907 gnd.n4624 gnd.n4623 9.3005
R9908 gnd.n4620 gnd.n4605 9.3005
R9909 gnd.n4617 gnd.n4616 9.3005
R9910 gnd.n4615 gnd.n4606 9.3005
R9911 gnd.n4614 gnd.n4613 9.3005
R9912 gnd.n4610 gnd.n4608 9.3005
R9913 gnd.n4607 gnd.n4587 9.3005
R9914 gnd.n4854 gnd.n4586 9.3005
R9915 gnd.n4856 gnd.n4855 9.3005
R9916 gnd.n4644 gnd.n4643 9.3005
R9917 gnd.n4867 gnd.n4573 9.3005
R9918 gnd.n4874 gnd.n4574 9.3005
R9919 gnd.n4876 gnd.n4875 9.3005
R9920 gnd.n4877 gnd.n4554 9.3005
R9921 gnd.n4896 gnd.n4895 9.3005
R9922 gnd.n4898 gnd.n4546 9.3005
R9923 gnd.n4905 gnd.n4548 9.3005
R9924 gnd.n4906 gnd.n4543 9.3005
R9925 gnd.n4908 gnd.n4907 9.3005
R9926 gnd.n4544 gnd.n4529 9.3005
R9927 gnd.n4924 gnd.n4527 9.3005
R9928 gnd.n4928 gnd.n4927 9.3005
R9929 gnd.n4926 gnd.n4503 9.3005
R9930 gnd.n4963 gnd.n4502 9.3005
R9931 gnd.n4966 gnd.n4965 9.3005
R9932 gnd.n4499 gnd.n4498 9.3005
R9933 gnd.n4972 gnd.n4500 9.3005
R9934 gnd.n4974 gnd.n4973 9.3005
R9935 gnd.n4976 gnd.n4497 9.3005
R9936 gnd.n4979 gnd.n4978 9.3005
R9937 gnd.n4982 gnd.n4980 9.3005
R9938 gnd.n4984 gnd.n4983 9.3005
R9939 gnd.n4990 gnd.n4985 9.3005
R9940 gnd.n4989 gnd.n4988 9.3005
R9941 gnd.n4373 gnd.n4372 9.3005
R9942 gnd.n5056 gnd.n5055 9.3005
R9943 gnd.n5057 gnd.n4366 9.3005
R9944 gnd.n5065 gnd.n4365 9.3005
R9945 gnd.n5068 gnd.n5067 9.3005
R9946 gnd.n5070 gnd.n5069 9.3005
R9947 gnd.n5073 gnd.n4348 9.3005
R9948 gnd.n5071 gnd.n4346 9.3005
R9949 gnd.n5093 gnd.n4344 9.3005
R9950 gnd.n5095 gnd.n5094 9.3005
R9951 gnd.n4318 gnd.n4317 9.3005
R9952 gnd.n5141 gnd.n5140 9.3005
R9953 gnd.n5142 gnd.n4311 9.3005
R9954 gnd.n5150 gnd.n4310 9.3005
R9955 gnd.n5153 gnd.n5152 9.3005
R9956 gnd.n5155 gnd.n5154 9.3005
R9957 gnd.n5158 gnd.n4293 9.3005
R9958 gnd.n5156 gnd.n4291 9.3005
R9959 gnd.n5178 gnd.n4289 9.3005
R9960 gnd.n5180 gnd.n5179 9.3005
R9961 gnd.n4264 gnd.n4263 9.3005
R9962 gnd.n5230 gnd.n5229 9.3005
R9963 gnd.n5231 gnd.n4257 9.3005
R9964 gnd.n5239 gnd.n4256 9.3005
R9965 gnd.n5498 gnd.n5497 9.3005
R9966 gnd.n5500 gnd.n5499 9.3005
R9967 gnd.n5501 gnd.n4237 9.3005
R9968 gnd.n5525 gnd.n5524 9.3005
R9969 gnd.n4238 gnd.n4200 9.3005
R9970 gnd.n4865 gnd.n4864 9.3005
R9971 gnd.n5581 gnd.n4201 9.3005
R9972 gnd.n5580 gnd.n4203 9.3005
R9973 gnd.n5577 gnd.n4204 9.3005
R9974 gnd.n5576 gnd.n4205 9.3005
R9975 gnd.n5573 gnd.n4206 9.3005
R9976 gnd.n5572 gnd.n4207 9.3005
R9977 gnd.n5569 gnd.n4208 9.3005
R9978 gnd.n5568 gnd.n4209 9.3005
R9979 gnd.n5565 gnd.n4210 9.3005
R9980 gnd.n5564 gnd.n4211 9.3005
R9981 gnd.n5561 gnd.n4212 9.3005
R9982 gnd.n5560 gnd.n4213 9.3005
R9983 gnd.n5557 gnd.n4214 9.3005
R9984 gnd.n5556 gnd.n4215 9.3005
R9985 gnd.n5553 gnd.n4216 9.3005
R9986 gnd.n5552 gnd.n4217 9.3005
R9987 gnd.n5549 gnd.n4218 9.3005
R9988 gnd.n5548 gnd.n4219 9.3005
R9989 gnd.n5545 gnd.n4220 9.3005
R9990 gnd.n5544 gnd.n4221 9.3005
R9991 gnd.n5541 gnd.n4222 9.3005
R9992 gnd.n5540 gnd.n4223 9.3005
R9993 gnd.n5537 gnd.n4227 9.3005
R9994 gnd.n5536 gnd.n4228 9.3005
R9995 gnd.n5533 gnd.n4229 9.3005
R9996 gnd.n5532 gnd.n4230 9.3005
R9997 gnd.n5583 gnd.n5582 9.3005
R9998 gnd.n5034 gnd.n5018 9.3005
R9999 gnd.n5033 gnd.n5019 9.3005
R10000 gnd.n5032 gnd.n5020 9.3005
R10001 gnd.n5030 gnd.n5021 9.3005
R10002 gnd.n5029 gnd.n5022 9.3005
R10003 gnd.n5027 gnd.n5023 9.3005
R10004 gnd.n5026 gnd.n5024 9.3005
R10005 gnd.n4336 gnd.n4335 9.3005
R10006 gnd.n5103 gnd.n5102 9.3005
R10007 gnd.n5104 gnd.n4334 9.3005
R10008 gnd.n5121 gnd.n5105 9.3005
R10009 gnd.n5120 gnd.n5106 9.3005
R10010 gnd.n5119 gnd.n5107 9.3005
R10011 gnd.n5117 gnd.n5108 9.3005
R10012 gnd.n5116 gnd.n5109 9.3005
R10013 gnd.n5114 gnd.n5110 9.3005
R10014 gnd.n5113 gnd.n5111 9.3005
R10015 gnd.n4280 gnd.n4279 9.3005
R10016 gnd.n5188 gnd.n5187 9.3005
R10017 gnd.n5189 gnd.n4278 9.3005
R10018 gnd.n5210 gnd.n5190 9.3005
R10019 gnd.n5209 gnd.n5191 9.3005
R10020 gnd.n5208 gnd.n5192 9.3005
R10021 gnd.n5205 gnd.n5193 9.3005
R10022 gnd.n5204 gnd.n5194 9.3005
R10023 gnd.n5202 gnd.n5195 9.3005
R10024 gnd.n5201 gnd.n5196 9.3005
R10025 gnd.n5199 gnd.n5198 9.3005
R10026 gnd.n5197 gnd.n4232 9.3005
R10027 gnd.n4775 gnd.n4774 9.3005
R10028 gnd.n4665 gnd.n4664 9.3005
R10029 gnd.n4789 gnd.n4788 9.3005
R10030 gnd.n4790 gnd.n4663 9.3005
R10031 gnd.n4792 gnd.n4791 9.3005
R10032 gnd.n4653 gnd.n4652 9.3005
R10033 gnd.n4805 gnd.n4804 9.3005
R10034 gnd.n4806 gnd.n4651 9.3005
R10035 gnd.n4838 gnd.n4807 9.3005
R10036 gnd.n4837 gnd.n4808 9.3005
R10037 gnd.n4836 gnd.n4809 9.3005
R10038 gnd.n4835 gnd.n4810 9.3005
R10039 gnd.n4832 gnd.n4811 9.3005
R10040 gnd.n4831 gnd.n4812 9.3005
R10041 gnd.n4830 gnd.n4813 9.3005
R10042 gnd.n4828 gnd.n4814 9.3005
R10043 gnd.n4827 gnd.n4815 9.3005
R10044 gnd.n4824 gnd.n4816 9.3005
R10045 gnd.n4823 gnd.n4817 9.3005
R10046 gnd.n4822 gnd.n4818 9.3005
R10047 gnd.n4820 gnd.n4819 9.3005
R10048 gnd.n4519 gnd.n4518 9.3005
R10049 gnd.n4936 gnd.n4935 9.3005
R10050 gnd.n4937 gnd.n4517 9.3005
R10051 gnd.n4941 gnd.n4938 9.3005
R10052 gnd.n4940 gnd.n4939 9.3005
R10053 gnd.n4441 gnd.n4440 9.3005
R10054 gnd.n5016 gnd.n5015 9.3005
R10055 gnd.n4773 gnd.n4674 9.3005
R10056 gnd.n4676 gnd.n4675 9.3005
R10057 gnd.n4720 gnd.n4718 9.3005
R10058 gnd.n4721 gnd.n4717 9.3005
R10059 gnd.n4724 gnd.n4713 9.3005
R10060 gnd.n4725 gnd.n4712 9.3005
R10061 gnd.n4728 gnd.n4711 9.3005
R10062 gnd.n4729 gnd.n4710 9.3005
R10063 gnd.n4732 gnd.n4709 9.3005
R10064 gnd.n4733 gnd.n4708 9.3005
R10065 gnd.n4736 gnd.n4707 9.3005
R10066 gnd.n4737 gnd.n4706 9.3005
R10067 gnd.n4740 gnd.n4705 9.3005
R10068 gnd.n4741 gnd.n4704 9.3005
R10069 gnd.n4744 gnd.n4703 9.3005
R10070 gnd.n4745 gnd.n4702 9.3005
R10071 gnd.n4748 gnd.n4701 9.3005
R10072 gnd.n4749 gnd.n4700 9.3005
R10073 gnd.n4752 gnd.n4699 9.3005
R10074 gnd.n4753 gnd.n4698 9.3005
R10075 gnd.n4756 gnd.n4697 9.3005
R10076 gnd.n4757 gnd.n4696 9.3005
R10077 gnd.n4760 gnd.n4695 9.3005
R10078 gnd.n4762 gnd.n4694 9.3005
R10079 gnd.n4763 gnd.n4693 9.3005
R10080 gnd.n4764 gnd.n4692 9.3005
R10081 gnd.n4765 gnd.n4691 9.3005
R10082 gnd.n4772 gnd.n4771 9.3005
R10083 gnd.n4781 gnd.n4780 9.3005
R10084 gnd.n4782 gnd.n4668 9.3005
R10085 gnd.n4784 gnd.n4783 9.3005
R10086 gnd.n4659 gnd.n4658 9.3005
R10087 gnd.n4797 gnd.n4796 9.3005
R10088 gnd.n4798 gnd.n4657 9.3005
R10089 gnd.n4800 gnd.n4799 9.3005
R10090 gnd.n4646 gnd.n4645 9.3005
R10091 gnd.n4843 gnd.n4842 9.3005
R10092 gnd.n4844 gnd.n4600 9.3005
R10093 gnd.n4848 gnd.n4846 9.3005
R10094 gnd.n4847 gnd.n4579 9.3005
R10095 gnd.n4866 gnd.n4578 9.3005
R10096 gnd.n4869 gnd.n4868 9.3005
R10097 gnd.n4572 gnd.n4571 9.3005
R10098 gnd.n4880 gnd.n4878 9.3005
R10099 gnd.n4879 gnd.n4553 9.3005
R10100 gnd.n4897 gnd.n4552 9.3005
R10101 gnd.n4900 gnd.n4899 9.3005
R10102 gnd.n4547 gnd.n4542 9.3005
R10103 gnd.n4910 gnd.n4909 9.3005
R10104 gnd.n4545 gnd.n4525 9.3005
R10105 gnd.n4931 gnd.n4526 9.3005
R10106 gnd.n4930 gnd.n4929 9.3005
R10107 gnd.n4528 gnd.n4504 9.3005
R10108 gnd.n4962 gnd.n4961 9.3005
R10109 gnd.n4964 gnd.n4449 9.3005
R10110 gnd.n5011 gnd.n4450 9.3005
R10111 gnd.n5010 gnd.n4451 9.3005
R10112 gnd.n5009 gnd.n4452 9.3005
R10113 gnd.n4975 gnd.n4453 9.3005
R10114 gnd.n4977 gnd.n4471 9.3005
R10115 gnd.n4997 gnd.n4472 9.3005
R10116 gnd.n4996 gnd.n4473 9.3005
R10117 gnd.n4995 gnd.n4474 9.3005
R10118 gnd.n4986 gnd.n4475 9.3005
R10119 gnd.n4987 gnd.n4374 9.3005
R10120 gnd.n5053 gnd.n5052 9.3005
R10121 gnd.n5054 gnd.n4367 9.3005
R10122 gnd.n5064 gnd.n5063 9.3005
R10123 gnd.n5066 gnd.n4363 9.3005
R10124 gnd.n5076 gnd.n4364 9.3005
R10125 gnd.n5075 gnd.n5074 9.3005
R10126 gnd.n5072 gnd.n4342 9.3005
R10127 gnd.n5098 gnd.n4343 9.3005
R10128 gnd.n5097 gnd.n5096 9.3005
R10129 gnd.n4345 gnd.n4319 9.3005
R10130 gnd.n5138 gnd.n5137 9.3005
R10131 gnd.n5139 gnd.n4312 9.3005
R10132 gnd.n5149 gnd.n5148 9.3005
R10133 gnd.n5151 gnd.n4308 9.3005
R10134 gnd.n5161 gnd.n4309 9.3005
R10135 gnd.n5160 gnd.n5159 9.3005
R10136 gnd.n5157 gnd.n4287 9.3005
R10137 gnd.n5183 gnd.n4288 9.3005
R10138 gnd.n5182 gnd.n5181 9.3005
R10139 gnd.n4290 gnd.n4265 9.3005
R10140 gnd.n5227 gnd.n5226 9.3005
R10141 gnd.n5228 gnd.n4258 9.3005
R10142 gnd.n5238 gnd.n5237 9.3005
R10143 gnd.n5496 gnd.n4254 9.3005
R10144 gnd.n5504 gnd.n4255 9.3005
R10145 gnd.n5503 gnd.n5502 9.3005
R10146 gnd.n4236 gnd.n4235 9.3005
R10147 gnd.n5527 gnd.n5526 9.3005
R10148 gnd.n4670 gnd.n4669 9.3005
R10149 gnd.n2408 gnd.n2297 9.3005
R10150 gnd.n2368 gnd.n2308 9.3005
R10151 gnd.n2371 gnd.n2369 9.3005
R10152 gnd.n2372 gnd.n2307 9.3005
R10153 gnd.n2375 gnd.n2374 9.3005
R10154 gnd.n2376 gnd.n2306 9.3005
R10155 gnd.n2379 gnd.n2377 9.3005
R10156 gnd.n2380 gnd.n2305 9.3005
R10157 gnd.n2383 gnd.n2382 9.3005
R10158 gnd.n2384 gnd.n2304 9.3005
R10159 gnd.n2387 gnd.n2385 9.3005
R10160 gnd.n2388 gnd.n2303 9.3005
R10161 gnd.n2391 gnd.n2390 9.3005
R10162 gnd.n2392 gnd.n2302 9.3005
R10163 gnd.n2395 gnd.n2393 9.3005
R10164 gnd.n2396 gnd.n2301 9.3005
R10165 gnd.n2399 gnd.n2398 9.3005
R10166 gnd.n2400 gnd.n2300 9.3005
R10167 gnd.n2403 gnd.n2401 9.3005
R10168 gnd.n2404 gnd.n2299 9.3005
R10169 gnd.n2407 gnd.n2406 9.3005
R10170 gnd.n2367 gnd.n2366 9.3005
R10171 gnd.n3870 gnd.n1405 9.3005
R10172 gnd.n3873 gnd.n1404 9.3005
R10173 gnd.n3874 gnd.n1403 9.3005
R10174 gnd.n3877 gnd.n1402 9.3005
R10175 gnd.n3878 gnd.n1401 9.3005
R10176 gnd.n3881 gnd.n1400 9.3005
R10177 gnd.n3882 gnd.n1399 9.3005
R10178 gnd.n3885 gnd.n1398 9.3005
R10179 gnd.n3887 gnd.n1395 9.3005
R10180 gnd.n3890 gnd.n1394 9.3005
R10181 gnd.n3891 gnd.n1393 9.3005
R10182 gnd.n3894 gnd.n1392 9.3005
R10183 gnd.n3895 gnd.n1391 9.3005
R10184 gnd.n3898 gnd.n1390 9.3005
R10185 gnd.n3899 gnd.n1389 9.3005
R10186 gnd.n3902 gnd.n1388 9.3005
R10187 gnd.n3903 gnd.n1387 9.3005
R10188 gnd.n3906 gnd.n1386 9.3005
R10189 gnd.n3907 gnd.n1385 9.3005
R10190 gnd.n3910 gnd.n1384 9.3005
R10191 gnd.n3911 gnd.n1383 9.3005
R10192 gnd.n3914 gnd.n1382 9.3005
R10193 gnd.n3915 gnd.n1381 9.3005
R10194 gnd.n3916 gnd.n1380 9.3005
R10195 gnd.n1337 gnd.n1336 9.3005
R10196 gnd.n3922 gnd.n3921 9.3005
R10197 gnd.n2174 gnd.n2172 9.3005
R10198 gnd.n2176 gnd.n2175 9.3005
R10199 gnd.n2179 gnd.n2169 9.3005
R10200 gnd.n2183 gnd.n2182 9.3005
R10201 gnd.n2184 gnd.n2168 9.3005
R10202 gnd.n2186 gnd.n2185 9.3005
R10203 gnd.n2189 gnd.n2167 9.3005
R10204 gnd.n2193 gnd.n2192 9.3005
R10205 gnd.n2194 gnd.n2166 9.3005
R10206 gnd.n2196 gnd.n2195 9.3005
R10207 gnd.n2199 gnd.n2163 9.3005
R10208 gnd.n2203 gnd.n2202 9.3005
R10209 gnd.n2204 gnd.n2162 9.3005
R10210 gnd.n2206 gnd.n2205 9.3005
R10211 gnd.n2209 gnd.n2161 9.3005
R10212 gnd.n2213 gnd.n2212 9.3005
R10213 gnd.n2214 gnd.n2160 9.3005
R10214 gnd.n2216 gnd.n2215 9.3005
R10215 gnd.n2219 gnd.n2159 9.3005
R10216 gnd.n2223 gnd.n2222 9.3005
R10217 gnd.n2224 gnd.n2158 9.3005
R10218 gnd.n2226 gnd.n2225 9.3005
R10219 gnd.n2229 gnd.n2157 9.3005
R10220 gnd.n2233 gnd.n2232 9.3005
R10221 gnd.n2234 gnd.n2156 9.3005
R10222 gnd.n2236 gnd.n2235 9.3005
R10223 gnd.n2239 gnd.n2155 9.3005
R10224 gnd.n2243 gnd.n2242 9.3005
R10225 gnd.n2244 gnd.n2154 9.3005
R10226 gnd.n2246 gnd.n2245 9.3005
R10227 gnd.n2173 gnd.n1406 9.3005
R10228 gnd.n3997 gnd.n1217 9.3005
R10229 gnd.n3996 gnd.n1218 9.3005
R10230 gnd.n3995 gnd.n1219 9.3005
R10231 gnd.n1236 gnd.n1220 9.3005
R10232 gnd.n3985 gnd.n1237 9.3005
R10233 gnd.n3984 gnd.n1238 9.3005
R10234 gnd.n3983 gnd.n1239 9.3005
R10235 gnd.n1255 gnd.n1240 9.3005
R10236 gnd.n3973 gnd.n1256 9.3005
R10237 gnd.n3972 gnd.n1257 9.3005
R10238 gnd.n3971 gnd.n1258 9.3005
R10239 gnd.n1274 gnd.n1259 9.3005
R10240 gnd.n3961 gnd.n1275 9.3005
R10241 gnd.n3960 gnd.n1276 9.3005
R10242 gnd.n3959 gnd.n1277 9.3005
R10243 gnd.n1293 gnd.n1278 9.3005
R10244 gnd.n3949 gnd.n1294 9.3005
R10245 gnd.n3948 gnd.n1295 9.3005
R10246 gnd.n3947 gnd.n1296 9.3005
R10247 gnd.n1314 gnd.n1297 9.3005
R10248 gnd.n3937 gnd.n1315 9.3005
R10249 gnd.n3936 gnd.n1316 9.3005
R10250 gnd.n3935 gnd.n1317 9.3005
R10251 gnd.n1334 gnd.n1318 9.3005
R10252 gnd.n3925 gnd.n1335 9.3005
R10253 gnd.n3924 gnd.n3923 9.3005
R10254 gnd.n4047 gnd.n4046 9.3005
R10255 gnd.n4045 gnd.n1141 9.3005
R10256 gnd.n4044 gnd.n4043 9.3005
R10257 gnd.n1144 gnd.n1143 9.3005
R10258 gnd.n4033 gnd.n1161 9.3005
R10259 gnd.n4032 gnd.n1162 9.3005
R10260 gnd.n4031 gnd.n1163 9.3005
R10261 gnd.n1178 gnd.n1164 9.3005
R10262 gnd.n4021 gnd.n1179 9.3005
R10263 gnd.n4020 gnd.n1180 9.3005
R10264 gnd.n4019 gnd.n1181 9.3005
R10265 gnd.n1198 gnd.n1182 9.3005
R10266 gnd.n4009 gnd.n1199 9.3005
R10267 gnd.n4008 gnd.n1200 9.3005
R10268 gnd.n4007 gnd.n1201 9.3005
R10269 gnd.n1216 gnd.n1202 9.3005
R10270 gnd.n1142 gnd.n1140 9.3005
R10271 gnd.n4057 gnd.n4056 9.3005
R10272 gnd.n4060 gnd.n1125 9.3005
R10273 gnd.n4061 gnd.n1124 9.3005
R10274 gnd.n4064 gnd.n1123 9.3005
R10275 gnd.n4065 gnd.n1122 9.3005
R10276 gnd.n4068 gnd.n1121 9.3005
R10277 gnd.n4069 gnd.n1120 9.3005
R10278 gnd.n4072 gnd.n1119 9.3005
R10279 gnd.n4073 gnd.n1118 9.3005
R10280 gnd.n4076 gnd.n1117 9.3005
R10281 gnd.n4077 gnd.n1116 9.3005
R10282 gnd.n4080 gnd.n1115 9.3005
R10283 gnd.n4081 gnd.n1114 9.3005
R10284 gnd.n4084 gnd.n1113 9.3005
R10285 gnd.n4085 gnd.n1112 9.3005
R10286 gnd.n4088 gnd.n1111 9.3005
R10287 gnd.n4089 gnd.n1110 9.3005
R10288 gnd.n4092 gnd.n1109 9.3005
R10289 gnd.n4093 gnd.n1108 9.3005
R10290 gnd.n4096 gnd.n1107 9.3005
R10291 gnd.n4100 gnd.n1103 9.3005
R10292 gnd.n4101 gnd.n1102 9.3005
R10293 gnd.n4104 gnd.n1101 9.3005
R10294 gnd.n4105 gnd.n1100 9.3005
R10295 gnd.n4108 gnd.n1099 9.3005
R10296 gnd.n4109 gnd.n1098 9.3005
R10297 gnd.n4112 gnd.n1097 9.3005
R10298 gnd.n4113 gnd.n1096 9.3005
R10299 gnd.n4116 gnd.n1095 9.3005
R10300 gnd.n4117 gnd.n1094 9.3005
R10301 gnd.n4120 gnd.n1093 9.3005
R10302 gnd.n4121 gnd.n1092 9.3005
R10303 gnd.n4124 gnd.n1091 9.3005
R10304 gnd.n4125 gnd.n1090 9.3005
R10305 gnd.n4128 gnd.n1089 9.3005
R10306 gnd.n4129 gnd.n1088 9.3005
R10307 gnd.n4132 gnd.n1087 9.3005
R10308 gnd.n4133 gnd.n1086 9.3005
R10309 gnd.n4136 gnd.n1085 9.3005
R10310 gnd.n4138 gnd.n1082 9.3005
R10311 gnd.n4141 gnd.n1081 9.3005
R10312 gnd.n4142 gnd.n1080 9.3005
R10313 gnd.n4145 gnd.n1079 9.3005
R10314 gnd.n4146 gnd.n1078 9.3005
R10315 gnd.n4149 gnd.n1077 9.3005
R10316 gnd.n4150 gnd.n1076 9.3005
R10317 gnd.n4153 gnd.n1075 9.3005
R10318 gnd.n4154 gnd.n1074 9.3005
R10319 gnd.n4157 gnd.n1073 9.3005
R10320 gnd.n4158 gnd.n1072 9.3005
R10321 gnd.n4161 gnd.n1071 9.3005
R10322 gnd.n4162 gnd.n1070 9.3005
R10323 gnd.n4165 gnd.n1069 9.3005
R10324 gnd.n4167 gnd.n1068 9.3005
R10325 gnd.n4168 gnd.n1067 9.3005
R10326 gnd.n4169 gnd.n1066 9.3005
R10327 gnd.n4170 gnd.n1065 9.3005
R10328 gnd.n4097 gnd.n1104 9.3005
R10329 gnd.n4055 gnd.n1126 9.3005
R10330 gnd.n2361 gnd.n2360 9.3005
R10331 gnd.n2359 gnd.n2313 9.3005
R10332 gnd.n2358 gnd.n2357 9.3005
R10333 gnd.n2354 gnd.n2316 9.3005
R10334 gnd.n2353 gnd.n2350 9.3005
R10335 gnd.n2349 gnd.n2317 9.3005
R10336 gnd.n2348 gnd.n2347 9.3005
R10337 gnd.n2344 gnd.n2318 9.3005
R10338 gnd.n2343 gnd.n2340 9.3005
R10339 gnd.n2339 gnd.n2319 9.3005
R10340 gnd.n2338 gnd.n2337 9.3005
R10341 gnd.n2334 gnd.n2320 9.3005
R10342 gnd.n2333 gnd.n2330 9.3005
R10343 gnd.n2329 gnd.n2321 9.3005
R10344 gnd.n2328 gnd.n2327 9.3005
R10345 gnd.n2324 gnd.n2322 9.3005
R10346 gnd.n2323 gnd.n1129 9.3005
R10347 gnd.n2362 gnd.n2309 9.3005
R10348 gnd.n2364 gnd.n2363 9.3005
R10349 gnd.n2433 gnd.n1131 9.3005
R10350 gnd.n2436 gnd.n2434 9.3005
R10351 gnd.n2437 gnd.n1152 9.3005
R10352 gnd.n2439 gnd.n1153 9.3005
R10353 gnd.n2440 gnd.n1154 9.3005
R10354 gnd.n2443 gnd.n2441 9.3005
R10355 gnd.n2444 gnd.n1170 9.3005
R10356 gnd.n2446 gnd.n1171 9.3005
R10357 gnd.n2447 gnd.n1172 9.3005
R10358 gnd.n2450 gnd.n2448 9.3005
R10359 gnd.n2451 gnd.n1188 9.3005
R10360 gnd.n2453 gnd.n1189 9.3005
R10361 gnd.n2454 gnd.n1190 9.3005
R10362 gnd.n2457 gnd.n2455 9.3005
R10363 gnd.n2458 gnd.n1208 9.3005
R10364 gnd.n2460 gnd.n1209 9.3005
R10365 gnd.n2461 gnd.n1210 9.3005
R10366 gnd.n2464 gnd.n2462 9.3005
R10367 gnd.n2465 gnd.n1226 9.3005
R10368 gnd.n2467 gnd.n1227 9.3005
R10369 gnd.n2468 gnd.n1228 9.3005
R10370 gnd.n2471 gnd.n2469 9.3005
R10371 gnd.n2472 gnd.n1246 9.3005
R10372 gnd.n2474 gnd.n1247 9.3005
R10373 gnd.n2475 gnd.n1248 9.3005
R10374 gnd.n2478 gnd.n2476 9.3005
R10375 gnd.n2479 gnd.n1264 9.3005
R10376 gnd.n2481 gnd.n1265 9.3005
R10377 gnd.n2482 gnd.n1266 9.3005
R10378 gnd.n2485 gnd.n2483 9.3005
R10379 gnd.n2486 gnd.n1284 9.3005
R10380 gnd.n2488 gnd.n1285 9.3005
R10381 gnd.n2489 gnd.n1286 9.3005
R10382 gnd.n2492 gnd.n2490 9.3005
R10383 gnd.n2493 gnd.n1304 9.3005
R10384 gnd.n2494 gnd.n1305 9.3005
R10385 gnd.n2284 gnd.n1306 9.3005
R10386 gnd.n2507 gnd.n2285 9.3005
R10387 gnd.n2508 gnd.n1325 9.3005
R10388 gnd.n2512 gnd.n1326 9.3005
R10389 gnd.n2511 gnd.n1327 9.3005
R10390 gnd.n2510 gnd.n2509 9.3005
R10391 gnd.n4053 gnd.n1130 9.3005
R10392 gnd.n1132 gnd.n1131 9.3005
R10393 gnd.n2434 gnd.n1151 9.3005
R10394 gnd.n4039 gnd.n1152 9.3005
R10395 gnd.n4038 gnd.n1153 9.3005
R10396 gnd.n4037 gnd.n1154 9.3005
R10397 gnd.n2441 gnd.n1155 9.3005
R10398 gnd.n4027 gnd.n1170 9.3005
R10399 gnd.n4026 gnd.n1171 9.3005
R10400 gnd.n4025 gnd.n1172 9.3005
R10401 gnd.n2448 gnd.n1173 9.3005
R10402 gnd.n4015 gnd.n1188 9.3005
R10403 gnd.n4014 gnd.n1189 9.3005
R10404 gnd.n4013 gnd.n1190 9.3005
R10405 gnd.n2455 gnd.n1191 9.3005
R10406 gnd.n4003 gnd.n1208 9.3005
R10407 gnd.n4002 gnd.n1209 9.3005
R10408 gnd.n4001 gnd.n1210 9.3005
R10409 gnd.n2462 gnd.n1211 9.3005
R10410 gnd.n3991 gnd.n1226 9.3005
R10411 gnd.n3990 gnd.n1227 9.3005
R10412 gnd.n3989 gnd.n1228 9.3005
R10413 gnd.n2469 gnd.n1229 9.3005
R10414 gnd.n3979 gnd.n1246 9.3005
R10415 gnd.n3978 gnd.n1247 9.3005
R10416 gnd.n3977 gnd.n1248 9.3005
R10417 gnd.n2476 gnd.n1249 9.3005
R10418 gnd.n3967 gnd.n1264 9.3005
R10419 gnd.n3966 gnd.n1265 9.3005
R10420 gnd.n3965 gnd.n1266 9.3005
R10421 gnd.n2483 gnd.n1267 9.3005
R10422 gnd.n3955 gnd.n1284 9.3005
R10423 gnd.n3954 gnd.n1285 9.3005
R10424 gnd.n3953 gnd.n1286 9.3005
R10425 gnd.n2490 gnd.n1287 9.3005
R10426 gnd.n3943 gnd.n1304 9.3005
R10427 gnd.n3942 gnd.n1305 9.3005
R10428 gnd.n3941 gnd.n1306 9.3005
R10429 gnd.n2285 gnd.n1307 9.3005
R10430 gnd.n3931 gnd.n1325 9.3005
R10431 gnd.n3930 gnd.n1326 9.3005
R10432 gnd.n3929 gnd.n1327 9.3005
R10433 gnd.n2509 gnd.n1328 9.3005
R10434 gnd.n4053 gnd.n4052 9.3005
R10435 gnd.n5793 gnd.n5792 9.3005
R10436 gnd.n5794 gnd.n837 9.3005
R10437 gnd.n5796 gnd.n5795 9.3005
R10438 gnd.n833 gnd.n832 9.3005
R10439 gnd.n5803 gnd.n5802 9.3005
R10440 gnd.n5804 gnd.n831 9.3005
R10441 gnd.n5806 gnd.n5805 9.3005
R10442 gnd.n827 gnd.n826 9.3005
R10443 gnd.n5813 gnd.n5812 9.3005
R10444 gnd.n5814 gnd.n825 9.3005
R10445 gnd.n5816 gnd.n5815 9.3005
R10446 gnd.n821 gnd.n820 9.3005
R10447 gnd.n5823 gnd.n5822 9.3005
R10448 gnd.n5824 gnd.n819 9.3005
R10449 gnd.n5826 gnd.n5825 9.3005
R10450 gnd.n815 gnd.n814 9.3005
R10451 gnd.n5833 gnd.n5832 9.3005
R10452 gnd.n5834 gnd.n813 9.3005
R10453 gnd.n5836 gnd.n5835 9.3005
R10454 gnd.n809 gnd.n808 9.3005
R10455 gnd.n5843 gnd.n5842 9.3005
R10456 gnd.n5844 gnd.n807 9.3005
R10457 gnd.n5846 gnd.n5845 9.3005
R10458 gnd.n803 gnd.n802 9.3005
R10459 gnd.n5853 gnd.n5852 9.3005
R10460 gnd.n5854 gnd.n801 9.3005
R10461 gnd.n5856 gnd.n5855 9.3005
R10462 gnd.n797 gnd.n796 9.3005
R10463 gnd.n5863 gnd.n5862 9.3005
R10464 gnd.n5864 gnd.n795 9.3005
R10465 gnd.n5866 gnd.n5865 9.3005
R10466 gnd.n791 gnd.n790 9.3005
R10467 gnd.n5873 gnd.n5872 9.3005
R10468 gnd.n5874 gnd.n789 9.3005
R10469 gnd.n5876 gnd.n5875 9.3005
R10470 gnd.n785 gnd.n784 9.3005
R10471 gnd.n5883 gnd.n5882 9.3005
R10472 gnd.n5884 gnd.n783 9.3005
R10473 gnd.n5886 gnd.n5885 9.3005
R10474 gnd.n779 gnd.n778 9.3005
R10475 gnd.n5893 gnd.n5892 9.3005
R10476 gnd.n5894 gnd.n777 9.3005
R10477 gnd.n5896 gnd.n5895 9.3005
R10478 gnd.n773 gnd.n772 9.3005
R10479 gnd.n5903 gnd.n5902 9.3005
R10480 gnd.n5904 gnd.n771 9.3005
R10481 gnd.n5906 gnd.n5905 9.3005
R10482 gnd.n767 gnd.n766 9.3005
R10483 gnd.n5913 gnd.n5912 9.3005
R10484 gnd.n5914 gnd.n765 9.3005
R10485 gnd.n5916 gnd.n5915 9.3005
R10486 gnd.n761 gnd.n760 9.3005
R10487 gnd.n5923 gnd.n5922 9.3005
R10488 gnd.n5924 gnd.n759 9.3005
R10489 gnd.n5926 gnd.n5925 9.3005
R10490 gnd.n755 gnd.n754 9.3005
R10491 gnd.n5933 gnd.n5932 9.3005
R10492 gnd.n5934 gnd.n753 9.3005
R10493 gnd.n5936 gnd.n5935 9.3005
R10494 gnd.n749 gnd.n748 9.3005
R10495 gnd.n5943 gnd.n5942 9.3005
R10496 gnd.n5944 gnd.n747 9.3005
R10497 gnd.n5946 gnd.n5945 9.3005
R10498 gnd.n743 gnd.n742 9.3005
R10499 gnd.n5953 gnd.n5952 9.3005
R10500 gnd.n5954 gnd.n741 9.3005
R10501 gnd.n5956 gnd.n5955 9.3005
R10502 gnd.n737 gnd.n736 9.3005
R10503 gnd.n5963 gnd.n5962 9.3005
R10504 gnd.n5964 gnd.n735 9.3005
R10505 gnd.n5966 gnd.n5965 9.3005
R10506 gnd.n731 gnd.n730 9.3005
R10507 gnd.n5973 gnd.n5972 9.3005
R10508 gnd.n5974 gnd.n729 9.3005
R10509 gnd.n5976 gnd.n5975 9.3005
R10510 gnd.n725 gnd.n724 9.3005
R10511 gnd.n5983 gnd.n5982 9.3005
R10512 gnd.n5984 gnd.n723 9.3005
R10513 gnd.n5986 gnd.n5985 9.3005
R10514 gnd.n719 gnd.n718 9.3005
R10515 gnd.n5993 gnd.n5992 9.3005
R10516 gnd.n5994 gnd.n717 9.3005
R10517 gnd.n5996 gnd.n5995 9.3005
R10518 gnd.n713 gnd.n712 9.3005
R10519 gnd.n6003 gnd.n6002 9.3005
R10520 gnd.n6004 gnd.n711 9.3005
R10521 gnd.n6006 gnd.n6005 9.3005
R10522 gnd.n707 gnd.n706 9.3005
R10523 gnd.n6013 gnd.n6012 9.3005
R10524 gnd.n6014 gnd.n705 9.3005
R10525 gnd.n6016 gnd.n6015 9.3005
R10526 gnd.n701 gnd.n700 9.3005
R10527 gnd.n6023 gnd.n6022 9.3005
R10528 gnd.n6024 gnd.n699 9.3005
R10529 gnd.n6026 gnd.n6025 9.3005
R10530 gnd.n695 gnd.n694 9.3005
R10531 gnd.n6033 gnd.n6032 9.3005
R10532 gnd.n6034 gnd.n693 9.3005
R10533 gnd.n6036 gnd.n6035 9.3005
R10534 gnd.n689 gnd.n688 9.3005
R10535 gnd.n6043 gnd.n6042 9.3005
R10536 gnd.n6044 gnd.n687 9.3005
R10537 gnd.n6046 gnd.n6045 9.3005
R10538 gnd.n683 gnd.n682 9.3005
R10539 gnd.n6053 gnd.n6052 9.3005
R10540 gnd.n6054 gnd.n681 9.3005
R10541 gnd.n6056 gnd.n6055 9.3005
R10542 gnd.n677 gnd.n676 9.3005
R10543 gnd.n6063 gnd.n6062 9.3005
R10544 gnd.n6064 gnd.n675 9.3005
R10545 gnd.n6066 gnd.n6065 9.3005
R10546 gnd.n671 gnd.n670 9.3005
R10547 gnd.n6073 gnd.n6072 9.3005
R10548 gnd.n6074 gnd.n669 9.3005
R10549 gnd.n6076 gnd.n6075 9.3005
R10550 gnd.n665 gnd.n664 9.3005
R10551 gnd.n6083 gnd.n6082 9.3005
R10552 gnd.n6084 gnd.n663 9.3005
R10553 gnd.n6086 gnd.n6085 9.3005
R10554 gnd.n659 gnd.n658 9.3005
R10555 gnd.n6093 gnd.n6092 9.3005
R10556 gnd.n6094 gnd.n657 9.3005
R10557 gnd.n6096 gnd.n6095 9.3005
R10558 gnd.n653 gnd.n652 9.3005
R10559 gnd.n6103 gnd.n6102 9.3005
R10560 gnd.n6104 gnd.n651 9.3005
R10561 gnd.n6106 gnd.n6105 9.3005
R10562 gnd.n647 gnd.n646 9.3005
R10563 gnd.n6113 gnd.n6112 9.3005
R10564 gnd.n6116 gnd.n6115 9.3005
R10565 gnd.n641 gnd.n640 9.3005
R10566 gnd.n6123 gnd.n6122 9.3005
R10567 gnd.n6124 gnd.n639 9.3005
R10568 gnd.n6126 gnd.n6125 9.3005
R10569 gnd.n635 gnd.n634 9.3005
R10570 gnd.n6133 gnd.n6132 9.3005
R10571 gnd.n6134 gnd.n633 9.3005
R10572 gnd.n6136 gnd.n6135 9.3005
R10573 gnd.n629 gnd.n628 9.3005
R10574 gnd.n6143 gnd.n6142 9.3005
R10575 gnd.n6144 gnd.n627 9.3005
R10576 gnd.n6146 gnd.n6145 9.3005
R10577 gnd.n623 gnd.n622 9.3005
R10578 gnd.n6153 gnd.n6152 9.3005
R10579 gnd.n6154 gnd.n621 9.3005
R10580 gnd.n6156 gnd.n6155 9.3005
R10581 gnd.n617 gnd.n616 9.3005
R10582 gnd.n6163 gnd.n6162 9.3005
R10583 gnd.n6164 gnd.n615 9.3005
R10584 gnd.n6166 gnd.n6165 9.3005
R10585 gnd.n611 gnd.n610 9.3005
R10586 gnd.n6173 gnd.n6172 9.3005
R10587 gnd.n6174 gnd.n609 9.3005
R10588 gnd.n6176 gnd.n6175 9.3005
R10589 gnd.n605 gnd.n604 9.3005
R10590 gnd.n6183 gnd.n6182 9.3005
R10591 gnd.n6184 gnd.n603 9.3005
R10592 gnd.n6186 gnd.n6185 9.3005
R10593 gnd.n599 gnd.n598 9.3005
R10594 gnd.n6193 gnd.n6192 9.3005
R10595 gnd.n6194 gnd.n597 9.3005
R10596 gnd.n6196 gnd.n6195 9.3005
R10597 gnd.n593 gnd.n592 9.3005
R10598 gnd.n6203 gnd.n6202 9.3005
R10599 gnd.n6204 gnd.n591 9.3005
R10600 gnd.n6206 gnd.n6205 9.3005
R10601 gnd.n587 gnd.n586 9.3005
R10602 gnd.n6213 gnd.n6212 9.3005
R10603 gnd.n6214 gnd.n585 9.3005
R10604 gnd.n6216 gnd.n6215 9.3005
R10605 gnd.n581 gnd.n580 9.3005
R10606 gnd.n6223 gnd.n6222 9.3005
R10607 gnd.n6224 gnd.n579 9.3005
R10608 gnd.n6226 gnd.n6225 9.3005
R10609 gnd.n575 gnd.n574 9.3005
R10610 gnd.n6233 gnd.n6232 9.3005
R10611 gnd.n6234 gnd.n573 9.3005
R10612 gnd.n6236 gnd.n6235 9.3005
R10613 gnd.n569 gnd.n568 9.3005
R10614 gnd.n6243 gnd.n6242 9.3005
R10615 gnd.n6244 gnd.n567 9.3005
R10616 gnd.n6246 gnd.n6245 9.3005
R10617 gnd.n563 gnd.n562 9.3005
R10618 gnd.n6253 gnd.n6252 9.3005
R10619 gnd.n6254 gnd.n561 9.3005
R10620 gnd.n6256 gnd.n6255 9.3005
R10621 gnd.n557 gnd.n556 9.3005
R10622 gnd.n6263 gnd.n6262 9.3005
R10623 gnd.n6264 gnd.n555 9.3005
R10624 gnd.n6266 gnd.n6265 9.3005
R10625 gnd.n551 gnd.n550 9.3005
R10626 gnd.n6273 gnd.n6272 9.3005
R10627 gnd.n6274 gnd.n549 9.3005
R10628 gnd.n6276 gnd.n6275 9.3005
R10629 gnd.n545 gnd.n544 9.3005
R10630 gnd.n6283 gnd.n6282 9.3005
R10631 gnd.n6284 gnd.n543 9.3005
R10632 gnd.n6286 gnd.n6285 9.3005
R10633 gnd.n539 gnd.n538 9.3005
R10634 gnd.n6293 gnd.n6292 9.3005
R10635 gnd.n6294 gnd.n537 9.3005
R10636 gnd.n6296 gnd.n6295 9.3005
R10637 gnd.n533 gnd.n532 9.3005
R10638 gnd.n6303 gnd.n6302 9.3005
R10639 gnd.n6304 gnd.n531 9.3005
R10640 gnd.n6306 gnd.n6305 9.3005
R10641 gnd.n527 gnd.n526 9.3005
R10642 gnd.n6313 gnd.n6312 9.3005
R10643 gnd.n6314 gnd.n525 9.3005
R10644 gnd.n6318 gnd.n6315 9.3005
R10645 gnd.n6317 gnd.n6316 9.3005
R10646 gnd.n521 gnd.n520 9.3005
R10647 gnd.n6327 gnd.n6326 9.3005
R10648 gnd.n6114 gnd.n645 9.3005
R10649 gnd.n2523 gnd.n2522 9.3005
R10650 gnd.n2517 gnd.n2516 9.3005
R10651 gnd.n2528 gnd.n2527 9.3005
R10652 gnd.n2529 gnd.n2515 9.3005
R10653 gnd.n2532 gnd.n2531 9.3005
R10654 gnd.n2530 gnd.n2251 9.3005
R10655 gnd.n2564 gnd.n2252 9.3005
R10656 gnd.n2563 gnd.n2253 9.3005
R10657 gnd.n2562 gnd.n2254 9.3005
R10658 gnd.n2548 gnd.n2255 9.3005
R10659 gnd.n2549 gnd.n2547 9.3005
R10660 gnd.n2553 gnd.n2550 9.3005
R10661 gnd.n2552 gnd.n2551 9.3005
R10662 gnd.n2069 gnd.n2068 9.3005
R10663 gnd.n2648 gnd.n2647 9.3005
R10664 gnd.n2649 gnd.n2067 9.3005
R10665 gnd.n2653 gnd.n2650 9.3005
R10666 gnd.n2652 gnd.n2651 9.3005
R10667 gnd.n2044 gnd.n2043 9.3005
R10668 gnd.n2678 gnd.n2677 9.3005
R10669 gnd.n2679 gnd.n2042 9.3005
R10670 gnd.n2683 gnd.n2680 9.3005
R10671 gnd.n2682 gnd.n2681 9.3005
R10672 gnd.n2019 gnd.n2018 9.3005
R10673 gnd.n2708 gnd.n2707 9.3005
R10674 gnd.n2709 gnd.n2017 9.3005
R10675 gnd.n2713 gnd.n2710 9.3005
R10676 gnd.n2712 gnd.n2711 9.3005
R10677 gnd.n1994 gnd.n1993 9.3005
R10678 gnd.n2742 gnd.n2741 9.3005
R10679 gnd.n2743 gnd.n1992 9.3005
R10680 gnd.n2760 gnd.n2744 9.3005
R10681 gnd.n2759 gnd.n2745 9.3005
R10682 gnd.n2758 gnd.n2746 9.3005
R10683 gnd.n2749 gnd.n2747 9.3005
R10684 gnd.n2753 gnd.n2750 9.3005
R10685 gnd.n2752 gnd.n2751 9.3005
R10686 gnd.n1963 gnd.n1962 9.3005
R10687 gnd.n2916 gnd.n2915 9.3005
R10688 gnd.n2917 gnd.n1961 9.3005
R10689 gnd.n2921 gnd.n2918 9.3005
R10690 gnd.n2920 gnd.n2919 9.3005
R10691 gnd.n1936 gnd.n1935 9.3005
R10692 gnd.n2953 gnd.n2952 9.3005
R10693 gnd.n2954 gnd.n1934 9.3005
R10694 gnd.n2956 gnd.n2955 9.3005
R10695 gnd.n1915 gnd.n1914 9.3005
R10696 gnd.n2983 gnd.n2982 9.3005
R10697 gnd.n2984 gnd.n1913 9.3005
R10698 gnd.n2988 gnd.n2985 9.3005
R10699 gnd.n2987 gnd.n2986 9.3005
R10700 gnd.n1885 gnd.n1884 9.3005
R10701 gnd.n3034 gnd.n3033 9.3005
R10702 gnd.n3035 gnd.n1883 9.3005
R10703 gnd.n3039 gnd.n3036 9.3005
R10704 gnd.n3038 gnd.n3037 9.3005
R10705 gnd.n1866 gnd.n1865 9.3005
R10706 gnd.n3062 gnd.n3061 9.3005
R10707 gnd.n3063 gnd.n1864 9.3005
R10708 gnd.n3065 gnd.n3064 9.3005
R10709 gnd.n1838 gnd.n1837 9.3005
R10710 gnd.n3118 gnd.n3117 9.3005
R10711 gnd.n3119 gnd.n1836 9.3005
R10712 gnd.n3121 gnd.n3120 9.3005
R10713 gnd.n1815 gnd.n1814 9.3005
R10714 gnd.n3158 gnd.n3157 9.3005
R10715 gnd.n3159 gnd.n1813 9.3005
R10716 gnd.n3161 gnd.n3160 9.3005
R10717 gnd.n1792 gnd.n1791 9.3005
R10718 gnd.n3198 gnd.n3197 9.3005
R10719 gnd.n3199 gnd.n1790 9.3005
R10720 gnd.n3201 gnd.n3200 9.3005
R10721 gnd.n1770 gnd.n1769 9.3005
R10722 gnd.n3245 gnd.n3244 9.3005
R10723 gnd.n3246 gnd.n1768 9.3005
R10724 gnd.n3248 gnd.n3247 9.3005
R10725 gnd.n1752 gnd.n1751 9.3005
R10726 gnd.n3272 gnd.n3271 9.3005
R10727 gnd.n3273 gnd.n1750 9.3005
R10728 gnd.n3280 gnd.n3274 9.3005
R10729 gnd.n3279 gnd.n3275 9.3005
R10730 gnd.n3278 gnd.n3276 9.3005
R10731 gnd.n1716 gnd.n1715 9.3005
R10732 gnd.n3339 gnd.n3338 9.3005
R10733 gnd.n3340 gnd.n1714 9.3005
R10734 gnd.n3344 gnd.n3341 9.3005
R10735 gnd.n3343 gnd.n3342 9.3005
R10736 gnd.n1689 gnd.n1688 9.3005
R10737 gnd.n3390 gnd.n3389 9.3005
R10738 gnd.n3391 gnd.n1687 9.3005
R10739 gnd.n3398 gnd.n3392 9.3005
R10740 gnd.n3397 gnd.n3393 9.3005
R10741 gnd.n3396 gnd.n3394 9.3005
R10742 gnd.n1628 gnd.n1627 9.3005
R10743 gnd.n3578 gnd.n3577 9.3005
R10744 gnd.n3579 gnd.n1626 9.3005
R10745 gnd.n3581 gnd.n3580 9.3005
R10746 gnd.n1617 gnd.n1616 9.3005
R10747 gnd.n3600 gnd.n3599 9.3005
R10748 gnd.n3601 gnd.n1615 9.3005
R10749 gnd.n3603 gnd.n3602 9.3005
R10750 gnd.n1605 gnd.n1604 9.3005
R10751 gnd.n3621 gnd.n3620 9.3005
R10752 gnd.n3622 gnd.n1603 9.3005
R10753 gnd.n3624 gnd.n3623 9.3005
R10754 gnd.n1593 gnd.n1592 9.3005
R10755 gnd.n3642 gnd.n3641 9.3005
R10756 gnd.n3643 gnd.n1591 9.3005
R10757 gnd.n3645 gnd.n3644 9.3005
R10758 gnd.n1580 gnd.n1579 9.3005
R10759 gnd.n3663 gnd.n3662 9.3005
R10760 gnd.n3664 gnd.n1578 9.3005
R10761 gnd.n3672 gnd.n3665 9.3005
R10762 gnd.n3671 gnd.n3666 9.3005
R10763 gnd.n3670 gnd.n3668 9.3005
R10764 gnd.n3667 gnd.n493 9.3005
R10765 gnd.n6352 gnd.n494 9.3005
R10766 gnd.n6351 gnd.n495 9.3005
R10767 gnd.n6350 gnd.n496 9.3005
R10768 gnd.n509 gnd.n497 9.3005
R10769 gnd.n510 gnd.n499 9.3005
R10770 gnd.n511 gnd.n508 9.3005
R10771 gnd.n6336 gnd.n512 9.3005
R10772 gnd.n6335 gnd.n513 9.3005
R10773 gnd.n6334 gnd.n514 9.3005
R10774 gnd.n518 gnd.n515 9.3005
R10775 gnd.n6330 gnd.n519 9.3005
R10776 gnd.n6329 gnd.n6328 9.3005
R10777 gnd.n2521 gnd.n2519 9.3005
R10778 gnd.n5624 gnd.n1005 9.3005
R10779 gnd.n5625 gnd.n1004 9.3005
R10780 gnd.n5626 gnd.n1003 9.3005
R10781 gnd.n1002 gnd.n998 9.3005
R10782 gnd.n5632 gnd.n997 9.3005
R10783 gnd.n5633 gnd.n996 9.3005
R10784 gnd.n5634 gnd.n995 9.3005
R10785 gnd.n994 gnd.n990 9.3005
R10786 gnd.n5640 gnd.n989 9.3005
R10787 gnd.n5641 gnd.n988 9.3005
R10788 gnd.n5642 gnd.n987 9.3005
R10789 gnd.n986 gnd.n982 9.3005
R10790 gnd.n5648 gnd.n981 9.3005
R10791 gnd.n5649 gnd.n980 9.3005
R10792 gnd.n5650 gnd.n979 9.3005
R10793 gnd.n978 gnd.n974 9.3005
R10794 gnd.n5656 gnd.n973 9.3005
R10795 gnd.n5657 gnd.n972 9.3005
R10796 gnd.n5658 gnd.n971 9.3005
R10797 gnd.n970 gnd.n966 9.3005
R10798 gnd.n5664 gnd.n965 9.3005
R10799 gnd.n5665 gnd.n964 9.3005
R10800 gnd.n5666 gnd.n963 9.3005
R10801 gnd.n962 gnd.n958 9.3005
R10802 gnd.n5672 gnd.n957 9.3005
R10803 gnd.n5673 gnd.n956 9.3005
R10804 gnd.n5674 gnd.n955 9.3005
R10805 gnd.n954 gnd.n950 9.3005
R10806 gnd.n5680 gnd.n949 9.3005
R10807 gnd.n5681 gnd.n948 9.3005
R10808 gnd.n5682 gnd.n947 9.3005
R10809 gnd.n946 gnd.n942 9.3005
R10810 gnd.n5688 gnd.n941 9.3005
R10811 gnd.n5689 gnd.n940 9.3005
R10812 gnd.n5690 gnd.n939 9.3005
R10813 gnd.n938 gnd.n934 9.3005
R10814 gnd.n5696 gnd.n933 9.3005
R10815 gnd.n5697 gnd.n932 9.3005
R10816 gnd.n5698 gnd.n931 9.3005
R10817 gnd.n930 gnd.n926 9.3005
R10818 gnd.n5704 gnd.n925 9.3005
R10819 gnd.n5705 gnd.n924 9.3005
R10820 gnd.n5706 gnd.n923 9.3005
R10821 gnd.n922 gnd.n918 9.3005
R10822 gnd.n5712 gnd.n917 9.3005
R10823 gnd.n5713 gnd.n916 9.3005
R10824 gnd.n5714 gnd.n915 9.3005
R10825 gnd.n914 gnd.n910 9.3005
R10826 gnd.n5720 gnd.n909 9.3005
R10827 gnd.n5721 gnd.n908 9.3005
R10828 gnd.n5722 gnd.n907 9.3005
R10829 gnd.n906 gnd.n902 9.3005
R10830 gnd.n5728 gnd.n901 9.3005
R10831 gnd.n5729 gnd.n900 9.3005
R10832 gnd.n5730 gnd.n899 9.3005
R10833 gnd.n898 gnd.n894 9.3005
R10834 gnd.n5736 gnd.n893 9.3005
R10835 gnd.n5737 gnd.n892 9.3005
R10836 gnd.n5738 gnd.n891 9.3005
R10837 gnd.n890 gnd.n886 9.3005
R10838 gnd.n5744 gnd.n885 9.3005
R10839 gnd.n5745 gnd.n884 9.3005
R10840 gnd.n5746 gnd.n883 9.3005
R10841 gnd.n882 gnd.n878 9.3005
R10842 gnd.n5752 gnd.n877 9.3005
R10843 gnd.n5753 gnd.n876 9.3005
R10844 gnd.n5754 gnd.n875 9.3005
R10845 gnd.n874 gnd.n870 9.3005
R10846 gnd.n5760 gnd.n869 9.3005
R10847 gnd.n5761 gnd.n868 9.3005
R10848 gnd.n5762 gnd.n867 9.3005
R10849 gnd.n866 gnd.n862 9.3005
R10850 gnd.n5768 gnd.n861 9.3005
R10851 gnd.n5769 gnd.n860 9.3005
R10852 gnd.n5770 gnd.n859 9.3005
R10853 gnd.n858 gnd.n854 9.3005
R10854 gnd.n5776 gnd.n853 9.3005
R10855 gnd.n5777 gnd.n852 9.3005
R10856 gnd.n5778 gnd.n851 9.3005
R10857 gnd.n850 gnd.n846 9.3005
R10858 gnd.n5784 gnd.n845 9.3005
R10859 gnd.n5785 gnd.n844 9.3005
R10860 gnd.n5786 gnd.n843 9.3005
R10861 gnd.n842 gnd.n838 9.3005
R10862 gnd.n2520 gnd.n1006 9.3005
R10863 gnd.n6375 gnd.n452 9.3005
R10864 gnd.n2639 gnd.n2073 9.3005
R10865 gnd.n2642 gnd.n2641 9.3005
R10866 gnd.n2640 gnd.n2074 9.3005
R10867 gnd.n2051 gnd.n2050 9.3005
R10868 gnd.n2668 gnd.n2667 9.3005
R10869 gnd.n2669 gnd.n2048 9.3005
R10870 gnd.n2672 gnd.n2671 9.3005
R10871 gnd.n2670 gnd.n2049 9.3005
R10872 gnd.n2025 gnd.n2024 9.3005
R10873 gnd.n2698 gnd.n2697 9.3005
R10874 gnd.n2699 gnd.n2022 9.3005
R10875 gnd.n2702 gnd.n2701 9.3005
R10876 gnd.n2700 gnd.n2023 9.3005
R10877 gnd.n2001 gnd.n2000 9.3005
R10878 gnd.n2728 gnd.n2727 9.3005
R10879 gnd.n2729 gnd.n1998 9.3005
R10880 gnd.n2736 gnd.n2735 9.3005
R10881 gnd.n2734 gnd.n1999 9.3005
R10882 gnd.n2733 gnd.n2732 9.3005
R10883 gnd.n2731 gnd.n1978 9.3005
R10884 gnd.n2730 gnd.n1976 9.3005
R10885 gnd.n2896 gnd.n1975 9.3005
R10886 gnd.n2898 gnd.n2897 9.3005
R10887 gnd.n2899 gnd.n1973 9.3005
R10888 gnd.n2902 gnd.n2901 9.3005
R10889 gnd.n2900 gnd.n1974 9.3005
R10890 gnd.n1949 gnd.n1948 9.3005
R10891 gnd.n2935 gnd.n2934 9.3005
R10892 gnd.n2936 gnd.n1947 9.3005
R10893 gnd.n2938 gnd.n2937 9.3005
R10894 gnd.n1930 gnd.n1929 9.3005
R10895 gnd.n2964 gnd.n2963 9.3005
R10896 gnd.n2965 gnd.n1927 9.3005
R10897 gnd.n2968 gnd.n2967 9.3005
R10898 gnd.n2966 gnd.n1928 9.3005
R10899 gnd.n1901 gnd.n1900 9.3005
R10900 gnd.n3003 gnd.n3002 9.3005
R10901 gnd.n3004 gnd.n1898 9.3005
R10902 gnd.n3021 gnd.n3020 9.3005
R10903 gnd.n3019 gnd.n1899 9.3005
R10904 gnd.n3018 gnd.n3017 9.3005
R10905 gnd.n3016 gnd.n3005 9.3005
R10906 gnd.n3015 gnd.n3014 9.3005
R10907 gnd.n3013 gnd.n3009 9.3005
R10908 gnd.n3012 gnd.n3011 9.3005
R10909 gnd.n3010 gnd.n1853 9.3005
R10910 gnd.n3086 gnd.n1852 9.3005
R10911 gnd.n3088 gnd.n3087 9.3005
R10912 gnd.n3089 gnd.n1851 9.3005
R10913 gnd.n3091 gnd.n3090 9.3005
R10914 gnd.n1830 gnd.n1828 9.3005
R10915 gnd.n3141 gnd.n3140 9.3005
R10916 gnd.n3139 gnd.n1829 9.3005
R10917 gnd.n3138 gnd.n3137 9.3005
R10918 gnd.n1807 gnd.n1805 9.3005
R10919 gnd.n3181 gnd.n3180 9.3005
R10920 gnd.n3179 gnd.n1806 9.3005
R10921 gnd.n3178 gnd.n3177 9.3005
R10922 gnd.n1784 gnd.n1782 9.3005
R10923 gnd.n3230 gnd.n3229 9.3005
R10924 gnd.n3228 gnd.n1783 9.3005
R10925 gnd.n3227 gnd.n3226 9.3005
R10926 gnd.n3225 gnd.n1785 9.3005
R10927 gnd.n3224 gnd.n3223 9.3005
R10928 gnd.n3222 gnd.n3221 9.3005
R10929 gnd.n1734 gnd.n1733 9.3005
R10930 gnd.n3296 gnd.n3295 9.3005
R10931 gnd.n3297 gnd.n1731 9.3005
R10932 gnd.n3300 gnd.n3299 9.3005
R10933 gnd.n3298 gnd.n1732 9.3005
R10934 gnd.n1708 gnd.n1707 9.3005
R10935 gnd.n3351 gnd.n3350 9.3005
R10936 gnd.n3352 gnd.n1705 9.3005
R10937 gnd.n3363 gnd.n3362 9.3005
R10938 gnd.n3361 gnd.n1706 9.3005
R10939 gnd.n3360 gnd.n3359 9.3005
R10940 gnd.n3358 gnd.n3353 9.3005
R10941 gnd.n3357 gnd.n3356 9.3005
R10942 gnd.n1634 gnd.n1633 9.3005
R10943 gnd.n3568 gnd.n3567 9.3005
R10944 gnd.n3569 gnd.n1632 9.3005
R10945 gnd.n3571 gnd.n3570 9.3005
R10946 gnd.n1622 gnd.n1621 9.3005
R10947 gnd.n3590 gnd.n3589 9.3005
R10948 gnd.n3591 gnd.n1620 9.3005
R10949 gnd.n3593 gnd.n3592 9.3005
R10950 gnd.n1611 gnd.n1610 9.3005
R10951 gnd.n3611 gnd.n3610 9.3005
R10952 gnd.n3612 gnd.n1609 9.3005
R10953 gnd.n3614 gnd.n3613 9.3005
R10954 gnd.n1599 gnd.n1598 9.3005
R10955 gnd.n3632 gnd.n3631 9.3005
R10956 gnd.n3633 gnd.n1597 9.3005
R10957 gnd.n3635 gnd.n3634 9.3005
R10958 gnd.n1587 gnd.n1586 9.3005
R10959 gnd.n3653 gnd.n3652 9.3005
R10960 gnd.n3654 gnd.n1584 9.3005
R10961 gnd.n3657 gnd.n3656 9.3005
R10962 gnd.n3655 gnd.n1585 9.3005
R10963 gnd.n454 gnd.n453 9.3005
R10964 gnd.n6374 gnd.n6373 9.3005
R10965 gnd.n2638 gnd.n2637 9.3005
R10966 gnd.n2281 gnd.n2075 9.3005
R10967 gnd.n2410 gnd.n2409 9.3005
R10968 gnd.n2411 gnd.n2296 9.3005
R10969 gnd.n2414 gnd.n2413 9.3005
R10970 gnd.n2415 gnd.n2294 9.3005
R10971 gnd.n2417 gnd.n2416 9.3005
R10972 gnd.n2418 gnd.n2293 9.3005
R10973 gnd.n2421 gnd.n2420 9.3005
R10974 gnd.n2422 gnd.n2291 9.3005
R10975 gnd.n2424 gnd.n2423 9.3005
R10976 gnd.n2425 gnd.n2290 9.3005
R10977 gnd.n2428 gnd.n2427 9.3005
R10978 gnd.n2429 gnd.n2288 9.3005
R10979 gnd.n2431 gnd.n2430 9.3005
R10980 gnd.n2432 gnd.n2287 9.3005
R10981 gnd.n2499 gnd.n2498 9.3005
R10982 gnd.n2500 gnd.n2286 9.3005
R10983 gnd.n2503 gnd.n2502 9.3005
R10984 gnd.n2501 gnd.n2283 9.3005
R10985 gnd.n2537 gnd.n2282 9.3005
R10986 gnd.n2539 gnd.n2538 9.3005
R10987 gnd.n2540 gnd.n2151 9.3005
R10988 gnd.n2613 gnd.n2612 9.3005
R10989 gnd.n2611 gnd.n2610 9.3005
R10990 gnd.n2102 gnd.n2101 9.3005
R10991 gnd.n2605 gnd.n2604 9.3005
R10992 gnd.n2603 gnd.n2602 9.3005
R10993 gnd.n2110 gnd.n2109 9.3005
R10994 gnd.n2597 gnd.n2596 9.3005
R10995 gnd.n2595 gnd.n2594 9.3005
R10996 gnd.n2120 gnd.n2119 9.3005
R10997 gnd.n2589 gnd.n2588 9.3005
R10998 gnd.n2587 gnd.n2586 9.3005
R10999 gnd.n2128 gnd.n2127 9.3005
R11000 gnd.n2581 gnd.n2580 9.3005
R11001 gnd.n2579 gnd.n2578 9.3005
R11002 gnd.n2138 gnd.n2137 9.3005
R11003 gnd.n2573 gnd.n2572 9.3005
R11004 gnd.n2571 gnd.n2148 9.3005
R11005 gnd.n2570 gnd.n2150 9.3005
R11006 gnd.n2097 gnd.n2092 9.3005
R11007 gnd.n2543 gnd.n2542 9.3005
R11008 gnd.n2280 gnd.n2279 9.3005
R11009 gnd.n2278 gnd.n2144 9.3005
R11010 gnd.n2575 gnd.n2574 9.3005
R11011 gnd.n2577 gnd.n2576 9.3005
R11012 gnd.n2132 gnd.n2131 9.3005
R11013 gnd.n2583 gnd.n2582 9.3005
R11014 gnd.n2585 gnd.n2584 9.3005
R11015 gnd.n2124 gnd.n2123 9.3005
R11016 gnd.n2591 gnd.n2590 9.3005
R11017 gnd.n2593 gnd.n2592 9.3005
R11018 gnd.n2114 gnd.n2113 9.3005
R11019 gnd.n2599 gnd.n2598 9.3005
R11020 gnd.n2601 gnd.n2600 9.3005
R11021 gnd.n2106 gnd.n2105 9.3005
R11022 gnd.n2607 gnd.n2606 9.3005
R11023 gnd.n2609 gnd.n2608 9.3005
R11024 gnd.n2096 gnd.n2095 9.3005
R11025 gnd.n2615 gnd.n2614 9.3005
R11026 gnd.n2617 gnd.n2616 9.3005
R11027 gnd.n2618 gnd.n2090 9.3005
R11028 gnd.n2621 gnd.n2620 9.3005
R11029 gnd.n2622 gnd.n2086 9.3005
R11030 gnd.n2624 gnd.n2623 9.3005
R11031 gnd.n2625 gnd.n2085 9.3005
R11032 gnd.n2627 gnd.n2626 9.3005
R11033 gnd.n2628 gnd.n2082 9.3005
R11034 gnd.n2630 gnd.n2629 9.3005
R11035 gnd.n2631 gnd.n2081 9.3005
R11036 gnd.n2060 gnd.n2059 9.3005
R11037 gnd.n2659 gnd.n2658 9.3005
R11038 gnd.n2660 gnd.n2057 9.3005
R11039 gnd.n2663 gnd.n2662 9.3005
R11040 gnd.n2661 gnd.n2058 9.3005
R11041 gnd.n2035 gnd.n2034 9.3005
R11042 gnd.n2689 gnd.n2688 9.3005
R11043 gnd.n2690 gnd.n2032 9.3005
R11044 gnd.n2693 gnd.n2692 9.3005
R11045 gnd.n2691 gnd.n2033 9.3005
R11046 gnd.n2010 gnd.n2009 9.3005
R11047 gnd.n2719 gnd.n2718 9.3005
R11048 gnd.n2720 gnd.n2007 9.3005
R11049 gnd.n2723 gnd.n2722 9.3005
R11050 gnd.n2721 gnd.n2008 9.3005
R11051 gnd.n1985 gnd.n1984 9.3005
R11052 gnd.n2766 gnd.n2765 9.3005
R11053 gnd.n2767 gnd.n1982 9.3005
R11054 gnd.n2770 gnd.n2769 9.3005
R11055 gnd.n2768 gnd.n1983 9.3005
R11056 gnd.n1479 gnd.n1477 9.3005
R11057 gnd.n3792 gnd.n3791 9.3005
R11058 gnd.n3790 gnd.n1478 9.3005
R11059 gnd.n3789 gnd.n3788 9.3005
R11060 gnd.n3787 gnd.n1480 9.3005
R11061 gnd.n3786 gnd.n3785 9.3005
R11062 gnd.n3784 gnd.n1484 9.3005
R11063 gnd.n3783 gnd.n3782 9.3005
R11064 gnd.n3781 gnd.n1485 9.3005
R11065 gnd.n3780 gnd.n3779 9.3005
R11066 gnd.n3778 gnd.n1489 9.3005
R11067 gnd.n3777 gnd.n3776 9.3005
R11068 gnd.n3775 gnd.n1490 9.3005
R11069 gnd.n3774 gnd.n3773 9.3005
R11070 gnd.n3772 gnd.n1494 9.3005
R11071 gnd.n3771 gnd.n3770 9.3005
R11072 gnd.n3769 gnd.n1495 9.3005
R11073 gnd.n3768 gnd.n3767 9.3005
R11074 gnd.n3766 gnd.n1499 9.3005
R11075 gnd.n3765 gnd.n3764 9.3005
R11076 gnd.n3763 gnd.n1500 9.3005
R11077 gnd.n3762 gnd.n3761 9.3005
R11078 gnd.n3760 gnd.n1504 9.3005
R11079 gnd.n3759 gnd.n3758 9.3005
R11080 gnd.n3757 gnd.n1505 9.3005
R11081 gnd.n3756 gnd.n3755 9.3005
R11082 gnd.n3754 gnd.n1509 9.3005
R11083 gnd.n3753 gnd.n3752 9.3005
R11084 gnd.n3751 gnd.n1510 9.3005
R11085 gnd.n3750 gnd.n3749 9.3005
R11086 gnd.n3748 gnd.n1514 9.3005
R11087 gnd.n3747 gnd.n3746 9.3005
R11088 gnd.n3745 gnd.n1515 9.3005
R11089 gnd.n3744 gnd.n3743 9.3005
R11090 gnd.n3742 gnd.n1519 9.3005
R11091 gnd.n3741 gnd.n3740 9.3005
R11092 gnd.n3739 gnd.n1520 9.3005
R11093 gnd.n3738 gnd.n3737 9.3005
R11094 gnd.n3736 gnd.n1524 9.3005
R11095 gnd.n3735 gnd.n3734 9.3005
R11096 gnd.n3733 gnd.n1525 9.3005
R11097 gnd.n3732 gnd.n3731 9.3005
R11098 gnd.n3730 gnd.n1529 9.3005
R11099 gnd.n3729 gnd.n3728 9.3005
R11100 gnd.n3727 gnd.n1530 9.3005
R11101 gnd.n3726 gnd.n3725 9.3005
R11102 gnd.n3724 gnd.n1534 9.3005
R11103 gnd.n3723 gnd.n3722 9.3005
R11104 gnd.n3721 gnd.n1535 9.3005
R11105 gnd.n3720 gnd.n3719 9.3005
R11106 gnd.n3718 gnd.n1539 9.3005
R11107 gnd.n3717 gnd.n3716 9.3005
R11108 gnd.n3715 gnd.n1540 9.3005
R11109 gnd.n3714 gnd.n3713 9.3005
R11110 gnd.n3712 gnd.n1544 9.3005
R11111 gnd.n3711 gnd.n3710 9.3005
R11112 gnd.n3709 gnd.n1545 9.3005
R11113 gnd.n3708 gnd.n3707 9.3005
R11114 gnd.n3706 gnd.n1549 9.3005
R11115 gnd.n3705 gnd.n3704 9.3005
R11116 gnd.n3703 gnd.n1550 9.3005
R11117 gnd.n3702 gnd.n3701 9.3005
R11118 gnd.n3700 gnd.n1554 9.3005
R11119 gnd.n3699 gnd.n3698 9.3005
R11120 gnd.n3697 gnd.n1555 9.3005
R11121 gnd.n3696 gnd.n3695 9.3005
R11122 gnd.n3694 gnd.n1559 9.3005
R11123 gnd.n3693 gnd.n3692 9.3005
R11124 gnd.n3691 gnd.n1560 9.3005
R11125 gnd.n3690 gnd.n3689 9.3005
R11126 gnd.n3688 gnd.n1564 9.3005
R11127 gnd.n3687 gnd.n3686 9.3005
R11128 gnd.n3685 gnd.n1565 9.3005
R11129 gnd.n3684 gnd.n3683 9.3005
R11130 gnd.n3682 gnd.n1569 9.3005
R11131 gnd.n3681 gnd.n3680 9.3005
R11132 gnd.n3679 gnd.n1570 9.3005
R11133 gnd.n3678 gnd.n3677 9.3005
R11134 gnd.n462 gnd.n461 9.3005
R11135 gnd.n6369 gnd.n6368 9.3005
R11136 gnd.n2633 gnd.n2632 9.3005
R11137 gnd.n6365 gnd.n463 9.3005
R11138 gnd.n6364 gnd.n6363 9.3005
R11139 gnd.n6362 gnd.n466 9.3005
R11140 gnd.n6361 gnd.n6360 9.3005
R11141 gnd.n6359 gnd.n467 9.3005
R11142 gnd.n391 gnd.n389 9.3005
R11143 gnd.n6367 gnd.n6366 9.3005
R11144 gnd.n6387 gnd.n6386 9.3005
R11145 gnd.n438 gnd.n437 9.3005
R11146 gnd.n6393 gnd.n6392 9.3005
R11147 gnd.n6395 gnd.n6394 9.3005
R11148 gnd.n430 gnd.n429 9.3005
R11149 gnd.n6401 gnd.n6400 9.3005
R11150 gnd.n6403 gnd.n6402 9.3005
R11151 gnd.n420 gnd.n419 9.3005
R11152 gnd.n6409 gnd.n6408 9.3005
R11153 gnd.n6411 gnd.n6410 9.3005
R11154 gnd.n412 gnd.n411 9.3005
R11155 gnd.n6417 gnd.n6416 9.3005
R11156 gnd.n6419 gnd.n6418 9.3005
R11157 gnd.n402 gnd.n401 9.3005
R11158 gnd.n6425 gnd.n6424 9.3005
R11159 gnd.n6427 gnd.n6426 9.3005
R11160 gnd.n398 gnd.n396 9.3005
R11161 gnd.n6385 gnd.n6381 9.3005
R11162 gnd.n448 gnd.n447 9.3005
R11163 gnd.n6432 gnd.n6431 9.3005
R11164 gnd.n6430 gnd.n390 9.3005
R11165 gnd.n6429 gnd.n6428 9.3005
R11166 gnd.n397 gnd.n395 9.3005
R11167 gnd.n6423 gnd.n6422 9.3005
R11168 gnd.n6421 gnd.n6420 9.3005
R11169 gnd.n406 gnd.n405 9.3005
R11170 gnd.n6415 gnd.n6414 9.3005
R11171 gnd.n6413 gnd.n6412 9.3005
R11172 gnd.n416 gnd.n415 9.3005
R11173 gnd.n6407 gnd.n6406 9.3005
R11174 gnd.n6405 gnd.n6404 9.3005
R11175 gnd.n424 gnd.n423 9.3005
R11176 gnd.n6399 gnd.n6398 9.3005
R11177 gnd.n6397 gnd.n6396 9.3005
R11178 gnd.n434 gnd.n433 9.3005
R11179 gnd.n6391 gnd.n6390 9.3005
R11180 gnd.n6389 gnd.n6388 9.3005
R11181 gnd.n449 gnd.n444 9.3005
R11182 gnd.n6380 gnd.n6379 9.3005
R11183 gnd.n6378 gnd.n6377 9.3005
R11184 gnd.n6559 gnd.n6558 9.3005
R11185 gnd.n6560 gnd.n269 9.3005
R11186 gnd.n6563 gnd.n6562 9.3005
R11187 gnd.n6561 gnd.n270 9.3005
R11188 gnd.n244 gnd.n243 9.3005
R11189 gnd.n6594 gnd.n6593 9.3005
R11190 gnd.n6595 gnd.n241 9.3005
R11191 gnd.n6608 gnd.n6607 9.3005
R11192 gnd.n6606 gnd.n242 9.3005
R11193 gnd.n6605 gnd.n6604 9.3005
R11194 gnd.n6603 gnd.n6596 9.3005
R11195 gnd.n6602 gnd.n6601 9.3005
R11196 gnd.n6600 gnd.n6599 9.3005
R11197 gnd.n199 gnd.n198 9.3005
R11198 gnd.n6658 gnd.n6657 9.3005
R11199 gnd.n6659 gnd.n196 9.3005
R11200 gnd.n6666 gnd.n6665 9.3005
R11201 gnd.n6664 gnd.n197 9.3005
R11202 gnd.n6663 gnd.n6662 9.3005
R11203 gnd.n6661 gnd.n67 9.3005
R11204 gnd.n272 gnd.n271 9.3005
R11205 gnd.n7128 gnd.n68 9.3005
R11206 gnd.t269 gnd.n4349 9.24152
R11207 gnd.n4251 gnd.t77 9.24152
R11208 gnd.n5519 gnd.t178 9.24152
R11209 gnd.t38 gnd.t269 8.92286
R11210 gnd.n2932 gnd.n1951 8.92286
R11211 gnd.n2871 gnd.t70 8.92286
R11212 gnd.n3023 gnd.n1887 8.92286
R11213 gnd.n3076 gnd.n3075 8.92286
R11214 gnd.n3184 gnd.n1794 8.92286
R11215 gnd.n3215 gnd.n3214 8.92286
R11216 gnd.n3327 gnd.n3326 8.92286
R11217 gnd.n3494 gnd.n1676 8.92286
R11218 gnd.n5489 gnd.n5464 8.92171
R11219 gnd.n5457 gnd.n5432 8.92171
R11220 gnd.n5425 gnd.n5400 8.92171
R11221 gnd.n5394 gnd.n5369 8.92171
R11222 gnd.n5362 gnd.n5337 8.92171
R11223 gnd.n5330 gnd.n5305 8.92171
R11224 gnd.n5298 gnd.n5273 8.92171
R11225 gnd.n5267 gnd.n5242 8.92171
R11226 gnd.n3423 gnd.n3405 8.72777
R11227 gnd.n4993 gnd.t274 8.60421
R11228 gnd.n2645 gnd.t106 8.60421
R11229 gnd.n2705 gnd.t19 8.60421
R11230 gnd.n3618 gnd.t244 8.60421
R11231 gnd.t73 gnd.n3674 8.60421
R11232 gnd.n6322 gnd.n116 8.60421
R11233 gnd.n4413 gnd.n4401 8.43656
R11234 gnd.n42 gnd.n30 8.43656
R11235 gnd.t162 gnd.n1968 8.28555
R11236 gnd.n2999 gnd.n1905 8.28555
R11237 gnd.n3068 gnd.n3067 8.28555
R11238 gnd.n3163 gnd.n1811 8.28555
R11239 gnd.n3258 gnd.n1759 8.28555
R11240 gnd.t132 gnd.n1681 8.28555
R11241 gnd.n5490 gnd.n5462 8.14595
R11242 gnd.n5458 gnd.n5430 8.14595
R11243 gnd.n5426 gnd.n5398 8.14595
R11244 gnd.n5395 gnd.n5367 8.14595
R11245 gnd.n5363 gnd.n5335 8.14595
R11246 gnd.n5331 gnd.n5303 8.14595
R11247 gnd.n5299 gnd.n5271 8.14595
R11248 gnd.n5268 gnd.n5240 8.14595
R11249 gnd.n2408 gnd.n0 8.10675
R11250 gnd.n7129 gnd.n7128 8.10675
R11251 gnd.n5495 gnd.n5494 7.97301
R11252 gnd.t272 gnd.n4508 7.9669
R11253 gnd.n2557 gnd.n2555 7.9669
R11254 gnd.n6355 gnd.n470 7.9669
R11255 gnd.n7129 gnd.n66 7.78567
R11256 gnd.n6385 gnd.n447 7.75808
R11257 gnd.n6850 gnd.n6753 7.75808
R11258 gnd.n2571 gnd.n2570 7.75808
R11259 gnd.n2363 gnd.n2362 7.75808
R11260 gnd.n3000 gnd.n2999 7.64824
R11261 gnd.t186 gnd.n1860 7.64824
R11262 gnd.n3082 gnd.t306 7.64824
R11263 gnd.n3068 gnd.n1846 7.64824
R11264 gnd.n3135 gnd.n1811 7.64824
R11265 gnd.n3165 gnd.t304 7.64824
R11266 gnd.n3195 gnd.t263 7.64824
R11267 gnd.n3258 gnd.n1761 7.64824
R11268 gnd.t88 gnd.n3378 7.64824
R11269 gnd.n4438 gnd.n4437 7.53171
R11270 gnd.n4902 gnd.t267 7.32958
R11271 gnd.t106 gnd.n2644 7.32958
R11272 gnd.n2030 gnd.t19 7.32958
R11273 gnd.t244 gnd.n3617 7.32958
R11274 gnd.n3675 gnd.t73 7.32958
R11275 gnd.n1467 gnd.n1466 7.30353
R11276 gnd.n3422 gnd.n3421 7.30353
R11277 gnd.n4862 gnd.n4581 7.01093
R11278 gnd.n4584 gnd.n4582 7.01093
R11279 gnd.n4872 gnd.n4871 7.01093
R11280 gnd.n4883 gnd.n4565 7.01093
R11281 gnd.n4882 gnd.n4568 7.01093
R11282 gnd.n4893 gnd.n4556 7.01093
R11283 gnd.n4559 gnd.n4557 7.01093
R11284 gnd.n4903 gnd.n4902 7.01093
R11285 gnd.n4913 gnd.n4537 7.01093
R11286 gnd.n4912 gnd.n4540 7.01093
R11287 gnd.n4921 gnd.n4531 7.01093
R11288 gnd.n4933 gnd.n4521 7.01093
R11289 gnd.n4943 gnd.n4506 7.01093
R11290 gnd.n4959 gnd.n4958 7.01093
R11291 gnd.n4508 gnd.n4445 7.01093
R11292 gnd.n5013 gnd.n4446 7.01093
R11293 gnd.n5007 gnd.n5006 7.01093
R11294 gnd.n4495 gnd.n4457 7.01093
R11295 gnd.n4999 gnd.n4468 7.01093
R11296 gnd.n4486 gnd.n4481 7.01093
R11297 gnd.n4993 gnd.n4992 7.01093
R11298 gnd.n5039 gnd.n4384 7.01093
R11299 gnd.n5038 gnd.n5037 7.01093
R11300 gnd.n5050 gnd.n5049 7.01093
R11301 gnd.n4377 gnd.n4369 7.01093
R11302 gnd.n5079 gnd.n4357 7.01093
R11303 gnd.n5078 gnd.n4360 7.01093
R11304 gnd.n5089 gnd.n4349 7.01093
R11305 gnd.n4350 gnd.n4338 7.01093
R11306 gnd.n5100 gnd.n4339 7.01093
R11307 gnd.n5124 gnd.n4330 7.01093
R11308 gnd.n5123 gnd.n4321 7.01093
R11309 gnd.n5146 gnd.n5145 7.01093
R11310 gnd.n5164 gnd.n4302 7.01093
R11311 gnd.n5163 gnd.n4305 7.01093
R11312 gnd.n5174 gnd.n4294 7.01093
R11313 gnd.n4295 gnd.n4282 7.01093
R11314 gnd.n5185 gnd.n4283 7.01093
R11315 gnd.n5212 gnd.n4267 7.01093
R11316 gnd.n5224 gnd.n5223 7.01093
R11317 gnd.n5206 gnd.n4260 7.01093
R11318 gnd.n5235 gnd.n5234 7.01093
R11319 gnd.n5507 gnd.n4248 7.01093
R11320 gnd.n5506 gnd.n4251 7.01093
R11321 gnd.n5519 gnd.n4240 7.01093
R11322 gnd.n4241 gnd.n4233 7.01093
R11323 gnd.n5529 gnd.n1008 7.01093
R11324 gnd.n2893 gnd.n1471 7.01093
R11325 gnd.n2923 gnd.n1951 7.01093
R11326 gnd.t70 gnd.n1953 7.01093
R11327 gnd.n3031 gnd.n1887 7.01093
R11328 gnd.n3055 gnd.t186 7.01093
R11329 gnd.n3076 gnd.n1860 7.01093
R11330 gnd.n3195 gnd.n1794 7.01093
R11331 gnd.t263 gnd.n3194 7.01093
R11332 gnd.n3214 gnd.n1775 7.01093
R11333 gnd.n3494 gnd.n1675 7.01093
R11334 gnd.n4540 gnd.t268 6.69227
R11335 gnd.n4360 gnd.t38 6.69227
R11336 gnd.n5213 gnd.t264 6.69227
R11337 gnd.n2872 gnd.t323 6.69227
R11338 gnd.t190 gnd.n3311 6.69227
R11339 gnd.n3555 gnd.n3554 6.5566
R11340 gnd.n2782 gnd.n2781 6.5566
R11341 gnd.n3806 gnd.n3802 6.5566
R11342 gnd.n3433 gnd.n3432 6.5566
R11343 gnd.t81 gnd.n2893 6.37362
R11344 gnd.n2857 gnd.n1918 6.37362
R11345 gnd.n1881 gnd.t185 6.37362
R11346 gnd.n3114 gnd.n1841 6.37362
R11347 gnd.n3144 gnd.n1817 6.37362
R11348 gnd.n3204 gnd.t257 6.37362
R11349 gnd.n3285 gnd.n3284 6.37362
R11350 gnd.n2278 gnd.n2143 6.20656
R11351 gnd.n449 gnd.n443 6.20656
R11352 gnd.t210 gnd.n4969 6.05496
R11353 gnd.n4970 gnd.t288 6.05496
R11354 gnd.t325 gnd.n4384 6.05496
R11355 gnd.t294 gnd.n5134 6.05496
R11356 gnd.t314 gnd.t305 6.05496
R11357 gnd.t204 gnd.t250 6.05496
R11358 gnd.n5492 gnd.n5462 5.81868
R11359 gnd.n5460 gnd.n5430 5.81868
R11360 gnd.n5428 gnd.n5398 5.81868
R11361 gnd.n5397 gnd.n5367 5.81868
R11362 gnd.n5365 gnd.n5335 5.81868
R11363 gnd.n5333 gnd.n5303 5.81868
R11364 gnd.n5301 gnd.n5271 5.81868
R11365 gnd.n5270 gnd.n5240 5.81868
R11366 gnd.n2906 gnd.n2905 5.73631
R11367 gnd.n3042 gnd.n3041 5.73631
R11368 gnd.n3049 gnd.n1873 5.73631
R11369 gnd.n3067 gnd.t306 5.73631
R11370 gnd.t304 gnd.n3163 5.73631
R11371 gnd.n3203 gnd.n1788 5.73631
R11372 gnd.n3234 gnd.n1779 5.73631
R11373 gnd.n3372 gnd.n1693 5.73631
R11374 gnd.n3559 gnd.n351 5.62001
R11375 gnd.n3868 gnd.n1409 5.62001
R11376 gnd.n3868 gnd.n1410 5.62001
R11377 gnd.n3428 gnd.n351 5.62001
R11378 gnd.n4721 gnd.n4716 5.4308
R11379 gnd.n5537 gnd.n4226 5.4308
R11380 gnd.n5037 gnd.t266 5.41765
R11381 gnd.t293 gnd.n5060 5.41765
R11382 gnd.t214 gnd.n4314 5.41765
R11383 gnd.n5621 gnd.n1008 5.41765
R11384 gnd.n2980 gnd.t197 5.41765
R11385 gnd.n3282 gnd.t236 5.41765
R11386 gnd.t287 gnd.n2940 5.09899
R11387 gnd.n2973 gnd.n1922 5.09899
R11388 gnd.n3093 gnd.n1834 5.09899
R11389 gnd.n3125 gnd.n3124 5.09899
R11390 gnd.n1741 gnd.n1740 5.09899
R11391 gnd.t262 gnd.n1720 5.09899
R11392 gnd.n5490 gnd.n5489 5.04292
R11393 gnd.n5458 gnd.n5457 5.04292
R11394 gnd.n5426 gnd.n5425 5.04292
R11395 gnd.n5395 gnd.n5394 5.04292
R11396 gnd.n5363 gnd.n5362 5.04292
R11397 gnd.n5331 gnd.n5330 5.04292
R11398 gnd.n5299 gnd.n5298 5.04292
R11399 gnd.n5268 gnd.n5267 5.04292
R11400 gnd.n5000 gnd.t289 4.78034
R11401 gnd.n4339 gnd.t273 4.78034
R11402 gnd.t0 gnd.n1996 4.78034
R11403 gnd.n3584 gnd.t246 4.78034
R11404 gnd.n4442 gnd.n4439 4.74817
R11405 gnd.n4492 gnd.n4390 4.74817
R11406 gnd.n4479 gnd.n4389 4.74817
R11407 gnd.n4388 gnd.n4387 4.74817
R11408 gnd.n4488 gnd.n4439 4.74817
R11409 gnd.n4489 gnd.n4390 4.74817
R11410 gnd.n4491 gnd.n4389 4.74817
R11411 gnd.n4478 gnd.n4388 4.74817
R11412 gnd.n4437 gnd.n4436 4.74296
R11413 gnd.n66 gnd.n65 4.74296
R11414 gnd.n4413 gnd.n4412 4.7074
R11415 gnd.n4425 gnd.n4424 4.7074
R11416 gnd.n42 gnd.n41 4.7074
R11417 gnd.n54 gnd.n53 4.7074
R11418 gnd.n4437 gnd.n4425 4.65959
R11419 gnd.n66 gnd.n54 4.65959
R11420 gnd.n6497 gnd.n353 4.6132
R11421 gnd.n3869 gnd.n1408 4.6132
R11422 gnd.n2887 gnd.n1474 4.46168
R11423 gnd.n2881 gnd.n2880 4.46168
R11424 gnd.t187 gnd.n1890 4.46168
R11425 gnd.n2842 gnd.n2841 4.46168
R11426 gnd.n3058 gnd.n1868 4.46168
R11427 gnd.n3174 gnd.n1808 4.46168
R11428 gnd.n3242 gnd.n1772 4.46168
R11429 gnd.t261 gnd.n3241 4.46168
R11430 gnd.n3327 gnd.t113 4.46168
R11431 gnd.n3380 gnd.n1698 4.46168
R11432 gnd.n3401 gnd.n3400 4.46168
R11433 gnd.n3418 gnd.n3405 4.46111
R11434 gnd.n5475 gnd.n5471 4.38594
R11435 gnd.n5443 gnd.n5439 4.38594
R11436 gnd.n5411 gnd.n5407 4.38594
R11437 gnd.n5380 gnd.n5376 4.38594
R11438 gnd.n5348 gnd.n5344 4.38594
R11439 gnd.n5316 gnd.n5312 4.38594
R11440 gnd.n5284 gnd.n5280 4.38594
R11441 gnd.n5253 gnd.n5249 4.38594
R11442 gnd.n5486 gnd.n5464 4.26717
R11443 gnd.n5454 gnd.n5432 4.26717
R11444 gnd.n5422 gnd.n5400 4.26717
R11445 gnd.n5391 gnd.n5369 4.26717
R11446 gnd.n5359 gnd.n5337 4.26717
R11447 gnd.n5327 gnd.n5305 4.26717
R11448 gnd.n5295 gnd.n5273 4.26717
R11449 gnd.n5264 gnd.n5242 4.26717
R11450 gnd.n4944 gnd.t270 4.14303
R11451 gnd.n5174 gnd.t275 4.14303
R11452 gnd.n5494 gnd.n5493 4.08274
R11453 gnd.n3554 gnd.n3553 4.05904
R11454 gnd.n2783 gnd.n2782 4.05904
R11455 gnd.n3809 gnd.n3802 4.05904
R11456 gnd.n3434 gnd.n3433 4.05904
R11457 gnd.n19 gnd.n9 3.99943
R11458 gnd.n3919 gnd.n1350 3.82437
R11459 gnd.n2949 gnd.n2948 3.82437
R11460 gnd.n2971 gnd.t226 3.82437
R11461 gnd.n2993 gnd.n2992 3.82437
R11462 gnd.n3103 gnd.n3101 3.82437
R11463 gnd.n3115 gnd.t305 3.82437
R11464 gnd.n3155 gnd.t204 3.82437
R11465 gnd.n3154 gnd.n1819 3.82437
R11466 gnd.n3268 gnd.n3267 3.82437
R11467 gnd.t8 gnd.n3292 3.82437
R11468 gnd.n3318 gnd.n1718 3.82437
R11469 gnd.n6546 gnd.n284 3.82437
R11470 gnd.n5017 gnd.n4438 3.81325
R11471 gnd.n4425 gnd.n4413 3.72967
R11472 gnd.n54 gnd.n42 3.72967
R11473 gnd.n5494 gnd.n5366 3.70378
R11474 gnd.n19 gnd.n18 3.60163
R11475 gnd.n2675 gnd.t192 3.50571
R11476 gnd.t280 gnd.n3637 3.50571
R11477 gnd.n5485 gnd.n5466 3.49141
R11478 gnd.n5453 gnd.n5434 3.49141
R11479 gnd.n5421 gnd.n5402 3.49141
R11480 gnd.n5390 gnd.n5371 3.49141
R11481 gnd.n5358 gnd.n5339 3.49141
R11482 gnd.n5326 gnd.n5307 3.49141
R11483 gnd.n5294 gnd.n5275 3.49141
R11484 gnd.n5263 gnd.n5244 3.49141
R11485 gnd.n7020 gnd.n7017 3.29747
R11486 gnd.n7021 gnd.n7020 3.29747
R11487 gnd.n6515 gnd.n6514 3.29747
R11488 gnd.n6514 gnd.n6513 3.29747
R11489 gnd.n4138 gnd.n4137 3.29747
R11490 gnd.n4137 gnd.n4136 3.29747
R11491 gnd.n3887 gnd.n3886 3.29747
R11492 gnd.n3886 gnd.n3885 3.29747
R11493 gnd.n3945 gnd.n1302 3.18706
R11494 gnd.n2496 gnd.n1309 3.18706
R11495 gnd.n3939 gnd.n1312 3.18706
R11496 gnd.n2505 gnd.n1320 3.18706
R11497 gnd.n3933 gnd.n1323 3.18706
R11498 gnd.n2535 gnd.n2534 3.18706
R11499 gnd.n3927 gnd.n1332 3.18706
R11500 gnd.n2567 gnd.n2566 3.18706
R11501 gnd.n2887 gnd.t162 3.18706
R11502 gnd.n2913 gnd.t175 3.18706
R11503 gnd.n2913 gnd.t84 3.18706
R11504 gnd.n2930 gnd.n1953 3.18706
R11505 gnd.n2864 gnd.t260 3.18706
R11506 gnd.n2961 gnd.t260 3.18706
R11507 gnd.n3024 gnd.n1894 3.18706
R11508 gnd.n3074 gnd.n1855 3.18706
R11509 gnd.n3185 gnd.n1801 3.18706
R11510 gnd.n3251 gnd.n3250 3.18706
R11511 gnd.n3302 gnd.t307 3.18706
R11512 gnd.n3320 gnd.t307 3.18706
R11513 gnd.n3346 gnd.n1711 3.18706
R11514 gnd.n3387 gnd.t91 3.18706
R11515 gnd.t103 gnd.n1675 3.18706
R11516 gnd.n6346 gnd.n6345 3.18706
R11517 gnd.n6556 gnd.n274 3.18706
R11518 gnd.n6339 gnd.n6338 3.18706
R11519 gnd.n6565 gnd.n267 3.18706
R11520 gnd.n6581 gnd.n255 3.18706
R11521 gnd.n6569 gnd.n258 3.18706
R11522 gnd.n6591 gnd.n246 3.18706
R11523 gnd.n516 gnd.n239 3.18706
R11524 gnd.n4523 gnd.t270 2.8684
R11525 gnd.n3865 gnd.n1413 2.8684
R11526 gnd.n2904 gnd.t312 2.8684
R11527 gnd.t45 gnd.n3386 2.8684
R11528 gnd.n3565 gnd.n3562 2.8684
R11529 gnd.n4426 gnd.t10 2.82907
R11530 gnd.n4426 gnd.t194 2.82907
R11531 gnd.n4428 gnd.t295 2.82907
R11532 gnd.n4428 gnd.t50 2.82907
R11533 gnd.n4430 gnd.t202 2.82907
R11534 gnd.n4430 gnd.t12 2.82907
R11535 gnd.n4432 gnd.t217 2.82907
R11536 gnd.n4432 gnd.t184 2.82907
R11537 gnd.n4434 gnd.t297 2.82907
R11538 gnd.n4434 gnd.t7 2.82907
R11539 gnd.n4391 gnd.t203 2.82907
R11540 gnd.n4391 gnd.t49 2.82907
R11541 gnd.n4393 gnd.t239 2.82907
R11542 gnd.n4393 gnd.t240 2.82907
R11543 gnd.n4395 gnd.t311 2.82907
R11544 gnd.n4395 gnd.t277 2.82907
R11545 gnd.n4397 gnd.t249 2.82907
R11546 gnd.n4397 gnd.t183 2.82907
R11547 gnd.n4399 gnd.t320 2.82907
R11548 gnd.n4399 gnd.t256 2.82907
R11549 gnd.n4402 gnd.t252 2.82907
R11550 gnd.n4402 gnd.t32 2.82907
R11551 gnd.n4404 gnd.t230 2.82907
R11552 gnd.n4404 gnd.t48 2.82907
R11553 gnd.n4406 gnd.t189 2.82907
R11554 gnd.n4406 gnd.t308 2.82907
R11555 gnd.n4408 gnd.t207 2.82907
R11556 gnd.n4408 gnd.t37 2.82907
R11557 gnd.n4410 gnd.t196 2.82907
R11558 gnd.n4410 gnd.t51 2.82907
R11559 gnd.n4414 gnd.t220 2.82907
R11560 gnd.n4414 gnd.t317 2.82907
R11561 gnd.n4416 gnd.t223 2.82907
R11562 gnd.n4416 gnd.t59 2.82907
R11563 gnd.n4418 gnd.t27 2.82907
R11564 gnd.n4418 gnd.t283 2.82907
R11565 gnd.n4420 gnd.t276 2.82907
R11566 gnd.n4420 gnd.t43 2.82907
R11567 gnd.n4422 gnd.t329 2.82907
R11568 gnd.n4422 gnd.t241 2.82907
R11569 gnd.n63 gnd.t14 2.82907
R11570 gnd.n63 gnd.t213 2.82907
R11571 gnd.n61 gnd.t208 2.82907
R11572 gnd.n61 gnd.t309 2.82907
R11573 gnd.n59 gnd.t301 2.82907
R11574 gnd.n59 gnd.t188 2.82907
R11575 gnd.n57 gnd.t258 2.82907
R11576 gnd.n57 gnd.t205 2.82907
R11577 gnd.n55 gnd.t310 2.82907
R11578 gnd.n55 gnd.t282 2.82907
R11579 gnd.n28 gnd.t28 2.82907
R11580 gnd.n28 gnd.t296 2.82907
R11581 gnd.n26 gnd.t238 2.82907
R11582 gnd.n26 gnd.t302 2.82907
R11583 gnd.n24 gnd.t182 2.82907
R11584 gnd.n24 gnd.t284 2.82907
R11585 gnd.n22 gnd.t216 2.82907
R11586 gnd.n22 gnd.t209 2.82907
R11587 gnd.n20 gnd.t290 2.82907
R11588 gnd.n20 gnd.t16 2.82907
R11589 gnd.n39 gnd.t212 2.82907
R11590 gnd.n39 gnd.t201 2.82907
R11591 gnd.n37 gnd.t41 2.82907
R11592 gnd.n37 gnd.t255 2.82907
R11593 gnd.n35 gnd.t285 2.82907
R11594 gnd.n35 gnd.t44 2.82907
R11595 gnd.n33 gnd.t55 2.82907
R11596 gnd.n33 gnd.t18 2.82907
R11597 gnd.n31 gnd.t231 2.82907
R11598 gnd.n31 gnd.t286 2.82907
R11599 gnd.n51 gnd.t199 2.82907
R11600 gnd.n51 gnd.t292 2.82907
R11601 gnd.n49 gnd.t299 2.82907
R11602 gnd.n49 gnd.t330 2.82907
R11603 gnd.n47 gnd.t248 2.82907
R11604 gnd.n47 gnd.t34 2.82907
R11605 gnd.n45 gnd.t58 2.82907
R11606 gnd.n45 gnd.t56 2.82907
R11607 gnd.n43 gnd.t3 2.82907
R11608 gnd.n43 gnd.t259 2.82907
R11609 gnd.n5482 gnd.n5481 2.71565
R11610 gnd.n5450 gnd.n5449 2.71565
R11611 gnd.n5418 gnd.n5417 2.71565
R11612 gnd.n5387 gnd.n5386 2.71565
R11613 gnd.n5355 gnd.n5354 2.71565
R11614 gnd.n5323 gnd.n5322 2.71565
R11615 gnd.n5291 gnd.n5290 2.71565
R11616 gnd.n5260 gnd.n5259 2.71565
R11617 gnd.n2894 gnd.t81 2.54975
R11618 gnd.t84 gnd.n2912 2.54975
R11619 gnd.n2873 gnd.n2871 2.54975
R11620 gnd.n2941 gnd.t287 2.54975
R11621 gnd.n2850 gnd.n2849 2.54975
R11622 gnd.n2849 gnd.t35 2.54975
R11623 gnd.n3083 gnd.n3082 2.54975
R11624 gnd.n3165 gnd.n3164 2.54975
R11625 gnd.n3218 gnd.t57 2.54975
R11626 gnd.n3218 gnd.n3217 2.54975
R11627 gnd.n3312 gnd.t262 2.54975
R11628 gnd.n3348 gnd.n1710 2.54975
R11629 gnd.t113 gnd.n1703 2.54975
R11630 gnd.n3379 gnd.t88 2.54975
R11631 gnd.n3378 gnd.t91 2.54975
R11632 gnd.n5017 gnd.n4439 2.27742
R11633 gnd.n5017 gnd.n4390 2.27742
R11634 gnd.n5017 gnd.n4389 2.27742
R11635 gnd.n5017 gnd.n4388 2.27742
R11636 gnd.n4871 gnd.t125 2.23109
R11637 gnd.n4494 gnd.t289 2.23109
R11638 gnd.n3058 gnd.t234 2.23109
R11639 gnd.n3101 gnd.t314 2.23109
R11640 gnd.t250 gnd.n3154 2.23109
R11641 gnd.n1808 gnd.t218 2.23109
R11642 gnd.n5478 gnd.n5468 1.93989
R11643 gnd.n5446 gnd.n5436 1.93989
R11644 gnd.n5414 gnd.n5404 1.93989
R11645 gnd.n5383 gnd.n5373 1.93989
R11646 gnd.n5351 gnd.n5341 1.93989
R11647 gnd.n5319 gnd.n5309 1.93989
R11648 gnd.n5287 gnd.n5277 1.93989
R11649 gnd.n5256 gnd.n5246 1.93989
R11650 gnd.n2950 gnd.n1938 1.91244
R11651 gnd.n2990 gnd.n1903 1.91244
R11652 gnd.n3105 gnd.n3104 1.91244
R11653 gnd.n3134 gnd.n1831 1.91244
R11654 gnd.n3269 gnd.n1754 1.91244
R11655 gnd.n3336 gnd.n3335 1.91244
R11656 gnd.n3372 gnd.t132 1.91244
R11657 gnd.n3565 gnd.t138 1.91244
R11658 gnd.t242 gnd.n4882 1.59378
R11659 gnd.n5061 gnd.t293 1.59378
R11660 gnd.n4323 gnd.t214 1.59378
R11661 gnd.n2941 gnd.t323 1.59378
R11662 gnd.t278 gnd.n3023 1.59378
R11663 gnd.n3215 gnd.t327 1.59378
R11664 gnd.n3312 gnd.t190 1.59378
R11665 gnd.n3795 gnd.n3794 1.27512
R11666 gnd.n2924 gnd.n1957 1.27512
R11667 gnd.t226 gnd.n2970 1.27512
R11668 gnd.n3030 gnd.n1890 1.27512
R11669 gnd.n3057 gnd.n3055 1.27512
R11670 gnd.n3194 gnd.n1796 1.27512
R11671 gnd.n3241 gnd.n3240 1.27512
R11672 gnd.n3293 gnd.t8 1.27512
R11673 gnd.n3366 gnd.n3365 1.27512
R11674 gnd.n1684 gnd.n1683 1.27512
R11675 gnd.n4724 gnd.n4716 1.16414
R11676 gnd.n5540 gnd.n4226 1.16414
R11677 gnd.n5477 gnd.n5470 1.16414
R11678 gnd.n5445 gnd.n5438 1.16414
R11679 gnd.n5413 gnd.n5406 1.16414
R11680 gnd.n5382 gnd.n5375 1.16414
R11681 gnd.n5350 gnd.n5343 1.16414
R11682 gnd.n5318 gnd.n5311 1.16414
R11683 gnd.n5286 gnd.n5279 1.16414
R11684 gnd.n5255 gnd.n5248 1.16414
R11685 gnd.n6497 gnd.n6496 0.970197
R11686 gnd.n3869 gnd.n1406 0.970197
R11687 gnd.n5461 gnd.n5429 0.962709
R11688 gnd.n5493 gnd.n5461 0.962709
R11689 gnd.n5334 gnd.n5302 0.962709
R11690 gnd.n5366 gnd.n5334 0.962709
R11691 gnd.n4970 gnd.t210 0.956468
R11692 gnd.n5135 gnd.t294 0.956468
R11693 gnd.n4023 gnd.t195 0.956468
R11694 gnd.n3951 gnd.t31 0.956468
R11695 gnd.n2756 gnd.t29 0.956468
R11696 gnd.n3563 gnd.t321 0.956468
R11697 gnd.n6621 gnd.t2 0.956468
R11698 gnd.n7093 gnd.t200 0.956468
R11699 gnd.n2 gnd.n1 0.672012
R11700 gnd.n3 gnd.n2 0.672012
R11701 gnd.n4 gnd.n3 0.672012
R11702 gnd.n5 gnd.n4 0.672012
R11703 gnd.n6 gnd.n5 0.672012
R11704 gnd.n7 gnd.n6 0.672012
R11705 gnd.n8 gnd.n7 0.672012
R11706 gnd.n9 gnd.n8 0.672012
R11707 gnd.n11 gnd.n10 0.672012
R11708 gnd.n12 gnd.n11 0.672012
R11709 gnd.n13 gnd.n12 0.672012
R11710 gnd.n14 gnd.n13 0.672012
R11711 gnd.n15 gnd.n14 0.672012
R11712 gnd.n16 gnd.n15 0.672012
R11713 gnd.n17 gnd.n16 0.672012
R11714 gnd.n18 gnd.n17 0.672012
R11715 gnd.n2924 gnd.t116 0.637812
R11716 gnd.n2959 gnd.n2958 0.637812
R11717 gnd.n2980 gnd.n2979 0.637812
R11718 gnd.n2992 gnd.t229 0.637812
R11719 gnd.n3095 gnd.n3094 0.637812
R11720 gnd.n3145 gnd.n1824 0.637812
R11721 gnd.t23 gnd.n3268 0.637812
R11722 gnd.n3283 gnd.n3282 0.637812
R11723 gnd.n3303 gnd.n1728 0.637812
R11724 gnd gnd.n0 0.624033
R11725 gnd.n4436 gnd.n4435 0.573776
R11726 gnd.n4435 gnd.n4433 0.573776
R11727 gnd.n4433 gnd.n4431 0.573776
R11728 gnd.n4431 gnd.n4429 0.573776
R11729 gnd.n4429 gnd.n4427 0.573776
R11730 gnd.n4401 gnd.n4400 0.573776
R11731 gnd.n4400 gnd.n4398 0.573776
R11732 gnd.n4398 gnd.n4396 0.573776
R11733 gnd.n4396 gnd.n4394 0.573776
R11734 gnd.n4394 gnd.n4392 0.573776
R11735 gnd.n4412 gnd.n4411 0.573776
R11736 gnd.n4411 gnd.n4409 0.573776
R11737 gnd.n4409 gnd.n4407 0.573776
R11738 gnd.n4407 gnd.n4405 0.573776
R11739 gnd.n4405 gnd.n4403 0.573776
R11740 gnd.n4424 gnd.n4423 0.573776
R11741 gnd.n4423 gnd.n4421 0.573776
R11742 gnd.n4421 gnd.n4419 0.573776
R11743 gnd.n4419 gnd.n4417 0.573776
R11744 gnd.n4417 gnd.n4415 0.573776
R11745 gnd.n58 gnd.n56 0.573776
R11746 gnd.n60 gnd.n58 0.573776
R11747 gnd.n62 gnd.n60 0.573776
R11748 gnd.n64 gnd.n62 0.573776
R11749 gnd.n65 gnd.n64 0.573776
R11750 gnd.n23 gnd.n21 0.573776
R11751 gnd.n25 gnd.n23 0.573776
R11752 gnd.n27 gnd.n25 0.573776
R11753 gnd.n29 gnd.n27 0.573776
R11754 gnd.n30 gnd.n29 0.573776
R11755 gnd.n34 gnd.n32 0.573776
R11756 gnd.n36 gnd.n34 0.573776
R11757 gnd.n38 gnd.n36 0.573776
R11758 gnd.n40 gnd.n38 0.573776
R11759 gnd.n41 gnd.n40 0.573776
R11760 gnd.n46 gnd.n44 0.573776
R11761 gnd.n48 gnd.n46 0.573776
R11762 gnd.n50 gnd.n48 0.573776
R11763 gnd.n52 gnd.n50 0.573776
R11764 gnd.n53 gnd.n52 0.573776
R11765 gnd.n6849 gnd.n6848 0.532512
R11766 gnd.n2367 gnd.n2364 0.532512
R11767 gnd.n6883 gnd.n6882 0.497451
R11768 gnd.n3923 gnd.n3922 0.497451
R11769 gnd.n6551 gnd.n6550 0.497451
R11770 gnd.n1142 gnd.n1065 0.497451
R11771 gnd.n5197 gnd.n4230 0.486781
R11772 gnd.n4773 gnd.n4772 0.48678
R11773 gnd.n5514 gnd.n4184 0.480683
R11774 gnd.n4857 gnd.n4856 0.480683
R11775 gnd.n7130 gnd.n7129 0.4705
R11776 gnd.n6375 gnd.n6374 0.451719
R11777 gnd.n2638 gnd.n2075 0.451719
R11778 gnd.n2632 gnd.n2630 0.451719
R11779 gnd.n6368 gnd.n6367 0.451719
R11780 gnd.n5793 gnd.n838 0.416659
R11781 gnd.n6114 gnd.n6113 0.416659
R11782 gnd.n6328 gnd.n6327 0.416659
R11783 gnd.n2521 gnd.n2520 0.416659
R11784 gnd.n2575 gnd.n2143 0.388379
R11785 gnd.n5474 gnd.n5473 0.388379
R11786 gnd.n5442 gnd.n5441 0.388379
R11787 gnd.n5410 gnd.n5409 0.388379
R11788 gnd.n5379 gnd.n5378 0.388379
R11789 gnd.n5347 gnd.n5346 0.388379
R11790 gnd.n5315 gnd.n5314 0.388379
R11791 gnd.n5283 gnd.n5282 0.388379
R11792 gnd.n5252 gnd.n5251 0.388379
R11793 gnd.n6389 gnd.n443 0.388379
R11794 gnd.n7130 gnd.n19 0.374463
R11795 gnd gnd.n7130 0.367492
R11796 gnd.n4285 gnd.t264 0.319156
R11797 gnd.n3999 gnd.t36 0.319156
R11798 gnd.n3975 gnd.t222 0.319156
R11799 gnd.n6668 gnd.t17 0.319156
R11800 gnd.n7117 gnd.t40 0.319156
R11801 gnd.n4691 gnd.n4669 0.311721
R11802 gnd.n2541 gnd.n2540 0.302329
R11803 gnd.n6376 gnd.n271 0.302329
R11804 gnd.n7064 gnd.n6734 0.293183
R11805 gnd.n4054 gnd.n1129 0.293183
R11806 gnd.n5585 gnd.n5584 0.268793
R11807 gnd.n6435 gnd.n6434 0.258122
R11808 gnd.n7064 gnd.n7063 0.258122
R11809 gnd.n2245 gnd.n2091 0.258122
R11810 gnd.n4055 gnd.n4054 0.258122
R11811 gnd.n5584 gnd.n5583 0.241354
R11812 gnd.n353 gnd.n350 0.229039
R11813 gnd.n354 gnd.n353 0.229039
R11814 gnd.n1408 gnd.n1405 0.229039
R11815 gnd.n2173 gnd.n1408 0.229039
R11816 gnd.n4845 gnd.n4644 0.206293
R11817 gnd.n5491 gnd.n5463 0.155672
R11818 gnd.n5484 gnd.n5463 0.155672
R11819 gnd.n5484 gnd.n5483 0.155672
R11820 gnd.n5483 gnd.n5467 0.155672
R11821 gnd.n5476 gnd.n5467 0.155672
R11822 gnd.n5476 gnd.n5475 0.155672
R11823 gnd.n5459 gnd.n5431 0.155672
R11824 gnd.n5452 gnd.n5431 0.155672
R11825 gnd.n5452 gnd.n5451 0.155672
R11826 gnd.n5451 gnd.n5435 0.155672
R11827 gnd.n5444 gnd.n5435 0.155672
R11828 gnd.n5444 gnd.n5443 0.155672
R11829 gnd.n5427 gnd.n5399 0.155672
R11830 gnd.n5420 gnd.n5399 0.155672
R11831 gnd.n5420 gnd.n5419 0.155672
R11832 gnd.n5419 gnd.n5403 0.155672
R11833 gnd.n5412 gnd.n5403 0.155672
R11834 gnd.n5412 gnd.n5411 0.155672
R11835 gnd.n5396 gnd.n5368 0.155672
R11836 gnd.n5389 gnd.n5368 0.155672
R11837 gnd.n5389 gnd.n5388 0.155672
R11838 gnd.n5388 gnd.n5372 0.155672
R11839 gnd.n5381 gnd.n5372 0.155672
R11840 gnd.n5381 gnd.n5380 0.155672
R11841 gnd.n5364 gnd.n5336 0.155672
R11842 gnd.n5357 gnd.n5336 0.155672
R11843 gnd.n5357 gnd.n5356 0.155672
R11844 gnd.n5356 gnd.n5340 0.155672
R11845 gnd.n5349 gnd.n5340 0.155672
R11846 gnd.n5349 gnd.n5348 0.155672
R11847 gnd.n5332 gnd.n5304 0.155672
R11848 gnd.n5325 gnd.n5304 0.155672
R11849 gnd.n5325 gnd.n5324 0.155672
R11850 gnd.n5324 gnd.n5308 0.155672
R11851 gnd.n5317 gnd.n5308 0.155672
R11852 gnd.n5317 gnd.n5316 0.155672
R11853 gnd.n5300 gnd.n5272 0.155672
R11854 gnd.n5293 gnd.n5272 0.155672
R11855 gnd.n5293 gnd.n5292 0.155672
R11856 gnd.n5292 gnd.n5276 0.155672
R11857 gnd.n5285 gnd.n5276 0.155672
R11858 gnd.n5285 gnd.n5284 0.155672
R11859 gnd.n5269 gnd.n5241 0.155672
R11860 gnd.n5262 gnd.n5241 0.155672
R11861 gnd.n5262 gnd.n5261 0.155672
R11862 gnd.n5261 gnd.n5245 0.155672
R11863 gnd.n5254 gnd.n5245 0.155672
R11864 gnd.n5254 gnd.n5253 0.155672
R11865 gnd.n6550 gnd.n281 0.152939
R11866 gnd.n325 gnd.n281 0.152939
R11867 gnd.n326 gnd.n325 0.152939
R11868 gnd.n327 gnd.n326 0.152939
R11869 gnd.n328 gnd.n327 0.152939
R11870 gnd.n329 gnd.n328 0.152939
R11871 gnd.n330 gnd.n329 0.152939
R11872 gnd.n331 gnd.n330 0.152939
R11873 gnd.n332 gnd.n331 0.152939
R11874 gnd.n333 gnd.n332 0.152939
R11875 gnd.n334 gnd.n333 0.152939
R11876 gnd.n335 gnd.n334 0.152939
R11877 gnd.n336 gnd.n335 0.152939
R11878 gnd.n337 gnd.n336 0.152939
R11879 gnd.n338 gnd.n337 0.152939
R11880 gnd.n339 gnd.n338 0.152939
R11881 gnd.n340 gnd.n339 0.152939
R11882 gnd.n343 gnd.n340 0.152939
R11883 gnd.n344 gnd.n343 0.152939
R11884 gnd.n345 gnd.n344 0.152939
R11885 gnd.n346 gnd.n345 0.152939
R11886 gnd.n347 gnd.n346 0.152939
R11887 gnd.n348 gnd.n347 0.152939
R11888 gnd.n349 gnd.n348 0.152939
R11889 gnd.n350 gnd.n349 0.152939
R11890 gnd.n355 gnd.n354 0.152939
R11891 gnd.n356 gnd.n355 0.152939
R11892 gnd.n357 gnd.n356 0.152939
R11893 gnd.n358 gnd.n357 0.152939
R11894 gnd.n359 gnd.n358 0.152939
R11895 gnd.n360 gnd.n359 0.152939
R11896 gnd.n361 gnd.n360 0.152939
R11897 gnd.n362 gnd.n361 0.152939
R11898 gnd.n363 gnd.n362 0.152939
R11899 gnd.n366 gnd.n363 0.152939
R11900 gnd.n367 gnd.n366 0.152939
R11901 gnd.n368 gnd.n367 0.152939
R11902 gnd.n369 gnd.n368 0.152939
R11903 gnd.n370 gnd.n369 0.152939
R11904 gnd.n371 gnd.n370 0.152939
R11905 gnd.n372 gnd.n371 0.152939
R11906 gnd.n373 gnd.n372 0.152939
R11907 gnd.n374 gnd.n373 0.152939
R11908 gnd.n375 gnd.n374 0.152939
R11909 gnd.n376 gnd.n375 0.152939
R11910 gnd.n377 gnd.n376 0.152939
R11911 gnd.n378 gnd.n377 0.152939
R11912 gnd.n379 gnd.n378 0.152939
R11913 gnd.n380 gnd.n379 0.152939
R11914 gnd.n381 gnd.n380 0.152939
R11915 gnd.n382 gnd.n381 0.152939
R11916 gnd.n383 gnd.n382 0.152939
R11917 gnd.n384 gnd.n383 0.152939
R11918 gnd.n6436 gnd.n384 0.152939
R11919 gnd.n6436 gnd.n6435 0.152939
R11920 gnd.n6553 gnd.n6551 0.152939
R11921 gnd.n6553 gnd.n6552 0.152939
R11922 gnd.n6552 gnd.n252 0.152939
R11923 gnd.n6584 gnd.n252 0.152939
R11924 gnd.n6585 gnd.n6584 0.152939
R11925 gnd.n6586 gnd.n6585 0.152939
R11926 gnd.n6587 gnd.n6586 0.152939
R11927 gnd.n6587 gnd.n226 0.152939
R11928 gnd.n6624 gnd.n226 0.152939
R11929 gnd.n6625 gnd.n6624 0.152939
R11930 gnd.n6626 gnd.n6625 0.152939
R11931 gnd.n6626 gnd.n206 0.152939
R11932 gnd.n6648 gnd.n206 0.152939
R11933 gnd.n6649 gnd.n6648 0.152939
R11934 gnd.n6650 gnd.n6649 0.152939
R11935 gnd.n6651 gnd.n6650 0.152939
R11936 gnd.n99 gnd.n98 0.152939
R11937 gnd.n100 gnd.n99 0.152939
R11938 gnd.n101 gnd.n100 0.152939
R11939 gnd.n118 gnd.n101 0.152939
R11940 gnd.n119 gnd.n118 0.152939
R11941 gnd.n120 gnd.n119 0.152939
R11942 gnd.n121 gnd.n120 0.152939
R11943 gnd.n136 gnd.n121 0.152939
R11944 gnd.n137 gnd.n136 0.152939
R11945 gnd.n138 gnd.n137 0.152939
R11946 gnd.n139 gnd.n138 0.152939
R11947 gnd.n156 gnd.n139 0.152939
R11948 gnd.n157 gnd.n156 0.152939
R11949 gnd.n158 gnd.n157 0.152939
R11950 gnd.n159 gnd.n158 0.152939
R11951 gnd.n6882 gnd.n159 0.152939
R11952 gnd.n7127 gnd.n69 0.152939
R11953 gnd.n6812 gnd.n69 0.152939
R11954 gnd.n6813 gnd.n6812 0.152939
R11955 gnd.n6817 gnd.n6813 0.152939
R11956 gnd.n6818 gnd.n6817 0.152939
R11957 gnd.n6819 gnd.n6818 0.152939
R11958 gnd.n6819 gnd.n6810 0.152939
R11959 gnd.n6825 gnd.n6810 0.152939
R11960 gnd.n6826 gnd.n6825 0.152939
R11961 gnd.n6827 gnd.n6826 0.152939
R11962 gnd.n6827 gnd.n6808 0.152939
R11963 gnd.n6833 gnd.n6808 0.152939
R11964 gnd.n6834 gnd.n6833 0.152939
R11965 gnd.n6835 gnd.n6834 0.152939
R11966 gnd.n6835 gnd.n6806 0.152939
R11967 gnd.n6841 gnd.n6806 0.152939
R11968 gnd.n6842 gnd.n6841 0.152939
R11969 gnd.n6843 gnd.n6842 0.152939
R11970 gnd.n6843 gnd.n6804 0.152939
R11971 gnd.n6848 gnd.n6804 0.152939
R11972 gnd.n6764 gnd.n6734 0.152939
R11973 gnd.n6765 gnd.n6764 0.152939
R11974 gnd.n6765 gnd.n6760 0.152939
R11975 gnd.n6773 gnd.n6760 0.152939
R11976 gnd.n6774 gnd.n6773 0.152939
R11977 gnd.n6775 gnd.n6774 0.152939
R11978 gnd.n6775 gnd.n6758 0.152939
R11979 gnd.n6783 gnd.n6758 0.152939
R11980 gnd.n6784 gnd.n6783 0.152939
R11981 gnd.n6785 gnd.n6784 0.152939
R11982 gnd.n6785 gnd.n6756 0.152939
R11983 gnd.n6793 gnd.n6756 0.152939
R11984 gnd.n6794 gnd.n6793 0.152939
R11985 gnd.n6795 gnd.n6794 0.152939
R11986 gnd.n6795 gnd.n6754 0.152939
R11987 gnd.n6802 gnd.n6754 0.152939
R11988 gnd.n6803 gnd.n6802 0.152939
R11989 gnd.n6849 gnd.n6803 0.152939
R11990 gnd.n7054 gnd.n6883 0.152939
R11991 gnd.n7054 gnd.n7053 0.152939
R11992 gnd.n7053 gnd.n7052 0.152939
R11993 gnd.n7052 gnd.n6885 0.152939
R11994 gnd.n6886 gnd.n6885 0.152939
R11995 gnd.n6887 gnd.n6886 0.152939
R11996 gnd.n6888 gnd.n6887 0.152939
R11997 gnd.n6889 gnd.n6888 0.152939
R11998 gnd.n6890 gnd.n6889 0.152939
R11999 gnd.n6891 gnd.n6890 0.152939
R12000 gnd.n6892 gnd.n6891 0.152939
R12001 gnd.n6893 gnd.n6892 0.152939
R12002 gnd.n6894 gnd.n6893 0.152939
R12003 gnd.n6895 gnd.n6894 0.152939
R12004 gnd.n6896 gnd.n6895 0.152939
R12005 gnd.n6897 gnd.n6896 0.152939
R12006 gnd.n6898 gnd.n6897 0.152939
R12007 gnd.n6899 gnd.n6898 0.152939
R12008 gnd.n6900 gnd.n6899 0.152939
R12009 gnd.n6901 gnd.n6900 0.152939
R12010 gnd.n6902 gnd.n6901 0.152939
R12011 gnd.n6903 gnd.n6902 0.152939
R12012 gnd.n6904 gnd.n6903 0.152939
R12013 gnd.n6905 gnd.n6904 0.152939
R12014 gnd.n6906 gnd.n6905 0.152939
R12015 gnd.n6907 gnd.n6906 0.152939
R12016 gnd.n6908 gnd.n6907 0.152939
R12017 gnd.n6909 gnd.n6908 0.152939
R12018 gnd.n6910 gnd.n6909 0.152939
R12019 gnd.n6911 gnd.n6910 0.152939
R12020 gnd.n6912 gnd.n6911 0.152939
R12021 gnd.n6913 gnd.n6912 0.152939
R12022 gnd.n6914 gnd.n6913 0.152939
R12023 gnd.n6915 gnd.n6914 0.152939
R12024 gnd.n6916 gnd.n6915 0.152939
R12025 gnd.n6917 gnd.n6916 0.152939
R12026 gnd.n6977 gnd.n6917 0.152939
R12027 gnd.n6977 gnd.n6976 0.152939
R12028 gnd.n6976 gnd.n6975 0.152939
R12029 gnd.n6975 gnd.n6921 0.152939
R12030 gnd.n6922 gnd.n6921 0.152939
R12031 gnd.n6923 gnd.n6922 0.152939
R12032 gnd.n6924 gnd.n6923 0.152939
R12033 gnd.n6925 gnd.n6924 0.152939
R12034 gnd.n6926 gnd.n6925 0.152939
R12035 gnd.n6927 gnd.n6926 0.152939
R12036 gnd.n6928 gnd.n6927 0.152939
R12037 gnd.n6929 gnd.n6928 0.152939
R12038 gnd.n6930 gnd.n6929 0.152939
R12039 gnd.n6931 gnd.n6930 0.152939
R12040 gnd.n6932 gnd.n6931 0.152939
R12041 gnd.n6933 gnd.n6932 0.152939
R12042 gnd.n6934 gnd.n6933 0.152939
R12043 gnd.n6935 gnd.n6934 0.152939
R12044 gnd.n6936 gnd.n6935 0.152939
R12045 gnd.n6937 gnd.n6936 0.152939
R12046 gnd.n6937 gnd.n6735 0.152939
R12047 gnd.n7063 gnd.n6735 0.152939
R12048 gnd.n5616 gnd.n4184 0.152939
R12049 gnd.n5616 gnd.n5615 0.152939
R12050 gnd.n5615 gnd.n5614 0.152939
R12051 gnd.n5614 gnd.n4186 0.152939
R12052 gnd.n4187 gnd.n4186 0.152939
R12053 gnd.n4188 gnd.n4187 0.152939
R12054 gnd.n4189 gnd.n4188 0.152939
R12055 gnd.n4190 gnd.n4189 0.152939
R12056 gnd.n4191 gnd.n4190 0.152939
R12057 gnd.n4192 gnd.n4191 0.152939
R12058 gnd.n4193 gnd.n4192 0.152939
R12059 gnd.n4194 gnd.n4193 0.152939
R12060 gnd.n4195 gnd.n4194 0.152939
R12061 gnd.n4196 gnd.n4195 0.152939
R12062 gnd.n5586 gnd.n4196 0.152939
R12063 gnd.n5586 gnd.n5585 0.152939
R12064 gnd.n4858 gnd.n4857 0.152939
R12065 gnd.n4858 gnd.n4562 0.152939
R12066 gnd.n4886 gnd.n4562 0.152939
R12067 gnd.n4887 gnd.n4886 0.152939
R12068 gnd.n4888 gnd.n4887 0.152939
R12069 gnd.n4889 gnd.n4888 0.152939
R12070 gnd.n4889 gnd.n4534 0.152939
R12071 gnd.n4916 gnd.n4534 0.152939
R12072 gnd.n4917 gnd.n4916 0.152939
R12073 gnd.n4918 gnd.n4917 0.152939
R12074 gnd.n4918 gnd.n4512 0.152939
R12075 gnd.n4947 gnd.n4512 0.152939
R12076 gnd.n4948 gnd.n4947 0.152939
R12077 gnd.n4949 gnd.n4948 0.152939
R12078 gnd.n4950 gnd.n4949 0.152939
R12079 gnd.n4952 gnd.n4950 0.152939
R12080 gnd.n4952 gnd.n4951 0.152939
R12081 gnd.n4951 gnd.n4461 0.152939
R12082 gnd.n4462 gnd.n4461 0.152939
R12083 gnd.n4463 gnd.n4462 0.152939
R12084 gnd.n4482 gnd.n4463 0.152939
R12085 gnd.n4483 gnd.n4482 0.152939
R12086 gnd.n4483 gnd.n4381 0.152939
R12087 gnd.n5042 gnd.n4381 0.152939
R12088 gnd.n5043 gnd.n5042 0.152939
R12089 gnd.n5044 gnd.n5043 0.152939
R12090 gnd.n5045 gnd.n5044 0.152939
R12091 gnd.n5045 gnd.n4354 0.152939
R12092 gnd.n5082 gnd.n4354 0.152939
R12093 gnd.n5083 gnd.n5082 0.152939
R12094 gnd.n5084 gnd.n5083 0.152939
R12095 gnd.n5085 gnd.n5084 0.152939
R12096 gnd.n5085 gnd.n4327 0.152939
R12097 gnd.n5127 gnd.n4327 0.152939
R12098 gnd.n5128 gnd.n5127 0.152939
R12099 gnd.n5129 gnd.n5128 0.152939
R12100 gnd.n5130 gnd.n5129 0.152939
R12101 gnd.n5130 gnd.n4299 0.152939
R12102 gnd.n5167 gnd.n4299 0.152939
R12103 gnd.n5168 gnd.n5167 0.152939
R12104 gnd.n5169 gnd.n5168 0.152939
R12105 gnd.n5170 gnd.n5169 0.152939
R12106 gnd.n5170 gnd.n4272 0.152939
R12107 gnd.n5216 gnd.n4272 0.152939
R12108 gnd.n5217 gnd.n5216 0.152939
R12109 gnd.n5218 gnd.n5217 0.152939
R12110 gnd.n5219 gnd.n5218 0.152939
R12111 gnd.n5219 gnd.n4245 0.152939
R12112 gnd.n5510 gnd.n4245 0.152939
R12113 gnd.n5511 gnd.n5510 0.152939
R12114 gnd.n5512 gnd.n5511 0.152939
R12115 gnd.n5513 gnd.n5512 0.152939
R12116 gnd.n5514 gnd.n5513 0.152939
R12117 gnd.n4856 gnd.n4586 0.152939
R12118 gnd.n4607 gnd.n4586 0.152939
R12119 gnd.n4608 gnd.n4607 0.152939
R12120 gnd.n4614 gnd.n4608 0.152939
R12121 gnd.n4615 gnd.n4614 0.152939
R12122 gnd.n4616 gnd.n4615 0.152939
R12123 gnd.n4616 gnd.n4605 0.152939
R12124 gnd.n4624 gnd.n4605 0.152939
R12125 gnd.n4625 gnd.n4624 0.152939
R12126 gnd.n4626 gnd.n4625 0.152939
R12127 gnd.n4626 gnd.n4603 0.152939
R12128 gnd.n4634 gnd.n4603 0.152939
R12129 gnd.n4635 gnd.n4634 0.152939
R12130 gnd.n4636 gnd.n4635 0.152939
R12131 gnd.n4636 gnd.n4601 0.152939
R12132 gnd.n4644 gnd.n4601 0.152939
R12133 gnd.n5583 gnd.n4201 0.152939
R12134 gnd.n4203 gnd.n4201 0.152939
R12135 gnd.n4204 gnd.n4203 0.152939
R12136 gnd.n4205 gnd.n4204 0.152939
R12137 gnd.n4206 gnd.n4205 0.152939
R12138 gnd.n4207 gnd.n4206 0.152939
R12139 gnd.n4208 gnd.n4207 0.152939
R12140 gnd.n4209 gnd.n4208 0.152939
R12141 gnd.n4210 gnd.n4209 0.152939
R12142 gnd.n4211 gnd.n4210 0.152939
R12143 gnd.n4212 gnd.n4211 0.152939
R12144 gnd.n4213 gnd.n4212 0.152939
R12145 gnd.n4214 gnd.n4213 0.152939
R12146 gnd.n4215 gnd.n4214 0.152939
R12147 gnd.n4216 gnd.n4215 0.152939
R12148 gnd.n4217 gnd.n4216 0.152939
R12149 gnd.n4218 gnd.n4217 0.152939
R12150 gnd.n4219 gnd.n4218 0.152939
R12151 gnd.n4220 gnd.n4219 0.152939
R12152 gnd.n4221 gnd.n4220 0.152939
R12153 gnd.n4222 gnd.n4221 0.152939
R12154 gnd.n4223 gnd.n4222 0.152939
R12155 gnd.n4227 gnd.n4223 0.152939
R12156 gnd.n4228 gnd.n4227 0.152939
R12157 gnd.n4229 gnd.n4228 0.152939
R12158 gnd.n4230 gnd.n4229 0.152939
R12159 gnd.n5019 gnd.n5018 0.152939
R12160 gnd.n5020 gnd.n5019 0.152939
R12161 gnd.n5021 gnd.n5020 0.152939
R12162 gnd.n5022 gnd.n5021 0.152939
R12163 gnd.n5023 gnd.n5022 0.152939
R12164 gnd.n5024 gnd.n5023 0.152939
R12165 gnd.n5024 gnd.n4335 0.152939
R12166 gnd.n5103 gnd.n4335 0.152939
R12167 gnd.n5104 gnd.n5103 0.152939
R12168 gnd.n5105 gnd.n5104 0.152939
R12169 gnd.n5106 gnd.n5105 0.152939
R12170 gnd.n5107 gnd.n5106 0.152939
R12171 gnd.n5108 gnd.n5107 0.152939
R12172 gnd.n5109 gnd.n5108 0.152939
R12173 gnd.n5110 gnd.n5109 0.152939
R12174 gnd.n5111 gnd.n5110 0.152939
R12175 gnd.n5111 gnd.n4279 0.152939
R12176 gnd.n5188 gnd.n4279 0.152939
R12177 gnd.n5189 gnd.n5188 0.152939
R12178 gnd.n5190 gnd.n5189 0.152939
R12179 gnd.n5191 gnd.n5190 0.152939
R12180 gnd.n5192 gnd.n5191 0.152939
R12181 gnd.n5193 gnd.n5192 0.152939
R12182 gnd.n5194 gnd.n5193 0.152939
R12183 gnd.n5195 gnd.n5194 0.152939
R12184 gnd.n5196 gnd.n5195 0.152939
R12185 gnd.n5198 gnd.n5196 0.152939
R12186 gnd.n5198 gnd.n5197 0.152939
R12187 gnd.n4774 gnd.n4773 0.152939
R12188 gnd.n4774 gnd.n4664 0.152939
R12189 gnd.n4789 gnd.n4664 0.152939
R12190 gnd.n4790 gnd.n4789 0.152939
R12191 gnd.n4791 gnd.n4790 0.152939
R12192 gnd.n4791 gnd.n4652 0.152939
R12193 gnd.n4805 gnd.n4652 0.152939
R12194 gnd.n4806 gnd.n4805 0.152939
R12195 gnd.n4807 gnd.n4806 0.152939
R12196 gnd.n4808 gnd.n4807 0.152939
R12197 gnd.n4809 gnd.n4808 0.152939
R12198 gnd.n4810 gnd.n4809 0.152939
R12199 gnd.n4811 gnd.n4810 0.152939
R12200 gnd.n4812 gnd.n4811 0.152939
R12201 gnd.n4813 gnd.n4812 0.152939
R12202 gnd.n4814 gnd.n4813 0.152939
R12203 gnd.n4815 gnd.n4814 0.152939
R12204 gnd.n4816 gnd.n4815 0.152939
R12205 gnd.n4817 gnd.n4816 0.152939
R12206 gnd.n4818 gnd.n4817 0.152939
R12207 gnd.n4819 gnd.n4818 0.152939
R12208 gnd.n4819 gnd.n4518 0.152939
R12209 gnd.n4936 gnd.n4518 0.152939
R12210 gnd.n4937 gnd.n4936 0.152939
R12211 gnd.n4938 gnd.n4937 0.152939
R12212 gnd.n4939 gnd.n4938 0.152939
R12213 gnd.n4939 gnd.n4440 0.152939
R12214 gnd.n5016 gnd.n4440 0.152939
R12215 gnd.n4692 gnd.n4691 0.152939
R12216 gnd.n4693 gnd.n4692 0.152939
R12217 gnd.n4694 gnd.n4693 0.152939
R12218 gnd.n4695 gnd.n4694 0.152939
R12219 gnd.n4696 gnd.n4695 0.152939
R12220 gnd.n4697 gnd.n4696 0.152939
R12221 gnd.n4698 gnd.n4697 0.152939
R12222 gnd.n4699 gnd.n4698 0.152939
R12223 gnd.n4700 gnd.n4699 0.152939
R12224 gnd.n4701 gnd.n4700 0.152939
R12225 gnd.n4702 gnd.n4701 0.152939
R12226 gnd.n4703 gnd.n4702 0.152939
R12227 gnd.n4704 gnd.n4703 0.152939
R12228 gnd.n4705 gnd.n4704 0.152939
R12229 gnd.n4706 gnd.n4705 0.152939
R12230 gnd.n4707 gnd.n4706 0.152939
R12231 gnd.n4708 gnd.n4707 0.152939
R12232 gnd.n4709 gnd.n4708 0.152939
R12233 gnd.n4710 gnd.n4709 0.152939
R12234 gnd.n4711 gnd.n4710 0.152939
R12235 gnd.n4712 gnd.n4711 0.152939
R12236 gnd.n4713 gnd.n4712 0.152939
R12237 gnd.n4717 gnd.n4713 0.152939
R12238 gnd.n4718 gnd.n4717 0.152939
R12239 gnd.n4718 gnd.n4675 0.152939
R12240 gnd.n4772 gnd.n4675 0.152939
R12241 gnd.n2368 gnd.n2367 0.152939
R12242 gnd.n2369 gnd.n2368 0.152939
R12243 gnd.n2369 gnd.n2307 0.152939
R12244 gnd.n2375 gnd.n2307 0.152939
R12245 gnd.n2376 gnd.n2375 0.152939
R12246 gnd.n2377 gnd.n2376 0.152939
R12247 gnd.n2377 gnd.n2305 0.152939
R12248 gnd.n2383 gnd.n2305 0.152939
R12249 gnd.n2384 gnd.n2383 0.152939
R12250 gnd.n2385 gnd.n2384 0.152939
R12251 gnd.n2385 gnd.n2303 0.152939
R12252 gnd.n2391 gnd.n2303 0.152939
R12253 gnd.n2392 gnd.n2391 0.152939
R12254 gnd.n2393 gnd.n2392 0.152939
R12255 gnd.n2393 gnd.n2301 0.152939
R12256 gnd.n2399 gnd.n2301 0.152939
R12257 gnd.n2400 gnd.n2399 0.152939
R12258 gnd.n2401 gnd.n2400 0.152939
R12259 gnd.n2401 gnd.n2299 0.152939
R12260 gnd.n2407 gnd.n2299 0.152939
R12261 gnd.n3922 gnd.n1336 0.152939
R12262 gnd.n1380 gnd.n1336 0.152939
R12263 gnd.n1381 gnd.n1380 0.152939
R12264 gnd.n1382 gnd.n1381 0.152939
R12265 gnd.n1383 gnd.n1382 0.152939
R12266 gnd.n1384 gnd.n1383 0.152939
R12267 gnd.n1385 gnd.n1384 0.152939
R12268 gnd.n1386 gnd.n1385 0.152939
R12269 gnd.n1387 gnd.n1386 0.152939
R12270 gnd.n1388 gnd.n1387 0.152939
R12271 gnd.n1389 gnd.n1388 0.152939
R12272 gnd.n1390 gnd.n1389 0.152939
R12273 gnd.n1391 gnd.n1390 0.152939
R12274 gnd.n1392 gnd.n1391 0.152939
R12275 gnd.n1393 gnd.n1392 0.152939
R12276 gnd.n1394 gnd.n1393 0.152939
R12277 gnd.n1395 gnd.n1394 0.152939
R12278 gnd.n1398 gnd.n1395 0.152939
R12279 gnd.n1399 gnd.n1398 0.152939
R12280 gnd.n1400 gnd.n1399 0.152939
R12281 gnd.n1401 gnd.n1400 0.152939
R12282 gnd.n1402 gnd.n1401 0.152939
R12283 gnd.n1403 gnd.n1402 0.152939
R12284 gnd.n1404 gnd.n1403 0.152939
R12285 gnd.n1405 gnd.n1404 0.152939
R12286 gnd.n2174 gnd.n2173 0.152939
R12287 gnd.n2175 gnd.n2174 0.152939
R12288 gnd.n2175 gnd.n2169 0.152939
R12289 gnd.n2183 gnd.n2169 0.152939
R12290 gnd.n2184 gnd.n2183 0.152939
R12291 gnd.n2185 gnd.n2184 0.152939
R12292 gnd.n2185 gnd.n2167 0.152939
R12293 gnd.n2193 gnd.n2167 0.152939
R12294 gnd.n2194 gnd.n2193 0.152939
R12295 gnd.n2195 gnd.n2194 0.152939
R12296 gnd.n2195 gnd.n2163 0.152939
R12297 gnd.n2203 gnd.n2163 0.152939
R12298 gnd.n2204 gnd.n2203 0.152939
R12299 gnd.n2205 gnd.n2204 0.152939
R12300 gnd.n2205 gnd.n2161 0.152939
R12301 gnd.n2213 gnd.n2161 0.152939
R12302 gnd.n2214 gnd.n2213 0.152939
R12303 gnd.n2215 gnd.n2214 0.152939
R12304 gnd.n2215 gnd.n2159 0.152939
R12305 gnd.n2223 gnd.n2159 0.152939
R12306 gnd.n2224 gnd.n2223 0.152939
R12307 gnd.n2225 gnd.n2224 0.152939
R12308 gnd.n2225 gnd.n2157 0.152939
R12309 gnd.n2233 gnd.n2157 0.152939
R12310 gnd.n2234 gnd.n2233 0.152939
R12311 gnd.n2235 gnd.n2234 0.152939
R12312 gnd.n2235 gnd.n2155 0.152939
R12313 gnd.n2243 gnd.n2155 0.152939
R12314 gnd.n2244 gnd.n2243 0.152939
R12315 gnd.n2245 gnd.n2244 0.152939
R12316 gnd.n1258 gnd.n1257 0.152939
R12317 gnd.n1274 gnd.n1258 0.152939
R12318 gnd.n1275 gnd.n1274 0.152939
R12319 gnd.n1276 gnd.n1275 0.152939
R12320 gnd.n1277 gnd.n1276 0.152939
R12321 gnd.n1293 gnd.n1277 0.152939
R12322 gnd.n1294 gnd.n1293 0.152939
R12323 gnd.n1295 gnd.n1294 0.152939
R12324 gnd.n1296 gnd.n1295 0.152939
R12325 gnd.n1314 gnd.n1296 0.152939
R12326 gnd.n1315 gnd.n1314 0.152939
R12327 gnd.n1316 gnd.n1315 0.152939
R12328 gnd.n1317 gnd.n1316 0.152939
R12329 gnd.n1334 gnd.n1317 0.152939
R12330 gnd.n1335 gnd.n1334 0.152939
R12331 gnd.n3923 gnd.n1335 0.152939
R12332 gnd.n4046 gnd.n1142 0.152939
R12333 gnd.n4046 gnd.n4045 0.152939
R12334 gnd.n4045 gnd.n4044 0.152939
R12335 gnd.n4044 gnd.n1143 0.152939
R12336 gnd.n1161 gnd.n1143 0.152939
R12337 gnd.n1162 gnd.n1161 0.152939
R12338 gnd.n1163 gnd.n1162 0.152939
R12339 gnd.n1178 gnd.n1163 0.152939
R12340 gnd.n1179 gnd.n1178 0.152939
R12341 gnd.n1180 gnd.n1179 0.152939
R12342 gnd.n1181 gnd.n1180 0.152939
R12343 gnd.n1198 gnd.n1181 0.152939
R12344 gnd.n1199 gnd.n1198 0.152939
R12345 gnd.n1200 gnd.n1199 0.152939
R12346 gnd.n1201 gnd.n1200 0.152939
R12347 gnd.n1216 gnd.n1201 0.152939
R12348 gnd.n1066 gnd.n1065 0.152939
R12349 gnd.n1067 gnd.n1066 0.152939
R12350 gnd.n1068 gnd.n1067 0.152939
R12351 gnd.n1069 gnd.n1068 0.152939
R12352 gnd.n1070 gnd.n1069 0.152939
R12353 gnd.n1071 gnd.n1070 0.152939
R12354 gnd.n1072 gnd.n1071 0.152939
R12355 gnd.n1073 gnd.n1072 0.152939
R12356 gnd.n1074 gnd.n1073 0.152939
R12357 gnd.n1075 gnd.n1074 0.152939
R12358 gnd.n1076 gnd.n1075 0.152939
R12359 gnd.n1077 gnd.n1076 0.152939
R12360 gnd.n1078 gnd.n1077 0.152939
R12361 gnd.n1079 gnd.n1078 0.152939
R12362 gnd.n1080 gnd.n1079 0.152939
R12363 gnd.n1081 gnd.n1080 0.152939
R12364 gnd.n1082 gnd.n1081 0.152939
R12365 gnd.n1085 gnd.n1082 0.152939
R12366 gnd.n1086 gnd.n1085 0.152939
R12367 gnd.n1087 gnd.n1086 0.152939
R12368 gnd.n1088 gnd.n1087 0.152939
R12369 gnd.n1089 gnd.n1088 0.152939
R12370 gnd.n1090 gnd.n1089 0.152939
R12371 gnd.n1091 gnd.n1090 0.152939
R12372 gnd.n1092 gnd.n1091 0.152939
R12373 gnd.n1093 gnd.n1092 0.152939
R12374 gnd.n1094 gnd.n1093 0.152939
R12375 gnd.n1095 gnd.n1094 0.152939
R12376 gnd.n1096 gnd.n1095 0.152939
R12377 gnd.n1097 gnd.n1096 0.152939
R12378 gnd.n1098 gnd.n1097 0.152939
R12379 gnd.n1099 gnd.n1098 0.152939
R12380 gnd.n1100 gnd.n1099 0.152939
R12381 gnd.n1101 gnd.n1100 0.152939
R12382 gnd.n1102 gnd.n1101 0.152939
R12383 gnd.n1103 gnd.n1102 0.152939
R12384 gnd.n1104 gnd.n1103 0.152939
R12385 gnd.n1107 gnd.n1104 0.152939
R12386 gnd.n1108 gnd.n1107 0.152939
R12387 gnd.n1109 gnd.n1108 0.152939
R12388 gnd.n1110 gnd.n1109 0.152939
R12389 gnd.n1111 gnd.n1110 0.152939
R12390 gnd.n1112 gnd.n1111 0.152939
R12391 gnd.n1113 gnd.n1112 0.152939
R12392 gnd.n1114 gnd.n1113 0.152939
R12393 gnd.n1115 gnd.n1114 0.152939
R12394 gnd.n1116 gnd.n1115 0.152939
R12395 gnd.n1117 gnd.n1116 0.152939
R12396 gnd.n1118 gnd.n1117 0.152939
R12397 gnd.n1119 gnd.n1118 0.152939
R12398 gnd.n1120 gnd.n1119 0.152939
R12399 gnd.n1121 gnd.n1120 0.152939
R12400 gnd.n1122 gnd.n1121 0.152939
R12401 gnd.n1123 gnd.n1122 0.152939
R12402 gnd.n1124 gnd.n1123 0.152939
R12403 gnd.n1125 gnd.n1124 0.152939
R12404 gnd.n4056 gnd.n1125 0.152939
R12405 gnd.n4056 gnd.n4055 0.152939
R12406 gnd.n2322 gnd.n1129 0.152939
R12407 gnd.n2328 gnd.n2322 0.152939
R12408 gnd.n2329 gnd.n2328 0.152939
R12409 gnd.n2330 gnd.n2329 0.152939
R12410 gnd.n2330 gnd.n2320 0.152939
R12411 gnd.n2338 gnd.n2320 0.152939
R12412 gnd.n2339 gnd.n2338 0.152939
R12413 gnd.n2340 gnd.n2339 0.152939
R12414 gnd.n2340 gnd.n2318 0.152939
R12415 gnd.n2348 gnd.n2318 0.152939
R12416 gnd.n2349 gnd.n2348 0.152939
R12417 gnd.n2350 gnd.n2349 0.152939
R12418 gnd.n2350 gnd.n2316 0.152939
R12419 gnd.n2358 gnd.n2316 0.152939
R12420 gnd.n2359 gnd.n2358 0.152939
R12421 gnd.n2360 gnd.n2359 0.152939
R12422 gnd.n2360 gnd.n2309 0.152939
R12423 gnd.n2364 gnd.n2309 0.152939
R12424 gnd.n5794 gnd.n5793 0.152939
R12425 gnd.n5795 gnd.n5794 0.152939
R12426 gnd.n5795 gnd.n832 0.152939
R12427 gnd.n5803 gnd.n832 0.152939
R12428 gnd.n5804 gnd.n5803 0.152939
R12429 gnd.n5805 gnd.n5804 0.152939
R12430 gnd.n5805 gnd.n826 0.152939
R12431 gnd.n5813 gnd.n826 0.152939
R12432 gnd.n5814 gnd.n5813 0.152939
R12433 gnd.n5815 gnd.n5814 0.152939
R12434 gnd.n5815 gnd.n820 0.152939
R12435 gnd.n5823 gnd.n820 0.152939
R12436 gnd.n5824 gnd.n5823 0.152939
R12437 gnd.n5825 gnd.n5824 0.152939
R12438 gnd.n5825 gnd.n814 0.152939
R12439 gnd.n5833 gnd.n814 0.152939
R12440 gnd.n5834 gnd.n5833 0.152939
R12441 gnd.n5835 gnd.n5834 0.152939
R12442 gnd.n5835 gnd.n808 0.152939
R12443 gnd.n5843 gnd.n808 0.152939
R12444 gnd.n5844 gnd.n5843 0.152939
R12445 gnd.n5845 gnd.n5844 0.152939
R12446 gnd.n5845 gnd.n802 0.152939
R12447 gnd.n5853 gnd.n802 0.152939
R12448 gnd.n5854 gnd.n5853 0.152939
R12449 gnd.n5855 gnd.n5854 0.152939
R12450 gnd.n5855 gnd.n796 0.152939
R12451 gnd.n5863 gnd.n796 0.152939
R12452 gnd.n5864 gnd.n5863 0.152939
R12453 gnd.n5865 gnd.n5864 0.152939
R12454 gnd.n5865 gnd.n790 0.152939
R12455 gnd.n5873 gnd.n790 0.152939
R12456 gnd.n5874 gnd.n5873 0.152939
R12457 gnd.n5875 gnd.n5874 0.152939
R12458 gnd.n5875 gnd.n784 0.152939
R12459 gnd.n5883 gnd.n784 0.152939
R12460 gnd.n5884 gnd.n5883 0.152939
R12461 gnd.n5885 gnd.n5884 0.152939
R12462 gnd.n5885 gnd.n778 0.152939
R12463 gnd.n5893 gnd.n778 0.152939
R12464 gnd.n5894 gnd.n5893 0.152939
R12465 gnd.n5895 gnd.n5894 0.152939
R12466 gnd.n5895 gnd.n772 0.152939
R12467 gnd.n5903 gnd.n772 0.152939
R12468 gnd.n5904 gnd.n5903 0.152939
R12469 gnd.n5905 gnd.n5904 0.152939
R12470 gnd.n5905 gnd.n766 0.152939
R12471 gnd.n5913 gnd.n766 0.152939
R12472 gnd.n5914 gnd.n5913 0.152939
R12473 gnd.n5915 gnd.n5914 0.152939
R12474 gnd.n5915 gnd.n760 0.152939
R12475 gnd.n5923 gnd.n760 0.152939
R12476 gnd.n5924 gnd.n5923 0.152939
R12477 gnd.n5925 gnd.n5924 0.152939
R12478 gnd.n5925 gnd.n754 0.152939
R12479 gnd.n5933 gnd.n754 0.152939
R12480 gnd.n5934 gnd.n5933 0.152939
R12481 gnd.n5935 gnd.n5934 0.152939
R12482 gnd.n5935 gnd.n748 0.152939
R12483 gnd.n5943 gnd.n748 0.152939
R12484 gnd.n5944 gnd.n5943 0.152939
R12485 gnd.n5945 gnd.n5944 0.152939
R12486 gnd.n5945 gnd.n742 0.152939
R12487 gnd.n5953 gnd.n742 0.152939
R12488 gnd.n5954 gnd.n5953 0.152939
R12489 gnd.n5955 gnd.n5954 0.152939
R12490 gnd.n5955 gnd.n736 0.152939
R12491 gnd.n5963 gnd.n736 0.152939
R12492 gnd.n5964 gnd.n5963 0.152939
R12493 gnd.n5965 gnd.n5964 0.152939
R12494 gnd.n5965 gnd.n730 0.152939
R12495 gnd.n5973 gnd.n730 0.152939
R12496 gnd.n5974 gnd.n5973 0.152939
R12497 gnd.n5975 gnd.n5974 0.152939
R12498 gnd.n5975 gnd.n724 0.152939
R12499 gnd.n5983 gnd.n724 0.152939
R12500 gnd.n5984 gnd.n5983 0.152939
R12501 gnd.n5985 gnd.n5984 0.152939
R12502 gnd.n5985 gnd.n718 0.152939
R12503 gnd.n5993 gnd.n718 0.152939
R12504 gnd.n5994 gnd.n5993 0.152939
R12505 gnd.n5995 gnd.n5994 0.152939
R12506 gnd.n5995 gnd.n712 0.152939
R12507 gnd.n6003 gnd.n712 0.152939
R12508 gnd.n6004 gnd.n6003 0.152939
R12509 gnd.n6005 gnd.n6004 0.152939
R12510 gnd.n6005 gnd.n706 0.152939
R12511 gnd.n6013 gnd.n706 0.152939
R12512 gnd.n6014 gnd.n6013 0.152939
R12513 gnd.n6015 gnd.n6014 0.152939
R12514 gnd.n6015 gnd.n700 0.152939
R12515 gnd.n6023 gnd.n700 0.152939
R12516 gnd.n6024 gnd.n6023 0.152939
R12517 gnd.n6025 gnd.n6024 0.152939
R12518 gnd.n6025 gnd.n694 0.152939
R12519 gnd.n6033 gnd.n694 0.152939
R12520 gnd.n6034 gnd.n6033 0.152939
R12521 gnd.n6035 gnd.n6034 0.152939
R12522 gnd.n6035 gnd.n688 0.152939
R12523 gnd.n6043 gnd.n688 0.152939
R12524 gnd.n6044 gnd.n6043 0.152939
R12525 gnd.n6045 gnd.n6044 0.152939
R12526 gnd.n6045 gnd.n682 0.152939
R12527 gnd.n6053 gnd.n682 0.152939
R12528 gnd.n6054 gnd.n6053 0.152939
R12529 gnd.n6055 gnd.n6054 0.152939
R12530 gnd.n6055 gnd.n676 0.152939
R12531 gnd.n6063 gnd.n676 0.152939
R12532 gnd.n6064 gnd.n6063 0.152939
R12533 gnd.n6065 gnd.n6064 0.152939
R12534 gnd.n6065 gnd.n670 0.152939
R12535 gnd.n6073 gnd.n670 0.152939
R12536 gnd.n6074 gnd.n6073 0.152939
R12537 gnd.n6075 gnd.n6074 0.152939
R12538 gnd.n6075 gnd.n664 0.152939
R12539 gnd.n6083 gnd.n664 0.152939
R12540 gnd.n6084 gnd.n6083 0.152939
R12541 gnd.n6085 gnd.n6084 0.152939
R12542 gnd.n6085 gnd.n658 0.152939
R12543 gnd.n6093 gnd.n658 0.152939
R12544 gnd.n6094 gnd.n6093 0.152939
R12545 gnd.n6095 gnd.n6094 0.152939
R12546 gnd.n6095 gnd.n652 0.152939
R12547 gnd.n6103 gnd.n652 0.152939
R12548 gnd.n6104 gnd.n6103 0.152939
R12549 gnd.n6105 gnd.n6104 0.152939
R12550 gnd.n6105 gnd.n646 0.152939
R12551 gnd.n6113 gnd.n646 0.152939
R12552 gnd.n6115 gnd.n6114 0.152939
R12553 gnd.n6115 gnd.n640 0.152939
R12554 gnd.n6123 gnd.n640 0.152939
R12555 gnd.n6124 gnd.n6123 0.152939
R12556 gnd.n6125 gnd.n6124 0.152939
R12557 gnd.n6125 gnd.n634 0.152939
R12558 gnd.n6133 gnd.n634 0.152939
R12559 gnd.n6134 gnd.n6133 0.152939
R12560 gnd.n6135 gnd.n6134 0.152939
R12561 gnd.n6135 gnd.n628 0.152939
R12562 gnd.n6143 gnd.n628 0.152939
R12563 gnd.n6144 gnd.n6143 0.152939
R12564 gnd.n6145 gnd.n6144 0.152939
R12565 gnd.n6145 gnd.n622 0.152939
R12566 gnd.n6153 gnd.n622 0.152939
R12567 gnd.n6154 gnd.n6153 0.152939
R12568 gnd.n6155 gnd.n6154 0.152939
R12569 gnd.n6155 gnd.n616 0.152939
R12570 gnd.n6163 gnd.n616 0.152939
R12571 gnd.n6164 gnd.n6163 0.152939
R12572 gnd.n6165 gnd.n6164 0.152939
R12573 gnd.n6165 gnd.n610 0.152939
R12574 gnd.n6173 gnd.n610 0.152939
R12575 gnd.n6174 gnd.n6173 0.152939
R12576 gnd.n6175 gnd.n6174 0.152939
R12577 gnd.n6175 gnd.n604 0.152939
R12578 gnd.n6183 gnd.n604 0.152939
R12579 gnd.n6184 gnd.n6183 0.152939
R12580 gnd.n6185 gnd.n6184 0.152939
R12581 gnd.n6185 gnd.n598 0.152939
R12582 gnd.n6193 gnd.n598 0.152939
R12583 gnd.n6194 gnd.n6193 0.152939
R12584 gnd.n6195 gnd.n6194 0.152939
R12585 gnd.n6195 gnd.n592 0.152939
R12586 gnd.n6203 gnd.n592 0.152939
R12587 gnd.n6204 gnd.n6203 0.152939
R12588 gnd.n6205 gnd.n6204 0.152939
R12589 gnd.n6205 gnd.n586 0.152939
R12590 gnd.n6213 gnd.n586 0.152939
R12591 gnd.n6214 gnd.n6213 0.152939
R12592 gnd.n6215 gnd.n6214 0.152939
R12593 gnd.n6215 gnd.n580 0.152939
R12594 gnd.n6223 gnd.n580 0.152939
R12595 gnd.n6224 gnd.n6223 0.152939
R12596 gnd.n6225 gnd.n6224 0.152939
R12597 gnd.n6225 gnd.n574 0.152939
R12598 gnd.n6233 gnd.n574 0.152939
R12599 gnd.n6234 gnd.n6233 0.152939
R12600 gnd.n6235 gnd.n6234 0.152939
R12601 gnd.n6235 gnd.n568 0.152939
R12602 gnd.n6243 gnd.n568 0.152939
R12603 gnd.n6244 gnd.n6243 0.152939
R12604 gnd.n6245 gnd.n6244 0.152939
R12605 gnd.n6245 gnd.n562 0.152939
R12606 gnd.n6253 gnd.n562 0.152939
R12607 gnd.n6254 gnd.n6253 0.152939
R12608 gnd.n6255 gnd.n6254 0.152939
R12609 gnd.n6255 gnd.n556 0.152939
R12610 gnd.n6263 gnd.n556 0.152939
R12611 gnd.n6264 gnd.n6263 0.152939
R12612 gnd.n6265 gnd.n6264 0.152939
R12613 gnd.n6265 gnd.n550 0.152939
R12614 gnd.n6273 gnd.n550 0.152939
R12615 gnd.n6274 gnd.n6273 0.152939
R12616 gnd.n6275 gnd.n6274 0.152939
R12617 gnd.n6275 gnd.n544 0.152939
R12618 gnd.n6283 gnd.n544 0.152939
R12619 gnd.n6284 gnd.n6283 0.152939
R12620 gnd.n6285 gnd.n6284 0.152939
R12621 gnd.n6285 gnd.n538 0.152939
R12622 gnd.n6293 gnd.n538 0.152939
R12623 gnd.n6294 gnd.n6293 0.152939
R12624 gnd.n6295 gnd.n6294 0.152939
R12625 gnd.n6295 gnd.n532 0.152939
R12626 gnd.n6303 gnd.n532 0.152939
R12627 gnd.n6304 gnd.n6303 0.152939
R12628 gnd.n6305 gnd.n6304 0.152939
R12629 gnd.n6305 gnd.n526 0.152939
R12630 gnd.n6313 gnd.n526 0.152939
R12631 gnd.n6314 gnd.n6313 0.152939
R12632 gnd.n6315 gnd.n6314 0.152939
R12633 gnd.n6316 gnd.n6315 0.152939
R12634 gnd.n6316 gnd.n520 0.152939
R12635 gnd.n6327 gnd.n520 0.152939
R12636 gnd.n2522 gnd.n2521 0.152939
R12637 gnd.n2522 gnd.n2516 0.152939
R12638 gnd.n2528 gnd.n2516 0.152939
R12639 gnd.n2529 gnd.n2528 0.152939
R12640 gnd.n2531 gnd.n2529 0.152939
R12641 gnd.n2531 gnd.n2530 0.152939
R12642 gnd.n2530 gnd.n2252 0.152939
R12643 gnd.n2253 gnd.n2252 0.152939
R12644 gnd.n2254 gnd.n2253 0.152939
R12645 gnd.n2548 gnd.n2254 0.152939
R12646 gnd.n2549 gnd.n2548 0.152939
R12647 gnd.n2550 gnd.n2549 0.152939
R12648 gnd.n2551 gnd.n2550 0.152939
R12649 gnd.n2551 gnd.n2068 0.152939
R12650 gnd.n2648 gnd.n2068 0.152939
R12651 gnd.n2649 gnd.n2648 0.152939
R12652 gnd.n2650 gnd.n2649 0.152939
R12653 gnd.n2651 gnd.n2650 0.152939
R12654 gnd.n2651 gnd.n2043 0.152939
R12655 gnd.n2678 gnd.n2043 0.152939
R12656 gnd.n2679 gnd.n2678 0.152939
R12657 gnd.n2680 gnd.n2679 0.152939
R12658 gnd.n2681 gnd.n2680 0.152939
R12659 gnd.n2681 gnd.n2018 0.152939
R12660 gnd.n2708 gnd.n2018 0.152939
R12661 gnd.n2709 gnd.n2708 0.152939
R12662 gnd.n2710 gnd.n2709 0.152939
R12663 gnd.n2711 gnd.n2710 0.152939
R12664 gnd.n2711 gnd.n1993 0.152939
R12665 gnd.n2742 gnd.n1993 0.152939
R12666 gnd.n2743 gnd.n2742 0.152939
R12667 gnd.n2744 gnd.n2743 0.152939
R12668 gnd.n2745 gnd.n2744 0.152939
R12669 gnd.n2746 gnd.n2745 0.152939
R12670 gnd.n2749 gnd.n2746 0.152939
R12671 gnd.n2750 gnd.n2749 0.152939
R12672 gnd.n2751 gnd.n2750 0.152939
R12673 gnd.n2751 gnd.n1962 0.152939
R12674 gnd.n2916 gnd.n1962 0.152939
R12675 gnd.n2917 gnd.n2916 0.152939
R12676 gnd.n2918 gnd.n2917 0.152939
R12677 gnd.n2919 gnd.n2918 0.152939
R12678 gnd.n2919 gnd.n1935 0.152939
R12679 gnd.n2953 gnd.n1935 0.152939
R12680 gnd.n2954 gnd.n2953 0.152939
R12681 gnd.n2955 gnd.n2954 0.152939
R12682 gnd.n2955 gnd.n1914 0.152939
R12683 gnd.n2983 gnd.n1914 0.152939
R12684 gnd.n2984 gnd.n2983 0.152939
R12685 gnd.n2985 gnd.n2984 0.152939
R12686 gnd.n2986 gnd.n2985 0.152939
R12687 gnd.n2986 gnd.n1884 0.152939
R12688 gnd.n3034 gnd.n1884 0.152939
R12689 gnd.n3035 gnd.n3034 0.152939
R12690 gnd.n3036 gnd.n3035 0.152939
R12691 gnd.n3037 gnd.n3036 0.152939
R12692 gnd.n3037 gnd.n1865 0.152939
R12693 gnd.n3062 gnd.n1865 0.152939
R12694 gnd.n3063 gnd.n3062 0.152939
R12695 gnd.n3064 gnd.n3063 0.152939
R12696 gnd.n3064 gnd.n1837 0.152939
R12697 gnd.n3118 gnd.n1837 0.152939
R12698 gnd.n3119 gnd.n3118 0.152939
R12699 gnd.n3120 gnd.n3119 0.152939
R12700 gnd.n3120 gnd.n1814 0.152939
R12701 gnd.n3158 gnd.n1814 0.152939
R12702 gnd.n3159 gnd.n3158 0.152939
R12703 gnd.n3160 gnd.n3159 0.152939
R12704 gnd.n3160 gnd.n1791 0.152939
R12705 gnd.n3198 gnd.n1791 0.152939
R12706 gnd.n3199 gnd.n3198 0.152939
R12707 gnd.n3200 gnd.n3199 0.152939
R12708 gnd.n3200 gnd.n1769 0.152939
R12709 gnd.n3245 gnd.n1769 0.152939
R12710 gnd.n3246 gnd.n3245 0.152939
R12711 gnd.n3247 gnd.n3246 0.152939
R12712 gnd.n3247 gnd.n1751 0.152939
R12713 gnd.n3272 gnd.n1751 0.152939
R12714 gnd.n3273 gnd.n3272 0.152939
R12715 gnd.n3274 gnd.n3273 0.152939
R12716 gnd.n3275 gnd.n3274 0.152939
R12717 gnd.n3276 gnd.n3275 0.152939
R12718 gnd.n3276 gnd.n1715 0.152939
R12719 gnd.n3339 gnd.n1715 0.152939
R12720 gnd.n3340 gnd.n3339 0.152939
R12721 gnd.n3341 gnd.n3340 0.152939
R12722 gnd.n3342 gnd.n3341 0.152939
R12723 gnd.n3342 gnd.n1688 0.152939
R12724 gnd.n3390 gnd.n1688 0.152939
R12725 gnd.n3391 gnd.n3390 0.152939
R12726 gnd.n3392 gnd.n3391 0.152939
R12727 gnd.n3393 gnd.n3392 0.152939
R12728 gnd.n3394 gnd.n3393 0.152939
R12729 gnd.n3394 gnd.n1627 0.152939
R12730 gnd.n3578 gnd.n1627 0.152939
R12731 gnd.n3579 gnd.n3578 0.152939
R12732 gnd.n3580 gnd.n3579 0.152939
R12733 gnd.n3580 gnd.n1616 0.152939
R12734 gnd.n3600 gnd.n1616 0.152939
R12735 gnd.n3601 gnd.n3600 0.152939
R12736 gnd.n3602 gnd.n3601 0.152939
R12737 gnd.n3602 gnd.n1604 0.152939
R12738 gnd.n3621 gnd.n1604 0.152939
R12739 gnd.n3622 gnd.n3621 0.152939
R12740 gnd.n3623 gnd.n3622 0.152939
R12741 gnd.n3623 gnd.n1592 0.152939
R12742 gnd.n3642 gnd.n1592 0.152939
R12743 gnd.n3643 gnd.n3642 0.152939
R12744 gnd.n3644 gnd.n3643 0.152939
R12745 gnd.n3644 gnd.n1579 0.152939
R12746 gnd.n3663 gnd.n1579 0.152939
R12747 gnd.n3664 gnd.n3663 0.152939
R12748 gnd.n3665 gnd.n3664 0.152939
R12749 gnd.n3666 gnd.n3665 0.152939
R12750 gnd.n3668 gnd.n3666 0.152939
R12751 gnd.n3668 gnd.n3667 0.152939
R12752 gnd.n3667 gnd.n494 0.152939
R12753 gnd.n495 gnd.n494 0.152939
R12754 gnd.n496 gnd.n495 0.152939
R12755 gnd.n509 gnd.n496 0.152939
R12756 gnd.n510 gnd.n509 0.152939
R12757 gnd.n511 gnd.n510 0.152939
R12758 gnd.n512 gnd.n511 0.152939
R12759 gnd.n513 gnd.n512 0.152939
R12760 gnd.n514 gnd.n513 0.152939
R12761 gnd.n518 gnd.n514 0.152939
R12762 gnd.n519 gnd.n518 0.152939
R12763 gnd.n6328 gnd.n519 0.152939
R12764 gnd.n843 gnd.n838 0.152939
R12765 gnd.n844 gnd.n843 0.152939
R12766 gnd.n845 gnd.n844 0.152939
R12767 gnd.n850 gnd.n845 0.152939
R12768 gnd.n851 gnd.n850 0.152939
R12769 gnd.n852 gnd.n851 0.152939
R12770 gnd.n853 gnd.n852 0.152939
R12771 gnd.n858 gnd.n853 0.152939
R12772 gnd.n859 gnd.n858 0.152939
R12773 gnd.n860 gnd.n859 0.152939
R12774 gnd.n861 gnd.n860 0.152939
R12775 gnd.n866 gnd.n861 0.152939
R12776 gnd.n867 gnd.n866 0.152939
R12777 gnd.n868 gnd.n867 0.152939
R12778 gnd.n869 gnd.n868 0.152939
R12779 gnd.n874 gnd.n869 0.152939
R12780 gnd.n875 gnd.n874 0.152939
R12781 gnd.n876 gnd.n875 0.152939
R12782 gnd.n877 gnd.n876 0.152939
R12783 gnd.n882 gnd.n877 0.152939
R12784 gnd.n883 gnd.n882 0.152939
R12785 gnd.n884 gnd.n883 0.152939
R12786 gnd.n885 gnd.n884 0.152939
R12787 gnd.n890 gnd.n885 0.152939
R12788 gnd.n891 gnd.n890 0.152939
R12789 gnd.n892 gnd.n891 0.152939
R12790 gnd.n893 gnd.n892 0.152939
R12791 gnd.n898 gnd.n893 0.152939
R12792 gnd.n899 gnd.n898 0.152939
R12793 gnd.n900 gnd.n899 0.152939
R12794 gnd.n901 gnd.n900 0.152939
R12795 gnd.n906 gnd.n901 0.152939
R12796 gnd.n907 gnd.n906 0.152939
R12797 gnd.n908 gnd.n907 0.152939
R12798 gnd.n909 gnd.n908 0.152939
R12799 gnd.n914 gnd.n909 0.152939
R12800 gnd.n915 gnd.n914 0.152939
R12801 gnd.n916 gnd.n915 0.152939
R12802 gnd.n917 gnd.n916 0.152939
R12803 gnd.n922 gnd.n917 0.152939
R12804 gnd.n923 gnd.n922 0.152939
R12805 gnd.n924 gnd.n923 0.152939
R12806 gnd.n925 gnd.n924 0.152939
R12807 gnd.n930 gnd.n925 0.152939
R12808 gnd.n931 gnd.n930 0.152939
R12809 gnd.n932 gnd.n931 0.152939
R12810 gnd.n933 gnd.n932 0.152939
R12811 gnd.n938 gnd.n933 0.152939
R12812 gnd.n939 gnd.n938 0.152939
R12813 gnd.n940 gnd.n939 0.152939
R12814 gnd.n941 gnd.n940 0.152939
R12815 gnd.n946 gnd.n941 0.152939
R12816 gnd.n947 gnd.n946 0.152939
R12817 gnd.n948 gnd.n947 0.152939
R12818 gnd.n949 gnd.n948 0.152939
R12819 gnd.n954 gnd.n949 0.152939
R12820 gnd.n955 gnd.n954 0.152939
R12821 gnd.n956 gnd.n955 0.152939
R12822 gnd.n957 gnd.n956 0.152939
R12823 gnd.n962 gnd.n957 0.152939
R12824 gnd.n963 gnd.n962 0.152939
R12825 gnd.n964 gnd.n963 0.152939
R12826 gnd.n965 gnd.n964 0.152939
R12827 gnd.n970 gnd.n965 0.152939
R12828 gnd.n971 gnd.n970 0.152939
R12829 gnd.n972 gnd.n971 0.152939
R12830 gnd.n973 gnd.n972 0.152939
R12831 gnd.n978 gnd.n973 0.152939
R12832 gnd.n979 gnd.n978 0.152939
R12833 gnd.n980 gnd.n979 0.152939
R12834 gnd.n981 gnd.n980 0.152939
R12835 gnd.n986 gnd.n981 0.152939
R12836 gnd.n987 gnd.n986 0.152939
R12837 gnd.n988 gnd.n987 0.152939
R12838 gnd.n989 gnd.n988 0.152939
R12839 gnd.n994 gnd.n989 0.152939
R12840 gnd.n995 gnd.n994 0.152939
R12841 gnd.n996 gnd.n995 0.152939
R12842 gnd.n997 gnd.n996 0.152939
R12843 gnd.n1002 gnd.n997 0.152939
R12844 gnd.n1003 gnd.n1002 0.152939
R12845 gnd.n1004 gnd.n1003 0.152939
R12846 gnd.n1005 gnd.n1004 0.152939
R12847 gnd.n2520 gnd.n1005 0.152939
R12848 gnd.n2639 gnd.n2638 0.152939
R12849 gnd.n2641 gnd.n2639 0.152939
R12850 gnd.n2641 gnd.n2640 0.152939
R12851 gnd.n2640 gnd.n2050 0.152939
R12852 gnd.n2668 gnd.n2050 0.152939
R12853 gnd.n2669 gnd.n2668 0.152939
R12854 gnd.n2671 gnd.n2669 0.152939
R12855 gnd.n2671 gnd.n2670 0.152939
R12856 gnd.n2670 gnd.n2024 0.152939
R12857 gnd.n2698 gnd.n2024 0.152939
R12858 gnd.n2699 gnd.n2698 0.152939
R12859 gnd.n2701 gnd.n2699 0.152939
R12860 gnd.n2701 gnd.n2700 0.152939
R12861 gnd.n2700 gnd.n2000 0.152939
R12862 gnd.n2728 gnd.n2000 0.152939
R12863 gnd.n2729 gnd.n2728 0.152939
R12864 gnd.n2735 gnd.n2729 0.152939
R12865 gnd.n2735 gnd.n2734 0.152939
R12866 gnd.n2734 gnd.n2733 0.152939
R12867 gnd.n2733 gnd.n2731 0.152939
R12868 gnd.n2731 gnd.n2730 0.152939
R12869 gnd.n2730 gnd.n1975 0.152939
R12870 gnd.n2898 gnd.n1975 0.152939
R12871 gnd.n2899 gnd.n2898 0.152939
R12872 gnd.n2901 gnd.n2899 0.152939
R12873 gnd.n2901 gnd.n2900 0.152939
R12874 gnd.n2900 gnd.n1948 0.152939
R12875 gnd.n2935 gnd.n1948 0.152939
R12876 gnd.n2936 gnd.n2935 0.152939
R12877 gnd.n2937 gnd.n2936 0.152939
R12878 gnd.n2937 gnd.n1929 0.152939
R12879 gnd.n2964 gnd.n1929 0.152939
R12880 gnd.n2965 gnd.n2964 0.152939
R12881 gnd.n2967 gnd.n2965 0.152939
R12882 gnd.n2967 gnd.n2966 0.152939
R12883 gnd.n2966 gnd.n1900 0.152939
R12884 gnd.n3003 gnd.n1900 0.152939
R12885 gnd.n3004 gnd.n3003 0.152939
R12886 gnd.n3020 gnd.n3004 0.152939
R12887 gnd.n3020 gnd.n3019 0.152939
R12888 gnd.n3019 gnd.n3018 0.152939
R12889 gnd.n3018 gnd.n3005 0.152939
R12890 gnd.n3014 gnd.n3005 0.152939
R12891 gnd.n3014 gnd.n3013 0.152939
R12892 gnd.n3013 gnd.n3012 0.152939
R12893 gnd.n3012 gnd.n3010 0.152939
R12894 gnd.n3010 gnd.n1852 0.152939
R12895 gnd.n3088 gnd.n1852 0.152939
R12896 gnd.n3089 gnd.n3088 0.152939
R12897 gnd.n3090 gnd.n3089 0.152939
R12898 gnd.n3090 gnd.n1830 0.152939
R12899 gnd.n3140 gnd.n1830 0.152939
R12900 gnd.n3140 gnd.n3139 0.152939
R12901 gnd.n3139 gnd.n3138 0.152939
R12902 gnd.n3138 gnd.n1807 0.152939
R12903 gnd.n3180 gnd.n1807 0.152939
R12904 gnd.n3180 gnd.n3179 0.152939
R12905 gnd.n3179 gnd.n3178 0.152939
R12906 gnd.n3178 gnd.n1784 0.152939
R12907 gnd.n3229 gnd.n1784 0.152939
R12908 gnd.n3229 gnd.n3228 0.152939
R12909 gnd.n3228 gnd.n3227 0.152939
R12910 gnd.n3227 gnd.n1785 0.152939
R12911 gnd.n3223 gnd.n1785 0.152939
R12912 gnd.n3223 gnd.n3222 0.152939
R12913 gnd.n3222 gnd.n1733 0.152939
R12914 gnd.n3296 gnd.n1733 0.152939
R12915 gnd.n3297 gnd.n3296 0.152939
R12916 gnd.n3299 gnd.n3297 0.152939
R12917 gnd.n3299 gnd.n3298 0.152939
R12918 gnd.n3298 gnd.n1707 0.152939
R12919 gnd.n3351 gnd.n1707 0.152939
R12920 gnd.n3352 gnd.n3351 0.152939
R12921 gnd.n3362 gnd.n3352 0.152939
R12922 gnd.n3362 gnd.n3361 0.152939
R12923 gnd.n3361 gnd.n3360 0.152939
R12924 gnd.n3360 gnd.n3353 0.152939
R12925 gnd.n3356 gnd.n3353 0.152939
R12926 gnd.n3356 gnd.n1633 0.152939
R12927 gnd.n3568 gnd.n1633 0.152939
R12928 gnd.n3569 gnd.n3568 0.152939
R12929 gnd.n3570 gnd.n3569 0.152939
R12930 gnd.n3570 gnd.n1621 0.152939
R12931 gnd.n3590 gnd.n1621 0.152939
R12932 gnd.n3591 gnd.n3590 0.152939
R12933 gnd.n3592 gnd.n3591 0.152939
R12934 gnd.n3592 gnd.n1610 0.152939
R12935 gnd.n3611 gnd.n1610 0.152939
R12936 gnd.n3612 gnd.n3611 0.152939
R12937 gnd.n3613 gnd.n3612 0.152939
R12938 gnd.n3613 gnd.n1598 0.152939
R12939 gnd.n3632 gnd.n1598 0.152939
R12940 gnd.n3633 gnd.n3632 0.152939
R12941 gnd.n3634 gnd.n3633 0.152939
R12942 gnd.n3634 gnd.n1586 0.152939
R12943 gnd.n3653 gnd.n1586 0.152939
R12944 gnd.n3654 gnd.n3653 0.152939
R12945 gnd.n3656 gnd.n3654 0.152939
R12946 gnd.n3656 gnd.n3655 0.152939
R12947 gnd.n3655 gnd.n453 0.152939
R12948 gnd.n6374 gnd.n453 0.152939
R12949 gnd.n2409 gnd.n2296 0.152939
R12950 gnd.n2414 gnd.n2296 0.152939
R12951 gnd.n2415 gnd.n2414 0.152939
R12952 gnd.n2416 gnd.n2415 0.152939
R12953 gnd.n2416 gnd.n2293 0.152939
R12954 gnd.n2421 gnd.n2293 0.152939
R12955 gnd.n2422 gnd.n2421 0.152939
R12956 gnd.n2423 gnd.n2422 0.152939
R12957 gnd.n2423 gnd.n2290 0.152939
R12958 gnd.n2428 gnd.n2290 0.152939
R12959 gnd.n2429 gnd.n2428 0.152939
R12960 gnd.n2430 gnd.n2429 0.152939
R12961 gnd.n2430 gnd.n2287 0.152939
R12962 gnd.n2499 gnd.n2287 0.152939
R12963 gnd.n2500 gnd.n2499 0.152939
R12964 gnd.n2502 gnd.n2500 0.152939
R12965 gnd.n2502 gnd.n2501 0.152939
R12966 gnd.n2501 gnd.n2282 0.152939
R12967 gnd.n2539 gnd.n2282 0.152939
R12968 gnd.n2540 gnd.n2539 0.152939
R12969 gnd.n2630 gnd.n2082 0.152939
R12970 gnd.n2626 gnd.n2082 0.152939
R12971 gnd.n2626 gnd.n2625 0.152939
R12972 gnd.n2625 gnd.n2624 0.152939
R12973 gnd.n2624 gnd.n2086 0.152939
R12974 gnd.n2620 gnd.n2086 0.152939
R12975 gnd.n2632 gnd.n2631 0.152939
R12976 gnd.n2631 gnd.n2059 0.152939
R12977 gnd.n2659 gnd.n2059 0.152939
R12978 gnd.n2660 gnd.n2659 0.152939
R12979 gnd.n2662 gnd.n2660 0.152939
R12980 gnd.n2662 gnd.n2661 0.152939
R12981 gnd.n2661 gnd.n2034 0.152939
R12982 gnd.n2689 gnd.n2034 0.152939
R12983 gnd.n2690 gnd.n2689 0.152939
R12984 gnd.n2692 gnd.n2690 0.152939
R12985 gnd.n2692 gnd.n2691 0.152939
R12986 gnd.n2691 gnd.n2009 0.152939
R12987 gnd.n2719 gnd.n2009 0.152939
R12988 gnd.n2720 gnd.n2719 0.152939
R12989 gnd.n2722 gnd.n2720 0.152939
R12990 gnd.n2722 gnd.n2721 0.152939
R12991 gnd.n2721 gnd.n1984 0.152939
R12992 gnd.n2766 gnd.n1984 0.152939
R12993 gnd.n2767 gnd.n2766 0.152939
R12994 gnd.n2769 gnd.n2767 0.152939
R12995 gnd.n2769 gnd.n2768 0.152939
R12996 gnd.n2768 gnd.n1479 0.152939
R12997 gnd.n3791 gnd.n1479 0.152939
R12998 gnd.n3791 gnd.n3790 0.152939
R12999 gnd.n3790 gnd.n3789 0.152939
R13000 gnd.n3789 gnd.n1480 0.152939
R13001 gnd.n3785 gnd.n1480 0.152939
R13002 gnd.n3785 gnd.n3784 0.152939
R13003 gnd.n3784 gnd.n3783 0.152939
R13004 gnd.n3783 gnd.n1485 0.152939
R13005 gnd.n3779 gnd.n1485 0.152939
R13006 gnd.n3779 gnd.n3778 0.152939
R13007 gnd.n3778 gnd.n3777 0.152939
R13008 gnd.n3777 gnd.n1490 0.152939
R13009 gnd.n3773 gnd.n1490 0.152939
R13010 gnd.n3773 gnd.n3772 0.152939
R13011 gnd.n3772 gnd.n3771 0.152939
R13012 gnd.n3771 gnd.n1495 0.152939
R13013 gnd.n3767 gnd.n1495 0.152939
R13014 gnd.n3767 gnd.n3766 0.152939
R13015 gnd.n3766 gnd.n3765 0.152939
R13016 gnd.n3765 gnd.n1500 0.152939
R13017 gnd.n3761 gnd.n1500 0.152939
R13018 gnd.n3761 gnd.n3760 0.152939
R13019 gnd.n3760 gnd.n3759 0.152939
R13020 gnd.n3759 gnd.n1505 0.152939
R13021 gnd.n3755 gnd.n1505 0.152939
R13022 gnd.n3755 gnd.n3754 0.152939
R13023 gnd.n3754 gnd.n3753 0.152939
R13024 gnd.n3753 gnd.n1510 0.152939
R13025 gnd.n3749 gnd.n1510 0.152939
R13026 gnd.n3749 gnd.n3748 0.152939
R13027 gnd.n3748 gnd.n3747 0.152939
R13028 gnd.n3747 gnd.n1515 0.152939
R13029 gnd.n3743 gnd.n1515 0.152939
R13030 gnd.n3743 gnd.n3742 0.152939
R13031 gnd.n3742 gnd.n3741 0.152939
R13032 gnd.n3741 gnd.n1520 0.152939
R13033 gnd.n3737 gnd.n1520 0.152939
R13034 gnd.n3737 gnd.n3736 0.152939
R13035 gnd.n3736 gnd.n3735 0.152939
R13036 gnd.n3735 gnd.n1525 0.152939
R13037 gnd.n3731 gnd.n1525 0.152939
R13038 gnd.n3731 gnd.n3730 0.152939
R13039 gnd.n3730 gnd.n3729 0.152939
R13040 gnd.n3729 gnd.n1530 0.152939
R13041 gnd.n3725 gnd.n1530 0.152939
R13042 gnd.n3725 gnd.n3724 0.152939
R13043 gnd.n3724 gnd.n3723 0.152939
R13044 gnd.n3723 gnd.n1535 0.152939
R13045 gnd.n3719 gnd.n1535 0.152939
R13046 gnd.n3719 gnd.n3718 0.152939
R13047 gnd.n3718 gnd.n3717 0.152939
R13048 gnd.n3717 gnd.n1540 0.152939
R13049 gnd.n3713 gnd.n1540 0.152939
R13050 gnd.n3713 gnd.n3712 0.152939
R13051 gnd.n3712 gnd.n3711 0.152939
R13052 gnd.n3711 gnd.n1545 0.152939
R13053 gnd.n3707 gnd.n1545 0.152939
R13054 gnd.n3707 gnd.n3706 0.152939
R13055 gnd.n3706 gnd.n3705 0.152939
R13056 gnd.n3705 gnd.n1550 0.152939
R13057 gnd.n3701 gnd.n1550 0.152939
R13058 gnd.n3701 gnd.n3700 0.152939
R13059 gnd.n3700 gnd.n3699 0.152939
R13060 gnd.n3699 gnd.n1555 0.152939
R13061 gnd.n3695 gnd.n1555 0.152939
R13062 gnd.n3695 gnd.n3694 0.152939
R13063 gnd.n3694 gnd.n3693 0.152939
R13064 gnd.n3693 gnd.n1560 0.152939
R13065 gnd.n3689 gnd.n1560 0.152939
R13066 gnd.n3689 gnd.n3688 0.152939
R13067 gnd.n3688 gnd.n3687 0.152939
R13068 gnd.n3687 gnd.n1565 0.152939
R13069 gnd.n3683 gnd.n1565 0.152939
R13070 gnd.n3683 gnd.n3682 0.152939
R13071 gnd.n3682 gnd.n3681 0.152939
R13072 gnd.n3681 gnd.n1570 0.152939
R13073 gnd.n3677 gnd.n1570 0.152939
R13074 gnd.n3677 gnd.n462 0.152939
R13075 gnd.n6368 gnd.n462 0.152939
R13076 gnd.n6367 gnd.n463 0.152939
R13077 gnd.n6363 gnd.n463 0.152939
R13078 gnd.n6363 gnd.n6362 0.152939
R13079 gnd.n6362 gnd.n6361 0.152939
R13080 gnd.n6361 gnd.n467 0.152939
R13081 gnd.n467 gnd.n389 0.152939
R13082 gnd.n6559 gnd.n271 0.152939
R13083 gnd.n6560 gnd.n6559 0.152939
R13084 gnd.n6562 gnd.n6560 0.152939
R13085 gnd.n6562 gnd.n6561 0.152939
R13086 gnd.n6561 gnd.n243 0.152939
R13087 gnd.n6594 gnd.n243 0.152939
R13088 gnd.n6595 gnd.n6594 0.152939
R13089 gnd.n6607 gnd.n6595 0.152939
R13090 gnd.n6607 gnd.n6606 0.152939
R13091 gnd.n6606 gnd.n6605 0.152939
R13092 gnd.n6605 gnd.n6596 0.152939
R13093 gnd.n6601 gnd.n6596 0.152939
R13094 gnd.n6601 gnd.n6600 0.152939
R13095 gnd.n6600 gnd.n198 0.152939
R13096 gnd.n6658 gnd.n198 0.152939
R13097 gnd.n6659 gnd.n6658 0.152939
R13098 gnd.n6665 gnd.n6659 0.152939
R13099 gnd.n6665 gnd.n6664 0.152939
R13100 gnd.n6664 gnd.n6663 0.152939
R13101 gnd.n6663 gnd.n67 0.152939
R13102 gnd.n7128 gnd.n7127 0.145814
R13103 gnd.n2408 gnd.n2407 0.145814
R13104 gnd.n2409 gnd.n2408 0.145814
R13105 gnd.n7128 gnd.n67 0.145814
R13106 gnd.n2620 gnd.n2619 0.128549
R13107 gnd.n6433 gnd.n389 0.128549
R13108 gnd.n4438 gnd.n0 0.127478
R13109 gnd.n5018 gnd.n5017 0.0767195
R13110 gnd.n5017 gnd.n5016 0.0767195
R13111 gnd.n2619 gnd.n2091 0.063
R13112 gnd.n6434 gnd.n6433 0.063
R13113 gnd.n6434 gnd.n388 0.0538288
R13114 gnd.n7065 gnd.n7064 0.0538288
R13115 gnd.n4054 gnd.n4053 0.0538288
R13116 gnd.n2509 gnd.n2091 0.0538288
R13117 gnd.n5584 gnd.n4200 0.0477147
R13118 gnd.n4781 gnd.n4669 0.0442063
R13119 gnd.n4782 gnd.n4781 0.0442063
R13120 gnd.n4783 gnd.n4782 0.0442063
R13121 gnd.n4783 gnd.n4658 0.0442063
R13122 gnd.n4797 gnd.n4658 0.0442063
R13123 gnd.n4798 gnd.n4797 0.0442063
R13124 gnd.n4799 gnd.n4798 0.0442063
R13125 gnd.n4799 gnd.n4645 0.0442063
R13126 gnd.n4843 gnd.n4645 0.0442063
R13127 gnd.n4844 gnd.n4843 0.0442063
R13128 gnd.n505 gnd.n388 0.0344674
R13129 gnd.n506 gnd.n505 0.0344674
R13130 gnd.n506 gnd.n265 0.0344674
R13131 gnd.n265 gnd.n262 0.0344674
R13132 gnd.n263 gnd.n262 0.0344674
R13133 gnd.n6573 gnd.n263 0.0344674
R13134 gnd.n6574 gnd.n6573 0.0344674
R13135 gnd.n6574 gnd.n237 0.0344674
R13136 gnd.n237 gnd.n235 0.0344674
R13137 gnd.n6615 gnd.n235 0.0344674
R13138 gnd.n6616 gnd.n6615 0.0344674
R13139 gnd.n6616 gnd.n219 0.0344674
R13140 gnd.n219 gnd.n216 0.0344674
R13141 gnd.n217 gnd.n216 0.0344674
R13142 gnd.n6637 gnd.n217 0.0344674
R13143 gnd.n6638 gnd.n6637 0.0344674
R13144 gnd.n6638 gnd.n191 0.0344674
R13145 gnd.n6674 gnd.n191 0.0344674
R13146 gnd.n6674 gnd.n174 0.0344674
R13147 gnd.n6691 gnd.n174 0.0344674
R13148 gnd.n6692 gnd.n6691 0.0344674
R13149 gnd.n6692 gnd.n168 0.0344674
R13150 gnd.n6700 gnd.n168 0.0344674
R13151 gnd.n6701 gnd.n6700 0.0344674
R13152 gnd.n6701 gnd.n90 0.0344674
R13153 gnd.n91 gnd.n90 0.0344674
R13154 gnd.n92 gnd.n91 0.0344674
R13155 gnd.n6708 gnd.n92 0.0344674
R13156 gnd.n6708 gnd.n109 0.0344674
R13157 gnd.n110 gnd.n109 0.0344674
R13158 gnd.n111 gnd.n110 0.0344674
R13159 gnd.n6715 gnd.n111 0.0344674
R13160 gnd.n6715 gnd.n128 0.0344674
R13161 gnd.n129 gnd.n128 0.0344674
R13162 gnd.n130 gnd.n129 0.0344674
R13163 gnd.n6722 gnd.n130 0.0344674
R13164 gnd.n6722 gnd.n147 0.0344674
R13165 gnd.n148 gnd.n147 0.0344674
R13166 gnd.n149 gnd.n148 0.0344674
R13167 gnd.n6729 gnd.n149 0.0344674
R13168 gnd.n6729 gnd.n166 0.0344674
R13169 gnd.n7065 gnd.n166 0.0344674
R13170 gnd.n4846 gnd.n4579 0.0344674
R13171 gnd.n4053 gnd.n1131 0.0344674
R13172 gnd.n2434 gnd.n1131 0.0344674
R13173 gnd.n2434 gnd.n1152 0.0344674
R13174 gnd.n1153 gnd.n1152 0.0344674
R13175 gnd.n1154 gnd.n1153 0.0344674
R13176 gnd.n2441 gnd.n1154 0.0344674
R13177 gnd.n2441 gnd.n1170 0.0344674
R13178 gnd.n1171 gnd.n1170 0.0344674
R13179 gnd.n1172 gnd.n1171 0.0344674
R13180 gnd.n2448 gnd.n1172 0.0344674
R13181 gnd.n2448 gnd.n1188 0.0344674
R13182 gnd.n1189 gnd.n1188 0.0344674
R13183 gnd.n1190 gnd.n1189 0.0344674
R13184 gnd.n2455 gnd.n1190 0.0344674
R13185 gnd.n2455 gnd.n1208 0.0344674
R13186 gnd.n1209 gnd.n1208 0.0344674
R13187 gnd.n1210 gnd.n1209 0.0344674
R13188 gnd.n2462 gnd.n1210 0.0344674
R13189 gnd.n2462 gnd.n1226 0.0344674
R13190 gnd.n1227 gnd.n1226 0.0344674
R13191 gnd.n1228 gnd.n1227 0.0344674
R13192 gnd.n2469 gnd.n1228 0.0344674
R13193 gnd.n2469 gnd.n1246 0.0344674
R13194 gnd.n1247 gnd.n1246 0.0344674
R13195 gnd.n1248 gnd.n1247 0.0344674
R13196 gnd.n2476 gnd.n1248 0.0344674
R13197 gnd.n2476 gnd.n1264 0.0344674
R13198 gnd.n1265 gnd.n1264 0.0344674
R13199 gnd.n1266 gnd.n1265 0.0344674
R13200 gnd.n2483 gnd.n1266 0.0344674
R13201 gnd.n2483 gnd.n1284 0.0344674
R13202 gnd.n1285 gnd.n1284 0.0344674
R13203 gnd.n1286 gnd.n1285 0.0344674
R13204 gnd.n2490 gnd.n1286 0.0344674
R13205 gnd.n2490 gnd.n1304 0.0344674
R13206 gnd.n1305 gnd.n1304 0.0344674
R13207 gnd.n1306 gnd.n1305 0.0344674
R13208 gnd.n2285 gnd.n1306 0.0344674
R13209 gnd.n2285 gnd.n1325 0.0344674
R13210 gnd.n1326 gnd.n1325 0.0344674
R13211 gnd.n1327 gnd.n1326 0.0344674
R13212 gnd.n2509 gnd.n1327 0.0344674
R13213 gnd.n2618 gnd.n2617 0.0343753
R13214 gnd.n6432 gnd.n390 0.0343753
R13215 gnd.n2542 gnd.n2541 0.0296328
R13216 gnd.n6377 gnd.n6376 0.0296328
R13217 gnd.n4866 gnd.n4865 0.0269946
R13218 gnd.n4868 gnd.n4867 0.0269946
R13219 gnd.n4574 gnd.n4572 0.0269946
R13220 gnd.n4878 gnd.n4876 0.0269946
R13221 gnd.n4877 gnd.n4553 0.0269946
R13222 gnd.n4897 gnd.n4896 0.0269946
R13223 gnd.n4899 gnd.n4898 0.0269946
R13224 gnd.n4548 gnd.n4547 0.0269946
R13225 gnd.n4909 gnd.n4543 0.0269946
R13226 gnd.n4908 gnd.n4545 0.0269946
R13227 gnd.n4544 gnd.n4526 0.0269946
R13228 gnd.n4929 gnd.n4527 0.0269946
R13229 gnd.n4928 gnd.n4528 0.0269946
R13230 gnd.n4962 gnd.n4503 0.0269946
R13231 gnd.n4964 gnd.n4963 0.0269946
R13232 gnd.n4965 gnd.n4450 0.0269946
R13233 gnd.n4498 gnd.n4451 0.0269946
R13234 gnd.n4500 gnd.n4452 0.0269946
R13235 gnd.n4975 gnd.n4974 0.0269946
R13236 gnd.n4977 gnd.n4976 0.0269946
R13237 gnd.n4978 gnd.n4472 0.0269946
R13238 gnd.n4980 gnd.n4473 0.0269946
R13239 gnd.n4983 gnd.n4474 0.0269946
R13240 gnd.n4986 gnd.n4985 0.0269946
R13241 gnd.n4988 gnd.n4987 0.0269946
R13242 gnd.n5053 gnd.n4373 0.0269946
R13243 gnd.n5055 gnd.n5054 0.0269946
R13244 gnd.n5064 gnd.n4366 0.0269946
R13245 gnd.n5066 gnd.n5065 0.0269946
R13246 gnd.n5067 gnd.n4364 0.0269946
R13247 gnd.n5074 gnd.n5070 0.0269946
R13248 gnd.n5073 gnd.n5072 0.0269946
R13249 gnd.n5071 gnd.n4343 0.0269946
R13250 gnd.n5096 gnd.n4344 0.0269946
R13251 gnd.n5095 gnd.n4345 0.0269946
R13252 gnd.n5138 gnd.n4318 0.0269946
R13253 gnd.n5140 gnd.n5139 0.0269946
R13254 gnd.n5149 gnd.n4311 0.0269946
R13255 gnd.n5151 gnd.n5150 0.0269946
R13256 gnd.n5152 gnd.n4309 0.0269946
R13257 gnd.n5159 gnd.n5155 0.0269946
R13258 gnd.n5158 gnd.n5157 0.0269946
R13259 gnd.n5156 gnd.n4288 0.0269946
R13260 gnd.n5181 gnd.n4289 0.0269946
R13261 gnd.n5180 gnd.n4290 0.0269946
R13262 gnd.n5227 gnd.n4264 0.0269946
R13263 gnd.n5229 gnd.n5228 0.0269946
R13264 gnd.n5238 gnd.n4257 0.0269946
R13265 gnd.n5497 gnd.n4255 0.0269946
R13266 gnd.n5502 gnd.n5500 0.0269946
R13267 gnd.n5501 gnd.n4236 0.0269946
R13268 gnd.n5526 gnd.n5525 0.0269946
R13269 gnd.n2614 gnd.n2092 0.022519
R13270 gnd.n2613 gnd.n2096 0.022519
R13271 gnd.n2610 gnd.n2609 0.022519
R13272 gnd.n2606 gnd.n2102 0.022519
R13273 gnd.n2605 gnd.n2106 0.022519
R13274 gnd.n2602 gnd.n2601 0.022519
R13275 gnd.n2598 gnd.n2110 0.022519
R13276 gnd.n2597 gnd.n2114 0.022519
R13277 gnd.n2594 gnd.n2593 0.022519
R13278 gnd.n2590 gnd.n2120 0.022519
R13279 gnd.n2589 gnd.n2124 0.022519
R13280 gnd.n2586 gnd.n2585 0.022519
R13281 gnd.n2582 gnd.n2128 0.022519
R13282 gnd.n2581 gnd.n2132 0.022519
R13283 gnd.n2578 gnd.n2577 0.022519
R13284 gnd.n2574 gnd.n2138 0.022519
R13285 gnd.n2573 gnd.n2144 0.022519
R13286 gnd.n2279 gnd.n2148 0.022519
R13287 gnd.n2542 gnd.n2150 0.022519
R13288 gnd.n6428 gnd.n396 0.022519
R13289 gnd.n6427 gnd.n397 0.022519
R13290 gnd.n6424 gnd.n6423 0.022519
R13291 gnd.n6420 gnd.n402 0.022519
R13292 gnd.n6419 gnd.n406 0.022519
R13293 gnd.n6416 gnd.n6415 0.022519
R13294 gnd.n6412 gnd.n412 0.022519
R13295 gnd.n6411 gnd.n416 0.022519
R13296 gnd.n6408 gnd.n6407 0.022519
R13297 gnd.n6404 gnd.n420 0.022519
R13298 gnd.n6403 gnd.n424 0.022519
R13299 gnd.n6400 gnd.n6399 0.022519
R13300 gnd.n6396 gnd.n430 0.022519
R13301 gnd.n6395 gnd.n434 0.022519
R13302 gnd.n6392 gnd.n6391 0.022519
R13303 gnd.n6388 gnd.n438 0.022519
R13304 gnd.n6387 gnd.n444 0.022519
R13305 gnd.n6381 gnd.n6380 0.022519
R13306 gnd.n6377 gnd.n448 0.022519
R13307 gnd.n6376 gnd.n6375 0.0218415
R13308 gnd.n2541 gnd.n2075 0.0218415
R13309 gnd.n4846 gnd.n4845 0.0202011
R13310 gnd.n4845 gnd.n4844 0.0148637
R13311 gnd.n5495 gnd.n5239 0.0144266
R13312 gnd.n5496 gnd.n5495 0.0130679
R13313 gnd.n2617 gnd.n2092 0.0123564
R13314 gnd.n2614 gnd.n2613 0.0123564
R13315 gnd.n2610 gnd.n2096 0.0123564
R13316 gnd.n2609 gnd.n2102 0.0123564
R13317 gnd.n2606 gnd.n2605 0.0123564
R13318 gnd.n2602 gnd.n2106 0.0123564
R13319 gnd.n2601 gnd.n2110 0.0123564
R13320 gnd.n2598 gnd.n2597 0.0123564
R13321 gnd.n2594 gnd.n2114 0.0123564
R13322 gnd.n2593 gnd.n2120 0.0123564
R13323 gnd.n2590 gnd.n2589 0.0123564
R13324 gnd.n2586 gnd.n2124 0.0123564
R13325 gnd.n2585 gnd.n2128 0.0123564
R13326 gnd.n2582 gnd.n2581 0.0123564
R13327 gnd.n2578 gnd.n2132 0.0123564
R13328 gnd.n2577 gnd.n2138 0.0123564
R13329 gnd.n2574 gnd.n2573 0.0123564
R13330 gnd.n2148 gnd.n2144 0.0123564
R13331 gnd.n2279 gnd.n2150 0.0123564
R13332 gnd.n396 gnd.n390 0.0123564
R13333 gnd.n6428 gnd.n6427 0.0123564
R13334 gnd.n6424 gnd.n397 0.0123564
R13335 gnd.n6423 gnd.n402 0.0123564
R13336 gnd.n6420 gnd.n6419 0.0123564
R13337 gnd.n6416 gnd.n406 0.0123564
R13338 gnd.n6415 gnd.n412 0.0123564
R13339 gnd.n6412 gnd.n6411 0.0123564
R13340 gnd.n6408 gnd.n416 0.0123564
R13341 gnd.n6407 gnd.n420 0.0123564
R13342 gnd.n6404 gnd.n6403 0.0123564
R13343 gnd.n6400 gnd.n424 0.0123564
R13344 gnd.n6399 gnd.n430 0.0123564
R13345 gnd.n6396 gnd.n6395 0.0123564
R13346 gnd.n6392 gnd.n434 0.0123564
R13347 gnd.n6391 gnd.n438 0.0123564
R13348 gnd.n6388 gnd.n6387 0.0123564
R13349 gnd.n6381 gnd.n444 0.0123564
R13350 gnd.n6380 gnd.n448 0.0123564
R13351 gnd.n4865 gnd.n4579 0.00797283
R13352 gnd.n4867 gnd.n4866 0.00797283
R13353 gnd.n4868 gnd.n4574 0.00797283
R13354 gnd.n4876 gnd.n4572 0.00797283
R13355 gnd.n4878 gnd.n4877 0.00797283
R13356 gnd.n4896 gnd.n4553 0.00797283
R13357 gnd.n4898 gnd.n4897 0.00797283
R13358 gnd.n4899 gnd.n4548 0.00797283
R13359 gnd.n4547 gnd.n4543 0.00797283
R13360 gnd.n4909 gnd.n4908 0.00797283
R13361 gnd.n4545 gnd.n4544 0.00797283
R13362 gnd.n4527 gnd.n4526 0.00797283
R13363 gnd.n4929 gnd.n4928 0.00797283
R13364 gnd.n4528 gnd.n4503 0.00797283
R13365 gnd.n4963 gnd.n4962 0.00797283
R13366 gnd.n4965 gnd.n4964 0.00797283
R13367 gnd.n4498 gnd.n4450 0.00797283
R13368 gnd.n4500 gnd.n4451 0.00797283
R13369 gnd.n4974 gnd.n4452 0.00797283
R13370 gnd.n4976 gnd.n4975 0.00797283
R13371 gnd.n4978 gnd.n4977 0.00797283
R13372 gnd.n4980 gnd.n4472 0.00797283
R13373 gnd.n4983 gnd.n4473 0.00797283
R13374 gnd.n4985 gnd.n4474 0.00797283
R13375 gnd.n4988 gnd.n4986 0.00797283
R13376 gnd.n4987 gnd.n4373 0.00797283
R13377 gnd.n5055 gnd.n5053 0.00797283
R13378 gnd.n5054 gnd.n4366 0.00797283
R13379 gnd.n5065 gnd.n5064 0.00797283
R13380 gnd.n5067 gnd.n5066 0.00797283
R13381 gnd.n5070 gnd.n4364 0.00797283
R13382 gnd.n5074 gnd.n5073 0.00797283
R13383 gnd.n5072 gnd.n5071 0.00797283
R13384 gnd.n4344 gnd.n4343 0.00797283
R13385 gnd.n5096 gnd.n5095 0.00797283
R13386 gnd.n4345 gnd.n4318 0.00797283
R13387 gnd.n5140 gnd.n5138 0.00797283
R13388 gnd.n5139 gnd.n4311 0.00797283
R13389 gnd.n5150 gnd.n5149 0.00797283
R13390 gnd.n5152 gnd.n5151 0.00797283
R13391 gnd.n5155 gnd.n4309 0.00797283
R13392 gnd.n5159 gnd.n5158 0.00797283
R13393 gnd.n5157 gnd.n5156 0.00797283
R13394 gnd.n4289 gnd.n4288 0.00797283
R13395 gnd.n5181 gnd.n5180 0.00797283
R13396 gnd.n4290 gnd.n4264 0.00797283
R13397 gnd.n5229 gnd.n5227 0.00797283
R13398 gnd.n5228 gnd.n4257 0.00797283
R13399 gnd.n5239 gnd.n5238 0.00797283
R13400 gnd.n5497 gnd.n5496 0.00797283
R13401 gnd.n5500 gnd.n4255 0.00797283
R13402 gnd.n5502 gnd.n5501 0.00797283
R13403 gnd.n5525 gnd.n4236 0.00797283
R13404 gnd.n5526 gnd.n4200 0.00797283
R13405 gnd.n2619 gnd.n2618 0.00592005
R13406 gnd.n6433 gnd.n6432 0.00592005
R13407 gnd.n6651 gnd.n183 0.00417647
R13408 gnd.n6680 gnd.n183 0.00417647
R13409 gnd.n6681 gnd.n6680 0.00417647
R13410 gnd.n6682 gnd.n6681 0.00417647
R13411 gnd.n6684 gnd.n6682 0.00417647
R13412 gnd.n6684 gnd.n6683 0.00417647
R13413 gnd.n6683 gnd.n79 0.00417647
R13414 gnd.n80 gnd.n79 0.00417647
R13415 gnd.n81 gnd.n80 0.00417647
R13416 gnd.n98 gnd.n81 0.00417647
R13417 gnd.n1217 gnd.n1216 0.00417647
R13418 gnd.n1218 gnd.n1217 0.00417647
R13419 gnd.n1219 gnd.n1218 0.00417647
R13420 gnd.n1236 gnd.n1219 0.00417647
R13421 gnd.n1237 gnd.n1236 0.00417647
R13422 gnd.n1238 gnd.n1237 0.00417647
R13423 gnd.n1239 gnd.n1238 0.00417647
R13424 gnd.n1255 gnd.n1239 0.00417647
R13425 gnd.n1256 gnd.n1255 0.00417647
R13426 gnd.n1257 gnd.n1256 0.00417647
R13427 commonsourceibias.n25 commonsourceibias.t34 230.006
R13428 commonsourceibias.n91 commonsourceibias.t95 230.006
R13429 commonsourceibias.n218 commonsourceibias.t117 230.006
R13430 commonsourceibias.n154 commonsourceibias.t97 230.006
R13431 commonsourceibias.n322 commonsourceibias.t4 230.006
R13432 commonsourceibias.n281 commonsourceibias.t70 230.006
R13433 commonsourceibias.n483 commonsourceibias.t55 230.006
R13434 commonsourceibias.n419 commonsourceibias.t80 230.006
R13435 commonsourceibias.n70 commonsourceibias.t16 207.983
R13436 commonsourceibias.n136 commonsourceibias.t56 207.983
R13437 commonsourceibias.n263 commonsourceibias.t111 207.983
R13438 commonsourceibias.n199 commonsourceibias.t89 207.983
R13439 commonsourceibias.n368 commonsourceibias.t26 207.983
R13440 commonsourceibias.n402 commonsourceibias.t114 207.983
R13441 commonsourceibias.n529 commonsourceibias.t51 207.983
R13442 commonsourceibias.n465 commonsourceibias.t74 207.983
R13443 commonsourceibias.n10 commonsourceibias.t30 168.701
R13444 commonsourceibias.n63 commonsourceibias.t2 168.701
R13445 commonsourceibias.n57 commonsourceibias.t22 168.701
R13446 commonsourceibias.n16 commonsourceibias.t42 168.701
R13447 commonsourceibias.n49 commonsourceibias.t18 168.701
R13448 commonsourceibias.n43 commonsourceibias.t32 168.701
R13449 commonsourceibias.n19 commonsourceibias.t40 168.701
R13450 commonsourceibias.n21 commonsourceibias.t24 168.701
R13451 commonsourceibias.n23 commonsourceibias.t44 168.701
R13452 commonsourceibias.n26 commonsourceibias.t6 168.701
R13453 commonsourceibias.n1 commonsourceibias.t109 168.701
R13454 commonsourceibias.n129 commonsourceibias.t69 168.701
R13455 commonsourceibias.n123 commonsourceibias.t119 168.701
R13456 commonsourceibias.n7 commonsourceibias.t85 168.701
R13457 commonsourceibias.n115 commonsourceibias.t54 168.701
R13458 commonsourceibias.n109 commonsourceibias.t100 168.701
R13459 commonsourceibias.n85 commonsourceibias.t87 168.701
R13460 commonsourceibias.n87 commonsourceibias.t115 168.701
R13461 commonsourceibias.n89 commonsourceibias.t79 168.701
R13462 commonsourceibias.n92 commonsourceibias.t66 168.701
R13463 commonsourceibias.n219 commonsourceibias.t75 168.701
R13464 commonsourceibias.n216 commonsourceibias.t59 168.701
R13465 commonsourceibias.n214 commonsourceibias.t49 168.701
R13466 commonsourceibias.n212 commonsourceibias.t84 168.701
R13467 commonsourceibias.n236 commonsourceibias.t93 168.701
R13468 commonsourceibias.n242 commonsourceibias.t52 168.701
R13469 commonsourceibias.n209 commonsourceibias.t118 168.701
R13470 commonsourceibias.n250 commonsourceibias.t104 168.701
R13471 commonsourceibias.n256 commonsourceibias.t60 168.701
R13472 commonsourceibias.n203 commonsourceibias.t50 168.701
R13473 commonsourceibias.n139 commonsourceibias.t106 168.701
R13474 commonsourceibias.n192 commonsourceibias.t101 168.701
R13475 commonsourceibias.n186 commonsourceibias.t88 168.701
R13476 commonsourceibias.n145 commonsourceibias.t105 168.701
R13477 commonsourceibias.n178 commonsourceibias.t99 168.701
R13478 commonsourceibias.n172 commonsourceibias.t86 168.701
R13479 commonsourceibias.n148 commonsourceibias.t108 168.701
R13480 commonsourceibias.n150 commonsourceibias.t98 168.701
R13481 commonsourceibias.n152 commonsourceibias.t112 168.701
R13482 commonsourceibias.n155 commonsourceibias.t107 168.701
R13483 commonsourceibias.n323 commonsourceibias.t14 168.701
R13484 commonsourceibias.n320 commonsourceibias.t12 168.701
R13485 commonsourceibias.n318 commonsourceibias.t38 168.701
R13486 commonsourceibias.n316 commonsourceibias.t8 168.701
R13487 commonsourceibias.n340 commonsourceibias.t0 168.701
R13488 commonsourceibias.n346 commonsourceibias.t28 168.701
R13489 commonsourceibias.n348 commonsourceibias.t10 168.701
R13490 commonsourceibias.n355 commonsourceibias.t36 168.701
R13491 commonsourceibias.n361 commonsourceibias.t20 168.701
R13492 commonsourceibias.n308 commonsourceibias.t46 168.701
R13493 commonsourceibias.n267 commonsourceibias.t78 168.701
R13494 commonsourceibias.n395 commonsourceibias.t53 168.701
R13495 commonsourceibias.n389 commonsourceibias.t94 168.701
R13496 commonsourceibias.n382 commonsourceibias.t64 168.701
R13497 commonsourceibias.n380 commonsourceibias.t113 168.701
R13498 commonsourceibias.n282 commonsourceibias.t58 168.701
R13499 commonsourceibias.n279 commonsourceibias.t63 168.701
R13500 commonsourceibias.n277 commonsourceibias.t92 168.701
R13501 commonsourceibias.n275 commonsourceibias.t65 168.701
R13502 commonsourceibias.n299 commonsourceibias.t76 168.701
R13503 commonsourceibias.n484 commonsourceibias.t68 168.701
R13504 commonsourceibias.n481 commonsourceibias.t72 168.701
R13505 commonsourceibias.n479 commonsourceibias.t61 168.701
R13506 commonsourceibias.n477 commonsourceibias.t110 168.701
R13507 commonsourceibias.n501 commonsourceibias.t77 168.701
R13508 commonsourceibias.n507 commonsourceibias.t67 168.701
R13509 commonsourceibias.n509 commonsourceibias.t57 168.701
R13510 commonsourceibias.n516 commonsourceibias.t48 168.701
R13511 commonsourceibias.n522 commonsourceibias.t71 168.701
R13512 commonsourceibias.n469 commonsourceibias.t62 168.701
R13513 commonsourceibias.n420 commonsourceibias.t116 168.701
R13514 commonsourceibias.n417 commonsourceibias.t102 168.701
R13515 commonsourceibias.n415 commonsourceibias.t81 168.701
R13516 commonsourceibias.n413 commonsourceibias.t96 168.701
R13517 commonsourceibias.n437 commonsourceibias.t103 168.701
R13518 commonsourceibias.n443 commonsourceibias.t82 168.701
R13519 commonsourceibias.n445 commonsourceibias.t90 168.701
R13520 commonsourceibias.n452 commonsourceibias.t73 168.701
R13521 commonsourceibias.n458 commonsourceibias.t83 168.701
R13522 commonsourceibias.n405 commonsourceibias.t91 168.701
R13523 commonsourceibias.n27 commonsourceibias.n24 161.3
R13524 commonsourceibias.n29 commonsourceibias.n28 161.3
R13525 commonsourceibias.n31 commonsourceibias.n30 161.3
R13526 commonsourceibias.n32 commonsourceibias.n22 161.3
R13527 commonsourceibias.n34 commonsourceibias.n33 161.3
R13528 commonsourceibias.n36 commonsourceibias.n35 161.3
R13529 commonsourceibias.n37 commonsourceibias.n20 161.3
R13530 commonsourceibias.n39 commonsourceibias.n38 161.3
R13531 commonsourceibias.n41 commonsourceibias.n40 161.3
R13532 commonsourceibias.n42 commonsourceibias.n18 161.3
R13533 commonsourceibias.n45 commonsourceibias.n44 161.3
R13534 commonsourceibias.n46 commonsourceibias.n17 161.3
R13535 commonsourceibias.n48 commonsourceibias.n47 161.3
R13536 commonsourceibias.n50 commonsourceibias.n15 161.3
R13537 commonsourceibias.n52 commonsourceibias.n51 161.3
R13538 commonsourceibias.n53 commonsourceibias.n14 161.3
R13539 commonsourceibias.n55 commonsourceibias.n54 161.3
R13540 commonsourceibias.n56 commonsourceibias.n13 161.3
R13541 commonsourceibias.n59 commonsourceibias.n58 161.3
R13542 commonsourceibias.n60 commonsourceibias.n12 161.3
R13543 commonsourceibias.n62 commonsourceibias.n61 161.3
R13544 commonsourceibias.n64 commonsourceibias.n11 161.3
R13545 commonsourceibias.n66 commonsourceibias.n65 161.3
R13546 commonsourceibias.n68 commonsourceibias.n67 161.3
R13547 commonsourceibias.n69 commonsourceibias.n9 161.3
R13548 commonsourceibias.n93 commonsourceibias.n90 161.3
R13549 commonsourceibias.n95 commonsourceibias.n94 161.3
R13550 commonsourceibias.n97 commonsourceibias.n96 161.3
R13551 commonsourceibias.n98 commonsourceibias.n88 161.3
R13552 commonsourceibias.n100 commonsourceibias.n99 161.3
R13553 commonsourceibias.n102 commonsourceibias.n101 161.3
R13554 commonsourceibias.n103 commonsourceibias.n86 161.3
R13555 commonsourceibias.n105 commonsourceibias.n104 161.3
R13556 commonsourceibias.n107 commonsourceibias.n106 161.3
R13557 commonsourceibias.n108 commonsourceibias.n84 161.3
R13558 commonsourceibias.n111 commonsourceibias.n110 161.3
R13559 commonsourceibias.n112 commonsourceibias.n8 161.3
R13560 commonsourceibias.n114 commonsourceibias.n113 161.3
R13561 commonsourceibias.n116 commonsourceibias.n6 161.3
R13562 commonsourceibias.n118 commonsourceibias.n117 161.3
R13563 commonsourceibias.n119 commonsourceibias.n5 161.3
R13564 commonsourceibias.n121 commonsourceibias.n120 161.3
R13565 commonsourceibias.n122 commonsourceibias.n4 161.3
R13566 commonsourceibias.n125 commonsourceibias.n124 161.3
R13567 commonsourceibias.n126 commonsourceibias.n3 161.3
R13568 commonsourceibias.n128 commonsourceibias.n127 161.3
R13569 commonsourceibias.n130 commonsourceibias.n2 161.3
R13570 commonsourceibias.n132 commonsourceibias.n131 161.3
R13571 commonsourceibias.n134 commonsourceibias.n133 161.3
R13572 commonsourceibias.n135 commonsourceibias.n0 161.3
R13573 commonsourceibias.n262 commonsourceibias.n202 161.3
R13574 commonsourceibias.n261 commonsourceibias.n260 161.3
R13575 commonsourceibias.n259 commonsourceibias.n258 161.3
R13576 commonsourceibias.n257 commonsourceibias.n204 161.3
R13577 commonsourceibias.n255 commonsourceibias.n254 161.3
R13578 commonsourceibias.n253 commonsourceibias.n205 161.3
R13579 commonsourceibias.n252 commonsourceibias.n251 161.3
R13580 commonsourceibias.n249 commonsourceibias.n206 161.3
R13581 commonsourceibias.n248 commonsourceibias.n247 161.3
R13582 commonsourceibias.n246 commonsourceibias.n207 161.3
R13583 commonsourceibias.n245 commonsourceibias.n244 161.3
R13584 commonsourceibias.n243 commonsourceibias.n208 161.3
R13585 commonsourceibias.n241 commonsourceibias.n240 161.3
R13586 commonsourceibias.n239 commonsourceibias.n210 161.3
R13587 commonsourceibias.n238 commonsourceibias.n237 161.3
R13588 commonsourceibias.n235 commonsourceibias.n211 161.3
R13589 commonsourceibias.n234 commonsourceibias.n233 161.3
R13590 commonsourceibias.n232 commonsourceibias.n231 161.3
R13591 commonsourceibias.n230 commonsourceibias.n213 161.3
R13592 commonsourceibias.n229 commonsourceibias.n228 161.3
R13593 commonsourceibias.n227 commonsourceibias.n226 161.3
R13594 commonsourceibias.n225 commonsourceibias.n215 161.3
R13595 commonsourceibias.n224 commonsourceibias.n223 161.3
R13596 commonsourceibias.n222 commonsourceibias.n221 161.3
R13597 commonsourceibias.n220 commonsourceibias.n217 161.3
R13598 commonsourceibias.n156 commonsourceibias.n153 161.3
R13599 commonsourceibias.n158 commonsourceibias.n157 161.3
R13600 commonsourceibias.n160 commonsourceibias.n159 161.3
R13601 commonsourceibias.n161 commonsourceibias.n151 161.3
R13602 commonsourceibias.n163 commonsourceibias.n162 161.3
R13603 commonsourceibias.n165 commonsourceibias.n164 161.3
R13604 commonsourceibias.n166 commonsourceibias.n149 161.3
R13605 commonsourceibias.n168 commonsourceibias.n167 161.3
R13606 commonsourceibias.n170 commonsourceibias.n169 161.3
R13607 commonsourceibias.n171 commonsourceibias.n147 161.3
R13608 commonsourceibias.n174 commonsourceibias.n173 161.3
R13609 commonsourceibias.n175 commonsourceibias.n146 161.3
R13610 commonsourceibias.n177 commonsourceibias.n176 161.3
R13611 commonsourceibias.n179 commonsourceibias.n144 161.3
R13612 commonsourceibias.n181 commonsourceibias.n180 161.3
R13613 commonsourceibias.n182 commonsourceibias.n143 161.3
R13614 commonsourceibias.n184 commonsourceibias.n183 161.3
R13615 commonsourceibias.n185 commonsourceibias.n142 161.3
R13616 commonsourceibias.n188 commonsourceibias.n187 161.3
R13617 commonsourceibias.n189 commonsourceibias.n141 161.3
R13618 commonsourceibias.n191 commonsourceibias.n190 161.3
R13619 commonsourceibias.n193 commonsourceibias.n140 161.3
R13620 commonsourceibias.n195 commonsourceibias.n194 161.3
R13621 commonsourceibias.n197 commonsourceibias.n196 161.3
R13622 commonsourceibias.n198 commonsourceibias.n138 161.3
R13623 commonsourceibias.n367 commonsourceibias.n307 161.3
R13624 commonsourceibias.n366 commonsourceibias.n365 161.3
R13625 commonsourceibias.n364 commonsourceibias.n363 161.3
R13626 commonsourceibias.n362 commonsourceibias.n309 161.3
R13627 commonsourceibias.n360 commonsourceibias.n359 161.3
R13628 commonsourceibias.n358 commonsourceibias.n310 161.3
R13629 commonsourceibias.n357 commonsourceibias.n356 161.3
R13630 commonsourceibias.n354 commonsourceibias.n311 161.3
R13631 commonsourceibias.n353 commonsourceibias.n352 161.3
R13632 commonsourceibias.n351 commonsourceibias.n312 161.3
R13633 commonsourceibias.n350 commonsourceibias.n349 161.3
R13634 commonsourceibias.n347 commonsourceibias.n313 161.3
R13635 commonsourceibias.n345 commonsourceibias.n344 161.3
R13636 commonsourceibias.n343 commonsourceibias.n314 161.3
R13637 commonsourceibias.n342 commonsourceibias.n341 161.3
R13638 commonsourceibias.n339 commonsourceibias.n315 161.3
R13639 commonsourceibias.n338 commonsourceibias.n337 161.3
R13640 commonsourceibias.n336 commonsourceibias.n335 161.3
R13641 commonsourceibias.n334 commonsourceibias.n317 161.3
R13642 commonsourceibias.n333 commonsourceibias.n332 161.3
R13643 commonsourceibias.n331 commonsourceibias.n330 161.3
R13644 commonsourceibias.n329 commonsourceibias.n319 161.3
R13645 commonsourceibias.n328 commonsourceibias.n327 161.3
R13646 commonsourceibias.n326 commonsourceibias.n325 161.3
R13647 commonsourceibias.n324 commonsourceibias.n321 161.3
R13648 commonsourceibias.n301 commonsourceibias.n300 161.3
R13649 commonsourceibias.n298 commonsourceibias.n274 161.3
R13650 commonsourceibias.n297 commonsourceibias.n296 161.3
R13651 commonsourceibias.n295 commonsourceibias.n294 161.3
R13652 commonsourceibias.n293 commonsourceibias.n276 161.3
R13653 commonsourceibias.n292 commonsourceibias.n291 161.3
R13654 commonsourceibias.n290 commonsourceibias.n289 161.3
R13655 commonsourceibias.n288 commonsourceibias.n278 161.3
R13656 commonsourceibias.n287 commonsourceibias.n286 161.3
R13657 commonsourceibias.n285 commonsourceibias.n284 161.3
R13658 commonsourceibias.n283 commonsourceibias.n280 161.3
R13659 commonsourceibias.n377 commonsourceibias.n273 161.3
R13660 commonsourceibias.n401 commonsourceibias.n266 161.3
R13661 commonsourceibias.n400 commonsourceibias.n399 161.3
R13662 commonsourceibias.n398 commonsourceibias.n397 161.3
R13663 commonsourceibias.n396 commonsourceibias.n268 161.3
R13664 commonsourceibias.n394 commonsourceibias.n393 161.3
R13665 commonsourceibias.n392 commonsourceibias.n269 161.3
R13666 commonsourceibias.n391 commonsourceibias.n390 161.3
R13667 commonsourceibias.n388 commonsourceibias.n270 161.3
R13668 commonsourceibias.n387 commonsourceibias.n386 161.3
R13669 commonsourceibias.n385 commonsourceibias.n271 161.3
R13670 commonsourceibias.n384 commonsourceibias.n383 161.3
R13671 commonsourceibias.n381 commonsourceibias.n272 161.3
R13672 commonsourceibias.n379 commonsourceibias.n378 161.3
R13673 commonsourceibias.n528 commonsourceibias.n468 161.3
R13674 commonsourceibias.n527 commonsourceibias.n526 161.3
R13675 commonsourceibias.n525 commonsourceibias.n524 161.3
R13676 commonsourceibias.n523 commonsourceibias.n470 161.3
R13677 commonsourceibias.n521 commonsourceibias.n520 161.3
R13678 commonsourceibias.n519 commonsourceibias.n471 161.3
R13679 commonsourceibias.n518 commonsourceibias.n517 161.3
R13680 commonsourceibias.n515 commonsourceibias.n472 161.3
R13681 commonsourceibias.n514 commonsourceibias.n513 161.3
R13682 commonsourceibias.n512 commonsourceibias.n473 161.3
R13683 commonsourceibias.n511 commonsourceibias.n510 161.3
R13684 commonsourceibias.n508 commonsourceibias.n474 161.3
R13685 commonsourceibias.n506 commonsourceibias.n505 161.3
R13686 commonsourceibias.n504 commonsourceibias.n475 161.3
R13687 commonsourceibias.n503 commonsourceibias.n502 161.3
R13688 commonsourceibias.n500 commonsourceibias.n476 161.3
R13689 commonsourceibias.n499 commonsourceibias.n498 161.3
R13690 commonsourceibias.n497 commonsourceibias.n496 161.3
R13691 commonsourceibias.n495 commonsourceibias.n478 161.3
R13692 commonsourceibias.n494 commonsourceibias.n493 161.3
R13693 commonsourceibias.n492 commonsourceibias.n491 161.3
R13694 commonsourceibias.n490 commonsourceibias.n480 161.3
R13695 commonsourceibias.n489 commonsourceibias.n488 161.3
R13696 commonsourceibias.n487 commonsourceibias.n486 161.3
R13697 commonsourceibias.n485 commonsourceibias.n482 161.3
R13698 commonsourceibias.n464 commonsourceibias.n404 161.3
R13699 commonsourceibias.n463 commonsourceibias.n462 161.3
R13700 commonsourceibias.n461 commonsourceibias.n460 161.3
R13701 commonsourceibias.n459 commonsourceibias.n406 161.3
R13702 commonsourceibias.n457 commonsourceibias.n456 161.3
R13703 commonsourceibias.n455 commonsourceibias.n407 161.3
R13704 commonsourceibias.n454 commonsourceibias.n453 161.3
R13705 commonsourceibias.n451 commonsourceibias.n408 161.3
R13706 commonsourceibias.n450 commonsourceibias.n449 161.3
R13707 commonsourceibias.n448 commonsourceibias.n409 161.3
R13708 commonsourceibias.n447 commonsourceibias.n446 161.3
R13709 commonsourceibias.n444 commonsourceibias.n410 161.3
R13710 commonsourceibias.n442 commonsourceibias.n441 161.3
R13711 commonsourceibias.n440 commonsourceibias.n411 161.3
R13712 commonsourceibias.n439 commonsourceibias.n438 161.3
R13713 commonsourceibias.n436 commonsourceibias.n412 161.3
R13714 commonsourceibias.n435 commonsourceibias.n434 161.3
R13715 commonsourceibias.n433 commonsourceibias.n432 161.3
R13716 commonsourceibias.n431 commonsourceibias.n414 161.3
R13717 commonsourceibias.n430 commonsourceibias.n429 161.3
R13718 commonsourceibias.n428 commonsourceibias.n427 161.3
R13719 commonsourceibias.n426 commonsourceibias.n416 161.3
R13720 commonsourceibias.n425 commonsourceibias.n424 161.3
R13721 commonsourceibias.n423 commonsourceibias.n422 161.3
R13722 commonsourceibias.n421 commonsourceibias.n418 161.3
R13723 commonsourceibias.n80 commonsourceibias.n78 81.5057
R13724 commonsourceibias.n304 commonsourceibias.n302 81.5057
R13725 commonsourceibias.n80 commonsourceibias.n79 80.9324
R13726 commonsourceibias.n82 commonsourceibias.n81 80.9324
R13727 commonsourceibias.n77 commonsourceibias.n76 80.9324
R13728 commonsourceibias.n75 commonsourceibias.n74 80.9324
R13729 commonsourceibias.n73 commonsourceibias.n72 80.9324
R13730 commonsourceibias.n371 commonsourceibias.n370 80.9324
R13731 commonsourceibias.n373 commonsourceibias.n372 80.9324
R13732 commonsourceibias.n375 commonsourceibias.n374 80.9324
R13733 commonsourceibias.n306 commonsourceibias.n305 80.9324
R13734 commonsourceibias.n304 commonsourceibias.n303 80.9324
R13735 commonsourceibias.n71 commonsourceibias.n70 80.6037
R13736 commonsourceibias.n137 commonsourceibias.n136 80.6037
R13737 commonsourceibias.n264 commonsourceibias.n263 80.6037
R13738 commonsourceibias.n200 commonsourceibias.n199 80.6037
R13739 commonsourceibias.n369 commonsourceibias.n368 80.6037
R13740 commonsourceibias.n403 commonsourceibias.n402 80.6037
R13741 commonsourceibias.n530 commonsourceibias.n529 80.6037
R13742 commonsourceibias.n466 commonsourceibias.n465 80.6037
R13743 commonsourceibias.n65 commonsourceibias.n64 56.5617
R13744 commonsourceibias.n51 commonsourceibias.n50 56.5617
R13745 commonsourceibias.n42 commonsourceibias.n41 56.5617
R13746 commonsourceibias.n28 commonsourceibias.n27 56.5617
R13747 commonsourceibias.n131 commonsourceibias.n130 56.5617
R13748 commonsourceibias.n117 commonsourceibias.n116 56.5617
R13749 commonsourceibias.n108 commonsourceibias.n107 56.5617
R13750 commonsourceibias.n94 commonsourceibias.n93 56.5617
R13751 commonsourceibias.n221 commonsourceibias.n220 56.5617
R13752 commonsourceibias.n235 commonsourceibias.n234 56.5617
R13753 commonsourceibias.n244 commonsourceibias.n243 56.5617
R13754 commonsourceibias.n258 commonsourceibias.n257 56.5617
R13755 commonsourceibias.n194 commonsourceibias.n193 56.5617
R13756 commonsourceibias.n180 commonsourceibias.n179 56.5617
R13757 commonsourceibias.n171 commonsourceibias.n170 56.5617
R13758 commonsourceibias.n157 commonsourceibias.n156 56.5617
R13759 commonsourceibias.n325 commonsourceibias.n324 56.5617
R13760 commonsourceibias.n339 commonsourceibias.n338 56.5617
R13761 commonsourceibias.n349 commonsourceibias.n347 56.5617
R13762 commonsourceibias.n363 commonsourceibias.n362 56.5617
R13763 commonsourceibias.n397 commonsourceibias.n396 56.5617
R13764 commonsourceibias.n383 commonsourceibias.n381 56.5617
R13765 commonsourceibias.n284 commonsourceibias.n283 56.5617
R13766 commonsourceibias.n298 commonsourceibias.n297 56.5617
R13767 commonsourceibias.n486 commonsourceibias.n485 56.5617
R13768 commonsourceibias.n500 commonsourceibias.n499 56.5617
R13769 commonsourceibias.n510 commonsourceibias.n508 56.5617
R13770 commonsourceibias.n524 commonsourceibias.n523 56.5617
R13771 commonsourceibias.n422 commonsourceibias.n421 56.5617
R13772 commonsourceibias.n436 commonsourceibias.n435 56.5617
R13773 commonsourceibias.n446 commonsourceibias.n444 56.5617
R13774 commonsourceibias.n460 commonsourceibias.n459 56.5617
R13775 commonsourceibias.n56 commonsourceibias.n55 56.0773
R13776 commonsourceibias.n37 commonsourceibias.n36 56.0773
R13777 commonsourceibias.n122 commonsourceibias.n121 56.0773
R13778 commonsourceibias.n103 commonsourceibias.n102 56.0773
R13779 commonsourceibias.n230 commonsourceibias.n229 56.0773
R13780 commonsourceibias.n249 commonsourceibias.n248 56.0773
R13781 commonsourceibias.n185 commonsourceibias.n184 56.0773
R13782 commonsourceibias.n166 commonsourceibias.n165 56.0773
R13783 commonsourceibias.n334 commonsourceibias.n333 56.0773
R13784 commonsourceibias.n354 commonsourceibias.n353 56.0773
R13785 commonsourceibias.n388 commonsourceibias.n387 56.0773
R13786 commonsourceibias.n293 commonsourceibias.n292 56.0773
R13787 commonsourceibias.n495 commonsourceibias.n494 56.0773
R13788 commonsourceibias.n515 commonsourceibias.n514 56.0773
R13789 commonsourceibias.n431 commonsourceibias.n430 56.0773
R13790 commonsourceibias.n451 commonsourceibias.n450 56.0773
R13791 commonsourceibias.n70 commonsourceibias.n69 46.0096
R13792 commonsourceibias.n136 commonsourceibias.n135 46.0096
R13793 commonsourceibias.n263 commonsourceibias.n262 46.0096
R13794 commonsourceibias.n199 commonsourceibias.n198 46.0096
R13795 commonsourceibias.n368 commonsourceibias.n367 46.0096
R13796 commonsourceibias.n402 commonsourceibias.n401 46.0096
R13797 commonsourceibias.n529 commonsourceibias.n528 46.0096
R13798 commonsourceibias.n465 commonsourceibias.n464 46.0096
R13799 commonsourceibias.n58 commonsourceibias.n12 41.5458
R13800 commonsourceibias.n33 commonsourceibias.n32 41.5458
R13801 commonsourceibias.n124 commonsourceibias.n3 41.5458
R13802 commonsourceibias.n99 commonsourceibias.n98 41.5458
R13803 commonsourceibias.n226 commonsourceibias.n225 41.5458
R13804 commonsourceibias.n251 commonsourceibias.n205 41.5458
R13805 commonsourceibias.n187 commonsourceibias.n141 41.5458
R13806 commonsourceibias.n162 commonsourceibias.n161 41.5458
R13807 commonsourceibias.n330 commonsourceibias.n329 41.5458
R13808 commonsourceibias.n356 commonsourceibias.n310 41.5458
R13809 commonsourceibias.n390 commonsourceibias.n269 41.5458
R13810 commonsourceibias.n289 commonsourceibias.n288 41.5458
R13811 commonsourceibias.n491 commonsourceibias.n490 41.5458
R13812 commonsourceibias.n517 commonsourceibias.n471 41.5458
R13813 commonsourceibias.n427 commonsourceibias.n426 41.5458
R13814 commonsourceibias.n453 commonsourceibias.n407 41.5458
R13815 commonsourceibias.n48 commonsourceibias.n17 40.577
R13816 commonsourceibias.n44 commonsourceibias.n17 40.577
R13817 commonsourceibias.n114 commonsourceibias.n8 40.577
R13818 commonsourceibias.n110 commonsourceibias.n8 40.577
R13819 commonsourceibias.n237 commonsourceibias.n210 40.577
R13820 commonsourceibias.n241 commonsourceibias.n210 40.577
R13821 commonsourceibias.n177 commonsourceibias.n146 40.577
R13822 commonsourceibias.n173 commonsourceibias.n146 40.577
R13823 commonsourceibias.n341 commonsourceibias.n314 40.577
R13824 commonsourceibias.n345 commonsourceibias.n314 40.577
R13825 commonsourceibias.n379 commonsourceibias.n273 40.577
R13826 commonsourceibias.n300 commonsourceibias.n273 40.577
R13827 commonsourceibias.n502 commonsourceibias.n475 40.577
R13828 commonsourceibias.n506 commonsourceibias.n475 40.577
R13829 commonsourceibias.n438 commonsourceibias.n411 40.577
R13830 commonsourceibias.n442 commonsourceibias.n411 40.577
R13831 commonsourceibias.n62 commonsourceibias.n12 39.6083
R13832 commonsourceibias.n32 commonsourceibias.n31 39.6083
R13833 commonsourceibias.n128 commonsourceibias.n3 39.6083
R13834 commonsourceibias.n98 commonsourceibias.n97 39.6083
R13835 commonsourceibias.n225 commonsourceibias.n224 39.6083
R13836 commonsourceibias.n255 commonsourceibias.n205 39.6083
R13837 commonsourceibias.n191 commonsourceibias.n141 39.6083
R13838 commonsourceibias.n161 commonsourceibias.n160 39.6083
R13839 commonsourceibias.n329 commonsourceibias.n328 39.6083
R13840 commonsourceibias.n360 commonsourceibias.n310 39.6083
R13841 commonsourceibias.n394 commonsourceibias.n269 39.6083
R13842 commonsourceibias.n288 commonsourceibias.n287 39.6083
R13843 commonsourceibias.n490 commonsourceibias.n489 39.6083
R13844 commonsourceibias.n521 commonsourceibias.n471 39.6083
R13845 commonsourceibias.n426 commonsourceibias.n425 39.6083
R13846 commonsourceibias.n457 commonsourceibias.n407 39.6083
R13847 commonsourceibias.n26 commonsourceibias.n25 33.0515
R13848 commonsourceibias.n92 commonsourceibias.n91 33.0515
R13849 commonsourceibias.n155 commonsourceibias.n154 33.0515
R13850 commonsourceibias.n219 commonsourceibias.n218 33.0515
R13851 commonsourceibias.n323 commonsourceibias.n322 33.0515
R13852 commonsourceibias.n282 commonsourceibias.n281 33.0515
R13853 commonsourceibias.n484 commonsourceibias.n483 33.0515
R13854 commonsourceibias.n420 commonsourceibias.n419 33.0515
R13855 commonsourceibias.n25 commonsourceibias.n24 28.5514
R13856 commonsourceibias.n91 commonsourceibias.n90 28.5514
R13857 commonsourceibias.n218 commonsourceibias.n217 28.5514
R13858 commonsourceibias.n154 commonsourceibias.n153 28.5514
R13859 commonsourceibias.n322 commonsourceibias.n321 28.5514
R13860 commonsourceibias.n281 commonsourceibias.n280 28.5514
R13861 commonsourceibias.n483 commonsourceibias.n482 28.5514
R13862 commonsourceibias.n419 commonsourceibias.n418 28.5514
R13863 commonsourceibias.n69 commonsourceibias.n68 26.0455
R13864 commonsourceibias.n135 commonsourceibias.n134 26.0455
R13865 commonsourceibias.n262 commonsourceibias.n261 26.0455
R13866 commonsourceibias.n198 commonsourceibias.n197 26.0455
R13867 commonsourceibias.n367 commonsourceibias.n366 26.0455
R13868 commonsourceibias.n401 commonsourceibias.n400 26.0455
R13869 commonsourceibias.n528 commonsourceibias.n527 26.0455
R13870 commonsourceibias.n464 commonsourceibias.n463 26.0455
R13871 commonsourceibias.n55 commonsourceibias.n14 25.0767
R13872 commonsourceibias.n38 commonsourceibias.n37 25.0767
R13873 commonsourceibias.n121 commonsourceibias.n5 25.0767
R13874 commonsourceibias.n104 commonsourceibias.n103 25.0767
R13875 commonsourceibias.n231 commonsourceibias.n230 25.0767
R13876 commonsourceibias.n248 commonsourceibias.n207 25.0767
R13877 commonsourceibias.n184 commonsourceibias.n143 25.0767
R13878 commonsourceibias.n167 commonsourceibias.n166 25.0767
R13879 commonsourceibias.n335 commonsourceibias.n334 25.0767
R13880 commonsourceibias.n353 commonsourceibias.n312 25.0767
R13881 commonsourceibias.n387 commonsourceibias.n271 25.0767
R13882 commonsourceibias.n294 commonsourceibias.n293 25.0767
R13883 commonsourceibias.n496 commonsourceibias.n495 25.0767
R13884 commonsourceibias.n514 commonsourceibias.n473 25.0767
R13885 commonsourceibias.n432 commonsourceibias.n431 25.0767
R13886 commonsourceibias.n450 commonsourceibias.n409 25.0767
R13887 commonsourceibias.n51 commonsourceibias.n16 24.3464
R13888 commonsourceibias.n41 commonsourceibias.n19 24.3464
R13889 commonsourceibias.n117 commonsourceibias.n7 24.3464
R13890 commonsourceibias.n107 commonsourceibias.n85 24.3464
R13891 commonsourceibias.n234 commonsourceibias.n212 24.3464
R13892 commonsourceibias.n244 commonsourceibias.n209 24.3464
R13893 commonsourceibias.n180 commonsourceibias.n145 24.3464
R13894 commonsourceibias.n170 commonsourceibias.n148 24.3464
R13895 commonsourceibias.n338 commonsourceibias.n316 24.3464
R13896 commonsourceibias.n349 commonsourceibias.n348 24.3464
R13897 commonsourceibias.n383 commonsourceibias.n382 24.3464
R13898 commonsourceibias.n297 commonsourceibias.n275 24.3464
R13899 commonsourceibias.n499 commonsourceibias.n477 24.3464
R13900 commonsourceibias.n510 commonsourceibias.n509 24.3464
R13901 commonsourceibias.n435 commonsourceibias.n413 24.3464
R13902 commonsourceibias.n446 commonsourceibias.n445 24.3464
R13903 commonsourceibias.n65 commonsourceibias.n10 23.8546
R13904 commonsourceibias.n27 commonsourceibias.n26 23.8546
R13905 commonsourceibias.n131 commonsourceibias.n1 23.8546
R13906 commonsourceibias.n93 commonsourceibias.n92 23.8546
R13907 commonsourceibias.n220 commonsourceibias.n219 23.8546
R13908 commonsourceibias.n258 commonsourceibias.n203 23.8546
R13909 commonsourceibias.n194 commonsourceibias.n139 23.8546
R13910 commonsourceibias.n156 commonsourceibias.n155 23.8546
R13911 commonsourceibias.n324 commonsourceibias.n323 23.8546
R13912 commonsourceibias.n363 commonsourceibias.n308 23.8546
R13913 commonsourceibias.n397 commonsourceibias.n267 23.8546
R13914 commonsourceibias.n283 commonsourceibias.n282 23.8546
R13915 commonsourceibias.n485 commonsourceibias.n484 23.8546
R13916 commonsourceibias.n524 commonsourceibias.n469 23.8546
R13917 commonsourceibias.n421 commonsourceibias.n420 23.8546
R13918 commonsourceibias.n460 commonsourceibias.n405 23.8546
R13919 commonsourceibias.n64 commonsourceibias.n63 16.9689
R13920 commonsourceibias.n28 commonsourceibias.n23 16.9689
R13921 commonsourceibias.n130 commonsourceibias.n129 16.9689
R13922 commonsourceibias.n94 commonsourceibias.n89 16.9689
R13923 commonsourceibias.n221 commonsourceibias.n216 16.9689
R13924 commonsourceibias.n257 commonsourceibias.n256 16.9689
R13925 commonsourceibias.n193 commonsourceibias.n192 16.9689
R13926 commonsourceibias.n157 commonsourceibias.n152 16.9689
R13927 commonsourceibias.n325 commonsourceibias.n320 16.9689
R13928 commonsourceibias.n362 commonsourceibias.n361 16.9689
R13929 commonsourceibias.n396 commonsourceibias.n395 16.9689
R13930 commonsourceibias.n284 commonsourceibias.n279 16.9689
R13931 commonsourceibias.n486 commonsourceibias.n481 16.9689
R13932 commonsourceibias.n523 commonsourceibias.n522 16.9689
R13933 commonsourceibias.n422 commonsourceibias.n417 16.9689
R13934 commonsourceibias.n459 commonsourceibias.n458 16.9689
R13935 commonsourceibias.n50 commonsourceibias.n49 16.477
R13936 commonsourceibias.n43 commonsourceibias.n42 16.477
R13937 commonsourceibias.n116 commonsourceibias.n115 16.477
R13938 commonsourceibias.n109 commonsourceibias.n108 16.477
R13939 commonsourceibias.n236 commonsourceibias.n235 16.477
R13940 commonsourceibias.n243 commonsourceibias.n242 16.477
R13941 commonsourceibias.n179 commonsourceibias.n178 16.477
R13942 commonsourceibias.n172 commonsourceibias.n171 16.477
R13943 commonsourceibias.n340 commonsourceibias.n339 16.477
R13944 commonsourceibias.n347 commonsourceibias.n346 16.477
R13945 commonsourceibias.n381 commonsourceibias.n380 16.477
R13946 commonsourceibias.n299 commonsourceibias.n298 16.477
R13947 commonsourceibias.n501 commonsourceibias.n500 16.477
R13948 commonsourceibias.n508 commonsourceibias.n507 16.477
R13949 commonsourceibias.n437 commonsourceibias.n436 16.477
R13950 commonsourceibias.n444 commonsourceibias.n443 16.477
R13951 commonsourceibias.n57 commonsourceibias.n56 15.9852
R13952 commonsourceibias.n36 commonsourceibias.n21 15.9852
R13953 commonsourceibias.n123 commonsourceibias.n122 15.9852
R13954 commonsourceibias.n102 commonsourceibias.n87 15.9852
R13955 commonsourceibias.n229 commonsourceibias.n214 15.9852
R13956 commonsourceibias.n250 commonsourceibias.n249 15.9852
R13957 commonsourceibias.n186 commonsourceibias.n185 15.9852
R13958 commonsourceibias.n165 commonsourceibias.n150 15.9852
R13959 commonsourceibias.n333 commonsourceibias.n318 15.9852
R13960 commonsourceibias.n355 commonsourceibias.n354 15.9852
R13961 commonsourceibias.n389 commonsourceibias.n388 15.9852
R13962 commonsourceibias.n292 commonsourceibias.n277 15.9852
R13963 commonsourceibias.n494 commonsourceibias.n479 15.9852
R13964 commonsourceibias.n516 commonsourceibias.n515 15.9852
R13965 commonsourceibias.n430 commonsourceibias.n415 15.9852
R13966 commonsourceibias.n452 commonsourceibias.n451 15.9852
R13967 commonsourceibias.n73 commonsourceibias.n71 13.2057
R13968 commonsourceibias.n371 commonsourceibias.n369 13.2057
R13969 commonsourceibias.n532 commonsourceibias.n265 10.4122
R13970 commonsourceibias.n112 commonsourceibias.n83 9.50363
R13971 commonsourceibias.n377 commonsourceibias.n376 9.50363
R13972 commonsourceibias.n201 commonsourceibias.n137 8.7339
R13973 commonsourceibias.n467 commonsourceibias.n403 8.7339
R13974 commonsourceibias.n58 commonsourceibias.n57 8.60764
R13975 commonsourceibias.n33 commonsourceibias.n21 8.60764
R13976 commonsourceibias.n124 commonsourceibias.n123 8.60764
R13977 commonsourceibias.n99 commonsourceibias.n87 8.60764
R13978 commonsourceibias.n226 commonsourceibias.n214 8.60764
R13979 commonsourceibias.n251 commonsourceibias.n250 8.60764
R13980 commonsourceibias.n187 commonsourceibias.n186 8.60764
R13981 commonsourceibias.n162 commonsourceibias.n150 8.60764
R13982 commonsourceibias.n330 commonsourceibias.n318 8.60764
R13983 commonsourceibias.n356 commonsourceibias.n355 8.60764
R13984 commonsourceibias.n390 commonsourceibias.n389 8.60764
R13985 commonsourceibias.n289 commonsourceibias.n277 8.60764
R13986 commonsourceibias.n491 commonsourceibias.n479 8.60764
R13987 commonsourceibias.n517 commonsourceibias.n516 8.60764
R13988 commonsourceibias.n427 commonsourceibias.n415 8.60764
R13989 commonsourceibias.n453 commonsourceibias.n452 8.60764
R13990 commonsourceibias.n532 commonsourceibias.n531 8.46921
R13991 commonsourceibias.n49 commonsourceibias.n48 8.11581
R13992 commonsourceibias.n44 commonsourceibias.n43 8.11581
R13993 commonsourceibias.n115 commonsourceibias.n114 8.11581
R13994 commonsourceibias.n110 commonsourceibias.n109 8.11581
R13995 commonsourceibias.n237 commonsourceibias.n236 8.11581
R13996 commonsourceibias.n242 commonsourceibias.n241 8.11581
R13997 commonsourceibias.n178 commonsourceibias.n177 8.11581
R13998 commonsourceibias.n173 commonsourceibias.n172 8.11581
R13999 commonsourceibias.n341 commonsourceibias.n340 8.11581
R14000 commonsourceibias.n346 commonsourceibias.n345 8.11581
R14001 commonsourceibias.n380 commonsourceibias.n379 8.11581
R14002 commonsourceibias.n300 commonsourceibias.n299 8.11581
R14003 commonsourceibias.n502 commonsourceibias.n501 8.11581
R14004 commonsourceibias.n507 commonsourceibias.n506 8.11581
R14005 commonsourceibias.n438 commonsourceibias.n437 8.11581
R14006 commonsourceibias.n443 commonsourceibias.n442 8.11581
R14007 commonsourceibias.n63 commonsourceibias.n62 7.62397
R14008 commonsourceibias.n31 commonsourceibias.n23 7.62397
R14009 commonsourceibias.n129 commonsourceibias.n128 7.62397
R14010 commonsourceibias.n97 commonsourceibias.n89 7.62397
R14011 commonsourceibias.n224 commonsourceibias.n216 7.62397
R14012 commonsourceibias.n256 commonsourceibias.n255 7.62397
R14013 commonsourceibias.n192 commonsourceibias.n191 7.62397
R14014 commonsourceibias.n160 commonsourceibias.n152 7.62397
R14015 commonsourceibias.n328 commonsourceibias.n320 7.62397
R14016 commonsourceibias.n361 commonsourceibias.n360 7.62397
R14017 commonsourceibias.n395 commonsourceibias.n394 7.62397
R14018 commonsourceibias.n287 commonsourceibias.n279 7.62397
R14019 commonsourceibias.n489 commonsourceibias.n481 7.62397
R14020 commonsourceibias.n522 commonsourceibias.n521 7.62397
R14021 commonsourceibias.n425 commonsourceibias.n417 7.62397
R14022 commonsourceibias.n458 commonsourceibias.n457 7.62397
R14023 commonsourceibias.n265 commonsourceibias.n264 5.00473
R14024 commonsourceibias.n201 commonsourceibias.n200 5.00473
R14025 commonsourceibias.n531 commonsourceibias.n530 5.00473
R14026 commonsourceibias.n467 commonsourceibias.n466 5.00473
R14027 commonsourceibias commonsourceibias.n532 3.87639
R14028 commonsourceibias.n265 commonsourceibias.n201 3.72967
R14029 commonsourceibias.n531 commonsourceibias.n467 3.72967
R14030 commonsourceibias.n78 commonsourceibias.t7 2.82907
R14031 commonsourceibias.n78 commonsourceibias.t35 2.82907
R14032 commonsourceibias.n79 commonsourceibias.t25 2.82907
R14033 commonsourceibias.n79 commonsourceibias.t45 2.82907
R14034 commonsourceibias.n81 commonsourceibias.t33 2.82907
R14035 commonsourceibias.n81 commonsourceibias.t41 2.82907
R14036 commonsourceibias.n76 commonsourceibias.t43 2.82907
R14037 commonsourceibias.n76 commonsourceibias.t19 2.82907
R14038 commonsourceibias.n74 commonsourceibias.t3 2.82907
R14039 commonsourceibias.n74 commonsourceibias.t23 2.82907
R14040 commonsourceibias.n72 commonsourceibias.t17 2.82907
R14041 commonsourceibias.n72 commonsourceibias.t31 2.82907
R14042 commonsourceibias.n370 commonsourceibias.t47 2.82907
R14043 commonsourceibias.n370 commonsourceibias.t27 2.82907
R14044 commonsourceibias.n372 commonsourceibias.t37 2.82907
R14045 commonsourceibias.n372 commonsourceibias.t21 2.82907
R14046 commonsourceibias.n374 commonsourceibias.t29 2.82907
R14047 commonsourceibias.n374 commonsourceibias.t11 2.82907
R14048 commonsourceibias.n305 commonsourceibias.t9 2.82907
R14049 commonsourceibias.n305 commonsourceibias.t1 2.82907
R14050 commonsourceibias.n303 commonsourceibias.t13 2.82907
R14051 commonsourceibias.n303 commonsourceibias.t39 2.82907
R14052 commonsourceibias.n302 commonsourceibias.t5 2.82907
R14053 commonsourceibias.n302 commonsourceibias.t15 2.82907
R14054 commonsourceibias.n68 commonsourceibias.n10 0.738255
R14055 commonsourceibias.n134 commonsourceibias.n1 0.738255
R14056 commonsourceibias.n261 commonsourceibias.n203 0.738255
R14057 commonsourceibias.n197 commonsourceibias.n139 0.738255
R14058 commonsourceibias.n366 commonsourceibias.n308 0.738255
R14059 commonsourceibias.n400 commonsourceibias.n267 0.738255
R14060 commonsourceibias.n527 commonsourceibias.n469 0.738255
R14061 commonsourceibias.n463 commonsourceibias.n405 0.738255
R14062 commonsourceibias.n75 commonsourceibias.n73 0.573776
R14063 commonsourceibias.n77 commonsourceibias.n75 0.573776
R14064 commonsourceibias.n82 commonsourceibias.n80 0.573776
R14065 commonsourceibias.n306 commonsourceibias.n304 0.573776
R14066 commonsourceibias.n375 commonsourceibias.n373 0.573776
R14067 commonsourceibias.n373 commonsourceibias.n371 0.573776
R14068 commonsourceibias.n83 commonsourceibias.n77 0.287138
R14069 commonsourceibias.n83 commonsourceibias.n82 0.287138
R14070 commonsourceibias.n376 commonsourceibias.n306 0.287138
R14071 commonsourceibias.n376 commonsourceibias.n375 0.287138
R14072 commonsourceibias.n71 commonsourceibias.n9 0.285035
R14073 commonsourceibias.n137 commonsourceibias.n0 0.285035
R14074 commonsourceibias.n264 commonsourceibias.n202 0.285035
R14075 commonsourceibias.n200 commonsourceibias.n138 0.285035
R14076 commonsourceibias.n369 commonsourceibias.n307 0.285035
R14077 commonsourceibias.n403 commonsourceibias.n266 0.285035
R14078 commonsourceibias.n530 commonsourceibias.n468 0.285035
R14079 commonsourceibias.n466 commonsourceibias.n404 0.285035
R14080 commonsourceibias.n16 commonsourceibias.n14 0.246418
R14081 commonsourceibias.n38 commonsourceibias.n19 0.246418
R14082 commonsourceibias.n7 commonsourceibias.n5 0.246418
R14083 commonsourceibias.n104 commonsourceibias.n85 0.246418
R14084 commonsourceibias.n231 commonsourceibias.n212 0.246418
R14085 commonsourceibias.n209 commonsourceibias.n207 0.246418
R14086 commonsourceibias.n145 commonsourceibias.n143 0.246418
R14087 commonsourceibias.n167 commonsourceibias.n148 0.246418
R14088 commonsourceibias.n335 commonsourceibias.n316 0.246418
R14089 commonsourceibias.n348 commonsourceibias.n312 0.246418
R14090 commonsourceibias.n382 commonsourceibias.n271 0.246418
R14091 commonsourceibias.n294 commonsourceibias.n275 0.246418
R14092 commonsourceibias.n496 commonsourceibias.n477 0.246418
R14093 commonsourceibias.n509 commonsourceibias.n473 0.246418
R14094 commonsourceibias.n432 commonsourceibias.n413 0.246418
R14095 commonsourceibias.n445 commonsourceibias.n409 0.246418
R14096 commonsourceibias.n67 commonsourceibias.n9 0.189894
R14097 commonsourceibias.n67 commonsourceibias.n66 0.189894
R14098 commonsourceibias.n66 commonsourceibias.n11 0.189894
R14099 commonsourceibias.n61 commonsourceibias.n11 0.189894
R14100 commonsourceibias.n61 commonsourceibias.n60 0.189894
R14101 commonsourceibias.n60 commonsourceibias.n59 0.189894
R14102 commonsourceibias.n59 commonsourceibias.n13 0.189894
R14103 commonsourceibias.n54 commonsourceibias.n13 0.189894
R14104 commonsourceibias.n54 commonsourceibias.n53 0.189894
R14105 commonsourceibias.n53 commonsourceibias.n52 0.189894
R14106 commonsourceibias.n52 commonsourceibias.n15 0.189894
R14107 commonsourceibias.n47 commonsourceibias.n15 0.189894
R14108 commonsourceibias.n47 commonsourceibias.n46 0.189894
R14109 commonsourceibias.n46 commonsourceibias.n45 0.189894
R14110 commonsourceibias.n45 commonsourceibias.n18 0.189894
R14111 commonsourceibias.n40 commonsourceibias.n18 0.189894
R14112 commonsourceibias.n40 commonsourceibias.n39 0.189894
R14113 commonsourceibias.n39 commonsourceibias.n20 0.189894
R14114 commonsourceibias.n35 commonsourceibias.n20 0.189894
R14115 commonsourceibias.n35 commonsourceibias.n34 0.189894
R14116 commonsourceibias.n34 commonsourceibias.n22 0.189894
R14117 commonsourceibias.n30 commonsourceibias.n22 0.189894
R14118 commonsourceibias.n30 commonsourceibias.n29 0.189894
R14119 commonsourceibias.n29 commonsourceibias.n24 0.189894
R14120 commonsourceibias.n111 commonsourceibias.n84 0.189894
R14121 commonsourceibias.n106 commonsourceibias.n84 0.189894
R14122 commonsourceibias.n106 commonsourceibias.n105 0.189894
R14123 commonsourceibias.n105 commonsourceibias.n86 0.189894
R14124 commonsourceibias.n101 commonsourceibias.n86 0.189894
R14125 commonsourceibias.n101 commonsourceibias.n100 0.189894
R14126 commonsourceibias.n100 commonsourceibias.n88 0.189894
R14127 commonsourceibias.n96 commonsourceibias.n88 0.189894
R14128 commonsourceibias.n96 commonsourceibias.n95 0.189894
R14129 commonsourceibias.n95 commonsourceibias.n90 0.189894
R14130 commonsourceibias.n133 commonsourceibias.n0 0.189894
R14131 commonsourceibias.n133 commonsourceibias.n132 0.189894
R14132 commonsourceibias.n132 commonsourceibias.n2 0.189894
R14133 commonsourceibias.n127 commonsourceibias.n2 0.189894
R14134 commonsourceibias.n127 commonsourceibias.n126 0.189894
R14135 commonsourceibias.n126 commonsourceibias.n125 0.189894
R14136 commonsourceibias.n125 commonsourceibias.n4 0.189894
R14137 commonsourceibias.n120 commonsourceibias.n4 0.189894
R14138 commonsourceibias.n120 commonsourceibias.n119 0.189894
R14139 commonsourceibias.n119 commonsourceibias.n118 0.189894
R14140 commonsourceibias.n118 commonsourceibias.n6 0.189894
R14141 commonsourceibias.n113 commonsourceibias.n6 0.189894
R14142 commonsourceibias.n260 commonsourceibias.n202 0.189894
R14143 commonsourceibias.n260 commonsourceibias.n259 0.189894
R14144 commonsourceibias.n259 commonsourceibias.n204 0.189894
R14145 commonsourceibias.n254 commonsourceibias.n204 0.189894
R14146 commonsourceibias.n254 commonsourceibias.n253 0.189894
R14147 commonsourceibias.n253 commonsourceibias.n252 0.189894
R14148 commonsourceibias.n252 commonsourceibias.n206 0.189894
R14149 commonsourceibias.n247 commonsourceibias.n206 0.189894
R14150 commonsourceibias.n247 commonsourceibias.n246 0.189894
R14151 commonsourceibias.n246 commonsourceibias.n245 0.189894
R14152 commonsourceibias.n245 commonsourceibias.n208 0.189894
R14153 commonsourceibias.n240 commonsourceibias.n208 0.189894
R14154 commonsourceibias.n240 commonsourceibias.n239 0.189894
R14155 commonsourceibias.n239 commonsourceibias.n238 0.189894
R14156 commonsourceibias.n238 commonsourceibias.n211 0.189894
R14157 commonsourceibias.n233 commonsourceibias.n211 0.189894
R14158 commonsourceibias.n233 commonsourceibias.n232 0.189894
R14159 commonsourceibias.n232 commonsourceibias.n213 0.189894
R14160 commonsourceibias.n228 commonsourceibias.n213 0.189894
R14161 commonsourceibias.n228 commonsourceibias.n227 0.189894
R14162 commonsourceibias.n227 commonsourceibias.n215 0.189894
R14163 commonsourceibias.n223 commonsourceibias.n215 0.189894
R14164 commonsourceibias.n223 commonsourceibias.n222 0.189894
R14165 commonsourceibias.n222 commonsourceibias.n217 0.189894
R14166 commonsourceibias.n196 commonsourceibias.n138 0.189894
R14167 commonsourceibias.n196 commonsourceibias.n195 0.189894
R14168 commonsourceibias.n195 commonsourceibias.n140 0.189894
R14169 commonsourceibias.n190 commonsourceibias.n140 0.189894
R14170 commonsourceibias.n190 commonsourceibias.n189 0.189894
R14171 commonsourceibias.n189 commonsourceibias.n188 0.189894
R14172 commonsourceibias.n188 commonsourceibias.n142 0.189894
R14173 commonsourceibias.n183 commonsourceibias.n142 0.189894
R14174 commonsourceibias.n183 commonsourceibias.n182 0.189894
R14175 commonsourceibias.n182 commonsourceibias.n181 0.189894
R14176 commonsourceibias.n181 commonsourceibias.n144 0.189894
R14177 commonsourceibias.n176 commonsourceibias.n144 0.189894
R14178 commonsourceibias.n176 commonsourceibias.n175 0.189894
R14179 commonsourceibias.n175 commonsourceibias.n174 0.189894
R14180 commonsourceibias.n174 commonsourceibias.n147 0.189894
R14181 commonsourceibias.n169 commonsourceibias.n147 0.189894
R14182 commonsourceibias.n169 commonsourceibias.n168 0.189894
R14183 commonsourceibias.n168 commonsourceibias.n149 0.189894
R14184 commonsourceibias.n164 commonsourceibias.n149 0.189894
R14185 commonsourceibias.n164 commonsourceibias.n163 0.189894
R14186 commonsourceibias.n163 commonsourceibias.n151 0.189894
R14187 commonsourceibias.n159 commonsourceibias.n151 0.189894
R14188 commonsourceibias.n159 commonsourceibias.n158 0.189894
R14189 commonsourceibias.n158 commonsourceibias.n153 0.189894
R14190 commonsourceibias.n326 commonsourceibias.n321 0.189894
R14191 commonsourceibias.n327 commonsourceibias.n326 0.189894
R14192 commonsourceibias.n327 commonsourceibias.n319 0.189894
R14193 commonsourceibias.n331 commonsourceibias.n319 0.189894
R14194 commonsourceibias.n332 commonsourceibias.n331 0.189894
R14195 commonsourceibias.n332 commonsourceibias.n317 0.189894
R14196 commonsourceibias.n336 commonsourceibias.n317 0.189894
R14197 commonsourceibias.n337 commonsourceibias.n336 0.189894
R14198 commonsourceibias.n337 commonsourceibias.n315 0.189894
R14199 commonsourceibias.n342 commonsourceibias.n315 0.189894
R14200 commonsourceibias.n343 commonsourceibias.n342 0.189894
R14201 commonsourceibias.n344 commonsourceibias.n343 0.189894
R14202 commonsourceibias.n344 commonsourceibias.n313 0.189894
R14203 commonsourceibias.n350 commonsourceibias.n313 0.189894
R14204 commonsourceibias.n351 commonsourceibias.n350 0.189894
R14205 commonsourceibias.n352 commonsourceibias.n351 0.189894
R14206 commonsourceibias.n352 commonsourceibias.n311 0.189894
R14207 commonsourceibias.n357 commonsourceibias.n311 0.189894
R14208 commonsourceibias.n358 commonsourceibias.n357 0.189894
R14209 commonsourceibias.n359 commonsourceibias.n358 0.189894
R14210 commonsourceibias.n359 commonsourceibias.n309 0.189894
R14211 commonsourceibias.n364 commonsourceibias.n309 0.189894
R14212 commonsourceibias.n365 commonsourceibias.n364 0.189894
R14213 commonsourceibias.n365 commonsourceibias.n307 0.189894
R14214 commonsourceibias.n285 commonsourceibias.n280 0.189894
R14215 commonsourceibias.n286 commonsourceibias.n285 0.189894
R14216 commonsourceibias.n286 commonsourceibias.n278 0.189894
R14217 commonsourceibias.n290 commonsourceibias.n278 0.189894
R14218 commonsourceibias.n291 commonsourceibias.n290 0.189894
R14219 commonsourceibias.n291 commonsourceibias.n276 0.189894
R14220 commonsourceibias.n295 commonsourceibias.n276 0.189894
R14221 commonsourceibias.n296 commonsourceibias.n295 0.189894
R14222 commonsourceibias.n296 commonsourceibias.n274 0.189894
R14223 commonsourceibias.n301 commonsourceibias.n274 0.189894
R14224 commonsourceibias.n378 commonsourceibias.n272 0.189894
R14225 commonsourceibias.n384 commonsourceibias.n272 0.189894
R14226 commonsourceibias.n385 commonsourceibias.n384 0.189894
R14227 commonsourceibias.n386 commonsourceibias.n385 0.189894
R14228 commonsourceibias.n386 commonsourceibias.n270 0.189894
R14229 commonsourceibias.n391 commonsourceibias.n270 0.189894
R14230 commonsourceibias.n392 commonsourceibias.n391 0.189894
R14231 commonsourceibias.n393 commonsourceibias.n392 0.189894
R14232 commonsourceibias.n393 commonsourceibias.n268 0.189894
R14233 commonsourceibias.n398 commonsourceibias.n268 0.189894
R14234 commonsourceibias.n399 commonsourceibias.n398 0.189894
R14235 commonsourceibias.n399 commonsourceibias.n266 0.189894
R14236 commonsourceibias.n487 commonsourceibias.n482 0.189894
R14237 commonsourceibias.n488 commonsourceibias.n487 0.189894
R14238 commonsourceibias.n488 commonsourceibias.n480 0.189894
R14239 commonsourceibias.n492 commonsourceibias.n480 0.189894
R14240 commonsourceibias.n493 commonsourceibias.n492 0.189894
R14241 commonsourceibias.n493 commonsourceibias.n478 0.189894
R14242 commonsourceibias.n497 commonsourceibias.n478 0.189894
R14243 commonsourceibias.n498 commonsourceibias.n497 0.189894
R14244 commonsourceibias.n498 commonsourceibias.n476 0.189894
R14245 commonsourceibias.n503 commonsourceibias.n476 0.189894
R14246 commonsourceibias.n504 commonsourceibias.n503 0.189894
R14247 commonsourceibias.n505 commonsourceibias.n504 0.189894
R14248 commonsourceibias.n505 commonsourceibias.n474 0.189894
R14249 commonsourceibias.n511 commonsourceibias.n474 0.189894
R14250 commonsourceibias.n512 commonsourceibias.n511 0.189894
R14251 commonsourceibias.n513 commonsourceibias.n512 0.189894
R14252 commonsourceibias.n513 commonsourceibias.n472 0.189894
R14253 commonsourceibias.n518 commonsourceibias.n472 0.189894
R14254 commonsourceibias.n519 commonsourceibias.n518 0.189894
R14255 commonsourceibias.n520 commonsourceibias.n519 0.189894
R14256 commonsourceibias.n520 commonsourceibias.n470 0.189894
R14257 commonsourceibias.n525 commonsourceibias.n470 0.189894
R14258 commonsourceibias.n526 commonsourceibias.n525 0.189894
R14259 commonsourceibias.n526 commonsourceibias.n468 0.189894
R14260 commonsourceibias.n423 commonsourceibias.n418 0.189894
R14261 commonsourceibias.n424 commonsourceibias.n423 0.189894
R14262 commonsourceibias.n424 commonsourceibias.n416 0.189894
R14263 commonsourceibias.n428 commonsourceibias.n416 0.189894
R14264 commonsourceibias.n429 commonsourceibias.n428 0.189894
R14265 commonsourceibias.n429 commonsourceibias.n414 0.189894
R14266 commonsourceibias.n433 commonsourceibias.n414 0.189894
R14267 commonsourceibias.n434 commonsourceibias.n433 0.189894
R14268 commonsourceibias.n434 commonsourceibias.n412 0.189894
R14269 commonsourceibias.n439 commonsourceibias.n412 0.189894
R14270 commonsourceibias.n440 commonsourceibias.n439 0.189894
R14271 commonsourceibias.n441 commonsourceibias.n440 0.189894
R14272 commonsourceibias.n441 commonsourceibias.n410 0.189894
R14273 commonsourceibias.n447 commonsourceibias.n410 0.189894
R14274 commonsourceibias.n448 commonsourceibias.n447 0.189894
R14275 commonsourceibias.n449 commonsourceibias.n448 0.189894
R14276 commonsourceibias.n449 commonsourceibias.n408 0.189894
R14277 commonsourceibias.n454 commonsourceibias.n408 0.189894
R14278 commonsourceibias.n455 commonsourceibias.n454 0.189894
R14279 commonsourceibias.n456 commonsourceibias.n455 0.189894
R14280 commonsourceibias.n456 commonsourceibias.n406 0.189894
R14281 commonsourceibias.n461 commonsourceibias.n406 0.189894
R14282 commonsourceibias.n462 commonsourceibias.n461 0.189894
R14283 commonsourceibias.n462 commonsourceibias.n404 0.189894
R14284 commonsourceibias.n112 commonsourceibias.n111 0.170955
R14285 commonsourceibias.n113 commonsourceibias.n112 0.170955
R14286 commonsourceibias.n377 commonsourceibias.n301 0.170955
R14287 commonsourceibias.n378 commonsourceibias.n377 0.170955
R14288 CSoutput.n19 CSoutput.t137 184.661
R14289 CSoutput.n78 CSoutput.n77 165.8
R14290 CSoutput.n76 CSoutput.n0 165.8
R14291 CSoutput.n75 CSoutput.n74 165.8
R14292 CSoutput.n73 CSoutput.n72 165.8
R14293 CSoutput.n71 CSoutput.n2 165.8
R14294 CSoutput.n69 CSoutput.n68 165.8
R14295 CSoutput.n67 CSoutput.n3 165.8
R14296 CSoutput.n66 CSoutput.n65 165.8
R14297 CSoutput.n63 CSoutput.n4 165.8
R14298 CSoutput.n61 CSoutput.n60 165.8
R14299 CSoutput.n59 CSoutput.n5 165.8
R14300 CSoutput.n58 CSoutput.n57 165.8
R14301 CSoutput.n55 CSoutput.n6 165.8
R14302 CSoutput.n54 CSoutput.n53 165.8
R14303 CSoutput.n52 CSoutput.n51 165.8
R14304 CSoutput.n50 CSoutput.n8 165.8
R14305 CSoutput.n48 CSoutput.n47 165.8
R14306 CSoutput.n46 CSoutput.n9 165.8
R14307 CSoutput.n45 CSoutput.n44 165.8
R14308 CSoutput.n42 CSoutput.n10 165.8
R14309 CSoutput.n41 CSoutput.n40 165.8
R14310 CSoutput.n39 CSoutput.n38 165.8
R14311 CSoutput.n37 CSoutput.n12 165.8
R14312 CSoutput.n35 CSoutput.n34 165.8
R14313 CSoutput.n33 CSoutput.n13 165.8
R14314 CSoutput.n32 CSoutput.n31 165.8
R14315 CSoutput.n29 CSoutput.n14 165.8
R14316 CSoutput.n28 CSoutput.n27 165.8
R14317 CSoutput.n26 CSoutput.n25 165.8
R14318 CSoutput.n24 CSoutput.n16 165.8
R14319 CSoutput.n22 CSoutput.n21 165.8
R14320 CSoutput.n20 CSoutput.n17 165.8
R14321 CSoutput.n77 CSoutput.t138 162.194
R14322 CSoutput.n18 CSoutput.t126 120.501
R14323 CSoutput.n23 CSoutput.t128 120.501
R14324 CSoutput.n15 CSoutput.t139 120.501
R14325 CSoutput.n30 CSoutput.t129 120.501
R14326 CSoutput.n36 CSoutput.t130 120.501
R14327 CSoutput.n11 CSoutput.t124 120.501
R14328 CSoutput.n43 CSoutput.t136 120.501
R14329 CSoutput.n49 CSoutput.t133 120.501
R14330 CSoutput.n7 CSoutput.t127 120.501
R14331 CSoutput.n56 CSoutput.t123 120.501
R14332 CSoutput.n62 CSoutput.t134 120.501
R14333 CSoutput.n64 CSoutput.t135 120.501
R14334 CSoutput.n70 CSoutput.t125 120.501
R14335 CSoutput.n1 CSoutput.t120 120.501
R14336 CSoutput.n270 CSoutput.n268 103.469
R14337 CSoutput.n262 CSoutput.n260 103.469
R14338 CSoutput.n255 CSoutput.n253 103.469
R14339 CSoutput.n96 CSoutput.n94 103.469
R14340 CSoutput.n88 CSoutput.n86 103.469
R14341 CSoutput.n81 CSoutput.n79 103.469
R14342 CSoutput.n272 CSoutput.n271 103.111
R14343 CSoutput.n270 CSoutput.n269 103.111
R14344 CSoutput.n266 CSoutput.n265 103.111
R14345 CSoutput.n264 CSoutput.n263 103.111
R14346 CSoutput.n262 CSoutput.n261 103.111
R14347 CSoutput.n259 CSoutput.n258 103.111
R14348 CSoutput.n257 CSoutput.n256 103.111
R14349 CSoutput.n255 CSoutput.n254 103.111
R14350 CSoutput.n96 CSoutput.n95 103.111
R14351 CSoutput.n98 CSoutput.n97 103.111
R14352 CSoutput.n100 CSoutput.n99 103.111
R14353 CSoutput.n88 CSoutput.n87 103.111
R14354 CSoutput.n90 CSoutput.n89 103.111
R14355 CSoutput.n92 CSoutput.n91 103.111
R14356 CSoutput.n81 CSoutput.n80 103.111
R14357 CSoutput.n83 CSoutput.n82 103.111
R14358 CSoutput.n85 CSoutput.n84 103.111
R14359 CSoutput.n274 CSoutput.n273 103.111
R14360 CSoutput.n302 CSoutput.n300 81.5057
R14361 CSoutput.n290 CSoutput.n288 81.5057
R14362 CSoutput.n279 CSoutput.n277 81.5057
R14363 CSoutput.n338 CSoutput.n336 81.5057
R14364 CSoutput.n326 CSoutput.n324 81.5057
R14365 CSoutput.n315 CSoutput.n313 81.5057
R14366 CSoutput.n310 CSoutput.n309 80.9324
R14367 CSoutput.n308 CSoutput.n307 80.9324
R14368 CSoutput.n306 CSoutput.n305 80.9324
R14369 CSoutput.n304 CSoutput.n303 80.9324
R14370 CSoutput.n302 CSoutput.n301 80.9324
R14371 CSoutput.n298 CSoutput.n297 80.9324
R14372 CSoutput.n296 CSoutput.n295 80.9324
R14373 CSoutput.n294 CSoutput.n293 80.9324
R14374 CSoutput.n292 CSoutput.n291 80.9324
R14375 CSoutput.n290 CSoutput.n289 80.9324
R14376 CSoutput.n287 CSoutput.n286 80.9324
R14377 CSoutput.n285 CSoutput.n284 80.9324
R14378 CSoutput.n283 CSoutput.n282 80.9324
R14379 CSoutput.n281 CSoutput.n280 80.9324
R14380 CSoutput.n279 CSoutput.n278 80.9324
R14381 CSoutput.n338 CSoutput.n337 80.9324
R14382 CSoutput.n340 CSoutput.n339 80.9324
R14383 CSoutput.n342 CSoutput.n341 80.9324
R14384 CSoutput.n344 CSoutput.n343 80.9324
R14385 CSoutput.n346 CSoutput.n345 80.9324
R14386 CSoutput.n326 CSoutput.n325 80.9324
R14387 CSoutput.n328 CSoutput.n327 80.9324
R14388 CSoutput.n330 CSoutput.n329 80.9324
R14389 CSoutput.n332 CSoutput.n331 80.9324
R14390 CSoutput.n334 CSoutput.n333 80.9324
R14391 CSoutput.n315 CSoutput.n314 80.9324
R14392 CSoutput.n317 CSoutput.n316 80.9324
R14393 CSoutput.n319 CSoutput.n318 80.9324
R14394 CSoutput.n321 CSoutput.n320 80.9324
R14395 CSoutput.n323 CSoutput.n322 80.9324
R14396 CSoutput.n25 CSoutput.n24 48.1486
R14397 CSoutput.n69 CSoutput.n3 48.1486
R14398 CSoutput.n38 CSoutput.n37 48.1486
R14399 CSoutput.n42 CSoutput.n41 48.1486
R14400 CSoutput.n51 CSoutput.n50 48.1486
R14401 CSoutput.n55 CSoutput.n54 48.1486
R14402 CSoutput.n22 CSoutput.n17 46.462
R14403 CSoutput.n72 CSoutput.n71 46.462
R14404 CSoutput.n20 CSoutput.n19 44.9055
R14405 CSoutput.n29 CSoutput.n28 43.7635
R14406 CSoutput.n65 CSoutput.n63 43.7635
R14407 CSoutput.n35 CSoutput.n13 41.7396
R14408 CSoutput.n57 CSoutput.n5 41.7396
R14409 CSoutput.n44 CSoutput.n9 37.0171
R14410 CSoutput.n48 CSoutput.n9 37.0171
R14411 CSoutput.n76 CSoutput.n75 34.9932
R14412 CSoutput.n31 CSoutput.n13 32.2947
R14413 CSoutput.n61 CSoutput.n5 32.2947
R14414 CSoutput.n30 CSoutput.n29 29.6014
R14415 CSoutput.n63 CSoutput.n62 29.6014
R14416 CSoutput.n19 CSoutput.n18 28.4085
R14417 CSoutput.n18 CSoutput.n17 25.1176
R14418 CSoutput.n72 CSoutput.n1 25.1176
R14419 CSoutput.n43 CSoutput.n42 22.0922
R14420 CSoutput.n50 CSoutput.n49 22.0922
R14421 CSoutput.n77 CSoutput.n76 21.8586
R14422 CSoutput.n37 CSoutput.n36 18.9681
R14423 CSoutput.n56 CSoutput.n55 18.9681
R14424 CSoutput.n25 CSoutput.n15 17.6292
R14425 CSoutput.n64 CSoutput.n3 17.6292
R14426 CSoutput.n24 CSoutput.n23 15.844
R14427 CSoutput.n70 CSoutput.n69 15.844
R14428 CSoutput.n38 CSoutput.n11 14.5051
R14429 CSoutput.n54 CSoutput.n7 14.5051
R14430 CSoutput.n349 CSoutput.n78 11.4982
R14431 CSoutput.n41 CSoutput.n11 11.3811
R14432 CSoutput.n51 CSoutput.n7 11.3811
R14433 CSoutput.n23 CSoutput.n22 10.0422
R14434 CSoutput.n71 CSoutput.n70 10.0422
R14435 CSoutput.n267 CSoutput.n259 9.25285
R14436 CSoutput.n93 CSoutput.n85 9.25285
R14437 CSoutput.n312 CSoutput.n276 9.07337
R14438 CSoutput.n299 CSoutput.n287 8.98182
R14439 CSoutput.n335 CSoutput.n323 8.98182
R14440 CSoutput.n28 CSoutput.n15 8.25698
R14441 CSoutput.n65 CSoutput.n64 8.25698
R14442 CSoutput.n276 CSoutput.n275 7.12641
R14443 CSoutput.n102 CSoutput.n101 7.12641
R14444 CSoutput.n36 CSoutput.n35 6.91809
R14445 CSoutput.n57 CSoutput.n56 6.91809
R14446 CSoutput.n312 CSoutput.n311 6.02792
R14447 CSoutput.n348 CSoutput.n347 6.02792
R14448 CSoutput.n349 CSoutput.n102 5.48093
R14449 CSoutput.n311 CSoutput.n310 5.25266
R14450 CSoutput.n299 CSoutput.n298 5.25266
R14451 CSoutput.n347 CSoutput.n346 5.25266
R14452 CSoutput.n335 CSoutput.n334 5.25266
R14453 CSoutput.n275 CSoutput.n274 5.1449
R14454 CSoutput.n267 CSoutput.n266 5.1449
R14455 CSoutput.n101 CSoutput.n100 5.1449
R14456 CSoutput.n93 CSoutput.n92 5.1449
R14457 CSoutput.n193 CSoutput.n146 4.5005
R14458 CSoutput.n162 CSoutput.n146 4.5005
R14459 CSoutput.n157 CSoutput.n141 4.5005
R14460 CSoutput.n157 CSoutput.n143 4.5005
R14461 CSoutput.n157 CSoutput.n140 4.5005
R14462 CSoutput.n157 CSoutput.n144 4.5005
R14463 CSoutput.n157 CSoutput.n139 4.5005
R14464 CSoutput.n157 CSoutput.t140 4.5005
R14465 CSoutput.n157 CSoutput.n138 4.5005
R14466 CSoutput.n157 CSoutput.n145 4.5005
R14467 CSoutput.n157 CSoutput.n146 4.5005
R14468 CSoutput.n155 CSoutput.n141 4.5005
R14469 CSoutput.n155 CSoutput.n143 4.5005
R14470 CSoutput.n155 CSoutput.n140 4.5005
R14471 CSoutput.n155 CSoutput.n144 4.5005
R14472 CSoutput.n155 CSoutput.n139 4.5005
R14473 CSoutput.n155 CSoutput.t140 4.5005
R14474 CSoutput.n155 CSoutput.n138 4.5005
R14475 CSoutput.n155 CSoutput.n145 4.5005
R14476 CSoutput.n155 CSoutput.n146 4.5005
R14477 CSoutput.n154 CSoutput.n141 4.5005
R14478 CSoutput.n154 CSoutput.n143 4.5005
R14479 CSoutput.n154 CSoutput.n140 4.5005
R14480 CSoutput.n154 CSoutput.n144 4.5005
R14481 CSoutput.n154 CSoutput.n139 4.5005
R14482 CSoutput.n154 CSoutput.t140 4.5005
R14483 CSoutput.n154 CSoutput.n138 4.5005
R14484 CSoutput.n154 CSoutput.n145 4.5005
R14485 CSoutput.n154 CSoutput.n146 4.5005
R14486 CSoutput.n239 CSoutput.n141 4.5005
R14487 CSoutput.n239 CSoutput.n143 4.5005
R14488 CSoutput.n239 CSoutput.n140 4.5005
R14489 CSoutput.n239 CSoutput.n144 4.5005
R14490 CSoutput.n239 CSoutput.n139 4.5005
R14491 CSoutput.n239 CSoutput.t140 4.5005
R14492 CSoutput.n239 CSoutput.n138 4.5005
R14493 CSoutput.n239 CSoutput.n145 4.5005
R14494 CSoutput.n239 CSoutput.n146 4.5005
R14495 CSoutput.n237 CSoutput.n141 4.5005
R14496 CSoutput.n237 CSoutput.n143 4.5005
R14497 CSoutput.n237 CSoutput.n140 4.5005
R14498 CSoutput.n237 CSoutput.n144 4.5005
R14499 CSoutput.n237 CSoutput.n139 4.5005
R14500 CSoutput.n237 CSoutput.t140 4.5005
R14501 CSoutput.n237 CSoutput.n138 4.5005
R14502 CSoutput.n237 CSoutput.n145 4.5005
R14503 CSoutput.n235 CSoutput.n141 4.5005
R14504 CSoutput.n235 CSoutput.n143 4.5005
R14505 CSoutput.n235 CSoutput.n140 4.5005
R14506 CSoutput.n235 CSoutput.n144 4.5005
R14507 CSoutput.n235 CSoutput.n139 4.5005
R14508 CSoutput.n235 CSoutput.t140 4.5005
R14509 CSoutput.n235 CSoutput.n138 4.5005
R14510 CSoutput.n235 CSoutput.n145 4.5005
R14511 CSoutput.n165 CSoutput.n141 4.5005
R14512 CSoutput.n165 CSoutput.n143 4.5005
R14513 CSoutput.n165 CSoutput.n140 4.5005
R14514 CSoutput.n165 CSoutput.n144 4.5005
R14515 CSoutput.n165 CSoutput.n139 4.5005
R14516 CSoutput.n165 CSoutput.t140 4.5005
R14517 CSoutput.n165 CSoutput.n138 4.5005
R14518 CSoutput.n165 CSoutput.n145 4.5005
R14519 CSoutput.n165 CSoutput.n146 4.5005
R14520 CSoutput.n164 CSoutput.n141 4.5005
R14521 CSoutput.n164 CSoutput.n143 4.5005
R14522 CSoutput.n164 CSoutput.n140 4.5005
R14523 CSoutput.n164 CSoutput.n144 4.5005
R14524 CSoutput.n164 CSoutput.n139 4.5005
R14525 CSoutput.n164 CSoutput.t140 4.5005
R14526 CSoutput.n164 CSoutput.n138 4.5005
R14527 CSoutput.n164 CSoutput.n145 4.5005
R14528 CSoutput.n164 CSoutput.n146 4.5005
R14529 CSoutput.n168 CSoutput.n141 4.5005
R14530 CSoutput.n168 CSoutput.n143 4.5005
R14531 CSoutput.n168 CSoutput.n140 4.5005
R14532 CSoutput.n168 CSoutput.n144 4.5005
R14533 CSoutput.n168 CSoutput.n139 4.5005
R14534 CSoutput.n168 CSoutput.t140 4.5005
R14535 CSoutput.n168 CSoutput.n138 4.5005
R14536 CSoutput.n168 CSoutput.n145 4.5005
R14537 CSoutput.n168 CSoutput.n146 4.5005
R14538 CSoutput.n167 CSoutput.n141 4.5005
R14539 CSoutput.n167 CSoutput.n143 4.5005
R14540 CSoutput.n167 CSoutput.n140 4.5005
R14541 CSoutput.n167 CSoutput.n144 4.5005
R14542 CSoutput.n167 CSoutput.n139 4.5005
R14543 CSoutput.n167 CSoutput.t140 4.5005
R14544 CSoutput.n167 CSoutput.n138 4.5005
R14545 CSoutput.n167 CSoutput.n145 4.5005
R14546 CSoutput.n167 CSoutput.n146 4.5005
R14547 CSoutput.n150 CSoutput.n141 4.5005
R14548 CSoutput.n150 CSoutput.n143 4.5005
R14549 CSoutput.n150 CSoutput.n140 4.5005
R14550 CSoutput.n150 CSoutput.n144 4.5005
R14551 CSoutput.n150 CSoutput.n139 4.5005
R14552 CSoutput.n150 CSoutput.t140 4.5005
R14553 CSoutput.n150 CSoutput.n138 4.5005
R14554 CSoutput.n150 CSoutput.n145 4.5005
R14555 CSoutput.n150 CSoutput.n146 4.5005
R14556 CSoutput.n242 CSoutput.n141 4.5005
R14557 CSoutput.n242 CSoutput.n143 4.5005
R14558 CSoutput.n242 CSoutput.n140 4.5005
R14559 CSoutput.n242 CSoutput.n144 4.5005
R14560 CSoutput.n242 CSoutput.n139 4.5005
R14561 CSoutput.n242 CSoutput.t140 4.5005
R14562 CSoutput.n242 CSoutput.n138 4.5005
R14563 CSoutput.n242 CSoutput.n145 4.5005
R14564 CSoutput.n242 CSoutput.n146 4.5005
R14565 CSoutput.n229 CSoutput.n200 4.5005
R14566 CSoutput.n229 CSoutput.n206 4.5005
R14567 CSoutput.n187 CSoutput.n176 4.5005
R14568 CSoutput.n187 CSoutput.n178 4.5005
R14569 CSoutput.n187 CSoutput.n175 4.5005
R14570 CSoutput.n187 CSoutput.n179 4.5005
R14571 CSoutput.n187 CSoutput.n174 4.5005
R14572 CSoutput.n187 CSoutput.t132 4.5005
R14573 CSoutput.n187 CSoutput.n173 4.5005
R14574 CSoutput.n187 CSoutput.n180 4.5005
R14575 CSoutput.n229 CSoutput.n187 4.5005
R14576 CSoutput.n208 CSoutput.n176 4.5005
R14577 CSoutput.n208 CSoutput.n178 4.5005
R14578 CSoutput.n208 CSoutput.n175 4.5005
R14579 CSoutput.n208 CSoutput.n179 4.5005
R14580 CSoutput.n208 CSoutput.n174 4.5005
R14581 CSoutput.n208 CSoutput.t132 4.5005
R14582 CSoutput.n208 CSoutput.n173 4.5005
R14583 CSoutput.n208 CSoutput.n180 4.5005
R14584 CSoutput.n229 CSoutput.n208 4.5005
R14585 CSoutput.n186 CSoutput.n176 4.5005
R14586 CSoutput.n186 CSoutput.n178 4.5005
R14587 CSoutput.n186 CSoutput.n175 4.5005
R14588 CSoutput.n186 CSoutput.n179 4.5005
R14589 CSoutput.n186 CSoutput.n174 4.5005
R14590 CSoutput.n186 CSoutput.t132 4.5005
R14591 CSoutput.n186 CSoutput.n173 4.5005
R14592 CSoutput.n186 CSoutput.n180 4.5005
R14593 CSoutput.n229 CSoutput.n186 4.5005
R14594 CSoutput.n210 CSoutput.n176 4.5005
R14595 CSoutput.n210 CSoutput.n178 4.5005
R14596 CSoutput.n210 CSoutput.n175 4.5005
R14597 CSoutput.n210 CSoutput.n179 4.5005
R14598 CSoutput.n210 CSoutput.n174 4.5005
R14599 CSoutput.n210 CSoutput.t132 4.5005
R14600 CSoutput.n210 CSoutput.n173 4.5005
R14601 CSoutput.n210 CSoutput.n180 4.5005
R14602 CSoutput.n229 CSoutput.n210 4.5005
R14603 CSoutput.n176 CSoutput.n171 4.5005
R14604 CSoutput.n178 CSoutput.n171 4.5005
R14605 CSoutput.n175 CSoutput.n171 4.5005
R14606 CSoutput.n179 CSoutput.n171 4.5005
R14607 CSoutput.n174 CSoutput.n171 4.5005
R14608 CSoutput.t132 CSoutput.n171 4.5005
R14609 CSoutput.n173 CSoutput.n171 4.5005
R14610 CSoutput.n180 CSoutput.n171 4.5005
R14611 CSoutput.n232 CSoutput.n176 4.5005
R14612 CSoutput.n232 CSoutput.n178 4.5005
R14613 CSoutput.n232 CSoutput.n175 4.5005
R14614 CSoutput.n232 CSoutput.n179 4.5005
R14615 CSoutput.n232 CSoutput.n174 4.5005
R14616 CSoutput.n232 CSoutput.t132 4.5005
R14617 CSoutput.n232 CSoutput.n173 4.5005
R14618 CSoutput.n232 CSoutput.n180 4.5005
R14619 CSoutput.n230 CSoutput.n176 4.5005
R14620 CSoutput.n230 CSoutput.n178 4.5005
R14621 CSoutput.n230 CSoutput.n175 4.5005
R14622 CSoutput.n230 CSoutput.n179 4.5005
R14623 CSoutput.n230 CSoutput.n174 4.5005
R14624 CSoutput.n230 CSoutput.t132 4.5005
R14625 CSoutput.n230 CSoutput.n173 4.5005
R14626 CSoutput.n230 CSoutput.n180 4.5005
R14627 CSoutput.n230 CSoutput.n229 4.5005
R14628 CSoutput.n212 CSoutput.n176 4.5005
R14629 CSoutput.n212 CSoutput.n178 4.5005
R14630 CSoutput.n212 CSoutput.n175 4.5005
R14631 CSoutput.n212 CSoutput.n179 4.5005
R14632 CSoutput.n212 CSoutput.n174 4.5005
R14633 CSoutput.n212 CSoutput.t132 4.5005
R14634 CSoutput.n212 CSoutput.n173 4.5005
R14635 CSoutput.n212 CSoutput.n180 4.5005
R14636 CSoutput.n229 CSoutput.n212 4.5005
R14637 CSoutput.n184 CSoutput.n176 4.5005
R14638 CSoutput.n184 CSoutput.n178 4.5005
R14639 CSoutput.n184 CSoutput.n175 4.5005
R14640 CSoutput.n184 CSoutput.n179 4.5005
R14641 CSoutput.n184 CSoutput.n174 4.5005
R14642 CSoutput.n184 CSoutput.t132 4.5005
R14643 CSoutput.n184 CSoutput.n173 4.5005
R14644 CSoutput.n184 CSoutput.n180 4.5005
R14645 CSoutput.n229 CSoutput.n184 4.5005
R14646 CSoutput.n214 CSoutput.n176 4.5005
R14647 CSoutput.n214 CSoutput.n178 4.5005
R14648 CSoutput.n214 CSoutput.n175 4.5005
R14649 CSoutput.n214 CSoutput.n179 4.5005
R14650 CSoutput.n214 CSoutput.n174 4.5005
R14651 CSoutput.n214 CSoutput.t132 4.5005
R14652 CSoutput.n214 CSoutput.n173 4.5005
R14653 CSoutput.n214 CSoutput.n180 4.5005
R14654 CSoutput.n229 CSoutput.n214 4.5005
R14655 CSoutput.n183 CSoutput.n176 4.5005
R14656 CSoutput.n183 CSoutput.n178 4.5005
R14657 CSoutput.n183 CSoutput.n175 4.5005
R14658 CSoutput.n183 CSoutput.n179 4.5005
R14659 CSoutput.n183 CSoutput.n174 4.5005
R14660 CSoutput.n183 CSoutput.t132 4.5005
R14661 CSoutput.n183 CSoutput.n173 4.5005
R14662 CSoutput.n183 CSoutput.n180 4.5005
R14663 CSoutput.n229 CSoutput.n183 4.5005
R14664 CSoutput.n228 CSoutput.n176 4.5005
R14665 CSoutput.n228 CSoutput.n178 4.5005
R14666 CSoutput.n228 CSoutput.n175 4.5005
R14667 CSoutput.n228 CSoutput.n179 4.5005
R14668 CSoutput.n228 CSoutput.n174 4.5005
R14669 CSoutput.n228 CSoutput.t132 4.5005
R14670 CSoutput.n228 CSoutput.n173 4.5005
R14671 CSoutput.n228 CSoutput.n180 4.5005
R14672 CSoutput.n229 CSoutput.n228 4.5005
R14673 CSoutput.n227 CSoutput.n112 4.5005
R14674 CSoutput.n128 CSoutput.n112 4.5005
R14675 CSoutput.n123 CSoutput.n107 4.5005
R14676 CSoutput.n123 CSoutput.n109 4.5005
R14677 CSoutput.n123 CSoutput.n106 4.5005
R14678 CSoutput.n123 CSoutput.n110 4.5005
R14679 CSoutput.n123 CSoutput.n105 4.5005
R14680 CSoutput.n123 CSoutput.t131 4.5005
R14681 CSoutput.n123 CSoutput.n104 4.5005
R14682 CSoutput.n123 CSoutput.n111 4.5005
R14683 CSoutput.n123 CSoutput.n112 4.5005
R14684 CSoutput.n121 CSoutput.n107 4.5005
R14685 CSoutput.n121 CSoutput.n109 4.5005
R14686 CSoutput.n121 CSoutput.n106 4.5005
R14687 CSoutput.n121 CSoutput.n110 4.5005
R14688 CSoutput.n121 CSoutput.n105 4.5005
R14689 CSoutput.n121 CSoutput.t131 4.5005
R14690 CSoutput.n121 CSoutput.n104 4.5005
R14691 CSoutput.n121 CSoutput.n111 4.5005
R14692 CSoutput.n121 CSoutput.n112 4.5005
R14693 CSoutput.n120 CSoutput.n107 4.5005
R14694 CSoutput.n120 CSoutput.n109 4.5005
R14695 CSoutput.n120 CSoutput.n106 4.5005
R14696 CSoutput.n120 CSoutput.n110 4.5005
R14697 CSoutput.n120 CSoutput.n105 4.5005
R14698 CSoutput.n120 CSoutput.t131 4.5005
R14699 CSoutput.n120 CSoutput.n104 4.5005
R14700 CSoutput.n120 CSoutput.n111 4.5005
R14701 CSoutput.n120 CSoutput.n112 4.5005
R14702 CSoutput.n249 CSoutput.n107 4.5005
R14703 CSoutput.n249 CSoutput.n109 4.5005
R14704 CSoutput.n249 CSoutput.n106 4.5005
R14705 CSoutput.n249 CSoutput.n110 4.5005
R14706 CSoutput.n249 CSoutput.n105 4.5005
R14707 CSoutput.n249 CSoutput.t131 4.5005
R14708 CSoutput.n249 CSoutput.n104 4.5005
R14709 CSoutput.n249 CSoutput.n111 4.5005
R14710 CSoutput.n249 CSoutput.n112 4.5005
R14711 CSoutput.n247 CSoutput.n107 4.5005
R14712 CSoutput.n247 CSoutput.n109 4.5005
R14713 CSoutput.n247 CSoutput.n106 4.5005
R14714 CSoutput.n247 CSoutput.n110 4.5005
R14715 CSoutput.n247 CSoutput.n105 4.5005
R14716 CSoutput.n247 CSoutput.t131 4.5005
R14717 CSoutput.n247 CSoutput.n104 4.5005
R14718 CSoutput.n247 CSoutput.n111 4.5005
R14719 CSoutput.n245 CSoutput.n107 4.5005
R14720 CSoutput.n245 CSoutput.n109 4.5005
R14721 CSoutput.n245 CSoutput.n106 4.5005
R14722 CSoutput.n245 CSoutput.n110 4.5005
R14723 CSoutput.n245 CSoutput.n105 4.5005
R14724 CSoutput.n245 CSoutput.t131 4.5005
R14725 CSoutput.n245 CSoutput.n104 4.5005
R14726 CSoutput.n245 CSoutput.n111 4.5005
R14727 CSoutput.n131 CSoutput.n107 4.5005
R14728 CSoutput.n131 CSoutput.n109 4.5005
R14729 CSoutput.n131 CSoutput.n106 4.5005
R14730 CSoutput.n131 CSoutput.n110 4.5005
R14731 CSoutput.n131 CSoutput.n105 4.5005
R14732 CSoutput.n131 CSoutput.t131 4.5005
R14733 CSoutput.n131 CSoutput.n104 4.5005
R14734 CSoutput.n131 CSoutput.n111 4.5005
R14735 CSoutput.n131 CSoutput.n112 4.5005
R14736 CSoutput.n130 CSoutput.n107 4.5005
R14737 CSoutput.n130 CSoutput.n109 4.5005
R14738 CSoutput.n130 CSoutput.n106 4.5005
R14739 CSoutput.n130 CSoutput.n110 4.5005
R14740 CSoutput.n130 CSoutput.n105 4.5005
R14741 CSoutput.n130 CSoutput.t131 4.5005
R14742 CSoutput.n130 CSoutput.n104 4.5005
R14743 CSoutput.n130 CSoutput.n111 4.5005
R14744 CSoutput.n130 CSoutput.n112 4.5005
R14745 CSoutput.n134 CSoutput.n107 4.5005
R14746 CSoutput.n134 CSoutput.n109 4.5005
R14747 CSoutput.n134 CSoutput.n106 4.5005
R14748 CSoutput.n134 CSoutput.n110 4.5005
R14749 CSoutput.n134 CSoutput.n105 4.5005
R14750 CSoutput.n134 CSoutput.t131 4.5005
R14751 CSoutput.n134 CSoutput.n104 4.5005
R14752 CSoutput.n134 CSoutput.n111 4.5005
R14753 CSoutput.n134 CSoutput.n112 4.5005
R14754 CSoutput.n133 CSoutput.n107 4.5005
R14755 CSoutput.n133 CSoutput.n109 4.5005
R14756 CSoutput.n133 CSoutput.n106 4.5005
R14757 CSoutput.n133 CSoutput.n110 4.5005
R14758 CSoutput.n133 CSoutput.n105 4.5005
R14759 CSoutput.n133 CSoutput.t131 4.5005
R14760 CSoutput.n133 CSoutput.n104 4.5005
R14761 CSoutput.n133 CSoutput.n111 4.5005
R14762 CSoutput.n133 CSoutput.n112 4.5005
R14763 CSoutput.n116 CSoutput.n107 4.5005
R14764 CSoutput.n116 CSoutput.n109 4.5005
R14765 CSoutput.n116 CSoutput.n106 4.5005
R14766 CSoutput.n116 CSoutput.n110 4.5005
R14767 CSoutput.n116 CSoutput.n105 4.5005
R14768 CSoutput.n116 CSoutput.t131 4.5005
R14769 CSoutput.n116 CSoutput.n104 4.5005
R14770 CSoutput.n116 CSoutput.n111 4.5005
R14771 CSoutput.n116 CSoutput.n112 4.5005
R14772 CSoutput.n252 CSoutput.n107 4.5005
R14773 CSoutput.n252 CSoutput.n109 4.5005
R14774 CSoutput.n252 CSoutput.n106 4.5005
R14775 CSoutput.n252 CSoutput.n110 4.5005
R14776 CSoutput.n252 CSoutput.n105 4.5005
R14777 CSoutput.n252 CSoutput.t131 4.5005
R14778 CSoutput.n252 CSoutput.n104 4.5005
R14779 CSoutput.n252 CSoutput.n111 4.5005
R14780 CSoutput.n252 CSoutput.n112 4.5005
R14781 CSoutput.n275 CSoutput.n267 4.10845
R14782 CSoutput.n101 CSoutput.n93 4.10845
R14783 CSoutput.n273 CSoutput.t112 4.06363
R14784 CSoutput.n273 CSoutput.t85 4.06363
R14785 CSoutput.n271 CSoutput.t104 4.06363
R14786 CSoutput.n271 CSoutput.t91 4.06363
R14787 CSoutput.n269 CSoutput.t108 4.06363
R14788 CSoutput.n269 CSoutput.t73 4.06363
R14789 CSoutput.n268 CSoutput.t95 4.06363
R14790 CSoutput.n268 CSoutput.t96 4.06363
R14791 CSoutput.n265 CSoutput.t119 4.06363
R14792 CSoutput.n265 CSoutput.t113 4.06363
R14793 CSoutput.n263 CSoutput.t79 4.06363
R14794 CSoutput.n263 CSoutput.t109 4.06363
R14795 CSoutput.n261 CSoutput.t110 4.06363
R14796 CSoutput.n261 CSoutput.t75 4.06363
R14797 CSoutput.n260 CSoutput.t106 4.06363
R14798 CSoutput.n260 CSoutput.t102 4.06363
R14799 CSoutput.n258 CSoutput.t84 4.06363
R14800 CSoutput.n258 CSoutput.t117 4.06363
R14801 CSoutput.n256 CSoutput.t115 4.06363
R14802 CSoutput.n256 CSoutput.t97 4.06363
R14803 CSoutput.n254 CSoutput.t105 4.06363
R14804 CSoutput.n254 CSoutput.t118 4.06363
R14805 CSoutput.n253 CSoutput.t81 4.06363
R14806 CSoutput.n253 CSoutput.t93 4.06363
R14807 CSoutput.n94 CSoutput.t77 4.06363
R14808 CSoutput.n94 CSoutput.t78 4.06363
R14809 CSoutput.n95 CSoutput.t90 4.06363
R14810 CSoutput.n95 CSoutput.t88 4.06363
R14811 CSoutput.n97 CSoutput.t83 4.06363
R14812 CSoutput.n97 CSoutput.t76 4.06363
R14813 CSoutput.n99 CSoutput.t89 4.06363
R14814 CSoutput.n99 CSoutput.t103 4.06363
R14815 CSoutput.n86 CSoutput.t92 4.06363
R14816 CSoutput.n86 CSoutput.t107 4.06363
R14817 CSoutput.n87 CSoutput.t101 4.06363
R14818 CSoutput.n87 CSoutput.t82 4.06363
R14819 CSoutput.n89 CSoutput.t87 4.06363
R14820 CSoutput.n89 CSoutput.t98 4.06363
R14821 CSoutput.n91 CSoutput.t100 4.06363
R14822 CSoutput.n91 CSoutput.t86 4.06363
R14823 CSoutput.n79 CSoutput.t94 4.06363
R14824 CSoutput.n79 CSoutput.t74 4.06363
R14825 CSoutput.n80 CSoutput.t111 4.06363
R14826 CSoutput.n80 CSoutput.t80 4.06363
R14827 CSoutput.n82 CSoutput.t99 4.06363
R14828 CSoutput.n82 CSoutput.t72 4.06363
R14829 CSoutput.n84 CSoutput.t116 4.06363
R14830 CSoutput.n84 CSoutput.t114 4.06363
R14831 CSoutput.n44 CSoutput.n43 3.79402
R14832 CSoutput.n49 CSoutput.n48 3.79402
R14833 CSoutput.n311 CSoutput.n299 3.72967
R14834 CSoutput.n347 CSoutput.n335 3.72967
R14835 CSoutput.n349 CSoutput.n348 3.57343
R14836 CSoutput.n348 CSoutput.n312 3.04641
R14837 CSoutput.n309 CSoutput.t44 2.82907
R14838 CSoutput.n309 CSoutput.t2 2.82907
R14839 CSoutput.n307 CSoutput.t70 2.82907
R14840 CSoutput.n307 CSoutput.t60 2.82907
R14841 CSoutput.n305 CSoutput.t26 2.82907
R14842 CSoutput.n305 CSoutput.t35 2.82907
R14843 CSoutput.n303 CSoutput.t1 2.82907
R14844 CSoutput.n303 CSoutput.t67 2.82907
R14845 CSoutput.n301 CSoutput.t59 2.82907
R14846 CSoutput.n301 CSoutput.t15 2.82907
R14847 CSoutput.n300 CSoutput.t8 2.82907
R14848 CSoutput.n300 CSoutput.t69 2.82907
R14849 CSoutput.n297 CSoutput.t12 2.82907
R14850 CSoutput.n297 CSoutput.t22 2.82907
R14851 CSoutput.n295 CSoutput.t21 2.82907
R14852 CSoutput.n295 CSoutput.t7 2.82907
R14853 CSoutput.n293 CSoutput.t33 2.82907
R14854 CSoutput.n293 CSoutput.t11 2.82907
R14855 CSoutput.n291 CSoutput.t14 2.82907
R14856 CSoutput.n291 CSoutput.t20 2.82907
R14857 CSoutput.n289 CSoutput.t18 2.82907
R14858 CSoutput.n289 CSoutput.t31 2.82907
R14859 CSoutput.n288 CSoutput.t30 2.82907
R14860 CSoutput.n288 CSoutput.t13 2.82907
R14861 CSoutput.n286 CSoutput.t53 2.82907
R14862 CSoutput.n286 CSoutput.t24 2.82907
R14863 CSoutput.n284 CSoutput.t4 2.82907
R14864 CSoutput.n284 CSoutput.t40 2.82907
R14865 CSoutput.n282 CSoutput.t19 2.82907
R14866 CSoutput.n282 CSoutput.t32 2.82907
R14867 CSoutput.n280 CSoutput.t34 2.82907
R14868 CSoutput.n280 CSoutput.t65 2.82907
R14869 CSoutput.n278 CSoutput.t50 2.82907
R14870 CSoutput.n278 CSoutput.t0 2.82907
R14871 CSoutput.n277 CSoutput.t63 2.82907
R14872 CSoutput.n277 CSoutput.t10 2.82907
R14873 CSoutput.n336 CSoutput.t57 2.82907
R14874 CSoutput.n336 CSoutput.t68 2.82907
R14875 CSoutput.n337 CSoutput.t71 2.82907
R14876 CSoutput.n337 CSoutput.t48 2.82907
R14877 CSoutput.n339 CSoutput.t52 2.82907
R14878 CSoutput.n339 CSoutput.t62 2.82907
R14879 CSoutput.n341 CSoutput.t9 2.82907
R14880 CSoutput.n341 CSoutput.t42 2.82907
R14881 CSoutput.n343 CSoutput.t47 2.82907
R14882 CSoutput.n343 CSoutput.t58 2.82907
R14883 CSoutput.n345 CSoutput.t64 2.82907
R14884 CSoutput.n345 CSoutput.t51 2.82907
R14885 CSoutput.n324 CSoutput.t28 2.82907
R14886 CSoutput.n324 CSoutput.t45 2.82907
R14887 CSoutput.n325 CSoutput.t46 2.82907
R14888 CSoutput.n325 CSoutput.t36 2.82907
R14889 CSoutput.n327 CSoutput.t37 2.82907
R14890 CSoutput.n327 CSoutput.t29 2.82907
R14891 CSoutput.n329 CSoutput.t23 2.82907
R14892 CSoutput.n329 CSoutput.t16 2.82907
R14893 CSoutput.n331 CSoutput.t17 2.82907
R14894 CSoutput.n331 CSoutput.t38 2.82907
R14895 CSoutput.n333 CSoutput.t39 2.82907
R14896 CSoutput.n333 CSoutput.t3 2.82907
R14897 CSoutput.n313 CSoutput.t41 2.82907
R14898 CSoutput.n313 CSoutput.t5 2.82907
R14899 CSoutput.n314 CSoutput.t25 2.82907
R14900 CSoutput.n314 CSoutput.t66 2.82907
R14901 CSoutput.n316 CSoutput.t6 2.82907
R14902 CSoutput.n316 CSoutput.t55 2.82907
R14903 CSoutput.n318 CSoutput.t54 2.82907
R14904 CSoutput.n318 CSoutput.t43 2.82907
R14905 CSoutput.n320 CSoutput.t56 2.82907
R14906 CSoutput.n320 CSoutput.t27 2.82907
R14907 CSoutput.n322 CSoutput.t49 2.82907
R14908 CSoutput.n322 CSoutput.t61 2.82907
R14909 CSoutput.n75 CSoutput.n1 2.45513
R14910 CSoutput.n193 CSoutput.n191 2.251
R14911 CSoutput.n193 CSoutput.n190 2.251
R14912 CSoutput.n193 CSoutput.n189 2.251
R14913 CSoutput.n193 CSoutput.n188 2.251
R14914 CSoutput.n162 CSoutput.n161 2.251
R14915 CSoutput.n162 CSoutput.n160 2.251
R14916 CSoutput.n162 CSoutput.n159 2.251
R14917 CSoutput.n162 CSoutput.n158 2.251
R14918 CSoutput.n235 CSoutput.n234 2.251
R14919 CSoutput.n200 CSoutput.n198 2.251
R14920 CSoutput.n200 CSoutput.n197 2.251
R14921 CSoutput.n200 CSoutput.n196 2.251
R14922 CSoutput.n218 CSoutput.n200 2.251
R14923 CSoutput.n206 CSoutput.n205 2.251
R14924 CSoutput.n206 CSoutput.n204 2.251
R14925 CSoutput.n206 CSoutput.n203 2.251
R14926 CSoutput.n206 CSoutput.n202 2.251
R14927 CSoutput.n232 CSoutput.n172 2.251
R14928 CSoutput.n227 CSoutput.n225 2.251
R14929 CSoutput.n227 CSoutput.n224 2.251
R14930 CSoutput.n227 CSoutput.n223 2.251
R14931 CSoutput.n227 CSoutput.n222 2.251
R14932 CSoutput.n128 CSoutput.n127 2.251
R14933 CSoutput.n128 CSoutput.n126 2.251
R14934 CSoutput.n128 CSoutput.n125 2.251
R14935 CSoutput.n128 CSoutput.n124 2.251
R14936 CSoutput.n245 CSoutput.n244 2.251
R14937 CSoutput.n162 CSoutput.n142 2.2505
R14938 CSoutput.n157 CSoutput.n142 2.2505
R14939 CSoutput.n155 CSoutput.n142 2.2505
R14940 CSoutput.n154 CSoutput.n142 2.2505
R14941 CSoutput.n239 CSoutput.n142 2.2505
R14942 CSoutput.n237 CSoutput.n142 2.2505
R14943 CSoutput.n235 CSoutput.n142 2.2505
R14944 CSoutput.n165 CSoutput.n142 2.2505
R14945 CSoutput.n164 CSoutput.n142 2.2505
R14946 CSoutput.n168 CSoutput.n142 2.2505
R14947 CSoutput.n167 CSoutput.n142 2.2505
R14948 CSoutput.n150 CSoutput.n142 2.2505
R14949 CSoutput.n242 CSoutput.n142 2.2505
R14950 CSoutput.n242 CSoutput.n241 2.2505
R14951 CSoutput.n206 CSoutput.n177 2.2505
R14952 CSoutput.n187 CSoutput.n177 2.2505
R14953 CSoutput.n208 CSoutput.n177 2.2505
R14954 CSoutput.n186 CSoutput.n177 2.2505
R14955 CSoutput.n210 CSoutput.n177 2.2505
R14956 CSoutput.n177 CSoutput.n171 2.2505
R14957 CSoutput.n232 CSoutput.n177 2.2505
R14958 CSoutput.n230 CSoutput.n177 2.2505
R14959 CSoutput.n212 CSoutput.n177 2.2505
R14960 CSoutput.n184 CSoutput.n177 2.2505
R14961 CSoutput.n214 CSoutput.n177 2.2505
R14962 CSoutput.n183 CSoutput.n177 2.2505
R14963 CSoutput.n228 CSoutput.n177 2.2505
R14964 CSoutput.n228 CSoutput.n181 2.2505
R14965 CSoutput.n128 CSoutput.n108 2.2505
R14966 CSoutput.n123 CSoutput.n108 2.2505
R14967 CSoutput.n121 CSoutput.n108 2.2505
R14968 CSoutput.n120 CSoutput.n108 2.2505
R14969 CSoutput.n249 CSoutput.n108 2.2505
R14970 CSoutput.n247 CSoutput.n108 2.2505
R14971 CSoutput.n245 CSoutput.n108 2.2505
R14972 CSoutput.n131 CSoutput.n108 2.2505
R14973 CSoutput.n130 CSoutput.n108 2.2505
R14974 CSoutput.n134 CSoutput.n108 2.2505
R14975 CSoutput.n133 CSoutput.n108 2.2505
R14976 CSoutput.n116 CSoutput.n108 2.2505
R14977 CSoutput.n252 CSoutput.n108 2.2505
R14978 CSoutput.n252 CSoutput.n251 2.2505
R14979 CSoutput.n170 CSoutput.n163 2.25024
R14980 CSoutput.n170 CSoutput.n156 2.25024
R14981 CSoutput.n238 CSoutput.n170 2.25024
R14982 CSoutput.n170 CSoutput.n166 2.25024
R14983 CSoutput.n170 CSoutput.n169 2.25024
R14984 CSoutput.n170 CSoutput.n137 2.25024
R14985 CSoutput.n220 CSoutput.n217 2.25024
R14986 CSoutput.n220 CSoutput.n216 2.25024
R14987 CSoutput.n220 CSoutput.n215 2.25024
R14988 CSoutput.n220 CSoutput.n182 2.25024
R14989 CSoutput.n220 CSoutput.n219 2.25024
R14990 CSoutput.n221 CSoutput.n220 2.25024
R14991 CSoutput.n136 CSoutput.n129 2.25024
R14992 CSoutput.n136 CSoutput.n122 2.25024
R14993 CSoutput.n248 CSoutput.n136 2.25024
R14994 CSoutput.n136 CSoutput.n132 2.25024
R14995 CSoutput.n136 CSoutput.n135 2.25024
R14996 CSoutput.n136 CSoutput.n103 2.25024
R14997 CSoutput.n276 CSoutput.n102 1.95131
R14998 CSoutput.n237 CSoutput.n147 1.50111
R14999 CSoutput.n185 CSoutput.n171 1.50111
R15000 CSoutput.n247 CSoutput.n113 1.50111
R15001 CSoutput.n193 CSoutput.n192 1.501
R15002 CSoutput.n200 CSoutput.n199 1.501
R15003 CSoutput.n227 CSoutput.n226 1.501
R15004 CSoutput.n241 CSoutput.n152 1.12536
R15005 CSoutput.n241 CSoutput.n153 1.12536
R15006 CSoutput.n241 CSoutput.n240 1.12536
R15007 CSoutput.n201 CSoutput.n181 1.12536
R15008 CSoutput.n207 CSoutput.n181 1.12536
R15009 CSoutput.n209 CSoutput.n181 1.12536
R15010 CSoutput.n251 CSoutput.n118 1.12536
R15011 CSoutput.n251 CSoutput.n119 1.12536
R15012 CSoutput.n251 CSoutput.n250 1.12536
R15013 CSoutput.n241 CSoutput.n148 1.12536
R15014 CSoutput.n241 CSoutput.n149 1.12536
R15015 CSoutput.n241 CSoutput.n151 1.12536
R15016 CSoutput.n231 CSoutput.n181 1.12536
R15017 CSoutput.n211 CSoutput.n181 1.12536
R15018 CSoutput.n213 CSoutput.n181 1.12536
R15019 CSoutput.n251 CSoutput.n114 1.12536
R15020 CSoutput.n251 CSoutput.n115 1.12536
R15021 CSoutput.n251 CSoutput.n117 1.12536
R15022 CSoutput.n31 CSoutput.n30 0.669944
R15023 CSoutput.n62 CSoutput.n61 0.669944
R15024 CSoutput.n304 CSoutput.n302 0.573776
R15025 CSoutput.n306 CSoutput.n304 0.573776
R15026 CSoutput.n308 CSoutput.n306 0.573776
R15027 CSoutput.n310 CSoutput.n308 0.573776
R15028 CSoutput.n292 CSoutput.n290 0.573776
R15029 CSoutput.n294 CSoutput.n292 0.573776
R15030 CSoutput.n296 CSoutput.n294 0.573776
R15031 CSoutput.n298 CSoutput.n296 0.573776
R15032 CSoutput.n281 CSoutput.n279 0.573776
R15033 CSoutput.n283 CSoutput.n281 0.573776
R15034 CSoutput.n285 CSoutput.n283 0.573776
R15035 CSoutput.n287 CSoutput.n285 0.573776
R15036 CSoutput.n346 CSoutput.n344 0.573776
R15037 CSoutput.n344 CSoutput.n342 0.573776
R15038 CSoutput.n342 CSoutput.n340 0.573776
R15039 CSoutput.n340 CSoutput.n338 0.573776
R15040 CSoutput.n334 CSoutput.n332 0.573776
R15041 CSoutput.n332 CSoutput.n330 0.573776
R15042 CSoutput.n330 CSoutput.n328 0.573776
R15043 CSoutput.n328 CSoutput.n326 0.573776
R15044 CSoutput.n323 CSoutput.n321 0.573776
R15045 CSoutput.n321 CSoutput.n319 0.573776
R15046 CSoutput.n319 CSoutput.n317 0.573776
R15047 CSoutput.n317 CSoutput.n315 0.573776
R15048 CSoutput.n349 CSoutput.n252 0.53442
R15049 CSoutput.n272 CSoutput.n270 0.358259
R15050 CSoutput.n274 CSoutput.n272 0.358259
R15051 CSoutput.n264 CSoutput.n262 0.358259
R15052 CSoutput.n266 CSoutput.n264 0.358259
R15053 CSoutput.n257 CSoutput.n255 0.358259
R15054 CSoutput.n259 CSoutput.n257 0.358259
R15055 CSoutput.n100 CSoutput.n98 0.358259
R15056 CSoutput.n98 CSoutput.n96 0.358259
R15057 CSoutput.n92 CSoutput.n90 0.358259
R15058 CSoutput.n90 CSoutput.n88 0.358259
R15059 CSoutput.n85 CSoutput.n83 0.358259
R15060 CSoutput.n83 CSoutput.n81 0.358259
R15061 CSoutput.n21 CSoutput.n20 0.169105
R15062 CSoutput.n21 CSoutput.n16 0.169105
R15063 CSoutput.n26 CSoutput.n16 0.169105
R15064 CSoutput.n27 CSoutput.n26 0.169105
R15065 CSoutput.n27 CSoutput.n14 0.169105
R15066 CSoutput.n32 CSoutput.n14 0.169105
R15067 CSoutput.n33 CSoutput.n32 0.169105
R15068 CSoutput.n34 CSoutput.n33 0.169105
R15069 CSoutput.n34 CSoutput.n12 0.169105
R15070 CSoutput.n39 CSoutput.n12 0.169105
R15071 CSoutput.n40 CSoutput.n39 0.169105
R15072 CSoutput.n40 CSoutput.n10 0.169105
R15073 CSoutput.n45 CSoutput.n10 0.169105
R15074 CSoutput.n46 CSoutput.n45 0.169105
R15075 CSoutput.n47 CSoutput.n46 0.169105
R15076 CSoutput.n47 CSoutput.n8 0.169105
R15077 CSoutput.n52 CSoutput.n8 0.169105
R15078 CSoutput.n53 CSoutput.n52 0.169105
R15079 CSoutput.n53 CSoutput.n6 0.169105
R15080 CSoutput.n58 CSoutput.n6 0.169105
R15081 CSoutput.n59 CSoutput.n58 0.169105
R15082 CSoutput.n60 CSoutput.n59 0.169105
R15083 CSoutput.n60 CSoutput.n4 0.169105
R15084 CSoutput.n66 CSoutput.n4 0.169105
R15085 CSoutput.n67 CSoutput.n66 0.169105
R15086 CSoutput.n68 CSoutput.n67 0.169105
R15087 CSoutput.n68 CSoutput.n2 0.169105
R15088 CSoutput.n73 CSoutput.n2 0.169105
R15089 CSoutput.n74 CSoutput.n73 0.169105
R15090 CSoutput.n74 CSoutput.n0 0.169105
R15091 CSoutput.n78 CSoutput.n0 0.169105
R15092 CSoutput.n195 CSoutput.n194 0.0910737
R15093 CSoutput.n246 CSoutput.n243 0.0723685
R15094 CSoutput.n200 CSoutput.n195 0.0522944
R15095 CSoutput.n243 CSoutput.n242 0.0499135
R15096 CSoutput.n194 CSoutput.n193 0.0499135
R15097 CSoutput.n228 CSoutput.n227 0.0464294
R15098 CSoutput.n236 CSoutput.n233 0.0391444
R15099 CSoutput.n195 CSoutput.t141 0.023435
R15100 CSoutput.n243 CSoutput.t121 0.02262
R15101 CSoutput.n194 CSoutput.t122 0.02262
R15102 CSoutput CSoutput.n349 0.0052
R15103 CSoutput.n165 CSoutput.n148 0.00365111
R15104 CSoutput.n168 CSoutput.n149 0.00365111
R15105 CSoutput.n151 CSoutput.n150 0.00365111
R15106 CSoutput.n193 CSoutput.n152 0.00365111
R15107 CSoutput.n157 CSoutput.n153 0.00365111
R15108 CSoutput.n240 CSoutput.n154 0.00365111
R15109 CSoutput.n231 CSoutput.n230 0.00365111
R15110 CSoutput.n211 CSoutput.n184 0.00365111
R15111 CSoutput.n213 CSoutput.n183 0.00365111
R15112 CSoutput.n201 CSoutput.n200 0.00365111
R15113 CSoutput.n207 CSoutput.n187 0.00365111
R15114 CSoutput.n209 CSoutput.n186 0.00365111
R15115 CSoutput.n131 CSoutput.n114 0.00365111
R15116 CSoutput.n134 CSoutput.n115 0.00365111
R15117 CSoutput.n117 CSoutput.n116 0.00365111
R15118 CSoutput.n227 CSoutput.n118 0.00365111
R15119 CSoutput.n123 CSoutput.n119 0.00365111
R15120 CSoutput.n250 CSoutput.n120 0.00365111
R15121 CSoutput.n162 CSoutput.n152 0.00340054
R15122 CSoutput.n155 CSoutput.n153 0.00340054
R15123 CSoutput.n240 CSoutput.n239 0.00340054
R15124 CSoutput.n235 CSoutput.n148 0.00340054
R15125 CSoutput.n164 CSoutput.n149 0.00340054
R15126 CSoutput.n167 CSoutput.n151 0.00340054
R15127 CSoutput.n206 CSoutput.n201 0.00340054
R15128 CSoutput.n208 CSoutput.n207 0.00340054
R15129 CSoutput.n210 CSoutput.n209 0.00340054
R15130 CSoutput.n232 CSoutput.n231 0.00340054
R15131 CSoutput.n212 CSoutput.n211 0.00340054
R15132 CSoutput.n214 CSoutput.n213 0.00340054
R15133 CSoutput.n128 CSoutput.n118 0.00340054
R15134 CSoutput.n121 CSoutput.n119 0.00340054
R15135 CSoutput.n250 CSoutput.n249 0.00340054
R15136 CSoutput.n245 CSoutput.n114 0.00340054
R15137 CSoutput.n130 CSoutput.n115 0.00340054
R15138 CSoutput.n133 CSoutput.n117 0.00340054
R15139 CSoutput.n163 CSoutput.n157 0.00252698
R15140 CSoutput.n156 CSoutput.n154 0.00252698
R15141 CSoutput.n238 CSoutput.n237 0.00252698
R15142 CSoutput.n166 CSoutput.n164 0.00252698
R15143 CSoutput.n169 CSoutput.n167 0.00252698
R15144 CSoutput.n242 CSoutput.n137 0.00252698
R15145 CSoutput.n163 CSoutput.n162 0.00252698
R15146 CSoutput.n156 CSoutput.n155 0.00252698
R15147 CSoutput.n239 CSoutput.n238 0.00252698
R15148 CSoutput.n166 CSoutput.n165 0.00252698
R15149 CSoutput.n169 CSoutput.n168 0.00252698
R15150 CSoutput.n150 CSoutput.n137 0.00252698
R15151 CSoutput.n217 CSoutput.n187 0.00252698
R15152 CSoutput.n216 CSoutput.n186 0.00252698
R15153 CSoutput.n215 CSoutput.n171 0.00252698
R15154 CSoutput.n212 CSoutput.n182 0.00252698
R15155 CSoutput.n219 CSoutput.n214 0.00252698
R15156 CSoutput.n228 CSoutput.n221 0.00252698
R15157 CSoutput.n217 CSoutput.n206 0.00252698
R15158 CSoutput.n216 CSoutput.n208 0.00252698
R15159 CSoutput.n215 CSoutput.n210 0.00252698
R15160 CSoutput.n230 CSoutput.n182 0.00252698
R15161 CSoutput.n219 CSoutput.n184 0.00252698
R15162 CSoutput.n221 CSoutput.n183 0.00252698
R15163 CSoutput.n129 CSoutput.n123 0.00252698
R15164 CSoutput.n122 CSoutput.n120 0.00252698
R15165 CSoutput.n248 CSoutput.n247 0.00252698
R15166 CSoutput.n132 CSoutput.n130 0.00252698
R15167 CSoutput.n135 CSoutput.n133 0.00252698
R15168 CSoutput.n252 CSoutput.n103 0.00252698
R15169 CSoutput.n129 CSoutput.n128 0.00252698
R15170 CSoutput.n122 CSoutput.n121 0.00252698
R15171 CSoutput.n249 CSoutput.n248 0.00252698
R15172 CSoutput.n132 CSoutput.n131 0.00252698
R15173 CSoutput.n135 CSoutput.n134 0.00252698
R15174 CSoutput.n116 CSoutput.n103 0.00252698
R15175 CSoutput.n237 CSoutput.n236 0.0020275
R15176 CSoutput.n236 CSoutput.n235 0.0020275
R15177 CSoutput.n233 CSoutput.n171 0.0020275
R15178 CSoutput.n233 CSoutput.n232 0.0020275
R15179 CSoutput.n247 CSoutput.n246 0.0020275
R15180 CSoutput.n246 CSoutput.n245 0.0020275
R15181 CSoutput.n147 CSoutput.n146 0.00166668
R15182 CSoutput.n229 CSoutput.n185 0.00166668
R15183 CSoutput.n113 CSoutput.n112 0.00166668
R15184 CSoutput.n251 CSoutput.n113 0.00133328
R15185 CSoutput.n185 CSoutput.n181 0.00133328
R15186 CSoutput.n241 CSoutput.n147 0.00133328
R15187 CSoutput.n244 CSoutput.n136 0.001
R15188 CSoutput.n222 CSoutput.n136 0.001
R15189 CSoutput.n124 CSoutput.n104 0.001
R15190 CSoutput.n223 CSoutput.n104 0.001
R15191 CSoutput.n125 CSoutput.n105 0.001
R15192 CSoutput.n224 CSoutput.n105 0.001
R15193 CSoutput.n126 CSoutput.n106 0.001
R15194 CSoutput.n225 CSoutput.n106 0.001
R15195 CSoutput.n127 CSoutput.n107 0.001
R15196 CSoutput.n226 CSoutput.n107 0.001
R15197 CSoutput.n220 CSoutput.n172 0.001
R15198 CSoutput.n220 CSoutput.n218 0.001
R15199 CSoutput.n202 CSoutput.n173 0.001
R15200 CSoutput.n196 CSoutput.n173 0.001
R15201 CSoutput.n203 CSoutput.n174 0.001
R15202 CSoutput.n197 CSoutput.n174 0.001
R15203 CSoutput.n204 CSoutput.n175 0.001
R15204 CSoutput.n198 CSoutput.n175 0.001
R15205 CSoutput.n205 CSoutput.n176 0.001
R15206 CSoutput.n199 CSoutput.n176 0.001
R15207 CSoutput.n234 CSoutput.n170 0.001
R15208 CSoutput.n188 CSoutput.n170 0.001
R15209 CSoutput.n158 CSoutput.n138 0.001
R15210 CSoutput.n189 CSoutput.n138 0.001
R15211 CSoutput.n159 CSoutput.n139 0.001
R15212 CSoutput.n190 CSoutput.n139 0.001
R15213 CSoutput.n160 CSoutput.n140 0.001
R15214 CSoutput.n191 CSoutput.n140 0.001
R15215 CSoutput.n161 CSoutput.n141 0.001
R15216 CSoutput.n192 CSoutput.n141 0.001
R15217 CSoutput.n192 CSoutput.n142 0.001
R15218 CSoutput.n191 CSoutput.n143 0.001
R15219 CSoutput.n190 CSoutput.n144 0.001
R15220 CSoutput.n189 CSoutput.t140 0.001
R15221 CSoutput.n188 CSoutput.n145 0.001
R15222 CSoutput.n161 CSoutput.n143 0.001
R15223 CSoutput.n160 CSoutput.n144 0.001
R15224 CSoutput.n159 CSoutput.t140 0.001
R15225 CSoutput.n158 CSoutput.n145 0.001
R15226 CSoutput.n234 CSoutput.n146 0.001
R15227 CSoutput.n199 CSoutput.n177 0.001
R15228 CSoutput.n198 CSoutput.n178 0.001
R15229 CSoutput.n197 CSoutput.n179 0.001
R15230 CSoutput.n196 CSoutput.t132 0.001
R15231 CSoutput.n218 CSoutput.n180 0.001
R15232 CSoutput.n205 CSoutput.n178 0.001
R15233 CSoutput.n204 CSoutput.n179 0.001
R15234 CSoutput.n203 CSoutput.t132 0.001
R15235 CSoutput.n202 CSoutput.n180 0.001
R15236 CSoutput.n229 CSoutput.n172 0.001
R15237 CSoutput.n226 CSoutput.n108 0.001
R15238 CSoutput.n225 CSoutput.n109 0.001
R15239 CSoutput.n224 CSoutput.n110 0.001
R15240 CSoutput.n223 CSoutput.t131 0.001
R15241 CSoutput.n222 CSoutput.n111 0.001
R15242 CSoutput.n127 CSoutput.n109 0.001
R15243 CSoutput.n126 CSoutput.n110 0.001
R15244 CSoutput.n125 CSoutput.t131 0.001
R15245 CSoutput.n124 CSoutput.n111 0.001
R15246 CSoutput.n244 CSoutput.n112 0.001
R15247 vdd.n291 vdd.n255 756.745
R15248 vdd.n244 vdd.n208 756.745
R15249 vdd.n201 vdd.n165 756.745
R15250 vdd.n154 vdd.n118 756.745
R15251 vdd.n112 vdd.n76 756.745
R15252 vdd.n65 vdd.n29 756.745
R15253 vdd.n1106 vdd.n1070 756.745
R15254 vdd.n1153 vdd.n1117 756.745
R15255 vdd.n1016 vdd.n980 756.745
R15256 vdd.n1063 vdd.n1027 756.745
R15257 vdd.n927 vdd.n891 756.745
R15258 vdd.n974 vdd.n938 756.745
R15259 vdd.n1791 vdd.t128 640.208
R15260 vdd.n755 vdd.t113 640.208
R15261 vdd.n1765 vdd.t154 640.208
R15262 vdd.n747 vdd.t145 640.208
R15263 vdd.n2536 vdd.t96 640.208
R15264 vdd.n2256 vdd.t136 640.208
R15265 vdd.n622 vdd.t117 640.208
R15266 vdd.n2253 vdd.t121 640.208
R15267 vdd.n589 vdd.t125 640.208
R15268 vdd.n817 vdd.t132 640.208
R15269 vdd.n1320 vdd.t92 592.009
R15270 vdd.n1358 vdd.t139 592.009
R15271 vdd.n1254 vdd.t142 592.009
R15272 vdd.n1947 vdd.t88 592.009
R15273 vdd.n1584 vdd.t100 592.009
R15274 vdd.n1544 vdd.t107 592.009
R15275 vdd.n2908 vdd.t151 592.009
R15276 vdd.n405 vdd.t103 592.009
R15277 vdd.n365 vdd.t110 592.009
R15278 vdd.n557 vdd.t81 592.009
R15279 vdd.n2804 vdd.t85 592.009
R15280 vdd.n2711 vdd.t148 592.009
R15281 vdd.n292 vdd.n291 585
R15282 vdd.n290 vdd.n257 585
R15283 vdd.n289 vdd.n288 585
R15284 vdd.n260 vdd.n258 585
R15285 vdd.n283 vdd.n282 585
R15286 vdd.n281 vdd.n280 585
R15287 vdd.n264 vdd.n263 585
R15288 vdd.n275 vdd.n274 585
R15289 vdd.n273 vdd.n272 585
R15290 vdd.n268 vdd.n267 585
R15291 vdd.n245 vdd.n244 585
R15292 vdd.n243 vdd.n210 585
R15293 vdd.n242 vdd.n241 585
R15294 vdd.n213 vdd.n211 585
R15295 vdd.n236 vdd.n235 585
R15296 vdd.n234 vdd.n233 585
R15297 vdd.n217 vdd.n216 585
R15298 vdd.n228 vdd.n227 585
R15299 vdd.n226 vdd.n225 585
R15300 vdd.n221 vdd.n220 585
R15301 vdd.n202 vdd.n201 585
R15302 vdd.n200 vdd.n167 585
R15303 vdd.n199 vdd.n198 585
R15304 vdd.n170 vdd.n168 585
R15305 vdd.n193 vdd.n192 585
R15306 vdd.n191 vdd.n190 585
R15307 vdd.n174 vdd.n173 585
R15308 vdd.n185 vdd.n184 585
R15309 vdd.n183 vdd.n182 585
R15310 vdd.n178 vdd.n177 585
R15311 vdd.n155 vdd.n154 585
R15312 vdd.n153 vdd.n120 585
R15313 vdd.n152 vdd.n151 585
R15314 vdd.n123 vdd.n121 585
R15315 vdd.n146 vdd.n145 585
R15316 vdd.n144 vdd.n143 585
R15317 vdd.n127 vdd.n126 585
R15318 vdd.n138 vdd.n137 585
R15319 vdd.n136 vdd.n135 585
R15320 vdd.n131 vdd.n130 585
R15321 vdd.n113 vdd.n112 585
R15322 vdd.n111 vdd.n78 585
R15323 vdd.n110 vdd.n109 585
R15324 vdd.n81 vdd.n79 585
R15325 vdd.n104 vdd.n103 585
R15326 vdd.n102 vdd.n101 585
R15327 vdd.n85 vdd.n84 585
R15328 vdd.n96 vdd.n95 585
R15329 vdd.n94 vdd.n93 585
R15330 vdd.n89 vdd.n88 585
R15331 vdd.n66 vdd.n65 585
R15332 vdd.n64 vdd.n31 585
R15333 vdd.n63 vdd.n62 585
R15334 vdd.n34 vdd.n32 585
R15335 vdd.n57 vdd.n56 585
R15336 vdd.n55 vdd.n54 585
R15337 vdd.n38 vdd.n37 585
R15338 vdd.n49 vdd.n48 585
R15339 vdd.n47 vdd.n46 585
R15340 vdd.n42 vdd.n41 585
R15341 vdd.n1107 vdd.n1106 585
R15342 vdd.n1105 vdd.n1072 585
R15343 vdd.n1104 vdd.n1103 585
R15344 vdd.n1075 vdd.n1073 585
R15345 vdd.n1098 vdd.n1097 585
R15346 vdd.n1096 vdd.n1095 585
R15347 vdd.n1079 vdd.n1078 585
R15348 vdd.n1090 vdd.n1089 585
R15349 vdd.n1088 vdd.n1087 585
R15350 vdd.n1083 vdd.n1082 585
R15351 vdd.n1154 vdd.n1153 585
R15352 vdd.n1152 vdd.n1119 585
R15353 vdd.n1151 vdd.n1150 585
R15354 vdd.n1122 vdd.n1120 585
R15355 vdd.n1145 vdd.n1144 585
R15356 vdd.n1143 vdd.n1142 585
R15357 vdd.n1126 vdd.n1125 585
R15358 vdd.n1137 vdd.n1136 585
R15359 vdd.n1135 vdd.n1134 585
R15360 vdd.n1130 vdd.n1129 585
R15361 vdd.n1017 vdd.n1016 585
R15362 vdd.n1015 vdd.n982 585
R15363 vdd.n1014 vdd.n1013 585
R15364 vdd.n985 vdd.n983 585
R15365 vdd.n1008 vdd.n1007 585
R15366 vdd.n1006 vdd.n1005 585
R15367 vdd.n989 vdd.n988 585
R15368 vdd.n1000 vdd.n999 585
R15369 vdd.n998 vdd.n997 585
R15370 vdd.n993 vdd.n992 585
R15371 vdd.n1064 vdd.n1063 585
R15372 vdd.n1062 vdd.n1029 585
R15373 vdd.n1061 vdd.n1060 585
R15374 vdd.n1032 vdd.n1030 585
R15375 vdd.n1055 vdd.n1054 585
R15376 vdd.n1053 vdd.n1052 585
R15377 vdd.n1036 vdd.n1035 585
R15378 vdd.n1047 vdd.n1046 585
R15379 vdd.n1045 vdd.n1044 585
R15380 vdd.n1040 vdd.n1039 585
R15381 vdd.n928 vdd.n927 585
R15382 vdd.n926 vdd.n893 585
R15383 vdd.n925 vdd.n924 585
R15384 vdd.n896 vdd.n894 585
R15385 vdd.n919 vdd.n918 585
R15386 vdd.n917 vdd.n916 585
R15387 vdd.n900 vdd.n899 585
R15388 vdd.n911 vdd.n910 585
R15389 vdd.n909 vdd.n908 585
R15390 vdd.n904 vdd.n903 585
R15391 vdd.n975 vdd.n974 585
R15392 vdd.n973 vdd.n940 585
R15393 vdd.n972 vdd.n971 585
R15394 vdd.n943 vdd.n941 585
R15395 vdd.n966 vdd.n965 585
R15396 vdd.n964 vdd.n963 585
R15397 vdd.n947 vdd.n946 585
R15398 vdd.n958 vdd.n957 585
R15399 vdd.n956 vdd.n955 585
R15400 vdd.n951 vdd.n950 585
R15401 vdd.n3024 vdd.n330 515.122
R15402 vdd.n2906 vdd.n328 515.122
R15403 vdd.n515 vdd.n478 515.122
R15404 vdd.n2842 vdd.n479 515.122
R15405 vdd.n1942 vdd.n865 515.122
R15406 vdd.n1945 vdd.n1944 515.122
R15407 vdd.n1227 vdd.n1191 515.122
R15408 vdd.n1423 vdd.n1192 515.122
R15409 vdd.n269 vdd.t34 329.043
R15410 vdd.n222 vdd.t45 329.043
R15411 vdd.n179 vdd.t30 329.043
R15412 vdd.n132 vdd.t40 329.043
R15413 vdd.n90 vdd.t71 329.043
R15414 vdd.n43 vdd.t13 329.043
R15415 vdd.n1084 vdd.t69 329.043
R15416 vdd.n1131 vdd.t55 329.043
R15417 vdd.n994 vdd.t61 329.043
R15418 vdd.n1041 vdd.t48 329.043
R15419 vdd.n905 vdd.t11 329.043
R15420 vdd.n952 vdd.t70 329.043
R15421 vdd.n1320 vdd.t95 319.788
R15422 vdd.n1358 vdd.t141 319.788
R15423 vdd.n1254 vdd.t144 319.788
R15424 vdd.n1947 vdd.t90 319.788
R15425 vdd.n1584 vdd.t101 319.788
R15426 vdd.n1544 vdd.t108 319.788
R15427 vdd.n2908 vdd.t152 319.788
R15428 vdd.n405 vdd.t105 319.788
R15429 vdd.n365 vdd.t111 319.788
R15430 vdd.n557 vdd.t84 319.788
R15431 vdd.n2804 vdd.t87 319.788
R15432 vdd.n2711 vdd.t150 319.788
R15433 vdd.n1321 vdd.t94 303.69
R15434 vdd.n1359 vdd.t140 303.69
R15435 vdd.n1255 vdd.t143 303.69
R15436 vdd.n1948 vdd.t91 303.69
R15437 vdd.n1585 vdd.t102 303.69
R15438 vdd.n1545 vdd.t109 303.69
R15439 vdd.n2909 vdd.t153 303.69
R15440 vdd.n406 vdd.t106 303.69
R15441 vdd.n366 vdd.t112 303.69
R15442 vdd.n558 vdd.t83 303.69
R15443 vdd.n2805 vdd.t86 303.69
R15444 vdd.n2712 vdd.t149 303.69
R15445 vdd.n2479 vdd.n703 297.074
R15446 vdd.n2672 vdd.n599 297.074
R15447 vdd.n2609 vdd.n596 297.074
R15448 vdd.n2402 vdd.n704 297.074
R15449 vdd.n2217 vdd.n744 297.074
R15450 vdd.n2148 vdd.n2147 297.074
R15451 vdd.n1894 vdd.n840 297.074
R15452 vdd.n1990 vdd.n838 297.074
R15453 vdd.n2588 vdd.n597 297.074
R15454 vdd.n2675 vdd.n2674 297.074
R15455 vdd.n2251 vdd.n705 297.074
R15456 vdd.n2477 vdd.n706 297.074
R15457 vdd.n2145 vdd.n753 297.074
R15458 vdd.n751 vdd.n726 297.074
R15459 vdd.n1831 vdd.n841 297.074
R15460 vdd.n1988 vdd.n842 297.074
R15461 vdd.n2590 vdd.n597 185
R15462 vdd.n2673 vdd.n597 185
R15463 vdd.n2592 vdd.n2591 185
R15464 vdd.n2591 vdd.n595 185
R15465 vdd.n2593 vdd.n629 185
R15466 vdd.n2603 vdd.n629 185
R15467 vdd.n2594 vdd.n638 185
R15468 vdd.n638 vdd.n636 185
R15469 vdd.n2596 vdd.n2595 185
R15470 vdd.n2597 vdd.n2596 185
R15471 vdd.n2549 vdd.n637 185
R15472 vdd.n637 vdd.n633 185
R15473 vdd.n2548 vdd.n2547 185
R15474 vdd.n2547 vdd.n2546 185
R15475 vdd.n640 vdd.n639 185
R15476 vdd.n641 vdd.n640 185
R15477 vdd.n2539 vdd.n2538 185
R15478 vdd.n2540 vdd.n2539 185
R15479 vdd.n2535 vdd.n650 185
R15480 vdd.n650 vdd.n647 185
R15481 vdd.n2534 vdd.n2533 185
R15482 vdd.n2533 vdd.n2532 185
R15483 vdd.n652 vdd.n651 185
R15484 vdd.n660 vdd.n652 185
R15485 vdd.n2525 vdd.n2524 185
R15486 vdd.n2526 vdd.n2525 185
R15487 vdd.n2523 vdd.n661 185
R15488 vdd.n2374 vdd.n661 185
R15489 vdd.n2522 vdd.n2521 185
R15490 vdd.n2521 vdd.n2520 185
R15491 vdd.n663 vdd.n662 185
R15492 vdd.n664 vdd.n663 185
R15493 vdd.n2513 vdd.n2512 185
R15494 vdd.n2514 vdd.n2513 185
R15495 vdd.n2511 vdd.n673 185
R15496 vdd.n673 vdd.n670 185
R15497 vdd.n2510 vdd.n2509 185
R15498 vdd.n2509 vdd.n2508 185
R15499 vdd.n675 vdd.n674 185
R15500 vdd.n683 vdd.n675 185
R15501 vdd.n2501 vdd.n2500 185
R15502 vdd.n2502 vdd.n2501 185
R15503 vdd.n2499 vdd.n684 185
R15504 vdd.n690 vdd.n684 185
R15505 vdd.n2498 vdd.n2497 185
R15506 vdd.n2497 vdd.n2496 185
R15507 vdd.n686 vdd.n685 185
R15508 vdd.n687 vdd.n686 185
R15509 vdd.n2489 vdd.n2488 185
R15510 vdd.n2490 vdd.n2489 185
R15511 vdd.n2487 vdd.n696 185
R15512 vdd.n2395 vdd.n696 185
R15513 vdd.n2486 vdd.n2485 185
R15514 vdd.n2485 vdd.n2484 185
R15515 vdd.n698 vdd.n697 185
R15516 vdd.t198 vdd.n698 185
R15517 vdd.n2477 vdd.n2476 185
R15518 vdd.n2478 vdd.n2477 185
R15519 vdd.n2475 vdd.n706 185
R15520 vdd.n2474 vdd.n2473 185
R15521 vdd.n708 vdd.n707 185
R15522 vdd.n2260 vdd.n2259 185
R15523 vdd.n2262 vdd.n2261 185
R15524 vdd.n2264 vdd.n2263 185
R15525 vdd.n2266 vdd.n2265 185
R15526 vdd.n2268 vdd.n2267 185
R15527 vdd.n2270 vdd.n2269 185
R15528 vdd.n2272 vdd.n2271 185
R15529 vdd.n2274 vdd.n2273 185
R15530 vdd.n2276 vdd.n2275 185
R15531 vdd.n2278 vdd.n2277 185
R15532 vdd.n2280 vdd.n2279 185
R15533 vdd.n2282 vdd.n2281 185
R15534 vdd.n2284 vdd.n2283 185
R15535 vdd.n2286 vdd.n2285 185
R15536 vdd.n2288 vdd.n2287 185
R15537 vdd.n2290 vdd.n2289 185
R15538 vdd.n2292 vdd.n2291 185
R15539 vdd.n2294 vdd.n2293 185
R15540 vdd.n2296 vdd.n2295 185
R15541 vdd.n2298 vdd.n2297 185
R15542 vdd.n2300 vdd.n2299 185
R15543 vdd.n2302 vdd.n2301 185
R15544 vdd.n2304 vdd.n2303 185
R15545 vdd.n2306 vdd.n2305 185
R15546 vdd.n2308 vdd.n2307 185
R15547 vdd.n2310 vdd.n2309 185
R15548 vdd.n2312 vdd.n2311 185
R15549 vdd.n2314 vdd.n2313 185
R15550 vdd.n2316 vdd.n2315 185
R15551 vdd.n2318 vdd.n2317 185
R15552 vdd.n2320 vdd.n2319 185
R15553 vdd.n2321 vdd.n2251 185
R15554 vdd.n2471 vdd.n2251 185
R15555 vdd.n2676 vdd.n2675 185
R15556 vdd.n2677 vdd.n588 185
R15557 vdd.n2679 vdd.n2678 185
R15558 vdd.n2681 vdd.n586 185
R15559 vdd.n2683 vdd.n2682 185
R15560 vdd.n2684 vdd.n585 185
R15561 vdd.n2686 vdd.n2685 185
R15562 vdd.n2688 vdd.n583 185
R15563 vdd.n2690 vdd.n2689 185
R15564 vdd.n2691 vdd.n582 185
R15565 vdd.n2693 vdd.n2692 185
R15566 vdd.n2695 vdd.n580 185
R15567 vdd.n2697 vdd.n2696 185
R15568 vdd.n2698 vdd.n579 185
R15569 vdd.n2700 vdd.n2699 185
R15570 vdd.n2702 vdd.n578 185
R15571 vdd.n2703 vdd.n576 185
R15572 vdd.n2706 vdd.n2705 185
R15573 vdd.n577 vdd.n575 185
R15574 vdd.n2562 vdd.n2561 185
R15575 vdd.n2564 vdd.n2563 185
R15576 vdd.n2566 vdd.n2558 185
R15577 vdd.n2568 vdd.n2567 185
R15578 vdd.n2569 vdd.n2557 185
R15579 vdd.n2571 vdd.n2570 185
R15580 vdd.n2573 vdd.n2555 185
R15581 vdd.n2575 vdd.n2574 185
R15582 vdd.n2576 vdd.n2554 185
R15583 vdd.n2578 vdd.n2577 185
R15584 vdd.n2580 vdd.n2552 185
R15585 vdd.n2582 vdd.n2581 185
R15586 vdd.n2583 vdd.n2551 185
R15587 vdd.n2585 vdd.n2584 185
R15588 vdd.n2587 vdd.n2550 185
R15589 vdd.n2589 vdd.n2588 185
R15590 vdd.n2588 vdd.n484 185
R15591 vdd.n2674 vdd.n592 185
R15592 vdd.n2674 vdd.n2673 185
R15593 vdd.n2326 vdd.n594 185
R15594 vdd.n595 vdd.n594 185
R15595 vdd.n2327 vdd.n628 185
R15596 vdd.n2603 vdd.n628 185
R15597 vdd.n2329 vdd.n2328 185
R15598 vdd.n2328 vdd.n636 185
R15599 vdd.n2330 vdd.n635 185
R15600 vdd.n2597 vdd.n635 185
R15601 vdd.n2332 vdd.n2331 185
R15602 vdd.n2331 vdd.n633 185
R15603 vdd.n2333 vdd.n643 185
R15604 vdd.n2546 vdd.n643 185
R15605 vdd.n2335 vdd.n2334 185
R15606 vdd.n2334 vdd.n641 185
R15607 vdd.n2336 vdd.n649 185
R15608 vdd.n2540 vdd.n649 185
R15609 vdd.n2338 vdd.n2337 185
R15610 vdd.n2337 vdd.n647 185
R15611 vdd.n2339 vdd.n654 185
R15612 vdd.n2532 vdd.n654 185
R15613 vdd.n2341 vdd.n2340 185
R15614 vdd.n2340 vdd.n660 185
R15615 vdd.n2342 vdd.n659 185
R15616 vdd.n2526 vdd.n659 185
R15617 vdd.n2376 vdd.n2375 185
R15618 vdd.n2375 vdd.n2374 185
R15619 vdd.n2377 vdd.n666 185
R15620 vdd.n2520 vdd.n666 185
R15621 vdd.n2379 vdd.n2378 185
R15622 vdd.n2378 vdd.n664 185
R15623 vdd.n2380 vdd.n672 185
R15624 vdd.n2514 vdd.n672 185
R15625 vdd.n2382 vdd.n2381 185
R15626 vdd.n2381 vdd.n670 185
R15627 vdd.n2383 vdd.n677 185
R15628 vdd.n2508 vdd.n677 185
R15629 vdd.n2385 vdd.n2384 185
R15630 vdd.n2384 vdd.n683 185
R15631 vdd.n2386 vdd.n682 185
R15632 vdd.n2502 vdd.n682 185
R15633 vdd.n2388 vdd.n2387 185
R15634 vdd.n2387 vdd.n690 185
R15635 vdd.n2389 vdd.n689 185
R15636 vdd.n2496 vdd.n689 185
R15637 vdd.n2391 vdd.n2390 185
R15638 vdd.n2390 vdd.n687 185
R15639 vdd.n2392 vdd.n695 185
R15640 vdd.n2490 vdd.n695 185
R15641 vdd.n2394 vdd.n2393 185
R15642 vdd.n2395 vdd.n2394 185
R15643 vdd.n2325 vdd.n700 185
R15644 vdd.n2484 vdd.n700 185
R15645 vdd.n2324 vdd.n2323 185
R15646 vdd.n2323 vdd.t198 185
R15647 vdd.n2322 vdd.n705 185
R15648 vdd.n2478 vdd.n705 185
R15649 vdd.n1942 vdd.n1941 185
R15650 vdd.n1943 vdd.n1942 185
R15651 vdd.n866 vdd.n864 185
R15652 vdd.n1508 vdd.n864 185
R15653 vdd.n1511 vdd.n1510 185
R15654 vdd.n1510 vdd.n1509 185
R15655 vdd.n869 vdd.n868 185
R15656 vdd.n870 vdd.n869 185
R15657 vdd.n1497 vdd.n1496 185
R15658 vdd.n1498 vdd.n1497 185
R15659 vdd.n878 vdd.n877 185
R15660 vdd.n1489 vdd.n877 185
R15661 vdd.n1492 vdd.n1491 185
R15662 vdd.n1491 vdd.n1490 185
R15663 vdd.n881 vdd.n880 185
R15664 vdd.n888 vdd.n881 185
R15665 vdd.n1480 vdd.n1479 185
R15666 vdd.n1481 vdd.n1480 185
R15667 vdd.n890 vdd.n889 185
R15668 vdd.n889 vdd.n887 185
R15669 vdd.n1475 vdd.n1474 185
R15670 vdd.n1474 vdd.n1473 185
R15671 vdd.n1163 vdd.n1162 185
R15672 vdd.n1164 vdd.n1163 185
R15673 vdd.n1464 vdd.n1463 185
R15674 vdd.n1465 vdd.n1464 185
R15675 vdd.n1171 vdd.n1170 185
R15676 vdd.n1455 vdd.n1170 185
R15677 vdd.n1458 vdd.n1457 185
R15678 vdd.n1457 vdd.n1456 185
R15679 vdd.n1174 vdd.n1173 185
R15680 vdd.n1180 vdd.n1174 185
R15681 vdd.n1446 vdd.n1445 185
R15682 vdd.n1447 vdd.n1446 185
R15683 vdd.n1182 vdd.n1181 185
R15684 vdd.n1438 vdd.n1181 185
R15685 vdd.n1441 vdd.n1440 185
R15686 vdd.n1440 vdd.n1439 185
R15687 vdd.n1185 vdd.n1184 185
R15688 vdd.n1186 vdd.n1185 185
R15689 vdd.n1429 vdd.n1428 185
R15690 vdd.n1430 vdd.n1429 185
R15691 vdd.n1193 vdd.n1192 185
R15692 vdd.n1228 vdd.n1192 185
R15693 vdd.n1424 vdd.n1423 185
R15694 vdd.n1196 vdd.n1195 185
R15695 vdd.n1420 vdd.n1419 185
R15696 vdd.n1421 vdd.n1420 185
R15697 vdd.n1230 vdd.n1229 185
R15698 vdd.n1415 vdd.n1232 185
R15699 vdd.n1414 vdd.n1233 185
R15700 vdd.n1413 vdd.n1234 185
R15701 vdd.n1236 vdd.n1235 185
R15702 vdd.n1409 vdd.n1238 185
R15703 vdd.n1408 vdd.n1239 185
R15704 vdd.n1407 vdd.n1240 185
R15705 vdd.n1242 vdd.n1241 185
R15706 vdd.n1403 vdd.n1244 185
R15707 vdd.n1402 vdd.n1245 185
R15708 vdd.n1401 vdd.n1246 185
R15709 vdd.n1248 vdd.n1247 185
R15710 vdd.n1397 vdd.n1250 185
R15711 vdd.n1396 vdd.n1251 185
R15712 vdd.n1395 vdd.n1252 185
R15713 vdd.n1256 vdd.n1253 185
R15714 vdd.n1391 vdd.n1258 185
R15715 vdd.n1390 vdd.n1259 185
R15716 vdd.n1389 vdd.n1260 185
R15717 vdd.n1262 vdd.n1261 185
R15718 vdd.n1385 vdd.n1264 185
R15719 vdd.n1384 vdd.n1265 185
R15720 vdd.n1383 vdd.n1266 185
R15721 vdd.n1268 vdd.n1267 185
R15722 vdd.n1379 vdd.n1270 185
R15723 vdd.n1378 vdd.n1271 185
R15724 vdd.n1377 vdd.n1272 185
R15725 vdd.n1274 vdd.n1273 185
R15726 vdd.n1373 vdd.n1276 185
R15727 vdd.n1372 vdd.n1277 185
R15728 vdd.n1371 vdd.n1278 185
R15729 vdd.n1280 vdd.n1279 185
R15730 vdd.n1367 vdd.n1282 185
R15731 vdd.n1366 vdd.n1283 185
R15732 vdd.n1365 vdd.n1284 185
R15733 vdd.n1286 vdd.n1285 185
R15734 vdd.n1361 vdd.n1288 185
R15735 vdd.n1360 vdd.n1357 185
R15736 vdd.n1356 vdd.n1289 185
R15737 vdd.n1291 vdd.n1290 185
R15738 vdd.n1352 vdd.n1293 185
R15739 vdd.n1351 vdd.n1294 185
R15740 vdd.n1350 vdd.n1295 185
R15741 vdd.n1297 vdd.n1296 185
R15742 vdd.n1346 vdd.n1299 185
R15743 vdd.n1345 vdd.n1300 185
R15744 vdd.n1344 vdd.n1301 185
R15745 vdd.n1303 vdd.n1302 185
R15746 vdd.n1340 vdd.n1305 185
R15747 vdd.n1339 vdd.n1306 185
R15748 vdd.n1338 vdd.n1307 185
R15749 vdd.n1309 vdd.n1308 185
R15750 vdd.n1334 vdd.n1311 185
R15751 vdd.n1333 vdd.n1312 185
R15752 vdd.n1332 vdd.n1313 185
R15753 vdd.n1315 vdd.n1314 185
R15754 vdd.n1328 vdd.n1317 185
R15755 vdd.n1327 vdd.n1318 185
R15756 vdd.n1326 vdd.n1319 185
R15757 vdd.n1323 vdd.n1227 185
R15758 vdd.n1421 vdd.n1227 185
R15759 vdd.n1946 vdd.n1945 185
R15760 vdd.n1950 vdd.n859 185
R15761 vdd.n1613 vdd.n858 185
R15762 vdd.n1616 vdd.n1615 185
R15763 vdd.n1618 vdd.n1617 185
R15764 vdd.n1621 vdd.n1620 185
R15765 vdd.n1623 vdd.n1622 185
R15766 vdd.n1625 vdd.n1611 185
R15767 vdd.n1627 vdd.n1626 185
R15768 vdd.n1628 vdd.n1605 185
R15769 vdd.n1630 vdd.n1629 185
R15770 vdd.n1632 vdd.n1603 185
R15771 vdd.n1634 vdd.n1633 185
R15772 vdd.n1635 vdd.n1598 185
R15773 vdd.n1637 vdd.n1636 185
R15774 vdd.n1639 vdd.n1596 185
R15775 vdd.n1641 vdd.n1640 185
R15776 vdd.n1642 vdd.n1592 185
R15777 vdd.n1644 vdd.n1643 185
R15778 vdd.n1646 vdd.n1589 185
R15779 vdd.n1648 vdd.n1647 185
R15780 vdd.n1590 vdd.n1583 185
R15781 vdd.n1652 vdd.n1587 185
R15782 vdd.n1653 vdd.n1579 185
R15783 vdd.n1655 vdd.n1654 185
R15784 vdd.n1657 vdd.n1577 185
R15785 vdd.n1659 vdd.n1658 185
R15786 vdd.n1660 vdd.n1572 185
R15787 vdd.n1662 vdd.n1661 185
R15788 vdd.n1664 vdd.n1570 185
R15789 vdd.n1666 vdd.n1665 185
R15790 vdd.n1667 vdd.n1565 185
R15791 vdd.n1669 vdd.n1668 185
R15792 vdd.n1671 vdd.n1563 185
R15793 vdd.n1673 vdd.n1672 185
R15794 vdd.n1674 vdd.n1558 185
R15795 vdd.n1676 vdd.n1675 185
R15796 vdd.n1678 vdd.n1556 185
R15797 vdd.n1680 vdd.n1679 185
R15798 vdd.n1681 vdd.n1552 185
R15799 vdd.n1683 vdd.n1682 185
R15800 vdd.n1685 vdd.n1549 185
R15801 vdd.n1687 vdd.n1686 185
R15802 vdd.n1550 vdd.n1543 185
R15803 vdd.n1691 vdd.n1547 185
R15804 vdd.n1692 vdd.n1539 185
R15805 vdd.n1694 vdd.n1693 185
R15806 vdd.n1696 vdd.n1537 185
R15807 vdd.n1698 vdd.n1697 185
R15808 vdd.n1699 vdd.n1532 185
R15809 vdd.n1701 vdd.n1700 185
R15810 vdd.n1703 vdd.n1530 185
R15811 vdd.n1705 vdd.n1704 185
R15812 vdd.n1706 vdd.n1525 185
R15813 vdd.n1708 vdd.n1707 185
R15814 vdd.n1710 vdd.n1524 185
R15815 vdd.n1711 vdd.n1521 185
R15816 vdd.n1714 vdd.n1713 185
R15817 vdd.n1523 vdd.n1519 185
R15818 vdd.n1931 vdd.n1517 185
R15819 vdd.n1933 vdd.n1932 185
R15820 vdd.n1935 vdd.n1515 185
R15821 vdd.n1937 vdd.n1936 185
R15822 vdd.n1938 vdd.n865 185
R15823 vdd.n1944 vdd.n862 185
R15824 vdd.n1944 vdd.n1943 185
R15825 vdd.n873 vdd.n861 185
R15826 vdd.n1508 vdd.n861 185
R15827 vdd.n1507 vdd.n1506 185
R15828 vdd.n1509 vdd.n1507 185
R15829 vdd.n872 vdd.n871 185
R15830 vdd.n871 vdd.n870 185
R15831 vdd.n1500 vdd.n1499 185
R15832 vdd.n1499 vdd.n1498 185
R15833 vdd.n876 vdd.n875 185
R15834 vdd.n1489 vdd.n876 185
R15835 vdd.n1488 vdd.n1487 185
R15836 vdd.n1490 vdd.n1488 185
R15837 vdd.n883 vdd.n882 185
R15838 vdd.n888 vdd.n882 185
R15839 vdd.n1483 vdd.n1482 185
R15840 vdd.n1482 vdd.n1481 185
R15841 vdd.n886 vdd.n885 185
R15842 vdd.n887 vdd.n886 185
R15843 vdd.n1472 vdd.n1471 185
R15844 vdd.n1473 vdd.n1472 185
R15845 vdd.n1166 vdd.n1165 185
R15846 vdd.n1165 vdd.n1164 185
R15847 vdd.n1467 vdd.n1466 185
R15848 vdd.n1466 vdd.n1465 185
R15849 vdd.n1169 vdd.n1168 185
R15850 vdd.n1455 vdd.n1169 185
R15851 vdd.n1454 vdd.n1453 185
R15852 vdd.n1456 vdd.n1454 185
R15853 vdd.n1176 vdd.n1175 185
R15854 vdd.n1180 vdd.n1175 185
R15855 vdd.n1449 vdd.n1448 185
R15856 vdd.n1448 vdd.n1447 185
R15857 vdd.n1179 vdd.n1178 185
R15858 vdd.n1438 vdd.n1179 185
R15859 vdd.n1437 vdd.n1436 185
R15860 vdd.n1439 vdd.n1437 185
R15861 vdd.n1188 vdd.n1187 185
R15862 vdd.n1187 vdd.n1186 185
R15863 vdd.n1432 vdd.n1431 185
R15864 vdd.n1431 vdd.n1430 185
R15865 vdd.n1191 vdd.n1190 185
R15866 vdd.n1228 vdd.n1191 185
R15867 vdd.n746 vdd.n744 185
R15868 vdd.n2146 vdd.n744 185
R15869 vdd.n2068 vdd.n763 185
R15870 vdd.n763 vdd.t2 185
R15871 vdd.n2070 vdd.n2069 185
R15872 vdd.n2071 vdd.n2070 185
R15873 vdd.n2067 vdd.n762 185
R15874 vdd.n1770 vdd.n762 185
R15875 vdd.n2066 vdd.n2065 185
R15876 vdd.n2065 vdd.n2064 185
R15877 vdd.n765 vdd.n764 185
R15878 vdd.n766 vdd.n765 185
R15879 vdd.n2055 vdd.n2054 185
R15880 vdd.n2056 vdd.n2055 185
R15881 vdd.n2053 vdd.n776 185
R15882 vdd.n776 vdd.n773 185
R15883 vdd.n2052 vdd.n2051 185
R15884 vdd.n2051 vdd.n2050 185
R15885 vdd.n778 vdd.n777 185
R15886 vdd.n779 vdd.n778 185
R15887 vdd.n2043 vdd.n2042 185
R15888 vdd.n2044 vdd.n2043 185
R15889 vdd.n2041 vdd.n787 185
R15890 vdd.n792 vdd.n787 185
R15891 vdd.n2040 vdd.n2039 185
R15892 vdd.n2039 vdd.n2038 185
R15893 vdd.n789 vdd.n788 185
R15894 vdd.n798 vdd.n789 185
R15895 vdd.n2031 vdd.n2030 185
R15896 vdd.n2032 vdd.n2031 185
R15897 vdd.n2029 vdd.n799 185
R15898 vdd.n1871 vdd.n799 185
R15899 vdd.n2028 vdd.n2027 185
R15900 vdd.n2027 vdd.n2026 185
R15901 vdd.n801 vdd.n800 185
R15902 vdd.n802 vdd.n801 185
R15903 vdd.n2019 vdd.n2018 185
R15904 vdd.n2020 vdd.n2019 185
R15905 vdd.n2017 vdd.n811 185
R15906 vdd.n811 vdd.n808 185
R15907 vdd.n2016 vdd.n2015 185
R15908 vdd.n2015 vdd.n2014 185
R15909 vdd.n813 vdd.n812 185
R15910 vdd.n823 vdd.n813 185
R15911 vdd.n2006 vdd.n2005 185
R15912 vdd.n2007 vdd.n2006 185
R15913 vdd.n2004 vdd.n824 185
R15914 vdd.n824 vdd.n820 185
R15915 vdd.n2003 vdd.n2002 185
R15916 vdd.n2002 vdd.n2001 185
R15917 vdd.n826 vdd.n825 185
R15918 vdd.n827 vdd.n826 185
R15919 vdd.n1994 vdd.n1993 185
R15920 vdd.n1995 vdd.n1994 185
R15921 vdd.n1992 vdd.n836 185
R15922 vdd.n836 vdd.n833 185
R15923 vdd.n1991 vdd.n1990 185
R15924 vdd.n1990 vdd.n1989 185
R15925 vdd.n838 vdd.n837 185
R15926 vdd.n1726 vdd.n1725 185
R15927 vdd.n1727 vdd.n1723 185
R15928 vdd.n1723 vdd.n839 185
R15929 vdd.n1729 vdd.n1728 185
R15930 vdd.n1731 vdd.n1722 185
R15931 vdd.n1734 vdd.n1733 185
R15932 vdd.n1735 vdd.n1721 185
R15933 vdd.n1737 vdd.n1736 185
R15934 vdd.n1739 vdd.n1720 185
R15935 vdd.n1742 vdd.n1741 185
R15936 vdd.n1743 vdd.n1719 185
R15937 vdd.n1745 vdd.n1744 185
R15938 vdd.n1747 vdd.n1718 185
R15939 vdd.n1750 vdd.n1749 185
R15940 vdd.n1751 vdd.n1717 185
R15941 vdd.n1753 vdd.n1752 185
R15942 vdd.n1755 vdd.n1716 185
R15943 vdd.n1928 vdd.n1756 185
R15944 vdd.n1927 vdd.n1926 185
R15945 vdd.n1924 vdd.n1757 185
R15946 vdd.n1922 vdd.n1921 185
R15947 vdd.n1920 vdd.n1758 185
R15948 vdd.n1919 vdd.n1918 185
R15949 vdd.n1916 vdd.n1759 185
R15950 vdd.n1914 vdd.n1913 185
R15951 vdd.n1912 vdd.n1760 185
R15952 vdd.n1911 vdd.n1910 185
R15953 vdd.n1908 vdd.n1761 185
R15954 vdd.n1906 vdd.n1905 185
R15955 vdd.n1904 vdd.n1762 185
R15956 vdd.n1903 vdd.n1902 185
R15957 vdd.n1900 vdd.n1763 185
R15958 vdd.n1898 vdd.n1897 185
R15959 vdd.n1896 vdd.n1764 185
R15960 vdd.n1895 vdd.n1894 185
R15961 vdd.n2149 vdd.n2148 185
R15962 vdd.n2151 vdd.n2150 185
R15963 vdd.n2153 vdd.n2152 185
R15964 vdd.n2156 vdd.n2155 185
R15965 vdd.n2158 vdd.n2157 185
R15966 vdd.n2160 vdd.n2159 185
R15967 vdd.n2162 vdd.n2161 185
R15968 vdd.n2164 vdd.n2163 185
R15969 vdd.n2166 vdd.n2165 185
R15970 vdd.n2168 vdd.n2167 185
R15971 vdd.n2170 vdd.n2169 185
R15972 vdd.n2172 vdd.n2171 185
R15973 vdd.n2174 vdd.n2173 185
R15974 vdd.n2176 vdd.n2175 185
R15975 vdd.n2178 vdd.n2177 185
R15976 vdd.n2180 vdd.n2179 185
R15977 vdd.n2182 vdd.n2181 185
R15978 vdd.n2184 vdd.n2183 185
R15979 vdd.n2186 vdd.n2185 185
R15980 vdd.n2188 vdd.n2187 185
R15981 vdd.n2190 vdd.n2189 185
R15982 vdd.n2192 vdd.n2191 185
R15983 vdd.n2194 vdd.n2193 185
R15984 vdd.n2196 vdd.n2195 185
R15985 vdd.n2198 vdd.n2197 185
R15986 vdd.n2200 vdd.n2199 185
R15987 vdd.n2202 vdd.n2201 185
R15988 vdd.n2204 vdd.n2203 185
R15989 vdd.n2206 vdd.n2205 185
R15990 vdd.n2208 vdd.n2207 185
R15991 vdd.n2210 vdd.n2209 185
R15992 vdd.n2212 vdd.n2211 185
R15993 vdd.n2214 vdd.n2213 185
R15994 vdd.n2215 vdd.n745 185
R15995 vdd.n2217 vdd.n2216 185
R15996 vdd.n2218 vdd.n2217 185
R15997 vdd.n2147 vdd.n749 185
R15998 vdd.n2147 vdd.n2146 185
R15999 vdd.n1768 vdd.n750 185
R16000 vdd.t2 vdd.n750 185
R16001 vdd.n1769 vdd.n760 185
R16002 vdd.n2071 vdd.n760 185
R16003 vdd.n1772 vdd.n1771 185
R16004 vdd.n1771 vdd.n1770 185
R16005 vdd.n1773 vdd.n767 185
R16006 vdd.n2064 vdd.n767 185
R16007 vdd.n1775 vdd.n1774 185
R16008 vdd.n1774 vdd.n766 185
R16009 vdd.n1776 vdd.n774 185
R16010 vdd.n2056 vdd.n774 185
R16011 vdd.n1778 vdd.n1777 185
R16012 vdd.n1777 vdd.n773 185
R16013 vdd.n1779 vdd.n780 185
R16014 vdd.n2050 vdd.n780 185
R16015 vdd.n1781 vdd.n1780 185
R16016 vdd.n1780 vdd.n779 185
R16017 vdd.n1782 vdd.n785 185
R16018 vdd.n2044 vdd.n785 185
R16019 vdd.n1784 vdd.n1783 185
R16020 vdd.n1783 vdd.n792 185
R16021 vdd.n1785 vdd.n790 185
R16022 vdd.n2038 vdd.n790 185
R16023 vdd.n1787 vdd.n1786 185
R16024 vdd.n1786 vdd.n798 185
R16025 vdd.n1788 vdd.n796 185
R16026 vdd.n2032 vdd.n796 185
R16027 vdd.n1873 vdd.n1872 185
R16028 vdd.n1872 vdd.n1871 185
R16029 vdd.n1874 vdd.n803 185
R16030 vdd.n2026 vdd.n803 185
R16031 vdd.n1876 vdd.n1875 185
R16032 vdd.n1875 vdd.n802 185
R16033 vdd.n1877 vdd.n809 185
R16034 vdd.n2020 vdd.n809 185
R16035 vdd.n1879 vdd.n1878 185
R16036 vdd.n1878 vdd.n808 185
R16037 vdd.n1880 vdd.n814 185
R16038 vdd.n2014 vdd.n814 185
R16039 vdd.n1882 vdd.n1881 185
R16040 vdd.n1881 vdd.n823 185
R16041 vdd.n1883 vdd.n821 185
R16042 vdd.n2007 vdd.n821 185
R16043 vdd.n1885 vdd.n1884 185
R16044 vdd.n1884 vdd.n820 185
R16045 vdd.n1886 vdd.n828 185
R16046 vdd.n2001 vdd.n828 185
R16047 vdd.n1888 vdd.n1887 185
R16048 vdd.n1887 vdd.n827 185
R16049 vdd.n1889 vdd.n834 185
R16050 vdd.n1995 vdd.n834 185
R16051 vdd.n1891 vdd.n1890 185
R16052 vdd.n1890 vdd.n833 185
R16053 vdd.n1892 vdd.n840 185
R16054 vdd.n1989 vdd.n840 185
R16055 vdd.n3024 vdd.n3023 185
R16056 vdd.n3025 vdd.n3024 185
R16057 vdd.n325 vdd.n324 185
R16058 vdd.n3026 vdd.n325 185
R16059 vdd.n3029 vdd.n3028 185
R16060 vdd.n3028 vdd.n3027 185
R16061 vdd.n3030 vdd.n319 185
R16062 vdd.n319 vdd.n318 185
R16063 vdd.n3032 vdd.n3031 185
R16064 vdd.n3033 vdd.n3032 185
R16065 vdd.n314 vdd.n313 185
R16066 vdd.n3034 vdd.n314 185
R16067 vdd.n3037 vdd.n3036 185
R16068 vdd.n3036 vdd.n3035 185
R16069 vdd.n3038 vdd.n309 185
R16070 vdd.n309 vdd.n308 185
R16071 vdd.n3040 vdd.n3039 185
R16072 vdd.n3041 vdd.n3040 185
R16073 vdd.n303 vdd.n301 185
R16074 vdd.n3042 vdd.n303 185
R16075 vdd.n3045 vdd.n3044 185
R16076 vdd.n3044 vdd.n3043 185
R16077 vdd.n302 vdd.n300 185
R16078 vdd.n304 vdd.n302 185
R16079 vdd.n2881 vdd.n2880 185
R16080 vdd.n2882 vdd.n2881 185
R16081 vdd.n458 vdd.n457 185
R16082 vdd.n457 vdd.n456 185
R16083 vdd.n2876 vdd.n2875 185
R16084 vdd.n2875 vdd.n2874 185
R16085 vdd.n461 vdd.n460 185
R16086 vdd.n467 vdd.n461 185
R16087 vdd.n2865 vdd.n2864 185
R16088 vdd.n2866 vdd.n2865 185
R16089 vdd.n469 vdd.n468 185
R16090 vdd.n2857 vdd.n468 185
R16091 vdd.n2860 vdd.n2859 185
R16092 vdd.n2859 vdd.n2858 185
R16093 vdd.n472 vdd.n471 185
R16094 vdd.n473 vdd.n472 185
R16095 vdd.n2848 vdd.n2847 185
R16096 vdd.n2849 vdd.n2848 185
R16097 vdd.n480 vdd.n479 185
R16098 vdd.n516 vdd.n479 185
R16099 vdd.n2843 vdd.n2842 185
R16100 vdd.n483 vdd.n482 185
R16101 vdd.n2839 vdd.n2838 185
R16102 vdd.n2840 vdd.n2839 185
R16103 vdd.n518 vdd.n517 185
R16104 vdd.n522 vdd.n521 185
R16105 vdd.n2834 vdd.n523 185
R16106 vdd.n2833 vdd.n2832 185
R16107 vdd.n2831 vdd.n2830 185
R16108 vdd.n2829 vdd.n2828 185
R16109 vdd.n2827 vdd.n2826 185
R16110 vdd.n2825 vdd.n2824 185
R16111 vdd.n2823 vdd.n2822 185
R16112 vdd.n2821 vdd.n2820 185
R16113 vdd.n2819 vdd.n2818 185
R16114 vdd.n2817 vdd.n2816 185
R16115 vdd.n2815 vdd.n2814 185
R16116 vdd.n2813 vdd.n2812 185
R16117 vdd.n2811 vdd.n2810 185
R16118 vdd.n2809 vdd.n2808 185
R16119 vdd.n2807 vdd.n2806 185
R16120 vdd.n2798 vdd.n536 185
R16121 vdd.n2800 vdd.n2799 185
R16122 vdd.n2797 vdd.n2796 185
R16123 vdd.n2795 vdd.n2794 185
R16124 vdd.n2793 vdd.n2792 185
R16125 vdd.n2791 vdd.n2790 185
R16126 vdd.n2789 vdd.n2788 185
R16127 vdd.n2787 vdd.n2786 185
R16128 vdd.n2785 vdd.n2784 185
R16129 vdd.n2783 vdd.n2782 185
R16130 vdd.n2781 vdd.n2780 185
R16131 vdd.n2779 vdd.n2778 185
R16132 vdd.n2777 vdd.n2776 185
R16133 vdd.n2775 vdd.n2774 185
R16134 vdd.n2773 vdd.n2772 185
R16135 vdd.n2771 vdd.n2770 185
R16136 vdd.n2769 vdd.n2768 185
R16137 vdd.n2767 vdd.n2766 185
R16138 vdd.n2765 vdd.n2764 185
R16139 vdd.n2763 vdd.n2762 185
R16140 vdd.n2761 vdd.n2760 185
R16141 vdd.n2759 vdd.n2758 185
R16142 vdd.n2752 vdd.n556 185
R16143 vdd.n2754 vdd.n2753 185
R16144 vdd.n2751 vdd.n2750 185
R16145 vdd.n2749 vdd.n2748 185
R16146 vdd.n2747 vdd.n2746 185
R16147 vdd.n2745 vdd.n2744 185
R16148 vdd.n2743 vdd.n2742 185
R16149 vdd.n2741 vdd.n2740 185
R16150 vdd.n2739 vdd.n2738 185
R16151 vdd.n2737 vdd.n2736 185
R16152 vdd.n2735 vdd.n2734 185
R16153 vdd.n2733 vdd.n2732 185
R16154 vdd.n2731 vdd.n2730 185
R16155 vdd.n2729 vdd.n2728 185
R16156 vdd.n2727 vdd.n2726 185
R16157 vdd.n2725 vdd.n2724 185
R16158 vdd.n2723 vdd.n2722 185
R16159 vdd.n2721 vdd.n2720 185
R16160 vdd.n2719 vdd.n2718 185
R16161 vdd.n2717 vdd.n2716 185
R16162 vdd.n2715 vdd.n2714 185
R16163 vdd.n2710 vdd.n515 185
R16164 vdd.n2840 vdd.n515 185
R16165 vdd.n2907 vdd.n2906 185
R16166 vdd.n2911 vdd.n440 185
R16167 vdd.n2913 vdd.n2912 185
R16168 vdd.n2915 vdd.n438 185
R16169 vdd.n2917 vdd.n2916 185
R16170 vdd.n2918 vdd.n433 185
R16171 vdd.n2920 vdd.n2919 185
R16172 vdd.n2922 vdd.n431 185
R16173 vdd.n2924 vdd.n2923 185
R16174 vdd.n2925 vdd.n426 185
R16175 vdd.n2927 vdd.n2926 185
R16176 vdd.n2929 vdd.n424 185
R16177 vdd.n2931 vdd.n2930 185
R16178 vdd.n2932 vdd.n419 185
R16179 vdd.n2934 vdd.n2933 185
R16180 vdd.n2936 vdd.n417 185
R16181 vdd.n2938 vdd.n2937 185
R16182 vdd.n2939 vdd.n413 185
R16183 vdd.n2941 vdd.n2940 185
R16184 vdd.n2943 vdd.n410 185
R16185 vdd.n2945 vdd.n2944 185
R16186 vdd.n411 vdd.n404 185
R16187 vdd.n2949 vdd.n408 185
R16188 vdd.n2950 vdd.n400 185
R16189 vdd.n2952 vdd.n2951 185
R16190 vdd.n2954 vdd.n398 185
R16191 vdd.n2956 vdd.n2955 185
R16192 vdd.n2957 vdd.n393 185
R16193 vdd.n2959 vdd.n2958 185
R16194 vdd.n2961 vdd.n391 185
R16195 vdd.n2963 vdd.n2962 185
R16196 vdd.n2964 vdd.n386 185
R16197 vdd.n2966 vdd.n2965 185
R16198 vdd.n2968 vdd.n384 185
R16199 vdd.n2970 vdd.n2969 185
R16200 vdd.n2971 vdd.n379 185
R16201 vdd.n2973 vdd.n2972 185
R16202 vdd.n2975 vdd.n377 185
R16203 vdd.n2977 vdd.n2976 185
R16204 vdd.n2978 vdd.n373 185
R16205 vdd.n2980 vdd.n2979 185
R16206 vdd.n2982 vdd.n370 185
R16207 vdd.n2984 vdd.n2983 185
R16208 vdd.n371 vdd.n364 185
R16209 vdd.n2988 vdd.n368 185
R16210 vdd.n2989 vdd.n360 185
R16211 vdd.n2991 vdd.n2990 185
R16212 vdd.n2993 vdd.n358 185
R16213 vdd.n2995 vdd.n2994 185
R16214 vdd.n2996 vdd.n353 185
R16215 vdd.n2998 vdd.n2997 185
R16216 vdd.n3000 vdd.n351 185
R16217 vdd.n3002 vdd.n3001 185
R16218 vdd.n3003 vdd.n346 185
R16219 vdd.n3005 vdd.n3004 185
R16220 vdd.n3007 vdd.n344 185
R16221 vdd.n3009 vdd.n3008 185
R16222 vdd.n3010 vdd.n338 185
R16223 vdd.n3012 vdd.n3011 185
R16224 vdd.n3014 vdd.n337 185
R16225 vdd.n3015 vdd.n336 185
R16226 vdd.n3018 vdd.n3017 185
R16227 vdd.n3019 vdd.n334 185
R16228 vdd.n3020 vdd.n330 185
R16229 vdd.n2902 vdd.n328 185
R16230 vdd.n3025 vdd.n328 185
R16231 vdd.n2901 vdd.n327 185
R16232 vdd.n3026 vdd.n327 185
R16233 vdd.n2900 vdd.n326 185
R16234 vdd.n3027 vdd.n326 185
R16235 vdd.n446 vdd.n445 185
R16236 vdd.n445 vdd.n318 185
R16237 vdd.n2896 vdd.n317 185
R16238 vdd.n3033 vdd.n317 185
R16239 vdd.n2895 vdd.n316 185
R16240 vdd.n3034 vdd.n316 185
R16241 vdd.n2894 vdd.n315 185
R16242 vdd.n3035 vdd.n315 185
R16243 vdd.n449 vdd.n448 185
R16244 vdd.n448 vdd.n308 185
R16245 vdd.n2890 vdd.n307 185
R16246 vdd.n3041 vdd.n307 185
R16247 vdd.n2889 vdd.n306 185
R16248 vdd.n3042 vdd.n306 185
R16249 vdd.n2888 vdd.n305 185
R16250 vdd.n3043 vdd.n305 185
R16251 vdd.n455 vdd.n451 185
R16252 vdd.n455 vdd.n304 185
R16253 vdd.n2884 vdd.n2883 185
R16254 vdd.n2883 vdd.n2882 185
R16255 vdd.n454 vdd.n453 185
R16256 vdd.n456 vdd.n454 185
R16257 vdd.n2873 vdd.n2872 185
R16258 vdd.n2874 vdd.n2873 185
R16259 vdd.n463 vdd.n462 185
R16260 vdd.n467 vdd.n462 185
R16261 vdd.n2868 vdd.n2867 185
R16262 vdd.n2867 vdd.n2866 185
R16263 vdd.n466 vdd.n465 185
R16264 vdd.n2857 vdd.n466 185
R16265 vdd.n2856 vdd.n2855 185
R16266 vdd.n2858 vdd.n2856 185
R16267 vdd.n475 vdd.n474 185
R16268 vdd.n474 vdd.n473 185
R16269 vdd.n2851 vdd.n2850 185
R16270 vdd.n2850 vdd.n2849 185
R16271 vdd.n478 vdd.n477 185
R16272 vdd.n516 vdd.n478 185
R16273 vdd.n703 vdd.n702 185
R16274 vdd.n2469 vdd.n2468 185
R16275 vdd.n2467 vdd.n2252 185
R16276 vdd.n2471 vdd.n2252 185
R16277 vdd.n2466 vdd.n2465 185
R16278 vdd.n2464 vdd.n2463 185
R16279 vdd.n2462 vdd.n2461 185
R16280 vdd.n2460 vdd.n2459 185
R16281 vdd.n2458 vdd.n2457 185
R16282 vdd.n2456 vdd.n2455 185
R16283 vdd.n2454 vdd.n2453 185
R16284 vdd.n2452 vdd.n2451 185
R16285 vdd.n2450 vdd.n2449 185
R16286 vdd.n2448 vdd.n2447 185
R16287 vdd.n2446 vdd.n2445 185
R16288 vdd.n2444 vdd.n2443 185
R16289 vdd.n2442 vdd.n2441 185
R16290 vdd.n2440 vdd.n2439 185
R16291 vdd.n2438 vdd.n2437 185
R16292 vdd.n2436 vdd.n2435 185
R16293 vdd.n2434 vdd.n2433 185
R16294 vdd.n2432 vdd.n2431 185
R16295 vdd.n2430 vdd.n2429 185
R16296 vdd.n2428 vdd.n2427 185
R16297 vdd.n2426 vdd.n2425 185
R16298 vdd.n2424 vdd.n2423 185
R16299 vdd.n2422 vdd.n2421 185
R16300 vdd.n2420 vdd.n2419 185
R16301 vdd.n2418 vdd.n2417 185
R16302 vdd.n2416 vdd.n2415 185
R16303 vdd.n2414 vdd.n2413 185
R16304 vdd.n2412 vdd.n2411 185
R16305 vdd.n2410 vdd.n2409 185
R16306 vdd.n2407 vdd.n2406 185
R16307 vdd.n2405 vdd.n2404 185
R16308 vdd.n2403 vdd.n2402 185
R16309 vdd.n2609 vdd.n2608 185
R16310 vdd.n2611 vdd.n624 185
R16311 vdd.n2613 vdd.n2612 185
R16312 vdd.n2615 vdd.n621 185
R16313 vdd.n2617 vdd.n2616 185
R16314 vdd.n2619 vdd.n619 185
R16315 vdd.n2621 vdd.n2620 185
R16316 vdd.n2622 vdd.n618 185
R16317 vdd.n2624 vdd.n2623 185
R16318 vdd.n2626 vdd.n616 185
R16319 vdd.n2628 vdd.n2627 185
R16320 vdd.n2629 vdd.n615 185
R16321 vdd.n2631 vdd.n2630 185
R16322 vdd.n2633 vdd.n613 185
R16323 vdd.n2635 vdd.n2634 185
R16324 vdd.n2636 vdd.n612 185
R16325 vdd.n2638 vdd.n2637 185
R16326 vdd.n2640 vdd.n520 185
R16327 vdd.n2642 vdd.n2641 185
R16328 vdd.n2644 vdd.n610 185
R16329 vdd.n2646 vdd.n2645 185
R16330 vdd.n2647 vdd.n609 185
R16331 vdd.n2649 vdd.n2648 185
R16332 vdd.n2651 vdd.n607 185
R16333 vdd.n2653 vdd.n2652 185
R16334 vdd.n2654 vdd.n606 185
R16335 vdd.n2656 vdd.n2655 185
R16336 vdd.n2658 vdd.n604 185
R16337 vdd.n2660 vdd.n2659 185
R16338 vdd.n2661 vdd.n603 185
R16339 vdd.n2663 vdd.n2662 185
R16340 vdd.n2665 vdd.n602 185
R16341 vdd.n2666 vdd.n601 185
R16342 vdd.n2669 vdd.n2668 185
R16343 vdd.n2670 vdd.n599 185
R16344 vdd.n599 vdd.n484 185
R16345 vdd.n2607 vdd.n596 185
R16346 vdd.n2673 vdd.n596 185
R16347 vdd.n2606 vdd.n2605 185
R16348 vdd.n2605 vdd.n595 185
R16349 vdd.n2604 vdd.n626 185
R16350 vdd.n2604 vdd.n2603 185
R16351 vdd.n2358 vdd.n627 185
R16352 vdd.n636 vdd.n627 185
R16353 vdd.n2359 vdd.n634 185
R16354 vdd.n2597 vdd.n634 185
R16355 vdd.n2361 vdd.n2360 185
R16356 vdd.n2360 vdd.n633 185
R16357 vdd.n2362 vdd.n642 185
R16358 vdd.n2546 vdd.n642 185
R16359 vdd.n2364 vdd.n2363 185
R16360 vdd.n2363 vdd.n641 185
R16361 vdd.n2365 vdd.n648 185
R16362 vdd.n2540 vdd.n648 185
R16363 vdd.n2367 vdd.n2366 185
R16364 vdd.n2366 vdd.n647 185
R16365 vdd.n2368 vdd.n653 185
R16366 vdd.n2532 vdd.n653 185
R16367 vdd.n2370 vdd.n2369 185
R16368 vdd.n2369 vdd.n660 185
R16369 vdd.n2371 vdd.n658 185
R16370 vdd.n2526 vdd.n658 185
R16371 vdd.n2373 vdd.n2372 185
R16372 vdd.n2374 vdd.n2373 185
R16373 vdd.n2357 vdd.n665 185
R16374 vdd.n2520 vdd.n665 185
R16375 vdd.n2356 vdd.n2355 185
R16376 vdd.n2355 vdd.n664 185
R16377 vdd.n2354 vdd.n671 185
R16378 vdd.n2514 vdd.n671 185
R16379 vdd.n2353 vdd.n2352 185
R16380 vdd.n2352 vdd.n670 185
R16381 vdd.n2351 vdd.n676 185
R16382 vdd.n2508 vdd.n676 185
R16383 vdd.n2350 vdd.n2349 185
R16384 vdd.n2349 vdd.n683 185
R16385 vdd.n2348 vdd.n681 185
R16386 vdd.n2502 vdd.n681 185
R16387 vdd.n2347 vdd.n2346 185
R16388 vdd.n2346 vdd.n690 185
R16389 vdd.n2345 vdd.n688 185
R16390 vdd.n2496 vdd.n688 185
R16391 vdd.n2344 vdd.n2343 185
R16392 vdd.n2343 vdd.n687 185
R16393 vdd.n2255 vdd.n694 185
R16394 vdd.n2490 vdd.n694 185
R16395 vdd.n2397 vdd.n2396 185
R16396 vdd.n2396 vdd.n2395 185
R16397 vdd.n2398 vdd.n699 185
R16398 vdd.n2484 vdd.n699 185
R16399 vdd.n2400 vdd.n2399 185
R16400 vdd.n2399 vdd.t198 185
R16401 vdd.n2401 vdd.n704 185
R16402 vdd.n2478 vdd.n704 185
R16403 vdd.n2480 vdd.n2479 185
R16404 vdd.n2479 vdd.n2478 185
R16405 vdd.n2481 vdd.n701 185
R16406 vdd.n701 vdd.t198 185
R16407 vdd.n2483 vdd.n2482 185
R16408 vdd.n2484 vdd.n2483 185
R16409 vdd.n693 vdd.n692 185
R16410 vdd.n2395 vdd.n693 185
R16411 vdd.n2492 vdd.n2491 185
R16412 vdd.n2491 vdd.n2490 185
R16413 vdd.n2493 vdd.n691 185
R16414 vdd.n691 vdd.n687 185
R16415 vdd.n2495 vdd.n2494 185
R16416 vdd.n2496 vdd.n2495 185
R16417 vdd.n680 vdd.n679 185
R16418 vdd.n690 vdd.n680 185
R16419 vdd.n2504 vdd.n2503 185
R16420 vdd.n2503 vdd.n2502 185
R16421 vdd.n2505 vdd.n678 185
R16422 vdd.n683 vdd.n678 185
R16423 vdd.n2507 vdd.n2506 185
R16424 vdd.n2508 vdd.n2507 185
R16425 vdd.n669 vdd.n668 185
R16426 vdd.n670 vdd.n669 185
R16427 vdd.n2516 vdd.n2515 185
R16428 vdd.n2515 vdd.n2514 185
R16429 vdd.n2517 vdd.n667 185
R16430 vdd.n667 vdd.n664 185
R16431 vdd.n2519 vdd.n2518 185
R16432 vdd.n2520 vdd.n2519 185
R16433 vdd.n657 vdd.n656 185
R16434 vdd.n2374 vdd.n657 185
R16435 vdd.n2528 vdd.n2527 185
R16436 vdd.n2527 vdd.n2526 185
R16437 vdd.n2529 vdd.n655 185
R16438 vdd.n660 vdd.n655 185
R16439 vdd.n2531 vdd.n2530 185
R16440 vdd.n2532 vdd.n2531 185
R16441 vdd.n646 vdd.n645 185
R16442 vdd.n647 vdd.n646 185
R16443 vdd.n2542 vdd.n2541 185
R16444 vdd.n2541 vdd.n2540 185
R16445 vdd.n2543 vdd.n644 185
R16446 vdd.n644 vdd.n641 185
R16447 vdd.n2545 vdd.n2544 185
R16448 vdd.n2546 vdd.n2545 185
R16449 vdd.n632 vdd.n631 185
R16450 vdd.n633 vdd.n632 185
R16451 vdd.n2599 vdd.n2598 185
R16452 vdd.n2598 vdd.n2597 185
R16453 vdd.n2600 vdd.n630 185
R16454 vdd.n636 vdd.n630 185
R16455 vdd.n2602 vdd.n2601 185
R16456 vdd.n2603 vdd.n2602 185
R16457 vdd.n600 vdd.n598 185
R16458 vdd.n598 vdd.n595 185
R16459 vdd.n2672 vdd.n2671 185
R16460 vdd.n2673 vdd.n2672 185
R16461 vdd.n2145 vdd.n2144 185
R16462 vdd.n2146 vdd.n2145 185
R16463 vdd.n754 vdd.n752 185
R16464 vdd.n752 vdd.t2 185
R16465 vdd.n2060 vdd.n761 185
R16466 vdd.n2071 vdd.n761 185
R16467 vdd.n2061 vdd.n770 185
R16468 vdd.n1770 vdd.n770 185
R16469 vdd.n2063 vdd.n2062 185
R16470 vdd.n2064 vdd.n2063 185
R16471 vdd.n2059 vdd.n769 185
R16472 vdd.n769 vdd.n766 185
R16473 vdd.n2058 vdd.n2057 185
R16474 vdd.n2057 vdd.n2056 185
R16475 vdd.n772 vdd.n771 185
R16476 vdd.n773 vdd.n772 185
R16477 vdd.n2049 vdd.n2048 185
R16478 vdd.n2050 vdd.n2049 185
R16479 vdd.n2047 vdd.n782 185
R16480 vdd.n782 vdd.n779 185
R16481 vdd.n2046 vdd.n2045 185
R16482 vdd.n2045 vdd.n2044 185
R16483 vdd.n784 vdd.n783 185
R16484 vdd.n792 vdd.n784 185
R16485 vdd.n2037 vdd.n2036 185
R16486 vdd.n2038 vdd.n2037 185
R16487 vdd.n2035 vdd.n793 185
R16488 vdd.n798 vdd.n793 185
R16489 vdd.n2034 vdd.n2033 185
R16490 vdd.n2033 vdd.n2032 185
R16491 vdd.n795 vdd.n794 185
R16492 vdd.n1871 vdd.n795 185
R16493 vdd.n2025 vdd.n2024 185
R16494 vdd.n2026 vdd.n2025 185
R16495 vdd.n2023 vdd.n805 185
R16496 vdd.n805 vdd.n802 185
R16497 vdd.n2022 vdd.n2021 185
R16498 vdd.n2021 vdd.n2020 185
R16499 vdd.n807 vdd.n806 185
R16500 vdd.n808 vdd.n807 185
R16501 vdd.n2013 vdd.n2012 185
R16502 vdd.n2014 vdd.n2013 185
R16503 vdd.n2010 vdd.n816 185
R16504 vdd.n823 vdd.n816 185
R16505 vdd.n2009 vdd.n2008 185
R16506 vdd.n2008 vdd.n2007 185
R16507 vdd.n819 vdd.n818 185
R16508 vdd.n820 vdd.n819 185
R16509 vdd.n2000 vdd.n1999 185
R16510 vdd.n2001 vdd.n2000 185
R16511 vdd.n1998 vdd.n830 185
R16512 vdd.n830 vdd.n827 185
R16513 vdd.n1997 vdd.n1996 185
R16514 vdd.n1996 vdd.n1995 185
R16515 vdd.n832 vdd.n831 185
R16516 vdd.n833 vdd.n832 185
R16517 vdd.n1988 vdd.n1987 185
R16518 vdd.n1989 vdd.n1988 185
R16519 vdd.n2076 vdd.n726 185
R16520 vdd.n2218 vdd.n726 185
R16521 vdd.n2078 vdd.n2077 185
R16522 vdd.n2080 vdd.n2079 185
R16523 vdd.n2082 vdd.n2081 185
R16524 vdd.n2084 vdd.n2083 185
R16525 vdd.n2086 vdd.n2085 185
R16526 vdd.n2088 vdd.n2087 185
R16527 vdd.n2090 vdd.n2089 185
R16528 vdd.n2092 vdd.n2091 185
R16529 vdd.n2094 vdd.n2093 185
R16530 vdd.n2096 vdd.n2095 185
R16531 vdd.n2098 vdd.n2097 185
R16532 vdd.n2100 vdd.n2099 185
R16533 vdd.n2102 vdd.n2101 185
R16534 vdd.n2104 vdd.n2103 185
R16535 vdd.n2106 vdd.n2105 185
R16536 vdd.n2108 vdd.n2107 185
R16537 vdd.n2110 vdd.n2109 185
R16538 vdd.n2112 vdd.n2111 185
R16539 vdd.n2114 vdd.n2113 185
R16540 vdd.n2116 vdd.n2115 185
R16541 vdd.n2118 vdd.n2117 185
R16542 vdd.n2120 vdd.n2119 185
R16543 vdd.n2122 vdd.n2121 185
R16544 vdd.n2124 vdd.n2123 185
R16545 vdd.n2126 vdd.n2125 185
R16546 vdd.n2128 vdd.n2127 185
R16547 vdd.n2130 vdd.n2129 185
R16548 vdd.n2132 vdd.n2131 185
R16549 vdd.n2134 vdd.n2133 185
R16550 vdd.n2136 vdd.n2135 185
R16551 vdd.n2138 vdd.n2137 185
R16552 vdd.n2140 vdd.n2139 185
R16553 vdd.n2142 vdd.n2141 185
R16554 vdd.n2143 vdd.n753 185
R16555 vdd.n2075 vdd.n751 185
R16556 vdd.n2146 vdd.n751 185
R16557 vdd.n2074 vdd.n2073 185
R16558 vdd.n2073 vdd.t2 185
R16559 vdd.n2072 vdd.n758 185
R16560 vdd.n2072 vdd.n2071 185
R16561 vdd.n1852 vdd.n759 185
R16562 vdd.n1770 vdd.n759 185
R16563 vdd.n1853 vdd.n768 185
R16564 vdd.n2064 vdd.n768 185
R16565 vdd.n1855 vdd.n1854 185
R16566 vdd.n1854 vdd.n766 185
R16567 vdd.n1856 vdd.n775 185
R16568 vdd.n2056 vdd.n775 185
R16569 vdd.n1858 vdd.n1857 185
R16570 vdd.n1857 vdd.n773 185
R16571 vdd.n1859 vdd.n781 185
R16572 vdd.n2050 vdd.n781 185
R16573 vdd.n1861 vdd.n1860 185
R16574 vdd.n1860 vdd.n779 185
R16575 vdd.n1862 vdd.n786 185
R16576 vdd.n2044 vdd.n786 185
R16577 vdd.n1864 vdd.n1863 185
R16578 vdd.n1863 vdd.n792 185
R16579 vdd.n1865 vdd.n791 185
R16580 vdd.n2038 vdd.n791 185
R16581 vdd.n1867 vdd.n1866 185
R16582 vdd.n1866 vdd.n798 185
R16583 vdd.n1868 vdd.n797 185
R16584 vdd.n2032 vdd.n797 185
R16585 vdd.n1870 vdd.n1869 185
R16586 vdd.n1871 vdd.n1870 185
R16587 vdd.n1851 vdd.n804 185
R16588 vdd.n2026 vdd.n804 185
R16589 vdd.n1850 vdd.n1849 185
R16590 vdd.n1849 vdd.n802 185
R16591 vdd.n1848 vdd.n810 185
R16592 vdd.n2020 vdd.n810 185
R16593 vdd.n1847 vdd.n1846 185
R16594 vdd.n1846 vdd.n808 185
R16595 vdd.n1845 vdd.n815 185
R16596 vdd.n2014 vdd.n815 185
R16597 vdd.n1844 vdd.n1843 185
R16598 vdd.n1843 vdd.n823 185
R16599 vdd.n1842 vdd.n822 185
R16600 vdd.n2007 vdd.n822 185
R16601 vdd.n1841 vdd.n1840 185
R16602 vdd.n1840 vdd.n820 185
R16603 vdd.n1839 vdd.n829 185
R16604 vdd.n2001 vdd.n829 185
R16605 vdd.n1838 vdd.n1837 185
R16606 vdd.n1837 vdd.n827 185
R16607 vdd.n1836 vdd.n835 185
R16608 vdd.n1995 vdd.n835 185
R16609 vdd.n1835 vdd.n1834 185
R16610 vdd.n1834 vdd.n833 185
R16611 vdd.n1833 vdd.n841 185
R16612 vdd.n1989 vdd.n841 185
R16613 vdd.n1986 vdd.n842 185
R16614 vdd.n1985 vdd.n1984 185
R16615 vdd.n1982 vdd.n843 185
R16616 vdd.n1980 vdd.n1979 185
R16617 vdd.n1978 vdd.n844 185
R16618 vdd.n1977 vdd.n1976 185
R16619 vdd.n1974 vdd.n845 185
R16620 vdd.n1972 vdd.n1971 185
R16621 vdd.n1970 vdd.n846 185
R16622 vdd.n1969 vdd.n1968 185
R16623 vdd.n1966 vdd.n847 185
R16624 vdd.n1964 vdd.n1963 185
R16625 vdd.n1962 vdd.n848 185
R16626 vdd.n1961 vdd.n1960 185
R16627 vdd.n1958 vdd.n849 185
R16628 vdd.n1956 vdd.n1955 185
R16629 vdd.n1954 vdd.n850 185
R16630 vdd.n1953 vdd.n852 185
R16631 vdd.n1798 vdd.n853 185
R16632 vdd.n1801 vdd.n1800 185
R16633 vdd.n1803 vdd.n1802 185
R16634 vdd.n1805 vdd.n1797 185
R16635 vdd.n1808 vdd.n1807 185
R16636 vdd.n1809 vdd.n1796 185
R16637 vdd.n1811 vdd.n1810 185
R16638 vdd.n1813 vdd.n1795 185
R16639 vdd.n1816 vdd.n1815 185
R16640 vdd.n1817 vdd.n1794 185
R16641 vdd.n1819 vdd.n1818 185
R16642 vdd.n1821 vdd.n1793 185
R16643 vdd.n1824 vdd.n1823 185
R16644 vdd.n1825 vdd.n1790 185
R16645 vdd.n1828 vdd.n1827 185
R16646 vdd.n1830 vdd.n1789 185
R16647 vdd.n1832 vdd.n1831 185
R16648 vdd.n1831 vdd.n839 185
R16649 vdd.n291 vdd.n290 171.744
R16650 vdd.n290 vdd.n289 171.744
R16651 vdd.n289 vdd.n258 171.744
R16652 vdd.n282 vdd.n258 171.744
R16653 vdd.n282 vdd.n281 171.744
R16654 vdd.n281 vdd.n263 171.744
R16655 vdd.n274 vdd.n263 171.744
R16656 vdd.n274 vdd.n273 171.744
R16657 vdd.n273 vdd.n267 171.744
R16658 vdd.n244 vdd.n243 171.744
R16659 vdd.n243 vdd.n242 171.744
R16660 vdd.n242 vdd.n211 171.744
R16661 vdd.n235 vdd.n211 171.744
R16662 vdd.n235 vdd.n234 171.744
R16663 vdd.n234 vdd.n216 171.744
R16664 vdd.n227 vdd.n216 171.744
R16665 vdd.n227 vdd.n226 171.744
R16666 vdd.n226 vdd.n220 171.744
R16667 vdd.n201 vdd.n200 171.744
R16668 vdd.n200 vdd.n199 171.744
R16669 vdd.n199 vdd.n168 171.744
R16670 vdd.n192 vdd.n168 171.744
R16671 vdd.n192 vdd.n191 171.744
R16672 vdd.n191 vdd.n173 171.744
R16673 vdd.n184 vdd.n173 171.744
R16674 vdd.n184 vdd.n183 171.744
R16675 vdd.n183 vdd.n177 171.744
R16676 vdd.n154 vdd.n153 171.744
R16677 vdd.n153 vdd.n152 171.744
R16678 vdd.n152 vdd.n121 171.744
R16679 vdd.n145 vdd.n121 171.744
R16680 vdd.n145 vdd.n144 171.744
R16681 vdd.n144 vdd.n126 171.744
R16682 vdd.n137 vdd.n126 171.744
R16683 vdd.n137 vdd.n136 171.744
R16684 vdd.n136 vdd.n130 171.744
R16685 vdd.n112 vdd.n111 171.744
R16686 vdd.n111 vdd.n110 171.744
R16687 vdd.n110 vdd.n79 171.744
R16688 vdd.n103 vdd.n79 171.744
R16689 vdd.n103 vdd.n102 171.744
R16690 vdd.n102 vdd.n84 171.744
R16691 vdd.n95 vdd.n84 171.744
R16692 vdd.n95 vdd.n94 171.744
R16693 vdd.n94 vdd.n88 171.744
R16694 vdd.n65 vdd.n64 171.744
R16695 vdd.n64 vdd.n63 171.744
R16696 vdd.n63 vdd.n32 171.744
R16697 vdd.n56 vdd.n32 171.744
R16698 vdd.n56 vdd.n55 171.744
R16699 vdd.n55 vdd.n37 171.744
R16700 vdd.n48 vdd.n37 171.744
R16701 vdd.n48 vdd.n47 171.744
R16702 vdd.n47 vdd.n41 171.744
R16703 vdd.n1106 vdd.n1105 171.744
R16704 vdd.n1105 vdd.n1104 171.744
R16705 vdd.n1104 vdd.n1073 171.744
R16706 vdd.n1097 vdd.n1073 171.744
R16707 vdd.n1097 vdd.n1096 171.744
R16708 vdd.n1096 vdd.n1078 171.744
R16709 vdd.n1089 vdd.n1078 171.744
R16710 vdd.n1089 vdd.n1088 171.744
R16711 vdd.n1088 vdd.n1082 171.744
R16712 vdd.n1153 vdd.n1152 171.744
R16713 vdd.n1152 vdd.n1151 171.744
R16714 vdd.n1151 vdd.n1120 171.744
R16715 vdd.n1144 vdd.n1120 171.744
R16716 vdd.n1144 vdd.n1143 171.744
R16717 vdd.n1143 vdd.n1125 171.744
R16718 vdd.n1136 vdd.n1125 171.744
R16719 vdd.n1136 vdd.n1135 171.744
R16720 vdd.n1135 vdd.n1129 171.744
R16721 vdd.n1016 vdd.n1015 171.744
R16722 vdd.n1015 vdd.n1014 171.744
R16723 vdd.n1014 vdd.n983 171.744
R16724 vdd.n1007 vdd.n983 171.744
R16725 vdd.n1007 vdd.n1006 171.744
R16726 vdd.n1006 vdd.n988 171.744
R16727 vdd.n999 vdd.n988 171.744
R16728 vdd.n999 vdd.n998 171.744
R16729 vdd.n998 vdd.n992 171.744
R16730 vdd.n1063 vdd.n1062 171.744
R16731 vdd.n1062 vdd.n1061 171.744
R16732 vdd.n1061 vdd.n1030 171.744
R16733 vdd.n1054 vdd.n1030 171.744
R16734 vdd.n1054 vdd.n1053 171.744
R16735 vdd.n1053 vdd.n1035 171.744
R16736 vdd.n1046 vdd.n1035 171.744
R16737 vdd.n1046 vdd.n1045 171.744
R16738 vdd.n1045 vdd.n1039 171.744
R16739 vdd.n927 vdd.n926 171.744
R16740 vdd.n926 vdd.n925 171.744
R16741 vdd.n925 vdd.n894 171.744
R16742 vdd.n918 vdd.n894 171.744
R16743 vdd.n918 vdd.n917 171.744
R16744 vdd.n917 vdd.n899 171.744
R16745 vdd.n910 vdd.n899 171.744
R16746 vdd.n910 vdd.n909 171.744
R16747 vdd.n909 vdd.n903 171.744
R16748 vdd.n974 vdd.n973 171.744
R16749 vdd.n973 vdd.n972 171.744
R16750 vdd.n972 vdd.n941 171.744
R16751 vdd.n965 vdd.n941 171.744
R16752 vdd.n965 vdd.n964 171.744
R16753 vdd.n964 vdd.n946 171.744
R16754 vdd.n957 vdd.n946 171.744
R16755 vdd.n957 vdd.n956 171.744
R16756 vdd.n956 vdd.n950 171.744
R16757 vdd.n3017 vdd.n334 146.341
R16758 vdd.n3015 vdd.n3014 146.341
R16759 vdd.n3012 vdd.n338 146.341
R16760 vdd.n3008 vdd.n3007 146.341
R16761 vdd.n3005 vdd.n346 146.341
R16762 vdd.n3001 vdd.n3000 146.341
R16763 vdd.n2998 vdd.n353 146.341
R16764 vdd.n2994 vdd.n2993 146.341
R16765 vdd.n2991 vdd.n360 146.341
R16766 vdd.n371 vdd.n368 146.341
R16767 vdd.n2983 vdd.n2982 146.341
R16768 vdd.n2980 vdd.n373 146.341
R16769 vdd.n2976 vdd.n2975 146.341
R16770 vdd.n2973 vdd.n379 146.341
R16771 vdd.n2969 vdd.n2968 146.341
R16772 vdd.n2966 vdd.n386 146.341
R16773 vdd.n2962 vdd.n2961 146.341
R16774 vdd.n2959 vdd.n393 146.341
R16775 vdd.n2955 vdd.n2954 146.341
R16776 vdd.n2952 vdd.n400 146.341
R16777 vdd.n411 vdd.n408 146.341
R16778 vdd.n2944 vdd.n2943 146.341
R16779 vdd.n2941 vdd.n413 146.341
R16780 vdd.n2937 vdd.n2936 146.341
R16781 vdd.n2934 vdd.n419 146.341
R16782 vdd.n2930 vdd.n2929 146.341
R16783 vdd.n2927 vdd.n426 146.341
R16784 vdd.n2923 vdd.n2922 146.341
R16785 vdd.n2920 vdd.n433 146.341
R16786 vdd.n2916 vdd.n2915 146.341
R16787 vdd.n2913 vdd.n440 146.341
R16788 vdd.n2850 vdd.n478 146.341
R16789 vdd.n2850 vdd.n474 146.341
R16790 vdd.n2856 vdd.n474 146.341
R16791 vdd.n2856 vdd.n466 146.341
R16792 vdd.n2867 vdd.n466 146.341
R16793 vdd.n2867 vdd.n462 146.341
R16794 vdd.n2873 vdd.n462 146.341
R16795 vdd.n2873 vdd.n454 146.341
R16796 vdd.n2883 vdd.n454 146.341
R16797 vdd.n2883 vdd.n455 146.341
R16798 vdd.n455 vdd.n305 146.341
R16799 vdd.n306 vdd.n305 146.341
R16800 vdd.n307 vdd.n306 146.341
R16801 vdd.n448 vdd.n307 146.341
R16802 vdd.n448 vdd.n315 146.341
R16803 vdd.n316 vdd.n315 146.341
R16804 vdd.n317 vdd.n316 146.341
R16805 vdd.n445 vdd.n317 146.341
R16806 vdd.n445 vdd.n326 146.341
R16807 vdd.n327 vdd.n326 146.341
R16808 vdd.n328 vdd.n327 146.341
R16809 vdd.n2839 vdd.n483 146.341
R16810 vdd.n2839 vdd.n517 146.341
R16811 vdd.n523 vdd.n522 146.341
R16812 vdd.n2832 vdd.n2831 146.341
R16813 vdd.n2828 vdd.n2827 146.341
R16814 vdd.n2824 vdd.n2823 146.341
R16815 vdd.n2820 vdd.n2819 146.341
R16816 vdd.n2816 vdd.n2815 146.341
R16817 vdd.n2812 vdd.n2811 146.341
R16818 vdd.n2808 vdd.n2807 146.341
R16819 vdd.n2799 vdd.n2798 146.341
R16820 vdd.n2796 vdd.n2795 146.341
R16821 vdd.n2792 vdd.n2791 146.341
R16822 vdd.n2788 vdd.n2787 146.341
R16823 vdd.n2784 vdd.n2783 146.341
R16824 vdd.n2780 vdd.n2779 146.341
R16825 vdd.n2776 vdd.n2775 146.341
R16826 vdd.n2772 vdd.n2771 146.341
R16827 vdd.n2768 vdd.n2767 146.341
R16828 vdd.n2764 vdd.n2763 146.341
R16829 vdd.n2760 vdd.n2759 146.341
R16830 vdd.n2753 vdd.n2752 146.341
R16831 vdd.n2750 vdd.n2749 146.341
R16832 vdd.n2746 vdd.n2745 146.341
R16833 vdd.n2742 vdd.n2741 146.341
R16834 vdd.n2738 vdd.n2737 146.341
R16835 vdd.n2734 vdd.n2733 146.341
R16836 vdd.n2730 vdd.n2729 146.341
R16837 vdd.n2726 vdd.n2725 146.341
R16838 vdd.n2722 vdd.n2721 146.341
R16839 vdd.n2718 vdd.n2717 146.341
R16840 vdd.n2714 vdd.n515 146.341
R16841 vdd.n2848 vdd.n479 146.341
R16842 vdd.n2848 vdd.n472 146.341
R16843 vdd.n2859 vdd.n472 146.341
R16844 vdd.n2859 vdd.n468 146.341
R16845 vdd.n2865 vdd.n468 146.341
R16846 vdd.n2865 vdd.n461 146.341
R16847 vdd.n2875 vdd.n461 146.341
R16848 vdd.n2875 vdd.n457 146.341
R16849 vdd.n2881 vdd.n457 146.341
R16850 vdd.n2881 vdd.n302 146.341
R16851 vdd.n3044 vdd.n302 146.341
R16852 vdd.n3044 vdd.n303 146.341
R16853 vdd.n3040 vdd.n303 146.341
R16854 vdd.n3040 vdd.n309 146.341
R16855 vdd.n3036 vdd.n309 146.341
R16856 vdd.n3036 vdd.n314 146.341
R16857 vdd.n3032 vdd.n314 146.341
R16858 vdd.n3032 vdd.n319 146.341
R16859 vdd.n3028 vdd.n319 146.341
R16860 vdd.n3028 vdd.n325 146.341
R16861 vdd.n3024 vdd.n325 146.341
R16862 vdd.n1936 vdd.n1935 146.341
R16863 vdd.n1933 vdd.n1517 146.341
R16864 vdd.n1713 vdd.n1523 146.341
R16865 vdd.n1711 vdd.n1710 146.341
R16866 vdd.n1708 vdd.n1525 146.341
R16867 vdd.n1704 vdd.n1703 146.341
R16868 vdd.n1701 vdd.n1532 146.341
R16869 vdd.n1697 vdd.n1696 146.341
R16870 vdd.n1694 vdd.n1539 146.341
R16871 vdd.n1550 vdd.n1547 146.341
R16872 vdd.n1686 vdd.n1685 146.341
R16873 vdd.n1683 vdd.n1552 146.341
R16874 vdd.n1679 vdd.n1678 146.341
R16875 vdd.n1676 vdd.n1558 146.341
R16876 vdd.n1672 vdd.n1671 146.341
R16877 vdd.n1669 vdd.n1565 146.341
R16878 vdd.n1665 vdd.n1664 146.341
R16879 vdd.n1662 vdd.n1572 146.341
R16880 vdd.n1658 vdd.n1657 146.341
R16881 vdd.n1655 vdd.n1579 146.341
R16882 vdd.n1590 vdd.n1587 146.341
R16883 vdd.n1647 vdd.n1646 146.341
R16884 vdd.n1644 vdd.n1592 146.341
R16885 vdd.n1640 vdd.n1639 146.341
R16886 vdd.n1637 vdd.n1598 146.341
R16887 vdd.n1633 vdd.n1632 146.341
R16888 vdd.n1630 vdd.n1605 146.341
R16889 vdd.n1626 vdd.n1625 146.341
R16890 vdd.n1623 vdd.n1620 146.341
R16891 vdd.n1618 vdd.n1615 146.341
R16892 vdd.n1613 vdd.n859 146.341
R16893 vdd.n1431 vdd.n1191 146.341
R16894 vdd.n1431 vdd.n1187 146.341
R16895 vdd.n1437 vdd.n1187 146.341
R16896 vdd.n1437 vdd.n1179 146.341
R16897 vdd.n1448 vdd.n1179 146.341
R16898 vdd.n1448 vdd.n1175 146.341
R16899 vdd.n1454 vdd.n1175 146.341
R16900 vdd.n1454 vdd.n1169 146.341
R16901 vdd.n1466 vdd.n1169 146.341
R16902 vdd.n1466 vdd.n1165 146.341
R16903 vdd.n1472 vdd.n1165 146.341
R16904 vdd.n1472 vdd.n886 146.341
R16905 vdd.n1482 vdd.n886 146.341
R16906 vdd.n1482 vdd.n882 146.341
R16907 vdd.n1488 vdd.n882 146.341
R16908 vdd.n1488 vdd.n876 146.341
R16909 vdd.n1499 vdd.n876 146.341
R16910 vdd.n1499 vdd.n871 146.341
R16911 vdd.n1507 vdd.n871 146.341
R16912 vdd.n1507 vdd.n861 146.341
R16913 vdd.n1944 vdd.n861 146.341
R16914 vdd.n1420 vdd.n1196 146.341
R16915 vdd.n1420 vdd.n1229 146.341
R16916 vdd.n1233 vdd.n1232 146.341
R16917 vdd.n1235 vdd.n1234 146.341
R16918 vdd.n1239 vdd.n1238 146.341
R16919 vdd.n1241 vdd.n1240 146.341
R16920 vdd.n1245 vdd.n1244 146.341
R16921 vdd.n1247 vdd.n1246 146.341
R16922 vdd.n1251 vdd.n1250 146.341
R16923 vdd.n1253 vdd.n1252 146.341
R16924 vdd.n1259 vdd.n1258 146.341
R16925 vdd.n1261 vdd.n1260 146.341
R16926 vdd.n1265 vdd.n1264 146.341
R16927 vdd.n1267 vdd.n1266 146.341
R16928 vdd.n1271 vdd.n1270 146.341
R16929 vdd.n1273 vdd.n1272 146.341
R16930 vdd.n1277 vdd.n1276 146.341
R16931 vdd.n1279 vdd.n1278 146.341
R16932 vdd.n1283 vdd.n1282 146.341
R16933 vdd.n1285 vdd.n1284 146.341
R16934 vdd.n1357 vdd.n1288 146.341
R16935 vdd.n1290 vdd.n1289 146.341
R16936 vdd.n1294 vdd.n1293 146.341
R16937 vdd.n1296 vdd.n1295 146.341
R16938 vdd.n1300 vdd.n1299 146.341
R16939 vdd.n1302 vdd.n1301 146.341
R16940 vdd.n1306 vdd.n1305 146.341
R16941 vdd.n1308 vdd.n1307 146.341
R16942 vdd.n1312 vdd.n1311 146.341
R16943 vdd.n1314 vdd.n1313 146.341
R16944 vdd.n1318 vdd.n1317 146.341
R16945 vdd.n1319 vdd.n1227 146.341
R16946 vdd.n1429 vdd.n1192 146.341
R16947 vdd.n1429 vdd.n1185 146.341
R16948 vdd.n1440 vdd.n1185 146.341
R16949 vdd.n1440 vdd.n1181 146.341
R16950 vdd.n1446 vdd.n1181 146.341
R16951 vdd.n1446 vdd.n1174 146.341
R16952 vdd.n1457 vdd.n1174 146.341
R16953 vdd.n1457 vdd.n1170 146.341
R16954 vdd.n1464 vdd.n1170 146.341
R16955 vdd.n1464 vdd.n1163 146.341
R16956 vdd.n1474 vdd.n1163 146.341
R16957 vdd.n1474 vdd.n889 146.341
R16958 vdd.n1480 vdd.n889 146.341
R16959 vdd.n1480 vdd.n881 146.341
R16960 vdd.n1491 vdd.n881 146.341
R16961 vdd.n1491 vdd.n877 146.341
R16962 vdd.n1497 vdd.n877 146.341
R16963 vdd.n1497 vdd.n869 146.341
R16964 vdd.n1510 vdd.n869 146.341
R16965 vdd.n1510 vdd.n864 146.341
R16966 vdd.n1942 vdd.n864 146.341
R16967 vdd.n863 vdd.n839 141.707
R16968 vdd.n2840 vdd.n484 141.707
R16969 vdd.n1791 vdd.t131 127.284
R16970 vdd.n755 vdd.t115 127.284
R16971 vdd.n1765 vdd.t156 127.284
R16972 vdd.n747 vdd.t146 127.284
R16973 vdd.n2536 vdd.t98 127.284
R16974 vdd.n2536 vdd.t99 127.284
R16975 vdd.n2256 vdd.t138 127.284
R16976 vdd.n622 vdd.t119 127.284
R16977 vdd.n2253 vdd.t124 127.284
R16978 vdd.n589 vdd.t126 127.284
R16979 vdd.n817 vdd.t134 127.284
R16980 vdd.n817 vdd.t135 127.284
R16981 vdd.n22 vdd.n20 117.314
R16982 vdd.n17 vdd.n15 117.314
R16983 vdd.n27 vdd.n26 116.927
R16984 vdd.n24 vdd.n23 116.927
R16985 vdd.n22 vdd.n21 116.927
R16986 vdd.n17 vdd.n16 116.927
R16987 vdd.n19 vdd.n18 116.927
R16988 vdd.n27 vdd.n25 116.927
R16989 vdd.n1792 vdd.t130 111.188
R16990 vdd.n756 vdd.t116 111.188
R16991 vdd.n1766 vdd.t155 111.188
R16992 vdd.n748 vdd.t147 111.188
R16993 vdd.n2257 vdd.t137 111.188
R16994 vdd.n623 vdd.t120 111.188
R16995 vdd.n2254 vdd.t123 111.188
R16996 vdd.n590 vdd.t127 111.188
R16997 vdd.n2479 vdd.n701 99.5127
R16998 vdd.n2483 vdd.n701 99.5127
R16999 vdd.n2483 vdd.n693 99.5127
R17000 vdd.n2491 vdd.n693 99.5127
R17001 vdd.n2491 vdd.n691 99.5127
R17002 vdd.n2495 vdd.n691 99.5127
R17003 vdd.n2495 vdd.n680 99.5127
R17004 vdd.n2503 vdd.n680 99.5127
R17005 vdd.n2503 vdd.n678 99.5127
R17006 vdd.n2507 vdd.n678 99.5127
R17007 vdd.n2507 vdd.n669 99.5127
R17008 vdd.n2515 vdd.n669 99.5127
R17009 vdd.n2515 vdd.n667 99.5127
R17010 vdd.n2519 vdd.n667 99.5127
R17011 vdd.n2519 vdd.n657 99.5127
R17012 vdd.n2527 vdd.n657 99.5127
R17013 vdd.n2527 vdd.n655 99.5127
R17014 vdd.n2531 vdd.n655 99.5127
R17015 vdd.n2531 vdd.n646 99.5127
R17016 vdd.n2541 vdd.n646 99.5127
R17017 vdd.n2541 vdd.n644 99.5127
R17018 vdd.n2545 vdd.n644 99.5127
R17019 vdd.n2545 vdd.n632 99.5127
R17020 vdd.n2598 vdd.n632 99.5127
R17021 vdd.n2598 vdd.n630 99.5127
R17022 vdd.n2602 vdd.n630 99.5127
R17023 vdd.n2602 vdd.n598 99.5127
R17024 vdd.n2672 vdd.n598 99.5127
R17025 vdd.n2668 vdd.n599 99.5127
R17026 vdd.n2666 vdd.n2665 99.5127
R17027 vdd.n2663 vdd.n603 99.5127
R17028 vdd.n2659 vdd.n2658 99.5127
R17029 vdd.n2656 vdd.n606 99.5127
R17030 vdd.n2652 vdd.n2651 99.5127
R17031 vdd.n2649 vdd.n609 99.5127
R17032 vdd.n2645 vdd.n2644 99.5127
R17033 vdd.n2642 vdd.n2640 99.5127
R17034 vdd.n2638 vdd.n612 99.5127
R17035 vdd.n2634 vdd.n2633 99.5127
R17036 vdd.n2631 vdd.n615 99.5127
R17037 vdd.n2627 vdd.n2626 99.5127
R17038 vdd.n2624 vdd.n618 99.5127
R17039 vdd.n2620 vdd.n2619 99.5127
R17040 vdd.n2617 vdd.n621 99.5127
R17041 vdd.n2612 vdd.n2611 99.5127
R17042 vdd.n2399 vdd.n704 99.5127
R17043 vdd.n2399 vdd.n699 99.5127
R17044 vdd.n2396 vdd.n699 99.5127
R17045 vdd.n2396 vdd.n694 99.5127
R17046 vdd.n2343 vdd.n694 99.5127
R17047 vdd.n2343 vdd.n688 99.5127
R17048 vdd.n2346 vdd.n688 99.5127
R17049 vdd.n2346 vdd.n681 99.5127
R17050 vdd.n2349 vdd.n681 99.5127
R17051 vdd.n2349 vdd.n676 99.5127
R17052 vdd.n2352 vdd.n676 99.5127
R17053 vdd.n2352 vdd.n671 99.5127
R17054 vdd.n2355 vdd.n671 99.5127
R17055 vdd.n2355 vdd.n665 99.5127
R17056 vdd.n2373 vdd.n665 99.5127
R17057 vdd.n2373 vdd.n658 99.5127
R17058 vdd.n2369 vdd.n658 99.5127
R17059 vdd.n2369 vdd.n653 99.5127
R17060 vdd.n2366 vdd.n653 99.5127
R17061 vdd.n2366 vdd.n648 99.5127
R17062 vdd.n2363 vdd.n648 99.5127
R17063 vdd.n2363 vdd.n642 99.5127
R17064 vdd.n2360 vdd.n642 99.5127
R17065 vdd.n2360 vdd.n634 99.5127
R17066 vdd.n634 vdd.n627 99.5127
R17067 vdd.n2604 vdd.n627 99.5127
R17068 vdd.n2605 vdd.n2604 99.5127
R17069 vdd.n2605 vdd.n596 99.5127
R17070 vdd.n2469 vdd.n2252 99.5127
R17071 vdd.n2465 vdd.n2252 99.5127
R17072 vdd.n2463 vdd.n2462 99.5127
R17073 vdd.n2459 vdd.n2458 99.5127
R17074 vdd.n2455 vdd.n2454 99.5127
R17075 vdd.n2451 vdd.n2450 99.5127
R17076 vdd.n2447 vdd.n2446 99.5127
R17077 vdd.n2443 vdd.n2442 99.5127
R17078 vdd.n2439 vdd.n2438 99.5127
R17079 vdd.n2435 vdd.n2434 99.5127
R17080 vdd.n2431 vdd.n2430 99.5127
R17081 vdd.n2427 vdd.n2426 99.5127
R17082 vdd.n2423 vdd.n2422 99.5127
R17083 vdd.n2419 vdd.n2418 99.5127
R17084 vdd.n2415 vdd.n2414 99.5127
R17085 vdd.n2411 vdd.n2410 99.5127
R17086 vdd.n2406 vdd.n2405 99.5127
R17087 vdd.n2217 vdd.n745 99.5127
R17088 vdd.n2213 vdd.n2212 99.5127
R17089 vdd.n2209 vdd.n2208 99.5127
R17090 vdd.n2205 vdd.n2204 99.5127
R17091 vdd.n2201 vdd.n2200 99.5127
R17092 vdd.n2197 vdd.n2196 99.5127
R17093 vdd.n2193 vdd.n2192 99.5127
R17094 vdd.n2189 vdd.n2188 99.5127
R17095 vdd.n2185 vdd.n2184 99.5127
R17096 vdd.n2181 vdd.n2180 99.5127
R17097 vdd.n2177 vdd.n2176 99.5127
R17098 vdd.n2173 vdd.n2172 99.5127
R17099 vdd.n2169 vdd.n2168 99.5127
R17100 vdd.n2165 vdd.n2164 99.5127
R17101 vdd.n2161 vdd.n2160 99.5127
R17102 vdd.n2157 vdd.n2156 99.5127
R17103 vdd.n2152 vdd.n2151 99.5127
R17104 vdd.n1890 vdd.n840 99.5127
R17105 vdd.n1890 vdd.n834 99.5127
R17106 vdd.n1887 vdd.n834 99.5127
R17107 vdd.n1887 vdd.n828 99.5127
R17108 vdd.n1884 vdd.n828 99.5127
R17109 vdd.n1884 vdd.n821 99.5127
R17110 vdd.n1881 vdd.n821 99.5127
R17111 vdd.n1881 vdd.n814 99.5127
R17112 vdd.n1878 vdd.n814 99.5127
R17113 vdd.n1878 vdd.n809 99.5127
R17114 vdd.n1875 vdd.n809 99.5127
R17115 vdd.n1875 vdd.n803 99.5127
R17116 vdd.n1872 vdd.n803 99.5127
R17117 vdd.n1872 vdd.n796 99.5127
R17118 vdd.n1786 vdd.n796 99.5127
R17119 vdd.n1786 vdd.n790 99.5127
R17120 vdd.n1783 vdd.n790 99.5127
R17121 vdd.n1783 vdd.n785 99.5127
R17122 vdd.n1780 vdd.n785 99.5127
R17123 vdd.n1780 vdd.n780 99.5127
R17124 vdd.n1777 vdd.n780 99.5127
R17125 vdd.n1777 vdd.n774 99.5127
R17126 vdd.n1774 vdd.n774 99.5127
R17127 vdd.n1774 vdd.n767 99.5127
R17128 vdd.n1771 vdd.n767 99.5127
R17129 vdd.n1771 vdd.n760 99.5127
R17130 vdd.n760 vdd.n750 99.5127
R17131 vdd.n2147 vdd.n750 99.5127
R17132 vdd.n1725 vdd.n1723 99.5127
R17133 vdd.n1729 vdd.n1723 99.5127
R17134 vdd.n1733 vdd.n1731 99.5127
R17135 vdd.n1737 vdd.n1721 99.5127
R17136 vdd.n1741 vdd.n1739 99.5127
R17137 vdd.n1745 vdd.n1719 99.5127
R17138 vdd.n1749 vdd.n1747 99.5127
R17139 vdd.n1753 vdd.n1717 99.5127
R17140 vdd.n1756 vdd.n1755 99.5127
R17141 vdd.n1926 vdd.n1924 99.5127
R17142 vdd.n1922 vdd.n1758 99.5127
R17143 vdd.n1918 vdd.n1916 99.5127
R17144 vdd.n1914 vdd.n1760 99.5127
R17145 vdd.n1910 vdd.n1908 99.5127
R17146 vdd.n1906 vdd.n1762 99.5127
R17147 vdd.n1902 vdd.n1900 99.5127
R17148 vdd.n1898 vdd.n1764 99.5127
R17149 vdd.n1990 vdd.n836 99.5127
R17150 vdd.n1994 vdd.n836 99.5127
R17151 vdd.n1994 vdd.n826 99.5127
R17152 vdd.n2002 vdd.n826 99.5127
R17153 vdd.n2002 vdd.n824 99.5127
R17154 vdd.n2006 vdd.n824 99.5127
R17155 vdd.n2006 vdd.n813 99.5127
R17156 vdd.n2015 vdd.n813 99.5127
R17157 vdd.n2015 vdd.n811 99.5127
R17158 vdd.n2019 vdd.n811 99.5127
R17159 vdd.n2019 vdd.n801 99.5127
R17160 vdd.n2027 vdd.n801 99.5127
R17161 vdd.n2027 vdd.n799 99.5127
R17162 vdd.n2031 vdd.n799 99.5127
R17163 vdd.n2031 vdd.n789 99.5127
R17164 vdd.n2039 vdd.n789 99.5127
R17165 vdd.n2039 vdd.n787 99.5127
R17166 vdd.n2043 vdd.n787 99.5127
R17167 vdd.n2043 vdd.n778 99.5127
R17168 vdd.n2051 vdd.n778 99.5127
R17169 vdd.n2051 vdd.n776 99.5127
R17170 vdd.n2055 vdd.n776 99.5127
R17171 vdd.n2055 vdd.n765 99.5127
R17172 vdd.n2065 vdd.n765 99.5127
R17173 vdd.n2065 vdd.n762 99.5127
R17174 vdd.n2070 vdd.n762 99.5127
R17175 vdd.n2070 vdd.n763 99.5127
R17176 vdd.n763 vdd.n744 99.5127
R17177 vdd.n2588 vdd.n2587 99.5127
R17178 vdd.n2585 vdd.n2551 99.5127
R17179 vdd.n2581 vdd.n2580 99.5127
R17180 vdd.n2578 vdd.n2554 99.5127
R17181 vdd.n2574 vdd.n2573 99.5127
R17182 vdd.n2571 vdd.n2557 99.5127
R17183 vdd.n2567 vdd.n2566 99.5127
R17184 vdd.n2564 vdd.n2561 99.5127
R17185 vdd.n2705 vdd.n577 99.5127
R17186 vdd.n2703 vdd.n2702 99.5127
R17187 vdd.n2700 vdd.n579 99.5127
R17188 vdd.n2696 vdd.n2695 99.5127
R17189 vdd.n2693 vdd.n582 99.5127
R17190 vdd.n2689 vdd.n2688 99.5127
R17191 vdd.n2686 vdd.n585 99.5127
R17192 vdd.n2682 vdd.n2681 99.5127
R17193 vdd.n2679 vdd.n588 99.5127
R17194 vdd.n2323 vdd.n705 99.5127
R17195 vdd.n2323 vdd.n700 99.5127
R17196 vdd.n2394 vdd.n700 99.5127
R17197 vdd.n2394 vdd.n695 99.5127
R17198 vdd.n2390 vdd.n695 99.5127
R17199 vdd.n2390 vdd.n689 99.5127
R17200 vdd.n2387 vdd.n689 99.5127
R17201 vdd.n2387 vdd.n682 99.5127
R17202 vdd.n2384 vdd.n682 99.5127
R17203 vdd.n2384 vdd.n677 99.5127
R17204 vdd.n2381 vdd.n677 99.5127
R17205 vdd.n2381 vdd.n672 99.5127
R17206 vdd.n2378 vdd.n672 99.5127
R17207 vdd.n2378 vdd.n666 99.5127
R17208 vdd.n2375 vdd.n666 99.5127
R17209 vdd.n2375 vdd.n659 99.5127
R17210 vdd.n2340 vdd.n659 99.5127
R17211 vdd.n2340 vdd.n654 99.5127
R17212 vdd.n2337 vdd.n654 99.5127
R17213 vdd.n2337 vdd.n649 99.5127
R17214 vdd.n2334 vdd.n649 99.5127
R17215 vdd.n2334 vdd.n643 99.5127
R17216 vdd.n2331 vdd.n643 99.5127
R17217 vdd.n2331 vdd.n635 99.5127
R17218 vdd.n2328 vdd.n635 99.5127
R17219 vdd.n2328 vdd.n628 99.5127
R17220 vdd.n628 vdd.n594 99.5127
R17221 vdd.n2674 vdd.n594 99.5127
R17222 vdd.n2473 vdd.n708 99.5127
R17223 vdd.n2261 vdd.n2260 99.5127
R17224 vdd.n2265 vdd.n2264 99.5127
R17225 vdd.n2269 vdd.n2268 99.5127
R17226 vdd.n2273 vdd.n2272 99.5127
R17227 vdd.n2277 vdd.n2276 99.5127
R17228 vdd.n2281 vdd.n2280 99.5127
R17229 vdd.n2285 vdd.n2284 99.5127
R17230 vdd.n2289 vdd.n2288 99.5127
R17231 vdd.n2293 vdd.n2292 99.5127
R17232 vdd.n2297 vdd.n2296 99.5127
R17233 vdd.n2301 vdd.n2300 99.5127
R17234 vdd.n2305 vdd.n2304 99.5127
R17235 vdd.n2309 vdd.n2308 99.5127
R17236 vdd.n2313 vdd.n2312 99.5127
R17237 vdd.n2317 vdd.n2316 99.5127
R17238 vdd.n2319 vdd.n2251 99.5127
R17239 vdd.n2477 vdd.n698 99.5127
R17240 vdd.n2485 vdd.n698 99.5127
R17241 vdd.n2485 vdd.n696 99.5127
R17242 vdd.n2489 vdd.n696 99.5127
R17243 vdd.n2489 vdd.n686 99.5127
R17244 vdd.n2497 vdd.n686 99.5127
R17245 vdd.n2497 vdd.n684 99.5127
R17246 vdd.n2501 vdd.n684 99.5127
R17247 vdd.n2501 vdd.n675 99.5127
R17248 vdd.n2509 vdd.n675 99.5127
R17249 vdd.n2509 vdd.n673 99.5127
R17250 vdd.n2513 vdd.n673 99.5127
R17251 vdd.n2513 vdd.n663 99.5127
R17252 vdd.n2521 vdd.n663 99.5127
R17253 vdd.n2521 vdd.n661 99.5127
R17254 vdd.n2525 vdd.n661 99.5127
R17255 vdd.n2525 vdd.n652 99.5127
R17256 vdd.n2533 vdd.n652 99.5127
R17257 vdd.n2533 vdd.n650 99.5127
R17258 vdd.n2539 vdd.n650 99.5127
R17259 vdd.n2539 vdd.n640 99.5127
R17260 vdd.n2547 vdd.n640 99.5127
R17261 vdd.n2547 vdd.n637 99.5127
R17262 vdd.n2596 vdd.n637 99.5127
R17263 vdd.n2596 vdd.n638 99.5127
R17264 vdd.n638 vdd.n629 99.5127
R17265 vdd.n2591 vdd.n629 99.5127
R17266 vdd.n2591 vdd.n597 99.5127
R17267 vdd.n2141 vdd.n2140 99.5127
R17268 vdd.n2137 vdd.n2136 99.5127
R17269 vdd.n2133 vdd.n2132 99.5127
R17270 vdd.n2129 vdd.n2128 99.5127
R17271 vdd.n2125 vdd.n2124 99.5127
R17272 vdd.n2121 vdd.n2120 99.5127
R17273 vdd.n2117 vdd.n2116 99.5127
R17274 vdd.n2113 vdd.n2112 99.5127
R17275 vdd.n2109 vdd.n2108 99.5127
R17276 vdd.n2105 vdd.n2104 99.5127
R17277 vdd.n2101 vdd.n2100 99.5127
R17278 vdd.n2097 vdd.n2096 99.5127
R17279 vdd.n2093 vdd.n2092 99.5127
R17280 vdd.n2089 vdd.n2088 99.5127
R17281 vdd.n2085 vdd.n2084 99.5127
R17282 vdd.n2081 vdd.n2080 99.5127
R17283 vdd.n2077 vdd.n726 99.5127
R17284 vdd.n1834 vdd.n841 99.5127
R17285 vdd.n1834 vdd.n835 99.5127
R17286 vdd.n1837 vdd.n835 99.5127
R17287 vdd.n1837 vdd.n829 99.5127
R17288 vdd.n1840 vdd.n829 99.5127
R17289 vdd.n1840 vdd.n822 99.5127
R17290 vdd.n1843 vdd.n822 99.5127
R17291 vdd.n1843 vdd.n815 99.5127
R17292 vdd.n1846 vdd.n815 99.5127
R17293 vdd.n1846 vdd.n810 99.5127
R17294 vdd.n1849 vdd.n810 99.5127
R17295 vdd.n1849 vdd.n804 99.5127
R17296 vdd.n1870 vdd.n804 99.5127
R17297 vdd.n1870 vdd.n797 99.5127
R17298 vdd.n1866 vdd.n797 99.5127
R17299 vdd.n1866 vdd.n791 99.5127
R17300 vdd.n1863 vdd.n791 99.5127
R17301 vdd.n1863 vdd.n786 99.5127
R17302 vdd.n1860 vdd.n786 99.5127
R17303 vdd.n1860 vdd.n781 99.5127
R17304 vdd.n1857 vdd.n781 99.5127
R17305 vdd.n1857 vdd.n775 99.5127
R17306 vdd.n1854 vdd.n775 99.5127
R17307 vdd.n1854 vdd.n768 99.5127
R17308 vdd.n768 vdd.n759 99.5127
R17309 vdd.n2072 vdd.n759 99.5127
R17310 vdd.n2073 vdd.n2072 99.5127
R17311 vdd.n2073 vdd.n751 99.5127
R17312 vdd.n1984 vdd.n1982 99.5127
R17313 vdd.n1980 vdd.n844 99.5127
R17314 vdd.n1976 vdd.n1974 99.5127
R17315 vdd.n1972 vdd.n846 99.5127
R17316 vdd.n1968 vdd.n1966 99.5127
R17317 vdd.n1964 vdd.n848 99.5127
R17318 vdd.n1960 vdd.n1958 99.5127
R17319 vdd.n1956 vdd.n850 99.5127
R17320 vdd.n1798 vdd.n852 99.5127
R17321 vdd.n1803 vdd.n1800 99.5127
R17322 vdd.n1807 vdd.n1805 99.5127
R17323 vdd.n1811 vdd.n1796 99.5127
R17324 vdd.n1815 vdd.n1813 99.5127
R17325 vdd.n1819 vdd.n1794 99.5127
R17326 vdd.n1823 vdd.n1821 99.5127
R17327 vdd.n1828 vdd.n1790 99.5127
R17328 vdd.n1831 vdd.n1830 99.5127
R17329 vdd.n1988 vdd.n832 99.5127
R17330 vdd.n1996 vdd.n832 99.5127
R17331 vdd.n1996 vdd.n830 99.5127
R17332 vdd.n2000 vdd.n830 99.5127
R17333 vdd.n2000 vdd.n819 99.5127
R17334 vdd.n2008 vdd.n819 99.5127
R17335 vdd.n2008 vdd.n816 99.5127
R17336 vdd.n2013 vdd.n816 99.5127
R17337 vdd.n2013 vdd.n807 99.5127
R17338 vdd.n2021 vdd.n807 99.5127
R17339 vdd.n2021 vdd.n805 99.5127
R17340 vdd.n2025 vdd.n805 99.5127
R17341 vdd.n2025 vdd.n795 99.5127
R17342 vdd.n2033 vdd.n795 99.5127
R17343 vdd.n2033 vdd.n793 99.5127
R17344 vdd.n2037 vdd.n793 99.5127
R17345 vdd.n2037 vdd.n784 99.5127
R17346 vdd.n2045 vdd.n784 99.5127
R17347 vdd.n2045 vdd.n782 99.5127
R17348 vdd.n2049 vdd.n782 99.5127
R17349 vdd.n2049 vdd.n772 99.5127
R17350 vdd.n2057 vdd.n772 99.5127
R17351 vdd.n2057 vdd.n769 99.5127
R17352 vdd.n2063 vdd.n769 99.5127
R17353 vdd.n2063 vdd.n770 99.5127
R17354 vdd.n770 vdd.n761 99.5127
R17355 vdd.n761 vdd.n752 99.5127
R17356 vdd.n2145 vdd.n752 99.5127
R17357 vdd.n9 vdd.n7 98.9633
R17358 vdd.n2 vdd.n0 98.9633
R17359 vdd.n9 vdd.n8 98.6055
R17360 vdd.n11 vdd.n10 98.6055
R17361 vdd.n13 vdd.n12 98.6055
R17362 vdd.n6 vdd.n5 98.6055
R17363 vdd.n4 vdd.n3 98.6055
R17364 vdd.n2 vdd.n1 98.6055
R17365 vdd.t34 vdd.n267 85.8723
R17366 vdd.t45 vdd.n220 85.8723
R17367 vdd.t30 vdd.n177 85.8723
R17368 vdd.t40 vdd.n130 85.8723
R17369 vdd.t71 vdd.n88 85.8723
R17370 vdd.t13 vdd.n41 85.8723
R17371 vdd.t69 vdd.n1082 85.8723
R17372 vdd.t55 vdd.n1129 85.8723
R17373 vdd.t61 vdd.n992 85.8723
R17374 vdd.t48 vdd.n1039 85.8723
R17375 vdd.t11 vdd.n903 85.8723
R17376 vdd.t70 vdd.n950 85.8723
R17377 vdd.n2537 vdd.n2536 78.546
R17378 vdd.n2011 vdd.n817 78.546
R17379 vdd.n254 vdd.n253 75.1835
R17380 vdd.n252 vdd.n251 75.1835
R17381 vdd.n250 vdd.n249 75.1835
R17382 vdd.n164 vdd.n163 75.1835
R17383 vdd.n162 vdd.n161 75.1835
R17384 vdd.n160 vdd.n159 75.1835
R17385 vdd.n75 vdd.n74 75.1835
R17386 vdd.n73 vdd.n72 75.1835
R17387 vdd.n71 vdd.n70 75.1835
R17388 vdd.n1112 vdd.n1111 75.1835
R17389 vdd.n1114 vdd.n1113 75.1835
R17390 vdd.n1116 vdd.n1115 75.1835
R17391 vdd.n1022 vdd.n1021 75.1835
R17392 vdd.n1024 vdd.n1023 75.1835
R17393 vdd.n1026 vdd.n1025 75.1835
R17394 vdd.n933 vdd.n932 75.1835
R17395 vdd.n935 vdd.n934 75.1835
R17396 vdd.n937 vdd.n936 75.1835
R17397 vdd.n2472 vdd.n2471 72.8958
R17398 vdd.n2471 vdd.n2235 72.8958
R17399 vdd.n2471 vdd.n2236 72.8958
R17400 vdd.n2471 vdd.n2237 72.8958
R17401 vdd.n2471 vdd.n2238 72.8958
R17402 vdd.n2471 vdd.n2239 72.8958
R17403 vdd.n2471 vdd.n2240 72.8958
R17404 vdd.n2471 vdd.n2241 72.8958
R17405 vdd.n2471 vdd.n2242 72.8958
R17406 vdd.n2471 vdd.n2243 72.8958
R17407 vdd.n2471 vdd.n2244 72.8958
R17408 vdd.n2471 vdd.n2245 72.8958
R17409 vdd.n2471 vdd.n2246 72.8958
R17410 vdd.n2471 vdd.n2247 72.8958
R17411 vdd.n2471 vdd.n2248 72.8958
R17412 vdd.n2471 vdd.n2249 72.8958
R17413 vdd.n2471 vdd.n2250 72.8958
R17414 vdd.n593 vdd.n484 72.8958
R17415 vdd.n2680 vdd.n484 72.8958
R17416 vdd.n587 vdd.n484 72.8958
R17417 vdd.n2687 vdd.n484 72.8958
R17418 vdd.n584 vdd.n484 72.8958
R17419 vdd.n2694 vdd.n484 72.8958
R17420 vdd.n581 vdd.n484 72.8958
R17421 vdd.n2701 vdd.n484 72.8958
R17422 vdd.n2704 vdd.n484 72.8958
R17423 vdd.n2560 vdd.n484 72.8958
R17424 vdd.n2565 vdd.n484 72.8958
R17425 vdd.n2559 vdd.n484 72.8958
R17426 vdd.n2572 vdd.n484 72.8958
R17427 vdd.n2556 vdd.n484 72.8958
R17428 vdd.n2579 vdd.n484 72.8958
R17429 vdd.n2553 vdd.n484 72.8958
R17430 vdd.n2586 vdd.n484 72.8958
R17431 vdd.n1724 vdd.n839 72.8958
R17432 vdd.n1730 vdd.n839 72.8958
R17433 vdd.n1732 vdd.n839 72.8958
R17434 vdd.n1738 vdd.n839 72.8958
R17435 vdd.n1740 vdd.n839 72.8958
R17436 vdd.n1746 vdd.n839 72.8958
R17437 vdd.n1748 vdd.n839 72.8958
R17438 vdd.n1754 vdd.n839 72.8958
R17439 vdd.n1925 vdd.n839 72.8958
R17440 vdd.n1923 vdd.n839 72.8958
R17441 vdd.n1917 vdd.n839 72.8958
R17442 vdd.n1915 vdd.n839 72.8958
R17443 vdd.n1909 vdd.n839 72.8958
R17444 vdd.n1907 vdd.n839 72.8958
R17445 vdd.n1901 vdd.n839 72.8958
R17446 vdd.n1899 vdd.n839 72.8958
R17447 vdd.n1893 vdd.n839 72.8958
R17448 vdd.n2218 vdd.n727 72.8958
R17449 vdd.n2218 vdd.n728 72.8958
R17450 vdd.n2218 vdd.n729 72.8958
R17451 vdd.n2218 vdd.n730 72.8958
R17452 vdd.n2218 vdd.n731 72.8958
R17453 vdd.n2218 vdd.n732 72.8958
R17454 vdd.n2218 vdd.n733 72.8958
R17455 vdd.n2218 vdd.n734 72.8958
R17456 vdd.n2218 vdd.n735 72.8958
R17457 vdd.n2218 vdd.n736 72.8958
R17458 vdd.n2218 vdd.n737 72.8958
R17459 vdd.n2218 vdd.n738 72.8958
R17460 vdd.n2218 vdd.n739 72.8958
R17461 vdd.n2218 vdd.n740 72.8958
R17462 vdd.n2218 vdd.n741 72.8958
R17463 vdd.n2218 vdd.n742 72.8958
R17464 vdd.n2218 vdd.n743 72.8958
R17465 vdd.n2471 vdd.n2470 72.8958
R17466 vdd.n2471 vdd.n2219 72.8958
R17467 vdd.n2471 vdd.n2220 72.8958
R17468 vdd.n2471 vdd.n2221 72.8958
R17469 vdd.n2471 vdd.n2222 72.8958
R17470 vdd.n2471 vdd.n2223 72.8958
R17471 vdd.n2471 vdd.n2224 72.8958
R17472 vdd.n2471 vdd.n2225 72.8958
R17473 vdd.n2471 vdd.n2226 72.8958
R17474 vdd.n2471 vdd.n2227 72.8958
R17475 vdd.n2471 vdd.n2228 72.8958
R17476 vdd.n2471 vdd.n2229 72.8958
R17477 vdd.n2471 vdd.n2230 72.8958
R17478 vdd.n2471 vdd.n2231 72.8958
R17479 vdd.n2471 vdd.n2232 72.8958
R17480 vdd.n2471 vdd.n2233 72.8958
R17481 vdd.n2471 vdd.n2234 72.8958
R17482 vdd.n2610 vdd.n484 72.8958
R17483 vdd.n625 vdd.n484 72.8958
R17484 vdd.n2618 vdd.n484 72.8958
R17485 vdd.n620 vdd.n484 72.8958
R17486 vdd.n2625 vdd.n484 72.8958
R17487 vdd.n617 vdd.n484 72.8958
R17488 vdd.n2632 vdd.n484 72.8958
R17489 vdd.n614 vdd.n484 72.8958
R17490 vdd.n2639 vdd.n484 72.8958
R17491 vdd.n2643 vdd.n484 72.8958
R17492 vdd.n611 vdd.n484 72.8958
R17493 vdd.n2650 vdd.n484 72.8958
R17494 vdd.n608 vdd.n484 72.8958
R17495 vdd.n2657 vdd.n484 72.8958
R17496 vdd.n605 vdd.n484 72.8958
R17497 vdd.n2664 vdd.n484 72.8958
R17498 vdd.n2667 vdd.n484 72.8958
R17499 vdd.n2218 vdd.n725 72.8958
R17500 vdd.n2218 vdd.n724 72.8958
R17501 vdd.n2218 vdd.n723 72.8958
R17502 vdd.n2218 vdd.n722 72.8958
R17503 vdd.n2218 vdd.n721 72.8958
R17504 vdd.n2218 vdd.n720 72.8958
R17505 vdd.n2218 vdd.n719 72.8958
R17506 vdd.n2218 vdd.n718 72.8958
R17507 vdd.n2218 vdd.n717 72.8958
R17508 vdd.n2218 vdd.n716 72.8958
R17509 vdd.n2218 vdd.n715 72.8958
R17510 vdd.n2218 vdd.n714 72.8958
R17511 vdd.n2218 vdd.n713 72.8958
R17512 vdd.n2218 vdd.n712 72.8958
R17513 vdd.n2218 vdd.n711 72.8958
R17514 vdd.n2218 vdd.n710 72.8958
R17515 vdd.n2218 vdd.n709 72.8958
R17516 vdd.n1983 vdd.n839 72.8958
R17517 vdd.n1981 vdd.n839 72.8958
R17518 vdd.n1975 vdd.n839 72.8958
R17519 vdd.n1973 vdd.n839 72.8958
R17520 vdd.n1967 vdd.n839 72.8958
R17521 vdd.n1965 vdd.n839 72.8958
R17522 vdd.n1959 vdd.n839 72.8958
R17523 vdd.n1957 vdd.n839 72.8958
R17524 vdd.n851 vdd.n839 72.8958
R17525 vdd.n1799 vdd.n839 72.8958
R17526 vdd.n1804 vdd.n839 72.8958
R17527 vdd.n1806 vdd.n839 72.8958
R17528 vdd.n1812 vdd.n839 72.8958
R17529 vdd.n1814 vdd.n839 72.8958
R17530 vdd.n1820 vdd.n839 72.8958
R17531 vdd.n1822 vdd.n839 72.8958
R17532 vdd.n1829 vdd.n839 72.8958
R17533 vdd.n1422 vdd.n1421 66.2847
R17534 vdd.n1421 vdd.n1197 66.2847
R17535 vdd.n1421 vdd.n1198 66.2847
R17536 vdd.n1421 vdd.n1199 66.2847
R17537 vdd.n1421 vdd.n1200 66.2847
R17538 vdd.n1421 vdd.n1201 66.2847
R17539 vdd.n1421 vdd.n1202 66.2847
R17540 vdd.n1421 vdd.n1203 66.2847
R17541 vdd.n1421 vdd.n1204 66.2847
R17542 vdd.n1421 vdd.n1205 66.2847
R17543 vdd.n1421 vdd.n1206 66.2847
R17544 vdd.n1421 vdd.n1207 66.2847
R17545 vdd.n1421 vdd.n1208 66.2847
R17546 vdd.n1421 vdd.n1209 66.2847
R17547 vdd.n1421 vdd.n1210 66.2847
R17548 vdd.n1421 vdd.n1211 66.2847
R17549 vdd.n1421 vdd.n1212 66.2847
R17550 vdd.n1421 vdd.n1213 66.2847
R17551 vdd.n1421 vdd.n1214 66.2847
R17552 vdd.n1421 vdd.n1215 66.2847
R17553 vdd.n1421 vdd.n1216 66.2847
R17554 vdd.n1421 vdd.n1217 66.2847
R17555 vdd.n1421 vdd.n1218 66.2847
R17556 vdd.n1421 vdd.n1219 66.2847
R17557 vdd.n1421 vdd.n1220 66.2847
R17558 vdd.n1421 vdd.n1221 66.2847
R17559 vdd.n1421 vdd.n1222 66.2847
R17560 vdd.n1421 vdd.n1223 66.2847
R17561 vdd.n1421 vdd.n1224 66.2847
R17562 vdd.n1421 vdd.n1225 66.2847
R17563 vdd.n1421 vdd.n1226 66.2847
R17564 vdd.n863 vdd.n860 66.2847
R17565 vdd.n1614 vdd.n863 66.2847
R17566 vdd.n1619 vdd.n863 66.2847
R17567 vdd.n1624 vdd.n863 66.2847
R17568 vdd.n1612 vdd.n863 66.2847
R17569 vdd.n1631 vdd.n863 66.2847
R17570 vdd.n1604 vdd.n863 66.2847
R17571 vdd.n1638 vdd.n863 66.2847
R17572 vdd.n1597 vdd.n863 66.2847
R17573 vdd.n1645 vdd.n863 66.2847
R17574 vdd.n1591 vdd.n863 66.2847
R17575 vdd.n1586 vdd.n863 66.2847
R17576 vdd.n1656 vdd.n863 66.2847
R17577 vdd.n1578 vdd.n863 66.2847
R17578 vdd.n1663 vdd.n863 66.2847
R17579 vdd.n1571 vdd.n863 66.2847
R17580 vdd.n1670 vdd.n863 66.2847
R17581 vdd.n1564 vdd.n863 66.2847
R17582 vdd.n1677 vdd.n863 66.2847
R17583 vdd.n1557 vdd.n863 66.2847
R17584 vdd.n1684 vdd.n863 66.2847
R17585 vdd.n1551 vdd.n863 66.2847
R17586 vdd.n1546 vdd.n863 66.2847
R17587 vdd.n1695 vdd.n863 66.2847
R17588 vdd.n1538 vdd.n863 66.2847
R17589 vdd.n1702 vdd.n863 66.2847
R17590 vdd.n1531 vdd.n863 66.2847
R17591 vdd.n1709 vdd.n863 66.2847
R17592 vdd.n1712 vdd.n863 66.2847
R17593 vdd.n1522 vdd.n863 66.2847
R17594 vdd.n1934 vdd.n863 66.2847
R17595 vdd.n1516 vdd.n863 66.2847
R17596 vdd.n2841 vdd.n2840 66.2847
R17597 vdd.n2840 vdd.n485 66.2847
R17598 vdd.n2840 vdd.n486 66.2847
R17599 vdd.n2840 vdd.n487 66.2847
R17600 vdd.n2840 vdd.n488 66.2847
R17601 vdd.n2840 vdd.n489 66.2847
R17602 vdd.n2840 vdd.n490 66.2847
R17603 vdd.n2840 vdd.n491 66.2847
R17604 vdd.n2840 vdd.n492 66.2847
R17605 vdd.n2840 vdd.n493 66.2847
R17606 vdd.n2840 vdd.n494 66.2847
R17607 vdd.n2840 vdd.n495 66.2847
R17608 vdd.n2840 vdd.n496 66.2847
R17609 vdd.n2840 vdd.n497 66.2847
R17610 vdd.n2840 vdd.n498 66.2847
R17611 vdd.n2840 vdd.n499 66.2847
R17612 vdd.n2840 vdd.n500 66.2847
R17613 vdd.n2840 vdd.n501 66.2847
R17614 vdd.n2840 vdd.n502 66.2847
R17615 vdd.n2840 vdd.n503 66.2847
R17616 vdd.n2840 vdd.n504 66.2847
R17617 vdd.n2840 vdd.n505 66.2847
R17618 vdd.n2840 vdd.n506 66.2847
R17619 vdd.n2840 vdd.n507 66.2847
R17620 vdd.n2840 vdd.n508 66.2847
R17621 vdd.n2840 vdd.n509 66.2847
R17622 vdd.n2840 vdd.n510 66.2847
R17623 vdd.n2840 vdd.n511 66.2847
R17624 vdd.n2840 vdd.n512 66.2847
R17625 vdd.n2840 vdd.n513 66.2847
R17626 vdd.n2840 vdd.n514 66.2847
R17627 vdd.n2905 vdd.n329 66.2847
R17628 vdd.n2914 vdd.n329 66.2847
R17629 vdd.n439 vdd.n329 66.2847
R17630 vdd.n2921 vdd.n329 66.2847
R17631 vdd.n432 vdd.n329 66.2847
R17632 vdd.n2928 vdd.n329 66.2847
R17633 vdd.n425 vdd.n329 66.2847
R17634 vdd.n2935 vdd.n329 66.2847
R17635 vdd.n418 vdd.n329 66.2847
R17636 vdd.n2942 vdd.n329 66.2847
R17637 vdd.n412 vdd.n329 66.2847
R17638 vdd.n407 vdd.n329 66.2847
R17639 vdd.n2953 vdd.n329 66.2847
R17640 vdd.n399 vdd.n329 66.2847
R17641 vdd.n2960 vdd.n329 66.2847
R17642 vdd.n392 vdd.n329 66.2847
R17643 vdd.n2967 vdd.n329 66.2847
R17644 vdd.n385 vdd.n329 66.2847
R17645 vdd.n2974 vdd.n329 66.2847
R17646 vdd.n378 vdd.n329 66.2847
R17647 vdd.n2981 vdd.n329 66.2847
R17648 vdd.n372 vdd.n329 66.2847
R17649 vdd.n367 vdd.n329 66.2847
R17650 vdd.n2992 vdd.n329 66.2847
R17651 vdd.n359 vdd.n329 66.2847
R17652 vdd.n2999 vdd.n329 66.2847
R17653 vdd.n352 vdd.n329 66.2847
R17654 vdd.n3006 vdd.n329 66.2847
R17655 vdd.n345 vdd.n329 66.2847
R17656 vdd.n3013 vdd.n329 66.2847
R17657 vdd.n3016 vdd.n329 66.2847
R17658 vdd.n333 vdd.n329 66.2847
R17659 vdd.n334 vdd.n333 52.4337
R17660 vdd.n3016 vdd.n3015 52.4337
R17661 vdd.n3013 vdd.n3012 52.4337
R17662 vdd.n3008 vdd.n345 52.4337
R17663 vdd.n3006 vdd.n3005 52.4337
R17664 vdd.n3001 vdd.n352 52.4337
R17665 vdd.n2999 vdd.n2998 52.4337
R17666 vdd.n2994 vdd.n359 52.4337
R17667 vdd.n2992 vdd.n2991 52.4337
R17668 vdd.n368 vdd.n367 52.4337
R17669 vdd.n2983 vdd.n372 52.4337
R17670 vdd.n2981 vdd.n2980 52.4337
R17671 vdd.n2976 vdd.n378 52.4337
R17672 vdd.n2974 vdd.n2973 52.4337
R17673 vdd.n2969 vdd.n385 52.4337
R17674 vdd.n2967 vdd.n2966 52.4337
R17675 vdd.n2962 vdd.n392 52.4337
R17676 vdd.n2960 vdd.n2959 52.4337
R17677 vdd.n2955 vdd.n399 52.4337
R17678 vdd.n2953 vdd.n2952 52.4337
R17679 vdd.n408 vdd.n407 52.4337
R17680 vdd.n2944 vdd.n412 52.4337
R17681 vdd.n2942 vdd.n2941 52.4337
R17682 vdd.n2937 vdd.n418 52.4337
R17683 vdd.n2935 vdd.n2934 52.4337
R17684 vdd.n2930 vdd.n425 52.4337
R17685 vdd.n2928 vdd.n2927 52.4337
R17686 vdd.n2923 vdd.n432 52.4337
R17687 vdd.n2921 vdd.n2920 52.4337
R17688 vdd.n2916 vdd.n439 52.4337
R17689 vdd.n2914 vdd.n2913 52.4337
R17690 vdd.n2906 vdd.n2905 52.4337
R17691 vdd.n2842 vdd.n2841 52.4337
R17692 vdd.n517 vdd.n485 52.4337
R17693 vdd.n523 vdd.n486 52.4337
R17694 vdd.n2831 vdd.n487 52.4337
R17695 vdd.n2827 vdd.n488 52.4337
R17696 vdd.n2823 vdd.n489 52.4337
R17697 vdd.n2819 vdd.n490 52.4337
R17698 vdd.n2815 vdd.n491 52.4337
R17699 vdd.n2811 vdd.n492 52.4337
R17700 vdd.n2807 vdd.n493 52.4337
R17701 vdd.n2799 vdd.n494 52.4337
R17702 vdd.n2795 vdd.n495 52.4337
R17703 vdd.n2791 vdd.n496 52.4337
R17704 vdd.n2787 vdd.n497 52.4337
R17705 vdd.n2783 vdd.n498 52.4337
R17706 vdd.n2779 vdd.n499 52.4337
R17707 vdd.n2775 vdd.n500 52.4337
R17708 vdd.n2771 vdd.n501 52.4337
R17709 vdd.n2767 vdd.n502 52.4337
R17710 vdd.n2763 vdd.n503 52.4337
R17711 vdd.n2759 vdd.n504 52.4337
R17712 vdd.n2753 vdd.n505 52.4337
R17713 vdd.n2749 vdd.n506 52.4337
R17714 vdd.n2745 vdd.n507 52.4337
R17715 vdd.n2741 vdd.n508 52.4337
R17716 vdd.n2737 vdd.n509 52.4337
R17717 vdd.n2733 vdd.n510 52.4337
R17718 vdd.n2729 vdd.n511 52.4337
R17719 vdd.n2725 vdd.n512 52.4337
R17720 vdd.n2721 vdd.n513 52.4337
R17721 vdd.n2717 vdd.n514 52.4337
R17722 vdd.n1936 vdd.n1516 52.4337
R17723 vdd.n1934 vdd.n1933 52.4337
R17724 vdd.n1523 vdd.n1522 52.4337
R17725 vdd.n1712 vdd.n1711 52.4337
R17726 vdd.n1709 vdd.n1708 52.4337
R17727 vdd.n1704 vdd.n1531 52.4337
R17728 vdd.n1702 vdd.n1701 52.4337
R17729 vdd.n1697 vdd.n1538 52.4337
R17730 vdd.n1695 vdd.n1694 52.4337
R17731 vdd.n1547 vdd.n1546 52.4337
R17732 vdd.n1686 vdd.n1551 52.4337
R17733 vdd.n1684 vdd.n1683 52.4337
R17734 vdd.n1679 vdd.n1557 52.4337
R17735 vdd.n1677 vdd.n1676 52.4337
R17736 vdd.n1672 vdd.n1564 52.4337
R17737 vdd.n1670 vdd.n1669 52.4337
R17738 vdd.n1665 vdd.n1571 52.4337
R17739 vdd.n1663 vdd.n1662 52.4337
R17740 vdd.n1658 vdd.n1578 52.4337
R17741 vdd.n1656 vdd.n1655 52.4337
R17742 vdd.n1587 vdd.n1586 52.4337
R17743 vdd.n1647 vdd.n1591 52.4337
R17744 vdd.n1645 vdd.n1644 52.4337
R17745 vdd.n1640 vdd.n1597 52.4337
R17746 vdd.n1638 vdd.n1637 52.4337
R17747 vdd.n1633 vdd.n1604 52.4337
R17748 vdd.n1631 vdd.n1630 52.4337
R17749 vdd.n1626 vdd.n1612 52.4337
R17750 vdd.n1624 vdd.n1623 52.4337
R17751 vdd.n1619 vdd.n1618 52.4337
R17752 vdd.n1614 vdd.n1613 52.4337
R17753 vdd.n1945 vdd.n860 52.4337
R17754 vdd.n1423 vdd.n1422 52.4337
R17755 vdd.n1229 vdd.n1197 52.4337
R17756 vdd.n1233 vdd.n1198 52.4337
R17757 vdd.n1235 vdd.n1199 52.4337
R17758 vdd.n1239 vdd.n1200 52.4337
R17759 vdd.n1241 vdd.n1201 52.4337
R17760 vdd.n1245 vdd.n1202 52.4337
R17761 vdd.n1247 vdd.n1203 52.4337
R17762 vdd.n1251 vdd.n1204 52.4337
R17763 vdd.n1253 vdd.n1205 52.4337
R17764 vdd.n1259 vdd.n1206 52.4337
R17765 vdd.n1261 vdd.n1207 52.4337
R17766 vdd.n1265 vdd.n1208 52.4337
R17767 vdd.n1267 vdd.n1209 52.4337
R17768 vdd.n1271 vdd.n1210 52.4337
R17769 vdd.n1273 vdd.n1211 52.4337
R17770 vdd.n1277 vdd.n1212 52.4337
R17771 vdd.n1279 vdd.n1213 52.4337
R17772 vdd.n1283 vdd.n1214 52.4337
R17773 vdd.n1285 vdd.n1215 52.4337
R17774 vdd.n1357 vdd.n1216 52.4337
R17775 vdd.n1290 vdd.n1217 52.4337
R17776 vdd.n1294 vdd.n1218 52.4337
R17777 vdd.n1296 vdd.n1219 52.4337
R17778 vdd.n1300 vdd.n1220 52.4337
R17779 vdd.n1302 vdd.n1221 52.4337
R17780 vdd.n1306 vdd.n1222 52.4337
R17781 vdd.n1308 vdd.n1223 52.4337
R17782 vdd.n1312 vdd.n1224 52.4337
R17783 vdd.n1314 vdd.n1225 52.4337
R17784 vdd.n1318 vdd.n1226 52.4337
R17785 vdd.n1422 vdd.n1196 52.4337
R17786 vdd.n1232 vdd.n1197 52.4337
R17787 vdd.n1234 vdd.n1198 52.4337
R17788 vdd.n1238 vdd.n1199 52.4337
R17789 vdd.n1240 vdd.n1200 52.4337
R17790 vdd.n1244 vdd.n1201 52.4337
R17791 vdd.n1246 vdd.n1202 52.4337
R17792 vdd.n1250 vdd.n1203 52.4337
R17793 vdd.n1252 vdd.n1204 52.4337
R17794 vdd.n1258 vdd.n1205 52.4337
R17795 vdd.n1260 vdd.n1206 52.4337
R17796 vdd.n1264 vdd.n1207 52.4337
R17797 vdd.n1266 vdd.n1208 52.4337
R17798 vdd.n1270 vdd.n1209 52.4337
R17799 vdd.n1272 vdd.n1210 52.4337
R17800 vdd.n1276 vdd.n1211 52.4337
R17801 vdd.n1278 vdd.n1212 52.4337
R17802 vdd.n1282 vdd.n1213 52.4337
R17803 vdd.n1284 vdd.n1214 52.4337
R17804 vdd.n1288 vdd.n1215 52.4337
R17805 vdd.n1289 vdd.n1216 52.4337
R17806 vdd.n1293 vdd.n1217 52.4337
R17807 vdd.n1295 vdd.n1218 52.4337
R17808 vdd.n1299 vdd.n1219 52.4337
R17809 vdd.n1301 vdd.n1220 52.4337
R17810 vdd.n1305 vdd.n1221 52.4337
R17811 vdd.n1307 vdd.n1222 52.4337
R17812 vdd.n1311 vdd.n1223 52.4337
R17813 vdd.n1313 vdd.n1224 52.4337
R17814 vdd.n1317 vdd.n1225 52.4337
R17815 vdd.n1319 vdd.n1226 52.4337
R17816 vdd.n860 vdd.n859 52.4337
R17817 vdd.n1615 vdd.n1614 52.4337
R17818 vdd.n1620 vdd.n1619 52.4337
R17819 vdd.n1625 vdd.n1624 52.4337
R17820 vdd.n1612 vdd.n1605 52.4337
R17821 vdd.n1632 vdd.n1631 52.4337
R17822 vdd.n1604 vdd.n1598 52.4337
R17823 vdd.n1639 vdd.n1638 52.4337
R17824 vdd.n1597 vdd.n1592 52.4337
R17825 vdd.n1646 vdd.n1645 52.4337
R17826 vdd.n1591 vdd.n1590 52.4337
R17827 vdd.n1586 vdd.n1579 52.4337
R17828 vdd.n1657 vdd.n1656 52.4337
R17829 vdd.n1578 vdd.n1572 52.4337
R17830 vdd.n1664 vdd.n1663 52.4337
R17831 vdd.n1571 vdd.n1565 52.4337
R17832 vdd.n1671 vdd.n1670 52.4337
R17833 vdd.n1564 vdd.n1558 52.4337
R17834 vdd.n1678 vdd.n1677 52.4337
R17835 vdd.n1557 vdd.n1552 52.4337
R17836 vdd.n1685 vdd.n1684 52.4337
R17837 vdd.n1551 vdd.n1550 52.4337
R17838 vdd.n1546 vdd.n1539 52.4337
R17839 vdd.n1696 vdd.n1695 52.4337
R17840 vdd.n1538 vdd.n1532 52.4337
R17841 vdd.n1703 vdd.n1702 52.4337
R17842 vdd.n1531 vdd.n1525 52.4337
R17843 vdd.n1710 vdd.n1709 52.4337
R17844 vdd.n1713 vdd.n1712 52.4337
R17845 vdd.n1522 vdd.n1517 52.4337
R17846 vdd.n1935 vdd.n1934 52.4337
R17847 vdd.n1516 vdd.n865 52.4337
R17848 vdd.n2841 vdd.n483 52.4337
R17849 vdd.n522 vdd.n485 52.4337
R17850 vdd.n2832 vdd.n486 52.4337
R17851 vdd.n2828 vdd.n487 52.4337
R17852 vdd.n2824 vdd.n488 52.4337
R17853 vdd.n2820 vdd.n489 52.4337
R17854 vdd.n2816 vdd.n490 52.4337
R17855 vdd.n2812 vdd.n491 52.4337
R17856 vdd.n2808 vdd.n492 52.4337
R17857 vdd.n2798 vdd.n493 52.4337
R17858 vdd.n2796 vdd.n494 52.4337
R17859 vdd.n2792 vdd.n495 52.4337
R17860 vdd.n2788 vdd.n496 52.4337
R17861 vdd.n2784 vdd.n497 52.4337
R17862 vdd.n2780 vdd.n498 52.4337
R17863 vdd.n2776 vdd.n499 52.4337
R17864 vdd.n2772 vdd.n500 52.4337
R17865 vdd.n2768 vdd.n501 52.4337
R17866 vdd.n2764 vdd.n502 52.4337
R17867 vdd.n2760 vdd.n503 52.4337
R17868 vdd.n2752 vdd.n504 52.4337
R17869 vdd.n2750 vdd.n505 52.4337
R17870 vdd.n2746 vdd.n506 52.4337
R17871 vdd.n2742 vdd.n507 52.4337
R17872 vdd.n2738 vdd.n508 52.4337
R17873 vdd.n2734 vdd.n509 52.4337
R17874 vdd.n2730 vdd.n510 52.4337
R17875 vdd.n2726 vdd.n511 52.4337
R17876 vdd.n2722 vdd.n512 52.4337
R17877 vdd.n2718 vdd.n513 52.4337
R17878 vdd.n2714 vdd.n514 52.4337
R17879 vdd.n2905 vdd.n440 52.4337
R17880 vdd.n2915 vdd.n2914 52.4337
R17881 vdd.n439 vdd.n433 52.4337
R17882 vdd.n2922 vdd.n2921 52.4337
R17883 vdd.n432 vdd.n426 52.4337
R17884 vdd.n2929 vdd.n2928 52.4337
R17885 vdd.n425 vdd.n419 52.4337
R17886 vdd.n2936 vdd.n2935 52.4337
R17887 vdd.n418 vdd.n413 52.4337
R17888 vdd.n2943 vdd.n2942 52.4337
R17889 vdd.n412 vdd.n411 52.4337
R17890 vdd.n407 vdd.n400 52.4337
R17891 vdd.n2954 vdd.n2953 52.4337
R17892 vdd.n399 vdd.n393 52.4337
R17893 vdd.n2961 vdd.n2960 52.4337
R17894 vdd.n392 vdd.n386 52.4337
R17895 vdd.n2968 vdd.n2967 52.4337
R17896 vdd.n385 vdd.n379 52.4337
R17897 vdd.n2975 vdd.n2974 52.4337
R17898 vdd.n378 vdd.n373 52.4337
R17899 vdd.n2982 vdd.n2981 52.4337
R17900 vdd.n372 vdd.n371 52.4337
R17901 vdd.n367 vdd.n360 52.4337
R17902 vdd.n2993 vdd.n2992 52.4337
R17903 vdd.n359 vdd.n353 52.4337
R17904 vdd.n3000 vdd.n2999 52.4337
R17905 vdd.n352 vdd.n346 52.4337
R17906 vdd.n3007 vdd.n3006 52.4337
R17907 vdd.n345 vdd.n338 52.4337
R17908 vdd.n3014 vdd.n3013 52.4337
R17909 vdd.n3017 vdd.n3016 52.4337
R17910 vdd.n333 vdd.n330 52.4337
R17911 vdd.t181 vdd.t79 51.4683
R17912 vdd.n250 vdd.n248 42.0461
R17913 vdd.n160 vdd.n158 42.0461
R17914 vdd.n71 vdd.n69 42.0461
R17915 vdd.n1112 vdd.n1110 42.0461
R17916 vdd.n1022 vdd.n1020 42.0461
R17917 vdd.n933 vdd.n931 42.0461
R17918 vdd.n296 vdd.n295 41.6884
R17919 vdd.n206 vdd.n205 41.6884
R17920 vdd.n117 vdd.n116 41.6884
R17921 vdd.n1158 vdd.n1157 41.6884
R17922 vdd.n1068 vdd.n1067 41.6884
R17923 vdd.n979 vdd.n978 41.6884
R17924 vdd.n1322 vdd.n1321 41.1157
R17925 vdd.n1360 vdd.n1359 41.1157
R17926 vdd.n1256 vdd.n1255 41.1157
R17927 vdd.n2910 vdd.n2909 41.1157
R17928 vdd.n2949 vdd.n406 41.1157
R17929 vdd.n2988 vdd.n366 41.1157
R17930 vdd.n2667 vdd.n2666 39.2114
R17931 vdd.n2664 vdd.n2663 39.2114
R17932 vdd.n2659 vdd.n605 39.2114
R17933 vdd.n2657 vdd.n2656 39.2114
R17934 vdd.n2652 vdd.n608 39.2114
R17935 vdd.n2650 vdd.n2649 39.2114
R17936 vdd.n2645 vdd.n611 39.2114
R17937 vdd.n2643 vdd.n2642 39.2114
R17938 vdd.n2639 vdd.n2638 39.2114
R17939 vdd.n2634 vdd.n614 39.2114
R17940 vdd.n2632 vdd.n2631 39.2114
R17941 vdd.n2627 vdd.n617 39.2114
R17942 vdd.n2625 vdd.n2624 39.2114
R17943 vdd.n2620 vdd.n620 39.2114
R17944 vdd.n2618 vdd.n2617 39.2114
R17945 vdd.n2612 vdd.n625 39.2114
R17946 vdd.n2610 vdd.n2609 39.2114
R17947 vdd.n2470 vdd.n703 39.2114
R17948 vdd.n2465 vdd.n2219 39.2114
R17949 vdd.n2462 vdd.n2220 39.2114
R17950 vdd.n2458 vdd.n2221 39.2114
R17951 vdd.n2454 vdd.n2222 39.2114
R17952 vdd.n2450 vdd.n2223 39.2114
R17953 vdd.n2446 vdd.n2224 39.2114
R17954 vdd.n2442 vdd.n2225 39.2114
R17955 vdd.n2438 vdd.n2226 39.2114
R17956 vdd.n2434 vdd.n2227 39.2114
R17957 vdd.n2430 vdd.n2228 39.2114
R17958 vdd.n2426 vdd.n2229 39.2114
R17959 vdd.n2422 vdd.n2230 39.2114
R17960 vdd.n2418 vdd.n2231 39.2114
R17961 vdd.n2414 vdd.n2232 39.2114
R17962 vdd.n2410 vdd.n2233 39.2114
R17963 vdd.n2405 vdd.n2234 39.2114
R17964 vdd.n2213 vdd.n743 39.2114
R17965 vdd.n2209 vdd.n742 39.2114
R17966 vdd.n2205 vdd.n741 39.2114
R17967 vdd.n2201 vdd.n740 39.2114
R17968 vdd.n2197 vdd.n739 39.2114
R17969 vdd.n2193 vdd.n738 39.2114
R17970 vdd.n2189 vdd.n737 39.2114
R17971 vdd.n2185 vdd.n736 39.2114
R17972 vdd.n2181 vdd.n735 39.2114
R17973 vdd.n2177 vdd.n734 39.2114
R17974 vdd.n2173 vdd.n733 39.2114
R17975 vdd.n2169 vdd.n732 39.2114
R17976 vdd.n2165 vdd.n731 39.2114
R17977 vdd.n2161 vdd.n730 39.2114
R17978 vdd.n2157 vdd.n729 39.2114
R17979 vdd.n2152 vdd.n728 39.2114
R17980 vdd.n2148 vdd.n727 39.2114
R17981 vdd.n1724 vdd.n838 39.2114
R17982 vdd.n1730 vdd.n1729 39.2114
R17983 vdd.n1733 vdd.n1732 39.2114
R17984 vdd.n1738 vdd.n1737 39.2114
R17985 vdd.n1741 vdd.n1740 39.2114
R17986 vdd.n1746 vdd.n1745 39.2114
R17987 vdd.n1749 vdd.n1748 39.2114
R17988 vdd.n1754 vdd.n1753 39.2114
R17989 vdd.n1925 vdd.n1756 39.2114
R17990 vdd.n1924 vdd.n1923 39.2114
R17991 vdd.n1917 vdd.n1758 39.2114
R17992 vdd.n1916 vdd.n1915 39.2114
R17993 vdd.n1909 vdd.n1760 39.2114
R17994 vdd.n1908 vdd.n1907 39.2114
R17995 vdd.n1901 vdd.n1762 39.2114
R17996 vdd.n1900 vdd.n1899 39.2114
R17997 vdd.n1893 vdd.n1764 39.2114
R17998 vdd.n2586 vdd.n2585 39.2114
R17999 vdd.n2581 vdd.n2553 39.2114
R18000 vdd.n2579 vdd.n2578 39.2114
R18001 vdd.n2574 vdd.n2556 39.2114
R18002 vdd.n2572 vdd.n2571 39.2114
R18003 vdd.n2567 vdd.n2559 39.2114
R18004 vdd.n2565 vdd.n2564 39.2114
R18005 vdd.n2560 vdd.n577 39.2114
R18006 vdd.n2704 vdd.n2703 39.2114
R18007 vdd.n2701 vdd.n2700 39.2114
R18008 vdd.n2696 vdd.n581 39.2114
R18009 vdd.n2694 vdd.n2693 39.2114
R18010 vdd.n2689 vdd.n584 39.2114
R18011 vdd.n2687 vdd.n2686 39.2114
R18012 vdd.n2682 vdd.n587 39.2114
R18013 vdd.n2680 vdd.n2679 39.2114
R18014 vdd.n2675 vdd.n593 39.2114
R18015 vdd.n2472 vdd.n706 39.2114
R18016 vdd.n2235 vdd.n708 39.2114
R18017 vdd.n2261 vdd.n2236 39.2114
R18018 vdd.n2265 vdd.n2237 39.2114
R18019 vdd.n2269 vdd.n2238 39.2114
R18020 vdd.n2273 vdd.n2239 39.2114
R18021 vdd.n2277 vdd.n2240 39.2114
R18022 vdd.n2281 vdd.n2241 39.2114
R18023 vdd.n2285 vdd.n2242 39.2114
R18024 vdd.n2289 vdd.n2243 39.2114
R18025 vdd.n2293 vdd.n2244 39.2114
R18026 vdd.n2297 vdd.n2245 39.2114
R18027 vdd.n2301 vdd.n2246 39.2114
R18028 vdd.n2305 vdd.n2247 39.2114
R18029 vdd.n2309 vdd.n2248 39.2114
R18030 vdd.n2313 vdd.n2249 39.2114
R18031 vdd.n2317 vdd.n2250 39.2114
R18032 vdd.n2473 vdd.n2472 39.2114
R18033 vdd.n2260 vdd.n2235 39.2114
R18034 vdd.n2264 vdd.n2236 39.2114
R18035 vdd.n2268 vdd.n2237 39.2114
R18036 vdd.n2272 vdd.n2238 39.2114
R18037 vdd.n2276 vdd.n2239 39.2114
R18038 vdd.n2280 vdd.n2240 39.2114
R18039 vdd.n2284 vdd.n2241 39.2114
R18040 vdd.n2288 vdd.n2242 39.2114
R18041 vdd.n2292 vdd.n2243 39.2114
R18042 vdd.n2296 vdd.n2244 39.2114
R18043 vdd.n2300 vdd.n2245 39.2114
R18044 vdd.n2304 vdd.n2246 39.2114
R18045 vdd.n2308 vdd.n2247 39.2114
R18046 vdd.n2312 vdd.n2248 39.2114
R18047 vdd.n2316 vdd.n2249 39.2114
R18048 vdd.n2319 vdd.n2250 39.2114
R18049 vdd.n593 vdd.n588 39.2114
R18050 vdd.n2681 vdd.n2680 39.2114
R18051 vdd.n587 vdd.n585 39.2114
R18052 vdd.n2688 vdd.n2687 39.2114
R18053 vdd.n584 vdd.n582 39.2114
R18054 vdd.n2695 vdd.n2694 39.2114
R18055 vdd.n581 vdd.n579 39.2114
R18056 vdd.n2702 vdd.n2701 39.2114
R18057 vdd.n2705 vdd.n2704 39.2114
R18058 vdd.n2561 vdd.n2560 39.2114
R18059 vdd.n2566 vdd.n2565 39.2114
R18060 vdd.n2559 vdd.n2557 39.2114
R18061 vdd.n2573 vdd.n2572 39.2114
R18062 vdd.n2556 vdd.n2554 39.2114
R18063 vdd.n2580 vdd.n2579 39.2114
R18064 vdd.n2553 vdd.n2551 39.2114
R18065 vdd.n2587 vdd.n2586 39.2114
R18066 vdd.n1725 vdd.n1724 39.2114
R18067 vdd.n1731 vdd.n1730 39.2114
R18068 vdd.n1732 vdd.n1721 39.2114
R18069 vdd.n1739 vdd.n1738 39.2114
R18070 vdd.n1740 vdd.n1719 39.2114
R18071 vdd.n1747 vdd.n1746 39.2114
R18072 vdd.n1748 vdd.n1717 39.2114
R18073 vdd.n1755 vdd.n1754 39.2114
R18074 vdd.n1926 vdd.n1925 39.2114
R18075 vdd.n1923 vdd.n1922 39.2114
R18076 vdd.n1918 vdd.n1917 39.2114
R18077 vdd.n1915 vdd.n1914 39.2114
R18078 vdd.n1910 vdd.n1909 39.2114
R18079 vdd.n1907 vdd.n1906 39.2114
R18080 vdd.n1902 vdd.n1901 39.2114
R18081 vdd.n1899 vdd.n1898 39.2114
R18082 vdd.n1894 vdd.n1893 39.2114
R18083 vdd.n2151 vdd.n727 39.2114
R18084 vdd.n2156 vdd.n728 39.2114
R18085 vdd.n2160 vdd.n729 39.2114
R18086 vdd.n2164 vdd.n730 39.2114
R18087 vdd.n2168 vdd.n731 39.2114
R18088 vdd.n2172 vdd.n732 39.2114
R18089 vdd.n2176 vdd.n733 39.2114
R18090 vdd.n2180 vdd.n734 39.2114
R18091 vdd.n2184 vdd.n735 39.2114
R18092 vdd.n2188 vdd.n736 39.2114
R18093 vdd.n2192 vdd.n737 39.2114
R18094 vdd.n2196 vdd.n738 39.2114
R18095 vdd.n2200 vdd.n739 39.2114
R18096 vdd.n2204 vdd.n740 39.2114
R18097 vdd.n2208 vdd.n741 39.2114
R18098 vdd.n2212 vdd.n742 39.2114
R18099 vdd.n745 vdd.n743 39.2114
R18100 vdd.n2470 vdd.n2469 39.2114
R18101 vdd.n2463 vdd.n2219 39.2114
R18102 vdd.n2459 vdd.n2220 39.2114
R18103 vdd.n2455 vdd.n2221 39.2114
R18104 vdd.n2451 vdd.n2222 39.2114
R18105 vdd.n2447 vdd.n2223 39.2114
R18106 vdd.n2443 vdd.n2224 39.2114
R18107 vdd.n2439 vdd.n2225 39.2114
R18108 vdd.n2435 vdd.n2226 39.2114
R18109 vdd.n2431 vdd.n2227 39.2114
R18110 vdd.n2427 vdd.n2228 39.2114
R18111 vdd.n2423 vdd.n2229 39.2114
R18112 vdd.n2419 vdd.n2230 39.2114
R18113 vdd.n2415 vdd.n2231 39.2114
R18114 vdd.n2411 vdd.n2232 39.2114
R18115 vdd.n2406 vdd.n2233 39.2114
R18116 vdd.n2402 vdd.n2234 39.2114
R18117 vdd.n2611 vdd.n2610 39.2114
R18118 vdd.n625 vdd.n621 39.2114
R18119 vdd.n2619 vdd.n2618 39.2114
R18120 vdd.n620 vdd.n618 39.2114
R18121 vdd.n2626 vdd.n2625 39.2114
R18122 vdd.n617 vdd.n615 39.2114
R18123 vdd.n2633 vdd.n2632 39.2114
R18124 vdd.n614 vdd.n612 39.2114
R18125 vdd.n2640 vdd.n2639 39.2114
R18126 vdd.n2644 vdd.n2643 39.2114
R18127 vdd.n611 vdd.n609 39.2114
R18128 vdd.n2651 vdd.n2650 39.2114
R18129 vdd.n608 vdd.n606 39.2114
R18130 vdd.n2658 vdd.n2657 39.2114
R18131 vdd.n605 vdd.n603 39.2114
R18132 vdd.n2665 vdd.n2664 39.2114
R18133 vdd.n2668 vdd.n2667 39.2114
R18134 vdd.n753 vdd.n709 39.2114
R18135 vdd.n2140 vdd.n710 39.2114
R18136 vdd.n2136 vdd.n711 39.2114
R18137 vdd.n2132 vdd.n712 39.2114
R18138 vdd.n2128 vdd.n713 39.2114
R18139 vdd.n2124 vdd.n714 39.2114
R18140 vdd.n2120 vdd.n715 39.2114
R18141 vdd.n2116 vdd.n716 39.2114
R18142 vdd.n2112 vdd.n717 39.2114
R18143 vdd.n2108 vdd.n718 39.2114
R18144 vdd.n2104 vdd.n719 39.2114
R18145 vdd.n2100 vdd.n720 39.2114
R18146 vdd.n2096 vdd.n721 39.2114
R18147 vdd.n2092 vdd.n722 39.2114
R18148 vdd.n2088 vdd.n723 39.2114
R18149 vdd.n2084 vdd.n724 39.2114
R18150 vdd.n2080 vdd.n725 39.2114
R18151 vdd.n1983 vdd.n842 39.2114
R18152 vdd.n1982 vdd.n1981 39.2114
R18153 vdd.n1975 vdd.n844 39.2114
R18154 vdd.n1974 vdd.n1973 39.2114
R18155 vdd.n1967 vdd.n846 39.2114
R18156 vdd.n1966 vdd.n1965 39.2114
R18157 vdd.n1959 vdd.n848 39.2114
R18158 vdd.n1958 vdd.n1957 39.2114
R18159 vdd.n851 vdd.n850 39.2114
R18160 vdd.n1799 vdd.n1798 39.2114
R18161 vdd.n1804 vdd.n1803 39.2114
R18162 vdd.n1807 vdd.n1806 39.2114
R18163 vdd.n1812 vdd.n1811 39.2114
R18164 vdd.n1815 vdd.n1814 39.2114
R18165 vdd.n1820 vdd.n1819 39.2114
R18166 vdd.n1823 vdd.n1822 39.2114
R18167 vdd.n1829 vdd.n1828 39.2114
R18168 vdd.n2077 vdd.n725 39.2114
R18169 vdd.n2081 vdd.n724 39.2114
R18170 vdd.n2085 vdd.n723 39.2114
R18171 vdd.n2089 vdd.n722 39.2114
R18172 vdd.n2093 vdd.n721 39.2114
R18173 vdd.n2097 vdd.n720 39.2114
R18174 vdd.n2101 vdd.n719 39.2114
R18175 vdd.n2105 vdd.n718 39.2114
R18176 vdd.n2109 vdd.n717 39.2114
R18177 vdd.n2113 vdd.n716 39.2114
R18178 vdd.n2117 vdd.n715 39.2114
R18179 vdd.n2121 vdd.n714 39.2114
R18180 vdd.n2125 vdd.n713 39.2114
R18181 vdd.n2129 vdd.n712 39.2114
R18182 vdd.n2133 vdd.n711 39.2114
R18183 vdd.n2137 vdd.n710 39.2114
R18184 vdd.n2141 vdd.n709 39.2114
R18185 vdd.n1984 vdd.n1983 39.2114
R18186 vdd.n1981 vdd.n1980 39.2114
R18187 vdd.n1976 vdd.n1975 39.2114
R18188 vdd.n1973 vdd.n1972 39.2114
R18189 vdd.n1968 vdd.n1967 39.2114
R18190 vdd.n1965 vdd.n1964 39.2114
R18191 vdd.n1960 vdd.n1959 39.2114
R18192 vdd.n1957 vdd.n1956 39.2114
R18193 vdd.n852 vdd.n851 39.2114
R18194 vdd.n1800 vdd.n1799 39.2114
R18195 vdd.n1805 vdd.n1804 39.2114
R18196 vdd.n1806 vdd.n1796 39.2114
R18197 vdd.n1813 vdd.n1812 39.2114
R18198 vdd.n1814 vdd.n1794 39.2114
R18199 vdd.n1821 vdd.n1820 39.2114
R18200 vdd.n1822 vdd.n1790 39.2114
R18201 vdd.n1830 vdd.n1829 39.2114
R18202 vdd.n1949 vdd.n1948 37.2369
R18203 vdd.n1652 vdd.n1585 37.2369
R18204 vdd.n1691 vdd.n1545 37.2369
R18205 vdd.n2758 vdd.n558 37.2369
R18206 vdd.n2806 vdd.n2805 37.2369
R18207 vdd.n2713 vdd.n2712 37.2369
R18208 vdd.n1991 vdd.n837 31.6883
R18209 vdd.n2216 vdd.n746 31.6883
R18210 vdd.n2149 vdd.n749 31.6883
R18211 vdd.n1895 vdd.n1892 31.6883
R18212 vdd.n2403 vdd.n2401 31.6883
R18213 vdd.n2608 vdd.n2607 31.6883
R18214 vdd.n2480 vdd.n702 31.6883
R18215 vdd.n2671 vdd.n2670 31.6883
R18216 vdd.n2590 vdd.n2589 31.6883
R18217 vdd.n2676 vdd.n592 31.6883
R18218 vdd.n2322 vdd.n2321 31.6883
R18219 vdd.n2476 vdd.n2475 31.6883
R18220 vdd.n1987 vdd.n1986 31.6883
R18221 vdd.n2144 vdd.n2143 31.6883
R18222 vdd.n2076 vdd.n2075 31.6883
R18223 vdd.n1833 vdd.n1832 31.6883
R18224 vdd.n1826 vdd.n1792 30.449
R18225 vdd.n757 vdd.n756 30.449
R18226 vdd.n1767 vdd.n1766 30.449
R18227 vdd.n2154 vdd.n748 30.449
R18228 vdd.n2258 vdd.n2257 30.449
R18229 vdd.n2614 vdd.n623 30.449
R18230 vdd.n2408 vdd.n2254 30.449
R18231 vdd.n591 vdd.n590 30.449
R18232 vdd.n1421 vdd.n1228 22.6735
R18233 vdd.n1943 vdd.n863 22.6735
R18234 vdd.n2840 vdd.n516 22.6735
R18235 vdd.n3025 vdd.n329 22.6735
R18236 vdd.n1432 vdd.n1190 19.3944
R18237 vdd.n1432 vdd.n1188 19.3944
R18238 vdd.n1436 vdd.n1188 19.3944
R18239 vdd.n1436 vdd.n1178 19.3944
R18240 vdd.n1449 vdd.n1178 19.3944
R18241 vdd.n1449 vdd.n1176 19.3944
R18242 vdd.n1453 vdd.n1176 19.3944
R18243 vdd.n1453 vdd.n1168 19.3944
R18244 vdd.n1467 vdd.n1168 19.3944
R18245 vdd.n1467 vdd.n1166 19.3944
R18246 vdd.n1471 vdd.n1166 19.3944
R18247 vdd.n1471 vdd.n885 19.3944
R18248 vdd.n1483 vdd.n885 19.3944
R18249 vdd.n1483 vdd.n883 19.3944
R18250 vdd.n1487 vdd.n883 19.3944
R18251 vdd.n1487 vdd.n875 19.3944
R18252 vdd.n1500 vdd.n875 19.3944
R18253 vdd.n1500 vdd.n872 19.3944
R18254 vdd.n1506 vdd.n872 19.3944
R18255 vdd.n1506 vdd.n873 19.3944
R18256 vdd.n873 vdd.n862 19.3944
R18257 vdd.n1356 vdd.n1291 19.3944
R18258 vdd.n1352 vdd.n1291 19.3944
R18259 vdd.n1352 vdd.n1351 19.3944
R18260 vdd.n1351 vdd.n1350 19.3944
R18261 vdd.n1350 vdd.n1297 19.3944
R18262 vdd.n1346 vdd.n1297 19.3944
R18263 vdd.n1346 vdd.n1345 19.3944
R18264 vdd.n1345 vdd.n1344 19.3944
R18265 vdd.n1344 vdd.n1303 19.3944
R18266 vdd.n1340 vdd.n1303 19.3944
R18267 vdd.n1340 vdd.n1339 19.3944
R18268 vdd.n1339 vdd.n1338 19.3944
R18269 vdd.n1338 vdd.n1309 19.3944
R18270 vdd.n1334 vdd.n1309 19.3944
R18271 vdd.n1334 vdd.n1333 19.3944
R18272 vdd.n1333 vdd.n1332 19.3944
R18273 vdd.n1332 vdd.n1315 19.3944
R18274 vdd.n1328 vdd.n1315 19.3944
R18275 vdd.n1328 vdd.n1327 19.3944
R18276 vdd.n1327 vdd.n1326 19.3944
R18277 vdd.n1391 vdd.n1390 19.3944
R18278 vdd.n1390 vdd.n1389 19.3944
R18279 vdd.n1389 vdd.n1262 19.3944
R18280 vdd.n1385 vdd.n1262 19.3944
R18281 vdd.n1385 vdd.n1384 19.3944
R18282 vdd.n1384 vdd.n1383 19.3944
R18283 vdd.n1383 vdd.n1268 19.3944
R18284 vdd.n1379 vdd.n1268 19.3944
R18285 vdd.n1379 vdd.n1378 19.3944
R18286 vdd.n1378 vdd.n1377 19.3944
R18287 vdd.n1377 vdd.n1274 19.3944
R18288 vdd.n1373 vdd.n1274 19.3944
R18289 vdd.n1373 vdd.n1372 19.3944
R18290 vdd.n1372 vdd.n1371 19.3944
R18291 vdd.n1371 vdd.n1280 19.3944
R18292 vdd.n1367 vdd.n1280 19.3944
R18293 vdd.n1367 vdd.n1366 19.3944
R18294 vdd.n1366 vdd.n1365 19.3944
R18295 vdd.n1365 vdd.n1286 19.3944
R18296 vdd.n1361 vdd.n1286 19.3944
R18297 vdd.n1424 vdd.n1195 19.3944
R18298 vdd.n1419 vdd.n1195 19.3944
R18299 vdd.n1419 vdd.n1230 19.3944
R18300 vdd.n1415 vdd.n1230 19.3944
R18301 vdd.n1415 vdd.n1414 19.3944
R18302 vdd.n1414 vdd.n1413 19.3944
R18303 vdd.n1413 vdd.n1236 19.3944
R18304 vdd.n1409 vdd.n1236 19.3944
R18305 vdd.n1409 vdd.n1408 19.3944
R18306 vdd.n1408 vdd.n1407 19.3944
R18307 vdd.n1407 vdd.n1242 19.3944
R18308 vdd.n1403 vdd.n1242 19.3944
R18309 vdd.n1403 vdd.n1402 19.3944
R18310 vdd.n1402 vdd.n1401 19.3944
R18311 vdd.n1401 vdd.n1248 19.3944
R18312 vdd.n1397 vdd.n1248 19.3944
R18313 vdd.n1397 vdd.n1396 19.3944
R18314 vdd.n1396 vdd.n1395 19.3944
R18315 vdd.n1648 vdd.n1583 19.3944
R18316 vdd.n1648 vdd.n1589 19.3944
R18317 vdd.n1643 vdd.n1589 19.3944
R18318 vdd.n1643 vdd.n1642 19.3944
R18319 vdd.n1642 vdd.n1641 19.3944
R18320 vdd.n1641 vdd.n1596 19.3944
R18321 vdd.n1636 vdd.n1596 19.3944
R18322 vdd.n1636 vdd.n1635 19.3944
R18323 vdd.n1635 vdd.n1634 19.3944
R18324 vdd.n1634 vdd.n1603 19.3944
R18325 vdd.n1629 vdd.n1603 19.3944
R18326 vdd.n1629 vdd.n1628 19.3944
R18327 vdd.n1628 vdd.n1627 19.3944
R18328 vdd.n1627 vdd.n1611 19.3944
R18329 vdd.n1622 vdd.n1611 19.3944
R18330 vdd.n1622 vdd.n1621 19.3944
R18331 vdd.n1617 vdd.n1616 19.3944
R18332 vdd.n1950 vdd.n858 19.3944
R18333 vdd.n1687 vdd.n1543 19.3944
R18334 vdd.n1687 vdd.n1549 19.3944
R18335 vdd.n1682 vdd.n1549 19.3944
R18336 vdd.n1682 vdd.n1681 19.3944
R18337 vdd.n1681 vdd.n1680 19.3944
R18338 vdd.n1680 vdd.n1556 19.3944
R18339 vdd.n1675 vdd.n1556 19.3944
R18340 vdd.n1675 vdd.n1674 19.3944
R18341 vdd.n1674 vdd.n1673 19.3944
R18342 vdd.n1673 vdd.n1563 19.3944
R18343 vdd.n1668 vdd.n1563 19.3944
R18344 vdd.n1668 vdd.n1667 19.3944
R18345 vdd.n1667 vdd.n1666 19.3944
R18346 vdd.n1666 vdd.n1570 19.3944
R18347 vdd.n1661 vdd.n1570 19.3944
R18348 vdd.n1661 vdd.n1660 19.3944
R18349 vdd.n1660 vdd.n1659 19.3944
R18350 vdd.n1659 vdd.n1577 19.3944
R18351 vdd.n1654 vdd.n1577 19.3944
R18352 vdd.n1654 vdd.n1653 19.3944
R18353 vdd.n1938 vdd.n1937 19.3944
R18354 vdd.n1937 vdd.n1515 19.3944
R18355 vdd.n1932 vdd.n1931 19.3944
R18356 vdd.n1714 vdd.n1519 19.3944
R18357 vdd.n1714 vdd.n1521 19.3944
R18358 vdd.n1524 vdd.n1521 19.3944
R18359 vdd.n1707 vdd.n1524 19.3944
R18360 vdd.n1707 vdd.n1706 19.3944
R18361 vdd.n1706 vdd.n1705 19.3944
R18362 vdd.n1705 vdd.n1530 19.3944
R18363 vdd.n1700 vdd.n1530 19.3944
R18364 vdd.n1700 vdd.n1699 19.3944
R18365 vdd.n1699 vdd.n1698 19.3944
R18366 vdd.n1698 vdd.n1537 19.3944
R18367 vdd.n1693 vdd.n1537 19.3944
R18368 vdd.n1693 vdd.n1692 19.3944
R18369 vdd.n1428 vdd.n1193 19.3944
R18370 vdd.n1428 vdd.n1184 19.3944
R18371 vdd.n1441 vdd.n1184 19.3944
R18372 vdd.n1441 vdd.n1182 19.3944
R18373 vdd.n1445 vdd.n1182 19.3944
R18374 vdd.n1445 vdd.n1173 19.3944
R18375 vdd.n1458 vdd.n1173 19.3944
R18376 vdd.n1458 vdd.n1171 19.3944
R18377 vdd.n1463 vdd.n1171 19.3944
R18378 vdd.n1463 vdd.n1162 19.3944
R18379 vdd.n1475 vdd.n1162 19.3944
R18380 vdd.n1475 vdd.n890 19.3944
R18381 vdd.n1479 vdd.n890 19.3944
R18382 vdd.n1479 vdd.n880 19.3944
R18383 vdd.n1492 vdd.n880 19.3944
R18384 vdd.n1492 vdd.n878 19.3944
R18385 vdd.n1496 vdd.n878 19.3944
R18386 vdd.n1496 vdd.n868 19.3944
R18387 vdd.n1511 vdd.n868 19.3944
R18388 vdd.n1511 vdd.n866 19.3944
R18389 vdd.n1941 vdd.n866 19.3944
R18390 vdd.n2851 vdd.n477 19.3944
R18391 vdd.n2851 vdd.n475 19.3944
R18392 vdd.n2855 vdd.n475 19.3944
R18393 vdd.n2855 vdd.n465 19.3944
R18394 vdd.n2868 vdd.n465 19.3944
R18395 vdd.n2868 vdd.n463 19.3944
R18396 vdd.n2872 vdd.n463 19.3944
R18397 vdd.n2872 vdd.n453 19.3944
R18398 vdd.n2884 vdd.n453 19.3944
R18399 vdd.n2884 vdd.n451 19.3944
R18400 vdd.n2888 vdd.n451 19.3944
R18401 vdd.n2889 vdd.n2888 19.3944
R18402 vdd.n2890 vdd.n2889 19.3944
R18403 vdd.n2890 vdd.n449 19.3944
R18404 vdd.n2894 vdd.n449 19.3944
R18405 vdd.n2895 vdd.n2894 19.3944
R18406 vdd.n2896 vdd.n2895 19.3944
R18407 vdd.n2896 vdd.n446 19.3944
R18408 vdd.n2900 vdd.n446 19.3944
R18409 vdd.n2901 vdd.n2900 19.3944
R18410 vdd.n2902 vdd.n2901 19.3944
R18411 vdd.n2945 vdd.n404 19.3944
R18412 vdd.n2945 vdd.n410 19.3944
R18413 vdd.n2940 vdd.n410 19.3944
R18414 vdd.n2940 vdd.n2939 19.3944
R18415 vdd.n2939 vdd.n2938 19.3944
R18416 vdd.n2938 vdd.n417 19.3944
R18417 vdd.n2933 vdd.n417 19.3944
R18418 vdd.n2933 vdd.n2932 19.3944
R18419 vdd.n2932 vdd.n2931 19.3944
R18420 vdd.n2931 vdd.n424 19.3944
R18421 vdd.n2926 vdd.n424 19.3944
R18422 vdd.n2926 vdd.n2925 19.3944
R18423 vdd.n2925 vdd.n2924 19.3944
R18424 vdd.n2924 vdd.n431 19.3944
R18425 vdd.n2919 vdd.n431 19.3944
R18426 vdd.n2919 vdd.n2918 19.3944
R18427 vdd.n2918 vdd.n2917 19.3944
R18428 vdd.n2917 vdd.n438 19.3944
R18429 vdd.n2912 vdd.n438 19.3944
R18430 vdd.n2912 vdd.n2911 19.3944
R18431 vdd.n2984 vdd.n364 19.3944
R18432 vdd.n2984 vdd.n370 19.3944
R18433 vdd.n2979 vdd.n370 19.3944
R18434 vdd.n2979 vdd.n2978 19.3944
R18435 vdd.n2978 vdd.n2977 19.3944
R18436 vdd.n2977 vdd.n377 19.3944
R18437 vdd.n2972 vdd.n377 19.3944
R18438 vdd.n2972 vdd.n2971 19.3944
R18439 vdd.n2971 vdd.n2970 19.3944
R18440 vdd.n2970 vdd.n384 19.3944
R18441 vdd.n2965 vdd.n384 19.3944
R18442 vdd.n2965 vdd.n2964 19.3944
R18443 vdd.n2964 vdd.n2963 19.3944
R18444 vdd.n2963 vdd.n391 19.3944
R18445 vdd.n2958 vdd.n391 19.3944
R18446 vdd.n2958 vdd.n2957 19.3944
R18447 vdd.n2957 vdd.n2956 19.3944
R18448 vdd.n2956 vdd.n398 19.3944
R18449 vdd.n2951 vdd.n398 19.3944
R18450 vdd.n2951 vdd.n2950 19.3944
R18451 vdd.n3020 vdd.n3019 19.3944
R18452 vdd.n3019 vdd.n3018 19.3944
R18453 vdd.n3018 vdd.n336 19.3944
R18454 vdd.n337 vdd.n336 19.3944
R18455 vdd.n3011 vdd.n337 19.3944
R18456 vdd.n3011 vdd.n3010 19.3944
R18457 vdd.n3010 vdd.n3009 19.3944
R18458 vdd.n3009 vdd.n344 19.3944
R18459 vdd.n3004 vdd.n344 19.3944
R18460 vdd.n3004 vdd.n3003 19.3944
R18461 vdd.n3003 vdd.n3002 19.3944
R18462 vdd.n3002 vdd.n351 19.3944
R18463 vdd.n2997 vdd.n351 19.3944
R18464 vdd.n2997 vdd.n2996 19.3944
R18465 vdd.n2996 vdd.n2995 19.3944
R18466 vdd.n2995 vdd.n358 19.3944
R18467 vdd.n2990 vdd.n358 19.3944
R18468 vdd.n2990 vdd.n2989 19.3944
R18469 vdd.n2847 vdd.n480 19.3944
R18470 vdd.n2847 vdd.n471 19.3944
R18471 vdd.n2860 vdd.n471 19.3944
R18472 vdd.n2860 vdd.n469 19.3944
R18473 vdd.n2864 vdd.n469 19.3944
R18474 vdd.n2864 vdd.n460 19.3944
R18475 vdd.n2876 vdd.n460 19.3944
R18476 vdd.n2876 vdd.n458 19.3944
R18477 vdd.n2880 vdd.n458 19.3944
R18478 vdd.n2880 vdd.n300 19.3944
R18479 vdd.n3045 vdd.n300 19.3944
R18480 vdd.n3045 vdd.n301 19.3944
R18481 vdd.n3039 vdd.n301 19.3944
R18482 vdd.n3039 vdd.n3038 19.3944
R18483 vdd.n3038 vdd.n3037 19.3944
R18484 vdd.n3037 vdd.n313 19.3944
R18485 vdd.n3031 vdd.n313 19.3944
R18486 vdd.n3031 vdd.n3030 19.3944
R18487 vdd.n3030 vdd.n3029 19.3944
R18488 vdd.n3029 vdd.n324 19.3944
R18489 vdd.n3023 vdd.n324 19.3944
R18490 vdd.n2800 vdd.n536 19.3944
R18491 vdd.n2800 vdd.n2797 19.3944
R18492 vdd.n2797 vdd.n2794 19.3944
R18493 vdd.n2794 vdd.n2793 19.3944
R18494 vdd.n2793 vdd.n2790 19.3944
R18495 vdd.n2790 vdd.n2789 19.3944
R18496 vdd.n2789 vdd.n2786 19.3944
R18497 vdd.n2786 vdd.n2785 19.3944
R18498 vdd.n2785 vdd.n2782 19.3944
R18499 vdd.n2782 vdd.n2781 19.3944
R18500 vdd.n2781 vdd.n2778 19.3944
R18501 vdd.n2778 vdd.n2777 19.3944
R18502 vdd.n2777 vdd.n2774 19.3944
R18503 vdd.n2774 vdd.n2773 19.3944
R18504 vdd.n2773 vdd.n2770 19.3944
R18505 vdd.n2770 vdd.n2769 19.3944
R18506 vdd.n2769 vdd.n2766 19.3944
R18507 vdd.n2766 vdd.n2765 19.3944
R18508 vdd.n2765 vdd.n2762 19.3944
R18509 vdd.n2762 vdd.n2761 19.3944
R18510 vdd.n2843 vdd.n482 19.3944
R18511 vdd.n2838 vdd.n482 19.3944
R18512 vdd.n521 vdd.n518 19.3944
R18513 vdd.n2834 vdd.n2833 19.3944
R18514 vdd.n2833 vdd.n2830 19.3944
R18515 vdd.n2830 vdd.n2829 19.3944
R18516 vdd.n2829 vdd.n2826 19.3944
R18517 vdd.n2826 vdd.n2825 19.3944
R18518 vdd.n2825 vdd.n2822 19.3944
R18519 vdd.n2822 vdd.n2821 19.3944
R18520 vdd.n2821 vdd.n2818 19.3944
R18521 vdd.n2818 vdd.n2817 19.3944
R18522 vdd.n2817 vdd.n2814 19.3944
R18523 vdd.n2814 vdd.n2813 19.3944
R18524 vdd.n2813 vdd.n2810 19.3944
R18525 vdd.n2810 vdd.n2809 19.3944
R18526 vdd.n2754 vdd.n556 19.3944
R18527 vdd.n2754 vdd.n2751 19.3944
R18528 vdd.n2751 vdd.n2748 19.3944
R18529 vdd.n2748 vdd.n2747 19.3944
R18530 vdd.n2747 vdd.n2744 19.3944
R18531 vdd.n2744 vdd.n2743 19.3944
R18532 vdd.n2743 vdd.n2740 19.3944
R18533 vdd.n2740 vdd.n2739 19.3944
R18534 vdd.n2739 vdd.n2736 19.3944
R18535 vdd.n2736 vdd.n2735 19.3944
R18536 vdd.n2735 vdd.n2732 19.3944
R18537 vdd.n2732 vdd.n2731 19.3944
R18538 vdd.n2731 vdd.n2728 19.3944
R18539 vdd.n2728 vdd.n2727 19.3944
R18540 vdd.n2727 vdd.n2724 19.3944
R18541 vdd.n2724 vdd.n2723 19.3944
R18542 vdd.n2720 vdd.n2719 19.3944
R18543 vdd.n2716 vdd.n2715 19.3944
R18544 vdd.n1360 vdd.n1356 19.0066
R18545 vdd.n1652 vdd.n1583 19.0066
R18546 vdd.n2949 vdd.n404 19.0066
R18547 vdd.n2758 vdd.n556 19.0066
R18548 vdd.n1792 vdd.n1791 16.0975
R18549 vdd.n756 vdd.n755 16.0975
R18550 vdd.n1321 vdd.n1320 16.0975
R18551 vdd.n1359 vdd.n1358 16.0975
R18552 vdd.n1255 vdd.n1254 16.0975
R18553 vdd.n1948 vdd.n1947 16.0975
R18554 vdd.n1585 vdd.n1584 16.0975
R18555 vdd.n1545 vdd.n1544 16.0975
R18556 vdd.n1766 vdd.n1765 16.0975
R18557 vdd.n748 vdd.n747 16.0975
R18558 vdd.n2257 vdd.n2256 16.0975
R18559 vdd.n2909 vdd.n2908 16.0975
R18560 vdd.n406 vdd.n405 16.0975
R18561 vdd.n366 vdd.n365 16.0975
R18562 vdd.n558 vdd.n557 16.0975
R18563 vdd.n2805 vdd.n2804 16.0975
R18564 vdd.n623 vdd.n622 16.0975
R18565 vdd.n2254 vdd.n2253 16.0975
R18566 vdd.n2712 vdd.n2711 16.0975
R18567 vdd.n590 vdd.n589 16.0975
R18568 vdd.t79 vdd.n2218 15.4182
R18569 vdd.n2471 vdd.t181 15.4182
R18570 vdd.n28 vdd.n27 14.5458
R18571 vdd.n1989 vdd.n839 14.5112
R18572 vdd.n2673 vdd.n484 14.5112
R18573 vdd.n292 vdd.n257 13.1884
R18574 vdd.n245 vdd.n210 13.1884
R18575 vdd.n202 vdd.n167 13.1884
R18576 vdd.n155 vdd.n120 13.1884
R18577 vdd.n113 vdd.n78 13.1884
R18578 vdd.n66 vdd.n31 13.1884
R18579 vdd.n1107 vdd.n1072 13.1884
R18580 vdd.n1154 vdd.n1119 13.1884
R18581 vdd.n1017 vdd.n982 13.1884
R18582 vdd.n1064 vdd.n1029 13.1884
R18583 vdd.n928 vdd.n893 13.1884
R18584 vdd.n975 vdd.n940 13.1884
R18585 vdd.n1391 vdd.n1256 12.9944
R18586 vdd.n1395 vdd.n1256 12.9944
R18587 vdd.n1691 vdd.n1543 12.9944
R18588 vdd.n1692 vdd.n1691 12.9944
R18589 vdd.n2988 vdd.n364 12.9944
R18590 vdd.n2989 vdd.n2988 12.9944
R18591 vdd.n2806 vdd.n536 12.9944
R18592 vdd.n2809 vdd.n2806 12.9944
R18593 vdd.n293 vdd.n255 12.8005
R18594 vdd.n288 vdd.n259 12.8005
R18595 vdd.n246 vdd.n208 12.8005
R18596 vdd.n241 vdd.n212 12.8005
R18597 vdd.n203 vdd.n165 12.8005
R18598 vdd.n198 vdd.n169 12.8005
R18599 vdd.n156 vdd.n118 12.8005
R18600 vdd.n151 vdd.n122 12.8005
R18601 vdd.n114 vdd.n76 12.8005
R18602 vdd.n109 vdd.n80 12.8005
R18603 vdd.n67 vdd.n29 12.8005
R18604 vdd.n62 vdd.n33 12.8005
R18605 vdd.n1108 vdd.n1070 12.8005
R18606 vdd.n1103 vdd.n1074 12.8005
R18607 vdd.n1155 vdd.n1117 12.8005
R18608 vdd.n1150 vdd.n1121 12.8005
R18609 vdd.n1018 vdd.n980 12.8005
R18610 vdd.n1013 vdd.n984 12.8005
R18611 vdd.n1065 vdd.n1027 12.8005
R18612 vdd.n1060 vdd.n1031 12.8005
R18613 vdd.n929 vdd.n891 12.8005
R18614 vdd.n924 vdd.n895 12.8005
R18615 vdd.n976 vdd.n938 12.8005
R18616 vdd.n971 vdd.n942 12.8005
R18617 vdd.n287 vdd.n260 12.0247
R18618 vdd.n240 vdd.n213 12.0247
R18619 vdd.n197 vdd.n170 12.0247
R18620 vdd.n150 vdd.n123 12.0247
R18621 vdd.n108 vdd.n81 12.0247
R18622 vdd.n61 vdd.n34 12.0247
R18623 vdd.n1102 vdd.n1075 12.0247
R18624 vdd.n1149 vdd.n1122 12.0247
R18625 vdd.n1012 vdd.n985 12.0247
R18626 vdd.n1059 vdd.n1032 12.0247
R18627 vdd.n923 vdd.n896 12.0247
R18628 vdd.n970 vdd.n943 12.0247
R18629 vdd.n1430 vdd.n1186 11.337
R18630 vdd.n1439 vdd.n1186 11.337
R18631 vdd.n1439 vdd.n1438 11.337
R18632 vdd.n1447 vdd.n1180 11.337
R18633 vdd.n1456 vdd.n1455 11.337
R18634 vdd.n1473 vdd.n1164 11.337
R18635 vdd.n1481 vdd.n887 11.337
R18636 vdd.n1490 vdd.n1489 11.337
R18637 vdd.n1498 vdd.n870 11.337
R18638 vdd.n1509 vdd.n870 11.337
R18639 vdd.n1509 vdd.n1508 11.337
R18640 vdd.n2849 vdd.n473 11.337
R18641 vdd.n2858 vdd.n473 11.337
R18642 vdd.n2858 vdd.n2857 11.337
R18643 vdd.n2866 vdd.n467 11.337
R18644 vdd.n2882 vdd.n456 11.337
R18645 vdd.n3043 vdd.n304 11.337
R18646 vdd.n3041 vdd.n308 11.337
R18647 vdd.n3035 vdd.n3034 11.337
R18648 vdd.n3033 vdd.n318 11.337
R18649 vdd.n3027 vdd.n318 11.337
R18650 vdd.n3027 vdd.n3026 11.337
R18651 vdd.n284 vdd.n283 11.249
R18652 vdd.n237 vdd.n236 11.249
R18653 vdd.n194 vdd.n193 11.249
R18654 vdd.n147 vdd.n146 11.249
R18655 vdd.n105 vdd.n104 11.249
R18656 vdd.n58 vdd.n57 11.249
R18657 vdd.n1099 vdd.n1098 11.249
R18658 vdd.n1146 vdd.n1145 11.249
R18659 vdd.n1009 vdd.n1008 11.249
R18660 vdd.n1056 vdd.n1055 11.249
R18661 vdd.n920 vdd.n919 11.249
R18662 vdd.n967 vdd.n966 11.249
R18663 vdd.n2146 vdd.t4 11.1103
R18664 vdd.n2478 vdd.t196 11.1103
R18665 vdd.n1228 vdd.t93 10.7702
R18666 vdd.t104 vdd.n3025 10.7702
R18667 vdd.n269 vdd.n268 10.7238
R18668 vdd.n222 vdd.n221 10.7238
R18669 vdd.n179 vdd.n178 10.7238
R18670 vdd.n132 vdd.n131 10.7238
R18671 vdd.n90 vdd.n89 10.7238
R18672 vdd.n43 vdd.n42 10.7238
R18673 vdd.n1084 vdd.n1083 10.7238
R18674 vdd.n1131 vdd.n1130 10.7238
R18675 vdd.n994 vdd.n993 10.7238
R18676 vdd.n1041 vdd.n1040 10.7238
R18677 vdd.n905 vdd.n904 10.7238
R18678 vdd.n952 vdd.n951 10.7238
R18679 vdd.n1992 vdd.n1991 10.6151
R18680 vdd.n1993 vdd.n1992 10.6151
R18681 vdd.n1993 vdd.n825 10.6151
R18682 vdd.n2003 vdd.n825 10.6151
R18683 vdd.n2004 vdd.n2003 10.6151
R18684 vdd.n2005 vdd.n2004 10.6151
R18685 vdd.n2005 vdd.n812 10.6151
R18686 vdd.n2016 vdd.n812 10.6151
R18687 vdd.n2017 vdd.n2016 10.6151
R18688 vdd.n2018 vdd.n2017 10.6151
R18689 vdd.n2018 vdd.n800 10.6151
R18690 vdd.n2028 vdd.n800 10.6151
R18691 vdd.n2029 vdd.n2028 10.6151
R18692 vdd.n2030 vdd.n2029 10.6151
R18693 vdd.n2030 vdd.n788 10.6151
R18694 vdd.n2040 vdd.n788 10.6151
R18695 vdd.n2041 vdd.n2040 10.6151
R18696 vdd.n2042 vdd.n2041 10.6151
R18697 vdd.n2042 vdd.n777 10.6151
R18698 vdd.n2052 vdd.n777 10.6151
R18699 vdd.n2053 vdd.n2052 10.6151
R18700 vdd.n2054 vdd.n2053 10.6151
R18701 vdd.n2054 vdd.n764 10.6151
R18702 vdd.n2066 vdd.n764 10.6151
R18703 vdd.n2067 vdd.n2066 10.6151
R18704 vdd.n2069 vdd.n2067 10.6151
R18705 vdd.n2069 vdd.n2068 10.6151
R18706 vdd.n2068 vdd.n746 10.6151
R18707 vdd.n2216 vdd.n2215 10.6151
R18708 vdd.n2215 vdd.n2214 10.6151
R18709 vdd.n2214 vdd.n2211 10.6151
R18710 vdd.n2211 vdd.n2210 10.6151
R18711 vdd.n2210 vdd.n2207 10.6151
R18712 vdd.n2207 vdd.n2206 10.6151
R18713 vdd.n2206 vdd.n2203 10.6151
R18714 vdd.n2203 vdd.n2202 10.6151
R18715 vdd.n2202 vdd.n2199 10.6151
R18716 vdd.n2199 vdd.n2198 10.6151
R18717 vdd.n2198 vdd.n2195 10.6151
R18718 vdd.n2195 vdd.n2194 10.6151
R18719 vdd.n2194 vdd.n2191 10.6151
R18720 vdd.n2191 vdd.n2190 10.6151
R18721 vdd.n2190 vdd.n2187 10.6151
R18722 vdd.n2187 vdd.n2186 10.6151
R18723 vdd.n2186 vdd.n2183 10.6151
R18724 vdd.n2183 vdd.n2182 10.6151
R18725 vdd.n2182 vdd.n2179 10.6151
R18726 vdd.n2179 vdd.n2178 10.6151
R18727 vdd.n2178 vdd.n2175 10.6151
R18728 vdd.n2175 vdd.n2174 10.6151
R18729 vdd.n2174 vdd.n2171 10.6151
R18730 vdd.n2171 vdd.n2170 10.6151
R18731 vdd.n2170 vdd.n2167 10.6151
R18732 vdd.n2167 vdd.n2166 10.6151
R18733 vdd.n2166 vdd.n2163 10.6151
R18734 vdd.n2163 vdd.n2162 10.6151
R18735 vdd.n2162 vdd.n2159 10.6151
R18736 vdd.n2159 vdd.n2158 10.6151
R18737 vdd.n2158 vdd.n2155 10.6151
R18738 vdd.n2153 vdd.n2150 10.6151
R18739 vdd.n2150 vdd.n2149 10.6151
R18740 vdd.n1892 vdd.n1891 10.6151
R18741 vdd.n1891 vdd.n1889 10.6151
R18742 vdd.n1889 vdd.n1888 10.6151
R18743 vdd.n1888 vdd.n1886 10.6151
R18744 vdd.n1886 vdd.n1885 10.6151
R18745 vdd.n1885 vdd.n1883 10.6151
R18746 vdd.n1883 vdd.n1882 10.6151
R18747 vdd.n1882 vdd.n1880 10.6151
R18748 vdd.n1880 vdd.n1879 10.6151
R18749 vdd.n1879 vdd.n1877 10.6151
R18750 vdd.n1877 vdd.n1876 10.6151
R18751 vdd.n1876 vdd.n1874 10.6151
R18752 vdd.n1874 vdd.n1873 10.6151
R18753 vdd.n1873 vdd.n1788 10.6151
R18754 vdd.n1788 vdd.n1787 10.6151
R18755 vdd.n1787 vdd.n1785 10.6151
R18756 vdd.n1785 vdd.n1784 10.6151
R18757 vdd.n1784 vdd.n1782 10.6151
R18758 vdd.n1782 vdd.n1781 10.6151
R18759 vdd.n1781 vdd.n1779 10.6151
R18760 vdd.n1779 vdd.n1778 10.6151
R18761 vdd.n1778 vdd.n1776 10.6151
R18762 vdd.n1776 vdd.n1775 10.6151
R18763 vdd.n1775 vdd.n1773 10.6151
R18764 vdd.n1773 vdd.n1772 10.6151
R18765 vdd.n1772 vdd.n1769 10.6151
R18766 vdd.n1769 vdd.n1768 10.6151
R18767 vdd.n1768 vdd.n749 10.6151
R18768 vdd.n1726 vdd.n837 10.6151
R18769 vdd.n1727 vdd.n1726 10.6151
R18770 vdd.n1728 vdd.n1727 10.6151
R18771 vdd.n1728 vdd.n1722 10.6151
R18772 vdd.n1734 vdd.n1722 10.6151
R18773 vdd.n1735 vdd.n1734 10.6151
R18774 vdd.n1736 vdd.n1735 10.6151
R18775 vdd.n1736 vdd.n1720 10.6151
R18776 vdd.n1742 vdd.n1720 10.6151
R18777 vdd.n1743 vdd.n1742 10.6151
R18778 vdd.n1744 vdd.n1743 10.6151
R18779 vdd.n1744 vdd.n1718 10.6151
R18780 vdd.n1750 vdd.n1718 10.6151
R18781 vdd.n1751 vdd.n1750 10.6151
R18782 vdd.n1752 vdd.n1751 10.6151
R18783 vdd.n1752 vdd.n1716 10.6151
R18784 vdd.n1928 vdd.n1716 10.6151
R18785 vdd.n1928 vdd.n1927 10.6151
R18786 vdd.n1927 vdd.n1757 10.6151
R18787 vdd.n1921 vdd.n1757 10.6151
R18788 vdd.n1921 vdd.n1920 10.6151
R18789 vdd.n1920 vdd.n1919 10.6151
R18790 vdd.n1919 vdd.n1759 10.6151
R18791 vdd.n1913 vdd.n1759 10.6151
R18792 vdd.n1913 vdd.n1912 10.6151
R18793 vdd.n1912 vdd.n1911 10.6151
R18794 vdd.n1911 vdd.n1761 10.6151
R18795 vdd.n1905 vdd.n1761 10.6151
R18796 vdd.n1905 vdd.n1904 10.6151
R18797 vdd.n1904 vdd.n1903 10.6151
R18798 vdd.n1903 vdd.n1763 10.6151
R18799 vdd.n1897 vdd.n1896 10.6151
R18800 vdd.n1896 vdd.n1895 10.6151
R18801 vdd.n2401 vdd.n2400 10.6151
R18802 vdd.n2400 vdd.n2398 10.6151
R18803 vdd.n2398 vdd.n2397 10.6151
R18804 vdd.n2397 vdd.n2255 10.6151
R18805 vdd.n2344 vdd.n2255 10.6151
R18806 vdd.n2345 vdd.n2344 10.6151
R18807 vdd.n2347 vdd.n2345 10.6151
R18808 vdd.n2348 vdd.n2347 10.6151
R18809 vdd.n2350 vdd.n2348 10.6151
R18810 vdd.n2351 vdd.n2350 10.6151
R18811 vdd.n2353 vdd.n2351 10.6151
R18812 vdd.n2354 vdd.n2353 10.6151
R18813 vdd.n2356 vdd.n2354 10.6151
R18814 vdd.n2357 vdd.n2356 10.6151
R18815 vdd.n2372 vdd.n2357 10.6151
R18816 vdd.n2372 vdd.n2371 10.6151
R18817 vdd.n2371 vdd.n2370 10.6151
R18818 vdd.n2370 vdd.n2368 10.6151
R18819 vdd.n2368 vdd.n2367 10.6151
R18820 vdd.n2367 vdd.n2365 10.6151
R18821 vdd.n2365 vdd.n2364 10.6151
R18822 vdd.n2364 vdd.n2362 10.6151
R18823 vdd.n2362 vdd.n2361 10.6151
R18824 vdd.n2361 vdd.n2359 10.6151
R18825 vdd.n2359 vdd.n2358 10.6151
R18826 vdd.n2358 vdd.n626 10.6151
R18827 vdd.n2606 vdd.n626 10.6151
R18828 vdd.n2607 vdd.n2606 10.6151
R18829 vdd.n2468 vdd.n702 10.6151
R18830 vdd.n2468 vdd.n2467 10.6151
R18831 vdd.n2467 vdd.n2466 10.6151
R18832 vdd.n2466 vdd.n2464 10.6151
R18833 vdd.n2464 vdd.n2461 10.6151
R18834 vdd.n2461 vdd.n2460 10.6151
R18835 vdd.n2460 vdd.n2457 10.6151
R18836 vdd.n2457 vdd.n2456 10.6151
R18837 vdd.n2456 vdd.n2453 10.6151
R18838 vdd.n2453 vdd.n2452 10.6151
R18839 vdd.n2452 vdd.n2449 10.6151
R18840 vdd.n2449 vdd.n2448 10.6151
R18841 vdd.n2448 vdd.n2445 10.6151
R18842 vdd.n2445 vdd.n2444 10.6151
R18843 vdd.n2444 vdd.n2441 10.6151
R18844 vdd.n2441 vdd.n2440 10.6151
R18845 vdd.n2440 vdd.n2437 10.6151
R18846 vdd.n2437 vdd.n2436 10.6151
R18847 vdd.n2436 vdd.n2433 10.6151
R18848 vdd.n2433 vdd.n2432 10.6151
R18849 vdd.n2432 vdd.n2429 10.6151
R18850 vdd.n2429 vdd.n2428 10.6151
R18851 vdd.n2428 vdd.n2425 10.6151
R18852 vdd.n2425 vdd.n2424 10.6151
R18853 vdd.n2424 vdd.n2421 10.6151
R18854 vdd.n2421 vdd.n2420 10.6151
R18855 vdd.n2420 vdd.n2417 10.6151
R18856 vdd.n2417 vdd.n2416 10.6151
R18857 vdd.n2416 vdd.n2413 10.6151
R18858 vdd.n2413 vdd.n2412 10.6151
R18859 vdd.n2412 vdd.n2409 10.6151
R18860 vdd.n2407 vdd.n2404 10.6151
R18861 vdd.n2404 vdd.n2403 10.6151
R18862 vdd.n2481 vdd.n2480 10.6151
R18863 vdd.n2482 vdd.n2481 10.6151
R18864 vdd.n2482 vdd.n692 10.6151
R18865 vdd.n2492 vdd.n692 10.6151
R18866 vdd.n2493 vdd.n2492 10.6151
R18867 vdd.n2494 vdd.n2493 10.6151
R18868 vdd.n2494 vdd.n679 10.6151
R18869 vdd.n2504 vdd.n679 10.6151
R18870 vdd.n2505 vdd.n2504 10.6151
R18871 vdd.n2506 vdd.n2505 10.6151
R18872 vdd.n2506 vdd.n668 10.6151
R18873 vdd.n2516 vdd.n668 10.6151
R18874 vdd.n2517 vdd.n2516 10.6151
R18875 vdd.n2518 vdd.n2517 10.6151
R18876 vdd.n2518 vdd.n656 10.6151
R18877 vdd.n2528 vdd.n656 10.6151
R18878 vdd.n2529 vdd.n2528 10.6151
R18879 vdd.n2530 vdd.n2529 10.6151
R18880 vdd.n2530 vdd.n645 10.6151
R18881 vdd.n2542 vdd.n645 10.6151
R18882 vdd.n2543 vdd.n2542 10.6151
R18883 vdd.n2544 vdd.n2543 10.6151
R18884 vdd.n2544 vdd.n631 10.6151
R18885 vdd.n2599 vdd.n631 10.6151
R18886 vdd.n2600 vdd.n2599 10.6151
R18887 vdd.n2601 vdd.n2600 10.6151
R18888 vdd.n2601 vdd.n600 10.6151
R18889 vdd.n2671 vdd.n600 10.6151
R18890 vdd.n2670 vdd.n2669 10.6151
R18891 vdd.n2669 vdd.n601 10.6151
R18892 vdd.n602 vdd.n601 10.6151
R18893 vdd.n2662 vdd.n602 10.6151
R18894 vdd.n2662 vdd.n2661 10.6151
R18895 vdd.n2661 vdd.n2660 10.6151
R18896 vdd.n2660 vdd.n604 10.6151
R18897 vdd.n2655 vdd.n604 10.6151
R18898 vdd.n2655 vdd.n2654 10.6151
R18899 vdd.n2654 vdd.n2653 10.6151
R18900 vdd.n2653 vdd.n607 10.6151
R18901 vdd.n2648 vdd.n607 10.6151
R18902 vdd.n2648 vdd.n2647 10.6151
R18903 vdd.n2647 vdd.n2646 10.6151
R18904 vdd.n2646 vdd.n610 10.6151
R18905 vdd.n2641 vdd.n610 10.6151
R18906 vdd.n2641 vdd.n520 10.6151
R18907 vdd.n2637 vdd.n520 10.6151
R18908 vdd.n2637 vdd.n2636 10.6151
R18909 vdd.n2636 vdd.n2635 10.6151
R18910 vdd.n2635 vdd.n613 10.6151
R18911 vdd.n2630 vdd.n613 10.6151
R18912 vdd.n2630 vdd.n2629 10.6151
R18913 vdd.n2629 vdd.n2628 10.6151
R18914 vdd.n2628 vdd.n616 10.6151
R18915 vdd.n2623 vdd.n616 10.6151
R18916 vdd.n2623 vdd.n2622 10.6151
R18917 vdd.n2622 vdd.n2621 10.6151
R18918 vdd.n2621 vdd.n619 10.6151
R18919 vdd.n2616 vdd.n619 10.6151
R18920 vdd.n2616 vdd.n2615 10.6151
R18921 vdd.n2613 vdd.n624 10.6151
R18922 vdd.n2608 vdd.n624 10.6151
R18923 vdd.n2589 vdd.n2550 10.6151
R18924 vdd.n2584 vdd.n2550 10.6151
R18925 vdd.n2584 vdd.n2583 10.6151
R18926 vdd.n2583 vdd.n2582 10.6151
R18927 vdd.n2582 vdd.n2552 10.6151
R18928 vdd.n2577 vdd.n2552 10.6151
R18929 vdd.n2577 vdd.n2576 10.6151
R18930 vdd.n2576 vdd.n2575 10.6151
R18931 vdd.n2575 vdd.n2555 10.6151
R18932 vdd.n2570 vdd.n2555 10.6151
R18933 vdd.n2570 vdd.n2569 10.6151
R18934 vdd.n2569 vdd.n2568 10.6151
R18935 vdd.n2568 vdd.n2558 10.6151
R18936 vdd.n2563 vdd.n2558 10.6151
R18937 vdd.n2563 vdd.n2562 10.6151
R18938 vdd.n2562 vdd.n575 10.6151
R18939 vdd.n2706 vdd.n575 10.6151
R18940 vdd.n2706 vdd.n576 10.6151
R18941 vdd.n578 vdd.n576 10.6151
R18942 vdd.n2699 vdd.n578 10.6151
R18943 vdd.n2699 vdd.n2698 10.6151
R18944 vdd.n2698 vdd.n2697 10.6151
R18945 vdd.n2697 vdd.n580 10.6151
R18946 vdd.n2692 vdd.n580 10.6151
R18947 vdd.n2692 vdd.n2691 10.6151
R18948 vdd.n2691 vdd.n2690 10.6151
R18949 vdd.n2690 vdd.n583 10.6151
R18950 vdd.n2685 vdd.n583 10.6151
R18951 vdd.n2685 vdd.n2684 10.6151
R18952 vdd.n2684 vdd.n2683 10.6151
R18953 vdd.n2683 vdd.n586 10.6151
R18954 vdd.n2678 vdd.n2677 10.6151
R18955 vdd.n2677 vdd.n2676 10.6151
R18956 vdd.n2324 vdd.n2322 10.6151
R18957 vdd.n2325 vdd.n2324 10.6151
R18958 vdd.n2393 vdd.n2325 10.6151
R18959 vdd.n2393 vdd.n2392 10.6151
R18960 vdd.n2392 vdd.n2391 10.6151
R18961 vdd.n2391 vdd.n2389 10.6151
R18962 vdd.n2389 vdd.n2388 10.6151
R18963 vdd.n2388 vdd.n2386 10.6151
R18964 vdd.n2386 vdd.n2385 10.6151
R18965 vdd.n2385 vdd.n2383 10.6151
R18966 vdd.n2383 vdd.n2382 10.6151
R18967 vdd.n2382 vdd.n2380 10.6151
R18968 vdd.n2380 vdd.n2379 10.6151
R18969 vdd.n2379 vdd.n2377 10.6151
R18970 vdd.n2377 vdd.n2376 10.6151
R18971 vdd.n2376 vdd.n2342 10.6151
R18972 vdd.n2342 vdd.n2341 10.6151
R18973 vdd.n2341 vdd.n2339 10.6151
R18974 vdd.n2339 vdd.n2338 10.6151
R18975 vdd.n2338 vdd.n2336 10.6151
R18976 vdd.n2336 vdd.n2335 10.6151
R18977 vdd.n2335 vdd.n2333 10.6151
R18978 vdd.n2333 vdd.n2332 10.6151
R18979 vdd.n2332 vdd.n2330 10.6151
R18980 vdd.n2330 vdd.n2329 10.6151
R18981 vdd.n2329 vdd.n2327 10.6151
R18982 vdd.n2327 vdd.n2326 10.6151
R18983 vdd.n2326 vdd.n592 10.6151
R18984 vdd.n2475 vdd.n2474 10.6151
R18985 vdd.n2474 vdd.n707 10.6151
R18986 vdd.n2259 vdd.n707 10.6151
R18987 vdd.n2262 vdd.n2259 10.6151
R18988 vdd.n2263 vdd.n2262 10.6151
R18989 vdd.n2266 vdd.n2263 10.6151
R18990 vdd.n2267 vdd.n2266 10.6151
R18991 vdd.n2270 vdd.n2267 10.6151
R18992 vdd.n2271 vdd.n2270 10.6151
R18993 vdd.n2274 vdd.n2271 10.6151
R18994 vdd.n2275 vdd.n2274 10.6151
R18995 vdd.n2278 vdd.n2275 10.6151
R18996 vdd.n2279 vdd.n2278 10.6151
R18997 vdd.n2282 vdd.n2279 10.6151
R18998 vdd.n2283 vdd.n2282 10.6151
R18999 vdd.n2286 vdd.n2283 10.6151
R19000 vdd.n2287 vdd.n2286 10.6151
R19001 vdd.n2290 vdd.n2287 10.6151
R19002 vdd.n2291 vdd.n2290 10.6151
R19003 vdd.n2294 vdd.n2291 10.6151
R19004 vdd.n2295 vdd.n2294 10.6151
R19005 vdd.n2298 vdd.n2295 10.6151
R19006 vdd.n2299 vdd.n2298 10.6151
R19007 vdd.n2302 vdd.n2299 10.6151
R19008 vdd.n2303 vdd.n2302 10.6151
R19009 vdd.n2306 vdd.n2303 10.6151
R19010 vdd.n2307 vdd.n2306 10.6151
R19011 vdd.n2310 vdd.n2307 10.6151
R19012 vdd.n2311 vdd.n2310 10.6151
R19013 vdd.n2314 vdd.n2311 10.6151
R19014 vdd.n2315 vdd.n2314 10.6151
R19015 vdd.n2320 vdd.n2318 10.6151
R19016 vdd.n2321 vdd.n2320 10.6151
R19017 vdd.n2476 vdd.n697 10.6151
R19018 vdd.n2486 vdd.n697 10.6151
R19019 vdd.n2487 vdd.n2486 10.6151
R19020 vdd.n2488 vdd.n2487 10.6151
R19021 vdd.n2488 vdd.n685 10.6151
R19022 vdd.n2498 vdd.n685 10.6151
R19023 vdd.n2499 vdd.n2498 10.6151
R19024 vdd.n2500 vdd.n2499 10.6151
R19025 vdd.n2500 vdd.n674 10.6151
R19026 vdd.n2510 vdd.n674 10.6151
R19027 vdd.n2511 vdd.n2510 10.6151
R19028 vdd.n2512 vdd.n2511 10.6151
R19029 vdd.n2512 vdd.n662 10.6151
R19030 vdd.n2522 vdd.n662 10.6151
R19031 vdd.n2523 vdd.n2522 10.6151
R19032 vdd.n2524 vdd.n2523 10.6151
R19033 vdd.n2524 vdd.n651 10.6151
R19034 vdd.n2534 vdd.n651 10.6151
R19035 vdd.n2535 vdd.n2534 10.6151
R19036 vdd.n2538 vdd.n2535 10.6151
R19037 vdd.n2548 vdd.n639 10.6151
R19038 vdd.n2549 vdd.n2548 10.6151
R19039 vdd.n2595 vdd.n2549 10.6151
R19040 vdd.n2595 vdd.n2594 10.6151
R19041 vdd.n2594 vdd.n2593 10.6151
R19042 vdd.n2593 vdd.n2592 10.6151
R19043 vdd.n2592 vdd.n2590 10.6151
R19044 vdd.n1987 vdd.n831 10.6151
R19045 vdd.n1997 vdd.n831 10.6151
R19046 vdd.n1998 vdd.n1997 10.6151
R19047 vdd.n1999 vdd.n1998 10.6151
R19048 vdd.n1999 vdd.n818 10.6151
R19049 vdd.n2009 vdd.n818 10.6151
R19050 vdd.n2010 vdd.n2009 10.6151
R19051 vdd.n2012 vdd.n806 10.6151
R19052 vdd.n2022 vdd.n806 10.6151
R19053 vdd.n2023 vdd.n2022 10.6151
R19054 vdd.n2024 vdd.n2023 10.6151
R19055 vdd.n2024 vdd.n794 10.6151
R19056 vdd.n2034 vdd.n794 10.6151
R19057 vdd.n2035 vdd.n2034 10.6151
R19058 vdd.n2036 vdd.n2035 10.6151
R19059 vdd.n2036 vdd.n783 10.6151
R19060 vdd.n2046 vdd.n783 10.6151
R19061 vdd.n2047 vdd.n2046 10.6151
R19062 vdd.n2048 vdd.n2047 10.6151
R19063 vdd.n2048 vdd.n771 10.6151
R19064 vdd.n2058 vdd.n771 10.6151
R19065 vdd.n2059 vdd.n2058 10.6151
R19066 vdd.n2062 vdd.n2059 10.6151
R19067 vdd.n2062 vdd.n2061 10.6151
R19068 vdd.n2061 vdd.n2060 10.6151
R19069 vdd.n2060 vdd.n754 10.6151
R19070 vdd.n2144 vdd.n754 10.6151
R19071 vdd.n2143 vdd.n2142 10.6151
R19072 vdd.n2142 vdd.n2139 10.6151
R19073 vdd.n2139 vdd.n2138 10.6151
R19074 vdd.n2138 vdd.n2135 10.6151
R19075 vdd.n2135 vdd.n2134 10.6151
R19076 vdd.n2134 vdd.n2131 10.6151
R19077 vdd.n2131 vdd.n2130 10.6151
R19078 vdd.n2130 vdd.n2127 10.6151
R19079 vdd.n2127 vdd.n2126 10.6151
R19080 vdd.n2126 vdd.n2123 10.6151
R19081 vdd.n2123 vdd.n2122 10.6151
R19082 vdd.n2122 vdd.n2119 10.6151
R19083 vdd.n2119 vdd.n2118 10.6151
R19084 vdd.n2118 vdd.n2115 10.6151
R19085 vdd.n2115 vdd.n2114 10.6151
R19086 vdd.n2114 vdd.n2111 10.6151
R19087 vdd.n2111 vdd.n2110 10.6151
R19088 vdd.n2110 vdd.n2107 10.6151
R19089 vdd.n2107 vdd.n2106 10.6151
R19090 vdd.n2106 vdd.n2103 10.6151
R19091 vdd.n2103 vdd.n2102 10.6151
R19092 vdd.n2102 vdd.n2099 10.6151
R19093 vdd.n2099 vdd.n2098 10.6151
R19094 vdd.n2098 vdd.n2095 10.6151
R19095 vdd.n2095 vdd.n2094 10.6151
R19096 vdd.n2094 vdd.n2091 10.6151
R19097 vdd.n2091 vdd.n2090 10.6151
R19098 vdd.n2090 vdd.n2087 10.6151
R19099 vdd.n2087 vdd.n2086 10.6151
R19100 vdd.n2086 vdd.n2083 10.6151
R19101 vdd.n2083 vdd.n2082 10.6151
R19102 vdd.n2079 vdd.n2078 10.6151
R19103 vdd.n2078 vdd.n2076 10.6151
R19104 vdd.n1835 vdd.n1833 10.6151
R19105 vdd.n1836 vdd.n1835 10.6151
R19106 vdd.n1838 vdd.n1836 10.6151
R19107 vdd.n1839 vdd.n1838 10.6151
R19108 vdd.n1841 vdd.n1839 10.6151
R19109 vdd.n1842 vdd.n1841 10.6151
R19110 vdd.n1844 vdd.n1842 10.6151
R19111 vdd.n1845 vdd.n1844 10.6151
R19112 vdd.n1847 vdd.n1845 10.6151
R19113 vdd.n1848 vdd.n1847 10.6151
R19114 vdd.n1850 vdd.n1848 10.6151
R19115 vdd.n1851 vdd.n1850 10.6151
R19116 vdd.n1869 vdd.n1851 10.6151
R19117 vdd.n1869 vdd.n1868 10.6151
R19118 vdd.n1868 vdd.n1867 10.6151
R19119 vdd.n1867 vdd.n1865 10.6151
R19120 vdd.n1865 vdd.n1864 10.6151
R19121 vdd.n1864 vdd.n1862 10.6151
R19122 vdd.n1862 vdd.n1861 10.6151
R19123 vdd.n1861 vdd.n1859 10.6151
R19124 vdd.n1859 vdd.n1858 10.6151
R19125 vdd.n1858 vdd.n1856 10.6151
R19126 vdd.n1856 vdd.n1855 10.6151
R19127 vdd.n1855 vdd.n1853 10.6151
R19128 vdd.n1853 vdd.n1852 10.6151
R19129 vdd.n1852 vdd.n758 10.6151
R19130 vdd.n2074 vdd.n758 10.6151
R19131 vdd.n2075 vdd.n2074 10.6151
R19132 vdd.n1986 vdd.n1985 10.6151
R19133 vdd.n1985 vdd.n843 10.6151
R19134 vdd.n1979 vdd.n843 10.6151
R19135 vdd.n1979 vdd.n1978 10.6151
R19136 vdd.n1978 vdd.n1977 10.6151
R19137 vdd.n1977 vdd.n845 10.6151
R19138 vdd.n1971 vdd.n845 10.6151
R19139 vdd.n1971 vdd.n1970 10.6151
R19140 vdd.n1970 vdd.n1969 10.6151
R19141 vdd.n1969 vdd.n847 10.6151
R19142 vdd.n1963 vdd.n847 10.6151
R19143 vdd.n1963 vdd.n1962 10.6151
R19144 vdd.n1962 vdd.n1961 10.6151
R19145 vdd.n1961 vdd.n849 10.6151
R19146 vdd.n1955 vdd.n849 10.6151
R19147 vdd.n1955 vdd.n1954 10.6151
R19148 vdd.n1954 vdd.n1953 10.6151
R19149 vdd.n1953 vdd.n853 10.6151
R19150 vdd.n1801 vdd.n853 10.6151
R19151 vdd.n1802 vdd.n1801 10.6151
R19152 vdd.n1802 vdd.n1797 10.6151
R19153 vdd.n1808 vdd.n1797 10.6151
R19154 vdd.n1809 vdd.n1808 10.6151
R19155 vdd.n1810 vdd.n1809 10.6151
R19156 vdd.n1810 vdd.n1795 10.6151
R19157 vdd.n1816 vdd.n1795 10.6151
R19158 vdd.n1817 vdd.n1816 10.6151
R19159 vdd.n1818 vdd.n1817 10.6151
R19160 vdd.n1818 vdd.n1793 10.6151
R19161 vdd.n1824 vdd.n1793 10.6151
R19162 vdd.n1825 vdd.n1824 10.6151
R19163 vdd.n1827 vdd.n1789 10.6151
R19164 vdd.n1832 vdd.n1789 10.6151
R19165 vdd.n280 vdd.n262 10.4732
R19166 vdd.n233 vdd.n215 10.4732
R19167 vdd.n190 vdd.n172 10.4732
R19168 vdd.n143 vdd.n125 10.4732
R19169 vdd.n101 vdd.n83 10.4732
R19170 vdd.n54 vdd.n36 10.4732
R19171 vdd.n1095 vdd.n1077 10.4732
R19172 vdd.n1142 vdd.n1124 10.4732
R19173 vdd.n1005 vdd.n987 10.4732
R19174 vdd.n1052 vdd.n1034 10.4732
R19175 vdd.n916 vdd.n898 10.4732
R19176 vdd.n963 vdd.n945 10.4732
R19177 vdd.t18 vdd.n888 10.3167
R19178 vdd.n2874 vdd.t38 10.3167
R19179 vdd.n1465 vdd.t14 10.09
R19180 vdd.n3042 vdd.t51 10.09
R19181 vdd.n279 vdd.n264 9.69747
R19182 vdd.n232 vdd.n217 9.69747
R19183 vdd.n189 vdd.n174 9.69747
R19184 vdd.n142 vdd.n127 9.69747
R19185 vdd.n100 vdd.n85 9.69747
R19186 vdd.n53 vdd.n38 9.69747
R19187 vdd.n1094 vdd.n1079 9.69747
R19188 vdd.n1141 vdd.n1126 9.69747
R19189 vdd.n1004 vdd.n989 9.69747
R19190 vdd.n1051 vdd.n1036 9.69747
R19191 vdd.n915 vdd.n900 9.69747
R19192 vdd.n962 vdd.n947 9.69747
R19193 vdd.n1929 vdd.n1928 9.67831
R19194 vdd.n2836 vdd.n520 9.67831
R19195 vdd.n2707 vdd.n2706 9.67831
R19196 vdd.n1953 vdd.n1952 9.67831
R19197 vdd.n295 vdd.n294 9.45567
R19198 vdd.n248 vdd.n247 9.45567
R19199 vdd.n205 vdd.n204 9.45567
R19200 vdd.n158 vdd.n157 9.45567
R19201 vdd.n116 vdd.n115 9.45567
R19202 vdd.n69 vdd.n68 9.45567
R19203 vdd.n1110 vdd.n1109 9.45567
R19204 vdd.n1157 vdd.n1156 9.45567
R19205 vdd.n1020 vdd.n1019 9.45567
R19206 vdd.n1067 vdd.n1066 9.45567
R19207 vdd.n931 vdd.n930 9.45567
R19208 vdd.n978 vdd.n977 9.45567
R19209 vdd.n1689 vdd.n1543 9.3005
R19210 vdd.n1688 vdd.n1687 9.3005
R19211 vdd.n1549 vdd.n1548 9.3005
R19212 vdd.n1682 vdd.n1553 9.3005
R19213 vdd.n1681 vdd.n1554 9.3005
R19214 vdd.n1680 vdd.n1555 9.3005
R19215 vdd.n1559 vdd.n1556 9.3005
R19216 vdd.n1675 vdd.n1560 9.3005
R19217 vdd.n1674 vdd.n1561 9.3005
R19218 vdd.n1673 vdd.n1562 9.3005
R19219 vdd.n1566 vdd.n1563 9.3005
R19220 vdd.n1668 vdd.n1567 9.3005
R19221 vdd.n1667 vdd.n1568 9.3005
R19222 vdd.n1666 vdd.n1569 9.3005
R19223 vdd.n1573 vdd.n1570 9.3005
R19224 vdd.n1661 vdd.n1574 9.3005
R19225 vdd.n1660 vdd.n1575 9.3005
R19226 vdd.n1659 vdd.n1576 9.3005
R19227 vdd.n1580 vdd.n1577 9.3005
R19228 vdd.n1654 vdd.n1581 9.3005
R19229 vdd.n1653 vdd.n1582 9.3005
R19230 vdd.n1652 vdd.n1651 9.3005
R19231 vdd.n1650 vdd.n1583 9.3005
R19232 vdd.n1649 vdd.n1648 9.3005
R19233 vdd.n1589 vdd.n1588 9.3005
R19234 vdd.n1643 vdd.n1593 9.3005
R19235 vdd.n1642 vdd.n1594 9.3005
R19236 vdd.n1641 vdd.n1595 9.3005
R19237 vdd.n1599 vdd.n1596 9.3005
R19238 vdd.n1636 vdd.n1600 9.3005
R19239 vdd.n1635 vdd.n1601 9.3005
R19240 vdd.n1634 vdd.n1602 9.3005
R19241 vdd.n1606 vdd.n1603 9.3005
R19242 vdd.n1629 vdd.n1607 9.3005
R19243 vdd.n1628 vdd.n1608 9.3005
R19244 vdd.n1627 vdd.n1609 9.3005
R19245 vdd.n1611 vdd.n1610 9.3005
R19246 vdd.n1622 vdd.n854 9.3005
R19247 vdd.n1691 vdd.n1690 9.3005
R19248 vdd.n1715 vdd.n1714 9.3005
R19249 vdd.n1521 vdd.n1520 9.3005
R19250 vdd.n1526 vdd.n1524 9.3005
R19251 vdd.n1707 vdd.n1527 9.3005
R19252 vdd.n1706 vdd.n1528 9.3005
R19253 vdd.n1705 vdd.n1529 9.3005
R19254 vdd.n1533 vdd.n1530 9.3005
R19255 vdd.n1700 vdd.n1534 9.3005
R19256 vdd.n1699 vdd.n1535 9.3005
R19257 vdd.n1698 vdd.n1536 9.3005
R19258 vdd.n1540 vdd.n1537 9.3005
R19259 vdd.n1693 vdd.n1541 9.3005
R19260 vdd.n1692 vdd.n1542 9.3005
R19261 vdd.n1937 vdd.n1514 9.3005
R19262 vdd.n1939 vdd.n1938 9.3005
R19263 vdd.n1476 vdd.n1475 9.3005
R19264 vdd.n1477 vdd.n890 9.3005
R19265 vdd.n1479 vdd.n1478 9.3005
R19266 vdd.n880 vdd.n879 9.3005
R19267 vdd.n1493 vdd.n1492 9.3005
R19268 vdd.n1494 vdd.n878 9.3005
R19269 vdd.n1496 vdd.n1495 9.3005
R19270 vdd.n868 vdd.n867 9.3005
R19271 vdd.n1512 vdd.n1511 9.3005
R19272 vdd.n1513 vdd.n866 9.3005
R19273 vdd.n1941 vdd.n1940 9.3005
R19274 vdd.n271 vdd.n270 9.3005
R19275 vdd.n266 vdd.n265 9.3005
R19276 vdd.n277 vdd.n276 9.3005
R19277 vdd.n279 vdd.n278 9.3005
R19278 vdd.n262 vdd.n261 9.3005
R19279 vdd.n285 vdd.n284 9.3005
R19280 vdd.n287 vdd.n286 9.3005
R19281 vdd.n259 vdd.n256 9.3005
R19282 vdd.n294 vdd.n293 9.3005
R19283 vdd.n224 vdd.n223 9.3005
R19284 vdd.n219 vdd.n218 9.3005
R19285 vdd.n230 vdd.n229 9.3005
R19286 vdd.n232 vdd.n231 9.3005
R19287 vdd.n215 vdd.n214 9.3005
R19288 vdd.n238 vdd.n237 9.3005
R19289 vdd.n240 vdd.n239 9.3005
R19290 vdd.n212 vdd.n209 9.3005
R19291 vdd.n247 vdd.n246 9.3005
R19292 vdd.n181 vdd.n180 9.3005
R19293 vdd.n176 vdd.n175 9.3005
R19294 vdd.n187 vdd.n186 9.3005
R19295 vdd.n189 vdd.n188 9.3005
R19296 vdd.n172 vdd.n171 9.3005
R19297 vdd.n195 vdd.n194 9.3005
R19298 vdd.n197 vdd.n196 9.3005
R19299 vdd.n169 vdd.n166 9.3005
R19300 vdd.n204 vdd.n203 9.3005
R19301 vdd.n134 vdd.n133 9.3005
R19302 vdd.n129 vdd.n128 9.3005
R19303 vdd.n140 vdd.n139 9.3005
R19304 vdd.n142 vdd.n141 9.3005
R19305 vdd.n125 vdd.n124 9.3005
R19306 vdd.n148 vdd.n147 9.3005
R19307 vdd.n150 vdd.n149 9.3005
R19308 vdd.n122 vdd.n119 9.3005
R19309 vdd.n157 vdd.n156 9.3005
R19310 vdd.n92 vdd.n91 9.3005
R19311 vdd.n87 vdd.n86 9.3005
R19312 vdd.n98 vdd.n97 9.3005
R19313 vdd.n100 vdd.n99 9.3005
R19314 vdd.n83 vdd.n82 9.3005
R19315 vdd.n106 vdd.n105 9.3005
R19316 vdd.n108 vdd.n107 9.3005
R19317 vdd.n80 vdd.n77 9.3005
R19318 vdd.n115 vdd.n114 9.3005
R19319 vdd.n45 vdd.n44 9.3005
R19320 vdd.n40 vdd.n39 9.3005
R19321 vdd.n51 vdd.n50 9.3005
R19322 vdd.n53 vdd.n52 9.3005
R19323 vdd.n36 vdd.n35 9.3005
R19324 vdd.n59 vdd.n58 9.3005
R19325 vdd.n61 vdd.n60 9.3005
R19326 vdd.n33 vdd.n30 9.3005
R19327 vdd.n68 vdd.n67 9.3005
R19328 vdd.n2758 vdd.n2757 9.3005
R19329 vdd.n2761 vdd.n555 9.3005
R19330 vdd.n2762 vdd.n554 9.3005
R19331 vdd.n2765 vdd.n553 9.3005
R19332 vdd.n2766 vdd.n552 9.3005
R19333 vdd.n2769 vdd.n551 9.3005
R19334 vdd.n2770 vdd.n550 9.3005
R19335 vdd.n2773 vdd.n549 9.3005
R19336 vdd.n2774 vdd.n548 9.3005
R19337 vdd.n2777 vdd.n547 9.3005
R19338 vdd.n2778 vdd.n546 9.3005
R19339 vdd.n2781 vdd.n545 9.3005
R19340 vdd.n2782 vdd.n544 9.3005
R19341 vdd.n2785 vdd.n543 9.3005
R19342 vdd.n2786 vdd.n542 9.3005
R19343 vdd.n2789 vdd.n541 9.3005
R19344 vdd.n2790 vdd.n540 9.3005
R19345 vdd.n2793 vdd.n539 9.3005
R19346 vdd.n2794 vdd.n538 9.3005
R19347 vdd.n2797 vdd.n537 9.3005
R19348 vdd.n2801 vdd.n2800 9.3005
R19349 vdd.n2802 vdd.n536 9.3005
R19350 vdd.n2806 vdd.n2803 9.3005
R19351 vdd.n2809 vdd.n535 9.3005
R19352 vdd.n2810 vdd.n534 9.3005
R19353 vdd.n2813 vdd.n533 9.3005
R19354 vdd.n2814 vdd.n532 9.3005
R19355 vdd.n2817 vdd.n531 9.3005
R19356 vdd.n2818 vdd.n530 9.3005
R19357 vdd.n2821 vdd.n529 9.3005
R19358 vdd.n2822 vdd.n528 9.3005
R19359 vdd.n2825 vdd.n527 9.3005
R19360 vdd.n2826 vdd.n526 9.3005
R19361 vdd.n2829 vdd.n525 9.3005
R19362 vdd.n2830 vdd.n524 9.3005
R19363 vdd.n2833 vdd.n519 9.3005
R19364 vdd.n482 vdd.n481 9.3005
R19365 vdd.n2844 vdd.n2843 9.3005
R19366 vdd.n2847 vdd.n2846 9.3005
R19367 vdd.n471 vdd.n470 9.3005
R19368 vdd.n2861 vdd.n2860 9.3005
R19369 vdd.n2862 vdd.n469 9.3005
R19370 vdd.n2864 vdd.n2863 9.3005
R19371 vdd.n460 vdd.n459 9.3005
R19372 vdd.n2877 vdd.n2876 9.3005
R19373 vdd.n2878 vdd.n458 9.3005
R19374 vdd.n2880 vdd.n2879 9.3005
R19375 vdd.n300 vdd.n298 9.3005
R19376 vdd.n2845 vdd.n480 9.3005
R19377 vdd.n3046 vdd.n3045 9.3005
R19378 vdd.n301 vdd.n299 9.3005
R19379 vdd.n3039 vdd.n310 9.3005
R19380 vdd.n3038 vdd.n311 9.3005
R19381 vdd.n3037 vdd.n312 9.3005
R19382 vdd.n320 vdd.n313 9.3005
R19383 vdd.n3031 vdd.n321 9.3005
R19384 vdd.n3030 vdd.n322 9.3005
R19385 vdd.n3029 vdd.n323 9.3005
R19386 vdd.n331 vdd.n324 9.3005
R19387 vdd.n3023 vdd.n3022 9.3005
R19388 vdd.n3019 vdd.n332 9.3005
R19389 vdd.n3018 vdd.n335 9.3005
R19390 vdd.n339 vdd.n336 9.3005
R19391 vdd.n340 vdd.n337 9.3005
R19392 vdd.n3011 vdd.n341 9.3005
R19393 vdd.n3010 vdd.n342 9.3005
R19394 vdd.n3009 vdd.n343 9.3005
R19395 vdd.n347 vdd.n344 9.3005
R19396 vdd.n3004 vdd.n348 9.3005
R19397 vdd.n3003 vdd.n349 9.3005
R19398 vdd.n3002 vdd.n350 9.3005
R19399 vdd.n354 vdd.n351 9.3005
R19400 vdd.n2997 vdd.n355 9.3005
R19401 vdd.n2996 vdd.n356 9.3005
R19402 vdd.n2995 vdd.n357 9.3005
R19403 vdd.n361 vdd.n358 9.3005
R19404 vdd.n2990 vdd.n362 9.3005
R19405 vdd.n2989 vdd.n363 9.3005
R19406 vdd.n2988 vdd.n2987 9.3005
R19407 vdd.n2986 vdd.n364 9.3005
R19408 vdd.n2985 vdd.n2984 9.3005
R19409 vdd.n370 vdd.n369 9.3005
R19410 vdd.n2979 vdd.n374 9.3005
R19411 vdd.n2978 vdd.n375 9.3005
R19412 vdd.n2977 vdd.n376 9.3005
R19413 vdd.n380 vdd.n377 9.3005
R19414 vdd.n2972 vdd.n381 9.3005
R19415 vdd.n2971 vdd.n382 9.3005
R19416 vdd.n2970 vdd.n383 9.3005
R19417 vdd.n387 vdd.n384 9.3005
R19418 vdd.n2965 vdd.n388 9.3005
R19419 vdd.n2964 vdd.n389 9.3005
R19420 vdd.n2963 vdd.n390 9.3005
R19421 vdd.n394 vdd.n391 9.3005
R19422 vdd.n2958 vdd.n395 9.3005
R19423 vdd.n2957 vdd.n396 9.3005
R19424 vdd.n2956 vdd.n397 9.3005
R19425 vdd.n401 vdd.n398 9.3005
R19426 vdd.n2951 vdd.n402 9.3005
R19427 vdd.n2950 vdd.n403 9.3005
R19428 vdd.n2949 vdd.n2948 9.3005
R19429 vdd.n2947 vdd.n404 9.3005
R19430 vdd.n2946 vdd.n2945 9.3005
R19431 vdd.n410 vdd.n409 9.3005
R19432 vdd.n2940 vdd.n414 9.3005
R19433 vdd.n2939 vdd.n415 9.3005
R19434 vdd.n2938 vdd.n416 9.3005
R19435 vdd.n420 vdd.n417 9.3005
R19436 vdd.n2933 vdd.n421 9.3005
R19437 vdd.n2932 vdd.n422 9.3005
R19438 vdd.n2931 vdd.n423 9.3005
R19439 vdd.n427 vdd.n424 9.3005
R19440 vdd.n2926 vdd.n428 9.3005
R19441 vdd.n2925 vdd.n429 9.3005
R19442 vdd.n2924 vdd.n430 9.3005
R19443 vdd.n434 vdd.n431 9.3005
R19444 vdd.n2919 vdd.n435 9.3005
R19445 vdd.n2918 vdd.n436 9.3005
R19446 vdd.n2917 vdd.n437 9.3005
R19447 vdd.n441 vdd.n438 9.3005
R19448 vdd.n2912 vdd.n442 9.3005
R19449 vdd.n2911 vdd.n443 9.3005
R19450 vdd.n2907 vdd.n2904 9.3005
R19451 vdd.n3021 vdd.n3020 9.3005
R19452 vdd.n2852 vdd.n2851 9.3005
R19453 vdd.n2853 vdd.n475 9.3005
R19454 vdd.n2855 vdd.n2854 9.3005
R19455 vdd.n465 vdd.n464 9.3005
R19456 vdd.n2869 vdd.n2868 9.3005
R19457 vdd.n2870 vdd.n463 9.3005
R19458 vdd.n2872 vdd.n2871 9.3005
R19459 vdd.n453 vdd.n452 9.3005
R19460 vdd.n2885 vdd.n2884 9.3005
R19461 vdd.n2886 vdd.n451 9.3005
R19462 vdd.n2888 vdd.n2887 9.3005
R19463 vdd.n2889 vdd.n450 9.3005
R19464 vdd.n2891 vdd.n2890 9.3005
R19465 vdd.n2892 vdd.n449 9.3005
R19466 vdd.n2894 vdd.n2893 9.3005
R19467 vdd.n2895 vdd.n447 9.3005
R19468 vdd.n2897 vdd.n2896 9.3005
R19469 vdd.n2898 vdd.n446 9.3005
R19470 vdd.n2900 vdd.n2899 9.3005
R19471 vdd.n2901 vdd.n444 9.3005
R19472 vdd.n2903 vdd.n2902 9.3005
R19473 vdd.n477 vdd.n476 9.3005
R19474 vdd.n2710 vdd.n2709 9.3005
R19475 vdd.n2715 vdd.n2708 9.3005
R19476 vdd.n2724 vdd.n572 9.3005
R19477 vdd.n2727 vdd.n571 9.3005
R19478 vdd.n2728 vdd.n570 9.3005
R19479 vdd.n2731 vdd.n569 9.3005
R19480 vdd.n2732 vdd.n568 9.3005
R19481 vdd.n2735 vdd.n567 9.3005
R19482 vdd.n2736 vdd.n566 9.3005
R19483 vdd.n2739 vdd.n565 9.3005
R19484 vdd.n2740 vdd.n564 9.3005
R19485 vdd.n2743 vdd.n563 9.3005
R19486 vdd.n2744 vdd.n562 9.3005
R19487 vdd.n2747 vdd.n561 9.3005
R19488 vdd.n2748 vdd.n560 9.3005
R19489 vdd.n2751 vdd.n559 9.3005
R19490 vdd.n2755 vdd.n2754 9.3005
R19491 vdd.n2756 vdd.n556 9.3005
R19492 vdd.n1951 vdd.n1950 9.3005
R19493 vdd.n1946 vdd.n857 9.3005
R19494 vdd.n1433 vdd.n1432 9.3005
R19495 vdd.n1434 vdd.n1188 9.3005
R19496 vdd.n1436 vdd.n1435 9.3005
R19497 vdd.n1178 vdd.n1177 9.3005
R19498 vdd.n1450 vdd.n1449 9.3005
R19499 vdd.n1451 vdd.n1176 9.3005
R19500 vdd.n1453 vdd.n1452 9.3005
R19501 vdd.n1168 vdd.n1167 9.3005
R19502 vdd.n1468 vdd.n1467 9.3005
R19503 vdd.n1469 vdd.n1166 9.3005
R19504 vdd.n1471 vdd.n1470 9.3005
R19505 vdd.n885 vdd.n884 9.3005
R19506 vdd.n1484 vdd.n1483 9.3005
R19507 vdd.n1485 vdd.n883 9.3005
R19508 vdd.n1487 vdd.n1486 9.3005
R19509 vdd.n875 vdd.n874 9.3005
R19510 vdd.n1501 vdd.n1500 9.3005
R19511 vdd.n1502 vdd.n872 9.3005
R19512 vdd.n1506 vdd.n1505 9.3005
R19513 vdd.n1504 vdd.n873 9.3005
R19514 vdd.n1503 vdd.n862 9.3005
R19515 vdd.n1190 vdd.n1189 9.3005
R19516 vdd.n1326 vdd.n1325 9.3005
R19517 vdd.n1327 vdd.n1316 9.3005
R19518 vdd.n1329 vdd.n1328 9.3005
R19519 vdd.n1330 vdd.n1315 9.3005
R19520 vdd.n1332 vdd.n1331 9.3005
R19521 vdd.n1333 vdd.n1310 9.3005
R19522 vdd.n1335 vdd.n1334 9.3005
R19523 vdd.n1336 vdd.n1309 9.3005
R19524 vdd.n1338 vdd.n1337 9.3005
R19525 vdd.n1339 vdd.n1304 9.3005
R19526 vdd.n1341 vdd.n1340 9.3005
R19527 vdd.n1342 vdd.n1303 9.3005
R19528 vdd.n1344 vdd.n1343 9.3005
R19529 vdd.n1345 vdd.n1298 9.3005
R19530 vdd.n1347 vdd.n1346 9.3005
R19531 vdd.n1348 vdd.n1297 9.3005
R19532 vdd.n1350 vdd.n1349 9.3005
R19533 vdd.n1351 vdd.n1292 9.3005
R19534 vdd.n1353 vdd.n1352 9.3005
R19535 vdd.n1354 vdd.n1291 9.3005
R19536 vdd.n1356 vdd.n1355 9.3005
R19537 vdd.n1360 vdd.n1287 9.3005
R19538 vdd.n1362 vdd.n1361 9.3005
R19539 vdd.n1363 vdd.n1286 9.3005
R19540 vdd.n1365 vdd.n1364 9.3005
R19541 vdd.n1366 vdd.n1281 9.3005
R19542 vdd.n1368 vdd.n1367 9.3005
R19543 vdd.n1369 vdd.n1280 9.3005
R19544 vdd.n1371 vdd.n1370 9.3005
R19545 vdd.n1372 vdd.n1275 9.3005
R19546 vdd.n1374 vdd.n1373 9.3005
R19547 vdd.n1375 vdd.n1274 9.3005
R19548 vdd.n1377 vdd.n1376 9.3005
R19549 vdd.n1378 vdd.n1269 9.3005
R19550 vdd.n1380 vdd.n1379 9.3005
R19551 vdd.n1381 vdd.n1268 9.3005
R19552 vdd.n1383 vdd.n1382 9.3005
R19553 vdd.n1384 vdd.n1263 9.3005
R19554 vdd.n1386 vdd.n1385 9.3005
R19555 vdd.n1387 vdd.n1262 9.3005
R19556 vdd.n1389 vdd.n1388 9.3005
R19557 vdd.n1390 vdd.n1257 9.3005
R19558 vdd.n1392 vdd.n1391 9.3005
R19559 vdd.n1393 vdd.n1256 9.3005
R19560 vdd.n1395 vdd.n1394 9.3005
R19561 vdd.n1396 vdd.n1249 9.3005
R19562 vdd.n1398 vdd.n1397 9.3005
R19563 vdd.n1399 vdd.n1248 9.3005
R19564 vdd.n1401 vdd.n1400 9.3005
R19565 vdd.n1402 vdd.n1243 9.3005
R19566 vdd.n1404 vdd.n1403 9.3005
R19567 vdd.n1405 vdd.n1242 9.3005
R19568 vdd.n1407 vdd.n1406 9.3005
R19569 vdd.n1408 vdd.n1237 9.3005
R19570 vdd.n1410 vdd.n1409 9.3005
R19571 vdd.n1411 vdd.n1236 9.3005
R19572 vdd.n1413 vdd.n1412 9.3005
R19573 vdd.n1414 vdd.n1231 9.3005
R19574 vdd.n1416 vdd.n1415 9.3005
R19575 vdd.n1417 vdd.n1230 9.3005
R19576 vdd.n1419 vdd.n1418 9.3005
R19577 vdd.n1195 vdd.n1194 9.3005
R19578 vdd.n1425 vdd.n1424 9.3005
R19579 vdd.n1324 vdd.n1323 9.3005
R19580 vdd.n1428 vdd.n1427 9.3005
R19581 vdd.n1184 vdd.n1183 9.3005
R19582 vdd.n1442 vdd.n1441 9.3005
R19583 vdd.n1443 vdd.n1182 9.3005
R19584 vdd.n1445 vdd.n1444 9.3005
R19585 vdd.n1173 vdd.n1172 9.3005
R19586 vdd.n1459 vdd.n1458 9.3005
R19587 vdd.n1460 vdd.n1171 9.3005
R19588 vdd.n1463 vdd.n1462 9.3005
R19589 vdd.n1461 vdd.n1162 9.3005
R19590 vdd.n1426 vdd.n1193 9.3005
R19591 vdd.n1086 vdd.n1085 9.3005
R19592 vdd.n1081 vdd.n1080 9.3005
R19593 vdd.n1092 vdd.n1091 9.3005
R19594 vdd.n1094 vdd.n1093 9.3005
R19595 vdd.n1077 vdd.n1076 9.3005
R19596 vdd.n1100 vdd.n1099 9.3005
R19597 vdd.n1102 vdd.n1101 9.3005
R19598 vdd.n1074 vdd.n1071 9.3005
R19599 vdd.n1109 vdd.n1108 9.3005
R19600 vdd.n1133 vdd.n1132 9.3005
R19601 vdd.n1128 vdd.n1127 9.3005
R19602 vdd.n1139 vdd.n1138 9.3005
R19603 vdd.n1141 vdd.n1140 9.3005
R19604 vdd.n1124 vdd.n1123 9.3005
R19605 vdd.n1147 vdd.n1146 9.3005
R19606 vdd.n1149 vdd.n1148 9.3005
R19607 vdd.n1121 vdd.n1118 9.3005
R19608 vdd.n1156 vdd.n1155 9.3005
R19609 vdd.n996 vdd.n995 9.3005
R19610 vdd.n991 vdd.n990 9.3005
R19611 vdd.n1002 vdd.n1001 9.3005
R19612 vdd.n1004 vdd.n1003 9.3005
R19613 vdd.n987 vdd.n986 9.3005
R19614 vdd.n1010 vdd.n1009 9.3005
R19615 vdd.n1012 vdd.n1011 9.3005
R19616 vdd.n984 vdd.n981 9.3005
R19617 vdd.n1019 vdd.n1018 9.3005
R19618 vdd.n1043 vdd.n1042 9.3005
R19619 vdd.n1038 vdd.n1037 9.3005
R19620 vdd.n1049 vdd.n1048 9.3005
R19621 vdd.n1051 vdd.n1050 9.3005
R19622 vdd.n1034 vdd.n1033 9.3005
R19623 vdd.n1057 vdd.n1056 9.3005
R19624 vdd.n1059 vdd.n1058 9.3005
R19625 vdd.n1031 vdd.n1028 9.3005
R19626 vdd.n1066 vdd.n1065 9.3005
R19627 vdd.n907 vdd.n906 9.3005
R19628 vdd.n902 vdd.n901 9.3005
R19629 vdd.n913 vdd.n912 9.3005
R19630 vdd.n915 vdd.n914 9.3005
R19631 vdd.n898 vdd.n897 9.3005
R19632 vdd.n921 vdd.n920 9.3005
R19633 vdd.n923 vdd.n922 9.3005
R19634 vdd.n895 vdd.n892 9.3005
R19635 vdd.n930 vdd.n929 9.3005
R19636 vdd.n954 vdd.n953 9.3005
R19637 vdd.n949 vdd.n948 9.3005
R19638 vdd.n960 vdd.n959 9.3005
R19639 vdd.n962 vdd.n961 9.3005
R19640 vdd.n945 vdd.n944 9.3005
R19641 vdd.n968 vdd.n967 9.3005
R19642 vdd.n970 vdd.n969 9.3005
R19643 vdd.n942 vdd.n939 9.3005
R19644 vdd.n977 vdd.n976 9.3005
R19645 vdd.n1438 vdd.t47 8.95635
R19646 vdd.t29 vdd.n3033 8.95635
R19647 vdd.n276 vdd.n275 8.92171
R19648 vdd.n229 vdd.n228 8.92171
R19649 vdd.n186 vdd.n185 8.92171
R19650 vdd.n139 vdd.n138 8.92171
R19651 vdd.n97 vdd.n96 8.92171
R19652 vdd.n50 vdd.n49 8.92171
R19653 vdd.n1091 vdd.n1090 8.92171
R19654 vdd.n1138 vdd.n1137 8.92171
R19655 vdd.n1001 vdd.n1000 8.92171
R19656 vdd.n1048 vdd.n1047 8.92171
R19657 vdd.n912 vdd.n911 8.92171
R19658 vdd.n959 vdd.n958 8.92171
R19659 vdd.n207 vdd.n117 8.81535
R19660 vdd.n1069 vdd.n979 8.81535
R19661 vdd.n1465 vdd.t25 8.72962
R19662 vdd.t27 vdd.n3042 8.72962
R19663 vdd.n888 vdd.t63 8.50289
R19664 vdd.n1943 vdd.t89 8.50289
R19665 vdd.n516 vdd.t82 8.50289
R19666 vdd.n2874 vdd.t41 8.50289
R19667 vdd.n28 vdd.n14 8.42249
R19668 vdd.n3048 vdd.n3047 8.16225
R19669 vdd.n1161 vdd.n1160 8.16225
R19670 vdd.n272 vdd.n266 8.14595
R19671 vdd.n225 vdd.n219 8.14595
R19672 vdd.n182 vdd.n176 8.14595
R19673 vdd.n135 vdd.n129 8.14595
R19674 vdd.n93 vdd.n87 8.14595
R19675 vdd.n46 vdd.n40 8.14595
R19676 vdd.n1087 vdd.n1081 8.14595
R19677 vdd.n1134 vdd.n1128 8.14595
R19678 vdd.n997 vdd.n991 8.14595
R19679 vdd.n1044 vdd.n1038 8.14595
R19680 vdd.n908 vdd.n902 8.14595
R19681 vdd.n955 vdd.n949 8.14595
R19682 vdd.n2537 vdd.n639 8.11757
R19683 vdd.n2011 vdd.n2010 8.11757
R19684 vdd.n1989 vdd.n833 7.70933
R19685 vdd.n1995 vdd.n833 7.70933
R19686 vdd.n2001 vdd.n827 7.70933
R19687 vdd.n2001 vdd.n820 7.70933
R19688 vdd.n2007 vdd.n820 7.70933
R19689 vdd.n2007 vdd.n823 7.70933
R19690 vdd.n2014 vdd.n808 7.70933
R19691 vdd.n2020 vdd.n808 7.70933
R19692 vdd.n2026 vdd.n802 7.70933
R19693 vdd.n2032 vdd.n798 7.70933
R19694 vdd.n2038 vdd.n792 7.70933
R19695 vdd.n2050 vdd.n779 7.70933
R19696 vdd.n2056 vdd.n773 7.70933
R19697 vdd.n2056 vdd.n766 7.70933
R19698 vdd.n2064 vdd.n766 7.70933
R19699 vdd.n2071 vdd.t2 7.70933
R19700 vdd.n2146 vdd.t2 7.70933
R19701 vdd.n2478 vdd.t198 7.70933
R19702 vdd.n2484 vdd.t198 7.70933
R19703 vdd.n2490 vdd.n687 7.70933
R19704 vdd.n2496 vdd.n687 7.70933
R19705 vdd.n2496 vdd.n690 7.70933
R19706 vdd.n2502 vdd.n683 7.70933
R19707 vdd.n2514 vdd.n670 7.70933
R19708 vdd.n2520 vdd.n664 7.70933
R19709 vdd.n2526 vdd.n660 7.70933
R19710 vdd.n2532 vdd.n647 7.70933
R19711 vdd.n2540 vdd.n647 7.70933
R19712 vdd.n2546 vdd.n641 7.70933
R19713 vdd.n2546 vdd.n633 7.70933
R19714 vdd.n2597 vdd.n633 7.70933
R19715 vdd.n2597 vdd.n636 7.70933
R19716 vdd.n2603 vdd.n595 7.70933
R19717 vdd.n2673 vdd.n595 7.70933
R19718 vdd.n271 vdd.n268 7.3702
R19719 vdd.n224 vdd.n221 7.3702
R19720 vdd.n181 vdd.n178 7.3702
R19721 vdd.n134 vdd.n131 7.3702
R19722 vdd.n92 vdd.n89 7.3702
R19723 vdd.n45 vdd.n42 7.3702
R19724 vdd.n1086 vdd.n1083 7.3702
R19725 vdd.n1133 vdd.n1130 7.3702
R19726 vdd.n996 vdd.n993 7.3702
R19727 vdd.n1043 vdd.n1040 7.3702
R19728 vdd.n907 vdd.n904 7.3702
R19729 vdd.n954 vdd.n951 7.3702
R19730 vdd.n1361 vdd.n1360 6.98232
R19731 vdd.n1653 vdd.n1652 6.98232
R19732 vdd.n2950 vdd.n2949 6.98232
R19733 vdd.n2761 vdd.n2758 6.98232
R19734 vdd.n1498 vdd.t10 6.68904
R19735 vdd.n2857 vdd.t12 6.68904
R19736 vdd.t49 vdd.n887 6.46231
R19737 vdd.n2882 vdd.t16 6.46231
R19738 vdd.n1456 vdd.t31 6.23558
R19739 vdd.t20 vdd.n308 6.23558
R19740 vdd.n3048 vdd.n297 6.22547
R19741 vdd.n1160 vdd.n1159 6.22547
R19742 vdd.n2026 vdd.t185 6.00885
R19743 vdd.n2526 vdd.t178 6.00885
R19744 vdd.n823 vdd.t133 5.89549
R19745 vdd.t97 vdd.n641 5.89549
R19746 vdd.n272 vdd.n271 5.81868
R19747 vdd.n225 vdd.n224 5.81868
R19748 vdd.n182 vdd.n181 5.81868
R19749 vdd.n135 vdd.n134 5.81868
R19750 vdd.n93 vdd.n92 5.81868
R19751 vdd.n46 vdd.n45 5.81868
R19752 vdd.n1087 vdd.n1086 5.81868
R19753 vdd.n1134 vdd.n1133 5.81868
R19754 vdd.n997 vdd.n996 5.81868
R19755 vdd.n1044 vdd.n1043 5.81868
R19756 vdd.n908 vdd.n907 5.81868
R19757 vdd.n955 vdd.n954 5.81868
R19758 vdd.t129 vdd.n827 5.78212
R19759 vdd.n1770 vdd.t114 5.78212
R19760 vdd.n2395 vdd.t122 5.78212
R19761 vdd.n636 vdd.t118 5.78212
R19762 vdd.n2154 vdd.n2153 5.77611
R19763 vdd.n1897 vdd.n1767 5.77611
R19764 vdd.n2408 vdd.n2407 5.77611
R19765 vdd.n2614 vdd.n2613 5.77611
R19766 vdd.n2678 vdd.n591 5.77611
R19767 vdd.n2318 vdd.n2258 5.77611
R19768 vdd.n2079 vdd.n757 5.77611
R19769 vdd.n1827 vdd.n1826 5.77611
R19770 vdd.n1323 vdd.n1322 5.62474
R19771 vdd.n1949 vdd.n1946 5.62474
R19772 vdd.n2910 vdd.n2907 5.62474
R19773 vdd.n2713 vdd.n2710 5.62474
R19774 vdd.t183 vdd.n779 5.44203
R19775 vdd.n683 vdd.t179 5.44203
R19776 vdd.n1180 vdd.t31 5.10193
R19777 vdd.t175 vdd.n802 5.10193
R19778 vdd.n792 vdd.t9 5.10193
R19779 vdd.t6 vdd.n670 5.10193
R19780 vdd.n660 vdd.t173 5.10193
R19781 vdd.n3035 vdd.t20 5.10193
R19782 vdd.n275 vdd.n266 5.04292
R19783 vdd.n228 vdd.n219 5.04292
R19784 vdd.n185 vdd.n176 5.04292
R19785 vdd.n138 vdd.n129 5.04292
R19786 vdd.n96 vdd.n87 5.04292
R19787 vdd.n49 vdd.n40 5.04292
R19788 vdd.n1090 vdd.n1081 5.04292
R19789 vdd.n1137 vdd.n1128 5.04292
R19790 vdd.n1000 vdd.n991 5.04292
R19791 vdd.n1047 vdd.n1038 5.04292
R19792 vdd.n911 vdd.n902 5.04292
R19793 vdd.n958 vdd.n949 5.04292
R19794 vdd.n1473 vdd.t49 4.8752
R19795 vdd.t76 vdd.t176 4.8752
R19796 vdd.t191 vdd.t186 4.8752
R19797 vdd.t189 vdd.t78 4.8752
R19798 vdd.t194 vdd.t77 4.8752
R19799 vdd.t16 vdd.n304 4.8752
R19800 vdd.n2155 vdd.n2154 4.83952
R19801 vdd.n1767 vdd.n1763 4.83952
R19802 vdd.n2409 vdd.n2408 4.83952
R19803 vdd.n2615 vdd.n2614 4.83952
R19804 vdd.n591 vdd.n586 4.83952
R19805 vdd.n2315 vdd.n2258 4.83952
R19806 vdd.n2082 vdd.n757 4.83952
R19807 vdd.n1826 vdd.n1825 4.83952
R19808 vdd.n1621 vdd.n855 4.74817
R19809 vdd.n1616 vdd.n856 4.74817
R19810 vdd.n1518 vdd.n1515 4.74817
R19811 vdd.n1930 vdd.n1519 4.74817
R19812 vdd.n1932 vdd.n1518 4.74817
R19813 vdd.n1931 vdd.n1930 4.74817
R19814 vdd.n2838 vdd.n2837 4.74817
R19815 vdd.n2835 vdd.n2834 4.74817
R19816 vdd.n2835 vdd.n521 4.74817
R19817 vdd.n2837 vdd.n518 4.74817
R19818 vdd.n2720 vdd.n573 4.74817
R19819 vdd.n2716 vdd.n574 4.74817
R19820 vdd.n2719 vdd.n574 4.74817
R19821 vdd.n2723 vdd.n573 4.74817
R19822 vdd.n1617 vdd.n855 4.74817
R19823 vdd.n858 vdd.n856 4.74817
R19824 vdd.n297 vdd.n296 4.7074
R19825 vdd.n207 vdd.n206 4.7074
R19826 vdd.n1159 vdd.n1158 4.7074
R19827 vdd.n1069 vdd.n1068 4.7074
R19828 vdd.n1489 vdd.t10 4.64847
R19829 vdd.n2866 vdd.t12 4.64847
R19830 vdd.n2032 vdd.t192 4.53511
R19831 vdd.n2520 vdd.t0 4.53511
R19832 vdd.n2064 vdd.t74 4.30838
R19833 vdd.n2490 vdd.t7 4.30838
R19834 vdd.n276 vdd.n264 4.26717
R19835 vdd.n229 vdd.n217 4.26717
R19836 vdd.n186 vdd.n174 4.26717
R19837 vdd.n139 vdd.n127 4.26717
R19838 vdd.n97 vdd.n85 4.26717
R19839 vdd.n50 vdd.n38 4.26717
R19840 vdd.n1091 vdd.n1079 4.26717
R19841 vdd.n1138 vdd.n1126 4.26717
R19842 vdd.n1001 vdd.n989 4.26717
R19843 vdd.n1048 vdd.n1036 4.26717
R19844 vdd.n912 vdd.n900 4.26717
R19845 vdd.n959 vdd.n947 4.26717
R19846 vdd.n297 vdd.n207 4.10845
R19847 vdd.n1159 vdd.n1069 4.10845
R19848 vdd.n253 vdd.t57 4.06363
R19849 vdd.n253 vdd.t21 4.06363
R19850 vdd.n251 vdd.t23 4.06363
R19851 vdd.n251 vdd.t44 4.06363
R19852 vdd.n249 vdd.t46 4.06363
R19853 vdd.n249 vdd.t62 4.06363
R19854 vdd.n163 vdd.t52 4.06363
R19855 vdd.n163 vdd.t73 4.06363
R19856 vdd.n161 vdd.t17 4.06363
R19857 vdd.n161 vdd.t36 4.06363
R19858 vdd.n159 vdd.t42 4.06363
R19859 vdd.n159 vdd.t53 4.06363
R19860 vdd.n74 vdd.t58 4.06363
R19861 vdd.n74 vdd.t33 4.06363
R19862 vdd.n72 vdd.t72 4.06363
R19863 vdd.n72 vdd.t28 4.06363
R19864 vdd.n70 vdd.t65 4.06363
R19865 vdd.n70 vdd.t39 4.06363
R19866 vdd.n1111 vdd.t24 4.06363
R19867 vdd.n1111 vdd.t68 4.06363
R19868 vdd.n1113 vdd.t67 4.06363
R19869 vdd.n1113 vdd.t56 4.06363
R19870 vdd.n1115 vdd.t43 4.06363
R19871 vdd.n1115 vdd.t22 4.06363
R19872 vdd.n1021 vdd.t19 4.06363
R19873 vdd.n1021 vdd.t64 4.06363
R19874 vdd.n1023 vdd.t59 4.06363
R19875 vdd.n1023 vdd.t50 4.06363
R19876 vdd.n1025 vdd.t35 4.06363
R19877 vdd.n1025 vdd.t15 4.06363
R19878 vdd.n932 vdd.t37 4.06363
R19879 vdd.n932 vdd.t66 4.06363
R19880 vdd.n934 vdd.t26 4.06363
R19881 vdd.n934 vdd.t54 4.06363
R19882 vdd.n936 vdd.t32 4.06363
R19883 vdd.n936 vdd.t60 4.06363
R19884 vdd.n26 vdd.t163 3.9605
R19885 vdd.n26 vdd.t162 3.9605
R19886 vdd.n23 vdd.t170 3.9605
R19887 vdd.n23 vdd.t169 3.9605
R19888 vdd.n21 vdd.t171 3.9605
R19889 vdd.n21 vdd.t164 3.9605
R19890 vdd.n20 vdd.t166 3.9605
R19891 vdd.n20 vdd.t167 3.9605
R19892 vdd.n15 vdd.t165 3.9605
R19893 vdd.n15 vdd.t168 3.9605
R19894 vdd.n16 vdd.t157 3.9605
R19895 vdd.n16 vdd.t158 3.9605
R19896 vdd.n18 vdd.t161 3.9605
R19897 vdd.n18 vdd.t160 3.9605
R19898 vdd.n25 vdd.t159 3.9605
R19899 vdd.n25 vdd.t172 3.9605
R19900 vdd.n7 vdd.t195 3.61217
R19901 vdd.n7 vdd.t1 3.61217
R19902 vdd.n8 vdd.t190 3.61217
R19903 vdd.n8 vdd.t180 3.61217
R19904 vdd.n10 vdd.t199 3.61217
R19905 vdd.n10 vdd.t8 3.61217
R19906 vdd.n12 vdd.t182 3.61217
R19907 vdd.n12 vdd.t197 3.61217
R19908 vdd.n5 vdd.t5 3.61217
R19909 vdd.n5 vdd.t80 3.61217
R19910 vdd.n3 vdd.t75 3.61217
R19911 vdd.n3 vdd.t3 3.61217
R19912 vdd.n1 vdd.t184 3.61217
R19913 vdd.n1 vdd.t187 3.61217
R19914 vdd.n0 vdd.t193 3.61217
R19915 vdd.n0 vdd.t177 3.61217
R19916 vdd.n280 vdd.n279 3.49141
R19917 vdd.n233 vdd.n232 3.49141
R19918 vdd.n190 vdd.n189 3.49141
R19919 vdd.n143 vdd.n142 3.49141
R19920 vdd.n101 vdd.n100 3.49141
R19921 vdd.n54 vdd.n53 3.49141
R19922 vdd.n1095 vdd.n1094 3.49141
R19923 vdd.n1142 vdd.n1141 3.49141
R19924 vdd.n1005 vdd.n1004 3.49141
R19925 vdd.n1052 vdd.n1051 3.49141
R19926 vdd.n916 vdd.n915 3.49141
R19927 vdd.n963 vdd.n962 3.49141
R19928 vdd.n1770 vdd.t74 3.40145
R19929 vdd.n2218 vdd.t4 3.40145
R19930 vdd.n2471 vdd.t196 3.40145
R19931 vdd.n2395 vdd.t7 3.40145
R19932 vdd.n1871 vdd.t192 3.17472
R19933 vdd.n2374 vdd.t0 3.17472
R19934 vdd.n1490 vdd.t63 2.83463
R19935 vdd.n1508 vdd.t89 2.83463
R19936 vdd.n2849 vdd.t82 2.83463
R19937 vdd.n467 vdd.t41 2.83463
R19938 vdd.n283 vdd.n262 2.71565
R19939 vdd.n236 vdd.n215 2.71565
R19940 vdd.n193 vdd.n172 2.71565
R19941 vdd.n146 vdd.n125 2.71565
R19942 vdd.n104 vdd.n83 2.71565
R19943 vdd.n57 vdd.n36 2.71565
R19944 vdd.n1098 vdd.n1077 2.71565
R19945 vdd.n1145 vdd.n1124 2.71565
R19946 vdd.n1008 vdd.n987 2.71565
R19947 vdd.n1055 vdd.n1034 2.71565
R19948 vdd.n919 vdd.n898 2.71565
R19949 vdd.n966 vdd.n945 2.71565
R19950 vdd.t25 vdd.n1164 2.6079
R19951 vdd.n2020 vdd.t175 2.6079
R19952 vdd.n2044 vdd.t9 2.6079
R19953 vdd.n2508 vdd.t6 2.6079
R19954 vdd.n2532 vdd.t173 2.6079
R19955 vdd.n3043 vdd.t27 2.6079
R19956 vdd.n2538 vdd.n2537 2.49806
R19957 vdd.n2012 vdd.n2011 2.49806
R19958 vdd.n270 vdd.n269 2.4129
R19959 vdd.n223 vdd.n222 2.4129
R19960 vdd.n180 vdd.n179 2.4129
R19961 vdd.n133 vdd.n132 2.4129
R19962 vdd.n91 vdd.n90 2.4129
R19963 vdd.n44 vdd.n43 2.4129
R19964 vdd.n1085 vdd.n1084 2.4129
R19965 vdd.n1132 vdd.n1131 2.4129
R19966 vdd.n995 vdd.n994 2.4129
R19967 vdd.n1042 vdd.n1041 2.4129
R19968 vdd.n906 vdd.n905 2.4129
R19969 vdd.n953 vdd.n952 2.4129
R19970 vdd.n1447 vdd.t47 2.38117
R19971 vdd.n3034 vdd.t29 2.38117
R19972 vdd.n1929 vdd.n1518 2.27742
R19973 vdd.n1930 vdd.n1929 2.27742
R19974 vdd.n2836 vdd.n2835 2.27742
R19975 vdd.n2837 vdd.n2836 2.27742
R19976 vdd.n2707 vdd.n574 2.27742
R19977 vdd.n2707 vdd.n573 2.27742
R19978 vdd.n1952 vdd.n855 2.27742
R19979 vdd.n1952 vdd.n856 2.27742
R19980 vdd.n2044 vdd.t183 2.2678
R19981 vdd.n2508 vdd.t179 2.2678
R19982 vdd.t186 vdd.n773 2.04107
R19983 vdd.n690 vdd.t189 2.04107
R19984 vdd.n284 vdd.n260 1.93989
R19985 vdd.n237 vdd.n213 1.93989
R19986 vdd.n194 vdd.n170 1.93989
R19987 vdd.n147 vdd.n123 1.93989
R19988 vdd.n105 vdd.n81 1.93989
R19989 vdd.n58 vdd.n34 1.93989
R19990 vdd.n1099 vdd.n1075 1.93989
R19991 vdd.n1146 vdd.n1122 1.93989
R19992 vdd.n1009 vdd.n985 1.93989
R19993 vdd.n1056 vdd.n1032 1.93989
R19994 vdd.n920 vdd.n896 1.93989
R19995 vdd.n967 vdd.n943 1.93989
R19996 vdd.n1995 vdd.t129 1.92771
R19997 vdd.n2071 vdd.t114 1.92771
R19998 vdd.n2484 vdd.t122 1.92771
R19999 vdd.n2603 vdd.t118 1.92771
R20000 vdd.n1871 vdd.t185 1.70098
R20001 vdd.n798 vdd.t76 1.70098
R20002 vdd.t77 vdd.n664 1.70098
R20003 vdd.n2374 vdd.t178 1.70098
R20004 vdd.n1455 vdd.t14 1.24752
R20005 vdd.t51 vdd.n3041 1.24752
R20006 vdd.n295 vdd.n255 1.16414
R20007 vdd.n288 vdd.n287 1.16414
R20008 vdd.n248 vdd.n208 1.16414
R20009 vdd.n241 vdd.n240 1.16414
R20010 vdd.n205 vdd.n165 1.16414
R20011 vdd.n198 vdd.n197 1.16414
R20012 vdd.n158 vdd.n118 1.16414
R20013 vdd.n151 vdd.n150 1.16414
R20014 vdd.n116 vdd.n76 1.16414
R20015 vdd.n109 vdd.n108 1.16414
R20016 vdd.n69 vdd.n29 1.16414
R20017 vdd.n62 vdd.n61 1.16414
R20018 vdd.n1110 vdd.n1070 1.16414
R20019 vdd.n1103 vdd.n1102 1.16414
R20020 vdd.n1157 vdd.n1117 1.16414
R20021 vdd.n1150 vdd.n1149 1.16414
R20022 vdd.n1020 vdd.n980 1.16414
R20023 vdd.n1013 vdd.n1012 1.16414
R20024 vdd.n1067 vdd.n1027 1.16414
R20025 vdd.n1060 vdd.n1059 1.16414
R20026 vdd.n931 vdd.n891 1.16414
R20027 vdd.n924 vdd.n923 1.16414
R20028 vdd.n978 vdd.n938 1.16414
R20029 vdd.n971 vdd.n970 1.16414
R20030 vdd.n2038 vdd.t176 1.13415
R20031 vdd.n2514 vdd.t194 1.13415
R20032 vdd.n1481 vdd.t18 1.02079
R20033 vdd.t133 vdd.t174 1.02079
R20034 vdd.t188 vdd.t97 1.02079
R20035 vdd.t38 vdd.n456 1.02079
R20036 vdd.n1326 vdd.n1322 0.970197
R20037 vdd.n1950 vdd.n1949 0.970197
R20038 vdd.n2911 vdd.n2910 0.970197
R20039 vdd.n2715 vdd.n2713 0.970197
R20040 vdd.n2014 vdd.t174 0.794056
R20041 vdd.n2050 vdd.t191 0.794056
R20042 vdd.n2502 vdd.t78 0.794056
R20043 vdd.n2540 vdd.t188 0.794056
R20044 vdd.n1160 vdd.n28 0.74827
R20045 vdd vdd.n3048 0.740437
R20046 vdd.n1430 vdd.t93 0.567326
R20047 vdd.n3026 vdd.t104 0.567326
R20048 vdd.n1940 vdd.n1939 0.537085
R20049 vdd.n2845 vdd.n2844 0.537085
R20050 vdd.n3022 vdd.n3021 0.537085
R20051 vdd.n2904 vdd.n2903 0.537085
R20052 vdd.n2709 vdd.n476 0.537085
R20053 vdd.n1503 vdd.n857 0.537085
R20054 vdd.n1324 vdd.n1189 0.537085
R20055 vdd.n1426 vdd.n1425 0.537085
R20056 vdd.n4 vdd.n2 0.459552
R20057 vdd.n11 vdd.n9 0.459552
R20058 vdd.n293 vdd.n292 0.388379
R20059 vdd.n259 vdd.n257 0.388379
R20060 vdd.n246 vdd.n245 0.388379
R20061 vdd.n212 vdd.n210 0.388379
R20062 vdd.n203 vdd.n202 0.388379
R20063 vdd.n169 vdd.n167 0.388379
R20064 vdd.n156 vdd.n155 0.388379
R20065 vdd.n122 vdd.n120 0.388379
R20066 vdd.n114 vdd.n113 0.388379
R20067 vdd.n80 vdd.n78 0.388379
R20068 vdd.n67 vdd.n66 0.388379
R20069 vdd.n33 vdd.n31 0.388379
R20070 vdd.n1108 vdd.n1107 0.388379
R20071 vdd.n1074 vdd.n1072 0.388379
R20072 vdd.n1155 vdd.n1154 0.388379
R20073 vdd.n1121 vdd.n1119 0.388379
R20074 vdd.n1018 vdd.n1017 0.388379
R20075 vdd.n984 vdd.n982 0.388379
R20076 vdd.n1065 vdd.n1064 0.388379
R20077 vdd.n1031 vdd.n1029 0.388379
R20078 vdd.n929 vdd.n928 0.388379
R20079 vdd.n895 vdd.n893 0.388379
R20080 vdd.n976 vdd.n975 0.388379
R20081 vdd.n942 vdd.n940 0.388379
R20082 vdd.n19 vdd.n17 0.387128
R20083 vdd.n24 vdd.n22 0.387128
R20084 vdd.n6 vdd.n4 0.358259
R20085 vdd.n13 vdd.n11 0.358259
R20086 vdd.n252 vdd.n250 0.358259
R20087 vdd.n254 vdd.n252 0.358259
R20088 vdd.n296 vdd.n254 0.358259
R20089 vdd.n162 vdd.n160 0.358259
R20090 vdd.n164 vdd.n162 0.358259
R20091 vdd.n206 vdd.n164 0.358259
R20092 vdd.n73 vdd.n71 0.358259
R20093 vdd.n75 vdd.n73 0.358259
R20094 vdd.n117 vdd.n75 0.358259
R20095 vdd.n1158 vdd.n1116 0.358259
R20096 vdd.n1116 vdd.n1114 0.358259
R20097 vdd.n1114 vdd.n1112 0.358259
R20098 vdd.n1068 vdd.n1026 0.358259
R20099 vdd.n1026 vdd.n1024 0.358259
R20100 vdd.n1024 vdd.n1022 0.358259
R20101 vdd.n979 vdd.n937 0.358259
R20102 vdd.n937 vdd.n935 0.358259
R20103 vdd.n935 vdd.n933 0.358259
R20104 vdd.n14 vdd.n6 0.334552
R20105 vdd.n14 vdd.n13 0.334552
R20106 vdd.n27 vdd.n19 0.21707
R20107 vdd.n27 vdd.n24 0.21707
R20108 vdd.n294 vdd.n256 0.155672
R20109 vdd.n286 vdd.n256 0.155672
R20110 vdd.n286 vdd.n285 0.155672
R20111 vdd.n285 vdd.n261 0.155672
R20112 vdd.n278 vdd.n261 0.155672
R20113 vdd.n278 vdd.n277 0.155672
R20114 vdd.n277 vdd.n265 0.155672
R20115 vdd.n270 vdd.n265 0.155672
R20116 vdd.n247 vdd.n209 0.155672
R20117 vdd.n239 vdd.n209 0.155672
R20118 vdd.n239 vdd.n238 0.155672
R20119 vdd.n238 vdd.n214 0.155672
R20120 vdd.n231 vdd.n214 0.155672
R20121 vdd.n231 vdd.n230 0.155672
R20122 vdd.n230 vdd.n218 0.155672
R20123 vdd.n223 vdd.n218 0.155672
R20124 vdd.n204 vdd.n166 0.155672
R20125 vdd.n196 vdd.n166 0.155672
R20126 vdd.n196 vdd.n195 0.155672
R20127 vdd.n195 vdd.n171 0.155672
R20128 vdd.n188 vdd.n171 0.155672
R20129 vdd.n188 vdd.n187 0.155672
R20130 vdd.n187 vdd.n175 0.155672
R20131 vdd.n180 vdd.n175 0.155672
R20132 vdd.n157 vdd.n119 0.155672
R20133 vdd.n149 vdd.n119 0.155672
R20134 vdd.n149 vdd.n148 0.155672
R20135 vdd.n148 vdd.n124 0.155672
R20136 vdd.n141 vdd.n124 0.155672
R20137 vdd.n141 vdd.n140 0.155672
R20138 vdd.n140 vdd.n128 0.155672
R20139 vdd.n133 vdd.n128 0.155672
R20140 vdd.n115 vdd.n77 0.155672
R20141 vdd.n107 vdd.n77 0.155672
R20142 vdd.n107 vdd.n106 0.155672
R20143 vdd.n106 vdd.n82 0.155672
R20144 vdd.n99 vdd.n82 0.155672
R20145 vdd.n99 vdd.n98 0.155672
R20146 vdd.n98 vdd.n86 0.155672
R20147 vdd.n91 vdd.n86 0.155672
R20148 vdd.n68 vdd.n30 0.155672
R20149 vdd.n60 vdd.n30 0.155672
R20150 vdd.n60 vdd.n59 0.155672
R20151 vdd.n59 vdd.n35 0.155672
R20152 vdd.n52 vdd.n35 0.155672
R20153 vdd.n52 vdd.n51 0.155672
R20154 vdd.n51 vdd.n39 0.155672
R20155 vdd.n44 vdd.n39 0.155672
R20156 vdd.n1109 vdd.n1071 0.155672
R20157 vdd.n1101 vdd.n1071 0.155672
R20158 vdd.n1101 vdd.n1100 0.155672
R20159 vdd.n1100 vdd.n1076 0.155672
R20160 vdd.n1093 vdd.n1076 0.155672
R20161 vdd.n1093 vdd.n1092 0.155672
R20162 vdd.n1092 vdd.n1080 0.155672
R20163 vdd.n1085 vdd.n1080 0.155672
R20164 vdd.n1156 vdd.n1118 0.155672
R20165 vdd.n1148 vdd.n1118 0.155672
R20166 vdd.n1148 vdd.n1147 0.155672
R20167 vdd.n1147 vdd.n1123 0.155672
R20168 vdd.n1140 vdd.n1123 0.155672
R20169 vdd.n1140 vdd.n1139 0.155672
R20170 vdd.n1139 vdd.n1127 0.155672
R20171 vdd.n1132 vdd.n1127 0.155672
R20172 vdd.n1019 vdd.n981 0.155672
R20173 vdd.n1011 vdd.n981 0.155672
R20174 vdd.n1011 vdd.n1010 0.155672
R20175 vdd.n1010 vdd.n986 0.155672
R20176 vdd.n1003 vdd.n986 0.155672
R20177 vdd.n1003 vdd.n1002 0.155672
R20178 vdd.n1002 vdd.n990 0.155672
R20179 vdd.n995 vdd.n990 0.155672
R20180 vdd.n1066 vdd.n1028 0.155672
R20181 vdd.n1058 vdd.n1028 0.155672
R20182 vdd.n1058 vdd.n1057 0.155672
R20183 vdd.n1057 vdd.n1033 0.155672
R20184 vdd.n1050 vdd.n1033 0.155672
R20185 vdd.n1050 vdd.n1049 0.155672
R20186 vdd.n1049 vdd.n1037 0.155672
R20187 vdd.n1042 vdd.n1037 0.155672
R20188 vdd.n930 vdd.n892 0.155672
R20189 vdd.n922 vdd.n892 0.155672
R20190 vdd.n922 vdd.n921 0.155672
R20191 vdd.n921 vdd.n897 0.155672
R20192 vdd.n914 vdd.n897 0.155672
R20193 vdd.n914 vdd.n913 0.155672
R20194 vdd.n913 vdd.n901 0.155672
R20195 vdd.n906 vdd.n901 0.155672
R20196 vdd.n977 vdd.n939 0.155672
R20197 vdd.n969 vdd.n939 0.155672
R20198 vdd.n969 vdd.n968 0.155672
R20199 vdd.n968 vdd.n944 0.155672
R20200 vdd.n961 vdd.n944 0.155672
R20201 vdd.n961 vdd.n960 0.155672
R20202 vdd.n960 vdd.n948 0.155672
R20203 vdd.n953 vdd.n948 0.155672
R20204 vdd.n1715 vdd.n1520 0.152939
R20205 vdd.n1526 vdd.n1520 0.152939
R20206 vdd.n1527 vdd.n1526 0.152939
R20207 vdd.n1528 vdd.n1527 0.152939
R20208 vdd.n1529 vdd.n1528 0.152939
R20209 vdd.n1533 vdd.n1529 0.152939
R20210 vdd.n1534 vdd.n1533 0.152939
R20211 vdd.n1535 vdd.n1534 0.152939
R20212 vdd.n1536 vdd.n1535 0.152939
R20213 vdd.n1540 vdd.n1536 0.152939
R20214 vdd.n1541 vdd.n1540 0.152939
R20215 vdd.n1542 vdd.n1541 0.152939
R20216 vdd.n1690 vdd.n1542 0.152939
R20217 vdd.n1690 vdd.n1689 0.152939
R20218 vdd.n1689 vdd.n1688 0.152939
R20219 vdd.n1688 vdd.n1548 0.152939
R20220 vdd.n1553 vdd.n1548 0.152939
R20221 vdd.n1554 vdd.n1553 0.152939
R20222 vdd.n1555 vdd.n1554 0.152939
R20223 vdd.n1559 vdd.n1555 0.152939
R20224 vdd.n1560 vdd.n1559 0.152939
R20225 vdd.n1561 vdd.n1560 0.152939
R20226 vdd.n1562 vdd.n1561 0.152939
R20227 vdd.n1566 vdd.n1562 0.152939
R20228 vdd.n1567 vdd.n1566 0.152939
R20229 vdd.n1568 vdd.n1567 0.152939
R20230 vdd.n1569 vdd.n1568 0.152939
R20231 vdd.n1573 vdd.n1569 0.152939
R20232 vdd.n1574 vdd.n1573 0.152939
R20233 vdd.n1575 vdd.n1574 0.152939
R20234 vdd.n1576 vdd.n1575 0.152939
R20235 vdd.n1580 vdd.n1576 0.152939
R20236 vdd.n1581 vdd.n1580 0.152939
R20237 vdd.n1582 vdd.n1581 0.152939
R20238 vdd.n1651 vdd.n1582 0.152939
R20239 vdd.n1651 vdd.n1650 0.152939
R20240 vdd.n1650 vdd.n1649 0.152939
R20241 vdd.n1649 vdd.n1588 0.152939
R20242 vdd.n1593 vdd.n1588 0.152939
R20243 vdd.n1594 vdd.n1593 0.152939
R20244 vdd.n1595 vdd.n1594 0.152939
R20245 vdd.n1599 vdd.n1595 0.152939
R20246 vdd.n1600 vdd.n1599 0.152939
R20247 vdd.n1601 vdd.n1600 0.152939
R20248 vdd.n1602 vdd.n1601 0.152939
R20249 vdd.n1606 vdd.n1602 0.152939
R20250 vdd.n1607 vdd.n1606 0.152939
R20251 vdd.n1608 vdd.n1607 0.152939
R20252 vdd.n1609 vdd.n1608 0.152939
R20253 vdd.n1610 vdd.n1609 0.152939
R20254 vdd.n1610 vdd.n854 0.152939
R20255 vdd.n1939 vdd.n1514 0.152939
R20256 vdd.n1477 vdd.n1476 0.152939
R20257 vdd.n1478 vdd.n1477 0.152939
R20258 vdd.n1478 vdd.n879 0.152939
R20259 vdd.n1493 vdd.n879 0.152939
R20260 vdd.n1494 vdd.n1493 0.152939
R20261 vdd.n1495 vdd.n1494 0.152939
R20262 vdd.n1495 vdd.n867 0.152939
R20263 vdd.n1512 vdd.n867 0.152939
R20264 vdd.n1513 vdd.n1512 0.152939
R20265 vdd.n1940 vdd.n1513 0.152939
R20266 vdd.n524 vdd.n519 0.152939
R20267 vdd.n525 vdd.n524 0.152939
R20268 vdd.n526 vdd.n525 0.152939
R20269 vdd.n527 vdd.n526 0.152939
R20270 vdd.n528 vdd.n527 0.152939
R20271 vdd.n529 vdd.n528 0.152939
R20272 vdd.n530 vdd.n529 0.152939
R20273 vdd.n531 vdd.n530 0.152939
R20274 vdd.n532 vdd.n531 0.152939
R20275 vdd.n533 vdd.n532 0.152939
R20276 vdd.n534 vdd.n533 0.152939
R20277 vdd.n535 vdd.n534 0.152939
R20278 vdd.n2803 vdd.n535 0.152939
R20279 vdd.n2803 vdd.n2802 0.152939
R20280 vdd.n2802 vdd.n2801 0.152939
R20281 vdd.n2801 vdd.n537 0.152939
R20282 vdd.n538 vdd.n537 0.152939
R20283 vdd.n539 vdd.n538 0.152939
R20284 vdd.n540 vdd.n539 0.152939
R20285 vdd.n541 vdd.n540 0.152939
R20286 vdd.n542 vdd.n541 0.152939
R20287 vdd.n543 vdd.n542 0.152939
R20288 vdd.n544 vdd.n543 0.152939
R20289 vdd.n545 vdd.n544 0.152939
R20290 vdd.n546 vdd.n545 0.152939
R20291 vdd.n547 vdd.n546 0.152939
R20292 vdd.n548 vdd.n547 0.152939
R20293 vdd.n549 vdd.n548 0.152939
R20294 vdd.n550 vdd.n549 0.152939
R20295 vdd.n551 vdd.n550 0.152939
R20296 vdd.n552 vdd.n551 0.152939
R20297 vdd.n553 vdd.n552 0.152939
R20298 vdd.n554 vdd.n553 0.152939
R20299 vdd.n555 vdd.n554 0.152939
R20300 vdd.n2757 vdd.n555 0.152939
R20301 vdd.n2757 vdd.n2756 0.152939
R20302 vdd.n2756 vdd.n2755 0.152939
R20303 vdd.n2755 vdd.n559 0.152939
R20304 vdd.n560 vdd.n559 0.152939
R20305 vdd.n561 vdd.n560 0.152939
R20306 vdd.n562 vdd.n561 0.152939
R20307 vdd.n563 vdd.n562 0.152939
R20308 vdd.n564 vdd.n563 0.152939
R20309 vdd.n565 vdd.n564 0.152939
R20310 vdd.n566 vdd.n565 0.152939
R20311 vdd.n567 vdd.n566 0.152939
R20312 vdd.n568 vdd.n567 0.152939
R20313 vdd.n569 vdd.n568 0.152939
R20314 vdd.n570 vdd.n569 0.152939
R20315 vdd.n571 vdd.n570 0.152939
R20316 vdd.n572 vdd.n571 0.152939
R20317 vdd.n2844 vdd.n481 0.152939
R20318 vdd.n2846 vdd.n2845 0.152939
R20319 vdd.n2846 vdd.n470 0.152939
R20320 vdd.n2861 vdd.n470 0.152939
R20321 vdd.n2862 vdd.n2861 0.152939
R20322 vdd.n2863 vdd.n2862 0.152939
R20323 vdd.n2863 vdd.n459 0.152939
R20324 vdd.n2877 vdd.n459 0.152939
R20325 vdd.n2878 vdd.n2877 0.152939
R20326 vdd.n2879 vdd.n2878 0.152939
R20327 vdd.n2879 vdd.n298 0.152939
R20328 vdd.n3046 vdd.n299 0.152939
R20329 vdd.n310 vdd.n299 0.152939
R20330 vdd.n311 vdd.n310 0.152939
R20331 vdd.n312 vdd.n311 0.152939
R20332 vdd.n320 vdd.n312 0.152939
R20333 vdd.n321 vdd.n320 0.152939
R20334 vdd.n322 vdd.n321 0.152939
R20335 vdd.n323 vdd.n322 0.152939
R20336 vdd.n331 vdd.n323 0.152939
R20337 vdd.n3022 vdd.n331 0.152939
R20338 vdd.n3021 vdd.n332 0.152939
R20339 vdd.n335 vdd.n332 0.152939
R20340 vdd.n339 vdd.n335 0.152939
R20341 vdd.n340 vdd.n339 0.152939
R20342 vdd.n341 vdd.n340 0.152939
R20343 vdd.n342 vdd.n341 0.152939
R20344 vdd.n343 vdd.n342 0.152939
R20345 vdd.n347 vdd.n343 0.152939
R20346 vdd.n348 vdd.n347 0.152939
R20347 vdd.n349 vdd.n348 0.152939
R20348 vdd.n350 vdd.n349 0.152939
R20349 vdd.n354 vdd.n350 0.152939
R20350 vdd.n355 vdd.n354 0.152939
R20351 vdd.n356 vdd.n355 0.152939
R20352 vdd.n357 vdd.n356 0.152939
R20353 vdd.n361 vdd.n357 0.152939
R20354 vdd.n362 vdd.n361 0.152939
R20355 vdd.n363 vdd.n362 0.152939
R20356 vdd.n2987 vdd.n363 0.152939
R20357 vdd.n2987 vdd.n2986 0.152939
R20358 vdd.n2986 vdd.n2985 0.152939
R20359 vdd.n2985 vdd.n369 0.152939
R20360 vdd.n374 vdd.n369 0.152939
R20361 vdd.n375 vdd.n374 0.152939
R20362 vdd.n376 vdd.n375 0.152939
R20363 vdd.n380 vdd.n376 0.152939
R20364 vdd.n381 vdd.n380 0.152939
R20365 vdd.n382 vdd.n381 0.152939
R20366 vdd.n383 vdd.n382 0.152939
R20367 vdd.n387 vdd.n383 0.152939
R20368 vdd.n388 vdd.n387 0.152939
R20369 vdd.n389 vdd.n388 0.152939
R20370 vdd.n390 vdd.n389 0.152939
R20371 vdd.n394 vdd.n390 0.152939
R20372 vdd.n395 vdd.n394 0.152939
R20373 vdd.n396 vdd.n395 0.152939
R20374 vdd.n397 vdd.n396 0.152939
R20375 vdd.n401 vdd.n397 0.152939
R20376 vdd.n402 vdd.n401 0.152939
R20377 vdd.n403 vdd.n402 0.152939
R20378 vdd.n2948 vdd.n403 0.152939
R20379 vdd.n2948 vdd.n2947 0.152939
R20380 vdd.n2947 vdd.n2946 0.152939
R20381 vdd.n2946 vdd.n409 0.152939
R20382 vdd.n414 vdd.n409 0.152939
R20383 vdd.n415 vdd.n414 0.152939
R20384 vdd.n416 vdd.n415 0.152939
R20385 vdd.n420 vdd.n416 0.152939
R20386 vdd.n421 vdd.n420 0.152939
R20387 vdd.n422 vdd.n421 0.152939
R20388 vdd.n423 vdd.n422 0.152939
R20389 vdd.n427 vdd.n423 0.152939
R20390 vdd.n428 vdd.n427 0.152939
R20391 vdd.n429 vdd.n428 0.152939
R20392 vdd.n430 vdd.n429 0.152939
R20393 vdd.n434 vdd.n430 0.152939
R20394 vdd.n435 vdd.n434 0.152939
R20395 vdd.n436 vdd.n435 0.152939
R20396 vdd.n437 vdd.n436 0.152939
R20397 vdd.n441 vdd.n437 0.152939
R20398 vdd.n442 vdd.n441 0.152939
R20399 vdd.n443 vdd.n442 0.152939
R20400 vdd.n2904 vdd.n443 0.152939
R20401 vdd.n2852 vdd.n476 0.152939
R20402 vdd.n2853 vdd.n2852 0.152939
R20403 vdd.n2854 vdd.n2853 0.152939
R20404 vdd.n2854 vdd.n464 0.152939
R20405 vdd.n2869 vdd.n464 0.152939
R20406 vdd.n2870 vdd.n2869 0.152939
R20407 vdd.n2871 vdd.n2870 0.152939
R20408 vdd.n2871 vdd.n452 0.152939
R20409 vdd.n2885 vdd.n452 0.152939
R20410 vdd.n2886 vdd.n2885 0.152939
R20411 vdd.n2887 vdd.n2886 0.152939
R20412 vdd.n2887 vdd.n450 0.152939
R20413 vdd.n2891 vdd.n450 0.152939
R20414 vdd.n2892 vdd.n2891 0.152939
R20415 vdd.n2893 vdd.n2892 0.152939
R20416 vdd.n2893 vdd.n447 0.152939
R20417 vdd.n2897 vdd.n447 0.152939
R20418 vdd.n2898 vdd.n2897 0.152939
R20419 vdd.n2899 vdd.n2898 0.152939
R20420 vdd.n2899 vdd.n444 0.152939
R20421 vdd.n2903 vdd.n444 0.152939
R20422 vdd.n2709 vdd.n2708 0.152939
R20423 vdd.n1951 vdd.n857 0.152939
R20424 vdd.n1433 vdd.n1189 0.152939
R20425 vdd.n1434 vdd.n1433 0.152939
R20426 vdd.n1435 vdd.n1434 0.152939
R20427 vdd.n1435 vdd.n1177 0.152939
R20428 vdd.n1450 vdd.n1177 0.152939
R20429 vdd.n1451 vdd.n1450 0.152939
R20430 vdd.n1452 vdd.n1451 0.152939
R20431 vdd.n1452 vdd.n1167 0.152939
R20432 vdd.n1468 vdd.n1167 0.152939
R20433 vdd.n1469 vdd.n1468 0.152939
R20434 vdd.n1470 vdd.n1469 0.152939
R20435 vdd.n1470 vdd.n884 0.152939
R20436 vdd.n1484 vdd.n884 0.152939
R20437 vdd.n1485 vdd.n1484 0.152939
R20438 vdd.n1486 vdd.n1485 0.152939
R20439 vdd.n1486 vdd.n874 0.152939
R20440 vdd.n1501 vdd.n874 0.152939
R20441 vdd.n1502 vdd.n1501 0.152939
R20442 vdd.n1505 vdd.n1502 0.152939
R20443 vdd.n1505 vdd.n1504 0.152939
R20444 vdd.n1504 vdd.n1503 0.152939
R20445 vdd.n1425 vdd.n1194 0.152939
R20446 vdd.n1418 vdd.n1194 0.152939
R20447 vdd.n1418 vdd.n1417 0.152939
R20448 vdd.n1417 vdd.n1416 0.152939
R20449 vdd.n1416 vdd.n1231 0.152939
R20450 vdd.n1412 vdd.n1231 0.152939
R20451 vdd.n1412 vdd.n1411 0.152939
R20452 vdd.n1411 vdd.n1410 0.152939
R20453 vdd.n1410 vdd.n1237 0.152939
R20454 vdd.n1406 vdd.n1237 0.152939
R20455 vdd.n1406 vdd.n1405 0.152939
R20456 vdd.n1405 vdd.n1404 0.152939
R20457 vdd.n1404 vdd.n1243 0.152939
R20458 vdd.n1400 vdd.n1243 0.152939
R20459 vdd.n1400 vdd.n1399 0.152939
R20460 vdd.n1399 vdd.n1398 0.152939
R20461 vdd.n1398 vdd.n1249 0.152939
R20462 vdd.n1394 vdd.n1249 0.152939
R20463 vdd.n1394 vdd.n1393 0.152939
R20464 vdd.n1393 vdd.n1392 0.152939
R20465 vdd.n1392 vdd.n1257 0.152939
R20466 vdd.n1388 vdd.n1257 0.152939
R20467 vdd.n1388 vdd.n1387 0.152939
R20468 vdd.n1387 vdd.n1386 0.152939
R20469 vdd.n1386 vdd.n1263 0.152939
R20470 vdd.n1382 vdd.n1263 0.152939
R20471 vdd.n1382 vdd.n1381 0.152939
R20472 vdd.n1381 vdd.n1380 0.152939
R20473 vdd.n1380 vdd.n1269 0.152939
R20474 vdd.n1376 vdd.n1269 0.152939
R20475 vdd.n1376 vdd.n1375 0.152939
R20476 vdd.n1375 vdd.n1374 0.152939
R20477 vdd.n1374 vdd.n1275 0.152939
R20478 vdd.n1370 vdd.n1275 0.152939
R20479 vdd.n1370 vdd.n1369 0.152939
R20480 vdd.n1369 vdd.n1368 0.152939
R20481 vdd.n1368 vdd.n1281 0.152939
R20482 vdd.n1364 vdd.n1281 0.152939
R20483 vdd.n1364 vdd.n1363 0.152939
R20484 vdd.n1363 vdd.n1362 0.152939
R20485 vdd.n1362 vdd.n1287 0.152939
R20486 vdd.n1355 vdd.n1287 0.152939
R20487 vdd.n1355 vdd.n1354 0.152939
R20488 vdd.n1354 vdd.n1353 0.152939
R20489 vdd.n1353 vdd.n1292 0.152939
R20490 vdd.n1349 vdd.n1292 0.152939
R20491 vdd.n1349 vdd.n1348 0.152939
R20492 vdd.n1348 vdd.n1347 0.152939
R20493 vdd.n1347 vdd.n1298 0.152939
R20494 vdd.n1343 vdd.n1298 0.152939
R20495 vdd.n1343 vdd.n1342 0.152939
R20496 vdd.n1342 vdd.n1341 0.152939
R20497 vdd.n1341 vdd.n1304 0.152939
R20498 vdd.n1337 vdd.n1304 0.152939
R20499 vdd.n1337 vdd.n1336 0.152939
R20500 vdd.n1336 vdd.n1335 0.152939
R20501 vdd.n1335 vdd.n1310 0.152939
R20502 vdd.n1331 vdd.n1310 0.152939
R20503 vdd.n1331 vdd.n1330 0.152939
R20504 vdd.n1330 vdd.n1329 0.152939
R20505 vdd.n1329 vdd.n1316 0.152939
R20506 vdd.n1325 vdd.n1316 0.152939
R20507 vdd.n1325 vdd.n1324 0.152939
R20508 vdd.n1427 vdd.n1426 0.152939
R20509 vdd.n1427 vdd.n1183 0.152939
R20510 vdd.n1442 vdd.n1183 0.152939
R20511 vdd.n1443 vdd.n1442 0.152939
R20512 vdd.n1444 vdd.n1443 0.152939
R20513 vdd.n1444 vdd.n1172 0.152939
R20514 vdd.n1459 vdd.n1172 0.152939
R20515 vdd.n1460 vdd.n1459 0.152939
R20516 vdd.n1462 vdd.n1460 0.152939
R20517 vdd.n1462 vdd.n1461 0.152939
R20518 vdd.n1929 vdd.n1514 0.110256
R20519 vdd.n2836 vdd.n481 0.110256
R20520 vdd.n2708 vdd.n2707 0.110256
R20521 vdd.n1952 vdd.n1951 0.110256
R20522 vdd.n1476 vdd.n1161 0.0695946
R20523 vdd.n3047 vdd.n298 0.0695946
R20524 vdd.n3047 vdd.n3046 0.0695946
R20525 vdd.n1461 vdd.n1161 0.0695946
R20526 vdd.n1929 vdd.n1715 0.0431829
R20527 vdd.n1952 vdd.n854 0.0431829
R20528 vdd.n2836 vdd.n519 0.0431829
R20529 vdd.n2707 vdd.n572 0.0431829
R20530 vdd vdd.n28 0.00833333
R20531 a_n1996_n452.n86 a_n1996_n452.t60 512.366
R20532 a_n1996_n452.n76 a_n1996_n452.t51 512.366
R20533 a_n1996_n452.n87 a_n1996_n452.t45 512.366
R20534 a_n1996_n452.n84 a_n1996_n452.t68 512.366
R20535 a_n1996_n452.n77 a_n1996_n452.t57 512.366
R20536 a_n1996_n452.n85 a_n1996_n452.t56 512.366
R20537 a_n1996_n452.n82 a_n1996_n452.t64 512.366
R20538 a_n1996_n452.n78 a_n1996_n452.t49 512.366
R20539 a_n1996_n452.n83 a_n1996_n452.t50 512.366
R20540 a_n1996_n452.n80 a_n1996_n452.t53 512.366
R20541 a_n1996_n452.n79 a_n1996_n452.t62 512.366
R20542 a_n1996_n452.n81 a_n1996_n452.t44 512.366
R20543 a_n1996_n452.n24 a_n1996_n452.t71 539.01
R20544 a_n1996_n452.n91 a_n1996_n452.t54 512.366
R20545 a_n1996_n452.n90 a_n1996_n452.t58 512.366
R20546 a_n1996_n452.n64 a_n1996_n452.t48 512.366
R20547 a_n1996_n452.n89 a_n1996_n452.t63 512.366
R20548 a_n1996_n452.n52 a_n1996_n452.t19 533.058
R20549 a_n1996_n452.n26 a_n1996_n452.t5 539.01
R20550 a_n1996_n452.n94 a_n1996_n452.t3 512.366
R20551 a_n1996_n452.n93 a_n1996_n452.t7 512.366
R20552 a_n1996_n452.n53 a_n1996_n452.t11 512.366
R20553 a_n1996_n452.n92 a_n1996_n452.t17 512.366
R20554 a_n1996_n452.n16 a_n1996_n452.t21 539.01
R20555 a_n1996_n452.n72 a_n1996_n452.t9 512.366
R20556 a_n1996_n452.n73 a_n1996_n452.t25 512.366
R20557 a_n1996_n452.n67 a_n1996_n452.t15 512.366
R20558 a_n1996_n452.n74 a_n1996_n452.t13 512.366
R20559 a_n1996_n452.n20 a_n1996_n452.t66 539.01
R20560 a_n1996_n452.n69 a_n1996_n452.t67 512.366
R20561 a_n1996_n452.n70 a_n1996_n452.t46 512.366
R20562 a_n1996_n452.n68 a_n1996_n452.t52 512.366
R20563 a_n1996_n452.n71 a_n1996_n452.t61 512.366
R20564 a_n1996_n452.n4 a_n1996_n452.n51 70.1674
R20565 a_n1996_n452.n6 a_n1996_n452.n49 70.1674
R20566 a_n1996_n452.n8 a_n1996_n452.n47 70.1674
R20567 a_n1996_n452.n11 a_n1996_n452.n45 70.1674
R20568 a_n1996_n452.n37 a_n1996_n452.n22 70.3058
R20569 a_n1996_n452.n31 a_n1996_n452.n34 70.1674
R20570 a_n1996_n452.n34 a_n1996_n452.n53 20.9683
R20571 a_n1996_n452.n33 a_n1996_n452.n32 75.0448
R20572 a_n1996_n452.n93 a_n1996_n452.n33 11.2134
R20573 a_n1996_n452.n25 a_n1996_n452.n26 44.8194
R20574 a_n1996_n452.n52 a_n1996_n452.n31 70.3058
R20575 a_n1996_n452.n23 a_n1996_n452.n36 70.1674
R20576 a_n1996_n452.n36 a_n1996_n452.n64 20.9683
R20577 a_n1996_n452.n35 a_n1996_n452.n23 75.0448
R20578 a_n1996_n452.n90 a_n1996_n452.n35 11.2134
R20579 a_n1996_n452.n21 a_n1996_n452.n24 44.8194
R20580 a_n1996_n452.n13 a_n1996_n452.n43 70.3058
R20581 a_n1996_n452.n17 a_n1996_n452.n40 70.3058
R20582 a_n1996_n452.n39 a_n1996_n452.n18 70.1674
R20583 a_n1996_n452.n39 a_n1996_n452.n68 20.9683
R20584 a_n1996_n452.n18 a_n1996_n452.n38 75.0448
R20585 a_n1996_n452.n70 a_n1996_n452.n38 11.2134
R20586 a_n1996_n452.n19 a_n1996_n452.n20 44.8194
R20587 a_n1996_n452.n42 a_n1996_n452.n14 70.1674
R20588 a_n1996_n452.n42 a_n1996_n452.n67 20.9683
R20589 a_n1996_n452.n14 a_n1996_n452.n41 75.0448
R20590 a_n1996_n452.n73 a_n1996_n452.n41 11.2134
R20591 a_n1996_n452.n15 a_n1996_n452.n16 44.8194
R20592 a_n1996_n452.n81 a_n1996_n452.n45 20.9683
R20593 a_n1996_n452.n44 a_n1996_n452.n12 75.0448
R20594 a_n1996_n452.n44 a_n1996_n452.n79 11.2134
R20595 a_n1996_n452.n12 a_n1996_n452.n80 161.3
R20596 a_n1996_n452.n83 a_n1996_n452.n47 20.9683
R20597 a_n1996_n452.n46 a_n1996_n452.n9 75.0448
R20598 a_n1996_n452.n46 a_n1996_n452.n78 11.2134
R20599 a_n1996_n452.n9 a_n1996_n452.n82 161.3
R20600 a_n1996_n452.n85 a_n1996_n452.n49 20.9683
R20601 a_n1996_n452.n48 a_n1996_n452.n7 75.0448
R20602 a_n1996_n452.n48 a_n1996_n452.n77 11.2134
R20603 a_n1996_n452.n7 a_n1996_n452.n84 161.3
R20604 a_n1996_n452.n87 a_n1996_n452.n51 20.9683
R20605 a_n1996_n452.n50 a_n1996_n452.n5 75.0448
R20606 a_n1996_n452.n50 a_n1996_n452.n76 11.2134
R20607 a_n1996_n452.n5 a_n1996_n452.n86 161.3
R20608 a_n1996_n452.n3 a_n1996_n452.n62 81.3764
R20609 a_n1996_n452.n1 a_n1996_n452.n57 81.3764
R20610 a_n1996_n452.n0 a_n1996_n452.n54 81.3764
R20611 a_n1996_n452.n3 a_n1996_n452.n63 80.9324
R20612 a_n1996_n452.n3 a_n1996_n452.n61 80.9324
R20613 a_n1996_n452.n2 a_n1996_n452.n60 80.9324
R20614 a_n1996_n452.n2 a_n1996_n452.n59 80.9324
R20615 a_n1996_n452.n1 a_n1996_n452.n58 80.9324
R20616 a_n1996_n452.n1 a_n1996_n452.n56 80.9324
R20617 a_n1996_n452.n0 a_n1996_n452.n55 80.9324
R20618 a_n1996_n452.n30 a_n1996_n452.t20 74.6477
R20619 a_n1996_n452.n27 a_n1996_n452.t22 74.6477
R20620 a_n1996_n452.n29 a_n1996_n452.t6 74.2899
R20621 a_n1996_n452.n28 a_n1996_n452.t24 74.2897
R20622 a_n1996_n452.n30 a_n1996_n452.n96 70.6783
R20623 a_n1996_n452.n28 a_n1996_n452.n66 70.6783
R20624 a_n1996_n452.n27 a_n1996_n452.n65 70.6783
R20625 a_n1996_n452.n97 a_n1996_n452.n30 70.6782
R20626 a_n1996_n452.n86 a_n1996_n452.n76 48.2005
R20627 a_n1996_n452.t65 a_n1996_n452.n51 533.335
R20628 a_n1996_n452.n84 a_n1996_n452.n77 48.2005
R20629 a_n1996_n452.t70 a_n1996_n452.n49 533.335
R20630 a_n1996_n452.n82 a_n1996_n452.n78 48.2005
R20631 a_n1996_n452.t59 a_n1996_n452.n47 533.335
R20632 a_n1996_n452.n80 a_n1996_n452.n79 48.2005
R20633 a_n1996_n452.t55 a_n1996_n452.n45 533.335
R20634 a_n1996_n452.n91 a_n1996_n452.n90 48.2005
R20635 a_n1996_n452.n89 a_n1996_n452.n36 20.9683
R20636 a_n1996_n452.n94 a_n1996_n452.n93 48.2005
R20637 a_n1996_n452.n92 a_n1996_n452.n34 20.9683
R20638 a_n1996_n452.n73 a_n1996_n452.n72 48.2005
R20639 a_n1996_n452.n74 a_n1996_n452.n42 20.9683
R20640 a_n1996_n452.n70 a_n1996_n452.n69 48.2005
R20641 a_n1996_n452.n71 a_n1996_n452.n39 20.9683
R20642 a_n1996_n452.n37 a_n1996_n452.t69 533.058
R20643 a_n1996_n452.t23 a_n1996_n452.n43 533.058
R20644 a_n1996_n452.t47 a_n1996_n452.n40 533.058
R20645 a_n1996_n452.n2 a_n1996_n452.n1 32.0139
R20646 a_n1996_n452.n87 a_n1996_n452.n50 35.3134
R20647 a_n1996_n452.n85 a_n1996_n452.n48 35.3134
R20648 a_n1996_n452.n83 a_n1996_n452.n46 35.3134
R20649 a_n1996_n452.n81 a_n1996_n452.n44 35.3134
R20650 a_n1996_n452.n35 a_n1996_n452.n64 35.3134
R20651 a_n1996_n452.n33 a_n1996_n452.n53 35.3134
R20652 a_n1996_n452.n67 a_n1996_n452.n41 35.3134
R20653 a_n1996_n452.n68 a_n1996_n452.n38 35.3134
R20654 a_n1996_n452.n31 a_n1996_n452.n3 23.891
R20655 a_n1996_n452.n19 a_n1996_n452.n10 12.046
R20656 a_n1996_n452.n22 a_n1996_n452.n88 11.8414
R20657 a_n1996_n452.n95 a_n1996_n452.n25 10.5365
R20658 a_n1996_n452.n75 a_n1996_n452.n28 9.50122
R20659 a_n1996_n452.n88 a_n1996_n452.n4 7.47588
R20660 a_n1996_n452.n12 a_n1996_n452.n10 7.47588
R20661 a_n1996_n452.n75 a_n1996_n452.n13 6.70126
R20662 a_n1996_n452.n29 a_n1996_n452.n95 5.65783
R20663 a_n1996_n452.n88 a_n1996_n452.n75 5.3452
R20664 a_n1996_n452.n31 a_n1996_n452.n21 3.95126
R20665 a_n1996_n452.n15 a_n1996_n452.n17 3.95126
R20666 a_n1996_n452.n96 a_n1996_n452.t12 3.61217
R20667 a_n1996_n452.n96 a_n1996_n452.t18 3.61217
R20668 a_n1996_n452.n66 a_n1996_n452.t16 3.61217
R20669 a_n1996_n452.n66 a_n1996_n452.t14 3.61217
R20670 a_n1996_n452.n65 a_n1996_n452.t10 3.61217
R20671 a_n1996_n452.n65 a_n1996_n452.t26 3.61217
R20672 a_n1996_n452.t4 a_n1996_n452.n97 3.61217
R20673 a_n1996_n452.n97 a_n1996_n452.t8 3.61217
R20674 a_n1996_n452.n62 a_n1996_n452.t41 2.82907
R20675 a_n1996_n452.n62 a_n1996_n452.t43 2.82907
R20676 a_n1996_n452.n63 a_n1996_n452.t28 2.82907
R20677 a_n1996_n452.n63 a_n1996_n452.t29 2.82907
R20678 a_n1996_n452.n61 a_n1996_n452.t2 2.82907
R20679 a_n1996_n452.n61 a_n1996_n452.t30 2.82907
R20680 a_n1996_n452.n60 a_n1996_n452.t32 2.82907
R20681 a_n1996_n452.n60 a_n1996_n452.t33 2.82907
R20682 a_n1996_n452.n59 a_n1996_n452.t39 2.82907
R20683 a_n1996_n452.n59 a_n1996_n452.t35 2.82907
R20684 a_n1996_n452.n57 a_n1996_n452.t40 2.82907
R20685 a_n1996_n452.n57 a_n1996_n452.t37 2.82907
R20686 a_n1996_n452.n58 a_n1996_n452.t1 2.82907
R20687 a_n1996_n452.n58 a_n1996_n452.t0 2.82907
R20688 a_n1996_n452.n56 a_n1996_n452.t36 2.82907
R20689 a_n1996_n452.n56 a_n1996_n452.t27 2.82907
R20690 a_n1996_n452.n55 a_n1996_n452.t38 2.82907
R20691 a_n1996_n452.n55 a_n1996_n452.t34 2.82907
R20692 a_n1996_n452.n54 a_n1996_n452.t31 2.82907
R20693 a_n1996_n452.n54 a_n1996_n452.t42 2.82907
R20694 a_n1996_n452.n95 a_n1996_n452.n10 1.30542
R20695 a_n1996_n452.n7 a_n1996_n452.n8 1.04595
R20696 a_n1996_n452.n24 a_n1996_n452.n91 13.657
R20697 a_n1996_n452.n89 a_n1996_n452.n37 21.4216
R20698 a_n1996_n452.n26 a_n1996_n452.n94 13.657
R20699 a_n1996_n452.n92 a_n1996_n452.n52 21.4216
R20700 a_n1996_n452.n72 a_n1996_n452.n16 13.657
R20701 a_n1996_n452.n43 a_n1996_n452.n74 21.4216
R20702 a_n1996_n452.n69 a_n1996_n452.n20 13.657
R20703 a_n1996_n452.n40 a_n1996_n452.n71 21.4216
R20704 a_n1996_n452.n3 a_n1996_n452.n2 1.3324
R20705 a_n1996_n452.n1 a_n1996_n452.n0 0.888431
R20706 a_n1996_n452.n32 a_n1996_n452.n25 0.758076
R20707 a_n1996_n452.n23 a_n1996_n452.n21 0.758076
R20708 a_n1996_n452.n23 a_n1996_n452.n22 0.758076
R20709 a_n1996_n452.n19 a_n1996_n452.n18 0.758076
R20710 a_n1996_n452.n18 a_n1996_n452.n17 0.758076
R20711 a_n1996_n452.n15 a_n1996_n452.n14 0.758076
R20712 a_n1996_n452.n14 a_n1996_n452.n13 0.758076
R20713 a_n1996_n452.n12 a_n1996_n452.n11 0.758076
R20714 a_n1996_n452.n9 a_n1996_n452.n8 0.758076
R20715 a_n1996_n452.n7 a_n1996_n452.n6 0.758076
R20716 a_n1996_n452.n5 a_n1996_n452.n4 0.758076
R20717 a_n1996_n452.n32 a_n1996_n452.n31 0.720197
R20718 a_n1996_n452.n30 a_n1996_n452.n29 0.716017
R20719 a_n1996_n452.n28 a_n1996_n452.n27 0.716017
R20720 a_n1996_n452.n9 a_n1996_n452.n11 0.67853
R20721 a_n1996_n452.n5 a_n1996_n452.n6 0.67853
R20722 a_n1986_8322.n6 a_n1986_8322.t14 74.6477
R20723 a_n1986_8322.n1 a_n1986_8322.t1 74.6477
R20724 a_n1986_8322.n16 a_n1986_8322.t10 74.6474
R20725 a_n1986_8322.n14 a_n1986_8322.t3 74.2899
R20726 a_n1986_8322.n7 a_n1986_8322.t12 74.2899
R20727 a_n1986_8322.n8 a_n1986_8322.t15 74.2899
R20728 a_n1986_8322.n11 a_n1986_8322.t16 74.2899
R20729 a_n1986_8322.n4 a_n1986_8322.t0 74.2899
R20730 a_n1986_8322.n16 a_n1986_8322.n15 70.6783
R20731 a_n1986_8322.n6 a_n1986_8322.n5 70.6783
R20732 a_n1986_8322.n10 a_n1986_8322.n9 70.6783
R20733 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R20734 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R20735 a_n1986_8322.n18 a_n1986_8322.n17 70.6782
R20736 a_n1986_8322.n12 a_n1986_8322.n4 22.7556
R20737 a_n1986_8322.n13 a_n1986_8322.t20 9.94227
R20738 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R20739 a_n1986_8322.n14 a_n1986_8322.n13 5.83671
R20740 a_n1986_8322.n13 a_n1986_8322.n12 5.3452
R20741 a_n1986_8322.n15 a_n1986_8322.t8 3.61217
R20742 a_n1986_8322.n15 a_n1986_8322.t5 3.61217
R20743 a_n1986_8322.n5 a_n1986_8322.t18 3.61217
R20744 a_n1986_8322.n5 a_n1986_8322.t17 3.61217
R20745 a_n1986_8322.n9 a_n1986_8322.t13 3.61217
R20746 a_n1986_8322.n9 a_n1986_8322.t19 3.61217
R20747 a_n1986_8322.n0 a_n1986_8322.t9 3.61217
R20748 a_n1986_8322.n0 a_n1986_8322.t4 3.61217
R20749 a_n1986_8322.n2 a_n1986_8322.t7 3.61217
R20750 a_n1986_8322.n2 a_n1986_8322.t6 3.61217
R20751 a_n1986_8322.n18 a_n1986_8322.t2 3.61217
R20752 a_n1986_8322.t11 a_n1986_8322.n18 3.61217
R20753 a_n1986_8322.n11 a_n1986_8322.n10 0.358259
R20754 a_n1986_8322.n10 a_n1986_8322.n8 0.358259
R20755 a_n1986_8322.n7 a_n1986_8322.n6 0.358259
R20756 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R20757 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R20758 a_n1986_8322.n17 a_n1986_8322.n14 0.358259
R20759 a_n1986_8322.n17 a_n1986_8322.n16 0.358259
R20760 a_n1986_8322.n8 a_n1986_8322.n7 0.101793
R20761 a_n1986_8322.t23 a_n1986_8322.t22 0.0788333
R20762 a_n1986_8322.t21 a_n1986_8322.t23 0.0631667
R20763 a_n1986_8322.t20 a_n1986_8322.t21 0.0471944
R20764 a_n1986_8322.t20 a_n1986_8322.t22 0.0453889
R20765 a_n1808_13878.n5 a_n1808_13878.n3 98.9633
R20766 a_n1808_13878.n2 a_n1808_13878.n0 98.7517
R20767 a_n1808_13878.n2 a_n1808_13878.n1 98.6055
R20768 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R20769 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R20770 a_n1808_13878.n7 a_n1808_13878.n6 98.6054
R20771 a_n1808_13878.n9 a_n1808_13878.t13 74.6477
R20772 a_n1808_13878.n14 a_n1808_13878.t14 74.2899
R20773 a_n1808_13878.n11 a_n1808_13878.t15 74.2899
R20774 a_n1808_13878.n10 a_n1808_13878.t12 74.2899
R20775 a_n1808_13878.n13 a_n1808_13878.n12 70.6783
R20776 a_n1808_13878.n9 a_n1808_13878.n8 70.6783
R20777 a_n1808_13878.n16 a_n1808_13878.n15 13.5694
R20778 a_n1808_13878.n15 a_n1808_13878.n7 11.5762
R20779 a_n1808_13878.n15 a_n1808_13878.n14 6.2408
R20780 a_n1808_13878.n1 a_n1808_13878.t6 3.61217
R20781 a_n1808_13878.n1 a_n1808_13878.t1 3.61217
R20782 a_n1808_13878.n0 a_n1808_13878.t0 3.61217
R20783 a_n1808_13878.n0 a_n1808_13878.t2 3.61217
R20784 a_n1808_13878.n6 a_n1808_13878.t7 3.61217
R20785 a_n1808_13878.n6 a_n1808_13878.t8 3.61217
R20786 a_n1808_13878.n4 a_n1808_13878.t10 3.61217
R20787 a_n1808_13878.n4 a_n1808_13878.t3 3.61217
R20788 a_n1808_13878.n3 a_n1808_13878.t5 3.61217
R20789 a_n1808_13878.n3 a_n1808_13878.t9 3.61217
R20790 a_n1808_13878.n12 a_n1808_13878.t18 3.61217
R20791 a_n1808_13878.n12 a_n1808_13878.t19 3.61217
R20792 a_n1808_13878.n8 a_n1808_13878.t16 3.61217
R20793 a_n1808_13878.n8 a_n1808_13878.t17 3.61217
R20794 a_n1808_13878.n17 a_n1808_13878.t4 3.61217
R20795 a_n1808_13878.t11 a_n1808_13878.n17 3.61217
R20796 a_n1808_13878.n7 a_n1808_13878.n5 0.358259
R20797 a_n1808_13878.n10 a_n1808_13878.n9 0.358259
R20798 a_n1808_13878.n13 a_n1808_13878.n11 0.358259
R20799 a_n1808_13878.n14 a_n1808_13878.n13 0.358259
R20800 a_n1808_13878.n16 a_n1808_13878.n2 0.146627
R20801 a_n1808_13878.n11 a_n1808_13878.n10 0.101793
R20802 diffpairibias.n0 diffpairibias.t27 436.822
R20803 diffpairibias.n27 diffpairibias.t24 435.479
R20804 diffpairibias.n26 diffpairibias.t21 435.479
R20805 diffpairibias.n25 diffpairibias.t22 435.479
R20806 diffpairibias.n24 diffpairibias.t26 435.479
R20807 diffpairibias.n23 diffpairibias.t20 435.479
R20808 diffpairibias.n0 diffpairibias.t23 435.479
R20809 diffpairibias.n1 diffpairibias.t28 435.479
R20810 diffpairibias.n2 diffpairibias.t25 435.479
R20811 diffpairibias.n3 diffpairibias.t29 435.479
R20812 diffpairibias.n13 diffpairibias.t14 377.536
R20813 diffpairibias.n13 diffpairibias.t0 376.193
R20814 diffpairibias.n14 diffpairibias.t10 376.193
R20815 diffpairibias.n15 diffpairibias.t12 376.193
R20816 diffpairibias.n16 diffpairibias.t6 376.193
R20817 diffpairibias.n17 diffpairibias.t2 376.193
R20818 diffpairibias.n18 diffpairibias.t16 376.193
R20819 diffpairibias.n19 diffpairibias.t4 376.193
R20820 diffpairibias.n20 diffpairibias.t18 376.193
R20821 diffpairibias.n21 diffpairibias.t8 376.193
R20822 diffpairibias.n4 diffpairibias.t15 113.368
R20823 diffpairibias.n4 diffpairibias.t1 112.698
R20824 diffpairibias.n5 diffpairibias.t11 112.698
R20825 diffpairibias.n6 diffpairibias.t13 112.698
R20826 diffpairibias.n7 diffpairibias.t7 112.698
R20827 diffpairibias.n8 diffpairibias.t3 112.698
R20828 diffpairibias.n9 diffpairibias.t17 112.698
R20829 diffpairibias.n10 diffpairibias.t5 112.698
R20830 diffpairibias.n11 diffpairibias.t19 112.698
R20831 diffpairibias.n12 diffpairibias.t9 112.698
R20832 diffpairibias.n22 diffpairibias.n21 4.77242
R20833 diffpairibias.n22 diffpairibias.n12 4.30807
R20834 diffpairibias.n23 diffpairibias.n22 4.13945
R20835 diffpairibias.n21 diffpairibias.n20 1.34352
R20836 diffpairibias.n20 diffpairibias.n19 1.34352
R20837 diffpairibias.n19 diffpairibias.n18 1.34352
R20838 diffpairibias.n18 diffpairibias.n17 1.34352
R20839 diffpairibias.n17 diffpairibias.n16 1.34352
R20840 diffpairibias.n16 diffpairibias.n15 1.34352
R20841 diffpairibias.n15 diffpairibias.n14 1.34352
R20842 diffpairibias.n14 diffpairibias.n13 1.34352
R20843 diffpairibias.n3 diffpairibias.n2 1.34352
R20844 diffpairibias.n2 diffpairibias.n1 1.34352
R20845 diffpairibias.n1 diffpairibias.n0 1.34352
R20846 diffpairibias.n24 diffpairibias.n23 1.34352
R20847 diffpairibias.n25 diffpairibias.n24 1.34352
R20848 diffpairibias.n26 diffpairibias.n25 1.34352
R20849 diffpairibias.n27 diffpairibias.n26 1.34352
R20850 diffpairibias.n28 diffpairibias.n27 0.862419
R20851 diffpairibias diffpairibias.n28 0.684875
R20852 diffpairibias.n12 diffpairibias.n11 0.672012
R20853 diffpairibias.n11 diffpairibias.n10 0.672012
R20854 diffpairibias.n10 diffpairibias.n9 0.672012
R20855 diffpairibias.n9 diffpairibias.n8 0.672012
R20856 diffpairibias.n8 diffpairibias.n7 0.672012
R20857 diffpairibias.n7 diffpairibias.n6 0.672012
R20858 diffpairibias.n6 diffpairibias.n5 0.672012
R20859 diffpairibias.n5 diffpairibias.n4 0.672012
R20860 diffpairibias.n28 diffpairibias.n3 0.190907
R20861 minus.n43 minus.t24 322.512
R20862 minus.n9 minus.t8 322.512
R20863 minus.n66 minus.t5 297.12
R20864 minus.n64 minus.t6 297.12
R20865 minus.n36 minus.t22 297.12
R20866 minus.n58 minus.t18 297.12
R20867 minus.n38 minus.t19 297.12
R20868 minus.n52 minus.t14 297.12
R20869 minus.n40 minus.t15 297.12
R20870 minus.n46 minus.t9 297.12
R20871 minus.n42 minus.t23 297.12
R20872 minus.n8 minus.t7 297.12
R20873 minus.n12 minus.t11 297.12
R20874 minus.n14 minus.t10 297.12
R20875 minus.n18 minus.t12 297.12
R20876 minus.n20 minus.t17 297.12
R20877 minus.n24 minus.t16 297.12
R20878 minus.n26 minus.t21 297.12
R20879 minus.n30 minus.t20 297.12
R20880 minus.n32 minus.t13 297.12
R20881 minus.n72 minus.t4 243.255
R20882 minus.n71 minus.n69 224.169
R20883 minus.n71 minus.n70 223.454
R20884 minus.n45 minus.n44 161.3
R20885 minus.n46 minus.n41 161.3
R20886 minus.n48 minus.n47 161.3
R20887 minus.n49 minus.n40 161.3
R20888 minus.n51 minus.n50 161.3
R20889 minus.n52 minus.n39 161.3
R20890 minus.n54 minus.n53 161.3
R20891 minus.n55 minus.n38 161.3
R20892 minus.n57 minus.n56 161.3
R20893 minus.n58 minus.n37 161.3
R20894 minus.n60 minus.n59 161.3
R20895 minus.n61 minus.n36 161.3
R20896 minus.n63 minus.n62 161.3
R20897 minus.n64 minus.n35 161.3
R20898 minus.n65 minus.n34 161.3
R20899 minus.n67 minus.n66 161.3
R20900 minus.n33 minus.n32 161.3
R20901 minus.n31 minus.n0 161.3
R20902 minus.n30 minus.n29 161.3
R20903 minus.n28 minus.n1 161.3
R20904 minus.n27 minus.n26 161.3
R20905 minus.n25 minus.n2 161.3
R20906 minus.n24 minus.n23 161.3
R20907 minus.n22 minus.n3 161.3
R20908 minus.n21 minus.n20 161.3
R20909 minus.n19 minus.n4 161.3
R20910 minus.n18 minus.n17 161.3
R20911 minus.n16 minus.n5 161.3
R20912 minus.n15 minus.n14 161.3
R20913 minus.n13 minus.n6 161.3
R20914 minus.n12 minus.n11 161.3
R20915 minus.n10 minus.n7 161.3
R20916 minus.n44 minus.n43 45.0031
R20917 minus.n10 minus.n9 45.0031
R20918 minus.n66 minus.n65 41.6278
R20919 minus.n32 minus.n31 41.6278
R20920 minus.n64 minus.n63 37.246
R20921 minus.n45 minus.n42 37.246
R20922 minus.n8 minus.n7 37.246
R20923 minus.n30 minus.n1 37.246
R20924 minus.n59 minus.n36 32.8641
R20925 minus.n47 minus.n46 32.8641
R20926 minus.n13 minus.n12 32.8641
R20927 minus.n26 minus.n25 32.8641
R20928 minus.n68 minus.n67 31.8206
R20929 minus.n58 minus.n57 28.4823
R20930 minus.n51 minus.n40 28.4823
R20931 minus.n14 minus.n5 28.4823
R20932 minus.n24 minus.n3 28.4823
R20933 minus.n53 minus.n38 24.1005
R20934 minus.n53 minus.n52 24.1005
R20935 minus.n19 minus.n18 24.1005
R20936 minus.n20 minus.n19 24.1005
R20937 minus.n70 minus.t3 19.8005
R20938 minus.n70 minus.t1 19.8005
R20939 minus.n69 minus.t2 19.8005
R20940 minus.n69 minus.t0 19.8005
R20941 minus.n57 minus.n38 19.7187
R20942 minus.n52 minus.n51 19.7187
R20943 minus.n18 minus.n5 19.7187
R20944 minus.n20 minus.n3 19.7187
R20945 minus.n43 minus.n42 15.6319
R20946 minus.n9 minus.n8 15.6319
R20947 minus.n59 minus.n58 15.3369
R20948 minus.n47 minus.n40 15.3369
R20949 minus.n14 minus.n13 15.3369
R20950 minus.n25 minus.n24 15.3369
R20951 minus.n68 minus.n33 12.0819
R20952 minus minus.n73 11.4968
R20953 minus.n63 minus.n36 10.955
R20954 minus.n46 minus.n45 10.955
R20955 minus.n12 minus.n7 10.955
R20956 minus.n26 minus.n1 10.955
R20957 minus.n65 minus.n64 6.57323
R20958 minus.n31 minus.n30 6.57323
R20959 minus.n73 minus.n72 4.80222
R20960 minus.n73 minus.n68 0.972091
R20961 minus.n72 minus.n71 0.716017
R20962 minus.n67 minus.n34 0.189894
R20963 minus.n35 minus.n34 0.189894
R20964 minus.n62 minus.n35 0.189894
R20965 minus.n62 minus.n61 0.189894
R20966 minus.n61 minus.n60 0.189894
R20967 minus.n60 minus.n37 0.189894
R20968 minus.n56 minus.n37 0.189894
R20969 minus.n56 minus.n55 0.189894
R20970 minus.n55 minus.n54 0.189894
R20971 minus.n54 minus.n39 0.189894
R20972 minus.n50 minus.n39 0.189894
R20973 minus.n50 minus.n49 0.189894
R20974 minus.n49 minus.n48 0.189894
R20975 minus.n48 minus.n41 0.189894
R20976 minus.n44 minus.n41 0.189894
R20977 minus.n11 minus.n10 0.189894
R20978 minus.n11 minus.n6 0.189894
R20979 minus.n15 minus.n6 0.189894
R20980 minus.n16 minus.n15 0.189894
R20981 minus.n17 minus.n16 0.189894
R20982 minus.n17 minus.n4 0.189894
R20983 minus.n21 minus.n4 0.189894
R20984 minus.n22 minus.n21 0.189894
R20985 minus.n23 minus.n22 0.189894
R20986 minus.n23 minus.n2 0.189894
R20987 minus.n27 minus.n2 0.189894
R20988 minus.n28 minus.n27 0.189894
R20989 minus.n29 minus.n28 0.189894
R20990 minus.n29 minus.n0 0.189894
R20991 minus.n33 minus.n0 0.189894
R20992 outputibias.n27 outputibias.n1 289.615
R20993 outputibias.n58 outputibias.n32 289.615
R20994 outputibias.n90 outputibias.n64 289.615
R20995 outputibias.n122 outputibias.n96 289.615
R20996 outputibias.n28 outputibias.n27 185
R20997 outputibias.n26 outputibias.n25 185
R20998 outputibias.n5 outputibias.n4 185
R20999 outputibias.n20 outputibias.n19 185
R21000 outputibias.n18 outputibias.n17 185
R21001 outputibias.n9 outputibias.n8 185
R21002 outputibias.n12 outputibias.n11 185
R21003 outputibias.n59 outputibias.n58 185
R21004 outputibias.n57 outputibias.n56 185
R21005 outputibias.n36 outputibias.n35 185
R21006 outputibias.n51 outputibias.n50 185
R21007 outputibias.n49 outputibias.n48 185
R21008 outputibias.n40 outputibias.n39 185
R21009 outputibias.n43 outputibias.n42 185
R21010 outputibias.n91 outputibias.n90 185
R21011 outputibias.n89 outputibias.n88 185
R21012 outputibias.n68 outputibias.n67 185
R21013 outputibias.n83 outputibias.n82 185
R21014 outputibias.n81 outputibias.n80 185
R21015 outputibias.n72 outputibias.n71 185
R21016 outputibias.n75 outputibias.n74 185
R21017 outputibias.n123 outputibias.n122 185
R21018 outputibias.n121 outputibias.n120 185
R21019 outputibias.n100 outputibias.n99 185
R21020 outputibias.n115 outputibias.n114 185
R21021 outputibias.n113 outputibias.n112 185
R21022 outputibias.n104 outputibias.n103 185
R21023 outputibias.n107 outputibias.n106 185
R21024 outputibias.n0 outputibias.t10 178.945
R21025 outputibias.n133 outputibias.t8 177.018
R21026 outputibias.n132 outputibias.t11 177.018
R21027 outputibias.n0 outputibias.t9 177.018
R21028 outputibias.t7 outputibias.n10 147.661
R21029 outputibias.t1 outputibias.n41 147.661
R21030 outputibias.t3 outputibias.n73 147.661
R21031 outputibias.t5 outputibias.n105 147.661
R21032 outputibias.n128 outputibias.t6 132.363
R21033 outputibias.n128 outputibias.t0 130.436
R21034 outputibias.n129 outputibias.t2 130.436
R21035 outputibias.n130 outputibias.t4 130.436
R21036 outputibias.n27 outputibias.n26 104.615
R21037 outputibias.n26 outputibias.n4 104.615
R21038 outputibias.n19 outputibias.n4 104.615
R21039 outputibias.n19 outputibias.n18 104.615
R21040 outputibias.n18 outputibias.n8 104.615
R21041 outputibias.n11 outputibias.n8 104.615
R21042 outputibias.n58 outputibias.n57 104.615
R21043 outputibias.n57 outputibias.n35 104.615
R21044 outputibias.n50 outputibias.n35 104.615
R21045 outputibias.n50 outputibias.n49 104.615
R21046 outputibias.n49 outputibias.n39 104.615
R21047 outputibias.n42 outputibias.n39 104.615
R21048 outputibias.n90 outputibias.n89 104.615
R21049 outputibias.n89 outputibias.n67 104.615
R21050 outputibias.n82 outputibias.n67 104.615
R21051 outputibias.n82 outputibias.n81 104.615
R21052 outputibias.n81 outputibias.n71 104.615
R21053 outputibias.n74 outputibias.n71 104.615
R21054 outputibias.n122 outputibias.n121 104.615
R21055 outputibias.n121 outputibias.n99 104.615
R21056 outputibias.n114 outputibias.n99 104.615
R21057 outputibias.n114 outputibias.n113 104.615
R21058 outputibias.n113 outputibias.n103 104.615
R21059 outputibias.n106 outputibias.n103 104.615
R21060 outputibias.n63 outputibias.n31 95.6354
R21061 outputibias.n63 outputibias.n62 94.6732
R21062 outputibias.n95 outputibias.n94 94.6732
R21063 outputibias.n127 outputibias.n126 94.6732
R21064 outputibias.n11 outputibias.t7 52.3082
R21065 outputibias.n42 outputibias.t1 52.3082
R21066 outputibias.n74 outputibias.t3 52.3082
R21067 outputibias.n106 outputibias.t5 52.3082
R21068 outputibias.n12 outputibias.n10 15.6674
R21069 outputibias.n43 outputibias.n41 15.6674
R21070 outputibias.n75 outputibias.n73 15.6674
R21071 outputibias.n107 outputibias.n105 15.6674
R21072 outputibias.n13 outputibias.n9 12.8005
R21073 outputibias.n44 outputibias.n40 12.8005
R21074 outputibias.n76 outputibias.n72 12.8005
R21075 outputibias.n108 outputibias.n104 12.8005
R21076 outputibias.n17 outputibias.n16 12.0247
R21077 outputibias.n48 outputibias.n47 12.0247
R21078 outputibias.n80 outputibias.n79 12.0247
R21079 outputibias.n112 outputibias.n111 12.0247
R21080 outputibias.n20 outputibias.n7 11.249
R21081 outputibias.n51 outputibias.n38 11.249
R21082 outputibias.n83 outputibias.n70 11.249
R21083 outputibias.n115 outputibias.n102 11.249
R21084 outputibias.n21 outputibias.n5 10.4732
R21085 outputibias.n52 outputibias.n36 10.4732
R21086 outputibias.n84 outputibias.n68 10.4732
R21087 outputibias.n116 outputibias.n100 10.4732
R21088 outputibias.n25 outputibias.n24 9.69747
R21089 outputibias.n56 outputibias.n55 9.69747
R21090 outputibias.n88 outputibias.n87 9.69747
R21091 outputibias.n120 outputibias.n119 9.69747
R21092 outputibias.n31 outputibias.n30 9.45567
R21093 outputibias.n62 outputibias.n61 9.45567
R21094 outputibias.n94 outputibias.n93 9.45567
R21095 outputibias.n126 outputibias.n125 9.45567
R21096 outputibias.n30 outputibias.n29 9.3005
R21097 outputibias.n3 outputibias.n2 9.3005
R21098 outputibias.n24 outputibias.n23 9.3005
R21099 outputibias.n22 outputibias.n21 9.3005
R21100 outputibias.n7 outputibias.n6 9.3005
R21101 outputibias.n16 outputibias.n15 9.3005
R21102 outputibias.n14 outputibias.n13 9.3005
R21103 outputibias.n61 outputibias.n60 9.3005
R21104 outputibias.n34 outputibias.n33 9.3005
R21105 outputibias.n55 outputibias.n54 9.3005
R21106 outputibias.n53 outputibias.n52 9.3005
R21107 outputibias.n38 outputibias.n37 9.3005
R21108 outputibias.n47 outputibias.n46 9.3005
R21109 outputibias.n45 outputibias.n44 9.3005
R21110 outputibias.n93 outputibias.n92 9.3005
R21111 outputibias.n66 outputibias.n65 9.3005
R21112 outputibias.n87 outputibias.n86 9.3005
R21113 outputibias.n85 outputibias.n84 9.3005
R21114 outputibias.n70 outputibias.n69 9.3005
R21115 outputibias.n79 outputibias.n78 9.3005
R21116 outputibias.n77 outputibias.n76 9.3005
R21117 outputibias.n125 outputibias.n124 9.3005
R21118 outputibias.n98 outputibias.n97 9.3005
R21119 outputibias.n119 outputibias.n118 9.3005
R21120 outputibias.n117 outputibias.n116 9.3005
R21121 outputibias.n102 outputibias.n101 9.3005
R21122 outputibias.n111 outputibias.n110 9.3005
R21123 outputibias.n109 outputibias.n108 9.3005
R21124 outputibias.n28 outputibias.n3 8.92171
R21125 outputibias.n59 outputibias.n34 8.92171
R21126 outputibias.n91 outputibias.n66 8.92171
R21127 outputibias.n123 outputibias.n98 8.92171
R21128 outputibias.n29 outputibias.n1 8.14595
R21129 outputibias.n60 outputibias.n32 8.14595
R21130 outputibias.n92 outputibias.n64 8.14595
R21131 outputibias.n124 outputibias.n96 8.14595
R21132 outputibias.n31 outputibias.n1 5.81868
R21133 outputibias.n62 outputibias.n32 5.81868
R21134 outputibias.n94 outputibias.n64 5.81868
R21135 outputibias.n126 outputibias.n96 5.81868
R21136 outputibias.n131 outputibias.n130 5.20947
R21137 outputibias.n29 outputibias.n28 5.04292
R21138 outputibias.n60 outputibias.n59 5.04292
R21139 outputibias.n92 outputibias.n91 5.04292
R21140 outputibias.n124 outputibias.n123 5.04292
R21141 outputibias.n131 outputibias.n127 4.42209
R21142 outputibias.n14 outputibias.n10 4.38594
R21143 outputibias.n45 outputibias.n41 4.38594
R21144 outputibias.n77 outputibias.n73 4.38594
R21145 outputibias.n109 outputibias.n105 4.38594
R21146 outputibias.n132 outputibias.n131 4.28454
R21147 outputibias.n25 outputibias.n3 4.26717
R21148 outputibias.n56 outputibias.n34 4.26717
R21149 outputibias.n88 outputibias.n66 4.26717
R21150 outputibias.n120 outputibias.n98 4.26717
R21151 outputibias.n24 outputibias.n5 3.49141
R21152 outputibias.n55 outputibias.n36 3.49141
R21153 outputibias.n87 outputibias.n68 3.49141
R21154 outputibias.n119 outputibias.n100 3.49141
R21155 outputibias.n21 outputibias.n20 2.71565
R21156 outputibias.n52 outputibias.n51 2.71565
R21157 outputibias.n84 outputibias.n83 2.71565
R21158 outputibias.n116 outputibias.n115 2.71565
R21159 outputibias.n17 outputibias.n7 1.93989
R21160 outputibias.n48 outputibias.n38 1.93989
R21161 outputibias.n80 outputibias.n70 1.93989
R21162 outputibias.n112 outputibias.n102 1.93989
R21163 outputibias.n130 outputibias.n129 1.9266
R21164 outputibias.n129 outputibias.n128 1.9266
R21165 outputibias.n133 outputibias.n132 1.92658
R21166 outputibias.n134 outputibias.n133 1.29913
R21167 outputibias.n16 outputibias.n9 1.16414
R21168 outputibias.n47 outputibias.n40 1.16414
R21169 outputibias.n79 outputibias.n72 1.16414
R21170 outputibias.n111 outputibias.n104 1.16414
R21171 outputibias.n127 outputibias.n95 0.962709
R21172 outputibias.n95 outputibias.n63 0.962709
R21173 outputibias.n13 outputibias.n12 0.388379
R21174 outputibias.n44 outputibias.n43 0.388379
R21175 outputibias.n76 outputibias.n75 0.388379
R21176 outputibias.n108 outputibias.n107 0.388379
R21177 outputibias.n134 outputibias.n0 0.337251
R21178 outputibias outputibias.n134 0.302375
R21179 outputibias.n30 outputibias.n2 0.155672
R21180 outputibias.n23 outputibias.n2 0.155672
R21181 outputibias.n23 outputibias.n22 0.155672
R21182 outputibias.n22 outputibias.n6 0.155672
R21183 outputibias.n15 outputibias.n6 0.155672
R21184 outputibias.n15 outputibias.n14 0.155672
R21185 outputibias.n61 outputibias.n33 0.155672
R21186 outputibias.n54 outputibias.n33 0.155672
R21187 outputibias.n54 outputibias.n53 0.155672
R21188 outputibias.n53 outputibias.n37 0.155672
R21189 outputibias.n46 outputibias.n37 0.155672
R21190 outputibias.n46 outputibias.n45 0.155672
R21191 outputibias.n93 outputibias.n65 0.155672
R21192 outputibias.n86 outputibias.n65 0.155672
R21193 outputibias.n86 outputibias.n85 0.155672
R21194 outputibias.n85 outputibias.n69 0.155672
R21195 outputibias.n78 outputibias.n69 0.155672
R21196 outputibias.n78 outputibias.n77 0.155672
R21197 outputibias.n125 outputibias.n97 0.155672
R21198 outputibias.n118 outputibias.n97 0.155672
R21199 outputibias.n118 outputibias.n117 0.155672
R21200 outputibias.n117 outputibias.n101 0.155672
R21201 outputibias.n110 outputibias.n101 0.155672
R21202 outputibias.n110 outputibias.n109 0.155672
R21203 output.n41 output.n15 289.615
R21204 output.n72 output.n46 289.615
R21205 output.n104 output.n78 289.615
R21206 output.n136 output.n110 289.615
R21207 output.n77 output.n45 197.26
R21208 output.n77 output.n76 196.298
R21209 output.n109 output.n108 196.298
R21210 output.n141 output.n140 196.298
R21211 output.n42 output.n41 185
R21212 output.n40 output.n39 185
R21213 output.n19 output.n18 185
R21214 output.n34 output.n33 185
R21215 output.n32 output.n31 185
R21216 output.n23 output.n22 185
R21217 output.n26 output.n25 185
R21218 output.n73 output.n72 185
R21219 output.n71 output.n70 185
R21220 output.n50 output.n49 185
R21221 output.n65 output.n64 185
R21222 output.n63 output.n62 185
R21223 output.n54 output.n53 185
R21224 output.n57 output.n56 185
R21225 output.n105 output.n104 185
R21226 output.n103 output.n102 185
R21227 output.n82 output.n81 185
R21228 output.n97 output.n96 185
R21229 output.n95 output.n94 185
R21230 output.n86 output.n85 185
R21231 output.n89 output.n88 185
R21232 output.n137 output.n136 185
R21233 output.n135 output.n134 185
R21234 output.n114 output.n113 185
R21235 output.n129 output.n128 185
R21236 output.n127 output.n126 185
R21237 output.n118 output.n117 185
R21238 output.n121 output.n120 185
R21239 output.t17 output.n24 147.661
R21240 output.t18 output.n55 147.661
R21241 output.t19 output.n87 147.661
R21242 output.t16 output.n119 147.661
R21243 output.n41 output.n40 104.615
R21244 output.n40 output.n18 104.615
R21245 output.n33 output.n18 104.615
R21246 output.n33 output.n32 104.615
R21247 output.n32 output.n22 104.615
R21248 output.n25 output.n22 104.615
R21249 output.n72 output.n71 104.615
R21250 output.n71 output.n49 104.615
R21251 output.n64 output.n49 104.615
R21252 output.n64 output.n63 104.615
R21253 output.n63 output.n53 104.615
R21254 output.n56 output.n53 104.615
R21255 output.n104 output.n103 104.615
R21256 output.n103 output.n81 104.615
R21257 output.n96 output.n81 104.615
R21258 output.n96 output.n95 104.615
R21259 output.n95 output.n85 104.615
R21260 output.n88 output.n85 104.615
R21261 output.n136 output.n135 104.615
R21262 output.n135 output.n113 104.615
R21263 output.n128 output.n113 104.615
R21264 output.n128 output.n127 104.615
R21265 output.n127 output.n117 104.615
R21266 output.n120 output.n117 104.615
R21267 output.n1 output.t1 77.056
R21268 output.n14 output.t2 76.6694
R21269 output.n1 output.n0 72.7095
R21270 output.n3 output.n2 72.7095
R21271 output.n5 output.n4 72.7095
R21272 output.n7 output.n6 72.7095
R21273 output.n9 output.n8 72.7095
R21274 output.n11 output.n10 72.7095
R21275 output.n13 output.n12 72.7095
R21276 output.n25 output.t17 52.3082
R21277 output.n56 output.t18 52.3082
R21278 output.n88 output.t19 52.3082
R21279 output.n120 output.t16 52.3082
R21280 output.n26 output.n24 15.6674
R21281 output.n57 output.n55 15.6674
R21282 output.n89 output.n87 15.6674
R21283 output.n121 output.n119 15.6674
R21284 output.n27 output.n23 12.8005
R21285 output.n58 output.n54 12.8005
R21286 output.n90 output.n86 12.8005
R21287 output.n122 output.n118 12.8005
R21288 output.n31 output.n30 12.0247
R21289 output.n62 output.n61 12.0247
R21290 output.n94 output.n93 12.0247
R21291 output.n126 output.n125 12.0247
R21292 output.n34 output.n21 11.249
R21293 output.n65 output.n52 11.249
R21294 output.n97 output.n84 11.249
R21295 output.n129 output.n116 11.249
R21296 output.n35 output.n19 10.4732
R21297 output.n66 output.n50 10.4732
R21298 output.n98 output.n82 10.4732
R21299 output.n130 output.n114 10.4732
R21300 output.n39 output.n38 9.69747
R21301 output.n70 output.n69 9.69747
R21302 output.n102 output.n101 9.69747
R21303 output.n134 output.n133 9.69747
R21304 output.n45 output.n44 9.45567
R21305 output.n76 output.n75 9.45567
R21306 output.n108 output.n107 9.45567
R21307 output.n140 output.n139 9.45567
R21308 output.n44 output.n43 9.3005
R21309 output.n17 output.n16 9.3005
R21310 output.n38 output.n37 9.3005
R21311 output.n36 output.n35 9.3005
R21312 output.n21 output.n20 9.3005
R21313 output.n30 output.n29 9.3005
R21314 output.n28 output.n27 9.3005
R21315 output.n75 output.n74 9.3005
R21316 output.n48 output.n47 9.3005
R21317 output.n69 output.n68 9.3005
R21318 output.n67 output.n66 9.3005
R21319 output.n52 output.n51 9.3005
R21320 output.n61 output.n60 9.3005
R21321 output.n59 output.n58 9.3005
R21322 output.n107 output.n106 9.3005
R21323 output.n80 output.n79 9.3005
R21324 output.n101 output.n100 9.3005
R21325 output.n99 output.n98 9.3005
R21326 output.n84 output.n83 9.3005
R21327 output.n93 output.n92 9.3005
R21328 output.n91 output.n90 9.3005
R21329 output.n139 output.n138 9.3005
R21330 output.n112 output.n111 9.3005
R21331 output.n133 output.n132 9.3005
R21332 output.n131 output.n130 9.3005
R21333 output.n116 output.n115 9.3005
R21334 output.n125 output.n124 9.3005
R21335 output.n123 output.n122 9.3005
R21336 output.n42 output.n17 8.92171
R21337 output.n73 output.n48 8.92171
R21338 output.n105 output.n80 8.92171
R21339 output.n137 output.n112 8.92171
R21340 output output.n141 8.15037
R21341 output.n43 output.n15 8.14595
R21342 output.n74 output.n46 8.14595
R21343 output.n106 output.n78 8.14595
R21344 output.n138 output.n110 8.14595
R21345 output.n45 output.n15 5.81868
R21346 output.n76 output.n46 5.81868
R21347 output.n108 output.n78 5.81868
R21348 output.n140 output.n110 5.81868
R21349 output.n43 output.n42 5.04292
R21350 output.n74 output.n73 5.04292
R21351 output.n106 output.n105 5.04292
R21352 output.n138 output.n137 5.04292
R21353 output.n28 output.n24 4.38594
R21354 output.n59 output.n55 4.38594
R21355 output.n91 output.n87 4.38594
R21356 output.n123 output.n119 4.38594
R21357 output.n39 output.n17 4.26717
R21358 output.n70 output.n48 4.26717
R21359 output.n102 output.n80 4.26717
R21360 output.n134 output.n112 4.26717
R21361 output.n0 output.t12 3.9605
R21362 output.n0 output.t15 3.9605
R21363 output.n2 output.t5 3.9605
R21364 output.n2 output.t4 3.9605
R21365 output.n4 output.t10 3.9605
R21366 output.n4 output.t14 3.9605
R21367 output.n6 output.t3 3.9605
R21368 output.n6 output.t6 3.9605
R21369 output.n8 output.t7 3.9605
R21370 output.n8 output.t13 3.9605
R21371 output.n10 output.t0 3.9605
R21372 output.n10 output.t8 3.9605
R21373 output.n12 output.t11 3.9605
R21374 output.n12 output.t9 3.9605
R21375 output.n38 output.n19 3.49141
R21376 output.n69 output.n50 3.49141
R21377 output.n101 output.n82 3.49141
R21378 output.n133 output.n114 3.49141
R21379 output.n35 output.n34 2.71565
R21380 output.n66 output.n65 2.71565
R21381 output.n98 output.n97 2.71565
R21382 output.n130 output.n129 2.71565
R21383 output.n31 output.n21 1.93989
R21384 output.n62 output.n52 1.93989
R21385 output.n94 output.n84 1.93989
R21386 output.n126 output.n116 1.93989
R21387 output.n30 output.n23 1.16414
R21388 output.n61 output.n54 1.16414
R21389 output.n93 output.n86 1.16414
R21390 output.n125 output.n118 1.16414
R21391 output.n141 output.n109 0.962709
R21392 output.n109 output.n77 0.962709
R21393 output.n27 output.n26 0.388379
R21394 output.n58 output.n57 0.388379
R21395 output.n90 output.n89 0.388379
R21396 output.n122 output.n121 0.388379
R21397 output.n14 output.n13 0.387128
R21398 output.n13 output.n11 0.387128
R21399 output.n11 output.n9 0.387128
R21400 output.n9 output.n7 0.387128
R21401 output.n7 output.n5 0.387128
R21402 output.n5 output.n3 0.387128
R21403 output.n3 output.n1 0.387128
R21404 output.n44 output.n16 0.155672
R21405 output.n37 output.n16 0.155672
R21406 output.n37 output.n36 0.155672
R21407 output.n36 output.n20 0.155672
R21408 output.n29 output.n20 0.155672
R21409 output.n29 output.n28 0.155672
R21410 output.n75 output.n47 0.155672
R21411 output.n68 output.n47 0.155672
R21412 output.n68 output.n67 0.155672
R21413 output.n67 output.n51 0.155672
R21414 output.n60 output.n51 0.155672
R21415 output.n60 output.n59 0.155672
R21416 output.n107 output.n79 0.155672
R21417 output.n100 output.n79 0.155672
R21418 output.n100 output.n99 0.155672
R21419 output.n99 output.n83 0.155672
R21420 output.n92 output.n83 0.155672
R21421 output.n92 output.n91 0.155672
R21422 output.n139 output.n111 0.155672
R21423 output.n132 output.n111 0.155672
R21424 output.n132 output.n131 0.155672
R21425 output.n131 output.n115 0.155672
R21426 output.n124 output.n115 0.155672
R21427 output.n124 output.n123 0.155672
R21428 output output.n14 0.126227
C0 commonsourceibias diffpairibias 0.064336f
C1 minus plus 9.175731f
C2 CSoutput commonsourceibias 42.3358f
C3 minus commonsourceibias 0.332601f
C4 plus commonsourceibias 0.278362f
C5 output outputibias 2.34152f
C6 vdd output 7.23429f
C7 CSoutput output 6.13881f
C8 CSoutput outputibias 0.032386f
C9 vdd CSoutput 67.6707f
C10 minus diffpairibias 3.4e-19
C11 commonsourceibias output 0.006808f
C12 vdd plus 0.066355f
C13 CSoutput minus 2.72666f
C14 plus diffpairibias 3.42e-19
C15 commonsourceibias outputibias 0.003832f
C16 CSoutput plus 0.856333f
C17 vdd commonsourceibias 0.004218f
C18 diffpairibias gnd 60.00273f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.145027p
C22 plus gnd 33.4462f
C23 minus gnd 27.49025f
C24 CSoutput gnd 0.108285p
C25 vdd gnd 0.345061p
C26 output.t1 gnd 0.464308f
C27 output.t12 gnd 0.044422f
C28 output.t15 gnd 0.044422f
C29 output.n0 gnd 0.364624f
C30 output.n1 gnd 0.614102f
C31 output.t5 gnd 0.044422f
C32 output.t4 gnd 0.044422f
C33 output.n2 gnd 0.364624f
C34 output.n3 gnd 0.350265f
C35 output.t10 gnd 0.044422f
C36 output.t14 gnd 0.044422f
C37 output.n4 gnd 0.364624f
C38 output.n5 gnd 0.350265f
C39 output.t3 gnd 0.044422f
C40 output.t6 gnd 0.044422f
C41 output.n6 gnd 0.364624f
C42 output.n7 gnd 0.350265f
C43 output.t7 gnd 0.044422f
C44 output.t13 gnd 0.044422f
C45 output.n8 gnd 0.364624f
C46 output.n9 gnd 0.350265f
C47 output.t0 gnd 0.044422f
C48 output.t8 gnd 0.044422f
C49 output.n10 gnd 0.364624f
C50 output.n11 gnd 0.350265f
C51 output.t11 gnd 0.044422f
C52 output.t9 gnd 0.044422f
C53 output.n12 gnd 0.364624f
C54 output.n13 gnd 0.350265f
C55 output.t2 gnd 0.462979f
C56 output.n14 gnd 0.28994f
C57 output.n15 gnd 0.015803f
C58 output.n16 gnd 0.011243f
C59 output.n17 gnd 0.006041f
C60 output.n18 gnd 0.01428f
C61 output.n19 gnd 0.006397f
C62 output.n20 gnd 0.011243f
C63 output.n21 gnd 0.006041f
C64 output.n22 gnd 0.01428f
C65 output.n23 gnd 0.006397f
C66 output.n24 gnd 0.048111f
C67 output.t17 gnd 0.023274f
C68 output.n25 gnd 0.01071f
C69 output.n26 gnd 0.008435f
C70 output.n27 gnd 0.006041f
C71 output.n28 gnd 0.267512f
C72 output.n29 gnd 0.011243f
C73 output.n30 gnd 0.006041f
C74 output.n31 gnd 0.006397f
C75 output.n32 gnd 0.01428f
C76 output.n33 gnd 0.01428f
C77 output.n34 gnd 0.006397f
C78 output.n35 gnd 0.006041f
C79 output.n36 gnd 0.011243f
C80 output.n37 gnd 0.011243f
C81 output.n38 gnd 0.006041f
C82 output.n39 gnd 0.006397f
C83 output.n40 gnd 0.01428f
C84 output.n41 gnd 0.030913f
C85 output.n42 gnd 0.006397f
C86 output.n43 gnd 0.006041f
C87 output.n44 gnd 0.025987f
C88 output.n45 gnd 0.097665f
C89 output.n46 gnd 0.015803f
C90 output.n47 gnd 0.011243f
C91 output.n48 gnd 0.006041f
C92 output.n49 gnd 0.01428f
C93 output.n50 gnd 0.006397f
C94 output.n51 gnd 0.011243f
C95 output.n52 gnd 0.006041f
C96 output.n53 gnd 0.01428f
C97 output.n54 gnd 0.006397f
C98 output.n55 gnd 0.048111f
C99 output.t18 gnd 0.023274f
C100 output.n56 gnd 0.01071f
C101 output.n57 gnd 0.008435f
C102 output.n58 gnd 0.006041f
C103 output.n59 gnd 0.267512f
C104 output.n60 gnd 0.011243f
C105 output.n61 gnd 0.006041f
C106 output.n62 gnd 0.006397f
C107 output.n63 gnd 0.01428f
C108 output.n64 gnd 0.01428f
C109 output.n65 gnd 0.006397f
C110 output.n66 gnd 0.006041f
C111 output.n67 gnd 0.011243f
C112 output.n68 gnd 0.011243f
C113 output.n69 gnd 0.006041f
C114 output.n70 gnd 0.006397f
C115 output.n71 gnd 0.01428f
C116 output.n72 gnd 0.030913f
C117 output.n73 gnd 0.006397f
C118 output.n74 gnd 0.006041f
C119 output.n75 gnd 0.025987f
C120 output.n76 gnd 0.09306f
C121 output.n77 gnd 1.65264f
C122 output.n78 gnd 0.015803f
C123 output.n79 gnd 0.011243f
C124 output.n80 gnd 0.006041f
C125 output.n81 gnd 0.01428f
C126 output.n82 gnd 0.006397f
C127 output.n83 gnd 0.011243f
C128 output.n84 gnd 0.006041f
C129 output.n85 gnd 0.01428f
C130 output.n86 gnd 0.006397f
C131 output.n87 gnd 0.048111f
C132 output.t19 gnd 0.023274f
C133 output.n88 gnd 0.01071f
C134 output.n89 gnd 0.008435f
C135 output.n90 gnd 0.006041f
C136 output.n91 gnd 0.267512f
C137 output.n92 gnd 0.011243f
C138 output.n93 gnd 0.006041f
C139 output.n94 gnd 0.006397f
C140 output.n95 gnd 0.01428f
C141 output.n96 gnd 0.01428f
C142 output.n97 gnd 0.006397f
C143 output.n98 gnd 0.006041f
C144 output.n99 gnd 0.011243f
C145 output.n100 gnd 0.011243f
C146 output.n101 gnd 0.006041f
C147 output.n102 gnd 0.006397f
C148 output.n103 gnd 0.01428f
C149 output.n104 gnd 0.030913f
C150 output.n105 gnd 0.006397f
C151 output.n106 gnd 0.006041f
C152 output.n107 gnd 0.025987f
C153 output.n108 gnd 0.09306f
C154 output.n109 gnd 0.713089f
C155 output.n110 gnd 0.015803f
C156 output.n111 gnd 0.011243f
C157 output.n112 gnd 0.006041f
C158 output.n113 gnd 0.01428f
C159 output.n114 gnd 0.006397f
C160 output.n115 gnd 0.011243f
C161 output.n116 gnd 0.006041f
C162 output.n117 gnd 0.01428f
C163 output.n118 gnd 0.006397f
C164 output.n119 gnd 0.048111f
C165 output.t16 gnd 0.023274f
C166 output.n120 gnd 0.01071f
C167 output.n121 gnd 0.008435f
C168 output.n122 gnd 0.006041f
C169 output.n123 gnd 0.267512f
C170 output.n124 gnd 0.011243f
C171 output.n125 gnd 0.006041f
C172 output.n126 gnd 0.006397f
C173 output.n127 gnd 0.01428f
C174 output.n128 gnd 0.01428f
C175 output.n129 gnd 0.006397f
C176 output.n130 gnd 0.006041f
C177 output.n131 gnd 0.011243f
C178 output.n132 gnd 0.011243f
C179 output.n133 gnd 0.006041f
C180 output.n134 gnd 0.006397f
C181 output.n135 gnd 0.01428f
C182 output.n136 gnd 0.030913f
C183 output.n137 gnd 0.006397f
C184 output.n138 gnd 0.006041f
C185 output.n139 gnd 0.025987f
C186 output.n140 gnd 0.09306f
C187 output.n141 gnd 1.67353f
C188 outputibias.t9 gnd 0.11477f
C189 outputibias.t10 gnd 0.115567f
C190 outputibias.n0 gnd 0.130108f
C191 outputibias.n1 gnd 0.001372f
C192 outputibias.n2 gnd 9.76e-19
C193 outputibias.n3 gnd 5.24e-19
C194 outputibias.n4 gnd 0.001239f
C195 outputibias.n5 gnd 5.55e-19
C196 outputibias.n6 gnd 9.76e-19
C197 outputibias.n7 gnd 5.24e-19
C198 outputibias.n8 gnd 0.001239f
C199 outputibias.n9 gnd 5.55e-19
C200 outputibias.n10 gnd 0.004176f
C201 outputibias.t7 gnd 0.00202f
C202 outputibias.n11 gnd 9.3e-19
C203 outputibias.n12 gnd 7.32e-19
C204 outputibias.n13 gnd 5.24e-19
C205 outputibias.n14 gnd 0.02322f
C206 outputibias.n15 gnd 9.76e-19
C207 outputibias.n16 gnd 5.24e-19
C208 outputibias.n17 gnd 5.55e-19
C209 outputibias.n18 gnd 0.001239f
C210 outputibias.n19 gnd 0.001239f
C211 outputibias.n20 gnd 5.55e-19
C212 outputibias.n21 gnd 5.24e-19
C213 outputibias.n22 gnd 9.76e-19
C214 outputibias.n23 gnd 9.76e-19
C215 outputibias.n24 gnd 5.24e-19
C216 outputibias.n25 gnd 5.55e-19
C217 outputibias.n26 gnd 0.001239f
C218 outputibias.n27 gnd 0.002683f
C219 outputibias.n28 gnd 5.55e-19
C220 outputibias.n29 gnd 5.24e-19
C221 outputibias.n30 gnd 0.002256f
C222 outputibias.n31 gnd 0.005781f
C223 outputibias.n32 gnd 0.001372f
C224 outputibias.n33 gnd 9.76e-19
C225 outputibias.n34 gnd 5.24e-19
C226 outputibias.n35 gnd 0.001239f
C227 outputibias.n36 gnd 5.55e-19
C228 outputibias.n37 gnd 9.76e-19
C229 outputibias.n38 gnd 5.24e-19
C230 outputibias.n39 gnd 0.001239f
C231 outputibias.n40 gnd 5.55e-19
C232 outputibias.n41 gnd 0.004176f
C233 outputibias.t1 gnd 0.00202f
C234 outputibias.n42 gnd 9.3e-19
C235 outputibias.n43 gnd 7.32e-19
C236 outputibias.n44 gnd 5.24e-19
C237 outputibias.n45 gnd 0.02322f
C238 outputibias.n46 gnd 9.76e-19
C239 outputibias.n47 gnd 5.24e-19
C240 outputibias.n48 gnd 5.55e-19
C241 outputibias.n49 gnd 0.001239f
C242 outputibias.n50 gnd 0.001239f
C243 outputibias.n51 gnd 5.55e-19
C244 outputibias.n52 gnd 5.24e-19
C245 outputibias.n53 gnd 9.76e-19
C246 outputibias.n54 gnd 9.76e-19
C247 outputibias.n55 gnd 5.24e-19
C248 outputibias.n56 gnd 5.55e-19
C249 outputibias.n57 gnd 0.001239f
C250 outputibias.n58 gnd 0.002683f
C251 outputibias.n59 gnd 5.55e-19
C252 outputibias.n60 gnd 5.24e-19
C253 outputibias.n61 gnd 0.002256f
C254 outputibias.n62 gnd 0.005197f
C255 outputibias.n63 gnd 0.121892f
C256 outputibias.n64 gnd 0.001372f
C257 outputibias.n65 gnd 9.76e-19
C258 outputibias.n66 gnd 5.24e-19
C259 outputibias.n67 gnd 0.001239f
C260 outputibias.n68 gnd 5.55e-19
C261 outputibias.n69 gnd 9.76e-19
C262 outputibias.n70 gnd 5.24e-19
C263 outputibias.n71 gnd 0.001239f
C264 outputibias.n72 gnd 5.55e-19
C265 outputibias.n73 gnd 0.004176f
C266 outputibias.t3 gnd 0.00202f
C267 outputibias.n74 gnd 9.3e-19
C268 outputibias.n75 gnd 7.32e-19
C269 outputibias.n76 gnd 5.24e-19
C270 outputibias.n77 gnd 0.02322f
C271 outputibias.n78 gnd 9.76e-19
C272 outputibias.n79 gnd 5.24e-19
C273 outputibias.n80 gnd 5.55e-19
C274 outputibias.n81 gnd 0.001239f
C275 outputibias.n82 gnd 0.001239f
C276 outputibias.n83 gnd 5.55e-19
C277 outputibias.n84 gnd 5.24e-19
C278 outputibias.n85 gnd 9.76e-19
C279 outputibias.n86 gnd 9.76e-19
C280 outputibias.n87 gnd 5.24e-19
C281 outputibias.n88 gnd 5.55e-19
C282 outputibias.n89 gnd 0.001239f
C283 outputibias.n90 gnd 0.002683f
C284 outputibias.n91 gnd 5.55e-19
C285 outputibias.n92 gnd 5.24e-19
C286 outputibias.n93 gnd 0.002256f
C287 outputibias.n94 gnd 0.005197f
C288 outputibias.n95 gnd 0.064513f
C289 outputibias.n96 gnd 0.001372f
C290 outputibias.n97 gnd 9.76e-19
C291 outputibias.n98 gnd 5.24e-19
C292 outputibias.n99 gnd 0.001239f
C293 outputibias.n100 gnd 5.55e-19
C294 outputibias.n101 gnd 9.76e-19
C295 outputibias.n102 gnd 5.24e-19
C296 outputibias.n103 gnd 0.001239f
C297 outputibias.n104 gnd 5.55e-19
C298 outputibias.n105 gnd 0.004176f
C299 outputibias.t5 gnd 0.00202f
C300 outputibias.n106 gnd 9.3e-19
C301 outputibias.n107 gnd 7.32e-19
C302 outputibias.n108 gnd 5.24e-19
C303 outputibias.n109 gnd 0.02322f
C304 outputibias.n110 gnd 9.76e-19
C305 outputibias.n111 gnd 5.24e-19
C306 outputibias.n112 gnd 5.55e-19
C307 outputibias.n113 gnd 0.001239f
C308 outputibias.n114 gnd 0.001239f
C309 outputibias.n115 gnd 5.55e-19
C310 outputibias.n116 gnd 5.24e-19
C311 outputibias.n117 gnd 9.76e-19
C312 outputibias.n118 gnd 9.76e-19
C313 outputibias.n119 gnd 5.24e-19
C314 outputibias.n120 gnd 5.55e-19
C315 outputibias.n121 gnd 0.001239f
C316 outputibias.n122 gnd 0.002683f
C317 outputibias.n123 gnd 5.55e-19
C318 outputibias.n124 gnd 5.24e-19
C319 outputibias.n125 gnd 0.002256f
C320 outputibias.n126 gnd 0.005197f
C321 outputibias.n127 gnd 0.084814f
C322 outputibias.t4 gnd 0.108319f
C323 outputibias.t2 gnd 0.108319f
C324 outputibias.t0 gnd 0.108319f
C325 outputibias.t6 gnd 0.109238f
C326 outputibias.n128 gnd 0.134674f
C327 outputibias.n129 gnd 0.07244f
C328 outputibias.n130 gnd 0.079818f
C329 outputibias.n131 gnd 0.164901f
C330 outputibias.t11 gnd 0.11477f
C331 outputibias.n132 gnd 0.067481f
C332 outputibias.t8 gnd 0.11477f
C333 outputibias.n133 gnd 0.065115f
C334 outputibias.n134 gnd 0.029159f
C335 minus.n0 gnd 0.031825f
C336 minus.n1 gnd 0.007222f
C337 minus.n2 gnd 0.031825f
C338 minus.n3 gnd 0.007222f
C339 minus.n4 gnd 0.031825f
C340 minus.n5 gnd 0.007222f
C341 minus.n6 gnd 0.031825f
C342 minus.n7 gnd 0.007222f
C343 minus.t8 gnd 0.465911f
C344 minus.t7 gnd 0.45014f
C345 minus.n8 gnd 0.20529f
C346 minus.n9 gnd 0.186481f
C347 minus.n10 gnd 0.135844f
C348 minus.n11 gnd 0.031825f
C349 minus.t11 gnd 0.45014f
C350 minus.n12 gnd 0.199967f
C351 minus.n13 gnd 0.007222f
C352 minus.t10 gnd 0.45014f
C353 minus.n14 gnd 0.199967f
C354 minus.n15 gnd 0.031825f
C355 minus.n16 gnd 0.031825f
C356 minus.n17 gnd 0.031825f
C357 minus.t12 gnd 0.45014f
C358 minus.n18 gnd 0.199967f
C359 minus.n19 gnd 0.007222f
C360 minus.t17 gnd 0.45014f
C361 minus.n20 gnd 0.199967f
C362 minus.n21 gnd 0.031825f
C363 minus.n22 gnd 0.031825f
C364 minus.n23 gnd 0.031825f
C365 minus.t16 gnd 0.45014f
C366 minus.n24 gnd 0.199967f
C367 minus.n25 gnd 0.007222f
C368 minus.t21 gnd 0.45014f
C369 minus.n26 gnd 0.199967f
C370 minus.n27 gnd 0.031825f
C371 minus.n28 gnd 0.031825f
C372 minus.n29 gnd 0.031825f
C373 minus.t20 gnd 0.45014f
C374 minus.n30 gnd 0.199967f
C375 minus.n31 gnd 0.007222f
C376 minus.t13 gnd 0.45014f
C377 minus.n32 gnd 0.199672f
C378 minus.n33 gnd 0.367718f
C379 minus.n34 gnd 0.031825f
C380 minus.t5 gnd 0.45014f
C381 minus.t6 gnd 0.45014f
C382 minus.n35 gnd 0.031825f
C383 minus.t22 gnd 0.45014f
C384 minus.n36 gnd 0.199967f
C385 minus.n37 gnd 0.031825f
C386 minus.t18 gnd 0.45014f
C387 minus.t19 gnd 0.45014f
C388 minus.n38 gnd 0.199967f
C389 minus.n39 gnd 0.031825f
C390 minus.t14 gnd 0.45014f
C391 minus.t15 gnd 0.45014f
C392 minus.n40 gnd 0.199967f
C393 minus.n41 gnd 0.031825f
C394 minus.t9 gnd 0.45014f
C395 minus.t23 gnd 0.45014f
C396 minus.n42 gnd 0.20529f
C397 minus.t24 gnd 0.465911f
C398 minus.n43 gnd 0.186481f
C399 minus.n44 gnd 0.135844f
C400 minus.n45 gnd 0.007222f
C401 minus.n46 gnd 0.199967f
C402 minus.n47 gnd 0.007222f
C403 minus.n48 gnd 0.031825f
C404 minus.n49 gnd 0.031825f
C405 minus.n50 gnd 0.031825f
C406 minus.n51 gnd 0.007222f
C407 minus.n52 gnd 0.199967f
C408 minus.n53 gnd 0.007222f
C409 minus.n54 gnd 0.031825f
C410 minus.n55 gnd 0.031825f
C411 minus.n56 gnd 0.031825f
C412 minus.n57 gnd 0.007222f
C413 minus.n58 gnd 0.199967f
C414 minus.n59 gnd 0.007222f
C415 minus.n60 gnd 0.031825f
C416 minus.n61 gnd 0.031825f
C417 minus.n62 gnd 0.031825f
C418 minus.n63 gnd 0.007222f
C419 minus.n64 gnd 0.199967f
C420 minus.n65 gnd 0.007222f
C421 minus.n66 gnd 0.199672f
C422 minus.n67 gnd 0.994453f
C423 minus.n68 gnd 1.49713f
C424 minus.t2 gnd 0.009811f
C425 minus.t0 gnd 0.009811f
C426 minus.n69 gnd 0.03226f
C427 minus.t3 gnd 0.009811f
C428 minus.t1 gnd 0.009811f
C429 minus.n70 gnd 0.031818f
C430 minus.n71 gnd 0.271554f
C431 minus.t4 gnd 0.054606f
C432 minus.n72 gnd 0.148185f
C433 minus.n73 gnd 1.96997f
C434 diffpairibias.t27 gnd 0.090128f
C435 diffpairibias.t23 gnd 0.08996f
C436 diffpairibias.n0 gnd 0.105991f
C437 diffpairibias.t28 gnd 0.08996f
C438 diffpairibias.n1 gnd 0.051736f
C439 diffpairibias.t25 gnd 0.08996f
C440 diffpairibias.n2 gnd 0.051736f
C441 diffpairibias.t29 gnd 0.08996f
C442 diffpairibias.n3 gnd 0.041084f
C443 diffpairibias.t15 gnd 0.086371f
C444 diffpairibias.t1 gnd 0.085993f
C445 diffpairibias.n4 gnd 0.13579f
C446 diffpairibias.t11 gnd 0.085993f
C447 diffpairibias.n5 gnd 0.072463f
C448 diffpairibias.t13 gnd 0.085993f
C449 diffpairibias.n6 gnd 0.072463f
C450 diffpairibias.t7 gnd 0.085993f
C451 diffpairibias.n7 gnd 0.072463f
C452 diffpairibias.t3 gnd 0.085993f
C453 diffpairibias.n8 gnd 0.072463f
C454 diffpairibias.t17 gnd 0.085993f
C455 diffpairibias.n9 gnd 0.072463f
C456 diffpairibias.t5 gnd 0.085993f
C457 diffpairibias.n10 gnd 0.072463f
C458 diffpairibias.t19 gnd 0.085993f
C459 diffpairibias.n11 gnd 0.072463f
C460 diffpairibias.t9 gnd 0.085993f
C461 diffpairibias.n12 gnd 0.102883f
C462 diffpairibias.t14 gnd 0.086899f
C463 diffpairibias.t0 gnd 0.086748f
C464 diffpairibias.n13 gnd 0.094648f
C465 diffpairibias.t10 gnd 0.086748f
C466 diffpairibias.n14 gnd 0.052262f
C467 diffpairibias.t12 gnd 0.086748f
C468 diffpairibias.n15 gnd 0.052262f
C469 diffpairibias.t6 gnd 0.086748f
C470 diffpairibias.n16 gnd 0.052262f
C471 diffpairibias.t2 gnd 0.086748f
C472 diffpairibias.n17 gnd 0.052262f
C473 diffpairibias.t16 gnd 0.086748f
C474 diffpairibias.n18 gnd 0.052262f
C475 diffpairibias.t4 gnd 0.086748f
C476 diffpairibias.n19 gnd 0.052262f
C477 diffpairibias.t18 gnd 0.086748f
C478 diffpairibias.n20 gnd 0.052262f
C479 diffpairibias.t8 gnd 0.086748f
C480 diffpairibias.n21 gnd 0.061849f
C481 diffpairibias.n22 gnd 0.233513f
C482 diffpairibias.t20 gnd 0.08996f
C483 diffpairibias.n23 gnd 0.051747f
C484 diffpairibias.t26 gnd 0.08996f
C485 diffpairibias.n24 gnd 0.051736f
C486 diffpairibias.t22 gnd 0.08996f
C487 diffpairibias.n25 gnd 0.051736f
C488 diffpairibias.t21 gnd 0.08996f
C489 diffpairibias.n26 gnd 0.051736f
C490 diffpairibias.t24 gnd 0.08996f
C491 diffpairibias.n27 gnd 0.04729f
C492 diffpairibias.n28 gnd 0.047711f
C493 a_n1808_13878.t4 gnd 0.185683f
C494 a_n1808_13878.t0 gnd 0.185683f
C495 a_n1808_13878.t2 gnd 0.185683f
C496 a_n1808_13878.n0 gnd 1.46364f
C497 a_n1808_13878.t6 gnd 0.185683f
C498 a_n1808_13878.t1 gnd 0.185683f
C499 a_n1808_13878.n1 gnd 1.46209f
C500 a_n1808_13878.n2 gnd 2.04299f
C501 a_n1808_13878.t5 gnd 0.185683f
C502 a_n1808_13878.t9 gnd 0.185683f
C503 a_n1808_13878.n3 gnd 1.46451f
C504 a_n1808_13878.t10 gnd 0.185683f
C505 a_n1808_13878.t3 gnd 0.185683f
C506 a_n1808_13878.n4 gnd 1.46209f
C507 a_n1808_13878.n5 gnd 1.31424f
C508 a_n1808_13878.t7 gnd 0.185683f
C509 a_n1808_13878.t8 gnd 0.185683f
C510 a_n1808_13878.n6 gnd 1.46209f
C511 a_n1808_13878.n7 gnd 1.80499f
C512 a_n1808_13878.t13 gnd 1.73864f
C513 a_n1808_13878.t16 gnd 0.185683f
C514 a_n1808_13878.t17 gnd 0.185683f
C515 a_n1808_13878.n8 gnd 1.30795f
C516 a_n1808_13878.n9 gnd 1.46144f
C517 a_n1808_13878.t12 gnd 1.73518f
C518 a_n1808_13878.n10 gnd 0.735417f
C519 a_n1808_13878.t15 gnd 1.73518f
C520 a_n1808_13878.n11 gnd 0.735417f
C521 a_n1808_13878.t18 gnd 0.185683f
C522 a_n1808_13878.t19 gnd 0.185683f
C523 a_n1808_13878.n12 gnd 1.30795f
C524 a_n1808_13878.n13 gnd 0.742539f
C525 a_n1808_13878.t14 gnd 1.73518f
C526 a_n1808_13878.n14 gnd 1.73174f
C527 a_n1808_13878.n15 gnd 2.52099f
C528 a_n1808_13878.n16 gnd 3.70273f
C529 a_n1808_13878.n17 gnd 1.46209f
C530 a_n1808_13878.t11 gnd 0.185683f
C531 a_n1986_8322.t22 gnd 38.652897f
C532 a_n1986_8322.t20 gnd 28.1251f
C533 a_n1986_8322.t23 gnd 19.258501f
C534 a_n1986_8322.t21 gnd 38.652897f
C535 a_n1986_8322.t2 gnd 0.093486f
C536 a_n1986_8322.t1 gnd 0.875352f
C537 a_n1986_8322.t9 gnd 0.093486f
C538 a_n1986_8322.t4 gnd 0.093486f
C539 a_n1986_8322.n0 gnd 0.658513f
C540 a_n1986_8322.n1 gnd 0.735791f
C541 a_n1986_8322.t7 gnd 0.093486f
C542 a_n1986_8322.t6 gnd 0.093486f
C543 a_n1986_8322.n2 gnd 0.658513f
C544 a_n1986_8322.n3 gnd 0.373846f
C545 a_n1986_8322.t0 gnd 0.873609f
C546 a_n1986_8322.n4 gnd 1.39826f
C547 a_n1986_8322.t14 gnd 0.875352f
C548 a_n1986_8322.t18 gnd 0.093486f
C549 a_n1986_8322.t17 gnd 0.093486f
C550 a_n1986_8322.n5 gnd 0.658513f
C551 a_n1986_8322.n6 gnd 0.735791f
C552 a_n1986_8322.t12 gnd 0.873609f
C553 a_n1986_8322.n7 gnd 0.37026f
C554 a_n1986_8322.t15 gnd 0.873609f
C555 a_n1986_8322.n8 gnd 0.37026f
C556 a_n1986_8322.t13 gnd 0.093486f
C557 a_n1986_8322.t19 gnd 0.093486f
C558 a_n1986_8322.n9 gnd 0.658513f
C559 a_n1986_8322.n10 gnd 0.373846f
C560 a_n1986_8322.t16 gnd 0.873609f
C561 a_n1986_8322.n11 gnd 0.871879f
C562 a_n1986_8322.n12 gnd 1.58991f
C563 a_n1986_8322.n13 gnd 3.44798f
C564 a_n1986_8322.t3 gnd 0.873609f
C565 a_n1986_8322.n14 gnd 0.766135f
C566 a_n1986_8322.t10 gnd 0.875349f
C567 a_n1986_8322.t8 gnd 0.093486f
C568 a_n1986_8322.t5 gnd 0.093486f
C569 a_n1986_8322.n15 gnd 0.658513f
C570 a_n1986_8322.n16 gnd 0.735793f
C571 a_n1986_8322.n17 gnd 0.373844f
C572 a_n1986_8322.n18 gnd 0.658514f
C573 a_n1986_8322.t11 gnd 0.093486f
C574 a_n1996_n452.n0 gnd 0.822727f
C575 a_n1996_n452.n1 gnd 3.34433f
C576 a_n1996_n452.n2 gnd 3.17111f
C577 a_n1996_n452.n3 gnd 3.91594f
C578 a_n1996_n452.n4 gnd 0.527811f
C579 a_n1996_n452.n5 gnd 0.205584f
C580 a_n1996_n452.n6 gnd 0.151417f
C581 a_n1996_n452.n7 gnd 0.237979f
C582 a_n1996_n452.n8 gnd 0.183812f
C583 a_n1996_n452.n9 gnd 0.205584f
C584 a_n1996_n452.n10 gnd 1.00969f
C585 a_n1996_n452.n11 gnd 0.151417f
C586 a_n1996_n452.n12 gnd 0.581979f
C587 a_n1996_n452.n13 gnd 0.433746f
C588 a_n1996_n452.n14 gnd 0.21667f
C589 a_n1996_n452.n15 gnd 0.494132f
C590 a_n1996_n452.n16 gnd 0.283464f
C591 a_n1996_n452.n17 gnd 0.439964f
C592 a_n1996_n452.n18 gnd 0.21667f
C593 a_n1996_n452.n19 gnd 0.734001f
C594 a_n1996_n452.n20 gnd 0.283464f
C595 a_n1996_n452.n21 gnd 0.494132f
C596 a_n1996_n452.n22 gnd 0.666675f
C597 a_n1996_n452.n23 gnd 0.21667f
C598 a_n1996_n452.n24 gnd 0.283464f
C599 a_n1996_n452.n25 gnd 0.641354f
C600 a_n1996_n452.n26 gnd 0.283464f
C601 a_n1996_n452.n27 gnd 1.18284f
C602 a_n1996_n452.n28 gnd 1.92214f
C603 a_n1996_n452.n29 gnd 1.14844f
C604 a_n1996_n452.n30 gnd 1.78382f
C605 a_n1996_n452.n31 gnd 3.22512f
C606 a_n1996_n452.n32 gnd 0.108335f
C607 a_n1996_n452.n33 gnd 0.008389f
C608 a_n1996_n452.n35 gnd 0.008389f
C609 a_n1996_n452.n37 gnd 0.286629f
C610 a_n1996_n452.n38 gnd 0.008389f
C611 a_n1996_n452.n40 gnd 0.286629f
C612 a_n1996_n452.n41 gnd 0.008389f
C613 a_n1996_n452.n43 gnd 0.286629f
C614 a_n1996_n452.n44 gnd 0.008389f
C615 a_n1996_n452.n45 gnd 0.286221f
C616 a_n1996_n452.n46 gnd 0.008389f
C617 a_n1996_n452.n47 gnd 0.286221f
C618 a_n1996_n452.n48 gnd 0.008389f
C619 a_n1996_n452.n49 gnd 0.286221f
C620 a_n1996_n452.n50 gnd 0.008389f
C621 a_n1996_n452.n51 gnd 0.286221f
C622 a_n1996_n452.n52 gnd 0.286629f
C623 a_n1996_n452.t8 gnd 0.150285f
C624 a_n1996_n452.t5 gnd 0.713776f
C625 a_n1996_n452.t3 gnd 0.699053f
C626 a_n1996_n452.t7 gnd 0.699053f
C627 a_n1996_n452.t11 gnd 0.699053f
C628 a_n1996_n452.n53 gnd 0.307348f
C629 a_n1996_n452.t19 gnd 0.710611f
C630 a_n1996_n452.t31 gnd 0.116888f
C631 a_n1996_n452.t42 gnd 0.116888f
C632 a_n1996_n452.n54 gnd 1.03516f
C633 a_n1996_n452.t38 gnd 0.116888f
C634 a_n1996_n452.t34 gnd 0.116888f
C635 a_n1996_n452.n55 gnd 1.03287f
C636 a_n1996_n452.t36 gnd 0.116888f
C637 a_n1996_n452.t27 gnd 0.116888f
C638 a_n1996_n452.n56 gnd 1.03287f
C639 a_n1996_n452.t40 gnd 0.116888f
C640 a_n1996_n452.t37 gnd 0.116888f
C641 a_n1996_n452.n57 gnd 1.03516f
C642 a_n1996_n452.t1 gnd 0.116888f
C643 a_n1996_n452.t0 gnd 0.116888f
C644 a_n1996_n452.n58 gnd 1.03287f
C645 a_n1996_n452.t39 gnd 0.116888f
C646 a_n1996_n452.t35 gnd 0.116888f
C647 a_n1996_n452.n59 gnd 1.03287f
C648 a_n1996_n452.t32 gnd 0.116888f
C649 a_n1996_n452.t33 gnd 0.116888f
C650 a_n1996_n452.n60 gnd 1.03287f
C651 a_n1996_n452.t2 gnd 0.116888f
C652 a_n1996_n452.t30 gnd 0.116888f
C653 a_n1996_n452.n61 gnd 1.03287f
C654 a_n1996_n452.t41 gnd 0.116888f
C655 a_n1996_n452.t43 gnd 0.116888f
C656 a_n1996_n452.n62 gnd 1.03516f
C657 a_n1996_n452.t28 gnd 0.116888f
C658 a_n1996_n452.t29 gnd 0.116888f
C659 a_n1996_n452.n63 gnd 1.03287f
C660 a_n1996_n452.t71 gnd 0.713776f
C661 a_n1996_n452.t54 gnd 0.699053f
C662 a_n1996_n452.t58 gnd 0.699053f
C663 a_n1996_n452.t48 gnd 0.699053f
C664 a_n1996_n452.n64 gnd 0.307348f
C665 a_n1996_n452.t63 gnd 0.699053f
C666 a_n1996_n452.t69 gnd 0.710611f
C667 a_n1996_n452.t22 gnd 1.40719f
C668 a_n1996_n452.t10 gnd 0.150285f
C669 a_n1996_n452.t26 gnd 0.150285f
C670 a_n1996_n452.n65 gnd 1.05861f
C671 a_n1996_n452.t16 gnd 0.150285f
C672 a_n1996_n452.t14 gnd 0.150285f
C673 a_n1996_n452.n66 gnd 1.05861f
C674 a_n1996_n452.t24 gnd 1.40439f
C675 a_n1996_n452.t15 gnd 0.699053f
C676 a_n1996_n452.n67 gnd 0.307348f
C677 a_n1996_n452.t13 gnd 0.699053f
C678 a_n1996_n452.t9 gnd 0.699053f
C679 a_n1996_n452.t52 gnd 0.699053f
C680 a_n1996_n452.n68 gnd 0.307348f
C681 a_n1996_n452.t61 gnd 0.699053f
C682 a_n1996_n452.t67 gnd 0.699053f
C683 a_n1996_n452.t66 gnd 0.713776f
C684 a_n1996_n452.n69 gnd 0.309974f
C685 a_n1996_n452.t46 gnd 0.699053f
C686 a_n1996_n452.n70 gnd 0.303445f
C687 a_n1996_n452.n71 gnd 0.309974f
C688 a_n1996_n452.t47 gnd 0.710611f
C689 a_n1996_n452.t21 gnd 0.713776f
C690 a_n1996_n452.n72 gnd 0.309974f
C691 a_n1996_n452.t25 gnd 0.699053f
C692 a_n1996_n452.n73 gnd 0.303445f
C693 a_n1996_n452.n74 gnd 0.309974f
C694 a_n1996_n452.t23 gnd 0.710611f
C695 a_n1996_n452.n75 gnd 1.13585f
C696 a_n1996_n452.t51 gnd 0.699053f
C697 a_n1996_n452.n76 gnd 0.303445f
C698 a_n1996_n452.t57 gnd 0.699053f
C699 a_n1996_n452.n77 gnd 0.303445f
C700 a_n1996_n452.t49 gnd 0.699053f
C701 a_n1996_n452.n78 gnd 0.303445f
C702 a_n1996_n452.t62 gnd 0.699053f
C703 a_n1996_n452.n79 gnd 0.303445f
C704 a_n1996_n452.t53 gnd 0.699053f
C705 a_n1996_n452.n80 gnd 0.297934f
C706 a_n1996_n452.t44 gnd 0.699053f
C707 a_n1996_n452.n81 gnd 0.307348f
C708 a_n1996_n452.t55 gnd 0.710766f
C709 a_n1996_n452.t64 gnd 0.699053f
C710 a_n1996_n452.n82 gnd 0.297934f
C711 a_n1996_n452.t50 gnd 0.699053f
C712 a_n1996_n452.n83 gnd 0.307348f
C713 a_n1996_n452.t59 gnd 0.710766f
C714 a_n1996_n452.t68 gnd 0.699053f
C715 a_n1996_n452.n84 gnd 0.297934f
C716 a_n1996_n452.t56 gnd 0.699053f
C717 a_n1996_n452.n85 gnd 0.307348f
C718 a_n1996_n452.t70 gnd 0.710766f
C719 a_n1996_n452.t60 gnd 0.699053f
C720 a_n1996_n452.n86 gnd 0.297934f
C721 a_n1996_n452.t45 gnd 0.699053f
C722 a_n1996_n452.n87 gnd 0.307348f
C723 a_n1996_n452.t65 gnd 0.710766f
C724 a_n1996_n452.n88 gnd 1.34296f
C725 a_n1996_n452.n89 gnd 0.309974f
C726 a_n1996_n452.n90 gnd 0.303445f
C727 a_n1996_n452.n91 gnd 0.309974f
C728 a_n1996_n452.t17 gnd 0.699053f
C729 a_n1996_n452.n92 gnd 0.309974f
C730 a_n1996_n452.n93 gnd 0.303445f
C731 a_n1996_n452.n94 gnd 0.309974f
C732 a_n1996_n452.n95 gnd 0.789588f
C733 a_n1996_n452.t6 gnd 1.40439f
C734 a_n1996_n452.t20 gnd 1.40719f
C735 a_n1996_n452.t12 gnd 0.150285f
C736 a_n1996_n452.t18 gnd 0.150285f
C737 a_n1996_n452.n96 gnd 1.05861f
C738 a_n1996_n452.n97 gnd 1.05861f
C739 a_n1996_n452.t4 gnd 0.150285f
C740 vdd.t193 gnd 0.032948f
C741 vdd.t177 gnd 0.032948f
C742 vdd.n0 gnd 0.259864f
C743 vdd.t184 gnd 0.032948f
C744 vdd.t187 gnd 0.032948f
C745 vdd.n1 gnd 0.259435f
C746 vdd.n2 gnd 0.239248f
C747 vdd.t75 gnd 0.032948f
C748 vdd.t3 gnd 0.032948f
C749 vdd.n3 gnd 0.259435f
C750 vdd.n4 gnd 0.120997f
C751 vdd.t5 gnd 0.032948f
C752 vdd.t80 gnd 0.032948f
C753 vdd.n5 gnd 0.259435f
C754 vdd.n6 gnd 0.113533f
C755 vdd.t195 gnd 0.032948f
C756 vdd.t1 gnd 0.032948f
C757 vdd.n7 gnd 0.259864f
C758 vdd.t190 gnd 0.032948f
C759 vdd.t180 gnd 0.032948f
C760 vdd.n8 gnd 0.259435f
C761 vdd.n9 gnd 0.239248f
C762 vdd.t199 gnd 0.032948f
C763 vdd.t8 gnd 0.032948f
C764 vdd.n10 gnd 0.259435f
C765 vdd.n11 gnd 0.120997f
C766 vdd.t182 gnd 0.032948f
C767 vdd.t197 gnd 0.032948f
C768 vdd.n12 gnd 0.259435f
C769 vdd.n13 gnd 0.113533f
C770 vdd.n14 gnd 0.080266f
C771 vdd.t165 gnd 0.018304f
C772 vdd.t168 gnd 0.018304f
C773 vdd.n15 gnd 0.168483f
C774 vdd.t157 gnd 0.018304f
C775 vdd.t158 gnd 0.018304f
C776 vdd.n16 gnd 0.16799f
C777 vdd.n17 gnd 0.292355f
C778 vdd.t161 gnd 0.018304f
C779 vdd.t160 gnd 0.018304f
C780 vdd.n18 gnd 0.16799f
C781 vdd.n19 gnd 0.120951f
C782 vdd.t166 gnd 0.018304f
C783 vdd.t167 gnd 0.018304f
C784 vdd.n20 gnd 0.168483f
C785 vdd.t171 gnd 0.018304f
C786 vdd.t164 gnd 0.018304f
C787 vdd.n21 gnd 0.16799f
C788 vdd.n22 gnd 0.292355f
C789 vdd.t170 gnd 0.018304f
C790 vdd.t169 gnd 0.018304f
C791 vdd.n23 gnd 0.16799f
C792 vdd.n24 gnd 0.120951f
C793 vdd.t159 gnd 0.018304f
C794 vdd.t172 gnd 0.018304f
C795 vdd.n25 gnd 0.16799f
C796 vdd.t163 gnd 0.018304f
C797 vdd.t162 gnd 0.018304f
C798 vdd.n26 gnd 0.16799f
C799 vdd.n27 gnd 18.392f
C800 vdd.n28 gnd 6.85872f
C801 vdd.n29 gnd 0.004992f
C802 vdd.n30 gnd 0.004633f
C803 vdd.n31 gnd 0.002563f
C804 vdd.n32 gnd 0.005884f
C805 vdd.n33 gnd 0.002489f
C806 vdd.n34 gnd 0.002636f
C807 vdd.n35 gnd 0.004633f
C808 vdd.n36 gnd 0.002489f
C809 vdd.n37 gnd 0.005884f
C810 vdd.n38 gnd 0.002636f
C811 vdd.n39 gnd 0.004633f
C812 vdd.n40 gnd 0.002489f
C813 vdd.n41 gnd 0.004413f
C814 vdd.n42 gnd 0.004426f
C815 vdd.t13 gnd 0.012641f
C816 vdd.n43 gnd 0.028127f
C817 vdd.n44 gnd 0.146377f
C818 vdd.n45 gnd 0.002489f
C819 vdd.n46 gnd 0.002636f
C820 vdd.n47 gnd 0.005884f
C821 vdd.n48 gnd 0.005884f
C822 vdd.n49 gnd 0.002636f
C823 vdd.n50 gnd 0.002489f
C824 vdd.n51 gnd 0.004633f
C825 vdd.n52 gnd 0.004633f
C826 vdd.n53 gnd 0.002489f
C827 vdd.n54 gnd 0.002636f
C828 vdd.n55 gnd 0.005884f
C829 vdd.n56 gnd 0.005884f
C830 vdd.n57 gnd 0.002636f
C831 vdd.n58 gnd 0.002489f
C832 vdd.n59 gnd 0.004633f
C833 vdd.n60 gnd 0.004633f
C834 vdd.n61 gnd 0.002489f
C835 vdd.n62 gnd 0.002636f
C836 vdd.n63 gnd 0.005884f
C837 vdd.n64 gnd 0.005884f
C838 vdd.n65 gnd 0.013911f
C839 vdd.n66 gnd 0.002563f
C840 vdd.n67 gnd 0.002489f
C841 vdd.n68 gnd 0.011974f
C842 vdd.n69 gnd 0.008359f
C843 vdd.t65 gnd 0.029287f
C844 vdd.t39 gnd 0.029287f
C845 vdd.n70 gnd 0.201279f
C846 vdd.n71 gnd 0.158275f
C847 vdd.t72 gnd 0.029287f
C848 vdd.t28 gnd 0.029287f
C849 vdd.n72 gnd 0.201279f
C850 vdd.n73 gnd 0.127727f
C851 vdd.t58 gnd 0.029287f
C852 vdd.t33 gnd 0.029287f
C853 vdd.n74 gnd 0.201279f
C854 vdd.n75 gnd 0.127727f
C855 vdd.n76 gnd 0.004992f
C856 vdd.n77 gnd 0.004633f
C857 vdd.n78 gnd 0.002563f
C858 vdd.n79 gnd 0.005884f
C859 vdd.n80 gnd 0.002489f
C860 vdd.n81 gnd 0.002636f
C861 vdd.n82 gnd 0.004633f
C862 vdd.n83 gnd 0.002489f
C863 vdd.n84 gnd 0.005884f
C864 vdd.n85 gnd 0.002636f
C865 vdd.n86 gnd 0.004633f
C866 vdd.n87 gnd 0.002489f
C867 vdd.n88 gnd 0.004413f
C868 vdd.n89 gnd 0.004426f
C869 vdd.t71 gnd 0.012641f
C870 vdd.n90 gnd 0.028127f
C871 vdd.n91 gnd 0.146377f
C872 vdd.n92 gnd 0.002489f
C873 vdd.n93 gnd 0.002636f
C874 vdd.n94 gnd 0.005884f
C875 vdd.n95 gnd 0.005884f
C876 vdd.n96 gnd 0.002636f
C877 vdd.n97 gnd 0.002489f
C878 vdd.n98 gnd 0.004633f
C879 vdd.n99 gnd 0.004633f
C880 vdd.n100 gnd 0.002489f
C881 vdd.n101 gnd 0.002636f
C882 vdd.n102 gnd 0.005884f
C883 vdd.n103 gnd 0.005884f
C884 vdd.n104 gnd 0.002636f
C885 vdd.n105 gnd 0.002489f
C886 vdd.n106 gnd 0.004633f
C887 vdd.n107 gnd 0.004633f
C888 vdd.n108 gnd 0.002489f
C889 vdd.n109 gnd 0.002636f
C890 vdd.n110 gnd 0.005884f
C891 vdd.n111 gnd 0.005884f
C892 vdd.n112 gnd 0.013911f
C893 vdd.n113 gnd 0.002563f
C894 vdd.n114 gnd 0.002489f
C895 vdd.n115 gnd 0.011974f
C896 vdd.n116 gnd 0.008097f
C897 vdd.n117 gnd 0.09503f
C898 vdd.n118 gnd 0.004992f
C899 vdd.n119 gnd 0.004633f
C900 vdd.n120 gnd 0.002563f
C901 vdd.n121 gnd 0.005884f
C902 vdd.n122 gnd 0.002489f
C903 vdd.n123 gnd 0.002636f
C904 vdd.n124 gnd 0.004633f
C905 vdd.n125 gnd 0.002489f
C906 vdd.n126 gnd 0.005884f
C907 vdd.n127 gnd 0.002636f
C908 vdd.n128 gnd 0.004633f
C909 vdd.n129 gnd 0.002489f
C910 vdd.n130 gnd 0.004413f
C911 vdd.n131 gnd 0.004426f
C912 vdd.t40 gnd 0.012641f
C913 vdd.n132 gnd 0.028127f
C914 vdd.n133 gnd 0.146377f
C915 vdd.n134 gnd 0.002489f
C916 vdd.n135 gnd 0.002636f
C917 vdd.n136 gnd 0.005884f
C918 vdd.n137 gnd 0.005884f
C919 vdd.n138 gnd 0.002636f
C920 vdd.n139 gnd 0.002489f
C921 vdd.n140 gnd 0.004633f
C922 vdd.n141 gnd 0.004633f
C923 vdd.n142 gnd 0.002489f
C924 vdd.n143 gnd 0.002636f
C925 vdd.n144 gnd 0.005884f
C926 vdd.n145 gnd 0.005884f
C927 vdd.n146 gnd 0.002636f
C928 vdd.n147 gnd 0.002489f
C929 vdd.n148 gnd 0.004633f
C930 vdd.n149 gnd 0.004633f
C931 vdd.n150 gnd 0.002489f
C932 vdd.n151 gnd 0.002636f
C933 vdd.n152 gnd 0.005884f
C934 vdd.n153 gnd 0.005884f
C935 vdd.n154 gnd 0.013911f
C936 vdd.n155 gnd 0.002563f
C937 vdd.n156 gnd 0.002489f
C938 vdd.n157 gnd 0.011974f
C939 vdd.n158 gnd 0.008359f
C940 vdd.t42 gnd 0.029287f
C941 vdd.t53 gnd 0.029287f
C942 vdd.n159 gnd 0.201279f
C943 vdd.n160 gnd 0.158275f
C944 vdd.t17 gnd 0.029287f
C945 vdd.t36 gnd 0.029287f
C946 vdd.n161 gnd 0.201279f
C947 vdd.n162 gnd 0.127727f
C948 vdd.t52 gnd 0.029287f
C949 vdd.t73 gnd 0.029287f
C950 vdd.n163 gnd 0.201279f
C951 vdd.n164 gnd 0.127727f
C952 vdd.n165 gnd 0.004992f
C953 vdd.n166 gnd 0.004633f
C954 vdd.n167 gnd 0.002563f
C955 vdd.n168 gnd 0.005884f
C956 vdd.n169 gnd 0.002489f
C957 vdd.n170 gnd 0.002636f
C958 vdd.n171 gnd 0.004633f
C959 vdd.n172 gnd 0.002489f
C960 vdd.n173 gnd 0.005884f
C961 vdd.n174 gnd 0.002636f
C962 vdd.n175 gnd 0.004633f
C963 vdd.n176 gnd 0.002489f
C964 vdd.n177 gnd 0.004413f
C965 vdd.n178 gnd 0.004426f
C966 vdd.t30 gnd 0.012641f
C967 vdd.n179 gnd 0.028127f
C968 vdd.n180 gnd 0.146377f
C969 vdd.n181 gnd 0.002489f
C970 vdd.n182 gnd 0.002636f
C971 vdd.n183 gnd 0.005884f
C972 vdd.n184 gnd 0.005884f
C973 vdd.n185 gnd 0.002636f
C974 vdd.n186 gnd 0.002489f
C975 vdd.n187 gnd 0.004633f
C976 vdd.n188 gnd 0.004633f
C977 vdd.n189 gnd 0.002489f
C978 vdd.n190 gnd 0.002636f
C979 vdd.n191 gnd 0.005884f
C980 vdd.n192 gnd 0.005884f
C981 vdd.n193 gnd 0.002636f
C982 vdd.n194 gnd 0.002489f
C983 vdd.n195 gnd 0.004633f
C984 vdd.n196 gnd 0.004633f
C985 vdd.n197 gnd 0.002489f
C986 vdd.n198 gnd 0.002636f
C987 vdd.n199 gnd 0.005884f
C988 vdd.n200 gnd 0.005884f
C989 vdd.n201 gnd 0.013911f
C990 vdd.n202 gnd 0.002563f
C991 vdd.n203 gnd 0.002489f
C992 vdd.n204 gnd 0.011974f
C993 vdd.n205 gnd 0.008097f
C994 vdd.n206 gnd 0.056533f
C995 vdd.n207 gnd 0.203704f
C996 vdd.n208 gnd 0.004992f
C997 vdd.n209 gnd 0.004633f
C998 vdd.n210 gnd 0.002563f
C999 vdd.n211 gnd 0.005884f
C1000 vdd.n212 gnd 0.002489f
C1001 vdd.n213 gnd 0.002636f
C1002 vdd.n214 gnd 0.004633f
C1003 vdd.n215 gnd 0.002489f
C1004 vdd.n216 gnd 0.005884f
C1005 vdd.n217 gnd 0.002636f
C1006 vdd.n218 gnd 0.004633f
C1007 vdd.n219 gnd 0.002489f
C1008 vdd.n220 gnd 0.004413f
C1009 vdd.n221 gnd 0.004426f
C1010 vdd.t45 gnd 0.012641f
C1011 vdd.n222 gnd 0.028127f
C1012 vdd.n223 gnd 0.146377f
C1013 vdd.n224 gnd 0.002489f
C1014 vdd.n225 gnd 0.002636f
C1015 vdd.n226 gnd 0.005884f
C1016 vdd.n227 gnd 0.005884f
C1017 vdd.n228 gnd 0.002636f
C1018 vdd.n229 gnd 0.002489f
C1019 vdd.n230 gnd 0.004633f
C1020 vdd.n231 gnd 0.004633f
C1021 vdd.n232 gnd 0.002489f
C1022 vdd.n233 gnd 0.002636f
C1023 vdd.n234 gnd 0.005884f
C1024 vdd.n235 gnd 0.005884f
C1025 vdd.n236 gnd 0.002636f
C1026 vdd.n237 gnd 0.002489f
C1027 vdd.n238 gnd 0.004633f
C1028 vdd.n239 gnd 0.004633f
C1029 vdd.n240 gnd 0.002489f
C1030 vdd.n241 gnd 0.002636f
C1031 vdd.n242 gnd 0.005884f
C1032 vdd.n243 gnd 0.005884f
C1033 vdd.n244 gnd 0.013911f
C1034 vdd.n245 gnd 0.002563f
C1035 vdd.n246 gnd 0.002489f
C1036 vdd.n247 gnd 0.011974f
C1037 vdd.n248 gnd 0.008359f
C1038 vdd.t46 gnd 0.029287f
C1039 vdd.t62 gnd 0.029287f
C1040 vdd.n249 gnd 0.201279f
C1041 vdd.n250 gnd 0.158275f
C1042 vdd.t23 gnd 0.029287f
C1043 vdd.t44 gnd 0.029287f
C1044 vdd.n251 gnd 0.201279f
C1045 vdd.n252 gnd 0.127727f
C1046 vdd.t57 gnd 0.029287f
C1047 vdd.t21 gnd 0.029287f
C1048 vdd.n253 gnd 0.201279f
C1049 vdd.n254 gnd 0.127727f
C1050 vdd.n255 gnd 0.004992f
C1051 vdd.n256 gnd 0.004633f
C1052 vdd.n257 gnd 0.002563f
C1053 vdd.n258 gnd 0.005884f
C1054 vdd.n259 gnd 0.002489f
C1055 vdd.n260 gnd 0.002636f
C1056 vdd.n261 gnd 0.004633f
C1057 vdd.n262 gnd 0.002489f
C1058 vdd.n263 gnd 0.005884f
C1059 vdd.n264 gnd 0.002636f
C1060 vdd.n265 gnd 0.004633f
C1061 vdd.n266 gnd 0.002489f
C1062 vdd.n267 gnd 0.004413f
C1063 vdd.n268 gnd 0.004426f
C1064 vdd.t34 gnd 0.012641f
C1065 vdd.n269 gnd 0.028127f
C1066 vdd.n270 gnd 0.146377f
C1067 vdd.n271 gnd 0.002489f
C1068 vdd.n272 gnd 0.002636f
C1069 vdd.n273 gnd 0.005884f
C1070 vdd.n274 gnd 0.005884f
C1071 vdd.n275 gnd 0.002636f
C1072 vdd.n276 gnd 0.002489f
C1073 vdd.n277 gnd 0.004633f
C1074 vdd.n278 gnd 0.004633f
C1075 vdd.n279 gnd 0.002489f
C1076 vdd.n280 gnd 0.002636f
C1077 vdd.n281 gnd 0.005884f
C1078 vdd.n282 gnd 0.005884f
C1079 vdd.n283 gnd 0.002636f
C1080 vdd.n284 gnd 0.002489f
C1081 vdd.n285 gnd 0.004633f
C1082 vdd.n286 gnd 0.004633f
C1083 vdd.n287 gnd 0.002489f
C1084 vdd.n288 gnd 0.002636f
C1085 vdd.n289 gnd 0.005884f
C1086 vdd.n290 gnd 0.005884f
C1087 vdd.n291 gnd 0.013911f
C1088 vdd.n292 gnd 0.002563f
C1089 vdd.n293 gnd 0.002489f
C1090 vdd.n294 gnd 0.011974f
C1091 vdd.n295 gnd 0.008097f
C1092 vdd.n296 gnd 0.056533f
C1093 vdd.n297 gnd 0.220485f
C1094 vdd.n298 gnd 0.006991f
C1095 vdd.n299 gnd 0.009097f
C1096 vdd.n300 gnd 0.007322f
C1097 vdd.n301 gnd 0.007322f
C1098 vdd.n302 gnd 0.009097f
C1099 vdd.n303 gnd 0.009097f
C1100 vdd.n304 gnd 0.664689f
C1101 vdd.n305 gnd 0.009097f
C1102 vdd.n306 gnd 0.009097f
C1103 vdd.n307 gnd 0.009097f
C1104 vdd.n308 gnd 0.720467f
C1105 vdd.n309 gnd 0.009097f
C1106 vdd.n310 gnd 0.009097f
C1107 vdd.n311 gnd 0.009097f
C1108 vdd.n312 gnd 0.009097f
C1109 vdd.n313 gnd 0.007322f
C1110 vdd.n314 gnd 0.009097f
C1111 vdd.t20 gnd 0.464817f
C1112 vdd.n315 gnd 0.009097f
C1113 vdd.n316 gnd 0.009097f
C1114 vdd.n317 gnd 0.009097f
C1115 vdd.n318 gnd 0.929634f
C1116 vdd.n319 gnd 0.009097f
C1117 vdd.n320 gnd 0.009097f
C1118 vdd.n321 gnd 0.009097f
C1119 vdd.n322 gnd 0.009097f
C1120 vdd.n323 gnd 0.009097f
C1121 vdd.n324 gnd 0.007322f
C1122 vdd.n325 gnd 0.009097f
C1123 vdd.n326 gnd 0.009097f
C1124 vdd.n327 gnd 0.009097f
C1125 vdd.n328 gnd 0.022169f
C1126 vdd.n329 gnd 2.22183f
C1127 vdd.n330 gnd 0.022678f
C1128 vdd.n331 gnd 0.009097f
C1129 vdd.n332 gnd 0.009097f
C1130 vdd.n334 gnd 0.009097f
C1131 vdd.n335 gnd 0.009097f
C1132 vdd.n336 gnd 0.007322f
C1133 vdd.n337 gnd 0.007322f
C1134 vdd.n338 gnd 0.009097f
C1135 vdd.n339 gnd 0.009097f
C1136 vdd.n340 gnd 0.009097f
C1137 vdd.n341 gnd 0.009097f
C1138 vdd.n342 gnd 0.009097f
C1139 vdd.n343 gnd 0.009097f
C1140 vdd.n344 gnd 0.007322f
C1141 vdd.n346 gnd 0.009097f
C1142 vdd.n347 gnd 0.009097f
C1143 vdd.n348 gnd 0.009097f
C1144 vdd.n349 gnd 0.009097f
C1145 vdd.n350 gnd 0.009097f
C1146 vdd.n351 gnd 0.007322f
C1147 vdd.n353 gnd 0.009097f
C1148 vdd.n354 gnd 0.009097f
C1149 vdd.n355 gnd 0.009097f
C1150 vdd.n356 gnd 0.009097f
C1151 vdd.n357 gnd 0.009097f
C1152 vdd.n358 gnd 0.007322f
C1153 vdd.n360 gnd 0.009097f
C1154 vdd.n361 gnd 0.009097f
C1155 vdd.n362 gnd 0.009097f
C1156 vdd.n363 gnd 0.009097f
C1157 vdd.n364 gnd 0.006114f
C1158 vdd.t112 gnd 0.111913f
C1159 vdd.t111 gnd 0.119604f
C1160 vdd.t110 gnd 0.146157f
C1161 vdd.n365 gnd 0.187352f
C1162 vdd.n366 gnd 0.158142f
C1163 vdd.n368 gnd 0.009097f
C1164 vdd.n369 gnd 0.009097f
C1165 vdd.n370 gnd 0.007322f
C1166 vdd.n371 gnd 0.009097f
C1167 vdd.n373 gnd 0.009097f
C1168 vdd.n374 gnd 0.009097f
C1169 vdd.n375 gnd 0.009097f
C1170 vdd.n376 gnd 0.009097f
C1171 vdd.n377 gnd 0.007322f
C1172 vdd.n379 gnd 0.009097f
C1173 vdd.n380 gnd 0.009097f
C1174 vdd.n381 gnd 0.009097f
C1175 vdd.n382 gnd 0.009097f
C1176 vdd.n383 gnd 0.009097f
C1177 vdd.n384 gnd 0.007322f
C1178 vdd.n386 gnd 0.009097f
C1179 vdd.n387 gnd 0.009097f
C1180 vdd.n388 gnd 0.009097f
C1181 vdd.n389 gnd 0.009097f
C1182 vdd.n390 gnd 0.009097f
C1183 vdd.n391 gnd 0.007322f
C1184 vdd.n393 gnd 0.009097f
C1185 vdd.n394 gnd 0.009097f
C1186 vdd.n395 gnd 0.009097f
C1187 vdd.n396 gnd 0.009097f
C1188 vdd.n397 gnd 0.009097f
C1189 vdd.n398 gnd 0.007322f
C1190 vdd.n400 gnd 0.009097f
C1191 vdd.n401 gnd 0.009097f
C1192 vdd.n402 gnd 0.009097f
C1193 vdd.n403 gnd 0.009097f
C1194 vdd.n404 gnd 0.007248f
C1195 vdd.t106 gnd 0.111913f
C1196 vdd.t105 gnd 0.119604f
C1197 vdd.t103 gnd 0.146157f
C1198 vdd.n405 gnd 0.187352f
C1199 vdd.n406 gnd 0.158142f
C1200 vdd.n408 gnd 0.009097f
C1201 vdd.n409 gnd 0.009097f
C1202 vdd.n410 gnd 0.007322f
C1203 vdd.n411 gnd 0.009097f
C1204 vdd.n413 gnd 0.009097f
C1205 vdd.n414 gnd 0.009097f
C1206 vdd.n415 gnd 0.009097f
C1207 vdd.n416 gnd 0.009097f
C1208 vdd.n417 gnd 0.007322f
C1209 vdd.n419 gnd 0.009097f
C1210 vdd.n420 gnd 0.009097f
C1211 vdd.n421 gnd 0.009097f
C1212 vdd.n422 gnd 0.009097f
C1213 vdd.n423 gnd 0.009097f
C1214 vdd.n424 gnd 0.007322f
C1215 vdd.n426 gnd 0.009097f
C1216 vdd.n427 gnd 0.009097f
C1217 vdd.n428 gnd 0.009097f
C1218 vdd.n429 gnd 0.009097f
C1219 vdd.n430 gnd 0.009097f
C1220 vdd.n431 gnd 0.007322f
C1221 vdd.n433 gnd 0.009097f
C1222 vdd.n434 gnd 0.009097f
C1223 vdd.n435 gnd 0.009097f
C1224 vdd.n436 gnd 0.009097f
C1225 vdd.n437 gnd 0.009097f
C1226 vdd.n438 gnd 0.007322f
C1227 vdd.n440 gnd 0.009097f
C1228 vdd.n441 gnd 0.009097f
C1229 vdd.n442 gnd 0.009097f
C1230 vdd.n443 gnd 0.009097f
C1231 vdd.n444 gnd 0.009097f
C1232 vdd.n445 gnd 0.009097f
C1233 vdd.n446 gnd 0.007322f
C1234 vdd.n447 gnd 0.009097f
C1235 vdd.n448 gnd 0.009097f
C1236 vdd.n449 gnd 0.007322f
C1237 vdd.n450 gnd 0.009097f
C1238 vdd.n451 gnd 0.007322f
C1239 vdd.n452 gnd 0.009097f
C1240 vdd.n453 gnd 0.007322f
C1241 vdd.n454 gnd 0.009097f
C1242 vdd.n455 gnd 0.009097f
C1243 vdd.n456 gnd 0.506651f
C1244 vdd.t16 gnd 0.464817f
C1245 vdd.n457 gnd 0.009097f
C1246 vdd.n458 gnd 0.007322f
C1247 vdd.n459 gnd 0.009097f
C1248 vdd.n460 gnd 0.007322f
C1249 vdd.n461 gnd 0.009097f
C1250 vdd.t41 gnd 0.464817f
C1251 vdd.n462 gnd 0.009097f
C1252 vdd.n463 gnd 0.007322f
C1253 vdd.n464 gnd 0.009097f
C1254 vdd.n465 gnd 0.007322f
C1255 vdd.n466 gnd 0.009097f
C1256 vdd.t12 gnd 0.464817f
C1257 vdd.n467 gnd 0.581022f
C1258 vdd.n468 gnd 0.009097f
C1259 vdd.n469 gnd 0.007322f
C1260 vdd.n470 gnd 0.009097f
C1261 vdd.n471 gnd 0.007322f
C1262 vdd.n472 gnd 0.009097f
C1263 vdd.n473 gnd 0.929634f
C1264 vdd.n474 gnd 0.009097f
C1265 vdd.n475 gnd 0.007322f
C1266 vdd.n476 gnd 0.022169f
C1267 vdd.n477 gnd 0.006077f
C1268 vdd.n478 gnd 0.022169f
C1269 vdd.t82 gnd 0.464817f
C1270 vdd.n479 gnd 0.022169f
C1271 vdd.n480 gnd 0.006077f
C1272 vdd.n481 gnd 0.007823f
C1273 vdd.n482 gnd 0.007322f
C1274 vdd.n483 gnd 0.009097f
C1275 vdd.n484 gnd 6.40518f
C1276 vdd.n515 gnd 0.022678f
C1277 vdd.n516 gnd 1.27825f
C1278 vdd.n517 gnd 0.009097f
C1279 vdd.n518 gnd 0.007322f
C1280 vdd.n519 gnd 0.005822f
C1281 vdd.n520 gnd 0.014864f
C1282 vdd.n521 gnd 0.007322f
C1283 vdd.n522 gnd 0.009097f
C1284 vdd.n523 gnd 0.009097f
C1285 vdd.n524 gnd 0.009097f
C1286 vdd.n525 gnd 0.009097f
C1287 vdd.n526 gnd 0.009097f
C1288 vdd.n527 gnd 0.009097f
C1289 vdd.n528 gnd 0.009097f
C1290 vdd.n529 gnd 0.009097f
C1291 vdd.n530 gnd 0.009097f
C1292 vdd.n531 gnd 0.009097f
C1293 vdd.n532 gnd 0.009097f
C1294 vdd.n533 gnd 0.009097f
C1295 vdd.n534 gnd 0.009097f
C1296 vdd.n535 gnd 0.009097f
C1297 vdd.n536 gnd 0.006114f
C1298 vdd.n537 gnd 0.009097f
C1299 vdd.n538 gnd 0.009097f
C1300 vdd.n539 gnd 0.009097f
C1301 vdd.n540 gnd 0.009097f
C1302 vdd.n541 gnd 0.009097f
C1303 vdd.n542 gnd 0.009097f
C1304 vdd.n543 gnd 0.009097f
C1305 vdd.n544 gnd 0.009097f
C1306 vdd.n545 gnd 0.009097f
C1307 vdd.n546 gnd 0.009097f
C1308 vdd.n547 gnd 0.009097f
C1309 vdd.n548 gnd 0.009097f
C1310 vdd.n549 gnd 0.009097f
C1311 vdd.n550 gnd 0.009097f
C1312 vdd.n551 gnd 0.009097f
C1313 vdd.n552 gnd 0.009097f
C1314 vdd.n553 gnd 0.009097f
C1315 vdd.n554 gnd 0.009097f
C1316 vdd.n555 gnd 0.009097f
C1317 vdd.n556 gnd 0.007248f
C1318 vdd.t83 gnd 0.111913f
C1319 vdd.t84 gnd 0.119604f
C1320 vdd.t81 gnd 0.146157f
C1321 vdd.n557 gnd 0.187352f
C1322 vdd.n558 gnd 0.15741f
C1323 vdd.n559 gnd 0.009097f
C1324 vdd.n560 gnd 0.009097f
C1325 vdd.n561 gnd 0.009097f
C1326 vdd.n562 gnd 0.009097f
C1327 vdd.n563 gnd 0.009097f
C1328 vdd.n564 gnd 0.009097f
C1329 vdd.n565 gnd 0.009097f
C1330 vdd.n566 gnd 0.009097f
C1331 vdd.n567 gnd 0.009097f
C1332 vdd.n568 gnd 0.009097f
C1333 vdd.n569 gnd 0.009097f
C1334 vdd.n570 gnd 0.009097f
C1335 vdd.n571 gnd 0.009097f
C1336 vdd.n572 gnd 0.005822f
C1337 vdd.n575 gnd 0.006186f
C1338 vdd.n576 gnd 0.006186f
C1339 vdd.n577 gnd 0.006186f
C1340 vdd.n578 gnd 0.006186f
C1341 vdd.n579 gnd 0.006186f
C1342 vdd.n580 gnd 0.006186f
C1343 vdd.n582 gnd 0.006186f
C1344 vdd.n583 gnd 0.006186f
C1345 vdd.n585 gnd 0.006186f
C1346 vdd.n586 gnd 0.004503f
C1347 vdd.n588 gnd 0.006186f
C1348 vdd.t127 gnd 0.249964f
C1349 vdd.t126 gnd 0.255869f
C1350 vdd.t125 gnd 0.163186f
C1351 vdd.n589 gnd 0.088193f
C1352 vdd.n590 gnd 0.050026f
C1353 vdd.n591 gnd 0.00884f
C1354 vdd.n592 gnd 0.014457f
C1355 vdd.n594 gnd 0.006186f
C1356 vdd.n595 gnd 0.632151f
C1357 vdd.n596 gnd 0.013704f
C1358 vdd.n597 gnd 0.013704f
C1359 vdd.n598 gnd 0.006186f
C1360 vdd.n599 gnd 0.014678f
C1361 vdd.n600 gnd 0.006186f
C1362 vdd.n601 gnd 0.006186f
C1363 vdd.n602 gnd 0.006186f
C1364 vdd.n603 gnd 0.006186f
C1365 vdd.n604 gnd 0.006186f
C1366 vdd.n606 gnd 0.006186f
C1367 vdd.n607 gnd 0.006186f
C1368 vdd.n609 gnd 0.006186f
C1369 vdd.n610 gnd 0.006186f
C1370 vdd.n612 gnd 0.006186f
C1371 vdd.n613 gnd 0.006186f
C1372 vdd.n615 gnd 0.006186f
C1373 vdd.n616 gnd 0.006186f
C1374 vdd.n618 gnd 0.006186f
C1375 vdd.n619 gnd 0.006186f
C1376 vdd.n621 gnd 0.006186f
C1377 vdd.t120 gnd 0.249964f
C1378 vdd.t119 gnd 0.255869f
C1379 vdd.t117 gnd 0.163186f
C1380 vdd.n622 gnd 0.088193f
C1381 vdd.n623 gnd 0.050026f
C1382 vdd.n624 gnd 0.006186f
C1383 vdd.n626 gnd 0.006186f
C1384 vdd.n627 gnd 0.006186f
C1385 vdd.t118 gnd 0.316076f
C1386 vdd.n628 gnd 0.006186f
C1387 vdd.n629 gnd 0.006186f
C1388 vdd.n630 gnd 0.006186f
C1389 vdd.n631 gnd 0.006186f
C1390 vdd.n632 gnd 0.006186f
C1391 vdd.n633 gnd 0.632151f
C1392 vdd.n634 gnd 0.006186f
C1393 vdd.n635 gnd 0.006186f
C1394 vdd.n636 gnd 0.553133f
C1395 vdd.n637 gnd 0.006186f
C1396 vdd.n638 gnd 0.006186f
C1397 vdd.n639 gnd 0.005458f
C1398 vdd.n640 gnd 0.006186f
C1399 vdd.n641 gnd 0.557781f
C1400 vdd.n642 gnd 0.006186f
C1401 vdd.n643 gnd 0.006186f
C1402 vdd.n644 gnd 0.006186f
C1403 vdd.n645 gnd 0.006186f
C1404 vdd.n646 gnd 0.006186f
C1405 vdd.n647 gnd 0.632151f
C1406 vdd.n648 gnd 0.006186f
C1407 vdd.n649 gnd 0.006186f
C1408 vdd.t97 gnd 0.283539f
C1409 vdd.t188 gnd 0.074371f
C1410 vdd.n650 gnd 0.006186f
C1411 vdd.n651 gnd 0.006186f
C1412 vdd.n652 gnd 0.006186f
C1413 vdd.t173 gnd 0.316076f
C1414 vdd.n653 gnd 0.006186f
C1415 vdd.n654 gnd 0.006186f
C1416 vdd.n655 gnd 0.006186f
C1417 vdd.n656 gnd 0.006186f
C1418 vdd.n657 gnd 0.006186f
C1419 vdd.t178 gnd 0.316076f
C1420 vdd.n658 gnd 0.006186f
C1421 vdd.n659 gnd 0.006186f
C1422 vdd.n660 gnd 0.525243f
C1423 vdd.n661 gnd 0.006186f
C1424 vdd.n662 gnd 0.006186f
C1425 vdd.n663 gnd 0.006186f
C1426 vdd.n664 gnd 0.385798f
C1427 vdd.n665 gnd 0.006186f
C1428 vdd.n666 gnd 0.006186f
C1429 vdd.t0 gnd 0.316076f
C1430 vdd.n667 gnd 0.006186f
C1431 vdd.n668 gnd 0.006186f
C1432 vdd.n669 gnd 0.006186f
C1433 vdd.n670 gnd 0.525243f
C1434 vdd.n671 gnd 0.006186f
C1435 vdd.n672 gnd 0.006186f
C1436 vdd.t77 gnd 0.269594f
C1437 vdd.t194 gnd 0.246353f
C1438 vdd.n673 gnd 0.006186f
C1439 vdd.n674 gnd 0.006186f
C1440 vdd.n675 gnd 0.006186f
C1441 vdd.t179 gnd 0.316076f
C1442 vdd.n676 gnd 0.006186f
C1443 vdd.n677 gnd 0.006186f
C1444 vdd.t6 gnd 0.316076f
C1445 vdd.n678 gnd 0.006186f
C1446 vdd.n679 gnd 0.006186f
C1447 vdd.n680 gnd 0.006186f
C1448 vdd.t78 gnd 0.232409f
C1449 vdd.n681 gnd 0.006186f
C1450 vdd.n682 gnd 0.006186f
C1451 vdd.n683 gnd 0.539188f
C1452 vdd.n684 gnd 0.006186f
C1453 vdd.n685 gnd 0.006186f
C1454 vdd.n686 gnd 0.006186f
C1455 vdd.n687 gnd 0.632151f
C1456 vdd.n688 gnd 0.006186f
C1457 vdd.n689 gnd 0.006186f
C1458 vdd.t189 gnd 0.283539f
C1459 vdd.n690 gnd 0.399743f
C1460 vdd.n691 gnd 0.006186f
C1461 vdd.n692 gnd 0.006186f
C1462 vdd.n693 gnd 0.006186f
C1463 vdd.t7 gnd 0.316076f
C1464 vdd.n694 gnd 0.006186f
C1465 vdd.n695 gnd 0.006186f
C1466 vdd.n696 gnd 0.006186f
C1467 vdd.n697 gnd 0.006186f
C1468 vdd.n698 gnd 0.006186f
C1469 vdd.t198 gnd 0.632151f
C1470 vdd.n699 gnd 0.006186f
C1471 vdd.n700 gnd 0.006186f
C1472 vdd.t122 gnd 0.316076f
C1473 vdd.n701 gnd 0.006186f
C1474 vdd.n702 gnd 0.014678f
C1475 vdd.n703 gnd 0.014678f
C1476 vdd.t196 gnd 0.594966f
C1477 vdd.n704 gnd 0.013704f
C1478 vdd.n705 gnd 0.013704f
C1479 vdd.n706 gnd 0.014678f
C1480 vdd.n707 gnd 0.006186f
C1481 vdd.n708 gnd 0.006186f
C1482 vdd.t4 gnd 0.594966f
C1483 vdd.n726 gnd 0.014678f
C1484 vdd.n744 gnd 0.013704f
C1485 vdd.n745 gnd 0.006186f
C1486 vdd.n746 gnd 0.013704f
C1487 vdd.t147 gnd 0.249964f
C1488 vdd.t146 gnd 0.255869f
C1489 vdd.t145 gnd 0.163186f
C1490 vdd.n747 gnd 0.088193f
C1491 vdd.n748 gnd 0.050026f
C1492 vdd.n749 gnd 0.014457f
C1493 vdd.n750 gnd 0.006186f
C1494 vdd.t2 gnd 0.632151f
C1495 vdd.n751 gnd 0.013704f
C1496 vdd.n752 gnd 0.006186f
C1497 vdd.n753 gnd 0.014678f
C1498 vdd.n754 gnd 0.006186f
C1499 vdd.t116 gnd 0.249964f
C1500 vdd.t115 gnd 0.255869f
C1501 vdd.t113 gnd 0.163186f
C1502 vdd.n755 gnd 0.088193f
C1503 vdd.n756 gnd 0.050026f
C1504 vdd.n757 gnd 0.00884f
C1505 vdd.n758 gnd 0.006186f
C1506 vdd.n759 gnd 0.006186f
C1507 vdd.t114 gnd 0.316076f
C1508 vdd.n760 gnd 0.006186f
C1509 vdd.n761 gnd 0.006186f
C1510 vdd.n762 gnd 0.006186f
C1511 vdd.n763 gnd 0.006186f
C1512 vdd.n764 gnd 0.006186f
C1513 vdd.n765 gnd 0.006186f
C1514 vdd.n766 gnd 0.632151f
C1515 vdd.n767 gnd 0.006186f
C1516 vdd.n768 gnd 0.006186f
C1517 vdd.t74 gnd 0.316076f
C1518 vdd.n769 gnd 0.006186f
C1519 vdd.n770 gnd 0.006186f
C1520 vdd.n771 gnd 0.006186f
C1521 vdd.n772 gnd 0.006186f
C1522 vdd.n773 gnd 0.399743f
C1523 vdd.n774 gnd 0.006186f
C1524 vdd.n775 gnd 0.006186f
C1525 vdd.n776 gnd 0.006186f
C1526 vdd.n777 gnd 0.006186f
C1527 vdd.n778 gnd 0.006186f
C1528 vdd.n779 gnd 0.539188f
C1529 vdd.n780 gnd 0.006186f
C1530 vdd.n781 gnd 0.006186f
C1531 vdd.t186 gnd 0.283539f
C1532 vdd.t191 gnd 0.232409f
C1533 vdd.n782 gnd 0.006186f
C1534 vdd.n783 gnd 0.006186f
C1535 vdd.n784 gnd 0.006186f
C1536 vdd.t9 gnd 0.316076f
C1537 vdd.n785 gnd 0.006186f
C1538 vdd.n786 gnd 0.006186f
C1539 vdd.t183 gnd 0.316076f
C1540 vdd.n787 gnd 0.006186f
C1541 vdd.n788 gnd 0.006186f
C1542 vdd.n789 gnd 0.006186f
C1543 vdd.t176 gnd 0.246353f
C1544 vdd.n790 gnd 0.006186f
C1545 vdd.n791 gnd 0.006186f
C1546 vdd.n792 gnd 0.525243f
C1547 vdd.n793 gnd 0.006186f
C1548 vdd.n794 gnd 0.006186f
C1549 vdd.n795 gnd 0.006186f
C1550 vdd.t192 gnd 0.316076f
C1551 vdd.n796 gnd 0.006186f
C1552 vdd.n797 gnd 0.006186f
C1553 vdd.t76 gnd 0.269594f
C1554 vdd.n798 gnd 0.385798f
C1555 vdd.n799 gnd 0.006186f
C1556 vdd.n800 gnd 0.006186f
C1557 vdd.n801 gnd 0.006186f
C1558 vdd.n802 gnd 0.525243f
C1559 vdd.n803 gnd 0.006186f
C1560 vdd.n804 gnd 0.006186f
C1561 vdd.t185 gnd 0.316076f
C1562 vdd.n805 gnd 0.006186f
C1563 vdd.n806 gnd 0.006186f
C1564 vdd.n807 gnd 0.006186f
C1565 vdd.n808 gnd 0.632151f
C1566 vdd.n809 gnd 0.006186f
C1567 vdd.n810 gnd 0.006186f
C1568 vdd.t175 gnd 0.316076f
C1569 vdd.n811 gnd 0.006186f
C1570 vdd.n812 gnd 0.006186f
C1571 vdd.n813 gnd 0.006186f
C1572 vdd.t174 gnd 0.074371f
C1573 vdd.n814 gnd 0.006186f
C1574 vdd.n815 gnd 0.006186f
C1575 vdd.n816 gnd 0.006186f
C1576 vdd.t134 gnd 0.255869f
C1577 vdd.t132 gnd 0.163186f
C1578 vdd.t135 gnd 0.255869f
C1579 vdd.n817 gnd 0.143809f
C1580 vdd.n818 gnd 0.006186f
C1581 vdd.n819 gnd 0.006186f
C1582 vdd.n820 gnd 0.632151f
C1583 vdd.n821 gnd 0.006186f
C1584 vdd.n822 gnd 0.006186f
C1585 vdd.t133 gnd 0.283539f
C1586 vdd.n823 gnd 0.557781f
C1587 vdd.n824 gnd 0.006186f
C1588 vdd.n825 gnd 0.006186f
C1589 vdd.n826 gnd 0.006186f
C1590 vdd.n827 gnd 0.553133f
C1591 vdd.n828 gnd 0.006186f
C1592 vdd.n829 gnd 0.006186f
C1593 vdd.n830 gnd 0.006186f
C1594 vdd.n831 gnd 0.006186f
C1595 vdd.n832 gnd 0.006186f
C1596 vdd.n833 gnd 0.632151f
C1597 vdd.n834 gnd 0.006186f
C1598 vdd.n835 gnd 0.006186f
C1599 vdd.t129 gnd 0.316076f
C1600 vdd.n836 gnd 0.006186f
C1601 vdd.n837 gnd 0.014678f
C1602 vdd.n838 gnd 0.014678f
C1603 vdd.n839 gnd 6.40518f
C1604 vdd.n840 gnd 0.013704f
C1605 vdd.n841 gnd 0.013704f
C1606 vdd.n842 gnd 0.014678f
C1607 vdd.n843 gnd 0.006186f
C1608 vdd.n844 gnd 0.006186f
C1609 vdd.n845 gnd 0.006186f
C1610 vdd.n846 gnd 0.006186f
C1611 vdd.n847 gnd 0.006186f
C1612 vdd.n848 gnd 0.006186f
C1613 vdd.n849 gnd 0.006186f
C1614 vdd.n850 gnd 0.006186f
C1615 vdd.n852 gnd 0.006186f
C1616 vdd.n853 gnd 0.006186f
C1617 vdd.n854 gnd 0.005822f
C1618 vdd.n857 gnd 0.022678f
C1619 vdd.n858 gnd 0.007322f
C1620 vdd.n859 gnd 0.009097f
C1621 vdd.n861 gnd 0.009097f
C1622 vdd.n862 gnd 0.006077f
C1623 vdd.t89 gnd 0.464817f
C1624 vdd.n863 gnd 6.73985f
C1625 vdd.n864 gnd 0.009097f
C1626 vdd.n865 gnd 0.022678f
C1627 vdd.n866 gnd 0.007322f
C1628 vdd.n867 gnd 0.009097f
C1629 vdd.n868 gnd 0.007322f
C1630 vdd.n869 gnd 0.009097f
C1631 vdd.n870 gnd 0.929634f
C1632 vdd.n871 gnd 0.009097f
C1633 vdd.n872 gnd 0.007322f
C1634 vdd.n873 gnd 0.007322f
C1635 vdd.n874 gnd 0.009097f
C1636 vdd.n875 gnd 0.007322f
C1637 vdd.n876 gnd 0.009097f
C1638 vdd.t10 gnd 0.464817f
C1639 vdd.n877 gnd 0.009097f
C1640 vdd.n878 gnd 0.007322f
C1641 vdd.n879 gnd 0.009097f
C1642 vdd.n880 gnd 0.007322f
C1643 vdd.n881 gnd 0.009097f
C1644 vdd.t63 gnd 0.464817f
C1645 vdd.n882 gnd 0.009097f
C1646 vdd.n883 gnd 0.007322f
C1647 vdd.n884 gnd 0.009097f
C1648 vdd.n885 gnd 0.007322f
C1649 vdd.n886 gnd 0.009097f
C1650 vdd.n887 gnd 0.729763f
C1651 vdd.n888 gnd 0.771597f
C1652 vdd.t18 gnd 0.464817f
C1653 vdd.n889 gnd 0.009097f
C1654 vdd.n890 gnd 0.007322f
C1655 vdd.n891 gnd 0.004992f
C1656 vdd.n892 gnd 0.004633f
C1657 vdd.n893 gnd 0.002563f
C1658 vdd.n894 gnd 0.005884f
C1659 vdd.n895 gnd 0.002489f
C1660 vdd.n896 gnd 0.002636f
C1661 vdd.n897 gnd 0.004633f
C1662 vdd.n898 gnd 0.002489f
C1663 vdd.n899 gnd 0.005884f
C1664 vdd.n900 gnd 0.002636f
C1665 vdd.n901 gnd 0.004633f
C1666 vdd.n902 gnd 0.002489f
C1667 vdd.n903 gnd 0.004413f
C1668 vdd.n904 gnd 0.004426f
C1669 vdd.t11 gnd 0.012641f
C1670 vdd.n905 gnd 0.028127f
C1671 vdd.n906 gnd 0.146377f
C1672 vdd.n907 gnd 0.002489f
C1673 vdd.n908 gnd 0.002636f
C1674 vdd.n909 gnd 0.005884f
C1675 vdd.n910 gnd 0.005884f
C1676 vdd.n911 gnd 0.002636f
C1677 vdd.n912 gnd 0.002489f
C1678 vdd.n913 gnd 0.004633f
C1679 vdd.n914 gnd 0.004633f
C1680 vdd.n915 gnd 0.002489f
C1681 vdd.n916 gnd 0.002636f
C1682 vdd.n917 gnd 0.005884f
C1683 vdd.n918 gnd 0.005884f
C1684 vdd.n919 gnd 0.002636f
C1685 vdd.n920 gnd 0.002489f
C1686 vdd.n921 gnd 0.004633f
C1687 vdd.n922 gnd 0.004633f
C1688 vdd.n923 gnd 0.002489f
C1689 vdd.n924 gnd 0.002636f
C1690 vdd.n925 gnd 0.005884f
C1691 vdd.n926 gnd 0.005884f
C1692 vdd.n927 gnd 0.013911f
C1693 vdd.n928 gnd 0.002563f
C1694 vdd.n929 gnd 0.002489f
C1695 vdd.n930 gnd 0.011974f
C1696 vdd.n931 gnd 0.008359f
C1697 vdd.t37 gnd 0.029287f
C1698 vdd.t66 gnd 0.029287f
C1699 vdd.n932 gnd 0.201279f
C1700 vdd.n933 gnd 0.158275f
C1701 vdd.t26 gnd 0.029287f
C1702 vdd.t54 gnd 0.029287f
C1703 vdd.n934 gnd 0.201279f
C1704 vdd.n935 gnd 0.127727f
C1705 vdd.t32 gnd 0.029287f
C1706 vdd.t60 gnd 0.029287f
C1707 vdd.n936 gnd 0.201279f
C1708 vdd.n937 gnd 0.127727f
C1709 vdd.n938 gnd 0.004992f
C1710 vdd.n939 gnd 0.004633f
C1711 vdd.n940 gnd 0.002563f
C1712 vdd.n941 gnd 0.005884f
C1713 vdd.n942 gnd 0.002489f
C1714 vdd.n943 gnd 0.002636f
C1715 vdd.n944 gnd 0.004633f
C1716 vdd.n945 gnd 0.002489f
C1717 vdd.n946 gnd 0.005884f
C1718 vdd.n947 gnd 0.002636f
C1719 vdd.n948 gnd 0.004633f
C1720 vdd.n949 gnd 0.002489f
C1721 vdd.n950 gnd 0.004413f
C1722 vdd.n951 gnd 0.004426f
C1723 vdd.t70 gnd 0.012641f
C1724 vdd.n952 gnd 0.028127f
C1725 vdd.n953 gnd 0.146377f
C1726 vdd.n954 gnd 0.002489f
C1727 vdd.n955 gnd 0.002636f
C1728 vdd.n956 gnd 0.005884f
C1729 vdd.n957 gnd 0.005884f
C1730 vdd.n958 gnd 0.002636f
C1731 vdd.n959 gnd 0.002489f
C1732 vdd.n960 gnd 0.004633f
C1733 vdd.n961 gnd 0.004633f
C1734 vdd.n962 gnd 0.002489f
C1735 vdd.n963 gnd 0.002636f
C1736 vdd.n964 gnd 0.005884f
C1737 vdd.n965 gnd 0.005884f
C1738 vdd.n966 gnd 0.002636f
C1739 vdd.n967 gnd 0.002489f
C1740 vdd.n968 gnd 0.004633f
C1741 vdd.n969 gnd 0.004633f
C1742 vdd.n970 gnd 0.002489f
C1743 vdd.n971 gnd 0.002636f
C1744 vdd.n972 gnd 0.005884f
C1745 vdd.n973 gnd 0.005884f
C1746 vdd.n974 gnd 0.013911f
C1747 vdd.n975 gnd 0.002563f
C1748 vdd.n976 gnd 0.002489f
C1749 vdd.n977 gnd 0.011974f
C1750 vdd.n978 gnd 0.008097f
C1751 vdd.n979 gnd 0.09503f
C1752 vdd.n980 gnd 0.004992f
C1753 vdd.n981 gnd 0.004633f
C1754 vdd.n982 gnd 0.002563f
C1755 vdd.n983 gnd 0.005884f
C1756 vdd.n984 gnd 0.002489f
C1757 vdd.n985 gnd 0.002636f
C1758 vdd.n986 gnd 0.004633f
C1759 vdd.n987 gnd 0.002489f
C1760 vdd.n988 gnd 0.005884f
C1761 vdd.n989 gnd 0.002636f
C1762 vdd.n990 gnd 0.004633f
C1763 vdd.n991 gnd 0.002489f
C1764 vdd.n992 gnd 0.004413f
C1765 vdd.n993 gnd 0.004426f
C1766 vdd.t61 gnd 0.012641f
C1767 vdd.n994 gnd 0.028127f
C1768 vdd.n995 gnd 0.146377f
C1769 vdd.n996 gnd 0.002489f
C1770 vdd.n997 gnd 0.002636f
C1771 vdd.n998 gnd 0.005884f
C1772 vdd.n999 gnd 0.005884f
C1773 vdd.n1000 gnd 0.002636f
C1774 vdd.n1001 gnd 0.002489f
C1775 vdd.n1002 gnd 0.004633f
C1776 vdd.n1003 gnd 0.004633f
C1777 vdd.n1004 gnd 0.002489f
C1778 vdd.n1005 gnd 0.002636f
C1779 vdd.n1006 gnd 0.005884f
C1780 vdd.n1007 gnd 0.005884f
C1781 vdd.n1008 gnd 0.002636f
C1782 vdd.n1009 gnd 0.002489f
C1783 vdd.n1010 gnd 0.004633f
C1784 vdd.n1011 gnd 0.004633f
C1785 vdd.n1012 gnd 0.002489f
C1786 vdd.n1013 gnd 0.002636f
C1787 vdd.n1014 gnd 0.005884f
C1788 vdd.n1015 gnd 0.005884f
C1789 vdd.n1016 gnd 0.013911f
C1790 vdd.n1017 gnd 0.002563f
C1791 vdd.n1018 gnd 0.002489f
C1792 vdd.n1019 gnd 0.011974f
C1793 vdd.n1020 gnd 0.008359f
C1794 vdd.t19 gnd 0.029287f
C1795 vdd.t64 gnd 0.029287f
C1796 vdd.n1021 gnd 0.201279f
C1797 vdd.n1022 gnd 0.158275f
C1798 vdd.t59 gnd 0.029287f
C1799 vdd.t50 gnd 0.029287f
C1800 vdd.n1023 gnd 0.201279f
C1801 vdd.n1024 gnd 0.127727f
C1802 vdd.t35 gnd 0.029287f
C1803 vdd.t15 gnd 0.029287f
C1804 vdd.n1025 gnd 0.201279f
C1805 vdd.n1026 gnd 0.127727f
C1806 vdd.n1027 gnd 0.004992f
C1807 vdd.n1028 gnd 0.004633f
C1808 vdd.n1029 gnd 0.002563f
C1809 vdd.n1030 gnd 0.005884f
C1810 vdd.n1031 gnd 0.002489f
C1811 vdd.n1032 gnd 0.002636f
C1812 vdd.n1033 gnd 0.004633f
C1813 vdd.n1034 gnd 0.002489f
C1814 vdd.n1035 gnd 0.005884f
C1815 vdd.n1036 gnd 0.002636f
C1816 vdd.n1037 gnd 0.004633f
C1817 vdd.n1038 gnd 0.002489f
C1818 vdd.n1039 gnd 0.004413f
C1819 vdd.n1040 gnd 0.004426f
C1820 vdd.t48 gnd 0.012641f
C1821 vdd.n1041 gnd 0.028127f
C1822 vdd.n1042 gnd 0.146377f
C1823 vdd.n1043 gnd 0.002489f
C1824 vdd.n1044 gnd 0.002636f
C1825 vdd.n1045 gnd 0.005884f
C1826 vdd.n1046 gnd 0.005884f
C1827 vdd.n1047 gnd 0.002636f
C1828 vdd.n1048 gnd 0.002489f
C1829 vdd.n1049 gnd 0.004633f
C1830 vdd.n1050 gnd 0.004633f
C1831 vdd.n1051 gnd 0.002489f
C1832 vdd.n1052 gnd 0.002636f
C1833 vdd.n1053 gnd 0.005884f
C1834 vdd.n1054 gnd 0.005884f
C1835 vdd.n1055 gnd 0.002636f
C1836 vdd.n1056 gnd 0.002489f
C1837 vdd.n1057 gnd 0.004633f
C1838 vdd.n1058 gnd 0.004633f
C1839 vdd.n1059 gnd 0.002489f
C1840 vdd.n1060 gnd 0.002636f
C1841 vdd.n1061 gnd 0.005884f
C1842 vdd.n1062 gnd 0.005884f
C1843 vdd.n1063 gnd 0.013911f
C1844 vdd.n1064 gnd 0.002563f
C1845 vdd.n1065 gnd 0.002489f
C1846 vdd.n1066 gnd 0.011974f
C1847 vdd.n1067 gnd 0.008097f
C1848 vdd.n1068 gnd 0.056533f
C1849 vdd.n1069 gnd 0.203704f
C1850 vdd.n1070 gnd 0.004992f
C1851 vdd.n1071 gnd 0.004633f
C1852 vdd.n1072 gnd 0.002563f
C1853 vdd.n1073 gnd 0.005884f
C1854 vdd.n1074 gnd 0.002489f
C1855 vdd.n1075 gnd 0.002636f
C1856 vdd.n1076 gnd 0.004633f
C1857 vdd.n1077 gnd 0.002489f
C1858 vdd.n1078 gnd 0.005884f
C1859 vdd.n1079 gnd 0.002636f
C1860 vdd.n1080 gnd 0.004633f
C1861 vdd.n1081 gnd 0.002489f
C1862 vdd.n1082 gnd 0.004413f
C1863 vdd.n1083 gnd 0.004426f
C1864 vdd.t69 gnd 0.012641f
C1865 vdd.n1084 gnd 0.028127f
C1866 vdd.n1085 gnd 0.146377f
C1867 vdd.n1086 gnd 0.002489f
C1868 vdd.n1087 gnd 0.002636f
C1869 vdd.n1088 gnd 0.005884f
C1870 vdd.n1089 gnd 0.005884f
C1871 vdd.n1090 gnd 0.002636f
C1872 vdd.n1091 gnd 0.002489f
C1873 vdd.n1092 gnd 0.004633f
C1874 vdd.n1093 gnd 0.004633f
C1875 vdd.n1094 gnd 0.002489f
C1876 vdd.n1095 gnd 0.002636f
C1877 vdd.n1096 gnd 0.005884f
C1878 vdd.n1097 gnd 0.005884f
C1879 vdd.n1098 gnd 0.002636f
C1880 vdd.n1099 gnd 0.002489f
C1881 vdd.n1100 gnd 0.004633f
C1882 vdd.n1101 gnd 0.004633f
C1883 vdd.n1102 gnd 0.002489f
C1884 vdd.n1103 gnd 0.002636f
C1885 vdd.n1104 gnd 0.005884f
C1886 vdd.n1105 gnd 0.005884f
C1887 vdd.n1106 gnd 0.013911f
C1888 vdd.n1107 gnd 0.002563f
C1889 vdd.n1108 gnd 0.002489f
C1890 vdd.n1109 gnd 0.011974f
C1891 vdd.n1110 gnd 0.008359f
C1892 vdd.t24 gnd 0.029287f
C1893 vdd.t68 gnd 0.029287f
C1894 vdd.n1111 gnd 0.201279f
C1895 vdd.n1112 gnd 0.158275f
C1896 vdd.t67 gnd 0.029287f
C1897 vdd.t56 gnd 0.029287f
C1898 vdd.n1113 gnd 0.201279f
C1899 vdd.n1114 gnd 0.127727f
C1900 vdd.t43 gnd 0.029287f
C1901 vdd.t22 gnd 0.029287f
C1902 vdd.n1115 gnd 0.201279f
C1903 vdd.n1116 gnd 0.127727f
C1904 vdd.n1117 gnd 0.004992f
C1905 vdd.n1118 gnd 0.004633f
C1906 vdd.n1119 gnd 0.002563f
C1907 vdd.n1120 gnd 0.005884f
C1908 vdd.n1121 gnd 0.002489f
C1909 vdd.n1122 gnd 0.002636f
C1910 vdd.n1123 gnd 0.004633f
C1911 vdd.n1124 gnd 0.002489f
C1912 vdd.n1125 gnd 0.005884f
C1913 vdd.n1126 gnd 0.002636f
C1914 vdd.n1127 gnd 0.004633f
C1915 vdd.n1128 gnd 0.002489f
C1916 vdd.n1129 gnd 0.004413f
C1917 vdd.n1130 gnd 0.004426f
C1918 vdd.t55 gnd 0.012641f
C1919 vdd.n1131 gnd 0.028127f
C1920 vdd.n1132 gnd 0.146377f
C1921 vdd.n1133 gnd 0.002489f
C1922 vdd.n1134 gnd 0.002636f
C1923 vdd.n1135 gnd 0.005884f
C1924 vdd.n1136 gnd 0.005884f
C1925 vdd.n1137 gnd 0.002636f
C1926 vdd.n1138 gnd 0.002489f
C1927 vdd.n1139 gnd 0.004633f
C1928 vdd.n1140 gnd 0.004633f
C1929 vdd.n1141 gnd 0.002489f
C1930 vdd.n1142 gnd 0.002636f
C1931 vdd.n1143 gnd 0.005884f
C1932 vdd.n1144 gnd 0.005884f
C1933 vdd.n1145 gnd 0.002636f
C1934 vdd.n1146 gnd 0.002489f
C1935 vdd.n1147 gnd 0.004633f
C1936 vdd.n1148 gnd 0.004633f
C1937 vdd.n1149 gnd 0.002489f
C1938 vdd.n1150 gnd 0.002636f
C1939 vdd.n1151 gnd 0.005884f
C1940 vdd.n1152 gnd 0.005884f
C1941 vdd.n1153 gnd 0.013911f
C1942 vdd.n1154 gnd 0.002563f
C1943 vdd.n1155 gnd 0.002489f
C1944 vdd.n1156 gnd 0.011974f
C1945 vdd.n1157 gnd 0.008097f
C1946 vdd.n1158 gnd 0.056533f
C1947 vdd.n1159 gnd 0.220485f
C1948 vdd.n1160 gnd 1.85301f
C1949 vdd.n1161 gnd 0.536555f
C1950 vdd.n1162 gnd 0.007322f
C1951 vdd.n1163 gnd 0.009097f
C1952 vdd.n1164 gnd 0.571725f
C1953 vdd.n1165 gnd 0.009097f
C1954 vdd.n1166 gnd 0.007322f
C1955 vdd.n1167 gnd 0.009097f
C1956 vdd.n1168 gnd 0.007322f
C1957 vdd.n1169 gnd 0.009097f
C1958 vdd.t14 gnd 0.464817f
C1959 vdd.t25 gnd 0.464817f
C1960 vdd.n1170 gnd 0.009097f
C1961 vdd.n1171 gnd 0.007322f
C1962 vdd.n1172 gnd 0.009097f
C1963 vdd.n1173 gnd 0.007322f
C1964 vdd.n1174 gnd 0.009097f
C1965 vdd.t31 gnd 0.464817f
C1966 vdd.n1175 gnd 0.009097f
C1967 vdd.n1176 gnd 0.007322f
C1968 vdd.n1177 gnd 0.009097f
C1969 vdd.n1178 gnd 0.007322f
C1970 vdd.n1179 gnd 0.009097f
C1971 vdd.t47 gnd 0.464817f
C1972 vdd.n1180 gnd 0.673985f
C1973 vdd.n1181 gnd 0.009097f
C1974 vdd.n1182 gnd 0.007322f
C1975 vdd.n1183 gnd 0.009097f
C1976 vdd.n1184 gnd 0.007322f
C1977 vdd.n1185 gnd 0.009097f
C1978 vdd.n1186 gnd 0.929634f
C1979 vdd.n1187 gnd 0.009097f
C1980 vdd.n1188 gnd 0.007322f
C1981 vdd.n1189 gnd 0.022169f
C1982 vdd.n1190 gnd 0.006077f
C1983 vdd.n1191 gnd 0.022169f
C1984 vdd.t93 gnd 0.464817f
C1985 vdd.n1192 gnd 0.022169f
C1986 vdd.n1193 gnd 0.006077f
C1987 vdd.n1194 gnd 0.009097f
C1988 vdd.n1195 gnd 0.007322f
C1989 vdd.n1196 gnd 0.009097f
C1990 vdd.n1227 gnd 0.022678f
C1991 vdd.n1228 gnd 1.37121f
C1992 vdd.n1229 gnd 0.009097f
C1993 vdd.n1230 gnd 0.007322f
C1994 vdd.n1231 gnd 0.009097f
C1995 vdd.n1232 gnd 0.009097f
C1996 vdd.n1233 gnd 0.009097f
C1997 vdd.n1234 gnd 0.009097f
C1998 vdd.n1235 gnd 0.009097f
C1999 vdd.n1236 gnd 0.007322f
C2000 vdd.n1237 gnd 0.009097f
C2001 vdd.n1238 gnd 0.009097f
C2002 vdd.n1239 gnd 0.009097f
C2003 vdd.n1240 gnd 0.009097f
C2004 vdd.n1241 gnd 0.009097f
C2005 vdd.n1242 gnd 0.007322f
C2006 vdd.n1243 gnd 0.009097f
C2007 vdd.n1244 gnd 0.009097f
C2008 vdd.n1245 gnd 0.009097f
C2009 vdd.n1246 gnd 0.009097f
C2010 vdd.n1247 gnd 0.009097f
C2011 vdd.n1248 gnd 0.007322f
C2012 vdd.n1249 gnd 0.009097f
C2013 vdd.n1250 gnd 0.009097f
C2014 vdd.n1251 gnd 0.009097f
C2015 vdd.n1252 gnd 0.009097f
C2016 vdd.n1253 gnd 0.009097f
C2017 vdd.t143 gnd 0.111913f
C2018 vdd.t144 gnd 0.119604f
C2019 vdd.t142 gnd 0.146157f
C2020 vdd.n1254 gnd 0.187352f
C2021 vdd.n1255 gnd 0.158142f
C2022 vdd.n1256 gnd 0.015668f
C2023 vdd.n1257 gnd 0.009097f
C2024 vdd.n1258 gnd 0.009097f
C2025 vdd.n1259 gnd 0.009097f
C2026 vdd.n1260 gnd 0.009097f
C2027 vdd.n1261 gnd 0.009097f
C2028 vdd.n1262 gnd 0.007322f
C2029 vdd.n1263 gnd 0.009097f
C2030 vdd.n1264 gnd 0.009097f
C2031 vdd.n1265 gnd 0.009097f
C2032 vdd.n1266 gnd 0.009097f
C2033 vdd.n1267 gnd 0.009097f
C2034 vdd.n1268 gnd 0.007322f
C2035 vdd.n1269 gnd 0.009097f
C2036 vdd.n1270 gnd 0.009097f
C2037 vdd.n1271 gnd 0.009097f
C2038 vdd.n1272 gnd 0.009097f
C2039 vdd.n1273 gnd 0.009097f
C2040 vdd.n1274 gnd 0.007322f
C2041 vdd.n1275 gnd 0.009097f
C2042 vdd.n1276 gnd 0.009097f
C2043 vdd.n1277 gnd 0.009097f
C2044 vdd.n1278 gnd 0.009097f
C2045 vdd.n1279 gnd 0.009097f
C2046 vdd.n1280 gnd 0.007322f
C2047 vdd.n1281 gnd 0.009097f
C2048 vdd.n1282 gnd 0.009097f
C2049 vdd.n1283 gnd 0.009097f
C2050 vdd.n1284 gnd 0.009097f
C2051 vdd.n1285 gnd 0.009097f
C2052 vdd.n1286 gnd 0.007322f
C2053 vdd.n1287 gnd 0.009097f
C2054 vdd.n1288 gnd 0.009097f
C2055 vdd.n1289 gnd 0.009097f
C2056 vdd.n1290 gnd 0.009097f
C2057 vdd.n1291 gnd 0.007322f
C2058 vdd.n1292 gnd 0.009097f
C2059 vdd.n1293 gnd 0.009097f
C2060 vdd.n1294 gnd 0.009097f
C2061 vdd.n1295 gnd 0.009097f
C2062 vdd.n1296 gnd 0.009097f
C2063 vdd.n1297 gnd 0.007322f
C2064 vdd.n1298 gnd 0.009097f
C2065 vdd.n1299 gnd 0.009097f
C2066 vdd.n1300 gnd 0.009097f
C2067 vdd.n1301 gnd 0.009097f
C2068 vdd.n1302 gnd 0.009097f
C2069 vdd.n1303 gnd 0.007322f
C2070 vdd.n1304 gnd 0.009097f
C2071 vdd.n1305 gnd 0.009097f
C2072 vdd.n1306 gnd 0.009097f
C2073 vdd.n1307 gnd 0.009097f
C2074 vdd.n1308 gnd 0.009097f
C2075 vdd.n1309 gnd 0.007322f
C2076 vdd.n1310 gnd 0.009097f
C2077 vdd.n1311 gnd 0.009097f
C2078 vdd.n1312 gnd 0.009097f
C2079 vdd.n1313 gnd 0.009097f
C2080 vdd.n1314 gnd 0.009097f
C2081 vdd.n1315 gnd 0.007322f
C2082 vdd.n1316 gnd 0.009097f
C2083 vdd.n1317 gnd 0.009097f
C2084 vdd.n1318 gnd 0.009097f
C2085 vdd.n1319 gnd 0.009097f
C2086 vdd.t94 gnd 0.111913f
C2087 vdd.t95 gnd 0.119604f
C2088 vdd.t92 gnd 0.146157f
C2089 vdd.n1320 gnd 0.187352f
C2090 vdd.n1321 gnd 0.158142f
C2091 vdd.n1322 gnd 0.012008f
C2092 vdd.n1323 gnd 0.003478f
C2093 vdd.n1324 gnd 0.022678f
C2094 vdd.n1325 gnd 0.009097f
C2095 vdd.n1326 gnd 0.003844f
C2096 vdd.n1327 gnd 0.007322f
C2097 vdd.n1328 gnd 0.007322f
C2098 vdd.n1329 gnd 0.009097f
C2099 vdd.n1330 gnd 0.009097f
C2100 vdd.n1331 gnd 0.009097f
C2101 vdd.n1332 gnd 0.007322f
C2102 vdd.n1333 gnd 0.007322f
C2103 vdd.n1334 gnd 0.007322f
C2104 vdd.n1335 gnd 0.009097f
C2105 vdd.n1336 gnd 0.009097f
C2106 vdd.n1337 gnd 0.009097f
C2107 vdd.n1338 gnd 0.007322f
C2108 vdd.n1339 gnd 0.007322f
C2109 vdd.n1340 gnd 0.007322f
C2110 vdd.n1341 gnd 0.009097f
C2111 vdd.n1342 gnd 0.009097f
C2112 vdd.n1343 gnd 0.009097f
C2113 vdd.n1344 gnd 0.007322f
C2114 vdd.n1345 gnd 0.007322f
C2115 vdd.n1346 gnd 0.007322f
C2116 vdd.n1347 gnd 0.009097f
C2117 vdd.n1348 gnd 0.009097f
C2118 vdd.n1349 gnd 0.009097f
C2119 vdd.n1350 gnd 0.007322f
C2120 vdd.n1351 gnd 0.007322f
C2121 vdd.n1352 gnd 0.007322f
C2122 vdd.n1353 gnd 0.009097f
C2123 vdd.n1354 gnd 0.009097f
C2124 vdd.n1355 gnd 0.009097f
C2125 vdd.n1356 gnd 0.007248f
C2126 vdd.n1357 gnd 0.009097f
C2127 vdd.t140 gnd 0.111913f
C2128 vdd.t141 gnd 0.119604f
C2129 vdd.t139 gnd 0.146157f
C2130 vdd.n1358 gnd 0.187352f
C2131 vdd.n1359 gnd 0.158142f
C2132 vdd.n1360 gnd 0.015668f
C2133 vdd.n1361 gnd 0.004979f
C2134 vdd.n1362 gnd 0.009097f
C2135 vdd.n1363 gnd 0.009097f
C2136 vdd.n1364 gnd 0.009097f
C2137 vdd.n1365 gnd 0.007322f
C2138 vdd.n1366 gnd 0.007322f
C2139 vdd.n1367 gnd 0.007322f
C2140 vdd.n1368 gnd 0.009097f
C2141 vdd.n1369 gnd 0.009097f
C2142 vdd.n1370 gnd 0.009097f
C2143 vdd.n1371 gnd 0.007322f
C2144 vdd.n1372 gnd 0.007322f
C2145 vdd.n1373 gnd 0.007322f
C2146 vdd.n1374 gnd 0.009097f
C2147 vdd.n1375 gnd 0.009097f
C2148 vdd.n1376 gnd 0.009097f
C2149 vdd.n1377 gnd 0.007322f
C2150 vdd.n1378 gnd 0.007322f
C2151 vdd.n1379 gnd 0.007322f
C2152 vdd.n1380 gnd 0.009097f
C2153 vdd.n1381 gnd 0.009097f
C2154 vdd.n1382 gnd 0.009097f
C2155 vdd.n1383 gnd 0.007322f
C2156 vdd.n1384 gnd 0.007322f
C2157 vdd.n1385 gnd 0.007322f
C2158 vdd.n1386 gnd 0.009097f
C2159 vdd.n1387 gnd 0.009097f
C2160 vdd.n1388 gnd 0.009097f
C2161 vdd.n1389 gnd 0.007322f
C2162 vdd.n1390 gnd 0.007322f
C2163 vdd.n1391 gnd 0.006114f
C2164 vdd.n1392 gnd 0.009097f
C2165 vdd.n1393 gnd 0.009097f
C2166 vdd.n1394 gnd 0.009097f
C2167 vdd.n1395 gnd 0.006114f
C2168 vdd.n1396 gnd 0.007322f
C2169 vdd.n1397 gnd 0.007322f
C2170 vdd.n1398 gnd 0.009097f
C2171 vdd.n1399 gnd 0.009097f
C2172 vdd.n1400 gnd 0.009097f
C2173 vdd.n1401 gnd 0.007322f
C2174 vdd.n1402 gnd 0.007322f
C2175 vdd.n1403 gnd 0.007322f
C2176 vdd.n1404 gnd 0.009097f
C2177 vdd.n1405 gnd 0.009097f
C2178 vdd.n1406 gnd 0.009097f
C2179 vdd.n1407 gnd 0.007322f
C2180 vdd.n1408 gnd 0.007322f
C2181 vdd.n1409 gnd 0.007322f
C2182 vdd.n1410 gnd 0.009097f
C2183 vdd.n1411 gnd 0.009097f
C2184 vdd.n1412 gnd 0.009097f
C2185 vdd.n1413 gnd 0.007322f
C2186 vdd.n1414 gnd 0.007322f
C2187 vdd.n1415 gnd 0.007322f
C2188 vdd.n1416 gnd 0.009097f
C2189 vdd.n1417 gnd 0.009097f
C2190 vdd.n1418 gnd 0.009097f
C2191 vdd.n1419 gnd 0.007322f
C2192 vdd.n1420 gnd 0.009097f
C2193 vdd.n1421 gnd 2.22183f
C2194 vdd.n1423 gnd 0.022678f
C2195 vdd.n1424 gnd 0.006077f
C2196 vdd.n1425 gnd 0.022678f
C2197 vdd.n1426 gnd 0.022169f
C2198 vdd.n1427 gnd 0.009097f
C2199 vdd.n1428 gnd 0.007322f
C2200 vdd.n1429 gnd 0.009097f
C2201 vdd.n1430 gnd 0.488058f
C2202 vdd.n1431 gnd 0.009097f
C2203 vdd.n1432 gnd 0.007322f
C2204 vdd.n1433 gnd 0.009097f
C2205 vdd.n1434 gnd 0.009097f
C2206 vdd.n1435 gnd 0.009097f
C2207 vdd.n1436 gnd 0.007322f
C2208 vdd.n1437 gnd 0.009097f
C2209 vdd.n1438 gnd 0.832023f
C2210 vdd.n1439 gnd 0.929634f
C2211 vdd.n1440 gnd 0.009097f
C2212 vdd.n1441 gnd 0.007322f
C2213 vdd.n1442 gnd 0.009097f
C2214 vdd.n1443 gnd 0.009097f
C2215 vdd.n1444 gnd 0.009097f
C2216 vdd.n1445 gnd 0.007322f
C2217 vdd.n1446 gnd 0.009097f
C2218 vdd.n1447 gnd 0.562429f
C2219 vdd.n1448 gnd 0.009097f
C2220 vdd.n1449 gnd 0.007322f
C2221 vdd.n1450 gnd 0.009097f
C2222 vdd.n1451 gnd 0.009097f
C2223 vdd.n1452 gnd 0.009097f
C2224 vdd.n1453 gnd 0.007322f
C2225 vdd.n1454 gnd 0.009097f
C2226 vdd.n1455 gnd 0.515947f
C2227 vdd.n1456 gnd 0.720467f
C2228 vdd.n1457 gnd 0.009097f
C2229 vdd.n1458 gnd 0.007322f
C2230 vdd.n1459 gnd 0.009097f
C2231 vdd.n1460 gnd 0.009097f
C2232 vdd.n1461 gnd 0.006991f
C2233 vdd.n1462 gnd 0.009097f
C2234 vdd.n1463 gnd 0.007322f
C2235 vdd.n1464 gnd 0.009097f
C2236 vdd.n1465 gnd 0.771597f
C2237 vdd.n1466 gnd 0.009097f
C2238 vdd.n1467 gnd 0.007322f
C2239 vdd.n1468 gnd 0.009097f
C2240 vdd.n1469 gnd 0.009097f
C2241 vdd.n1470 gnd 0.009097f
C2242 vdd.n1471 gnd 0.007322f
C2243 vdd.n1472 gnd 0.009097f
C2244 vdd.t49 gnd 0.464817f
C2245 vdd.n1473 gnd 0.664689f
C2246 vdd.n1474 gnd 0.009097f
C2247 vdd.n1475 gnd 0.007322f
C2248 vdd.n1476 gnd 0.006991f
C2249 vdd.n1477 gnd 0.009097f
C2250 vdd.n1478 gnd 0.009097f
C2251 vdd.n1479 gnd 0.007322f
C2252 vdd.n1480 gnd 0.009097f
C2253 vdd.n1481 gnd 0.506651f
C2254 vdd.n1482 gnd 0.009097f
C2255 vdd.n1483 gnd 0.007322f
C2256 vdd.n1484 gnd 0.009097f
C2257 vdd.n1485 gnd 0.009097f
C2258 vdd.n1486 gnd 0.009097f
C2259 vdd.n1487 gnd 0.007322f
C2260 vdd.n1488 gnd 0.009097f
C2261 vdd.n1489 gnd 0.655392f
C2262 vdd.n1490 gnd 0.581022f
C2263 vdd.n1491 gnd 0.009097f
C2264 vdd.n1492 gnd 0.007322f
C2265 vdd.n1493 gnd 0.009097f
C2266 vdd.n1494 gnd 0.009097f
C2267 vdd.n1495 gnd 0.009097f
C2268 vdd.n1496 gnd 0.007322f
C2269 vdd.n1497 gnd 0.009097f
C2270 vdd.n1498 gnd 0.739059f
C2271 vdd.n1499 gnd 0.009097f
C2272 vdd.n1500 gnd 0.007322f
C2273 vdd.n1501 gnd 0.009097f
C2274 vdd.n1502 gnd 0.009097f
C2275 vdd.n1503 gnd 0.022169f
C2276 vdd.n1504 gnd 0.009097f
C2277 vdd.n1505 gnd 0.009097f
C2278 vdd.n1506 gnd 0.007322f
C2279 vdd.n1507 gnd 0.009097f
C2280 vdd.n1508 gnd 0.581022f
C2281 vdd.n1509 gnd 0.929634f
C2282 vdd.n1510 gnd 0.009097f
C2283 vdd.n1511 gnd 0.007322f
C2284 vdd.n1512 gnd 0.009097f
C2285 vdd.n1513 gnd 0.009097f
C2286 vdd.n1514 gnd 0.007823f
C2287 vdd.n1515 gnd 0.007322f
C2288 vdd.n1517 gnd 0.009097f
C2289 vdd.n1519 gnd 0.007322f
C2290 vdd.n1520 gnd 0.009097f
C2291 vdd.n1521 gnd 0.007322f
C2292 vdd.n1523 gnd 0.009097f
C2293 vdd.n1524 gnd 0.007322f
C2294 vdd.n1525 gnd 0.009097f
C2295 vdd.n1526 gnd 0.009097f
C2296 vdd.n1527 gnd 0.009097f
C2297 vdd.n1528 gnd 0.009097f
C2298 vdd.n1529 gnd 0.009097f
C2299 vdd.n1530 gnd 0.007322f
C2300 vdd.n1532 gnd 0.009097f
C2301 vdd.n1533 gnd 0.009097f
C2302 vdd.n1534 gnd 0.009097f
C2303 vdd.n1535 gnd 0.009097f
C2304 vdd.n1536 gnd 0.009097f
C2305 vdd.n1537 gnd 0.007322f
C2306 vdd.n1539 gnd 0.009097f
C2307 vdd.n1540 gnd 0.009097f
C2308 vdd.n1541 gnd 0.009097f
C2309 vdd.n1542 gnd 0.009097f
C2310 vdd.n1543 gnd 0.006114f
C2311 vdd.t109 gnd 0.111913f
C2312 vdd.t108 gnd 0.119604f
C2313 vdd.t107 gnd 0.146157f
C2314 vdd.n1544 gnd 0.187352f
C2315 vdd.n1545 gnd 0.15741f
C2316 vdd.n1547 gnd 0.009097f
C2317 vdd.n1548 gnd 0.009097f
C2318 vdd.n1549 gnd 0.007322f
C2319 vdd.n1550 gnd 0.009097f
C2320 vdd.n1552 gnd 0.009097f
C2321 vdd.n1553 gnd 0.009097f
C2322 vdd.n1554 gnd 0.009097f
C2323 vdd.n1555 gnd 0.009097f
C2324 vdd.n1556 gnd 0.007322f
C2325 vdd.n1558 gnd 0.009097f
C2326 vdd.n1559 gnd 0.009097f
C2327 vdd.n1560 gnd 0.009097f
C2328 vdd.n1561 gnd 0.009097f
C2329 vdd.n1562 gnd 0.009097f
C2330 vdd.n1563 gnd 0.007322f
C2331 vdd.n1565 gnd 0.009097f
C2332 vdd.n1566 gnd 0.009097f
C2333 vdd.n1567 gnd 0.009097f
C2334 vdd.n1568 gnd 0.009097f
C2335 vdd.n1569 gnd 0.009097f
C2336 vdd.n1570 gnd 0.007322f
C2337 vdd.n1572 gnd 0.009097f
C2338 vdd.n1573 gnd 0.009097f
C2339 vdd.n1574 gnd 0.009097f
C2340 vdd.n1575 gnd 0.009097f
C2341 vdd.n1576 gnd 0.009097f
C2342 vdd.n1577 gnd 0.007322f
C2343 vdd.n1579 gnd 0.009097f
C2344 vdd.n1580 gnd 0.009097f
C2345 vdd.n1581 gnd 0.009097f
C2346 vdd.n1582 gnd 0.009097f
C2347 vdd.n1583 gnd 0.007248f
C2348 vdd.t102 gnd 0.111913f
C2349 vdd.t101 gnd 0.119604f
C2350 vdd.t100 gnd 0.146157f
C2351 vdd.n1584 gnd 0.187352f
C2352 vdd.n1585 gnd 0.15741f
C2353 vdd.n1587 gnd 0.009097f
C2354 vdd.n1588 gnd 0.009097f
C2355 vdd.n1589 gnd 0.007322f
C2356 vdd.n1590 gnd 0.009097f
C2357 vdd.n1592 gnd 0.009097f
C2358 vdd.n1593 gnd 0.009097f
C2359 vdd.n1594 gnd 0.009097f
C2360 vdd.n1595 gnd 0.009097f
C2361 vdd.n1596 gnd 0.007322f
C2362 vdd.n1598 gnd 0.009097f
C2363 vdd.n1599 gnd 0.009097f
C2364 vdd.n1600 gnd 0.009097f
C2365 vdd.n1601 gnd 0.009097f
C2366 vdd.n1602 gnd 0.009097f
C2367 vdd.n1603 gnd 0.007322f
C2368 vdd.n1605 gnd 0.009097f
C2369 vdd.n1606 gnd 0.009097f
C2370 vdd.n1607 gnd 0.009097f
C2371 vdd.n1608 gnd 0.009097f
C2372 vdd.n1609 gnd 0.009097f
C2373 vdd.n1610 gnd 0.009097f
C2374 vdd.n1611 gnd 0.007322f
C2375 vdd.n1613 gnd 0.009097f
C2376 vdd.n1615 gnd 0.009097f
C2377 vdd.n1616 gnd 0.007322f
C2378 vdd.n1617 gnd 0.007322f
C2379 vdd.n1618 gnd 0.009097f
C2380 vdd.n1620 gnd 0.009097f
C2381 vdd.n1621 gnd 0.007322f
C2382 vdd.n1622 gnd 0.007322f
C2383 vdd.n1623 gnd 0.009097f
C2384 vdd.n1625 gnd 0.009097f
C2385 vdd.n1626 gnd 0.009097f
C2386 vdd.n1627 gnd 0.007322f
C2387 vdd.n1628 gnd 0.007322f
C2388 vdd.n1629 gnd 0.007322f
C2389 vdd.n1630 gnd 0.009097f
C2390 vdd.n1632 gnd 0.009097f
C2391 vdd.n1633 gnd 0.009097f
C2392 vdd.n1634 gnd 0.007322f
C2393 vdd.n1635 gnd 0.007322f
C2394 vdd.n1636 gnd 0.007322f
C2395 vdd.n1637 gnd 0.009097f
C2396 vdd.n1639 gnd 0.009097f
C2397 vdd.n1640 gnd 0.009097f
C2398 vdd.n1641 gnd 0.007322f
C2399 vdd.n1642 gnd 0.007322f
C2400 vdd.n1643 gnd 0.007322f
C2401 vdd.n1644 gnd 0.009097f
C2402 vdd.n1646 gnd 0.009097f
C2403 vdd.n1647 gnd 0.009097f
C2404 vdd.n1648 gnd 0.007322f
C2405 vdd.n1649 gnd 0.009097f
C2406 vdd.n1650 gnd 0.009097f
C2407 vdd.n1651 gnd 0.009097f
C2408 vdd.n1652 gnd 0.014936f
C2409 vdd.n1653 gnd 0.004979f
C2410 vdd.n1654 gnd 0.007322f
C2411 vdd.n1655 gnd 0.009097f
C2412 vdd.n1657 gnd 0.009097f
C2413 vdd.n1658 gnd 0.009097f
C2414 vdd.n1659 gnd 0.007322f
C2415 vdd.n1660 gnd 0.007322f
C2416 vdd.n1661 gnd 0.007322f
C2417 vdd.n1662 gnd 0.009097f
C2418 vdd.n1664 gnd 0.009097f
C2419 vdd.n1665 gnd 0.009097f
C2420 vdd.n1666 gnd 0.007322f
C2421 vdd.n1667 gnd 0.007322f
C2422 vdd.n1668 gnd 0.007322f
C2423 vdd.n1669 gnd 0.009097f
C2424 vdd.n1671 gnd 0.009097f
C2425 vdd.n1672 gnd 0.009097f
C2426 vdd.n1673 gnd 0.007322f
C2427 vdd.n1674 gnd 0.007322f
C2428 vdd.n1675 gnd 0.007322f
C2429 vdd.n1676 gnd 0.009097f
C2430 vdd.n1678 gnd 0.009097f
C2431 vdd.n1679 gnd 0.009097f
C2432 vdd.n1680 gnd 0.007322f
C2433 vdd.n1681 gnd 0.007322f
C2434 vdd.n1682 gnd 0.007322f
C2435 vdd.n1683 gnd 0.009097f
C2436 vdd.n1685 gnd 0.009097f
C2437 vdd.n1686 gnd 0.009097f
C2438 vdd.n1687 gnd 0.007322f
C2439 vdd.n1688 gnd 0.009097f
C2440 vdd.n1689 gnd 0.009097f
C2441 vdd.n1690 gnd 0.009097f
C2442 vdd.n1691 gnd 0.014936f
C2443 vdd.n1692 gnd 0.006114f
C2444 vdd.n1693 gnd 0.007322f
C2445 vdd.n1694 gnd 0.009097f
C2446 vdd.n1696 gnd 0.009097f
C2447 vdd.n1697 gnd 0.009097f
C2448 vdd.n1698 gnd 0.007322f
C2449 vdd.n1699 gnd 0.007322f
C2450 vdd.n1700 gnd 0.007322f
C2451 vdd.n1701 gnd 0.009097f
C2452 vdd.n1703 gnd 0.009097f
C2453 vdd.n1704 gnd 0.009097f
C2454 vdd.n1705 gnd 0.007322f
C2455 vdd.n1706 gnd 0.007322f
C2456 vdd.n1707 gnd 0.007322f
C2457 vdd.n1708 gnd 0.009097f
C2458 vdd.n1710 gnd 0.009097f
C2459 vdd.n1711 gnd 0.009097f
C2460 vdd.n1713 gnd 0.009097f
C2461 vdd.n1714 gnd 0.007322f
C2462 vdd.n1715 gnd 0.005822f
C2463 vdd.n1716 gnd 0.006186f
C2464 vdd.n1717 gnd 0.006186f
C2465 vdd.n1718 gnd 0.006186f
C2466 vdd.n1719 gnd 0.006186f
C2467 vdd.n1720 gnd 0.006186f
C2468 vdd.n1721 gnd 0.006186f
C2469 vdd.n1722 gnd 0.006186f
C2470 vdd.n1723 gnd 0.006186f
C2471 vdd.n1725 gnd 0.006186f
C2472 vdd.n1726 gnd 0.006186f
C2473 vdd.n1727 gnd 0.006186f
C2474 vdd.n1728 gnd 0.006186f
C2475 vdd.n1729 gnd 0.006186f
C2476 vdd.n1731 gnd 0.006186f
C2477 vdd.n1733 gnd 0.006186f
C2478 vdd.n1734 gnd 0.006186f
C2479 vdd.n1735 gnd 0.006186f
C2480 vdd.n1736 gnd 0.006186f
C2481 vdd.n1737 gnd 0.006186f
C2482 vdd.n1739 gnd 0.006186f
C2483 vdd.n1741 gnd 0.006186f
C2484 vdd.n1742 gnd 0.006186f
C2485 vdd.n1743 gnd 0.006186f
C2486 vdd.n1744 gnd 0.006186f
C2487 vdd.n1745 gnd 0.006186f
C2488 vdd.n1747 gnd 0.006186f
C2489 vdd.n1749 gnd 0.006186f
C2490 vdd.n1750 gnd 0.006186f
C2491 vdd.n1751 gnd 0.006186f
C2492 vdd.n1752 gnd 0.006186f
C2493 vdd.n1753 gnd 0.006186f
C2494 vdd.n1755 gnd 0.006186f
C2495 vdd.n1756 gnd 0.006186f
C2496 vdd.n1757 gnd 0.006186f
C2497 vdd.n1758 gnd 0.006186f
C2498 vdd.n1759 gnd 0.006186f
C2499 vdd.n1760 gnd 0.006186f
C2500 vdd.n1761 gnd 0.006186f
C2501 vdd.n1762 gnd 0.006186f
C2502 vdd.n1763 gnd 0.004503f
C2503 vdd.n1764 gnd 0.006186f
C2504 vdd.t155 gnd 0.249964f
C2505 vdd.t156 gnd 0.255869f
C2506 vdd.t154 gnd 0.163186f
C2507 vdd.n1765 gnd 0.088193f
C2508 vdd.n1766 gnd 0.050026f
C2509 vdd.n1767 gnd 0.00884f
C2510 vdd.n1768 gnd 0.006186f
C2511 vdd.n1769 gnd 0.006186f
C2512 vdd.n1770 gnd 0.376502f
C2513 vdd.n1771 gnd 0.006186f
C2514 vdd.n1772 gnd 0.006186f
C2515 vdd.n1773 gnd 0.006186f
C2516 vdd.n1774 gnd 0.006186f
C2517 vdd.n1775 gnd 0.006186f
C2518 vdd.n1776 gnd 0.006186f
C2519 vdd.n1777 gnd 0.006186f
C2520 vdd.n1778 gnd 0.006186f
C2521 vdd.n1779 gnd 0.006186f
C2522 vdd.n1780 gnd 0.006186f
C2523 vdd.n1781 gnd 0.006186f
C2524 vdd.n1782 gnd 0.006186f
C2525 vdd.n1783 gnd 0.006186f
C2526 vdd.n1784 gnd 0.006186f
C2527 vdd.n1785 gnd 0.006186f
C2528 vdd.n1786 gnd 0.006186f
C2529 vdd.n1787 gnd 0.006186f
C2530 vdd.n1788 gnd 0.006186f
C2531 vdd.n1789 gnd 0.006186f
C2532 vdd.n1790 gnd 0.006186f
C2533 vdd.t130 gnd 0.249964f
C2534 vdd.t131 gnd 0.255869f
C2535 vdd.t128 gnd 0.163186f
C2536 vdd.n1791 gnd 0.088193f
C2537 vdd.n1792 gnd 0.050026f
C2538 vdd.n1793 gnd 0.006186f
C2539 vdd.n1794 gnd 0.006186f
C2540 vdd.n1795 gnd 0.006186f
C2541 vdd.n1796 gnd 0.006186f
C2542 vdd.n1797 gnd 0.006186f
C2543 vdd.n1798 gnd 0.006186f
C2544 vdd.n1800 gnd 0.006186f
C2545 vdd.n1801 gnd 0.006186f
C2546 vdd.n1802 gnd 0.006186f
C2547 vdd.n1803 gnd 0.006186f
C2548 vdd.n1805 gnd 0.006186f
C2549 vdd.n1807 gnd 0.006186f
C2550 vdd.n1808 gnd 0.006186f
C2551 vdd.n1809 gnd 0.006186f
C2552 vdd.n1810 gnd 0.006186f
C2553 vdd.n1811 gnd 0.006186f
C2554 vdd.n1813 gnd 0.006186f
C2555 vdd.n1815 gnd 0.006186f
C2556 vdd.n1816 gnd 0.006186f
C2557 vdd.n1817 gnd 0.006186f
C2558 vdd.n1818 gnd 0.006186f
C2559 vdd.n1819 gnd 0.006186f
C2560 vdd.n1821 gnd 0.006186f
C2561 vdd.n1823 gnd 0.006186f
C2562 vdd.n1824 gnd 0.006186f
C2563 vdd.n1825 gnd 0.004503f
C2564 vdd.n1826 gnd 0.00884f
C2565 vdd.n1827 gnd 0.004776f
C2566 vdd.n1828 gnd 0.006186f
C2567 vdd.n1830 gnd 0.006186f
C2568 vdd.n1831 gnd 0.014678f
C2569 vdd.n1832 gnd 0.014678f
C2570 vdd.n1833 gnd 0.013704f
C2571 vdd.n1834 gnd 0.006186f
C2572 vdd.n1835 gnd 0.006186f
C2573 vdd.n1836 gnd 0.006186f
C2574 vdd.n1837 gnd 0.006186f
C2575 vdd.n1838 gnd 0.006186f
C2576 vdd.n1839 gnd 0.006186f
C2577 vdd.n1840 gnd 0.006186f
C2578 vdd.n1841 gnd 0.006186f
C2579 vdd.n1842 gnd 0.006186f
C2580 vdd.n1843 gnd 0.006186f
C2581 vdd.n1844 gnd 0.006186f
C2582 vdd.n1845 gnd 0.006186f
C2583 vdd.n1846 gnd 0.006186f
C2584 vdd.n1847 gnd 0.006186f
C2585 vdd.n1848 gnd 0.006186f
C2586 vdd.n1849 gnd 0.006186f
C2587 vdd.n1850 gnd 0.006186f
C2588 vdd.n1851 gnd 0.006186f
C2589 vdd.n1852 gnd 0.006186f
C2590 vdd.n1853 gnd 0.006186f
C2591 vdd.n1854 gnd 0.006186f
C2592 vdd.n1855 gnd 0.006186f
C2593 vdd.n1856 gnd 0.006186f
C2594 vdd.n1857 gnd 0.006186f
C2595 vdd.n1858 gnd 0.006186f
C2596 vdd.n1859 gnd 0.006186f
C2597 vdd.n1860 gnd 0.006186f
C2598 vdd.n1861 gnd 0.006186f
C2599 vdd.n1862 gnd 0.006186f
C2600 vdd.n1863 gnd 0.006186f
C2601 vdd.n1864 gnd 0.006186f
C2602 vdd.n1865 gnd 0.006186f
C2603 vdd.n1866 gnd 0.006186f
C2604 vdd.n1867 gnd 0.006186f
C2605 vdd.n1868 gnd 0.006186f
C2606 vdd.n1869 gnd 0.006186f
C2607 vdd.n1870 gnd 0.006186f
C2608 vdd.n1871 gnd 0.199871f
C2609 vdd.n1872 gnd 0.006186f
C2610 vdd.n1873 gnd 0.006186f
C2611 vdd.n1874 gnd 0.006186f
C2612 vdd.n1875 gnd 0.006186f
C2613 vdd.n1876 gnd 0.006186f
C2614 vdd.n1877 gnd 0.006186f
C2615 vdd.n1878 gnd 0.006186f
C2616 vdd.n1879 gnd 0.006186f
C2617 vdd.n1880 gnd 0.006186f
C2618 vdd.n1881 gnd 0.006186f
C2619 vdd.n1882 gnd 0.006186f
C2620 vdd.n1883 gnd 0.006186f
C2621 vdd.n1884 gnd 0.006186f
C2622 vdd.n1885 gnd 0.006186f
C2623 vdd.n1886 gnd 0.006186f
C2624 vdd.n1887 gnd 0.006186f
C2625 vdd.n1888 gnd 0.006186f
C2626 vdd.n1889 gnd 0.006186f
C2627 vdd.n1890 gnd 0.006186f
C2628 vdd.n1891 gnd 0.006186f
C2629 vdd.n1892 gnd 0.013704f
C2630 vdd.n1894 gnd 0.014678f
C2631 vdd.n1895 gnd 0.014678f
C2632 vdd.n1896 gnd 0.006186f
C2633 vdd.n1897 gnd 0.004776f
C2634 vdd.n1898 gnd 0.006186f
C2635 vdd.n1900 gnd 0.006186f
C2636 vdd.n1902 gnd 0.006186f
C2637 vdd.n1903 gnd 0.006186f
C2638 vdd.n1904 gnd 0.006186f
C2639 vdd.n1905 gnd 0.006186f
C2640 vdd.n1906 gnd 0.006186f
C2641 vdd.n1908 gnd 0.006186f
C2642 vdd.n1910 gnd 0.006186f
C2643 vdd.n1911 gnd 0.006186f
C2644 vdd.n1912 gnd 0.006186f
C2645 vdd.n1913 gnd 0.006186f
C2646 vdd.n1914 gnd 0.006186f
C2647 vdd.n1916 gnd 0.006186f
C2648 vdd.n1918 gnd 0.006186f
C2649 vdd.n1919 gnd 0.006186f
C2650 vdd.n1920 gnd 0.006186f
C2651 vdd.n1921 gnd 0.006186f
C2652 vdd.n1922 gnd 0.006186f
C2653 vdd.n1924 gnd 0.006186f
C2654 vdd.n1926 gnd 0.006186f
C2655 vdd.n1927 gnd 0.006186f
C2656 vdd.n1928 gnd 0.018451f
C2657 vdd.n1929 gnd 0.546958f
C2658 vdd.n1931 gnd 0.007322f
C2659 vdd.n1932 gnd 0.007322f
C2660 vdd.n1933 gnd 0.009097f
C2661 vdd.n1935 gnd 0.009097f
C2662 vdd.n1936 gnd 0.009097f
C2663 vdd.n1937 gnd 0.007322f
C2664 vdd.n1938 gnd 0.006077f
C2665 vdd.n1939 gnd 0.022678f
C2666 vdd.n1940 gnd 0.022169f
C2667 vdd.n1941 gnd 0.006077f
C2668 vdd.n1942 gnd 0.022169f
C2669 vdd.n1943 gnd 1.27825f
C2670 vdd.n1944 gnd 0.022169f
C2671 vdd.n1945 gnd 0.022678f
C2672 vdd.n1946 gnd 0.003478f
C2673 vdd.t91 gnd 0.111913f
C2674 vdd.t90 gnd 0.119604f
C2675 vdd.t88 gnd 0.146157f
C2676 vdd.n1947 gnd 0.187352f
C2677 vdd.n1948 gnd 0.15741f
C2678 vdd.n1949 gnd 0.011275f
C2679 vdd.n1950 gnd 0.003844f
C2680 vdd.n1951 gnd 0.007823f
C2681 vdd.n1952 gnd 0.546958f
C2682 vdd.n1953 gnd 0.018451f
C2683 vdd.n1954 gnd 0.006186f
C2684 vdd.n1955 gnd 0.006186f
C2685 vdd.n1956 gnd 0.006186f
C2686 vdd.n1958 gnd 0.006186f
C2687 vdd.n1960 gnd 0.006186f
C2688 vdd.n1961 gnd 0.006186f
C2689 vdd.n1962 gnd 0.006186f
C2690 vdd.n1963 gnd 0.006186f
C2691 vdd.n1964 gnd 0.006186f
C2692 vdd.n1966 gnd 0.006186f
C2693 vdd.n1968 gnd 0.006186f
C2694 vdd.n1969 gnd 0.006186f
C2695 vdd.n1970 gnd 0.006186f
C2696 vdd.n1971 gnd 0.006186f
C2697 vdd.n1972 gnd 0.006186f
C2698 vdd.n1974 gnd 0.006186f
C2699 vdd.n1976 gnd 0.006186f
C2700 vdd.n1977 gnd 0.006186f
C2701 vdd.n1978 gnd 0.006186f
C2702 vdd.n1979 gnd 0.006186f
C2703 vdd.n1980 gnd 0.006186f
C2704 vdd.n1982 gnd 0.006186f
C2705 vdd.n1984 gnd 0.006186f
C2706 vdd.n1985 gnd 0.006186f
C2707 vdd.n1986 gnd 0.014678f
C2708 vdd.n1987 gnd 0.013704f
C2709 vdd.n1988 gnd 0.013704f
C2710 vdd.n1989 gnd 0.911042f
C2711 vdd.n1990 gnd 0.013704f
C2712 vdd.n1991 gnd 0.013704f
C2713 vdd.n1992 gnd 0.006186f
C2714 vdd.n1993 gnd 0.006186f
C2715 vdd.n1994 gnd 0.006186f
C2716 vdd.n1995 gnd 0.395095f
C2717 vdd.n1996 gnd 0.006186f
C2718 vdd.n1997 gnd 0.006186f
C2719 vdd.n1998 gnd 0.006186f
C2720 vdd.n1999 gnd 0.006186f
C2721 vdd.n2000 gnd 0.006186f
C2722 vdd.n2001 gnd 0.632151f
C2723 vdd.n2002 gnd 0.006186f
C2724 vdd.n2003 gnd 0.006186f
C2725 vdd.n2004 gnd 0.006186f
C2726 vdd.n2005 gnd 0.006186f
C2727 vdd.n2006 gnd 0.006186f
C2728 vdd.n2007 gnd 0.632151f
C2729 vdd.n2008 gnd 0.006186f
C2730 vdd.n2009 gnd 0.006186f
C2731 vdd.n2010 gnd 0.005458f
C2732 vdd.n2011 gnd 0.017919f
C2733 vdd.n2012 gnd 0.003821f
C2734 vdd.n2013 gnd 0.006186f
C2735 vdd.n2014 gnd 0.348613f
C2736 vdd.n2015 gnd 0.006186f
C2737 vdd.n2016 gnd 0.006186f
C2738 vdd.n2017 gnd 0.006186f
C2739 vdd.n2018 gnd 0.006186f
C2740 vdd.n2019 gnd 0.006186f
C2741 vdd.n2020 gnd 0.422984f
C2742 vdd.n2021 gnd 0.006186f
C2743 vdd.n2022 gnd 0.006186f
C2744 vdd.n2023 gnd 0.006186f
C2745 vdd.n2024 gnd 0.006186f
C2746 vdd.n2025 gnd 0.006186f
C2747 vdd.n2026 gnd 0.562429f
C2748 vdd.n2027 gnd 0.006186f
C2749 vdd.n2028 gnd 0.006186f
C2750 vdd.n2029 gnd 0.006186f
C2751 vdd.n2030 gnd 0.006186f
C2752 vdd.n2031 gnd 0.006186f
C2753 vdd.n2032 gnd 0.502003f
C2754 vdd.n2033 gnd 0.006186f
C2755 vdd.n2034 gnd 0.006186f
C2756 vdd.n2035 gnd 0.006186f
C2757 vdd.n2036 gnd 0.006186f
C2758 vdd.n2037 gnd 0.006186f
C2759 vdd.n2038 gnd 0.362557f
C2760 vdd.n2039 gnd 0.006186f
C2761 vdd.n2040 gnd 0.006186f
C2762 vdd.n2041 gnd 0.006186f
C2763 vdd.n2042 gnd 0.006186f
C2764 vdd.n2043 gnd 0.006186f
C2765 vdd.n2044 gnd 0.199871f
C2766 vdd.n2045 gnd 0.006186f
C2767 vdd.n2046 gnd 0.006186f
C2768 vdd.n2047 gnd 0.006186f
C2769 vdd.n2048 gnd 0.006186f
C2770 vdd.n2049 gnd 0.006186f
C2771 vdd.n2050 gnd 0.348613f
C2772 vdd.n2051 gnd 0.006186f
C2773 vdd.n2052 gnd 0.006186f
C2774 vdd.n2053 gnd 0.006186f
C2775 vdd.n2054 gnd 0.006186f
C2776 vdd.n2055 gnd 0.006186f
C2777 vdd.n2056 gnd 0.632151f
C2778 vdd.n2057 gnd 0.006186f
C2779 vdd.n2058 gnd 0.006186f
C2780 vdd.n2059 gnd 0.006186f
C2781 vdd.n2060 gnd 0.006186f
C2782 vdd.n2061 gnd 0.006186f
C2783 vdd.n2062 gnd 0.006186f
C2784 vdd.n2063 gnd 0.006186f
C2785 vdd.n2064 gnd 0.492706f
C2786 vdd.n2065 gnd 0.006186f
C2787 vdd.n2066 gnd 0.006186f
C2788 vdd.n2067 gnd 0.006186f
C2789 vdd.n2068 gnd 0.006186f
C2790 vdd.n2069 gnd 0.006186f
C2791 vdd.n2070 gnd 0.006186f
C2792 vdd.n2071 gnd 0.395095f
C2793 vdd.n2072 gnd 0.006186f
C2794 vdd.n2073 gnd 0.006186f
C2795 vdd.n2074 gnd 0.006186f
C2796 vdd.n2075 gnd 0.014457f
C2797 vdd.n2076 gnd 0.013924f
C2798 vdd.n2077 gnd 0.006186f
C2799 vdd.n2078 gnd 0.006186f
C2800 vdd.n2079 gnd 0.004776f
C2801 vdd.n2080 gnd 0.006186f
C2802 vdd.n2081 gnd 0.006186f
C2803 vdd.n2082 gnd 0.004503f
C2804 vdd.n2083 gnd 0.006186f
C2805 vdd.n2084 gnd 0.006186f
C2806 vdd.n2085 gnd 0.006186f
C2807 vdd.n2086 gnd 0.006186f
C2808 vdd.n2087 gnd 0.006186f
C2809 vdd.n2088 gnd 0.006186f
C2810 vdd.n2089 gnd 0.006186f
C2811 vdd.n2090 gnd 0.006186f
C2812 vdd.n2091 gnd 0.006186f
C2813 vdd.n2092 gnd 0.006186f
C2814 vdd.n2093 gnd 0.006186f
C2815 vdd.n2094 gnd 0.006186f
C2816 vdd.n2095 gnd 0.006186f
C2817 vdd.n2096 gnd 0.006186f
C2818 vdd.n2097 gnd 0.006186f
C2819 vdd.n2098 gnd 0.006186f
C2820 vdd.n2099 gnd 0.006186f
C2821 vdd.n2100 gnd 0.006186f
C2822 vdd.n2101 gnd 0.006186f
C2823 vdd.n2102 gnd 0.006186f
C2824 vdd.n2103 gnd 0.006186f
C2825 vdd.n2104 gnd 0.006186f
C2826 vdd.n2105 gnd 0.006186f
C2827 vdd.n2106 gnd 0.006186f
C2828 vdd.n2107 gnd 0.006186f
C2829 vdd.n2108 gnd 0.006186f
C2830 vdd.n2109 gnd 0.006186f
C2831 vdd.n2110 gnd 0.006186f
C2832 vdd.n2111 gnd 0.006186f
C2833 vdd.n2112 gnd 0.006186f
C2834 vdd.n2113 gnd 0.006186f
C2835 vdd.n2114 gnd 0.006186f
C2836 vdd.n2115 gnd 0.006186f
C2837 vdd.n2116 gnd 0.006186f
C2838 vdd.n2117 gnd 0.006186f
C2839 vdd.n2118 gnd 0.006186f
C2840 vdd.n2119 gnd 0.006186f
C2841 vdd.n2120 gnd 0.006186f
C2842 vdd.n2121 gnd 0.006186f
C2843 vdd.n2122 gnd 0.006186f
C2844 vdd.n2123 gnd 0.006186f
C2845 vdd.n2124 gnd 0.006186f
C2846 vdd.n2125 gnd 0.006186f
C2847 vdd.n2126 gnd 0.006186f
C2848 vdd.n2127 gnd 0.006186f
C2849 vdd.n2128 gnd 0.006186f
C2850 vdd.n2129 gnd 0.006186f
C2851 vdd.n2130 gnd 0.006186f
C2852 vdd.n2131 gnd 0.006186f
C2853 vdd.n2132 gnd 0.006186f
C2854 vdd.n2133 gnd 0.006186f
C2855 vdd.n2134 gnd 0.006186f
C2856 vdd.n2135 gnd 0.006186f
C2857 vdd.n2136 gnd 0.006186f
C2858 vdd.n2137 gnd 0.006186f
C2859 vdd.n2138 gnd 0.006186f
C2860 vdd.n2139 gnd 0.006186f
C2861 vdd.n2140 gnd 0.006186f
C2862 vdd.n2141 gnd 0.006186f
C2863 vdd.n2142 gnd 0.006186f
C2864 vdd.n2143 gnd 0.014678f
C2865 vdd.n2144 gnd 0.013704f
C2866 vdd.n2145 gnd 0.013704f
C2867 vdd.n2146 gnd 0.771597f
C2868 vdd.n2147 gnd 0.013704f
C2869 vdd.n2148 gnd 0.014678f
C2870 vdd.n2149 gnd 0.013924f
C2871 vdd.n2150 gnd 0.006186f
C2872 vdd.n2151 gnd 0.006186f
C2873 vdd.n2152 gnd 0.006186f
C2874 vdd.n2153 gnd 0.004776f
C2875 vdd.n2154 gnd 0.00884f
C2876 vdd.n2155 gnd 0.004503f
C2877 vdd.n2156 gnd 0.006186f
C2878 vdd.n2157 gnd 0.006186f
C2879 vdd.n2158 gnd 0.006186f
C2880 vdd.n2159 gnd 0.006186f
C2881 vdd.n2160 gnd 0.006186f
C2882 vdd.n2161 gnd 0.006186f
C2883 vdd.n2162 gnd 0.006186f
C2884 vdd.n2163 gnd 0.006186f
C2885 vdd.n2164 gnd 0.006186f
C2886 vdd.n2165 gnd 0.006186f
C2887 vdd.n2166 gnd 0.006186f
C2888 vdd.n2167 gnd 0.006186f
C2889 vdd.n2168 gnd 0.006186f
C2890 vdd.n2169 gnd 0.006186f
C2891 vdd.n2170 gnd 0.006186f
C2892 vdd.n2171 gnd 0.006186f
C2893 vdd.n2172 gnd 0.006186f
C2894 vdd.n2173 gnd 0.006186f
C2895 vdd.n2174 gnd 0.006186f
C2896 vdd.n2175 gnd 0.006186f
C2897 vdd.n2176 gnd 0.006186f
C2898 vdd.n2177 gnd 0.006186f
C2899 vdd.n2178 gnd 0.006186f
C2900 vdd.n2179 gnd 0.006186f
C2901 vdd.n2180 gnd 0.006186f
C2902 vdd.n2181 gnd 0.006186f
C2903 vdd.n2182 gnd 0.006186f
C2904 vdd.n2183 gnd 0.006186f
C2905 vdd.n2184 gnd 0.006186f
C2906 vdd.n2185 gnd 0.006186f
C2907 vdd.n2186 gnd 0.006186f
C2908 vdd.n2187 gnd 0.006186f
C2909 vdd.n2188 gnd 0.006186f
C2910 vdd.n2189 gnd 0.006186f
C2911 vdd.n2190 gnd 0.006186f
C2912 vdd.n2191 gnd 0.006186f
C2913 vdd.n2192 gnd 0.006186f
C2914 vdd.n2193 gnd 0.006186f
C2915 vdd.n2194 gnd 0.006186f
C2916 vdd.n2195 gnd 0.006186f
C2917 vdd.n2196 gnd 0.006186f
C2918 vdd.n2197 gnd 0.006186f
C2919 vdd.n2198 gnd 0.006186f
C2920 vdd.n2199 gnd 0.006186f
C2921 vdd.n2200 gnd 0.006186f
C2922 vdd.n2201 gnd 0.006186f
C2923 vdd.n2202 gnd 0.006186f
C2924 vdd.n2203 gnd 0.006186f
C2925 vdd.n2204 gnd 0.006186f
C2926 vdd.n2205 gnd 0.006186f
C2927 vdd.n2206 gnd 0.006186f
C2928 vdd.n2207 gnd 0.006186f
C2929 vdd.n2208 gnd 0.006186f
C2930 vdd.n2209 gnd 0.006186f
C2931 vdd.n2210 gnd 0.006186f
C2932 vdd.n2211 gnd 0.006186f
C2933 vdd.n2212 gnd 0.006186f
C2934 vdd.n2213 gnd 0.006186f
C2935 vdd.n2214 gnd 0.006186f
C2936 vdd.n2215 gnd 0.006186f
C2937 vdd.n2216 gnd 0.014678f
C2938 vdd.n2217 gnd 0.014678f
C2939 vdd.n2218 gnd 0.771597f
C2940 vdd.t79 gnd 2.74242f
C2941 vdd.t181 gnd 2.74242f
C2942 vdd.n2251 gnd 0.014678f
C2943 vdd.n2252 gnd 0.006186f
C2944 vdd.t123 gnd 0.249964f
C2945 vdd.t124 gnd 0.255869f
C2946 vdd.t121 gnd 0.163186f
C2947 vdd.n2253 gnd 0.088193f
C2948 vdd.n2254 gnd 0.050026f
C2949 vdd.n2255 gnd 0.006186f
C2950 vdd.t137 gnd 0.249964f
C2951 vdd.t138 gnd 0.255869f
C2952 vdd.t136 gnd 0.163186f
C2953 vdd.n2256 gnd 0.088193f
C2954 vdd.n2257 gnd 0.050026f
C2955 vdd.n2258 gnd 0.00884f
C2956 vdd.n2259 gnd 0.006186f
C2957 vdd.n2260 gnd 0.006186f
C2958 vdd.n2261 gnd 0.006186f
C2959 vdd.n2262 gnd 0.006186f
C2960 vdd.n2263 gnd 0.006186f
C2961 vdd.n2264 gnd 0.006186f
C2962 vdd.n2265 gnd 0.006186f
C2963 vdd.n2266 gnd 0.006186f
C2964 vdd.n2267 gnd 0.006186f
C2965 vdd.n2268 gnd 0.006186f
C2966 vdd.n2269 gnd 0.006186f
C2967 vdd.n2270 gnd 0.006186f
C2968 vdd.n2271 gnd 0.006186f
C2969 vdd.n2272 gnd 0.006186f
C2970 vdd.n2273 gnd 0.006186f
C2971 vdd.n2274 gnd 0.006186f
C2972 vdd.n2275 gnd 0.006186f
C2973 vdd.n2276 gnd 0.006186f
C2974 vdd.n2277 gnd 0.006186f
C2975 vdd.n2278 gnd 0.006186f
C2976 vdd.n2279 gnd 0.006186f
C2977 vdd.n2280 gnd 0.006186f
C2978 vdd.n2281 gnd 0.006186f
C2979 vdd.n2282 gnd 0.006186f
C2980 vdd.n2283 gnd 0.006186f
C2981 vdd.n2284 gnd 0.006186f
C2982 vdd.n2285 gnd 0.006186f
C2983 vdd.n2286 gnd 0.006186f
C2984 vdd.n2287 gnd 0.006186f
C2985 vdd.n2288 gnd 0.006186f
C2986 vdd.n2289 gnd 0.006186f
C2987 vdd.n2290 gnd 0.006186f
C2988 vdd.n2291 gnd 0.006186f
C2989 vdd.n2292 gnd 0.006186f
C2990 vdd.n2293 gnd 0.006186f
C2991 vdd.n2294 gnd 0.006186f
C2992 vdd.n2295 gnd 0.006186f
C2993 vdd.n2296 gnd 0.006186f
C2994 vdd.n2297 gnd 0.006186f
C2995 vdd.n2298 gnd 0.006186f
C2996 vdd.n2299 gnd 0.006186f
C2997 vdd.n2300 gnd 0.006186f
C2998 vdd.n2301 gnd 0.006186f
C2999 vdd.n2302 gnd 0.006186f
C3000 vdd.n2303 gnd 0.006186f
C3001 vdd.n2304 gnd 0.006186f
C3002 vdd.n2305 gnd 0.006186f
C3003 vdd.n2306 gnd 0.006186f
C3004 vdd.n2307 gnd 0.006186f
C3005 vdd.n2308 gnd 0.006186f
C3006 vdd.n2309 gnd 0.006186f
C3007 vdd.n2310 gnd 0.006186f
C3008 vdd.n2311 gnd 0.006186f
C3009 vdd.n2312 gnd 0.006186f
C3010 vdd.n2313 gnd 0.006186f
C3011 vdd.n2314 gnd 0.006186f
C3012 vdd.n2315 gnd 0.004503f
C3013 vdd.n2316 gnd 0.006186f
C3014 vdd.n2317 gnd 0.006186f
C3015 vdd.n2318 gnd 0.004776f
C3016 vdd.n2319 gnd 0.006186f
C3017 vdd.n2320 gnd 0.006186f
C3018 vdd.n2321 gnd 0.014678f
C3019 vdd.n2322 gnd 0.013704f
C3020 vdd.n2323 gnd 0.006186f
C3021 vdd.n2324 gnd 0.006186f
C3022 vdd.n2325 gnd 0.006186f
C3023 vdd.n2326 gnd 0.006186f
C3024 vdd.n2327 gnd 0.006186f
C3025 vdd.n2328 gnd 0.006186f
C3026 vdd.n2329 gnd 0.006186f
C3027 vdd.n2330 gnd 0.006186f
C3028 vdd.n2331 gnd 0.006186f
C3029 vdd.n2332 gnd 0.006186f
C3030 vdd.n2333 gnd 0.006186f
C3031 vdd.n2334 gnd 0.006186f
C3032 vdd.n2335 gnd 0.006186f
C3033 vdd.n2336 gnd 0.006186f
C3034 vdd.n2337 gnd 0.006186f
C3035 vdd.n2338 gnd 0.006186f
C3036 vdd.n2339 gnd 0.006186f
C3037 vdd.n2340 gnd 0.006186f
C3038 vdd.n2341 gnd 0.006186f
C3039 vdd.n2342 gnd 0.006186f
C3040 vdd.n2343 gnd 0.006186f
C3041 vdd.n2344 gnd 0.006186f
C3042 vdd.n2345 gnd 0.006186f
C3043 vdd.n2346 gnd 0.006186f
C3044 vdd.n2347 gnd 0.006186f
C3045 vdd.n2348 gnd 0.006186f
C3046 vdd.n2349 gnd 0.006186f
C3047 vdd.n2350 gnd 0.006186f
C3048 vdd.n2351 gnd 0.006186f
C3049 vdd.n2352 gnd 0.006186f
C3050 vdd.n2353 gnd 0.006186f
C3051 vdd.n2354 gnd 0.006186f
C3052 vdd.n2355 gnd 0.006186f
C3053 vdd.n2356 gnd 0.006186f
C3054 vdd.n2357 gnd 0.006186f
C3055 vdd.n2358 gnd 0.006186f
C3056 vdd.n2359 gnd 0.006186f
C3057 vdd.n2360 gnd 0.006186f
C3058 vdd.n2361 gnd 0.006186f
C3059 vdd.n2362 gnd 0.006186f
C3060 vdd.n2363 gnd 0.006186f
C3061 vdd.n2364 gnd 0.006186f
C3062 vdd.n2365 gnd 0.006186f
C3063 vdd.n2366 gnd 0.006186f
C3064 vdd.n2367 gnd 0.006186f
C3065 vdd.n2368 gnd 0.006186f
C3066 vdd.n2369 gnd 0.006186f
C3067 vdd.n2370 gnd 0.006186f
C3068 vdd.n2371 gnd 0.006186f
C3069 vdd.n2372 gnd 0.006186f
C3070 vdd.n2373 gnd 0.006186f
C3071 vdd.n2374 gnd 0.199871f
C3072 vdd.n2375 gnd 0.006186f
C3073 vdd.n2376 gnd 0.006186f
C3074 vdd.n2377 gnd 0.006186f
C3075 vdd.n2378 gnd 0.006186f
C3076 vdd.n2379 gnd 0.006186f
C3077 vdd.n2380 gnd 0.006186f
C3078 vdd.n2381 gnd 0.006186f
C3079 vdd.n2382 gnd 0.006186f
C3080 vdd.n2383 gnd 0.006186f
C3081 vdd.n2384 gnd 0.006186f
C3082 vdd.n2385 gnd 0.006186f
C3083 vdd.n2386 gnd 0.006186f
C3084 vdd.n2387 gnd 0.006186f
C3085 vdd.n2388 gnd 0.006186f
C3086 vdd.n2389 gnd 0.006186f
C3087 vdd.n2390 gnd 0.006186f
C3088 vdd.n2391 gnd 0.006186f
C3089 vdd.n2392 gnd 0.006186f
C3090 vdd.n2393 gnd 0.006186f
C3091 vdd.n2394 gnd 0.006186f
C3092 vdd.n2395 gnd 0.376502f
C3093 vdd.n2396 gnd 0.006186f
C3094 vdd.n2397 gnd 0.006186f
C3095 vdd.n2398 gnd 0.006186f
C3096 vdd.n2399 gnd 0.006186f
C3097 vdd.n2400 gnd 0.006186f
C3098 vdd.n2401 gnd 0.013704f
C3099 vdd.n2402 gnd 0.014678f
C3100 vdd.n2403 gnd 0.014678f
C3101 vdd.n2404 gnd 0.006186f
C3102 vdd.n2405 gnd 0.006186f
C3103 vdd.n2406 gnd 0.006186f
C3104 vdd.n2407 gnd 0.004776f
C3105 vdd.n2408 gnd 0.00884f
C3106 vdd.n2409 gnd 0.004503f
C3107 vdd.n2410 gnd 0.006186f
C3108 vdd.n2411 gnd 0.006186f
C3109 vdd.n2412 gnd 0.006186f
C3110 vdd.n2413 gnd 0.006186f
C3111 vdd.n2414 gnd 0.006186f
C3112 vdd.n2415 gnd 0.006186f
C3113 vdd.n2416 gnd 0.006186f
C3114 vdd.n2417 gnd 0.006186f
C3115 vdd.n2418 gnd 0.006186f
C3116 vdd.n2419 gnd 0.006186f
C3117 vdd.n2420 gnd 0.006186f
C3118 vdd.n2421 gnd 0.006186f
C3119 vdd.n2422 gnd 0.006186f
C3120 vdd.n2423 gnd 0.006186f
C3121 vdd.n2424 gnd 0.006186f
C3122 vdd.n2425 gnd 0.006186f
C3123 vdd.n2426 gnd 0.006186f
C3124 vdd.n2427 gnd 0.006186f
C3125 vdd.n2428 gnd 0.006186f
C3126 vdd.n2429 gnd 0.006186f
C3127 vdd.n2430 gnd 0.006186f
C3128 vdd.n2431 gnd 0.006186f
C3129 vdd.n2432 gnd 0.006186f
C3130 vdd.n2433 gnd 0.006186f
C3131 vdd.n2434 gnd 0.006186f
C3132 vdd.n2435 gnd 0.006186f
C3133 vdd.n2436 gnd 0.006186f
C3134 vdd.n2437 gnd 0.006186f
C3135 vdd.n2438 gnd 0.006186f
C3136 vdd.n2439 gnd 0.006186f
C3137 vdd.n2440 gnd 0.006186f
C3138 vdd.n2441 gnd 0.006186f
C3139 vdd.n2442 gnd 0.006186f
C3140 vdd.n2443 gnd 0.006186f
C3141 vdd.n2444 gnd 0.006186f
C3142 vdd.n2445 gnd 0.006186f
C3143 vdd.n2446 gnd 0.006186f
C3144 vdd.n2447 gnd 0.006186f
C3145 vdd.n2448 gnd 0.006186f
C3146 vdd.n2449 gnd 0.006186f
C3147 vdd.n2450 gnd 0.006186f
C3148 vdd.n2451 gnd 0.006186f
C3149 vdd.n2452 gnd 0.006186f
C3150 vdd.n2453 gnd 0.006186f
C3151 vdd.n2454 gnd 0.006186f
C3152 vdd.n2455 gnd 0.006186f
C3153 vdd.n2456 gnd 0.006186f
C3154 vdd.n2457 gnd 0.006186f
C3155 vdd.n2458 gnd 0.006186f
C3156 vdd.n2459 gnd 0.006186f
C3157 vdd.n2460 gnd 0.006186f
C3158 vdd.n2461 gnd 0.006186f
C3159 vdd.n2462 gnd 0.006186f
C3160 vdd.n2463 gnd 0.006186f
C3161 vdd.n2464 gnd 0.006186f
C3162 vdd.n2465 gnd 0.006186f
C3163 vdd.n2466 gnd 0.006186f
C3164 vdd.n2467 gnd 0.006186f
C3165 vdd.n2468 gnd 0.006186f
C3166 vdd.n2469 gnd 0.006186f
C3167 vdd.n2471 gnd 0.771597f
C3168 vdd.n2473 gnd 0.006186f
C3169 vdd.n2474 gnd 0.006186f
C3170 vdd.n2475 gnd 0.014678f
C3171 vdd.n2476 gnd 0.013704f
C3172 vdd.n2477 gnd 0.013704f
C3173 vdd.n2478 gnd 0.771597f
C3174 vdd.n2479 gnd 0.013704f
C3175 vdd.n2480 gnd 0.013704f
C3176 vdd.n2481 gnd 0.006186f
C3177 vdd.n2482 gnd 0.006186f
C3178 vdd.n2483 gnd 0.006186f
C3179 vdd.n2484 gnd 0.395095f
C3180 vdd.n2485 gnd 0.006186f
C3181 vdd.n2486 gnd 0.006186f
C3182 vdd.n2487 gnd 0.006186f
C3183 vdd.n2488 gnd 0.006186f
C3184 vdd.n2489 gnd 0.006186f
C3185 vdd.n2490 gnd 0.492706f
C3186 vdd.n2491 gnd 0.006186f
C3187 vdd.n2492 gnd 0.006186f
C3188 vdd.n2493 gnd 0.006186f
C3189 vdd.n2494 gnd 0.006186f
C3190 vdd.n2495 gnd 0.006186f
C3191 vdd.n2496 gnd 0.632151f
C3192 vdd.n2497 gnd 0.006186f
C3193 vdd.n2498 gnd 0.006186f
C3194 vdd.n2499 gnd 0.006186f
C3195 vdd.n2500 gnd 0.006186f
C3196 vdd.n2501 gnd 0.006186f
C3197 vdd.n2502 gnd 0.348613f
C3198 vdd.n2503 gnd 0.006186f
C3199 vdd.n2504 gnd 0.006186f
C3200 vdd.n2505 gnd 0.006186f
C3201 vdd.n2506 gnd 0.006186f
C3202 vdd.n2507 gnd 0.006186f
C3203 vdd.n2508 gnd 0.199871f
C3204 vdd.n2509 gnd 0.006186f
C3205 vdd.n2510 gnd 0.006186f
C3206 vdd.n2511 gnd 0.006186f
C3207 vdd.n2512 gnd 0.006186f
C3208 vdd.n2513 gnd 0.006186f
C3209 vdd.n2514 gnd 0.362557f
C3210 vdd.n2515 gnd 0.006186f
C3211 vdd.n2516 gnd 0.006186f
C3212 vdd.n2517 gnd 0.006186f
C3213 vdd.n2518 gnd 0.006186f
C3214 vdd.n2519 gnd 0.006186f
C3215 vdd.n2520 gnd 0.502003f
C3216 vdd.n2521 gnd 0.006186f
C3217 vdd.n2522 gnd 0.006186f
C3218 vdd.n2523 gnd 0.006186f
C3219 vdd.n2524 gnd 0.006186f
C3220 vdd.n2525 gnd 0.006186f
C3221 vdd.n2526 gnd 0.562429f
C3222 vdd.n2527 gnd 0.006186f
C3223 vdd.n2528 gnd 0.006186f
C3224 vdd.n2529 gnd 0.006186f
C3225 vdd.n2530 gnd 0.006186f
C3226 vdd.n2531 gnd 0.006186f
C3227 vdd.n2532 gnd 0.422984f
C3228 vdd.n2533 gnd 0.006186f
C3229 vdd.n2534 gnd 0.006186f
C3230 vdd.n2535 gnd 0.006186f
C3231 vdd.t98 gnd 0.255869f
C3232 vdd.t96 gnd 0.163186f
C3233 vdd.t99 gnd 0.255869f
C3234 vdd.n2536 gnd 0.143809f
C3235 vdd.n2537 gnd 0.017919f
C3236 vdd.n2538 gnd 0.003821f
C3237 vdd.n2539 gnd 0.006186f
C3238 vdd.n2540 gnd 0.348613f
C3239 vdd.n2541 gnd 0.006186f
C3240 vdd.n2542 gnd 0.006186f
C3241 vdd.n2543 gnd 0.006186f
C3242 vdd.n2544 gnd 0.006186f
C3243 vdd.n2545 gnd 0.006186f
C3244 vdd.n2546 gnd 0.632151f
C3245 vdd.n2547 gnd 0.006186f
C3246 vdd.n2548 gnd 0.006186f
C3247 vdd.n2549 gnd 0.006186f
C3248 vdd.n2550 gnd 0.006186f
C3249 vdd.n2551 gnd 0.006186f
C3250 vdd.n2552 gnd 0.006186f
C3251 vdd.n2554 gnd 0.006186f
C3252 vdd.n2555 gnd 0.006186f
C3253 vdd.n2557 gnd 0.006186f
C3254 vdd.n2558 gnd 0.006186f
C3255 vdd.n2561 gnd 0.006186f
C3256 vdd.n2562 gnd 0.006186f
C3257 vdd.n2563 gnd 0.006186f
C3258 vdd.n2564 gnd 0.006186f
C3259 vdd.n2566 gnd 0.006186f
C3260 vdd.n2567 gnd 0.006186f
C3261 vdd.n2568 gnd 0.006186f
C3262 vdd.n2569 gnd 0.006186f
C3263 vdd.n2570 gnd 0.006186f
C3264 vdd.n2571 gnd 0.006186f
C3265 vdd.n2573 gnd 0.006186f
C3266 vdd.n2574 gnd 0.006186f
C3267 vdd.n2575 gnd 0.006186f
C3268 vdd.n2576 gnd 0.006186f
C3269 vdd.n2577 gnd 0.006186f
C3270 vdd.n2578 gnd 0.006186f
C3271 vdd.n2580 gnd 0.006186f
C3272 vdd.n2581 gnd 0.006186f
C3273 vdd.n2582 gnd 0.006186f
C3274 vdd.n2583 gnd 0.006186f
C3275 vdd.n2584 gnd 0.006186f
C3276 vdd.n2585 gnd 0.006186f
C3277 vdd.n2587 gnd 0.006186f
C3278 vdd.n2588 gnd 0.014678f
C3279 vdd.n2589 gnd 0.014678f
C3280 vdd.n2590 gnd 0.013704f
C3281 vdd.n2591 gnd 0.006186f
C3282 vdd.n2592 gnd 0.006186f
C3283 vdd.n2593 gnd 0.006186f
C3284 vdd.n2594 gnd 0.006186f
C3285 vdd.n2595 gnd 0.006186f
C3286 vdd.n2596 gnd 0.006186f
C3287 vdd.n2597 gnd 0.632151f
C3288 vdd.n2598 gnd 0.006186f
C3289 vdd.n2599 gnd 0.006186f
C3290 vdd.n2600 gnd 0.006186f
C3291 vdd.n2601 gnd 0.006186f
C3292 vdd.n2602 gnd 0.006186f
C3293 vdd.n2603 gnd 0.395095f
C3294 vdd.n2604 gnd 0.006186f
C3295 vdd.n2605 gnd 0.006186f
C3296 vdd.n2606 gnd 0.006186f
C3297 vdd.n2607 gnd 0.014457f
C3298 vdd.n2608 gnd 0.013924f
C3299 vdd.n2609 gnd 0.014678f
C3300 vdd.n2611 gnd 0.006186f
C3301 vdd.n2612 gnd 0.006186f
C3302 vdd.n2613 gnd 0.004776f
C3303 vdd.n2614 gnd 0.00884f
C3304 vdd.n2615 gnd 0.004503f
C3305 vdd.n2616 gnd 0.006186f
C3306 vdd.n2617 gnd 0.006186f
C3307 vdd.n2619 gnd 0.006186f
C3308 vdd.n2620 gnd 0.006186f
C3309 vdd.n2621 gnd 0.006186f
C3310 vdd.n2622 gnd 0.006186f
C3311 vdd.n2623 gnd 0.006186f
C3312 vdd.n2624 gnd 0.006186f
C3313 vdd.n2626 gnd 0.006186f
C3314 vdd.n2627 gnd 0.006186f
C3315 vdd.n2628 gnd 0.006186f
C3316 vdd.n2629 gnd 0.006186f
C3317 vdd.n2630 gnd 0.006186f
C3318 vdd.n2631 gnd 0.006186f
C3319 vdd.n2633 gnd 0.006186f
C3320 vdd.n2634 gnd 0.006186f
C3321 vdd.n2635 gnd 0.006186f
C3322 vdd.n2636 gnd 0.006186f
C3323 vdd.n2637 gnd 0.006186f
C3324 vdd.n2638 gnd 0.006186f
C3325 vdd.n2640 gnd 0.006186f
C3326 vdd.n2641 gnd 0.006186f
C3327 vdd.n2642 gnd 0.006186f
C3328 vdd.n2644 gnd 0.006186f
C3329 vdd.n2645 gnd 0.006186f
C3330 vdd.n2646 gnd 0.006186f
C3331 vdd.n2647 gnd 0.006186f
C3332 vdd.n2648 gnd 0.006186f
C3333 vdd.n2649 gnd 0.006186f
C3334 vdd.n2651 gnd 0.006186f
C3335 vdd.n2652 gnd 0.006186f
C3336 vdd.n2653 gnd 0.006186f
C3337 vdd.n2654 gnd 0.006186f
C3338 vdd.n2655 gnd 0.006186f
C3339 vdd.n2656 gnd 0.006186f
C3340 vdd.n2658 gnd 0.006186f
C3341 vdd.n2659 gnd 0.006186f
C3342 vdd.n2660 gnd 0.006186f
C3343 vdd.n2661 gnd 0.006186f
C3344 vdd.n2662 gnd 0.006186f
C3345 vdd.n2663 gnd 0.006186f
C3346 vdd.n2665 gnd 0.006186f
C3347 vdd.n2666 gnd 0.006186f
C3348 vdd.n2668 gnd 0.006186f
C3349 vdd.n2669 gnd 0.006186f
C3350 vdd.n2670 gnd 0.014678f
C3351 vdd.n2671 gnd 0.013704f
C3352 vdd.n2672 gnd 0.013704f
C3353 vdd.n2673 gnd 0.911042f
C3354 vdd.n2674 gnd 0.013704f
C3355 vdd.n2675 gnd 0.014678f
C3356 vdd.n2676 gnd 0.013924f
C3357 vdd.n2677 gnd 0.006186f
C3358 vdd.n2678 gnd 0.004776f
C3359 vdd.n2679 gnd 0.006186f
C3360 vdd.n2681 gnd 0.006186f
C3361 vdd.n2682 gnd 0.006186f
C3362 vdd.n2683 gnd 0.006186f
C3363 vdd.n2684 gnd 0.006186f
C3364 vdd.n2685 gnd 0.006186f
C3365 vdd.n2686 gnd 0.006186f
C3366 vdd.n2688 gnd 0.006186f
C3367 vdd.n2689 gnd 0.006186f
C3368 vdd.n2690 gnd 0.006186f
C3369 vdd.n2691 gnd 0.006186f
C3370 vdd.n2692 gnd 0.006186f
C3371 vdd.n2693 gnd 0.006186f
C3372 vdd.n2695 gnd 0.006186f
C3373 vdd.n2696 gnd 0.006186f
C3374 vdd.n2697 gnd 0.006186f
C3375 vdd.n2698 gnd 0.006186f
C3376 vdd.n2699 gnd 0.006186f
C3377 vdd.n2700 gnd 0.006186f
C3378 vdd.n2702 gnd 0.006186f
C3379 vdd.n2703 gnd 0.006186f
C3380 vdd.n2705 gnd 0.006186f
C3381 vdd.n2706 gnd 0.014864f
C3382 vdd.n2707 gnd 0.550544f
C3383 vdd.n2708 gnd 0.007823f
C3384 vdd.n2709 gnd 0.022678f
C3385 vdd.n2710 gnd 0.003478f
C3386 vdd.t149 gnd 0.111913f
C3387 vdd.t150 gnd 0.119604f
C3388 vdd.t148 gnd 0.146157f
C3389 vdd.n2711 gnd 0.187352f
C3390 vdd.n2712 gnd 0.15741f
C3391 vdd.n2713 gnd 0.011275f
C3392 vdd.n2714 gnd 0.009097f
C3393 vdd.n2715 gnd 0.003844f
C3394 vdd.n2716 gnd 0.007322f
C3395 vdd.n2717 gnd 0.009097f
C3396 vdd.n2718 gnd 0.009097f
C3397 vdd.n2719 gnd 0.007322f
C3398 vdd.n2720 gnd 0.007322f
C3399 vdd.n2721 gnd 0.009097f
C3400 vdd.n2722 gnd 0.009097f
C3401 vdd.n2723 gnd 0.007322f
C3402 vdd.n2724 gnd 0.007322f
C3403 vdd.n2725 gnd 0.009097f
C3404 vdd.n2726 gnd 0.009097f
C3405 vdd.n2727 gnd 0.007322f
C3406 vdd.n2728 gnd 0.007322f
C3407 vdd.n2729 gnd 0.009097f
C3408 vdd.n2730 gnd 0.009097f
C3409 vdd.n2731 gnd 0.007322f
C3410 vdd.n2732 gnd 0.007322f
C3411 vdd.n2733 gnd 0.009097f
C3412 vdd.n2734 gnd 0.009097f
C3413 vdd.n2735 gnd 0.007322f
C3414 vdd.n2736 gnd 0.007322f
C3415 vdd.n2737 gnd 0.009097f
C3416 vdd.n2738 gnd 0.009097f
C3417 vdd.n2739 gnd 0.007322f
C3418 vdd.n2740 gnd 0.007322f
C3419 vdd.n2741 gnd 0.009097f
C3420 vdd.n2742 gnd 0.009097f
C3421 vdd.n2743 gnd 0.007322f
C3422 vdd.n2744 gnd 0.007322f
C3423 vdd.n2745 gnd 0.009097f
C3424 vdd.n2746 gnd 0.009097f
C3425 vdd.n2747 gnd 0.007322f
C3426 vdd.n2748 gnd 0.007322f
C3427 vdd.n2749 gnd 0.009097f
C3428 vdd.n2750 gnd 0.009097f
C3429 vdd.n2751 gnd 0.007322f
C3430 vdd.n2752 gnd 0.009097f
C3431 vdd.n2753 gnd 0.009097f
C3432 vdd.n2754 gnd 0.007322f
C3433 vdd.n2755 gnd 0.009097f
C3434 vdd.n2756 gnd 0.009097f
C3435 vdd.n2757 gnd 0.009097f
C3436 vdd.n2758 gnd 0.014936f
C3437 vdd.n2759 gnd 0.009097f
C3438 vdd.n2760 gnd 0.009097f
C3439 vdd.n2761 gnd 0.004979f
C3440 vdd.n2762 gnd 0.007322f
C3441 vdd.n2763 gnd 0.009097f
C3442 vdd.n2764 gnd 0.009097f
C3443 vdd.n2765 gnd 0.007322f
C3444 vdd.n2766 gnd 0.007322f
C3445 vdd.n2767 gnd 0.009097f
C3446 vdd.n2768 gnd 0.009097f
C3447 vdd.n2769 gnd 0.007322f
C3448 vdd.n2770 gnd 0.007322f
C3449 vdd.n2771 gnd 0.009097f
C3450 vdd.n2772 gnd 0.009097f
C3451 vdd.n2773 gnd 0.007322f
C3452 vdd.n2774 gnd 0.007322f
C3453 vdd.n2775 gnd 0.009097f
C3454 vdd.n2776 gnd 0.009097f
C3455 vdd.n2777 gnd 0.007322f
C3456 vdd.n2778 gnd 0.007322f
C3457 vdd.n2779 gnd 0.009097f
C3458 vdd.n2780 gnd 0.009097f
C3459 vdd.n2781 gnd 0.007322f
C3460 vdd.n2782 gnd 0.007322f
C3461 vdd.n2783 gnd 0.009097f
C3462 vdd.n2784 gnd 0.009097f
C3463 vdd.n2785 gnd 0.007322f
C3464 vdd.n2786 gnd 0.007322f
C3465 vdd.n2787 gnd 0.009097f
C3466 vdd.n2788 gnd 0.009097f
C3467 vdd.n2789 gnd 0.007322f
C3468 vdd.n2790 gnd 0.007322f
C3469 vdd.n2791 gnd 0.009097f
C3470 vdd.n2792 gnd 0.009097f
C3471 vdd.n2793 gnd 0.007322f
C3472 vdd.n2794 gnd 0.007322f
C3473 vdd.n2795 gnd 0.009097f
C3474 vdd.n2796 gnd 0.009097f
C3475 vdd.n2797 gnd 0.007322f
C3476 vdd.n2798 gnd 0.009097f
C3477 vdd.n2799 gnd 0.009097f
C3478 vdd.n2800 gnd 0.007322f
C3479 vdd.n2801 gnd 0.009097f
C3480 vdd.n2802 gnd 0.009097f
C3481 vdd.n2803 gnd 0.009097f
C3482 vdd.t86 gnd 0.111913f
C3483 vdd.t87 gnd 0.119604f
C3484 vdd.t85 gnd 0.146157f
C3485 vdd.n2804 gnd 0.187352f
C3486 vdd.n2805 gnd 0.15741f
C3487 vdd.n2806 gnd 0.014936f
C3488 vdd.n2807 gnd 0.009097f
C3489 vdd.n2808 gnd 0.009097f
C3490 vdd.n2809 gnd 0.006114f
C3491 vdd.n2810 gnd 0.007322f
C3492 vdd.n2811 gnd 0.009097f
C3493 vdd.n2812 gnd 0.009097f
C3494 vdd.n2813 gnd 0.007322f
C3495 vdd.n2814 gnd 0.007322f
C3496 vdd.n2815 gnd 0.009097f
C3497 vdd.n2816 gnd 0.009097f
C3498 vdd.n2817 gnd 0.007322f
C3499 vdd.n2818 gnd 0.007322f
C3500 vdd.n2819 gnd 0.009097f
C3501 vdd.n2820 gnd 0.009097f
C3502 vdd.n2821 gnd 0.007322f
C3503 vdd.n2822 gnd 0.007322f
C3504 vdd.n2823 gnd 0.009097f
C3505 vdd.n2824 gnd 0.009097f
C3506 vdd.n2825 gnd 0.007322f
C3507 vdd.n2826 gnd 0.007322f
C3508 vdd.n2827 gnd 0.009097f
C3509 vdd.n2828 gnd 0.009097f
C3510 vdd.n2829 gnd 0.007322f
C3511 vdd.n2830 gnd 0.007322f
C3512 vdd.n2831 gnd 0.009097f
C3513 vdd.n2832 gnd 0.009097f
C3514 vdd.n2833 gnd 0.007322f
C3515 vdd.n2834 gnd 0.007322f
C3516 vdd.n2836 gnd 0.550544f
C3517 vdd.n2838 gnd 0.007322f
C3518 vdd.n2839 gnd 0.009097f
C3519 vdd.n2840 gnd 6.73985f
C3520 vdd.n2842 gnd 0.022678f
C3521 vdd.n2843 gnd 0.006077f
C3522 vdd.n2844 gnd 0.022678f
C3523 vdd.n2845 gnd 0.022169f
C3524 vdd.n2846 gnd 0.009097f
C3525 vdd.n2847 gnd 0.007322f
C3526 vdd.n2848 gnd 0.009097f
C3527 vdd.n2849 gnd 0.581022f
C3528 vdd.n2850 gnd 0.009097f
C3529 vdd.n2851 gnd 0.007322f
C3530 vdd.n2852 gnd 0.009097f
C3531 vdd.n2853 gnd 0.009097f
C3532 vdd.n2854 gnd 0.009097f
C3533 vdd.n2855 gnd 0.007322f
C3534 vdd.n2856 gnd 0.009097f
C3535 vdd.n2857 gnd 0.739059f
C3536 vdd.n2858 gnd 0.929634f
C3537 vdd.n2859 gnd 0.009097f
C3538 vdd.n2860 gnd 0.007322f
C3539 vdd.n2861 gnd 0.009097f
C3540 vdd.n2862 gnd 0.009097f
C3541 vdd.n2863 gnd 0.009097f
C3542 vdd.n2864 gnd 0.007322f
C3543 vdd.n2865 gnd 0.009097f
C3544 vdd.n2866 gnd 0.655392f
C3545 vdd.n2867 gnd 0.009097f
C3546 vdd.n2868 gnd 0.007322f
C3547 vdd.n2869 gnd 0.009097f
C3548 vdd.n2870 gnd 0.009097f
C3549 vdd.n2871 gnd 0.009097f
C3550 vdd.n2872 gnd 0.007322f
C3551 vdd.n2873 gnd 0.009097f
C3552 vdd.t38 gnd 0.464817f
C3553 vdd.n2874 gnd 0.771597f
C3554 vdd.n2875 gnd 0.009097f
C3555 vdd.n2876 gnd 0.007322f
C3556 vdd.n2877 gnd 0.009097f
C3557 vdd.n2878 gnd 0.009097f
C3558 vdd.n2879 gnd 0.009097f
C3559 vdd.n2880 gnd 0.007322f
C3560 vdd.n2881 gnd 0.009097f
C3561 vdd.n2882 gnd 0.729763f
C3562 vdd.n2883 gnd 0.009097f
C3563 vdd.n2884 gnd 0.007322f
C3564 vdd.n2885 gnd 0.009097f
C3565 vdd.n2886 gnd 0.009097f
C3566 vdd.n2887 gnd 0.009097f
C3567 vdd.n2888 gnd 0.007322f
C3568 vdd.n2889 gnd 0.007322f
C3569 vdd.n2890 gnd 0.007322f
C3570 vdd.n2891 gnd 0.009097f
C3571 vdd.n2892 gnd 0.009097f
C3572 vdd.n2893 gnd 0.009097f
C3573 vdd.n2894 gnd 0.007322f
C3574 vdd.n2895 gnd 0.007322f
C3575 vdd.n2896 gnd 0.007322f
C3576 vdd.n2897 gnd 0.009097f
C3577 vdd.n2898 gnd 0.009097f
C3578 vdd.n2899 gnd 0.009097f
C3579 vdd.n2900 gnd 0.007322f
C3580 vdd.n2901 gnd 0.007322f
C3581 vdd.n2902 gnd 0.006077f
C3582 vdd.n2903 gnd 0.022169f
C3583 vdd.n2904 gnd 0.022678f
C3584 vdd.n2906 gnd 0.022678f
C3585 vdd.n2907 gnd 0.003478f
C3586 vdd.t153 gnd 0.111913f
C3587 vdd.t152 gnd 0.119604f
C3588 vdd.t151 gnd 0.146157f
C3589 vdd.n2908 gnd 0.187352f
C3590 vdd.n2909 gnd 0.158142f
C3591 vdd.n2910 gnd 0.012008f
C3592 vdd.n2911 gnd 0.003844f
C3593 vdd.n2912 gnd 0.007322f
C3594 vdd.n2913 gnd 0.009097f
C3595 vdd.n2915 gnd 0.009097f
C3596 vdd.n2916 gnd 0.009097f
C3597 vdd.n2917 gnd 0.007322f
C3598 vdd.n2918 gnd 0.007322f
C3599 vdd.n2919 gnd 0.007322f
C3600 vdd.n2920 gnd 0.009097f
C3601 vdd.n2922 gnd 0.009097f
C3602 vdd.n2923 gnd 0.009097f
C3603 vdd.n2924 gnd 0.007322f
C3604 vdd.n2925 gnd 0.007322f
C3605 vdd.n2926 gnd 0.007322f
C3606 vdd.n2927 gnd 0.009097f
C3607 vdd.n2929 gnd 0.009097f
C3608 vdd.n2930 gnd 0.009097f
C3609 vdd.n2931 gnd 0.007322f
C3610 vdd.n2932 gnd 0.007322f
C3611 vdd.n2933 gnd 0.007322f
C3612 vdd.n2934 gnd 0.009097f
C3613 vdd.n2936 gnd 0.009097f
C3614 vdd.n2937 gnd 0.009097f
C3615 vdd.n2938 gnd 0.007322f
C3616 vdd.n2939 gnd 0.007322f
C3617 vdd.n2940 gnd 0.007322f
C3618 vdd.n2941 gnd 0.009097f
C3619 vdd.n2943 gnd 0.009097f
C3620 vdd.n2944 gnd 0.009097f
C3621 vdd.n2945 gnd 0.007322f
C3622 vdd.n2946 gnd 0.009097f
C3623 vdd.n2947 gnd 0.009097f
C3624 vdd.n2948 gnd 0.009097f
C3625 vdd.n2949 gnd 0.015668f
C3626 vdd.n2950 gnd 0.004979f
C3627 vdd.n2951 gnd 0.007322f
C3628 vdd.n2952 gnd 0.009097f
C3629 vdd.n2954 gnd 0.009097f
C3630 vdd.n2955 gnd 0.009097f
C3631 vdd.n2956 gnd 0.007322f
C3632 vdd.n2957 gnd 0.007322f
C3633 vdd.n2958 gnd 0.007322f
C3634 vdd.n2959 gnd 0.009097f
C3635 vdd.n2961 gnd 0.009097f
C3636 vdd.n2962 gnd 0.009097f
C3637 vdd.n2963 gnd 0.007322f
C3638 vdd.n2964 gnd 0.007322f
C3639 vdd.n2965 gnd 0.007322f
C3640 vdd.n2966 gnd 0.009097f
C3641 vdd.n2968 gnd 0.009097f
C3642 vdd.n2969 gnd 0.009097f
C3643 vdd.n2970 gnd 0.007322f
C3644 vdd.n2971 gnd 0.007322f
C3645 vdd.n2972 gnd 0.007322f
C3646 vdd.n2973 gnd 0.009097f
C3647 vdd.n2975 gnd 0.009097f
C3648 vdd.n2976 gnd 0.009097f
C3649 vdd.n2977 gnd 0.007322f
C3650 vdd.n2978 gnd 0.007322f
C3651 vdd.n2979 gnd 0.007322f
C3652 vdd.n2980 gnd 0.009097f
C3653 vdd.n2982 gnd 0.009097f
C3654 vdd.n2983 gnd 0.009097f
C3655 vdd.n2984 gnd 0.007322f
C3656 vdd.n2985 gnd 0.009097f
C3657 vdd.n2986 gnd 0.009097f
C3658 vdd.n2987 gnd 0.009097f
C3659 vdd.n2988 gnd 0.015668f
C3660 vdd.n2989 gnd 0.006114f
C3661 vdd.n2990 gnd 0.007322f
C3662 vdd.n2991 gnd 0.009097f
C3663 vdd.n2993 gnd 0.009097f
C3664 vdd.n2994 gnd 0.009097f
C3665 vdd.n2995 gnd 0.007322f
C3666 vdd.n2996 gnd 0.007322f
C3667 vdd.n2997 gnd 0.007322f
C3668 vdd.n2998 gnd 0.009097f
C3669 vdd.n3000 gnd 0.009097f
C3670 vdd.n3001 gnd 0.009097f
C3671 vdd.n3002 gnd 0.007322f
C3672 vdd.n3003 gnd 0.007322f
C3673 vdd.n3004 gnd 0.007322f
C3674 vdd.n3005 gnd 0.009097f
C3675 vdd.n3007 gnd 0.009097f
C3676 vdd.n3008 gnd 0.009097f
C3677 vdd.n3009 gnd 0.007322f
C3678 vdd.n3010 gnd 0.007322f
C3679 vdd.n3011 gnd 0.007322f
C3680 vdd.n3012 gnd 0.009097f
C3681 vdd.n3014 gnd 0.009097f
C3682 vdd.n3015 gnd 0.009097f
C3683 vdd.n3017 gnd 0.009097f
C3684 vdd.n3018 gnd 0.007322f
C3685 vdd.n3019 gnd 0.007322f
C3686 vdd.n3020 gnd 0.006077f
C3687 vdd.n3021 gnd 0.022678f
C3688 vdd.n3022 gnd 0.022169f
C3689 vdd.n3023 gnd 0.006077f
C3690 vdd.n3024 gnd 0.022169f
C3691 vdd.n3025 gnd 1.37121f
C3692 vdd.t104 gnd 0.464817f
C3693 vdd.n3026 gnd 0.488058f
C3694 vdd.n3027 gnd 0.929634f
C3695 vdd.n3028 gnd 0.009097f
C3696 vdd.n3029 gnd 0.007322f
C3697 vdd.n3030 gnd 0.007322f
C3698 vdd.n3031 gnd 0.007322f
C3699 vdd.n3032 gnd 0.009097f
C3700 vdd.n3033 gnd 0.832023f
C3701 vdd.t29 gnd 0.464817f
C3702 vdd.n3034 gnd 0.562429f
C3703 vdd.n3035 gnd 0.673985f
C3704 vdd.n3036 gnd 0.009097f
C3705 vdd.n3037 gnd 0.007322f
C3706 vdd.n3038 gnd 0.007322f
C3707 vdd.n3039 gnd 0.007322f
C3708 vdd.n3040 gnd 0.009097f
C3709 vdd.n3041 gnd 0.515947f
C3710 vdd.t51 gnd 0.464817f
C3711 vdd.n3042 gnd 0.771597f
C3712 vdd.t27 gnd 0.464817f
C3713 vdd.n3043 gnd 0.571725f
C3714 vdd.n3044 gnd 0.009097f
C3715 vdd.n3045 gnd 0.007322f
C3716 vdd.n3046 gnd 0.006991f
C3717 vdd.n3047 gnd 0.536555f
C3718 vdd.n3048 gnd 1.84238f
C3719 CSoutput.n0 gnd 0.037112f
C3720 CSoutput.t120 gnd 0.245489f
C3721 CSoutput.n1 gnd 0.11085f
C3722 CSoutput.n2 gnd 0.037112f
C3723 CSoutput.t125 gnd 0.245489f
C3724 CSoutput.n3 gnd 0.029414f
C3725 CSoutput.n4 gnd 0.037112f
C3726 CSoutput.t134 gnd 0.245489f
C3727 CSoutput.n5 gnd 0.025364f
C3728 CSoutput.n6 gnd 0.037112f
C3729 CSoutput.t123 gnd 0.245489f
C3730 CSoutput.t127 gnd 0.245489f
C3731 CSoutput.n7 gnd 0.109642f
C3732 CSoutput.n8 gnd 0.037112f
C3733 CSoutput.t133 gnd 0.245489f
C3734 CSoutput.n9 gnd 0.024183f
C3735 CSoutput.n10 gnd 0.037112f
C3736 CSoutput.t136 gnd 0.245489f
C3737 CSoutput.t124 gnd 0.245489f
C3738 CSoutput.n11 gnd 0.109642f
C3739 CSoutput.n12 gnd 0.037112f
C3740 CSoutput.t130 gnd 0.245489f
C3741 CSoutput.n13 gnd 0.025364f
C3742 CSoutput.n14 gnd 0.037112f
C3743 CSoutput.t129 gnd 0.245489f
C3744 CSoutput.t139 gnd 0.245489f
C3745 CSoutput.n15 gnd 0.109642f
C3746 CSoutput.n16 gnd 0.037112f
C3747 CSoutput.t128 gnd 0.245489f
C3748 CSoutput.n17 gnd 0.02709f
C3749 CSoutput.t137 gnd 0.293365f
C3750 CSoutput.t126 gnd 0.245489f
C3751 CSoutput.n18 gnd 0.13997f
C3752 CSoutput.n19 gnd 0.13582f
C3753 CSoutput.n20 gnd 0.157567f
C3754 CSoutput.n21 gnd 0.037112f
C3755 CSoutput.n22 gnd 0.030974f
C3756 CSoutput.n23 gnd 0.109642f
C3757 CSoutput.n24 gnd 0.029858f
C3758 CSoutput.n25 gnd 0.029414f
C3759 CSoutput.n26 gnd 0.037112f
C3760 CSoutput.n27 gnd 0.037112f
C3761 CSoutput.n28 gnd 0.030736f
C3762 CSoutput.n29 gnd 0.026096f
C3763 CSoutput.n30 gnd 0.112083f
C3764 CSoutput.n31 gnd 0.026455f
C3765 CSoutput.n32 gnd 0.037112f
C3766 CSoutput.n33 gnd 0.037112f
C3767 CSoutput.n34 gnd 0.037112f
C3768 CSoutput.n35 gnd 0.030409f
C3769 CSoutput.n36 gnd 0.109642f
C3770 CSoutput.n37 gnd 0.029081f
C3771 CSoutput.n38 gnd 0.030191f
C3772 CSoutput.n39 gnd 0.037112f
C3773 CSoutput.n40 gnd 0.037112f
C3774 CSoutput.n41 gnd 0.030968f
C3775 CSoutput.n42 gnd 0.028305f
C3776 CSoutput.n43 gnd 0.109642f
C3777 CSoutput.n44 gnd 0.029022f
C3778 CSoutput.n45 gnd 0.037112f
C3779 CSoutput.n46 gnd 0.037112f
C3780 CSoutput.n47 gnd 0.037112f
C3781 CSoutput.n48 gnd 0.029022f
C3782 CSoutput.n49 gnd 0.109642f
C3783 CSoutput.n50 gnd 0.028305f
C3784 CSoutput.n51 gnd 0.030968f
C3785 CSoutput.n52 gnd 0.037112f
C3786 CSoutput.n53 gnd 0.037112f
C3787 CSoutput.n54 gnd 0.030191f
C3788 CSoutput.n55 gnd 0.029081f
C3789 CSoutput.n56 gnd 0.109642f
C3790 CSoutput.n57 gnd 0.030409f
C3791 CSoutput.n58 gnd 0.037112f
C3792 CSoutput.n59 gnd 0.037112f
C3793 CSoutput.n60 gnd 0.037112f
C3794 CSoutput.n61 gnd 0.026455f
C3795 CSoutput.n62 gnd 0.112083f
C3796 CSoutput.n63 gnd 0.026096f
C3797 CSoutput.t135 gnd 0.245489f
C3798 CSoutput.n64 gnd 0.109642f
C3799 CSoutput.n65 gnd 0.030736f
C3800 CSoutput.n66 gnd 0.037112f
C3801 CSoutput.n67 gnd 0.037112f
C3802 CSoutput.n68 gnd 0.037112f
C3803 CSoutput.n69 gnd 0.029858f
C3804 CSoutput.n70 gnd 0.109642f
C3805 CSoutput.n71 gnd 0.030974f
C3806 CSoutput.n72 gnd 0.02709f
C3807 CSoutput.n73 gnd 0.037112f
C3808 CSoutput.n74 gnd 0.037112f
C3809 CSoutput.n75 gnd 0.028094f
C3810 CSoutput.n76 gnd 0.016685f
C3811 CSoutput.t138 gnd 0.275824f
C3812 CSoutput.n77 gnd 0.137018f
C3813 CSoutput.n78 gnd 0.560535f
C3814 CSoutput.t94 gnd 0.046292f
C3815 CSoutput.t74 gnd 0.046292f
C3816 CSoutput.n79 gnd 0.358409f
C3817 CSoutput.t111 gnd 0.046292f
C3818 CSoutput.t80 gnd 0.046292f
C3819 CSoutput.n80 gnd 0.35777f
C3820 CSoutput.n81 gnd 0.363136f
C3821 CSoutput.t99 gnd 0.046292f
C3822 CSoutput.t72 gnd 0.046292f
C3823 CSoutput.n82 gnd 0.35777f
C3824 CSoutput.n83 gnd 0.178938f
C3825 CSoutput.t116 gnd 0.046292f
C3826 CSoutput.t114 gnd 0.046292f
C3827 CSoutput.n84 gnd 0.35777f
C3828 CSoutput.n85 gnd 0.328131f
C3829 CSoutput.t92 gnd 0.046292f
C3830 CSoutput.t107 gnd 0.046292f
C3831 CSoutput.n86 gnd 0.358409f
C3832 CSoutput.t101 gnd 0.046292f
C3833 CSoutput.t82 gnd 0.046292f
C3834 CSoutput.n87 gnd 0.35777f
C3835 CSoutput.n88 gnd 0.363136f
C3836 CSoutput.t87 gnd 0.046292f
C3837 CSoutput.t98 gnd 0.046292f
C3838 CSoutput.n89 gnd 0.35777f
C3839 CSoutput.n90 gnd 0.178938f
C3840 CSoutput.t100 gnd 0.046292f
C3841 CSoutput.t86 gnd 0.046292f
C3842 CSoutput.n91 gnd 0.35777f
C3843 CSoutput.n92 gnd 0.266842f
C3844 CSoutput.n93 gnd 0.336486f
C3845 CSoutput.t77 gnd 0.046292f
C3846 CSoutput.t78 gnd 0.046292f
C3847 CSoutput.n94 gnd 0.358409f
C3848 CSoutput.t90 gnd 0.046292f
C3849 CSoutput.t88 gnd 0.046292f
C3850 CSoutput.n95 gnd 0.35777f
C3851 CSoutput.n96 gnd 0.363136f
C3852 CSoutput.t83 gnd 0.046292f
C3853 CSoutput.t76 gnd 0.046292f
C3854 CSoutput.n97 gnd 0.35777f
C3855 CSoutput.n98 gnd 0.178938f
C3856 CSoutput.t89 gnd 0.046292f
C3857 CSoutput.t103 gnd 0.046292f
C3858 CSoutput.n99 gnd 0.35777f
C3859 CSoutput.n100 gnd 0.266842f
C3860 CSoutput.n101 gnd 0.376105f
C3861 CSoutput.n102 gnd 6.72714f
C3862 CSoutput.n104 gnd 0.656506f
C3863 CSoutput.n105 gnd 0.49238f
C3864 CSoutput.n106 gnd 0.656506f
C3865 CSoutput.n107 gnd 0.656506f
C3866 CSoutput.n108 gnd 1.76752f
C3867 CSoutput.n109 gnd 0.656506f
C3868 CSoutput.n110 gnd 0.656506f
C3869 CSoutput.t131 gnd 0.820633f
C3870 CSoutput.n111 gnd 0.656506f
C3871 CSoutput.n112 gnd 0.656506f
C3872 CSoutput.n116 gnd 0.656506f
C3873 CSoutput.n120 gnd 0.656506f
C3874 CSoutput.n121 gnd 0.656506f
C3875 CSoutput.n123 gnd 0.656506f
C3876 CSoutput.n128 gnd 0.656506f
C3877 CSoutput.n130 gnd 0.656506f
C3878 CSoutput.n131 gnd 0.656506f
C3879 CSoutput.n133 gnd 0.656506f
C3880 CSoutput.n134 gnd 0.656506f
C3881 CSoutput.n136 gnd 0.656506f
C3882 CSoutput.t121 gnd 10.970099f
C3883 CSoutput.n138 gnd 0.656506f
C3884 CSoutput.n139 gnd 0.49238f
C3885 CSoutput.n140 gnd 0.656506f
C3886 CSoutput.n141 gnd 0.656506f
C3887 CSoutput.n142 gnd 1.76752f
C3888 CSoutput.n143 gnd 0.656506f
C3889 CSoutput.n144 gnd 0.656506f
C3890 CSoutput.t140 gnd 0.820633f
C3891 CSoutput.n145 gnd 0.656506f
C3892 CSoutput.n146 gnd 0.656506f
C3893 CSoutput.n150 gnd 0.656506f
C3894 CSoutput.n154 gnd 0.656506f
C3895 CSoutput.n155 gnd 0.656506f
C3896 CSoutput.n157 gnd 0.656506f
C3897 CSoutput.n162 gnd 0.656506f
C3898 CSoutput.n164 gnd 0.656506f
C3899 CSoutput.n165 gnd 0.656506f
C3900 CSoutput.n167 gnd 0.656506f
C3901 CSoutput.n168 gnd 0.656506f
C3902 CSoutput.n170 gnd 0.656506f
C3903 CSoutput.n171 gnd 0.49238f
C3904 CSoutput.n173 gnd 0.656506f
C3905 CSoutput.n174 gnd 0.49238f
C3906 CSoutput.n175 gnd 0.656506f
C3907 CSoutput.n176 gnd 0.656506f
C3908 CSoutput.n177 gnd 1.76752f
C3909 CSoutput.n178 gnd 0.656506f
C3910 CSoutput.n179 gnd 0.656506f
C3911 CSoutput.t132 gnd 0.820633f
C3912 CSoutput.n180 gnd 0.656506f
C3913 CSoutput.n181 gnd 1.76752f
C3914 CSoutput.n183 gnd 0.656506f
C3915 CSoutput.n184 gnd 0.656506f
C3916 CSoutput.n186 gnd 0.656506f
C3917 CSoutput.n187 gnd 0.656506f
C3918 CSoutput.t141 gnd 10.791401f
C3919 CSoutput.t122 gnd 10.970099f
C3920 CSoutput.n193 gnd 2.05956f
C3921 CSoutput.n194 gnd 8.38989f
C3922 CSoutput.n195 gnd 8.740951f
C3923 CSoutput.n200 gnd 2.23106f
C3924 CSoutput.n206 gnd 0.656506f
C3925 CSoutput.n208 gnd 0.656506f
C3926 CSoutput.n210 gnd 0.656506f
C3927 CSoutput.n212 gnd 0.656506f
C3928 CSoutput.n214 gnd 0.656506f
C3929 CSoutput.n220 gnd 0.656506f
C3930 CSoutput.n227 gnd 1.20444f
C3931 CSoutput.n228 gnd 1.20444f
C3932 CSoutput.n229 gnd 0.656506f
C3933 CSoutput.n230 gnd 0.656506f
C3934 CSoutput.n232 gnd 0.49238f
C3935 CSoutput.n233 gnd 0.421679f
C3936 CSoutput.n235 gnd 0.49238f
C3937 CSoutput.n236 gnd 0.421679f
C3938 CSoutput.n237 gnd 0.49238f
C3939 CSoutput.n239 gnd 0.656506f
C3940 CSoutput.n241 gnd 1.76752f
C3941 CSoutput.n242 gnd 2.05956f
C3942 CSoutput.n243 gnd 7.71654f
C3943 CSoutput.n245 gnd 0.49238f
C3944 CSoutput.n246 gnd 1.26692f
C3945 CSoutput.n247 gnd 0.49238f
C3946 CSoutput.n249 gnd 0.656506f
C3947 CSoutput.n251 gnd 1.76752f
C3948 CSoutput.n252 gnd 3.84994f
C3949 CSoutput.t81 gnd 0.046292f
C3950 CSoutput.t93 gnd 0.046292f
C3951 CSoutput.n253 gnd 0.358409f
C3952 CSoutput.t105 gnd 0.046292f
C3953 CSoutput.t118 gnd 0.046292f
C3954 CSoutput.n254 gnd 0.35777f
C3955 CSoutput.n255 gnd 0.363136f
C3956 CSoutput.t115 gnd 0.046292f
C3957 CSoutput.t97 gnd 0.046292f
C3958 CSoutput.n256 gnd 0.35777f
C3959 CSoutput.n257 gnd 0.178938f
C3960 CSoutput.t84 gnd 0.046292f
C3961 CSoutput.t117 gnd 0.046292f
C3962 CSoutput.n258 gnd 0.35777f
C3963 CSoutput.n259 gnd 0.328131f
C3964 CSoutput.t106 gnd 0.046292f
C3965 CSoutput.t102 gnd 0.046292f
C3966 CSoutput.n260 gnd 0.358409f
C3967 CSoutput.t110 gnd 0.046292f
C3968 CSoutput.t75 gnd 0.046292f
C3969 CSoutput.n261 gnd 0.35777f
C3970 CSoutput.n262 gnd 0.363136f
C3971 CSoutput.t79 gnd 0.046292f
C3972 CSoutput.t109 gnd 0.046292f
C3973 CSoutput.n263 gnd 0.35777f
C3974 CSoutput.n264 gnd 0.178938f
C3975 CSoutput.t119 gnd 0.046292f
C3976 CSoutput.t113 gnd 0.046292f
C3977 CSoutput.n265 gnd 0.35777f
C3978 CSoutput.n266 gnd 0.266842f
C3979 CSoutput.n267 gnd 0.336486f
C3980 CSoutput.t95 gnd 0.046292f
C3981 CSoutput.t96 gnd 0.046292f
C3982 CSoutput.n268 gnd 0.358409f
C3983 CSoutput.t108 gnd 0.046292f
C3984 CSoutput.t73 gnd 0.046292f
C3985 CSoutput.n269 gnd 0.35777f
C3986 CSoutput.n270 gnd 0.363136f
C3987 CSoutput.t104 gnd 0.046292f
C3988 CSoutput.t91 gnd 0.046292f
C3989 CSoutput.n271 gnd 0.35777f
C3990 CSoutput.n272 gnd 0.178938f
C3991 CSoutput.t112 gnd 0.046292f
C3992 CSoutput.t85 gnd 0.046292f
C3993 CSoutput.n273 gnd 0.357769f
C3994 CSoutput.n274 gnd 0.266843f
C3995 CSoutput.n275 gnd 0.376105f
C3996 CSoutput.n276 gnd 9.67674f
C3997 CSoutput.t63 gnd 0.040506f
C3998 CSoutput.t10 gnd 0.040506f
C3999 CSoutput.n277 gnd 0.35912f
C4000 CSoutput.t50 gnd 0.040506f
C4001 CSoutput.t0 gnd 0.040506f
C4002 CSoutput.n278 gnd 0.357922f
C4003 CSoutput.n279 gnd 0.333516f
C4004 CSoutput.t34 gnd 0.040506f
C4005 CSoutput.t65 gnd 0.040506f
C4006 CSoutput.n280 gnd 0.357922f
C4007 CSoutput.n281 gnd 0.164408f
C4008 CSoutput.t19 gnd 0.040506f
C4009 CSoutput.t32 gnd 0.040506f
C4010 CSoutput.n282 gnd 0.357922f
C4011 CSoutput.n283 gnd 0.164408f
C4012 CSoutput.t4 gnd 0.040506f
C4013 CSoutput.t40 gnd 0.040506f
C4014 CSoutput.n284 gnd 0.357922f
C4015 CSoutput.n285 gnd 0.164408f
C4016 CSoutput.t53 gnd 0.040506f
C4017 CSoutput.t24 gnd 0.040506f
C4018 CSoutput.n286 gnd 0.357922f
C4019 CSoutput.n287 gnd 0.303241f
C4020 CSoutput.t30 gnd 0.040506f
C4021 CSoutput.t13 gnd 0.040506f
C4022 CSoutput.n288 gnd 0.35912f
C4023 CSoutput.t18 gnd 0.040506f
C4024 CSoutput.t31 gnd 0.040506f
C4025 CSoutput.n289 gnd 0.357922f
C4026 CSoutput.n290 gnd 0.333516f
C4027 CSoutput.t14 gnd 0.040506f
C4028 CSoutput.t20 gnd 0.040506f
C4029 CSoutput.n291 gnd 0.357922f
C4030 CSoutput.n292 gnd 0.164408f
C4031 CSoutput.t33 gnd 0.040506f
C4032 CSoutput.t11 gnd 0.040506f
C4033 CSoutput.n293 gnd 0.357922f
C4034 CSoutput.n294 gnd 0.164408f
C4035 CSoutput.t21 gnd 0.040506f
C4036 CSoutput.t7 gnd 0.040506f
C4037 CSoutput.n295 gnd 0.357922f
C4038 CSoutput.n296 gnd 0.164408f
C4039 CSoutput.t12 gnd 0.040506f
C4040 CSoutput.t22 gnd 0.040506f
C4041 CSoutput.n297 gnd 0.357922f
C4042 CSoutput.n298 gnd 0.249606f
C4043 CSoutput.n299 gnd 0.314831f
C4044 CSoutput.t8 gnd 0.040506f
C4045 CSoutput.t69 gnd 0.040506f
C4046 CSoutput.n300 gnd 0.35912f
C4047 CSoutput.t59 gnd 0.040506f
C4048 CSoutput.t15 gnd 0.040506f
C4049 CSoutput.n301 gnd 0.357922f
C4050 CSoutput.n302 gnd 0.333516f
C4051 CSoutput.t1 gnd 0.040506f
C4052 CSoutput.t67 gnd 0.040506f
C4053 CSoutput.n303 gnd 0.357922f
C4054 CSoutput.n304 gnd 0.164408f
C4055 CSoutput.t26 gnd 0.040506f
C4056 CSoutput.t35 gnd 0.040506f
C4057 CSoutput.n305 gnd 0.357922f
C4058 CSoutput.n306 gnd 0.164408f
C4059 CSoutput.t70 gnd 0.040506f
C4060 CSoutput.t60 gnd 0.040506f
C4061 CSoutput.n307 gnd 0.357922f
C4062 CSoutput.n308 gnd 0.164408f
C4063 CSoutput.t44 gnd 0.040506f
C4064 CSoutput.t2 gnd 0.040506f
C4065 CSoutput.n309 gnd 0.357922f
C4066 CSoutput.n310 gnd 0.249606f
C4067 CSoutput.n311 gnd 0.338079f
C4068 CSoutput.n312 gnd 10.3251f
C4069 CSoutput.t41 gnd 0.040506f
C4070 CSoutput.t5 gnd 0.040506f
C4071 CSoutput.n313 gnd 0.35912f
C4072 CSoutput.t25 gnd 0.040506f
C4073 CSoutput.t66 gnd 0.040506f
C4074 CSoutput.n314 gnd 0.357922f
C4075 CSoutput.n315 gnd 0.333516f
C4076 CSoutput.t6 gnd 0.040506f
C4077 CSoutput.t55 gnd 0.040506f
C4078 CSoutput.n316 gnd 0.357922f
C4079 CSoutput.n317 gnd 0.164408f
C4080 CSoutput.t54 gnd 0.040506f
C4081 CSoutput.t43 gnd 0.040506f
C4082 CSoutput.n318 gnd 0.357922f
C4083 CSoutput.n319 gnd 0.164408f
C4084 CSoutput.t56 gnd 0.040506f
C4085 CSoutput.t27 gnd 0.040506f
C4086 CSoutput.n320 gnd 0.357922f
C4087 CSoutput.n321 gnd 0.164408f
C4088 CSoutput.t49 gnd 0.040506f
C4089 CSoutput.t61 gnd 0.040506f
C4090 CSoutput.n322 gnd 0.357922f
C4091 CSoutput.n323 gnd 0.303241f
C4092 CSoutput.t28 gnd 0.040506f
C4093 CSoutput.t45 gnd 0.040506f
C4094 CSoutput.n324 gnd 0.35912f
C4095 CSoutput.t46 gnd 0.040506f
C4096 CSoutput.t36 gnd 0.040506f
C4097 CSoutput.n325 gnd 0.357922f
C4098 CSoutput.n326 gnd 0.333516f
C4099 CSoutput.t37 gnd 0.040506f
C4100 CSoutput.t29 gnd 0.040506f
C4101 CSoutput.n327 gnd 0.357922f
C4102 CSoutput.n328 gnd 0.164408f
C4103 CSoutput.t23 gnd 0.040506f
C4104 CSoutput.t16 gnd 0.040506f
C4105 CSoutput.n329 gnd 0.357922f
C4106 CSoutput.n330 gnd 0.164408f
C4107 CSoutput.t17 gnd 0.040506f
C4108 CSoutput.t38 gnd 0.040506f
C4109 CSoutput.n331 gnd 0.357922f
C4110 CSoutput.n332 gnd 0.164408f
C4111 CSoutput.t39 gnd 0.040506f
C4112 CSoutput.t3 gnd 0.040506f
C4113 CSoutput.n333 gnd 0.357922f
C4114 CSoutput.n334 gnd 0.249606f
C4115 CSoutput.n335 gnd 0.314831f
C4116 CSoutput.t57 gnd 0.040506f
C4117 CSoutput.t68 gnd 0.040506f
C4118 CSoutput.n336 gnd 0.35912f
C4119 CSoutput.t71 gnd 0.040506f
C4120 CSoutput.t48 gnd 0.040506f
C4121 CSoutput.n337 gnd 0.357922f
C4122 CSoutput.n338 gnd 0.333516f
C4123 CSoutput.t52 gnd 0.040506f
C4124 CSoutput.t62 gnd 0.040506f
C4125 CSoutput.n339 gnd 0.357922f
C4126 CSoutput.n340 gnd 0.164408f
C4127 CSoutput.t9 gnd 0.040506f
C4128 CSoutput.t42 gnd 0.040506f
C4129 CSoutput.n341 gnd 0.357922f
C4130 CSoutput.n342 gnd 0.164408f
C4131 CSoutput.t47 gnd 0.040506f
C4132 CSoutput.t58 gnd 0.040506f
C4133 CSoutput.n343 gnd 0.357922f
C4134 CSoutput.n344 gnd 0.164408f
C4135 CSoutput.t64 gnd 0.040506f
C4136 CSoutput.t51 gnd 0.040506f
C4137 CSoutput.n345 gnd 0.357922f
C4138 CSoutput.n346 gnd 0.249606f
C4139 CSoutput.n347 gnd 0.338079f
C4140 CSoutput.n348 gnd 5.82483f
C4141 CSoutput.n349 gnd 11.4197f
C4142 commonsourceibias.n0 gnd 0.012299f
C4143 commonsourceibias.t56 gnd 0.18623f
C4144 commonsourceibias.t109 gnd 0.172196f
C4145 commonsourceibias.n1 gnd 0.068706f
C4146 commonsourceibias.n2 gnd 0.009217f
C4147 commonsourceibias.t69 gnd 0.172196f
C4148 commonsourceibias.n3 gnd 0.007456f
C4149 commonsourceibias.n4 gnd 0.009217f
C4150 commonsourceibias.t119 gnd 0.172196f
C4151 commonsourceibias.n5 gnd 0.008898f
C4152 commonsourceibias.n6 gnd 0.009217f
C4153 commonsourceibias.t85 gnd 0.172196f
C4154 commonsourceibias.n7 gnd 0.068706f
C4155 commonsourceibias.t54 gnd 0.172196f
C4156 commonsourceibias.n8 gnd 0.007444f
C4157 commonsourceibias.n9 gnd 0.012299f
C4158 commonsourceibias.t16 gnd 0.18623f
C4159 commonsourceibias.t30 gnd 0.172196f
C4160 commonsourceibias.n10 gnd 0.068706f
C4161 commonsourceibias.n11 gnd 0.009217f
C4162 commonsourceibias.t2 gnd 0.172196f
C4163 commonsourceibias.n12 gnd 0.007456f
C4164 commonsourceibias.n13 gnd 0.009217f
C4165 commonsourceibias.t22 gnd 0.172196f
C4166 commonsourceibias.n14 gnd 0.008898f
C4167 commonsourceibias.n15 gnd 0.009217f
C4168 commonsourceibias.t42 gnd 0.172196f
C4169 commonsourceibias.n16 gnd 0.068706f
C4170 commonsourceibias.t18 gnd 0.172196f
C4171 commonsourceibias.n17 gnd 0.007444f
C4172 commonsourceibias.n18 gnd 0.009217f
C4173 commonsourceibias.t32 gnd 0.172196f
C4174 commonsourceibias.t40 gnd 0.172196f
C4175 commonsourceibias.n19 gnd 0.068706f
C4176 commonsourceibias.n20 gnd 0.009217f
C4177 commonsourceibias.t24 gnd 0.172196f
C4178 commonsourceibias.n21 gnd 0.068706f
C4179 commonsourceibias.n22 gnd 0.009217f
C4180 commonsourceibias.t44 gnd 0.172196f
C4181 commonsourceibias.n23 gnd 0.068706f
C4182 commonsourceibias.n24 gnd 0.046399f
C4183 commonsourceibias.t6 gnd 0.172196f
C4184 commonsourceibias.t34 gnd 0.194303f
C4185 commonsourceibias.n25 gnd 0.079733f
C4186 commonsourceibias.n26 gnd 0.082545f
C4187 commonsourceibias.n27 gnd 0.01136f
C4188 commonsourceibias.n28 gnd 0.012567f
C4189 commonsourceibias.n29 gnd 0.009217f
C4190 commonsourceibias.n30 gnd 0.009217f
C4191 commonsourceibias.n31 gnd 0.012485f
C4192 commonsourceibias.n32 gnd 0.007456f
C4193 commonsourceibias.n33 gnd 0.01264f
C4194 commonsourceibias.n34 gnd 0.009217f
C4195 commonsourceibias.n35 gnd 0.009217f
C4196 commonsourceibias.n36 gnd 0.012717f
C4197 commonsourceibias.n37 gnd 0.010966f
C4198 commonsourceibias.n38 gnd 0.008898f
C4199 commonsourceibias.n39 gnd 0.009217f
C4200 commonsourceibias.n40 gnd 0.009217f
C4201 commonsourceibias.n41 gnd 0.011274f
C4202 commonsourceibias.n42 gnd 0.012653f
C4203 commonsourceibias.n43 gnd 0.068706f
C4204 commonsourceibias.n44 gnd 0.012568f
C4205 commonsourceibias.n45 gnd 0.009217f
C4206 commonsourceibias.n46 gnd 0.009217f
C4207 commonsourceibias.n47 gnd 0.009217f
C4208 commonsourceibias.n48 gnd 0.012568f
C4209 commonsourceibias.n49 gnd 0.068706f
C4210 commonsourceibias.n50 gnd 0.012653f
C4211 commonsourceibias.n51 gnd 0.011274f
C4212 commonsourceibias.n52 gnd 0.009217f
C4213 commonsourceibias.n53 gnd 0.009217f
C4214 commonsourceibias.n54 gnd 0.009217f
C4215 commonsourceibias.n55 gnd 0.010966f
C4216 commonsourceibias.n56 gnd 0.012717f
C4217 commonsourceibias.n57 gnd 0.068706f
C4218 commonsourceibias.n58 gnd 0.01264f
C4219 commonsourceibias.n59 gnd 0.009217f
C4220 commonsourceibias.n60 gnd 0.009217f
C4221 commonsourceibias.n61 gnd 0.009217f
C4222 commonsourceibias.n62 gnd 0.012485f
C4223 commonsourceibias.n63 gnd 0.068706f
C4224 commonsourceibias.n64 gnd 0.012567f
C4225 commonsourceibias.n65 gnd 0.01136f
C4226 commonsourceibias.n66 gnd 0.009217f
C4227 commonsourceibias.n67 gnd 0.009217f
C4228 commonsourceibias.n68 gnd 0.009349f
C4229 commonsourceibias.n69 gnd 0.009666f
C4230 commonsourceibias.n70 gnd 0.082208f
C4231 commonsourceibias.n71 gnd 0.091197f
C4232 commonsourceibias.t17 gnd 0.019889f
C4233 commonsourceibias.t31 gnd 0.019889f
C4234 commonsourceibias.n72 gnd 0.175743f
C4235 commonsourceibias.n73 gnd 0.151855f
C4236 commonsourceibias.t3 gnd 0.019889f
C4237 commonsourceibias.t23 gnd 0.019889f
C4238 commonsourceibias.n74 gnd 0.175743f
C4239 commonsourceibias.n75 gnd 0.080726f
C4240 commonsourceibias.t43 gnd 0.019889f
C4241 commonsourceibias.t19 gnd 0.019889f
C4242 commonsourceibias.n76 gnd 0.175743f
C4243 commonsourceibias.n77 gnd 0.067443f
C4244 commonsourceibias.t7 gnd 0.019889f
C4245 commonsourceibias.t35 gnd 0.019889f
C4246 commonsourceibias.n78 gnd 0.176331f
C4247 commonsourceibias.t25 gnd 0.019889f
C4248 commonsourceibias.t45 gnd 0.019889f
C4249 commonsourceibias.n79 gnd 0.175743f
C4250 commonsourceibias.n80 gnd 0.16376f
C4251 commonsourceibias.t33 gnd 0.019889f
C4252 commonsourceibias.t41 gnd 0.019889f
C4253 commonsourceibias.n81 gnd 0.175743f
C4254 commonsourceibias.n82 gnd 0.067443f
C4255 commonsourceibias.n83 gnd 0.081666f
C4256 commonsourceibias.n84 gnd 0.009217f
C4257 commonsourceibias.t100 gnd 0.172196f
C4258 commonsourceibias.t87 gnd 0.172196f
C4259 commonsourceibias.n85 gnd 0.068706f
C4260 commonsourceibias.n86 gnd 0.009217f
C4261 commonsourceibias.t115 gnd 0.172196f
C4262 commonsourceibias.n87 gnd 0.068706f
C4263 commonsourceibias.n88 gnd 0.009217f
C4264 commonsourceibias.t79 gnd 0.172196f
C4265 commonsourceibias.n89 gnd 0.068706f
C4266 commonsourceibias.n90 gnd 0.046399f
C4267 commonsourceibias.t66 gnd 0.172196f
C4268 commonsourceibias.t95 gnd 0.194303f
C4269 commonsourceibias.n91 gnd 0.079733f
C4270 commonsourceibias.n92 gnd 0.082545f
C4271 commonsourceibias.n93 gnd 0.01136f
C4272 commonsourceibias.n94 gnd 0.012567f
C4273 commonsourceibias.n95 gnd 0.009217f
C4274 commonsourceibias.n96 gnd 0.009217f
C4275 commonsourceibias.n97 gnd 0.012485f
C4276 commonsourceibias.n98 gnd 0.007456f
C4277 commonsourceibias.n99 gnd 0.01264f
C4278 commonsourceibias.n100 gnd 0.009217f
C4279 commonsourceibias.n101 gnd 0.009217f
C4280 commonsourceibias.n102 gnd 0.012717f
C4281 commonsourceibias.n103 gnd 0.010966f
C4282 commonsourceibias.n104 gnd 0.008898f
C4283 commonsourceibias.n105 gnd 0.009217f
C4284 commonsourceibias.n106 gnd 0.009217f
C4285 commonsourceibias.n107 gnd 0.011274f
C4286 commonsourceibias.n108 gnd 0.012653f
C4287 commonsourceibias.n109 gnd 0.068706f
C4288 commonsourceibias.n110 gnd 0.012568f
C4289 commonsourceibias.n111 gnd 0.009172f
C4290 commonsourceibias.n112 gnd 0.066626f
C4291 commonsourceibias.n113 gnd 0.009172f
C4292 commonsourceibias.n114 gnd 0.012568f
C4293 commonsourceibias.n115 gnd 0.068706f
C4294 commonsourceibias.n116 gnd 0.012653f
C4295 commonsourceibias.n117 gnd 0.011274f
C4296 commonsourceibias.n118 gnd 0.009217f
C4297 commonsourceibias.n119 gnd 0.009217f
C4298 commonsourceibias.n120 gnd 0.009217f
C4299 commonsourceibias.n121 gnd 0.010966f
C4300 commonsourceibias.n122 gnd 0.012717f
C4301 commonsourceibias.n123 gnd 0.068706f
C4302 commonsourceibias.n124 gnd 0.01264f
C4303 commonsourceibias.n125 gnd 0.009217f
C4304 commonsourceibias.n126 gnd 0.009217f
C4305 commonsourceibias.n127 gnd 0.009217f
C4306 commonsourceibias.n128 gnd 0.012485f
C4307 commonsourceibias.n129 gnd 0.068706f
C4308 commonsourceibias.n130 gnd 0.012567f
C4309 commonsourceibias.n131 gnd 0.01136f
C4310 commonsourceibias.n132 gnd 0.009217f
C4311 commonsourceibias.n133 gnd 0.009217f
C4312 commonsourceibias.n134 gnd 0.009349f
C4313 commonsourceibias.n135 gnd 0.009666f
C4314 commonsourceibias.n136 gnd 0.082208f
C4315 commonsourceibias.n137 gnd 0.05322f
C4316 commonsourceibias.n138 gnd 0.012299f
C4317 commonsourceibias.t89 gnd 0.18623f
C4318 commonsourceibias.t106 gnd 0.172196f
C4319 commonsourceibias.n139 gnd 0.068706f
C4320 commonsourceibias.n140 gnd 0.009217f
C4321 commonsourceibias.t101 gnd 0.172196f
C4322 commonsourceibias.n141 gnd 0.007456f
C4323 commonsourceibias.n142 gnd 0.009217f
C4324 commonsourceibias.t88 gnd 0.172196f
C4325 commonsourceibias.n143 gnd 0.008898f
C4326 commonsourceibias.n144 gnd 0.009217f
C4327 commonsourceibias.t105 gnd 0.172196f
C4328 commonsourceibias.n145 gnd 0.068706f
C4329 commonsourceibias.t99 gnd 0.172196f
C4330 commonsourceibias.n146 gnd 0.007444f
C4331 commonsourceibias.n147 gnd 0.009217f
C4332 commonsourceibias.t86 gnd 0.172196f
C4333 commonsourceibias.t108 gnd 0.172196f
C4334 commonsourceibias.n148 gnd 0.068706f
C4335 commonsourceibias.n149 gnd 0.009217f
C4336 commonsourceibias.t98 gnd 0.172196f
C4337 commonsourceibias.n150 gnd 0.068706f
C4338 commonsourceibias.n151 gnd 0.009217f
C4339 commonsourceibias.t112 gnd 0.172196f
C4340 commonsourceibias.n152 gnd 0.068706f
C4341 commonsourceibias.n153 gnd 0.046399f
C4342 commonsourceibias.t107 gnd 0.172196f
C4343 commonsourceibias.t97 gnd 0.194303f
C4344 commonsourceibias.n154 gnd 0.079733f
C4345 commonsourceibias.n155 gnd 0.082545f
C4346 commonsourceibias.n156 gnd 0.01136f
C4347 commonsourceibias.n157 gnd 0.012567f
C4348 commonsourceibias.n158 gnd 0.009217f
C4349 commonsourceibias.n159 gnd 0.009217f
C4350 commonsourceibias.n160 gnd 0.012485f
C4351 commonsourceibias.n161 gnd 0.007456f
C4352 commonsourceibias.n162 gnd 0.01264f
C4353 commonsourceibias.n163 gnd 0.009217f
C4354 commonsourceibias.n164 gnd 0.009217f
C4355 commonsourceibias.n165 gnd 0.012717f
C4356 commonsourceibias.n166 gnd 0.010966f
C4357 commonsourceibias.n167 gnd 0.008898f
C4358 commonsourceibias.n168 gnd 0.009217f
C4359 commonsourceibias.n169 gnd 0.009217f
C4360 commonsourceibias.n170 gnd 0.011274f
C4361 commonsourceibias.n171 gnd 0.012653f
C4362 commonsourceibias.n172 gnd 0.068706f
C4363 commonsourceibias.n173 gnd 0.012568f
C4364 commonsourceibias.n174 gnd 0.009217f
C4365 commonsourceibias.n175 gnd 0.009217f
C4366 commonsourceibias.n176 gnd 0.009217f
C4367 commonsourceibias.n177 gnd 0.012568f
C4368 commonsourceibias.n178 gnd 0.068706f
C4369 commonsourceibias.n179 gnd 0.012653f
C4370 commonsourceibias.n180 gnd 0.011274f
C4371 commonsourceibias.n181 gnd 0.009217f
C4372 commonsourceibias.n182 gnd 0.009217f
C4373 commonsourceibias.n183 gnd 0.009217f
C4374 commonsourceibias.n184 gnd 0.010966f
C4375 commonsourceibias.n185 gnd 0.012717f
C4376 commonsourceibias.n186 gnd 0.068706f
C4377 commonsourceibias.n187 gnd 0.01264f
C4378 commonsourceibias.n188 gnd 0.009217f
C4379 commonsourceibias.n189 gnd 0.009217f
C4380 commonsourceibias.n190 gnd 0.009217f
C4381 commonsourceibias.n191 gnd 0.012485f
C4382 commonsourceibias.n192 gnd 0.068706f
C4383 commonsourceibias.n193 gnd 0.012567f
C4384 commonsourceibias.n194 gnd 0.01136f
C4385 commonsourceibias.n195 gnd 0.009217f
C4386 commonsourceibias.n196 gnd 0.009217f
C4387 commonsourceibias.n197 gnd 0.009349f
C4388 commonsourceibias.n198 gnd 0.009666f
C4389 commonsourceibias.n199 gnd 0.082208f
C4390 commonsourceibias.n200 gnd 0.027976f
C4391 commonsourceibias.n201 gnd 0.147064f
C4392 commonsourceibias.n202 gnd 0.012299f
C4393 commonsourceibias.t50 gnd 0.172196f
C4394 commonsourceibias.n203 gnd 0.068706f
C4395 commonsourceibias.n204 gnd 0.009217f
C4396 commonsourceibias.t60 gnd 0.172196f
C4397 commonsourceibias.n205 gnd 0.007456f
C4398 commonsourceibias.n206 gnd 0.009217f
C4399 commonsourceibias.t104 gnd 0.172196f
C4400 commonsourceibias.n207 gnd 0.008898f
C4401 commonsourceibias.n208 gnd 0.009217f
C4402 commonsourceibias.t118 gnd 0.172196f
C4403 commonsourceibias.n209 gnd 0.068706f
C4404 commonsourceibias.t52 gnd 0.172196f
C4405 commonsourceibias.n210 gnd 0.007444f
C4406 commonsourceibias.n211 gnd 0.009217f
C4407 commonsourceibias.t93 gnd 0.172196f
C4408 commonsourceibias.t84 gnd 0.172196f
C4409 commonsourceibias.n212 gnd 0.068706f
C4410 commonsourceibias.n213 gnd 0.009217f
C4411 commonsourceibias.t49 gnd 0.172196f
C4412 commonsourceibias.n214 gnd 0.068706f
C4413 commonsourceibias.n215 gnd 0.009217f
C4414 commonsourceibias.t59 gnd 0.172196f
C4415 commonsourceibias.n216 gnd 0.068706f
C4416 commonsourceibias.n217 gnd 0.046399f
C4417 commonsourceibias.t75 gnd 0.172196f
C4418 commonsourceibias.t117 gnd 0.194303f
C4419 commonsourceibias.n218 gnd 0.079733f
C4420 commonsourceibias.n219 gnd 0.082545f
C4421 commonsourceibias.n220 gnd 0.01136f
C4422 commonsourceibias.n221 gnd 0.012567f
C4423 commonsourceibias.n222 gnd 0.009217f
C4424 commonsourceibias.n223 gnd 0.009217f
C4425 commonsourceibias.n224 gnd 0.012485f
C4426 commonsourceibias.n225 gnd 0.007456f
C4427 commonsourceibias.n226 gnd 0.01264f
C4428 commonsourceibias.n227 gnd 0.009217f
C4429 commonsourceibias.n228 gnd 0.009217f
C4430 commonsourceibias.n229 gnd 0.012717f
C4431 commonsourceibias.n230 gnd 0.010966f
C4432 commonsourceibias.n231 gnd 0.008898f
C4433 commonsourceibias.n232 gnd 0.009217f
C4434 commonsourceibias.n233 gnd 0.009217f
C4435 commonsourceibias.n234 gnd 0.011274f
C4436 commonsourceibias.n235 gnd 0.012653f
C4437 commonsourceibias.n236 gnd 0.068706f
C4438 commonsourceibias.n237 gnd 0.012568f
C4439 commonsourceibias.n238 gnd 0.009217f
C4440 commonsourceibias.n239 gnd 0.009217f
C4441 commonsourceibias.n240 gnd 0.009217f
C4442 commonsourceibias.n241 gnd 0.012568f
C4443 commonsourceibias.n242 gnd 0.068706f
C4444 commonsourceibias.n243 gnd 0.012653f
C4445 commonsourceibias.n244 gnd 0.011274f
C4446 commonsourceibias.n245 gnd 0.009217f
C4447 commonsourceibias.n246 gnd 0.009217f
C4448 commonsourceibias.n247 gnd 0.009217f
C4449 commonsourceibias.n248 gnd 0.010966f
C4450 commonsourceibias.n249 gnd 0.012717f
C4451 commonsourceibias.n250 gnd 0.068706f
C4452 commonsourceibias.n251 gnd 0.01264f
C4453 commonsourceibias.n252 gnd 0.009217f
C4454 commonsourceibias.n253 gnd 0.009217f
C4455 commonsourceibias.n254 gnd 0.009217f
C4456 commonsourceibias.n255 gnd 0.012485f
C4457 commonsourceibias.n256 gnd 0.068706f
C4458 commonsourceibias.n257 gnd 0.012567f
C4459 commonsourceibias.n258 gnd 0.01136f
C4460 commonsourceibias.n259 gnd 0.009217f
C4461 commonsourceibias.n260 gnd 0.009217f
C4462 commonsourceibias.n261 gnd 0.009349f
C4463 commonsourceibias.n262 gnd 0.009666f
C4464 commonsourceibias.t111 gnd 0.18623f
C4465 commonsourceibias.n263 gnd 0.082208f
C4466 commonsourceibias.n264 gnd 0.027976f
C4467 commonsourceibias.n265 gnd 0.517265f
C4468 commonsourceibias.n266 gnd 0.012299f
C4469 commonsourceibias.t114 gnd 0.18623f
C4470 commonsourceibias.t78 gnd 0.172196f
C4471 commonsourceibias.n267 gnd 0.068706f
C4472 commonsourceibias.n268 gnd 0.009217f
C4473 commonsourceibias.t53 gnd 0.172196f
C4474 commonsourceibias.n269 gnd 0.007456f
C4475 commonsourceibias.n270 gnd 0.009217f
C4476 commonsourceibias.t94 gnd 0.172196f
C4477 commonsourceibias.n271 gnd 0.008898f
C4478 commonsourceibias.n272 gnd 0.009217f
C4479 commonsourceibias.t113 gnd 0.172196f
C4480 commonsourceibias.n273 gnd 0.007444f
C4481 commonsourceibias.n274 gnd 0.009217f
C4482 commonsourceibias.t76 gnd 0.172196f
C4483 commonsourceibias.t65 gnd 0.172196f
C4484 commonsourceibias.n275 gnd 0.068706f
C4485 commonsourceibias.n276 gnd 0.009217f
C4486 commonsourceibias.t92 gnd 0.172196f
C4487 commonsourceibias.n277 gnd 0.068706f
C4488 commonsourceibias.n278 gnd 0.009217f
C4489 commonsourceibias.t63 gnd 0.172196f
C4490 commonsourceibias.n279 gnd 0.068706f
C4491 commonsourceibias.n280 gnd 0.046399f
C4492 commonsourceibias.t58 gnd 0.172196f
C4493 commonsourceibias.t70 gnd 0.194303f
C4494 commonsourceibias.n281 gnd 0.079733f
C4495 commonsourceibias.n282 gnd 0.082545f
C4496 commonsourceibias.n283 gnd 0.01136f
C4497 commonsourceibias.n284 gnd 0.012567f
C4498 commonsourceibias.n285 gnd 0.009217f
C4499 commonsourceibias.n286 gnd 0.009217f
C4500 commonsourceibias.n287 gnd 0.012485f
C4501 commonsourceibias.n288 gnd 0.007456f
C4502 commonsourceibias.n289 gnd 0.01264f
C4503 commonsourceibias.n290 gnd 0.009217f
C4504 commonsourceibias.n291 gnd 0.009217f
C4505 commonsourceibias.n292 gnd 0.012717f
C4506 commonsourceibias.n293 gnd 0.010966f
C4507 commonsourceibias.n294 gnd 0.008898f
C4508 commonsourceibias.n295 gnd 0.009217f
C4509 commonsourceibias.n296 gnd 0.009217f
C4510 commonsourceibias.n297 gnd 0.011274f
C4511 commonsourceibias.n298 gnd 0.012653f
C4512 commonsourceibias.n299 gnd 0.068706f
C4513 commonsourceibias.n300 gnd 0.012568f
C4514 commonsourceibias.n301 gnd 0.009172f
C4515 commonsourceibias.t5 gnd 0.019889f
C4516 commonsourceibias.t15 gnd 0.019889f
C4517 commonsourceibias.n302 gnd 0.176331f
C4518 commonsourceibias.t13 gnd 0.019889f
C4519 commonsourceibias.t39 gnd 0.019889f
C4520 commonsourceibias.n303 gnd 0.175743f
C4521 commonsourceibias.n304 gnd 0.16376f
C4522 commonsourceibias.t9 gnd 0.019889f
C4523 commonsourceibias.t1 gnd 0.019889f
C4524 commonsourceibias.n305 gnd 0.175743f
C4525 commonsourceibias.n306 gnd 0.067443f
C4526 commonsourceibias.n307 gnd 0.012299f
C4527 commonsourceibias.t46 gnd 0.172196f
C4528 commonsourceibias.n308 gnd 0.068706f
C4529 commonsourceibias.n309 gnd 0.009217f
C4530 commonsourceibias.t20 gnd 0.172196f
C4531 commonsourceibias.n310 gnd 0.007456f
C4532 commonsourceibias.n311 gnd 0.009217f
C4533 commonsourceibias.t36 gnd 0.172196f
C4534 commonsourceibias.n312 gnd 0.008898f
C4535 commonsourceibias.n313 gnd 0.009217f
C4536 commonsourceibias.t28 gnd 0.172196f
C4537 commonsourceibias.n314 gnd 0.007444f
C4538 commonsourceibias.n315 gnd 0.009217f
C4539 commonsourceibias.t0 gnd 0.172196f
C4540 commonsourceibias.t8 gnd 0.172196f
C4541 commonsourceibias.n316 gnd 0.068706f
C4542 commonsourceibias.n317 gnd 0.009217f
C4543 commonsourceibias.t38 gnd 0.172196f
C4544 commonsourceibias.n318 gnd 0.068706f
C4545 commonsourceibias.n319 gnd 0.009217f
C4546 commonsourceibias.t12 gnd 0.172196f
C4547 commonsourceibias.n320 gnd 0.068706f
C4548 commonsourceibias.n321 gnd 0.046399f
C4549 commonsourceibias.t14 gnd 0.172196f
C4550 commonsourceibias.t4 gnd 0.194303f
C4551 commonsourceibias.n322 gnd 0.079733f
C4552 commonsourceibias.n323 gnd 0.082545f
C4553 commonsourceibias.n324 gnd 0.01136f
C4554 commonsourceibias.n325 gnd 0.012567f
C4555 commonsourceibias.n326 gnd 0.009217f
C4556 commonsourceibias.n327 gnd 0.009217f
C4557 commonsourceibias.n328 gnd 0.012485f
C4558 commonsourceibias.n329 gnd 0.007456f
C4559 commonsourceibias.n330 gnd 0.01264f
C4560 commonsourceibias.n331 gnd 0.009217f
C4561 commonsourceibias.n332 gnd 0.009217f
C4562 commonsourceibias.n333 gnd 0.012717f
C4563 commonsourceibias.n334 gnd 0.010966f
C4564 commonsourceibias.n335 gnd 0.008898f
C4565 commonsourceibias.n336 gnd 0.009217f
C4566 commonsourceibias.n337 gnd 0.009217f
C4567 commonsourceibias.n338 gnd 0.011274f
C4568 commonsourceibias.n339 gnd 0.012653f
C4569 commonsourceibias.n340 gnd 0.068706f
C4570 commonsourceibias.n341 gnd 0.012568f
C4571 commonsourceibias.n342 gnd 0.009217f
C4572 commonsourceibias.n343 gnd 0.009217f
C4573 commonsourceibias.n344 gnd 0.009217f
C4574 commonsourceibias.n345 gnd 0.012568f
C4575 commonsourceibias.n346 gnd 0.068706f
C4576 commonsourceibias.n347 gnd 0.012653f
C4577 commonsourceibias.t10 gnd 0.172196f
C4578 commonsourceibias.n348 gnd 0.068706f
C4579 commonsourceibias.n349 gnd 0.011274f
C4580 commonsourceibias.n350 gnd 0.009217f
C4581 commonsourceibias.n351 gnd 0.009217f
C4582 commonsourceibias.n352 gnd 0.009217f
C4583 commonsourceibias.n353 gnd 0.010966f
C4584 commonsourceibias.n354 gnd 0.012717f
C4585 commonsourceibias.n355 gnd 0.068706f
C4586 commonsourceibias.n356 gnd 0.01264f
C4587 commonsourceibias.n357 gnd 0.009217f
C4588 commonsourceibias.n358 gnd 0.009217f
C4589 commonsourceibias.n359 gnd 0.009217f
C4590 commonsourceibias.n360 gnd 0.012485f
C4591 commonsourceibias.n361 gnd 0.068706f
C4592 commonsourceibias.n362 gnd 0.012567f
C4593 commonsourceibias.n363 gnd 0.01136f
C4594 commonsourceibias.n364 gnd 0.009217f
C4595 commonsourceibias.n365 gnd 0.009217f
C4596 commonsourceibias.n366 gnd 0.009349f
C4597 commonsourceibias.n367 gnd 0.009666f
C4598 commonsourceibias.t26 gnd 0.18623f
C4599 commonsourceibias.n368 gnd 0.082208f
C4600 commonsourceibias.n369 gnd 0.091197f
C4601 commonsourceibias.t47 gnd 0.019889f
C4602 commonsourceibias.t27 gnd 0.019889f
C4603 commonsourceibias.n370 gnd 0.175743f
C4604 commonsourceibias.n371 gnd 0.151855f
C4605 commonsourceibias.t37 gnd 0.019889f
C4606 commonsourceibias.t21 gnd 0.019889f
C4607 commonsourceibias.n372 gnd 0.175743f
C4608 commonsourceibias.n373 gnd 0.080726f
C4609 commonsourceibias.t29 gnd 0.019889f
C4610 commonsourceibias.t11 gnd 0.019889f
C4611 commonsourceibias.n374 gnd 0.175743f
C4612 commonsourceibias.n375 gnd 0.067443f
C4613 commonsourceibias.n376 gnd 0.081666f
C4614 commonsourceibias.n377 gnd 0.066626f
C4615 commonsourceibias.n378 gnd 0.009172f
C4616 commonsourceibias.n379 gnd 0.012568f
C4617 commonsourceibias.n380 gnd 0.068706f
C4618 commonsourceibias.n381 gnd 0.012653f
C4619 commonsourceibias.t64 gnd 0.172196f
C4620 commonsourceibias.n382 gnd 0.068706f
C4621 commonsourceibias.n383 gnd 0.011274f
C4622 commonsourceibias.n384 gnd 0.009217f
C4623 commonsourceibias.n385 gnd 0.009217f
C4624 commonsourceibias.n386 gnd 0.009217f
C4625 commonsourceibias.n387 gnd 0.010966f
C4626 commonsourceibias.n388 gnd 0.012717f
C4627 commonsourceibias.n389 gnd 0.068706f
C4628 commonsourceibias.n390 gnd 0.01264f
C4629 commonsourceibias.n391 gnd 0.009217f
C4630 commonsourceibias.n392 gnd 0.009217f
C4631 commonsourceibias.n393 gnd 0.009217f
C4632 commonsourceibias.n394 gnd 0.012485f
C4633 commonsourceibias.n395 gnd 0.068706f
C4634 commonsourceibias.n396 gnd 0.012567f
C4635 commonsourceibias.n397 gnd 0.01136f
C4636 commonsourceibias.n398 gnd 0.009217f
C4637 commonsourceibias.n399 gnd 0.009217f
C4638 commonsourceibias.n400 gnd 0.009349f
C4639 commonsourceibias.n401 gnd 0.009666f
C4640 commonsourceibias.n402 gnd 0.082208f
C4641 commonsourceibias.n403 gnd 0.05322f
C4642 commonsourceibias.n404 gnd 0.012299f
C4643 commonsourceibias.t91 gnd 0.172196f
C4644 commonsourceibias.n405 gnd 0.068706f
C4645 commonsourceibias.n406 gnd 0.009217f
C4646 commonsourceibias.t83 gnd 0.172196f
C4647 commonsourceibias.n407 gnd 0.007456f
C4648 commonsourceibias.n408 gnd 0.009217f
C4649 commonsourceibias.t73 gnd 0.172196f
C4650 commonsourceibias.n409 gnd 0.008898f
C4651 commonsourceibias.n410 gnd 0.009217f
C4652 commonsourceibias.t82 gnd 0.172196f
C4653 commonsourceibias.n411 gnd 0.007444f
C4654 commonsourceibias.n412 gnd 0.009217f
C4655 commonsourceibias.t103 gnd 0.172196f
C4656 commonsourceibias.t96 gnd 0.172196f
C4657 commonsourceibias.n413 gnd 0.068706f
C4658 commonsourceibias.n414 gnd 0.009217f
C4659 commonsourceibias.t81 gnd 0.172196f
C4660 commonsourceibias.n415 gnd 0.068706f
C4661 commonsourceibias.n416 gnd 0.009217f
C4662 commonsourceibias.t102 gnd 0.172196f
C4663 commonsourceibias.n417 gnd 0.068706f
C4664 commonsourceibias.n418 gnd 0.046399f
C4665 commonsourceibias.t116 gnd 0.172196f
C4666 commonsourceibias.t80 gnd 0.194303f
C4667 commonsourceibias.n419 gnd 0.079733f
C4668 commonsourceibias.n420 gnd 0.082545f
C4669 commonsourceibias.n421 gnd 0.01136f
C4670 commonsourceibias.n422 gnd 0.012567f
C4671 commonsourceibias.n423 gnd 0.009217f
C4672 commonsourceibias.n424 gnd 0.009217f
C4673 commonsourceibias.n425 gnd 0.012485f
C4674 commonsourceibias.n426 gnd 0.007456f
C4675 commonsourceibias.n427 gnd 0.01264f
C4676 commonsourceibias.n428 gnd 0.009217f
C4677 commonsourceibias.n429 gnd 0.009217f
C4678 commonsourceibias.n430 gnd 0.012717f
C4679 commonsourceibias.n431 gnd 0.010966f
C4680 commonsourceibias.n432 gnd 0.008898f
C4681 commonsourceibias.n433 gnd 0.009217f
C4682 commonsourceibias.n434 gnd 0.009217f
C4683 commonsourceibias.n435 gnd 0.011274f
C4684 commonsourceibias.n436 gnd 0.012653f
C4685 commonsourceibias.n437 gnd 0.068706f
C4686 commonsourceibias.n438 gnd 0.012568f
C4687 commonsourceibias.n439 gnd 0.009217f
C4688 commonsourceibias.n440 gnd 0.009217f
C4689 commonsourceibias.n441 gnd 0.009217f
C4690 commonsourceibias.n442 gnd 0.012568f
C4691 commonsourceibias.n443 gnd 0.068706f
C4692 commonsourceibias.n444 gnd 0.012653f
C4693 commonsourceibias.t90 gnd 0.172196f
C4694 commonsourceibias.n445 gnd 0.068706f
C4695 commonsourceibias.n446 gnd 0.011274f
C4696 commonsourceibias.n447 gnd 0.009217f
C4697 commonsourceibias.n448 gnd 0.009217f
C4698 commonsourceibias.n449 gnd 0.009217f
C4699 commonsourceibias.n450 gnd 0.010966f
C4700 commonsourceibias.n451 gnd 0.012717f
C4701 commonsourceibias.n452 gnd 0.068706f
C4702 commonsourceibias.n453 gnd 0.01264f
C4703 commonsourceibias.n454 gnd 0.009217f
C4704 commonsourceibias.n455 gnd 0.009217f
C4705 commonsourceibias.n456 gnd 0.009217f
C4706 commonsourceibias.n457 gnd 0.012485f
C4707 commonsourceibias.n458 gnd 0.068706f
C4708 commonsourceibias.n459 gnd 0.012567f
C4709 commonsourceibias.n460 gnd 0.01136f
C4710 commonsourceibias.n461 gnd 0.009217f
C4711 commonsourceibias.n462 gnd 0.009217f
C4712 commonsourceibias.n463 gnd 0.009349f
C4713 commonsourceibias.n464 gnd 0.009666f
C4714 commonsourceibias.t74 gnd 0.18623f
C4715 commonsourceibias.n465 gnd 0.082208f
C4716 commonsourceibias.n466 gnd 0.027976f
C4717 commonsourceibias.n467 gnd 0.147064f
C4718 commonsourceibias.n468 gnd 0.012299f
C4719 commonsourceibias.t62 gnd 0.172196f
C4720 commonsourceibias.n469 gnd 0.068706f
C4721 commonsourceibias.n470 gnd 0.009217f
C4722 commonsourceibias.t71 gnd 0.172196f
C4723 commonsourceibias.n471 gnd 0.007456f
C4724 commonsourceibias.n472 gnd 0.009217f
C4725 commonsourceibias.t48 gnd 0.172196f
C4726 commonsourceibias.n473 gnd 0.008898f
C4727 commonsourceibias.n474 gnd 0.009217f
C4728 commonsourceibias.t67 gnd 0.172196f
C4729 commonsourceibias.n475 gnd 0.007444f
C4730 commonsourceibias.n476 gnd 0.009217f
C4731 commonsourceibias.t77 gnd 0.172196f
C4732 commonsourceibias.t110 gnd 0.172196f
C4733 commonsourceibias.n477 gnd 0.068706f
C4734 commonsourceibias.n478 gnd 0.009217f
C4735 commonsourceibias.t61 gnd 0.172196f
C4736 commonsourceibias.n479 gnd 0.068706f
C4737 commonsourceibias.n480 gnd 0.009217f
C4738 commonsourceibias.t72 gnd 0.172196f
C4739 commonsourceibias.n481 gnd 0.068706f
C4740 commonsourceibias.n482 gnd 0.046399f
C4741 commonsourceibias.t68 gnd 0.172196f
C4742 commonsourceibias.t55 gnd 0.194303f
C4743 commonsourceibias.n483 gnd 0.079733f
C4744 commonsourceibias.n484 gnd 0.082545f
C4745 commonsourceibias.n485 gnd 0.01136f
C4746 commonsourceibias.n486 gnd 0.012567f
C4747 commonsourceibias.n487 gnd 0.009217f
C4748 commonsourceibias.n488 gnd 0.009217f
C4749 commonsourceibias.n489 gnd 0.012485f
C4750 commonsourceibias.n490 gnd 0.007456f
C4751 commonsourceibias.n491 gnd 0.01264f
C4752 commonsourceibias.n492 gnd 0.009217f
C4753 commonsourceibias.n493 gnd 0.009217f
C4754 commonsourceibias.n494 gnd 0.012717f
C4755 commonsourceibias.n495 gnd 0.010966f
C4756 commonsourceibias.n496 gnd 0.008898f
C4757 commonsourceibias.n497 gnd 0.009217f
C4758 commonsourceibias.n498 gnd 0.009217f
C4759 commonsourceibias.n499 gnd 0.011274f
C4760 commonsourceibias.n500 gnd 0.012653f
C4761 commonsourceibias.n501 gnd 0.068706f
C4762 commonsourceibias.n502 gnd 0.012568f
C4763 commonsourceibias.n503 gnd 0.009217f
C4764 commonsourceibias.n504 gnd 0.009217f
C4765 commonsourceibias.n505 gnd 0.009217f
C4766 commonsourceibias.n506 gnd 0.012568f
C4767 commonsourceibias.n507 gnd 0.068706f
C4768 commonsourceibias.n508 gnd 0.012653f
C4769 commonsourceibias.t57 gnd 0.172196f
C4770 commonsourceibias.n509 gnd 0.068706f
C4771 commonsourceibias.n510 gnd 0.011274f
C4772 commonsourceibias.n511 gnd 0.009217f
C4773 commonsourceibias.n512 gnd 0.009217f
C4774 commonsourceibias.n513 gnd 0.009217f
C4775 commonsourceibias.n514 gnd 0.010966f
C4776 commonsourceibias.n515 gnd 0.012717f
C4777 commonsourceibias.n516 gnd 0.068706f
C4778 commonsourceibias.n517 gnd 0.01264f
C4779 commonsourceibias.n518 gnd 0.009217f
C4780 commonsourceibias.n519 gnd 0.009217f
C4781 commonsourceibias.n520 gnd 0.009217f
C4782 commonsourceibias.n521 gnd 0.012485f
C4783 commonsourceibias.n522 gnd 0.068706f
C4784 commonsourceibias.n523 gnd 0.012567f
C4785 commonsourceibias.n524 gnd 0.01136f
C4786 commonsourceibias.n525 gnd 0.009217f
C4787 commonsourceibias.n526 gnd 0.009217f
C4788 commonsourceibias.n527 gnd 0.009349f
C4789 commonsourceibias.n528 gnd 0.009666f
C4790 commonsourceibias.t51 gnd 0.18623f
C4791 commonsourceibias.n529 gnd 0.082208f
C4792 commonsourceibias.n530 gnd 0.027976f
C4793 commonsourceibias.n531 gnd 0.194274f
C4794 commonsourceibias.n532 gnd 5.09694f
C4795 a_n5644_8799.t26 gnd 0.111879f
C4796 a_n5644_8799.t21 gnd 0.111879f
C4797 a_n5644_8799.t20 gnd 0.111879f
C4798 a_n5644_8799.n0 gnd 0.990799f
C4799 a_n5644_8799.t7 gnd 0.143844f
C4800 a_n5644_8799.t8 gnd 0.143844f
C4801 a_n5644_8799.n1 gnd 1.13452f
C4802 a_n5644_8799.t5 gnd 0.143844f
C4803 a_n5644_8799.t1 gnd 0.143844f
C4804 a_n5644_8799.n2 gnd 1.13265f
C4805 a_n5644_8799.n3 gnd 1.01812f
C4806 a_n5644_8799.t31 gnd 0.143844f
C4807 a_n5644_8799.t9 gnd 0.143844f
C4808 a_n5644_8799.n4 gnd 1.13265f
C4809 a_n5644_8799.n5 gnd 2.94695f
C4810 a_n5644_8799.t3 gnd 0.143844f
C4811 a_n5644_8799.t0 gnd 0.143844f
C4812 a_n5644_8799.n6 gnd 1.13452f
C4813 a_n5644_8799.t2 gnd 0.143844f
C4814 a_n5644_8799.t4 gnd 0.143844f
C4815 a_n5644_8799.n7 gnd 1.13265f
C4816 a_n5644_8799.n8 gnd 1.01811f
C4817 a_n5644_8799.t6 gnd 0.143844f
C4818 a_n5644_8799.t10 gnd 0.143844f
C4819 a_n5644_8799.n9 gnd 1.13265f
C4820 a_n5644_8799.n10 gnd 1.80867f
C4821 a_n5644_8799.n11 gnd 5.67846f
C4822 a_n5644_8799.n12 gnd 0.051846f
C4823 a_n5644_8799.t71 gnd 0.596445f
C4824 a_n5644_8799.n13 gnd 0.266384f
C4825 a_n5644_8799.n14 gnd 0.051846f
C4826 a_n5644_8799.n15 gnd 0.011765f
C4827 a_n5644_8799.t38 gnd 0.596445f
C4828 a_n5644_8799.n16 gnd 0.16507f
C4829 a_n5644_8799.t58 gnd 0.596445f
C4830 a_n5644_8799.t49 gnd 0.607734f
C4831 a_n5644_8799.n17 gnd 0.250039f
C4832 a_n5644_8799.n18 gnd 0.263347f
C4833 a_n5644_8799.n19 gnd 0.011765f
C4834 a_n5644_8799.t73 gnd 0.596445f
C4835 a_n5644_8799.n20 gnd 0.266384f
C4836 a_n5644_8799.n21 gnd 0.051846f
C4837 a_n5644_8799.n22 gnd 0.051846f
C4838 a_n5644_8799.n23 gnd 0.051846f
C4839 a_n5644_8799.n24 gnd 0.263667f
C4840 a_n5644_8799.t48 gnd 0.596445f
C4841 a_n5644_8799.n25 gnd 0.263667f
C4842 a_n5644_8799.n26 gnd 0.011765f
C4843 a_n5644_8799.n27 gnd 0.051846f
C4844 a_n5644_8799.n28 gnd 0.051846f
C4845 a_n5644_8799.n29 gnd 0.051846f
C4846 a_n5644_8799.n30 gnd 0.011765f
C4847 a_n5644_8799.t37 gnd 0.596445f
C4848 a_n5644_8799.n31 gnd 0.263347f
C4849 a_n5644_8799.t36 gnd 0.596445f
C4850 a_n5644_8799.n32 gnd 0.26095f
C4851 a_n5644_8799.n33 gnd 0.295016f
C4852 a_n5644_8799.n34 gnd 0.051846f
C4853 a_n5644_8799.t75 gnd 0.596445f
C4854 a_n5644_8799.n35 gnd 0.266384f
C4855 a_n5644_8799.n36 gnd 0.051846f
C4856 a_n5644_8799.n37 gnd 0.011765f
C4857 a_n5644_8799.t45 gnd 0.596445f
C4858 a_n5644_8799.n38 gnd 0.16507f
C4859 a_n5644_8799.t64 gnd 0.596445f
C4860 a_n5644_8799.t54 gnd 0.607734f
C4861 a_n5644_8799.n39 gnd 0.250039f
C4862 a_n5644_8799.n40 gnd 0.263347f
C4863 a_n5644_8799.n41 gnd 0.011765f
C4864 a_n5644_8799.t77 gnd 0.596445f
C4865 a_n5644_8799.n42 gnd 0.266384f
C4866 a_n5644_8799.n43 gnd 0.051846f
C4867 a_n5644_8799.n44 gnd 0.051846f
C4868 a_n5644_8799.n45 gnd 0.051846f
C4869 a_n5644_8799.n46 gnd 0.263667f
C4870 a_n5644_8799.t53 gnd 0.596445f
C4871 a_n5644_8799.n47 gnd 0.263667f
C4872 a_n5644_8799.n48 gnd 0.011765f
C4873 a_n5644_8799.n49 gnd 0.051846f
C4874 a_n5644_8799.n50 gnd 0.051846f
C4875 a_n5644_8799.n51 gnd 0.051846f
C4876 a_n5644_8799.n52 gnd 0.011765f
C4877 a_n5644_8799.t41 gnd 0.596445f
C4878 a_n5644_8799.n53 gnd 0.263347f
C4879 a_n5644_8799.t43 gnd 0.596445f
C4880 a_n5644_8799.n54 gnd 0.26095f
C4881 a_n5644_8799.n55 gnd 0.130362f
C4882 a_n5644_8799.n56 gnd 0.897033f
C4883 a_n5644_8799.n57 gnd 0.051846f
C4884 a_n5644_8799.t62 gnd 0.596445f
C4885 a_n5644_8799.n58 gnd 0.266384f
C4886 a_n5644_8799.n59 gnd 0.051846f
C4887 a_n5644_8799.n60 gnd 0.011765f
C4888 a_n5644_8799.t70 gnd 0.596445f
C4889 a_n5644_8799.n61 gnd 0.16507f
C4890 a_n5644_8799.t67 gnd 0.596445f
C4891 a_n5644_8799.t35 gnd 0.607734f
C4892 a_n5644_8799.n62 gnd 0.250039f
C4893 a_n5644_8799.n63 gnd 0.263347f
C4894 a_n5644_8799.n64 gnd 0.011765f
C4895 a_n5644_8799.t44 gnd 0.596445f
C4896 a_n5644_8799.n65 gnd 0.266384f
C4897 a_n5644_8799.n66 gnd 0.051846f
C4898 a_n5644_8799.n67 gnd 0.051846f
C4899 a_n5644_8799.n68 gnd 0.051846f
C4900 a_n5644_8799.n69 gnd 0.263667f
C4901 a_n5644_8799.t50 gnd 0.596445f
C4902 a_n5644_8799.n70 gnd 0.263667f
C4903 a_n5644_8799.n71 gnd 0.011765f
C4904 a_n5644_8799.n72 gnd 0.051846f
C4905 a_n5644_8799.n73 gnd 0.051846f
C4906 a_n5644_8799.n74 gnd 0.051846f
C4907 a_n5644_8799.n75 gnd 0.011765f
C4908 a_n5644_8799.t39 gnd 0.596445f
C4909 a_n5644_8799.n76 gnd 0.263347f
C4910 a_n5644_8799.t79 gnd 0.596445f
C4911 a_n5644_8799.n77 gnd 0.26095f
C4912 a_n5644_8799.n78 gnd 0.130362f
C4913 a_n5644_8799.n79 gnd 1.4561f
C4914 a_n5644_8799.n80 gnd 0.051846f
C4915 a_n5644_8799.t56 gnd 0.596445f
C4916 a_n5644_8799.t55 gnd 0.596445f
C4917 a_n5644_8799.t42 gnd 0.596445f
C4918 a_n5644_8799.n81 gnd 0.266384f
C4919 a_n5644_8799.n82 gnd 0.051846f
C4920 a_n5644_8799.t72 gnd 0.596445f
C4921 a_n5644_8799.t57 gnd 0.596445f
C4922 a_n5644_8799.n83 gnd 0.051846f
C4923 a_n5644_8799.t47 gnd 0.596445f
C4924 a_n5644_8799.n84 gnd 0.266384f
C4925 a_n5644_8799.t65 gnd 0.607734f
C4926 a_n5644_8799.n85 gnd 0.250039f
C4927 a_n5644_8799.t74 gnd 0.596445f
C4928 a_n5644_8799.n86 gnd 0.263347f
C4929 a_n5644_8799.n87 gnd 0.011765f
C4930 a_n5644_8799.n88 gnd 0.16507f
C4931 a_n5644_8799.n89 gnd 0.051846f
C4932 a_n5644_8799.n90 gnd 0.051846f
C4933 a_n5644_8799.n91 gnd 0.011765f
C4934 a_n5644_8799.n92 gnd 0.263667f
C4935 a_n5644_8799.n93 gnd 0.263667f
C4936 a_n5644_8799.n94 gnd 0.011765f
C4937 a_n5644_8799.n95 gnd 0.051846f
C4938 a_n5644_8799.n96 gnd 0.051846f
C4939 a_n5644_8799.n97 gnd 0.051846f
C4940 a_n5644_8799.n98 gnd 0.011765f
C4941 a_n5644_8799.n99 gnd 0.263347f
C4942 a_n5644_8799.n100 gnd 0.26095f
C4943 a_n5644_8799.n101 gnd 0.295016f
C4944 a_n5644_8799.n102 gnd 0.051846f
C4945 a_n5644_8799.t60 gnd 0.596445f
C4946 a_n5644_8799.t59 gnd 0.596445f
C4947 a_n5644_8799.t51 gnd 0.596445f
C4948 a_n5644_8799.n103 gnd 0.266384f
C4949 a_n5644_8799.n104 gnd 0.051846f
C4950 a_n5644_8799.t76 gnd 0.596445f
C4951 a_n5644_8799.t63 gnd 0.596445f
C4952 a_n5644_8799.n105 gnd 0.051846f
C4953 a_n5644_8799.t52 gnd 0.596445f
C4954 a_n5644_8799.n106 gnd 0.266384f
C4955 a_n5644_8799.t68 gnd 0.607734f
C4956 a_n5644_8799.n107 gnd 0.250039f
C4957 a_n5644_8799.t32 gnd 0.596445f
C4958 a_n5644_8799.n108 gnd 0.263347f
C4959 a_n5644_8799.n109 gnd 0.011765f
C4960 a_n5644_8799.n110 gnd 0.16507f
C4961 a_n5644_8799.n111 gnd 0.051846f
C4962 a_n5644_8799.n112 gnd 0.051846f
C4963 a_n5644_8799.n113 gnd 0.011765f
C4964 a_n5644_8799.n114 gnd 0.263667f
C4965 a_n5644_8799.n115 gnd 0.263667f
C4966 a_n5644_8799.n116 gnd 0.011765f
C4967 a_n5644_8799.n117 gnd 0.051846f
C4968 a_n5644_8799.n118 gnd 0.051846f
C4969 a_n5644_8799.n119 gnd 0.051846f
C4970 a_n5644_8799.n120 gnd 0.011765f
C4971 a_n5644_8799.n121 gnd 0.263347f
C4972 a_n5644_8799.n122 gnd 0.26095f
C4973 a_n5644_8799.n123 gnd 0.130362f
C4974 a_n5644_8799.n124 gnd 0.897033f
C4975 a_n5644_8799.n125 gnd 0.051846f
C4976 a_n5644_8799.t78 gnd 0.596445f
C4977 a_n5644_8799.t40 gnd 0.596445f
C4978 a_n5644_8799.t61 gnd 0.596445f
C4979 a_n5644_8799.n126 gnd 0.266384f
C4980 a_n5644_8799.n127 gnd 0.051846f
C4981 a_n5644_8799.t33 gnd 0.596445f
C4982 a_n5644_8799.t69 gnd 0.596445f
C4983 a_n5644_8799.n128 gnd 0.051846f
C4984 a_n5644_8799.t46 gnd 0.596445f
C4985 a_n5644_8799.n129 gnd 0.266384f
C4986 a_n5644_8799.t34 gnd 0.607734f
C4987 a_n5644_8799.n130 gnd 0.250039f
C4988 a_n5644_8799.t66 gnd 0.596445f
C4989 a_n5644_8799.n131 gnd 0.263347f
C4990 a_n5644_8799.n132 gnd 0.011765f
C4991 a_n5644_8799.n133 gnd 0.16507f
C4992 a_n5644_8799.n134 gnd 0.051846f
C4993 a_n5644_8799.n135 gnd 0.051846f
C4994 a_n5644_8799.n136 gnd 0.011765f
C4995 a_n5644_8799.n137 gnd 0.263667f
C4996 a_n5644_8799.n138 gnd 0.263667f
C4997 a_n5644_8799.n139 gnd 0.011765f
C4998 a_n5644_8799.n140 gnd 0.051846f
C4999 a_n5644_8799.n141 gnd 0.051846f
C5000 a_n5644_8799.n142 gnd 0.051846f
C5001 a_n5644_8799.n143 gnd 0.011765f
C5002 a_n5644_8799.n144 gnd 0.263347f
C5003 a_n5644_8799.n145 gnd 0.26095f
C5004 a_n5644_8799.n146 gnd 0.130362f
C5005 a_n5644_8799.n147 gnd 1.13032f
C5006 a_n5644_8799.n148 gnd 12.2154f
C5007 a_n5644_8799.n149 gnd 4.36511f
C5008 a_n5644_8799.t17 gnd 0.111879f
C5009 a_n5644_8799.t18 gnd 0.111879f
C5010 a_n5644_8799.n150 gnd 0.990799f
C5011 a_n5644_8799.t13 gnd 0.111879f
C5012 a_n5644_8799.t14 gnd 0.111879f
C5013 a_n5644_8799.n151 gnd 0.988601f
C5014 a_n5644_8799.n152 gnd 0.787466f
C5015 a_n5644_8799.t12 gnd 0.111879f
C5016 a_n5644_8799.t27 gnd 0.111879f
C5017 a_n5644_8799.n153 gnd 0.988601f
C5018 a_n5644_8799.n154 gnd 0.740399f
C5019 a_n5644_8799.t28 gnd 0.111879f
C5020 a_n5644_8799.t23 gnd 0.111879f
C5021 a_n5644_8799.n155 gnd 0.988601f
C5022 a_n5644_8799.n156 gnd 0.386686f
C5023 a_n5644_8799.t25 gnd 0.111879f
C5024 a_n5644_8799.t11 gnd 0.111879f
C5025 a_n5644_8799.n157 gnd 0.988601f
C5026 a_n5644_8799.n158 gnd 2.70455f
C5027 a_n5644_8799.t24 gnd 0.111879f
C5028 a_n5644_8799.t22 gnd 0.111879f
C5029 a_n5644_8799.n159 gnd 0.990799f
C5030 a_n5644_8799.t15 gnd 0.111879f
C5031 a_n5644_8799.t19 gnd 0.111879f
C5032 a_n5644_8799.n160 gnd 0.9886f
C5033 a_n5644_8799.n161 gnd 0.787468f
C5034 a_n5644_8799.t29 gnd 0.111879f
C5035 a_n5644_8799.t16 gnd 0.111879f
C5036 a_n5644_8799.n162 gnd 0.9886f
C5037 a_n5644_8799.n163 gnd 2.46205f
C5038 a_n5644_8799.n164 gnd 0.78747f
C5039 a_n5644_8799.n165 gnd 0.988597f
C5040 a_n5644_8799.t30 gnd 0.111879f
C5041 a_n3827_n3924.n0 gnd 1.70953f
C5042 a_n3827_n3924.n1 gnd 0.682769f
C5043 a_n3827_n3924.n2 gnd 1.24153f
C5044 a_n3827_n3924.n3 gnd 1.20073f
C5045 a_n3827_n3924.n4 gnd 1.70952f
C5046 a_n3827_n3924.n5 gnd 0.682766f
C5047 a_n3827_n3924.n6 gnd 1.54211f
C5048 a_n3827_n3924.n7 gnd 2.34829f
C5049 a_n3827_n3924.n8 gnd 1.67197f
C5050 a_n3827_n3924.n9 gnd 1.67197f
C5051 a_n3827_n3924.n10 gnd 2.84498f
C5052 a_n3827_n3924.n11 gnd 0.900148f
C5053 a_n3827_n3924.t4 gnd 0.091917f
C5054 a_n3827_n3924.t2 gnd 0.091917f
C5055 a_n3827_n3924.n12 gnd 0.750696f
C5056 a_n3827_n3924.t25 gnd 0.955301f
C5057 a_n3827_n3924.t38 gnd 0.091917f
C5058 a_n3827_n3924.t31 gnd 0.091917f
C5059 a_n3827_n3924.n13 gnd 0.750697f
C5060 a_n3827_n3924.t29 gnd 0.091917f
C5061 a_n3827_n3924.t28 gnd 0.091917f
C5062 a_n3827_n3924.n14 gnd 0.750697f
C5063 a_n3827_n3924.t32 gnd 0.091917f
C5064 a_n3827_n3924.t40 gnd 0.091917f
C5065 a_n3827_n3924.n15 gnd 0.750697f
C5066 a_n3827_n3924.t33 gnd 0.091917f
C5067 a_n3827_n3924.t24 gnd 0.091917f
C5068 a_n3827_n3924.n16 gnd 0.750697f
C5069 a_n3827_n3924.t39 gnd 0.955305f
C5070 a_n3827_n3924.t48 gnd 0.955305f
C5071 a_n3827_n3924.t6 gnd 0.091917f
C5072 a_n3827_n3924.t45 gnd 0.091917f
C5073 a_n3827_n3924.n17 gnd 0.750697f
C5074 a_n3827_n3924.t7 gnd 0.091917f
C5075 a_n3827_n3924.t5 gnd 0.091917f
C5076 a_n3827_n3924.n18 gnd 0.750697f
C5077 a_n3827_n3924.t13 gnd 0.091917f
C5078 a_n3827_n3924.t3 gnd 0.091917f
C5079 a_n3827_n3924.n19 gnd 0.750697f
C5080 a_n3827_n3924.t18 gnd 0.091917f
C5081 a_n3827_n3924.t12 gnd 0.091917f
C5082 a_n3827_n3924.n20 gnd 0.750697f
C5083 a_n3827_n3924.t22 gnd 0.955305f
C5084 a_n3827_n3924.t17 gnd 0.091917f
C5085 a_n3827_n3924.t19 gnd 0.091917f
C5086 a_n3827_n3924.n21 gnd 0.750696f
C5087 a_n3827_n3924.t46 gnd 0.091917f
C5088 a_n3827_n3924.t21 gnd 0.091917f
C5089 a_n3827_n3924.n22 gnd 0.750696f
C5090 a_n3827_n3924.t11 gnd 0.955301f
C5091 a_n3827_n3924.t23 gnd 0.955301f
C5092 a_n3827_n3924.t30 gnd 0.091917f
C5093 a_n3827_n3924.t42 gnd 0.091917f
C5094 a_n3827_n3924.n23 gnd 0.750696f
C5095 a_n3827_n3924.t35 gnd 0.091917f
C5096 a_n3827_n3924.t41 gnd 0.091917f
C5097 a_n3827_n3924.n24 gnd 0.750696f
C5098 a_n3827_n3924.t26 gnd 0.091917f
C5099 a_n3827_n3924.t36 gnd 0.091917f
C5100 a_n3827_n3924.n25 gnd 0.750696f
C5101 a_n3827_n3924.t34 gnd 0.091917f
C5102 a_n3827_n3924.t27 gnd 0.091917f
C5103 a_n3827_n3924.n26 gnd 0.750696f
C5104 a_n3827_n3924.t37 gnd 0.955301f
C5105 a_n3827_n3924.n27 gnd 0.862207f
C5106 a_n3827_n3924.t9 gnd 1.18864f
C5107 a_n3827_n3924.t0 gnd 1.18694f
C5108 a_n3827_n3924.t44 gnd 1.18694f
C5109 a_n3827_n3924.t10 gnd 1.18694f
C5110 a_n3827_n3924.t14 gnd 1.18694f
C5111 a_n3827_n3924.t16 gnd 1.18694f
C5112 a_n3827_n3924.t49 gnd 1.18694f
C5113 a_n3827_n3924.t8 gnd 1.18694f
C5114 a_n3827_n3924.t15 gnd 1.19019f
C5115 a_n3827_n3924.t47 gnd 1.18694f
C5116 a_n3827_n3924.n28 gnd 0.862207f
C5117 a_n3827_n3924.t20 gnd 0.955301f
C5118 a_n3827_n3924.t43 gnd 0.091917f
C5119 a_n3827_n3924.n29 gnd 0.750693f
C5120 a_n3827_n3924.t1 gnd 0.091917f
C5121 plus.n0 gnd 0.023253f
C5122 plus.t14 gnd 0.328886f
C5123 plus.n1 gnd 0.023253f
C5124 plus.t15 gnd 0.328886f
C5125 plus.t9 gnd 0.328886f
C5126 plus.n2 gnd 0.146102f
C5127 plus.n3 gnd 0.023253f
C5128 plus.t5 gnd 0.328886f
C5129 plus.t6 gnd 0.328886f
C5130 plus.n4 gnd 0.146102f
C5131 plus.n5 gnd 0.023253f
C5132 plus.t19 gnd 0.328886f
C5133 plus.t20 gnd 0.328886f
C5134 plus.n6 gnd 0.146102f
C5135 plus.n7 gnd 0.023253f
C5136 plus.t16 gnd 0.328886f
C5137 plus.t11 gnd 0.328886f
C5138 plus.n8 gnd 0.149991f
C5139 plus.t13 gnd 0.340409f
C5140 plus.n9 gnd 0.136249f
C5141 plus.n10 gnd 0.099252f
C5142 plus.n11 gnd 0.005277f
C5143 plus.n12 gnd 0.146102f
C5144 plus.n13 gnd 0.005277f
C5145 plus.n14 gnd 0.023253f
C5146 plus.n15 gnd 0.023253f
C5147 plus.n16 gnd 0.023253f
C5148 plus.n17 gnd 0.005277f
C5149 plus.n18 gnd 0.146102f
C5150 plus.n19 gnd 0.005277f
C5151 plus.n20 gnd 0.023253f
C5152 plus.n21 gnd 0.023253f
C5153 plus.n22 gnd 0.023253f
C5154 plus.n23 gnd 0.005277f
C5155 plus.n24 gnd 0.146102f
C5156 plus.n25 gnd 0.005277f
C5157 plus.n26 gnd 0.023253f
C5158 plus.n27 gnd 0.023253f
C5159 plus.n28 gnd 0.023253f
C5160 plus.n29 gnd 0.005277f
C5161 plus.n30 gnd 0.146102f
C5162 plus.n31 gnd 0.005277f
C5163 plus.n32 gnd 0.145887f
C5164 plus.n33 gnd 0.262676f
C5165 plus.n34 gnd 0.023253f
C5166 plus.n35 gnd 0.005277f
C5167 plus.t10 gnd 0.328886f
C5168 plus.n36 gnd 0.023253f
C5169 plus.n37 gnd 0.005277f
C5170 plus.t7 gnd 0.328886f
C5171 plus.n38 gnd 0.023253f
C5172 plus.n39 gnd 0.005277f
C5173 plus.t23 gnd 0.328886f
C5174 plus.n40 gnd 0.023253f
C5175 plus.n41 gnd 0.005277f
C5176 plus.t22 gnd 0.328886f
C5177 plus.t18 gnd 0.340409f
C5178 plus.t17 gnd 0.328886f
C5179 plus.n42 gnd 0.149991f
C5180 plus.n43 gnd 0.136249f
C5181 plus.n44 gnd 0.099252f
C5182 plus.n45 gnd 0.023253f
C5183 plus.n46 gnd 0.146102f
C5184 plus.n47 gnd 0.005277f
C5185 plus.t21 gnd 0.328886f
C5186 plus.n48 gnd 0.146102f
C5187 plus.n49 gnd 0.023253f
C5188 plus.n50 gnd 0.023253f
C5189 plus.n51 gnd 0.023253f
C5190 plus.n52 gnd 0.146102f
C5191 plus.n53 gnd 0.005277f
C5192 plus.t8 gnd 0.328886f
C5193 plus.n54 gnd 0.146102f
C5194 plus.n55 gnd 0.023253f
C5195 plus.n56 gnd 0.023253f
C5196 plus.n57 gnd 0.023253f
C5197 plus.n58 gnd 0.146102f
C5198 plus.n59 gnd 0.005277f
C5199 plus.t12 gnd 0.328886f
C5200 plus.n60 gnd 0.146102f
C5201 plus.n61 gnd 0.023253f
C5202 plus.n62 gnd 0.023253f
C5203 plus.n63 gnd 0.023253f
C5204 plus.n64 gnd 0.146102f
C5205 plus.n65 gnd 0.005277f
C5206 plus.t24 gnd 0.328886f
C5207 plus.n66 gnd 0.145887f
C5208 plus.n67 gnd 0.71725f
C5209 plus.n68 gnd 1.08466f
C5210 plus.t1 gnd 0.040141f
C5211 plus.t3 gnd 0.007168f
C5212 plus.t4 gnd 0.007168f
C5213 plus.n69 gnd 0.023247f
C5214 plus.n70 gnd 0.180471f
C5215 plus.t2 gnd 0.007168f
C5216 plus.t0 gnd 0.007168f
C5217 plus.n71 gnd 0.023247f
C5218 plus.n72 gnd 0.135466f
C5219 plus.n73 gnd 2.59716f
.ends

